

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gD7l84kB+WAh1ATog3H36h0/cMgn9QL5jGe9p9PjvP7N+FJAVvGVlrxcgBw6dZaWDNZqNANQuRFv
ZSE8fsSCFg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YQUcxim/tlzHeVlJ7otHN7u41KO3Yg5DFb1yF4GCsbXGLtUvWNlkFjY+UPIlgYImR4Zo4dTHJQ+j
3BaUNSUOqAVzT9CfyUelv2YD2ZTfAtzIe1Mboyb3+StKnuzxnZmIhVPiZlowdW5lQ1r7BjDPOsge
ztxOfUTbvYcTUE1ABIE=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eu4MFD/NMz3pssr62VCh1XDd9mthYydX9VaOq3lWUwHi5/7e5dl2SAWHtYwTnBgGPY+jCcMycJhy
WSlkhQxVj5BsMm2aAItwXFvH2mSbjlPggtI0/+DNGQ4x8LQSFLTDYnnQbBrHlJymsS+/asMkXACD
SJ2tF8LF5tMhAlMPZZ0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rNAzbNlIFUMjdhvgzZ2FokzvR4AuFtV+1AHGDKa9QgeBsZ1e0Fom48uKbJ9iakvqUoUcKKAvRzeY
OBkbx9P7Imx0gvIgzFsgiVw23cBYWOhbhSqVb7mef9aKx8yeF8T48n7gKldUkwBHIPeqaayRI9/Q
HCZO+k2+HCjRZE6L/Gzd+IOdEVUFOg3NtWFPk2JFkfZkxs8X7Vg/xxtvH7uvp+/EbVyiMbnwDT/p
NSqOyA+rJwBJYD3xRIPTFDI83XJLCF+1i4E8hyu7Y0F9MtjKugqEHwAG+JK3jde00nzNNaeLVUQ1
OfFMZJpkk0Cg66d2cvJY/G11oPkmvTq/JZ4+5g==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
apuTRT8aJu0TR7Ciy6ONiGK4AT7TUEiokS4gFf1g+kDg6PdKk9VRun4HKszIadRtahjPQo0of9uS
yvu3GS4EQo+Y+T116wnAIXnZSa8EQaEsDkziOI+rCvXv8IgaPYN8Cq0aRlASFL7IHOWNI49V0c0A
FIG/+5U7ZyNQFCVwuE4gCgK/pA6apm5kY4FGJft/EdZ5YAbR/nCTzK4P53+XsKHrtGfw+/MthFWz
tI0OtloKqc7laKZWKOVFqWq8Qmq7UL6utFODtxEQqzczH+q+Gw4rkUyOosIY+cbB67hX+GlmXXEF
jMwvUcen9t6c+wiH6rmBDcUIiuUHHz6q+jCwJQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dfDj35aI8y6zqcW/IHFxmCDw2mpyex25qQAUnsL+tIRxivv/85PqpCOrf3b7NWnwUKMrsxtw+JBY
mtlPsVxQKR1gn6VkaHwbEgwxXXxFe71Z+1nWQhfF8Nt55jGvq1joWKMrurSV7Mo+HkvHMSszXj3v
8ElD0S6sN91oml0nObejOhxzHf0ybK+sGag+CFA7aBr4k4rYglf7AzOYrPl3nNoCkyrFDQFa46/w
SXJm/os7zUHbsDI5GGUH3BU+NktHZV6GK3iyhtHTwrMgDtpGk6vKHMKULM1Gjv9g1/jp9Ao4cUhr
bCVOXM1v2e8A3564rmh3if78zTzCKamPRAB5Ig==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
AabbJR4gDsagM2rIXw5Cn9uasvL139Xven0Guy7rKn0iaTEmkK+paytaenytgrdHoRHwbySTa9CX
t02I4JMTAXYAl2yp8oPTpOHDlQszmnJVuU9sQYamRISTL9iMiuOSRLwhQWQk/d1R97dRhu66nv8X
z70k19ZAnOwZdHIl463RUtOAlGKRhAPgF0qpQqbQfiVXWWI0GUQOcA8/vRFR71fXHssiMkunQWdS
0gkE3KcL3Vmaw4/Xd8sOIPjlSjQhFE/6CDE+/0vzEBO9tMRUTRm5DXk7r52acq+xgQIzvfnp8zX1
NqoR92848mLib5kz6AI82wxHRjD+czT2Cy9O61JRLIc8x4MHcsAF+6TQHdL2MPek2rnrGCYHu8Q5
whOsgxnV47gviX8bSC+7omvFaKu8La8FXFYNDYyKEebnal9J8iEnAIjzUoaToEjbFCcqR6kCkSEd
g4f8165aphjdf38/tIKOpKjHZXi4Ig7xmEVzeOl4yZzPidYDnVjQ/SjiAWuU9NAGb8+q30FQ9MIn
oWtmgyDAG6F32kn8Bnn2PyftIyAw1YpBZci6y6CmwqPLnxJCo8lL5pS33Ezqyfc/d2pXRkvHmTSV
gUFTBuT0Ot/u/8iJKlpCqbY+lJraxUyh8bPuJYkf7zSpNKuiHwWClWSpfT9/IWyPhKdSYqTR0sBM
z1iWks1WTZXgwIkycE9uXQ+4RDIPWotGN8vb86c2KqOQZvUdi9F1+AUD0sIOZ33sWVnRBIQyFp8z
tAwS3dTD8kY9i5LXFM7LkpX+SRbjy4MrNrInZ2I4rJ4HEDr1/u0YR1UaRreb+bxEHq+eX17nhc2j
YQQE/X2m5H5z7WTLgmn2t+q8XZgtkOPjt7TpjkmF6smugFNyVuR3CD6mNU1YvbixcLDqiVB/v1p2
PmapsShPqKnlap1jEhgLzVU8/xbvdCzyDsQ59K1/XY7doUviRkbnMWnD4JvSqDYKek8FsvMbgxq0
imGgLVYO+3yyE1yVZgzTeZ+o6PXDVEtPKYncc/PMcCGS7Hk8xnqEZYVmWktrORe6tLdJ1Do/5gtC
SnwriwGcUh+XsZpJE/06K2jaFVrD1LjaM2FoHfd1w8QS5Xjbl3IhPcod4Yqn8iF15c7avHhkUFGd
oGMblffeaBKwcF46z9LM4x0vdkrw5szW9u5ZLOdOmVlgbHWKjEE288jDQ423bVoytCgqiW9A5HVR
m9yOqq9TXOEsXxM4Vlhz7XNRY+shH/UrUloVD/4a4zDM10uNYTiEBXxUzObhiEfEnvDRAounymk/
yRUu5C52BC1Zl9IpC+91TP7heFYijJ82kiiOniNwbvTUz6wIuVMtcNaIEZbdX756lwbh/HET/Q4O
aReIvlExz2Gk58UwtTJjsJ/bZAqRRH3LSlTJjFuv+skXzfpQ9MVQ9MDmlKiI5/n+AMeRXpu718fw
AdgQ5CurmOYJi7Y3K+qJ/gdKE3+LDSb/+4784wN/Ipi0kU5dlQ7zyIeaEQkbWIR6o0v5Udi5schp
pkHJPwODb1WbMntNtddFc2Y4+dseffTzGLSwHx3TJvLmftfRQvkEcknLGTDTj/M/R/4DqVw/G5S3
ZAiJkNmL52iM0ySFNCBcFZ3EJmm7Q2PxPIs2kxFxQMDN4/srusa26KA2XbyQ47h8wYLTW1pdzgnD
kq7HdR0fUUeVioZoNSk0+sKlC9m5X+Em2Qg28OE0yTWVqaXQsG3sVRSmLiL4HguCvvI8WusZcBZf
R3cT4NzSBBsHxpwmhAOzxVhhOqYQzTRO5HvIdurIN9bJs/poH+hbDREpYuzmB5fSHOJK+OqQQH8q
+TDesKve1ksN1F0M8TvSW5tRijIxm3yu06P1oxNqPoX/U0TwAdb721ikmRm7UfUIWYNo3MUPonRU
nOWigDlbtG11HDKw+Sp2e25oW8QUJacZygWLE2tKBtDnLmiIqnv4g7nlhkeJurrHV5GYuFGLTwSJ
OVGihajasb4bnIN1Z2zTyNcCW3XcXDiuuqtz4MU5PKr5n1Bi71oIvCny8EwDZrmuyD1ozTcNV/7H
1eH6YgtIHd4odvO66pLAdQw4iPsurov+vRBQWryhyPnaolE+KkxlYNTRIZB5zAHhiR4SP6ZGwcmb
fIBInA+QN6gPvx8LmAzmowX0iGAVsDUEhJOdxCvEnchFALH5j4dYN/qEDcs8BsLtlsfj+8mbJH6U
pzf9/sLRahnD4oKNU1nZ2IGwawhDdG+9eIDDkV5kB8aQwyDmq8mWtCGAa9K8vmNwNLr+O+SMrmjO
I4ypK58jVD4R/wnEJJB4EvW5PZcPXZc9g4Pqr6wqp949ofSVRCofcB81vZ2tXjQCJe58xqjQX5G5
Je1FQ6Z63uUwzJMjODyPhNbt0QtrvqPUqH0eHYsLOHXQD9NBZ0y9wMuXxBrIy6CEl+iekEHxcv0b
7E9N5I6CXSGx09StYsyFsGsvFCsmXgfU9yiemDGSXsqk6tDBQrvYeeKxtcg0Jt19TCJHm14TplZF
Y4dVOavA2CXYefoVuz4ek1Z3aIGEsXbBldkxJsDlnaL/EOy3r3lLgZEV+UhoGooow8OV0f87VXO+
SAbT6ZdL3SA7RBT6gl0Rr/FIwFrfhPnZWgTgVJCwKkZLIY+V4KDHXEZCTaHkBsQSDxRGNTPfUgya
I2s7eU72EIzdSVGG5mIAVaC2EdX3cD4V3w8nnWx+eOCSFrLoCFJKiahr8vS0z3NYGhuzat3Bdqj/
UB60U7BQ99/Gy2rSlczfp2VPTMLeUyPU36CdujCAwlORxzZU3TmuOKE0h+kurB4litNDoGVgoX8T
fpopmMaNSUegAW5l4PPqaKa2nMezHF8hXT1Y7RR6DMM8IGmbe9py3sapB2VsFJO4c4p/o1elprWV
ttNGwU3bBZqdikTcmXqMlxv1TC+22mfD4WE6S5aPCebM+Zpl0WPKO3UpsjStXhs9lXDhm0Efqs3J
uHw/w5fhGeF9kSDJYukZKP5VWfv6scvsjOPjEMqMwXDuVENWAXIUO7tDr5hFFG9oz5gdlpe+C6MC
M9hLIQx4AsTvmimgp8UYJflonuLiKyOLOWcIo/peBNGrXh7z7nRwFqwC7/hH9RWyLKkAscVKJO6V
mJxvq328/PupiyiBzPA6Hfvbc7K7Fji9dMrsvNT65o6Ad59umv/fMYZJ74VQy7ClL33ZiUYbabSa
Oyn1k8sfzxW+T+/I4zttq2oyKvZBgFbh2lkDXEbSeWA0dkrpcqZ+qDuGX8iXacdEdzLKaQri1A5M
tDemIjf8sk/ChzVnAibETue/HqJwhFP7uFzDh9xcxfThd99Yx4AICPND4B8gqwNOxSMp5Z00KGwc
GUhlshzKE4JINksZSts8BR16eUyQTzakNp01u0PHYq8FWVOFQi/LOTiw4R4RPvF5oAW5HE210nft
cOH7kBCxaxCNAuSTnHd9WrpOEGs65+Buuq1todnh2HHzXolk6Ejit87RibzmP7uakjykoAUsycBa
BSuqpQjJNafxWqLL/3eoIpjHyIgmh1Ogen2NV5MQbwnue5vk+WtiXFgC+I19lwQoPNZbgxZn6R13
x49OPjq6i/z2zhvEzS/ILIufQhABsWft+AaaNLzNZnD/Cr7mWKE95AqengTTfMI/Qi7E3G1CK6gx
kKoxS/jNiuFNMawMCejdx9pw3PZ5ri9EYe9oInpO81Cp+JIHvd5VIB3lePGz+ew5fRbhMw/7zav5
y4VieCNR743znngmq1WJoRcZ/VTsk9Yei82rV8a+05VZHV2hshQCXUr7QJiG2OCm6qxwgRIPQmtC
r2dBcIR7UzxpRigc8h0dj/IuBdqr6MmDKjubeTMaG3Gq0uHni0T6adQm9T64hWQQZJZjU3nfszsH
5UYgx02EexkMyCMy97yzhsH6cx7VjObyER+AbyFL4BCzm/4bZ5KPM+idPqnlY24D+PaEaEHQpzer
GXJU6vtKkcYU5swooJklTFrz4O4k919G4bIJk+KR3MwIU/SBikk5UcbV0Yr3LGQhxEqHVX/MPmjg
kGAfSBzbQ5XF+i01BnK7752JXTyFpijPaZrtjyKciwpcS32RSvePnEFQvEZ7sCLjDT6HXfoNFb53
gPibWmHHwQzw0r53HVJr7Ql7VOay3UdqKpLjJOLqM69Z3JuYmXNXraL3oSNV5ONMysSsQVW7xxrk
VATCGEe1VrUNU+JPfinBtQq3YF/4dQ8l3Ckz1zfbw178BbvXQWNv5zZ3l/tS56I79KZTTWSiW9iH
/Ij6g4/mCuNk4Um1vh9rxLHkxF+zWGnTZVMb3b54FnrdaKDjUmRU1R+/9s4186+18wID2RK2UIgg
a0lHOumnHX+NFwVoJ4IFa0tfnl/bJvX+UPKlOYKnUO5sC7GJzLrwzeKyFlEHGy9Rva1RWuQQUVoV
jNkOpcg71OlsEeWMJHLJxugJFL1pdeJG+EAUxWifK0lf9sbhK7sUgnAeflSSQzlIhnI0bJupqZU/
SJnWBTKcQYTsjQ2Xe3Iti3IWsucSSSUbcw3RvxJkfZaE4uUzz38BseTPj1jlhg5Kg4ZeIJvAfnHM
xf9CUZ2LGxpo0fAvCFLc//RnUxvfmUWeV3wpBnPCQlYgXSTxZ/nny3tn/T4gtZ4AWSsyJt6Dddro
Vi7JYPHQafbohWWCS3KEeTtZTVlmdrCR5m3SfNyfPQFayTv49YQ131ZIhcYiZxXtTo08wQF/L2F4
dVHjtQlbI1cWyfJJhqMk7kVbKSzRE/cFrQbBCSaUGiL64m5F3f75y0gCpXE5rLADzs4O3efl6vZh
wleVX+znuoJKpgvQ9UkdnEWBqwm6JBECXAThB0MJzHMIP7fJPMD88aFycG23bXv+/z9UmJm6JWK9
alHOvAqjuWOMwgQedt1ZdRbeuBpKC4KmjEOR4zMNqDaS5ZYbEpKefWSWCTBfmdayNC6ZQesrr7dj
Ay5yNesigPbejauW+SyZ/aCxsylkHoKHt9lYFYOtaDxMLOkZ+XLfVvCKzq+EIdi8aosMTqrrU8FK
l2Ke0krzX72py+Xgm/aiUztqTA5r5iDb7VxKAK4zyQAgX0+6olMK3UGAFDDuaBMk6WEsAiDRH7P+
faw7qmrTirBz/Ttv81vBjQhgLnpfyZ7lg/tGECZS1wA74RuLmZRbNf63RThPE1AEWywE8PSfb2bn
HYhLPse6IWashIRIPbe3eEJXzUwyP5eJioJTHGbrYz0bhP8Wyk+thpOEBN15gYlpsqmgw0RDqZ0S
4ws9l3HLrMRApuoo1VlbXXcVU2XpuBZMCG8M9aGhcM7DWeusEOx0Hdt3vpdfTbcRyQUY+3DIc0D1
p+aSArVwU7OmQLxbBgAiMuELKfeCnRiRhy3KdFuvWSS+22mc2+B0d6VETp3HxHW9gpZ7efXSdd+C
D99wqT95jyd0UyxGopshjVKMdp6eirRtbDgpTmbYTF/D31+p+bJOJUuARSp3k9aA/iv065iapLe9
2aajum506K8wUb9gVGn3/nwCFaCkabSGJyEktickNnEr826ie7Ph9s/clEuwotfr/VcKyWxi02wn
9Pw+mkbyG2frRaMoPqENOl/zXV9Cg10rwc3iboWwYxGfIZgnsY24IfquRtBmwlC3Vy1JQddeKajc
Jc+C0c9FdA8mI78vrNHYQFIQ6KMFDjsojy4VxayJzlunwhJxrgsF4eHtXEelR3T7AT/u/3lKJxYr
0IoWrZTCWAqfhMGNJaU+STwVC2E1KEbNKVbMg5ixiJGU406OEnoYH9I8mXb8MmSNFkZHJF10gw2m
+KWbZcFY4hO1XJzASV0yhYRAu6c1/JQRnTxGYdEXKLH6GIyLbyq76EtoNkW3KGPrBKlovfKC/cBW
JeMRKtXadkxAJOPO1V2Pyo5zOoLhVxyj5RtlKRfxjjblCh4w1CE2LhrZQrrwcL+dPi5gucPHZVTa
AyjioMrNI06sVs13/7LtACbZSpUrSdQYmKYNWTmEVjqsXz4HRVu1ncInbld2OyfPFQUJBoO25Exd
Jcy+7o7EATTBxM0SOn/OBr876RJAeoX7FET4amJ3oHC66ullLGI4oBVxDsua1GtSKF+bMVd3amEb
vriUvUenN8UWnpbtYDCbKEMRFayXWP2dv0w+6PdAaxhEYOwqyeGvVEf03XbJuV/nTQNbn1gbW6lk
cTO4Iq07eJDQbZw89+XgdlweGDqiAsKJE1T3a3cs+e33JQGsECMpmcw9OE6MTCzgTxLnpnUrb9Yy
JesnTGvD60T57rn1RMqYjGK2qtLkQU21KutgSzjOd3o++VPLNAelYaSVP5/EGrzRosTRUKU+Bk93
WFPb3MdBWYCBC99zezHv3YhU2/2okPdrxbS5ZR3g8PHHtGzxtjU9+VHk6aqDa/nIW9OzOFrhxXFD
PjQGiGv7pUz7Ldh+R0neTduhBDEamh2zLn8tlik3IkI+wTvCQA490NZxJlFsg1RCILI7s0a7J9bV
xGQWxvWIF30Oh5ehXDXTL/ZMiQUMzRjup07BpXRILGLlurzlBaSJ4MoLqtHDaxvea+yxHkdl0eDE
zo3VEbFlyWjjsYp23NC1IyAeQGOw5Z1tRwphLh5su5e6Uqr+Iar1gmRxayAB5ogpENjKL1sAnpR7
J4PL5Rq0eFatu8g7nlCYOPZPJIiIZE9tD9wcnC1IFB8Ri4Z6KPuTKptWFjDefWSsTc65BVPHRNUc
xROfxLWz8ggKOvYF1/fLj04zRGMqzJdvALXOsaPlBdEBXZdlOmU1sYj/D+T9k80lQkSIbmgMLuaa
AxocJMeVt4qwMEF3GWoKTgjKZNQvjY0n+bDHRqOE5/gsZUnfNWlokZjR6Cak6yG2vMU+ctaFohi9
c5K64gLec7qj0STnp5rmqR2buIuKqct5MWbonBaOLaUQeu/ZQ3lz5iNMrB4LBLEPh4iQ6uwxYcR9
uAu6NV0wvvascqK/ZVjNhZyQAGeISSZga1/w37tqEzy7RlWupErQ/GQ1+Ka8lpDndhpUXiNku8/2
KVNpPwI6s1TtY4MKFuvqmiuOvWdDL/Vo5pro78uqcPmRtmM0BgAy1wN+V5aI1l/NbiRNCJDo7qm3
tdEUC+psMModgkU=
`protect end_protected

