

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bx24XPMbQl0ZuYgzgnvmK2UJsn5v5rHRrHaBzymEsRVRAjuRN3xRCY+goyOwSGiaL5BZpex2sDSK
2sd0nljSnw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CSRfZVLMWm0HJLEB7NOFzWrGIhgXL0zMCnVPoqKjG5Ur0+RK898D8TnT1vzg0/m9z9AJo34CsLar
7ajBwWmQaStI2T7HakgiApYlcuC6de1XuIEH3rZRMj/RWcjpTLbgkrbMj7lCzKzQdvZHARVRsJHt
n6KxqqDLGxMs1/m4zV8=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YDR4T6HZUUPDmkJ3uEF/8DG9RH1KIm/Soi0XWVOdqKCDBSgk2PKH3QgKdeu/Ygc+E4sEfsdQ97ZX
ZNKLn57bC8vQMoMyVXHXP/gB1IkATHDtiORbiLIN6gz0rbLre/0AWJ4pnD6+ix+zJ2ZtVx7uSjJD
UeDwmSaYOZQhEg4QN3w=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b5TzJrebbTGq/pRucwAvmRYTRYSTXLJ31UHhj7qPdtWGaTRXaKbjtJHLK6r2fdEku+xRcQgb4iwR
VR2WDz2dfhkKseFS1Yxa2DFJTK597UszihjnkRHDocjQO3cUY+io6Cbq8kFDe4t/wEf721IVy63Z
z1z8RoAbpBZZGG1+seGG0kHDtkTe8wOMD9mRo2qsutfBPBsV5sK8/fmf9Y9E2sAlYwKjVvsGOjpr
dIS4pkfWNQ1UbQXn1WlPTe4wXcRDxSDWm2NMDLpVsB7PHxXe/ma6En4gcBeXFN40LqU3TWcyfbF4
Fgd267nviONJrvDRA6uaiECsHX40iXKsaxsGyQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LoXyfjLEjXF6IqzWN8H3K7nR07wwyqyXVISYV16h6KsboFmbDcRTEPo0gH2rwN+AX6fpfnjiQCDi
qZVj+jq+3Jpyaex4T6xZDGqASKvTFZ53Vog5975jRBzfQilhyEnt1jyw4Z0UhtEM8LILdgabJqA8
cXdC2MS8KixvDgzWP6ABnTAwC9pDqbLUIqs+coqVvcy1nM4qt9WlS3/X4SHWNrmKgZ5d/HUtKouY
9yGUMGTi2nl4U+Zd7UaI2yJjVCW8JLst+BTCam4lPyVXo4ebpoEbDK6tTwa5DlOxI45b/ZooNuYE
Rpmlrdz/peCtaLTTS4+P11HF/WIAxGHuvcXpOg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
splRKPjEH+uTzvqD2tjFWmYXGYcB4TmcJH8LhGT8ueKKhMoa+orNkr7mpiSfxGo4nOfb4ddB5A74
rXupMEGR44uXFXmGFms0uV3Mo+LAVOswYWiSib2qqWdsJAVPQV+uS8kwf1pFIhgSfyhJYccE2+LN
qen4ppn5nmwPuAnPwhqNoxWgV6I1SCeKHMvOOim/bGhWBFyFuI4F9GeL1p+BC2DYSvijB6DHJgjd
lmuMd4WuXe78W//Vv2jhHriZx5nGgRFuRWE3VBR/38AWtMEOOrO4ijdAV2GyHZrphPmDHXfSwU6z
9JSFgLsD3Pd9zxwPDkqCeFOIFV991nTMDEBaMg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16112)
`protect data_block
ZaAS219W6bcUidr2opI6O7MIiXTm/68NNm8SzK3+iEVJFgZ8sprbVwYZB43pd58WezpfAPEl2VC5
eNjqUQK5sgI1E1cDCU1Rz9Cn1o3xAx7vrEvRNEkz5SQaum1iiQB/Sn2kPIUN64Ir+NZNGjw63fNk
N96VFKfY6YiJLEkY4guX9w5LUr8XYzCf0hKYO1xf8lT72tJz1ZApmz+7Gjq/MMglrh53q1t4aKNA
i01EFJYaTiLvzhMkXYCZZtp2HokceehGGpI8ks7L+sR4yFxDBHfdZawVvPX7ERjb+VGr3aQXdxok
yO2y2QBMyK33V5Ue00NIsf1NIdzQFBDMQUMrg7QikIp3mi7ZhQWa8qUsz9YMI4APq1dtGauKV0Hb
Cs3y5Fi3f0gI5rM42ZkVH5iVNomMnzge6zKhWP28fujOqQjVkxxwreF0S9ob3DvoQ8Z6w2cIDDt2
pAImE+YoQvwWFXIZ8o1a6SyiqSKj6Awju8bIPoVlYOyX5tgSEjkDvS7epSDvdT35RiOTD2+M+PU3
HAVWn1k5qcCHU0GyUA/zC4eZ7GbTTXBVy9xKcAy/hS74ZtekV9zq3o4gLpf7IoIIVNrWULo9/jwE
U71vHfbQXwsgvoEl5vJ1V54OrHcYJAtmovZX5rda+xHx6wczb5PBq5ELEgi6ssEwEcDImusjw1yx
R/A3nD2S3LGYqWhXD+mA73cx2Fu7zuXAe8RvPdZI4qrMEk5P0q66HkEAi3nlPTRQ5TsOKmCmYyG4
cIxm+j7YHhb0wUUB0+LEDzZkLseDsp9+m1X1PbTk5B/rK8EGh44Xqs2wJ+tFFATpS64x37F5/Msr
GwLy329qVVKfjjQB1fmdIjHvR19yGtsJnfpEsYODfVuyp3Cr64mpehRuKPFpj8d8EK8KaT9ven+K
wtUuwx1VYXDLsR3oWthb7dLdZaXQJ5mKe4+UvDX11KG4VPVScTIpESKSS7NPxGdky9WGJp9TlDfv
OJoR1JVJvHXKO0wkBGKOJhq0gbQhR7eW3s12h7qO6RHxC69x6ZgcuOPy9fMT/L5RxLx908TF1lQ/
72zyoiKEQHzjtUUqmPooyTvJ3czZA1/BE1e8tsCzOC9s4CHueXHiZppDjx2ACWa14zBwDhqTKz8S
EqrnKomrCIeH7T4uJZBiLlJmvhpB7R7uY76wdtBW7+T22Dbv4V/RcvLAxq1ir3MzDYF0iACkMcXJ
HOdRkS2ABB0dAwctfG0GSzUIVjzLGe9GQffIKLKRAOh6W7Cw29Ffpn1Qc/qs8Rh+2smLdRfAPIEm
42BjTnsM5yNSzY4qz7/j4dnHrbtQF9MX/8RKV/ZMnbbc2DpLhU6WLuA0JZ/8soms7MmYeKF7FjUX
Yw2CzH+J70sWQ/de9M6Dx6qZm9EWDYLg5qwtVV46vAiTfdzAQF3ZTLGKdjI9KWgqiJf6zIU2Zk5e
HZG2bggjbcYDZUi9qgKVs/vskGgXDLHho5w2v3he2jYEVAr3SM8BzSdt89559OEPac2IK2OwGOJr
2Oitf+RBWFY5U6/IT4kct3viiPPS662iq3itSZ7n9+srKqRDPaCoATe8wHDcTcdN7LEQyV9OEri+
8pAcT/PLQZTTvKkgOo8zgMrwiHRmVAYvLe7pZou+1nSADiSvamZh9dtkCI9dnumfNGz2t7/z8BZ4
GO7ycPmM/QE4dvBL3PRKuFHLoeskzK9SVqS9Tudg7e1ORH+BMCAXhpdRlYQBTZESLKHdnci7bOWB
kONRQmC1/cnSfaI3NlZUV1H6UkBOWzmfelcDkmbPqA/YJ9ItotUev2zI1wxadrEAx/VQPlz2q0Nb
Y9SeFfrJLH8cCfjLAnmXwD0Iuic9alLPeHhI6iq8N9qSWz6TCpbiC1FSOUY62I7IYhGu1kD60zig
I2HLmyKJT3SbhdEmMTJQh48LFozN4FUGRD+MikKXnCDJOSS8H3O2ob6cJThqIacoDWhxzagmZ3L5
wnqHEzdPlFSlyC9mpYZYumriHfQjaZBQ5e/tgbS2YAH5eIwQs2fWluGrbyUua4ce3g1QQxYHgW0p
7swqFcrMTzk+xAWrxWJ9B+WzdLzudxqWKZETCAcQMa2rMQF5/KBV+TNkTHrRkzqTikJjiXUdSe/l
GhKtrsqeCGE4RGrviwpJXCrCNl7IbfdsLaQjovtTp4jCEuJk7LUYZvrTIjfsFvbXfiEvVpwmozq/
+2JglUH97YI2t/u0p9czH9jIkhruL+PUBlWlsXYvZLIegUu3utcaTXsI9Q7gH8Ytu47VzeOdmeH3
0IZH7XVyPZxINzAA1j7I18ThDYOZMG5Ndjx6b/voGXdoHxM9bRJYaOAXDu6mFC62Z4pvoC31GH52
s0/432ZbkYs+AxEs7R8F5ZNdRrj8adgGSgzyMLPRUtQlFwwkBtNTMp3d/wXk7HlAExTK4iChs5aU
tJOM8+JQH/w+11Xn69WHAL3LMjbNUUTn17QKG3iVJYl82+iSH23jeUXD2ccRxquntfJX4uMp84vL
0/q4lyKwfcXTofo84lduE1g+wT+JphcnrLryLUa0taWQmRmDJKjHX96SD8Nn+0MabXUF/RHgiWOL
hy1OywTVMBoT4QeYgh9fhJmhUYFTrEmihmTliyM2wQ4BRxfTjFE6QQLczpBH8TAzidlDvzVt2Gi/
emZO+jGnb3MekjCXYBRDVmR8P5VQuNREkbd6KZddI8mBdMzjOqgggkQyStfJPoHMmXw8Zx4tGEK4
h+t61iY5mRm0sy/ks8LfuDduyahM70FGV5c8O1bUTImr4y7NcNaO558m+nOvYxYS/B06XcBGOQa1
aTD75gDkKDouvazl65cB9veKt+d9YYn9b47MnNgUCt2TB1eHi8U7+KFNsO0/eB+8r6F6GLArlVEJ
uEPJiqQYiCQc5jtrBlibJzyd0TxwnZgGZox3mH/+rrahzvTwOvCge0Iu9vrJ5ws9ePEYlY6Yt8kC
7pQ7BteSYKbV8rLDwAVsznK07pwTEGutLGHkcGqYls//eEJOPChawPXvdgpSjU4FV2LPB6j9Nw+O
zsDVoHKs1YCjOHra9/37ZlLg/J4kCGMqL6PUOW6ddN1jxwBB9E76OAj8618IViEaOnPt+JH1LqAM
4mqe0d/j9TzaIuA5ekCJSY2a03Enjn7wgkcE+uLY994WIDi689fj4F3/LY9D/vKRlR/4gpCG8ydu
4PjogxFDh9t41dCNaIO/HPWCQSQEx682AaMqPdXB8rJnxCgcLu1axKi0to+gZ88yP4N/g9ojZnjy
QXersHu8oXu2Gv4NXIl3DX6cNka/qNL+f7J4LjvDoxxCmQWPBerD3YOynNjRewmjooqVowjryxkM
HlADt8a0VSip4l/rT9cGRgFjBpnNYQ5A64lItCRywapU5IsP+1j/5THpEUuHm+WJi2DsuIQZtGF5
Qez2M6sB07N95sF7Zc1ZD65UvN/Mr5l6E/tkj+pVlN0m2QUpJvSr4LPbmsZeBrvPhSLQfRgtMXrM
1gZOHFATE/EGLDTzQtkrJyOr6HL+eqoJUioI5Z+mPhdx6GFmdOTnxJdHzWC+tZZptvG1GQoHQRky
8CG6+LbLWlXLHgDxv6z8uKykPK/KGAI35NFaHgsJbdXzPnUit5PWneS9wagKLauDqzCYSNfYLU+Y
ppmE3hztVmvxyPuaWF/aWiHRBMIZWBN7HebswuqvZJHsGW20kkWF4ysPn+5+b9VREbj1hN0V9ZKh
nCbB09al2bDkVuxmTDnsMawDNUYla0sWI8ULI7D5mo5W3smN3Zl9FtPsoGrCPXTZQrBp4pwA2T4M
mHz6POW3qNTFeTNJ/qBJhLql9czAZBCDZxrZ6ZFOz9G3jgK1RdDFh8Qpe2SxeK6mO4kc54eB2q7t
Wu4OGXHH6jYQOPyju2El+ytbdGEpB66+pcdD8RNLD7p90Cmu4zza5RIWJm33NJ0oXzySyPWYJ84o
/I/brCK6dgAXOFllpa2/rkShvOO1AzV15MsJKNEXMkLnTk1CEyMH6YJocHwIgfw7WDOckvdMRVU9
ROGEQIVW4nfnCOqyaummcaIY50KYD33/qS2Rn1HUJrTQkQ3JiILrZt2aBJ9PbI9YSjWM7lqogEMm
ezr3a6AGl6NDtjYi3vSy4wM7BvCSZbQPM9vI2DQnNTuo/twq/VeCCY3/fX2gKWWHPqQ8Cxakf2N4
hTIvovNuTqeeYPyjT/1VqgMAY0BBPXBT/ZmNNmwNv2hG6exTNoPB7c3TbCITiXE53ytxaAZcyKHv
ERIn4Sr/MQTJ7n7Z0/JiS4IpD1tof1UnLxDzEfsSjqBJ3eB3CLl7LFMyfF984xnbr39b1sU89SzZ
7mZ+1O1FwjYV5gA8LTc+6ahDcFnBPNG6LDAHExcEjLl7cl3j0NhFa+XRvYWDRDePqFL7pQAEnRse
BRNAahpHh03KMaBNEZOWxEv82D9ygiIt7CVLJa9y/4SepzbuOR9Hj99FhjmMYdN6/bIIwAz3kQoj
6zy3Vtg6oz/2VFWYC5J46SeQtz2vo0rmjXhUudA6fzMRQQwpMBliIvaL+MpkwF6QjBFX9OMGPRmM
yQlunTia7uKln1Us0cecbCntjE9VkfKNvMOUlNsfn5F7FONsvBeKM6l9qX1nJkSCmJiySQKkAhtb
lLvbB0DK3yM6c2az8+OqTo7gv3wHPy4kMYqnZpV9Gu1++O1ZblezsDGjtrBdhuC/2WsR5Lmrih+L
vL9z6AdNZ05Cnlf85xRd75r4dQDOry6lAG+N40Y89WdUR+8h/gkB+nlDmRn0dSIC23CGuIQzY9+X
NemiRxmQKg8SMVdYOL0ncp1utVWaeybz4pAqIhX/dkitnWQ0eDIdNcVUOLvED3S+kECgeSCrnltB
UairwL7NxlWhsubeIhOYqxvxtPvC0PO0/X5JqVMGcljuyNK5D18tIH4xxvgrWUnZSGQ351wuTvbK
/vydZbT000WIkMpKbwV7wI4/ROZOAZz1vh7KrVR1596O/95zJ1wShCnCMl5gA/5Q29+sgVYyxPsS
QBxUzx2E+k/F3VvhUNBRuv+XLR0VjbojOREOKtk4eBILYgLwHJwqdv/dqNFnc8YOgsCUAzyCUqtS
4PuVDqIr2qE+zmAx2cwD49+LwGLwO9kyD9A136iC+GczX1+ijT1zotOfeuhm+gwgNs16dTe49j7c
hjvlIQ784KEnYxdZ334JCa4LR1g5TXhnQyBjs40RSMM3uqZp19n01QBPSjXBi/0L7pNQUbarthPD
Zmri1KK0AhNjK1rgV+aQojGxxs7qKhmZHi0Hu3h0Q8QfRasjTjP4G/F38Rc06iGiqdeZM0ymX+x4
Bs7dyhVeaiTmUkCcA0SG6G5yJIIftdZtZ+lid+IknWWyoG0/BDvNJo5nqm1kgvzH8ZSs5awBb+jG
mhH7FHy21opaHBmdGD/DjHzNgl0LFgYPpZ7SNGTUhQSz3bXT6oPRIi//v7EIGFGyxioZHxlDlBgM
hphDyAlOGUicg4AIIEAYqy15PrI8BcR6EDgFRIjGkEKG7l9F1FfEpWA/KFMk0/6A7CtJaBRMlntV
EQvQFHJOskRl6j1YVq3pliUjnYczCKkVAWpo7GY6emDdHH7N/2WxYDNbzpZS6TpA7C8Hx7JBo3Yz
5N66+B2EuC3PjtysGrxadcIiqvDUXSvW/R5EJ0o6e0QnfW8IKv1EocgJHrhMeRFUybWYs5ZsKPyU
+5VCqtXmDMU+6LxCd/6DBtV4TMoJs49wmdU0Rf0HqVq2zjHajAQbaecRRK/setuB99CDc8cDYsPn
SDFej5GR/7jIMK+UijTjsk/tIyRlKiDgrghgcstN7VfPQd2pcm+Ft5o1CXNBuXRtipINLSd+5xhO
qQUu1pgr9dVwrRbPY1bsfRaY+wgVhO4TbehINu05wVH8QffrCnvdyR0Y6IP5Q95eCjhL4B6kYCCc
i5PMc/l3QeHTXeMKBn/5jPAgLnwbYDrNT+oRzWmRIggOQFfdZSzX8TYJ4Q69h77sX8vQrQUUsUPa
3zleLR8ddYUUp7EqJmYmxy9D9F4EU5oud28/M0t+G1j0PRxaMZlTnSwOw9mXVuFQFcLpLKxGlFqW
HRT76BVuhnZMF3c59GG63eQaylsvHx/JBp4XJqJIFHqCHir5V7pDeKZfAmy9N+Rbw7zJKGN1PlnG
EtID3wfmeMmQaexIW0tMYgZHPrXOeYuxY78DS14Hsnad/evrel9J0lo8WheO+aS1B5PSsMh54nbA
8TOv/oG7lrEIHpaVQa265AqzA1AxTICGa+fiuGTFOjiUYwCiUlLRQnNhpI2u5lBnIJNjW7YuaRRA
GMJ4RdqyINceLAwcrlUc3rgTDNqkxmhn2pKF0qGH3Jriqu+NQAMjFEzdVwPM87CsIBdGI17MdLrT
dUlGcZaeCJBUhGUfxuPm1NC6f6mHIje+X7z0ylCVSH2WxVdApx7G3YiXehbAbmIPf2Gr1oaJveO+
5uRQ5wSrTXd9YtrQZSANSvYP/d2PGZhdSAyPsCMukETd+2Z+K1abjT9CwRHj2Hs80b162AGR/qXt
DU/GTZhwL89flfeGWd+fF+LLUPvQWz1vJoVbgz0B70wGh0v3FFIuW88ptTjj7x40QsC/1VdRHksL
Ep4keSv6/MjkKek/AIVsxd3Uutd+zK9sVLQWP/1s3+lVjz8fgXlau8r6/gb6suPHi+uXkSCJu4O2
zfIZhYksJWBHVT6E0LoqFeOP2YCRTpo3abcvwtP67vEJq/ZBb7FcRN389XbLmeWPGv2Hd7FM/2HF
SG2O9/Lqg0hn8XQ0y73WBYS/ShYx5Yx9rm4pFYV/pWzIfMv5FcYw6hq0+AdrUti+yBjQgKbIJnsX
slYaPE6bN77YEoByJ5BgTCIcDmi/AgpSzuF+gm9qx4ViVu09Aj67dXq0uikHXmMSYfCEDjYq4xyR
BKpGyWtySQdOdn06FXQfkAbPlTFkzxBNBa2yRPkzsE3V5l9hKJ4R4Dv1kphd9JGItzWT/FAgEKwY
X36cXdzgfh1uBKwBnLmEm5IFbhj4Cr60DKTVUIoaF6GJfQkpUBzdtJ54CAWVIq5N1PxbwS3QEQ08
G4EIZiV7ZSIAS50YJhwipfZsNUCJR+hODXP1vlb3rBJEkXNkdbzL7n2duAVV41ziQ4P26QLF4qI0
3hGf3l3rPychZTdWxaiVqfdXbN1hxJc/Vtsbl7v3FEz5+6g//kWKm9mqGtmZN36mEiUPrYMII35o
p5YVlYozoyhiezTHKzL7RaaFu9bPXRSNSwTxyEZFDCGldXNKnC1rXaJbf2YfzlhJxpDxrjsYl4L9
RcTLu0kAmAGvxRBSbhBAuB92V4hhCfb0BqumvFLZJS1a2Oq2rxeWaGFa+sOqYsFjvHEAW1Df2Jqi
jJedQDG+eyAgL39AU/Cf233cp3Vt/vSi13dNZrPY1jh9gemW7N7HQLlEzaJ5eRtzd5ROJt/JfLnY
w86Dy2K+xRzJ+0BTvpJV7ijdrou8gsiLb8hGU8moW6ODIm3NqnninEKmJ1reJbX4wQlij6cLITjF
G9+VTGSWK0pJiAPxiqwewBfSluS4XyvwUKO5M7HLn6bVglgZKuzU0Mxo3dtRjQnimNZum8Id66Zv
pHbskR0RSCnA1Xe946sudG0uQW/MzybBWTNCHTG26EYor5WJWIId8jHtltQGQz4Csk69d5fHrJ9o
5eVcjIjlvI8sw4dU62+oMBOAiBQVrbPsQC22USvbDqbScv2xh29Ea+C+ZWW8nxwe5fNsQMXYFaLY
KScypBWRaCo5Jz7+pNctNMi9ozDIqP0CPtj+RIF4Y4Zm0DhmuLD9j8BFlrN6ZQlde/GKmy7j01nm
xDJB9YXTsGfCNncZSTH9Uz8XNLcH5ebHSoH9Y7tvWhGRccXpSXUy4MPqlu/zRnRDrn5JP0EFg9nS
Q3s/q1tYZOzb+r+VpelC62wO5/WmaWi68a+JDItamf/gRJxlDm5jb8ZTVQI9V3D2624WZzM1mqGC
SYvSEIHco7s9rwK6RJ3wkMHAHzyYfTP90hPzJM4gB8MjNqIY7qktJUZDzCGum3TZ+hVIg/Icy9kM
l9q+IHuOo+LtlbzqqIjk7Q1FdoBnDORm1GK7cV/9oRBwhtIMz9g2T4ZLSymmJbEyMYZQI17C0xIL
/BhfJ1NgaUBnSTqZPsEOPW8TEGHHkLBcuHm2Eheg9Q92wr+/z8Ux8u8Fg2z+DLIE8verlamfSmnf
GEKhtmGB3+GHuyWemuyMYRlBw9pgULIAtqLcLY6iu0Ixr2MvKH9Img8Z8qWQwjXmIP5SJ6Wb+AXB
iTJN+qOAAJwvi1bT4++MKxG9px7Ag+ehxYyKfQJdqTXnf6hzJmmNN8jNVP8P1OZb67VRO93aIOlz
I8MHiwsZZkzQqw38XSkwhJYkm7bJtlOEkz6QtkAPV2KeK17665QQrKSVlrauuT/pJtTSlQPBkxQT
18OStf9WtJUhm0Wws/fDRn6B/BhGXsVgwAoFJttNZqTBJj9xuftaKkktrPOsBRbJzPTMbZLXA1Yg
LN48lXTMl3Y+++klRmb+pOVSMApbqayn9onyeM8Tj0xlqr3P6dBWjKVritPvs9aGdmGoQSZd2bko
5eZKGiU3uVStsGj5VvlhfNVH+BMiL5FcUaCHCuYI3dkEJsDXiCecTjpiJSnDDTLy28BMYGizM5xy
oyT35mba0lE23LGPl4ejhVzu9IwjWzRmBwEYl4bscffdGWvLAi39MxOGByPCe2it9y1VZJqxf32w
vlw/IpGJfMI7mmfpwfTC1/hR2Qdy4rg0IyHMS60KIvv2fztrP14IEET7bXR97IwzSgryTXywAkKv
4KfUGq7sV59G66mTib1AA0H9MdgInaSasXoWV1nxoJEiBWQUFkMmu36GfbRBGqyIizlNdvWw1cBL
qygH6/CllsbzHmA7NZo0qrkTv+hsLEomW9tm6W7gdIL4gJ4qHoQmc0nyVq6VCctvbTyZ/6b2haCb
UyffkpYo9QLDLiaB4LiOxhcqnm+L9NgZO+oTcwN8eAJbJKrCMZXNtWZMpE9zPTIv8i6cmMgefXGs
opIuDt43cN0qJKKBBWficOdeu1lntEhVyckob8Dh5jJOB2A+SiZQcAzBT2lwJLw9I1tZzxgiRQUI
Vo1nWPKTYg1EZO9e+pG0lBQOBOefEv1+3sRSPvSHp3lv4rjNJiZWd+69/h9OJ52BqMonlO7rQohu
CcY/4RpJMX58mOHpeSciewgAQzlNGtDEzdMSKv5ADMNEcQGDq/ZTk1ODFrNOaEYsyEMKHMteX7yV
boAtQLDlKXeQ5aXp+hleAfPihzIzeXjuvIeVvutHjihYAg9p8P2TmAZuVIOgL5Pg3jV8YLcubp5B
Aj+tVw0mVjt1VKUNXzm7c766ExFNM5KfX+REhAauYI3X3lXT8UvgVRtEev2nbhYzWmoXE72ckyal
F7vHrgM1FKOrWFbzq0nrmbcut05s4VAy04XNdAhQ7WSW+oy++D1CQFbIvbVkNX9MnbFvIfEEwO36
jechBYuNXwB2+1M8yO6jD+gx7t9wVfftP8zUlXWHRjyBGUFRzL4KM0f1xspLoDK8LHeunx3ReEje
Gglu7ukTmMQvPdtWipdyIMqZoYFtaLC2ud4+i37LbPla57b4ir2Y77zRB1lyivJxCtIan5vXHGhu
FSaNcER5EZrMSPS+8Mqutw6RVwbKOuLpZKyvXIlSmolTZh8f1GKd4XLoLExRJcaeVltj96NP4avW
Tn/j49l+ULd9wkqesroFYMrRtqOm7wzLr4VW6IAIWlX9a3h7T71WGMx1+JD/2P8XMyfGY/73IdmX
tGvz4k9a4dv9zZouGVY782Rq4ILnrCJmdsYFdG0uIRW2U9BM5dwqnDsXn/THs3THEoFk3mRs5Zgm
aLxXZdiVyc5GIhGmKQzPiHuOdT/BkcvztBD0Wz5aDeBovBNOwGZDhVFS4RT8maLsZ5tkLBt4leDb
iln5Fw9ixn31e/mESPLw61h7CtuSoQDop/29XiWGQ8m5kJx9YGkrETiKIcyY+AwPdGFYdr+4+H1C
kIpTftv8cXNhDnZnEkjJDA1sv0q0O76VdJ3CuEAElbEL8C4aL9kSx44scXq8hnWoZgMmUDiQl4Xf
7yHfrwF1SOZ4cIKnKIWpjVaUR34kGYKErSlCR9j/OLsSQvUS8HyLTk4GKVpjd/jg4MVzcu+TesVO
jc3XhYris9mtbPeGnIyVclFLnb4RkuhRYqV0wg9JZ3dsVXBmhq6PUkNJVATLapH/a03H2cpChfSR
oR1xnlwue5bVU7pbikTQ2+ncfN3oM4CkcipVM6zqB3kcHph8zQsxhUTe9o5V22hnTDEOW5+nkxKM
D6cPg1vttwZLJDujnNfW09zj/W9SwUVlX9HpoXJC80ccwwqTUk9ySixGi96ZNeeQ9g3+2nFIeF9U
ajS5b35syN7Yx8F2N0ajAgWtL8WP5DuXi8g1G+LK4rl5bFK6BDMXLdlxagl523r9cHBo2uKXTpvc
qo7QjrlRZPrQT5Ek5IKtJg9w6Io1dt74XdAZsPDr0a2l/VR6tSnQjETFiWSqFtlwdFAr09XphTvQ
KXvMQtI+RYlgvHc7KUKNhdBWGBKuJw956RihthPz2KQnvPPdixlNcShc/d0A0Z+jC1i65q5oM2qU
V+m1Cp7Gb1zz+CYn2FDUzf94iUQtdzIH5BsPBrpxqBI6y0/dNsXMhYh/eOStyt9fz2F8jVO2BTY1
4GEhzkcO1S/TzLxZa7cj8wb2TsSLyCGOAHlQ6G5Hz+sxUsQY2ffXt8LGv+r08OHGdTw4Ijphxgh0
eYxMRsWw8tU3720hjK8yCDsm6bz1hd+ywigfGxVdZbh5NvL7J8ndL+AsWmvp2b5uvHWKs8gdrO93
vf+0NVJ/wjACSDXAfuwzVq31PzB0UySyFqJQq2T2JzDaGaoTwfK7ZVjOitVPMkICzDvcgveSta8r
LwKZpkSp8jw4vJZ10ru7WBLA0RrsVIH4/SVgjtBkaVmkSfJ8UiCBXKAvUSjIBdoTKKclF//NF970
rzvNRpqgMbP165u6FdUONHwkd3kaIsxDjTnfigqZ97r7Cut5fHC1PLmFIgY68wDFBdpj5as+X5to
/dsj+NlHu92cu+QcfQIxrmsCBNsPtBvHCc3VHRkJ/GOrISQpj2IHHA6JA9S5CP/B3zjQssXxjgnF
2MLOIh1UJVMzcJD/IaNfYucPrvpI+RjR4bmrQ05h7dcNRx8cg3v1omWmjxaU/miLt0RoUazilARO
JFlAbk7Lgcq9tsFJNcSHnvsspUmf/8r/J1p3FEHPObhsVqATHWIbgCs8TYp6KO/8w3gEAwHm2Eb5
Q6guZwJ9kC2YhE2vEcVheCS24VDwUMmMCVZBTjpf611bQvFZOzaiZGMPKmT53NwuEnsyLzX355M4
5PiMyeuIIC9VqInNY+W3HMet5B1+nJWptFi88rAyqAF+zagM4V/tODJXG0Ge0ZytE/LTM0MjIvit
FEBwT6bvh4Xq7u6zMGj8ppBy1dfDWckr6Qcmr59dYgtpBlb0XlFKIRuH1odm6nUxAnTb/lAe8n2R
wq8sJYDUeMeGBF/dLCpJTK3QkrC85zVQ1ucunkT8VG1yIwYYKfeANUhUd/lhdUP9rjA9yTkHNAL4
CsJAGiH2FlI/8A6NodVomRgQ5P5I9gJ5nm2gbBQ7/gE+4Da24hMDD/6uHdhVMbbNV2rSNMnjO6Cd
yhV9BCVoxqx6OT7r1Vjqw5oY3W4gKCQu8AP0i0LZVZzwznLMN00uc253lQ2R2gUJnUnbe5LgL41a
gCpGLQCDaISzS09ynw0yBiUxN6RFDannBI4IffTJ4ZP5+VF0XZbVCP5MrmVORn1RsNbRqjeYdGmQ
paPQM5rstG7y48NwBzO1vOg+YmMQrhW6wrKilNAv6XX5RME/Qdjcw6WhHlT/IN5r6gRAJeovovfo
cF75j/wRxwXPaAYPZj91L+nqWr77h5HPKCwgPU4YJnyr2PBZ8jO5E7ZS+wco0tOqSYSYsg4P10wD
3m0wQ4ENu5fwH/otanwJ21RhJRTE60VbZ7ht/n/nvsdmR1UsbR1PJe8Mv3bXJx5YzZDADVMovgBM
wyzMRye3n8FoHXZrIcVN6YjRzGviHOdnHfpnGtgtYemvNUt6IeM3h3TIhh8kVUwGU8tjVmm57FI5
zGZtSrr1AQnyh890LbqRKuZ753JJbxQctipQ+Na4vXzaEHqqPmXDoG9EM9JfeWvJh9oBIDwZ6vKD
cLjMZHxqbGll/D9YOKYXMYCoF9HKew1ojEsd2GLQ1vLH+xIJZfTAq/PHAZsbJjuznL2zIUOwEIeP
ncZ8hdyEEoGq3dyhQ30dmht4RhpWsZtB4QhVqJp2EQBGjPm2prpOhXnjuNw8Lilv7RgOAt5R+Avj
n+6y6ly/d7cR/iAPqU+T4V7GbF+d1f2TNVPpDS6LwSpltNAVVTdKFw3kwxtmgNWxCPvUCTtIbbzW
ajKRki6B1+kDR5MmS5GCDU4hvQOh7Q1Kt3U1Db9PyuDx47MLV4QXHpkVVdluwj39XN2IYz98At4/
K4GCrhQYRowAx0baV5gkJELdsLyKT8PCuZHodsY7CgVeL52mh2uWyb/RF5pG/L3HAp7KB3EwydIF
GquLw2pbE88uRSLgaB4LyhvSjTNf7bZx3YBD9mVjJfEhHf5a0Ka6KBTr91u3peYe0iXtOHlzGtkG
7OgUyYI/XdFgbr6BZWjf5K9Y2EJnF3qVCZbbqLBWSjvBtIP6C1+yegcG0NC+IyWjf8sjPoAmrwHB
clnMOEiBujuasxX1pFd+G+g7Mvgp4ZmDmYCcfj4ZJP5GKOnD/y2r03lulpFYzz5VoriXUj/RrMm8
7Uw7mMq0CthEN+Xon2O+/mYE8G/BGtQr/ozVsO/ulGU2IA0NGLDzWXJL+s3KBaa8DASz33MkC3hZ
+bkZPqfTcTA7ir16XnJ0t3UDq4lWRJYi1xZKI1UPKjPtkAaGu64xQtj/RAVaf7wxZk6N3jXj6Gv2
EJ37UG0OoqLyC7UB4SdnpiXGxJGv9aUMPRhNFeYTLBwCzfOcXNikmI8zUbtCfzsBdkmRwhIVmulY
Z9uz3r79gU1+jaLBx0fzO0YKV3Kq5mtyf8a44o/2i09d6nHTICTCR9i4YNfGLTdRVvHpbh9arcl6
uY7eiNTQSMXWl0N2IB04QCkqY1tleEmziIrjT/1YRQB/fbcFAo+pM5U6jwaBNLB2gpxMvYKMOew5
iQjKyAyG0UW1IPyC36OBuggv1mFs/S8jtqIUfbzXEmih24rmaSRclVcmjHSpcrXSy+DCDJQi+bEU
gi5VUYRQCN1Ij6ZfH5pScfOY02I22PFKluTJ4lRCegphKhb47YuZyzvBd0nuKfZC09Gib4uzJb/Z
JI+KXMiYtVnlfcvIdzeNMfgDfCa3/vkQYzNBE6cZV/MEkpxvNm97wsfV5cxVtYrD3Id4J//Ftncg
TJOjJo7HBReoKyKHFtOwKUyRXc1BJpuhb+b7nyPb+tAPSuwD0F51HhdlJV8fTfqzxaPCgcO2Q8wM
i1/zwpUWwDzXi0Y8SQ6yFBq1sA/PkvMurLSnSLkfbIY2d3kLpzAvia0aZDv6oMFVpNYBulaUG4zF
zWhntWlafWisOhQ8smtFFyR6COzqW5Ch1NUR+uCxQFPVsI5iRfjIhUXHaYHv/CtgsRLprVpKQXaK
cU1iT1ayTmsTxVhfTU1Afow1bncJ3UitcFIt6w9hep81mS17qY3rGZZMAl9+JzoEcEfdqGId99Ot
ebQzs4S2WW+S2a06AMQx3FNGKVgXOqaLi2cnfOhGgJaiBJ1hZ/+s9utnwTyYNU3/HmWl5x3KnYOT
U7fkatVO/nd4w9CcIVVagAVwZLkfqeXH4lLsU/dX/kE9ZvtjJHNW9l/GbWTLww1c3LXqPkoJ3YIT
/wUoJNpaJ+VmcFk6SeehDSGAzfODYNTE1hxjNQfayF6iZ26p53W3/M+FYI+RX2c04fS9/X0FYYCD
dXCEqDLEJ4dLhB8LqZPMPgyFeXbvCeBTDqtfvBOliM/c5a7Xq2yz9ng9PkBozDygoj5ibPx8HGeO
HoYLENuUlykWzAe+eY9pdkN4hPoWXJstUBPRtthKuFX0qJnQC/jS3P1GrldOZlHO902Xy7NffpBw
0bIxPmyIiJtVP+Nj5fkRBres1XiHefgP20frADFvjo0+1WB/ppISR5JTOsR+BX2/n0xLX2P9lSn1
+mPPsZujNY76LlsHPJpqyVGOp2n3iiSw7Y3rwpLj6QUc8SKD0SeIch/EVi9IudOzSxHdnAmnhyez
zEZ9hbU0kHJK+UeWvCzaytAJaRUVqYQ6zD4mZ/RufCKgYeEHZofabighwp9nWsKTL9Ms2t2FlvSj
Msy08a8VouPvGao+pYornLpmXndMtEEep1sOYoiRjY2IFdpM2kG+81KISSrE5ZRLgx/F6b0qeEW/
WiAEAauY3W2z8pD9UZEjsVoIcMmI9IkpgYI8XEW9fA1+0IE8OnG8T3YyHk1zZniJdOq6f0b8FdF7
1GI++KGqS0Un2YN/BKHeG48KCE8J8EVCchJ0P+eel97wdbni7Toqw2xI2BrLhTkNHqXIch6GQyJG
SSJBWmr8Y6BWLrtw0YaMF3IOdpjulQEmop64Ty7ja8/3HC8kw/loRV+WpYzTv7KXJxY9qVbdoJ4Z
jqZ1QwHvrlL0vFw8jMgtFb05zRKJs6faHJFhf64gefDgeGDwERUr/6qdwuUesj6rXjPKMUz/qaJm
tI0GeK7Syq/2toSKeDkqwIE7ELp8dcvzKcCJw+MbzHabBLHmZWqb4J2hhW1HlcFyDCb7ww47xv57
m3a2s+aKF6Ee/PueOTA85bUsrZ2JIlwOsauE1EffBs1FIz52Uhts4KK0nnzapU4R8ublYR4ElA8s
INY5NgR4OSZheYB91Ubn6D3ShibUoyK0lFS+NurCQKvalAoWocSDSJrjirdVpqqzW87OpdIcoiJj
M5jJ6MhPfPjhuZFOcf/ijfQYWHGJPYN3oFi5ATsrcVAp1W9+sSU9ksON4onpDt4hMGvxGz96ND3r
AZ+9/UTFI4vU9lh+CusLjeAAmlsn7jrvV69hgvrz5svj8YFAMCj6ofvS912UMAu7YV8p781SNXra
glXNYnKskFO97rQA4UpxcFOZhrXTSi6TOrrKJzs9UM46g+mCtrtks7wFgx0PEF4PktGn2i4CRwy+
PaM+SLhhUUDpjLxo8s7J19Dw8K77qXrxkWm2IT3j658nrHaDQfp9YR8r2l/qTE5IIAJh4m+uCGK/
MqH1fEFV6GMZDM3xhr/4PZYuRSu4iXAJyDQmtfQSx8SefsfDTjz9BBrQ0h0u8Ik++QQYC2hDa8Fz
lQ7uwmeL/YDJifsI/qYWYQ7sLWuiNlxaoH0oiir9zu7rlNGG9tFzJJT6NKD+u5W3+jO4czZf+C25
KxV3o9h63b7vzZRDu3bxyUFl1JlYMgh8pr8/gFwJz/+eQIopkZ0LuXPmGKRpGSz7doxIh1JHvzox
s5Jr9W3vBNDH3P8O8tVxCMbiIs3s8lR7HoN4061S/QHWaGCOAl2eCopVpJ21GG4VZjKYBwultqyM
ZbMjEycKp4njbN4Guh/wih/1kvQv6oy9M73lysmwjPrKd5eTupYl5ZtLBrQzhRuZ6oTvye9HYMMu
nlw8ZsrOwierVY3LO57Hf7+O5BFKpPMgoP1ya7w4JHrUHtrMErvwU2bEOEjsRrEfWze8U8Iybm0p
XU13VKwodWQs6N+8DHewW3Uhh5a1GTHw8MLkXgoaov2MF1lOIYgmZtmpJCc0h8f/1BED+yy98+pp
V6sCyP+5lQ60ogv1Mt23jPtit+3gfUnKeSjbKW0ozeMK/SSgrk5F8vrywVXdxUyrM7353jzUqwO9
YQ9yHssvHGcy8ZQEB1bHY51dwMMeVwmH2ygyuPaLfXe07K9qZ8ouOLOBdkeIMyTWDly/BQWtDk6w
uZdv01F//IrPPODC0oBKl4rvgcnMHyA2VuN9Flgmy8n1Ir5qkSBcO2u2BrX71TUo/9zLNGT6ddrh
iWONmedFM47VyaFeaqO/f+CEvDnDnou6vulXbeqm0Qi/QNtL6mhQF4pGTv774hj6Bg04jGeo1lSG
An5WkPqivaDpDABuCD2p/sdzjZyPHw+BSvXV40HCBIB7iGprzSnsoYzGKa+VCNxfGswv/7m+3Grz
KU68gm1w16kXmiZvvlUzeahHzEmUJeTP8MXQVu6Z0i8LEUzVfquZQqVM3TMHk1j0hyzud8upuF/F
dX3Zha/HupMCQ2PbS0x79tm9iM/32ThN6rWjc+wvx8F+81W5JRcAhhrhB/ekrDXXxhKZHzB388A8
2txAfcjPR4VEB4qzBLJGk34KdgJm6FuoD1FYf3RyTGLI3rXHSJ5ZQNtaQQlNhrKIjnSzGULEzK13
buOZ6vQBd5flD21Ftfsg+47iSTxWT4miUnJPNW7HDu9dFsiDtFBWGVlH6rgsO7lxFUzkioE6OoYz
32vWGjp8H+c8U+Kd5O+x3LGJZlYtiSxPxAACk22jFvs20yajhlVLkmyNlr6KLTjZ2rOB3xqSaJB/
D6hULZqnmEnEOi53rdy4k8UPKMFijiSGdiQ1v69qlVR+H4GREOeAuiQVTxNQ08Cqr/dYBxcVq5Id
EvxqnsbUksGkJyX7uYaWZfT4tpbdXupfWiEyw3eNrQLH7GY+/UpsCIXw1Av0+iYvVclvI4vUPHYr
s0BA4mPLA+fQAfOagxvE8vXuFyYe3WSi/0jWkWfFDeP0oZxGQI/Vfk0QwOKAuaub/OoHZ8R/OxHR
BBJSHUOFmZPu9Yyywk0bSaY5yeuGGeIWvftv7Ow8XwHMbSFy0wZDx1c7mBK/LLbN1vTqbnwe/6g4
nvP4+4bdwQM+5/JtW/tG0o/+xHWZ84qPrIoCsLncKCyH2QAVIKYnJr9NVlBBOAKRTQtwlpi8NVQ6
+A7nH8SC65eej4Lf16G0s9+45i7+s3gcNGFdaecTblHPDNKiwoCj9jYq3Gqmzpa1ZfXi0FvwWmM0
2d+7JVNgpRvDIMnbRJdEhjOv5rv3FugTkOOR12ntIlxBtu7hg7zQbYXYdRTo1rjYLI8jM4CdyPp6
ECPwTkAk+yIlRoqjvVsZz9VBpgdgtf3Z9FJh9aQTW6ZBXCm+wTfs8tIwfJPWr99wbYQbEtoFgh7N
G2hf4DN04usibWQ09/TClrpUkI+CndlyVQ1TZM1Zwe9SvnZLmNsxobkIfBrcY/eSMhU5OHnE8k/+
ftcb4T46E+BY1Fh3nMm/7L65CWJmTEwleNwafoNiC4J1QGhHtQvyF/snqch6dQ2u5v9obnGffPgA
0Q9+nbKqlXWeR2jtBaF8e5STBlq97mp7jPJcRvFQuSpqo4wIiNxWb7hgODdMkrPmqevX40v4TiCO
9EjXtDHONGvunoLxxFqUFIfcn4yq5PkQjAmS6/Ko5xFhciSu0XZ3LLnPO3mtzQCvAa6cIgH8JSQw
WpSn8YEDr6o6gA786Y3qjcqD4wlwO/UFZFxdyED19adZf2mMgYcj09816uhh0Tk1pUr9IT8GL9HF
iJqAj+lYeFwEanDLatE7B7Dv7BAFJ3a4UrCzSL4nLZgEFu414pTw1/A/GI1INhdgVcLiiDbcu1EW
zE/rWZPr1f9OL7xW72WqRIY3tPovZ6eDlMie1vHg9wum1dL2tNZ2ku/uCo+2mdMG+sm04ggDwK+n
uxEN9JtIDRgG/wjHZ5sT5Axv3AX5/uCpszj2FWYHLaOUCBFlkusQNi5sJnXcf7bKaAKYW1/aAaZ9
92usXupN4rAccokX7UJrRSkNv7c11n4Hc6tq/YKcTVg9gvJVpqrJP3uosZopZ1hvQOt/M6sdRdSC
WEPVLZaxbzt3PeRyUunFvQLEB5GHmzt+h30cqxGvgwyfdPuLZiBLovxFkWMYGQKpNVz58x/kjRfM
FYio2lKBw74wiq7TnGp1ydp9Hw+5YAzLYEGMyYhEa1ewH3+0+V1UX/WoOMDl2bGHfiSrbffRuPih
0hwO+21FlLBVZDpB5hBKg07jwjgNZiEE3hA04yAjxBat8rY58PmlAA7VRRvZPBtqD9KX9w2pt5RR
bVe4xq1/p4c1H77qHmzw5KZwgF7cPRo6UkA3kP6AuUR10m6f4UaTMU+uIN91GUtsDAICF/11U3Xj
jrFiUxAjXV1pgGZlF1iLPq0QQQCQkmjC+AHZutCuVBDCCTkxwisTECjoZC4nsoriRxpgfw5HjJsP
Lq7K7Egy9HzRc3RiNhhEzdf/XY7eQwH78YO4PlqynRVcVbXvtjQhsfXuZLlHhGD+lIM80Gx56xq8
yhQ2tmIP2RHUO95wys/cYBxSsiLQex/9zRUKnJZktAGekeG26Tl/F3ppq5kk096sfeJj3bxxHCoe
BhZFwR8r3GqLQJ5iUDW9/bHHd4N6yBoiNEPrTlIhG2xjByIzKOvQFtVTzU8UsTVuVdzr+wbCAuak
5SWDzxIcMqOG8f45FAFgll5FD7piv7eKJ9UEJiV2jtVzrYlniKJ7YJJJYbhy8jq+BfhtPWomn5Mo
FOjesyIm9cwBXp3ITRAIVGWBZdfBaa0g+J/AKZJfZb3JdJu97F8AiB+/Lw3IYJ5xlg6SYVVXsDWd
0tV6Xe3B43iAss6Innnfo6jjhXmRc2LkAcz/M+FLhmXUJncU/JGXMSrLIx8e7uIthLwd7r1kEcF4
l4QfbirbmMM0INuufpA136rDwz//KJTvTQxjJgDLXxME7Q8h7AmQjVgbmFM0QmXSYFqm5wP4kYrx
CgjGx2np3SCCmtRt/SYpcez50m3WobjKTybvdzP/hu0vnZVPxRyGxFJgHmhHo92LuoubWvbZgHjW
8VOTjjfi1l46m+M0ulg0cmLVJENriUkdDEQiVDk9u3WXbjbs44Q+7VKXReoprMozuwh7O4iBNLye
6WJPPq8XvqW04l3Oj6LSUDujChPzQ2KstSt3BEfP7nxrSeX3bztcEfnB1VhLI5KidQo5xuQ4Hxf0
9rzCSISosJjwRFVzD1IykD2iyYUUTxffy4WL4aYkkYI1fMIR8bqPBziUoVtVsVB8NXC+8bPGkVvN
Qlu1tPQimuAQK6xS72NnYMJjPdn0rTjL6TKHmOsmkRl8ke+h+GvEEapZ52hbkPtoQPrwp/KQ+2uU
j2bk1MJCT140Cv5mSoQFvhejHPXl3t842tRwyDgj8NutRP4S6tJwuwtxc+Z/P4LPI6T4huqzLC2Q
DGk2KcIjJ9u5w84wi1NX2JDASYfQ8PRyLPoplr1cmRagBLXAgcXFjLsKQlUSBycfWQRwUMC/h05I
u32vmQlCjozI6/J/mWyHX1jpS8vi77tTmiNv/cjw++ZiDFyN28w720VCU/8FYx1fQ86cFruPLGA5
c5cpkfd77joy2FUgyuIzBrfLBE6xzm9snhUXL9MgZYaigLUBfLnb+W5FfzV9MNVP1xiStvNvEAui
oPeISB1ukjBq1rdVOwu+GXVNOxd6fSJT4BbQqwirwKns5ECgRNr6RkWaptE8/vlcGVblBXfkJjFy
5Cgp4JDqPJgMOQdlTuh/MOANOY/DGwxWn5Xlv4LBiyXsUAn0EwWoiInt5iGwoCBUh3mB80aqKnVh
1XnwYZYeTtO3yNbRJybmVVPieJssn7QQUWP/PyfnptvOfpRnIFmgHUDQXJftKjxJmpUN+pH4b6K1
T9IVHHUK8clEiiyHYD6oY5EdZ9XkXOaAAFAscnieqnfeku+dF2V3pV/wma3iMGC5NgOKuWHwdsRd
m5gGWA3VjutgeeUV2pvktLzHdl3erQB6xEye2I2BxFB+pnN9/DqsUOFYXgXi348mEpIGFLffGpQO
S2BUBxE3tbHQ7agDAQ0PI/KioxuiFshwo5mYsdsPnGjc9KM9DD9v6TyzCWnW1+WVqJngtpJnwzGd
dWNOvERfPgsu2wlgV8+kKxpNIgO7mk7vwXVOFnJkClKRcZHqHRWqMC84R2JS7NLQilN5mV9/ed8m
7AceJgvoSCkK9539UzX9uxEyypDKm8OB47g7QU9Cnhi+1wxfBdl+7yM/RzHxx16U5IKaaqdyHbIw
5AI6l8rJJr5s+ESB+YZtk+WFGpA2idxDUg1Hri8T8qeFex8HrA/EdQBY/SUfBwmZe7SAY+wn7E3Y
6C8sKc0GmagiSTwTj1w1HKc6C0Cp+OTCGgpnEDKS1Zj0WC9SMWeJYXBDg5QwNAxneTnnA1RzYEmc
MTDx4V0VqxaOEYhRFHJoMyzdr4xyvB6GR9djixTQvXGpnaksdftaz7mWh37eNHwSS+lsVzom2+5n
Yz8OWc6YOhDLFgGxF2UksyjKzSz+OpVAdUMWGb3tWfIfIkOA+B7XiyoGaqAl+53/GmRZ1dnMT1dI
s8uGxbZgGNCb9mwCOQJ4Lcb8guQOYUBhjuj+eYMZW2hJQqMtDAz8JZNe1Clgav/R5IDWniY6SIse
jxHawVqC/bKEABgFha9Vmlo4SRDAmf9WVypqmf/n5dpSFEiWzrtBDOMSk42R6jRASjvnfuEssdxd
ZIdwRBqqSf5IUbQdHM6dzFSSoDWZNIio4se4yvhWR+HuDMBI0KxU4QuzWJQ4Yod5pKgZ2gSOVycU
GpEwvzzPrm3WD+JpxgLNgHcmcwoBPjybUkhHgHYUR7SIANWudpyD8K8WVmmHzEI4vvaNhkRdQpW0
T2GFMTidkr2cwATRncVFK4HlwgTo3Q/KIpFTfpPtff/Jcr7QLABI4MVfvORmN/4MQRNnnYRNYeiZ
7THECYaLqsLdD0KIPsSKu2+vAkeqdvIVxrXq+1rB31yv9t8NFO51usK/alLpSCWYiAhxyLLAmLNx
9GWYEnLu1YQOjGwbvHlGem/iRHULUutxVtUD0uQMZoSfzuV7ieApUveX9dYcWHrNXSuTiJPjBiPj
pwiqaS5kCzn4+z9190mQLL1WtEaGKqOTS2V/cQ/SNQ9UT9bPvtRUKg45o9oICMu/TqL5i5uk6c5X
MS20Ma/eM/84DQ+fP2Y9+yEBEX/beaHruZWQ+maLtr8g4b7BwAHhsXrtspDUI592U/jOxtxGGcSN
HQhuui/1+Eb674ihmIZEMRMTUH4yXCz/TzBmCW99R9uL7zoXmGTDMnViujEzc5DatLlg6w0Bm5tw
v9W3dH3UKjhR18p5S5KC5oR/6yhQC9xOLGdGMnt+4A4djvhB3Eby99QrJjbJMLsb5ux/JR+hBvN9
KdnE01nttPe7aLJacUB/P4oKpbVFFO+1IjV/9OjLHqjnZWRpFOtiLAYx8IvLmPTEOW7pHLe4vUrR
DHroMEBy4LdZGFsd35EeDT17K139du6ZT6s1zqWSkc0hmSaBpANajUh7EuiBly2LXjLegQeBzazY
2S9qCTBmFBBjlzwlt1kaGWnp9ZiFtPHuaNeIZHn2Xr5VVIWB4TPeyjv5pjWNO9EpsZBJJBupFcPJ
bwAEFWvZhBDjvjlD2J300jiNSHTJw/sQ5GgUOKthmVU0ZtbTq14=
`protect end_protected

