

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U7hExZJod/vUi3z5N4RSr1wa48P7uP/A8O0jgaKOZBD7WNfzo6GmQd7doggkH00XJgs7nLyNvPm0
0zWCfXninQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k253ey4kkVql4FDzRxE0SZp0nnUl5fXV3ls/4mgbh/6ghGRjfZ71MsiTZ71s3tpy77tZHD0rpNoh
xUysBr1hFwWkTjAISVTsWyokKm82DELzMzaI0lqt04f7kevY+q4XugjttAECZCOOrrnUQb5ODPuL
TN/5/7rekkgE3das7WY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WoA52aV8kh0bkIXA7aISXPgNn7kpio3O4wNzPv7z4wZK/v9qsQ4Fa+1FXV0tZ0D+Si1URd5Yt8PQ
TB8Mp2LGBm7aAfzTAAqLpPZr3KRYlBsnuQptgQwkquHJi1BcDR3dhZHYw2oUKeYXBoZJ80Dg1iyE
mKNc2EAX8dBe7hH745fnWjhDqr0z4schwVFz8IHUPGI/WDdrXtDdyYzuiWdux2vjC9Gao0MkqalL
zCFAkEPTT0xtWcvaccmMU2ICHf+NVjiwhEmFT/vt1jXBw7quncqpEDMuzTHteQFztMFqsgBfXXAR
/Q4rfhaHiuQ7xUCcTEngpAsL2ypgKweMgL0LDw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yb4xLqu3x9ghRLjHN7QkYl0tDMsZMeJQgGEQuxDwwPb+acIMCaRAm0LVh6gbF0arOSlfOKBs+X6I
1sCY01AUXvqPtXEUt+RvllN5odbTYkY9f5RujZ5aQ9olezUe3+JLEML7oIeJ23v82E3q5lEn2hpd
Yirga3+XXZGIeEC2Q5F3LdU1PK/hOr/QQAn7r3cfSPSRAYJBv2q0KFRrpHEdaRVBAVRTnMADnWqM
+83djfdVuwjO+GhXELQ+rhNH9dkL0cqvHYfgIcRG0rYfPORpbXH4Uiizi44H6tpqRpTeCgmUfW/1
kW3FxovGX7M2+iedny4BJan5eJXy8iA1/NmnQw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pj6m4D23BtF6RtOvVlnmIzux1ocpf3A3ahzdQxUHuwpW9nlstiQd0oSmGGaiF66UD31sHUT6dfQd
yKhb6vxivgHto8LAAEiyTiUmNTH/c41wB3zGzcZFasAPOJZMvUysBGURofn88ip4eLF52/qIKVON
l8AKPEa6atmUOWXPGRix1yyvpjUnvxZ+wFAbBvP0ZsReS6AW7b6zRE+vUOJaMz0EaWEMMRdw3vLT
W/hp9Ruis3IsgHsdn6M611ZJnxSa2tuwXuWdXURUJzFjnTsi2R7EoD0bDJINDuh7T6iiDjBFdO8L
a4ER9/C3EG6IOxU+oP2sYgSHnI7dLthCIjJ+rw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B2bb9hbJCVaDRqGS393PhTqcBLIIS3eowUvDjLX1RVvD9vYwfdlG9rjfAUVzitJwz5TOhOabACyb
mMpxy7hxgVO56ex26Ce3uZlntRRrSfXZFQT0ENioLNV+BxEHrr7uipCant7HxRFrLFt9nR5wi4m9
ZZq5zS207DucLy0jTX0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eqzUQVv3z3gvc1IAF6D1gFpnG3jJXG9SSewyb0B7YFlkq+2WoV55oUnb7Smo54ZcwqBR15BnF2xS
jlkL+wI6xvjzAFZaDFixez8MkTdRnrNZscyGLFWOHz7RNKwEpAxAm7RSsBEcZUaS6x+lEu8Fai/i
gBi8OQLkjYbSnKt8sfNmpRhCWxhkRR0QylraXCBqvJVR8s/2S9YSm3zj5TqvYxlJahDh9O3V0iE2
aVTZ//VjzAQrgKQboTMB5R+3O0GmOfi7O8vgrOvK/PiOq6kVyAYEvce5/1FU9VRi8AQk3Hi7BRZM
1pWTxx+bC6qDX+NQvgu8HPGpHmqeqS/CQlftQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506800)
`protect data_block
YJlYUITjEbMzco72x/wW/x2fqTwAXwo+x/aKq15E0LMf9bSP5+VI2aCzLoTylIBCGJFEn1Mtj66s
DacYQVtTWQT6+b9GWO682SMGROAd2ikKHjf6ZbRiH4JYYotck8QoQpM9/1ow5KqgNjmznYslld5X
KOS9EjsuM1BLAj3PEW3FqfVQTq1ZRzJIFrg2wCuKoQz8WyCMmvarYIWYvZD3TKG8NqKTAjUvbutf
anUhiGcw12/AN2WvBl+7WKtAb64EfQWFGuuuvRG99vL3/JJUr3SgH2yngnZnjjQq1kB7fbm9o2Wg
7RfHeNy/s7PVLg+4A5l/OHXZMfDkI1iBCcCbay0tIsud1kM4PJ8L8ECqmisYb5Nha6CaTKWzq1Ox
5G40By/ebB23Xv4pPA+uaQaeKR35rON7CY7/qJlZ5nYEbDHxyIWVfLOK+o/xBSrWLeGwdktRsSv+
h83M1YsLczJpL9yNQ54CKHSgdcUGMA683+dOPLtmrnMb1NuPCgHRa2oxmLreGhLF2mKIykDjySuM
h6MyQkU/f6BB6QhXTNdR0Nab93TMgz4D3eTeR0V8e4VuqJuAboibYrIWPdn5QqGaqlIf1R/XDONV
eunKxlwKI4g8zEoU1wqENQGJa1gigwFcgck3v7YqlHnMtwDenQAOKJIpqicMlqmOs0wEnOCIYvZ/
Q8B/nBlHfq907jrvzHbqzOSZIlb1tT/PSCe4JA58LotOkSRCllJPXXkWdEZCbAsKkskt72NVweyr
kpI1ecLDMgYZ6jelv027NA1gSx6fPRsjz4ZTn+uba/XxasVmIaWf/8A+JBhSXKiroTIz4xkek4Ff
fY+O6h+nTFX9qe0qNdevOz+wAIwZGpG90EL5soQia1+eeAPUyWLMqON3U9evPsl8f8HsHCJuD9uA
tDpeczmJYf1sBXA+fo91uKCv1v9ci5KAxm2JVTL6WskBCrjXzi72yK/lzFYMzs5uvtQdnvCWD224
FPL63fAy7+yOHKscH9YGg0smVXKmCsSF6G11vutdZ3M7HcKcnUmS0m7twQ4MfqIzP52xNecZSqMe
QZEl4QDwzSdfGTKCtPi+FyuMcMdw6ySAfT2u+z+lFr9ZwjH3bka2m6yqCOCJKKrZgAwQ2F7DW7ue
LL8qrMTPLqIfqAdmDo2RQna0XcA1mQLwJMiNalp6xmT66CkcbJdiLmG0dog4b43r2SXmlIknrghQ
6LzpfjXa1m3Z3jD3O1Yxmlz/kRIAQfIeQRAjLTiHpH/QWpsZcnYGO55k8NKmb/r4IF1/b2FoYXWz
u0i07YmhtXIGnz3BNzuaLc3CxajfqqZcCXOQ/SuZR8Utg8JDmTPRuYq38F0Ua4wbvFAr+gQpfPsH
1Sq7IzCpfeoY1c0m/jszvoH2+Qnn1UeOZXoi+pRQb7vdTsfOY4Pj/djVpWC0tiOhXUWb0AgT+HsB
DasR/V4nrnyE8SxHaLWhjbc32trd67gWh39+kMY3HE6pM6Sty97vRkBXWNPPHide3zFDtJLfPTrQ
kHzuAG6p/l829Ph6+b2zdlV4HgvgYwWu3HGD/ANfQ9HZIQwSOcLzLDmFaK9UzgWeOWfj/9Lo3gNl
cNM23DB1n9gDroZ0Ziu0VqcOmclgZEpZ5RzBzohbtK71coZeHOZCLuY3kSr1KkNgd2PheJpilyAf
nChOau4Rwri/lE1wxeBt44hLtZE3jonrnaCdwJMpNn/uXjI3BOEoBHRu8xbhx2gSbcfDnCy+CBZa
+uKGTA7aR8HWnyAuSpmS20VR/IXbwYBok3v8ZzDw3IBA/lM/CTw+G8CUH4T3KZ227+pf0IAfOZTY
20QmIbh78A8XKvzcZ73n3X5hFaSbowO2BsQtuINPQPO/DXSdWtekIvQTL9fg9AnwcAnEE3I3w60S
HeR8dhb5Va3yKkSCvudM5lNJAnab60zkUqdSKjY2do5Mv0+BS4gthO01c6yuNia3QS9T5TjaBQn0
U0AXTeZX617eg9ql35HOrwtX703At1fgcMdKmj4nr13Qz5YZAnCiMQJRON78at4sbJPpkAott0Zi
eiFEe4efPxc2m84/uPiCMSfRfM2bqP0Ga2dei4roVRzIsOqeA+QSOaRBkI2T8icvVLGBtV1PZqLJ
e6DlsXeGQ3E53WMBklxq6VMTtlUn4zxk8ccWxCdlLhBTIFr1fCX90kCgsOJCL/+/W7o6uDLH5grK
oFcv6a63rvNXNn93NO4Tmf6bvRohzM3L8BtakAFwYf5selH4CKGBxD+3lYDRv6VQS4Z2SXQczhY2
iJEPMHtVxkAjwrI7yatBqtYPtyGB1GGYfl8N/8LCe6qow3MOSc4pxEA68vLijTbqsTjV//3z8h3P
tk2CWygE9cEpIhRveF/NAAHW8hzhlQiLqYYKjrM9FzIcJKnlZM0vcP3OkI0VatMGhIVV2Qvx9e6C
oIbt4+o2GefHZQQ770Hm4rde9V4TXzag8XC40Z0x7SNDO7xvlvmVWS3nA9/TePJrErOHQ9uTVrvZ
s3W1Ro8d/alBuLvTrWz1psRSyZ1l5JS/marJRd+j9zPrWHLzARfkoCv+3zCoseZk5RQXsTyeELT1
ufTAX52X+c4W0uQdK3aLrI5h4RLuT2zR5ITa0DyGcYY3c4oBYfDphFNQS9frf6Higv7EzHhl0iAO
GQMA8J4fR8kLO/Tif5XCYMxWUqUs5RBst/o0f9jJB7MBltxmTDnbdDfnl7MawJxmj9LzFMKcQFjl
qD78haKMuDIVtVaCMg7VGBruzC389mqbw/2+XZOTwkw2Odpu/2IZk/AYfr+GJ711ozNDWAWII//k
HdOpo3yTyL/bpWQfXB6Ll3wjbaHI42DgJJgvZMHDRC2rjas7TQFWw3IEpmEtcjDRwMpdIsdok7AS
1ybd7z2wpVlDl4cB2qzU+A6Wo8E3gQx6EsHSj/Qaf+T53cw3NXEHFGlpq41QmO/gbWv/nrgu3hTm
gLj/duuAKya+ZA9048p4K2wAu5CYuF5XjXthRqXq+0rlPr2tYjR9b+eGSXyyxcBFAIxYQvnyuwGI
jHrtLHiSpw5Y1g8MR8NuvTwSJfX3a3AR3i+0YlR2ewbHhHvo+PtiYpzIQvCVZAP5FQPc8DLAH9pB
63t81TL+bkuFg8jo8lNxuAfs8Jte99nvBwr3cUbggSc/vqMoOpdsWp4A2wm6z2seFGj4K/1ec+eO
M/U1Bott85AsQ5wbEFRxg3MpWCCojN2snNr1Y4Yu69OSL3ETzV7sUimkRs/NTelJ6D13thMpii6H
NobyrdHLOTTx6MTcZjXt1LIn5B6rJSZkO6/JxFh674z49wQKzSpL8psEGeArV4RXB+aA8iWo1w6E
bcyO67MlPfVKsxYzPnc6GIpzPlHg2GHf25BVuQRf7VHdi3WgvfWysZMdJ63DM0avT2Bjtt6yJKfa
Ce/w0/dmJdIWGNEHl947uyT6an+aW5mI/P8hKjK/4aha4N7RVQEt3tZZOz4RUQ6HWeA5kptKHztj
sJEv7S67U9Q6Yd964oA0ylhnhzi9LWerU8z7oaTuPc2xskBdNwoTD528lQd3pam7ym8y/C4VSCOs
ssyYAqGetM81JM9pBksuuSw7ijKCyrZGeoOnf/YgKOUyzW3jJf51SXoMOPQ7ovEsezfbEBWZ+SSp
Y+/4q4xWqK6QD6fyAzaIx42ZwPxOZcJNj5TiHgvzO/qKW3V1mSS3aliE4zgQSeIVqcYc+rLmIAm/
3hiVLhh1OxkfOK0UFHtsjSb8YaKES5gI99tkmX7D9KO9oQp7tq9NW6t8aPS2n6zWCmA8FyP6H+Y/
l95ljO1V3MbgZKZbDkTOzufQEmE7xAuU4PHQ81j90TrQESX7xmAqhIDelqpI2TLANwrqu6+E8ENE
VdV6OgZB/LIGQ78+VpKZkc+4reolSrKTyif/p5UokcJXA/DJVFO4YWS53dT+ID3NIKo+EYQ1e7IB
9XiqQl6u/T4qLCr5taFgutbZXo2Ly/jqIsBU+SjLAnmMpip3rJHogrd4y5c3le2aj6odCrqnV88N
tYGBZ21UlRjt4IkdOfeqenBDdtpiRSMvijly5nj4pDytiSSL4svQuAWJSOP9QW8q3na6OOneCaJr
AKQuF3d4RPqbpW7MA6pkSZDUCycTvKtF4BDeBK0NwlW4jejUgsz7tMeQJMca1GlVduNsh9kvDG2C
pCfGapdFReZZnQ77PsVdoQhkKF5gyIMqmu/8JraAhr9pm/2zKyRge34YkxaaikAJalxdNG29l8HS
qZiBXfQCwvgdVjXfSSD9kP/F4qVGrQ2Zs2NI5H3rGd7+nK7p4j2UT+cSo+NvanQrjgLLtqmWVbhN
DwdBEcgQxaWVEIHE99VTJ2a1Q77hlSRLq0ljVoY4SKrn0buc2gUCKG0asvNAYd0ltEpptv7xeWml
FxwxGtJPGmDLszxWfKhdq7UIwzsR3HbJYmiiXzysOOOTClVLhkWTl2ccUyxroLw6ui/HoGVTT9CN
+zainQ1HiG6Fztnmc7XvsLywfug435LxN33tOXVIy1xYWs/cqGA0NPFKVfTwHdmacjBANzKwQVUe
9X4IhTVSMD4by7P94crI3tDEWbl1WEO9w0iNihhAwZpr6QjwtvXZOWc5JiQoUJLbOqhZISluZCyc
gJpd+ZA9kevFheuXlGykq42RD4/d8LUqPkqKmuRXANI8hzBIyWboBZmVq4nf9LcY2ZWSMMjKp5zy
q2Jf5NFrGXEXMGdEsUcxoZLVsnLoM+VfHNypedfK/9SpBCdgKmZrEwz970JN4TmgXxGcodx9WZE4
lcZrrGXBfBEPsHnpcgQPjh/JKhdm3UZJMKtRBqBGRNFPTmDg6AwleTsDLXcRJx4P3kyVk++5vXU+
JGrHU+nfbRRsxOcY14U/BA1SWrErb2hciKYC9VHyYUlUk3w49AAi44H4Spz8oBT/LwPoPrgbvi8+
sPdPdf2epR8rn/b78KRgdAfNiPkEYIHWTSTXcTRBWCmwGIFurPvZQzKNdM+s6rKYAjjBAC5Y1xfm
qMsutkM+TVtoN1kJMWb/C+HMiMjgmqx3KgPeoNjA6T56IMJL3g5zHBE13GZvAXAPE6XjHDyHsYLG
TjVdH3jVDWgA8yqfMBs4KbGwUNA8mPgDDKhkyYazu7ahX14VlibMrz2a8GmaKcBFnfHy3o8T9hHU
OnpCXURWJJuBiGgBIZgnaXWazwiq/29V+z96baS82N2/dRCmsArBeqWP5ElM+fhkR525s+lahk/g
vRBqZ7fMa7jZqrPtWIEG6DS6oeT6xZ4W754ahKAJ26H3apl5Jbh+I4difvFRETwe6ABZRYEH13qW
x0NstZBcJ0BfzoBuYvylekhRyrT8NddTbhrzOk5nz4xlJs36kZFXvLJnp+jpUyG2MYFQQo8ele/1
KiSB2a+F+sXrgEArgJJ0FZlC5aB2cm6AlmQc6DcPltZBtUBayaaKyEHCaoS6hZmv0lS/EEd2hee4
m5eGtQkOuRqY007HLj4b0SgBs4xEWRuCyX3D4y2eIayAhXqKRk1ynlepL69WJE+0j7nP7lbOXFnV
bxeR3HVljf289QzPXPP+ZLsvixtjgw0gQPRqH+YbMZyyqEJmsSx1yTHvH+OxeLVV/3l3aXL+fkVy
5rwBzcipRrRj+ndwgNbRWsdCYp62b218Kbdj/c69n0io9QzFywakAhc98Iioqy8CuDFkMCToCiMn
phJPwftGczMWnqZ7YoWxDM6GR5aqNq/tMYT3SJ6owFlFQzZvON/v/LnoNKtoIDAqTOyVQ6igAt98
WHoW7P4KvFTqDqvbMEznzf+Sa+ymjt5vmug8YZSoDJN2JCw56TJVOYyoG/laEvLIjeBwXss6bz3O
AkEQuwkdIjHSdO9pfp0IRjSCFtxRn3xGMfEYInQW1462bJrFOkfKDSlb/PpPTrljBQ4UtkP1l1Jg
NUvVxAHRWp6/i5/DafeG0NzTmC2fiALEZpBn20yOvF8MOnsiMBMLtGpCbPZJbq6BQUAqxpJ6+d9S
OW4oE+l8SBaKzCOHQTJRXqrrpWbwbRq/DugHL8+7KMxN6N67I9YaHL0MuYn/ZfXIRFDBAVF4P57u
sl7JJMKZyrcy9kztCXLcAw/iLt4LZE6hUPvRaRuEGfJZw3JfN0CTLhgxbpnulWVArI15sDYQCqTI
Ht2yTAjO4u/4ZiQXlm4oIL7sQOUvB0OpG7528CfZMHYbI9NxSwTocqdjeqriT+28ps8VRt7a55B3
XDAZSg2dXHSAp29mQtZapm7BrMM1WbOSgl8vQtkZAk6XJlUPyZ4CuYLbCbyhyH72eV6ujLBXsK9O
eo4X1f2RWXNWQmkncb6miSejF50aRgRb037kUKWdDaYy7eUB0f0eGwO66/DScMOdsaNC8yij0CjZ
lFlYPMBlo7R/pabN4s4fY824/52N//wZYvIIMPC3C3e8dvgB8EjgdmwABfpR8/ODP6QgG2edkF3d
JeUfzTX90W6u7YPdz/5q7rarcooe1NaHR37ShK2r0NwmJjM/CoifCG0pCM/3aidtQtffwES2/8V7
BPuZXp5EGt1v5PLNASU4oS6tiDqkN5t7/aHybZpsEr7J29QKYKtNbdCK0j6KW0sH4xEJqdlqY8/1
PDL4INH/rzwDAYVTj8bsQScXHJJoeQ3JNzYfrErelxICnXHq5njZ8pgQ7BqUNnh/mDxen85Gnvbk
fAk23zgV8aHmrgb23lTbNWoY/TuT+cRm+7nPAcQ6U9oe+ECPXlnSEqSZ5nM72ac30RiooFfk5qJ1
qVe0CBz9oUHTnPwGyCJA1O1yiPDiKEZQYhR7LUQflm+3I5EDDD/SvWyRt91kYEyzDmN5g08wBkmf
S6hp5BVG3H3dNfjb+uJVCo7U2LM57B6Fz5iGaqIeF3GqlLDKKocnQrXETZceSokJGsobTiBvm2fS
kbT2WS96lqETEco91IdJN6fKDsyclWvZdCrZKv1f3RHmRGfW/2ch3nLIH5y1dHgkVyPZJQNVvPjw
k0NPE3q4h5vBj0cJmzKG9H3kgji6bKnJLZ3kw2934/sjXajoRvGwD3CIMBkGO0zTAuoeeBqW6pPb
XKHN1VTTMoizNoUaCvj1achvIHAscfU3wmDcM5Jf6l48cfFxK8fsQgJaCCkkSEza85AcaK/Jfwsq
H96lWQecpY49JXrhT5A7njyOcMcuvoduCkkrfEvK1Fa9+XuEpPKTBbqWIaVUfKKmK4mIFU0X7jEG
Zoq5W94fL5+vuRpgCzsyC24oF4lt1tUbT2+Vq1MkARxOeDC2PnmJKROIlVPB0B/lf/opz4+Rm79d
HiXb5Onxn0SJF+xpqF69Y1GIMKg4VQQdABX/VhwLtHUVw/6eXoAcspefQkLdCd3fTICzRsLHt5RK
C01lJb/GVoOWUyTt/WgUfbJCfn98e8x/553HuhYJrVe9ZC7uLO8h6ybuS7LargGk9Rt5S2VPN5T+
qbMjKwcZ/cWPtbO6JXg9L+IEdV5gh9lwuJNKLFG7ngT+O5N1mwfaBrw3D/5MNAsu60SzuMntGpMc
e8LsBw2TsCzO3zTRk5nqQEM6bpiWgRHccvnBfaFZW8b6kfs3225Xa35hVxofVtAnGF59O4VqSNCx
ATB39ByQSl5klk/I7gOBDCOaY6g9NzbIFreTBtCGHYrP+HdndwN9tW2QaZ6pTRD97fiWTSiNBbfu
v0b6K20wZEaSz3rhTD1PPFrh5eEHbq4oPFkCbkmwfxDeRiszmdoHfmlUw/7VzeNBQ22iLPNxYieJ
LVjrhzKUWtvvMZ8xEb/hFUPlb2DZ/MwcnDjf2kLLWjh5wCHqOzq4qAkFUs+Y6xpJ84S370GHJNN/
JsYKvVJQKMID5Lj0a0qs6P8wElhNFlTG1oTCpa4xUtWAHNSvDUewH63hpoaiHRjA2AJWEHG/CvSD
WGmU5Hws8cCWDDr1XV3eWYKb1XBa3EPD8BwaPLC4XcZYho9tMZdEgWwHAu4IjiwJdxsNe8gSk8X6
5oJhELpkmpRMoiV9wsGZqMj+eS9WcGabFi9kdyPZGSFBQ6UNCSvbTQaOySQe0g0+DhCjKSqv2QJF
lWxc/XZgKFA/iVkP16TdeMqkJXwjBCHZYIFP+6Ph4yLTXTT3L7fLX7FDZMM1YlewFsWRN7lo6IYj
ERc6zXYzvKGf1dk2J+bUQ9m0z7J6lFbOneqUYNkRJSApttwgni3mh0nNSc2w5t415/MpvEIe0ttC
7QAI9snixLYDtmpJlClFrlPwuWCZzHxJ1HpdgtSeIk1i4scsCtyh27fXheY82zRJ48UZ23uy8xNW
8a093d0yf845r6hnXnKZH9VaOocikt7m32QFV7cNiKeWGvGF1/P9SqN0NC07oZFfSzfMMVal/Qhb
1rK4ggOse6aWUXFkVe14YMj0mOOlRQcusxZ+0d8xggraA80lRiwOXCLNZqDfWBi8a7rpDr4daAZO
2Iyaqcu3OsBUwwhv8o3nmIsUQuGnq0MhB1sEbHd/DuX/mlsMk2UR2Xkb0+XuHVvJGK6VUCPGUDZz
nOcgSk562Uuete7dpLaVx4QF9Y7nJCshmaVbWhxh5Ht51oGUu6tRChYxVaRAvVxr/HV09lT3FygM
nc8mCGN/8SoFWAkESfdAMKVoBY2MyOhPhaRNFU5pCUleZlmBnOKTWbCZ1iVWx1vymJncrGvzUseZ
8S5AgJD1CBIdp/yF5p9RsED1z+xylDVV26U8lAmG03juJUiY4QlxoYyqhf8srGPAV0FxZmhroEsw
8nBtEVVOjbZKmuckNfZrpN/W/1UUjKn99gqKQ3jSxJpuGSZH+sULOysBuQhKCYk64QA2PppsTnSi
5m41p1HeqC1YwPs1+NwnMS199lZL3ek9yJ3ke+5iITjNFvmwDiKPPLBkBqs7FPj9e6/R7CLuDNVi
3ayfvB7Hc3XKJ7c/J381aocFMTMi3r0gRRPxOsflFcPk4rNDa/xBMZF/KCOHTTkyh2bVDTSbqP/y
4yJfDTm1ymDTKE5fkk7CiD5grGeywLV62dMiX+L/cUZKeqMVznd/RHI1a/dEw/UkTI3GvVSWGdC+
C7XxxCNB00xMwRN/enJiDHNFcRnEtR8F4yvXQgUUNN3mbi8y3iVLPFuDBSTZpcsBm8LayCFxK/rR
4g9N3aRoULTllCWaEY6LTMHWDUF90hFfhNxzukzfEqQin47IETqxRF4P/sjGTu37w4dvMQ4DQ/H8
rryJ3RcYDKVFCLB0knYezoNRsVmsM4F++Cn0k5tn9iXCkksH/dy0iIZWHegDdNGfl+6dGwtx0RMG
h1vMMzGB3LCrPPHZvKBkgNewNmA/XQL+UeZs28LPL3OBju6NeG1rHST2Mc0PantFjC6zC62/tphU
yVj66Z9Vik60F3IekVWB8tTX5YQNu1A7/QOFgplsJKYL8+rzo15IBNLIrVFhEScpm2wZngMCOmRC
8tCWWbdBVav8myUSjqf7zX+Jn8M02Zb2A5uwhG5B4ZGHjBdwN56WZ51OhMwXel4eR9ldjN9u5XX6
PAm5y2cIuyzWYyxSUf3LlAoWQw3rx09grtMuvFdZzNPjF9G3YiV0bSJStib6MyWAxp+3H2UEc3t6
Wc4/N22X8PymVKUXgugiBiMeAYgw31rWR/DyGT8GLY6YFqiA6N6UQ6VAx9E9RKFICS0h3WHqAre/
3hvoeIfGFZMuyGYShc81PqOMFsklBQDmtS6y6LWfkGoHXlg5TTTiLS0QjxOeYpQMI5yOiYIQYran
WPsphZN+LnS8YwG2Xukj5QW6HDz+66dVL8PNlNvJd8cDuoDaXvsxEipRRZcuX+9m6rX1uvkf56J5
6VEOmw9ri/3Uhv6flzHG9qKeE8YeGHHX+kuSo6HKqMEZ+C4Lr+BbMNdYhMwdAzWI6z98vKxx5PjF
O2jgCzrlQOFXXg5k2buujuF6/pAgaBWTLjmGcqzm2DAw/v3b5/HBnZFw8t7/ssfh57PKoYtFs0oS
lAK8rGYKQhBFr7AycYEmn6xsuZkeig1Prsm8AGakAMrt5uAFFcX35Y4VfZVvYOSoNC2vG3Zpsuz9
G+1wBbhXK+oMX6noSh5UZU2ftqk+En5waodlTvQxHjZF/TV1IfQzgrdR7r9DQGpT1WAMlm8p8G+x
3bcWZuETi9rvw+qkqBOhgFare5QxO73N9Rwv4qevpYtu4eAJORdh5K6PkN8rCUyWFwOO9hCbo9rL
NOPAldRGHqBOUPJ5f5vqHzMOUvNui8qLgc0IgJS7oFA7cc5/6vBw9HD5XdWCUwYL93OMuC6N5c9Z
swrxO9ISrs27BUI8cqkeA7e6jc7ezEHGNt/MhC66yGHLzSxa6ohIRLXydR3CN9M/5xRunGHchU5x
TkYbpsjEJYQTjJg7Gqd/MxIiTf274Ox+hEwFN/bml5dLA45qIT/kMbBKffbvD4l8yqQWGj6bvpfF
MZqvTVITZ1iPgDQGGvO7NJVaN1nOXVkQQedgBLa3lMf/6e4HirVPBPtbQhInsSFQVofTTTc6R33q
qgEr5WBzr0+QQBROtWN+kWo8TsiGgpspjupYpxAQ6bgzMApNJMup9RzaQOiTWV+2NQN3vCR05f7p
6SrnYjDINwWM6NOAvgX7me7Z4+3jnvVMavjEsg6vOM1v379mx6EGaiYhPr6tMkbrs8k03/Mgaw3e
Eb5bIzzhUs42rnq9ORz9uIypoMcWQaDS13B69mTWwOCdiWJvP2P3Nj8KgW74iUEFdofFIPZOAMko
ySyfVMfoV4LL/xmGw6iTV718bohLTVooRRA03PzxPXZyw1/P6xmhZova2pLNdwa1Bn7p/BRqDymV
7634WnctBrs5dU8RcsrGAYHPU2APbat56QlwfzjmECFAJba53ERbMHqNffGjWKKUmdl7RHgaL/JM
rYeCJXpbDitni6Psp04jq8Y2nIrIVf/Cke9VkiLRMegCRmd1PErJ6eqgpSGukVgfmR//cRPSpDDn
dOXrMjJQLOXClcxMk06AcgB8KPQuso/Hg54uIG7grompRvCL2NabqrDAc6URLQZ+4tWIxdGrSKLV
jMcIxEVDeQ6mrpmeVA+Zpp8CowN1GpIq6MOHuZUPpriqy3e28gTx6ejfLXmrdmJLwG746sV/VVFf
WAMwArRi2VG2R5yQhK7OF90LPGoYNz9RmL0eQleRg10kSEQUUVlZ0bz1bDQ8a+sFZv/v93gTZnz1
fgQ+kZvnwre/0XIk5hjr8KLZ87Mba2eyPTpnsMr1hv6yd53uuhImzK3cVNrsphFlfZBasgRnFfY8
YhhKuuEPnPpjwAkfampBEESpg/NZQm9bNbvyJ8dxgYbzf03TcCH1W3GorjoY+Gu80ofPnPlK31KO
cFHRtKPFS+KQl/zg9uw5koh1kZtlqeXQbL5BJjqYnUGu9NWZlZmOYGbIoDCpTB0Boc9oboYIfLfv
vp2q2fD8SoXHXqQzV+kdi8M/U139kO1WfeznxuMDODnDkGdLZQxkh4e2QnJsJ1c3pqiR+UA6GQyN
RzPFD942cBmtn1uQzgkuAe/s/kyJRpf7Ja4OmkSH5sKQTkmS/E01kCv2cOVldeU6mpbsYj2WZOoW
eAS+o3jCuvG5CIid4AkFiXsDpsgJQwKTnHZDNXJ8B2xQ/uz7xKowReJRP1f83YGdexBgm9/EOCiA
cbHJqrp7f1se91MAdPnGaEGm8HAq2pA48CwGaIcmsDNiJK2tAvK2gGtKTOMf6Ta7Ms6RNyTyibgv
fzIEVGEwAE+gRr3hntOsONiT1Un4VUD5itqfAfufGyVkrgfGzIk954esSsefEA353XXezO8Skh9V
dLUBvXWWa7RDg6EZpKcxwCf5+HvpyCesCwTFFR2jXEWpWr2uFN4r9LLyd39KI9fsqZ9VwUuZp5IM
BA+Nsp+ZjESJ1+oBqajD5hFSFqUv8BkA0BQU6X1raoJVplMUVUYj7oG1QSDmlVszwD+RFzHQl/jK
g5bDd86B2b3f8Y6wlftoTO9RuoznmcV/io9ufo9/kG6rz5KXXnKoKIHfwdddbV5i8ibCDtLDaEQw
C+aadtywcgPAnZ9F+JA4UiEHjVlqIJFPTPWXlpwlcIHFNA/Kihupr0DQKDhzcqUDv4Y1VTjlWhRD
Gd9L+cEGxVLXeH6a9fMY1+jndNDRHfcrnH4ary/6O86DRePaZ+oGIb39ImnjwOadbLgzn6EKnapa
8KaAP63+WNQ3BPXdixXfUi3K7jFarTvYbNSWJF402+afu+3tJV1IAPiENxysKx1dtRelX6tEQl07
m39kuYF0rWMeesUuuJyzD4t37gyG1FrF4MsKv2vgTiE08RRrzdZP1pYwq8cYOvlZuMM5qHjJD71+
C5Xwd5CPzq559ihixWDp3WiY246Ypt4eR58gBLSEAkQ4wE7sSu0Wxnyima5jh9CW8HXZOgTUNki7
Li47O6WJ5PO9igaOP9YVPE7GGR3l0BkpwidjndEWIiRuTOV2D/q0zvnkbdqbm++hznNL2ETmjndA
6j21KNcxnsYsUsTn/eJlEKArCaRO3E9718l0OA5hWMYhlhSt9IkOt0Cci6njqEoGew7yHdGZue1v
FvRcjQJnHo8QFFz32xMiDlwCLzSTt5As5/4Io5ElLCvjzcRWD3INhjoaMIC3uS4qYz8rsyq5Bu0y
iqqY5boGtfx8gSrqFWSWm6xcGgk/dPMVdeev8h71YrQWF7jRohUQur4oOHAIWzNsnJ+7Eh52cq93
4kSTVQWwz4rYeuB14iWVpvl1z+Fa0xIFCoUMpcsWFozOdvMKB5jhshyAgDBp0v8fZrYq+iceyJMN
JC0WybiQGVwEHkL2ciqYaWy1sajlnmG6ASI855WjGCAC6pEDLMmDBFuj/jqIYZcRMKKruis/BWEK
7DsbWO87cj3az6v4HuhAYpC1JA0n0Yz6JmzzhOrtsttQfUng9rzRD/G48oEI0dBjRf1QhE7I2zfY
eMU2OESkt8BL6XRRFhOXsTNl7uZFgh1Zlr5yscDewzazzDOjzl8f+SiojZmx4tH5WTdCHsbwASlo
8Dx/fo5yVsjlrY+ynBjfVpNEfkOm+idKHb9YZu9y8KBJxhcR6ZNMQjJBpgS1gNl+1kfFJQTiN341
E9eRx6xgXfrd4171S0VOSCHqxQiscXir5fc2ZOq8lNcrYRVCZxOqSFcHBDDX27AXh/QKEChu1vG9
qrCFNT7NSTrrJJGwPgjmhq1M0jYjj6dPFz0v5DPE7Kfzc1iswIGuyowhpwjj7XaNtpNhgyi9lhOm
HyRoz3M2DuaZbk4Bz3WmAVaAiKIKTCt9dRieNIgryIXZlON6KiQPQf8YwKgWWTa5SPsoTQNeQr78
c0HOoYrZR6L9Kmdxl//84SOREBj3Z1VnP1uwfRmcMlySeNboWNRvq5wnmQGhWhD9d6lL1tL8njB9
5ByNb7u8ci7Pnw8wCfG8jts2NDwP7cMlkFW6BFRjrqGLc4QC9GjdUEvCh8MIBEHTOdMaGRBSC1RL
LOzuncGu0SPJSZnpE9vxU0JclL/HnMo4miwoqWAaPr+L5XjYKG3o52swJfgoVfsxRnFalU9kbuLz
gxQEWVvGqilR2uzE5cW2Ngv3u3D215schout/RmzWMk0vnyEAvW886pZUFwRQaQi+kcEd3Rqx4Er
rxHBUjyg5gnEqH57t4jh06RER5QyiCHqklkfiho/x+E5rxl/CFidEl4QyBdUZifCTxTcC4qqDzWl
7dsXlYK2EdR0+QNB88DIoBK643woe8YT3GdodPxcsFbs9J30icmrw+NpEOjk2R7VqpCV1jhxaiB0
QM+qhuqAwQ46/dE2dUd4DBOYmmopS6w/AMdgtvv/kSTlax3mnoQsYTpuQTqwzbvVsotweCZW/Ye3
NCpuDthf3udihzuWx/HlgvNzXeRUvROxjpr2ZNsow+rPHA9FsuWbDE3+U/SLGSNuwt/IC8VphIfH
GV0j5HTxj5B557kruf2CuhB5thjIJ7W+Cc5RFGnctGH8vqcBGd1elYdQwbt1+AQv091+F95ESj3n
EiSqiSKmkm8bSDVXh0z5KQ/XvYuzdpQXjo67FyipJoqTc8JIp39wDsbllpYmbIFbjpMmNDBUH3yy
jwJVMnth9R2O4VcNs7j4lzl/1W12mfPvzJqYG9UwflulgshkzQIdYmcgXEtdbnbQLyhw46ASwhiF
BlyMdqSPRIoE+Jl1fUU09bMwp+G6Ma23T/FwTbA6eyQH/RM/NbGh5Y2TOGwnMi2fsa9xFfXOkbfv
Xw62tv0g0B5A7gKASTuTzBjFHQUIGW5s1z2mbOwB8Z/kLbB+Bw+OiDRYgIzCrVUCGZT4tdM3no/+
vwQZG7GAIe41NtmNYxuEqvVqi0zZycIHJB7FXhnjCMGqi1TLu+g+IYfAqoyK1r4l6Y8xNcdsl0n+
pT3OQ7PYWeaMj4WZQ0h71+pT8ExbfHuKx4s52lWz/9i3202x5V6ttby4pIc2D6QwdhrEI9efq9Q2
lvrN+FiDG0MeZfY51/P39xwbx6WUjrswVtqIarr7Eg3RdTTtXZLKBoFDVpU/mIabZigAGeuRpVVu
BvW6aEBomTC+FBfyaeQMY2Q8OqmeDL69zzIvJbSXL9rWrPcZ9STZhKGFACtH3ZPwYgFLnSieG1Uk
3sMc8Z2ZBTabDyKDzQbuxCZShNvr9gYP+MkY+8Wcs96eciPLfjZtVycB4K3bfmuA8FsMhAWYzlcb
TOcRwcjzddUy3NdcWx7xxSW/DHgCFsvceo3T2myAeUOtULMAAvp4WE4jUrdWTtHx/7MAVXXufKZ5
YpEeoDDyTJMySCj9GkilkxuAZ94agQ/DpvJtiNUIDyVwgJNr6he8kvc3PTTgnyL0N5t/uO40XIe/
RZk2NEBStnHPvuIpBLnWm+2v23u0NxBwRPl8+R+9rIs3FD07ZhtkSViyvP8pEucRu/q7gjr4lQUu
vLIDzE8OnEDOpxnA+tJfAQEO4k+X2I9QEEA9+m/mbllXdpnAsRyfTcDcW3g4qgr1zkl3ApJOBubf
r+lXNeuPA/VvzOJl7aqOuO5eKg332y0DuOyI3qRd65STLPV6Dxd2F71AuFFwNX2afJW7DtBcCTUD
0Z3uteK2Z+3jPRGdY3UMwR+l5pO0Wwnf6+ht77TBisI3isU/1S1MVTTm0lTAZ02IIL3f7oNl1vae
hUrLVc9gLB7D75odwwdXo3aZzkCYUxZmtMBcu/zHqvvhOFLwBDMk4QokKAhn/0rw+42hvjr+WeGO
aoy9COT4E5SnMeUxDYnL8+fhr+KeUVPgDNuDvbnkq5/R7eL3yAjLtq6DB7k0yY3EeS13nNnmQY9Y
Tou/cpW0eOYYMQUx9sE3Jau4sESVLTkHqEE7SKGZWw2cH2v1hFNmKeIkJdjlS49dRnH8lTQVYUmA
0dJQRWnB99nJiRr4cYhYxl/eP9Z11a4qVWpio8XSxloCItvsUCMKdteQpBWJP+jRpkCDPkkW5W2w
nkytXcAnvFkhvt/hTxPbJfQcURFRx86dUjOI9hR9Pn9ywEYBO6kjxtZEeSDGsLqRYY+WuXdtn50d
rAJH8J0zoFemfNTvaukfoJ0VWrClCb897GEJNJtumd33W6vUV9+aj98jppeBvfEDsku+Bq3/etdl
Up1Xe5JvY9Ap1EFqN//XYLxXKn1IbKoWcVLGbmwIl0T1R412I7X8GsbnpuN8NV6duTazivEOAByH
SMzRMV9LH76+9AzGRMD3pRefuOD7sRKkaeUOIGaotFh2Ypm3JezAW5k4o4ybw8MVXTEKvc7WFNWH
vE5+c3XoIkBjTmvHWALQvGiN96x4QaPvildTR6SjnB65q7XXKHLwcAMwz4iqg58WQij+rKxwep0B
Jgvynz6ybfOqIY6UDiPZYrwYOyFVMDN2q1qc77mldAdoFZ95fJIi9cLWEqPAsaphKVDZIHn6YvGJ
TofBEvDaDut//RKXT5uM4eLBUEWu23UJATeVQ9EVVCkxgEkNVB7bWsyauaeSU/UmIrTEzQnmbH0H
tLZU5pRkWAguc365A61av+ZveRq8URZV/mupBgweDxFEpM7yEDFWF3lgOddDrAx5xY/r9vhf/IMJ
/rvjx/HCzPCA126C0jt0fpY5diNoEqkkZzpro5KBJV1+KVFI3yio6fqa9V0R+pnmLNG4vZ21PfKn
o6A+2ms5mSmFRpx1NItPVlIejUIzRM2cWi/AgD32B8XhG4BFm5f0cPA2ecAzOftvUZMYnShR6BIy
hSWPC9+cbKgsm+XiPFSfIMuRzkkI712IB11FNq2xm01FJ8DWdljJpQeu0bY35IVDhpGehCTQFyUF
tr1NeorTdUl4kbUnUUENZLoGtvBhSV5GNzvDFJA7dyP80cLusPDitCQeKiPKZC8tTreSZ42Ae/FG
p1KaTvuKdKrCsNKja9WZ6ixfBpTerU0mZ87xV3jb6UXoLI94gfk1E9ClehvuaA0zEoWgea7hl5EY
14XVKgAlyyvgkHOQUsWMt0IssYOQuaxS2DW/Vv8Y6TYb6zSNZ/pEkwQkcZJkYwn1cVUqJxk1mX+T
l4iAKMBzgUsMNNvTuEbNrlOoi5iL7ivSu4xVJ/rYLTneirP73NQV2RdK8s7jlXMy7MyNIGh6QGZE
GLp3qEjahtuDYu1ys4AQj7lzUsCIwgcUqJl6jtaKRbITKEEabFy+G8SmLZ0IofSIll5Gbl7jJxIH
BvQV49Xx7K5R9UQjRdopVLkOuqLOGBBh6fKMyYl7wkytwWAUAbJaAGME6K41Cozzn3G3YgouPNLo
gcW6ZXcEktgwBz5pxB+aW7at4cx6bMhFcanfBkjR0tTaKz8J9KrwvJYhjMiAaXaBjkdRYwimcwYZ
GbmfQ4KfEpEet6R3TCRPkF824FBmG3jxLz0OYxhv1yEwvwpPBKjMuuFjmzzvgWa436bdlr47Iexy
63c43sd2FusLBPZNNSRmYpBCAwCWISaV7TvJgDdsqCo4iG6ESmaKzWjtoh/xnVXKJvSLubKrCV47
d37aVMF80mJdwfv3DBleLykNMOvWgZxiP0lzd563qTeZYLteSPk+mym5O8JYIaisghgXf0AicVas
jHQoQuAPRtgnfQqUCFG/mBlz0eHTBTeu3yGULrS6DUPMXgfwaPw4o8FxV3RpvjO8oMYBJCWv7Xt6
fgMCQgSW4GALuR19ZSdse4fQXoo4iP0pvXBk5AQepKsPcBqfJ6ngGu6IsJaYW0hsuT03AXu8SMrY
quBCXHuz3DoBxcdkpt9Mo2/ygq3PTmPMRVg9Mv8QQlbTAncptHXT4AYraMG4NV0go97myubQxX1y
zkb0zCb6yUOa1vK1YbWgvE2iA4XoNhzZUVOeyof0uhExKyS0EfoH+dSA7tqg8kAr9pE9RtwihqcV
hPhbypm7sgNDU8LjTPhaE5Z6VYfNHzR8MLA9Tp0VFPCQD3/+xrlSEhkFa/N2eS+DE5CE8IbqCScO
0KUYh8fWqxJGrN0yKk7Bt63pRJTiNawG/Q0165UruW0p+EefZfUVJ8LH1uoclZHpWhjMaZWlSWCZ
2DBLwFkGpOVmUamGHxlkpaVF5Q4ZpbAUtnR9t0o89hf8BkXToE/QWHXJTLOu2pGiHmc3h+wQCbmH
MruvlJAoggcvTgJXZyd3PHMbmS/2OmlpJs/wW82L9DxuqukqWtGyPHKcFdyAWo4YUbtABH4rObVs
eMbEagCB6tk/be/CJX8YqbO7qvMIaHtyhDJtI7vhh9cjLXJ9pgCZ00t3JfaDt2zG9fcTTVylWZTl
hb2KamaFyKtNsqdWISJ1DqhIZhIuDvqGzxZkYTgbx6Ej0lRKCprLRy2HmtPBIQha2tc5IjaPZHGR
mZKwAPL4vBp8j9sHe86N2CfcGAv3pg3rkcxo5b80BqoZK7Sfb5P+toTHhoXJyA2LI6aCgWb+LgDL
x80wDsTbfH0r1EKK4upX29AfVhrjcI2pL/psd4b+GnkB0HkMDvL7h8JQDQfUhVbFXa5ggiXc57zM
2R/k3uD7TUr+tCA+hLQ5K7+qIxpH+VXhg2D4c44hkXdG4wdUEvssU78bu1BnOCVfQp5Abhiwo2fi
Cygeb4cjlWoWFGcQa0vjk5OxMi6DKo5/hd5CMSmMmy6UFAix0TV3HscvkahX2nmaRIvBHcNG3kp5
athOXkM4DZUmM/wXGFXQnoe4iOQIrtAU4skoXnGct9xKGvGkntoDRBh1JBdHHXa8uBgaQfT7cyLt
qLr3C+cmBPQWL86qmSIcRuHL1c/NaO17rHozq5VZVAbXt013Qedid5F9fBNjiZC70wzty/X2hjrC
dvAYgQl+W9bR8Q4ugwXuCtyGg8mPeqiuvLFBzcL1qeQc+QoOSlwChN+r5a8MQ++bOR24a48HBmVp
I99puJ+vPcK1jIodLSFNJ+n4hlZ3Nk2JgipKhao7R7alVZa1hgKc4Wn0HXiA3UHjpIWL3Rj5az3s
u9CMKDSx3kVGAC+weSvKJyOlgRD3G/5QQiXLgKVIJJddajpW4brP1Qy1WkN+i0viRxa6D9PRpncQ
aKqrHa1Z3gUD4NDSNedbfLuPaVv/nGTJZJe4C7HdhQmaY0X9YETH26q0ZzJhnh9aSNIej/6y1jxh
fOiu/uur5tn4zPjQfS+whqu0sP9Om0PT5NYZPcaqt4NRkhdXsA6/t2hopPzA0vunZze9vMRfAFpx
4L8L4SPQcJBrrflNbqHj3lncnK5JObT/BPMuzmDZ0GeXHxpNhxzfgCG9vemaxvBRfzaNvJ8n+NJX
etEJ6Ko0/anWtEgrEuO3WfVu0+nEVSeTUT3QSBWLIg6WFPq2Y0McdKN1GEeaFpgWDZ97wSzWibaZ
eEr9zX9velrJR1rYssmU7zrdfsevaolxk2SSNmZAnea6hQCkZm05GlHrXQMNS4YNTMu9rGn2FzZI
PZT2vBFtQccjLTOdF8HbsA2U5wHrIWHcrA2RrZWVbKgS+sWq73Aan4QSR5cUFk4ZfnV+/fHHg2t/
Cjhi8Kz4raanmKTzH2FHz7AXGAgN2kP3YXTQuu/FrV9hhRI2muCyqTwU9jmAgucbZkZkbeun1sLZ
1de2SOaHoPGjoNDFObwLBpIZKf2b54CS65H8VE4BmLhFqOwcM/gnsCl7K006O6SB/vw1hWipb7Cy
L7+mx4thgjIvB/JJ1ikBwjElNEqkJyNSm+KuTXO7unGqXUs3zpbfvZhcGIeEtNBn30dQYOFEjkmc
P9znlgaoROxvAfIe0dhrTFand3iyUvm0GNfrYPD8n5UcVDqLnv/9JvmdD7QmnC5xl8fthm6Ped8T
cdXB+0u/DVx8M/w7aETUktYamli4EXHWV2MDdd4IPG/3+meIOsD7QWrkrIBtftbPBCY+abaXD7k5
ksxNNdKMFQskFvcOPX15lXS6Vd5MaSIjmRo4qdZvmkrjBdHtdfkhduJVovGGffQFyIFddG0/vN8J
SAXU1aifDqFchPLQT7Y/wHRoHxoyHur1vR3hSs8TfMxTLhZhqxjCrrEP4XSYQMUPxIbZVW+6FyAU
9V9XaMW42bcQm3PFwHFoEAPS19alkUsTkdNQbLBCja3wV3hkvLmxF9iG/QHIAVCDeMhDvZjw/5Ds
D3J+/Ke1RgBjLlo+uXmcASCeL+XbAO9rU/ClGuZhGsbuBKYkUbYp9J9cIh0NOjs55OZDjz7j4bUc
B0SA6f+ic4MoSIzWEVfXkYQPgMw4XYKcccEvN67vEgbKIodd0KbZ3SPHhXYsMU/Ey3gun5rZUttO
OWhUg3REKhTYVrtFQxC1GBqzQDKCRuDXpb36PT0lT65YSpGm3qumCI/RN9sEoKuLYnVk+6WJWlg/
p9iU7McHyH9zFHtM2SyfezaoxvbUUKhvtzywMTxQ7rPXeukR5Vv2aucjfT4kET4rIOKEKhOG/TiS
ID0q6jVsTs7XOhnwhtV3b4e7ZMvwT3+B7uRBzFah7KflOtRbTAeFMi1XVAxyQYcOXbbVayKZ1vPd
IXqceyF5Nz7340BhXwA9A2gTJW8c5inLrmwPkPyeZKEyVQIp3BsVAJAmlbgahK6ETJZKvR8p8mhN
0PtoLa8WyuYp5Ec3hQPiPu1Ib1FPbtvI4e9yqFyu0LBSOWG+698UFcLHQYxUzDUxnbtCWlGMCsVq
dsVBuJ+545gx7Kt34lT//Ik0UaWCJx2jJm55xGdNGxwxyO72KGbr8II49VVkfCgod0QZPB0rN4PA
C7oSHDA2jSPvdYNTyI2qE1VAynWnMwI7GsFHFfxQ59x3b8ORL9n2G8ITF/O6O3d5kEA66AFKSwK6
Ach78cAadK3VjL+8QqTRoSzmh273WdZS8Rg9pEbHGQ49Dh9I1lDfBlmEpkM/2qbOL7+fgqDWgxaG
kSX1zsEeWMRc7t0lOsXfehcOIX9Yt61OR7eqlL5OJvCfzdw5EfnMSpXZzgd4CzKLm74gPuhocOpg
NsxMTJzEL64nQZjN8rJjGx58JnIqIaC5GSCpyzncfrBVGH7GM4JziQC1OpXZYMIgH29td96ECiN+
9dEjlUo0mlyfPp/K3KoXbUbAa/jOkU2Ww7OWTHmTHAH1I7JhzlQvuw0KtROI21asr3sDt5CdsHXl
XYyMa3lQMyiftk613nPHFam9GqMwYV/yTRLiP9jXU5+NPVAjaYVWQupIzg9Ri2cFT4HbX6E4PtQp
DsuYaYtwKGor4SsScJYBsBlP3owJ2rRmIYMUjk8xXPVHxHte9O4b0sp34SfArq6dU/TZljrXlf9n
3sC0bukJyHGwojU8KWT9s8vALSYiTrBmxdZee6eHQ/5Svq4EjnHjjoJTfpyFVc+pL1IUmN6FFEVh
BfcmMuJTCWqCQSbcewoXsr5BJVUveVtRWn+lKGMVsE3XyKXf6ySGr5c7FV1Sj2Uaic1vWpyj/DJq
naFAOGcm/ODZrsRyKidee66zpbMeVmDtkpgEVl0RCCxoNrSDe6dsKSKPGtfZ7osrUCJCH46lzhkN
KiNlFeSSJcZT1YdDWj/tVgh1kAowEozXGALXTP+xTzkalaUURdsBQs9/v2UmeJvS2yG9SJ7R0TTl
6MaNiqQ4EJ/KYZvAJcCvJ8J2yCup817kPfiqj7HSEedHbuxDJKdpuh5l1xE6W//WKe5hdUu1RO8v
k6H1EG/SDcuELb1xFMp3xHSnV+Fhkk4nBqBZ9Fj7khmufJXiHIhIWyvS7SY5k5AI9e3DkXeeKmrd
fzQfOk1rKxiQqu0SH/RS8AJgQWJoFo5XZnB16yhptJgbG/iecyt+x1V7k7ZBulqMk8gx7qGsSmGH
htbeOe/969oxeSmXsHGwVP3CFQfsC9MAHqUZ7EDIfZtAZTAuPrsyrPBF1Z7BJhhZrn9Ih0s1XQuQ
mQdePd3oz65u4k3157SSPg70vIZnguFayG4g/qS1NAknq4CdFw3u03vlIJnc3XmaBJoHbGi509bs
ye1InTGITc63cFvAIsRDUzaLBEgpHROBPSQo7kEZRAZQjt7/cYzqOhDHtZdF+B+NV79C0RjRYo+N
4BsPlB9WuUlLS3gWCpyenYikPxsPIaaOsGBSKtNjykJu4yz9azGYhVv6XVr3Ps3lTGjyfGO+LkLA
BCIvK8N/tQryoOlaf55L6yJc+hRPerfF+XhXZbV0/3FPwvimeeR6qq1Hl+K2M6o2hO6HuKpSxBvp
PKElM+Q5J39xrtj6djElyuLgoEpaaiWsTx6m/SA3MTB7BinLMSucZt8dpWWF6rz7IfqdstSiIZSo
nUKKox6cwTr6LeAMoZNg6WSd2baozUXFQ6EPdtZl+rsDDypjOLW8b5c4TUq41MyiC/3LQ28uylXR
5g1M5aZ3SDgaaamtXJsoG+yyh2FY24JYmO2EOLqg8WItKyuhPGxIZ2FBWbkVnxPM2Robr1pOKCrn
bnTRP6BRhFDLW01H7hOAI1N1oSZkGNgfhDjB8wV0rK8YQlfdOtSm//e1QjC5gsZuPeRc3/rlFXu8
uDNjsTSnFUbv3m3wZI5P8lEQgtVUeNoi1TeinE/a2dVbNQMHUIdK/MdysAp3PFZKU955V3ntsU/h
DQ5dAOrigmAnjqOFkfaGupV/cEhnfkCBuSawaesEeV+xdgpzcvTFxYyFHEcvxHjnqvRjgGjQD13P
Or1FdpqDZd4fIWyYAInrddRQNKt39Qxe15bHZXq9NUPRYRfKxNt3avn15t7hJBbpJ0UHq5BK++rR
bMLRlNqdvmMtrUIqcW7nrcbhv+G2k/QABbK7POBr/yU/1WoNWfh86O+D4cV/HeahIRey434A7MXT
4PhGt3f/d9BvM6rKq9IZJ5+5jb6Ab40wqCEaCyA+YAVuWGCCCFCuaIka8qCjdZTKGDLCrAM/MjMl
aLvwfm84piJB7t7Y4tfGR9faEb0Vl+1feqik3jX8OnZ6nuIQi8gAZCjq3oaMX3CZYyAn92HMoJQ+
PFOWLkEtUE/gcdnevdwL0XNEutb7xaoCTiZzxK4+rxo+NXVg9qu7xq5cUeHTJpjliRhOh8dsy4gy
AO/i0mQGA2EyKNXN/492Ml6JctQOSGfTlKzd5jmfiAbtDY/vC9iJrNlgmGHe8l9egbPFZrRE8lAd
C5ldNb8oaMeAC5e6LmzSDMOWtYcN07z2mosn6h7IgmgMQncrFGU6MOYE2FjSZ9r8X1tOabH+zmk/
Hs3LhS4e52cQGY8YytPJOERY9KFbJZ3QOLo/we2lzd1SaWs5OGVfkFkgyp0Zyg89OuCZhpwrIhiy
oyxB7+Shgwm1OIFHwycfv96IpD6XsK/mGjZQKsF8Q3tjKitzFrG3iIdE/yPfMpORsXBw4TL42giu
qQVSAfq4XWLPibix8YsiBtuDmVkK8myFIOO10YNHeem6Chws3DhE++sV4PGx8vNAom0e4w9WtgHH
tYC6UirGqrPLmiIiDsMVaV7juYns6vghy3WILXr0h2FFqj7CGKlbSQA39B5P5DXy5bOvYJVBVdkW
PC5h1UOwWXgr/TNF+dTzXHcJAS/JKeqoJLsTdwChlBFmepUpGWyidOKsOX+K5HhGDlIhStZDv6og
llqOuSEbOPfKnd04LXhoufOpKKHNQIas1fVyF4T7IeoGLk/XuExoW2KePspt6eOHawUpVG6FkyZk
V5gtCD7pQOwMowyhCnOICXM+3/4IKyKCoGPgtQ51YQpv8Q3thTub8ubObXEhDgaizPwwDq8MO1Ow
AUgXrolmcsJGtyrQiNo/8mfXJRg6qZ60DT6LdK5b9vaD/Lj4Wh/G6iFzA7oo9CbP88kcOOHDZD1g
8DusoMxp8hXHx36+EG2zICxacwc76k/dwAqisJiG0/ji9j6nxNxu3fUp7Z/H3//m3U7Zdd03Ob0w
mbAr8KEmP3AFH/sjie/9jQGBxSsAjHImcDuBU+P5ZIjm/Xg0pyTYlBEhqFlVE0d9NTinAifzN3jg
d18G8ZE96QQ26gYYxbPysZhb9um5AnCj8k/n5pp7V+3GJnsM5C1l6xLJ2AJ0ctEBvB3HpQOSrYcw
FIyhfAiHU3i/yZ7G+ZAAzLHmsFQ9xyXcShAdmn3uKgNQhPQ0f5S5+kBF0iR0mfZmTCgr9zHafXgC
YUNcjRBRn/G3rQ3+SzWc4E7xn1Iks3DtGmDfALboKEbq/ZkI/pXbtB2cCQhuBG4agmxMOTeFnmth
jPr71fc+r7hDo4WadfOnerRFm5FQMq3RohOYQanMwecF7X8cBomWMEhyypDHQ20elZ8fRwIZ7Hxy
d9tab/G266SvhzpJ8yzf60Xdm3hqk69kLtJae7AP8jze+DNB6WYP14tgx+NlRrMwSNTc+PisZgtQ
cddHdYdrJzwBG2GOO4iKTDevcO9jwLUjfEJSfF0FwTP4tDzI1SzORf01eGIVu2UX+H8vO6KFgNgV
KyfSG1iMr7qK5hjh3hfAYE2wtJ6hjt+cxoWssZcjfjCy4nLmjMTgoUlvZfK9cyp7rLlsmSRpNlaY
mH6xM2z3t8O5JwSOoZFnpNKXuY96c6qSwyl6S+Rgl8Axc7vQuFVflYKzG8Ev/JIA8B17m8my79Yz
y6Ic3EBN9uZ16I1ZsolcAPUxuY5hOLpvIPKw7DZIpn/l1Q0DMEJYv1rlWI/uN0eiZ21Lq8vmibfx
Se3/tStqiUZlzWZEBHeXc+Xs9vR0NA/sAupoMlKZnJ+ziJNutfG43m5gfdK6tm+RqIx44jo9DVYs
X8EBDbWMOH6DC/2oNj5Km5HopGbQddf7a/dAIcV9tdCDTga4XPCxQcqJBS62k6A2O5dLy5fw77rn
QVOsSSYVmXqMKzc7tcdnpnxdIe7cL7ACGtwGi7kmSVfl7Gl+NtG5PDKQI9xxO3HULia+tKFi/rRy
mqzuBuwYlBi8sWz8MKSoUmn+IcuN9Bjlg+aYPUh4RhMAqCqK0eQa6ZyPpsyuovlLZSLmm0q3lde6
D08hoRErQw/hJGsQu4JbcNYnUjQc2Y4VIMV7BMu/D4kyhAtinp/vBi5Nq4sq+naDGjH4/IvWLxPE
/G75PPKjKWCSe/dy9UkJJtXQPg3dWsKRxtkyLBBCDo8FlBb2CBQd4NLRA4hB1XMGLzW9RmTdFB/8
u3SfR2zI5N76js0MltrzayTAU1MZwJDEtfbdAvComOZSmGzGx7eO1Zamj3jQ1GGe1Q0C2Co6LfRJ
3I3LvtJ9OekevCaZXD6kwKsTQGhSSts/pjWLV5+9cuU+jrnwBP25402cgZNw26ZnWRluFwmfKVOG
Ob4UURyBNjsnGz+PscrjLCWYnFgSPy3EI7+gEMPhqs8frL6PcKNcAuHdUcin5mesffeKxTNsPclh
T63nYbt1BDrnR+ZuneXfrqMwWAyQYZo+orj8wYJiXE9wF6G9z2e5sEhGCFZwDeX24R878g+wdCda
sPALyEVTJWg+gtJtrKRZUQqvIqfcMi+fMo4ooIW3hYXIjgxbHfknzV0b7EqRnfr28WWMsZNjMG1J
D8GcQF9aW5du9ueXKl+9A0tEm6ytNqqixo/KcVXVfeyiTbSrXVMLOaOCXEndfJ6KKLV6VEqHZEAZ
L48q+qrmLdr9VPbzktoEqyl3EAQGlHx327xISM89OmkcT4wFb+T7Vh3uTnjGQYaLCIb+jrAwWR6r
bY0j8gwYcVhdnzMrMn5Y3cpt6YLdn4T7yCvAJRI/M/cUUuyriVSU7SScvV9WRmi3FoOfs+E3GMPP
YoYLc4pbyLgbuj4it4JI0u/V2beQUqQPC8RNkoe5z61R/rdkOmos5lDh2ry50jcm2lv380uklsfP
+KN0Q2+ENXXvkMbK+s40YWDy8ANNCE4Im6F1hfdVHxXZgEn8Q1WOpxWv9nuj9rIYwRd2aJu3vTKg
zvWpYF2u435KYNZMHM48pLTq0Xq9eRe5OfYmm9vaQL78vd7VwB5FHTPylfh02Yakl5hXhSIKCQVC
DofL8Pmxx0CQHnJA6+ZlU1wopJdwWqhWpCT7gcY+fC5VLvM/Fl0CfjilNB+W2VS9WOpxn7wNBT/t
G9kbWAjxST1g3g8WDA4dI/VBEqZ7fLb+BFrcMANhJjEiJ+yUCdhNWSNC6rZbzv+m7Pgb/zHiekTF
IR8S1KxgbRbO9vNopJ7TMbDsv6InbFw9W0ShEu7ArDcUp5UQHomcz8MvAIEjmxq3pVK6vnUbjnNi
zG9RoMcAFo52FkV9hC+JwAOePVp2Kato5iECCMLJDRUwoD2lPh+Ard+WSZwTLEA0Cx3cYynQ6EtM
Hsn4TMBCqia7ThkZ7FvL+6dqi030zg6dVQP2nhxusj9e0g/KcBZ2PQfXxOYG+KtyGD1WHxD+2R5r
vbsin12ZVtt+dnL6Wunks1ahZcUsnd5bMNmdr8h/ULqOpidXZ70RSh4nZT9mzyYWRgzoUd+d4BGm
8Qh5BR25hAETaGrYZjTbb+PRefq4Btp9/BLeyqfR7yDa+wExDccLOA1PwjoaWYPnbJDVd4GbkdNa
Sy8dv0OlSeH0QVTyO5EY285/vHFfntyJ+2/hFncE7Qv7gApMYHGWK/5yVWLPfgF9bt9SuHeEh1hg
VK7O4O2qs1LQ3QmDUh0o2jh+fy46+RWMvP+S/S5ISmCny2n5hQnm4WRfbCBIC/XxK49NJM59zulf
g0fdNbXUdYZxZPaHzph9zX9I1qG+UPt6iBQGvXFIJKt5Ng2L1M4f9z9SLdK5ymwG9iVntBwhgQgi
ENefq/F4UvO3HvdrqFOOlcp23kVYM7kwefyONQ2XTZDiOJZzNHiUxwDluqflvGl3JSnH5eTKNPGa
fPXuHu/q38QEFOpnF2a8RJwNhWK8otaF1ju47cAQZIyPtBUY9g0sfA80w9Wrlye7fQkUFn35Ztxv
fzmt53/OLwqIOJFFrGGjHVwE/eJ/UdR5+PErICGppz+bee318fjrufJMPhihHBAzQIdAoLnsfJs9
JhIrr+N11NX5wc0dns6b/36GuWpZz/u6utOf4DGrxDM7D4gkH+nwKxqEP/zl8oJK4pDQXa0hi8tn
gmm1RMhuf5Ez8EkZk9rSJsEVAgVfabWujtannXSe5qZPy3VIIxyPsHzFvYuDAVHVLrd6naRXNEvs
jSIy8IVW+FgXV5w1Ph4boiQoNQjdokTirhAbu7Om+FFalrOfgW2SOG5AVSR+WgpPJGVn6Ac1GBQR
BuHdUP6Wck0dHp8FmR1GfMHfBafITTs6Dq9CiadI63cF6Qbnwl+9HNiZA1fhdVXaR/BGGiY9kBTf
CMrTi+MhDY4XQeHDPz3iFlnIGCmevHaUmNk3eEqkzK4hmmLZGptgf6yGvWMOfVhHm5s215HiYQ9J
+9HTWDmkdN0tMFz2ZErHuZQ6Z1/zo27/zA85SetYbueRpR4PX2Dhc6HEmmEQ7zRogDz4TYA+oPLP
b9tUCqVA+AeBWwCDv3/hIRQBch9YYu/LNYl441AxMSmCwaNKtIIM7gUKw5kJaf9Y7IBPUAflrTsv
2wk11+cWYIeRAMxxmBAhgE/iquhBFVQZLz+6nojDySkpML3c3Z0qeenBgWG2wG0sc6zTUiGLMC/f
F0U9yTMFYRjkMMTFz7FlzTSx+DYdoe4GRlD4VFPpHd5sseotMVbx9CXPd/bjySADl/ajn6EGiu+j
gltNFVcVQSWk1fc5el12lQSYmpXlzfFFy/7hTVP+J0zi2rvd+yu66FqAPeyYD9Iu9jDLMWImE3cp
JLhT4rbdhbEYc7GOp0j5dnNHTxZvBUZxe61GFYkyqX+v3Yv6SHo/vjQnLQYxJ/nyJ59lBYz0KXmX
frFiGuxGjkL97C+fzg5RwbAAJwVPN0UMBKYgvy1qlgrLDzibfGDYvf/0s/mKqeCewgbGEGQKqR0O
P3s6xPG90AN6sgpGmHhhUVQ9fVfVc2UIV/rRwRUGrUFsFPgfAgp8YBGIhp8TyYj63XFterlQeGjl
acaUv6E2r0Wdl+VVgCrBD33iyRrxMD7g4fePEwhg3OT+GA0+3doS9QJYe12xonkgfEsPM4GgvP+C
q4m6IZn4nwIs6OSau+vJX7WJvQGw/7qm25AUxagmJ3xhf8TbHKo1vNaiovU0QSkjGQgX2JEVMfFv
MUajsg0pqRligNjrmURx/+tjgHqg4MYa/9eh6IcXjdj4VK/h/J/yWythz4uzuOqeg8z2rVWwk3BN
G9J1KoPqUSq50tqQGB4Xg2NebUXj29VsTVvjBraJGw7KvKM7wJYXuD2LNSdRk6/q22CT/tR5fwZk
1SsVPxOoEhbE7YeRiH4YfPWfUt7M5u0595kwNor9Yh7JcHxUFRIkslLoij2Vrdn2pv8o+lHaW8Qd
cppqdv2fdtAZ06kDBrYZ5qQD8GUpJq0I8LeYXwwOZEDbkpA4GMGHuV+YiTzs86DhlowtlwnBzLFF
pJr4K/YZSeDh9uYFKe7n6zPh1Y5cCHB0vvxOoOSxZUUQTiLUPfCUNBBSbOx4jLgB0PTJi4P15e2Z
1SJxb0dG2VZIM7EV1aOdDwtFQQakPox9+rqqXk032DJRUIJ3KjqWOZD/L8bTLKxQ0NLzVvx8F6uY
tBuxl008gwdHT4MMLE+dLABmnws1ozTbGpO8pQE1iBlWYpUsmROtq9RcCJUmPNd9L6Z7r4bZqeVX
LbyFjYvVQJOTSYBVux1uLt6nQMdpuZPUakzxID/5B/RiEc5oSfRyzWY31vIu1NMz0ThSkg/GFUOx
x/fB0LhYbXQigfdUmmE4jhga8tN4ItPcXKGLhM1WI6t6XRlC6I5/A93yspO0ygovdZFUB8/0cYWb
aiHvA2WYnirxvZwxtmdrSEYlO4GPKz1LQJcg5sL6I1PC/d3nskVO2K8IJ1nJPCJpS4h/rAQ7aGkB
rhkU21pM17F+u9H5wgsezxGLvrPq3kax9EsFERpGBeFEay/Iw4bLRrqUryCyl1uLwPrjrbvWbv3W
pGp24s+ArWtL7KUGMgY7Ip5ddkWqfZdW0Wy6hXZ3cE63oFn+RcBLYCa4P2pnRLvbEuATtUBDxPyA
pA1szRkJy0lyWavwcRWwtoSbCmDI9dE3trwi0DS1dm8i8tSyAR1egxD+lPkNS5yeAVV9fXHPgR0F
0CFUzkuyEo45E5AVP681/DrbQfZtigYNqoXUBTUhUKzdnE4C4hP+MVEyu+Yr6hc0tfJ8JFjbuba0
n93VYId/gAapLe/QEswYfOh9owOwiF9yYHFWCZ6D4kJohUrC/AfofjwQdPlmXT6ktZbHJYMV3r0R
244a70RY/d9J/sMTHXkAwJv4KNVr+6036eRl9GK3FD7Yv9eesQL5qMdFLYSmhK578egGwUafj00L
bspx2MjWogKOgvDQNp7QyA2EopNG47RMkyADMCBrR4fZZC8KCxvAH3S3bwvGpUC8KVReuk2MKCqy
oMSEAt3WtB7NXL6SHb92knPW66v+OMstxyWOiKlxWUQz5Q4W/nXVv1jAC4c0YIxbOlbNyfvTzB+e
vsBIgopKInRecgnnLg4AAUUPP+mLASYs2hgG7lNKX/oRdFlIVLDLQQOONd+9X1WYEtBLOjxFz1oB
BzXOlnLmPHBXjDUjFrB/gNxjY+EoLUpJffpGhGfOY0tt9w0c5l7aj6IqwTFtg4RbK+uLNakUZW+d
YkM5tq/hUoAkuujavh2NOt9WMTeEDgftbah+tR81ZoHwu6GlsBqMDZ2X3UGV6+srfrS0Wn099mO7
lPL7x9iPFZDpVsGFCTIwRphda7YyaTqjT7nriyf4OGyUWJKyRdcRlLosstfyx3MozA/D+hqPeRh0
vtngfdAYtZNxybgHYzwf3Lh9OMgKB0NkPuj71Zd3zJhyu1Y0i5S33UT5a0tZ6qDuyOOdTtVKEZ6e
Eda04ceJ9lOaVH19YDRPX8lWICbHe91XGaWuQgibRo6qttPn9oUauDAQNEF/3Q0s7yYA2Iolreua
voC30v/WxFR8AXue9QXUwGD5HnlHNrBAZ19O+UjrqHnph1k2HcOu34c4e1UEgZrEhZA1LQngTf+h
7N0sBILb+XCo7eH11GILHMWdJDK4Ox+VuBnpwEyIWqim2NSWfvufb2jdy3w9dkSM4sLHLoUh1nPG
aYwKslnHw3gIFm7bSbP6tgBkoVXjXy83qddkSjR76H+7lZEV7XxrcAy72pCbLJh/Cw5vZg0uFUiI
018CY62aZ0ssN3RlPKozLXhN1T3f2K4D315KO+P/zwEN6R5QelL22treFfJE/5Kp9YZTeUGq/Jd+
Cg+Qm+dT6J5SBpxEQKNmbMxx3jTb2CSSLAn66eXtTYsGUT21KEuZ82f/0mtKa2arLotMhoyhSeXL
LYyZ9JfvEJ4RpPFh84jYBHUQ8+3XAMBPuuPt+c0NpX1ErgQX87Jzr+YXaAQKtkbL/ZkvpYm9/5Rg
f3gW6z5VIr8zq2WLwgtJXSIu5L1yH+bZcS3eNqRmS6srftyaUvy9Tg5BjjU1Uvf+jkxzRggxnPmE
Qt4MiuOougWZndyP5dlx8XbpJNrqCq25EGmB75OLcl3XGiczb8q6CEkWAGQUFKirnPJjuyynJ5K0
RALJ/HrSZDq4bqDK5nyIj3RlJRa4HjyOKwU2M55/BFrWQaD3H7VOuwmNwrv+SWxdUb+ODMYbVRXg
01tdF2k/AN507sircGWo7mXjFNHRYL6VCEWHlXxsAuP9GNwsD7iUyvUblZf985WUn+ZrTZ8g18Em
qKtxw5HrhX2R9FKB/VaclvX/muwa6GdmWJzleidicpKlN2LtfsBM3PDX/eVqCHRRnJTDExcbbnvJ
IbXTUSoeGdPhYzcy5cenOp2/6ljgb7ldIRvPBtkne9P974/EFsVlS16XzceB2DCWz+RSwkLlN1P2
JrfCvePchEpd4k5xj2qx+TKimJqjmhSkSal+VtahiagOvclzVqAkzU6SkxLk3UVo6SE+WmDbJb5C
oSjtC0xAXTEGsczvpdbnxTgboxjkp9VkgulGfFHe4zzYSVJUocTGssEPgeywVaxjRLNYn/YubZQg
aRMR+is9PttaC2hzRAepQH/H/AjQdG1zOUvNDIDcERSp/wMwVd4dpxT3QTEMY6Zdsh+3vax9wKFy
LWQkrrbya1HwNoKBs1i2SVi+6BWDOUC05BIQjtxISMrOcAUjMjZhLauQ/aBzvn36PX7nezxTjNLj
EepZRvW5XzIr2+Lj1404VOF6MdnLUiR8VcVijn2PVJcm45CR/mTjBhEDiH0mGpUovDAvv8VJZPgl
3JwhlpeOJbyZw6GBEOol27PDyDyRt84t4kUrtlBTWTRvRgY2Qa6nNEXQQ+qZdD+9HzhxUo+H4AJN
iC0L5uh/w/p5hnSR7+l5V1I8FmqV78+9CS21hAOO8718uIXQYZxsF9AwrUPN1XECkWzfdH0SfzD/
uQGwdr14fmb/Wxa7DFdUOyiAzHgk5CrSonZflOki8hWkCl9NlYhPNscQzl2ISZ3P7FHks6/zy9UQ
WSHeKK1bH9JJsSMQUdLsouP52R27+22SSAakgMYRy+Gll9jEsy0y7ntfi+tCPaHHpHfh+2mPAWPm
qwbkCDCWy/RG2ChjfDLSwIX+dM0KpQpVN9ICr+cFuCIRiEuzM4Ec7lF2X06DJrNp8/3aodNidF1w
nDovNksD7LyZvAyq7tEFhjSnWOoO+WVTQaCrOFOrDYksubTUnUWIgRmL/fWVC4bAV507nlWoMAaj
WRX3IEClaY8vpKJcxHPWq4ns9ibNcGJ/9LFndv6/e3KNbOymRbxunlmS2QXBjn/ygR4EQdqSj56t
F5WmoRad327mWSC7CT0WuVjW8HhKuxczlWxlCRhGVWzfiz6MaWclOVqU689Hmzjl/g+zYarmYpuc
7crWwnvsPies+ExEy6hThtx/0c0SnLHEPxGJSWSqt64sIhW7LJk097Ym+0jhTNXqL3J/pANBGPGR
CIRVfwlMRR00ej+nGFS4yv4V+RwNuzmAuqtuRmE45ZRsJkW7gknOMcyurkDWXcAI7Oh91vLQrhZq
463zoDjrsUalTzq6XCikN9occ+zFi+B6KN91o+SuSkL8NDxDB/2q3B/jPjWs2ArG7ryQ9t7GvIXN
Q7eEh73w0qmuiOKc3Y1sxMJ77oI3nr5iG4DwZgELkjj78RYg9tCznBNZOu0+d018eGIiK1MKqfPl
O3vJUtNvJLpAsrC+s1pOj0F2pFcpyIbeahr8nWBa1jQ79SoJQxjY6//vhpwfd93m9IZctWDIRUki
I8+ennkGEj8I9485aaEIdPTOYzAzA8zJcXkgMCOS63SF5lUy0dmbS4WuHf39YD2bLYs6uQSACIrN
fxxyXheuO/JKsuYDrdBzM7VkaMJWDQqARxzmxFaPX4t7vZQKVKlVQjP66q8WMP6+8HRU4mAIb+f8
2OKofBPIg6B3LH1vWAQlFbNHGZ4N6cfeCmyr2OI9vqIam+c0u1xB4nhuZIYsobI71j05CZU6d5eL
rqyTB4eVHTUk1/ljFNF+iAvUnQizUsPbcfK+zByS0Hs6uEg1qiVs0SnP+YJ5g0RrdnaJqPlOsDRl
hDXL6/Pfo5SY7S+hC/NhWlTKZKgMPZIVgnuSP4I4xWbTmR287y1lLKHGFgygNI5rKChypx6WcGMn
8pnVR/Jf1MA/48CTamAGIJICIVSTi1EYOFPxKYRdtIXq2tLfdwXwTBMdAKFHFBZexJ42Pk/6UV79
z33F2Y9plZSKsOa3Yoe29CvPUh3TiNi7U5LT29rQl12a176T7tnoTPERjRk+LaJU0rhtcmYQDsBg
SaKnUXBI52exlEM4XoWsdPbQwrxtqQuRClj/Reum5ZTlFVV/rbL+uhhtVQhE33H2uaRkqwRnr24u
jqAdf8h3eexbIeusmMypuC5JRd6Qujd85qOumMhZAWnohpMyUmYfb+OaGZibUG3Q9QN0JcFbqC+x
NJfkJXAdDnhWp3Bejx2N6Y1vBpwZpdQua684QwBgnwLE/8MoaarUai+cRq593KDTB8WvrA+ef1Yt
GtuGsJXiiLmSTkfz0ShDg71/YTo9QdKqcmjmvLxqfPHKbYbXbJCZY9KYEsWIn1VIJDaFoJv7yvZo
0SSh31MlzAo4vfq4gDO8Sy/vI5ZMDHr3YIO9pxfY1auzQysBBpZrJP1Pys50tjSJFrk+PSJlcv7C
Ur5iitXCdBiQm0n8WmuHa3yGH15/OHMhEYMy1BLvHcbwBZKXeKbQki7dHTWq7RcUebx0lVErRua0
qtX4GwZndd1fE93Hg90ESyp02iECzHOrHWghG6cPphFQTKfo23pAz0tNNzPeXaZjnRJ22ZKgx99j
W/PCLMbtspxP5XAT8elHIY2vRzqN0bTk2gTrDoyyd5hBTto1PNaWUAY9TKbfTfLnQUV0zaX2z4Zn
kzml3z6OrWdofxw20eQViDL0LCsUxUH7BqGvx3oCa8RaQDFOne6jeESpuBqeUVgV87vw6lcrBcvz
MWjDHi9WlABEXE4x/uN9rkc4m0o+aCGe6bbOTJVRdcnVXUKPfPkTqOr/6BYiDn9pi0djXwZ5F8cO
gdiq9LVvKC2EOpmF7/Kmesn/uBJULMSCS4MEKQ8eDssyaM1JyZgANfAQX7v8annMGQkamsv2A2PJ
41xQCsh8qYjUNy3ge3h6zbZss5CSnONpMZIesO6lti/+2Y/++EO652JWLR01LcbXuxiQDTkuWET/
7k5TfoC/upLoia8oRmIHVU6LTtqhnwFOXQlmv9PgB3QXt70q2kyJEs7YnqCtyjl9HzvxjW+nMyyv
LG4W7NaDlrJYGXDfwi7njFDFfbGXMeYDOOw1uLbdDSDzAgmut7qjoIUz5IklF+ni5J81l4n8aTDm
atAqa3jyIYP3rCMhJBWzcKsMO02MhVQSlu2nLboIJ5eI22W63gxZNs6IJ7rjxHwcQSJdsl/TY6x5
vcL2I/ly7I8E+u+8BntNyMj9yvPC2L2P0SMyo/2GhC5mIUo1lhBF7yFR8FjmEez/V8MOuKBxXVnk
tykqmrWx7IAm0AaQgR16pQFOvSe/RkS/o8nba/QXJ28qevJnt+PC+VF0ZlKciCTnYG2rSfo17NKm
peHcDuu9lpB0Rn1btsI8pDSU2WwZjYt9u2VJXReXZ1vH1u/SfcjPCBttzL9axbc0DQCG5Dw4XAAV
LJ4Gj6CHtjFmxwo5Xp5pTMNf9qn2jrIXub9iXRu3g6QVXzf8PcfBCqD5uSzvTvlZjvNMCA0dhipK
KE3ze42Qbn/3H2cmDkqEGlWiCv7lNqHbLoTKhuvhUnaaOmRRfsB7YsIpUG9vNteHHgQGMMPHBv9K
vO4H2MAyNitJmk4eaBGi/9CvNvIDKRT1vFUm2/yGjpeuDIYomXa3qOja1hADAuRItFtPc2g83zmU
2EKd4gqLNf6QzGJHPbOfXywSlqVqcXpyLr9iYPl+TKmxEOibhYDxvnAZpLZKEhNPOMPaOYt8Lj1a
WvODKU2vHF5xG8EnDDYimqM6A5zTckkgRrMfoKE5WJmz9PfYAK+DE5XLdgyVGykaxw5x7gX+MJOY
H2nO4ZLfxGlsLRoB7ctOCmCFxfU7oYy1sddcPEFIHQQAyppDL4o3IPjbswB2yFPbfFL5yGUQ2pzh
4rdUC8xASZ/PuMsbGG1B0Wuy/SYMgtvSaO9aJfSkB/w7GA8xjdXd3GZA6IqL5d082LyAYdhFY6m3
6110mPqPVcLSchARTKFchH6LcE0caHkI2L/NMLWNyASOPhfMjS7zHFHNU/N0BLUNssLytcqkbadH
GEi+SoZMt7HN7tXefBbDIk7lw+16oQhI8o2EBtS+zfD2Jj9oGN7o1smDzSIatPTooEMGRlO079fd
clt/VdvEyNO1jj53lKE4F4zuc5+y7fK5SdQp9EAkNdp4XrwC5pSMf/iCIjSy0AXjJVUnHT13V1F8
2n4WXJT/FOpDxZYExrW51brvk5H4sp4Vv+5h9k54jnRsvMhsftNyhv+GuqXjdjwJFDt0xRetEfy3
tR7UMRmn81Ya5jsgUca1mXHDAwounY2wq90QZEnv/sxDT3nA7AjnG+GH7Xxkz/2hbbnHyBMEKz1u
fQwEQovBgOoyVnhr9g+eKd/tARDUZruy3uQbr7BVlwYT++4L0gsyZFZNP2ijk5ww0YuXQ2WbIAHp
MgnWLsCYClHhfql1DjLKs5ABCtFATN37Un7qe9R8czMAigzAtLzVi/3RILv1PrWBIQkbx+C/uPzy
IUgSMt8HBqjkNsxSgTXwBAhaGz53UrTJj0GaMpNpdhalA1wl7wthuPJRyE2NXU0XB61sxvvT/7Aj
iYKmNMWdr0PyiREu1E3w7oaYgp/Bhxij43MXVIKpHpqvHmBUF5IUONnoWOe2VniUdM78PghSwXtU
1O52WWaFV7cNA9S+aA8UYqefjDGTXuZhLjJRnPMk7Mb3m/+ShH8ICmpkBfzdE0YmxTmt1izO6rkX
K60oJURKcGP8o/e2UEfgKpQCwigOXt7xN0G4l78FhHNtFKaWCaJEwilAxqg8kTfEjB4qLTO2G8Bt
OTrQq3lpIonZfq2RTy0YYrrbVALMNUcfad8zF83G9P31nWgIH6Syz6Gd/d8wTdp9t09wZZoifjAm
gyGBIYLqrVZ+G9wjKGl+gRy5PtDaOnGBfDxT9kow00fTZOMEVzFAN8AwDipV0H5yHg0xfN+iDAjP
oPqDD7q/r5stqQopOYAEtjCOof8Mr4xTJ43cGhojwHBpccQ0ij24JDZZ6+3W8rdx6p/qPzzfMfDt
tWdC08e57tC4j3ep2fYEfj0R2FkEc230pRQAzUmPRrqaIRQQG1lBowec4RPPik9QvOCHY71H7jBa
GLdrvffq1urpWp50N5dBz7nMHB83IS7yCr53wEKSYrK1HyDdrLm5Fs5FLqbgE+OAbyaDtG9TIAac
LuHzA+lRROSQluZDCfJeXUV8znC9Ys4Y/JM49AO0jBR2+ciQMnqhu+84KfxKsTLQ0gIiCZt5QrKX
TiK4DO90KASD8eKInsY/OGowCx7saCSfcoD1Ll/gC7jwee0hN/tXjSfU6T9/Uil7OtTFVlZ2l8ZN
G7jZN0MxHJ+qpIHLvLHO6VzreD9BIs+r7vUKUFwSTFeJ9WAopliWswB1LIVSt3JYa73/tbRco4Ua
o5m1O6kUrVl21z4ETZMKBxPxKnraSs4f+UkaeJE+tEk3Xi0LQhnQbiWFof2pcABcde0Hu7puCosz
AYUbab0LrBma3xS7sKPmTfQLqD76FE/HohLdhn8NOctVEoCacUs6xMkwxvmcnZwNScl0Z+ch6Djc
oR14pfW9z1ElDqLD+T7gsbAwidnBNNK8W8cjLvTKAXmwVFtghlzxmLENevWcy3Y2kTAJ+Mp4eYW7
5/waCT462Guy73ioiLOQOisH3s6Oe3oe6pOI6HjYdQ67/HskUtwxWjCatg3D5StjMrnak/nxxYfw
KYjDens9tWCK1RK+l3BfqqeE7bJguwjqOEmoFsfSC04xZ0idhlZcSw7ybcsNaEA/PGOXOK2Rl3ep
x4kz+hCvXwr0nukML9CGwrD2O2svbB2hWXr6QXZjVwtr6WkAohyFbOJhY42KR6RhcVmsOgiyG81I
joyf2Z7a81fh/cHQw7EryMC0pWs52/kQEPjUxqD1vXxo/La2FY88ReMZ57YyWMV3seTo7KDAMdpt
CDNkKRGoYW8MLbedG/WnBV/KlrOw4m+6vST//8eR6Oq7bDlY3ugwqxob4EckYszAyYPYgO66/oCf
fHNIjUby85rB48uCaDFvwxSI/F1k5+OaM2s4Eu8KhqXqp6rEiszmF6nKn6y8TC5l0VFtwzAqvfMi
ExZ4UFi06xIPRCZmYIc1XWjenPiQMWEoZjgEOhSo9SKEGTm/u8fE7h+Sx1INYHbVu78kqDfMCFg3
Q3qtRIe6NQ+mSjr3ujGTDbcHX18JY1WE4KkncdgEerD1ZuxtjDePN1hlih4EX4LjRRvzA8pTbvEY
Ise4h+tdt4pHDK8r/fwzFH4P1Z5xfzk71h/BDtp8OzzgbCOGc6uqvAStLLGeX9COBBDOWbn4Z/Rs
rIpdiN4f+sh2IUxC4HYdd1oGoenUfQoQlHIArmYEbOHOROhSEhnykHZlG4F86DAQ6bzJBm1DPx16
vGStfwiRs3iVPdXRaIR+abRp8rOK6PBWsJYdPJwhOlbcohaf1lFL0ymvpkW7YfOs1Y4MPf1Wgcel
WBc7tRxDDdz1BorEZHoQW4GFqGxqYvU8Ep1c3PGJbymuKt06JKYFkLtxSQaL6u3Cz0fu4NIFnY7k
flE2bomK96QMuh8vUT68RigvDGS1UyPeDtsL1kc/Re/e2O2vy9jx+sUWj7GVcFzy0UJzAtx3Cg+Y
4+L22I21VKGUTGv5wC4pYGkcqgHW82rBd25fFocqdab1tiwzpFf05cGh62wPbfHxFpfSywz6IeF5
Zx1ALNoe8QcjukMVRM8UU58BJ3B3EOKcZWIt95RNUTjtfHttNOgRVcqHMVaU6ZC5kmMiV5f2gLL3
n6zly5a/Sc0Bvi197Q+T/hrRQGaUpr171VQdlrD6j2j7JSjyhztOWJEFYpdZDUgLKPSoJhw4O3bx
Rix1yG5PqaPngKOqlNuHkfzdYg2hXE2fKpR4moSqWgc8Wa592CDX1085wEfruWrgTj3Pigl4ipeA
kvLQ2DPLrRws/HVLR6uWKVa5fiEB+aq3qOR6YcfyBSd5TzDyW7Kwg7fw5UME3IlRwpoYmIMosOFQ
3qMoCnB3vMfg4N+iCdA+bTfRwZh8qQzQPAnjzXOOFTLCT0HKRSlwkenAFWEl1Ij5lkMzxtmTzgii
lnS57dMveB8Vz9KemQEmy4+b6EM4UBpLAQtBJTDazRyZbvBGvaQSOJiQCQZbCHzNV24a0Hf41sZT
a7uKDgr5Hh1EgKPybS713WH3tUO8Gq/6qidH8K9XqJuPpI3eFgMyGYaKbqhORIpTZec/z1MiLIOs
disvXIY8rjV3QJIIhMLruK47EyYGeLlGUfpGPba2bolIZR6QTNG5A1fvYX1OHnFVUBflAIsIFbT0
TcarWtirvbZrNIJ2JwQyj0cijvgVkjF+6nE48v6V59tgUK5Ol6E7kcCuwHd/MuqOoowfS1/ydlFZ
mJM1N1LRU5B7zS0GOG9eIK0qzMGkqnAiXaAE8tAdhlEiqbGnNxYD5kTa/a7KNqZbBzOlzWOODG9X
5SrJfzNlFSIQ0g2LTg2dwOcIDASsgz0Ph9dlxC3qUAXIBDN16q8eQdl4EMgAhS/nHTljvNR0Xjw+
SeylfkOxA83X4YUaAVcqu3blNGUVWygin0+wASxpusJF7C2lT5PAuzxFLSkj8tMzz69H6nWs9/WC
WzardQgmts8M2tvEzqHXRFK5i8Z+MAUKUUB01S6P8zvwoBUV1HC0UtoW5rE3e9iqM1OOXYBiQQ91
jiMpiS+lI7gjDafgF2NTE++UPEz//9C6wr+anGFW4ETBJek6QggfjG52pUhAVHxZvldhaaRMVWFu
+iNdxr9gPNkJ8wf51tW7eTDl/x0QtAbyf1EO/CegQo5eoTGxuq6uZ9NNWDSCyGxEPngpnd0Qwszr
itFL8VuaRYA0/E2cR9kla8Hemd4wyjcOaWeI/O1emngNo3/3FwQQWtkrJ5eFGlsioDQG+qyUEkWV
gqanXZ/iyc9gnid/aKvolvh/GXmAXkxejU81MwG+nmuyR2+zm5hs9GqE7ZUVGHHwTOnVTqd1xbKC
LJ6kqRT1d2t55wrVQjDgX9bxlIfbthrHRLcGiwKF7IsM5AG4DN+chjXKHDRSYg00sRaXPOFvqBlZ
+lR6dA7r1WpHDK3dw7Zxplk/dPDXPQMk4ybhopNPqzqvVZG/K3DyyTF6OmMrR9Qb1ekCOjhpL08m
CM7Oat81AXjpV2DypMkP81/Rt+eCrnZDYSL4H8TevLK3GpHnmkr7as0BU4EaiM296zIGwtmS0XTP
5V3mrijnTL3m7b88brGOKXh8DgzGJvsJrzf0gxCnhzpWPbrEBvmrt/IcAoB6K94+lP8tKHWLmEnx
CG4aTWroxSjZ5pg97oTLjgPATS2HKR37HE+4tkvSItQMgxT9BKwmbOTwQ6V7Ou/0bfPfV4Adr3GI
9F+i89kzkqLTDBAzri0YWwRnOTmDMW4F4v+oV7RI0cgd1K8Q1AsBzg2CU1xnY7R5266V2RIIX6qc
Qk+wjp1SMaq4e7whanu18XlZW6HhLlXefgWY3+R5xqmUXaeVdI9stMetVVe8to2SkiJLzWd2VcaY
uWOx3Tf19elm0fGmGqbr1xark/uU/a4f1JUrpxPV4SarVsUcy85jIouK3Tah5XCWylUmWyTfvjkB
VZ7rSKFrWdJYIESe7tKDIfvmsdLPfCsQKg/fg/IwCWqO5AE+Ey6YHAvKUyArBUhqV2kM60VyBCLw
rkPrwaHQyR41aCBGb8/cFhGe28dsqwwlOSqIYwu2NO0umpp6wBr6Hug+XTCYHfo6FzNw1Xt1lxRD
d0jSpc66Du6aIscNpjUUSWtxvxKVsYmdTfsn7DvIRooNzYUtXRGGdObj6jS8DU4EEGvYTxwjmaMV
9g1Scq8CqE3za9S+l4ZeJNkN1qZaZWRenO51hBIvjnDa5mQA3vjXlSL/L1vcZsRMS9s9ty+8VVrj
zP1EGNahDK/3zL/UUNr5w+O+g+5RiJ67x7LMhKwc2s6GyE3PJryuPZvM6Be2DSeDJLtQLguZGsF9
PuepjfZPqHx6/Nejz5Z7Vd2GcwOiGmhIqTMlHqu7nUAJ0UHlOr/n0lhp7BMf/8qMzAVqu39p2ozA
OisSRdlklXfSB3e8uzrrE0dPnkkBhuEE+wmoLw5VfDU2XVLI2ZPcpJzs76kJ+VIGMvAsIAJI+bNv
e2iJ0cpiTGSzZBXiv6piK6HUeZsJm7jpyQ7xmBbqgv2pwYiOFXtu5YnTjwT/5d7D80eO5cUNE9+a
y4Mlg3voc2b1cihXMrgexj5K/VFlxm2CvnMEfG490sFVcklp1mXkQkcVPJx7tIJXnOx9d4PZbZMC
XA9/H84RaIr4CJWEe3uCAQ8oBVQKmiQaX4KdO0vVUW5h54uBZ1+iysIsyl2u0SLUBBmBdLHFHKEt
pENyKsdqqPBdpetn99QjjaU4XYbvI4f+/3WOhJ8+W9DdnJ70Y4s9qAyMwG0R53HSvg+d9ycxTJL2
mR7wEnakppxE9KKg++urntR8duY6l8we16B55xDoIHsQh5ZTQ4i+XOg+SX5p2QN6OGT65OS7snfy
RIFvAgVZU1jxyYnoRtsTfuiRO2k6wCZ5aHZhwvBZELTxgTdV2U34J+Q3Cj1MT2VHtPDxu4WdjQ94
WrQ0C54xUhgNXflvRnOFkaLOVF+vw5iD8zsBDo8TEWrgedsPl7njYe3MxA79ARMfMwgtbKoEI4hF
pzvYjDTX5k0I0rJwU7gRvvXr1NBXhunb/T9QDdsniWn0ssIRaZJbUkoXlwC5yHr1rfLRFzqs6SSE
7l9DP+BCXAUHe0YETGzPRVeNx43n/JUzEdRn/aMvQppQ6va9E8SOyNJ/tRCvAupyV57CpucbzfBD
0onYaeXF22Up7gDKtWGsxhjJGbYj7XdVpBMhGPkPgyXSSKj7mXqdcIpiakjdWnNAhGu/gCvNJHh6
dZtnln1h/BczP2pf/Ng2wG8QRmANfGUBgAmGwiuG/kZ21lG679a1Zqd/Y1igtmp4xPFX0yxcA1+1
KUiaDrOTwxUFaoylTfieaa1fYsT5+bHk2IwaLlOMM67akJB2jh4VH27+jdj4jlR5SLRRR9As9j8s
zI1TkbXZ0aijCwTpc3QfzoklRab8Xg0G555gqiu5vsYfSi/yp6ugwXJONfRaq1ebwCR3Li73845l
ZS1gFAkSehpokxmqP6tlHmDXvkkSsAxgNbNt7mOILBdhO7nMl8WxPAZzJZRcQdXEqxWA8mz3d1tc
J1LwclTMufnFdYnOC5tRsAH9BjXfSrWqramGoVQVJq48Gd6k4CYpN5ONavhr6+JLOVC2S9mOMQBb
6RYulqh60HtQ9q30LHK9DqlKP15TZNJoZFAqxkPymQESidwZKWb0feN6kuJmzQAuyqiWPRWBj+gn
RSBq3SKBi4iJt4SxypszXsaMcOyR6c/2e40BnZx3oWOZyqn0Q12xgZ7SuS4bnGRlr/+l33DJpUsI
r6VQbJ3yOiIBGm9a7pb587ym510Xd/lEIQRmpWjDKyYT77nM9PvPXtXMOEOTeI/L74jgMtz+PkWD
OGpwokr2/ig8MEfE3vRP1v03z0m/tbzElGfpNb46HtsPf6xDNIT5kSgSCG+IHO1Kq4h2cd7ZwGWe
I6g5pWgdIRuxJsoAQs//SGYi9bRLDbzHBqtihtsuBIkaL/a9y0WxK3iPK6NROBUSVupSHMAUi8RJ
NhS3vXwxfFr7AwJCGDKp4GzL7LX7PNI/ybTBJdHMpS2SKihaVMtHqN1jLcnXf+bSehIACIqoiMtB
1krSi3K2g6djj0q+SXjBu3dq3TWw9tX9g6R5Mbzx+uGNHVYmH3159JQRKYUmxR5KMVqQh1RvfURi
fPxh4ofXZz5buuNYluKNItWflzNoyjK3nLyVnPEGeFK7fhDoSOVh20pqBbJ/MetakzLVbC4FbSEV
mN3A12j/ZqFzELfmdNLLVs+UTpPSc3Vp7XKD4MOiGiRLBBhx36EaBH/QWm3wIbfGIGCN8MKeTiT3
9ljP5DJkbpBRGP/vE8Ii2Q6DmqaRye9o3AkZOzjhyD6EYxkXU+St7wefQDCbyDcPzp640rj6E8ag
y7TwA5KXezcVWH4HYYpAuVcb7WXhtiozlyUvBafJ8k1weHkdOE0ZgS6QuGcm/PHVJEhn9NQl6Xz5
jQ+VEbPqD5WcHmtg5wmZD70r9gFuUg8P619Hz64ZOD75Hi9YahUXJVap2LMizHaMzlAt8ttrXige
nWSGCsBDIaAv7ARLj72uJH5OrLIHk19h2FWDDB/QSQb2Ue7+4+gID84RgrvPgVkMB4Kozt86oBAw
Zym5zlH/HYge2IhGiOn0JD3RjelteNTW2ricXlvq+cSs8BQGbUEk96PFCvgYlxPaI2m269PIuO6v
FoU3lyjaDdL6J+mOUzILaCB/XhpuuIsB89lMNdj3Ecy+3TALajmq23KnbEb7CJMJfj7W/rzldAvV
kgs4A/n5eLvvpM5giuUvYCEMSUT0C97Ub8AMNGoU9soaM1I17GEZ2Et3sAbFfFNv7vBI05MNxfXn
IZQ+MUiuK9B5WvrXgDS+HLYFl62G50B4UP2J7j/cNlRIPXtGPswO/8hifsbEvk4Fa3MDR2z8x2u/
uLiAU05sf3daSCGovW9isznHCVbF1PACETihEeLPiPYP/c9KEHIYo+8ahlZFJ7UMaBaz9rI1u+Nl
6ZHJaT0gc7j4xzC2HU8uCQBas/mxXTRK+kTwNcOILcx1X7wuNHeQFOiA3z6oOtgqB9NwAb9oClKu
nJHMIQTsaLn1OyvUYoLQY5vb/SqBpIOb1OzJCJ3gHYhMk6tdojGFHFszgCh3QR/HxjFGmLVHroz3
41IgnkhUNFI7ZPg2VJSCQLGmynccickWxJQGtL/T162Bq5uXigKMdO1k5dBe68YuRyIR4KdZZ+Ac
LO4Md3wWSYkVAOaSveLnLkYrLn3LBn9AEIWSIw+hekt9NpQPDWxwbwzTVoors7NUgBPOQEFvIQLI
T+UrxadMG/E6w2zN3l0t5a3hWHUQniheyRZIGZw687UqD1ZruoJvHWi14wiux1xY3CkJRmKY0bqT
VMfAaV+7WaiR07dOT+KoEpu49VTSJ09lw6Wmym35nqXw0IGCfD+sKjTMPOr8B51Jcg+jqG+AzlzD
fmWcgvYP8MFNorEL3nylStQ3oHQUxB2VRme63UX2Rp90ehKa5FzC1LgQLRDooqFGvVgEQel2xEmc
YmDXLGZbtzqJmSmR83e8ZJIHJPPKn2R6X8d8otmtlWdUWIZXTzSxK11cvzWTwImaxGQYCchbJPBP
AnthhhWNtGSIRj3bOdDxwDDGvMiuVjkiqT/JSy5ZOxDbwHJAwGEifzn8X65oH21qMv2Enh5wtJPr
5krUamnGnG/0aU/Qjbk9e64wd7iCrpJ2rPbsBSHcofwB1soi5ghd6xuQEG/G6GZ7f17QiXeBzHES
6TMeHq/WlM+AsFPqNBQrTVV2Jk+wfr31AUhdXADp9OcYzHE49HZnyMVzK0orpeqMCvpS5AdmbtKj
5rifh8FlQyFBzYzfPrl0tVUjcWVXO6dP+9zd0TWN7Pwz+LB8/CVI825Pzeg8V9nqoNn8rAeTqt9r
fSiue4MmE2YaeIsVvkYjExnKkK1p76Vx4UsINo0Vl+j6hhTQ9jCi6STn+1wDRl5rO/wmCPwpHn5H
UR3guYrXprw6cg5lZ7Ton0pT1jv8U0YCAvDXBXK1GyxZJUjpPMuGWC9trrW6CXaxRzq9jz1SZScV
WQRwTVtahCnAFhJI/b9SpPfXOHgGjxm1wKCXd0hnIxfNiUUngBuqyptVClwXHcjlaC7sM49eKMEi
rVhxeIgEprlYDDcBlKQfazVpVv85CHPLTJUH6pczzzVg2mqJ6YLXItLGS/ETVxFikxIN5oculyYb
pE3pEQwUZ+vEybZfkw3fMv5VQZkYv+syKVxTv3ou1YiTsRAMU08Ly37bC/XD4/ObswyYjmayqw9T
a8MWNinOtWsY6urpFr3FD4RR1WcEbGDZjxKgugkq27uvC9eQPi1gHcvir/AqrFWkAuIYIk//YduY
1BkIamImU42Em4odv5+3b1lf/4pdDy8fxSZn+jlgksOal/nfTMqrG8UvAUJSHGV1/AbXODfl3nVA
gvrrQuv75pXDeTGpgEjRH8AMQIqY90exHK9FG4bVW2T2jeK/HR/T5pcuTw6dADUrKEMLhcUtU0TS
wPJOoWmau8ffTIl3UsZjCwPviKVQZEmy5GSipF0xrWvsSCfVTkrrclBkhC1GvPkY/EotZG4nv0EX
O38PRAlPmRB70Dfv9EuXEfljM2lu+kBNUZ1qxKqe46Y4YDO1IlK1zDzApS4XUMz8zfPq+8Os4Uvi
FweJ3oUBsvZW/pBEaUlfh6ywo8fJ4KOPujwudy6gpkMWBp1y7CY2cCtPVeWBlVYQcEtfHnTcugsd
NcIKgOsmlTM9V8ilM+kus0Btzw30tV1N62OSdRthD9sVVdZADxtVzGpOU6hIXzmI94GIWwoQ3vrL
6cx+Rh65nbM+Rh6D7xwr4vTIopR7IOIw3F4yauDOK+a0MBtEt8fxGGbCEQw8cPk8VlMORROOa0Eo
hZdm3MMX9tEn1Qy/XMS6BsWNq7U2+bRLLHuwDnkbVVlcQiGY3fJHVs/7YtTgjQ9ZrWeMzWjXgvXm
fhV+r9y1TscheQQ8bBHBQv/NDThURD/uZrksrKs+eJsRr4dwcUFgQXXre2nH5oTypV9qWgmpYI/8
g51NdEceKbezpR5EtFeK5OAERmEEv3NBVyjTJlNCQcoBThsEC5cfZArNS8IkYacFEDa8tK0rnIux
5dpK0EE3mTlUUchIJWnLHr/630LfMaWnB6HVeuXoBX5kJnBHK3OeeXP6QXkxo59gbuLZxUPhJvcw
tUn7ZPUcODo+pzMmkX69YgE/xdU4cTZ0I1C4eY30iQMJq/AjCl1IQbvkSGbFYcYXKogzcWeJJ7gU
mmQUGhwsWEToD/9WzBbDXjUMIMUSh91O8XyrZoMv//5NZ0E4+bSqu8MK4mVNMXvStFtC+l18HYoc
d3mdCtJAtvE7+r6OxZ6K+WUT8V9AO94VG5UPt36WXqHcJ+74VhkEti7cGMWrfe2yYiYfwVsrXZAf
W20iTxCjMg41tG3pCWr2hbICIhZTQzByZmr8nOcacZYXE4nkcbE7bZHBaSmrCif1ufDhicAu80hz
w97KL0giu/EL6scKcm3Q0oOY5zLiL1YbX28YYNrgmkkjWm/VcJ3VgwppnAVqwfy3aGTSlX0i2JIG
bb0CLl6V+8pzZLV7zJ66VPvqIjooLI3U04P17fLIkFaKQO4LLkAsfehAQHeee/TVm2Ch5O/ekbNP
kordQnLdwXFz69iMVgTrVZ/Vs7GxUbbyxB9OxlVJ/D34ba+z0HW1hoIvkLUKRF7R3ZJBwkHHeHEz
q55zaJpUaaxiebHiIBbAaoHmmHKf2vblL4IxFxLJXZ1gvNO2QyOs/KahHg7MYlsEIosSyDrjzomq
bhbfCjBNHsrXGA3Kz20ofF/1vR5cjL6lOQjYKh/6KwzIt+2iWVvoO5terMezuYzLOonJ28iJ4lft
Cnsu8WXix3Uixot35psUO7JWJPCmM1Jt2L6nGhbi3MezF8l6Zt8iScDYKPrr+9iVXVn2vS/S3GVk
JljD0g6jJOt5/JGZr1bfvuJoM8sCOmbwRjOeb8ol6wt6z2yVpJSnTGB/EZFv3YYnWThyu7VDLV8/
fWeOPaCVHS5NuUlk5ghkVmWVlWRxS1f4MZTbV5YxBsPjlo7T2/Rkewp5T5GB0JEwKn21L2UKAKf0
CYp/Y8Er8ITKQEsJovXGmoYwVg2o4/qySNer3jia8lsQC9VLRHbAqC2IidxMspDs5vx4otcHdS8V
tZLIYNE5jYomSuA4yRb34/8kLtT07CHj+6ueOCaXz6aNhKsX+JUsBTfqEee45h/jBvgra1Z2k2E5
auYNzxcLJg9JgfgyVYghMbLodFofUlW8fCMQa156BjtSjmMjF0mWvJKqQ4cEzyyCpYG318aAO4np
kaeN+We4UOFo72gmesUiUpn3Md76GtS3Jgw77pY/vkZvZBCP35qJoPGY1WcZYVq5xcMps3QKMYne
L0bF+Fa9jdPnsbHKXeNQsDQaWPtlpNI289WLpZcDDQTvBrdqfREl3bObWi95Pog4xjK3Hdf5Fqxt
qBrvyFzymp9K9plfpTESeNwLZid1DpMxQsXW+od+5vK8WqwLL0eqSSHB48eDAlwXqkh9EuNQag/3
aJmPOMGjTHQvqk6Njv6fNwrmgZQGRmmVjXpBY0T7F5W+KnW7XmDKErX4aboY1NK2vwPeuZxhysIP
8CcrYoJ/eGagGwyjmu4fKA9wL2upt7oc9A15ZpAL8lBhq3xtvBzo4mh+WBlFzoFZgE3YolmCT5QH
XREU/UzNdv8ffxLc/KbcquGgcCZcj/VMIbSgGLjAxfYejB+OSlMlXEyaZECYam8zZOf0u7Z9Yfsa
kQag2LngOispxJQRPr8hwcw3LrMm+NrtAHYepkhUpxXoGCUJD1g1R6gRLAAWlltq2cPOIupwkZ2w
yDbMbryemiiyy8bsE15t5KLzRBds+IKh7CbHJOY6r4cxViyjVjPXz78tWK65IcqAlUFDx+ZG2vn0
tBpjusLYwlv547VgnU8uR0ovP0sNqoogxMqaBRkp+34MEmKw+CvBUt0W7wcTuLW9kltQp0D7J/KC
33J+/q7O8+Xw156PpJAuq+svn7c8/lpCtO/NpwvuMHl4uc4cdR5Fpv7zq//LoM96MdH0uIXFzQcL
ycPndun1u7lKJvsQ9gYIMT3bRj/PQd6h9GFpHJHkFstVeqob0wgAzukkWdPxXeeg1MX9lLXxpM1G
8lqVe66YPvevuURjolV4KilJz7n8bKQ7xODeaYDSZyT3Y2Q9SzsgOuEVdZRNl3G4x750e/oCyZs6
rBKVl46qMJ+6bdHnlpt0DALNVsE/A243FDYbNSjusFWVmeFmY0JduMUiYjVL+nT9v20IvW94cIoU
GqIU65v6wUPZY2jUzX9jmiuKfWhEkDS28aMJ72b6eVoFFLWxUd8X0tys711UR619bwg0SYhEdb69
Cb+06lXbdapfB8tVuMatNJeoUz8XMKeeQLan4As4WZtp4f975LoD6BHqbuyiAsSQMPQb4P5DXf9I
6l1nacjXualc7sl1TQ4KGcjizrqTum/SmiEtqUM7+HiS5iN6t3txdGS+XXWHWgABeyVq5fpVrFam
IJTWRLIbyl8jpjBINUep5W7hH/Y8XGJdERz9uXw87/r+TdZKjTLw1Ux0iiLlwWQl8AgIGQr0axiz
GY0dbyWhz46hPJ3TxOkQ7fVc2s7n0yFSb3NV+y9EHIuTNrW63iMe2mhz3p6RrnoUCT0pbhFkQWsd
kEObo/wsg+S3/FBl7PJDoB79Cz8lzBxufm2lC5TAOh5XRNBtoE/SQ92u/hVAgG1u2g6tGw8ma87D
RNGUxkoZffr+C1HevUJey3r/nxSSl9EvPuHcz+x3hS3aGKuca/6YZ3SkypktfdiewK7ezjNzc6pA
o02xBK8X789AsIzMn9Momy6237sWssqt3cJbznNI9mV5biO6Yp9cuzgiaSq45+qMMJpYOXrf0ZmJ
oSM+I3cia3lQ4KpYgQw7q/8yjrJt4YmkP4wi9ge+dMvym05gqHlImi2LsYmXyCJXz0aIrICnj9kl
8z3YEE6P+ht4OJLJI/o6/WVOt5s+tTPxRys+LhH07y/dEoDOwcvK096roxmFyOTnU2eSToypwF1l
StEr3A1H9vjiILRjXOCCg8F5m0Z0vmOXgLduudVCValdXK4i2WZyCDzN0xJjyP+G40ARB9ou9a2a
98Mdhg40wuOt3EhtrOPAE9djOBEZ2GUaszvrxHWCTC/FCtjX1Yp6mIrsbEqxLHehUtY3AQICLjd9
raOP6b8gIz0tWOQkG+MdkUunrIVmOhTY+51Hm2MxYs57sARlQ78ULp2M/dBL7S0jHLawI8WOw4Ge
/QR6Rz0qAtpXgisrZa3r8NiESSBFeOHZy5UYfPN1vEr5sDXVqoGqpcRKgjWFRjZZaYUFA+TptBE3
hkVysKoez/MZxpScGd9PCI+/ULxLU+fuZMET2R48CHOeHyHrFnDk3h2xPJG2X+Uivyg/k+ebP4GY
j7KK5syQpYmx8eGQ8IYqB6C14lJuyFxa2ATtCIhLM4vZDWbiU87X7sQDxMgR268ErOt2zdcFiWYl
PEPbsE0O2fUK12SIK7GDB8OjMuN0JW/LNMT21HmrjOgzncvHppSoaF0P0TJz8LBg8GWXI/QE0Z2f
73zL5vbgV9f3Jy3r6dKtrucsmpJzYLZqm6DwvtukB7oivXmYe7jEEX12M6Q7qOlDex8/AISE0fgW
33/0il7hQFz82W+i4BB/PxSmyK+wLVIbjDnHX7TNQULLrWxfG0nXM/V9D3wEJ900+QPq7REJauuX
+PsxQsBGelRHXhbpT+Apb7V3DbpFDMZDtfACpzepoDFM6L0yZXIjrjiD7ZKrZNC8rVERrub/ftMD
kY6PAD/0wOWx9fWR2Og2ctOaKO0O5TEnO4SIO7TsEsEX1qR5k+knY5RtKHmmqPdsyARkK7Gv7lcT
LU06L860e6ZHgk7TAARmXwcqtKEex+IIwwDwSta1kad66fMgD2YEERJSDiiLuWkTYQU5wwgaX8XV
1KCvRmaWyAy9MbR4t2YlOSH9e4lAwhXfmzehrzkQZ0nU6mcyUTc11JP/DrJIjflhWKDgMlISUYPl
ATgCN/BOxwMNKT+VygkOFQQI4T1pJ3IQKyuGSaAuh50j9qLb5TMdMS73MwigCZqnXicKacB28WpH
h8iaheJsJy8TH6VbXcc1V3oUd1ohNf8t2q5W0bhwxW70Y6mpqomoSoKQy2MLEUNn9ZcIv2mKKpwP
fzThFssHt9iPndc6kLrY21d4ujzsVTpJdQtt7p5q3Bkfu8zloOfzozra9cfdIcgbr7CtTsV90/pD
2rLVukTe7xyKCq5ZzZaX8gV4QF6d+0Zh2pfMlK6rXJmDTEfTJ9C3UFRi3QNC4Har/OViJTNHdSNN
50moaSGnbnpEssXCSnk0iR9ECMQOW0Mx1+ytyel+pL0XxZpQuVSgIM2FyOnvqOBEIe7o4bIW1E4U
HtHuo179uFtqkf9KgwiSuCisfubSawDixhYzExP0Qnn5htwex03AxWv8FX3ii2AmP3fujoXbqrPh
6V4APjOXQF3XSfs7FUBRENVs/NlI1Y/xOQE1yUg34eflQCNpL8HUKMZjOonB/xVIMJDtWm11ojdA
Vmmk9oVwxb2D2p98gOTdZnGxLS0KSwQlMpO8AbFjzCRYDZDqLmCPvYkIz20FQWdAaqShu0nlnIsI
Q9NxCzmauAqTkXA8wozutwjckR57VuZsxx5fFUbob3De50gCoPRkl8USyaDXGcf1LYd3BPINIASA
Q+k6Ks/jddbP6ukkrAmAyUCzTmE0GQLK5cfDlouxLMt62VjvBvC5l1rCZR9WJhzEmbRvGT9fgZz2
mngDElo2mOkNJPJo4bPk0HmfgKFqMHlvCS/0L9JNMrDTVur8i50oAm50K62kfDZHtT79EFIWz7OQ
Ut7K3wyDIiQpW3EYhmMAbYTOMOZAV1lHPnDt1/M4d9Bh115wj533wMRzvmFaiwItwQIAMIeLB9+4
ciRs0L1uPIxOI2iide3DmglQ3Deyyv0rLmyjKjf83CpI4Rx1PNIfTRusJin3T64v6PHHojOBoGse
FB92jGhXG08UW2WAnxsR7QRz/+W419u64y88bAsKrDXaBRN8RPZuczqH4hJjjW+c37a2Ew/wer4B
qZTxD0J7pqycUAPZCu6vY2LfViAJkSnd7+gYTwUFZpOxKPm5lG8XuBkYm4yE/M0gyDdb1Rmzj8ww
Z7FCYtbCU6agqghJjRb6PBVgCt568u92l8CrzNAD/n56zbnygO6xf8H58BWnvh1bBqIkZf4CPq/Q
Pp5OHZFUNRxiSl4VQds4PQdp5UK87vFnlvjuvmFiKDYsmzAUJkbksRDEbMgIbMFpaIZTj/opO3N0
My6o4RUm5nfXk5Qx9TcYnkKLNzGRZuLaaj04ESR0hTgBUAOLGfViW3VK16qYeQsgaghohj5d2lHM
a/8fztJFRn6txbV2RpMfB9SD5Yxm6rHf2JM45X8Hux0Cw1mzsu1FwbSJtUqGFrMaC9ER1TnpWkdO
AzkzqOvISGWPJQswee3DqYuj6yhw20awT4APjhiZTQiirSKQkN1ry1fuJImxVpbStKRwFByB3CaV
XK8ZSbyIn7Qm5TOhom7ucI4o+g803kNflBrkIDFRWdu/u77Oe17Vc7vTLuEJK03ho3kmgzIN689g
GwinyOZwtbR8zI6TQHdBju7CfDx27H8rN4okgOb2Lc2QaOQeBaszGbZIWvvnR4LrjaZKQZ9l3Jj0
mZbFknPsnIDdgYnUYtwbNWfjXx1InZK5Z8Tli+p7Rj5yOBulVyX5MiOxPeDKMwZbZ0izM4DWQ5Td
iLOe1DKzpigJuvgdeDIXf+QI/w3uhBz436JwSEjpwb7MaUdvB0ABwiRy4fmoNogPTFFcOkja/r+K
XEG/6PuY0LQKqfv1RfO10bPbojYrBlySdZXu0HeCGbX5nITyjH8patr6ytsBhVLf6p0yHVuuYFAi
XgDSqK/xdFE8IkSsvfiZPCVXGCGyWlM3HQ2BgPiEMgB56t6sOVdSLBHmReK0oWbFmwemCIPC1dMQ
6epz87VVKc+z9FSZQecPIbXBb7abn9Vm0C0gwfM8cHPyRT43gvYD0W/l/ytGBDGhipN2RJUx0ERg
99vMrM8CZwho687msWR5aRtfIo7MumTi4CfVoKovwEJyfIEeBTRocDsW56zFmrNKEJ3fRy1nyXrG
zsDFz6Ga49TnytL80/U/GSs2Q0wqV/Ln2NOzUOF5u34DaLdEQbxAV2SVQhoE4xY2KB2sNsrdxqe9
rFYW8BeyQlvxHIytO8dBY8xenYuAIkvCFIsdmAM+/7bo6vEZxpUg7w6sCZaSaX6ZLI4Wai3dJPgF
j99wUeQTJuLR37GJ3z6Qd0USxEjGwr/j8LhmaSywL1KtHuAGPiyAS6+SmT6zEX7AJhPYTtkl5djF
ZgyLsL6IxHpDui6p+pakJfEF99a56+9D6CoCnSP9dk8aQ+TGfp0+NNmKkFpQm/s2KQntcL0fie1z
YpGUGOlCLssD+AkMmPArV+TmYqnML2BfqopcCZaYzLcG6UIh8nOmn1kkpvDgFKNg+b/jIqwaalui
+2b1GkUALTMubWfXtH4y86Y0gwdF+4DkwC8F959ytHtZUaHq3FdIpE/rOGyWR0R5+bGDWW4EiQyf
DcQYI8uNsVkJD5FQCf7eYbdgcXNluR7fOwwFHekRyg4bmKJM7lSKAdMEqP8+7Bz7/z9T85da++la
JVz2ROOS7J9peFmfEMO68T6OzHjhH03qT+bUDdXyqNeyRXFKWeSCcJnl58lrnzEOzLCZSJqLSUNm
zKsnY8TUeD/Mh0/8SZLKTTCAWSuZCN6ZWJ3jb6/O5h+mcY6NWCj3ITLjQkhNlm4/Lj1uvId5j7/1
BwuhFWcA15wiyaiXNw1kea4YKYwgRJOWW13KeqQ165HJwRYfUmBjYsWQQ2iL6gFQvBbDFfhfHID8
esxbCf44Ucbd9+b37yuh9YgslDFuZNrX/LEWIetQDgLW0C7ZRSrsncmyZLg9nw2HOTu9NNCsKdIS
6BowgcPV66O6+9WlofpjYjMW/aGxgH94YUBVLZVgEuJV+xd/ZKdt11nzr7dY3Y3Cv41GZMwOS5rp
KNfc4we6z87gavwFP5UWGrQizlgQ4VVof0HNnoNLINfpg7yErOC3foTqAdRGkfgMeNIDa20JWQ8j
OvhSzEGIXzQtZAgNZ/BtnYG7kpzoojCGGOrSw0D31KrnUGMFT8AwLcXQdPXHaKXuHfGaX3F6WlHP
cARRI/pUJb7fGMHKAkQVpSu5vKVAvergi0GL+G5DdQ8yxGA0xbkHzR0GRqujQtQ4o6mA0o3/UoNW
RvhfynJk0fJVGspqMGTEN2met0uP/8jIOqLfcs8aPPrMGBdjb8aBeKAQQ8HUomR4eZ4XubvV0xI/
c3gA0vwtSl0lqHNJH3XFkgrXZq2Cx/UDJi7FijXUf6DbiMCYk/UBgORilLlHtpX1j3XfAiOcZ9mR
HracI1M44seFPfSdkvMmu4jI9qGAI/gzFE+lVq3zi1yNDH2xBmCeZQxMcCdnKDLpU3jhBlMClrXw
XUNwJNJm3FdXZ/bDxketCh2ZKQsTpK3I+mA5l2vm0he8KfmNX6iAoF/iHcWiiDNkVR4GitCWXLhv
A9yzzQkUB/83rWCOGcL9a5xpWQvfGBvbXcIpI6y04oS72vSIIMM8mqebJCUPEBCxKIeMBwVbXeSO
bVjY/fhp0jZe+Cvi87xZUIfw3NR/6obwDMZY3Ptapu/89dnsuJrAmtZBfE1uMDCulPc5N9vCIpmg
DtjuraxWX3g3ie25K2o7/sTn/p+gQ0B4+K0fWRywxLTKGmX8XYaqhr+CUlUNwfsQLXflsgr9dvvW
SNhrO5H9MParKuZRJQvzJ15r6T92+SnHFHalQveMuh6zIrJf20zP6MOQmF8RYT91kd4+zNnDOcEV
DrQP7NOqSIHriEQpmNF7T3+fFTm08QfvmTh82J1j4DnEaSsLh6al1WJYQ4AotBEEua2zFyGDQTEe
BWhgWT6JptDcUdSoXmBqFI5zMvKXn64RTE3jbiTBO+5oAmEytFLKRK4qYrey0V/mFfB82Q8Ml4bK
QaZ9lIi3YwmE+JwRNkyHcLNKhEeZ7fSYQudWogJRV5OTu2vdaiB3wTt8EzMS5sPYt08yc5HgeZj9
GLdqw00IJxL5YARdIJKpqhBVRDVYd/rwvQOgUO4VHc0R+pKuzvCepi6V/qrN7hRQh7fLzsv8G+cd
ZvVt9Xg1HntL8Bt6rBd9qbhAmn+3bdjdNifvudfF1uwIDxHg0oIPD+w/I66uDB5ShsRX3Bi1ETAx
7WEuCk9gVDNkAGWTcZsDdhEPQlnEW08ljFrNAwOAp2Xw6pNnDpe2K1mnIMVm9/FFeK9dz9mghwCY
FkmKtID+HwYyuuNPXhYBdU5K2iIQ77hrFwqQ+UPddQvw7FzA1Qk1QjdoKPMu6xVyKhHJacbzWEY6
9QGl6UTR4eDYvjNTPos0D01NUfQpDjhueVfnFhAiJYIPWxL4FzENolcLUi/H6GfXwY0Kk9KmOHeF
R2Zz7pYpbOEW46HyqwSqE5fOWB3UKfOewRnzaIv0Kq12q83gsWtIgUUQGh+Oi1Pt3jnmzgR6MDUX
rW1qkF/eynrfY/xZZ+pf04QuDXQFQshezoSS0pFYbxGhec44djPFkZcY6bN9AF61tZ22ZUuRzJ/b
P1/DoPRsnBi/2Mjm/3OuGAffftYLTkfkVTOjYT0P/mt5ICRCNba3Bxb+8TXVS+0nGoan6/xV2G7Y
FjaTPncMUfMN5XtcAjlK+uCLzWiozlKskLCdfNhaZyYKc2tez1zYtyCB5W3F91VN7sEzBcDOfDCV
MnKVVJWPszOjf93eBuQK3e2itZlTdrXEBmAKlOxqwxgduHFbplHWdqINCUftheR21i1xV3JCjHnD
6Gm+QDxGumos/FTPf0Hb1EJM0UD+5Uyq3STO5CY5uvNAQPUFe9Veur+x925ck9eq5VFKIu4DaSWw
KgPlUVJ1erNgLmezEwJ5cONXn5lxpRRzAm2GVUmWwNuQGc/kiXEKrD2sd4XXUicKu8iPeDQJCH8E
McKOvYQ2FjL1VT652qHpKHG8JhNtQpJ0nT+v4dz1P7CSvePnThEtaGv0iDzMEWUIcWa3mP6JIhyE
O9h4EutE/Arkz9ROWNEb12M4Ww+03kn0BD+bHC5GAtIsOq8knUZvmi6W66b77wKcWvQkWR1HQm/S
QrOPiFvVXqugI3SXBwewNeNdQgB0NOb1HZL7BRFPGgA4FmN0hvaUHiw62MoMl3wT8Ui6SPdmK4t8
gQG5o8Mp0wPyyV6rM0FsylmE4d3wqNovUPlOxdBVmrZhtbR2ZDKqA+H5uqXigui7ifUAVA9BrGHP
krOjuY8GmX4rN3s5hP+PFWr4/LtP4/mH4qeVLdHU4w2mIFNZNMh57/QFapE0C+QmxviQBQb5HJIi
UCjSbzj+wGFi2tCDrFhP/V5ioTCTMCdvY0D3Wbtf0qsQeSbNtic4h+laZ5FAzpCoX4mCRI5/r46V
TXxsC7MxN+4rCa1UOspgVeRklKn7LgRDgY+QVdSPLdrwE+NdsdkprMdXCRqPA96TrxRKVcxamxb3
/EhMAoEM0/jEF11qNtc/Ies7c5SS66DHkOTyDb/tuBKekOrrlfidA2/e7Q6xAKEsGE4suLadFLRE
SelTyrPox0bRA7KG1FkheTFGUQQEGD30yoRHmEpbJ+kdpyp6WgzqHAwOetAJ90EHJdfbtNDzTKYR
Cm5tZkD+cdYG84Mgu+Myqud+oIK9/sbbs+9g8wSa8iJxc4IryhlpKHZiNFW7PLxdm+NsRoDSPl2y
RirN9EFvgY86I0G5W+ZU/DoGqPt6TP3HVzTwi5nZlb9Bs2KZRksSKC5hDzBxW5D9GnKzWExH5AcX
GvKOwn7scDgwP9t9QgQ7/2SzfjjitR0aVptU9I9Pwxn5NVZ65ezPn0MRdxxUP6dKcilCKRlyWFkK
3ij4t+RowtVT6S8LrpxdtARHpV8ci36eIJuKxh9tvNdmVK4cdOW/oXNzDtmuR+jKNxL2WbsjiGZD
GvSJqJlJeF+nGCh7b8yfLs+O4pyRMu4LK3+RWkIsGHJq5a0iRDgTGbWaAdCAKAenUUMPiyJPyxJ6
rWjSpB1uFtHrR/7yzTX9tMOO8W9fz+TNclYFnooAoaGiPW5mppLtNrq9AkULK8+Lywkwrwcu5fiI
4Sshhk5l0Y84UnBy2B5/KdM5VcBDcy/rxTbX5N7Hm7JQTsV44jZ2WhTsGfWekGQ+5Juc0ozsvu7W
IJJFxWITRQ4e0XVPnSomGPwXbpqlcJUTspyhi/dgPbPxQihbqVwcg2eoe4fzT46i7hWiEUyLiKXv
Xxg7XBz/5t6bkI/drsu8DT51k+b3qMEXSuZR4YrtxGiOhb6UwsYqWhoe4q8PiNMZB5EhwCTFvHZj
oqPSx629OKh8R/pWMxd/sRPecMi0l73KIoufGA937Cp/q/f1D4mVuQgQKMASzsCNnR2lN1Oufuxu
DKYvOE1XnW67s90/qtkF9Bb8KIi2hoWJdTZ+/h5h8MB6z+NiyQ2hQOyGDwR7r9ssqhY/xCSP7Ohu
DNFljQvoK1XS79Ju12fwRvbtzfPKyIZ6ts+5u3epX2/rRng7K+EFK33Zf67w3uzz5oxP00CdeANV
nb+tBb/VIU4vYncHIiVu3KF8WyiuSDrNiFk9uGQC4hljR42aEXMV0AMSdv5dEt+zjMqmMlEAoPG5
IAaEI0ScOuNCbNN7cA1kQLEOcb23gLFrioKuBq5Xlhxha8B/AuhxtaC7+FKaa4OOqddJCMGAx9pb
J/dNS3iztTSYfRwvwtK1neURp98d7Z7yE6Fupj1ORvpISLKNn8zLYjfA0pgPBmSuo0QMmJ1xjJg+
m7wVTHzyQU76eUS9JXsVZPkwZr+fz1n8ILzCdG7NWN5e59XNJ3VHXF4/T/w0Ve8JnE7tMrau80gE
e2oeavXRcYWqaLyS3Pe0U7uNcguPg1ik2srL0rdM2mPYmR9Z1O4e8aNMIZXRh09UNBkphsNQXg5X
7medWkMgBRiWApSJYJIlq05G1WyRhby2+4BRjKg/dDYCCEfE1F8vE5eJp6L1vdP2Au8FLPWvtgnc
rLoQPc2ywHjUp3kIhPmAYr4NGlc4ywJdyNmKgbMOLV++k02PEoPd+NZXcic1ov5GUzd1DcSXKdaZ
8FM3GRa8+hzQ4RWufQqrv+RuofGmUMG051U98YradtKcD7RkFY22bVoABCk5Jz9CiKFhmooRLgma
yA3P3PME6XDWzpfUclHaRVTN2fz4r2rgcAyybBJU8lzPk+xpJp5pDViFQlqAerH+Xlo5Wtod6ngp
h6Nrhh7qYSJ+Ioho0eEgTOOZPX+XaDsf1wHKuQkkY1VmNe7kI4IvepFwOji0VzfWUGb4R3g2V9Cs
/szMEQu3eEpnd7dai19UEF+xPQPDL/Bf2YZM0E9eOQ8LcAO5JrPy9It+AbkMIqjqPD/qae1JdE9z
720UNw57K0sdrPSrLN3g4BfNvTaxAFQWFlgPeLJQk+MGCWMy831b67/O5sWiBOlYoJeYA2GBDmz6
/ngxz/1dY/114p2dcH8z1ksqkxkKDlQTg9zY0pXt5/BSsJLQ6I16TnDZId2YkBKijTT8x54d0bqj
ZMFBS1z0VrqXOpwwzMdRSwaj4w1nUH03jLauiumWTro4Tv6Dm0Z52sVVAbVFNjSPFad2hAgmTb+2
RTmQMdDsFReBuGxgIHsb7YPu7G1fDcGXz+rBdZjoaW4tK7rbufK1Gfk4CeOSM43TYnqR9HmNCeZ6
nKZD1YUCEU5HJyi4PZsOms48NjfDh3jfeRlJ+hn7H/AoAN3A/ZMe2jwXsrJbRBIin1z+jRmyVrSh
Zr96AdVmdJ5X+1whlnSnCyTnRVegHBv9CKbK+g2svu9ZMPzJ+P0HbTbFp1aJCKS4j9M69K/JuVzG
2XbE4IH2+2lWn5EctV+m8WkLbPdCzqWWlGJss3r1VaREnsBFelb4HOIG5ODDx+zSyCTT/k2OCC4z
j4TGFbkejxqgzyVv7y9z46gjndbhLq61pzhcCOLuV3F2f2K4YkevPiQ2qFsEKoRLrDR9MmVuU2jH
zHG22IvTNaHNFtXSZ2EwYsx7lpo9ZpPUTpOJfpyX8P1Tr1fwkAW2PBmZG62Dgk61wyOxjklHfiwR
Sr6+nEWngcJaG8HeGHDga0GC4c4hc68nnwpF7SiWwmx479vSaMJ+MZFtnQDmC+b1/pL5YGmKG/WJ
CsBHTYCt8qiC2sOTf2Unso7eVfvIx4vCVSWlnE0JenCyvaCo4OnAQcs+t4FaaAZsP3GTDXfUh0+Z
hoAZNSmaIAqXOmPrwnkEwrMDICAT0GutpIxQtwXrImnU7419p43mpP+JU3ukJZmwmR5wUqHuKeZB
406MpdDjXjo6mMRvZxSVmcIWOSeYWiuAjKhBVxxkt2AEOLwgYzPusFxMS4kpRuIxF3KzlzfUyhjI
pK+AJnpxP6l8xrSMA7TjH7Nnyoyw6dQU45+JPPmATDG8PuC2yAvqVvc5lXNTkENPjMjYzV/i5f92
0soiFpJJL5f6drlyyRyaJEsBlRaV+TFN3qEX2Ibr49nlUyUGb69FuAuNaVCimy5SLqoI/PBCnXa1
Rf872tQEQPYVgpk3YOsGSfOEn9zU+TbJT9lGRo95Meej/sXqXE2/XK8833q0gtrOon6QHDU9Z428
oA4eFBdxE4s+Tvo4GoH61j3LCFkXkWxjQz8mqpAS28PEDStIEj81FP9IZrlYTmilgj5aHTGxALKz
7LX+9bqF0sQJXYN2+IsEUnAnT+vOQw9ebMqP6J4RBczTbLtmb2PiASOmNBVjQxo7ON2JH+9l2gH7
Jg7kZroOlC84HM1WXrkWEtUgMSQd49bOsmC29fo2EUYPpGtXXGsKFw8Rf1KmLdghpFJChkfBcHSh
prZIWR9oh9ZbhG6pdnzaX4EfuCPRlwPPNzmoKRyHZ5ApsjnTg2fUDAaWrd4XZhh2CasVNXSEoKhP
O+yCgifFpDkP/vB5Iejwdyo8f436vIhRXly7GWrKjUE125Y7D2XanqWnuv+gVdr84ukYzSTDtka5
2QIFCluXdU3dzx7GQ6E0Kn5nkwTFPnu3HIp/HRelOfVE+4G0PLW4NcyjHJCfPTl9VDBSvO6oIJHN
XW5VvYcMKjzslRpTMMShcc3H8oFmRfsdgYA2FsrOoTL6t4PfOv+PPmPxsKta6Kk+VDvmHNq182fs
SLvQTR63xvH5f70C/Uz3q8yPFgH2jDCBlwa5kaNUScsaIRzBciVXybVU5+RSK0JLCOQcBz+Bs9vz
FBNVw3DwMyrS1qBwZKAPnlaf8CaDcazCst+nbQ6sNB9RbspMMtt4dLFfGRXZeH6xUQi3x60m45sN
0381Ly5jnQ+Jdk1wUTjzzpQlqLmlDRC1GTdNHJoNaPFZwknUKu9RD/ZaedzZEpyYu1DoLwps8D5n
B16SGxwCEfMBmounb4rqajMgmBGaoia8eQ5qWhIfCQZhdNG8zX7yqhFNtBKfHWjKSGRG4OswSAAf
gX30rH66R1nzG7zhfTRdAuZrle4Ei1/jCiYMc06eDYlFQE1m/9/9zyi7I08nMQuI/s3GMhwPVLQf
OucH3Qu9sNmuaYBiQ1H0ASPzO43u+llzniOzwB2nWSAa/Uc0HWKAa8SFRo3W9v1vU+6WMu73cGLt
/scSZv23qS11CaK4KyRONd9jckOZjPL8Kyixe82yCrzbU98vTd10txV71/pYJkCsSOD8kSHGOqif
SeYnKO9reZWmOKMcqeGNJPjgiVqG2qHSKgGiyKss62QG8tWQ2u/FsQY749Q/90wxxdv9TJI6CJ5h
4XFXu5G6CGa5NV3NmTGmQBWll3nbb/Ha001wt5cMNb4qvVBVwIiq4TyKYLcgeQqIoH4dCWC30wU0
ly3wv2epknyuLygouJUJQQZnQH+TcUUZcppffq2Cri1FysT3VJa9zziGpQqOcKWY+D/h7qLoADNU
Lkj0Gm4RgG88CIq3yDfb2MUFcmqW/flJYBaYocE8Dx+6HVz7BcDB/3lV3hbDjhYKuLiBxQheXlW/
nMCxeY5fIlKubF2AHGieZPdReGu8+vXxD1VaOD9HDiV+HaQut24jvtYoyuLnmDtrA+IwqvuEXGqw
FzCGRgxxQenuoSAt8OlLTc5vs9PdwPQPYNrZM7Q06cAoM/HW+OYYM5XdLPccK9si7//ps2jkKNBj
Cfu4ofAfEIze73Jlp327MB/4hE8qbVCTKFVWoNBHWw0UjD2+BZi7nB37kkDK5pAwruJjypeJaUXb
w9Kagyw0wlAENklcN5/rKMRnM6t7ggN5BEOryD+RGDANGXoN1exGd/nn//7LnmyazP48frCSYAKF
xRPdGELbLclwGLftdcDda407j4EJ7026TVwBSIFmKhEQefcF/h7/rDgxbvfWOJ5rDqPU04ocpQDp
iS42WhxvkgHF8k9mwTNmKmbH09Wt8ZpEHvGXPkyGRnkgEA5lu8odpqkipwmkkzgFivgONTEBFlZS
4y0H1JikmxZNu8kA8uxcPtQ3KMyjuSwe1BcNjgLTTk5s9YcnkymvQ9RW0KeFp9Mg0YAwjtAou/zX
V/ZLbTj8QsMsWD4Ne+Dejv5GRR+PXwHvrXO0Z+17Eq2XmTvX/cC7kx9iaz3hQjh7NP9Wyr3hnS+C
CmgxbbAoNXznZRB7Xsdnxfeq62sL12c2UuLWMiglqmvWp88IeRZyUVXdoopcEC43p8pESCgBb010
mwpzvGcLso21N4TL4DHwCuF96AUIz0IesXxMJ3Kx2H9S7/fS/+o/+EuvaTS3khjdPp7do0H980bJ
m+xDB/cZIyQjgAQBfoNqpU/Yojm55BMPhlRFQ+dCETHI11yZ/CdF4b/kVXe2x7qUKP9aVRnrWKqC
AIikaXdbCgs0Zq3wSvYsaX8gabzl+KapKC2QNmg0/jCscmEX+280mCtbX43YCy7cNUK7E6EoKm7p
WNt3BXcLj9HAxPcFFft0F+UnpMMVr2QBjMBCF1rgxEbRzY2VVO3tUrTjMRJQVH8ZllChRcuMi3sP
/N1A3rr0avBvci2/5GvXrn8xjHYX8X3m3SbqzpydMqj887y63ulfoK9iNVm8Km9LBtnzIbMMU35V
g76exdOQGKxzBotEwNmyX6utXHLaQrD9iMLHNQRKs5mDT+VNYw2Z69eUEQXfEgEkGNaY/6px5zre
HGBNXK4EcMrmyknvXy+vsy/eYBD6SYlc8D68mt4BmDohyrs6vD88UYaMApOO9t4+G2uMthSZ8yBg
51Chw5/CZ5RciOkbMNYQO/AvMEOAVC40ny2EYSqvai85A0hWXzgiJLdxd64sqzcNxHkTPMmhTfP4
he60tvuf26ePdBADq4FECp5Fu5iT1jfOcxUqt5ojkSJPEyyv1CTSIK2SQimivLSkMIn0NHY7f39e
gnAGi06z7p+iAfZUAuDUukPTl1zYaO6hQLW28Hd0OFEzUKAtdP7v2Zk3NbuLqu2eLEc7liT5BVj4
34qGOONZHtqo0TwvL1WYAL47d5u/+4/Bok0G90hzox+4Vy0Ct/EK7oQItuSmY1Vv3b1YJiC55scT
cvVEHAUJES8ZfD2GevkfsgKT3U5sfFcttnJwIrgabCVGxjdUcj3MFkW7/zlYzyVtaXmYATLCdL6w
iXx54SbjLgqbhfrLiTbwTMzB+6I7HqwODuyCkurZVJrJT4UFjxIj1SGj8UHY47X3wL8DAa1RKd/Q
+IJk2daz3CAYJBvh42bE7bUGoFMk+/SNjGZbNAD1uSdP4vwtF+xuCnUOAG+NybGvEouUF270IzTI
w79yn6fx30HVZ9yi+QlEgwI7h+WaRaDYFsQXa8fD4HyHgmxqkZhKI/T4YA7caktTBnwVbtliUrG1
v3rayjxDlix+su93KV3sP4aut5QXwKdTdt1ftwZPQYR0knt1A7fzqIEdA6Z8zyPefqOTMq9MrCpJ
aqwiCcevUzvr3rSK5OL3Br69M5VU2MnqmLvWz/S+AyxAhyu4jyW/v4/+mMSOpOcgWHtjSXUw2+2D
nr+oV4z4cY/D1QXthJxpvBVzuFEqQjjwEdutIxIEb2o9eOMuu+J4WU/TlTqSWRGD8rGgdnpC4i/D
6O3iOCBD0a4j0KViRrYSC50TubiOgl0xJc387OA35DDgH2+R1CcSeWTVZa8UmUbYQCW+z4Eyiu7V
z8p/MKWn988BA0zT5swDC8uVd1/tNWRGfjvnakw04mF7Ukh+ZdVMP1a6nS/iKxVURcYIBEfSNSP8
44pRRH2bZ6AGAaFfsQuw1i26lb/2JS7Dn2/A/2dGsqi6Z0UJiZIr6+WNopcOnGLELObUr9p7km/z
4qR1NhW7gAL11kVtvindlxULoEU1MQyT5qAndjMx1wYePyFpahCkAGVnHZWdF0qdRyjHLOUSZsFR
biyv7aZFwWwi0dfT6RlDj9FnHvA2eAnavMJT3EHTdldrt4AUMxkpMs7U0WsnpC+mbtn4qZVASKs2
zRct1d9MFAZdvEnLNbucnVDtHbRYR4r8D4ECjvGGxYcIyKe5NeiKKQt6oSNWSGTuqilfOOYGnUci
AwMVqyNPSX3i0r3chMu/q6L+xAA2i25/dyeKkDr4I85rM5orBZvCV+uY/UgEboTOq5vJSA3fF6yd
ies8esLHirdmqxqL55BnV6bGYW0z8NHJ5ZYHJiQjK43L5Iwo1AlmY1FPXzwR1JRhO9Jtm/6i/2Eh
Pos3Q9zHrn43ugPpPsIi3jlL/IO+lMU8H1OkE169ZLaxuuGCCwSmVxxYXhbmG32/jXRBMn13QU+B
tiyKCzVGl91H+0oUvRhCdV8VHEG4ux8wreKGgeT89lapFXATtsFApZ5rqDW3/IgRJcxYhkMe8ufj
DU1aYk7aUfGDW5D5DeZdMgkpGrAI/IcTWpZN+CYuNAtsuQV61iu5YWB85T7nE4RvYbtsAFyuVo5k
qbAfFLi3c6v66pxEt5NfIDIQ/rwfR6FHYP0k5I5G5bxky1co5DinYjgg+QWnMDssR3FEiVcgWa3j
O0ZM40p+jDg3qtb8swifPGiOeb5rLb/m9hwwXUpSm3dVRl1HXE/LWHxWiHIKJR1b+enN8Zngj1zP
0EgPrmqed81Ja1SWbv2eG+0W2c+wOOK5CVboG2UW9iKDKb3ov8/E4oACvgOoouXwRQa+JNg2TwGC
ctVMtQd313tba6EJ4/poKW0kC11B+BllFOmeAlZ/qoH6X9RnYDt1gv3R0z2clDRTl+s/A8ZSEZuU
sAlSOZyxl1RRvWzS5Tt0nllY01z7LftHOn6o4G0hJeSn4yuWI36d5z8wBA+UjcrgHP9RQS5OFQO/
X2fMO7jgX7/JVTkKrf5xOGVp9AbqJtYLQM3PeVB2kASLyC+gvttT6do9bS60BAFOwYePlgK0NuG4
FBplKHSvGws+8jvIILG/txi/Pxy8eFI6iGJtaqgTUx3EvXhSxzXQP1vsGErHDR05yHjn0PsI+abX
ZP2ng7h0Ua2SCW1I1nHTvHd/KDjTTMGAJPSBXshjUIweAJHH0Nkyi1Uz2vr7fiDj6v7ykQL9idnc
sVJTNQkXtdyT6r8WRyDqHn9+dx/0dWc/QwJE30ijRe4GW4T2t9bi6sIR9BTjfCCjhaIu5k5hcEt7
PJkJwrbXV+Ve/wFaiixOW5rad+gRkjiMEYm7zNhhNWz1goX17iiNJWirbn4nXSOMNvxrHZdLKvYS
GWDYVpTpdWZioJj33UBjmEJNdzRmTh3AgilImz03s2ua+TbgDBTNX2iSmPeoimAD8JlTpV+KYS9D
P2NRMMxxFPjRigqF0SzP69dRGc/KubQQyCFM/TXD615mkUEWIw3HDyw8SOA5j+qE+iyQLRnNtB7u
7tGJRIJ48gw2PMHyCoPlUJXaEZ6qhJEfXpMA0XJ2uE8fHNva2n02aorm6IhD9uNHrNVtgpT3FupT
LIB6cWYlNTlGD6eg+XdTlvCDMEXW7fua36qmfcRYbe45cFxkRZmNwlCE9pTP7Vt0JZokqz1hcUmm
scGPnGUU02zWi0knJ7sB1/TSqKAEmLuLYCT1mdNx/rbsjTksUbctSokuX4bPZQvxvETgneR8yAJq
+v5kvfWoYasMrvPXItvvl7vqvP0xWHqBDjXmu5mUrhBFPjZNey87RSEQvOqZYw6SMTsRCRKjtqjE
jc5n0bFDoKtkyZGKs9Sr7XpMHsSCPqW/NIW6Ms9eAszea6B5VmkIKECBe5xoaG5OmfkRw1ISN0jq
bPhtP6V4MY/dP5eQVz/K8lzamBJDiOfA3GEoBSz4g81e47AAjdly3a9y82232nWqkuO9HfuU1e80
bZ7O2e/UFZc/QVAyUUbpm/1ejYMhdVaK1N5wuv0y6/NGVQNVwdrLi1+T1ueYoVLvjquJgPb1Q6Xk
7MON+JSyc5sBAuezeesd2ntj9nPrrWtKUi4rA4CwNBlfR6xHQlUWLsgNapIJGSwHacJ3jrNcATuD
4Qr9gTFCd4BXlsoL4Ajjh41QBHO/SEcfUvJcBR68XaAlxzNkAOkZBBgPKN3V6/y1CEVQ2n/YImHa
DbrhbX/AJWjOoy47+m9L1MSB2i/0+fPDHgFrlxul8hc4rKo/kj6Fx+scCgTp33+L+cBwyFg60Xs/
fxFMpX7qatO4ASHT+RzqfUkYQ1CUVfTOAzkH8mORW2WN/IcoGUwYgbZImug+wajL2ka2OXtm2RNS
hXLX8kN+uo3vZO+DjxUdSee4/7ofWQfGERvV47cA7Kas+TxMWhPuv/JfI5sFLjP2xtnsgdCeTi1v
ZzhqkXeFZlD6QIz47thLWbQny8JrLjg+7gTCtGcjXrgOS58gynq55pbPmYNa4sep90SnMs4B4n3y
iP2shBUp/iQu0QWrN87hHmEe/f7SUjHpCoZ3dXbBrbPlkvC4c+ObT07uEVsVvHQjF51THsHxe/Hk
h5gkv8he++p+SpJpDoGLqBOBJN4MlHIhcbpr1pGbk0mXTRX8rE3pNWtN/7lXZTuA4Oi32BWLN+34
lsBgf/pF940X3hPdpusnuaNHGrfcouTRL09TrtKnXWSfSjcSB5v21z6Av7WtraSF43EG3umANgFT
vsyFxvFTjNL6UsKhmRs1yCECWvu5q/z2f2sjxvLqx2+0Uk0SDvTwd2q+MLelznqkgAFIbqSDrXl1
b0FpDQVvXOFFFS+tXlLKiLzmpUzil0kA7A1ZfpxIPqcZOVz9Pw+kT7u994eD33bf4JIu9s/RGwGW
cFCeAmZ+RpxGPavzsnbW9GY1OqJ2zm2Hy9VhH1QKM8bOQ6RPN/K70vJ7dwbuyHbZS5mt8Shgh6tO
aI8n+FOD32O67oly3wUIKRgC6qOLZZKBmPEL1y8aZq2UISrQzbN7A0M4uv+nF6K5AHWprrTH62WU
IbRkOGccmFjT8oxkz2iK9N3kcMnLSP7+YdI6qGqRwuLeCEw9WfCY1FPGgzBQOiMMsu5M3j7bDIJv
kIj7rOJwShqxnTMK8AWUx4LBLe0VN62ul91hsnteyi11L4WhzwGfASeH9rQr7Mk3SvSWcoXYFshv
uzNYyphRcwhzd+9ySGua7O/Ho+qNzr50vSILqBhoc1Q3dbV0lW/heeCGEXP1BxdZAybmpCzndl2+
eUK3y19C+rvYjwpcfATmeSlQuLhYCI+vD3XEMphyr0PT2kjNs9MXjMJ9k5O80CGLwRB8LGM8BZ3e
cdF+9lbFdXlCB0o2/81T6BMMtmx96wOg/HF8VvPDPTh/ix4wbvu2bA7Gu5rpV1qicXxwgSI8SYTq
s8c07Fxyoxr50t1YEazvWWXmT5YVriFdhXwAjLAI+L4uHLBEobmPnIidZP+4GOxlv/yh8ZzGGdJt
iv9Y/N2zCs8/5tBHgi+iV4+Z7ZQgob1fiYnCHU6n9BPNbh3sOlGSMmF4y1LKwd7CjdOD9WJvjQSO
7vrvRxL4BfldyG2O/+qS35cEnGBMDbpbBPYCAfL6L7U9gx46Z8Tkz4epnLc/1VvV8LAxnqGxQL7X
2XXuhae44misB+Un7f1YAtVN9S/DI3VJr1o1VNuwl5oQI6rmBFcOlG5st6Rf1UGdvwA6L0GXOgD2
URVr+9qsQNVQeli5uxMt3NH1LHE1XWE8vw/+xRaUiD9qCBi8wRefzDHdvwKQ1rPCZQLeL9RKBeUG
dosVHiOuCCUGGcQZAGBanGFjx/wMaVB2rF3+3DWJ8+Czc/I2OvqWwut/SUcE0eeRh23u5bVrGq+I
vb823ST8Ov84Occiq9SgrRCXb2nvPMVdKj/1dCMSS4HqWGulD2ZNKVzxpN0umrWk9+aSpBQTcPc1
cTjaBLolNJiN9S7s6ZHAFDPOr5gnkNc+EJ6QaQnPB/2sAs9VhjD6aoGRuC1RvkuZZLPL5zfmprQ9
CxiF9+M0/mrvRsfAaRioYUM8Pd1jGnUJXIh37a+CP51hKlMo/Yo0bx58fGQYGqxIF+OOXp8LNnGK
Qtnht6bAbnMCmdBd2T+PjJW8HHBuuonv6togNATcsFUO0hOHE+eLCexhVCa+EbTpRpEl901vg+qi
ag3Cc2gCUKQScFSVDKwyVyuW4YMITa3QV1yjEUA/Fv7Gt+APbLP27m0a866isNntvEX5atPtqZW6
QpLdMfhwvJQzg+bl9YYqMRU25OsJUaoIto4gabhpdeBm995du52T1fe4Yj7dbZgLQlS3Ft7JJbjE
J8mP7/m1GRkyQs5gBUPg3Yk1d/NUTQOfJQdarJcrxLMqvnClarDCYix+uAtoHbS2iGLWlw9+1pKi
wpmnNc/MESOGuenX4NsQPu1hZqpsLeuQKdha4ARL45H5PixVZ7VrHArAjNA/koJyP+d1N+yrak4e
EYrhhodeT9gpporcflSNVEEDEpf+91cntXrvN/3IiQHYNOzYMjGyR0KL8loxGBjsbbF67caq+r8A
NWVKbypafrf+xRs8kvPYvSUVfr+H07fa1LuhNxCkyUmv/x4pVrhSseo5s5OzWskqaqwzBir3bPvV
7bv31QggiW4/XWooGRiqwX8mEk4hMYXISLXcm6n1BSQ3pMd9oe/t6VViGHZD+yexYCSlHsQC9Pzz
U/itqakPZuHJE4PokpA8b8zd0m23qLqhP8upXRA76iP8Ovad+UyjZ9LSqpS8bs9gSiLUw2P02w0a
nXVz78Oa8tFH7ojrmsYHOTADoT7NgN5X+Im1YjapggusziNvpu+udr7h3Xx4s5b6MPV0zXfTq2At
EtL+iXV0Z/uda6/M5f0EKMOov8OzOKQaFvb6k7f3rVVWL3QockzOqjC/E1YPxOpAiSyYDltBy5QP
R61RZ0wPWQoMBVBOSlRrko4PqYoW6aivxMSLwP0TBS6L2OhutvHQ23TOcA7JgM0J3vpPkmDVGLMH
C4ssFtOa0kgovpa6Sm6YP9kcvMG2W3qbSZrhCNphcdgTUhGRrvULzq5EgJKbYZICRiP4SZEBFPfB
ZAlRPNJ5awmZpM5WOnrnvwK+Q609nFU81s3w2u4Km24SWbE0zieSlcdFctn5pEnc9dolsBO+qqwv
fXqy84ftuMr0phBp1EIxuxHW4n9Nhq4Or/7ntg2IiefiJX67+4uFiqZ/qB8HWUCpZ4o+fJDPLAUf
GeqeLmMam7tmOzMm0uwro0YdDmSNTSmOoWu7ZYyTcRDQqGsAL2qOL0FevbKfhrKMl6Sc0HqvnVag
0nYika3JTJqkWQudiJTnv7zHKhxfOlHzSVp9VAxN1JqxBJvBJadifRJkYbx7AC9A5ExSNM8vTO1N
drQaaRv6MYaLsasXfycKFgi1PWi9xMSvMyrHhWInEA4aUNXs0SKF8oJsEU3t+vHyzSQyA+q5MoPR
NuAkkyBDe9hcR5PfhUii7a4XNSut+ZOOeGAKCD0h4OURcEjKZS9JZWpw0vkA4Bct2WOxeHCRDOzo
VB7rWFE5SPBjUxmjqSnRbhzN0caszZs59OHRFQWaahS+8W64ojjYish5ca1vQ88rvtw6ezVlGDIC
66RAy+6VJx9w8zpIWrqunndblYzSG+qr+rl7mcPvCiqgqfal6b7aRWBRhBtN6yvQMfUd1F64QlQS
NijemKLgu6vl3/zaL0Vg1Va7Ab89Lj0f7+b8cIeDf5OhmhIsKni0k7CySBQ+Gmx0cbA3yed5AQ1Z
nMTq6BPpXkwwtMG6K+QbmicASqi3E0TaQcxqFsh4wercklia98R5rFuY1xObAp+yj3ptikbdHu+8
/gBq9I1M6DuEA2dB4+yeInau9ZU25cjH1lerQgaB6IiKHzBJuZH183OHrXIj5TYpsV6Prp7UjZct
saKkrcKuEYg8WVY6QHZ+wBWfqPlkdoUrRF3cshLyD3z7xY0kF36v2zSnpjjviyHz6iU+gByFdPXC
KouJL+ILQq7NQEDToxgEJuH/gJGHhFTq6YOwiFRLcYdNsV0nwx02f0eEx4UUahIhf/fkOzFagzAB
4MH3uFHry8euuAuxdFI0IYUOCNgLJ86wCX9br3w+/TGm6fbYk0E+kKTqj3WJw8bsmo9A4/gJvbB/
E9OScmEumPE0f/t32dr2+D81tW6mK/xPKAovBFIl/l89kmHh5cjQ0rkXnEz7MRqTt5cSKjXd455i
XMeKsrbyyI7ACEw29gJ9ldICCxpzS2/j9uaKcnH6mGclXW7VpTnW9wAdPN4qSAfAZZS/GrslIEwe
THdjTBqVfqhJimo8dKAnEoGYDvBKXvNeZPFBhCW2AeuZLtp2F5cOPipLGBVVE460QZxDxncOn15Y
PK+HhpW0n+WCjYgev2w2TWgw5aRMcP6CGOy9pB4jHns2oHMK3Llk3B3v7F+5t3M2MM4iABY5STBS
rDcOqxvsoT0uWjs0a3oNno1dNkao1h1mZ5iu69CA9B0h6j9aIwmnJgnVLwgobABNwBZlPTWKcJb4
5O0KbZ74CScH15PDie5vs6WHJzS6+Wl++k9+rKG0uVimFsT0bVCXtepOls52VWXXJq2hEJXlVO9J
lIH4rIzeWHtmNZJxoaAcwHmEx6LUA7ZYN7SQk+zCmEjruyJghrBC0fFZfqZnt6mIONzDPc4tyrpN
ZlL6yPJLYh6GgvhWNLeDx1/GD0lFs7iXWHou13xJrPoVg/ef/KHN490qvEQ3xsVDwo0pAd/k6jfS
OTU8qICgtmKTS2Hs59d1Ysha11/ELx9QbmQzRDeP+4nWOsPoKu+7CH6KLhJqbxGjL1mfFt83f/+R
wxjBpJ576t6x2+yfJLMqAVYKH38IytGHjuQ7KODaLwoP15j64IGgZ12PipB7ahtWkk7oue2LPL2e
6Y/3lsTr1GjEP1iFmX0gfzejcXd1Btz3G+Fm/nf2+hDblUsTWoc3KWd6rvwpEnyzAVULQHiHknpK
oe0Pl/yb1vckbQdr1THW7cJoaLvh7FSma28Y0fbybDStoSpy93tJquTo/wLMrlYhlv48mgDNRlBy
UsRKHtKdyCqyUqs5zQXO3WZkIvU4JuRdUkwlMeojTeR6m99aFSe23VE+EWs6tQpapq+Pdis4sx1R
lQUbozOolt18p+zYRuH4QKxseRBpiFuyAVP6CjBZjiaiM+6Q/7uEkAy1ILxInvuQN7qFjhuevQyH
kHPUWpdAKlHTXmmIrR0AZtEJqDUc6TcVjCAaY4uG7JoVp1u0CyDlhqQG55CAOin6Km/sv5hFT9nx
HbauSc0D6JB45eXMh+qiJCjQUT/1JJgv5DepLt0ECoxr202u1XqTRt8D3z+cg1r6nPBhvDJkSonS
/p2ucyn9H017fszb9boc8j9rg2+PsEKcaXMCzzJRT3m2fxLkyzjlvCg6vwUwz3QW3Xh7R9wMeF7N
JsobpGZjuZesLECxoOAoOkPnTZvmgbfjbyYHcfiqdcaYW3R20+yA1QjFhBlBG7B1X9AiutFA7I+E
KukGdhbi6DCNBapCjipptOr2WGL/4SilFzxlTEI73Q3xK6DmUY7dzzwTu8X7alJl9joYHZ28qvnk
F42KC8kw84Eybgjd3a2GKl4xxKq4637EdXEIQ5YcmMh6qZ9w4+967Gu4ojhbb/6kAR+kAVK2osB4
XBO1fUe7eM9ah19iQvLo/CfNkO4beagnlgwaBg7CrIdgfOdMmffnBfecT5if74/rdRQLovRPvMRw
72rCduWq951gmGMOywk5fLvr0LLS6kMsqDhH2pLxlT6Ij57UGrdXP6g8yHpjMsvviEo837nXLUU/
Lbqofuh8pQ/oy0BVoNPFiVCiAj6bLCS6R5FHe9qrU6GML2mCC4Z97AzOdFOesYyHnQrep8HISlCC
1KOQ/ZNwzynKnpht/mVBquSLgAsstJVDa1v/RvC0tHpQVAStUa1oVngoc5kERseBbUP1LTnSLci0
I3gielOmJNLu3xJk/G1f70Cq5frVmS4qYwlz02VradAMeDe1Mg8RWITf7BKTZMFpJS4QIALKnzl5
9pA9VI+5bIlWMIuT5mKiuSmIw1XsmaNVICteL9X5pxX3HiwM4tzFlVFP8EkXnfz//pPKlYZmcffG
EujmBJq/5OMQlgOW3m4E2SKSCcyViu7GRJgt7NmoiPxEZXhLSCbaYCgRMBdWOgzfGlbLZYibxtr2
p72pj2dNZt2QJa9tQ6P43ePuPRHVgVRy757j4InnHDH3cUfyIqGWa0EJJMmYIxeY9vNi8pL0xmXT
dZXz6vElUm+ILWL/y/+EBFziIR8EYIqH1O9uvNf4HIscMtkvAa5eoqgP93nfgxQ6fo8wNEIb5JQm
wBNj5jfPkuLkavYn3OxkWR/kQDrp7dUc6W9lHkml6bJW1/z6ZJ5/UFHhMXKA/DGz9LVK/21qKDzo
+IAZ+B7CZJ+v4Jhea+Bu0oMKu9/W8y+uBtmwSBW++386sP6AQggpsDvJ4kR9Uob+JHASvqW/LuKO
cNNyxEFKVZywUWUbxEyMUx8hemu/ASswSj/Dc6ogboyhZzAlNKWsbf774ydeIWpZYSztI0V5VZEg
G+t8ihOqvyHbmIL8rCExyXKDzV/PJYqHH+je4usTxYxshs6y1WDoXmlR46MRKPMZqyddWMnG3cxG
bm5w5dZQ+MHrXN/jjEFRMJ8iSKO4nqV+Ww+weIYofmGfTWKO/OprWUlqjV7k34HLL57PYunq9ePk
dfOdfxuYkEpsc8MveXKhEPvDxHnLocqKAQkuNdBHZsku6htdfd/YeY9h9EeiKo6xPwUGkUW92QOa
nyrsJRMGrO1ed+FGmFL3Wvi1SH79y6nfSRMQD2PWb64rQKA9qYQcJisFrMRrUvTF/DSXnTanNaPg
T25Vf0jbdF879iBkOqTu65DBK7WNy5xe7IayMVKfNIcVE2x1a3VZhUTT0qD8SEyVL0sP6mH3aVtb
9Nc8MU1gOCvxbzglt1eE3UkmfGoBc/s1psIfOxpHT6BEdL9sUnjrZvxO74JPMsbHEElQDY8vyvAu
EYg/BS6xL++8RDcAaudXjsAlj7jtzQUcq0rK0/6dpbchT0wZyzWY4NYzL+8dQJvrYUJI9xSDcEdq
AShFyWEdIR88Yrebec6rXQrzsIKyllw15DCTzZxaRTH1KtcOYG1t0eRDojhkubFmIZRC4zSRVnKy
OYapqt/KuQhXaajWnW8sttbTN4QukCzGKnXY1g8eZ7AYX/PbD8XQ44psq27+fK8rsQA3sHFFKgym
CEH1x3sm/6/rlwdr0HSZXMVTne7G1C66KY3F3q/7B5tqzfdF9k7HhQVKwtZ9FnS64LLuRwdgAxrr
OsvKAmNF/gPez9lVvu5e4/UXL40qt94PtPSKaun1w9RJH1AbXXTZ2i2QYKsXPMnVCwTI1DlXWwXI
CkbNnfAAEZGq+4mv5Np0YSXiVmQwKuZVGSxV9oHPQCiJQ0jdtho2ORVmcRYJZxgTpkm62hyEKL/u
crskhUcE/EL0LsSq7P/rsVbfdNJmWizcFM4djo2V5+Jx/7kzEs1R0T7yC9f5LSh8vmK7Epemqeyq
VdypS+tL+ROj74Q9q4LI05hMVeMYCq9RbHMP0xVjwFobx3veQQGI2zYoccJ71VSKsKG5mqjDP9PW
XcABTIN6YKwINXVU2Q36/PIBIXjnyp/T9AfJVx/Bo5UdTLo9NsD5yZ2A7DWS3E7ePxyduDdiobKA
iBPDXdf5zBEsaDn2pXmOIspYVJoY9d62bxjbI5nO5dAGfRCFGwR04xLNOXy6uQ2JdilBALjahp4f
YEz4Xypu9aC74A2qCq/SN0lf49XNokWXhU4JxVk3tpmY10aYUj8UoI22WB5PcxCpAlHi9tLb7Vcp
5HY9VzEehpkIVSder009Pui7UzaKPISqxGAbLdqcbNyeIY8u4SmJrL6j2SjtrAFslqYFAr3GXQvN
HjgNYn4CfV7V1+lgeinvwzUayETCn2U1ACudBU4uCZ5V5EUBCXehFDbgub8SF8kFus0oESJLItPh
ghpbMS8UagiVMyIpIELjscKbXnvSAIX84ksioeRWTpiu03WXaMGZZXKhtYv7rz2ocE0iNxJ97HOl
bSONOdnM/velOzpMy+Us4UxjV+WjhBmlF05baAIMt5tR1E7guAfUxJpi+tdJrEeygFh/BTFaeFkM
Ite+NjKTBDjdcjdz2P7Qkz7gbDJKBZ/+oS39hTR3jzDyqlK5jGkDi8+4s5BRBYwwvnYXbu1ng7GD
aYh5f+MbYaMEoNwTy3lIw3M/1qw1P0paxTjLzO5s83acumu2JVII9G7399bYTCEZgM7h2/XpMGN7
bWrL6nMSGOEC55T7Xw/+Qt+MN4UxrONz5aM2yiVt4TbLx0bj2MjcMZ20LTq9Vpwl7OTx3xPPL9tI
AfFiAvYLheeXwOSW/1+QbsJakUqS3vXxTnDsoRWLm1nkS7qqOsvb835Khszep84JzMNKH03EEG87
PZISGo8ri07TA1FYZDdayUL2nJiwswYWY39HtvPtlEYiJxw1m+YFh2OlkGINeDabn3/nGfvhfLvS
RPjJVMZy/xkcDcM1+l1KO5wI9tc3kiXskG3QyQ2w8TREc5nvCse6UwvJmlDQKVRZrNbimdqX0ID/
YCL98fDvPVkfrHDxgHBePlvCVGyfxqIDiZCJiuNCT3bTw8ruLD+rZN+jJKTV186tvsYAL3Xkf11t
ra+vua/iRLXpi/o6q5EQLrZPV7IFPAeCiM5s8eW2tvKHHaOfvhpP4Ke5twChZ21Of08Gcsf333sJ
qPI6mFaqsdD4M14qJ100UqSpNvu68yJimygkFENTMvFdvstpSrnHYuXR3HeLWzRMMpuxnQPW7ykQ
GafjjRzklhP8Wsp/dSZ4l7Isktop9/S1zyCzQC3Hg1bJUe30vcbO3xkr0+xaKdNJrsYwqzTilavN
j8teODQICm9JVasqyqkDcoGovwMDlvmS5g9XduT3OlxmUe/7yWsC3Lz+oM7guCuqtW43jpzGX3E5
9D4GlXSU4yGOAs7dRsceUnnqXdJXkFLMkkWRZNce6eS5B1Tj/zDK5/9v/Uc6inKIxkAkeVJ+yzMJ
r/3n+QJh3dpOtKBWHHH0806EeWbwfgMC03SkDyD259Mzytd4jtQYyyj95Pqw69hU9dzUXuTjx5/e
NXU4JO/27swKwXpND1kwqmjKd39P2ggYQRKGjNGU5XHOEGl2c09E2CMHSxWuLhUbFq8rTXx6RQaF
SO21PHTTFBN4hIF/VigMT9a81h0XBxZCFreH8Vkahu+6Zt/tC9cAPdxoFSC7l54jyG9vDSX61Wlz
lvv8E4UvjLj3b7cR8fXVSFrcsS07roujfXlvM8mRQRhdEKo3whufYxqnWPbxjZB00q6zVzSCXAKl
tQLzGTitYAV2tbNkt+Ae9IeSN13fhQ3w1UK/eL56DfoGryhQYPFsgJoJ+PSaQo0ewm6JLV8EOfkJ
zOw7Ttuvecp+lYTB72YS5HI4luQxhS/67zjlZa+wzGY3+Sa3tEokfdA25HAy/duH5FXkUUuVniga
OpiG/IMQWS2K/1DhIdF/v4Tn1zFaM4TlyHf9TOqRusnMLdMqIsNs2CRHxaWCinxqrqM2SZ+kBpdG
mAsG2QFQrz0PAglE4aq+ZNYzt009yc0p0TH3AvMml7p8INRu1Ns478VefBbP5MdSFJyqS3MiSNUb
Cwb90hGpRPopnQYT8rXWUit5ZD5+CMEo3aWsklL84UVGOw13nLT5AZaYJFo+S/K17MBV3AdESUh+
hBUpOe0ap3Q8W8TEGCQwpopMzDOBD08SBMyiWGYhjyopZjPoP1ygZOnJ5UCtQoY+M+DWdLxmBNXI
LM+GnajdlO3JJciCHPTzv5PtYGUlPC4j0tGOuHU1SzV/CAkmRY0m87d7Liy6PVR9bEDt5HIdCa3X
LgxcGZowd3KdP6Tw2cs4E8snqTPtWSCy0gNLDjY5+Y2bNIMPpHmSwjHmA2tPcHnT71nDBIdeC4fg
O2oNE26Pd/vFni51pBwmDUWSLOB/fG90ue2T/XBBjNjg0BgVNvqlnvv20mGmOOjopVfFFhFtSzV2
rgAnitJWHDQdoKuPQIJ3+6wUFHR/R4rdAblAs3p+kfc8UuB2ot162BUw/ooLoDM6xiU0n9YMqXlj
QQMWZ4RFUAssLc/1RCbL8on4cIfxk2Kc6rEcPDZETze7bJCKaKRGAmgmjM0FVSFblUBuKuyLMWh9
UFMe+WPE+L731YvMBstrHB+NB3h2Oci0qtffY658OJZaTlK/u0oI0KQ68pxcCBK7MvIVXkNrvGlJ
r0bd/e7Qou30vXPdYsHLjnxabpofaRxVG4P08220aX/FQXs8gd/z1qum7x6RGPHWuat/rRujZtmx
M8ZwnmySqI0s9ice7WLFWrEFQh2DbDxjXpGvO2ZpJlqarXa+d6T7nVTVZ2C0X1d66iAqPc3wvd6c
Ii2UTmV2YygTk4KbpCEIIGqRt5MEl7h35HmSlYH5PqXT2Ig5EfQeHoiz7PQ7VH9EV2upidJ3UmU5
CxEHzC4qIPALQHDhgYyTIjD8xCJk6rI0uR060h2eQCNGExU7Xka000wIQvGiB7RZBQojf4Y6WbAV
MYxrc974c1JgheqTgCsY6ZRbnPyVNZF21S7i1bKD83WD7ELv5Mrp7EuuYDesz5A3cZJp7kpC7TYz
1ZzNhkHhJVgsTNgDlTPdAszl+okSBtkc9TZupCFsxzDdFRbr+0zXaquV0cnL96HthhEhOWDdYlDp
9hmLiV6zcfaiiPngEFPrMQ9tbiFWbC0mdsiPSBDeVBevWZbn/4i4NIuI2Ha6OnYz7Ec7UBheDpq7
nhs3SSeyIcwicOmdfbISr4OPxvG5wdLj0FR9IG7y9WcaPo0W/BAj1MEo6cqQczxdiXDWc8upv3zy
pPhL+/D9ewUwUuZARLtFfHA76Dcpi8ggkAjFQ41foUIW6FFkZbA4zWvcsLuaVhWhELeUwy8oHMKW
Eq+IvhnrCNFrLK4YOtWE1ZxT2sFRXp0S3qgxJ3VEtgr2fCY+J095HVtPk9zUqJiO0tWyTcRlTmDA
uQZPqbpCfKsjPdop2A53L8B4I2dfmwC+djwYiX1zjDliA1vgqNYR/HRUsx+lCl5JorcN6cIqu5bx
QSf2hVxUoOcivQUTeej0+GyAok7d0P+mU5ZprW2iFYYzF6R48dL+rSp/ZsADjlpZQG5KZRkrn6cl
IpS/TF9yFAKvd5uuGI4zlNkVXR+A0j72xiYSI4Egy5Hc7wVgRXXebel9pSBKmN6UkQMQnBkjD/I4
ukVeEIWsNxhVvrlySzyKHwIyZ/F6+dhnoW7ghqLWEd6w27RV3nLUljz5dq3rh0/XSaWO731H+9CJ
B+pe8CM8myRIBbrAIeoDdHrTx0GVbJOSUttqaXlV51ADdROkmb+FTj2sYXlBgJ/r1JnegjIq16M2
579vGmQsgcIK61cT+R9LTA5kCdOS2n9iyUAbUOQD70syE2awycSdBTKtrJv1pDchxyE4qGgOwGu+
74Iz1uVStIv2SZf8c7cQ3oZNAhpHAsEGAMiWjVt8Sdd/3xu55LDUm254pWtO5lnSBUF5zYltqyS8
aFxRP395qujsDomYll0mH+chpHES+atctrW68RF7lVTQW2zjPceCkRJ457z5SChAvLd7P9SuEyWb
H1P3GGIE7wf9c+6HiAGCivdLasBqM+B2r+7X/izEfVhzSFHM5XCQWtXkV9XMw64Z8Y/3J4G4+Y4F
W4DCv+3kI+8TH04FevDCK8NsYeiX3obLiP0QGlwQYr6mBaY3bbuaK54VGQ78TzJR1xFCwL20xQ35
QPqie94t1NL75DRz/iCAK1AkdGOVHPdq5iyxqGMnljDQ2sjClUqx1B6J8PkSM7JtJCZjL3zidF5D
zrATkLpP4csrQmBz7zmNFuE0D62+co6rA5Pn4PpZa/zsyW/aY+0brAZ7IzdVEj3wgX43k8w53WIB
WQm1eRe3uzOId8B1iX15DSsL3Kzajj8g85ZB8nvyI5SX9lIsFb6g6k8o5T9B4E7VG9H4paDLHbRG
NU4okh05T2mxzcWUCDwXSrIjRQTNfCJ2YzdSfhmHOgF3QNdRRGe2PBn4aJ/nmQeQHDVDIaiNMsNp
ueDbJGPAunx2NPv9T3pcyPUnpmEM9hBK+4NEMZXFvGBlnfVfBOTOjknXM1zkG97YyS1hTTFQdeS6
2ivsZfRFucHs7QuJX1kIYtt9r4TkpFPzkDo/XZVNwBfoCwEccm/u8YsN9atnCIGLdmfhuLob4NGP
I6r+rbUd+IWFp+ZtdvMi2lTDXWAHqTfyOnBnAD3X7lFY/yvNEwtruyufTyTvgwEfTvXLSms0DcWr
vAL76XX5TCmpJKgBguppz9lWh32sFmNWC/WXLrG7Amyy/eFt2rksUWIbujtcFI+IAUc8AFBrqkRN
yKfJHuhHBIZazNadPEAYof4GRdZA1vzGiumHlHN+c2X87enT5Ho6Q2WYT6lVlkggG1YwYr8Ykn9n
hn8n+oq6L7mwZm2SBKdXdpUYwZomyiC8UpLsp9YrYh4mzKZgbR3gemO47KlsMlrRDbsDKfa7RQJU
Tx8lRuw0v9i09bi2f1KHgglL6RuCqxOQYztzrXfqqrntwsQLW9QmbdD4X2eVarAngjIGejVfWuIU
F5LpydilumIN5q4FtQhmKtnyehxEyjGB/ZWPlRzjhNHNtWQEqqkf1FZRqeqJitDqd3JypYrY0V6v
cU5Bb/yYUTbWEejMIzQxdKV45Aec2kwYO9lJ3wftN8rR2AuJLSDFJ6Pa0VuPewv7SWuQR42DxPG9
vvn/6x/rV9tGKjW+dUsq3WABGKWOp4Fq5hCPuay0pK0DXJAMV+wl7xYbWkZjUrAWVqFAu6wVEo+f
rkwTVHYpedR+R3AsrVZMgxnCxlBJE3nZdn1W/TDDosiFxIvzk6AHCbScNiIL8FyMSzDvJK7A5m8l
JoFbzNtvRxMw+bho2YOcR8B6NNilE42DgNAKYqHZr3x6z5UCgis6HraDw1dey02dZW9Z93rIHHNX
MXhAyqnH94BLCg6t4Qs551a9VXDrcxqEWPING1RdNfcBESraKb3gSbvDkWJDtEbyuOmJX3OH9hY8
0XYlnAePFtnvqs98Djf8d60u+Sx2do5M5zqOU6jSKfvd+SvPwLBld1UfBv8yzBIvfN+w19TEN64B
XeVjRKw8ac+Q4x6IszRFxl9u7Yef17sJpFi+6kNmeqWEkGrIqxiNHlKTwYS3zOFVdsShnBsEiH63
TJEMu2DAB5M30MrtCNGz32ab3YxT6YWx1Rp8no8vGW6+MNbEIiYKJAvauTFqr+U7jimPJEnRSB9r
HfLjgtPI4rfdTDsTiGoIzPFwkJJd5x8ug7twAg/KyY4GDfrFVU5o5J5yGC5ZIz6vsBMUZxhAh8RH
oLOfnRYVcKwdDMWmeWa0BdRI1aU3PL7rGW9IHSCpA5EqQ/pFp4qignYT1t06CjoFclzyGAoOvSTT
qZFyWDsbkcKONvNV0sftRmORMAg6NFjmNswKWzvT/x4FdOkEWHR81u2dVLWJAkeXBUj9tU3uVxQ7
uwTDttJqVv8cb+IHOxIYqq6HOGQ/t1/1GlrIMuCBHNwwdpP+60Ums3LAl2odYR/ZhU9XMgQsZvP4
PRjv39ADqf1bwKvDqT4oNzFOd2qAxNkgjPZ0JhxbQbMC1GvAv/WCelI/CeSEPkmN244u60+9je3O
+Yb3PALjvQgMkgnzkelfAd+HVnukgGKuCYQBOgSTfF4mQIk18L6W0TWsbL1CdUOQLmJRSFffd/9K
ivzALFAijo73eMtDp4m+UmoEHLJ1wBET+N18RDfrccKO4ZsL2NeUW4SeLYZEnEyeKqvdIagj7NgZ
KWK+N9avUQAbFJqwKXt8E3XawpRwTOHLs35pMWsAYKdomC/12gX6sPc/muUNHVUhYLyYLsOQBovy
UH7Uuh+JrqEysnx2NlWN96QToTh4TDx5wrdPPCzIkuH4Rbu5+V3zQfDIv9nqbYkY1dvreHGxzWup
mjTloNyj+injSvKNI5vxLA8xAQ3Dps2jqKLhX58kBdIgTartFpla8ZK9AprN2B4zvsPMftjph62z
kyNXZFi4KGg4LNKx3jzLi8q85Gt029/pIAtxvx+DRve4nlrqEMsFOGfGFTId+6QT3GQxWG9AdDo9
uL51YL1a+Ng2as3W3TI/2xYBjvuC6CI1ZM2M8KIqLNHmO1vdt42TCIQ/HkSM7pjUYP9pruI09bdZ
4y9+tLcUR1VG9NDX9SeygHTduebv62Vn/Qlj+y90XsTuibkt0xrDj8S2hFxRvzj4WCpRKL5HDwzX
mev29DscWJSio5uEmlsTjI6c9jU8PTqTrQ/FfFGtlIESJ7IUzLlk6P0tG9KRS7cYQp+SPr0JjFhz
bdMh8O/sK+cMqrHhT+V2BTreYYjUd9yCXOAsg1rTGPATAJdma/moCVRTznSVUCM59DxAp588lsdM
xLVXrRLUCnUkvxLCFA53gWQ7JB36R/VCMTrMakRKYcMCECB6tCQmkvoZdJWZ7pbpF5W9iEBcKHHN
hKq0r75BgOH56H6hyM+0RusDorDKj2HcWDZ87PknMfHvvIPqdVbFcpNtzKaH5YDlKQv6dvEcKF+g
w+YsLluvlmMuE6ivRE5e1KPz0mG2hhar/z9mNralIFQrHciLT5woQBeGmCTqadhfrA910VYG3Huz
1j9XuqniNMHXQ2jwuAOiU8kXY/3G+vlsn6stajYfiUB/rEwNx9wNTGHkH/tr6z334YvLZiTvp7Kx
doQFoHZnhYD1XhbWxBF/Pbvo+PNXTFYkgRw1SKQgeUuggWq+qYcfLkq9v7VD+KrcIRo4aM72aol6
GR94NfP2e9RSqmnDATMzpfQG0dbK45KmRRJ7Kq5TJ20PjfuXsEWgSZK/2PjmH/bXELYf/86YfkBD
WVz5mavjDxit0+a01BjjsphlSI7KxxwTz8VGk+Qo/JUxtHyHA3VL2A+nvc98s9/fjRmQsK5dNYkp
1PsH84IxXewJhhSo+z/YdSiREXv1g1KjiEIYZe3d++b6lHT+jhXfewIgl6CnXT9xv7z2JZJzz0DJ
v/xgwcT96sb+CB5N6jXQommeD4oL1UfDef7fYYrW2GRfvl9r4Z+ptafW/5bH5wIgmkSR96yhyhI0
JLreCHbijZei/R8iXYbqNm83QR6Aw4F850WQXuZp/ZRVbUa1skS9WyOM1yGRLZcQ9US0BuSdc1UD
/FcYLYxw06dVocTNlLbxLP/yn57cjWe5enDRSmAtu7y8Hh7LlOo1jO+6mDkNeOfOjohihbCo/pw2
vf8wOyvugiUfF+cNne26WyKAEKkZBVaIcvU4AmkLtydK2krpAv4IACw+MFnQzKwe1I5V4VRRj5Hs
mZoF4thDaGdpO6dCFcFZ2jlEvyx/sZaveDZJW2ePjE9ZYEtB9dJ5uwlPcaovzj9vYlVS79nMmTWj
T5pH40GaZQtT9nxMwpypK/z2/ix5ITUvhuW0DAYrq1WY2ilcLZfbcgN6zvlsmn4qoNyWzMFoHyj6
88b4x8w+/ImcEKKVRUYXUzQcqLiqVxakc1PxWNHS+/iztEe60XUpN3teSrZHT+TOq70zUTxtt1Vm
9b6w+Y++n6q6TJ3d7OGfnwqzHIkIaxN6KFQX2U3yH3PNshWC6tpwp2WwRmFQg8NAUjV2ndiGwGQ6
o1M3HDCu1qkaQU6C9jGBR9319SLeaEsTSZus0zKxaNlxGciCvDS3Y2Pj593VE+79QZKnP87/QfuZ
bjKwUwrwkBhQpzr6kXo6NNLhcn7Ek9owLRLSi7Fi0kTMtt2LSJ6A8yhbCHXaA2ZoaKZiR0cUq/XO
WvLxlkMn1ta5M1bkBQEoMFj9u+Ntta6EuORZmyIC2zgjBwfPP8KcWixSA9AcN2Nmj1l9HRlwYn3M
s1C/zV5KORvgOF5bsZGPatrqL5L+eDJetTJqlvgxbJqkiBYi9moBUhKIUzprrhNnERTqrtwWkTWs
+CL3aLSdewlS3K30/JmMAaFF0nAUlmFJZPsGbCL+FYWC/xf4OPwvnOnP0PF6oyS/y2A74K4mWsOB
FeQ3HPrrnKZnlazvDfKtrg+Dw4qZzx0PFgwzRWvlSzY2rprLme6JZpCyrksS3cEJDe/am/O+TJg/
px9OX9UeTkqStLt8mMKYOky0+hX5yBNmwqVyZsv9sEsZQyttexzDa4zSBfWUss6Psw3NTNuj0uPs
NFk2zMh7TDbqro+ErUW4kAfXyV8rvrQw8+olD9fUmlDaAs32y6jTpUbS1CmNDMKxB2Fe+3jotYw3
0fdxeb/0ymhv2vWPIfDt5/HGWQuG4XF9ZhtsltH41UHIMZLz8hh3wT79qvN2sTGqYsog/lIskfvB
UdIjF99WmwK/AXotZgGKg9JvKm+idySuG0AhSGL596pXCC76jAbFuURWQemt5iC3umuQuWZEY9ML
5Ylx9agHZBufEgH0inrJ7ACMR/Apye6YJ12STmvV9Qso4w+uW6jvOdpfSu7KEriF5HnNyU7X10N7
lo46NbmYN5bbkgEFWrQEZDZzmT5ZYjqAk46M7rhB7RPClO5vHntvcx63LIienIhY17zLfaF5Zz25
M6nCAqq/L4awp7yrRKAmdp+KdibpiUEMBOUt1R+FyzzbJs+H4carlXG+fE50ydiJfM/Wxoh28Ana
jJDv3K8LW3C5IggSA++RjdGDOMqZHSR/R3kihwStu3ZLk/tNU6FJLu5eE7mxAZujBl+p66W7S4fm
QieGm6CIzkOGZolsK4HaKSVnFpkmfxw4Vymo6XN3bhWpQQsByXSx7HFZN+H0xoKDYViOIylTZ/ep
NqYy6fT+nwanlSA/TYg1Zocb0+qfNvXLbOv00hA3gPE9Plfvxeoe70L3atzbXdONkoCuvSWt1dtI
oS7sb/6HuXmSPlqIxTPpuxG0fF4dHU6jrWj5yBropGPEER0BncJnPhP5qIlntYzFClVuNC0vNFzH
TTMOoewU7j6Zqp9/8nRFp12J267YmFl9b/WjMuzqKMOozNIdeMZSbgd/qYiYTNd89/zGfmdj6n4Q
iap34x6rCiL6a+THT35S3u4QwUAgBkXlJ+4DQiSphKPxIvoq2L3wIK97T8qL8NFkILK15mT3lHLJ
eZYGMDJZOJcK3uMsr4WDI9OnGqoXsb89op7AhwsizBGxttOt553KRZoCWb6NK+n+J2V8DX6RXbWa
P8E0eUqMvPk7G/TDm0e0e2vEmlMiQel1j+DtFMD98sXRedk77cgA/RkRv5nIS4dHrGe8/4/nBnsJ
pEbZunNG2cYfE6RO3qtyip2DbgeFvEkqUb1Muu0+kQBPexoUTAQTu44oU4kx4qOcNzN+79u8QkaK
Tcx7bwD65Q4EAlBcXWpxV6Q9t2GhJQ3y2C1WENEuy+oWjkg3NQAxIzu43yZN3ntZPmhwpEUAynL8
RB4APOkUGR3F34cOHwmGzRdUoiQlmhaF70FHnfmzS0u9XhSY+0/4sh1n4nP347kj8SWT7s3jVDwR
hY8o+wg/tw5BIgxsF5ISIzMfq/YAqC6zM5HAH4pQKo8xrYRl6veqgf5LdMhoQ2Ahx9xR25Jelfsz
zUBk9SuaXiTOjKEVD6lj0bAxw4mCEAnJYZcZTgfErUOLLx0hnjQxlLIFW5qggI4Z647nD+HbIXaW
DBxsPiBY2KPSnNIvCKBbi3A6KZNXLIvSfufC4/FnnJJDXdU9+sJwptEbk+YX7jTWiG/ULyv3/znt
BkNxbYRXddvaJNUsZnC0rGcOEasIeG8mAx8zikNCyOp4TfnThGbnZ9M3r46GNyTLqPK5chQUfGuu
qvpR5ArDjvwHKoVHqdqtWctMS4iHRjo017aMffu5rFkOOFR6Dq5WDEQZkGhoMNpAXwePRJ7Quun9
ifzYF7iiuwkrE96vzU9RML7/6BMspmdKLTEanqaBVnc0ve4DpjGr96jbaF7IzuC0sUHMC9XB4apy
nLg71ekmh/urG41s9ssuYmPe1yEVQaQAveDSBZAajrCrpJ7UkIMdKHN8xKhe3NcwF44pHwqgt9tZ
eYc2bkTaI3NPHUWJGOUkWmttjyzhMkMYLXhz/fkG5lSfBTzTBHFPa/m4awYbIH/Jvgsw2o7nA3yC
eoIqb3aQFRbrXR6Q3MPoZUz3a7F9gmRwZhvO4zfhoqHjo1Z4/oXx0sYgYpxP8Q5x64asw7l/cKxh
TDOG6KmYyYSSdRNuLIzHrnJ2duXOdVDV6GAB35jMuM+PB7bw7wPwYQz9vc2h7RlCC61nw0wZokHE
dBViUDaGQku5MP4y1nyaoojJAQDqSlmRj0e5aCu4E7qJqdeEJIPsuI1WQE1kkxpgwHWF9Nur19e3
Tu2cMlaZVejaMibeE3XiEeAHufCq+Ku38eiyWTfUG3vyC8G6+chd6d8WYZdq1tU6ILw70+C+mbf9
UYwuB/+rf6KfthkqoQzh5SvI9F8+GvVQBdYMf+93uEzwKDiFzXqE6avh/RIGJSNAhPdCMw7zLsTv
hqGZLH6ZtFMnQ60js/rLbIdQGJM8B1Ve+ejyq8sC4pv2QALHhQ6i1hOdN5Qafd11peMoF8RYhmr3
9zMBYeON5fQICK5rsIdqTLJS73/JG2/yNc0tWN7Jqchj6mJI/Er1m3yHos6w5Zi3C/CLcDPl8IuH
5Dqzj9qk/b9waUyD97mn1d3/69tfHy/KYjUtfbRb9vxN6DlKC6xj5+kHQkhUyHhcS5wkjbXLj2Ua
VvxmoobGzC7BRtHZqJdwEDbj9RZVssXO591EDZ2eO9+c+wlf9W47fw7F/oM0hcEHFUlk4qAe5KIS
xCgUumtntaIt5Dvsr938p0FSjeC9Ab8Zqy1IKSYpxQT6ej71L+TRa5UqLpUf59IzStuGqlRn0fjM
8P473weA4692rh/u6TC/0Jo/1BmIRiHwvV3dCqfJKLuNFe09rILF5nH5DmfvyavdIqxN1C7hCtWr
VhZQTQBHBPyMlNbq9nfoyzvKIMX57jHtVQT5Pd7Z3Kcr6v7uF0eVXEH+xeQg0BUHQKLOP/hTy68I
+rPOwZgN95OXyEYi351xh7ILBmMM31yhCCt1BeRV92+KBXxi8cz/RrO7OMR9bOfmv4eQNMjF0LHP
UZ4VKnz0OGn6U6nuygTQlQClvcB2+8Tt3t7DRNFiGAAYx645vJYcCV4SbQuf2Ie8FLwdPCP/LUb8
tDlvkAWkVzXItuzI85FxBmBfuWWMgcJjsRyuuiRDz9AfUmNnrOijxfMYVrwiwVcDRktGCy3SC6dt
Xt4Yu14y9HqNQnr1DIu62pb+zClgJpCg1rfX0sLVVyF8TxLm5iiIim7ZqTPA3MlKpHrKzLtDu9+N
HtnxhAHNM8DTbfuK1BcHMwYrYs595wQUAaUQOHBqCKwib7H51gvlJsUjlQQlV7IwB3jUtyQ3dxKD
2JK0tYzWy7A0RFyTxaUvpzNQJllzujg5zLVm08Uj8a3Zedsfc47sIlcHfpiAgXzkGNWlq7MZQ6jG
vYu/doJ6ZZrZkBpUTkbVpCqu/xJ1KY2HO7GFFYvVR2sgEG3DHp6iYGoJ5AB70RiUCkOa71enLOlM
WMjMYzVb5m+EelJZJnNff9XVasWxp/3BC1U/ascvGXL1jXnzisK3kv987kUb3MMsLfa0Z0iCaq+2
jWGj9+5gdRRMel2RXsLraVbYZ31TxB8E0TZATWxLTMj+bsI+hTTCTWhAHW6SB/puAcetjBT/I2IA
ltzi0MiNleor5D6IZmKMCUPeEIRvZerVDwuabNOECSuAREwsuqkHYD8gfFHBkWaFcvckhwJntcps
ur+0n6/0Av7KTH6PzyDjLqBYQLnnyV+ljD0iNEjX8Tm3OCg2X+rdDJInPQK9UInHtMJ8ynYSudox
n7MX+ERHmChzKZFxPLCBrkycuVdV0UnQR7t5XEwykFCNGWARvHM+HAWq1uu5MFyUBYfzcaMKgMlL
dnnkqetgQjekqG3cJWby75bhLnfcJQ2G/53KsqGfpIz8YkopMV9BLyik4nMkcnTYTnHiTX0CYY6v
JWhyZ9peTiv5tqulMkyOOQvoorWotVyJG1WP2+sMWVAg4dEuHeAtx5b6PHIiH/NB6sdzSgBrSOSV
z0p6msLqxY2EvUnICL402j+n+8i8UNOVoSmMR8U01NudxfNIko+3A2J5U8xTZEuyJedfVLY+f2MI
iq96C6q6wX2x/NsUNtc3UMIy7Mj9AfmbJBK0EaEIH23yozY0wbJKTMQeA+PVlLs+pJsoKthNAWdo
cvJv7QcM7cRUYJXUHfMWapqd7QFC9eAI5WVt6swsOvZKeKZJnzEpJU9a2/n1kBClj30FWKUH7Mgc
/lcV7Cbg+rm8bImBm+9QkL/zc/76wo4Xa6o7cmjh8aYojd55pDq+DCmL9LDCow/PAG9oVdijyb+u
Uo5x5t7TmxxiY4x2iH0gFm0PVGpl+y4llSt1JpyQo/95DID+GKsr+k/+P6IRy9aRlkLZtoAb/eaL
4xyxDRkDJz6vn6InWLnBsjh1b0cVgMh/tD48yJ3gptQ1FQZ8ckP3XXJdnjuDs66/CJqjOFVXCZTV
JY4XFplYppW5eaS7FT10gBXDtHd8aDV51JnvMs+YTGhUjMEVUK06TI45lAZM6XA2TLsHF7kiBxTo
e8cFJIxjpAYbY+gPaK7ZQjwN5jdB2gbeI/S3Wh2w0qTG5KNPOT1/PWrj5y9tffyAtc4a3WrmdUvF
/FbTFszQ4YleIOlfG5OBSr4uT+8lWGvJoofZ68/noPIN9pXt7Ga/qNtzymulBYNZgS5BqFf8iSar
HgRQz5XphZFjdoysK/W8/TNdfRqgh8eEzus92lse5rIoB5SS+qpmhmKf+2q1Qax6PjHwu5hj24hF
2ngVzS2O4ickb4QTWg15/P7CmVib5rHaCrtdYZkuSp/rN5D9oUcwhKKgYduA80zNHeAqJGDK0f+b
r0m52gvCXD3d0UatscD8pYp1XLro1ynCzGEdRMRnxeCmyLGNP9n/1XfIGUw/2v7bQoX5oH5A0WnP
LwnZs/mlHWWslM/P+02l6HxQG3Yz2DLljMR/cnKPZha13lWyB0sgl0Cs81FY1V8FPXyRUkXiG/zz
FHvQHgQXYsWPBqloD0d1a27AA8zZS4IKF/w+icKV7fggIKgDybHDatUWU8I2QFGgR40u8U6b+f1d
ncOeZ4WCGcwkJRH/ozukxjPpgOKYf/arcp/07Lwo1C+NQB3fUDfhLDuwbW+B9fhTgQxw3lCKJgjp
+u8a7r2ddD69U+HzlDvbYx3DNdkU6jP+zRrO6PXfx5/FXyq+MyJ0LddQSw3D4aQMYvU8WFI3NAFM
NItuWzvEPXfnDPJyZI8C/TykiWfdEXcQ6s8EwyAO4qEjxO0OlqGL04mqMTYIpye/Q7Oqg9f6Ihjp
WL/VlCBpNUNLkyZYjsSryVjnwOTA6AjH1pfWQkrUcDi58jKxvR0G+tahuLMRgN/Jbk/hrsb9CDfA
57fzXTrfqAlJT9tBANCpUbp/31W6GZCu9WNViUon5gOcqILhjOZIYmxgQNmZbNLUsOKnqf7x8G14
vdmBfNLLXuvQpQdQUKk62hKO9k/aP0u7XgNz2NrwJzFdco1grM+ReyF9qWJRFqhuO1deH+QRXkoP
SlKi58j/9FWyYBkpW2/Tch0FQGHkPhotIWrioA1WGJwd3LLz1PyjOQYMhv+9R5sMjLyD3Aqumt7h
/fed2ZMd4/SbBBj1xsGpi3KSH78XFyrIiCLmGVpczJGYMor4tGbbx+z5oo2CrUGlWC7TKw+KRJ2T
klMK0laivA6jpCDOZ7DIIyUAJi8xRicMm1Ldl0AK3uNqaN2pJm5HMhcr2UAhdRrV2V/cEEkdJ/ZY
MpuX2p8pRFntGe2B8nX88rbWS+Y7SowTfVaZVmfP5qgvoCFraHCrfOyok+A5SH0/jmUbfh4HKie6
HVR4SNQjnMOkVqNs7DwfjmvJJJXDj5N5vs+1ZwPHZ3rrZJ+v7+UICQDXTzpn1ZJZn1SJC14gefRc
yKnAHGLtJ8EYFNZ6QRVjM/MIMIjy0rsUiGHqfQ1C8XykXpmJUzH04YDqdDcGVXSGFhes3taqhik7
C0lGzAMeIfzewBK379+UmL175R9J6oJ2VLumAUTkUdb1Qcpr/wVvpDTRuVZcGRIoVTWEsq+b5mbO
ro++9G5KqC6x89fG+f7/Y4u7F8xQPI+JrgUadzJNGh8uzFEcPjyPHvK1l3eOScaQWLY+MblcjKcz
YExkjVcbI8D+YolRSHwJdsrr1cwV6ZH3LZKCqh/ouXECYRkpd8GIzmGa0UOC70QVHkJ1SpUHtYMF
WJgxPOUbsAh355wOvqhhP6fI+Raq4+K26xncPy30s813jdS3LrnVcGR8pmfmz8xrRyAZiWQNTQvo
0itsjlh1vicpPv4C7sB2SEd6B3qYDeyZKG8ADNkw+VYby0hSLilfjZFq/zVz7tTsjomsgRLH8fKo
1U2Img7sbIEHQWOZB41NQr1JxMzUtIlWu/J56ExL9A4b/rjYvB6BTtZmtyULs6BurCVkcEGflXG+
ghRUPebjPUkqUzNhh9zxvh4N0ltTTk1tCKMYj+vhWIokSbsjKSswNDnF6Z78vJWaaFNdy/en4nId
XRiDc1keBk4+HC94bT9A39LHmduo+wWbgTPSpWK4Hoz99xCeQQPEJfTU5nqWbXnirKL2GnjEHTf4
Q+RDJ0bM4QUov2x1TEvrLUewcI1MesFWupRv8dFhpgkBUljHcV4vWzxRCnv0Uy9Z8j7iVHGpod8z
LSghY0ud17Ei24iu1unfwK6hr6iD/7g8jqzksCymp/zKQxePZe3/HcsD35aYP55fJhbbyqo74NAu
7jMmSN4cnBnMk7nHSi+jD9MFJhhYGszuMgahvBxWvcYVjd6+6VTEw1VlhpqsK302zQRDCddeA3/8
tud4GP9rGif52ngQXM6xNrWN3HxtUkQLyco/rvcg3ElKehhbqWpbab78z5oLM2Z4VasqIP3M5g+y
8+jU/Q85MT4wRQqAYoTsdvIwWADO2T6PrzA8oNR0tJM+DqgrEDbNf5+RWgKPn/GUq69hXIHs2aKH
5cor1oIrO8F8+cv9UWZMVyIpMa6L+nvCpinN9Tp8NpcmYVBdbacxYHOTvil2JvNBgQQFw2GuE+7r
mN0B4326UmBzp5huPVvYPyuDgi7mVb1xsZhFPqWDukJG89EUdEpICuBWyyQZItgfEZB1xxCPZiGz
HdyMIHf8STyvnTEPk/WvCxazqsvi9sfz6QmCSZAekfBG/Bs3VRz+QbSAd/sLkl+uJJsKiuiGCeoq
fhKt1eiQZmG1Uy0g1A+yN0fRZzxV71Z4gI/2ZriFTrsVQ42/TazH59Pu1HLduoIKFcGt8wi/RKM9
sbBnPFnFoXEIfekyPdD+7v+Mlfw4VHCFE0yaiFm8pa7HmPi9HzQ4Zq2jTvnIWEGrRf5LLK2n5ybS
6V9x9OaNSQ0zOV88fbC7JIeMcpfDzk4aMT+M7bwTvV4Em4/KXpUrsaAKXoMqvNqKz10Yg3Yf82vw
77BgtwRhq/YsRi5FsvIYEKhAl1Wpk1ZsLKQhj2XGfU2TR8HoezSmPj0iynviAOR8Xlm4WydRFi6t
EE81d2oO5V1VltDkXRsyU0LQlbDbh3coBrJ4m2JXPgJTuMckS/MtTP6IOHxEzqxeiySekGnM9CdG
1GaezkCLnS3Nwt3SPOXMYLE1wmHy8PRgqcrQzWYuoxq/Jln2rhuFTzHudtI7PCR46+Cg9StGAFlD
ckcDEu6lDSBe33cQrOhEO9/mHTBUpxaHrOfcRzmWE1Q2uGT1XZn5078KyZmMfsA41++pFbOO9g8M
SOVZYSIIH0ZTvS9lNaExwsp1vzmN3iL7NCkgLrbKrwqNwuvJ/qmwCCtocjcthQ/60euxVs9eEUN1
1/X702IrLljZpSjyAcniVOFZxrqktexWfMiz9NbWwK+lkQ74Y60aOxfNWsZMFlJnoAIorW3azMZI
FaYQdIrdCXYeC6ua+DVMVoQvTNXgM1Y99RkCcPlmodfut/hWZkKSpielXIyAF5FyFD8kc32RWIK6
ma0VjNiw6k4uxurSKLDZnBlu4rzMbA8M/V3xGgXBWxaCklhT+UoZrZICCjRqmyjj5glEcCx9G/rs
902HSaoIJag+QA5JPkaZwAejSRWgTd/jET2IJ4fwVw1pHQiwlvJKbpNhRgrR+ezyhofcyU6mXGjU
cZxkEazzOPMXgjvVcmuFSVp1QRas0Is3dIn5Y5NdcsJtM9sRg677Cf3PVWvTiHYiFsgsAWLv1/jz
XDlHeid5ui69+V4FUHiPILhlGXqBQ0RYs7nwjGNOtgAf9Mlow1S+Xb3GYFD7My/cFS/l5BneIMi4
CEvxbFxPuXEsROeZ5+umTyMxCJ1X0k9VkjPCEz+Tg/z84EIxYQE7liajh2xF+eJ844Y3iy+8atxG
kg2CN/sulxJyGTgdZT0dWCybMfjbWTmTBrB8/NzPMDoo70bKAlL+fno7QttLAuMXhDXxddMsEJ2r
fe2LOjxp5ruqm0pRQkBGpcUqGEXszVeqqGUCstklbLwxS5HSC5h0TgBcEZ1zd9qA42/UbUBZVZzf
HmQpaZRSc5aT0CdxqfWjMe+XS0pOFgIwfngriHynhcCLkQ+Lec6ZDApIK94CPjMqJ2zIhe9CUoze
rpxaHl5O3Jc+KUgy1XM7R1wpDl1OMEOPe9GqYdkHabsi8YXfIEQ8F4A04xNUWafx5UlFEM6xbCSl
meq2DLGEKm3buDb8TOQinqRhHwnHGAjqIDZeVYAeQYy5giUu5QUFYDxzU6jw7HISfEjm0dDgdN1J
bKYMBi7vgHojM+Kz0gsYObyIIv8X5SXUrr/S6BWBGCZ3calAW29Q04dk1EqlbLa3H8ZSCVR/8RDL
PIwBqsS3PHSi3JqZUCna3GdTv2XSI5aAGE2p480W0NFzuYifoUbmxewfY7K5lMv3+NqQ2pQh6pc5
CjlAXvDa7FOgaEoBcmD/FTFnzE6p3mOP8G9KAHl4890qPVe5xJtR25ngfMnnVnlZCTXsDoFleFcm
Npb/z0T+ZBde2WYBHlZna33VbnUr/Cn4rlWSZTdmKyemWE3ptJw77hF3akqdUwMXwWaYHKnc/dty
Ksqh32FxOjbx/pM2W1wnEi9JnyXA91VTftINGdlxLRtzClfLz8atT1Veau6iBK7sEh0WzUdJwNyj
SCAS5TaF1mNwxC6/Z1vds3FY7GZhb3E18Y97LWeua8jwRxY/+B+hxCwl/XZLsza9GhHH6P1xTkZ6
U/IBn0maVWU1Fqtc1faoT+jPdMhoAj/H8kf47d08m3kwWvB9BGbVBm2z0ZhO8mCymTaMdq2luHBo
V8r8B+daKS2D1cQ5rm8FcdD2LBNqPJMpFYh/x3ip4o7wsBAanjbDDD3J3R+VBuiM6m9ETwhWep6d
n7irRqaxuaGoOuRgcKDOzpH7zEL0p3mf5gn1rxDtYdTBoIMhE3/kSaf3uZ/I5yHyPiKzwJNpvbUg
8X+v+JeF+GXEwm4gAYpz1zoOxOz4g1CfKIPdHNsijr2ErH2YijcOnCztQxalv61RJlOvFxGBPQlW
nnyOUueB9YaXpAQ0J6qpNBh9GWSWHONhPVT14QYc4TNrtsyhVaWQK1f6LQ+q/MkWfuOWoyiLQWVh
iASjaA6WERYnqsYcmN5wqIlRQtYLpolL7HVchbfmYBV8+pqgea2mEI87cWyRNScbZtB+dgSAtGHy
SqgW6lfzEtHBIZwm6eEFtZU2TPKBO5wPFIMyDrmgd/c5CLivnD4QpI8xw/ohRmVHDbjLCDXJBEoV
lE9FsX9knJlaTzMI30ISDUqM8i43hAJtsVed5ujiMi4R4T8tcEzqo64YHEkZmSVv2BgkRLuFOcTf
iV9FTKbIke3dw0KkOVzd3l7jYcy+K9xIcKJpuW/4h6TxOTpUXGm4onngYVtVkRWvxHQya2e/CmI8
NJTyErNXFDfTpqhc9+dcm+ppeZv+QCT9AbtWGmldOd0cS2ooFZnKCjetTeuDDMhz44iJQRVIpgpI
frbh+J4FpNBCgq8b1CNZ3KhLRk4+Mn8MsPSnm32JQKUbFAwOugMOceUaQ1ZrxJbgRoXUUKO3+fZ/
WRBD/VxLbvyahP27Mdzdnt3FGQlMve9kznQ7qs9QkOQkjjSw0l2/DzbywaNhQAN6Nnc0ejNRUYMO
KH5p9T5WijGvhNKqp1rF9Rq9grm+qRK7pFEQaLbwfPJTMX4M1V0Y39M010FnWTjRyRB1WwXH1Hbe
aPjj0+F8QZ8yTF9WdDeui+FJ8QatR5GJcF2MZaV2y4br6rJkyvU/cqQXcGjPKKhJfb2qG6dhYDQ9
Pk193vY9x8hgQZDPwHv/QKd0Q3PSH8f+AQAiKTbHpzQz8Nk9tHASP9D72vRBUy3Vuyyamqg20iFw
Xe4vvb7ULTIVigNsRUmlJ3f7Jx4W3TRUd+ELR4fbr3Rfde9QOVtKpu6WaLmt4R+va1eXLAk30DOC
piSI/kd8nuA+ujX+Y6Ovy/ddSvFOKyFcZtEDit12arDSyQHFHYrlzWLB+exBX6vg6crRHKvK68L/
gkRr9khNrRJlV+FEiuzlnbaqaGuSeRV16meyaZzT6iwb7/Pq1cRsJD/7b0KBz6nLYPWvkpNtairN
SOQwjZwsZDqWS7gmmsbvIwU1E7v6mPFYOFDqrkU0Vxnzq27b6+VhlcSwGcPMmfKIGcl1I1+++r/C
jny5DoynenB2fWMo9q2YTlVv82z1KiOiomJQ93FkGUI4Dt8+GvHVy2fBiie5mRi3yhghkBk8CtNS
/xMcWBXmX/6Sx9U43ldo6bE+quZVu8gTBzk++CoGKcbzJiCBZ2fKZ+l6ZzWlcbw0uP1hIYwkjNTq
iX3L4pGH6PWo8AHTQH69i+XvEByz8u3FKRKzMg534lnPkZanLauiysefGXS0xmMwJpzvP8682fR/
G7VLkCF1CqjlysCu6qwAxGJZOxunqL+0PJkpPawvTaRMzkdBq56w11Cp287BJ8ReXrkv8LVRDOgt
mL2pKmkWpGEZNdIwlocZ9y5Pe5xXwCjBGuDiJFYdVMJ5lFZgiJJ/lPpjCK6zreMzHdTDmES+zYqT
1rg1zmk64oOR2ibsx3j5mYA8kdi0p6hFhjO35sznA37VAOgrUPekaYDF/1lzyPBQijT5HXHjIfPP
76sEoA40FPAc0IE/GGRXOh2FyB55gTSCybkDxsaQpLkaaViZkWN8h4O5di8WUIjeNM/HqnrocdFr
q/prs2hmMPECsVi/qwkRxdIrH6WSHuzgH9nOYimIrMC5nM/daEN/B9v/xowP1S0YvdOqhZsHi9G9
A2atRCau0Dk+HRIAfq+etGQ4YSJmSKtwvNik8AqIzgLzzRp/FlpDeH6+Gr6TDUwIsht+E9lc7Ol2
l0pEAH0Oj6jtWmzwfiVmM2Oz0MM5hH0HTm+z1RuvN9lcpTdIBwAPVVM7+5TfCx3wK7wsDkGx2WtZ
Po6mmy37WWR+ENEZ9NJnIBLUTcWQvbrFiorvHZ57So1kCpF/F+PflOW62GOZPl5pKi+Js+r1HbGP
nXt+UHW+A4/Js12tGBb5Jhy8nAAw/qBaz9P7sy4ZXqWzwPbXFOCmJVu1WsTqE0ekBAJ6zxf9M48y
7gCUVq1N1pb3hpbW09jGaZPlE/mP0+pMiTw5zIUCsPC9VM1BxW2GUI9FnS1+GfxJYWL7ylSIxCrk
otinnfwd2VKcRfoJcGp7DfNWhiZzLBgszDYOKfsEVkBAF8OJVX9dM2swfp8jr/7Q+MmkzMnHEwOp
mEbro9y+/h7aytob2lm2FLgWt4ig0NCtkkXRk8Q0e7veFOeFAhnoVoL06v11ppBun7O5HlB6LT6q
u1wvqTO2Z80cpHCts87a9JfPYVyXRgPM6iiFaMKj5Rd58DiNu8FPtbX3oyvnLHSH+7WGPymD0CSX
AdF3qOic5Jhcnhqa9d7OChiW9+vdMThnBBbQ4yB2B3Xs14sc9/eVL6I69GTLJD7fFG0vboUG/Fs7
aYdjb6No7hpowPDpDR/Hu7QMRxUaRixIGn6uMg7l5At1BJselgcz9MDctL+NMHP0/hHfYRhk+XtW
4elm/ZIRXuufn3y0bw2o/RreezkGMzKhQ92TERjDuVI/hlCVUeILpRCzv/O+WQvclN/pN6DlxsGa
ymDKB+4FbWHiBbxDSiNE3w+kJ//TyFKUGZ/YPFYFb/fuFdbbiOy9M1uZlb381qmoaJfk8C3psjWe
Aujnr2RLosb4R7J9f7HQMX93V3qEdIwNVmqvkS8vLpbOxzvBYrmWSghoTEHPM0SXIMfOP4yBuPan
L39EFG7tZwoH8wkuTBC2olOeDYYn24RnbyKFL2vtaGoBXH1UOn2eyZa1npE9IPxpCeRezwm2Vybz
6zoPtbuRdXM6orE+cQ0Zhg3JlFp8iYg9VbzrXWWqa1ggbQripFi/ZUwqWQXZkS77XN2A1nDQFhTn
39mZ++CE9JY9iVTgIS/8FKweybGBXc0vD6NVUIu13DmEazaBlbZSxROutDFnps9s5oeY1F4aba5b
xH3IBak3kMbB2N6gC42UCC5kMDlzD5tozo+OsZQJcpzRv/KOajOF1yyeLv17cBU2iIMC4SPlh6Gw
NmHhUxmkv//BG2RnI2LhnDJvAcDywiBTGROMkuY7qR4k2O4esFy7l5ZNNoQbtUXKLXXc89QzOD1D
WmsncxVO9ecWbtmnmLGW8GB7mXDHzmStj8fdPJJ9i2OdzthhiIzesgMNiPKK4yDdNBU05Ls/oktt
nRZ/qxK9yCywEE20+vndByipxkq7Dg3aUGlcDyoT/2NLeP48uvTNawG9JIhTmZaxMiEP1HVIMNAR
NmktSTyIfQd5xuDCCDxuOSJmlPFZ/QfjPElSdQWB2cNDdak/XyfEgfcvtIIifWrMpYuoDROKUtWQ
SLlk0rXTA1k2902s3EMO/n4K1P2cHocXBm9kMd424Iz2dEwZw37m5pvpNR7CD3paMDbYblW+hy24
Hk0F0fIKh/jA4eOCU+79Eswks6Lt4OXdP5QqPFTIXit/AzMA3pZ7RfTkx5q9aIHM0LEcLDsh42zV
wnV968d6ISqsS6R33SyU5h7HDBri4PWUCPr7G0kN2mOyi8h37CkeajC+HqBxzT5W498/S/PwJU7x
CToH7PSN9X8ZnUlfMA8ODw8nKWuxnRWa0KnMTEcY8hbnz6JnD1qG+HaDnDhALi1gat0oXoMWTFmi
XuaJ5tihmBxkhWQVJDiNi2jPHpjJvxSNsBXmKtM1NCS2PmJiyNGaxwZ8bjDveX8j4/8uPaKiVSAV
G1emn3I3xlLDFeCL23+nfa3Q5F+X8F917dOK9Xy3KCcDE9IcFkIUCnhEN2oWkjHzfby4J1nhCaIF
O1ANpFJ3JU4Y1/IEwAQ1Q73caQ8HNnQOpXrn2G5PnuLhUfZpZlyKA7t0dN3yoEahA89URWSMJho+
HRtGEcKCHa+cXQV+msRuowmlu40y0DdfHJkrpXiFYHw8IP3Dp0Jb+XgbTD3u30cClgh9JsKAiJPa
AP4jHGNeTpmaX5URiIiOIqGlY9mjSdLyMreRmqCAIAfMMjUZh0m9So6d07k24EE4uobplVuAPJc+
3FzUDJ/PN0fH3ZCvwSoa3lZtTHV2Vv4z2v91v3o+zKKCS2yLs465qR4tMmUvXa7naA2DbGOGJWMi
g0R995BqbtIxpcZtMCOP1EpARBQCtTQidBFOwb+hRokfv7JcCkyJtzkLEegR1V7Y6qcGD5ce1qlG
zLfLDNwz0X46TVsdk9rEfE55P8q5RWMbOIJEFUWRRSI/FQuRCAuCyhhCOcUPDozLPg+nhI0m2jLB
7E9KWivFcfyTw4khUyp7bhVxs6MsQNfK5RW/gIVHNUVV1s8PQn/QGoYcxRwHvFwWgge7sHkNqnQt
v6EfUfsIcmttwwlkPcodgHU4TQKymSlmnr+2gijahH1jSRctL1fhOt6f//s7mJHf1V+Os6xHlQGN
A8oW4AI3h91yxCvrapgFQRrNQR7BwAvni6gFsh0fZZ5AHmnnhO3jB7QJrVxNDF9dehwwjJazuuFa
094tA8DsZ2UK0TnhJkED+0VROSCB3Hf3tdBLMs9WQibhIlayoMaW26Cjp0uN8y+vUdJD7DyMjnW5
d0GlqRvPi7WUr6t2RVrQOgjryfKf4vMbCnwKGBgLnUezf319+xIJXVqCFzbcWxGQUUkFiVTGwmjG
ENyb9QGnvNlti/ClfVDx+cECaVRGRbG9lHO2Qbch4i/kNHJkCb6LXCbE9IJezgXSZyNduP+FR5kD
DL/55aG6LAPCjkcc3LRz5QzBp8koKchFyey69l1jk4dZJaRMo6AKmZlnjqokhazU4XgpACvnoopK
/7c/XMQMMExWa1uDRQlNYc+cxvhhty76QmFmAS4xx5h+qgFkCyY/J+5JunJMNL/QlivlahIF+3by
KK4O/mYA8ZT0drKgB40G3gEFi1jUf6ZnK8RqKiuZscKGJWoRQY/9EtIIfXtKEQ1BBcL4DJ7Qa9fb
3tV4Cgly7vXihmVU+61lF3pq+C/8qfa10YfZ8ZF5Y2HKwufw5/ASKin677FBOc7TAXR00XvU4Wjq
O/fgzQf3xb/pe3SHJaGwKM8d4NotdGM4KagwhhWWF7V9z3CWwYzKlPLqfALJwV9KxZhwcayV/ubM
tEqlA7kjS+zyx6p7e6/m1/GPzIfkFN29SCjxp7MIJTzdmbUjNOY4ZovBOGMs96pQ0i6qryCvMD84
Dg63bctcmfi0eDxNetyKEBJkhEBTAY0hfgDepWT8ZKtKI9T4Q8EWWMG24/OO1MPYPRMMwXzyK1Wq
qJj/DPTjzLsPJBoBq0KOjaRIUQl3uMnrBWI15Iqbv+zz3JkkpdFWRnDDhq4z7/HkTYcH7Crhwe2D
qW13Rrz2ezvn/9DESmJsLggwlYEUqrxzTZvaZHfxVNIo1qZLvUuCT6t29BxYJ1wb7Zwm+4NuPrMg
xKtzcTIwJ5HgjNO3yaaXM4dyYaqIu7Gp3IuNAa4GmDc+VR0eDfwtIMgtVDuCfaa2meheq/BSoiyH
VsV8rOlNs3Tf1o6+lZh6JfnTeoIrM10S+l0WBp/0JUmoscO779Td1T1NGN/nmE8s9sd18JfZRBeu
2itC3hQR6Nxc3PdQvRf3eNJAUA3EXMxzFURrRpK9Dp/JPKMkj7dwi4S9+LKVHGS07pF4RiFCMAYH
aaSJINe4s4ER9d0HVmjMU7xWwLhUsqP00g51jmXnV6nIOerEGbVJdUrO/2WuDFjbp3PlYIvoa5ZK
AY1M3w7w517jlCqu0vscmdiDOPpU5CtogQYxL04R1p3kUjKfKAc4dTrwKu8GYGAIztnHK/jdIEGp
e/j/cO1ILy/tWWygGC6Ffmq0wz6UuzVg6ZKHibQtHnwVIsBHj+uxRMk638gLU/r6wRN1IZlH13P3
tzli7sreHsPWFIcXwiTM98J6ilTotdTNzR3ytEALknIEBYUllk8Gh7bDK8FBAXmLrdlvEL2RCa3x
swstplp3uwKd7dIGsQ9bVfUWR2aSnVD78k/KaNuiJ04OtAtrCb7pqeRxx0kL2bYJOa6+OONS1eWu
J7SPFY5fguEmWqBfi1MEZ1d+vNUKd3dX7mC5kgmQirUKVAN0litzOtGVW53lAIxnUyxoiEL0zxtF
cX29osEyG3NVFRV+8g8CnL9mgW/Q38RSzMdzzshQFsi8X8AH8emI/GtFWZKSeeJfkI7gM/O4M4Z3
+jDX7P8+hDXz0Kfd+wpoAMcEukA9L+UAkR7aZ+11eQduxHNS/6yU9TJRmlyONbyzhcj9iCPCa9qW
uWQHiHXRBNobmb6LCMHLVpfh/9uxnf2Khs5Z5xNcC8G3jP8QPNookhfPS90/HP/3XFxZzGZmd6U0
tR3beOl05Q2RPbPdlU/V+CEmNNCb+oEjqlifuEw6bvL4d0VfdfMZ6n3uej4BDtTiMkrB8owC33Vw
DC2+rHQJ6eNIKEfPQYiYKJ05ytcbwxHQvFUPbEOrcSQLDDKqzzcHDgS/tL7F7yCNQUeRYTBSAYah
gd6i1jHncTk1r60ESet4jVLQx5LmrOZQNjrKGwaKWpvAlho1lPDCeS/G01EMS/4QXpmq0egzVFE1
FddxpL2WfMjkBuhrP7UhK3S07+wqZCRiNV1Sqxi30Z6uutnzQkKZhoBz54EIuvA7n7PYx6EFYQNM
0T4nsw+n4eyaMs8HZQ+N2OIooYt/myzHCRmQJ2GZEqe/sW3cUt1Xu80TNilPKGkap6uzGxe9gPw0
VKQRJ/0ayyduTQb92Qufw0I17jvyC6yEPaPe0JpSDjPGLrU4hZwgqsZPlsz2ccDd1EtPlAzIs82L
dcxW5K89H7aL9wyMMm565dd2C/qIULUtC46fFOZJdXPXhDAalEqKTNHShVBCDSpGQl59VBIOECzU
Cd5ZnPu7J7efSxsDvaMp2oaROL8FEg+iSrjADKwzqHFLhMPfMs5O037/Obp2j4gU2TEiB33U62YG
iuiKOwYM00BGICVALySzzVOwGXvtSzwXyhl/NUQPcrLoeM5QKEFcORsYI/cgmsyhxN1b9hmjTf3a
P6K6WDsdYK6zA2j2ke2b8P2VvscHjiKWyV0kVkgSLO4G748zgdHKRYu7wzLp4d3BKpP9DcIen9Ai
UVvN4Vg1ZVyseOjvB8Z8j6Bsg1Um2zVUav9g4OICQyDh+GIvPXSXTv2CR2bWvV13/MDZFbVOhpsh
9mHjgorfbyP9imXQT+kewKrXiTNpJJeok9G46uZKrWlcQX0NVY5JM1JHOS0K46qEaoTv8u7qmPYr
AaZ0ldoSVlwix45iVBqUWOblz4L2kDn96MfkhcMOyGSp6bOVTKp3fCXrqWoODYyVwcw2Ds+irOnT
9DQH/pe/DsICVtw6ROe3dD1VobjxX6tsZZByovfPhBscxub4EH6TkyBsIPYwqz5qVrJj+++iDZCs
V1E9uqpvQ7T0/nik3OcUfs1Sxg7AfYCOnUz9ZdcThJyxA9Vkth1MBNObur2WbozqjW711g4hJhx+
roX2sBA0Gb35CaST1QiuGwp/CzeU1bwTlW0CpBuwuzmj+XPzxbyZqOAY1jiEbPbiJqfxjd4qxES3
Pj+TNEQGOZjcptkyTHCeVmzp/GU7KA0k+8nMsV7mNrONLtWDo2grYcEG9YTL+u+m/Pkr0WOA4eom
eOPaXHaETwcQbDhK33nVcej5byzxMERpfiraQudX5cR5M9wIxDXzKAxCmwAehnS10jMWnK32qyDq
lJHboympZM0x9wumJ9xhpUB1as8dUMwHncx9vnfvFQLL74PgqMhaYzWjTSU4oUZlIs7IXY7uLbwA
H8WSRB3q0W4JJ/xvjm1gnILmyf0pMlRaXdENImUTzyhfTOGUn+qrnMb/06zTE1TxrqVrM3S+AjNq
qYcCsX939TQ22wff7aKqNiSFaNDg8xtCjUYakCaHVJo/KCq7FUDZ6QnkWGi+ob8cwd/6v4AoMLCN
YvcIYKpHO4LogHk0B2R5PFWkeUvyG70ugKA4Tb8T24IW0sn9VFMVs4zxOgkq7wuyyRZEZL05c8zh
W9jIDq6kwe1Ercvj8lnx6RWrBiV2ULVEHVIP5WvZbzvlsCWH72GJ+SKFdtA/GjnBLXBCyit/G2d8
lNY203L9H3hhZJasAVQt2kQ6qutAztuRuyCT2YCw9v/ZbaF5KSs0nXVmdiIZhCKsku+OlJMHZVFu
7kSss/hsYq1uRkdePsrnwwvZzMmpknD521KIgPxc6B0SlGGlrTKX6Al3AcrmhdoRtfrxfuprFpf0
qQyw/+eiBW0AfHHsi4MUfL/AsnLAzNPqaPbj9eyNe8hON5as+uNw9Zu7BUhCo0IbqTs/B0G4cCBM
FDc4Qy0pl/feviaGqsowOgAe6Oj5q3FyvXec+fbJW8MD+EuJuYcGEtazTzGPWc7/lFEl4F/HHbT6
/PplLsyart0Xi5AYSANxDFl81aLpQFJsp4rCJU9StgrudkvXAUfu25wId1JwhC7X+DEMthw7gdf6
f1kOnP72zPeVrUcpB1E5dPJAeqoFHkrzDC5EuI/iN/OU72qULo88zELdkdMpIYpuPu2t3bps7AJJ
FDMg+kDSvY3pXzqGCGQYTYQwdkZw4NEkvNYVfWoh1yH1AxUMo8BXVK/EPGd2hAwGju9WmGERlbVm
QsXeSs4wvS9vwTbRBUWWNJdoMv0IthN0pjmcI5t1H1+Kz5G+yMr910tCK5g/3lu2a4watqfUcIlm
lX8CmYN5mnuTy9NfXOxePBG7sudlcN8kXiVosYOr16hfuJ0ZrfxgqwmdNV5pQCNe5S36HGb/AMN4
Xj5nPfQPJ7Bp2FhYL5geQJnc4dKPoVYTBUMh+nf6g3uhuGHJlOFNFr01ox/UnJdXtqVtMO6I2IR9
50ufe6rvoevzX9PZnUFOQhKd9YFGyFhbwutxRIT2Io1xLgmBmoPBxq4MKJBjcmOygzz68Gu06xNQ
UuqDOniK99ELlPNy+mdLefRsx9np6GDZ6R8mpbL0EWX+N4fnW5+jQD+UBZYoO2c8DAjdaKaRjcJl
oSniaOSLHIyqwLVnLam+90Bk2Qx2IaQ4g/SrxDsxrr1gRcJiugAm0O00v8X+aiN3cIf7ccLcjTI/
ZOSnietGPnmfOL9JKHZ4K7MWi05qEmp3HfxLAEIItSMvCmQDRtGxiz1F+s5s4ADo9JLW4a3gmJAQ
lMFnSYLVBTPpS2cdHyBykcO1ljQ5O0UVN0QQKHt2V3NvKVCNWXyqkJESvIxuTp5Kog7Zhx/3UdCi
yj8qpjWurN+m1Fkcv4eSUYspkm8CoSlyJq6vFMmQ4hYKVmjIHCWw5XdxP5xh9MT6Pym8Y3wV+zXI
vvleqJBIGDQP4hjs771A1DSs8/BwVgJGYRBLU7X4TPh6D5CwrqdTctMGlTBSqNZ/Dq9dFvEKrqSn
WPCW0++86iepl/0JFhYiFAzB2G0ITIkrE7exjnN1+hKAOiFsm4RnrW6oySZ0u9JOL8XKG1E4oJUS
Opy25rDCxbSTR+GPyfgTZOy7UxXRbrLAng7r/8bdg1IukIwHuO5maf9fpRwvwqSAQ2C2pa9mbOBj
Msy5LJdSr+7ntU1udh1Yd9ckj3Maq3m9eHSALqTnUpBaEqxWhm3bfiy659Qo46gUKU/FOhh4Pi9G
owU8uOhw3TfaJoEGH9tmjlrzabEzY+w0eVI3qRqmuOPVOJILPNobGC9jhclnC0+vCrAFnf8meDCv
4LcsIXg5VTAkthVO+HHpm1viLyPtd9U0WODCpp+vdeUYWnWpUIvloFYwYBZz8+b1au19XqhK9w1m
KWnYGdlnuKppCamXGsU8TXLEyC4myMwoydjOtks5Wbnqnqtq6ysvrR3jp+ciK7xJNWE08v4Pe4zR
C7R2hZWhODk47ovigjy3pxNGhExSSoIBFbyGk/Vi7n9hOaZUrpm+uUHBrAvxVIiwjzOdnax1W/73
HzwJjv3yHbLVJKyNAMTuWDkoZaNUh5w3j54X1x4Gdrcv4BeLwU8RENfjuNdjgZ3DbbnCJ4Kp5JH0
Z0tEeWlMoOf11VL46uZewx5aqIoC6/01LN26tdLvgsVO0fdf1GQjAOlvfF3/VC8iAt8EyGzPTb5E
LBhvcxmJbuEFevZZ63lShgaMd12Vy2QSgKnkNxYVNmb0JYBrvMRN20PbEvk3x+5WxbZpJ7E5yNSN
4WYMap3Sk54Hp1GsfoE1PU5cJoOXLwaMhbvwO4zs3mqcPEMVGqcRQDcbV+kctWQ4ZtWii2sLPrK7
IRHl2RLnpG9DtKkgLf+BF/MI79/zFqSaenUnOQWq4zzBIBQIALzgS6yE02+IaCeucZB2WO2QEHkc
QgRo1zlopUivs1kWRaFAyE0nW56ZHx9TkCg4JNQsSk9gUheOaaGiODNvi8klPRQN4rnJHKKvCvYZ
ns3+0yB968DUa0inuOvbzGSpCgyg8ew9AXwFsEtaFyjZdXy7OtdxqJPOywD6jaM43wCnpf/lySdK
nGit08l/DRLBlkRCjgmy90sgb8Qwocnw8Ipr7DhejZHXoyRWPDiE+ltbmGRRBetPTWXgCGVNAb3j
KT6lRTh5nM8r0Jgjdvj44KHltqNnYkD8vPvcwJXyHFM5wsm1zkzr8EZ8RTsu/wmUN+1ismCbG1n9
lOJjgYjRKXpjhex+v7+AesPX9fA5z8V+BdkIykYemCuoIkyf5CHKNCpVk6oFaOqs9Iq3aun4YGum
GGaZtgWOUjv5UNScmj8Q0g/LKrzIDKCgag7M07+BDhNS/NY9vNuSFk+Jf0H7ZNVS3bYhtT557epi
dP+7foJknxzN3wsGGSdWms//KbkP8B8A1pc3jWS3Lt1Vvspd3u5MzUK1I131GsftKc3z9lxUyZNY
/Db01Wp5v6577v5CTftRZVsTxCeJ5bZXNmbUXOMbKlsl9CnI7RlEzkZbwCctfynbkHtay9PJExE6
A58l4t77+3csybNsOPWe7NKxD95AZ43C4vPkWhGeVoQIhrOXEy/kCp63WDPa54agA/Z6NABj95Gg
nWvz99YrR8IwRy3jA/kwpTRCdkrgWroaVyECalcugKGo+tKhxLusKcALAugDOAjJdMxJmS54sfNN
nMOm8RliQGBpce792vAtMcoMoWwtX+IMchvoXyhAk9kFkx+c/ny9KoBkCnqFDFLfog/8476wErW2
3qoYddv+VT6w36hiRKDs6X3D5Na6OlZ0SRTytTf/qfpvovE09qmXJnJbA8M5KV709351iQuEPu4b
T5pfjm4Exi/nq+Nr0N31GoVEH9ndppwgjvzZHC8WA4ZvF2pyTvl4h6jJbjdIVFr+BLYKxc7gX6jy
4DiZIQqqUt4fJ+iUjRHKcUmIcChMIwfIlwmajND6KxsY/aXyZZLZParqPJA2Wtr2ucquxzSS2Tc8
iGcw6JFWrVgG6MOs38Neo37aiHNemt5N2fNZGqIay4TwwAc1/ry2bKWkxSDz+pi6FI/UArRO65nC
pIU3VJ2Qa3BogBjGi5avmwuSpieYjQS4JSAEHnWDWr6zP0C5DuIBkzAlF2b4gRxiX4CLBhlnXmJK
AxCM1clhWSd8L5p4V0hbEZFA0gdJ34hsdoAEX/pZn7o95lU9oKzzVIU9AsFrAK0xKO3L0lxYYm7t
4Y6I+9fFyx8EauQutzkjFUGR/4Q2IrqU7LobLSujndXnljrcxXKnoxYm3TTdxKnd8yv7zgI77S78
tWoOroi4tBxGs4cikKTpJZs9cdZj5SC4S5O8TaeR7FYEDFad7dQCP/jcc/Dg+FMLld8Klzv8ECk0
ejfPSej7kOGn0Ck4BMeXknCLb2y318eEOp++7SxYvQgG8Ssr9k59IoCjWRHVMRGRn0VghuwfMg8g
CogPmHScWZivqUcKbJShW/4Ll7/fsEHw324KJ9xRhctKEATKGlUwiDWPSH/BTggt3PJLkcUzsL7x
olo5dg/m4Oo6LXzBb5pIeUWaeSdVTlSd4klNeGSXihNabLQ5236Yyf1Fb0L7FVvlKIDig3eteP5P
P6RoKfW+Z/G6/dl8wa03ySQwdJOOJczVp+EAYNIzwO2Ch/dzo9f8NmPvygt7IuRNffW/p/uM+oro
ot4Dq6nCTLvT+LehFC0y9IGMCzqQiSrWRgeASPtLii5EU0ZVT1JS5TLw/Bo+V1WJ0AJfYnN2ao9E
qFYz6pHvkAveYYcdbFbsD1xg7YMpsoky8oYzeGGq2G+cWYlLq0VW8gY928FrN8Po9Lm4t0ETV3LG
/Hj6P/f1Ep7yrIlholR8zcXCx+jj2SbZg3sdhGOIwnCmYZHVlG2RI0EykQ6pgI4KuefLkioLtwn/
PVcZa3awuzlcp1Pu3VBvdRo2k6qFz8Yo2WVmnSEH3AyMQ5BL9ep+l0hafSBP5slNzwVxxY1Hova/
GSDw1JeYZMEtG5G8chfutQP7qbZ1x8RPMOP99jZG1JAMtodqqW03u1szfebJRqtokb6d29GtdZTD
SaLRC7NyE/BbhbERp/qa4HF21DJ2TWp+wxOLHOYDDBx32WTH1/d7MJXKgd5cKrdJSU21GD0YfNk7
kzwddvEY8nlXXQCLCzofnjqZeTVCSJO56BtikURqR/wXoHSu7DoKEBDnm2K4BhCCJL/xgoN1KEoe
oUdijV6XcdHMaQGBNfB49TcjZVz8EKS3NXX50QpFfw+GDym5jr3NF1ijzQicPWpYDJCjZK2LXbUM
BhsdDxBM6D2LK+bplb5UGX7Yfx/Riy+L5/pC7Cj0q6sBHwiANvmSHEnKQQHOwv+cR2eELnjO6ac0
HFj66NgVmHEUncarR6nKdybmVyNH2mXSmb3yXLGcMI7w4lSOzrPFIiIeoqStbkGVsH+QUu9HHZoD
NuCitGI4pQUj8M9wuW5zsIIIy4Z+yaNby8F0lIxRSZGNGCWQ9kTQN07XAduOWTypQNAQauq9onmD
STygoQU2RxYaDnjwDzBMFngVYashdU/IfLgoamA9Grkpzv1OMfoZJWlPkuHswiVfds7KW820Jt9A
jS6HYVaZjHcFW162PEi4tsTyu0GHPG4cN2A/pPaWLC1U+bfZcYdJNiU76522dfb9tSatKxInZvpq
SEQ0k3mZP1YXgGpiKvAxjTjifpATLMnQMSMMwJ3/xXuS1+VrcQ59wwRyaqiWvuXwUyzFXeAMkgHJ
P5nOgcMRT1i1tjBm7YcTKhypVNKRCcupxeqpGGjbZZnYKgbG8RE/wypyH/m0GHnHlgR25XjcipOi
OHf2RCu/ERTH4mrBd8CPx+DHmxalr0976nxm+e2NFyp0wRNqn8EMDNMQtdVs9JD9BwfBxuGYJJPO
wKfhFa7u1uClUMBpNXNsf9Yyoz1AwVAEpM8CoFJuzF6X67vdQasnKs9z3QMpT+vZmREVhRIcFlXf
8dJVOV5T2S526yap0GA4nabVzB1GihpgaBJmb8Qt/PnNIZ9Ew8xD8KTzlx44bv/ItscfvRH8IyGF
IxQ0r7YGfNzRsrAxyYmZZ5xxq+4ey4G0c77UNb+Vp/4SCcn7wBaw2f1x9rmtNyl2bFkLuZZhiSsr
dM9sGvIZxBrdHJ1NZGIxQ1OaVQnompukZZj3UaEI1KoqXnvBwCWBzhDaIR+y9fZQuzctS/ptI01+
5XPlsbmKm8hrdWDvyEEFwN7SS+prPvlTzXedFEhp9ite1gwGnEHy8VKDVVu7Ni6TQvz2b5CLmMKL
2cnq/2WFWiy4TmDu1l/O/d0VfLn1i9wiDMhcnnA60yGWlxdRuC/phRM8Ba+Su6ndftWZbb4JOB3b
Ny90/oxayVQGfBRi0T6mc8DnhNcgHQV/ceDhYKyEN/I1IKPMoqV0jHYPXyKEIrPqdjWLL2kUvWG5
3wCOOL4F0mp+WBwUiFjHtaVh1j7wTZ0zP6txEGdTJjvZhfhBJ5Wb4VIfb1Dc1cOZXhmH5JprJ+Ym
qFeM8lvjmOSLitdWBoKnTet91GSd0h1J8A2wJqLHDRbsAb6GtM9Q3ORoxUFY5s01XJcayjhdglGT
c03ZzgwJ2ecO0TDAd2Ua2rwjxcyo6QMz05uqEh6LhscObam+W24zV3IbOjMiNiI0MGDbJ5SG08fT
7GVcdDGFe97+W2wG1TWYTvWFXbwwN1P74FpQccYOnHA3f3KumELJWJ73K/o1Dn/pIoyTXIInGVp6
aSW0t2cI2XyyoTz3v4xPkYdknCycZbPXG+BPuZF+iyRsDNjc2zmSFxhgf/N79bYI+XbmG0WPXCq0
1ywSde0oMzBWtYEUeshAkmzpN6rn/aYexrZeWxWt3C9lYiewnF1R9c3EYux/hZfHWeIVXS5p/fVy
P3QwPCuAHk4RYhDP/XmRyJADP7lyNKsDTF0/mDyL50oKNXqkXsDFfFvEb9qBoD3cMj6uf1ueYWnW
yOAi976weW0mIsMABY9Kndo6j10OGVFkjYBFLN/vLcGiyVvHaoQBkpQXTGQ8lCiqJB/bOtHc1RRo
FOWnxNfNDIMJtacrWgum9uTHJpmnpjLJRzzNkUdLpmOSqk0VcfBSahuzBD8yseaQQupbl6/PVx0l
FEa4dnB0T3jgWUmQ+1M05HPdrnfo3MRCaIJ75nTas2q+Uu9XFOLZvLY0milqBSudbA9fM0bBKr40
PmCrfw9ckE/c9Qix6syKPPbHL/NYSCeFYTenvL0/jRBcTwxuM+KzylqBrvidQQ8+RqN9aMVhmmN4
vhe3ni+i4oI//ROt+2JhxV1MPXsZN4xoiEWHh5drSrV3arCXFAVLBEY6T2QBEKjNQ64XcW2kx96I
fhOp5S0zUtM2w9qWa5Ie+9gsrnrC6ciih0fXee2GC0IOku3/9RIaetB7cVmsxTJ/oBF4ZbqYPeQR
MyvExQ9c3lE5yrYvf96V9XdH0nHnYqX+ls2MVDkmwbNnaZ/aRhpxxJ1JvHyey7LPpuyv7gddEpgv
7pI88jGM7hXAKIXRdTrGpL6GhrNF9axi7yar8ePgLNnSnOeBY+HsXvaxLJ4py5TdeUjssqA+TlDM
XQxL7R/5KyuVB6ALERwBMgJIZ2ArBwlTEkKXbOskn/xOt+HIPNJotJup8QHlSmgbTZ8C5IkC6Yk+
aM5TFhO5kWDQmccfrcCWkzLTkJCtVRg5Eb+GrbEkzwH3HtSKA3w0U2ecyM1vLjLsMQ9lVh5KE+37
A93IClJDSJYivKPAJm+/yNWSWq41Mix1CS5Jgls+VVRAQ7ZkU2G9k72QfCXksWQMYlzoSVy8nDUT
nOD0rUeXXmK0KRu5vm5I5OQO4wYUW0DJ/V0B9MGoEK3SlIO2RAnJTV51LAagd0v/xg1a5g1BbrqT
PUVMvxgDCr3+eL3qLT74476EoJpJ8Eg285pdgxbRery6JNSrigiOA94BqQDquNib7be7tz5tuY0k
+Nv7VKNnRlzNiwezXVJ5BNe3xz4HWUPQudnh7cKPapzRvXX6w9rFBrGwXakXIudwpQWa5psFfOEo
+tznZxXOIunkw4jdfrIHfhjy5WuNgXNF/SZyyBh2rhKiscRxijF0QoQkRgc+yLSjwZQjbVwfQsip
jPtMH5upLssVhpXG9G1QNR5Mwo2DY1AeiMJJNX6xSQYMhVsR7K2RJigWYLU29Cf/YcvHUbBBatj9
aqCCnniDZaJpnAobR0f1NIIM+SBrkYTxYNB02aLS3+51sHZHSKSwCvBYHgRTIhw2TlWTzwfMAMHw
5rX9MDh0GFRuThKv68xRzSguanzvul5TzAqvtbUJRxzkwWbIxwi6fleLFoNyWv4hTcpNXlurqkQn
Wn6RYQeOsxNHG81SexJGVZPBixiwg2MY3OZHaCX3Hk2mxPAb6xAAxsefHhks1zgfhnW9Vvgs/QjK
s73MaDCLX8+YyQ+L79kXMXI7vEweQa+UMhItGosjuob1efhPk5dsxV93g4X1KABEbZ40vETkxPpC
gDZf04oNJ8usIE+XZ9LdDONmgt8T7RUSVbVvB0sdtb/J9e4Y3YBHBVN0L0E6IO0tn+IV26MTrfbu
+/mFu7UJptZ2e2rECanj0KTj2aZng5UdqDpyyk7rGV5MT71todHOha3Q/nNGb4xJ2buk6bdPY27T
LPMec4KlnfESonuMq70p3L8UGEQ8YXXoi06k45f+I8ny6B+dZkKVy/eQ7j79FPx8ZyjxIuGS5ON9
KxLfcNcR42dhX+J1PAp1sZ7YAheDlhgwzDmtD7bwdJkY8KjZUkYLfrqlEI2BXa/3V9tx0eer8um8
StBL+iXIPi5xo8l/432YxeyIStBJIOohdtwPsY9ZK5A7lS3Ia0H3afLWxUWd+IJxZkODDxQXoNYY
NSN4g1TFVJK6Ego3Sq3gk5XKvhLKgC0hE70j7wLFVeaTtTuBBNYOb3f23gY8DMKgqBfBmrBo3/WT
CwCnbtiuPfvF8yQIB1dIa3ZivWWA66X2XHC/9Kr3+wQfk5g4X9y0CL/MRVksN5d1AhEno31m/CVX
eyA4iM1jnSvHXTfbSnfy2oTvVRrVh5/os7CfR8eOyG+IRPMqpevszFqp/NGM9TTzuqKyMV2AjXyW
DW0OjwDl4Phk7SWv7ZD23QVeUI+057apBCheWisbYjWhcyEeU/+nA86H6jNtGJNCP29AFUxBEGIq
zjXs1IXv1iRym1dBWtrGdD8j9j0jTafuJLyXjljUTKs6+RBqlKGtC8SGOmpMK1raT+793lXRk1Ua
1/lFk7itmDV+EYgY95E5809v+jSMTKDa4SWnMEfWPFklIZb1TKAFtZXjk/td8youkNaDqfR/X+T+
1w5EI6XlJ62ErSWV3yaED1I9AI2BQefZATFurlEjbMcbBCyXTgBYgS2zb4kGnhCR8Y1wgxQEfRoA
8uBRjRwvNSDtLubkAJQfkwq4irVlhRuRCidFqABj3ogVw1Bk5CjFFh8Uy4zL4NMDfkQ+9114HCMC
2meRDk+DHfx1Nu4eiKFWRYRhOY54yUzlWORAjLYf8chHU4AmUzwWH/PTwqnMdhrU4B+l+RLS7+pX
jAMFQc4FwRrLvO+6t8kEBOMGozJUATNAbYJk5ZzRxmxjm31yuBPzeg/Seu6qvc2k3CSA51w2i0QG
GrEcgY7VMMQpuJxELHCdZamtSmfeE4hDaBjczMu3seeIx9UZVHc/hAr416YxBUb4SbabiB5lVLtB
y6SIjWkNr7J0qFOFL7PprI81F3EQSGQv2L56aWKdJJxQtZ0N7ZxAeZT8GuTYx7dPxIOmgqIA9FwB
7cJ0okJbYgOFDsHlry8oSmxqAatzn24QoAyLXEdIlyhwpfbdVNy085JCgbdBm+kls/LRaeKMzQr4
ZcbUFvuL37JopLU1BP/LTajeN07RxnDFOo+IZFH28Wpx2Vf+jcWjFtwT0iOtaZErtOWmSZff0Odf
O2ViS6hIzZ4mi7VZe/qKcg+UAGS4TjgOn8Yhfw5iaD+wJHFpv1hEZzvFrmMI/MLSXvBxMKA1i9oe
iMU2y9YO57pysqlbwUz8mg6eXLLK2zMyzzAQZJEozzKr0QFNDn74D3WEOQf9nMGem9bHl3VLeDqe
DoMtR9W9/hPilsrmDnenZTlmraG2Zj4eej5DCC/Ec8teVOszJieyOUYy7rRMnrjzHnKc0w4Ti4aZ
GGGADzwlbKV03uCWtkusytAMVFkcw4+UJ37Vks2pwZzVx+CnqPRj5meksSSmLYVxMNWz2S0OYQmL
oNgQFpTgLoZYe79Qi9kBd65R/82srz89QDUEjfccq1dS/iyLIi1INGBgF8TCNaA/53Ihj8o/yZXr
wKBc9eBcmuDuC5bMaII+XaWw+s7bbXAJEjEOZ5tANf+FR7VlVH/1Li/Vc9MQWbXcIBlkmmjmVka/
ZvmiPvVcGODbBj68/6qoqHfVrq82q+MUDZtATHcgNyfAAIZxSDDsowhsN/X9WSs6mKBUgj19tU0t
9zQI3KdkWDxp7Pt04nCTid5772ixxnSDZUuDRHsyssHpeFXbPNLmL829QeX/fK0h1Yw65TYe6hdR
/c2F9OVVKZWzPqpeVaIgANLsCX/7pI4X+g0CezAWf+gB9Zr4747EFUvq0TtSSFmXMYt/uBF+IBR7
UKC57riqL7ePhVS8VicKoSwBGRR0X/IJovlQJPSq+7RRhD3wM/WUvTv1P+zyYE/TKxx3gmm15z/b
Pnt1p2vYMo+/1CfpQjZDB1qvZvRyRW1B1Fh0wIRcIoamexJ1a84PjCaym9OsUPnsUtTtQ0fSleCu
8BFmlvm9/KtkuU/gHJdUWvazBedICvG+3w1Y3jOUHD8SIZLQJfEuhGlNbnmHf5pZxdVvz1FDHmv1
zLLX3SZv6YbwIhHWezxB3KFsohItqif1NBSrGSZbuHTAdmboLXW/ldGH0iB/oLeD4V13TmG5JeD4
3Kd5uBD9yP/XdKtdhKih8wjUlRK9J0kL/LGooGYgmm5TJ5JisxsRRYO8/tkJqJRWLifXZwWM8iWh
pgbDA86sKjWrqi5+Ehip4UMUu4RlChOMKynRQElQs3mMeLWyLsjO2uUKVUqlEg2tNwXFZvtag7NB
028iMukM7ZB9eR0mWxizOknloPxNbpufHyAZO95fVeOwC6yOiT39HtuG9fL7CWH3vSkviqOcis7M
zI2fTTRiXM5vcLZDSBl8bzBzf9JhatxUA92sYAv4IwaGlVGX3Mpvknzg2BWGL6G5dX3yeKNJlSed
5MWsoCjMPvKR8vv/h0kAz91BvlJThUhKIcP6OryxcMfPCNw9NUJQ66iMo6UxsuNgz9j3Bl1MrWLm
raJMUrCfaBfCxs5okeLNL4WGEAfsRz8a/JgGoABZ0TkanfavnSYGq65JsHxv1FKxzuYetY/k50Ts
RA2wYVoSGQu1ltpEBCN0AcARdzcdLsm6/GsyOZVL5ywQuHrQLbVw59di0n2SwK+OEoZZJ5ikBIn+
/5kq+xzcbBfzScraTwtEu9Esc0BQEsKZ2jggm7g+ONvFc4YnxquVAK1Blf3UBf5pqvb+Zd2qaKZh
ivr9J4nnmrZWLcw9DndMGKYsIq4urx4xG+ucLaF9fR0O4TyUX7JaS1YHkF0WlJFr7cwUispsEVff
H2u96mW3gqJ4k4lQitFiihmgkKrxEcmZRyJEzucl75F0nEsl9D9Hm9uD7+9X8msSxJxujmUNRILD
DLbhmcBILZMUrhfKexq6JXsJDNvEXdfPaCPEw9vLY4Z2nQCjvXoSgBPhU0NitvWF/Mh/4DxBwuC+
Fum/ZYxIK2Ta7vf+1ltoVmZTJQj41NRUulvY/iYQB7oyARbp7WwjZL2DtJciFR5i4EjnxXP75kgF
TvMVBQYKx+PQHyruO05kREEK2qiFEtz91BKXuM13/Pil5ZlovIeOzYTLu4jEr8L7mPvS95+RY9XC
ooTRy5a1g2HMlqCf+gVtLib+otYr98vKRAqSGbgh/iwIRx4Ph3Khif90giqDldCn0/p3XUOdAETr
Bg/wiPxI8geHGPmMDjIisg5PRqfHkgeCVH4DH4YOTvNQI0ZxxLJGiOdwP1r9/rzNfkMSV4flveQj
6Im5cGQ/vrFMXd5WTG0ytqeBWEU+fpE23Q1ztFeDuVh37aOqPNofPKAiEJr3/ZBdwk+IhXiM2Aup
EWZs6YvMWrTHx52BdNb7I5pbwGMd70t6RDRzLEHSUh71LI6KwvUxGi2gG3SsEeARKVHtzifZVtXw
tURwGZYg1MSL+X0EPBaj4i57ggFe3XZxGs1PZ/fQ4/QPBeMdzrGdNSNM0ra4NZOnbaQ/vTD6yPVh
YfVfinBiiJamzKqGqlSm0UXZ9/OYSqO5ksA443xD0bboq6c5k6aVQFsuQ73QVttRdoBBuPGbUmmh
AiplPhnWLVkAH0M2UTrBxkmkYTfzY1QpfMTI1JVTkWJimx1Ke0Qh4BGE9diz4lrKA8VhHjhzB9VX
Ag8ze2ihr2q2AAeUwCtxhr0LMdv4OK38dkuIWBj07aMc0fhQqn54x9toIFU9UOsa8ooxn7mqbuse
nGaW8/YzP1NKsRRxvKKAWEFcC2ODVKGGHzRiyOC0+7UfSdThh4D7sJIyxITfxSNbPzan6dbFz2jY
7dhV6UQPnSX4MQlEfEJFMf0iTQCkPzrPnn9kOj3WAhj71vEtoQSV1BET3TwdLk60nq6qTnVy/XxC
b2Or6A+CnLstd5rodqRhwa1xVsnyp7T7OlvkUC1jlBKXCE+2OZBHIHxF5DfUhkilauKLjr4wLC+b
2pavqh+kLb/nMh7tFgNmVU1/whVV9xYAGeKO/UUHmQfXAd8roGjjTq76U5ppbaQebsRU54tDV+jo
8thVrGobY89a/mMgQcP+UrSre+IA+Xa/XLXm2A2rPmog76E4cIws7dwuVzmCg98ZdCYMlcJltvbA
qxX55d4ja3wQh/17mt7Dq7ABuXS4drT1g+XA4cPLHdoWWE+fQVfsqXlo3qJSYRyR4Gx3CGX5Ts/z
vf07qTBKkrrzP9TTWizCTtPQir7YjZE7faKIqoFSWGJDM8sJ7FABAgK0onPTyO43EVqDQxmSDKM/
wMflsc+6PlqJ/eaAroPmYbS7Bx2t4+J91VjGm1M9hnF/PtuyFKVQYb+j+VfXi0sawEhB3C+Ke5Qk
N/oJI40cDVt4cKgDpJKM20gW61vavK8WidI6HLTFsSbArVi0gOPbS013OBPsZVYLki2YZJWuGOdc
h1a606HcJcbCaRVLZ5mYtg4yYTn4nATW7UX/aKEzFiYZjHMKveeunwgfEAjB0q1ygcMvVFYStaTF
V67oLAcYzRLkZbzeceioBLRoIGcZVf8RPK/DFLJoEGkSwSOJJ9UZuQf17eGLyt3RhkO56nredNjW
J7Vuvnxi6Hw9m7vSRNax7JxiSijUPzGYfhwQxdazEeppDeWyQurumTPblI1szdPxJKrGlf/inFnJ
yUimdPg1HD59iOAphWaf5qqCP9EQiB9td07L2tFqLi3KxZwraAOicDMZpiSkiX+9PuumeFpARwG6
lHkIzTVxwNH/COwM+ILrmRgSfHq3d/3Gt8p2yGxZUHFjIPvmiZa6RrkfHPFMy982WdNnaGoz4RYA
JJs5ZToQGpfdyhhpc6rGll44PaXT7H7+y90C61DMhajWahCkoCxO7F20XwmJfps+7inI2OwuXq4S
ev3RXId/nUnqRBXASffq1nIXj6HzAKsWHCfJbDwkYuVl70zWe6z5gdWeL/qKLPQEPUHg+j382Wmo
wvYWzLRKMUXU6bVWaLTq3s2qhK1KMR0EW7sXdnsVbW2yKOhRvje/TdRVq7115rgjNxUhuD73Vm9M
KIOaU5pXoQbw82s/GMfZYLyugA8cO1XJwBq3Tt4ivZDirRnJ+gwlQcfONB9pzatiIaprzlmx7M6m
zGF3eSUGNfqbN1t2SmxwDaU+v4SdGabHX0w/1rSEqhYyl6Ohmso2GYHF98VO9/+lXfaDnTQmu1Br
0dPIV8R75kUPl9gTkVi5l2oJdpmrrjlyOgrqDHMjDlG+z7W5iuuV3RDoIdgGeulBDGIuDULgmDBO
EfUPA1EJI4GC/mu+bEofWWVPJNt6ozq0IWZp01d+QgjtASTR7uURrRSeHzlZ0l+yDbx7zslzzKO5
gnh4vRAmYoJTQT7LHQZzlKFfvcZe7Kt6+lndObzzNaoFzhES1M6HXLOZCxgY2wqn4VF6zmlUGENJ
BITzU9xoAU6jF3Ac0ri/EpoQmu4ce/FgWpvaPfPFQNc53fXt72RPN2A+aTDZ2nsNJzZ4pqAe19wM
oWVShwkC52oRzNcUNevwAog7Xta6m1tmylnq1sMXtBeIPigyn/PAxTmAAwE0vMsvgHGjGKAeElDy
g3MsUjbZpIjRqnIdwUC5vtb9bl2Rf99dKzwLVCmtqJAhEaBEWdxUeNiTIKnk4LpYPt3RusgKQg/j
g1/+tHdFu66mlwR/ongggW9FaxpDfon9ZOj4JRvV+OJVjsyKYAsz8/KOwP6KWVDUWJKHrZIOiK2O
Y2Zq/BCj1c6R8kH51pReEwI/M3qh3XoLQuWSmcBDGqq3tfJs51T1o1wOQ4KCEgXX1HlHDISjEwqW
WOPnZEhWkfpZl2yiAm3nzgGG+cpckNj5foN3rIdJoJHWkIt6qTJae7AZba/op3a9mILoj3mVYm5x
fTpfX5dr4GvRyImIxf6WGLnmZewFnUYirA6xseiqgBALkLIyuYAGlK6K2YIbcvzUr35cHJkhFn2o
MrquB1vyDX8UM6Qtuz/qsqaU/Ioa/mpgRpFc/aBuvMhmjC6sFIKIbstlN0HSOPmEXmZAJtwfCoCM
jr5FLuQMqdRYb1kkBktKui0zR7Lo9nbO4tygn9JA4OyGG58GzUv2hMo9i6/VdR8/k1cwb3OXf9ZL
xNAe7v7xwP2gisYrfr9o2kD0PPVa96jV/GQrzOwDKJNrY6NdI8hPodBhZ26g93DAchydANegnu3m
0kUf2gefup7PFVhFsA0s9IDgavie+PZCUCtwzWNjQu1OS9AJhvxBJYWD8hBPPUc9rsXfTpWinvee
AzbK8D9iYxpwFLWiI8KoLmTZM7Xn/fYXhKKjWp7mYwgcG4X/3v24imFvJhtykoaoUGTqUBF8fO1r
JdX28y1AENrPeOPlHKNn8+z+IjIJae3SRiYMJPhOUsijZz3gRlglU1veMw3NGwDraVL59QCmMX7K
vN16sBm58x3+8kmijjW7nZL7OIu2BvcaSRkjVnmqBI7tTvyu7XR6DxzUDAVs03ashYQ5udqUDRgU
UZflk30qCyic92lzJCVN42B8jYMaOvOF9tjP8CfPvKc8D9fsxC4a74QMXMYG7jtoqbvtEAvJwBX4
GL9v539xCUYmS/Nio7WYIAl+8/AElvNFlJ+ZPZFAvm4Il+q+BaAyZHvm3GSBaaN2E1LihVDqgN4r
Q0tUm24DkA4C7QVFYBv+tQr/SQbnaB0zYQJt7FqMU7QWyyXuqW7Fjwors+VOAdMKeJHQmMHZNhjb
CKbwW73CIjic0aWh87WAg4aP+OemdOnpx0+iy2pnSCRsG/FqiZr7bkZpBJtAxshZdHYtFPuNCV6h
Fk1YB4lYftd130QuMVKXzBEGG88UASfvcas599SqKHSp0ys5OgaBPRsySiUKzDkhrCQqfh9y+12O
XADN3lcUxdMvxMj1S1o5D2J19gqHHW7WlZHcfXpv2ko1KgdmrkK4kK7E0ulAvbM7FKJ2YHe2j3t1
dnMoupxjPxY0EHH3VmirtW833hmabOSBsgNX3EUp49Cn8mAQcIrAY+8/4BtEHXoHLhhC0Ya95p5B
wGYRnB9GTyuFAmWbLDtCYUpuFJFqEy5cYHy9NmL8QOuDUWFIGIu20Nrjs3FTdJ703ykiJStQSe82
VltvZhfu6JH1hLI58dmjyJ2BuOtVTaseYwN0tEo6YEXQYsqZxfTR9m8ZE1NsFzTq8ZMW/uVUL6oU
ibiC/1GsdtRSrgFGugU9vvP614o35zqpFPC0qN7YfVc6+tARWOuJKR8JA0xzgzpOhXpXY5IoVQn/
4viRDOhU0d9bPPlhV1GrFmWXVY3fiBHdTMXggDnygNxVaQ3yN1NRd4+ZnsVqqqk0f9krIm0HXod2
CZgrDw9K5lUnKdFuiJLYuM6taa+Z3d8TG5bPCNd3TfpFzvdZRwqMN0AdqUw1v3ZkKsaNyQsIUfg5
aqaVqcePNHGXIpyNVU38l6N20rfRRcE4JhDYPYwiI3p6/GT/vbnfGv3qFHs+kUyC7eD1QMqXZ1Rf
0Gp8aZ7UzfYLjKhwjy589q5briKF1fvZKtN4ZJmBfkhRbzfUFXvzDMyLuGhSzQW7Xx9/60necBsA
RmV2jWlYNj/5WOtb18n7amrfu7hqo2gGIlyC9hlQjrI0Q9lA2lEHW5E7a41xY6eALy/zKxNlaR3d
PpXkkATGiGQgvm+oFmX1k7PYM7vF2YwHEFcAqw1+HEKnBeb3UTsv0chgBwMt9nOCp2f+YDiFfZkH
sgq1xPGiAPqOU1/t3C4P4dlt0P88BhcF+qA96zJNXUl1azm/lyiNvMBY0IWFqy33Uo4o55N5oODS
5uVqtQRIA0K9Avsh8ziK2CIsFkgDgGofPZK8FUFQt7xFnQitlmZ0IGDrVeAvHjzcxkszOzfpYiTk
0zXJLL3muQTg1gW6BcPimlA/EbjhCq0LIEZ7vkb71uJBmuocQi/FCdwwQ6v8zDzmE++osJrGSUdx
Fd+MjXPPx+dBdqAHjvvpoYPiDFjnmsyZqSEY5Jw0uV06WMOJM41LzS0JAoP9LgIYJWKxltvW5tSA
h47yZrA9+T2uNISLxgN8chVL+0Xk4/+ldlNi3lm/N7xkBim0Tw2/vR0cSe+ehlYTe1RFj4YzzMAE
7nja1mENcH6/nyqnEHifvmRiqhoV/gIKYcBEJYlJ1uG9vVgYbz5ktfEENkp1rq/K9xA2StUu0tP3
UKiJ2/1OawVYWW59UUKDZMzt/3MdWpLJYBEvctxgCPyKFDyrZ2CulJRIouXu2qzFea/RPkos/pZ2
ItxE5xuXrPytB2WaM575g4FWDsCgzaW3buxFM2KctBk/pb/UkLy3Kh1VZVaNCllctvNIan95UnTz
Oogk+bALaHM8c4JU/l63DS+EobeYqslWD0H0FzuTueUfLgrladiEi0GatarSsvdO19g9+xCj54GU
3T7vJXVsJMnrl4o6UfbeZX1bbcOE1b14FGIE5EDSG2kpILP8v+ILWgxPKTzQa8PwFSw7SmhX8xWm
5n4hAjvX6xa3Ee4PfkO3uTeFGRSJzOGLEAUqxBDpy6OROkBrKlM4QwF1ul10G9I4uDaFp/Z1yFr1
S46i00ZnzDGjNOeS/xnTEGkP/XGWJcUweWeuBbqoBgsu3PIuiGDi+tImduDGFB8A//3VD1xhknoz
MkKP3q1cMQFyWK/edc7wW3q5RMgJO0iIqcnOitngznv11Z3jUK48UtlGl/sM8RfpZwOedh7WVXM7
3eLC4H0weBRXyiso6dcxYZ53oAQEXcIQq8hG8U8diMqph8be6DXZs2jml+JVLeKBBMHrMQS5MRNa
931nBFG3V8d4hIBclbl3YH53r5eFY0d9gbWUpl1VFHVh+fI8AqXwCcx0fmJaOYjYPauu5vJbqAPU
QTfLib42IsN42nzFLpbTkNf0e2UNRFZQMV4EtfbREwCava31un3XX4VpnjP/mh8YP9jKK1fratgS
4jBvQQZkQKEiD64oLywMWTV9nBL5jvGVuNq+0uwIOUEp7dvMGv8OuxqGmSjNyDfUdyhuNUGmTXK/
S8vHBKy7pAtWsUhSWoR8hgZlt8jaXgPZaPwPCQS71kuwJhtm2mRCZ+EkGGKZtec4SDeANkuvGc4U
vq94CV3S51pBqlTdbc9LCw8YXXoryn1uZJQ2txRR4XkmoiciWjgNFtkuD0EMOlBAdJ29cIqvBsc0
N5TRWYd5OFqUaBN4QGMZ8oFK0pJZsDZiKD57kVI4UfsolP/8fLwekuueJtG43BTEGwx52NrrdIdX
92Ot01dFV68LkQ0bwlw47b77cPDQy4N1r7gxX/BAKGR/wrbOKVBRHAEXGGwcqhm2JZ7qulT4qTvF
MON9Fg+7jpEUZIb0OaTlu3If99LknOpFXJz+bQ9Ogw1bZROI/JiQs1MARPGkp6KgBYpZBwYFLKd0
wlfdp552cc9xOfOVLsrNoQDPuZj6ZrPeUN9kkocovTxmvxQxq7PonqOlhlEu1fB5XTmrT+QkLyRK
3iPX8RO8r9pQ120Ipa1ldcfVb7JsaUdVe1Wy8cWqIZ67odqqWksjmB/MvYPq5NQPEUYIA19nvA6i
ZsRxj0PCBh2rUFrg9OPS2389poW+SejRZyWvx+owHrU6QM1wmNdptPnvSTupYFitOd6nUe6qdNZT
F9dvyD1ErjQtwOEt/Ur5IHGBCPaUJrF7rSef08y26Qm6A4E2T2f2IUPy7nEf5ZrVO8RrjGJBDC5v
24bJs9YCHv7z0hqMD2DmgVHSxxOqlgiLvFQIXcoluYjk0rmRi50W9Ss6/T8ztjFR+wspMEnbrID7
ZMu3nGpUyf9fhX6MUL+tVX/OclGe6Wm5cxw0l2yz8jKNGCATTZ8PmOkjcfn9trFQN/+T4pi+rqjB
xekDMy+MkNDODXpMpSt/SWW7l+IZijv3RYVFzCKwg6OLuGAGb/wGjb4P4Qia88V31/bbWPlq139y
8tU85VaqQ8DcC7mIpu0/nLwdHfSbxGTcLV5z5JlxFn9rVd9kfBxpVlMtvuygE+2/egUgFrz9oE1w
LEhWeMCa9MaMiBLDRFn3yxb0sGKW1SsVSv9568zy8kOHYwiiUymvP4bySQeZvUX9ig4961JJZ6G9
lpWZma4UAcMDyewX5TWy9iuYJRjuAUx/Rqa36tE/wMYZ58uk+wJrQ4LFAYBY4aEuMHrK4oa4UU2y
muDvyKU/YputEqy4XFuVU+2Uq/Zz75t4z42JYg1JEBuxm/EHV38FTbg/4oEYMj6UUFByUfWosUcQ
0qlrZYlR4XHU2ZRr1XASjdkub27Z03qINv1SbY5sjXxO2lfri79ueSX0jQK0BjAne2I1dSy15VJj
jRe56uBegRKLW6vj2VgKUemIjGyljImlDkt2rjNzTpK+EkRvG45UuvhkYFaiFybEjAqOSZ0BActW
UnlccF4gInjGbkGCTsQMCRSHIm+o1IPSueFnmdvX+ok1XvL2dPdaf89UboCpaag20OSYNX9APjqM
MGa4x7nNsA/16aXNF/hY/6zohPZsCsDL6qgd96t5lY6rwOSOIf7N63CxNz9WJqJuIDizIzgnORAU
dXtwsqRifRLLhSbyryUmCoCqh6/1kTeBomPGtFchXtPZI4YLPm9Y0zZLvLJbNmM9tlF5qaMxf0QC
jATmYFgYPl8FNOZUymNAERjzMcDEKdn1alFOEZBb4xaNUDgJ+aILlnuqjwNWxZd79vh9cyoSEQdI
mQt5LSHQPcPpSDdftndypE8Hqmo2UZ3segUUHB6xLwwKFU3f/PitKMC3G0CFBVXYjfx9XBRRodWB
NnsLKObmdcDwDac5m4mQvZ2Yl4g+N1AV7FAnQA9yhb74LNkpRoqCAydhVfBAQqvqrdrnxkwxscQN
WsdTE+mZlWLvnxAJjvPz9JmJVgGgx1b66i0fA2npIUU5YaA2Md43K3+IJLmzBbTH+cYNMtC9RmRf
zevznHgiwJFXTBmjCY6A2hRMIlGa5PMkjtXp0N7+b7NSqlotQj/lQnvn73c4RxuAAv89PHyRKemc
DjoQoTDqyfCtz5PGuwa0wSilKz8DNzKY24VFD0t+lknQxx7+Zk4zB1562Og3AjXauuCw+giHNXQ8
hkWFQOZ0cHHshG3f0KDCIyTr34FHw8g6h3PP5+flZ74m0mHI9eFGLzTVHdeOMjmFarlGEynmHCP3
pcB+zS6wKrAfpUO7YPZrXbSP66dqD/l5lgKEWrN70x9jajHHSvFAPkJHCBG46hYyOK1fWWV7FVS6
JjJIBnCCDUc1J0/V3yVShjHXDKVQ/4UzWgbZya034Z646hkyEkCj7eoOhN8jy8NS8do/AEe2ulxS
1B3B+UW3Lfi8serOkfI90y3e0AGjq/N3TevIw+5y2i0rPwI5LXj/f6YhR7FC2HVf1fKcc4gE2ywl
GgtWzeBrJKMu7QHc+QwVxeohRAlJ5iIPqiS2vUcQWWO1ifIaqWU/7HoLGXE4SmUUAGGIT8KG39uB
n8jgJ1Y1WagoUj2nG3Mxrk8Z5rjaZ/jmXXxJoNRdjTErqKUlK+id8KjUoKtccx9yJ0gOtiJH+lf0
FFt4Y0OVDR4am2j/XKVztJDV7ePUOdhSv7E4rB1H7Wb1H5062u8w5edl50XHnvZLieRp/+hHOO7w
QjV/NeqySIRRBmi+IP34I84nx+7ffNHVWBumMk2jA3trKMXV8EX+h8nuchvkae86M7TuBDjSHvhB
YXWiDXg/hy5A3dvPrXONXZ2nCwjIF/k4lNv+NIAH53GRRn7S53ky/RjgL7sY/xdO+rGegV2Bw1zv
hiGU78gB9V0yVAUeGyU4LeXaiHkxFYtg7NWs45KtaSh04shfntB4Tjf8RL/bceeqASZrfNFTxA44
0HMXiR6DwozEKQ8pI4+s4zj2rLpsblHXpoOAUM+KNNpB4f3BwF34boeS6YqFDh9U8tWsB845D8Uu
h2059I1XVicJrhJT/EzGkSa1ZZ41bkMi+Pi2+u4nEY7irqAKf+QXi/fXFFFnZ44oECzRUakq+1IX
i1t5LwWltpqZPW5+ejd4RqtWpCsOyb90JHf7q1E8AnFOZMKO1qWXy8WfVa3BWIVphLO6ido7d2I2
2zGNj/p5lZgIN/2BPKXBKXFwJNNkYlfId5Y4CSYWr7u8qZQpNDtY35xtxgEeSwMB4xI4Z7WtVqHE
BpErXIVvM84LYLUvxX6I3csTCP2fCjNiGygcDhCMMNKJI7wscOwclo2G4MXcGspI0vwdKpw39iBv
WPApZRDWOv4TWvZTH2DtT7HoJBfS+GIsVoe90FFy7vFqaPSEl94aMdpIJ/Liw6uemEw322itDvTA
crTuXPuX2M59gL4nbrmRRRgmcyYswtjB1bvL0B7jK7tzrNjn3tfOnpizYQEPvKXVRjJWrBDZGYQ+
KqD58HLH3cjxWgw5QgFZHSFu+siXlE8rnnmZ2qgpaJOJtW1brIOoEnGZ06wjGNgICeu2c8Qm/TOJ
AR7nL3cqS/H2azc6oNF1BQgApblaGx0BA857ZigfXkDx9L8EGqMieTOq5uRjcIwUBabBBSDctQHQ
Wj4KL9IjIUEVdC6KSbgI6wyHTXNqVzGDYqCliBCatgV7VYDyQ6xWQW78lXKwIvRimMZiBmQpU9HS
40/6LyC7G21BuF/hJpO+WQwHUkeGPK6pqThyOYm2lfyGW762VG8k3z/ZXdMpqj4BFuZp6eDDijjh
rz7yJxZ6+AWyUA2Glk+jKznmHSNcOV03yEN85wCUfub3LtSYtcYNXUx958JmSEMzt1pIpd4A/DWm
YYZk6dcAvVAwrYZpeTWO56V2kWlPlPRrWfy77iRyFZO6rN815xjuoH0KwmMUrOc1ASWX0K2BnBLq
PuRmp9x7eF0QR+HsX8CNZOhImdEbcU0/GtT3yeoVZc5bLV9DzPY2F8pGF1eg3fVNeWeHW3PwVOUJ
AbIqYUKMi6HJip/Q1RX32whICzxroUAke1ZqqGiCpXZfQEHA3V+LhS01RZwCHb5gtQ0Rf0pN6sp2
y0HGB4iT0r208x0qqMAFrbggU9LF410VGdG9q3vOG3C3KdvGmLKNfuurLV8ri+GpkYy1o+BcB5zx
P3/HnefOu5lol40Yzs+iUvEEEoDuk3lgbNUwn3NNHY9q5tvqE6bEqvL1Inp0uRH0BRn5aLAXda8b
WMheUdghiYA0vi7UY/pRqbr3+szQVIzduaXSm6cUd59OyEeykFskeJ+6IlWHc4pybKL68NwUAKrT
NshzBZ0Wtfby9iaukiqxmRLm5Bs8Wo5HhpapGQsVvXkmPoTNoG1zY//kbcptCnFqRW5oooBCNawa
NTwJlY4lkSRJ6tGTzoXjaqfrflaehmSy6c4fbEPoVecQDMd7tv24aa/0sdnf+BgBjUMGVEoSaQ46
iGJBRi+6hut+7+yFRFCUS3tWfLzWsLR3aDqphATIKutFk65du5ub43Rg5qFMetJ1mtophhmRAgQK
N64P+j/67huhGeEQB7eBFhl/8E7AIlvp2WvvA6SOODpE5VvheduzWpZ609RscrvEFl+T9MUG1oip
N6DPfXdmGgWgWYEU0dsZ82ic2M1l0S8tICCa6r7rLnR29rtnLG4cK2qg3nenGBqCLc/pCSvPN9+d
6wsjpJrjvP4xAEdA6szVG+1SulAc3QIV1eZSpP8D3N4vSJhV1c/ONcn5dLRKNYQ5U0uO0tPIIyKY
DuJA+FCnygCRC7L4O2RnBaWANPuslGycILqxD7FHYdAtbDlFha1QavksdLNZ1PYZaUraPQe84nW1
V1b2y8LYh1xPQvf9F1Tb1RhlqDTt8EyhO37+EKTJVen/7aMAEk7Umvrm7YeTYtwWrz2zxOnh9wvc
j33yy+O5uDiJXo0QwZ1s7dMLVyVKFOXoH1PApd9ezx2BAHgpikqdGiIFTAs86DVcB1KeY4QrGhuc
LKg2A2az/fI/y1M/jPoXYlBfLnUDL53w5rXwMYjqPToXTr4gzhK2Y006gRq1UdhRno4feNEcrbQF
HdLTegO5D4XPRvI/VPbHigrXQy9ti6dgHxHX7NhrmQrOQobTg/IkqcpmhWW4zixm8ah/KJdXTBu/
ptXf30neuBNwD+uvL/meFCpuj5jNFHjbRiY3wFNAbxAbb4nMeRSZmPSs7bkT3RxAws8Mk5fVMBM7
bI0+uiz1UxkO8pYgS6ITa/swZN0t1qHCq1HQCC2HvmuT+68SmpFpjc3eOw2vE7GGFNihFDijtXkv
y2qkR1yvKIqZlMajPDsM21WXDrJKIVm52C3AYmEhRfbjKxx89ppN1WuqQLsarh1yjo2p8uX3aVt6
dTsIf9WySdDu55z2K2nFPRMwJh5AnYYB28ZsV1Z1fmYzINxzewUNeaU3McgBOOAH076foMMXOcPY
Q/SpjbtUk7EDI6q1YTKHXjWc/Ji5bFmfsdCXnNcmmEDEFVRB6LqkkFOJkHJJQAy6JaPrpI6uqGUJ
GsIRPSL0eSmlu5VTQSAfYyfAI/PAAvPIHm/Mf6FuvPXtj7ZcRon6TF3KLE/McRTYOPhCrzkkWSMB
5H/yYucECuofECA18R17aFt4kgnn/4WfPoHsrh9zZWpT/RaOe7U2WzzAdQgTh8xNOGqoVssqCk7E
iXX9SluxDUk38dpazZ5mYfkqr7o+fwwXIk+Xkc0CPHTxl5Yydf4CkG0X5/GYUTQ6R8DGvVP0OnyK
gQIfz5J56YfnIayNAKU84udGN9/lBf9mdhpPQBoiz5KufyKaiMqvRIEO+qIdP1BFa+dJxfADmIUN
NuC2gZ0K3OUATvLefDTU/1woZVUG97Z5IeqODiYHnRkxuND1IXLeHuoHvodFG4jvaRkIPBXUlOJ1
kWyNWuAxyXrIDCnJ7v+swBxyIrpOWte0yiF/GQpPrHlzl4chTYpAkqOnMGo9LwGHNrxSyZ+OV6pn
vGasBUjzb5kvRj50G5sWyb4I1JREiqI9iJIYkpFBDz1ilOAP7YOR4lECkt+bpH+RRz9tyCoYaTRJ
BGQhQRjmrP0Tla8mb13ITkT9jmKJiy0iPawBiboT+4JdN83vmBi8Fd+Bno38+LaTelr3AODWeny+
t2EOsjbUGtrFEHx/fB1hvfL7a4ZfBZzkyXIkAieJad1HOX3L8tLt2fpEes6obWYdnAqJ6FjFxy7k
SNLFX3Aqlpy0Tr7kKJlTfc4uzz/KWGPKQ2GmTeJa2t31apwk94IxZ23IOMFCyk9ETiTMBE0dHbuA
QkaZYAOcR5OZYmqYeBEJDQAPhAplBr9m/cvN+6BmqXybKJd6duDzERGhqQjPsDDR48i2oLUtsNad
xKYThKPEWkiot4oSuSKB+0s0gOTiynGL5wSzhsz1soUCtOtVZ+hDKWU4SBjbF6VS9bEBKKPMuwS/
yTXfF2/RKwWfiQjsxim171jTEj7G9UoFARF0g2dlX4Q6z3GfmfzNvlJANNlgdtTFIw28ElMaDWX/
+lW9F6+91JIbOYGQjDAzo9NLkqJLPOMIWHA7uV8rqXavMq3zrwBUm/K61JnMnEaLYAkIYEvgsIU9
PLAMXN8aPPREsYqQYOALM+eYCfMKEYvn5BtLs11kDNG+jyoSRDnqaU1RKWS8kMpQceE+k/MK+QZE
ia/EqpEOybyvLOtUGH5PW5q6DyPBLj6N8MLaGkGtCq2dPzoN2zPVdT/picrxI3p8ijs6HJgPe4Wl
tj/H7dRZ/GgOVhv+zWeUjih8wR3y8UhGjxwDVmeZwqD5H3N6BivjgLs1wYpzueZwDW8j+rk4FH+v
5Baw+pBw4cWjHGj8l7Cug67ZHxco0xKXt/sIBgy5LX5/wIlj7oeDTAe+rgXZSj1cYeIGuEAV4wC8
c5u2iGiOK1SlceF+m6JnJ2WLcY7wkAdfE43AUa3ePqVfrf7yGC81s6NSyQ7ElHu1RgdBFs9i7gwr
X4bKzgh2ZhuBfOQmvMlfDYoJiK2nASi9tZmYVCIoA3JmG9C/WUwhjYeOIjxt6rbHf1VRFmR3DWMc
ulaJhP/INykmdmB5rcRIPHN8bObttO8kAnmgLisnIUDKlH/fUjKYkvrbxszB2YRmZLFGMylm5GFP
B/KNOG+K1jKNOYKgjIN45xF16Rrhn4pb0Lu4pNXn3kn0T5+gOscN3LvN3dFEClNacuCdvP9BlO0u
K/Hw0SfQZ5w+zi0QJJjSlcPhFpdi4seZPXIUBq+EMEnQ54FY9v+ae++Wih9FJJrjPtFBNqheDWyL
VR4isuL0Pz2SdfQQU9jEvIfqUvf/xHPm/Vu+cu6tDwL4r2qXJpZfJYG1Vx7aS1bsWaFArGBV6mXE
Cg+jXvTQGFVh7i1a3sPvIiL8ulETPzzKRozPzDpd7xxOEKHPGNJDClEyGW/T8wPhCBRdkaBBP2XT
sXP8ZNFjnkW2eUL8sPY1g7TT8aZvgq8amCTuDAJjfBBtJoFSgcSeHQse5s0GH2K/Apz3yVoUMSf0
NK2Y6SXRMz0RH+z6CUiaqLgn/YNBDkI3X07xpIutXcpyTtrBsSrYGX9ZBEi9cIAq7NBhfGY+BTDr
VddIJFaNEA2BHy8UZMQj0PwaKzzmCqAmtQkSBrB5lwMcOl4JxxwFa3k1HeK3z7yxGbsOx9wYi5pL
tMoTW23+f5OIFROlI/X0Byn5RJOf3NzAiHRMkqt4E9QO/lGdwvJq5k9EbDo8Px8EOgpDFPohJwoZ
53LKDQAXm6RODK0u7hLz9s3DPQzXxXZXXsxkxKN89dU1HhgySRVQNVudqgL5SLBThqx5OytuXEFv
mDcV1Qx6WooDGPX/8O55x0qqOelv561pP3q0E6cOlUE+CcbpE5gOpWuMqTePr4Bs+RVkRNZijPZm
EnNA7koveJs4o21VBZoG7bOp3WJUTUZsmM8lNXjjb57j/cTQTjw+NgloXSLpECtfONadVMQi5CsB
RjdVQNSHCXaGeQVj7mptXZVV9U8uMRCwCXBhmoGHtl0flbRZWEtDVsLgr2BzFmtkcfpMur6uQTMy
K7Fu0YzrHnNRGOZN/uKTWjq3zJkaorBIalq/jsiKTLnVjzi6sEBaHoRGBx3KcLzjPkplIOkxcru2
S49eRr9f88oR2z/zEoGVp4B0ht71K4+ZwH5m0aRnFVoZ8tum6CoPMunlNmM1jBjZzq16GxVq6PGS
ZRSYLirHaaJnGQJk7SsN3Y/n765ptA1dFwQpkXOOtpoQSWXctVY+F6HAj7m/kzmTYzG8WQGeLTb+
34k7q+cGy/9Ncs9+A5NokRjjOoGD83oBDvF/MDNuAO1epQRxvcGEWmGL5zYaJ6oiaJ1ftVT5IqTX
hXxaDX4MmBkfKdlD5Am9gpEim3Pse8Ox60JeyIcb1WRpNRPzuOcQlIgN1MsB0/rgHRaaJ/1DpZWN
2OqlyBsB6Uzupsh+g6aq6csjNZ/VDICqlewhUAMSaCnLL1Q2DfHSi2COTkA8mxCjciO8X+fiPhMT
1NULn1XIM2MHlhqyZntOXvCmSqOwelonr+1E4cCiiRkDsdNifMD/nMYbiuw0GgnhiXOPlibyf7Tb
q4fcsnXE1psIbcv3Co/Ft1oxMNObUYso6AaeDc+E/LOvVg7At3s6hk7xkZp/dIhZwDazLzIEmEhE
Anvk4FTm8FTCGVvoPD16AuesUofBERvilATTCCHi7fxcWLpMoi260PedIF0xTe71FzGjjKwjD8TU
RWRftBBYZFegydt87lGITKeMNlhnZt50NiWD510JSm2w3XyFVbxtTsDdbH76zJvUKbQnwJb2szns
6/SJ+KVjNoSCqzhQMfauU5lc2mLRiC/efvTpyrgr9/V+sRQU0+MrbusBRMvg0cYdjdDISPDOvvN7
wNrqRrgIjF65p9vL4jqeTKYd0YpnMFvqTejv+ZZi1P9oNTadblGFSoH44DvlmGJnlp0l0JQLhhi/
t3Gq2KtHq1rbDan/uA6QDcCrxLnKQtBh8MN+0Ty2FW2BkLeVavf10uSw9Dlz9TQgMeazDTaxGN9C
ZK25bhofJH1xUCpo336XdHGRKefbIAswkRgf1rhE3Kw19H9zstHWVS+Cou1HAnbeIFzKemQR84My
i2k96hyd9p7QEzAx7YhLBjUfBSCtVKD7pwmEQP5ffntIdqgPgb84lAkil5clRsG0wnlOT/kSVBBl
AoWNqTCcvtjlRC5q/RVlc2+iLwGFDBJ80l1z3mKQ/50WE2Zh8Ap6o+6vDChOE9wroCwj9shpitZ4
gAK28qwP+yXb4r/3pJVIPtNpgmTxyz7sUwpfMSJD/BOZ6X1CFzufr4iFJPvuztYnDJkDW/Y8YOJf
KwyAzFRwyOSNPv3VQBJ6Wq/LsH2csKycP7RvDwFpZmO+OeV4T+vBOMBgL3BXlWbMd8mNW2eiC3fX
riZcuJgMfQzBz0ulvzhWnwQdPidFlG6aHou/6/UIgPMvSivsIuCD901v1W4XilYONEeu2rvH7fXZ
iQ1gmdUTYHWW2AgaGnCrKjKCeSl2ZQL2uJTHHl55C+yl3/oi0pBKJH7lXcvy29NKsAE+siMaBSii
sMgN2aH5Na0EAG5kjEGOvI+8bjZy7Y3nQS7GG+dAmCLyo/CtKpon0PUNRCYazPCakk8N4CtmUUgN
T2aQYOiGiUhXFZGUtoPXKtJNEjOIcjTDZ4vWuFJyxcPhz1l81TqaGfxT0l80CyjRH3w07UQ9IBpL
A84aPciJ/RPddBBB0vL9MOC644QsSIy9eMJfqku8t1081orwAWLaAbHD3qSe4V+MdDGeOt642J+5
mCtNG2mP5GkYs11S+dWxsRcARZAPZsMbWdqCQe+hWyzLwezZ+NbszP6u95G8eAjOmkHT+FVI0ty1
EqX8FDfoiVYUqH5fZOW9FsOVRt12MWyRMyyhqaXOu6LzoHr4hH5kgSCQWe6/ZhvNrIbbkhZJncae
/92xAcK5hGQfDcYdAdKACpjVOlv5gcHHrsezSdRfFSG/Cs8PibLJ/Yh8rGm0cj354PjMTrvWcUmk
N7f5+AmAtoJWHuk3qIiA7874IOIFxd10qP6saMP9DuB2rX1FiWvOpgXEhI0Ua7gtWgFx1d9T8f9M
K5W5uh1oRtFDWl3OOA21meTHfIcX7/H/HT3kxR8i6asdA0Xi0h2019JdAj+xfxxmclz4LpSVjebc
ay+FUBbAVTsKbekGP112omVIxXOif64MNgTh/qXjBY2/vzlXJhxub6hCTiiA7XU2M4aLlB5pJVdZ
bPM6kfocMGpFy3Kf09GY/8XNw4BLYdtoXW+nRXRlvEFCivNaS+Z3CyzydjRrDl4lUBx4DZIQfjNS
X8gNV5NIqr5lZ/SLWFOxbEWy5D27opdtOqouF48qGGlNTcxjzXwNVRvYPTd2+Dz38H8Qj0OMwFw9
lxf+eJxLWL8DNc/o6rEuY+ru5qHd7J6VLtNXxpF9bMGJcMDUODQO6TYSZPlj6P6xtRis+Ux9Ocwg
MCmFMe4WGK0fUUIaBQ8GAtnNz5dAX0+zp8b7BXGunNyMhrUZmDCjBEpsukYwMbDmIWZp7nx9VJva
r6OGbwR84TwgI/THpx2/zh1MkYlTpLvdd4uUzBMFLrGR5GmInJN93+WvK/xbc8/v4jJfdSbisn+H
8tKhidgY02t1ayc9PjI6Bg6Z+5UVUca/xvsDcQbs5BQq2TDsQuWUKG1GXpHc/k81FdaJ4hm+xi8q
uUsQFQAUW8/5oTNauXoYCUttsLLk9+WsIQczAulKpegM3DKhoxHRnUjgGxSpuSQvQ8edmPx6jMVS
nmNa/OFqtP7lkyXTnlz613eIbM2G68M8uJ63BisAD4c5/kuZuc9JQZcuQ9fIAjyt3dWHfeLGIQBc
XPlC8JowLWCyTLzZprSeqazCkHsKcZrKxoTdmuSTJxc6pXE688rEXzeD9hPe21VrkkvafpOoIc/0
VV8gVCA4+eE5tBv3+q5bbo26pnuuJDvrvCmUlollAdsXTrhLENqCvwdS269SLSrACFyRFuc955R8
JJNA2eccMpVsHui9mUT2r8PixKdV16N2IAp329RWB8Qtg9ZnW0Y+jAcOEv3HWrwwasN/KmNpKoy7
q49QESyA5pkXa21SF18LLeU+bprwqxTvZnBYkZUpuF8m4CphgL2LOEqosoUHWMg6jXgoi6jp7DmI
iUE+s0rvM3a6P2tq7dWSIAr75EpI4Go8+jHD6Ao59qHZ/QjtjRHZFbELeBv4FNtSWiiWGQkFXtuf
N/mZs+9XRPGtSC9KAOfQPjTVoxEmStt+QxnH++/SXfdOn/C8GHFpsdIgjeHvhhtpvd+zS8dvGdmA
SPRf/FR83cFwXpzQR+oE0dL7DMSTjavYuGnHKaatylnZ3NDOpYB2WDgfK20DtZnf8Z4i9VrTFPd2
6hlXKcxbAZZrH0/t0mn94wYTW15kaNH59wIWzEjxt90rK9N/6nY+Md0bFCCFkJoOkwGILX4dNJS4
FMaA6La28RuNpVP50to/ehA9sYUhPQzZ2rse2QKbAX4Cs/SloDf8lFpeYb0xjcB2evOqykQgY6hQ
jFQSMPsGX/YZaSlixdj3nkhgiPmLNxExN2OOah3lVzCvnsIMvFG3kNE+hy1aJiuWx4pNoZj3RwdU
ABiHepyyeAnctMKG+ov4C4BIANnzpHP5Xf6XhdC5DV5Li0WW3SCgUGWmumfmUULfp2E6AKXQzk9S
1Iq3U2/dJmTTjup7cmEkHjCv2axxv88xaW+L2xxYjGkqk3SrpjoINZSJw1v+zWDS7QrSgamyglqg
cZV8W4B6b5zmkDRDUFO3eUI5f+GEJECmhgzMGds9zLj0MF9Zt0Uw7i6Tuk23u9rs6fC9Aw5bKBq6
xDyDI4oz96tNkaTrdaCHsO7/JXjmfJ6lnMFFKXA6t1qgm/C/mn4ojqB/0ribMXlN82F+M8aw2uzU
A3jUYj4GQ8pgzkayL2b/p7XnsgapJdp5rZMNZK8lHff8HazXT9M1asOhkQ81if1zg9WLT8nsmspu
L+bPKiKrT1ul5CR+l5Lj4/JfBk41LAs0U4gVSA6cVZFzZ3eCzsWfGMRLe1VLEIWSslDEVETngBRO
hEYhSgsigYDi7agaLC7V+56Ttt1MS0iALeQVWeexUWoqD/iu8nWsmpJR/QL7g1HJsu1FRn7SV2vM
iUY4fcb9d0jWEDZbH7N2bcHkBwe0lOdBOJSkDrQ8h2xgXQu1Cx1jutuzEPNnvc/UR/ql9nKrXSj5
/6HhGkP2wobUUY+iDBzCOf57uRvqHdbXzPBD0peY/3I8wXRE+ueUHw5lVJvaYFO3gor3ltDB+Dk2
bQAqw4cj5V+bO4BLRCSOc9jFX7D2R0384GxRvCigau9d+XufOwI/3CYzsZL1RsK2sYNdQGtxemPK
xCvuKYqwZycBtvjcX6okPtVoY8KFsmVDUFG4a6shDZAhejx6K6LiSMxbaxcqrJJR3E9xXd+q/v4U
V++laAKfUFKlBL37NN9QfnXXapeStaOhrUIpXnngV9jyPfOGl5bv5XruLlInOc5pAAOX4S29uwS7
2ItTY3ghWdcXc/viLbDom1p+AM6EclZYLY5tK2rjDHVrSUXvLRJH8Hj+3SW0bYzWgwZZjrNcuPk0
L2xdTTwWzzwHczH1CBXMJHAoXp8oGbXjpbqFoz9qx7L3gfxf99I05NTOW5CwZMHQsX/SOCyD4n5X
1QdLwBU1NQ1fz0oLn434dsVjeV8Go6EkKYKdMWSCCUTpX5280E4JCksJu7uobfyh51Ky7ljiKoMT
4E2FYIs8PpKYPcDdVHxNWIsn9AwI8SNmKfsVrMhHzNwSZ3csy/hUgL/WAajYirjpXwN7Y7giIgp1
8018bCB3Qlb7WO7rfKybTCkqRkH0IPXPt4x3SUGQJczh9eqP4T1i/t7vH5+opdzPgkIEuqGFKvF6
eqRQK2momZ7+0kNgVrCAtr/Hwwv3UAyRZAjWBbfDCF0rglOcbSlpJI3kTooLgVK2DH1nS+wpEm1X
8enKWBdEVR2weGPCAJswjPU2PxnUAbn2r3YFMvpwxI97D/sCu6aZp+lsIW3wxcyzuSSZWEIlSFB8
yiEDVbL/8Ypmdp7f4N4NH+mGCOlmfCuOmhYmdPWi3kDMb89UDaATUvhNXAiSmWuXlgt+VYGPx7UO
m80DsyfhtriUwKulET/49X3PH6SM/KZ3HqM4KnZAdkbnDtH/fTCYTkNOmqUtcQS6pLNEjwVh6d5X
u+9xKIjPUUtgbM96mA0ZsmD/2FqvzIZWJIn+ZCXjJQHSym6R7UjQlLmwpeQZspNRfuQOPz7gtD48
tP22LNGPuya/duPZHpx4lVshB86ZrUo30FH8xtULLMnaDNFLQ8/Zv1GUJ159HEElt9IPoDJ704SD
ta/bzOUlInrZsC/rrbKBYh/DynkzYYRPfdYq0OhmlOw1FPZysraejNBJWsoO+kL2cIjtm0WDJhiq
v+JJQEhLfXX/WnuI+h754NDotwW0BuNUPkcBjKmtGFdLnVsoHvueojgVJCHjysBDJcTxRZoZ/iWS
5nGQF/ehZRA2trjlizp/AJm2hGtmNKp0UIHi6vOhdTEeG6/yxcL58Bf/ZfbZMqbQ1eaLOOW7/g5v
lartw88hHDVAXx2uOFIiTIWb+m022rgrTBq1981nv8aAiFUrowyfAmBd4AgRmkKmbVGbGE02KfIa
pN50vDaO/lHlJc0leFrQclmdXXM3eyUj7imgGDpAla/ohOe61ISXZCdQb+rzhZeYI62ujUPqbJt4
QQQT4wwxblJ7Trsl7srkHzAL6crO2HeqRaBCvWwGH9UZwYaGeE1N4CY1O49RjxUewEPEGXQx8sRq
EhJ9fMTabwS1Xv/Rgn8M5sRNn/zC1R13Cn15smKeQMeFigGLlyDCpCe2q1paC8BcEqNC8lxI29of
9phNW5/+pzhfovscNvqM3zPdwEdQ5y3NFYrMmd2ZKeuSb/5cNQNnTQWs67kR59HRsJd/BJ0MQr6s
RMfdHJdQiXfzEJ99yvnTHLPYUDBoEM/Q8Ny4GBEs66k9NP8GtuyywVrZ/gkkTKg3ZNqnld50XTUy
8o6qOy03zGgLqZs7ByMDrxWSO8mKieVvLeL18Pmulsk1lUc+5JcBGlD5zDea++6rxtyl8b5ZsnPK
FzPHRLVvKLnFXSfexNz3ZjtbnbaiA9ZjOu/LGoJx+c1NrcJVA9AfzdMKBwv6hn39DPglbofLD1Lh
XV4vG8MBfPBiYA0D7blh5Ul8MMec7tzw3UnImG+UwypsyuxMwWsF5s/5c1CkOSeZ5VcobzUkA1gm
jVDi3JaHYBBDEtq82H+awn7WvaA1pdkOKTmNhzCrymWtzNCxKHfGyvSWmM8cEJwyFBrGvtOXfK65
NMP65KLkCxzzezzat3xujzZcOIMZnfoBH2UpFWbaewxdxAhbd+Ak9Oaf89BZsG/dtA0Zj7990Ck8
G6JkBe7HEv85m4EyFH1tuTZ+03sccc1X4LhsAKW5wdsGwGXoXRm3j0R19vUiJ0fv01awa4gOJzhu
hlOivwA5ndIbOK8bPxWvq4BqdWQkIXVXR1vpcFb9blZbfo52Drra+0DCQeCIJlCB/pBFQ2LDjgdy
vJ0eqiIAOpQEKdFEriLLhw5YxVtFBxyGiwIBKl5/8NLNv0/jVEZbxArIpVQujE9hNxU52zsIHGmS
tBZ26ECZIIb4KRqvGso7Vsnja4zykpyWH7zWaK9AdXcpfSK+z6Ju7Rpj3YbAQzAU1V+8dyhtytQ2
DoSlFNCO40kosj0zn7XGlNfgUPsIJbbFl0F37kUH1jsLBtB7nAgS/nC1gLyDMl7CzW8ucdK2QpO+
EUiDZmebcON/9lcmMMtsypYya/o/espbT02beFqfiWczmjaNFCZ5m/BKKvGRXpPA2+5ejuwzVVwv
u5SvzTcv5szAnVbS0Fb6/8OersICbPCY8AaqQzfe8G2HHdmGcfemA1ors38Agme/NDX27e/35ulV
Y8fSoHmt3KHBJ91zdVBdv7WwbJnFspbHgTpc/1crgJXoC+5OGSrqbts+SqdPRdbv9bWNvs3XcerM
ixQjZ9ET4as6k13dQlQhQoKV4sXwQN4KbycM5EyAdvuv/a5WHVm8JWovR2oDNu8fuXy9VTAXJpOq
aD882dWSWK9MI7TFuBiQQJ5DAfmJ3evnOmh3HGrPdENB77d06CR99Rw/4jgrdWoasamohixmcGEd
pLPO7djytFMsh2mg1GfbWxfHbElkwY8ZvrA7i5zN9Ngsq28K0mno5YqquYXVcch7XQyJMTJJRCwz
d4EKQMZGLInj776M5vhFKwtIZ3BqkWLITLG2Tc+nmqBZiEiZgYsYmp4NGmj+yRueAFKXGJ5t3vWB
/WyW04WBRM2sSBj2WWmAbAtJ7qkfeLoTR5pEgrtc9r5J2ZyQRQfq+Em40+onNfzjDN+g3MP3FJc+
DoyQJkI0rxFn1RMCGocTQjupvhphvBlOuwbIi2hxNH2NezKA6O5mk1u9j1ETCm2yNQPwpSU6+8lV
cTIQEa5zN2okDsiTz9t7A17LEsHjBblDUl2qr3i5qOk5K7SgE1ysBfB1XmGqT4rgj/u6RorJxU4m
XEYn4R9pvSGFKiApM/mTiPHqFcO619pKwCQw4ZZ5RVqiLSkSVoZioBJFArGpXnW5hq4R9Hxe5WVT
RUvlfe3AZ9QeEZhaHpl0Zs156JZfGRHQifncQMKwGdHmgX/fiu6r8dyGhW/rg2pIb9fdxBXxedFf
1ZZ2hdhfgKdYyucZvCPYMZxepc82GTLO0+bCqtO95IUM3sZ1zAmHT8wrZaQDPxmlUP/wImLze+0m
N5Mz0e7u++iQypeTK5lQzEB1Y0cYJM1TYoQaG0k/uvvfg/Gfk7EIpFqUG3HMxUMYtS2DMQmmhKZq
lSefF9JfQwUrrlKCX28Ynm7/tIAco2E89ZwvP8VRMJKov78e7gKZ/TnRXcHqnKngeUfz5mb87kCR
kPznKDquuo8v2NwPqsfB+CRbqV1gdb7pDTTkbcLdvOPXFhcBa+JMbNLyWm0AQENSamLcduhXlvOn
3c0rysWOoSwaqe/BN/HlI/cOgJjzhKDkU1JbJWgWb+4w34u2X1CXoIJ9+5tqRQbRtvgCzgunH57X
ImPxdrc8Is2917pjNLBTisuSbCgSPSpyWffWrFuviYEgjK6N+4400+UwNW8z+yjNh87JUfn8M6+b
w6GHTd5Ev7bYeKVK46fvk/Im6K1iU7Z6YF5OgZtxkO+UkkBaozQ9vKs6Jgrg1/6OQwzSngvXGAhu
r7ov83U8yFwbfv1fCJ25J3l227UiMRpp4DyhoyZRsfbqWCLKM7vUpnQiXZ/ghzcL/OkaQe2mDUnu
LE9WXAuV10tTlgVKz4tmd3GHtC264w7hnhnBnxOK3Pr1E7cNwz3C4W8+THZsQb86+bfnoX/PIgRP
+83iN/2XwcYMi8n7Finih7mQZDFybiAokfatIvsjpfseQ2Gw6fKefwaOla2orBDC9pmDFcMP4HA6
B+0NIqLKaQx2iigSNOuQF+7/Sijst895/Lon56qHFtW8Zr9Cu0o+AXKDhc4ASmDGWWrhGV3Hazt7
ZMNLKd3qRtcoGcRJemOJc0xTuB7Ofj3QgaPXauhhBxvYKVZIYURamPE9DA3mfRcYg3dQ2kjb2ZPd
cFqQ984eKI/RUqllVhWQK4BBhIvk6MsyGba1U36yofk+16NZVllZuwbHfA2Gdlw2LnXpW+GwNjEx
KCGdsaYkRgq/P0/tc3V+w4/XjD+UHOFhRlylHiEL83BUREIJYzCzPWeFAiA+1VHWIRZ+GPxgQOp0
/Y6c/3MF3hIEx6VMfq9xTQ1Jh7KhqoFm1om62jD0fy6LI+JihlPqRHjpyea8IjBmH8+FzIoD20uf
gn/33UiEuyYJyLSccAqU3f+LxMPV8vz1BBG69uaEzzMYQEmGHqV9ZwMBy661lGGcBrlvwn7FqqDf
o/IRNiBI6YzTJV7/Gxx8Rsu8UjhK0Cqq2Sash4C+tOiVKaNBan+y6JqBohwwIsWllSIlvwrDUh43
K8xI2qoBguHgtP6XjKaUPpljcqWJLK4WBOI79Tp4YM8SQkMeAKbZZIW/hBkOXC8JxMTPtAuGk1jL
EFbkQ7ChMeCmN71m4JFoicahGCZVJTbDaEC6ZrgFf11uo2h9O3xH2CJASwJV2gOoJ7KDg01NuRhm
c4DQs76TFcIY1tRuS3CNicemlPYZuQ9I5o4lq5K6JeK04l0+blqJI0veD0WscAwCtLKdhCXDydbC
qxBl8iaTdLWjApocgAoNKYOIay2Gar7r1CE47rh3+OEJdpYcdAbsw9P/+JJsPPx7KCTR4LtVASyO
Y5FE3qYljP2XZPlr93c16XbZgvr2I6G5iwrl5no6KEvlG3RaH5NMLpScS/7TpxGNE+eI/o+5xl69
wTzJbExgiaPIwoVtbZd3pIUHCqZ0RFu0GCyB27coYBV+5gOKhIqGMf3V+LMfEcfwhCy9ItH4gp2D
SKUQFJLN8BW41zjOB84SIkKHgSRDtwTxMY6EYBdfFBf86atRxM6/ERPwuQTYac+VyE1V4mdmi8OC
Y2elWoYGf+BBpe5vb5zUJRaCYENUw+4C6xB+nPskclYK3XQb+B1z6VIKGsV8UqrItE+n+NnzuPnH
Oe80vixou5qsxXGqqtWbVcE7zVOHaula2Hn/35e4tXjzzTclxYJXklmNxHUXLwO3FKniIdDucoIY
kiRgKywy9X4mq4ofJ8uK3TUbo+bYYE61aEdB/my/qrpQm6Fynb1IxBbWYDfcifE+uK/+10TmJ3if
F3Z+iNaqgvWsvEiVrTC1l4E6TzcTRmkw+iERtHypAr4B61D3iPssALmnGrAP4krjhOKIu5xpB//l
CehiXGnxNmXHFXOZKVRygn3h5YHhaPWCMFwGqdQvKmMGFABROnAk2J0Oi0Ep/97utIhe6/vw3F6D
BfEn1T+fizjlnObXAUDsIhR2mn2MDr8uqEttA3rOkGUs5osF0ChxpsP+uW/vUKpN7IeFxjXWhP2V
mmwdcgFzlWyTPyUInoGK6fH/VvKXzZhuwUVEOhgQm9gro7BFVxHrWta/Zqs8LlXmD91mjw9KqxnD
FcRXn6vPAWsEhWSPzlksu9s0Cl80IP6LPHVj0ufwuPU8Z+3510vsES3ltiNDIxTxC7jwl75MNU58
/axoUu2wvLmUzZwJ3x+laCE8g3dI64vfjq5gzprfHnuOn4pNLXf6YX8gpOBwon+Rg9/chhN9fb03
IGBgHsTDpVCVIesnAkIuFovpFj9PtUCNu0xG6R9hvFOYhFrA1xBICV2W8YhvP0+CZD4b0h38c4zO
PNM1TCgkTf/z4BbAvycReypK9Z2ApXTuSVzvinGoAZi2YITBh8Pk2dfYeNBgNj/71D1VZNdq4K6H
Yt2yDaQyAcpu836CpW+mBBv2MaUah7WPNIYy1mFo5/U04V5ePBUY1bh6ptBLjK2tEnut8h625N/c
R0WAGxfpBPbEm/bWs8/YjoApAvn+fy7KFj9m96fNSc4k6UwDIYfCOwRaGLRtY2t+vIb13EM7GxMp
OyDnVNUXk/ncV2dCWoyP6vZKGrYaxudCbLsHBF1Q5TQK/ZUwvaY7G9b3TX2UNWoKi+mTF7wozw6S
XgJDYW9ZCU5FjRr0b8VWpmVzqzQ4kkZOV7LN7NXOF7pIM/xxQK0qvtwFpJMnNNmpps1cNm2GVgpH
iwUHddnYwcQErWt2Tf9RGGVx1PskNNuxV2UuZNnJ4wqY2kBfOoo1vpnMbUv4ZuommRX6yZGQXU/b
4bK3cnzJemozJu1/+68vgXYxofhfnHemDlSCB2dwP0kIC/lpZyZGaKQt4woivES/gbppEpB+JyLZ
sAk+COdRDhE6FaPleDDwGqDM/XLpJs5wsEgj5HqT2RK1YZIjuk4rlBTtPkEJ+sf3+/r/wu2EmZUT
ZZpCdAaRsxrcWy1i0U1AKOa4NhdQ8cDGJ9zTPiyY6iSHtlfhgKPI4s7J0DyZSEp6BazM6m6rX/h0
qT2JapX++mZh/56VCG0TH3+3QaeXQ3TRWQZFYbtIlmPfZ8i+61ygVnPbIsQ/8PkvcyuvDfnfI1cV
xTgfie/AtLPUVIOQd5EgBPhhSPKaorEOUhTqAbfcGe/Aofhp39qdOICta+/0uHvP49Uee4dogJpx
96BQsw5CMFqA033gTj1+mNNm/GnMXaMrQWV6/oVGRv03KYzUVD7RE8trAgQvFBixb5k/2y96wHy0
puxxKIe7YFSBvyaYNZXDBYEfiZGN4PDvIJygALayOKjHWN35PCl/79JomiJU4TO2uFT8PFFtBjia
7XFKA5VErljcTnmZp416fzBAqnIe6mpYlg8nig+KwL0mjbaNEFELL9IRxWd4NQb1R8rkXKYt0Xki
E3ARAvEl/7zYHs7dx7xB/qRRN0ec7aKPPD+h/b3KOSADAaj5bPKlSHQB29JvBcFRhWcKT7CXzEFu
1Y4A/YclOWfAqU221TyKXQC58Qg04JjMekV975mF/jLPJO+6nBXeLHlye/oc7fuFgC8PD9sCYqbZ
AUj1NDK+bwI7lt009+dGyakP86Rq5LjPRtjLEbKpio8irrqaxKD7cYOmS7GrM5GoSK5TW2kCvUV2
M1+msR92CIscgMFwshi++HFaZfuAgkolM2l+bBNcYkdiUqr77x3MWV64EhkEE/uDcWiU5ysz4dov
SGM7PaCLfcvbciXZZNnf2GOs3fxY8WdMfuphC593dxd6n4GfXrAC9+mX4R3KsrabKXfi7oeCRL7a
V1zYdwT+kFfZ/p9xrufJxkbW/7OS+HKcKFgERBQlgFCViBeEyyw4A2OOl3fUd1Tv5ht2EKKllBmu
ZDQD16qMohD4wCdo3Hu9RSkKDfzduLhtymrzdD/SAFC7H1DhA7BkRRm9wLO0DNJcCZ/fsiO2BrN/
aD/ehcGCriP9IcGpa/spXFtjQNrtlBU8tiWH4xQf62NuMGjT8ZM/Dk2+PFEh779y21CC1ST8ZODt
bbMADL9w3+/dWSYRBvsP6fDYfZSeJuOc42Behl+J4LqM6Kx+qKkF2ylXASmTry6Du56rR2asySp9
oiw5mfp62ibGVfDiT3Q8zAW66oSKeMpMVO2ObVSSAw0JUt+AUducycL8qPp7pZ432pOXYUoEDeGM
yu6t3vU82aayoCpVUS+lUxBbGGJe3NzD0bVw1DFg+L5sEitBYfb0IRSTaDhQPD7GZMKZ/ATLw0l+
K7rVAfCURmmrnMuzmRlZtuS4f4sUeVdbrkyn8yoZhWXoY0HHT9tr9tXJ0GLopiqAYJOZI0SPf9NI
AFO0bmJYQnHoHGQ2UMpw/ZgJ4b2JIIyZAv49ovzs0NBGnLyE1gVfcfBloHqV6rDDSOC3cm0LtuLi
cQjtIWc073YkUtYnXYr7Wz6ZnKJP+Ua58hlGTpRhaS/wFyiC6DDS6FUZLIiBA9+1ANY4p43kyROE
Rzh7W/8p1j1m78mgMNLLmEYRmdC3I75Beip9Mn6t80d93tfoevnXymDQiRKFX9xhodbbk5j+ZLZO
E2/6JbS5AXLo6jCwv8M4/Cbtsg2ZEZ5hd5+m7VzgubRtyaDd14rwWi+soMWHRo9Z7dxTcmYyOCKD
gDw3lsNJ1D0rl09KxOqtd79N5nh3PK9Xe+dormRHXKA3IbcqwkejpSvH2Y7iO3rfSaW12tpH4MVu
OeMIGVA01YXlUP00iruLMEcNn1mpAMKA0rHKhT4sl3TpGXCZACx9jujIUo2yuovl4piPRNziCaf+
MBLigmOVrQTIx2UfSVyiRVINkRoVnZUx5TYzraE4ecfB2KbVNxt2vMC+8naVhW4e+BTtiMnXZ+E7
vLvIUgoe61bZnmobBsBNp7ZmgV5LwjK1A9mxoQn6gSOVhdS+o06B4mr7Qg62Ac3Maf5nUYukWb52
vPqSpfzw0LtIbMfwEhcU8WG48AxIzPhxB3XCOFmzXqyhhbeIbs26s8dEXtC9T/vtzu6FoPrOUIuP
6cyhNxNh6Y1GWYoHzzLOgVmJ/WWEmY8fKgJsFffNbhkZSzRBLsEx7WT0v/Ty/AIDqTSvvz8ZHS1A
ZRAcIKKkpb3RwiBYXVpV7bDG/GZ40NgVpLZU0wYviF8FqeDamKDWVXNDbrjhSZC8I3ZLzhVAsH0I
AGFmwg5QhPLwPG62gqySqACRO25P2zpBzch9PUvYAt8U4Eu2dAfgp0PWCu0JfLzY/dQ3p0cCrkTX
L711UkGZXZ0tx/sFQ7utao6MBipvBmMxLZ6qCMcKwJQIG0W162zab9MW/eiqYs5GLXX4A1/oC6To
Q+F43Ww8mcVTXG89g+fbDMXswv1FM+mL/8zjWrZN9UaneuFfOU4wl+CORZbEdQO7Mkt+ssAXy7GN
zhiVmoKiBM8mLKx63Ez2cek8nPruhobl0ANVuWYzU7lBuPo2rWOBLcMLKuybS6kgv8lUyjdaFw3W
yE4QXR8MU5oVN0Ljznr+KlSCMruuQHMtI2whYfx2zyxjFwtg63J4eBH6JaTuCNscNXn3pQ1nRYjZ
lEgdjKWLHxx4q+HIyyv29rsSkXoS5PqCNupIfF90ox8TkBs6kmAnpfGcfvrPN+onm38UkKlcyE/V
YOctPk3Grb+Omq6tIsiRBXCQD0Or1bokfGuVwBTMx9mfX8Tx0YRQ9SVmiTC1ahA8KrCv3QXBhjcl
DpCFDjZGTltROBpOErjXAiZrDyCnnHiWDs+v5UQpYafPkNzqAgdP2huN+XGK2QZHVQqnDIe9EaJ9
6+09YYuAAAoEGUfrq0hANFy2BYFYm4WEmBtrnnjw9DNOJVfDgk4LwZjn2b/JCHgFkXUXSZGNhsFk
vNEIgZk7ermN614W13g/DRR7HQS/WtzfNU6BQzK8ydTBw4MtD3bNPM+xiY24tmjXm3zwYZaKOaM0
PtTtDjc9ELO6vGeIHIG6u8lcnVy6muekWlg81G/qnWW/u2ykK5M1RZhYXyvH6+40o79ECX86roPU
m3bC/YPQMW0IvWeMvpLEo1NFXs5q8/nlSYtvd6zFq0W0orqOCHK8uHLOEwzX1UNsZwC4FHknM/x3
keFLv8HfVXwGjZStqvkrCu36cEMJCGJtCYeNWhm+0Q5tGKsD41/rcEwzPiTqve3xDnzbPXrDoWN9
YiPJHotAQYv8ZAFFtVeuds8OhW49Rh0pso45aXGIuEbPD0HmueglwvC9lavf5nDvWP/rXFpixnxi
tUf5G5FRlPQGnB/HJJWpU7HYFkeB3OWoCY4ELDkWLe3ByeXQWvyObcYh1EpCNqgJUfSefCyZ5t1b
UIIvLRz7uYUqN+qaJmDKHFe6lG5L721SCIV6WLi4pTavdCXvNoUvq6tvf+wmetkA0S29Ro+SnCQ6
L83o23VjALBkdY8zAflPeAic1W8/rybD9xsQlGTuAb5gx6sZKUSG+znGnFeJeEUI5mf0E7rTkgKs
Xmt/qGN0op3gm/1011tVj1jGHkrkfEdw+YKzjv7grJvgrj0ww5OcgNFnfUWBY+LJ1LfIOB5n9xAh
tQlYxlslqFCxudgbIVviBqD9pqhT8PguYWryYP2gA7QoLO57VTOj0pWEZZIW/7GEhj0XPXrLzjc8
w2n5ejtH2TxD0Yo/MzS58/zCEZHRDucMUgTuidXGJuICI9jaqKqQ/8/Q+yjHwJIKNWHmgAZSfKiq
1XRKi829geTwfjUqh0ltIk1jCrDq+Xk3U+eGnyyzAYGkegaEPzjpqnHrQNyuenqyab4XAfK/JNIK
YCKg/TkdBADZW+//nUbGe8SpGCRBx2DkGaoA8V9MkjReY2wj6DZqIYYkzIQpNoEDfYMYZSiFqqwu
S7WrOvsKpXnc9AdLdredEowCzrzD4e/B2LIWA/5DOlzGLzbKWCA5WHjRtHJo6rs0wXUm+LUKL4VD
IU8bRZmmOU9qGmlBUBjAEtVxvICYvtv1HRxSFKyIuNewD+INdOwNZ5LuaoI6AlUMtbTkPNvEWOZT
S4a/LCEzvfi/55lcdx91oJ7W7/D0AX+6oSlK7WHSBTL2TrSm9ki30OmCOSotDjT/w0VS4d731ENC
v9uZgQ5W4rVMHUWqScLbFKjfwajSx2Hl31e3+KcuQY1FXYzDXccOqD82vdJ1yMR7XROyZQ9il2Mk
2MkF+c4DsDH2kQej0o62fChJ3j8LKAojm2HIpMxGwnVOFbNcQUWzUnR3GCz7HXxulvgu+h2H1BIL
p8MD311byY5fZQ+3vrlGFV2XAd8RrbkkAth2ankOrJe1TMuco90H0vKbIbj4dk3Gy6tL4sfjJUkK
g5o8AW7/+3F4zwLuqzgGNgR0FNxlgGephVTtU5Sq6JKs7W3MZlf1ZRGacOQkTSYpQ6j6YFBliiJW
a1kuyddNprkqr+U9OLdXjEzH457lGFVmcZAuRV+NKBUWnJ6gH7pT+zPD+GHz9mT1Q9Dd1eDQlkvQ
vU80u6bc0YkkSxCA+5/t8Kr0/iIvjsBg5ROgD1pazJZqD0nv0jYRgAG7NnzN8+0oNx65j4lo8gum
FY7bs+PNB6e5+l3X7I8UM8Zyh/Zg/xDkFNJf+Kso4u7NtVcC4m34j5Q0+lNkuT7gb6vleQbx9Oby
WlqnF4cn9Cd8iVnwBwV7K5Yb/+pJqHRpJKQPL//HpGk2twk2MOQNUjfAWdj/S+ElUrOVE/k8x2lJ
wtMuVplHWJvEfP6futd6QJc6iNR3/Pew5EdVlpeVoAoh0kNwBbWLQuRb4lko+p3fxpZgHC3XGMXM
oKINcojzEtu3I344HGnp2ulCbG6RUiMBz8MgOhVDzmIH7JEsf5dTZFIWTyL516S4UAqIu07bxQpy
FeQHAmsRzF+AtYwfjPfY55bEzGfC0POdS2DGuDkc8bHOHRtz4p7OGsYmN7epxKgkDhHSOhOt4Fhe
SWMsNdP80ehNSVWbgzV3COWTJ5AJb/afc64zjTJPu2pNhxgamjZfix9eW5e6yTMx1FN2o8kmtLjz
QsnVSkK/j4UQ7t03zrUthsjj2Ud3mMdwDBrHOMsxT58f3keaBTTbUGiczr6kHFr7sOCIeKXgTWmh
xZTjxM7gp5dnrrwsRdfnDBB8rhRKgDg6trAjZ/XqkvNqzxfuEXyP6ErkUcnZ7JFXsw6sGgk2UUx9
C5+gsM37TKjne15rvFpaS3MOlIh/Ua3Ur35Zu2xXvUw91ewjjlLf+Fl6On2GSaTkIkX0jyJKGf0E
/LRkPFoQ64FfqP3FAoMiI7Ac7SXj7ajuMZqYlrYk80RMfvFYr216bM68vzkVMq8trhXC8xDvRCk6
2X+fA3eL1CjCl//RJ8UQSDWN+hn87CljxGsePR29YmROrl6bYCrH9eqXQ2E2n4FaCpqXh1WkwiPx
GLgbgEK9kwj1dnWpKBuiXpuoSEylMfJAqtCzNNfmAH9Foje+0XvRzXyZ7ILlDAAegOkJj8zmQobF
jfTf22wITiCpOyKTPhzx2MLksogjUeXX1rCN7MsFAUx67QJecW1V9rSpmDFOkIE5sBsVBy7IYCab
vICK1uU+lzM/oVNo8V2MpiBKGB/qgMwzHQnxciXdAM7F83e7MY6Ss2n8FD4Uqri0NPvAM+a+6wf7
tKkersO3N0dj3zX/gbcDqmd0ZAFd2iQQkbtBGyXgT0bRZ+8bkg+UNVnK27z7dAwjM4eIpte8i1Ex
8HNCZbxWN0SOfpsysxouO6JMnwdBnzKqyOXYqsGDHXeNKWPzOoGpA0T0pbkBQSvldLIN30mIHKKx
lg/OOmOuoMAH8Q+ih48ngaa5UDUe+8wO5rkHNktZioXr2Rkx5+dEB0ONrlQVXqKuLWcmDdOWgKTB
z8+EDv/fCdjbhnFftvA2qOq2xbAoYzeWUTYjRsXUzqVWHle6Gw+neKbw8ItJsDBo6hkZMO4Q2v25
m/rvgVuOC/dyKWHFZxwkzL7gR3ob7Q0bFkry3TaAdcnt1g1nDAw2efrBRDEcNEhc037g7asAEu6H
vq4IZb/AQQTuSzMn4V3GzHPiVXyZyCs0ybTUvQlIoy/TcW6wJh6li+Psa06kwBYCTHZs5aF67c57
uDToVV2olxcyHTE3rWKnBAQ7hU7oInb/ewP0g28l2d4dDI1zcP8B6U8jneLKfkCs9OEZqO7f3e4e
EwwC/OlkNro3dYQ2rXKCGDgrB10SJEldsCsLcIVTe6yRKcrgQEwvMGTnx4o82yU1r0AyE3wVxZxV
V2rUA6nBYdZw450RcxZQLqyR7eeVaSC1rSglX9rYgE2pmdM0eSekhkjnNcd3VJdFEMq5R2bEj63E
9F74O80IeB8nTgaxEleLJGMr1KLrrl2rOgRdN6JQ7AmVoWhmHjLmZSgfV9hgndk7rXuNxg108sW+
uVKiTY+oK6px/+N7U2/Lhu4swxISq81BgE0+aaoxJj8i8AwPRpQA253AcwC6xYKX+WAIp1c12N3q
i9/0it2AftvtIk5ULbv6sT6qWW4Xg7py9i2sZQukT0maBtwylOqYp1L3v2RRsqwyLl/3EXZ6ODJU
Tub3e4Cmx0nSvKpt7G1x0EO1UBBEoBo4HsPtFxY7okVPs3DqPYWA0kbcNFTF299PmUWuuQ+TjXAU
Zx6Q3x0VkthFKJQAr7NYOMyi8GE01ifky7t/s1q/Yeq/LNTZM7EIFVOWPyIyzGD8RJrF14/CSEQj
GtpzWCuKrz4aLYmVEtDd2QZJYHWFz36sc7rHZEZiCkIi9UewXs/efHsg58lxwLjlMqcYQxEoQe94
8jCKx0uvPteS5Hn7asn10MWQ3QBbqBCiJ5XQTDqtT0rSu+5TkBS9fio+kWnvV6erGDZ/fcEf6VAF
P4dsPlXRIpIOq+1pTQ94YaVePvSC+qonrbq1b4v37UWJ49ROMBlhY5oHr85fBbGZ79d4kYeJ7a5g
1VBAD/VDcOuT0KeYHkxgFS6PqMC0oyMYRSZBQ9CQCUMGALJltshjv1h00D4gsONtupUXJ1vuxwHe
inxwQNe3Z8bzU0PEh8pldKK1ua5IAXE9kdsocl4D8LPlewtnOyX55TNOGcRQkCPKBrqW+9c3YnpF
sPgNRtt4e6M1I5YPy5kh7FDfh2MQ3XS1W1bUWkXK+NYaqU0BNQQE4aSYIDv7uEYuy/CDDNGb6LJ5
GbU830UcoPypOwmLYXPAtYIaNLvlJDEvXlKN7qKpyOb9mRIyqqdKeultMr4S111vNjMw7eJhjXXp
BbQhqpCfuaeX+p7lRcr39isPUY9cX95l0it8H1mz3v3ZUvpNqaKo018/w31PGHkXwI5BBaccmyy+
cnqmzioker0+6EfHN2HRkjdwanj5lOCL8/+TvTcEbhn5+RmAPYXoCDsjQRLbTx/jmg817b6H31Am
N6t2+KOTfUeEZqKmSX7qnSr6z9SKitE5em0ACelW3fcnLTjS+D5hBQBVaMFaNkSf1Sb5CORDJam/
f9Z6Y9aHRU3kRybgRkztedAal9xtN2wCigcdDshZz/FuNJtVin1Zthnop5fLS4RlqEkUmRn8DOPc
y7t8WZW4HNBRdCp72gAX/uzy/v+5BRIe/e+ngBg6SQphQbV1hweGE7lgXlG1y753ZaD9QNQLoOUD
VoNhrzlgUCGJJ3YHhX0jSMOAPby7M+bokTo6iAiPxunIDpKIqXYYi6atCnYN7uFbBFCY1fMBol+1
ooO8DfbWiAZrnZvbv21dJQtsv0jzP+W5R9GAmCOnLZbLP47MH7oO3XgYZ8uZ4fYFrfqnzgqs3Mqq
GGsrP8xvR6N9hAlut2T9eiUV1+WmexKMDEsisQ+w8dYauhABuiqHAcAd/TWTcbLDOSLncqu+eFn5
xKjxA4UI/d0fbSYQtShyfFBbat4XHCXl27ErKO+wcX/dWAE0wZVQUkvbHgTaYqql7hpUKLGqtN9q
DFYsh/CtDAlTkQ5HsIH9DbWeQ3Lm7y9loEg6/PbtRVA3SngpFCNYhfWnAWuaz/P+4C/EcoP/nU1t
psgIdJDZXtDtoZIKxM6NGbdKTjNB5bwTbwYNSUAKL28bLzjX9uTNAT8QkheWyczUxOE4J19blPqa
SnPWWp8cl42J2fN4XZDvahdMKri8PbvuE2Gq+xo1nXMyYeQJ0dcVct65/di8U+8XpLrHwhHECpTp
m+3r5gHrEgvOu2rVty5zJxYl9WO6P16sh5eM26BEekU4OOmy9yYfv8D+FPaA5q5uVFFHdoso+plW
M4PO0Zoekm6Z6d6eI0JxMWkiARwMxUd+zNBA90TbPU77lfhmQbtLgOlBfPh3j9exwHboJgSKwCec
lctca0Vqpf1cCLl3Xg4n0APMXFpDYGhHfQOM1HoAAJlKzzfxlR+ooK6DNghS4oQx+vU2LmTE1MrE
H0fcaWhNkUbagRtaL1nVNt6JV9uyxVHKDWvuNYkYex+raZ3vg7nKmy78wJ2tD5lPct59d3isg9Fe
rtdJwxQyvYNMnmp6h3CupaqrtgAvlaW7QKE+kxaRCl0McKaZulN55L1g5VkHIMECvvJVxhbcAMcv
PfrSbJEsVUPilQmlOWvMekcpKuR0rH9fjj8uMPMo1p8EBRFvKOtBl0yqHasKSDDApnzhGkVswzKz
u2ztq/EzhRTdH0F/0fYiEd3/na+XQuBkQ7iSoLwoGgJx3d6omAQm4iJRAA+/165Acz3Tmp56xY1U
VTOfuLY6a9Pt/ZbFEsHXnFl1PsoNIYkobeZrlBBbtMAjzoDZPIPky9MZ6g9k1SLMqmCQSU0Ifi9q
zHWZ0whbOtunY9EA7e9mrtsH7wKKI+V6gwbt2rKWfIfz8Hv9oKGosf/APImYMYv3lCXiVCecPB1W
/VDZRTf4JKa7n9o6gzn5D72RNwI1qNCW7VW6k+CpYmhGDfcDRp0v3JkL5AD8pmO2qRq2luztUMZw
iS4GIfcnkImB5Bsnpk8R803kUJRJSpSq70Ppfad3kCZECV9ypCslTmyhBi+z5uYbQtZ/DSyQNMvY
sMvtMD+b9DS//5c8trax/vq+aTFwUy5rE+cHGSCWWTf7j+wOkAVXM/O1KTx0UJ48LOhmZR5YRuON
hE50SxOFgAFWjjcP4xvo2DS1vWaAMl7j5mvod44RtlxbHG6uJaatvN0WPTjgD0gIkvafIq5NiILI
Da042Ix4bqof66xRXUekPEu8xyACBkj40It8RAXN8ykq1HPWi2ITWsiQtbV5uTjjsiJxINPqm6Vr
q6ePOkI8N7WJOt28ZGNIAfMJZP+0epJfEqckPYNcmyw3siMaKhsrwQOIaFCm84FnYRXgAlqEbLlP
GgR0aoguP2cD56EExdwc6BbPHGMXSmP+dRow8Oxwd4lxSMCXaECMB8x1Szkbm5p9Fq4obN2jhcII
/frq2yBoHg1DmhV2RlX3hGojbZy3ZDQ31fQUSlwqrFjrbkjT0j86z1QIb3Q50cdseK/UXjIdoDha
hyWyp2ASBJ2cYfCtSJPb5s9/ccqYZ4t3CS6ff5gr9SdduTRApvrB+6DUCVO6tVwMJTxyiRviLx2D
0HhJCTFucyzUzhD88VrPfZqko4Iqq74png+OxqH7AYm2JSRURN7iIp5Qqg5toXugNWbLifKeQO/T
r0cy3iHYNHXjxbUCa4l/336Csef2MxfDOVfC7RHRkwFTnp6c6EV6zBlCzbk/YuH0eBjJANkKl1JR
xDElk8kgvIBReVJBEaqd4nerIc78oU0U4Se66yr61mth7m/2NLaVs74+y5fSYc5E3PMicPWPqJ+L
NyAlyeTm/7Oo8bJjJdmT13stVXn0iFHJzjY//cAIpB7cQj3BaPn7ojlQ3ISyNaLgHSKkxVnVkcJt
tOMdEC4+IEZTCS2VdZt9CdIdtgG5wmUvIe7/zSSmpe6T+LKNXQIuFXV61npT/6kBuOhGesXeeits
MTXq0Lc9LxSagMvHDP0zoSa46CwLciXkHaRHEWqGA6AZVHGqJvmsPoViu+csi1FKhjdFyhaqqnF4
XqfaloASqUfLVUxOOb9oMTCnLLKfhlBiaBB2/i964FvKygFGhbXRyU1tcqDFVnt0QIZR/me2nJqm
6UmFd1KcLW2Ffh7M2NnyBDGl8Pn+8ucu6o8ARMPBj1iHDI6iis1Wqm2ACrwy0iYh46nm3jlRweU3
ybEtrixt7x774YmNxpnEt6eTwv0l7orvtmdK+QMAhE3+m8D2niB+Eq35Av5hJbJQLf3IRIlFMhi6
3DfgYktAUNr0ZmMpumjtEyKPHtLRvAWfelzdDeZ49VkIt64pDwQFsHyCrWh8wwhtgeofW6+QOFKw
Eidc0hmkrF1LRBXc+fRo8jGYP9hDZgr01whztS4B+kYGIau+9TwBLRjmaRZl9u/+UtMCwjPD2CqQ
ciVKfb7E3hkc2oqRywANHGQijNDnGb+3xUZPGkrD5mxfj5ulO3SCjcAhbutEcL4X/Agq5a5qxlSO
ICRfUODuZco5Jf0ax/XgJ+UuP5XvgDsPY7pIwAcHHVaK/zcrhusFBLG/7oNRHNobPPAGH1c17fH/
a9YDtDL/tGPkxmFd3zh1f5H8z67VfoHTOSRfw3qkcEv2ordAFgOXKJeOtQu66FL/ryx/mJa4Xio+
1HTNd5OAgB0Ocxoi4qaVPbTlxGJHnthXThj1RbqRdhFOajGxF4d3+MshSpEmhOI0LxpqiYzm72/s
UviMZz9Tc2p6iLfmtBwTCpY3rVoDprjca9C2sbcuL3rUm7j/h5VQDOtwMl23PmymYDp46uvBpp0u
nYWmipSNfk/vuMS+d24fFzNuTQFGmDtnkTw/d5KjwvgJaMj3v7tnwmB1KByIQanxpwoh7Yyi4Ayq
7fs077bSZDtLXz3oEElvyDtglE8i3xNnQfJn83XBhBsXnfaGdTtvQ0+pu0Lh/yHy/B8N6fc7fzAp
pInbfhHkyPhWcf+4itAccZLpwP4U3pQNvWSL3oPdiUbXP4ehhcndqOiiQU3IoJ5knn1SYJ9WBwCw
pY06nLApSzepmHjXHZ6GhhzpbmRTW66PA/ZWcNJyqhlhs1/RhoTqsZAVbjLhzhof6VFVQpM404kN
ZD9W1R1UQNpGWhYI2NqSIeJ940chZvYUMh49tR0NJwfX6jWmHb/uP8hHNOxBmqU1rnET3RQMrz9P
ncnouJ+B6XJD2Wv/A1YL3yngVVKR5lTeMyXCE/4kHx9fpgcgJWthCOl2zJ0kRw50Yg0+71Anaw3f
8OPGdRO0xSD9Sh3Z4ECUZPwaBrSyHK4Tzx3DC2MLVzTR1fOZDnCkdCoFZnaCG5HiK4ZL/G5HtUmU
F6eK56FlGbmRAdOER9+v+2ZJagnFxCUo0vo+1tsPnYaScNYPRsiRCL11hffTVY/dKEjjPs9VSwJD
h7TfmhI3ldfFJZKWcipBzk6SXHZ3PwzABGZPxw0jjcoZsPgrYpJ//Vuze+tBh/Teamd1e9hDn5FV
8IiFVDHZFMQRdi4lFJVMu48hU7ctxejCDA8Ozmwr8VtKjiTOSuYpxZQ/aOYCo91YHjVu8VZGEfh7
RQ/6CyiJWw2U8hFAhyDCuDm2UXIYNPbK7Dpwi921GsNe9oFZd2gy6CYf3zRfKOT2RfnpBriQf5WI
NU1ooKM4FkZiGO/Pl5HD+ynfaeH0mAe6awcWQaqL8Kpr+qUoMoI706ei075Dc0CD5voDt3JrWiyv
TRuedO2JJQoAgzTrUjXfhZoKi1rTHOYbSoam7qVwFDH0W1G/SVxElGeuIFzat00A21ehUmhae5ft
Lz8zh+dKJifQTcwT3hn4GBQ5hysm9Px6SUFjWzxk1PyNvRRd8pFJvPPZz6OT+xsfTJ/ofZMGkRIi
HcBgjnk9lkERL17kND8swom1Z8r9+ZW2tSgQa7gNIJWCWcDQerk5xo2PJvpH9RUfDZL1Ci8fmR5V
uWC1FsFmyZy71oDyEc8U6cXKK3MRTsYS9WchUSiP6gnmc46ajEgssPVb+g4ZJLw4BFxKNtzTA2PO
tmMFtcQ/78dfPuUdtCNlazo4vLDj3nnFmskaxRdejqIOvj3NIAR9i3UchQHxbgWRHmniOszLv9+E
/6JxADwS1dEVt0YEIeUSVd+atf48sX533Nc2oAO883A/0J0RQgsqbLIl03N490SdtgqgMrRatBSJ
EB2wwJVB7zU5S3Lid9inNH1eZqjdDmigDYdsON5a3erDQRzl5EMTkeIrgShf4yRXKHuUKfp+xssG
u1L5+pAky/Q68g6t/q3arQdEbDztF6qgRJg/F6DlacgzzL9Lrbjd/capr6ujDgww7BRqiuh3XeVp
0RhMwrRxon+hwfIyFzUHdn69akEQUSTxGYCN/pu8KKxJGrqWSYH3/+Ga2bAWBPJQ14gGquI8cJLm
iABR/H/csikNKOGN50ryxjG8rYtu7pf4tL1GbL37n/9ZRYr8t5FeKlRZFzEpMM73Z5KFmpjJ0wqh
Mbqu1vU6CG0S1bX0JULE7KTR7K7MxuRfAI34nDwAz3ikoKNhJt1BIi40GChzYvsbibmvqH0RPE5Q
60ir5JmyGh0XtYT/kRbFu60MtYbjr/8RJJJgEx4ThiCDWf3E16206jBODC3PbgvbRGOMEsQXLucd
7zyG8GJeWw8fOpyEduTGFqMfGB0iQEMMOGBazAl06ptdn5sRtYEENHvDmgbztl+T/a+75gMwoDoL
UKI4SCEtFUnEy84rIJkvfOozpjF8fX17qB7R8+HIQRH+105/baQG6ioodxxUtJbvXXkCbdEytvQc
RbLKdR6KMeNT3S4NHCOg9gOmy0Ngs/N6WQSS7CCuKmpezh0DLpkxrJxVFoQrD70wy9NL4a09pDG+
8P8EZ19nMmQ1dm5jt8W96YnXc2o63IXfxSZsflYxr+rGoo+GpZV2uEZNXoOGhS8C9eQWkMD3b32W
wQmcS1oLEpyCiSE3gd4mFlf9VUF2vJDT78kmy5sWrco5SMtMy85xWn7UYy8a4SXe0d4fQaWDmlv1
iDOpzUFcdo2LqyNoXYYpxGFH8rLSkYK6qpMix25LMjmp+LHCBqwWg6smtiIGJF28wYwNlR9Yov2b
DtbImfXhhuKWKQcP0/P6x3Tlay/UTORahXmm2fQErLWlqPUcltSmlkIWaILpsdC7BzQtve+gaP/S
bKOVmh9lDQID3wim7rnVf0VkUJTmTeY+8RV4yNhnhkXNSGW+q1Z6WpNoqLRzKPsLVD6cXrJMFxlr
UH5//uYtQ76J/5Qh+5YmbC9onl1LyYsJEENaF1CzV1BPb/C+Nf5Nx7lwKjh9oGsZIoFK6/U47EJ/
nPzn1VvZbrqZ0nD/4sK+khiA3oJ8NLZbj9EajmeGJXbkClrgYF/L54asWDYMAOTg7wdyFkvBomSi
78JCsvPLDqZ/iKGJQWh4bNxonKoJ/TlAFK5MRNUbL0JPIYUvEbrR3GwBqEoQOxukrFcdOebl+Xck
Nw2Wu20BvnbGeOWYvc2h+vpnl9rQLet7zBJGkAFK8+skmRbLj2wRzRXEZ0rCFAhlUYpaoz+hK2v3
az0KM6CQsKxDMXoMtmECtVk5xtDe4vIva60x38WE2IEChffhP8oqQ+fFBCYrR7ydpO265y463Cip
b1az9r6vqiXB2m8k0I1noBkdem4khM016Q7Oe8KN0ePAqpwQNwgfcDVE45bN6KfCwNY8wbo5jrWr
hODKt38KezXKO8MxGBxwLlphh2CgWvF45Pm9MwtXdwBGY2ZR3pV12daAAH/+p+QcmW7YgCdEYh18
3I+aI2YbxFvteA9Yf7YKLuXXkBvBFiP85t/n1f85XuiLZ8fFKkvSlK3P1H0KJlMJ+rC6wsLDt4Zy
tWCu1W8IeHVNPMavRdCslownLZpQsYu1zrCJxK027ewXyxJClFit3Rjm00TAaMoOpKhoMGUhzOzz
TXPJrQLcdqvbez9bvm1BZbL7v92RNjB/NlDesr8tGFlEn8Cp/sI7+DbUQgvUTCfOKEJfaRMB7bzy
auBYO3ztlB8cP/3sBNH92+LysY1wEbxmfchgIb2J5weR7Ii7jJJ99qHtXurOmw98yPSjYJ/Z6cdH
JyQoiaWrLlKkQ9VSFdCqSO1ZeMuCP0xqOz1gkE+khRMwj7ZJ2Lv1pTAhh3aqoc+fPuLWW+GSWVDJ
Y4z6is55TvsqLqPBP9ollXY+fQNDDjuW/k/gCdJDS3+5olqX8ZjGmZhY2CxLbQeH6XJ3ayd+sJIw
1nlJ3esgwtsLUcIIFDtCI3h6MENA8cgL6mR0iMt27ObpaEi3Np27YtEEZR6lwuzheJ7g2DBA9Bmr
ZZBwAZSDsmX7xSiTNlhpRCc6/R9fiF5XW2JV+scqMaolC5Im7GN9yT5IZ9T4OFBwRFYcK7hQ+gQA
w09hPuQeqxZ1dCCylcv6+MciDSywBxDTTVsuughp7QDU8zAZPyxKMlZ7uGkstBbJQOHlhFz4H1uz
JPbPVJUdopB+/Wsg0jyaqRZZVJZGWp7QRE+eeDIjpI69QIl1wiSlNR9q8S9rSNJyqmS4tuoqwB+z
xadkLmSzOSsSmvWaPxPJsguQGtUW0SqxQ2NKrkWJNcJUdz1i+BrvA1lCTaevvwmHC1e6u5IOiriH
sWm6bqzX3143W4sL/Mxl9rYq3XREMo+XQZjPIiVPSCmVpqp2+DxdRRw1zXelcGJO2XKJm6F2PoxY
fb05EpbeRhgkH2t1U2YbtEfnLYD4tZ7aGQRzd46EFXfcAX/4fFeImn6lekrWGJxQ4l4GaUO3ff83
1cX3htTmvAMvwrQdRHOHF67bHjj8tONKgSdnVN1VuxPzLKmjZ21rhzYaHYZtiylWIwbCploT3agg
NFJbCS7A8ivPZ+pKY13MdBJ6ESVFOve/hMivA3RG1pshuiOuOh+m1TE0+/FSboXcN5JCgPFjjooK
7MX7EpHCQlCf/slr1NYt5qfZ4Pt4WYy1sFuU34Gci7zUmwxN39bOcI/rymxztva2osJWElmp72fm
3SSywS31IGBDu1nDrehKHknncOZsO4oxRCSNFL5860AYTt2bdcAwuBY0btlpRWT5ZkaJ1ZziwCJU
WwL97jyHe3g2ImI2JdGvPCNkkd9l8X6aWM/FE4o6o7Z2CWlcD9sIlmszLBgTGUYFK7G2vJjBxSgd
IrbyumQPBE2GIyYbOP09izT/XpKrUf5dzmDXRtOQNtxO5kEYzCtmqRdMaDhu5P2qIe2xTm7nCeTj
7JBiADDbCXERVDTCWHpF2FuRYhPoGD7sbN+vHbrP2ri9znArTUN+vzldkW4KTqUMIr67oBjyFs9V
RRW+T0NUKEUfRF3OJZonhtESpKHxguXV0pZ6ul3ozz6BezshDUO9K1JXxHDBLUtnhI1nPdmwdlhc
hX3Q9Asi8KVE+li0g1TBad6me7465xXyp57XQyk1BZUKabJlta6HTlEJz9dtWKUh/bdiB3DandzA
NDdZDDgm6zcUMPW9cM/2ab5LwxCJjHv+WkBvn6JRZhUVhHyu+Ywq5JuDNGYUWvtaHDN6nI+vX5Us
YpiIRg7JQNA1RMXOnNReEHO0CFi5JYZqAn0eSRpj1f7zvhmuVYUU6m6EGPHCdW+Mf18mQFDMICWE
xMeV9aoRwvgbqVvH+PCJ3+TZxdjhSeib+/VkqMe8Zxoju78ULmprGGlA7Cb3PRsILPxpYaNikM37
CJFrdDNjcifWN5nD0QjGpl7cIRuFYNpg52xFQ0MNSkgCY/VC4oJy9r0cvojoJ5zQtlX3dL9Y/RIF
Z1vRaBTTqlTirRBSZikzSveSwLc7Lsli+WXQ8LHPd+7qLNf/vIpafrmCNxSshjGPhg2PA1/zA02H
ET4uC08WchNUEwlD/wAGM1hvOV1aexg7hwFdqRJBq3rp3Jlnzz20G+pgC0uU14+fWkmxPtfzow7e
vlb/IPQzL9RvM9L8cuAvV4bwRud/661KB44t9Z2fUZLNvyArEKjTegvyTZVqjdnQiwXCIOhME2oo
0e/DpZ+q84vw532HZy6n305vMO4Zjwv6s5XajG0X1j+H+9tWFSAUNvazcULtzoqYey3GQZiWD3WJ
SsUyEqnON+hy0QcF2C6LypSnrfo3s6sYIU+GfambsnC5QUPXMH7HIxhYOCwnWbULK62AZEtwmi6+
R2CeTFyP5ZJQii5NpkyIF+f9pORZP5uPWe3WfN4C90OFoYNjffvjEVt83dJ+ClSC1/xtYqY2YAfq
Gx/KP4M84AcKwbsj1FJxh07NgxJMiREpVXl+QJklsfCvli6uEl75v35vdiJQK/y4UAhqZoHlIofS
bkGBIob4fz0xWMT/f3LF+0qQD4gzr44nqZwkwGksup/WMMyz5Ob5JmKestMWQOaMyjSEHGteFXHN
JKvBJrQ28wPPtEkX/V07U7TjFu7TM7cLDfdURmAiibLREZCNvmtuSi1w0W4pyY0CtlXkh+iff8z1
I8P4F4g3gLaSAzWSSP66W0tPt/zqwC34HHuCZzTZlGEcJAzYlK7Na9cSuB3jIkfh/yOlIjJfce5P
60jzrwon9vKdAKsraN7qoh2Bnoe8TO71g2MuPB79KIdUg2Gx9hnYcx4ostU9NuuKgtedoeBbhtbl
x8qtE8+t8qnC10iVNAqsTtifYQi+6oCaXZ6k+XtXK6QyPsR91NhUuK0pMiwZzh5cAUa/FrDk6Ryb
wu6VR8VgyhdQ4eVXt1lyV6dC7bp0MLOaM+w3J2J2LKGEMbd4PTH9Qwtl4jEGKZtQPSHhXH8gNKYp
4ML6vg++uAy25eyvs95PqJEpfOFTslqyrIGF19WD2le4Ta1EyminGQ0aNbcKxKufBZwHjSjtDyec
OvEwJI1beWvrFNDQaMfF7Zpc9/J2EDRUz3ub6hNbFQiW04cPGdW0o6t1HbTbEoCc0Ty9Iuar0n2X
UVyShEiKpf7Wk+x2GcBIhJWts0SgkO8v2jRxzRAjIz4QRGC8oitFRIvqk8rnDwI0gHyQcxn/PZy6
bGXxb9ALRyIOYpc6zbApLuFu4VPTN81wDfGC+U+hGQye0R9lT8tlv+zpzDZepEMOxV18Y/QpGIwX
sx1AH44w/wBR/8bDgxMI3Qu05IaEZOfAg8prjfNYh66CbPoSOA2b0BDxl1e6ItgIkrpxG5lGPFv/
LnryzBxI69KpBGpZJ5UbLcUJogyH8UOAbJ+VtgHxQagVN0cI/OCK0Ch6/Nqhbh3x9DlIff0SyTcR
8kMeNWNohY5zE1gDTLANQzBPxLIJsZflbjQQAuLA8a2CSFoY4+bXw542EtVJSQutRahcFowioTfY
gZNoOPC4/upcum7bY9BudtIyq13XljhO9oGLXbCia/19Hcsq4Mq352pGG0/dTo7RJjfMiBtZjnzG
gNLR+QE19z3Yh2dwbuhtFeiSeVZ2LbyXmeUqNzFqtizdoMSfDgHuLd2dVly4ZMJk0XGDBKaeKHjZ
WCJkLs5jf7TSMWYJ+isaTHas8usap/2pq0UIw8WotNmAo1mD4ltQk2q/Ru3Ce6u9986m9EFFsPIQ
pHkIHWaiu90rNmTcGAKy9Bteoz/TQPPXq6zlGUkgjlcVnsgAjBOmfj9gz14eY7YE+pVYAtXqxfE8
KJJRGRBM7ML/yn45pS7XWjGqMwRLyVirMkbYLa2+JFjjovk5QGASSMLWIZrrD6nOAiAOHETw8UPX
sxFcGwBM0H9TJGHj4vUz2ZHMw0NJbaBa3K0zprUsMP2jahpe/zhrJcJH6O+E7l9pQ4U1qZNA4lUd
83EVj2DorkluiwQUDy3uxEmGQypaHRYV5YuUkFekLeShErZR8Fhtt2TuQW+0SM4SpbHUpYPNfbTz
e0SkgCdruvOZnSglxq4ibvteWCbxWjIycIP3w13mUIrBVuZhmm2xCpMzPANwuvWBQ6O43efMkPfU
U3+yRIdY/wMrjDr5L/d8vXPcLgy6TkbWG59PDTjBHY9YCT1Jqg96WHWXuHNgTmbR9E78Bc/y1fig
jg8lO78egyGZF/eBh9XDCKcyx5kfRLX7p66pBXkmWhnW/CN0HoY0IkpucSwuIOfq3LdrbRlat98E
DDhJPn6ls0ST2Zh4nRz6tvwCwuGFnVhnWs1pST882wf6zdiVx1Z3de8WKha8fO7hbrJ4L92QjAw0
kIWLKtY23QBqYPK61fjkIA5xJ4kLCOdmOnksprjxbq3OV5jYItM67dEKLTGZ4SrNeOFcjvoThp7W
MPsdPs7NynGz2a2Si+HKilyhhGvjrwmx9g326rrqHTk0hb3QCsntyC+B9WdgqRApgbkXyGgVm3g4
lZMEzuGgE3x7lCtdI7kJyXh86suydSptDTh+9HRHR2NzfhBV7UEG6Ne5UY/X6T9NxlogZEcFPG+4
N62+7HwLVsHR8357G4Bk+JRCU8G/Es86GQK4J4bZiikTNCsgM07fzf1qktuCnDbFHVgQgb2aGHLR
Rki/uv3OpNW37XpeswO6cBQDuUMgzw+q7SO5FdF7H2950DNvLjzsknhPrLarNI03DCBQQBQcoDwG
gmfmt0zI3CrMcjldg3YcrHk1GouyT92WBEXuIlF4hP7xyOCxAL4r9PKRvlf3Fh1+BQfNBRth/h5F
4C90ET6QqcgpOeC8zgyXGaJ9EsUMVN9Z+pZWD0B+Bkdv75nn+wwCTUu1AFvc4GGCCGQvUWmfhMlp
RkIimYaF+uVbTRQnVXLtvacoepl0Wn5db025lb4Sww5QIFDa5rwegMDlPQsACRJziRACz8fOZJMZ
puiEuKIumdqd6VwJ+Nja4JPw37PftYkzlrLEcDalBn3/QZEBG9WV4Mi6xXAxA83CuR7Grdrzr/P3
+8zS1aIBTe2eEdLPRS8cup5iqAjSPjGqRTCBvy6At9v9vDP6Lsdjf2CtVVtkZSaGPYw7z43BVxxf
ciP9TeouaDaSIKQtFjV/AH+Mb5qrhTSwTgGC+KF+f0NuzVr+JBrlr5kIjvU5Nej5XQfzZadkRPl/
zh/N/z3d1D94W0C4JlqkwqoNJprJSF2z3gSXwkcwv8gwFhZVC7QsBX0TYpMWidIa82v2uHxVLOUe
odkuQgHPTQAwq4nBGEiU3IOk46esR0AU3+2RMHCaJmjTw1ns45LGrBHBbtABIJmiyimqmPYxNUwo
E0lwAfB5Gjq2aRb4B/z2RW10w4e0jqiXWGcCOMBMusFI9s3YAp506IhFw8in4EHw64XcrJ1Ku5mz
W/nwumdKwM/TQwL580Mb+0mJXxIt/0KH6a9WGxoKemMyw+/16EmpyoVBB3cY46ACgJgGwipcE/0H
B4+6QVmNqTnELpEH5/sTCCfSwmd1Wq5wjEbe+lLpG6nl49s9mAXHRlK94XKLZayC407KyPPh4mKC
UtQHwcqZWiRnK8/OaEuF3hJqONZAVj6zeeGbDo5QUGBA6wXQAPROMg8bX2XYgbeQg+eL/eEVBQxr
eH5ySV61RTRaNiDaT9SvdtgE4JBVZ/3SFd9MdpU/DZsOZeEdog6P4IsGOGAFhC+TgtB93y6gMw8n
n1iU1P/ZDtA5Y7FsMK50RYhE1JXe4gvCNRVxtKa0tz2EX/w8ix9AD4BCYAPCzztYtC2+YGK9XNf6
mnZE+spmmmG2SJeHl70EqQjvBb+RFTEuEplVN6bRL1dgsSmmGzxqxUYX8H0qOgN4EYONmPHzSVgN
lib2WcKOmSNmamnSzC0HmhWX8Tk3bae7x7V8uOrKyyCIvVFoBxqx/yCI/0AX22GP3vvZ04DeWkDy
9z5+4e4d7QPJ0ebAssRsCKtkmyy3iyr9GbeLR14E3mnjmcq3HBmtaNxlHjKdNARj6g7BnkUj1GoR
TXhW+y5T+VqJ6Oy2KNQk9WJI01VxBRYhdlGkXIRGwFjV6GNo+mIfa4di1omjgYGvy1EHVHC0QkMC
DnKFHySHlRKQ2YUGSdeD/n0JO/njty3xBhkZUAbVUECvKC9hm+DjcVpTq62QoxAwbkHWjGcQPsAc
7JnCzhPNLthlWFEempDA2BP+MWJC8AuTPQ9jkKN2/o+6QVtX2rQbooVJ9quHW2ZLdCJuh93T33oQ
YC319YwKJQAnyUzY5jrON0H2ebdrtI5CLN5xrUqsijSUw3u0Gv/lqj9PKN3aJ1Rn4gNPt1XDlkem
INx/AQk8UUsTjXGOrXv6Zx1wHhTnyZ/BMG742E9H8MmUbwnu3pPsDSEvr89nRTNsnenlP35SHHB8
/TGjOSrAbyhqU8XI36SK6LMckuGULkMRjmgrzmcN6hxBbxk/q2R3Bug3ur28fDXJJzpBXaGBUeSb
uadoUmeDB8DGQGAf67VuwhlvO5YceAdNQg5QShho+6XZBbJLJF1n2RKhSIU/QkRE4l9bmTXp/J2v
LgEJ8ED5jdMIVKy2D2y1CQ3ISafdNBjHQEIcnXttiHJMMNMHUjgKkd/SeCutSenMuS3SW3AIByFs
3aYmvZ6apZ+s3d9aHW34uWLAQQWZGdboAL8a497hgCWgTZJmp0hnAsYQ8hQNQ+8pLb3FYQP7Egs3
N1vrz97hZfujlkwPT6sctERv4Z37nRPSjNYqw58dig7hIxqR6cbJq/YoQP7/PJ3A40Lli45AVrmQ
rA+qnNO+Xsq0oHTJNAcbuudFAPuU/w3gtFRe3XklXBrzlm0VeEd+P76/X1rWOGwMJEgP9YVmb5aS
JCDt97aJXbvPxNWu8BuWnysjAU5hhYSeftJWTTRB6EfgHxlincwpe9EOaJvSW4zmESzBVBuOujlw
A5vvHLCOMYHOO9cGO4karLFNLhEk40zS1zIUj+klA6866SgAZd/zXYs8swZIZuosENOeF6ea9Wrn
l/J9Ls5kIrp25eLu+159pdiBFwnGPjhKkmG2GQSsxde4FT67HL2IIliecEQ4kWmYVEoesSVuxYUa
pQhb5DPewLRcOHWj2xLk96AYeEf/h59tylzmFmccXpkaeKZf8Va8a1PtBuiluT0qheO2tdBf3qte
6QE4S47fsWqDNHjPxCnDAwSwxIc9XBQ2bbd4/fgEfwYUlqxyTWjA36cb54GsMiMyayWyp5fLiHJM
WVFavYRGQ/lG9WvApHh6gzqfUqsOFi9BRsJKR14DGeOD1Dms0DE6Ln1gWn9j0nFE5sFsmojL/Zwh
Uw3v01DmOcHp/Rb1vVncbJPfzDUKOI6VAxCtUzomZeUVQzZvcCREC+5bL8s9nUr3aIOATal/Jncy
AjejAjN0NrfigdCshWrj5uBejxs+gbNhpuKv/tMxHo7ZNWotiETkQqx9vWSKA954p6KSkb1hK56p
3LTqZO3VhA20W0XAtxIOeGqbMK51eGElnau5OUocy4pNMyfnlwvcTORiu6322qpqtBXVqy7rOpFE
KodalNdjEMPJ527v64tfoGNsuWZeO6LzXQpfa/KL1JMil/Bvg5r0UZCQAUb4ZOExtPGG6wuD1cql
9XVemfF77J462yo/j+XigSSW0erzrQzgCHprg13WR4DOo7K6SH28gDP6xHiL12yA7ScJEAWsUGBu
WS/uLV62mLCzTebCLrfNEHVMvbHaTi8KhIzRiNWBn/XRR90MCe1naPqI3WwDmkFJ88QzXJwyMCZB
7S9cFmEDSTGGp5OO+BXSXfpzTsXezN8MVoQ1jVL6aVplu1AZgV0WBWRr1CBwZtKlxK5XNtwkRYqI
jkvlKfol6AOiF1+sR/qDQ9x6wRNyAWiDLK9nL4sMiRbYGHSaQ61Lq3ryQq5Kzo0DbwtajIhirutk
peU2RdXAJgCpUJGVOMJBbhUhjttiHilqKT/JPPw3SP8msXVt19CxuUtMxVB94hnRN26zlPp7VeS2
R/RDMOYDwkn9I/MuDGWS6m35d92p50u8Lmuctr2f2yPDlX8MZ0ESY/sYaonDPX2y6VJWfx9Y7Ebx
ejqhC9jbx2Eg7lGEGyd3CjfmuvyTN6oxwDmpm2wUNP/zxQctdzqgw/QqA/BhDh3DYw5M2Zmtg/Tf
uOiXpdBqmc65LGDOwG267gEjdF02vnnIAJak2tAT5GgV3ZdtsL9vODFlRXHitVviswGSYUnMXeiU
RklZ1yQ+RJm6ElrXpVXHFWTurz+QisaSZlHPSZkl3VePnaJOFZ5Kp6xZiNSK41WQSYR373uwQM6I
UQlYIj9ju01kgOcvlesqD7FjthceYK/4cSMNLv0OPeBeXvkRV/2tamGg5TxOi+ZwHnO6pfxoPWfa
RdZUnNBmoKl6tlFavvyaoRbrY/7EdfKeq2LTMVST8CjvIyRYa50z1jhhmJzefJyzo2Rm99jEG9YG
54qXe0ab4dZZVawQHg/izg9e6BWsPnLj87psOBWowXutTvdV1OVmfTT8inunK26k5vMG99Mw6dFE
/6fDukSsAzonf6gfuIlTlIF87ZK9VgwNa8WYLUFDA99OEW8ysv65tPGYzMIJ0KPptU1P75EkbpTc
5l4+znn6VE/7KdhEE29s/7LH23wyfY6jKzYfq0WyEZQKRW8CS4QPRydd88CZDAT8XngTTlDvTdsS
5i5bmpB88MUZh+PIvS8Q1V8+MMvDNZ6TptYmbt343mroSRV70Tm9KLEQhyaMcuL76CDvyf5G1rBF
cRjkCdTiEKsIvHuEcR3zYy1Ga7hroD8pb/lVDAqBHamH8EuXJnlbr7btY0HNHjhTGfXWfPoQodWu
bzS+HIT50KTdFCHimBNadJrpScJpdQKtTVuqPkGkJEdzCFhuZOSG1ttM1FG+wd0IYpkUeSk/bf1d
fLZbXzOY8VkWfooyWXsxICzPC4sFqloeerKhH/ZqJ+jfQYKurPVgSrlLyk2l6v5XpYoMtwgXSvE5
Fy1KVihtrclhiB/l0GRRYLqz8xtq2nNmk/GKZeOMQvGZ2gNEFHYv+BbIKzSo0nylXHc8L+ivYrJz
TZlXQqY3T4BpxKsJIGtmtfxoSe6N2xybrC12ui5K3yxyjBzWoZ73OIQ66ghyg8qQfa8faom5xrUE
2NobqNHwQnfAPDth+LfZMJaaWR7YVI8MbyHjbTUXywu+eY8NrKE/xJYCUK8fWnymOFNiudeDwknc
W147l98bkdp67vo0CaHv5oyIvTZ3tvasovI4cmau3ZQ4GB6qoLxbkTdKYcLCiQ5BuRPNKvqz1mFD
gHe3lLRSlHmYJEVxFL3fgWpD1jdKvmgHIYrAJ6dN2gJTVOP4IA17Oy/UJau1K1A+VfQfRRLXVy44
WZfd23JJh03OEz6YRcbJ8FKLywQKm9qSPRpRhIW0L39mjpj1rsSz81IShndXfuVkCeUfBUy2+pjJ
C8KdzppRFjh79eMjtDHSFAR3Q+cVpJE+PJZmc/HjOKRV2cbCbP1xVPoGzblQy9pDE1hEkcUMVUdG
83Gn/jw0kLCrgOHvUG44dWyIl4/of1HsU/Nis7HwJJ9AkfLWOLJvkkRPWOkPhuVq3DkuBBu22IIG
9Jm3lDKMu98RLIYtEVb8rglH7F6zs2hEINljN5FohpTpmc3xhlB3Xn0Mr4OQ4b5ZhBif3rVBCWzj
1AqINLh8EtyoJWGZ8KZouGEt9fZtDvsBR7H7crywXhgqq1jVvPjoT4gX2Rz9GqrnCnELQLKz/DUl
ACfJrUoevk/Pht7jMLTrzg08Fa22JFtfuP2ezh/Dfgdl5mH7Yw7Nu+tIsSWWEC4Xvwr4fwE8ACjm
reJxGIkIQOLFIqhha6rzvQmqdmL8hGLsGfoCCk4L/fRb59LAmqXKpcFwONUFLByRgtDs1RNe1LVy
QuHfkjM4vBuQnF3QM1/kwriXFN/Gw/t4383IhGF8vON45TaaK+q4pK4z/wpelpo79ls1yNyE0djI
GrYqRzJYkvaHT1Cs0N9IBdOQ+p0MFwCXnNIBoAdRc+M9DRO16rsIjkMZ84D1Vm5XQfSmypAHj736
VgdAF4hiwMm5eMJe3OEZOMYlWLuf+KsDx9tDnoEzzWsiPQfdYCuybOKAvJMaDKogcZ8MjegUnVqu
iONYVZvAB02AxGjQ/Se9sfn1N2b0SDbtuXJnjTkgskjT7lVI1+3BPp3aHLIUEr4YsWDG2OMIc51N
BotSJsaF4QvicionmCT8vQhqMn/e/q62+nlMLetYp7ZWA9OuthGTPsRnx/lL5ammmEWtRNjbuSUa
bzELROJPhx5RTJXLqOrdS7Wx29RPlSiC3qcIcq/v4oa61oMCxy5/zFGRmN0I/ZZD0TaZZcrUurE0
w4oAkatwLESg8/MHCHE7UV4lTMckyeCkXaAnfwnUKHUxbt5CGQqklfB7QI3INHI6lQYbe4ZybuQW
pU8lMDStiIJ0k2ZexvJc5Ck7FV9KUcNhYCrtfXgyBkDvN7VULuWzX8s6NkmPhpcgKJiaOmXlry1l
Uu4iyHdySH13m9KTUvR8Txl3pQpUzWsW0OSLTCTsjHvH2RBLvAHxsipVZC8vDTq70yWC0EmXfBo5
kuEl+/OgXwBNc7y9v/rvFnkJLlX8nWv4ZowKokb/oGKuQ1UmiNC1oAYLiJJCjwaJP+5473wo3lwU
uMRbnsNGD+H9wRpNr2JQlBCy/9oZhhGLNmTuPpeEbNc7eiqaubpMfNn7kinH4yV3DHFN5DwQxCTK
7/kiELbkcTmd6AMtlxpEpZgiBo+nhiEEGrFq76KPrhU5TmdtQu1BwsDBT6AP8hp2neRV57WUr/7T
LYeP9Z3wu8UNxVf5OpnD0uvuwL1+/nV3OcNkL9QBNvfQcLOPozPuYTD27ADB1d3UI3XKpgihEuUa
wnOlGNLetMrNI4XjygUGSC5Ai3OXsiIW7XZrUdtSOb3xdY6o5opocn9o/b/hckMYaR8DYPL3OzsQ
Z/XKt13Wy+j9oqiBfCVPEH/DrAQl/a5tU6LuYX/bM8LqlDfOtwDN8q7szBIGyN+wEizjmCh/YsVX
PHOp70wWyHZM9Piq60WdDjd0sNtMJU1k5QC3wtl71TB8Vm7QhVQC6Q04L4tDm86/nk88sP1xGCme
j0U6n0gLJCja4jKXSIs6vPJHdXJlcjUcaRmgJ0nXrCs/yU48ARAmyr81nr/ekD0DuRjCR1MWDCzo
Fqo7wvGe9fXG744/kNn0Xhxb/9SAGvbEpyIvEVgP0DWD2jrDR75SqlUxPIlZtJtmOmN+SDqs62Wa
ZjbhxzOmoMp6rMZ1gwxrKiUo2xdBJgAmAOxaUsrdPMgMLk5DOY3tO0Jh2m2Xwuwx/aG6G7wrjp+H
7paRLayZOkKWYqHn2IjJf46gxchve763FgrfizTGqtMVoGsJW+n+/VztW4OpkaM5CCz4jBKsPN6Z
3UYaDh3Qsa7D+HYW08PBjPiFgo46n04/MtTtJfXvM/zzOoQWFHUdLhJjcON/G2oQ5cSZlaYR4GSW
UJl28rpl7edm4VA60B8PWAabx3gSS2mxAOgwQ62GAGgeHyJZLVvQYBheuxwfTLAe4aoKPg1xz2mN
+kDuPnCeAZ+d0L8lb9dtQl4/931GpFuK/KrMGWfyAD6eP+YF1+WL8m31eh73tEo6qKcuerDZQoWK
HsEhwWIY/e5qNXyybc7oUBJ2IrNpm4jCV565Uq9VcRuDx+skV6msYh9vXSn3sE2vTtRo8xYXg+B9
qVVWKLQmVHqsERPgBhhgccvcF5x30ZVqOgoPyr40Qa7/ZhgABgsksS7VuWns6UlJge7vIWhO87Rp
ynlRr8m8tuNsPW1T1+dM2jpXoXJMYttXLV4Jx0l/O/t0XNb2Avum3jkSjcfjmjWWUL54mUG1ExMo
92qN3XLQ9tve/rSoFKKGjz4pdiEQV8sLYGvBwHP0G4lLtitNSgfHtWQ8K4XD6BpaQoi/GXSPH4h2
AQWbR/9ZvYdRDTQwXRF9B5JRU13YjOVNQmqixI/2kr7bJZeohCgCktJg2xQRDHLJBsgMYTEu69NQ
GCFXElHRAdKrEH/aD2Vd9OW2u6n7EyJMDM5lDWi6j68pB9eX81ywFCyuWg7laOxFivKLaafY/dLJ
0IhyCbeGUY7sxqpFjYP19LtvNbDM2g2GBxFemMSbyaY4MRxekYNRC3QI04A9xhArByy7lQnGEusm
Z7DP/X4DRUyiQCi/dsWZ8bBmSCKvkqrWe1+p4jUhG8S9qJhuVRjECI4F2UisrYHh8R07niZiz8dW
X4Y7viwEBM8jMoCuXS26ZJCxIwl3cwgmEKstyGegaPkYxK6cy/BOTFGtatxgSLhLl9ZZWBEkgKO8
YOt1ewkL/CWSDWkCefun7AFS7jpEwjqQHXei6PqJbSfYTqSjeL0TDu+ArjJ6pjTBn/f3yAl/bqWm
uAHnq8ZobuG31CwIcs3NTt9klmO8PpECOnOdBVdJCyJyH5XiWmjM0/Qz6VZmBBVyZx/E4d6GY1kL
tpg2R8V1irfCqEXb9ZF+jIXkTsdSLwYFPA07Q4VZYPCogMN+oYNxRF8/nxJMImQp8XGg1+WHp++4
85Ajdf8PoZOTNCm9+70cS/C70cJGZKOiZIuzdKG6Gwe8i3clFE23PWGH4IuZGej29Fn9K4gWyKmD
cvwAbcNqKf8B8SXf8kPIIeM8FoxxAcUdLcggfbjTp1vvWw9eHYxMzAJWVBKRwApaWFr6IxfvyBVR
xG2/ROpeVNKXipseMJF/CzX6/E6ilgr3YqPAynj/T1Cg7+z2aAKkXAeSmiZ1CKdQhjHQ3NtWqbmr
g/0moGoG3yE3fLLKtxk7VOAYyNXiE3KDcEmXOMaOBC16SSaNMnPcj/tpWwHoG+sp9w/7TPCvyztf
n7e2vXcWeNLdqUCEyl8GcqGiHUZgsU7GbeRR8d5yx5x9HkbZ/MSGmOGWEMpX/dAPcc2jGhlMgdFA
8akvV/tzmWzBSflwFb6xOfkZ1HHLjKcpdWdkL/92akBNi1FSTiUyXk1ya5SkrW7R+7h882PsRWZF
78dqIFKjTh1AS80Xk/o7awRHpOmIcc0MfmBDXTK+MCd/m19NuGBkcss/uVBu7xToiTkXdBCV/6RW
7I74EctJL3eg+yRDjjy2F+f6xxcez+wIbjb5VpX+blof0lEVIG3q73zreBMPjdW1Enl1F98rNHwO
3Eojiwr73LUbTpekMBQf/DmGliQlOmBAwte8rG+8cwJjFoFOj/KfWd+a7Zpsw+Gw6JknQNAQxoLe
VGIXvDlXM7yy8mw/X+sYdpq8LjJVZi9/KZwWlCHF3OZa8w3DXuDhWl2bNOQa1IIl5V8ee2+26PoX
sewX1beVWn1LMBBdpRFotLxcfprPHCDOxuaDzu013FQiDab3wWRwRG5DxYnwVmwz5dJVxeVtSiRW
Bbz9QLmnAx1pxRzbjEMTxfsKkJM2ofV54W0F1O2nSbGTOggv8QAqMtuUoNkctiKj/la1FdJhxOTI
fGUzxvf/bK7oyKSYuvRNGU1pPBnGHdl58PDhU1kjloDCyhSeAzlSaRCXShGAfVO8X1wgY8Hnad0T
g6Qfvk+34t6FZlD3hOfolmdKgkwZU5aDiT4PdRRk19CdApdcY1r09ZbdUbhIV7eOK5Gw2bkX11Sd
+ck9VA95S0pdgtQ/ucYUo9To/s4P+roq8T8UhgZ5UWqMcCoZdJiBA93sfaMeg28u6fZ/+ZT74nir
PHbeLBB2ULLccktJrbFspxTT7Vx7eWYUM2/E9hqtnazeF5Vqi4CVsDO1d/g8I49WW/68MSZv6DAQ
533VuEJNwqL1Jvkm84uceaE+iW201x6P0tjyyzfouWsVId8eIQt+ppg5cKdsD45W0UPOWFwty1jg
hq5KuT29ndXHPUKaDDVtrKDxa86II1rDEhtQduxZXwqlXeSj8sc98g6ebs08vCFtP0oce6eLlzgB
GZNAtkg8AFiAqPVT1jMiMNCkLUtrnWlKLRgHEbUC+qY0VhZUZLK0ATXy6r9ELYithEImCVUWYnY4
/fARRFGrcAxxMFkiDgw0vTYdBBMauETNd+h1J1+XChP6V0z+fwyHwBqlUpPwk10ckGdTIWGri3Qc
gZcwPrDZojsMlFfL6Dw4gxd+2OoJTyNgiJUZ8IJVJj+O8vWrEoaNWcsh97NN0aBcG2B+QHRqmRwh
lTyDgpvsC96IlMBkeZs8tFCKNE4b7ow+ea3X+9jPpWyxe7DwQ5NCZD84/t72uu4plxp0Wkbha8Va
gNzsZRK0m5yArzTj/iqY6zMkZgUInrCt7Q0JY0K8WiKDtWjk0V4iwfaBuLhircnpmDC3r1nlUETg
JN9J+85w3DLcyVLP+dOtWvyFvQqHoAK9lNMMcq2Z4XLiCCCMtGWVNbbwemYk0e8KlOMwuXKHFysp
wxa2fHFOzrHeY74pJGm7/0W5dFw0REkWJSrz0DMBw+grWKwX2W3NiacGJ6lIe8zjVOApzvsJJAJp
DHDgpxTSL/8nOtYuHgw08/h2wm1/bczE2IUw3z1AKgoB8B2/gaOfCDYBXYpJu/JgTvOSeS9+gbkq
XJ0ihJqF19/nE6GcE0C6Po6FsSbq9QDsddJWqPZ9Hb8rysSvXQiFU+8zAf0I01D3wsDRy9Pvq3lR
4K1XrSNTrv/6RQPnkUOT89WYX1MkGUJ4/CRjfy0tPtIHVlxKElkxOwLMIes9Dilqpdpic9I0OigS
RhVBWAQWlHAPhstJlqTzqZUleVmZRIGgau8ADHDF+famAo8f6ln6MalgrriDg/Yd/UuApTPP3n9Y
hwRQrT8NmTo2yYC26sFkpaR9Fgm0+W5RZ/tgGgb8HgHfGDX9fw6x2ZRNKBKCTUcS4FaPDuhQAUAE
li484IJV8ca3lZ4KngejcjoQKwb/9rKm9i67+3SJ2vXn+hEFXm1L5P25xzu40LCh+PAroZejXDtF
2OMDzBmbSHwdaKT8awgotXtCtyJig4kOd0uGlG7KUapMgUUBSqH9uVBMA7a07uGBhtAYcZcLDkkr
sByIxMy1i14wLzcBEm+L0gC654/wz2TFlcrT1E0RA4/ixA3FwystAYNjHEbu+QjrJ6uC3Wy7sFBE
VcJEP1nfCQcDTtb8c0WPwqPBuXhxNeFFJUqC0nN56zKMtsbfao+qMw602MmNqeKCqx2utRY9WZ7N
2zrbikrX1pkGvXHRQJgC/G45xZPPXWm8lXuvKA27I41yqTBtUhPyctYGV2rZPsPDlq05SxNnr8QJ
r8mn0Mh4tSctpVCOO1/hnv96Z27J9Y3bbrG5FXGZcunLDLqQ6HkaaOvKq7SOefU7cA9Rvt8UIxBc
iG8XQf/Sw84kF+nFlN8ZtRJwpQz/cqW4Pps6KXydGug3qZyltUUdS6Hgeugz3d7rWy2apva1hOnB
l9p9pk9cQFfbLuNwHD88NJZMWSc9Ynt0gD4scygXD121yJ3lc0asY/UYtfrL1HPxSzsb12Cfs/4K
xTjaS6rHdH0510p0hmJy0F2roX9faVt8yywR/PhLcP6c5pmBLna7tqWVmO5KU46CqJOJEqCc0j4G
GQsAwZaMppTFQFDvUcx4bXZNNvtNIeiXNiPEjcwICH9y9To+zYt6QQxRSbnz3QkJyL7M12b7QfOH
ZHRD3FfeeFPgkJCA1zyYvM91jwKvo0HwjbKPs/w4uhpfEZI91iq5fFo8PIHbLDNilhhKFV1UUnHA
z6UHfmkpTcS/nNupjiwCvwTY8nFZG5k3AxP4ZRNoloEJHOwWuvQNKAIQasVtiKR3xfnrxmtdg/JG
jAvU3mgGnTVrPC5uOiAQZjQYMoqmvMRZ6DNwNYo7WddStJbjT/p5z9U2MKLSn7mjHcH5Mc9mmyMB
VfkKJj0Ho9XvGQ8QQCzgjwuorJs49TP6Nza0ES2dOhMusN001+ufL6QjJnoIEf9Og+HeQLBFxWID
zQ4Sea/kATYrKaC+HEzi/KKrUJWlQXFMO0UaKnIgoJxjr85BxaSFS/I4bJam4zIRA655Jq41CA5e
UseCxcFmAunuqCn8f1YUQ0QItFeQyQ1Utxf659o94oxlV0ucjshAFjd+/HRTnPfmaKzAQ6TA52pz
HmYJ8iutNdohxlVrjT7rlC+LlijAn9IGqYqW/W7zkytcVzxftV2tMMDs+prEOyU87gDXtaX07NL1
FeaFiSgxp0SenUa2HSsGuBW6j+LDrtK9mJY8uU0s2J0IESmMLXJwDnQErr3bqAnq8LWQXmdAMo5N
YYNLJolbcLmTPhd4v9XejcPzxIY6rv4v3IAmbpJlWOmziL8gWT7Lktk9FOI86drOl+ZdHxM6vrMo
1U4KhLA1NSV6LnmVlK9fjNeyZ4ZJ0y4ASKYJkTw+BdSQmFLOoy3nJsdNf9+un+76je0qkRnrAyDN
0V4x0Jp1bN7gusU/xB9/rGxHx7FnZFeTjy5j010DsX9IqGbcUo+2g90t0UHsibSj8NE9LA7EVWbG
rK0FJZISwfsAkfWJI+Eiv4fMtalCflzT5pNSXjN+voLXuCzwPJcd5ea0BeKBIFARXp/ZFFD1/DHq
E7KgN08fjwYX7fcHSzp1wsFUT2d8lWF3VGSBFOCAon7EDX7GzCB++fYQcENQA4r2c1HacjYxUOcg
I2nd748vlCok4g8MiBoYyBsAbx/kEZauDNjVzmA2CBP86acNWPyk5queWq+0/lH5ynv7u9ZKOnRF
4SICM21j3EmVVS4OD/7aPbUWtNbIJSp3rLAOwsPET7NcRXW4IAUnMtpKe93CBfAEiqkPYpGwnc7N
JN/4FnkMagO6QjP6Jy/uT033bgwrT1W/pEnlIjkSaiPh/ZaQSk2Ez5W0eTLtIDJb8afKqhui++x7
TuXvsmZnfeCUgi54hFJ3YFXwQ2g5ZStuBQEtZebGRRBBbO5puf1UaWaKBlZsMfkG2nhNBu3NtfTR
3yITyz+lCF1biKMgdlWpbom/D6/n+5hTYh8N27S273kZ4YNG+1B0ORQDDVMz0zrz7EsXOMexBDwA
F5Y4R9/EMARGHBStgkqAyxGcXqULZDdMAnHNPuDMRghUNfU/J+WQ8A22dglxBAxh4+eQFsCRo7Mr
R8UAxiau4p7Gv7ExI/cgDjx5WvKuuLH/sBS3jTu7EMZLGnIIE1WFCsxFXheu60xLT2QBkDuPLdXM
bWA2UU5GmOUExUkEQ3D8743DDeBQ0xbsHT0BR9VcPBT81kaz4SllOjxcghmSH2BCYveZ6GdLWyNE
pnOua4vXh+qGHrdDBjbq6UzA/oXqxLNr+4IjT0lkrp8PKmPG5mH1aUa0bQKQyDW09J3HLZ5ikDzL
rR3vNGyOLsiDlXpL+GpksFz7rfQrPTYhuBkYIHADVmdwWuwprXaFKEr8ho6ex5aQidh0KGKN3u/M
MbOOOy6OxBRVPgSfWeqRoZAl1SbUB2I9kuJN9if+6Pn4WrV5WC75BXN09VbNDpGGcSbGS9WNVA/Z
i41y/8bO8c8BhnZOHm3i5zviK5fdf79NNd9FNZ09z/zXUZy0Zx8HUwViuR3QdCRFqVIxnj9bLhPt
XiBLRu9fZJgYspM2L1RxZqMaQ5qu4SoifEuUHArHJP4+FE0C+77/LEj9HNpru0jaVBe+OG/nxKbo
ILRxu+UtnQ1avH3E+uzfYHalYGYUAJN5M0ebfkj78z2jrHmAWxqEsB67XYCpxcCK4kcUe+jqxK7V
MFi/2KV37jSVmW/9ORBppXz8kVIpAJpn/Rn5jIRfENeXe/A7aK6iwCGs4eTA/zVzW8XBzEQBhwSB
ilwOiOwCaqyPhNlOk/ZOV0qYf6q236QpN4gCxnFOYr//z5JTZLUqdXGfBfdKyYUPpDokYD5e8B1d
gwyPg2MCzSEiRZ7JX6ne/zy2I6Mfsve01/g/I1+3AFEIE/JhP3XvetpVYFTtEe+Vqo24SxKZNBKL
tg/2CGzgOdGkjCDLyfwZQId2t5PI6Zc/cCw7vRncNRlOrAKGePPmUyTWQuzfGUfTk8TmlzQlo6ha
+aupM8VSDbSHZCkjJxze1ezCsX7K/zSQMhFb+JncAoRRuB/JiUFnTC12u9V6QTlienFIZkyJIcCq
gzDXNhKT+JqAlHron5sIxEtgQL5feuWVYnZ+6MmjT3SQVs12ro328A1tx1s1Z+a1hcdg5drrwZar
8FOJyJzHnSfnHjdEgIMdIaCciPZdATOOQQxIjsWLPSgAMaz7/MTUzpwBtuI+iA/WbN0jtRULUK8A
n4bQOy92tAQQjPIFrmN5oa1zcYbviLPCaSRudYnnYp2rEBbb4rUF1w0e5ZZr51xcGq3p3VDVc4jv
shPztGzQz+/cv5bo/i3G61lzMHKyXZbWYwkPPeQbcyEUhMbHdD6BxaIQIEkoec08pHcSXEw9wPn3
pKX6rudDEMvLOwahD5lfyS9hIcq3XaW5VeM6qH/D6sKgl5c/ExbwB+EPxva8tZ1OutXfqjYQCR+j
cTbJg9uI/DM+TQZFJPWoNkaq4J9bA4cgESnAPZsM/TtrXxy5K8oiXTJ2XCfskBksPL5X1MB9xE10
KuSKSG5K9oy4JSN9jycmkKyaIVlBE/PO0W0FvwENpPaXUVay4H20XMFzPAq5X1n0DKA6SWasujZx
QUq08lkAFT4SVDP9oNei5aoDeFZdSFmZkWrDFz2osnngeaBr0W1id82ZW+JyqW2BYu9y8b/sHrCV
8zUSXipjUkTR/9JO54PJNSNl+WHzxd0+tl0mFcG1nms7XcEvE5d0Zq0I9W0GSpGak+PMjnfmRAUt
vnNeMryTalp7eBk/FIFBAAJQbTJn84TK04xu4xJhIjFVAwkfsvEms2G7Yes8yNpmqmQwrpzCwZc6
7Xy4dDkuYWmfxI4pYfjZoM/GxXR5uXrfbchpdyosxnLLwh2J/mFDSH8W3+xcn66iwbgcYpcyGia5
eYPpRu6QhedcEkleEo+k65RWhfzv1bnwGuQkfmLPDiScR4l5fvzPMvfFcGxkfA68y22/RRJCRSXw
osPzfpxzhKrU/TIxSAqm/Cbfal2eUUvTjzX3gAJRlF4ORZVayqEI+BscAi5OXfW6/8a7DqEOun9E
8lDzu1UEJ+qKaQvXL1BzH60mVhaycYcmVi2cxB7rvf4sMpIQv/shhxSG702Jt7pPkE0ro4Kqnv2R
m6jeGLjIaf1AryGsf8xyid/XIGHOOnh7kZlCFUK4PRTWHRYOtO1KRxJuD6l6AfDTOv+eh4Vhz2LB
Im4mb025ZT/5xkYQWG1raw/aORFhRIUdOWJmLiB0JCmr1yawfmqBXW7tgqKB41tyRvGSk3lVCWnS
8VKOWFgZ3YU1MMvsHySb5ZQ35Jba6XM0VKpJWhusV+Nkr69NszJqq8eeLaugXZF+ocYkO1DYC5Fd
vnnf43U82+UBqvPPTQnCS7K69ncaPtZdgolJ30Zsy4Q80xjDSBJ8/oF7GTufLgo6xiidCD34YOaS
lQpRR/BTnpil9PICYYcz3Mp+4iXDU2TqWKchKO72V9+eSoIJfRQaCzOr+vliqYaD+MFurXHaFd9W
BfW2KqtgPfH9uGwzRMWY7zuKrR2D2id0mmDkbjrE9t/DtrfQjqmLK6uFsFz1awJWgE8YN0ByUBTz
F1LPqCtBiUhBtSTKi4Bl0H2E8P9DveOdVtzlyUWBqGMPKDDh7Kj7S+vtUja9KHBxnCmjxoVbJm5b
KlUG3wGYWvwargbxER7/MulzamSIr547rnISnqOUp2z4eaulOfdvew7zThYvlplwXX7WREDe9xcm
2b1OylbgkbKO1TjHgHha+LAvTOYzXUIlx1/miSe6An2W+4t7EeHWAUpEi1qG3zjtO7lG5YPh6Zgu
u1NKbi6C0JeTEDFFwqlCrQzXPfinxUyCTfLUHhivBdiUc0/+38hgVmMLgdGvWl/YlxP1e5hWPH91
bqc2Pk968+ei/cQzeui7feTJQMbCgdYH4Xf3ojQNq4Cp2dkoxnGmU/IyAeMgpyNPAEQ9GRnVztJ0
VFRLV/6QylbkmZXwjVytmfJlStWQXzhfPhOOatJP9P8iawG1bPU1qj52NGl507ubrGs6PALdsDlb
7ygJqcjmzpjbvbu0u8ivobcrdrftNsCT1v+NxR+h11aDDNTOVnGfttzxWr8eBDWxgkwFdLDFNOUv
PjTw7+1lgaH57P9BDi9FDoH9ujAaXR0uFTzjybufm8l9N7o5XnlwX/Jx5FisK3N7QSjVeD0WxMer
QErwBvJeW75uch4KhSIGDSw9EzV2hxgsP2lKwwnVUQkOB7hZXol7iEc6lwX5eCGSR8VA7CZ0Xsp6
5BnoWa4akOqQUbORZUpLqOebg7zSNAG50u7LAbP0Pay1l656dDxXhwrYJ5uj3EJuYP9CmPpOlK1W
a9zC6aBlnvB6zIfXJwkDz/MHvt6nyRr08eXiM6v7k0JrCLqzmE9YtUB7kyiJ99IKzE2pGD2bSMSD
DmzjSkUm8SCgR5NcXwwrgmn5dL7ArqCIS0QdoEQvekb0Y8FHQ5VFVH6JTQQGpN8QS5WyNznPsNe4
8KSQUy8IV6FLmuURPx59H2STu2oj2eajYeqi8PR8bHmp1lEBnrxHZ/w60B+8KdG1bpd8+XQ4TNf9
Z1Nnmr5qEl5YJRywy4EGYmI7j3Q2vByhHMvIq4mXv7vv6Nv4GEDcYbIf9nJJxJb/IhfQxdhHLFMp
7j7SFJrJ5J4JXtTEecrM3HGCTcFhZT4oANQrk2kbC46ragFT1fl8Bhb1LMoAUVdGsdETRCgE2SNy
FoSunaUsCNEWKW1M6Jv0hoz4NFgqtp9KCu4fGJyRAfp2gMLqd8OrpsZ1n2aXxUpzoGZuTFCKThmU
hA6Ycc7IEG58Tu+QlnDutM4j32YaAxsbwRUzrGk+SbgD46CfwI4LzgZdHFBj4RT+Hs9RnQPphxHQ
305h8jdh85sSgcAYNmyL5eLWhwCRN4NBKiPn5mSRBtZnGJAT61F+nPvUPKQ7+FYTxbkQwnsG4Ank
BXmWvpANhMmUGGLH8SMiTh7507Fyj7wcsw3Xyz1acd6AM95MY2UzovlQSV5fw46+O/s4AE+mBXD8
SEnKabhYAOWhhWUJjCFaqg4KD2A66kt1uo8g0R3iE3lcO1XyxOrdd76laL6m0EC31Sb7jWIUW8ZV
MQYj37FsX0uRCjh6eVZ7/bSkdR2U2+sYrH0CcO/27Ky9sFyP88cuw2jD0uL47BtyjPOKDPXCHrEo
zR2fCBwGk2wCVXsyY3WeOeXQCE4DUt5Eytk9MUI0+J86gwogA2sbCwJzmoEOI3p0iaIhBrRjXtOX
IHnxcgJhSxogdA2JNyRQ19hQwHIPZUKYqtiXS1GoePNetvTUE8XAysSeg/S4O6Cj1hbYXzTEWs8W
qB+/qmpQEH4TvPbQOKA+0Wk1GNgCH3hQBe3cwfY3NHU6AnhZD+ZHg2C4gjzOhc1j53yaiuaXRXeD
M1a6ccfmYF8CJf84uJxx8CDfhDZDx773fZpNV5KqANrEuTgZmSheI+Urz7Zn/xSzE3vkN8uRABWw
MfG+9joYuhl3KV0R39AGcEZBL1WFwcBQKZjhUc2nngRIuh9BIVTOR53SWW7AA4eIPzCWzxzfDR7O
PXtir3ceIEJ0IRzV3SJBKannWoiVlAcZxJPOIvk6t/2bnk59Gq5sxhtR1iBt/cHQTwbfnc8tsagQ
efSUUSDgfMaGSDoRXyzte6RDZivdqf24WF5/8vjV4niBKn2B4ZTH44Sf3EW1UCDdk8c4stQFo+du
VogRnvmYU6vXrI/wbXEKkHyI/HrcBd8ppIc/EKQWv2qQXOc9hirVhC1OO4L3u/Zch9Qm4SY2Zcpl
46q61Lv2UHlWbp/iUXgS5rsFyXTGqBms7rSgbILFgATyA+DaAqpMfNRl5s1XzyT/Jnh9cySwUiSR
aWkqVRJsLN1K1bGR6+TTPf7zJnZIrOKvWGjB6GW41860GqOrZGi+tjW3ZBKtfCKbkzJcXrJ0Zf51
1Eu3L4sXyMZp5JPYV5LZEUWasrkkhGOUNP6mFYHg4Q6KQm1sO5l/gvEBuJEjcazR0G/StSNQjndE
IAQcMxbIydfXPBFYYoFIyQJYX9OnZ255bP5bGz4DKsSJC9VADBEK61QW9KEB7Qq3L3cO3MHe6YT5
MUNuhO3Rq8B+m6y2LGGp/fAyRNhKBqnwUS0FtEboU6nFkU7HWNlOiJM39OsXHPnh26dqSUakM5Cj
UJ5T3td2XWZYKR7I7YWyxcAE1+hk906PmuSKKPEl16J6NqY97HHozD12xKEZJKwPtNZ8oW4GA504
1CirsANK8mkZ8+tOKUAAKyRPpBneA2rtE2g5+HoUtCECYiJesooqrJudhfqUo1FoF+TNPWYMpTKN
tnaHzR+W4S5IswKcntWq57mnQvq23+cKeOlTSNIwnxIzr3qIkP65aOZeWpuCldLHuflPSuG83nbl
4QV5Mg0K5f2mOESBoiOaYGcAf504xofRJMRi0jAoYSB6xDyEZFY/DWK3fk5Ya3zOjBBlbc3zi72L
jgEtMAjjQ8+RDslOHj+OLV7o+aRniGrcHv/wVr3SfvTHPoEfDk2B79faJbmJ/JheQ7bbDXHVlq2e
UBmVbzvLsFJBglhltUW1tlO1pbQpXXLf6OlCGZ/JMUIl0c3VqVIlOA2uCnGTfRSp555pSw7eHAO3
cUgIR7r2AjY2a1y0DtJ4E3wnBWtScQykj6sWBLrdSf56lWaJuhJqLkT1q8ro5yx1WJE/I7yRk2uY
uBSmZqK6tdON/H/RZOodwNyWafLgdG7bkYSMXzlULhSDEu6Hbuuda664xnOorgS2L17qTp0JycUO
XBW4jVeg006ZrQNd6AcnFFrA2qWSf6s9tuC4nJtI2pMpuzEEMsXj5T+MuKMXSINh49+n3SVJALqx
5yIrVAV6ZQCW/F5UxdLZtF9ZtGtW2T1hm7Z3j/mGL5Qfe88JMYH0MfXl7xH3/QP5xRV7MFO67zdQ
eqFWJ2EXNNvzVPlKKORsVUac1kbjfkII+d1usmCSOS3VILRaePsc8JrIUj5oirmgLUJMlgk8fQbK
B6bGKhVk9tiuAC2XbIyjiko1PgV/Xk6uSE90+MLuqKMYPeVTLUvyH/iBz7u4MFDvchw9FJpp7Ztx
ujLJjKjmooiJIXgK26OOpSytfkit5QvbosGzHKwmThB/qp4p5Ad999vwMde7ka6bumYbly2fKGU6
gWOJX6YJEV16j28cxTXLqZw/cHc/2tVwioO5BAy7l7IBZfuQsqpetgnlNWq+JBPWiNSRqhIK9CM9
Melmyf+C7VcGvh+4Gm3CRr8gEGUqZBlQM2avizaBhTHgpKa6p9FnpEPwtxcSoIz4woZ4vcvwGyUt
QCxFwqVbpEh6VjbRu3WvIJxaC6XQ4Q8h5u74VPcFCPB6kVAs6ZryBQS+aiFl2gtzZMxrq/l0CeLW
BCkXHNkjp4NvNH4HeHVtNhrYnxM5O7y4HK8VMp51RBQUOOxVOx1P6lZOlwWKutPebIE1p0satnte
QyEcZ7EuPtpf3Xx23MCTcXZlnnzi7scsTlQNSiDgvrC5nv2sAprC0TpMDv0VKobHf556E4INvsmM
JPMShf63EvoMad8icUZ2gvcuuzE0/PKyDV2BM7I2L2U/GAJNiO360Kkmm5Ni9jfxhJ2e98f9hRv0
IaDBiVbFChixZoD1WjQHKJ6orISV/497l8c11zhKyVeG1LXg7nkvmbYB1I4IhYbG9sjbYwljYjBg
1zsejWw7iFtva7a3D1vtbjpd9rfohjms1uXvI3jm5iB3XMYMTkmWXQzIoCgp2wbS447CKCxAlldf
H2LPMlJwAkg7H33o/LKDy2nJGSu3jyD4qqK8pLjxcHvbTpgA4p1XqYceTHkJ2wF5F+asCp8q5ipx
iax05yvf9/zWXqjB6XrkjXDImrJc1BLJXO4geGcubgbBRhMPbsQbq+/slALH5gFS7EnvNlfLFYQ9
pFjjdMeod74QMry52vbAtwGvpKADY6TVNY8bqOTQqoC4AOnVHfxkRrF5aNGF90/8BCfL1qpYsbHI
QXgVRqRl/5rU9pGVhgaowi5qwvUOsHXw3xFnJe+LaHYjN6TaUJLTleRbX3osBxp23DHzd24+zbPQ
hYaw39msCFsMdeRywDb/tIWbm5+c/T8xG7+olFvofx0TBzBlGAJXSB8Ne6PebNclY/q/WZaviCIy
laMSmo2WIu3MlVRA5PRoNj98nHe9HWpcRR16igIjMUmWj1U0iqEMtiLwQxtvVhtFVuQxqusswoJO
G5TE1PdA+xZVxGnPYP2R3fsmCHHvoY29PUHNYtf46grMNq7zquj3Rv23C+NR0VxX4QUB9Grfvp6+
UZjjgFbfryIdljONPVWR0eBkcJIZJ6oVGSsT1V544hQtNqojxaBOim93RRQTrosMwiZvuahfchBF
4d2tdMQSUKPA+7AvBcfT1thJDNZif6SXIrHbbUXzzzaULBT4MAvA3e4erA9QB+6yQqeuTvMngeUN
sJxtWf8pjpPrNBzELmuSzoEufgWfjKwzK+/cBH6qbcT+Kn8jeOdhKuDFoLVIys+5q4NJRkSZuaPb
3G8ns9vkE6npwn1FI66gHyOLno8gEIMCwC9Y7MIIhGOBGfADszfG7RtLnJB9/Eye8f6HEb5qAldp
dRSDXM4Tj1YUpAR6n9+TbAF6/DG/XhQv9Q2f4uaF3G8I9/X7Msnt7jfixVkCTDL6JlpeuT8sN3Um
VF54vcNOKvb6G1KtFwfUAqzo7TZIB7YgUFl2lmtGwEMuatHacrmLlDnfU+Dsa75gOqoIq4Ik5Tc9
FOOXgnMLjWxTpMy+dqyAZ5C9RmrdrAfpJZd8eJFkX9n+HEgFGOcAD+AyfIPbMV2sVi2LFNFBRCf/
tSGyiEyoyvjr+V12o1G/trvBhH9C51/emMhupTKLaMmjfBeK7RzBADmv9bXLcv32jye5wuuCPfk2
XpJlmqsViol+mBieVilJzMrDCpIA89cHcuT8u8tyur0/yoQKyaCUy/7Ua1KuzT5SrNUd2lIgHR6k
AIzsIYI+IB6UrxLV1RXD79tw/aMwfq8qIm2aSwSseidgodLBw6mAReW1oksfPh7hbsXnt/ZEkbCi
Yn44BFBexV/ItrYg/6eUww4k1tkivNIryiysJen2GSPWZStHVQASLIV+F81ODpEs9g9iHwcLFPzO
Q9RyU96drravTQ1fbjbt6ft52I6F2N+WIw44msajsMmYH7d07aPlxu4mg0s48KmjSD/Kf4IQUP7Y
CGcPVkUeKhAsFNdnLhsTezRaRMcrNL7x5wwems00asdD/P3+eMDBltMHUqOAr5K7+cKlhUsuIZAy
gpO0/PMTd1akdhHZdRZPU5FhBamBiVhx3K/cWLBGjYJaBn07zyt8SMnDLa58+hbRc5Re/77fchcN
XO0IYBLW46zvToNmdTZZjA9RQkdpPRLwhfmhxjBNDDytisdxKkl/MIbytbVjSgIGYRgZ4sBLtSXn
tjDeIUTD5ZqqYpp3bdbbjI8Vpg+bx/7SzH/67TBsYd5AX9T+VpHk0K7NV5AhlWrSUgNOGOFDwQvO
Kk/74cV4zesBYeOla4r97AvnT+AxzSY8N/BzXhf3rZd4DSzRBGweIZf76ir8WCEVsjZN+Fd035Qu
u2N02QUDyhE5w1GREAVc71ehYLUCr8evQ5OYRb/Ig14fcvTaLAhnsQiJ/7Vj+pRFGKZay8wRte+R
58Cy7HyRkubzXcnSlgIZD4/a/A820oUBe+r7zMwh9AhjmKB7gG6XB8p+syFFn6HBjlHH5+pBFsVU
odeK9D+M125Krq73wVWzjCbiRKPVHMeoW+rGIABCTgd/hrbbBZuUMdTa6gYob18NKyh7xxhCa+9/
SkYuPbKOlkRxNf+hk7MhBm/0FaAbVyo5aNDRRv7AVQNr71y0B66v2BBXG2JBNY8PU3HNDFVOyef0
BV13fxcEscRrQ11Ou/i3BUJ2PdtM7ACbovFOoI1e5v9ozQoOpjhmXAu+5odvSCwegNHyqSBjmauD
nyluZr0HpFrsl2eaFmr16pW7OpOXAadGO2aEJFlag9WNh4rW/K5Xbu9cbJ98q18KRZBrs8fXWqef
B9jNOv6jd5e1WFaxyPdEWAr9VcEvoxjt8ebGx86NivR0An7hz22+USAByaS4B9TZHwrgTW5ziC4+
VuzdG/5tKhJd8oyrako5CfV1JKR6Fzq5D5n/GIQoi+xYts8y5jnHEPE1GA/qseNKE2SYDgNYZoqw
3pI95QrDv0Ecd12uVdZiIBIjU00olaRhPHec71xf8/SQcEh0C6Qhf2c97rxe9fqv/2QwGhFJc7S9
TjT/tTJLeaztPg4NZY44gNxLAo9Tiex4ZGDitVVOW7uYq9FSFG7/yI/Qhge7JSL2DzXp5cfs9flV
hPuUpkY1Z7mE0b859lmTQeOcsbUwl8DDF9ydGo1U4gaxNGcYAvF2Z+igPUk+r9tCmRXRWOTIma7b
gjuFgpNYIGgXrKSez6mBMhzB6Btaqq7lQCXeXTwb3gu3hxnzTEdTIiEjzgJAljsXvqqm0Z/OemZE
qw/mtcom+MGyv/t0cZzE9LuLar0UKxHlnCEG6+QpQTJB46l3ShpMroJsdGwGKj9ZfiIII1mWxHB/
RHzL4gObXOq6X8h83JVRGyLKU3bNGMd2AgsU+IyIKObYmUBnf1D02bvx73I2/A6W+MmBog6wnJlK
TwquBc27N3ilAuM1CAFl1uONYbfC/xL5OwRa52nxErGuYsG8s37Sm+VlsJIpStj82cswfQA2Sm0A
Cd2s8Mkkz3lfHGtYUGIvT4nBgOI1FVjmyF71NYxtM6jP70rWKcY0QpLguCjRR/fxYL2tgUcp90UR
Grsmd9WVCjs7i/HwuUkk/bl1tbXnjfn2keGLBv9209k1eTxktA4tgxv8ZLjcVIysnItXnhPeyl8c
qMBaiIR6psZbk0UYjH/8gD2NBkSTqOcaUb7LMzFF2M5Rd/pwT1A0nShWqAP2RAvl5MuTXkg425Rg
MWM0zfhrv5YIn+qvYrVD2qXbeZtxRIvmbI00TkjP0mK3XSP6n2PkSpH9DDhQ6tNUGuAoA1nsi1q0
9gNpucifke+zruKOOwn6vqe4JwJgJYciz2UEO/JxZE1jmegHV17XZOqjP8/X8lSz6vsWMNfSQnND
r5k0p1mRM7RstSEd9a2PumZ36V9cVyejzviOMCl6MxF3Dazd/DxjHAdxKHaiQ7LpDKsF47q7sonl
XFuat82vF+TiPEhxxIf2g2H837exkWIZa7OWw78f+WqYpCnUsTNeHNFl/WSkY4OGF3wBZc9sr6WR
4UEaUGAfPHdBD/hvQCLGrFqDmUzNYAAiIaRCxtcRhQEzWZUwZRk/LqyPq/8VuEQ14D2WxN9uE7Yh
puJrxGoarVh5iL5DSKLVPYs+trwClb22DuK2pnYr9iJmvX+RgGHSk4DsCcaxEKpiD5W1aWtXLlah
Os4tgqqi16C0JADsimewJLZ7Fl38hFboZ1xPuwLYG8z/yUjZX1pZVjzGKuvUWD9tGqG3dWW99Jt7
b2ERpH6ztp+PoW/O2VZXATETDVRVQhM3fFGJ5KbOZrSyFPsWhHoQvmc/vrDfY+JskqYHYxXVbAMy
+eC+pR/SAiKga4smFyfOr5g/V3zhuZO0fDLtuzPdI4KfVLPuf2MaUcIEUYW9ar78xZWbxQgyWSzF
LeUTG+N2IxHBv3dD65kcIPyC2PZ1cKU8a+GtjeI0/3Gkb0VTTGh2V1MbYGen9K77Ucxv4BlVUIWo
fw9aIWEkc4vzbvwJ3p1UPQ2dbVQlEAWYz4VSGr6GtoPK0+zrxReljeQS3b9Z9UGu/A9nKk2k1X4q
7t45qvUkalQ9vxopj5v55cp80j3sWY+a6z0CYuVg3zrSEPPc/ZvBhggZ3b7VsTunPSUSEteWlB53
FReehQgVkMcGrZTU2nOFu5tHdJB1WaT8r2Gh7oYpj97j7bS3ARWbxKCUcVtuBG/sbbw6uFyk7Ic/
L2ROuhcsx/O3Q/WhP2ucZZmSjtx/M10eJqwlQHvABIJp88F8JUFYahmXEMBsGvsjAcS00WELaUef
jMRsoAiBw06Z9yKn/VCVMSIEGPwAXWoRZPaVbLapV+j9Ub0iO8T2h2BJADlTmmrgZY4YlgEvFbih
CJbu7zYs7ALQbedek2ZemSYLpt4LoJIUHuSxuXmcD10+I30uGFYtEOjhlu1wKjFDkQKO7uB036DT
Oq4W3Y4v4lhFpzGN5Rho3KTRyD9cGuI2eKyQhUAFdQcUxzQVlHVzbgQoi3XT7VvIPVWl8baKZZAL
+sABqq0i6JA/ORGQqbgsjkriUVb3nsBkYYmPaochgOmpDuZsW/vvdO9AHllaMzwHaaOQmoatpQ5S
GzsKF5RoJDeVbmK8FiE9wR15L3Z3Zop+ro6VZ5LkBT6IqQsCxJCOF9dn9p9L4aKZum39ZiLmJe+o
Sf4e2ZIlt+UdxLliyVF2YEHp87Hx3sE6JTCDJxpspzlYZYG0s2gUWhQLf88ocYcSDQ6CTy10Jmxh
+apyVuh5XsE24m46c+R2xp1JgiJLMHWJ59DOUGblUA1wBXKf8F1coqfJ5dri/N7PtC0KmBEGhvi4
8r32v80gXVphZbNtRRICXkjHQcp+cuciSwR7qmUSj/ns67GWbkpAROLBIdJQykb/s4/p2lAw/AAn
K/gxX8MZ/2GSp6zuaHWgEylPJ4WMzDWIsNuuL3V9xMVGopw350sdAsCTorZIZiDmuULymh745WBD
1Z72u3dsh/q+JSD78Cgkf5qg0RWTrw6Fyi8y84bg3tlk4GZmpZybJbmmFOUlqm8CZn7+y+3uBtLr
CYz1Ah8JRsyZRHSRTwk85liybcQb3rv2EJ/6MMYFJ0Hawq5UkwsLRD/1Dd0hiW4fgtV3kXwwwW89
CWuf3ihSPvdSM4q6FKriqUqAY/TE8yrDYfEBwcPOH6sJlpmJLxmh0KB3aKfkmv7WEyMUoYeF8e+V
zAgoI1LdcGONAXhHxcA4s69khc9VOV+Sd4OKloXbnnwCoqhQeadYPiG7uoupK646ofqWN9Bj1lpj
suvv1LV66IrmODKebPpvgB47ZT3IoNmgTk03f748c7CmXRZPVlHkQ5fdhiIIcu9Ts++zgjotY9aJ
HWHwqIrvGek8ngt+dz3O8Ke6L5JaYvdJ8I1DMleGumsmOUIweGI/GA9quzkmzAJdqh1uxHuU+zvx
iba4HV5KAnDWAoA5TviN9dtWE2nZRt4zuWMB+4Avut4L75c8h+oR3pmAjsFx2XarWgkEm1op0POw
qlFp9t25Xn+vxlV8OsurzaQoeazFKStpONBLYigElGsoFXDZXaiLG9V4SRqXyLW4P22voUx2lO7v
FG8pq2b3N7mk7Fy0Y/14jBzu9XvRR4GoaIMTM0qvZ+sHM6J29GtjDLGMHG6nWIQHWOZPM7f3rIty
J0f6ckWa126Kh5zAk5Z73g5N1HgucPv6adTWPZtUEFFFoAPioQoGMOR25ZC/zxO5k/MUDEcsjaql
2+hYITG6VCj553EOx+kc6tQIP/zvaBeMDpZhTiPBrpCawTAQiK/7dJoDXGwllgS1ejlAba2O26WC
HYQYI0cCsKRFBdDXJSWMdoEo+SldEK9HVDgPL/iSYz9j/JjazHcvtbQ3LazBp/moHWyB6BY8Lauh
zXXXF2lGN2lD5nqtdg8TnBTHyIhayBQBOMdmtHMmfbkTHakVywToRBx/S4VkQAuN+tsQgp/q0ia5
vdth6kcz7B8gFO/nXES/0An0tk5i7KXUe6/+oG0pz8yoeoCSl5YiD4m02a2XheDZaBFwZSUniHe0
KHAzBQe224kAq4cR67yYLYlZ5nqQS/TTjbRo4Cozwbkij3Sr3JXgsbvROcBcaIpxixKTNO7enAFA
8PeBve6N4Hj0Tecs12H9btG/QzZJT+ncoSZEQ5mUgpzvItgZ7lqtaDLNJzMV2YE709O+Wg/vzocD
evCUJEoRPQaLl7U71KD6yw3M62ZEOK3eH3rsQ29cyk5JEb8n4kPCLQHpO96LrIxXelwJr56b8pxz
5+mPu1PK5ON7TCVhIpqzbMjxpe3dtP0HCz9XsVAIMWAZKNAwF75sAMQK25S1M0pv52DVhcSD0uNv
rFEMlBFMzo2lTxjwis+52GVQw8R5vnZ0k9Jb1jURoPEbucLURfObtAZkVcqkLY6bKDXn2dUUoj1m
Y13UH9dRSqmwweHlvslm09P+n0zdgI8Skjp7t0aINXpMRYyuH3pVL48WrDzPwnyiVIkay4NyAC5n
REe+50zP3VeI2R1BWj3zdYVOH99kTGO3Fp68iQbTcGJzk4izTT2DCfCx3+S6MKJHX1gK/ZkeIwGE
Dy2VWt5cNeNefCPZp4RyTm/wZkpCK53ELqS1OvMSzX8jKAkcwDAsKX0nsNvml7Q3+lp4BOykS7oZ
qtCSmbYMmonHaDlD73jaIEEGTeL82lYAHt0IhK/NYcUOl5BlUccV5HwAeKDzuV5n+epfH/vBCyPK
KGr5uj5ITU+vVp5XdywXCMDQ3yJgc2HDWWcaXWWM9kyGBSDQX4v3VHwChNX4jju3dNc0a+Huqq4Q
xH0SyrJ8pYyVrKwiDwQzLjIeuwjLxHX5dTG2efSdkgNcXsuR6lVIyphesbNVuKrxt1DKfYousN30
Z6xSs1drfPoXCk5D9Ldk6XKsZs+pN+wLfJvx13+62I68c4wAMRTNmn0cYon3iKQwcr6NfAAZ+J0c
EytWIPABY+6K7r4A0uskImMjakiO3BZgazS+eb28uBN/hCq5WkCd6DBTzfALg89Etl0o//U8CQ3T
1kBadNFXKI/KrtM9Z8LWRk9t8xDzaji0r6+klPjJpGFVEVeb84ppRrQnZIH/hOjPdO0fmrohK539
2wd53EQ+73tdXSgvsIs4JQE3cOn2+Y/LwMIf5jjg4MEjEvd3iUqfAMyY1QHz5KF9WmjiHgbihbK2
9Vaut/3W1R+h9GXJKItaXGY/PNGj1uJCFg8fz0kBOR9JBG3rmO06cMdKAOQ2G7NdGYPpIV/2wkzK
CbapWPAFiGjo2o6EZZ1QFntC4aXpFYrZEtFiU9bc7uz5Qp/H2BntbTYqAA05aLWuYjF9i+y234oX
OXZWnqMISiJd/MFvoCqAWytV4K8scoC6kzv/RpWIswmabo7SqA+4D6YVe98pNxvSmM/ag90TaplO
rjhdvuM/YxwVYZsYMIVrHc5GQxq1JNUIbDNoAHBsYzvd54VrTtVw7y3oPbv2CsAJ60lLzYHuua6X
pIJi15QBKVlBcVKRbeowsAERlVNYAPqqTaOT5Z3KexwmPmW9YHDcaqmquJ6kQbVv50FM5v/XDx6q
351Vpi0DwiBrd9LLuQm9v7CZqJtuX2PbM2WT/OtdpkA05HJF/UEUOG0lpOVJk0E5QWH9L1M6Cj2C
H37dBVk58n931PavCoxT+cTRSjZKsj0f8mRm2w9OOSFeXkISAERaZw2oIxRb5hZP/KvcNwN73zeK
l/dpZIJiBfAjOllarhicqYijxgCyTEjaLnkJNg6z3nRwXSSyJcUMs2kLTpdMqtYioA+7z5tfxU1/
sEvI6sYVtPcEQj05JCyVQI2zjs8CMcIK8VsU+iK1gbG7b9OG+PixPBtrwKytJNaSFqpm5ARNbPcD
ndBYcgyQCWC0M7Rsn+IJNOA7p8wrshWl0+fAn4w62k+itPDv7f4aUHJR9JhIjKFGFfPq8JyRuOZ6
3ayz2kKkxfJIN3ZwL4KJr4rvuPedHABBx3zz7pKZrduLVwLhjI+54gBcizEL452ZAcZjoYehgFa8
me5QS/KnDS2PLgdgQpyroj0WX30gnXCvdX8mWnOj8P6BR6kCHut+5CUDmKRTvfgkju6xhSIwnwJn
+oWWzYo48jzTqP18BPcukafXxJQ63xyT/XZKbw4Q6LFu6YHJEYOb9J8LMoqGJw+yTaNHYKg/fZvw
BrbTP+s4mKDIVw0iSWcjqiXGGBhpOhYQZwEgPYrNELUPgsA+04ClzEVpSAcnVrvFz/AY7XfeLgHV
/2jHbdo3kFQ43VqJG71Fh5bVXYPFLVJNkzhD9LhdfDJ01m073ClvF98ztownr5ouOJeeZ3v/Lvde
ZcRoO1Aju4SrP6TxyYQfOwG2N41f48zhH72BRxixWTAj+m5qgWRSFlzlyJTqpQtP1TDNoVBmMsiD
UcHU5IY0Ml1b9voDcHl9W2ZAGfRiWbBxXVrhbJMfSu45rdk48RfsjQvxd8iDVRpspwe5bSu/Oov9
zsv8Dnj4J7wZjisCmLzC1KEmtUv2wGC1bSghRrazlwupYNIAwRXvXHXdCtJBjF2e2b5iRWvPT4vJ
HPEUdpU61A3qf94cXSyGvaiMkmazmvkoEEwtkeOienO/opO5D+p9e5ULo/oulgVs8S5jeyKnc96B
WAIznhWA2LRRWwGGaSZRlqPdH/ESmm53bcqvsWZZQR1yJJs1+35fxeCYT5LBdomzY0AJ0TE8XJB+
zKyRopMikci2LvhxfgH6DPH7Ih+e8+ovIY+gt7DKKcz6nYVdOg1sSPSJ/h1z/MLrEz9Ydskmozuu
5yy10mI6AJtjmZ4r1mPJZjUQATMMLuIESPL5iA8thjFIVdI307QM1TFPejejCNyKAKXEyubMBm95
uWSBGRDE45NGeWy9lD7VjspBRsoGOuyCEqd6mcml5tpqi+je2Vn4clSoZm38Rt0nXNfSrJ+sZKAe
7osvy42GZn7b4nHuHxPPqUdfzwDcOhkX4hS465bAwuxRcAcXZec7JLzBbKGygOnoBiKV/VCBl6ys
D0gkUwpBJUh+KXcMEbh/tXX0Jbn44nfU6tQHW5yx671huUXDQy7H6ZHHs2p4KO8wr6FyoQ8+DdL5
vdZZNyMY7s407JAMtgL1oADA3YimWwwL7EDuehr2FwnxPwlIjRIH05dnwz/md2lo42eIh7DiHSrd
J9fmJr2P9NP3eaC2cM1Uj04arI2S4nkdXWzyP08tyO/jLjOl8d1bIXrPiFxrNMDdRMkzmrlO+aBv
TBJJNijDsRWKvU4nOEgbycrIyrtBtgdy+VAv98y8VFhjRdrrQ2ri/3C+OaRC4nZXRUaxPnv56qA2
CrraZn+Waa4z3WA1YqiIXSu5mfH2AqRQLp/d4tRuWlx5+KFx8qDmEtOClG0LhLqUGnOOM880Jroc
3eLl5nSaZ2xjAfYBMg35oZqcMObpy7dBvdiH2c9iJ3AVtI/JeFvWKiW3rdD6MXr5RhUtq2Rz6Z3j
9o9s86BsVaLkIPp3aD6v/HH0NWrPevFJsABuX2JSiCYXD8pLQ3nYv5r+RiPpgcYdrYL//BVURC0u
GY+6B/saQm+GeigESQa1IDkUxm8LyqZN+rSOFG/hcw6XDTDGyTHv2dcZKeJ9iTwvuc9Un/PbiSAU
ak9TmbU/K1L9UZZHXvH2CSAesE32P4M7fJQeqavnpSAExhS6O9sWH6wLZ0zATUXVS1bPBsCRi2QK
rRwnc+1WJyW1YE3KVS5pfRlYaQXFb1nJQfhrn2xJz4eoaDG4qS/g0cBZmJwxH7CxXsTYe6pcVO4L
ihvC1/GA+5RxYZqATjXHPE522wWdTzxgmVqynDgbjHRyLiRSJYDQGf9hdjpFTIw6Wfr7UFDjrUrz
DNhjFSKehztdWttSGOXW0BuVARfyVuzAuWzeQrPODEHmiB2wRdHEnOCP30ZeJMgB+cgoUoAelj6i
B5n2PHphesJwIpfQYmh1K9TDWP0kHjt956ezkL88E09G3ZF0Uk4uPJxqqkXieuHXH0bsNGeMTWXp
DjX66a98rdH1HR0/YtPK5X1Zc7OoBb6EetDW0Q3hYjTdn5Fc+V9CGXOdDvsXPvU4KbnhrUMDCnur
hHvGKz5Yt0nS2mJMOQzqxDySE5So+uNccD73lw6HL7QpYcL/kIkNmQVZePYavXXgEEvQdsUQlA10
UY9wJ9nKNLyFMZGngeiBF+DjO85rFG83JzGhXkxalKwI8CzZZGUAr9rIwxIHQHDH0tUDzdb6HEPq
RtVDkdPE6GQqNh5h1q6a8+9bLesU9ntMRTAr6szZorxDhHSy/80Hg0AXzn5+D+dxcftl6p/S+RY0
UzrHFIgCLMpNEBr5G9315G7OfxadSgCHwyDNPS/hRGWL0lWiX2n1V6xojeq1MUbf6DijJHhLpDuH
dXXRLAOT9WvtHj4QLGaTCidXfsyUjADJf8By5D/FtpenW5+21/rEbEzhhoICyTLacQVfOxF2NJVN
wsxSGZTnFI+Bq56YuQGTZIhCJTr4Y+SJRyv1JlUFW71OsZX0ICiK2vVV9pfe2ewcgPLHSSU9Uoaj
uzqUAFA61MjKy8ITYrGzujcW/AfbZSDuKANFfWficdl4iCmdqCccLdF5O7OKrRtTr+Mr1Q4Cj/7F
wWjEkk5/+9fGu8Tk4kSpKVL0myb6WCxSGUAXc/MNe8aJJ0mRQzUNb1x5KBm9EoH7tuQAgIxS88LX
qcT8WCZUihEwmKtZqh7QwD9y88PORF9MWcdvgo8rTAsrdMnHdEewNPD1YMevty9a2+vOCuWlDxg3
6gnPj/d8MaZPL3pCZBZ2/LFWCvs/tLjxfX8Qrfkn7aWVr+u8vLXQnUdRkl9nrBQDvPLT18E4FxnG
DF3+y7aRrh2tp5/oH3sKNae+bHycNmZjeQT3nxOZeww7RXz0Yto+okyf45VB09yHm9n4fWFvxRVh
YGNNQ9MLRWoCnx4kzFqDuRyKg0plBvx3W4isYcv7TVzWz/LgoQHEAVKRgeyBT0by3nUum89MCHTx
A4eMKizmyin3psGbaDvJ3KP0KrmRR50uhpwOkAUmPyoZnChz/dYLzICDtWNW9Zk5ynNuh71UH11u
x75EhUJL6SkPc0h/h+F+ib8YGnu7xidMAM55x8Qol47kGcEmoBeZazTMmXoB+Y7bmc+eAXGxPLw0
N/9T5p9ghizFdIavD9IkKBKUZWMfWeJqFNyTQEiVShcAlP+iXWkcevwqWYUPXqFRWBrtdzPf+Yvc
Y/SlrXIyaAIH+yl+KaRaKQhOYtMzMXkiKqp1zM/h8dkbpbnmqQa5ySA5rDC9hXIylRQQ6FVzt/9a
VqLtLrivu0DJ8bsbj3263EBu60P8nBemBCBb80ZQ507dSO+oEuiu4Ke7htxyWObGp9vxOfJu8BRV
M/t9FO7Gbw+Yb5oBje/dfwH/65AFw99JLrC+V128Y8LwMpnURovYX427NHoj0AxvPNpKgB3U11a3
fKV4jhJynAAJBhXP7puZeRvltwaSCyugE4dXLVZJ0s5KltgLlBTvSoUSAI68MlrDQkZA7o7GQ/5a
UHDKOWwDlV3dxZzOV3SZ4s6p9f1Lm4tZBkiBVcrufaObIf4BAxh9zZrVOHqw88xcdLZdjdrgshQh
7SlWEGbvQrBIO5piGJuvKMbhivwybvYxMtn1WmWNG4iA2Zz7t56OoNXd6wHsCIG/Jul/tvGHynRY
pwseFmmXEzcW88yEA98E2iPvrWXipa94KjrEbp0NgRyJNi4DIW3Yz+zx9UBsJ/3FGDRuZ/SAAP1f
LyhdrHflfmDelJLEUF7E38/k+FcyHUjC/BYnBhngnWAPVYGDmKFcO6y7ozOPfwAL/j28NfN8jJ8k
fqguBK2gNtk2hTtSlIBrM+rpSFMssZ4WxhxFYUKOYq4HD3grPmVnzj+RxwMGyLF2dMx2WqXpvdPd
721vr1Bfd21dpsFtCre9NZ1IRIRYdnFGPN3u4XlbYgaCDri18Xbr/ONiji1vM/olFUh1fm5m1pPO
ZmO5d4tj+R8VQTVIGBSpLvnN1qAX2qNMkkHlQNkmnAi+fiPeVvMtOWlqEkKREDyW5h5fASj+1BC0
yTtZmSFzTnp6NlfuHOGzW2Q3HPbEwMjEB/FhIKysvvUqt1RQtzt4DjCIEKbcMe4KJrcm7NlAfLUz
9x+SjV/dGoMJUS4eoYbe6XhvXWBagAewwITtJKikYJ0FHrBWY5LueMy2WyoELKUkmaaiz1F64JRn
aofVKJjeeffyPJXssIdP2BY9tiFuuTMasXeX8eIIK8DSf72unlykcN3uDJXGBBAc9VNwAUYUDOf3
Oco2TjoQxNHmfrDhHnV3+U0euN8NMXazzmLqLSt8u41j+mNxBJZg3uWM9q3qqQUGlXntWjTpR/wj
V+8C5Ys2tlTnxRdq+2+oEZj6+K1/s2ovPbqp4M2W4XG95iTjLJRk4itXsYa/naCBRuE26q+ksfVN
cG5cs/6lpkobH6oKBO0ApZ4KN+jygqfeP2PPVqE7CL9uZeeQlj010UB+z1vJZMbQSk/j05XZj6Vc
fPMlj+SMcDuYQyGIUr5NG6LwGCSFwYtbvyhMdWgEoctH+ic/rd3dUJDbE2xHvl1s++RD0IjzfAOx
F/o+sm1NX1GOu5j5lb2YUejsdlgZMO+UGQTJsLvB5Ttu8BVe/7GouueSRtBaO5j+xRyM6pSbBmv0
lFwt24OHdNHWDWYZy2RqcKbUrpAe2kOQSj3FeRrw3vjLXG11htzSLz/7R0YvOKEKYmUQo23HyzJq
NEstWBRvUxn8SHptVo8Nul+LLX8fBk6I/TnSxan51u8LEJC7V3OCh+HyWIH8NZZcs1VJwBqwgjA7
Qq3DYIwEnYzKDB2ktDE+6IP2o5TCiC/ar3w+oRJrLtv4WmQoO6vL7N9W9pRLjs6QBwo0VT8YNChx
Ys5//Eb54J65/mSEexltBGs/OXwwbBG4cbkiYL7vEAZ+JzCpC4cWObrYeJvFPCGIXMmUb8EY2JU7
AoqemRJwOPyoeteiAZ/75gs05t/m6mLS4PjurXwOFcVh1e8xHcav8aybm0SufYBRd0cRXwt60+yC
8DQ/FN1mtNzl2OeLwEIXIhdDNQ1pZ9jkTNQx3IA00Z2TZLg/2W94WQgbFRX6xrVGC1XQoUSrzzMD
VCqImt5qbcYCFLMpd3wsScwfTUNPGqWvixkLslaWhNqYxxXTxJJ2Wmuvnzz3BPgbt0Gckly1uWo2
ZWhDuHyqC1BFHjTVQyR0/nvUyeGoRNVtTIC43hlYMlQaPbdRRHsWfv2e6A9HNVowwyw2PMP2oz1v
chfgB+BtEBlj5ZYUpILrB5vt3hp4AvIULNJ7iTiugXK1X5leSTr5vkCU+oAzxxAXlR7Q0xjA0PQ/
nsxZmctDCKPTkf61PE8X3qqep55TpFDEWGg4Uksj5x3EwMfjUYbMehixPixfHKBsvrLPkP0+gMrt
JzoqYCvbZN/YUlZebv8yehW9rVRMiei6FgljD28o2VuZdVtQ1RIq1iAuRyiauWsV++eNTCzfHJtt
0yTgqxJH/qfaBTr2s7EqpHEdpSfKhkIajkmWbDH13JU8QHHG72t5gfq1rCzd9hGI7xrgBmGFMvNL
uXGecfJlYQ/Enka1FRbWt7LiFk/t6xwypL/0eDeQ3dzcQIY7a62C6yp+RnjNjCp8MlzaurpBqNL8
mwPDFO6DIX/aN627JDC9X435e/VY18WPo2+zhIPMPFNe81QNDdeHer5HIr0DZvUQ0rH6HDyIBR/l
8dANTOHLAca9A4RlD6rA+tN68UZD/mATzhYwVavlfStEsbwmATZv+R5kFHK/jCJ4I2iNWRn3WsKQ
Y4lFtcJQ0m6FhzWHYwln/kY0wOueysmk68Rq5BtFTWfWA8wow+dFN0oVDeGHIY3+uP7DluV2aZIv
B5+vA2pzBZgIvXc/xFugTrQEqU9qnS1tiZavyEve/trPfN+wFtvSU4o0F27umME75W1NEw61KDsh
eoT5zocYlzNHVZKJfzrVEYetxbbE7muJLtls5LgVXaZIouaFuOc/f2epo77L2dmAcFgQ+Q7r5usV
7GZSDBPkpP0SNbGp5NMKCsNdOekfWt243SEM11TiVL26NhWlsTcH3/RzP7uMrH9wYbKtgT8TZtbp
ZuoHMrI45s08CyRjPHJN5VLXKc6p9fMl4tLGqGzdIUiVQbz+SI202+iNjMmPANJtl+Q9VwiCL2uP
2EKxJ5LXAxDgHcz/mOgF+lc5vz+YuduteGWTQmFl5xQA88ATJcPzmeJAnbVrHvbtHCiTNjMvgsg1
rMnL0BndS1R8y/QOQlchNdSdqKtYtzCDU7mZ9XZOrnk5L7j2dvMEm9xMtbE4YdHk+hbeax6YCLRb
hdvbQ31wNMnw9m9uhzMiwIjXqENuK8ZOjgo3vu2lfQGvpukJEip8UHIyRvI+OLk1+k0b/QxkMrUI
vV+/jyhhDFXvmydiis1gxLxRGLjg4uhFSpfmfC2YIVZVnqfky4rLFnP0X7M5RNoTDKwU8sMnadMD
L4l+VmH5aialARYZLmohS/R5vREG81Fk1o53ueaAHqCOaS1p/3z84jW5fKHVFqCrpLpbkV7k/v/d
91YSuopJeBHisFtUFgK3zX692ylevJPamAi4AOO8HlH/za1XWc0v833pfRonD89lsCtYtINp1BFO
PEO8o/FXxnqwbTNy6JpiRHlXT4yF2dhNO+PG3NclU1QMdYNAGIhIrCSLg5Y7LuJ1JRWFfsSvwBq3
SOdaF4HW6B78Yk8owCcU3lzQydT4N8oANhKKxICaCuZq4iIWbiLKBOG4+xXkwW+ZqbmJFampg12I
bn+lWqc0fikE8cVPKWt9GWTaQceq5AV4OHKdHfaZZr1k/62/sfTQNIj6yBp4ckR6NY5PDxrdFvyk
M007Yk2vYXWBUC0+VvZvgq+Bbs5lYgIRLhx7t3EsHWl848LlBoT3SFyM+GK4hP2+DuwfBL9Px2Ik
sKaz0sokARDINKZaGK/zxTra1+/Lt/3kMq27yqL525YEZgcj6H0MdmA46vV6a49fTJKQJOtiMCgz
h1YiVMM8e88Mxzy/2FRNQQwbwOjwA+V9A1LNBurkOVGTZiJTGyIiBRjJX8e1AxBAt16kuFcydjxv
xGf6nOwabwEp0LSwvB4KaZ3gRuhC/7CTXGAnixUmOcVjyqX5yv7Vo2//22l39pRXKVY2BZRmQ4hw
gwzN72dLUCNBgS2rSDJhJNUKjFDLfozg1MHf9XFsrBsUTpbN7DjCw43bmLYIq4YQ+IauD5d4Nl1t
L+Q+OSaKWKfxYwLHQDXTQYRH1iEfrWa9ljcVX5mDfb8ZGb3nHtWHDRvi/FzMKNMfX+aw4KEyf1Mx
Wcbr9yQG1TIEg8H2Qo9Jyo5TBE5bo7wV+BcSmdjI0vTXhKZ0jxtRwbDO7ERsRgUDfBzpUl4+NqQc
INAcWGti42JMy3P+OTXIP9pHF+dHTGqDhxUGKR+hx5BZZleH0i5SH8eu7tJ8Gvf/2r5DG6RdDq5A
noIG2Jkab+9FO/+CPdLl+H3T1x7ovn/pZV2QwQC4Mo+J9Vlb4AdvCmg+dRFU82LE0q0EP+iJSPji
VNc32mkzolinKX15+hJilL59pjttZ8MX0RDi5ubbaNlFf4rYcSdIS1WdpVd3fnMB8wrPqp4Udyl8
E6SF76L9ae/Gn1lr+rsszMNI7t08XJDy4ITSdexycuOIpzKouR7ArB9pQs62EYSiGxkr4qmjwU8D
EJYUeoFg6lXXetkdlJrFuhCIw1HVmvr2kIdLN1rMoiPLmOIT2AHLssfJ0zCh+34KxqbIvviR7+Zk
aFymP+qOJU/ZeI1udtA59JgIamLhAiH55FG/xWZ4W+7lPls0AksWDNj8/EbMlJlr+kkVGGKBTTL6
4SLKBZzJOWN9MvqvPNY8SE6lx5oCWu4/Nx1dXqPuurdLiHYDCQg/A63lYENwabKCZAn4s/OFkWMN
RNv/53Vo2c+V//E4qO2c7xWLrSKrGlAJlQCdPI9JFTbylJe+BFlMxjsEjiJ5x8WXj1v4fupIMu2a
I3HSeq11bjcxjFkT2JkBH9D8BbEM0dryvBAtmzsNaJMsc68+xBbUywx905D9f7Y5OTP7fHen+ksX
Jr/+HxD+VIs0DiNCe4zXJQv9Zo8+VrAU4ZPRambCnWZ/z9Byd8zFjtAQCtdmqjtHBNqlvaSOgovV
tH8+Lzp/v+/f8Upuwarp+azrPjYmZS8GqbRZ1HUMHHk7dPaz6Q7NNE3893EHbfj+RlYm6E5IvVty
XMj9wgbhg16s1ypw6Orii8AoQSpers5xpK8uebK4Q9FxMOiZgwejoVfROJOuXSV0vdVEI2JV5TDU
nWKPxr1kHoPKPEUi7bYfsd5zarR6S8NaVW0bw+rFEkirj/VHYmJzzAPK8ALA5hirJfgQj/qDbUWP
CZOby1DE7LOT1dnn0h/iGNYIcPz4Rr4u1nFGTZaI/fnn1kb+4yZQ37JSUnW3WhWz8SzQxGvIyZUD
0fdGKZ19HDpLsQMcbzQug9lDVsB89xa/EWhUfHwJ0sshTlrfAwgPdFB3+j64xXNrWjlLOpIjfct+
6GX6dMHy0X5KgtTebmbC8tIxKiCStkeqQ2dQaH6xHUEAnzYJXtSdXP0qsgU3MSqtQeT3sbSB3yAY
zStwl9o3M2bnvNuMAfsXIeTsk2aL5K5XoML3BISDToVl0MkB4fV/8432ZW9/Ou97toA8Li6j/kBW
srkRLmyzD1psSoYZC2Wd7Q4eRW5VX3RdLtc46rd57XTm0Gd55V9eYWSw+yZ64OetN+/HbSCp7Vbs
KbxxHmJhrhd3rkWrAfoIxROSZtYhQUPmIa2ffJRSozYMeq9++QBYvdRMy5G7Rlf4qkD2rbodU/tp
QQ47XpvKu3VbzB8M/LLWzeDrmMoVUpXKpKA/jm7zDFxseS7jCmQtbWvYZB2HofcFf5+m+30ZKwu9
WBAWce7OGEJqfn7wJ/bzJhjcGGBf4Wl1tbf8dJmokXESnGVArCVENccMoq/2UTEN5elxcPeApa5F
a7XIBlrbkdm+a+llsNkDqrYOJQpkNDf8ZVAwxlFD6Qn7oZJltqNE34AMHCRJNIEr4hvg6N7HAto8
wiRP5JiM9JUsLWb1vffPi9dAEWFBKSUvobgkVwfDsIdy5gtWV14phlQrX4wdYpznUWoYER+eZ5Du
JX3bWWyK21ugCLCdIWuLVHRxgOXpAQZ/4Hi/GMOnXlbBQgoiURuJtQNNMiCvv89m02yMnBSI/3cW
xi5Z5j7NKtRJEdhaCXj29eRcvmTGJOUFwqIs/zi5vo+SfHAaQuBsNtY1YdMB+YWdSYS/3U2iskg7
Z5JzGzWFFGlP/PnKxf9F8KYsSGekU1gyVKRVR3JbgIC1BYETCbv8eLDH1E7/nW6OYINOOnOOJN2E
viHinDGTnapxFnf9OiUkQVUsie1hTiKWXi+Z+Ib/r/dsqm9aXJGOO+oPiK57/zp/EmTHR3rJ4slL
j03Zv7mP9+HrqbBTlqWlze+We/34yJVIRwI9r9ZXNpCXBcgTawt1v93xcGyi2yuiZWZ6AjApFEI1
5qVw3kCHSNJn559oD/8qDPH2Zn3TDos8ryNfA02WIUMlw4FHXXFb2+o96J2kOPy9DNxMDTmHO/2D
q1M+NDsfnJFGUNgHV3goLU1xQfzh73sWMFOMDdkqX+11yRC5D+7YT7RHhcH1Xdrz11AJaWnRAV0M
pxd9cd/3nNf0bISfHKQsI6PM5WGMAYOyhzbd1II0koqsyI20sPP9+uPXdlo6wM9rmwr0CcOtBN1B
ARrQeTx00hbOj7qz7hE3g/E5jSXXgJf2qVG/pjew9o8eJOuDcKM2rXSSZkjRKHKjQ+OURxlqBAhD
dcwPcQ4C5hiil9MKkZ5BgEjrpVol/gtJ0rR/6lWKnymE1uWKrqPqVPaDnqyYtuIWQpXlJcmAfFhA
XDCnjU/4dMsUBOU1mO0n//rBkABm82cRXciPMfvlIbxwmgNWJ9tXtiUS1tZ2jHxjKfZK/9AwdjZf
Bffo9hG3nXqPEuociUeWVOL6KhfBoJWabh1yP9brSX29nQuDGM0LJboYZeAjGreqTGN79wJqHkkf
OtSuhXmXxAa4DW+GHpLFYRG2fVq1UfX8O+PlU41Rjy19EwvsEgBbRkQXvS8ZRp6gQp175/uOZ/v4
QxTuYMTkbVu/7feEEU4Yz10Qv2dEeSOVWRDhUIheefdLd+1Dh5RI1KpBm1KiMDOqorj62Flr4PYo
bx0+LsaQrN0IZ8q4tZ2RKBHzCff3N2P4q/m7JaZrzkty5P5KyCAOPlRWDPHyIRrMHS11p4zt7Rbx
W5QH5N6Zk31m+hqpGJbWveFcDI2mwkqF6iC/ZIBW9aDodtuBrikepIpWaTUmERDswrU8uvnEFIVi
RdBpIYsn+tjSBqt0l20yxpftAoakrRg+sTI40a1h0r8o9b+W96FWXZptTkFqvLyI1fimP2MLrZVk
cqmbX5s1yIIBG5kMr03XIIXC0+MovuLOc4GLeRnIeELD6+i++6S5SqFGnNRjg2veeNE7Bc7HVTqL
Q4gRLPCPyZA+z+iSoLvLLDSKlgQ9IM7zgn//AC7i3JR1jO6YGqQ78W/0+5E/U7B8uv5FTQUuSwZE
J2wS4/c3iCkGEU17X0s/+V/D12eUQvEqBRWKLrK7ojmhIQG7CJt14H6UlWSHEapqR/vG/QdYmdJX
WY/1ipcLLQWCdeCiMcuySqQayg2bRGr/k1oIehtGqGAPqvFX/BelvtjSe304ZY07Tt8jt+QE1NCS
p2HFyXeFJf6Pamg3lifEZlKS+ak1SqUT8x/UeZ+A9lftRW3Jd4ryCL4fhwlC/M5Fllce4KqvcxE0
QrDFF7pZlDi6vr49hGxkl5ExjDD4IXWKYMFlmssYQDt+xP3t3HROjoXKwiujZGwyX7vS2+IB7Lrp
aLjlUOFoVrBFsMxxVeiNAi7ujLkYfxWErfH3GAXrCmBGhE7HXgfxjEyX7KizyFpABX9QPlhbqrCM
l8yck8gxsVYOaH83LHLpHbcwlzgf+t1WnH3dYrkoh4DY8UiOZj6KlGvcLgSu6VILAFStFUdQENE2
JO5qp85HHZd+AKCTnmDgm6xsh5OV+XFxMM+kg9oHh5nRwoRGxc5cvkKiG+cg+edpc/FOwbOXd+dh
j6sZHGUI/C79DuDExpKcvhveTWs/K1IwzUJcSJ4vkdf5R3esjD504MEScIeWDkn8e3PpkSTZo2dA
ByKtQmFWFuEf35vOrxw7w2UYEd8dfgaOAF1m0ekuYiAqcJ7yA4QmsuvN+ReGjpQKpHpcq557djXi
tGaMV769vt3TKxzxlL2P8f+JkukwXzG1CJCucpcmAvMV4GaWx1FsMfLiiXwc8dGXhRG0BZRLOaYz
0b7W3YpS+g0WAF6ZOCd5olJsVRy8MBQNxYhbai0M1KpCjKr+1pBNUeotc0eHmlnmywyzbXWRPR5Q
5MAq9PcdTQwCIj2/gutYzI+6zHM0y68KpFIhgtSNp6G1CKJOlyRw5zc6iFs12ye2kCFNfIPsFYEe
XCQbJdJsE1seaH2UhBUy1EL4ZQ0zY8kn7Uuryp6YkN8MTprzgFR0mnXuEIUsUhnaVp66AItXVnVL
QVia2zitwf6xQZIbiKpybifExTYzkuCu/H3QBI1fMIoSR4TvK9T3FwbTSb5e/6RAn7dOcfp/bLiB
ojM+PCB5ubDdlvIXsf6Hh3B8tRYwg7SYxW3JS4OOsqY2toO0VZgDi5Eh7/E3yOZ0R4W9b+sop6Hy
1fSSX5UlP5lp/rB6RRTBrRMP0Mfg1qaxxaiemf4TCgumI6sV0bPcCIq0XnlYGpu+zpdvPLyQpxFc
TdhKnCdmqD5C/BlMLGAZ+zEOs3I1HxxJlVNAcfWrLD9Ch9SeSDnU9EMUKd6vyBYryOFFE29yWiMM
THC3paYNF/4v+kPu1uQDk3Mk3PZFImBbb313bdUyNLY1dtNgcX4+k0hL0xY6ubOdGjKzi3QOMkTf
OaoqtDwUMcmArzlykSf+jZg58vMC8IEfu5u0bYJiXgluTNlLvm13J/vRFMuO+2TKNJGlUQhX36yB
2/EwnAJ3HANOeKZmVnVqGps+/YGeAwfjUufReqKMyyGpz4Chyw9PYQ95dogKMoNb88l+NzMvlBFE
d7HCu4TWFqoKHCQDE+SzULLb/nIMg0BfgzOeL4PyxWwB0PqCALJfpz87jPYKLr8K665adTxH/K+R
pyEgk74N5eVSwy2c5ytU2EwWgGe6O4xUUvA7R+XNlOuZpChPd1e6kpdBXhvbXEBHOlqqDGjBdalU
9vKJ35t+Puwm1mJTaerMY5Rfb6gOb/FtHVwzm/KAjo27BMlAYnXEz4x6YttuME7jRHKsEekb8LPp
nqmHUmULaZHU4X1DV7tZFEsh0KJh/zHwD2V9aI5y0NosOSRBZtD+ghSPlsYcMeLB0szxtCFlNbAQ
t/l3RarkEOsKKnNABs4j+hNONDDpxnqYxIEcmDihv8rnNFhGWuDmMxVKXrhehc/DIRP7otome0za
mZUjA+s1Keh7ZbN1FgCyhGq6AUY2AJz+I8DN/jLAZCEbkIBKUSWxr4ipSUVDjbldmRkH05EBKrla
3sJSHtNFj2wsSzg2toVSGSMrfthFzX6kAVuhhnHnHeNl7GMChQ1xQ0TgtWhSXbmhWm47mH6wVMQb
p1GzL04ro5/T6B5I/wmclE3I0h4v//c69eZDhvzfbR1cZ1HEQqPLlG6Qt5HKxXxLk/rfhonHNtc7
G6as5rY/3VI1wS2D5zsBnVmvWNpbKQQB4yiSQRR8sb0hKe5JW2Vx7ok84c8103oUbvGzrydd6zUm
iTa5uhkF5MQjs766ZZGgKOe+Fc2lePh8cZk1FwJTNBVgh66+TdXINOjJHfC0A3fTD7lGJNfFMkMM
BHJZEpNaMbG/9VlSjTue8rgnnUdOd4v+Y86Xfr/B2+l/4O14oRhnbZ0nNPn7lNdRu8Yb40ul3+gY
NpGLER0hWv0r+NO8F88CMzrBBcZ+tp7FlXwEdk/mRVIZrwwWH66FNVMdqrjwoGEH/zUorjN0M83U
jjLCZkAHt7B17fqfSIfcB0F7Bx9HmfSwLYBSr+2p2x+awzGbyr9qegL0gNB7+93S9TX0oY6km4XF
zM1e4bu6kefBrV8UCVZD+8nrdOMCnweSEaWk+5mk5HzsKM2zT1slghPPhR6I+4grt4nUGCpMdclu
d9wr5g6v/DJu2yp8ITXQwmVWf922jXY3bCw5In7J1Gyg5j5UtRTJ16JUuwtShIsKKKFtLFrBMXBk
fh/gBiGFqEIC9KZEZsXOo1usygxdBgcqCcAmfRoK828h3MSQ9LKd7kqZECIQk03ytkCoPuUjXn9t
a+IvNuEgBqUcTAQOu4ZqtArGn7l7fdfJWITYKClTqRn1TkfnzqZQt2r5MW8KG4CyYHviy6uufJK+
SKBsXC/hs9WxyN87RYODQuyZOn5EweshOdYkYaTRXGG2yjAJRLeWCWoSFX/kgMmELCrH/UUxhc4c
vAOrT1/Os9uXoo0boBApwPDuqOXXYRehCXZV39FG4HqJs1LsEC95xSVUiOidzhZ8rB438NSHQW3E
XjDkugD0neDOFPqAxBoqGyKa+AB0+TIFKUJTM4izhM7DlCb+xVp79oAHWocDAXmbzQGN++5WVecT
U5Z2JpyYqkIMuwSOt2Jl2h0Fx4RZ3JFJnWTEt4LsIKIfHuToTrjAs7Gxo3SM3qDD8AN+WlfCWHhk
N5jHiX5pHmk58ehyZzkZIBxLGtC6qt8l3MEb9QjUWERqVWtfokw0JQw8x5Klo8cNCTM5MnHIDrq0
QacOhyekXeqVOBY9OX8ChR12vaRPa8TU/Yx1v3ok/dJKeR6xZTvfKAmNjJzeafubE+tifrr/6TpD
CqCQydTLQ5xgQ0OnPFoyaMjQVe8sOsiOyuKpF4MeXg0QEKAVGY8lwljxq24Qu/ZWvVfvYhkYWFVJ
XmoLlX50222vXjBIkHe+Dp7OkslheQ38fMY6BvVwErpeLukm0RUiEztXMkx42K1UoBEsVfsn28xC
1tIvg+2PQbWuKBkGRzaSFTvO0wjy2QQb/n++tZiHd7bx3QVGP4d2Y9nVztKK68ZE7TPQlygXUlNA
d1Vw6QBXiwDSiX1ZIo+bBY+O/c6Ng/Jow+USTelv7jFl0P24SbZaCx2uAh5ujC9QTqgpac17ZPXb
fjrayTCkEKTB0upTjhI7Glkj1L3UYSnrXuV8Mj6HuUC3MF/2PUx3DQag6rKiFmuD1r9s18JuhLHS
/rpbhrp6vhPbyjxUQLdkKzQlvg37OZ3Va7/A09d8wiwjquJVNlyhIGNMTtg8ygYIMDq5GCoLZdFV
cp2V4WfbWoPAUfjMk2kdU1iLtdgoQzWyK56+VAEmbT152/H2YEE4HL8vZX36xkALqt3fiqH/ULXJ
UOPCk+O0IWzyI1VhjZvmTB8PjR6t2X/mEc1ESljjqWkrkfZbtb32t/zHSA+zOUykj+tQeGqxwLsM
CNWadlG/3Li2OzFig3wbvVCg1JB887nUBSZLv6GZSODxh7BdJhM6v1YkkPClxOoD4ScWw04DSO05
8T1nSwcmANCEGGLT99UKaNb6pYX9WiRiL77nKVEE9VdZHNjtnW4+gKn/7oqVCcjRQVac6aCqp9n4
ZkO0xLSl5mNSVwyTGNKevMoih6P17djTkO+4LitWTnWGidn2W/ex68Mm1n4gyTL01FZRtcfLrqnL
C0HR7j5ET7hyjDls+mgHngzCUW8L/g4VGyYeBjhwgwFpXZ6XOQs1T3IW1KWaHqQuFl+tJJXp+oiX
E7p/dbiqjwZmE+djp0+swPV9B3v1rjUkzR5AhUe7utUz8pJs9PP+qzyodj8sQZANxGcjjbVm5SJK
2tTsSA6y/T9WgNOEi91AVXY69Zj7TRBR5TTr2p5/ysbBbc3MrabhT5HwxmYVhPpiafefkiSpbsKN
pdh4SIzY9eakISGxqZ6bmOIA+xlUJDUngkOomaaPCadOR2DNSsxM8KxC0297DIoGHevp/3xWbTSA
itZTVkCwXfQK9N0c5TLKsGnOEsFkHC6FA2b6KMyrMx68f76m84Filn/z8AFwcg1punrN6ylb6lue
6VcNdmLXb8l7n+izoKboXdURTRsM4qmo21HMBYdCHPg4q7yA8HjPjNbNWn7ZLbgj2nGcQ0xg4aJK
RgGYpAnuOMuMgGvhAmGkESkWrKXJ4+JQRkhzfe+5h1fsawA1bZU5xFhiXWdtSDMztR7z8pJoqNhr
wDaQv+YleCbvf2vEy9sfIAn1DG4yu6bcQiThx2tXA82z7BvwQA5po9iz8PRyyz4/56jY1fkyJOVk
FCS+IgapmcWdoXdmrD2Q2x5donAEFN+qLBL+YMadYI0Y2n8HWcK/k7k1vhjGZbDmoT7+RiW1AjcD
AkSafV4fN4nOnx1y7fd8ud6FEumN839wvEs6KgUJqZk+SV3YqNz7t5SC2fm1SxVkzBRidXndEmgB
+T3PLIiDWCOJy6f/0ACdSCHio1/vtrEH7ADPf+WOadlTRzhG8ilHpFXwhsekhJ1OQR2eTKGIUJQ4
PqmfENPgauw3JqLsXoQpPKRPLH4t/CQoZ8/kk7W6miFXlAwlJ/igP1eYxL3VnpdmQT12x2IaUdR+
PWcnaNgo68x7cwS+RdWo0BC4GvJqEAhi9vcKo1Mo1GQTPX8ha7SRxrd6jAGCzn7swPPtvB0Lgnrs
Qopbn1QloccbQGI2WsrpH8ntkfIfiKBW5sFBvn8D8NBOBKYlargaKB1B/24awmZ4XYGrF/ro/ge4
XKhK3hTrxaeqkMkM8Te6eRZuc+KDGF5xaaWGdN6cYTlrVsb+rdoKLlMZIsgbEnHvlSBSPNbuuaXu
vAhyvpM/PcEGGesmlzkWrLvmVBBeg/d3TcmPyL9WZqXIBrKvKIwz95fzmjiqrT/t53+wz8ssfHHp
z5nZ+v5uOX4MUrm5iubQmQ1bTi8Fobwxqt7j8DqQn2rkSJMsW2YbdHo29Zqvcy9/S9VD59hfimj0
ZOg6aYo26rDTL7UvGq+XkFywvp8ZuB7+oX0Cqm8gCiZHVAwLlM8OnXlbPVv+/ZIkQypw7ctBVdjw
G3YPmMX3b8/1K09PFjvTyk2G1W2/LMK08s8khHeDzAThTiHn11Zn0GJP6cpky+OrLYkdILro9tVT
Xb43HCzf7fXAusehg5Trmj9jnBsT8UekTdN8OjIIwJU8urkZw5oY0krSN7lqaxO9db9atWk1/C0C
mV95nvqaLQs/fIe9+5WrS4RcvHie+fkxnfNoL5xh93CyeIEmBw+29UiHpFRSlCvqtjY05A4u8NHN
HIDzg9k3hZzi51zmMnbVKChVmsMygl/XtTL4YuR9TZDA2unzICK/1CM4OwMzoCHxLBkv9CH7ulD5
lUfmwMWrz9TEjvo6j6R8/Bs7bBtLvEzs1NrN5ZAvABUQ8ABK9lrIJENGBi7IX6sUiIritOT4vb6/
EoMxhjGnH+8k2wXbcG3uhuyGTRikgld/3didES2LoNcyFl1xP3jqWCT31GfZqRj1tIURqUIEBQ15
iRjmeuaFVp4IHOXGd3j3UHDZSMVqfrOzl5BE05TOCK4dp2u5n2CsJ3Y25UMYhoiTBUsDdl3y89sk
MTJky8SbLNw+hqud61Pvt/p7BWtzy4+pCNQhA47iPxUIJAXwbowIX8t7Sj0fj8qit4/J/Nu+J23z
JeeSxYvTSTFnIqfV8vWUmPks40kuDsVCLp3cNFlEC7ZuvQ8nCcBcJOIg1U+gRdHrqasoQRQFebyA
F51SlaWi4NROVWrfyMK8kLokt/F3QC+nJ26Pvd3a3/SuBHQMeAZcp3J7tp4dZJRusu5JjWmBJ/jJ
FdI8XUy5ZLL3mcXrx7MFtg6ubxWr6P47dtgHQlBON1srjCJS7aNigXEoSmC3Itt9/Clbih9VPbQe
jCJsIGO2UUo6GWVr2TDpo46EMOJHnm6rTTg6/mdE6kP2OSxkIRd7mpiJnQICvmj9iHzVEOTpQqY4
WRvKS1ULtFFuWqdx/1y6H+YkDctSEtRp5/F59lflirW08MwP9q0ih6hLcdOw0HPbBlpLTAD2NtT+
hA6Qbde+5m+ZkZILV0jRc333O3dy2Dgg4HWkIP0Lsjo19ojRW5Xe1EXJ6VwPdHpnX6wXeTXHpHhx
s8hNYqX8Xvg1FlvzS6329bfV7mB0Ypty44AENcR2wHPQ/b7xb/yy2UcdrTN8747250G71tiuKAIX
FcVriQJsExv00b/hb+kQp5AzbFgNSOukEM/S866EoLKNir7lfxGlLtuXlpmcM0vZdFgh3pJUNYzx
zCtPOoUXMGjUOkt+UUfB/5yAgBn+WX9cff6ECdZuIZyMTBit3o3m1ZM1IiW/wX4B0v4Y+uYprIuj
u171u9bUpgeARBeFB24kSsByclLy2mIvvzYPlxekdBvNM9lWk4/eDaB4xr6Zlxsmnt1tWiBm18Bm
FpgsYVq7MZOhfuMI+scNh38U49j7NX+xXXj9BuehVGa6JrvdNpfkVOHb3O7vcK8wgQTRiMiOOsE4
esYuzyAao7Kuz8ji27zfhQXiXAzkuXDPsS8i7RsOwjr4mHZNcos+Ns546m0ENQ1J8EPhsBP11t2C
dJ4XRgotnap21J/2imJUDZiouvKBA8Cw1sWN/Kk9Cn56vZs0XSN9uzrDE9sG9l3r37weS3Xr5f7r
txZjumORSQBhRYkMxHNVTAkKobqAcwmSfLdwusKr6h7KwW198SlZXfCJU3581sZ1hR6Arq8MUrxh
tMNCkhDhNtcbgsQhnWSSYw2ruKX83EFpNlgx1lumbo+4SHM4S9QCjpveKajNPzic2mT/Y4EEEGJx
BllpVP4VV7aL4J1rFDGXrqeEBVeQYqdrln+tK5ygLJvS+YYjHQ1wZ70SOIPNtsOh5KaZXMqtDAS0
FKxCziV2a0mapelYx0jaxsHSez1EWbaAYBOfl2HSGtzXD4hw7DoO/IGUJKR40649AWcGIIPYEYh5
I9hyRU8uM6kMVrzCdfXFRnWElrMAxFq4P4J7lhM88KBLW4yPj1nKEfHPAZ8NmXXTDdPck9xVaSwt
hvyfmZxlyJ2Il7MgLXZConhS0NDijyRHmknQYHcT8rtccNd96M6bfFXOQEHSHX8DXXEfDssiM886
UxumDqWLgAq4TVVR05/o9xD1TskvR+lDXns00bcZCfkKUu9hC71ehWnYawq6KyYt75wuLTxugPji
6lRcQBMUVFiwit4Qish9zY3Oau6KX7N2f/lAiuEEllsP5c1Zt1kj4QyV7DfKdNUsb1KgoXlZCgXL
N038DEgHADy3dhEFa+0/yTbAYhwdKWnnt/X/eL7b4Ll+OiqLi8fhxk0IblSGM8e5QuNUuJx9g91q
D9j2XU2/B69fOmZ0amuaqLocCicTFM6DMbeJUZbohao7ufb5eJNI1wpM+tUF+LGe9gGblYwiaQyI
q77l+vRiW9URPBFZy0nlxF6pJn9jQUVbKldkN/4iBZgSo1d6Z9gU0CXqpa4a/BKtgcdqznOyoB1m
kV+mzlw9gixpGIS3Fy7bZoqw8JpuNGux9IW4X+DDkVwYvsLaqVlOgPpVSYxk5rt47wizN94GQeJz
B8HQzJpyOUW/OiHoz5FNcrIQ0BJQsPLxiV+pcJEX6yFXoI24KZVJuQJr+GHA34bs+GttC8b6QT4f
mgaNxM7UiOyKLLFjolDueQ78a/CPjkObK8kyuqOEokFrJn04rM4yXbpxvYCELD/J0BzctKgmdjRv
1vkKvpMw54NroNTabL2iVcccKURjoYI/fObzqr4Ris9wZmRQovPnhcMbVLgZV86fqpLRQZF5GlsK
buGRRP0lr7CFKH0xatYz24Sb++Hg7xZLRH6SROh7to9cohxY19H+Uou2AJOofLgIgy9efSdGDpvM
reGQV9VNW7qrBDnP4S3+sDJApQuuDrWm+9Su1oNYhoMPv2gW9t0QvMSqNdFaia+HZM8qzENWPP2n
R0uZZqyi0zz5Bss9Z1XdGjcT/5uLYwgW+PcCSD4Le1AqzDPqd95QAKTK+zgnyvyFAT8dJl3HGX83
F41heIL+26sKN+Q3+pSc06/XrBgTkcCTmcG9To5GdmsJi64lIqswiTo6c5dfMSzbko9I2z2W0wB2
j9MYSJx12jDs/vWyKIpMoCkh2czaiSo1neyGgiN0dv2X/DO1iyEO3uoE02dyY+6YvXgY+johMV4o
FiKDGoSHVda3mZ4MgdvnTC5gKCt038QyFpPrvKovmtx4JB5xx5eoqiX5UcN4vRmblORvaFTa2QS1
UbhlIVYm+K1K/E0U6QJCZwpOiBJJX0xHyI4zGUj/OOOFqMLG0ZVnOKcwvEYxb1yXgHAxXGFobIak
f++awoTp01X5bWeC+32nuQudOdRAwjRU7sdF0m6cTRz+xe9x0NMtR+8g7NwcwbdQeG5lxb+/dot9
NvJAcKsIUAK2WmvUfKtUr7sV86XJ8LDmZlWIZghDIc8p1xEkpVYFn8+qnBaubjEuaEWt5VbDpWyr
Nj1VTxD0Qh0FWLT6RRNfqcMCtMleHq/AUOpbevlM1xhC3Z3/4HRc+8Z/H1Vtni2l85chJbkuI47C
ZR5sTnPzH9E48G7y1YaNSLQ7fEZhvGrWXxU5iDQCdqI6t+ufTc1mz0qKD15QRcCcR0GFnGGwpZ3h
tzoYwR0luLkyjpDbEWRP+gBHyz4gIvpL2rBPM2W/TMSQnf2vFOLSZ7zGpgCbdn1Vov++uqtOJhS2
vKve23YoLtgzyeVadNvr6lNvJU1B86NXLLI2kLhGplUI3O0KDPNwZtvKGUvlW0nEhfYbW0Tlp1dC
PWdtsJpYKrrKnR9LsshHf0LIOH36jse8qARLgUyGapscAntkPfd2zrZg+5RlErTj3Llbuh29Iwe4
85nybtWWtDEXFFSauGBlP2Uhxf3iPWpYY9Q2eLbq5PGZqjTvytsjqD7eA2nGHW0Di4AFAHpWONRu
qBWjxyxHkKc+5vaBrqzmb8fWwHE4FAbSL2EONI5rlRArdFP/cdc0p3KXvp7t2zltzLBWhhc/LhNn
UERdCoNyDc9aN7g/uTL2yK/XMKljpahm6yW4G62GLSxwuXGTmwk/qbtvpJnhkNpa5DXdMWUiF2R1
h5Bo2kRqevm0uqjFb91uT3+t7aR+MJc42+94qLTC+2jNkZDQeKlHWi8hKcs/ozRlSzgyUqIQjLaA
pBM4BomtRby2P9Yv0nAjyfT/D8nADTdm+XKD3pv9o2o5BWcMo9PSSaahNAwV24QQxPs0aIFc/0vQ
UZ1181wvPDPcI/jlc/fgba5ZZEsuNwmNWIX2Sg9iuiGWy+nynadA8nwVKttYwa5lh6YB4tRaCV0t
lSpRtwzUOT79tHIrD3jx2FFvlhHGhQsXaGW/3plQ+JP0woxlVwxFZA+5Gn3OvSaJlQb9QzWQ5jZz
8dKp0m+errabIgHnWbqJ8Ktvuukwiq56i7TFSiFswUFhyH0GeAI6MPWEj8fxyQ8qQ0wQ39tfnuz+
0hLuuva/msbPsU9c6Da/fli4Qk0Y1GkdOYgydmbIT3O/Kq2UNZ6RCXP4B2elbgxJs5dzmZR0FOZW
GqgUUzNZLhMqwcnF80Z9ccxYy3LGTEuQnrVFnZVk2rg0ZukEDZwYcwSEfeksUXDHYoYBIpsj/GbT
cp7NuMXECzyMVvGBYsS6zB0IyAP4NARwygNfJNAidYlh7MreZDVUaOYNHba3QpaCWFxvb80r8Cbj
t/N0no0OpKO9XDk/Qne3zCJkA2G2Ob8XcN8wWkYjoP77vNeXx+fcJey8JwKmWYmwI0oTRLPBXhkE
IhDG+4zu+kse6tEzO8hROZ0ES9HklTtyooJIDNZrYu/alEk/yb3CDsPCT5qxmsMLpkr5lLdTVz2s
m4Mj9im4q4csejbgRrzNoQYdFjSFuEKG8gMiFkyREgVpnnWbOPaUWQNRiwfvG8RsL99xsvAv6ngQ
Msu0/6g33R7UWurce5wnIa5a6cTTqkrqnjE4kWAahZc3xvB9E4N6F3yvXf2O2VIJg2y6EfMp+aTu
bACOkAH95tIO5kGkXw2TKIf6L1V1eos4BmYSbnBvA0MctvoUPxGLRBXnVcGWB/d1zmkB5zSDHcK4
Gh/VnS0uHPjxcGYFhva/JrDc94wOMtk/ZsPIa48oJEVf6ZfqdM9sf9JbaL/Cl6Bumr4v0PImmoGS
OpZHrBwyr6XylggtukmmflvBZfr/48raAsH/WSTfMdHo4jNIqSV/ccLRg3vAKQAPJ4EaZ+b+wFnX
nhvCyBIaUMOODv7ewmnPFXgcL8o78hZb4L8KG3CcUN15Ply3nQpob8TQSaPtpvVVfooIHVg7dxcx
Ziq3f7v/px0a4tL9lYmyj45ci8Sk856iOkj1G8hc7td5ge1sZ5uIl4HYECk3FmY5sOev1D9VYQe2
m0D5S0929K03A9ueotyFz+EXqMm+mJxsDN38WBkYRuKucjK3VxG2d41XQqigw4f8weYd9HaaT/Gm
qAQIhCPjTWpDOqND21DodoUHmqJQnAFJpy43MoMPDdk+o+cal1p9CABsqp8rU9KchvbYQojB4oxu
qX81dxCAN2M1iStV23hanML+R9tYaiYfpa2vF5A+r5GlpydKiEdyO/I8UhjB04Ea4n+FFwYj6ogN
SwKK8ifJvgf7i3XOoOKA3Fv4JunpR0b1Kc+uS2IqgEyxM3x7jawPSAkxPbIqLjq5ysR4GpXOoUYQ
Ybct/BhvZSgvTY4ZwXcDAf4KSuygIl93VgcGMeoNrIJ77ClieLxFyuGHCukfDcsPwdQ0Ajw33St1
vAx6/yf4TDieR8sMHuKZty6ARKpHFWJMXigq2bvPSnZlA+CMbo8pz3mah7StM95JMIgkmD/zF1sa
xC1pyL2prEhn1XPYr9e3tu1jJqNZfZY2KaKrkSbz8Wnp3ZrNUsepYkJQ/ttSgEfu3Xxb7+7xT+s/
jQzxHYoXWVoJAA0X9cxaeir6AhXc2lV8epvNxiGbA+GW1RDfSGDsm6ryXRnzY9NVMiS5lH1xphro
YK0lT2ViVbqf2K/k7faCiENtmNsJHHZPc5+YxLAIvMdBvXQ1d/ieqDxz+iXUTxSwlhqTDVsdoHSQ
4fa9epHDlhRbfiRgQzwRo4tt387tDrINhIXlrFIVtjSCuwewJubbneVXeYmvAMmoXkzlinC277zd
8QCs31qB2X8p8waDnMYIF9W8NhShFZpo15MBeA+dK6N82CWWRd/gt1a1Djd+7JRu1c6ljGwmQ3t3
BwPaVfOcNcjqgnIFpYnz3lrZIE3LsorQ28ctn8ydhq5aIbVMDG19nWwRwTIlE20HiPVDZKrC7TKE
YW9QwN+wED7a8NHhWtTtWiILqgADIhccLsvxg86L8nOGTJJoW9HbPmxX1jS59vovXHB+PdTfPhxh
bVlqGWKHktbo4RgEry3htl8l0SsbFMxpLkFodDK7SJxXR92uHKXza6HI7cufWdH/uX+VGXP5nAYc
/H7SJsUmAcZucSlB5IpnpllbQfzdd6XfhR7fo+3PSj1S7AST5BKv8RpCyse/EPLhFlfPJrj5tY4X
7/cy5v6Kgku8l4qrp026wpeINVjyk/AzE3uPF+eR7xJzdIudmSXrvoT/3TStcSzSkuPaT+mYDkEt
eceGzH03djZZY4eP0N5e16nZO/6zFO6MEc0uoU2NlMLF6sdcuNnN+TkEBKWM3dnHxAhqzJI5G1u6
RVXwTgtnwMAvTmYN5Of7m4/qVH20g28CuhVSMUp+xTGEcrz6+c/Fe+YqH39hAAhk/ZNMOJFk97Sp
0/tl6T/nWiWFNltTCh61bO/aIS2petqzhRAJVYswdAM80JtN2w7d+7v1aAYkXQcjasGRWs1yZIIw
4Xp79h4H8epFg39Ipsj8rMi2lzOl9mcVXupcCPNOoU6h1okMN0crN9bGmLxs9nYS+CIcct3p8Jnj
MmVsb2WqN7mhTg/Txh7C6NXKDZwN7+G+XVY2SszRp9ZyH/c0cMKSbALJYuTcJcUUwS9z39yZS8le
uNWrium/kfRocvw166UU3HplF1n/4AHBqA2GzJMPxOLDr87ROGJQCORYxfoTp6qlXrC43c66g0Y0
jF8fonoBXCMliOc5OGrhFHQg4OBtYdFcw1iUcjLKLILj7URikGj0KTcrzs46gfgZD0WdyUFtCN6d
mM+2X80m9cYW/8n33im0YWzctLpCyPXZi2IFvNs9T8uwYgFKJVHvf3h/FhA2eLxBr/z3p68/BItO
vUmazh25VHLY8OtfamO5Mfx6dOk8Lufe/Ad6f+DNp7s+QA90S2rQiPgJ3rrUEYeiC/rVpvigjJ82
B1WH57bOBzPFhr5f2SF6R6Nmt4JcK2lSOmk4wWTGmG0uM7DLoVjg/rVALaM6j6kzD3u1wvEJXNKD
9iFRMKy6jKEWc0oHSTksMLAjUmbTxv2WqNhTD7lL5lU4W4rFa44Pm//cS/56rgZLYSxk9OGXL72/
BvhhPdHcGsWlRwmbxhzQ4DgiiAa7KJmuePTohdOmSpCxq8JmTT9Q69zi3pjeyulgM+rRkAW9odcs
upeJwk0V3P9H5E57BuT2rstIdqongw66hXZEIZ6646mfuJU68FIIk4J69oLXnNzLngnhZOVaqzyy
zpmqRCGrrZEvygOevEcWXtb4837pXf3L3kx2qk96db1l7yXePXDUjXcScR/gPMYrczzd32H+ar9z
DvSTXEAhfz9gS/sOLg4XzZ6F2M8lqwz37tXRvdXEQMX753GkprnOcp8zBRjyubhymgMw0yTURcIo
JD31nrroRdvswd+ZR3Xst1DIUouozDmn1i9awmOa5enRwzcr85H4GI6e1Irao4pexo7+ZHPcEF33
EBXL0jUEt5KmDXrB/1fuwHagMb+86C8Ml0HutNxSovNKnXwynAifnKROnjaSaUopnPJofUxMYoCA
emVW5O7mqp9asHOuYRl2A2Sz3moxCol7On5+zkhsoqBVj2t0F++LK7/IlyhYLLb6C62BaUpg+yeN
vUASeGK//dg42/M8sblJQ9s8eHTCsGyuZ2RadnPDFdBONbOfY/7V4c8eIzgV67uphW1or5x1H1sE
hbLEecIfaJNxlp/PId6LUxMg1tF/iJiQEXoXoxPv0EIioKUQ/HWOfd/SYnfbQWcNoZH1Rqtwk659
iV9gtyoRKOqY3ECNHGDrHShYGRCPEpg4jL/PihLhh8dDJF4Gzxm0pZydwNrsdiwjbWAkzurLxFaP
BB0BqUoF7aStWVMhsCgjCrHUeondW7KjxheaPZaOSKqZDSY67vGodLrO+srHyk/SLx7zNEyZHn5g
Jl29b4AmWylczIvjDHi3xNnK0JRREUKE/4Krnze7Fipr9e9r/7nbzThDqKzKAMUJwuSmWlkQ7fi7
0tRqeJG1WFm7PkjSz0eABSRgCzR9TAAB/Ap+WTW4Bcv4Rfp5hccRarX91CLns1tMoebLpqozH0Q/
oZwzBDruL4tqEoIB9C3+ufJoliTWBQU4wJhaTThdvhnlv865syETn2x5KpOWCFUBSPtLeYVxJaIq
VSRvGr8jw6O77wkhwvnxB0xmrCOFoaWJD9nSGXQQ3FCz5ApsosF3OlDx+MFQ3NU2QBhCs9X9U+XF
sEp5WWbUXJckEOuUVdvNYx1HxqVM/ct177tjeBeEZpRQWzEkN7ToQ+DzvstPEeESZq8sZYo8v2Vw
vwxQSkt31ZRKwFHCBd8qxCFBcKj4J1D1cIUJ+7NC/8nS1XYdvW/oFKQ+BAkK3N9yVnL8VlviSygg
bwP0RDF7OpJd8/2g6Djnz3LewLTjODCGELG5haBmR1B9q8QMbA6Vc4p+SB5Je7N5YqR1OJzy4XTo
Ys0YN2dvExeVQ2LxIQcj268GYcTY4qWzAol/OQGztszueKd2hIrY64hnPDvlFpaDE9RoXQwV9DPS
wJN7+9Esatcye+vcNNqh8Aap7A/s1FMWvWUU6CxYVoeEE8Wc7wlc89kMe1BdPV4rzY48Mo5VCzUP
v0vaIjVpNxtqf4PIkPxnfAi0oEgDURqF+Dd2LVG2xgh6sAm3zCvZLehT2orHsZqiIselxgFBOerx
FpnGa9WOKqLwRmM3+GioREeUYF60yIR5hVbRYDZc8ykaFA6TzG8EpZ1fFfluJPCXxFZi2csi1KIM
eQlpUpWZh5JrZ6iR3aRxr/ATNxGn/84kPPr2Jd+kTdlAmQSTA4NaXL+oa5DlnlXVgResG+ycLXnN
KvfWC9S8QfQe2gaCHmkhAD4DhMHd3O8iwxUiEpR1kqL5wDXDmVOK/OrpTU7qS4BE4oOaTiHJlYIJ
U5D4y9qyl1U8eckGpoAUymmkrJ71ew5BqYy3Gwnp07q1LOKXtxlVv3XlcqP4HP9/slNLpVGFwUiK
nfJd3BxAd7BYrOBhBWLA63OeE5FCGiMsNd3G/QzOoxqTWnEWSqSItS20DRFNpHoIn9dPq29Jo0PO
H2Ng/NsEL5dI1KlBiaLhB0CIN/OOE70LzmYBVIAe+iyFr8mJSaHsHs7wlvqLRbck6SlW82Vnhacm
lVbbnhCOkodAtClO74/WFBVh7Tpulf591UYo1SlnOoAkk8tfdpRdaN6G5YHfck0wK1C52Cy1idGu
OwUaSzOU8+mvS+6TZJbTIfqohsZ+ref9lmSQKWs2JwIy6sc8u38fwVgv5hesVQGmCS9TkmjyyUga
PQYUTuaXiL9YjnulDuulorcmU0EHQqQwIceELDMUM5wBwLW2ufkD7CMYY/Q8P49XfOWoj/qtL2Kg
mrWsW/tQmZQHAdoEYpNfnjto0LUjgMhKNMOjiVgL7d3NwQIDo0NC3XovIBRnBh61fSEfhtRRIQkn
86x2GJEVafwNP5Ph/6ZHNJmHukFr3q0aBtrsJwVI/n2MDDLUPmQAQc8sC3ysPpwlua197nbVTK7w
DY7I0TjZTMkabCeMkprPwl+6sgJox7bfS+iwbwC0rSvZfMsr6bZQ2+N+m4C33wVG1ohEfQoXbvh5
d4GBTLGXYTtzylJU7GXmBjZGgJm2HmrdtDzp9CtSYoGVEqQM35lyKAyPYGueJJ39Sg/0tECsO8M8
71+XWznVA3NKzErTvL4XWEejDw2JSViTHVydO4tFrV4/9NPG11EiEPhR0witwE1p8aVkJRz6KHoc
lWN+IgA/jXUCcGFK1/pK0hoQAspp6BtwoEycYNzIhIJQhKlKofPBodXfEVphaiwfYCCc1CwFtGXO
ovjMc0wkREsWGA8nu9zbw7YYtKCzIVOWP0g3DL1O/RNLVTvaFi+uz2RZyt03Q39Dou0oka4W+/mM
cRpYyRbFG/+9WiduWb71cRDuAaLMCh2nN9g9MnoYXHCEjScU7pHZgYBXePNOfTrjGh1Y+Yj2hpP9
rLi1W14+UDLGDtAOudvsf8/vdFtzcIp0uKBcRlwEXjJ0rNQuxpmDxx70Ojv/2UVHV5m0CSqMDWdc
kziRjyZcfpGJoBsTHEyQEC7wlqJVG7kW1eTYiiyxmg3BgcXe3T874y19JZdEwP/ZsaMfgHqaZoTn
Opc18As8SzxjEf2UTaL9iIu9hdhHxJTROnXCvaw9wVUoeNxb07qoBqjNKCRNxNS1smAG9NW5LSbr
LmPLxb4suoryyUiHgp/1Vv3laQZG26OU0pxzMbtpgJU895S/tIOy1ubuJ7y9hdRL7g9McEehMq9V
eHwYENbPUEAfKu15+7QdIdL+QJ1FzTM4sgy5Wi3RqXCPFCEBh+HC3RlvCGidiskTk3ldYXKKRe+w
9WpFHATM8QtqriaPBxMp2Xus3eAaBfalNTpEZnYPovmkO4C1wmqsaEVYHNZnIaq9YElD3goOkF8s
FI5H/JUNr8JxFuxShS0C/Nub3RvDra0BTqoJeK3DXAueqH1cF9JRIcSmrJd3AxloF+73Kxhw3Ejn
g/HiSQ88hZVuRTGLAJxXtNm9TNgzjAtu2f7P04d0ra2GpmBKRxROttZzLx4tU7fUVblum7AVWD34
tbj1+OALeALFW0lUFnKsP4rMn1fTO4ait86RYbiErEolj5B7wJQXCHuy1qxbPDKqwVQBTjYJtT0D
HPeNosoSuoR0oJj/oBaJGssf5BoZynJtfgQAi9WS25MnLBz2ZmQT+vcRbpMabXFetOCacNhULOlv
2MuwzJhj217uiYzQd8YMYaQDYRN43X7fGa1qh0jsImZrFWp3JKbK7bsqm739uElI0DR9MIToiDSk
kJYQuj0vPz6DArZ84fHvmiYhjmq3B4/zyJFIYvnbP//nvJDQDiU+l8XMsH3qME8dt/PAXl7SUole
C/bL3iFYc2QLl74xUrg8wx16pdhHd/ZNO+0+lyT/1yfRJ1Z+Umn/ZdXiM7B7ChJYiDEcBNKHwlrL
iYa24cn3SW1FIG3EgINk+tt717DtJIceFBSsB+z0NEIsX5KnujXIBHBXkp4v7koBjBdSxwOzXwvh
Guij0TgDYdW265ILnTNSoKI3dW4i16HaSv6xoeNK+7RURFsxrtqsg0FPB6u0ipPDTDVoANxp5/Ns
j6/8MQdIgavMJylEpspHtRZQOghXur/OVqv1g+HL9ytQ3YpRFHJ1yls12mRqoQLk9v96wF09CdZp
Yb18RAROpaWHwGaURKSCkBMPjYomoUm4gEFrmNTIbKRA6ByT3cEJ5mE1v2InLAhCIXxGmkGVebyP
WaXsH47NUWD5v7xYvKkfVJsYNQHE2NqJJETHXUaJmGfLrTnbk6MSlwvBM0J4vV0WWBvNMHypgfIA
GT+0CSE6EBdLQNIN3RtYsg0cWBO6ID7MT98PtKO9V4P66tDeSMX1ELwRga23hoIJG5EBtHk+7Mhr
YtEqlKAyOoHxHRrVkAfKt7MyP0BshlATXA9KQk6EJU7t9KeHi8qdMnJMffca5aLcl65+J5hs2NTA
+hv8Udlw5yUoU5m/Zq1+/x4sCd81eU9RMNeuaSCCv6Uowr0VCaAN9fUobG/OcM60pFWXdFuHpY6c
igAWkNNCdNtTzGqQY7zZXlpmHgAXaNUPSPgNFsFdvTOdaCINvA3H3QivqY7rknk+PfT6DIe8y3Jx
2kj/R5JV1jFwRTlt1dyjQxB09/WP2puT2Voq108jMgs7keKUG+HYermbNu/h0nPgahuiCI9ymnne
fHG2n+Ar9fcC297qc7vZBCtIIntyhrMc/P+VxnP4dVTvfFkX+MCqt9S23l/Ti8TNV3/qEuwt/UXM
zrDXgusmX1xBYcWy+71ykfblEyzrzTm+xcp/8OUhGBP9jrj6eeXDAbBB6x1qHUxxGtaKojIU7Hix
OrbngtQTGr90Gq8wWkA39SB8E0TCSdMxebgtDI10A2Q0sISTqOSx3tCZR8/lvosKth4vZJRqpXEj
7iKLv0gkICyrbpT7V3UoL8R//y1btaqzf31c0C+VxgESLc4DAwihU+Nq9IG+gzeT6LN6ogznDLnI
uis4KxTqOLF17vYf/vQZ2ODJhD6lsRH7/5anjXWAk0w0C5cdBwlIDcgAXh7bcgd5OsH7OkUUnl/E
n0dK3gFDBnQ0KvIioWmwLkI3dfF9ddVrpY2pwvh3YocKvo8qDMa3a5/301YwxwojBO3TrTAHuzr3
QiiC+lQCDa6ykDfI4psrlyrGuvVe7T4+oN5SMZf8VK6CO1f1dMZQ0WiOZHBLk6E7yEaNwCD1RmFd
iGh3rnF2TdG6Xj0idC+P0sZM38PdfYAmFBdB94WfWYOmjbBZqt1migZjAB7kZxYdqCMrCG3BtbHu
C3H80LxPLrRkpP++Am0ikOeUNZXCW4TgXm40e3PgclaIIufY6vNYAWLCOO0VC5oV3+GuMZqdeAQk
rBjacgHOjtMLaiFKnnDvJPrN/TDSQnjv5UhuV4e+KZ3p/uLWyfyP4NuQD4rFA3imhRVyPT53I1za
BFsX+wkx8cMd4yl55gdnR0q1IrVVOpd3fm1oclqGy59yKG4+A+bs03ptnaNFucdPDy3ImfemNy57
IaGKzhHAM+HubNcG3PLKw/f5mkpLPyvo2NtOuGlZJ9W0uWqj6ULp3Zhlhm4yjtKpw8wgHA+LV/iu
0hROWNVSKZL0SAR80QCqit6mw4t/D+lZ/uwEqYzHcYRdalKXXikctNle5bF8Vp1qwgnaKFnx6gl2
8gRNyOpDtDDLaiqtEymyNyfygApKAWLx4KMuAubMoJbn+i4pNC6JkT+rZhr1DlPrP6YcH8tHjPsW
+X0OebDWMtrtg1t+3L4z/QrxYBX7G7hHd88VTfy1+z9srFoeFkJoPnRzmT3SwhGXqG0upkU6CwFb
VG1u4OXxACYQENbsRbr8eMnJXj5B2PSeCJSq5z0jGKZLBGxdFT/s0PpsV9Ik76WjNQm/KZWKryUK
NTTyUlOg1TNNt1+VPMqc0vWZlMXsbjteKGZLrs2e/2eb3WmzuOtKmSMkB1Q03vL1mZXWtMapj4wY
g+R8DnqtLdMRNt9dFlyjb36XvMrYELW0MFOxjGIPCDq9icxE9I++bgTyksHchMJ/S2iVfSbtb9ep
psmYJFR78AcNbc1UkvoUWnAU+F/a+FF/SHfnlV/nL3wnQ7OrcMiWi6vlMo5mCKi/SqjRMIMaxGtd
AKTiomcajPqlg3qmkp8BibbEal861i+LU843LeFSJGu2/+FDqTwh7pfoIBj3Wbud8po8XMT3k0Vv
TIdIKdkANhPSFNUpDyAdG/EJ0PjuACIbYAfzEOnM3XnyeXIT2X12lDuUrC3/wc/57/IO1FEaRz9m
472pnSJGxTLCvyDA9q1J4/9vjKQm+tbCnsZaGx6Tj09EfTSQhCnM5xKD8lJCRFX4SUU+OpgHr28R
pkI6xqNj+dqt8rxT2WNqISVbfpSeMzElhKLK0pl8cUECK85ayLKXGjuPsKF4x9wlxFn2OVeY5tyT
w6wjkOokeVytFDEw6JcyQpQaTUqkP4OVZnQ4/hB+EbitT9nS5UbEbTZ5gLoRzDwVMzGYOFjPdPRj
vQ4s+z/4fk3e4O3Kw9Ko2uxt+CLLkQfLser2aBvlFtQ8gtO4WCpYtwnrTMK6EaKf2UeYwHF7QFmM
YncTiyFUthqQNVAgmNqDdZtBD353z2PqOjjJU9iD71B5PfxCu5UBhSeGsmyjL3wtC1F/EAn9GY3S
C5blh/GFlTbyPn1NZo417KdF4uGYmcyk5D2TYSBEuaVFYziPdo3sO87cS/TAwHnzQI7GaXTdEGOm
NDIO9pKYe6VS7Iu+jTLzKygKn1dC3/DtUgI616mJPTpVE790zjZlEGCniqs/CDECwexHpDYIH9mK
64dNGQrBEh1CFKBJ9ZOPjbOagdL7dMtaoltjJR0nuxCbvq9QTKcEI/U1cbOMV7eG8RCQeZciQIx0
OpydI8IBX5HBDHWhSlbg6Ep8WwUHCQ85IyPNH1qhYTG+tTjoyp+CcIuXB/airtdZl1F4MjOeYcyR
tsD4MrJwIi/IWWSlWlZICIziIcNBNV+1wmkdwhKWJV6sTvFk3X4QgFgb3CmCxACyBBsf06JNpQHz
djJflJURywmvAQ06rfuF0DyMyTiic7c42JrR3fDaCR58+Slumk0v1G33hGPTTbYDWsP5LHF+jANw
5HW5NPQFLbfOTrQ2/7upxZGM69VGkOXlOBA/o0RtAlyXDDuPLrE4DjwMPTvPxgfFwX1KGBlSthrQ
kp3uVlUqGJxryrqABE7YMnTALp8lHxNxr3GHCxMNmqELAw325OEPs1f4WfUsKzT1uJzfPAXGIf6S
vQ4wB7SuKwqg3XuxiHs5CIDNoHaOTfMTFDP17UARkB9ClbMdDmd1iKYXnytiu/wjcKp90h8hEebt
n35RC0GKcFVeFqHfTqKXuLmEyxg7+vKBJX/iKkB79JdH8jQ1nvpMwD9cIKz36l6Zr0Vn2ZgS0v0H
dalY2UiWkpLz2RNz9l+OI2L7WSGi7Yvetdrs+h9CfzFwXlv8q9MGNEimSwmRFMzVa2BIMGDq6tpV
Y9vPgN4aImLWJHHkgVrInZ2VA/fjkuly4qbju/idi0Z+5nHKKBG9YfgNsegX10ukmWujjd1Uc5zl
l3YOp2csthlRBEj0o0C4wRFi/r5ogXwYK8q15VvFv48bzDDmPAslhMt8uKM5VyCcnimZI+1k1CNy
jKyJ81rLAWusMupPHWIHb3VXKDN3uP2W45c4AgBnpMBRXLOEeVmJChsbAwhcWWGYTe7qup8m6wt6
BDKqgtMlfRvHtdCBTvqMlzXt3kWQU8CRaVG/gWeUp55ZpAzQLG7BhOhkUN65UQcdaL2RoXpbPM5T
Yxwfm2mFUc5c7HsoL6xOxtrxyhnq6Kiw0mQwCbtryc0+r8cquVw1VJU7+7ozwmYsP23WV6+6zUwE
8SP1TXn64uxwJtidkleWiUj2suIUBIfdaLYJUxzTfxm4Ne+Zq5MFp0lAnLt4c5IzP+xSc7RnsVyG
SZSU2fjRAWhqpyCS0GH2wj59Ip4ddBRUOKbBt2myJjCzFs9RKcuT1xEVQE/AyCiAekWDV0VeX7Be
X2cUBx5HbfbD3YqasvX/eFlgPFrQbrX9UEcBzeHv3rpdoRLrCZMN/i2L1mHBVKDnxaDFU31C4oO5
5NT0mYjSjhz0G49qpSZJ7K22Bx4bMzQir6+EzUPgI2Lfcdt7E6KjwPyOAKpMQzUc8KOg9rUJjK3z
yt5SC/EryO+/qC+w8YMATZyw0QCku2X7kckZuoanuMWTVn+0DngAjxOhCzBn/qwfuqbvTDG8ekJm
kkfWeDPpNEDG2xV8zVqs0DjT4OPQmN6Mo8dum1R9mqzsLGu3DjsdBlRQnf2/UA+VXvmA4vvBhDrB
1DxJseg1bQZqQFjXnIEKbbi/1irr6atdLaaej9n01BJuAjBIqwnWQ921tO59GTrzNXKWU0GI96p0
iyE/YBqHnNLnAZwoE/9HnxMS9N94NkTMvg4EqUTQiS6z6LsA2ilTBpgU2JYy0ZNkRkdGJ2j5wUwT
UdShDrTtX0J0/mKjh3ZKYKDD8nS/dN+fC7u9AqDk1RtJ8oG14+/HARgyRLONGXXmkcsOvuTENJdw
FVlQIW6u85HOuvWKJFu9a2RG6ZPtArI0UhEQcISS7e7UIn6BdA5v49MWVb56K/zZmVkKREN3wxFJ
lx/lfFc1L6Ikp6lYOxaCdPBW3TL0Q0PGl83WchnotUAQUmtoqszquPkd5eOfrM6OB6BF4WUPFyFB
F9USP4BhWqaunq308qxcZ1kb0rs+wTdbrNMP7E4lVdimg3p5lDoBpyM0XNwjRPgZDjb9C76eRg7x
Mp0mvKPUW66FtvCWtQ1wEnHugyD3aJsN3sYAsZM2WPfeXd2NnWjKZAHsitq14UVtuM442n/QKC9s
IpKjMBAidnyXnl+pfMokY6fs/0p++VkO09t+/SzxdUNIaJ2D7bkg9mj5u/B5a/KFG+R4KAGnJyJP
xW8UDAXKOGsp8amMdBKOdaTE99BFsbAOvXiBgpkFaXy/vYXYa98jwGDUQVUlYcCwRrGBUenww8hy
I5CL5/kV5JvlpTtmjIc9kPW2muPfBt/h1ad5sd93dFkkcZX4oQB/dqmFswj0d317X3FT+SmVYU0n
j27LOwibEPr3vGhFW1WeoLVfzlfSMq/yu90i0WxMA1Fbt/pV3R3Xid/4F/eOWvpo7OXL/+whF/Cr
KTUjRbHctArpGpr3QstPfR9u26+/r8lJD7Dt+Gm/VCXcGZoCJXq/194QvcYHNCMb0KNjfMsmQ2LM
Vrh5jf7iFqxSW7bNqt5guUZW9aZ5d82psypBLjXhIZydjRz+UD40SAzrwGWjTX18nDu4LQtiujpc
ySwABA1LSTiX9q3NYJ82HilJa4DkuSuWym8csKHq3R7N5x3+yMKbTQfpbP7mpZzOhebqLVrbQiNu
6RgIz11up2wd1v4nLYfg8kwEMotG6iyF1rkpmQUUPZy6Ct1GcogD/20VsZ+Ak/K9AlCDLnCRq46t
B8kXXzYP0V0SM15nLVuivjH08rkDgTx/s35WxnxoqKEMxj2SgBF6ZYcpzR0MdtAU+6QXE5xaDgwu
qEPyZGKPqlg7dBCa0Lb9fICRjjswkTj/YjCYl5/PI5tLRtqrXDMhb+Ztw9URRIGnCZppFinCpfwl
Kdn0y6iqI4LVx51hJAN61B4mSlu+DeeNBbz3YORtBZP2MNqsurM4eSmXVbVMC9ChLibgbFctIiD8
6du+sq/dG7H27AbVwNLeKXsHb+YGUR59fFDZPOO8blp2mZQ/XGNIusPeqcEb8Eu5vzBmH7Zi1s8t
rUd7x064bO8BjrbkClUEVo9EfTv7J5ABLMSUf78ieE2woWIMnNGQnteWJEBG32Dk4snnimzk6fPh
mPZ/ST9bkTUNh+CzA14QQGbIbuFVyEnOOFe+0j7rJTT8QDAvV/9vwIkhhbgF53OsVzPDH+KdDUb3
OzDDAsyH4L8HGP9WKUFcygzwTGZXJ7LIftS+LOQx0Qo74lGnU8Pdb9pFFiZe4tMPoOrIWmusCbD3
H2B4ve3VWs+PiUSgDHEHbRQ8t3/wfKc4x5MSJ0SUaSapbV3JR86dJjcWU2C1DXWtu62pwWeGFlJu
lfJwgl6gKfNV/EbafhPEw2Byodf7WVFOPFpGsBlm2JE1o09gUxv/cOvlTwvIJ8FNDgoYXRKOChYJ
jdyYmiuTmzB1qKeYavGjc++n0ryB4FrrcMYuhAXbw2ck8/+bMAbDpmobqV6CPb4hNIOi6liSLFmK
eiT8bI1HTCGJZkBi7rZLdVFNF/IBlkrpEqAlgbsH2X6jqIWJX9y3eIOGZsrRZ9fgnmpAIWmLmV6G
ixYhLnxeiPy67u4b6wcaXZhEnLIPpQPIsfV+KwFcd/IcoumtztChUaC7OjzcdYw8LvRpNetFdJTh
R0Vkz4NeNib7AS8LLwjD5w1IAb8jWG6X4USXE6cOOOI9bzFm5DiN80k8Buj4zo/nJ01xqi+AwKaC
ZSPp+b08Y+vMq37c1pgUzJIoFenTFlmDJ2I90r2cFLDbAjLQ1Xqc1hBmcsYoxlsVbE+pQtNvMaRj
xB9xUyVEmKMqceJsMfiKT0yAzRl8Hs37k+AggjTWJBoRi4wwpdTfaL1RNo34ORgWMBjL86fJNFO5
vh3As+JCjuMqgNcnHhVeDyzUQJmzzY94B4jT7EckdHYaVK1RQo9kt8atHYbpUuPwpZEIif6u/ez9
9Iw6xQxVDkkr0gs9RoTGzrT1n7OfEDJt7OPtkNoM1EZuwFjJ25UN5g/xazfSRmrTiLV4S1yyf/f+
J+6P1Wh5VL1Yg0TVBTynqlvx0iwY5gnwvwrf36tLZg1KTcGj8Od128L2nOv5UrhsBW+x37KwhgDi
cQ1HLXu5yn7nHDMSa41NTqPJc60nANagx6Aoi9gs2J8Twn53KCpflGK1AMCMBiAkykRVdHnbhQjt
agpAi4kwUOluJQqiFqmHrEAsaj2u5EbhAFUqc+5JBkLoUUMpikZcegj38RNMY+mqvz47TbZiqW93
ZVr/QiRBvs/cre4rnsR1XNZEnSrApGpKyjM/eyiCtNAvqmL89Qln/tnsO+itQBLge5bO05VlEPuy
R7GGHkI2JJZHsE7FaHxvaTF0v3u9MDCuzWv39BZx4tTlMVwnOdMoB0cjAelu6IpnvS7/805a25Kc
VIFe+qya4NtGPFfOb0cCHmOTGQnz/5V8znfdSLILiopm7iDtbbzMh4ZP8NJ3fecV6Ez5gIlpBYwv
Nw3ruP6rB0+oSLaAj6dd2Q5DJmp7l2wn9d2HzF22SP9gKXihYASTTEzfCQtIDrrkRHjYxZlHTl1U
yISaTeuKmIhe+6IZ2HxfDcz1EVTmBIuNmqQVMPoqdzk54MXd/AGU4Q0WA+lhgXfx/+KOxM040jhn
b0HywZf3s2dfG6AYLmcZp6Fsi32tuiX/q7a8CeUxF7jAl9jUgYUcxuBWbUOMmS0qfBiorXek7CVy
A1SCuDQ/M/jmfzRiM8R43JHJ/MA7ujVTKTEnPnAVMUKD9t8DUKpYt4riOBPmqcptYSaFwFzG9H3v
8aXZ5OpO+kKBGKTH5U7IlOSJmw5ZzKfucX6U/zPCyrf/3DQgcUps5yij8lA3poxSRTjOUlALbVp8
kWu/iO81TF8TDEYQgIU4itGXdNVtx29YjZnOyuPFk6znQ1GyxOzersBKgH76Y7Yr88Qn4GJN2p3B
W9/QziaN8PqYnIGTwevZ00mInGFbjur1VqPncpVC4aAT92FoK7ILax2XxqBd3ezPeZWWvUtsiQGZ
K8yErKnKAQQcCYzBqJ3wrM4Y0jYODnQcLA6zVSv2389zGKIAVzMN5Ka4F1FM/t1BI9VKzK0tsAI8
lCl8JloXK+O5RQlrk/zHj3cPHAK2eak0UAOyu9hjvq47ksQjJTEj9U/hc7e+Pz/RSRwUoQ/T+1r+
inspOvPAwHzqhQSen8qO7AAPAoJJspPw1fN1NvAuSs0UFU8ltPOnCgbkJCyI5Nl1RS1RADEKSabD
rU7g1UmL0Ge1N6aWdKDvAoUhmjI17Yqu7nZ30gScJ8DHJUiaDKlmDll35s7JvH8SLmHySXLI8HUQ
hYqM+9q/0LcojaHk+xd+N1xMqcWYijPkB5If45mVsux2udX6QhkIpR03sM++vE4evul+T0TGxb6a
1T3efNmi16g5KIdaQAU3mzIz2C5MJdjD0m2p93T0cfNdM0JSV4UB5GgesHI+bV2qx9slUoUyo8RO
afOortE6FjXZmYcR4RI/1Wr/X6CH0Z9vHV7GvEZIsZ474GLa/wmBmvmWUFwPzj6GdEU27zUn1oUt
MeOx/L3WKJvDdtHJ3awRCGrRXL9HT8Tfv7DyryW96HgXltITcnu5sVgs3UQMbSNjNI1n7PdFEXw4
SjYaUldHMDIAYqmIC/lqxcUuCiGWaQTwMPV6vTlm/b0LspNeg8W/neeYZXjNwDT+wcE6iuhalz0d
lXlgaariNZkKvFCx+qDl/dYo26ABvfpuHCiDOhKbqw9qgaB1qYup5NFgqHFfrAjON7ObltPENYVt
ckl5k0j9EuDx0On+ar9rRAaBEOh1uHrgxwy5wJqDnDiMQ97DQODbwjOBieaPIlBvUKxEOQ9/dyIU
RBFLPK/rPvFcznkTugUXqx5hjjxJrh44G5VyfusVX5WzNyL/2HBKdX3GRpgTmv9aagp8hM957oc1
yd5BtNYZZTik7SAmr33cZJTAq8P+GS/hIQZTPaz+mtJDbsXDpZxOZcZef2f9hEPuWnRn3YQVUyQO
IWydMiOB1GdOkz9eysgODCRPBGorR8hxMQPuxOicuVO878EGAcANaA0S+JuHmKBCpqDji7+OtBxs
Nvmgyt1FySg+zOsBVJuuIje/OqjR+EzWjOZQVDF+ZBk5PFriE+/mDXX8pFTRT5rgx0XyvJe/rS8i
lGOqTZnLUbLurPkwIu7f+a70joyAyR9XqDRi/vAunz9im/Gu69cQ0bZ/UD4F9+e95ACNOlDHaVMP
zkNLAujKkZnQXLZV63TggnV3/iKE7wfnfq+El09GfiKW0UIu/xPOdr+YFYE6ViNkuJYJxXOWvknI
c7sPpo3afOLgns7++5/ysH6Naiir+ij5QfqpF1aqAjWUpUhEQcuL4tofe52mwygfMAksMoVc+jS0
A4eroVstqCKlgUOBBqUiQm9DZ/2w524SbGXAaB8sgPJd15YwocUjP6Fx7zG8Scc8OmIAbWuYkM49
oq1JrJLv80GdY7YVlWQSpk2Cnw4cuyZ/elJMEL4RbHIaE5S0F1fOBfSyM9mUT4Rq/IF0pNDHJkcz
zA2W27AN1IUGlFuluTkDFuCTjt8NphsYe+d1Wz2xTcxlAUzQGGUUejMUSmQw4WqDmwRcZ5ezYpaT
adsyTyOb51aYI77M7ChR1sj8tU2RZMtsMz9CoPhAbhV1u3wglGxUOXk9NmLzqckcTxhVpMYc5PSH
7neB17Y5RB84UB7pxyOghDVa0/GomjXrR3Raw7NEqR+gKZ77pcjkX0ecgyvzmO1CS0Glz9uKmyo3
sYC5qR8g5J+YmfABWAHPn/ZEl0t8eECTZQYm+UoT4OAeYmDS3Z0VhqIQHdt9zJSFmIAj00gEaCx2
6JSFsOM/B18+DQABY2fAIFEhwrkhykoCCI74G0yKbSlnwrd97lfSiaqOxB8Mr36xcKF1gVzLmywd
gbuXbFvOKE76MFerX4sWvbhAlM6Sz/eFW37qjazJX6U67koop2r7Y3+twNtY4tvc4murptHrFz/G
mZcqG8jHGeRtt2lZMrL+Ou7WGadd5r2pT50ELtGoz1WChD3EBmwB9AGyJeV2lBtwPTq9oLt3CYEp
nnTME8c2W+tiGCWkLIr9Kl+SqilRTyIpPO/xvVrrgdgZqzUW2eEGy/XpaIq6kvLQUYGmlvN4fVHD
71M5nlH/C59ZrVtJS6nUo613wOc1VqZJF0r0J4VzsxYFrRzQ/o3j5J1Ft5CZaLJvjFj7qiQZwH4W
TAbhcHnDZeUXqevM9pBGyPL0sMgj+fcTbkgHlKvNLoUxP/7sGGWSdBE96cp4MvukXeoXw3NWU9rI
ZVNdeCEAqFvNH43UQe5cl4lox51IrXGEfryn38RbEpE1zMHs+GxPEhteyIlxa8QIPmtd/5oEOpEW
bGDTeJwQw4Nst/OybNnC/nPQRf9OF8odJsPnBdMFt7Hbny1vsCTiIwZ0jv3VGJjT4+tj9xCy8dLz
3mEwJC75W8+1NkqFkuz5wa+Pgs0PCWEt3SvcTHUH6b/s2L6xBz5TLQcFEfGdUdwa2G1umfMLh7NY
3UnbMymS3iddvXZhZ2pD3hTawa0gdGLX/rcfx2X6+vfGghpzf4/2SQzPOCa3VAZwRdKF9IUWeIKW
iZkLdprRSQO5eTnZfawe0406qH30cBmqYFD1Q/NBGQjwr8yVXGwZ4AEa7DznQFOcuoBtRYMcWTp/
0bKsWV9zXE41vQZGdUkF2Q5LoIomyHPh0F6l/AlLqCfCeXzOgmJUFi8/pK91/b1J03uXi+R4l4JZ
gUj3E5Fm1mRA06Tznyx4RYPVCeB5PNqvpMaCJjU0vFAd9ME9T5dG9RYgXFqvhalGZlso2AiNs5dW
wVYTWlTDM9FKm1/52yhkRdpDHmFPUWOYSGIF6Ovt5vZTm2hMU5BY/GITdOr55K6P8it8z60e3XCC
UhSm32a5YsDo7GOcuctFiX0wyWt1W7+3g99pBvxX6ajE+IRZRLzsxah4/r7y0iVo0Xly4JnaVgMf
rahpl0BDRkyWcEoMSLSrFgCFtVBnhnp86lCKKQiL+wRaov1eWNbt3kV6KogSX+97XPLmB49heEVh
ZcltWZM5cM9nfrbKPFCyVIz0Fb+9kNBNSTaYeBT0KEIKsgKXV7TF4FEkBvk/j2ZqGaxTvwefUf/g
7YHkusKZzqAxByNem3ktanEm9jA1MVO/7vUiXpyR3LMPjkzGnEcZuduMRnV7BGWeISCB/iRLSYHt
9WfEHB33diiObCXxmGF8urm36tlGsBCDEv1qmwrPOJagidr1HzmuGfp9draTKRgkLHF3EH+GVnK/
gB9jLmPA9RUceU1TOfhV3gdFdHEUHCSjesbjMpNIsFHCoYiLI1PsoIPYW5IJIiH48rYA7+H6SPAi
ZQ4NMam3LY/XKOoAmIM/X5UlSCcN7PVJbImnoAESNIDFw91G8vgiy9Y0DG0y6BupxCOh53+GRJWm
wgFrkHoXDdqbLR7NWNMUpEX5P/MRfcMEQCp3no4qKMD2VCBpuijnihkQ043N99PL7pR8zDCosKTz
vIRqzkUmOqTwCBQIxjt3qFpKqsNUPp9RFpIiUS7TwayE42UBZBoz+tOr3C0CoLpgLcpo/0+Lswk3
h9aAP3qD/RoD/KIydk8K52vi6o1PXzsznGzocrcLbLBb009L1aXvBqAtoaiHB/0aqbA0d0m086Rp
lVZsSj8cKqTkV6za1SoyEdqaGy7ePyqXmReyb0OajtmMXYZk0haL9rvI2Amt8ZUbWRSCJcv+wEzb
IVBERsZ8XP/Oy9A9h5BAOTSgsv/9Y7GqnLjIMHe7aObK1ix7a2H8WsyXNp5Pb4PqYsbBP6wAhTE+
OdawORZvTJwj4Xn/QNlFxob5vGNzy+lRpoK2drMDJJ/CPZQrjbxEuse7S3IBnqgfz3kc+ijKDErn
9i0lfxthczEb8OPpYRWQnsH8AwsFFOB3mg+r6BC+2gF3I9xxp1nnhWer3btcAPldobgRi1oyg8pW
CogzKb/taCGvNQb8Ddw6RlUKXHobPACltpmCUyz1vokoTRuWM4yz3y/+Kvcv0pKbBWyqG4RO7Kcs
NIebW2OL49+zssVD7Jd2FGUfcQ51y1GU8M/lWTUISG1WXck5jk61MlAqCZ68iYhGJQ/OnoInZNt+
jpwbFNz5GJjsj/xCUi/4tQz+HxGrh4CXVHzY9PIwz5XQwioWJpUAA3/x288NU2zn8OGB+OqFeht3
NRKs8zg2mRduYKc4BW2ZRUyqdxbC6BReQx9ny1UbRp7vqV4oo1mnUwHs9+6hDY24jo7Mfk3bDZ2n
duUAPm4wVHIW/O7DKrBCfzk4/cISqfSf+glaNU92kUfy7u7fvIXQ1U4S4p2KRxTchnnQyyE2Y3Mg
h5gQ3WGpJHgIJxKFZQNgsbv70ZIzp+HNIAWkgRVrDSUazoX1S71JesAV5CZhU0sZEXQMP/awceqO
5VPyavGcG40xKPch8HRLw0agVB5Q0LktT183+2Mtn28O//4MuVc24m4m/w0RnpxIT0Fz1mdgxrBi
1QSEyD4djhfIoEy/aRaVCankFx2nEwV4AWEECPxo0enYvQea3PRNDhJ6rGh/QYizpLQR2tYhZqdW
fN7zczHIAPuZarYpb/qt5fwLSw6cLpqtVUP/lJ49XOUFVFn2UJ4uuDexGJZJmRQYeSvbBf2Et7tI
IuzCKSXSOFwnnwfDagEzQVqmRRg0ZitBW2rx//XrJjYAFS2I/2Pl57xsL03sSlQw/Udjy552bVDy
cn41JaVyEv1AtGquu2nL5C2n9WY2u5CVzhzI/q095ioBROs9qIj/OPs4iwjA+HH9MzAKgdpGA4pB
VxaBk8WUefKX+IhbnNZdkAoruZ/FJSMt3Of93cDpBCIImv5/nQ4zOXf+RQK5q+/0+Uk6MzHyeRjE
lSQBnThs+b8oJe223i93+yyZiGXlvdil5g0GJe36Obo2209RywQWKXlWeu+lzqntPoQ9nnS0yExP
InwzwzvIs08iZKtQ/dmW15q8inaoPxAkW6+mfDFlfZyXyZdnjpQ6YeUctjR1wRBI/UAvNRSs90my
yzsByl+gxNn/Lu5Aln5DdqDyROUoRSEbCtBmC05vafnxMPYhOqyj6RrXF2Rwbmx+sHMQkDW6nPBJ
fO4vNL+puVm2c4PHitpDHiDDrTX31j+Xl0/xcCykIMYIAZly2fjyXOblyN/WREU2t3xxl7HA8EWt
Ud6UNOU0FAXn+8Hk1AfBAWweIF30aApAS0PpuIMKvpkBvFWmplipnvpkiWqePRmZbXxo+CNAI3zb
DuD2xBgBkQjMkVXh6q5lUJC7H6fIwiwR++1AlmPWc7jo9nMRx3zMPoyVRSDD2IIzkBqJe5yWIfmt
z6EhqAOPGDxeqkeZlJBdd9shepdeohwx4ihgXJKGpKpKWExQ4JFKulvIV1bD5ww8cLELJg+190ZW
powazCjUGU6RbTH7mgHk6pve7zwKKgI19KRzj5Cxkuv+6fSBebcyg+LHCCyZuEnKTi9w4DIeIqxz
v6l5+9ThzZP7FmAPYYgfOko0eViqkxN3UUVfzb76Xbr2llhyxhrpikzoXVc+Yk3stE4aXMaCvnsn
NvIyDOdyE5NHC8+qeV82bI3e/psbqG0xmyelpBWxKcwtJWupnCrD6DHFmEDeBVXJe/NjDQ0hLqHs
hWVaN+uy6ZbPyS8bT74fz4gKi1geB4NLKmUyQduuNbVMTzGBwu6jxXInZpSIeQEiz7nWbIJicnw9
/HjEKiq1sQnMcoiRi/1eg/GnoggvkGpedCS3HWQyxT9QACr/AJzGk2/3pIFbq7TmPEQoEsbp8phB
EGeaAW7nggks4F9XUjBob2bqCLGjtER7evZr2QNm+OwOX/W7I3vFe5qRUlwNRdPBb2WtuEOdlMNO
e3PxLwHHVGmXSAeTON4J/q37PdmKIoIy8xKLW1/1i84klDcZPQT+7gupIPvYYmsi2g+BqjysEb8Z
NZQaEVg4k/wx1RlfIvCr29H4TUoZRvo3aYGjhNjSdAElE1plBh8KJmU9ZHc9TerYaM+ce8yvij9Z
HeHakMFoHAPoAnF8o7GEKcBh/Ak1+2zPyjypK6vjikQX6gQim+VSc0S8oQi4sox2hJkhk9lTNNAz
vVpPH6jqGLuCd6A639FoEnXbf17tbyqUuzlzrHpySJggwdQBw+h4tzxgwXOvAkr1jcRPQKl1XmoU
4MhvwT9K36p5Tlvm6RmGp8TvZFJWRS0Su/nJ7Ddqqj1THtEfPPK/J1A60GMEvY6IGGoGMK8uY8Ri
9ReSwD1WpIZRi/i329nJN8JPsLUu7hBaADwnFlCRI4VjHAdUzqqg3sMwAZU0gZp5wZJNVJagkYE+
A2nnFLC0L5hrD2KCOYu1BffI4v9PlWCNhB64nD8z4gX9fgZdQd2nDjBL60n0I10cHR0A4+QdEZBd
syior2To5BU+mCzTw5/PALHwIL5wNnETxXf6kw6hnrASkfjBdQcnc39e2VquP//eYyWxzA6eOBpj
MHPsvYqsYrTpLPFqa5BsXcB2Z7FpFEasdxo7Ziz2QpllnyrlnQZgvIyfdwZIJ5fO4bnz6zTkSPDU
+FOiWdGVfHN5leixW/D4lEoL3K3vt6K8xZ7VY8KYDtEyP8ZZDmtXvWllBCfXqLfhntR2ZukXkkKO
la1U2xSWGvChblQvufFAfCdMOKHnxqaQxG8btagdopkyKW4LKzEB6rNy666SwQcfl6ecyF/J/G+V
Nx0+6jMBpgoikqTqECFdzfKrg0+V4x3qpd77VAtl6LIwe7JVy3RYNp6e3iNWsI2Bo4pbNvahJkB6
/FVjInNn4zgTp9jvjKMBeE/SudWQl7iEYaMi0QuPt1ge5wy+Nz1xHEQGbwi82KxqpwM7RZffu7Q+
TM1ZWs22byG1bGNVHn1eQR4VxFvXveIveoDJiCJQJVy1HUUBOI0FmIzfHsqMw4afVfZrG51+PND0
y50KFyxe6jZQTa6/S9t/95/5OSq1BVW7uSs2bfnyfkKO5E/X4puHYqpfk3sonwNPoH2hAiauWHFF
mkObUDnAhAqlxqdkcnkVni9Tc53WmSaIKCYWBqjmJqs6jPJVc6TpaIaaNGt/lfX+NKHptW41qjRJ
UmL4cB2O0E+pKVWZPoL6nFx7nMBLHocYVvCtNxsRnt4ClxkwCXWSz9soalUpL1/MJ0srpcnYKdvN
53SL12r9xbo1+dqGOZySwMBIgWbCLPyDEpucI8FFdoq7R4+5YwQWhJf3OKXvmgzQva+R+QMw0Bcn
WtUB3NIQkJnki4sHD1JN5Igrch3zhCKRi66V/VOpgoz7XJ3hlCsxclJZTmMhz5By4dvKMsG7NgOH
QI8plCv8oL2L9tjHzG1sT1Kf0xFTUjy8zX4XeSrzDMwNmtCbyrrs5z0eNwgdBl+q+GyjdZcQz7Vp
2pQ8fWIHTRbH5T+A6nFIbPMS0LHoXV7SW3WNRGPF08k7dL1V60j9fpnz5lxKqUfHwv2aGp1crbSE
gSGWkkm+iZotOwzb1lNvJO0PLFp50TZBt9pXB0wZkcNVPnZLXluzLgUUDWFeHiWvvUFxgPbL/6w2
aJ3oFKMX+s0nLZqHeRKYJVcEvp1sVHp9ByrVgtpDl3BtC1wMnT07xuNmhxfj7h7cX313kuCEx1EM
Nus7vj1g20R+3n9RnqQ/AZ6a+YsKsH9ooqmxtdl4iO63wx5C1tKGYtaudeYTiZlSo3hC1//r6vgt
K0WJYmUyWMYi/v+e4OEhGiJOMy+6XPDqndseHkajiLuaLvmAoLJ+CXNHh07gNq9h5qlHotBqtDtm
ry1eK58zG42PPPs9HSZuVVk7enI273Ee4eBxtfq5iEBZau9cbrFNmVumTOef/af8JuQqPZYR/aO7
GUzqek7JXgeqGBaiezu50CqTPb74DoHrk4PZRFyGPNfUWaM+nR+eiHqicc+KUnkbft93qazRzXAM
d9HOkgCAvU/vVAlWnbx8AqEp62Cl87DRb8YyqZ3NdFpRY061eAW321TFS56Ze7D1/JCT59Ombj21
KKSCSJwPjo2tlujKU73sc6MhQY7z4EeQevfFbRtXuZLqFbGOwKzrn+9iKg73yqPz5gvffd2LduKg
AlxKh2KnE+nY/d1vonknFc7yQRTo7m6DTHR4xwOM3xwmB9ZgR5NAikkSz2oGXd1d2v3An7TpjvJ3
dY48RKfnFe32VU0SvSpniisvjIuSafdXwj6SmY/4/f0PRVJ+MsCMPP5QPOiNBAbn6PSweB0dRiEg
z4GCUWLVcydFtvZ639WI5/+VqRRrGNkk4TRGigeyVQ3IoYSxS2txM1cVlm36Kmxd0RfQZSU7V3kT
eErPTWnloWbBBRTbcEkFkY6F09sSGSwby3LjJmJncErVlaXsUy9ztUE1bLIbehIr5mGjiTaI8LII
zlDV2EY/fAPAoDdoqn1Sl5+9QDro3htF0bmFf02BA6aIAbO0qoYxjKxvRIagFMyB9xDABRLscoKM
rjBH42Pb3xj0RI2G27ME1tRf753F6RN5oE1RihMP6c1lcJYvMpi308ElYLz0ztxa/72cFgammSym
aD2HpQyqitkOkQY1slYiwIh2SGslDE+W2+ZVosAkQQlwvDItXpNjd5zLUnDSSFFPYvMMoiQ0gmXk
tn7ICBovq5wTll/xTx8DshCU//L2PuEVfJ9/SBDfMIOn9sXTLsIcilESyspWKjshu4j7sy90zDIF
Z0FS8WImTILF8YLmCb4FTqG8jKuHGylCjdXHCSHo1bIJhHwOMwxSnbzipqwNVQfevj5d1AlqAWlS
MTC++2oI9YogqflwJs+QMyolYrDzv+Gc0Qpt47MQqsyWWzfNhxz2SZJILVzbcQKKBjshHGLY4sMm
ydllQIQCltFtXDfNCwJinurixZE6Q/3xm/74evZfJLXYSReJ60MTDCVTVUBEnJUdiTFwWO4n7MxJ
wumha8iGTntPr+wf5iy1n3P2+GL6jzAdluHSAnP+Znh+Xjv/R1w3h3PjbWDtzUwmxaS27vlFe2Mq
B+jDhrtsHe9sMFj4vjoLEbTwm1/KW2wrA0C/bTDgSsOfBF4JhuGpiTVP4yFH7fVY0z8IY6ny3v2w
8/1x9awEszsCZEYjAOm1oQrnqHXRXGBTCqkPA7G697+fVELzjigoy1C+YvNzno2ofiF9pZar0Eer
CBpreklgZJKKOEG0Vs45n2Z6+nYdADNimjPS4LRXwC7Qj/ZO8R/Wi4blTyM0IkRtZW5RqucswFAn
6+dqkuvoWLJgUXzcX+juVH+0pH/Xv6llphQTeyE0DaeDY7PkAgK9yBxSuQuUuXOsFxATDqaKJf0j
Nhi6yt/zXVI8FYLc+BXRN2TBREv/v74E8oWOtKEdIuFnSfoUir8zhpQ4AeC0wUeSQKcGnk+xUJY/
/zFxQVhePAiiOgy2cv1vM20BEjLCQzxR1NGrZnlhPzlPMUTFFZxaatKQSCVfRrRJtq7avlPP4v6W
inQ7hkJMsfiOsAIXOMn7/rGiwJu7iMxm2utWhSKuoekpLHDqs8fvRvSWFEYRgOUdwRBNGnH4dU6t
ExgvXzogYmiLVLouFqKS8E5CDoKLvdBHm758hfBSIv9nlz4MlQNlJmbP9dXNtjdWr7XWNkUT+Bru
c3xIfzeHdnPDOsNBTldK592BXskIbkc15VyIDizfEX/lcngRiOOgQ4kmfDaNAQHBDHTuXFJV4bQW
bSrXOpHFXdV8aVdTaXA/btlhtNuZy4MinAqOmmcwwhsSnwhE/c/XPmKCEuBNC4M+ueQi35PFE1wj
8zLNfdpuY5XPgr7WRwuUMeLxRljPAGXqWMtsdAeKK4bBxU8sp/KQ2PUxadmrI/rHnS08WSXe0L5d
nQxNUFowQdTF/InMOVkgHwzXVaJo0oHcgAVFbbtWHykkL0Ox3LMLgxh4uaY9yH7IYxM3noffgelO
HUCfH3e59i05Pg5tqJAsIi9X4AExDTM4fmpLcYhwcQjkEXMLFPiH3M6Wrbe2eqzfNUZjA8XhGvKm
p0DcLFSM/sal7AZppxr4OsgN8955J7m6GHbaXBzWEVqIeJlha3v6TMDDz2UwdjTRjmWke1xmbZNg
joggAh8e3fMVwR+Xc+H2rWVk4EGhcUGWBBNM0RqEDhhogT+OgWLjIILZtdrWYgh/KCrD36J652FL
Up24dPPC4bI6r2gcsbQ480W5h7DgNk8fmWy1L+QenwY0MVy+yL2lhuNLmHQAgIxi14P6b4AZCVh0
vtqbRXiVsQq6RLEFb3dCR8XEotHm+6IvF2KvOuCpHe3icatdKhvFcpM7tZHVaD76CN5yFrpWidlV
g2K4Xa8ZUQrkhWWtKNORO88qTJXfQ7XkJeKpzScznpIvquvH2M+CjCgB0USnQ1//tIjmXHbzO20p
ukv4F2ngWqFb7lOGC2VE0Y5c0dlYSxtiQk4/e8MmbYOVllt5uAgZhvGSWxLEmsZG/a2dpr2hdAtM
i1jqV0CXnPJ82+nEynCCZxi8r48h6KjqTUQ3Gu9PSK00nk0IHnhxJmG7ONKCGT5DiJh0kSadeCWs
pmo+vfrkAwv0z8daiSA0LIBEIYwebxY2NpOkyzxigRsJzh/j5tTMjcDymJujH1BKCl0/0NIL9ONk
TWl7ujKrDdLvXSrjoyEuWQGLX4ECeRGw0081Pj9rXzGmij2Dr1zsKTa1lQBt72l67pA4XchB7EcX
YkmpT/HE0gSbF3mTqRv0QSg6Mv7gypOZkpSY74FPhlvkIL0RT4k9REFuhrMcCPyu2gG5/aZjj/hy
OToNuzpF1oDTfxz0/xauj6ekncf8Uh01UXKp4+26QqIqYspj1gNICeu5RZ9VzcuPMGu+JySOSnee
48zfqUQ5gRJHvLmL7qAmgl0UoCCezugy1AWOmW4DdXM6yG6FHr86wUQZbhP5GvDX2LHetMuOG7NP
IoQYXK5VFNZP4vQQO9O8spslnYMf7WofEwR/sQ6QBPh1t4ATQjXr8sFYlSF4Gm92Q2V+aj5nuOoV
1cSoawPqp3F9s8vkFe5Wwfk5F+YcK91AQrFBSCi3R3oZ/OYBMw0Tq3VhAMoxRLWv/NM3ZAslCc4d
WAs85qZEZhIhEoTQh7DDk/sLfAYmEYQ9Bg5laoIa7+NRU62qr0P3MbSqWVTZm6NfsrLc8t7SLtuX
Y4pthFhvHjZ1tD8vH53SdXezOhQTPlHbM0dX0YQmdkskyjngz4CviDKqnmQuTy8ZRoxs+OKIcZ8I
hObAcEh0aeQJTLODnT3LFjkNPKOP9k1W+56lFbxEAbXNBI8AOTfeHL8FHcLEqRJskZ97+pomEUBW
OaHvjDO/pvwM0JCxMFD6Ya0lM+AsU6XjeC6QP3s7bv3gIKKVHDuslGFqCCOsXNtwccpf9oL4AyoM
JGa0Z4anK+MFr03HIoBULJKbaHW3AQ/t49KrsEqcm/CyIrhMXProWUKjQllYiHrdd7LpCzXeVKX4
rT/LcgIQFhCCU6tJ1W2yfqtuSFb9rvuwnrBz3B0vVkxSU2IfW2Uo7Jbo2yOPDt13C71d6/e4DvZH
9JkXjZN3ayn8zbJWWvglIGuI53VKaFAhWN9xTNixOTgb33mOZiZJIH37vsCKfsTpq3xVlEQeEFDi
EpG6htzkg78HhZJQcNnKWHGN2DVOQcbyqAa0QmO3hI8718Q8k0NsOuA0oOPgmbH/O0DM4cPa6hQh
IT2TgNRX6KVS9wOxqK1/Z4F3SNphONDWdICnE9MHUO/zahrq181WNG9l6mdgv9UCVnnJtHp6yJyB
engHcVh4T6FrPdlkM8QJUYhpsr+dC2CP38QcC6EOccMj481Vl26ZuuvqsBcJUOgg8XA3aeRryt1h
afAXtBVGAzJqmcCdksuSF0VLUcSh6M8CwES5XNePGh+Swr6LpEY1kbK/oBu25Cj/KrDAmlNPtnFk
kgSXYotl2tQldGY8ntqBXqeIG221YuG5o3sOgZepHVwW8pruqKUu0isZXiGbXX5njCl03RV3WRXG
VlkopBUTH3TjIa3M4SQnNX+sIqguLNpBwXeYrrwhlqaGAnxLL0zckQD51A49nPMIMYsEzH6TQn7P
E18LOeyrxmtBR3/yyKAG+4o1Nm3lVFoKGoAfD+XmWQAI8PNsLxNQrKA3Na/hXRDsN2V4rNP/jxdX
WU8OD3euq9tJGwHPjNODAxRUDG0yGFTUaQRYIY28+6FMZNZTpbKOY3W8g5ffNu8XjtypuUd0D3t2
QC1KmQBMTFWTsgbXJ4tqYyaZ9nh79gvqUa7wsc2FdWsViRydLEelTQ/OFpQPmNrXnsIWQENrLz0w
Qqa6wRw61TuKNFHtgf8oahRjXl0QayY1sG8D2zRmhg0Iq/9NHiabPWL5Sqby4e6nT76HmYILaz1v
tYEAU6Z0oiQ4o21dX8YITUr6mmIPexK3myTi+H3/IG0BdVpWJXlIlGANzp/G/pug+bwyaHK2GXGg
7+bHM9IMmDhz+Ko991/0oXnWcmDGEGVG3tBjLUs8rIFuweikIOqRyRvg7ipVYcSeB67s1GKG786G
O2wmiUbH0TsDFS/YB+erJKAK/b9arp1qEZL2ztc6u7rlxsDWhjwV+FByP9w8Xzhba6HHtIUdMPRK
a3sP7UMHkkFUbEzOQmDxZQD0Rcb39EyYYBQFyMwG4kaSsuH+ICc6XAfx5xvThHaWrzUoz/PluUZM
R7dQAIXrFqWxPNSteLBh1AHnWGVSOl/KBdL1dxTT735TmAgOD80onQQPluiv254TmYneCM84MUq2
8iq7J43UTpqz7W7YTZtAfGo3PZMcooqfc9NnPjr6+Egrap70u/SnbpOySM3TcscT6yWS2gRXyIGz
VRZWDRe1xoG6V/7uSfFvH/RU3iX88oHK0yXCgKSGyLbCQZgmU1eeIG2rN6BRFwAnKDxe1YJ9mgm4
XyNu6sYzoEzDvHG4LrN5D2noZJd6iFD3fUijuFuiUFA6srsXL5reBGSBfYqz0fKAk6MMGAULIkZ6
UYyGiJMveTEfTqvSXhHEHEFjEoPXYPc+Nj2u1cPaUTpUQ8FWeH/MTJe0y0kPwpZeudTXd0cbcasS
fO9+rDwJ6UTRAK8TUbcJxSrQnSZYgGg4ls2GZRYBBWcN1HrVDzMOAKZo8DjjKw6+AaKVyZU2vA8q
7Q5cemBrR9t6S4iWGDMupZ/gJfcn2UYUY4d5ZLarzkgSk6T97nISqiA3naJbWskhgPYu7HeWDO+z
DLe8Oc5b/17w9K+iERDYVFoVAQp9v3ChcbMoFgMCtJ4+IQ6BCG+rbwtxnEzSoXqSH7cr+i+qp9hi
BjJX5fm611igHDR4MykbMWRyF5yRwoBTqkOzNT9muwU4VOz5PTA5hXlYw4n36X7nrkPR128QOPec
CatRYQqSEFMuvRtOH38lcWGgh7SXvq3zNuYkDseWhPRQ6iUG81kSs6QtpxsQS0AA0hAP46eNWSs5
A8wPlTmoXVem9Bk4i8P+Fia81O2OJhiXbIF8stYnlSX1h4rz1fLOjE98RJq98uClDlbtF7u6+9Xq
ea7cTiUe9mpKu0KTHEEcJ8zcbZFUaSHo/8fZ+CNVm5QyZV4ajgvKkMVzi6meL24sAWGqFl2NVDVG
igRRqml3o5QI/xBqL6GW4YkXFup3nfZRblnoSRmmLtzi0bPn75KxWCuGDTTD+NQrnHzVYgtUEyZU
xdXsuYBm0PAnf5CqXbkt5iS5Vy/pZLds8HbPV0+dc0SiCGslE6oOsV5gqP0XiIuRZ5WL8m9dccsx
b+fBn/uMUNCgoU2gqeXsnh75ajy5/Fy13yEKBnkcwJik8eaTGnkLADApjl5A2PEk/qhlIUBgEdXB
arVb4xH63QXNT0FthfV/je0WCjFvGHMXbP1UXg/kGN2VdlNiFErFnz00Jq838eq1n9E3t2czoAGS
1UwhDQDWixtg4462U1/IarP2OxsAFW2zCDHIL4HkB9xYG6PlBC7dEGX0omP57NKzGdKR5KwwvZPZ
xBTlsFfpWJSnTRS2TvLypFgS/GG4dKTHunKUM+DGjVuW1Cz4hXKB6MVGOXPSWBf2EspSfotVKd7i
4EYtfWYnW1Ol85VWg/SArH4XGiJURqQg1W0oUBIBA7xEX6F/Qi8ccOwSESS4snvVhDHru+oR6eix
m5j/skHo3Rx7Wik+wV1s6/bmPtR2UNHF1qGs5t+rLmuKp+oUs+w7jlH87s2pbdgDDwqj95dLUj9a
x2LjNnuRbPloleZoOLWIIElNv0/+NCrYNa5mgkTY0fEoKvm6zQJiNEclPNJrfmYQJsbiCOI8Xglq
bkDREh/oEGr4vg1hbCL0+ewgxVcbbe3bWw7E6p+y7SieViEAx/faK32TOKX00lS0EV5e9ynB/d+i
QJ3pE5ncNhHMQ7WVQEbQeIe7fGq72klJWaALEECOpi1NcnaqCD+Y6ab1cYuTwO91F1xLQ+s0GpTq
yi4hS8xzElY6rwZgzE2Eg8hmUsJR3kPHNYSzxgeBKEFmNhHUBV79ujMP1f85/SmheHZJKIyRPvoz
bnnEZLOoQ3kSiUTvCyv85sIweBlCe/wjLrosHqQKn3UIFBDZLXtYzMcwhf4eMAy8upI0MjgNrz1b
r4513fVzrrPkoOzH42q448AQl2NJ38IW3qxGS+HNns/FZN+Mnjzpa1I33tha2H7KQ2AgTFVsHbHn
/O5WPL0pe9I1tJ0Rva/wLwI0uBksPELaHVwiSwctqR+PJPzm27FIFeDRHj5mCKbSLczgFcxmt3w9
OMAY9VmQXPNBo5ZrqZlgN0D3C48Y59WTR37aYhCddEFYQxHuoANLpAD00Sz5619yg09R85SM4NUJ
PPuHZ3YcGTpkOpH1lochz/ODCr95146RVWUZVyKP6cOQoRMwJYTVdSWL3OmekCF+tmvpY7wUhhnR
QezFWbJ/d6TlAUOolenSpEY9zN5vhhCe56Dl7D5Mv2ub6d0BpFwE/jk9f/hnLN6kFgNmxpjgaaP8
7yViE8vo+O13JV/vbED7L4tQ5v8tlQJFK0pyFGkQr650VvbOMOhWh3vgWRwrSrZX0lK5QPzvBVvL
jyiw07eG/xuFbTdvaActCAYR0+LM5PkNprRBoJgAc1w4qSJi57MpW/9/Ql11M5NDWRKwaigM4PRK
obj+3bvTb+rvwf81k8N055sLwvWZw82uf68B0HdvWTg+eGn0sC9gj9p8/RbkGPIYEJAZIw26amOP
xqK4ALIMtXIU7hyBlbgAYMOeRbAuEIlO8hnl10UFJX828FbIRqsTxgBrTQh8+2TCnvkAtDGiyAsb
BtUXqiV/uo6heKwZ/X0u2Pa1yLicJCmOpMcbxu8EbxPwW1Vwso364Hdtn33mO5fiMPdtPpI9quXV
96vA3NDJddgYXqbWrs4ahvIrlgHe8z+Or/8QsPatv7qiPKlg6WoZgWYfQbFbreXpE9ILaWuhs/xb
IPB+ZUuyarqJEMW43y8HM4Ob6QlE1yime40TMLX7LwoYuAGravcPCuK8m80XImMR2qpFpEYsfojO
XIJm5eoJ78g9xYN0IsLophH5SI6bubnAKmwEbY2+48AOJD983wYycultp1Sprl5HQKAexJ1vwrq6
ebv4DQnLfPJESWP1qhefGkMWNj1dMejn1uaNcI2MTFbdaxSGAcbehhzpM/zQTSafa0yqC2EBldkN
Oc/lwbJ90aGWcvuNqg3C07ADWu6JYneJfF/JCb8xygJoOk0u4dt+4fe8pMkypQioUT7Uap5mUzuY
duPAZzxTcXUSQK65fjH0od21GRWbbsCFRRai8jSwO69A0Z5keoYTHeqJL3KJ8dqVONOymPClcq2e
4R/IeA4nWVEj7ChJTL8LEMU0bYEfq6VsNUmyVXa1cVw3arlbDELXYb+xchW7afkOUUoYzIg2S+yD
DSi692+a6fG3M0BGcCXE7JtbsVp80UlxXuE+Xl6EX2Qqpdnriivd7m7SEaZ4RD71/3IcIldkO8un
Ju8c2cJm1sD/iHqr1bReV5wTzvqpRtZrwdgwpW7ewoYMiZpZVvAQMUvJX3m1Jg/dEEbasYgGnTk5
FFAbkQ4hN6U7IJWRLUnWsN9EmVdjqtKjbmN/3NtzSaaZAUZ99LV6Pkm03yAHXBZ4petSZlt/x+kC
i0W22kbkETSvbP9U6jF+drXloGXPncP+sX5g8pw5mSAAPJDWlVNmJ8iblReUC/e4Ef7SiEvavN1k
eYb4DFK7p8HSaxPirrf66hMzvnwfWcc+4Ay20zyvBzmW3XqC3wpK2+CEMeC3QeA1NmCbU2P4P5UQ
7eWTLZyHmP8BbTgVFRZEH1B7tCh77bM0UE8qryZHR6QACcb00Kl7Yh2F8OKSApSTJlhXH7bXGpIB
fLX+R4nOMEzj3bi76xPHLk7XXwjSMYRrJiUqVrNDblzYQ4Z8n5X8GmcuehPHKSyeV1dVP2esWPK7
ylDzXh9fzbCtf3gsEORaWaDWOLWMU6N79vHf8TNrtjrTANpsN5Oe7l9a6GTZazAS9xkE+y1lh1B9
38qdUNnldZuf7QcHGfY5R6pFxccYNu+xpcPLbsKIzGt4uwL5G0QpwXiToPCTimf7WAzXEAueHfLL
H6koCqgYV8vyPwOunsY5F2UoDwjK/U32O9TePamSK1msa7a6Fq2pImqG+sidk3SodGjdogMnsMuo
M30Icr0SCP6AaCMDBzmtlH9b9aja1Cdag3TIdSL0UKNaGyPZ3s5O0+TDCpZTz0ngYrRG3fNzreJP
yXPh50vzPn23ZRQ8eD5V7nccijGurkYeLcORcW3tMwIrUL4MzWpwf3fYDt87KM+RDOpz0AGqku8j
nbiHI0jM8ccr3PhTXBS43cALo3VuHMWkF0QDrsrQcVnd7cQEozIERjWY22QnLCh/ulATcQvv5y5a
v768UaLnMwvUscJtW+f/ve3wCHe0vdXnczaULYTD8p06TOEeVqxumgXZaLkL3JtAOpC8a+TWuqzc
Xm+muT7aNDyOhcJ7WZ0L9MehvsMtqj55wCB9KnE8GPNP3KZm9vg7TXk4Tj5Qyzg8OoRhcFpfuPiM
XEfULhDXoCF1MvhFoq+RhkN3SbwkIYc5Jg6ZEZyS/UOMkVxPG0l9GPHxJYp+2f8d3avqFaWiFtoO
60SWdWdMm1185ddqkUAqUaot/dD1ZM4thPGr7JZoQLITZDtrz7nAcoBAQ1+NyDRTdFxD0QbjTNs/
L5X2RUbIKJAVhcUMzoTaEiEi+3jva+G7Xhyj6ikmq/gh+eDj+viK4UYMUQp8120R1fsmM6ZN33Ol
yYRESaiX7sIPmMjKJ3yr9wyreTZrB3edrmCxCwZZYMgyt0WZnCCOkCoFnhwlZs+nkCSd016rFflW
JGrjD6vkleTLXX9vv1uT6+CZ6Utxy8Ys1vhUn+Xnp8K9jgDThWWlVoU6Lhc6RClQmQumRmGEka4h
KNk+eB6K30MKj9n7NrjzYilo6X2emdG9flcVd7HtGDfoA5y6pkxDJDX5PZL3ad5ZA8uBernb8C5x
vuAgfmLeEKJ0RutKD7P5o3IlqpzNL/yXCzW+KHiD00hGpEKghEZEoE7qEhQyQdvTAgD0TSDXoy+N
rxtnTWxBQvfIqoW6rJnQ0h+6S4s3+Ng5eYLIEyc/lndj76X5qUcphYpRWFUcFS6n1wB402rau4t6
3FCVu/Zjk2EZBKKJKDo5piFNcFWrk4c0IWdReWp3P8FhCaJlkzxlGQgMWJtn4iQU2XU2BPdY3Nnf
159LUr0wFZgY/QZU+uagkKoW5FN3WFhFIhxT+vOghSh2uk8PAG3vwaHTVaWOAPHAGnevw63YTatm
cm349J3Hv5p3pBBQ68TCdGrZoAPXjmeOeXmqBIlQtVU7RNhuye+zUPKzSBWtr3c9nOx5PfE7jL5s
scPKt6MC5e+6LfYMStAcsYlKFc45Oqizg9LUAQKW1jqzcmkCjhdL8yR5x2CiaES5NpJ+yeiI2SVs
KCsGfdoR9Sm5q5AeUHM6yKD59Ff8APTdpYQ+5vvlSOMO9VF05NHoWPAjpzWVWmnu0iTS4yXsEsHD
ZSiwGPXCR+lz3jVAVhfBi/j/+h7e2m4m3O4X6GIEKQbjN+kLfjgh7vrR0xHxXnMzMQnATSJS/+8Z
Jvib75op+Bv4uns1vbDMtGHfCiDShw/VX7MnqcWNTgx1usWglvmJ1wGYF0MT0UuBfRO410gDjumj
3rjEENZXowRRKs1XjD45DEKVOuoyRAglZV8jQEFsEv7145m3YaDYy5D1ENlUMkij42px+RmERcBy
yxtr4slnnPAMvt1gqpvH+tFld/vxxlErDDtn4RcPVd9RyPN0cgnueHCNqGtYn4ufO90vTuuKfDML
ldHnQiJSQMv+wvzPfpJUjD3pXePP4acyX2gKPxYo27dWDe3glYRTOCyiqyLaM3vIBgvexHsvAYb4
a9AsdXVXmrKc8OBfUkLkST2aaesCdPs1VRD/fCUTrn1+L+2TaykqqFBtqyDIZy0yKa0o8EHDoHTF
CiQ8ZQqzFlKlny+C4xapQKW1GnoOqzCOAHoTJP3z6ZH7Uz6Xf9qUBuvQIKp5hDpdH1laRpgBbtVU
LsPVYc4Uvg3MZCYpYgTuyW1KUQSvEwzFT9cqSwmG2slzzx2jBECCm+9uF70dGIp2GBlz5RUOQOR7
ekf5PHaxC8wYfOAuwlioMIe1VjDWuLC+OAZpLzBjxd6wGyrHIi26Lt8xy1Wgp3sYpV5uBCfSaq34
5xj4d+gnK5+8pz3gGuDi93RwO2VO6pg8SH4+SuyeJO2VyUICxKZf9hPGanawvMdkZyh6pvu/BA4A
K5Kg9MoCO6YQPjVVFIAwbfXb97j6O0WqvvlUXgenR0bPJoiexMV2lP0FNyEQamHM22RgGIDRlsf2
Dz7SjawarLg+cNbJErnwNsDuxOQeTIbY4zdKf3LXUHw8xhQOB24vbjshajqUTkd9TxmCEg9NPKOH
v1pBDyTtoFV1RBgNthZuVhoc2D0vdeuOhC6/vNei0ajTkL7Tm1s2Yg+Y0dcGnmcgoSvKlOOWaNd0
r0rwEnne3GP44VKJv/IJuqWeLlUZJGlRNU3IjlU6MIkkuGy+bm7S47tujb0nncQexqfvDl70wQ6N
vJaXqCjVt8u8ZknNiy8ortgrEGvsS6EgmGMw5s/bpvZ35I7dhNKMPAiHy6T0v/XYGOo2PByX8ZLI
3VPQWKvqBnUqlvv2O1Bp2CWKh1g59gnF5eMajOmpkFsEOULc5OYJ0Nov8oLj3nTKTgUiKoYZ5RMc
F3gqJ8OlEtq2/z9YETk1KNVTlRD7eUi05FQ7TTouVToMh3fg8pTsbat1n4+XEqa/LJh9QCUiKdaw
Crx7oo2d/eIvaa11bldNFRTsOAihizQKlGuzTPjYm7Rv1A8cC+RqJ51I9IBEJUS3e9bLmSEgR5Ri
Px01LTSXkZPjUHteXFhT1b9DEY2U2eU8ip75HlUErZWATWDHBw6Yso2b37pUwcINUN2ZTRtJjUgc
8tV/p+lX72pOTckeNO2+tPDmVHObEz/sNjt9OPDCgJsEP1+ZVhmyjGVic9RzHi9yl2COhquYSMKq
/vjdxpUPo4hKAjm4DmfKsDyCNN823HgKeT5k9x+e+QJjZrCfvZM0p1Gs9ov5xEYZuBwT0cixfSVP
TAaPTcTibaWddEXXgBZburAjJd2sknaODaLnImHMWsvsasnEgGmlAcFCPkzI5KJaeAt7GWO48uNE
OTSaCsFqNIBUo0Xrvx0QWHTOyiefFl1ZOyOUxpLGvWCioNofBnNIs0OXKl6X0XZSniNMjNMwmcfA
4SWIl2ByxYiLUgBiPXadL+Ona7EoSJx5GNyCsSrkUps7cdYGCEhqFcaCVgNGiRzIV4Xh+4upIkKe
tdbnyWbdmUIariyHmruuPbyqePWW2JzWYRX9EYs1eMXuqa5nmqhwWMYL0C3lwgZ/Mvs4v/yWtn3i
1SfQpfWMkMzd9cgEHeKbCLVkdLUewrXBliLzOAGMoPWehVfWrEhhiCUr3i3dwtTt5KpEgQzBVsjj
XPQDbEx/3r1c1zAtGQ0vJ9DiOVK/jCMjDmCGpjY7dzt2vFZql6dmY/kaE2ZubXsa6owsGTRDzH1H
1UxF2JXZIQqJyqSuH8b1nQpoBic142qsvzJpCb4/CR454/qTSPNoCIdXwBT9Jg7YqsUaI4U5baCF
kzRrz7XKBE/vpZNDcFFLuncnTxLBfQaSW4Hhn8tPdXgO9lGC97ca82fAb/iL44HdIzmVyIXqReF4
eIYuHru0NIe9rhHognQoAviad12MGy30+fGAJORWC9Q5dTFVyY7GR05845nKKzJDqURIcmW4V1BA
J8DVW2sDzluJjOUiYBMU4pkW4vv020qXQUhRoWrWuJOtXjF6r9KwSKCkWlzeVHR9qtiKD0PBKSMZ
I93e55kHkf/MHil+37l9DJ5jeKMtzbDt6DvBhbVa3aE8JOWSumuBKhLJFe5PXIEPFKs1k846NAoM
LHM3SwgrUtn7eOqW+tZqtQEEeMeTe0X42LhuAGjQWm594dTIEeGnqbbI3rRgKOr9EINqvGHpB6wX
svAMFuezQa+DHDth2VFcQhMSqAprtfzs2czTWb2Q3D0ahlPm7a4C5EM9qJPYPMhiLvWtLXaCj8/C
Wh8BFYrCJoD+FfyiHtKpARedLkluN0aCQwxhan302JPfPepftL/SEhQ7lhX80vWuPOv3J+b4riYx
bRZQJ6NrH8LmeyKnplkdBLhf1RXlMJN+Em3atvtczybStzsyuNwvXPD55OVPNi59NryDHinfJBLQ
tQdkfp++txARi+fExReo3E+Q7yPm2YULHow+oJknUV9fa2V0fvIjxFh73oAO/wSKP1rdQ06ss8Ji
yaD9cJTQ3J3QF1JXRkmB6tpYru7Kqu1m58djcJbFRTO9cjinLJIFDpQ1NXQjLQewexR844nC/os7
zDXNBhqaLl8PwUS8lhCIeb77WWXcBjkER3AKdmvKVP+buM5Yvq/qtxav3hjkp+qsUfcnRRnBL7dm
qRNmMQFzuWBvAuHfgVjCOp2lLTWpJENe/sM935PlRctVPB6SdBtZMULHG2B8CoCGOn8QJeBCKHby
L8CFp5G2TMW1O5g7Yzi9FTsnT7h/5byzBY4DPs87aCRLo9jzJ4jxmkFkde7B/NFR1oaH+fqwUYHA
pHuWNM2U4GkRoQnHcl7GYgHl5MAJkL+XB/ZWENXKETHnMZZU1V52utjOQC2QM7TVT7Tgfp4LY2J0
QVfUE1Z0ss0d25f18cE9TURaRit1RgL+rPpQSaSgjEJcIxLj/JNIuHlR7Bwd5J+BPAnyx4A/LhOe
cy+HsIvxkmMLhTyU53s3B5geL9NmFPRZPdRUqFFyPQe0OeqUCmdlX4pwpttxxW1QPLm9FIIo0/Xo
lXZXucl/863bdxJRP4f8iE41pueM8EIImx6zsxI771gkliTOhUF37YWnhgbgfPfwKhBoTS//AiDq
vNfpGEtFoI8QvYAIVRlZssbkTANFagGx9MsemSlEfPkYPQDIXpmp2ptY8vBQg38pdea8hsS1d1LH
oSNs+C7RRd5aQOTuT+B1JLgaIz8xuY9M4fHK2MPFbnI1LYVS0+7nL0ZqyzO2mdx3n4IPTSLGbIXe
aMYR4mnfzrbX2PsJbqxrbrMLwFdndxmteGljfUaLrgiJhJ/5wx+3abzaYGFTFkR7opjbGgkVj6iX
J0aaLMpTJrbLkNbSHj2wpaDCTBEd8mwdOKmrjbPEmC2Hp6wfv5tyNHSdI8LzQtUUXf3QMAS2zygI
/wVpzNRslVdwH+YM0FvM3g12yx9dun6dpd96efeGUPLKpft8+H5I8Y6F7IJOu5Gvvy0MvvfFS+sk
iHkSArMwQXX6nH+xQQwDuB5v2fVvihcF1vZbPFXqCXQyuTIdaBJHmKlSyO7nrz2s83TH+T8lgZCQ
EaWXPF4nn82dJIESG//qZCGr0cyffXAxoNAXOHe/PE8UHseOv6She5b0AdGPNNMrDYxy+eKaOVMp
Qbmoh+CUR9MhuaQzcGvHlEw7fD1lkKdOR4o7DC90Lf9vEN77EZDx6rUBo4+eTiYSlEryfm0HT/4C
thcsO6pAIxRvzx6AouPFDgLOpChAuL9Uz2Y9/PSSrfcpfzJsBv8NI21u97KBgnzH8KCoaFw5OKnm
Sq0bmSz86gbWQn24inpMu6E1tWIPcdy+f8xbQ3lFlkKxi2SYOGG09we3pzRNw0Vo2ilZvlfV7Ew/
58bH+WDH7z1Rg16qgcfTIhloThlvWYxLyuds/ArqIUSmvMWSQRSKKUEPMOMZ2HdHW/btGg6Ci79d
3WK7kNeRKDOx2cOk22wF8BC9znu1NCISe4iqkyV1azx7PL1hILZ5SL6OeenqCo7czmx8jr52Oyiq
8/IlhGgUlVHMOSfksfkD/pVBZGOd9XJVVQS/Ohko6WzV0MgEkUvO//XkQeeXyJnJW4Kc+9bEB8nq
i3a8MZccRjO4AY8aBeP7Bv+UkUaQ2YvSBAPKklLzBlUP2TjUHARs5NszxqvgD/kF492U33/eifPf
U/L7aon195rS+oyvEw6i9ccLCBRAmXQS0xRdSSI9ifj/ZdFUr3JsmgUiPf6D+plKvtSJqZ0EFu1u
ICfP6T0cQwXMmKWGQcYEusFV9aGTpLoNkXSzmycJeCQadyvxa56EmbtxhOC9JPet9mzPP1llQSur
2FhaPXx1vp/XSop+jTe7yyQKOBA/LSN9829qUxRC3mgydAR1dFnOEM3O60yFYo8eGFrYWVU66DQM
wxJkVPG+Tdlcku2/R2XNhP6w7fvmFlcpRTpM3oQ2a3rDtsExcbljHqxlpb92GKzOyPMx4672aJCU
PJYeUS8R8maHYNIyF3f3Vods1xHIlVTivbm+v+M5+ibcoHIvki1aw1yOJTpVfCHB8HXl6ubOv+zh
NFT/EtoYrvgpMJBgTrMwVw5CkpmZhGV65EZxV5OOSMXjD1o9Ph9d1cX8EStPJkSU+ROWfyGnmAZM
tuEV0y8an7hNTv9o/ZXNrEz72E3MMzV3PWG38zV1qujt0m+K8r2Y3Ihc2eE6FepNhbMIcgzsBzeB
5yG2oEbonVQV4YNaUhiIGWPYBvdskh48QuAESSFh0OEI8v4U2rrNh/vpvOodmjm+c+uXRMI+wInO
UZjhSyi0ZH2+gBtWBVq6+dpyDXQY2I7Bbj86VEFn7TiMSX5WznqVyaOdZbX/u7GSu5GxCzg/gIIv
XupbcC2yhrV4OxMsOsldllZp6We7t/YQ9V/QiCeCPzoCyQHEvvZa41pGPz+wjFXYXS1622HA1qhm
qb/VEjgYntG9SlNLrJ/SnfzmG/5+doQetaU8nuf5mpOi3usnjfhZRtypwtb2EgynS7UVhOZE7yvn
iVfZc25uNpv75wn0dznC57+kzWsT0pI1DfeJPStdnb5+yZ2pQGoJmafqfL6ISXcx1Xx0jt+WiaMN
GZSnFRkSmcwnRs2H1wKD2ipize7mHMtOgIlbaIAR3N36HpYGaxJGuQdR1iwbaWHz1QmRlAuG7Fa4
LsKNTwMO2YKyu49UBRrBWLZXzjdtgUAPWrn+I2roSdFET06LaO6PMnfr/MvpHKjhP3Qz6rgjDEUV
Hx66tbBAh0poleZmIMKR3vqnLzp4dt3e49iw/T/lFq0yB48a/P+rMGhA8nzTq42NDZKYu/Q1SHMv
NY/DFkNSlgKuzLNQpF7kLSiyItyQmOOla0iyajIAaEluM2KOXqbfy5lQSa8BCYybTl/e+r7oNqG7
LbZJ9VyHOL+HvsxI2Q6dVKYT1U4it7l3r/BE7Zg6IpCTh2/DGTznDnAB5Ot/+oEZh7eiUj6f5Rq+
M2d9eD+MRdqhshSLw21uqBiVFEw9aqJ7ugmiZeIOd31QNfmvmvJJ6Mg6x06vZ2XWebTeE5d1dhjl
YMG3O7xSnI3HWOX3gAWTdXfln5pFhvw7k/0K9SGQb5BWVKLuPEgicpuao+8Cgt2q1kFQFfbBpN/I
cPQ48hE+Cgkf9kGBzqMLeRvSYBvUu8xa4N/f4boB34yfYsiDkw5GfRpyL5UGpfrKqpKo/dsuFa6I
CmRz4fDRddzLizfkg5yIURE0R6M8v6MpDutSmfNsljGMmWsC5PRRHjigbWxC0wcnYNlO6tb9obbt
wdZWVr2ejW+x1fTaWR31FLqn6UvQU74zpn/76PwzeFcjbfyeKbIvhBZ9QtZbpiROuD2j1T+fBoJh
Y4jVHeYak19wN5lu6cft4LfgwznYymxKH9jeUraiFem237uLkAc4StokMPtPxD59/LxRQXWYX18h
WtToioemF2s4SUMhLcKmCOFJ69lJ3cCVmN3Fh1ppXGZku582Nh+s0mNEu9KzoLo+CeLDSqidIkgY
4JcdtsFzuEG3Cl7VeDZLkdDrNCioKJODBux5BeaQUOQ+6SnnmTyYs1UpJMsQYCUbW2qIO2nAoXZR
Z+PLENP/bJjG5DekuzTxq/L56dP5K9ZgTSfBnJ2XeRr8ahxpM/KHWDG8JSOvM4h8nUyG6eQtWpRv
fDz1haInZeet6yosnqpplASDfNhSvc51qIlYlA49sP4p7NZBwpLm1ny2rgj9eJepYJmlePrk6CUt
vSG8lv5cMEZ6Tq4DpC0P7UrAyFCWcoYKTN1VW49EFtj1kyqgOh8BJ9jVB0c0cUsVCuj7bECM+ial
SnlqsghOY13s6SNDb8zCCw8l/pujVitrENcGi/+LXzKXt+tMcbiK1FgWGpwGFx11AY3rkQB2y70J
udvobLl4rdMenx87ibRxsg2Z5nDipn6DUDl5jptfSRKQNoJadO3fK9Ca6nOeRUi4oBferS3liiMc
VS9pKi9Jggz3y6HgIXSKkpkfFToBnEA11B6wuB2njYLTIRBNI6IxOsRkZyvaSW0GtRNn2HH2JxN0
kSnfK5U95t76Y4qAJRNUuwPHaNMTmFymZ4x+V+4AvT8lUtoihEyWYdshMk0TdeDmvDFfoz3hkBPy
Lm7Fxg77QITuMuYBI7LvUSxOacKvTjysKEL8Ur+UNWUiB6XHzFsFCnszGSnclF0yb9vGPBmQLDiq
B5Qx2Y9QxZMeNHFRGkUHY42p1od21g4sHUco59Nkyqmrlb/Wta4mCk6GLzPhB8d5AFaD3BAO56qz
Mka4aK1tqFgan4sfbn31uabFpexqSx+Hq1mwK2qvK6Iw4t0csPna03PgSLXWyEDztU4q7c47cV7l
6sMSYLwXvAbWFh6eSH6PDUr5wAoyuFc/nYbbCUjnRJ9XBr3fpvnW2r5HTZjxwMPnwOs/yYaZ05zY
ELcFuVh1JI+hnypsXGYL9S26AHKkta+cvo1B+DtxVlHIBqKaVtRxHqPn4OGUIgKspA/kr+WtxMay
/C3rtYjBPFxS6REtFDKHcoERhyTsz/F4H7DlMgTEzFSF8/qRVmQ7EuhfjtWnbWcWD75KBQnuph8l
2cLVWD5EwXoTQTL4X/LJgx/au6ymYJYV9G8Vl1brQ5/I+Ll/OU2OyZvIaWZXTO5Nf47BEMvDsTSQ
qXlqAg33kLpgvdTNqcMue7eknYQeqckPy9Cu5lwk+0/RSU/9CmO6jwXwvyJMwuf2lbkFyKbtM8wE
SOvJU0FefiXlQiDeGp0uczjNd8UQA2CEm8YEH1mzEjT6jX6uTD3hslKEZKE2FWD6KD161/VkVZoM
cFvHq/WBOlZEdLVq9efJAefBS5db8iUJtBboFz0+ovcVObf10z3wdjsIPszwbvBwWy1RxpUUKzWh
h+oZhv4cXv8dHaMLdy17NyGE8u8Md6WCpMN0CWaFaX0OSyxqZWkzTWdxZMQq3Eb2HOA+5nNlbLwU
prF5U8wUVNYcYOrZJmboye9CbOtY85PaEnDhtDWhcPszAvPI5uyFVmAr4VjSNDoMeUAaPv+dsmtc
r65nrD+jHDzovbT8J9Gx+yfuI0hQmImuzF1+MiWTpI8AqThB3qDRJgmfQ16rhLMJlHO/bi+8XOBP
/8meuHDFrj3DQ1MoWYeq/mX8zTgxCei7D2ZBtW/BVS6MJrkLG7xT+0pERCYmPLkTyOsKU4zYLeTD
QjznNBfuSyjWpKvmOWAMVhcHVBctgIDA3/7RXcwocG8BaGNMZDMRdB0Eh9xem92jxt2i0JhbWC2I
MzdfpNoj4HZVx7jDwFFKKXhnmfgpIgl9hFOG5HuRfJ8lCMeKapw3YjWLA9re9Rcnrjn97xco0Ctt
qL4+lcMhud5DRvd4UwxVn/HXbOtxQklqA9H30ZEuZez+Pfg1K2YE7/QZ1d9CqS6gw3NCnKXrBG1U
JZJrBoS7YqDfyplrXAh1emTPUMt5uE+xOUgJ4KjqMAztatzRianU+8xt0sIreDV7oRKx5hJ1Rmbm
cPpVMIoW4egjuZeMYHlRn+yI/Z+KGPrJl9ZgH6u5sDYD9uey9TsYiLZZB0+XPhOlpsMXkE6PkbkV
CVqZ+8N5ZdUd4Xs9Bq+BldS/9HsRME5oXThEEF/PTIFESnR8YC2UQzcT0cyirMHfALu1zkXXvyF9
5iMlU1/oQ+qudiIv57uEwZPa14ZMCLVlrZ67gcxjJNQysNCFxr9GemSXq5LZovryyGjh//JeD4Oz
ZgxOxdvzUM+diPJKam4vtOkjaT7ig0ktkfVBgqWy7mgNjKW7PrCQA06xwXUofWX7vXDhSFezXb8J
G4XsneDK3+Uf7A6JuULm1mEs27yxY2fes3RxMnBnjnmxaEEDQ2pvQ2fAO9KEYt17Nq4V8rYvR2NT
/DrMF+vanJH8MlD+IDIOGL0JzPtXLgRzHn10E6JIsRichh4Kl640JKE/Es/Hqo3w+WAtji2vx0J1
6H5qqQAUyQYAmvKYMJeXt32JJuZ+OEbwdv6u29wNShjYyu3ApOSVUW3oIJkTj59OKyHkoIAA9+Km
3L0t1lbf/FVRFRWJuKnzCurGoR0k/xzWDiHtNwivjFUtvnZFnvcWYT2FvZN7PKGA2AcOr7VL0e3e
E2fRJComddEUlOwvxbJU8ZjzDcMd9gIWSfRnqDjhdXMnCAwgPX/xH1J9OwziIDxt/sVn3KDpKrFG
u2/GuRGbq7h1OmepO443CdK3GGcuEKrZKp1FUkCWpE82uzv3JOGpcL8w2Rs+xX1Lf0Fgkk3hEaJn
36bKlseZUvxK2s1mmTxgkzsmKuR3bjGhi8YszR6SJKOwv87viRta9zsu+B0Aejgm/jqBKrQYtYcn
HlJK8e0xLMRR+KsMUYGxkKyGq53P8VizqKIJmGyLUAIcBXWH4bwaGywzSPnPQcf9ADBiULslSuDV
jipUN9gV9KieWdxFlZdngfrOmPPV2YaCYe/tmkWHw9vP4i0Zm/C9aBRu1WJHrXIvw/mzfx3mSyDD
80mCjTEHIRIYh0MkEBUxm7g8BLvKahX/M9SNIn8mFRkxaOWF/TqzUMqlJJHSka3IN5aVcojXoqsU
n4HIYQzURpUrHqWM5fvxen5v8/op72HBHtQbpkNcuNwDqdYoXoNaNyBAyiRqlGgmrFcjEbJz6KTL
psPbE0EUH5nBn5gp/3RXugrfn8RFMXoy3N6Ozv7GwKwhMxsk4ZGeGufhEpIW8y4DYdVFrVASVBNa
IYzOA31sOZpX702hdOG9eCUatjhTCA/UFrQPc9tyAUryLdjYGM39Jjdt7yZkb2d/31gjOmajyrQ0
VpBCYRdHFTLRwb/q94CxbJqFOrbbSFVNHvB0ZfB3Yg1W0XAP3daenodZrFlOUYgsu+ZhslqmAX7+
ZTXzvMjzE86U/tzc6n87me+6EULZaG9MTR0NVL+sq8daeuihoJq//5w/y5ScTW+YaSuP3Vun/k0Q
r3E5SXvGVqIXr8Ug+nK6uESyNRoUhHupz+MgKl3yvhTPoT8cF4Mu1WjaC8yPQ1U8QrK4G65pia4g
+A4oHPzWQfnr4dGEQAvVQmjUDPVMj43Aq0VgjieEMz++ASoxi3vWkj00KqI51FIMkIP4wfApVeQT
HiNKnTS4ptS2Azem6yd28Lb22TJaz5J4bobIp61nl23OumfSvw9bVaW1VoeYDiid6TlBuLvBoYR5
Hi3jUgm1dX95nd6lNX49ldhod0ebIHAsjrWpJom+ADUw05yJHJzaX7bVF6RtGDySsL1L+fvLLa8f
ygB8h3l0v78ekMyoP+KY/Lyf5J9g6bWMBdUzrpqcroWG3KtwgrmSTumbrrLyDAE3TYQnfjQt5WgZ
V0MctNmTSCK9e+ARxGBG8lnZxNo83QySUTe4CAFvkAIcAH/Jw6lRQsYNqO8iA07RGE30bYzkiENY
aXvQjEJu6sZwsJHJ5EBcnYlMKhZcUkcw6ZtKFkuDgHGQwRFe+zLjYp8iDkp8HC4S3DpAHPDEMi2D
sPLOZtA4MqG46Sbl5IAJSHfoENXFxJ1W4eVqBgNn+oWyU2fEUElZfw2hD4NXrp3efYNWWztD3Tad
IXRO6yS/8EhkXwOldKiPEZzOhI8Gu4qvnGZ6z5LqtS+r7Yqhflck5111qPBbOFDXIYReK1tFD31Q
D7EKQ6R56+uR232e9HNkZl+rGuLlGFUcT+YuVgauHujeQxeLHS2845XuycYHD50+Cf+zcHGj++Lf
ejVEaWWh9YCTULSkeYJHqP6c2vQDDPSXy2Ja+5N7CZ39mWl/m81bcxLVSe/K/cmRRLN8OAKGWEBr
K/erTcveE8vHI9/YxO3UFxYog9WchMHe9VpC3hMmcMtPb0LfX9k16va5HZlrrNNYSTJ/pDPFp6hW
/OWehsMcmH/fZiqkyO0xM4BAmSDwzC327MX7+vKivWOYhzkqpm/WL9k2Z0H8FFiS4KLSbJzcB911
RhSVCjXEuoTWR9Jlkv6shnf3KEl1GY6EepN80aeP9KFRGwZSOzrbNNGmXVIWBontB7KP4eCeay1k
Z6liUTyRNxcodFMT3DbOMhMtw3KrnKKgMu6Ix9ATel1UQ86fU8YiGqeYsbmJvrcBKhx7kUFouAkV
NOwS8uBdoBUUGk6HHM5Ogyl8rolpfjWpKe7MAwIi8WbZrstfL9DLakycJP3GKiPFAqltHjo17RK6
5X5eGS/r6HrFXrO7yESACa5/1U7k+CBKTUITZQebWAK90cLqKrJCMii++/xjHBpzmVY6fSXST6XU
5qcTqlH+Ztq0bZ51Sz5MkMhFUJgcBM85DybCVcHAHdDuR53aOr9/zzRWNwRhCVA/ZbvGYxKQHGmJ
Mr6JV8uYZwXKEWeDUA+GztsgBnSYYlxT7VrSRR0EVtpddPJ0442hsGLfBnudRaDYDBj7lSFvnV9M
WbYMOkd9LXWS4hhRAjxVtOIC+5zyt0F2/7JpW0IlnknUxRFM4zc9lCJmGaoJPEV/FGrS5+DWB/k2
0zMp/tgUBzWS1nZcq+bDSSqQIXBKGS/9JqGJPrPfwTjfMSi+HzHH/kKx6taw8kvi3YqGXLr6oRDS
DaZpaoRV0aYQbnfkg++DlWmoH7IXhJs1gKQpOrQjC9g0j1kZG4nNE4hFHREsDoi8nchY2JcPNrQN
SnpZQhO1a6hgUcNSuv+pXozCh5e+zMjYy1MBPMRAkQ0uA0qqgW2IdIBYoIS0tbP3OoRmLwoJd16c
XMoaAuJa16qmbOXjbdm9UlRPaIvbHNlH5gL7J0fnaf9bDaD16wf75cwd+M5qZRZ1Kj065nbn0tRB
lHRCgMy/1Z+xJ8DUz4PSAQpNZetYhCf6b0C4EN5CZNssB9rJz4xUqLOQHFF5HW3DVv5M2TChg45K
b0PCLdE0Z0dOY4L7vA1+I5DXPjffanvitnQyWn90MO1bnfHUA2BjTeAhGvN44Y3rMCT9w6gH8LNp
r7h1ZNsOms+m1CrhumB6TUpJx5kmX7I9SVd7hZuY3zKxSMOV2pxNkHawbPptX1WauWbcqELgs4v5
/EyJO9d+JKqM0YyWnGa3ne4MOo5ZU4gooRUbZ9aoEZwQR8doycp3cT/t/sKVOoZUe8nOkK6f0B29
bX5ByBj3+gXm2Nja+WgVzCZnEjKVQaafs7/ZUmzkTNtosIn2DrbU9C92O+BdL7NOR1Lue7LaIRnj
7TSG2Q4Nf2LkISS+vraOwxXuCO+UBueNtkCLtzNfEiz+3UnU9PFSy8Z6lV4Fagw7v/u1jg1Ft/I/
24FPTG1VTKLqX1eSQr+nyaud6E4259DoelEQ9IucAv0PzMRgQrAM6DdcmvzGpIzpC7DFibCl99ml
/PZsiDoUrRYNSe93KDQXM4/oYl5aAbhloquhv2Jeq27FuZKB/9JCM0XNiETxRgD+COar2XArEB+t
HRQzZuGZcVhZXW0tt+B5ewdzfL3HjsRJ3BaJpLAOTm56/pvsY65vCuBILOQ51uhrnvWCheTGQVJc
tF6ruZC3f/7QaVVyjKfm8JPUwS4167SMvt1C5pphypKjLtKt/N0HZoTylkxp/b8bnAwS1Edkf7bV
BzPHYoM+dXGdAGUh9CaocXhfMa/yd6GPFUPkjKSlzFzjiG6u/MDgi9gL04p+XeEgrkImUpqD3yIL
S4qXecTV0DSz8o5JYTkdKp3DLb9RUQZ9craZkfzzDVdON26ruMKAGurD+yT55mqEtVwfuN40Gzqu
cRJ88LxYEY9RqH2EBMqPOqxsAPLkgxrnIjuFX93lACKPidw1slnB5FtwLEPayoF+69HEeKN8v4fz
DsDaXYXc1fYogMZ4WeMGLA6/+lfXAYRHP3KNWpaSaYoyZ4P7rIoZhK6VflzI3uJXXmwv/2dTz6FT
OW9BDTJp3D5Too6Nb9KqeAYdSSiXWToYjYq+mnjx4KAUkZCrYFAfk/AsuVhn7e6MlxkRxlcNzIm+
+ZTgQK5Sp+79bvWMwUAOKDXf9GNrvjHpZQqQEm5c63F56T3OXO2CXI1362yA4jHUHFxh1xyeZOA4
Si8pXVFODSZIwFM26jOXekIBvDV2WJwft7i603xMIcwHGhhRCGxLdlh5bMfcvU4jmCQLbHw1IocC
BEBPXKMZmpYTmlzMADkkcZK4MCgOAaV/rXFbevIiSubigy/s9rWiGjbCGZshVPBF8/xJJXg0MJcf
eCkPFfFHosJUstM3pSe9WK+TLJpgYH158nPHAUcFGB8QHcaZe3ZEXypsoj/f9ZNib2ECxS6iWfG/
SReR42SIfHvEnlkL7eV9t/xR7TuQZsqF2BBnoVdRzWHBDZf5FO9XwiW7TvM8EGQzsj0WUkDmybRm
LpLfLMcsmyghE9mij3PtKrC6VyyFfDfpVwuGJ/eINHed9hHRp5TTcNcBuxQrSfbLKMyapg9y6oo/
6UQobMqEYCOE4djafm2Rbbxp/0UfgiNHENm0W9HPe/ob5pQvjCPmgH3rf/Zm/G6ddu25q9YDOaQm
6tV9ilGxK2jBQCZ7Ro7NU2kWPzjyzBqJcJjXT7UmusbrCYW9Z/IeKGFecJ5Z5Xl8xPT9M5sPJnmY
2EIeI+sQSb0yhIGuNQc/Rkv7pDoAiwNDt8o+6RxszII+y5pGmzk5M024kwdFEDjzpVxBxO5fSN9e
LX1agUAyEjFMFf/d83RsK8fXeXMgf4DRLfFMQ/gayxGJsFtMjdb1z9OPOgSZZT41zHIsPMihGRW5
+JMcpgGXzLVQvscJXTnui0CwRq0FyFlDhiJ3AdbRoRbpXtUjNVGSJ6Mdfg1yAmA+c7CavdYctvRj
Sgly79hwRo9X8RFsHVlUIXFNkr32rVpIHUuYMLv7rqag2maehNJDZVxwmMEf986SCDnXzDKO2Tbq
l+PUqll+b9GFzW1Gs1LaJl879iazOGMo3l+ZVG3pHpkFwPlpiMmslZ52R00JIWMloISR9pnIs4JG
mqTZNWzAxarjyNHpxrI2Kb1yW/sio/J8RQ4Lr+BMJEjhOkx1dDTVpfXGmmkyeeV2gCxrcEFuyGXQ
heskNDuR13LZrvXL9tsO5ZRz4kOOC3aCHQFu0U69HnbO4dgu4nzasFIr8MheyVN6KhmxNMD3xS+R
5JhUy7TfXAouRKhOW5k3otPkIfnFvCVq1uLU8nSYHiYHvhCrdbgyxWduYnfmDcMk6jvA2ti7vlaI
6zln+i5AUoy+nElDxQRppCTQx1wPZeVAcgscXKASASMYOtzs5ZwLb9uC3w+MESB8pe0nlLDoL4Y6
CcQl0SbmyReDcVjoRmPsZpt6yo7D1Mvs/zrx/GFlGH+TTMhKMAxUnbVk+wKawySykKb1+ktnE52G
Gzi43FzS0GDme9zdOaO8lQOPewGH/ErKGaPkIzKCdAwQ+7qHsCoJdh4dhsLsk7vg04H2AbigfDSs
Ie7zFhfiesYGJGJqikhWotwOY35JO5HjmvsT9yAPU8NhMik1n9MnxBWqjFPD1s6nOtRsqs1R/euf
EbnaC5ecCBU/YjD+5Eb65EXxGfPysqExAbsd/XEelARTKNKMe97PWG+Gv1a0m5UWVGDYP/1OkSmz
Ub4cZi9qhNDRql6Urpbhoc8wB0HTNLhSNPdrp0mda6C18haBur8I/1UF7DiFMRjjjOKLu0TwkBCB
pQIE2usOy3ucFwYeWjA95kODTVaE6ghR//VfK7w+KmzqMbvHQ4M8BNCHgc6viTZ3MrcWDX/eNDBx
B9P6r3wwxgDfJkHESuUhXkNCopDfB2T5MMMizKVKbsnFI/tSUc7SLfuw115UqEpN+7KZZHTc1uFR
NsRfeUhmFth8NpPjQljGW8CZHouy5JmqV0sjkvX6bBaiUZNXnEXHO+J/9/8BpsQWLmTQLxZ1GRYX
1D84koWj6hIZoIBQRAMRNHFEpr5j+iWuu3jVk4j90Oz5VK8uyE/e+ujydT5pbq5WTfrQB4hvOHpl
dX5a70M9nMDe1yWvyBkMeMHFDCOMRJ/wPcw971SFK2oFPncALH40kJd8d+dlHRwJIElwMqQJH0In
yvHQRODJ5C1p8IdsYxhRh+kD9F+CNZsrLLhnoytit2zlFZ4oY+R1aPpt8/0Ad7PS0ckLpggJuaHD
eA3oh+yZ9pE8He5XOBtGitXMs4uG616J9daqs3D1+qDOh6R4kPXsZymlvpKfbrnPa7NK2TXxdYG2
OP0vBTXMkSmmu1o44gWGnDbsU/kQ7VdvLOWd+SW+dy1RzJxtVhdLiGonjANfl3+FnVf23w2mFNfK
5vmb/9Amuyfm9e8BAGpVGHDdnxr//+s/YWLU/PLusmNHM+xH7Njr3TFtAvpEdg6bEIcZz3yubVX6
XU7fGmqTmpF9s0ct/0LRfN8dk1tNgGhuYFgjFV1WdjMenAX2N0A2SB4hUAqkf9GZ/gilQkcVJZUl
lAt7dFcFvPanItayfQJD7H1y+YK6aY8KNcNlMQCQDZChNJePAHR7aamM93V042vKp3EAWC5CoVWv
lPfAIm/T7+6Zh8Hl4YAsNidfpgZWOuoMe0NBFgKUZzj8ZRSmgT8tFc7ke2DL8vP49iaJrt3GLiv6
i8rM+GotmNDbJZuKb50kBOzDdDK+ZOVAG4XTHsWQL+DDbk1jLS6vxi4+0r0+B9pYdFQ86mHuGgFt
3o8StVHtcECGK0nqk88SgiDoIrULlpKJcqnQ5frCMk2tyPW8gM857uPDlfiSxx8ir+Di9QOzdz2u
hRrwxphzhLPe6JMf0ONgzWbpvgdEVYsDpBn9F7FAayWDjHDKR6OdTcxmDn63f0Dg5ubVqmLN1g/G
E8aXiPxmFnVE/JBV3mwxP0LLkb5G/pzc90auydWfwg1gGs4XLdaoGrzIPKqk+s7USodghfmV5ED4
4W2qp6rHOp1mwaugUFamNjhrxwazP3fhvNJ0XRaHyG1vzsFTRDN0OUMr1ButhKzjcTkimWOBnVAB
/44jt5IAlrsfX4/ou2HzgGM8bog0yXizgpSJTzrV4bPdT5Rm7z9BJvS2nK6tnb2rXJEo3XFFzMiS
CAwxEkSzE2bgEIjDGHoX9N5Zrqmzg1tM7uhLkeMg3QPblkZ+zHJ8Mpr3nfpmosway+jXRxfZQpxl
rAQK2nJZqkdro8hXXU6900GrQDyQnV7BoUxoJFGwxc0UdmIu7Lnfyq2RqyYm6z1kyqUGYgd/mkNv
NbQK0ZTqnUfenHrTUf3gSu23MNpGEoMSE3ELnmz/7A/Y9hIEW0Pv97eet8yh2tHYTFT3AIPKOnzS
0vFWehhob32NFR9xsZYyVflS0mspGX6jpkur0tum6820tRgWfSU3dhcsNmEGs7154l3K6DY8k0u1
HW2Ix7OgphyFvINdjvjfemHMepvqm6CKgnBA1hRaG4H1FAh6Em0eu+RKI+YQxIXHwgTrPMDmV1ib
VU9zhTtoIYq8Ej8M3f50E4SwKrABA0KjzKmL6ScxjpsxVw/wc3LOJiVpAOcSWjNJFRAEyucnSL9l
5Bfa8hWy39x2rFeT5FYwUZ8ZpiGKVA4BsO2deXA88O+aUgSG7el4h7fTObgk49J0HLuvohSbxfFw
8EeMM8YpCNnjsgJy95XcKf47Av6BHImPDcSPlvOG9gUW4yUvOg2YgQnba9k5jPYZVhQzzmzLXTAK
Pu6a7R8m2cq+54D+xiVdH0D4RRtSsQlifjPMZ46XqT9dqpYhxzieFTSWMfqd1twH5WTPnwRHyusW
febrP1x9kc1BQmT0mvaluighVmexNdyqJePXTi5hFOgDUzC1Z5EVO5rmtvpgD0gdOspLqBSXT91p
OAf9/GgGpiV2ziGYegTo94nYlAfBUfFgl4Ep3Omdyv4gOS/nb0cyNQHGo7wK31YRXFjfJ6EE6PQL
vV7oWmUwiB3bm2uxZO7DvyCIXNV/wctMkupgNk3D6ywwktNwTcF247KDV0XMBgRS4kmntm8uUkPt
82vYQCcZ56FHlzGKdeHRLB+5DEdyrS5ZO1eLn5d6Pn/tf7/PSVRL/Dm/loIQr5IUVohOCQGOhCAL
hH0gsvCVITx9Iin8r3wW3+wiEUtwvGTaRz8DVJU1KV1z5e/+BBybiNGx3lwpLK31azj/3TfduSFa
SwLGdm+YYNd5XEijyDfwU64RoA4EzKM7uERu9coQaQ0pUUjCfCj02kyhn2tPIo507ytcSHNCslvt
vZPHOwG6mV+k5tDZk3y/R7SZ3eTfqOAvgrIRvLhzwt8gsEQYYY/P5CBK50DOhjQk0CAlqXB+1zvb
Mhb/pAH5bl/qSLMdPKmoDcFZ17jSi5YgeLkHKd5rUNILBb0cRhN8XALwCpr7uiLCQwd+j+TbYVEr
kumsGh9ChBQXHd4CYszw46pZ0Xn25w/NMQRrGpSn5J7Wn05Od2b+RacumfbECXHIu3uaMjeW1i0K
uMk7ZSsFW8w0APTM4lPH/qVRCrGnqS+U2/3goh+vVG7XPdib9GHtOj35jLT32siaUMNLmRVdvYYk
q30wAHFhyHUX5aSx+v40+Syq5buHGkZnJ+PMG3d+xzwFP0BGFgTxZYR/Hbp6YIFynOanpQdbQxxr
a/hQHF1uavW5YVs8Eh+f7M6Q9Xc23T30ad1tLvW7bOn0o/qpgGXOaV/khK3645pQkq3VaWFbbWNa
8wGoBt4IVDeYVJN10XmgZ/uE5WU++JA7ll1P1JkSzXokV8Wu2e/T8IjA6V9jNtoM09GBpiZx+10L
NKooXaG6GixGXDBh12cyFoR3UnTRuF7cP7vnjXBWY/Pz8iNkoP1kmzBsJauofJqzrFCkkzzUW5Mm
n1kLm7lLiVcOx+5RbBYN2oi4QnIDglqru36E2bRzIGDpDW7/vHEAIMoJTneFBCmKPUN83XS1Cx2R
bTfZklhK4pOerg3Sfk5pKVRAmni75APCTP/4HH5b7TSNDudb9HiJIzORg9yZusVNZPLtZjXvY7tH
JhMvwbg02ZCMIu7RbNmcfPwhz3m1XZWsXasc4aW2qDN4zz810/DmKrj62lM2cyVDRUv3vE7XTe71
kCOQXJC6NWmTtnkjLx2sMgJyHEbuzDh9SPvcZ0if7xRvye19CPML0R7ZRTXFk5kTkGkqOwQcRqz5
bQh3jYuwk0SqvBSAZczuYSrkQRm6arOUvqnTEjnpBg37OUwWilK/ovEwNID9wdbvSRDSgPT+uaxY
CrBw8oKj3jIcOYiO/+hyrgF+efcAzyv/OeTol2TlzDS+QWA6keYlz9IrGQKBNxGAKAXHAjoem9r2
whuXrq6lmYuGxy2WfbTDL+HFkMukrnWbSARojaxulSBIMgw7lgzq5DfVIpP6UFmuYISlmRZcqdwu
Y0mfennnGvmyP+PXxL1lTRscMuoQEYbSTWn+D0wVFlxRD3zym2NCfngfzFRfNyHfIATS48dJiHNG
6ZAP4ATZCLmwOVpoICV/YMsfZi8Ena9TOGi5GqsvSGDPRRdrIORJWSmQPjbOZEd11c7M+82icP2p
iXs5ma1UbbDIlJN/CJdpLfNBArjkHSWG05iTfIjI6hPhiY9EaXhiWVf3qhuH9L5Yk6zeHF/hBbVF
UKuRnh63PD78riOKdcc09PKXVfvG8skWiipz6n7Xq6GdPAIAWMwHHKUNd0s5b1voQghlIcOQ1ggT
zpgDRtPYL3humalzIcPQh7KQOH7NoCschTBkinOmyMKtk+lADF7y0zBOKxL/8FyVqH1LtBWNKXGl
RWqOeteKGKIHoMnBFuYi26GN04+Nzc01bUE14DRXLwPUh6eSZj5MHKHA/I08rVA5Ngdnyu9EgKyk
b2q3YF9axLizs7QGvn4Jw5CD2blAAaj12aVaqtfJfj6eTD5Uwg7Z7/NSitroxsXnaOtIx3ADkq5v
+1C9vRffO+32KyTv5q0J6jMdX5URywtiQWBzzIYnXoh/ThErosrVT3oGnig1mrhAlc3D3D7a/y/1
wX8ItqezMGi9OwiszGR/5r0vJ/t1554VtYeRFIRBylC5QueGnG4q/blRH7YjmKxueTFox3bFI/Sv
foXa0iG0R0WHZGp4ubTIx4PNYngrhLWE5sSNkuFrOEwFHp0w4zRj6rkMWCCQgcNQ7oQoSdtSZIH/
6J31CNBSuJEvMbJB2SqP8s2cgzmPymJuOEndCIEhvCMpMpI+aekujX8SvUExJ5q/8zu6vYBRaM8O
Ix61TC8Y0yq3TBjjbMVdUQFUHvXS54wUSRebelLDL1udy6wUSVveNSAdPIL00UHM9TzC5guX49lh
/AQJvok7RxLuVVkN9ge5+B2mPu1VRSoGGQmVMjm3Or2G3t6zkqf6STpSHAB8ZHmtnJXyKd9T1zY6
Vci4gcu0GVco4kqCiA1EsbrccL7j5bHHrYnvum9TkGyDpt8QKHu7QOmnWsqhBdaD29uCDp16UnVm
0/8zcwy8Rcz1UCtDeo+/Wsm/aufxv35XHAC0/R3xmXYuO/V9dPiXo/hyieO+r2DSYV6Pols/BCXK
UO9h56YcE4FfsBPKxpFQjwjpIpSXzwsN5TDSYGx/MdQpjla2/Hug7Worr30Ao0MSndhwqKEil0Yg
6zRC4uC9lMVd6hPGEKwDf92Wow0vJ2n9dRV2O0cJD4iLNE+0uJfcLPp5XY00vpoFLKdbli0YFz2q
196NN9o1DQ1Odh7vjfnZeVMBhQEdh30Bh3Jht0gmP637I7XtRwFU828QzxaCRjRERPdDplh4mTKy
Lagi7xrvqsRvL8nszZphGtNZzTzGwkeVtiA7LgiIoAf0dPq3K7ScJK5E5E0IfzthIFF2sGEEuPlg
twP4QI6kjzY2xC4b2E6A+taVOMOsd3L9CYpMKQ7pq3jNE1QUEOAqjm1hJ3LjFguvYrYkfcU2HQQr
29TOy7FlnR25hdJ8g9/76NLJ66wT7QKYhwF29UJglhQDIGOq3QaW8j3dI6Se9tEzeYbIAFjZh4DB
hxeosTRThQPrevZi26s+L+7elGTA5bRUWCdYeOZMF81KK3OnxzQfeCtqBbaHbIdsNxGujfPtNCwc
0fXASPHyGcQt+JDz+yw/cNFDqTiryfWaaMpHYYfy2oVRHu0nGx+EX9kDPfIizOu1Ai2jpEAtcoZ4
SpUoJnoSPkJIMIPQZAiZOsS+nTIpZQpQ5Trd4s9ezWIwbsxdpD6v69/MTaU78KxIQAeEJno5FQDL
oSqLZL4LqNblVX0Gg6JCcpPIueElVLj6LWbrvFawCisSRGCgobg0uM4D+zgnYzZKkvEEz0LgI0Kb
9V68DzVqEQjiWCyw+8C4EIr2KNylTDWk7X2cogp2OZvdYolLL/R5nxWXBvh3wB5oY8TI5tqHIfmm
jNlde5Frre8XPo3MJxcLeHGHjZy4W5S/b4W14Vvl2OGS5AtcpYM1Wq7mO8yCdC13gDYpkbKoDBcd
Smn4+ORXld/6dZK3UsJ6zSaC8xgae2ZgyU4HtQ/5WOHdw8lYUUkBZSseXgh4GP6xrMoCN11BVo50
dcm/OToXIilKCmFYiUMB99gam5RjkLde60zpHyQIE8m6gCjsGQo65IPCJOZ1n5bFYgG17gl3ftCd
bRuV6wjjdAqEG5519vlb1QWvzNS/qnq7zmcYPDv3Z5aX3xS0GYkwdNJKAPHFbIARzJ6eeqPrYGLj
UIx3mGzQyPw+03BaAheI4KjMYcBeQk7QYZ9TxLJY/PSTrRTg32LmqAf4EcRkE4n8okk0xjc2+Ea1
TDPswKqZq98Cx7pI9OB4HNUe7kbibbwOoIpL3iZQ5cJ/gL+A8z1Q79msAXCpfDkIcfXLHCB9+bQR
ffuKVg4GrbdKEW+ux4xgGeTRcR2QOxxN3lEdZIjaUkYvfbTrrK9RKqLtYcwLEtUfD1uBALcabcR/
mmspEOW29dKxGs9ojPoIwSeEZjOZGg/fLG4iW+r1zyDCgRB5MqCS8eRJ7fRJCZcgfbg0eRCF+SHo
mExHceyOmBWK1y3HiVm8iOnWLADYYB5lqxBG0mEs5OQngKbrZMJkSq/wK4x9p2VfWG64epUa2gsx
bYSyVb0vx2v4W4PZPicrdAR0UnpQwP43y+fYnP+0ltOmSnyFO6kldy7oFtJiXNsBDc5Bo9i5kwiS
jKPQ8OywwrZxEVo1Sqe85km92FF+W3+DC1BZLyYKjJDRJy07koF0VxC/2Zw2z54+Vgtzv00sUxDe
DT6i5mPG4qaBBJ1W8B2GQc4mXHWfBeDa8gOTzhc36cPOOvoisxoDSi5Nkt5xSDWK40AypgFDiqSd
JE5CKpIFwwjlcLQ2o2ASApYe0aAT1bYKvcIWQfX/Iyo0XeJHcDRxeTJXH7Iq5CO8Px4P7h5qOFvk
s2f5IRqss2ftw2TInTYeQRej9PogH7pIwCD/B5OnAfqCbOiOCYUtV9ykHNEk19+7n9avZYZfycXL
4OSQLt9GMmsKi6rCKfpZkn4fZAd4jqHJTFvHxVtGO842DSRa48s3y6O5rKUih1FsudnJrWWwusQk
1w0/SNUEEhu9/5ryWbHdzZNfwmFlkQdJ8yIK0TO+hMtbPwhVv3vQk086tj4mzXVsZUh/BtJbxWyN
/ZV9TgWgMlCsP8ppR59Y+3Ql0CM+k3W4gVZhprGbl68NWnq54WgFSvIDAA7eJyUcI9ZnRvhiFYhG
8gBs4gmydshQyAN4fMkS8qENYWhdGUE5C7upKRqeYRLfDgbivFyrEuekIWgzxyHtcMeyR6kyDO7E
PkbPQGKXIrrxEB14Cigx4V8YOEu0B7IMmusFd8ES012vnXk3dGHs5/fJP+jIBgPUNhue6SBQFaB+
7bIwthtR41I2q3esQdCSFTUbODRxMgUTLeVhTIXCo9BPqbjLOYNkqFUjVJqSJBG0e1YUQbKCR/WJ
8IWJuVNqqBtxCQiNjVvWaSIZmYmD5dVn8MIIEJnUygCBSDDkqFrBgJ2mhUoV5kcuruFCpvqXvSVO
dTinAf29HxLJ/3PyCxKvoq1rq0L7U77yPPyuFmQZj2dl7D84LSNTm6vNCb8JqUPZnmJ6MSi1cJWj
3T8Fl0X52yVFCroiN2jite/Bw2Bmwlf5LJwknkfY4LJsT9m+73k2+Lc2S6eeetDYrh1BQh4DN50I
gHk7MAAzuRa02jgxIQ24f3tL5dxIKc92sgHlsKWhT+JzcXb9ne2oyimNqeK7ajoYBqwxYepRkZFa
htgH86/rAqppohLEcRGGrcWwU/SyKKaL+8uku2X+3vXYSqlgN+GAreku92nxtu9wqnx7xUqJerdH
y+soifY7JO9YgL/TvdvYreGuP+lDDwyjUuog1Kge2w3CfHJXZ55eaqhLJpPVx4W9Gk+MP+IedCGC
ZEB8UiUYitC4CllaPIPs1b4v6jQDHwlFI3in1lk8SEM+M2KCxNLQp7uv2q9FAZF9LsIGlxPJRmhG
aPqlFP5TBJsRZTWfgLJfOZKYTFOluNbqZCPlEp+hIjV31DiCNlH/IOj+bHaB1FYFncyN05p19WX8
micw1Uqh2Gd6xPM32/v32DUQSMLdS8SdwqG+R6yyQxd+XbvVkOrhJYU4jL/XXfh7VZRTGB9xRsZa
NK7c1/StwgHrA+SaeQiduRMYIBO+2YM/Qibfd0DzuFaGKNgydq9PiYz43xTyKHCqXHkT6FEoj1zg
/p/l8wZfG1POc15IwOHN02tqGI26P3sE7Ku3qfYsPKpWALufK9w1DR6XAlXtAqjhUsVZBYoxEV+c
a1CQFk1yGVHjm5xXJRG9MtYaPAPJ8jtVuI4KwY2884XH3m0EzOQbZU3gWQgZDCV7JaFFM55EkG3x
bkKoMo2lkZuLS4M9k7wwiY9fQVeuDByhfiap40qOn4lbiSQryMrsMzF9h2s9uMtDeqf9LoN4VcEU
2kkJYsPGN09/SsMR9JqGUTUaAbi0MFZC51XJ7+344ZQqqT3MVj6wr2RcNunHsEAJfJi10K+csWzO
+af6oMo/G71eJ9TfFZMVmygoZI/EXSXE87crj9HuLwAtvLjU/EDgLFh/5LLqHVSZf0zGJbpjrm2s
fJXw3zq1XUyJjSEodee4QYNgqIGle1ZmVofdKiXa/67onthp8dkFTS1w/qWiotDBgAZKVE4uQfiS
ZVLfsApd3WIJY3AkJoPDNzazm1tl/PLvn8AEQDpk88KlNVDWPhvNy9Po/OwWXa0jTnmb0AXUyzMl
nN+OCyVT3yYqvHm7MAoR4dA8T8le9tJkHhe27ieSMOUYuxNroOWcqPNVTvdudxsKJ9qLE6ySU2K7
L81+9eQb6LdrE183ILnhycxHt4Q7x06Zz4KvlkRusyaXLJo72atXWDoU9kjbIHKetcKed1nCeCHy
zo9eGpSEpXF5YT9sstmfZ2G8Naz16fW+LfgwOMnsUugUoLUO7Gx1meSnWRBsC0AbzpJvmblXn+72
aJ0ff3RBe+NUm8RSloYHolDdWD+FQ5NsHi5MDVS/MZvrJ+66cjgHbi5S7lFrR6uB/2aaBGBx782O
+yJ2RXxmjYwAE6CjOY1oiF6Z9OlXUV5AIUWJ35NcmxSolCKgYAYFo6+mzdnqHyCu0iBuMgSCEzMx
pQlIBKVOtsC8NmXeKr2d2XrfWNC2sZgs+7w1ggSMgQGy7SWcgMIIoKpLyswzvibRD93twTyq5GXR
MNmqcdRSBevbmlSYdT2hb/pGufI9E9zvs4+ioWw277Mna8vAZ1pz3i0y0CNo0bB/OMVhEJ6KUrdk
CHnqeFe/ELZNpKYjJgU5Yg56kOXtFwiDxDj26ur6bn6a5PzDKiztZ1BdN1JihDA4IvUn2m7YPIwz
k2jqEP+1Ik435tJkfXrmOa+l5by+5F8VYIRUvdVepPW15uSoHRHR+u2iIPY931tKmQRfbyMVXAHv
VQ5X8vVp6VsAUQeoEssxxTCJV1rg8ZDZhsSI4PDljDIluez4faU1wEqDUVRT1/kMQOiTazm53QMY
RPDGhDAaKx5AZTlaccZgcNFOf4IQxg1/yI4QSFEw9Fk+4JYOAXn2TQU1C6fbuuMBdGmIRGLy8oXO
UiBvtxeH/sh3ngG4CXCdqs6keDhDeejcTRZMgTiYmZzIGJeS9dNDd/xPHDpiIwSa1Nwqaq5E5esm
HXekH0dgNtenmYW7KKzCOPeDEHqzNwZ+GE2Ksx6a+VAr7SYTWGwQuZChKfVUFBX6rs8Ls/inPsxY
DXqlnd2iKv5pjy5tSq0+P4KwKA85MLgw95BUWtRny6wlH9oZv6flpzJcTFVAVDZPIKG8z3tnolfV
//r8oQab0AFjTxJvFoa59xHwzIoJLECiWzVs2WzyYy1+wf6R78eQlyRfFyKOiCLKc4VanTgwd6rh
SIT/UzO6D8Qko60+oDzVeVsxvf5M+DKG34KvPxVpSf0Mux/+VUgEhjg5G0ZP1+KW2zb1xjynSQpI
66d0MjyVU3WlwHw2llBjyVRInaCuOMwJb/xReFt8YvQ0WJU3ycU/9plrFSqjLkWRNC50Nmrq+QG1
mo2leVoRO1AYlNY+3H20RS+i8Gxib7ZGZWToHHBH+TWD1Fe2Hai0vPieyL0PbGZwHwvUcUr9JVFE
j42Jr8ayny33pt5yVmbOAzHz2I/CBPNE9idblbk+CDja65Mb3sY3ee4x/3wRqzrKJBPdPn2cYFEW
Wvit/Ck214Ji/ExEOTjU0gJzukgzCQm0OrRXFRHTxbf5y2P27wSTD+nIno5sbPD6YxU1RW8R/qjs
yPAgzskUAfG7AZOhF9r2QmfrISM9jcdCd/FRxFoGY1/rlLri5f7fOQSDfHNIi+p1oOwu6WZHnajy
EvPCyi7bulJUBt+m4sfMaVxMwmCdjP3G/9ePLDhugAtATjYg7kNt5N5ElRjwwLnFW3xj7SvJfq5b
DE3917Vd2fZSljv9QTGgcwsWLrIdRJ4KYnzuaxSj1jN0LlPLVNd/dhtt862KqBVtLle4/Q4fsGaQ
NviWCaY6EAWq2IK+6EoCzZH403aVEget/r+dxgaKn+27GCGj7i60xsFa55tEmXYcJzUVx8U3ZGd5
UZuSVxvTPKUCWmh5hmlmsxXvGhdgzRLN/mZ1xLW5spJLgi5M3lZJPENyTKmgGEdwtP9i+FmUIPRR
5J3uJLnWzZ2zOTgaIR4kUn5UrmINJqpeJbrPY8XWsZ7svsvZ+GTFDWCKe5RElozGrrmb3GX7e4FC
oHI1T7oHikTrrXNSwg++71A6ciMVBE6RAWK9XS+wzJakObR/1s6Geyd7L6ApZqMPfTcCGTKxguus
H3d4PYeJVrNOU2xIxZRKVE2keeL9jpxALxnTPYea4Qyuiii/cOTUxIotIUtAKSOyaeW7H0HEtdex
gp6jJudMufnXjkkY1k89mKpx7n3W9Urql1SA4BRWYiYNxtqjwUk9IuVgYXhtm9E4gmKngkJzUUAc
bS0NnGmo7YKkXbIzOlVsCMyTp7gwhtZ+wDbS4lauqEvB2dLuAWheZLTLIFPQ68qNhs1lzieHbPgC
Rc5fIIRDQeojmTNzcELRnroM1VwazWtfCPNxT1Uhf/N+2EC+qq8jFRqWjNW7DBu5aP1995lHgwrq
mBL+1ZGCMrYlq6bBXZ/aynge92xRO7OfBTMWbtmDZUxaL4uXu/1fiXTH+CdWMns1TTqTu1ndAgBa
UEE9Ca24ugFRIxeGpvPUm9yjWeDDi6Yr6vOOHC7GHoDRrK9sVB2cwwQFWy1X3opMtTaylAT0HS5M
SXNMLxX0DUMqfg1129dp3SNuLKo9rQ3cUVTKTsqmKvoYdEK3dlWqeNSfgVCsepnVLVDFJxV+4nZk
gHTZps9cauNbnoefa5UQgzOg1ZBgYBOVXhHk31ZtQ02DGyd8yyabqtN9cD5o7jZpgHU3bDzGQtD+
C8sjTvojHTeNMVllolalP4jES8jCNs5wGDdOOrbFZPhF3o1GqI03mDiS+8APEZi7UV9Xw3cpFZLR
/LJVOQKRxeRU6ypXDezJeF7QL5Q9EoMmQA2KMHzzyWGAeNIyT94OOo32K3+w4Yz7JVL0JMoLNPU8
3Lg3u/+RK0HzxMgQxsAXPii2LmrkYM//ZKkzF2LteFKD/PdZKFTjz9AhEMZtWE/SVy8M8jxtk6Uq
LjyZPSKwSI2Kw0NkeOoJFeH/W94Wr3xcuplab39VO7itxiBuDaQYZ0kU3+ET044Six1GgfM/6Vhl
Ea+NxV2iWazoPQiMFwBtLwvbefF16DRekWkpRC0cHGk6OiNuAUYwSOX1P49Swg5O3yoLTXrxBwBH
ov6E5vNPDnFLKhH89y8Uo5Rg7BwofbpbWU7yCge6AwHu6Q6aYr/A+UndAi5DQ3AWCDcLESGHZsqO
yJ2vTg2ZiOj0mojNi66o3RZYiJKquREJTKElFAEG0S//USDsaqnK1sDgjejwZDLzwN+IrnO3l2Ir
GPbxOTXEZThhTw+JNUa4cTWxUotfLJVMFEc+I2lPNdrJaRFGZYYnnnVRbBgGwSxy59b7WrJBoeqe
AdjZrDZ+GVJ0GlXnJpXGBn3rWTY/rrnMEFp/TaPhR031Xo3KU55wv+/PfZYLID7zjFcU7YfxiGXY
TklWGAAKJ+kNloHzNBd8O6SszmWNeX5KTNFB5vRnr+m7Of/TIcE85MqpWOZ9ReGeX4ELO4FGUEhA
6OgTJ9qqh2ZyC75PVcdKtJ88JgQbFm6mI/Gsf3piUiVRsSs9PKl/n5i6k5Wq4aC+eWvnG3K6WPyC
ZOTlEFiA8cU3jQeeVifekSK/hBzhBqvclfY/a91Qdo+ar9/ljzT7EiazPXBLr5S661QMxZtOb2ob
kqjtPgUKYlFPpBDwi2Vs2iAtUKvDfBDu088n3vHaAUZkCLBDifUMmZfZNOqE2PUDkt5Hs9Cdqp27
4tqL0axA96R4//O2o56l0Zzvy+3ZEQsZ7uEj/ELv631op5F2tT0SOt7IeUpCAVZi+PTZTc5G4FJO
38xB7NWNP7HTldrdU4xiOl3qKAcr52vZCPiR3C+OkRD5X9xgqG08bTNq8uP7fbixVrAEwVkZKsTM
bqkwzSinlkPZfqaissKQFdqYs0L9B9U8fnL3c42PG8mlJQ+bi2asdR+/cMyJ2z6pCNR2jxTEOkn0
xb9XtyfgUfXi1qfmbWVyee8YHTrYIedxY1t24zkmxLbRfs9CJcml+nq9NPVq/w3rMaM1UJ54gHMi
trnou8J31EV0MQSeKJSuSvxJwYCpnSKzP9qNX1hu8Da7EimifclR4TpgT/VteCgk06bmEDT8qqA0
n/gOkFK0goxsKhtj37yzyhNMpqo7pOwE7uDMXV5rs7hrf6Y2ITbrb6l8uCy2T0z2Ykz9HHMybwJ0
wYe+mMat0jxLDbJ+MDMC5p+hR5TauBY/vdYI9QPPBb30jG5w86IhAoMAkOIR5+irjhd33uJlJlzU
VesNvJZC7iBorKKUHgSbQ7j+rH6rr79gkfUfdp7XZgc6Yu5Dz8ySv97nPFszCYEiNhG4VxJe5Cq3
QVk/yd+Wdq1vOgL8C4TeF3UG0s6ljdU9pD1z8r5wEEBGn4eyc7zUnwsjmbWSSyOXOofPAOlryTMU
dRSAXNgZDAWvG+L1gV+0OnPqgsnlGENWT/MWuR0UApTDtwhAWmYfG/C/UcTk+H6DysZ2BUvImXqj
+CT1uFkqSC55Jw7Wp5BNIN8ayi6B2DBwI3wf9c2bOLTFP/yf0sX3mO/sjBDsfrJK51mTSu7eFBzV
6xJf0uOw/GOFC+xngCjFLFafBE6KHgSG5w34bHjUIxE8B+JZ8Fyrmxq6Xe5NcTJpvs5qE5ir+xYC
sLS5GfZo55jZ+IAhOOte5+74vioH54ns9ZqkdAj5Ko6HOJWpDtDX/xAysBvgUIgVU3DPqIKDTTg+
+cqe11nUrOt2Gv7lbSOBALN4+5zQb9ljlcZvztCmSZHfrihi+gqjfrag5CsxmuvKtzPGfBNayj8S
oxgH+Xy9yBYZEWE26qc31567j6vNlw40T1RZQ5PfgP5O4O1L46GSgtw2wwbtDOE4b7zVYWKNmfNs
pI/NiSp5KJkIugy/7irxe5399vnrctMICBF7v2dRToujTZDVWZFAToFplgWFq/J2Ir5eUD9W8y3L
s1aApwgJ6FWU9SyCtHwl7r7etGaIpPzWVR6jLBKr32ugGy2LXZ55cVb9GVg2sylFK+c3E7hd0vks
I1un9KwPvTKQGujVL+3OUGcRMbRQIQ+MsuO6ClRMP3siBUcuh17IbXFX6zf5FSqTapctXSRJ60I1
bCh1/bLij438ywRGo47ob1L7vtycX7meOIrMtXdMaSQ6TG/9Ux040RLNTeSYGk57FfV0nbyraFvC
Te2vv9QQOt1RMbgEBVznCAALVQLl16yVR9WItuW7EbeWBJgJ4JNMBjHwxqsuLcpBPSWSi8LNUK7L
jtXdgAX49T/9PB4taKakQ1RlzWTovSnMv/6Mn0OgCWLaBeiPxZcjCMRpvPsnPPXeEl+xJJczwhaU
1nBFbaqHMqKsW7OCjlsK8wBNSWyS708flrsSbVonNrGsHAxi2sE+Pogq1kiJqu3IVjQIU9TBvvKf
qHmfEMLvAH55vHdttATj7LJiiVz2e/j3yYRYck6DxLu35dkLV2Mpvf28JqkjFaXCz7U+ZiUu0aWP
ogRvexUhvfCGFiOCr6H7Ie5L+q1Q57MJW5Mvgzp0fGaODvE2b6TEEkR/bank2YUj1DxlSSbHd3Jw
Jmgp7pMoT/PZHAoNW1tTDIeH6kApAPe0bWX+JklI/lCxSEJHurhIZBNQZ8c9JbHifF9j1OSLKlfD
i1GxoRDd3yr6PwHpGnvoTBPiGx006lh7mecTQhXCj5WJ4u3mZZTDjgS5hx4CIxz4uN5xVVBOErSz
gyetLOKdQjEM2r7BhUi5+ajt8D/gw0ido18lQifonDrsPG0Wf3H/MWcig4wHDE1wIbfilnOpOyjd
oGL8KP9FZd8WpLoUbwwy1+NYNzJmPlkAI2ZhGlLPsGY3T54fuJj6ewilK3c2Z8bw9POE/kiIpyuJ
ysbVJO8JuExy7zZ7/gaLlttZPduQRE/Ny2ET5ARPiquoy8wnsmhbE4qqs9xkVFBKXPRvgGXsk7AP
nndaZE3cHzhnU7a80ZUJlBj0Aa60MxP5efBjJPRx/FTxPHP3ipo8Py3VCVW0MoiKDjlkqc7s1wcr
jgpV6HAHpW1E+eK+8TjDlO/9XZm7wJL9Rjzq04NW+1j2ibK9MEs5gRJeo962UsDoRoGVQ0KyNaX/
S651pJBKZwEf3zLZ0lB/zfyYVa0JSfSfXoY6FXVBTI+A7PUM9NRY0vUaK4cG2KokMH4eX4GpFCvf
9zTQ6G9TtwYVqE/BYsp6qUvXZ0eD9GgdPULeZqzDzCL9ZIMl/dJkDhzVFj6K1tXYqVZ6b5I6HCGA
quPqX/uYowayHS65Ou10PQumneFhZJnYP4+UmTstq+HZhLPLsIlNRQ4ZZiWjojVCUsCFI4EDO04a
EDgFF1n/dmRnFl3/8LNFIUbZc3IF6bboC0cnxWp8eLFVeUPvaBBS6nxeMXdsv1N7PJ7Y5BaRTWGn
yOOlUd3HKbLWB2kXnOhP4RTRLZV8e/PB4BfbgG2Ant/M1sbxFJ4eVkltSD+7GQ+SQaCPGHJSXEH4
t2CMLwE1QWR435R9AxyWp3zA10EwsZSVN/AjYCX0P+vKvRTRuHHXjC60UZPcA7pPfgtkIaWtxSvc
MG4Y0+UE3VMnPeFhZRDImN8+9UChNgdbSBArps3Ci6y61lcqmHwXs2pLWEg2yJMwExWX10P0vhLF
4eJHMqVSA2GSH3Q27Xx3XfNsZz6dUfOYyK1mI58KtGnCOuKZUjvzYVx8aBgGnPAqrhk/EQzjdZn2
zjYTExYzfYEEnj69li1x0uIUZ/vBa/uZLMvhH0smoOkeyLvnHMmw/TzaNib0j8XyPFB1OMdgOJu2
WBCR59qPcWa4zA5e27kzrlTQgsho5CuBT7qx+S/EpCtC9T3XD1ys1KxUA8WPHzgDKbtq9Jmlx3XS
nJEcY68d1h6CH1n1a77SGLoLufSOgQfjrhtY0bb2SRUD+pCZesN/X5Kk5Wp9paK3IZjY5luf/rK/
eAw5Xm5o7+rES/MaXtfSZepVBSz2Fmk0PkJGHF505M0I4zmYpL/iNm5JrWEmRZuM3eGvPISyvA+H
eVZy+lqlLXFlZEn060qug0SDM7kLsZwpqCPH0ssdVocyYnm4txSxo4KoWf47AF/LrYWS75PMcf8g
rkhUGbLfLWhUV2t5+R1/Dx3plXZburQ+oukC2JAuITgpxQqo2nzfZj2O6XMi7OKOEeF5j1WvtWTh
gflebhzWejQdh8Qy31D+hfS07wcpKPHEyc3tarTfHUQ0g1XXuQD+DJQoaJkNs076nMiiSqJT8mgP
929LR/G0tWAmxm+NkCftsgEJtxhuk8AX1XkJi360ewbrYVgaDNTUlX8OCHk3OGyozqKBe7erRDUU
2Y9UdH85mp4tc9Uxqqv9P7HX+c6YkP/iL5Lthj4z66CXKPny5NaSaSpEDChEc6Gf7Wns6ZDqcDaf
HU3mWy3yqBhsGRvSlympM/Y76N6AvWfSUG+rrN3qv8IEkgqC8NmvPhrObgriwa8rtEHIp5RgHsr3
l/4kcDOo8S219W1AAuoDSJhmHQgGCCFVieq8FWyZbtazjsAR0F3HDI63ebslMdASE7qLY/faXiL1
2oGjpl9lHBxKn1FRGX+bR4dw1T5wSbf134O+l2dbcV0hnzuj2DzqcGBjKYHBd9wA4FPwFDpOmbU0
lycxhhDlr2k+2bm/PVZFFvGXt0+8QMZczL7B/fcPdvMfu7GU7SZnXpSG6HXSENu+BZ1vFHjVZhRm
Tm3fSQ/BLpJTT3I6mcw4W3j7cTYLvbThH7+uUmMQF99D/3Mq3kkP4LNqfo/bbCVeKLZbB86dqsXX
L85ki+7TBaTqW7OEPvjTatxP+FdiqGiKZ8zbpQk4bymKneVpStgDC/f72OMXAb1Fg3BBrHU6ZNRC
aoHhJaS2t5MmP3JBAj3z1ctl2EyKDLtZIwNx0GyEulAi235Iy3ByH0ZIc1hnzhyLkOfjWHkIZeCt
zRIyWf4tUryrqznxik1G2cH5dGqlR2Gc4ELbl3ce2GBAHXJ2hO5uLXafiVFIX9bkcn1CTn8+nNiX
zv3hiDp66gwuEzcRgYUNiP6mmA4HT4c6aIpiC8/t+I186k8UPu63bLmwmnbtZZf4QhCtaHeMif/R
6OVClmr2chxLVSioNBBFTkVGgpXRnx34QDsuNhYELMoal3msnIz5PEMkYGae4pxCM21jWkp1/63J
Rej25Ywj+1rLdMsLqEDIBR5iFtN++ArdEV0Y+BHvAN7eln3s7NdAHsCRv2LraKwFd9V2IfVsRnCX
2ewk4+NtPbJJpsNi+3vhk7wfpFe22EtA1D16IYRJFI6J2z/7hTMXbeCc1jBcEAy5uZyziGAy/zOQ
yoBpk8QLAizMzYwpi/ccWnJiPHtPLSs/cpFKvroJnqm2jLUgJoRFfHchGJAqgamWMRTL/YF/JaaV
SZmM8OKXgeNAkaeGLrSwF2OrLpKXrFxcRflTrUl7fbEveN0GGW0ph6AWtf0u9Y+nRfj/yTBWDfEY
kHnV81QQAhyatFsBOF+XnS2HGdWyf2i5/2OqE+lXeXiVAIydjczTgSi3odjlq/Izx1KLIqcTZWM3
JRZprRNpkhl2ACgCvaJ6hcr11BIYcdyh4wc8l/o409vC0wrZCEM9BUihUotTtJtTavL7b35GOCsK
nanky2m9RI2mMprFjpT5P+T0jCZAbCqe/l8UsdSWz6kkyisgnQKWj4Kv6JR91CxY05SHBd148r2t
h1XUDxmFFYtZR0RXZQPi3CWKg0MvDL/9+JqYm2zgVqcKTRqYrgDqi0plNsZ4GQOXHYBp0pq08rke
1oBMVScEARrIsA4+iPZiVaelJmYlG29wTyvGUsYXnPI7heL+ns/DG7lfziSR+q+AWJg1jknHIeXb
7wJdTizrJuLxodoObvzTniW9iDq5wiYAFv8CdIIBhM83Y7m7f5Z4qr4KwWmiZ2hjlvm+aIVUYP4b
lZG4BxbQ0kGn90y3woikzoerjTzwinj40z61LpEU8PCN+Qn5i50pV3fLo2KfM1zjGJJ2sprWvbLz
pnMl7AzydFFCTZ5FtgnW8QZzSCd10pvgD4ICyPoAfMLZVw/vc67GLuMs7mN+DR+QGyOs4F3f1VH4
/vQGnaBmeCwswCveau8ETjdWYYCXT7vV9HljK/lA4eKaqFiR189+fbxyy849mPs3ZHjiMHOUezVi
+FYbhE9O/J4MRRkdKFIz9jzdY1jIQ1urwSrAtAV+5H6uKMOy75hATlBct0oANWdDF5phKSgJQ6y1
g5Qqm6+EPYg8Unr+P3b7II+GIHueV07JMckqbB2P1VI8EBUSP6S3CDry50iU92mYhVRHUaq2d6uk
0AYBtCT4VBPinfWALsUtExKBohVC0IFHa7QGzQtswQK11dQ2GBc/9M9EY+Jt+3IoS1rNWu0KobTM
xsTtn4LamIC5Vuv7qHDUEe+zqHy1Mp/dgSKEfP5QLFTyhV2PW7lNMNNZvA60YtDiNspK4ht9dup/
NqcdZDpv09aZp6TA+PA3NItGClclBQv+/MtXaart3a34TTRYR6BrN49BsBpy8ZuCnKMJ//IACj3G
+HNy+QqEY6W6llJIFbKrVX2XyIRsKCKjJ7UEiPH9lBtb511v1qAs72zr+bbfOGx/AdmJLl1aaaKa
YOO/ZIA17nuLu4qPTzJIO2V5Vh3SLLXYCNGE1GdK7G/tTslmXJc49K6yZjvxYM7zolC/DEkDPWnk
ipirloJv21Y2x4OcETscYfkpmHI6BrF6tcveibvZ/90xYAOVTqvGPPjyaSxeSqjYxGJ/T1LD1iYL
AGBwliRPA4fpbmp0q7pX/G+75PEzyBLfBqx3N6GtJclFM5nh9wmhT4SEdYncPbrZ4Ebt+bbmniop
T6+cy5MtQJDQR8eNoc++msk2EuneSXa1bK1agpmHj/10kJ2whuNIcCmGjtTbblapV7b0Pomi96g2
KKWCujnSWSwgpN8LwWtMuzUAUCeQRRzVgHJ7xALkQXZdwxiaM+GaAuT4aShnDDApRtigu5V1y5lB
/pz4UCmX+J/ro1LJ6GsgDg1FsXrI8KqINxrMbfYrWWlbw5LsA6Lj9GtPZUGsbP+vT4Z3tqpbuya5
4TyDi4PUpvfKps7SNxNZI7bqoyB2D8TwYJRPIWrmhrzYQjZjm9QzZ9fLf/tNLDMwKzCX4bZtH4nF
eoDmFicXt8ZBPh7InfXhi4Kivlf8rm1pDvGABUyZYLil3yyfgypEIVWOr6RlvokTG2OByUvKatjg
iv+zuitVMMcwCnhlx4mHPNqf10wszFEuom9AYA/oO3FpnsMPtP+eNTKLiLoru3DNJFVZJDS1AIGl
fRKnUjAilQv6eNB7DsLeOTF/ONcTXGfTzi3V/G2dH/aJbHqe9RXoUACdKXFOKbh71c/CrMCYnRrw
pMyldkW3WnP3EkOMRfsrW5VHDmtUm27W6Mo6e/xHCHRZHR3m/smDnnMDdno8ph8UkiWpyPCybTqm
8hCU/1EycIJdbaLMGmofPFBxLLskMawGXNIysehkgEmlGHOrkjAFRRbd4AeATWsYPIWSFCL0X2zp
yyIIMmY+J23O56t48MLQd9tQUfBL9/bNLzEjG1FuB9pDGH5gAYJ4V0bkDodCmLoM4Izgql5gpJFc
IHA8vIUOiyvhPp7ot/tQbMLpX97jmqVwFRTa4pW/pvvyH24Vody0kMnQaXre1/Z5xrDk/xkmjb5V
1L+JxOwVa+zp5J+4pDb1b5nTTmCpkVwFf0c7B75Ff4nbG6q2CSvMZvY6eENQTLrxTt214qqjaNPZ
sr+8R5cgO3P3uZ39PcZzEkDjaS5xvp80lU2mzz6fnqLaA5STZe5RYtGPRDvZF3mcfBE0OsBxXtcW
5V9dHyDyh+Dfceft1LVllQpUcPFPaOBgU0kLUEjKUq+eXITNBP73vNB2ToG61HKpIkMlCLMpNKob
NUt97qF4W+DCFJSRHt+00yKoIqQhG5ktMzzvGv4H7gfnF29ZY9j6ASjiArk09F+ite88DVo3uyrn
mRDWkh+br0m4bIzy8yIY44h/fZPzJsx3zwdp3F66XAC3xQgWrRTHxxuDS+1mQSegVKzaMy0opw24
o5do3U+9kISiGgMK6Cv/CPz5MZRJWDr1wy03ym7QqPZBMd3GlV5GLla69Gc12FF74viyp2ypp9Tc
RI7cu4RJZHZ/tMuhwu04sbEdAIB1K8hr9JVUNrShyxhFDpDtsRN5yvRnizMqy5xxHff4bPRCcoM0
nWHnU7c+FtZMSmNEhb1WxlLvyjvV8g905epjpXihTo1lSlCQSkxS4BOHAd/ZDxG8fgduSKvr/l7S
/z0a61ytuZ5t4YrjqBChU3uyTi0YbPDePIM2o3WyPX8LfZqLW4lsosn0NWLSsDUGUDuK3f3xkDgZ
6lACCeJSNtktBRjgjMQbCKGU3vX1f+rEvw3c58ysBsVjHTiCGhJoTcSTuzc3Jm7oPSjKCO4zBk6k
Ko8nCyFYj/6ls2y/I1VRT64AAahbJU7F6m8LYaCNBvThndEG+tzks+WubRSL7/WO6CXtDPq0wWjG
49MX1GlV3DbRwNgbpJKh4vnckADDVFq7TAFlbU8OUlHF5EQJXZUSnUm8orcnRJvscHK06XgshSsP
XN4Z8y642VTIDfa8SS00hslRuoMbtb/x32D+D7OHlw/r3lgwYjIZTmHyYkzmeTNx61x8QfdNXjEe
ASla9S2o8ZNTFGIbCpp8dkSn3raE0GCOVQiTOj1o5Nh3xju2xnZn91ilFjrtfwpMPOIpEOcEZ/ge
LtsUZmtZ2fhp5TW0J0iC/K3by/9EQ1dZyXLzFDopUG5gEUY03G/uIwMxwrkLor3ejZ9pYbP8fhFR
wHVhgFEIULLOSxu6CPjIKmg3C0nEeWXJ475dJ6jFvkRyomxZHHnZUD7QadF3rR0eGvpj/UtRVFFv
/iCFyH2t6o3YzurT6ONuksEhVdCZJ/vA4VrrRCPxQ+jE4YgssZRevA9A7/VtIdR+DeKF7Gd7s5Je
/HvYIJXOZ05RaBhtS9xexe7IGIwfepFRRFOndOpLxpNLxvUIqIq7xqhyuJx/in7pTIi5xjbRgg0l
M0Er8J0fQuOxQE9jQllg7JJMTXVBWYGhouXVWm1W5M/XXQvdpxruaI8Mg+OIpT7Ijx4FYLUsmv2Q
3T2LEpaqcg6pRa8+VMYA3vqxwunZyMnrMwBzL3F6H0opsFn9vJIagQyVbnF/Ny3APhH7ehx2wuHa
UMNrCokVhdlj8Pv02zo6XZZLx6V1P2fWrz/awcpKWxOXm9rd3DzFStj/sX1PKOK/AfAVtE7s9vci
GNxx6P/tsFQ8ReNsl3QrMKKXR5IwpLfLh5UV7eboNedjvQZeOeL60rcuLffGyo7gTYYgPaw7UsXi
89PfI01RdGcAFm2NGizVL7sFLpAk+luBzEda5GXMEqY4PIdvAo7YT+miFg1QLxWbSz/OHziilDhs
qadmHKpCX3EWr/wcb6fTyRuKX7Gxpd3bNZy9quum8LMtL3ofg9Q19Gwdp9SAOFWLTIg62J4hMmIS
kV7znmgeq4+5HkElm23r0vRzH4XrV/AUnqNe9yClRvgQeE6sc2AeQz0l1zJBRuP2Avpg+WUuEErb
ZwdWhCTsWlGq245oJWIrxSv7JvYQXou+mATKZ+G0Lg6PAN4/yVnQe5vvyjWYqasRK/6X6RYfQtou
p5GwCHWaZWpPDKpPoB0CyLJUJGBbJiVsQtvqPB6sAUQew1K8h+eLDtQKYHpdwYHV1VdT0qpX3LLW
bDvPM3/2RNUrnHAzqhgBCxT6z5bgQmOX6ExmfTGFVTUU+BSemE8hW/JSRFEv4f92IycXxpokeutK
MxfcwLNc3OeoXMFtXd9n4IY7M7XjsQnpT27nOT0nbeGPnsAA6F/7qtXDv8+lUM9EfMBk7wVWSeUZ
jaejWwz8AdH0UaeO/b8jOjb+akwcrmAVjsWTnidrm9C79mezShdxMhhPIvvuQImCPrQkVDmaf4rB
0b3FOgg3g2NM16qkbT3+4jbILTMwvoDMAYgVVe7HJ4W2Qh6edAUcIdJEvG4ERvLPerWwmH+K6EgJ
/DmLKIq1HTihD2JnWbJwjSb76M7Xdr8pKUcO1FVOfi8RGDelllEbeBPpRenJ3YIs1R2VbYT4g5XJ
J3/UsEOrRLwXVnPklpVv2yRHZJeVXopnsiirDvf8aeMsZOnjUOoHMEJAGg2TOyZgiMc3R8/iewuK
rN3D7DwuJ1cr7SDfvUf+wiaOyG+VE532u2qQtRcsMtc4TNEBzRwVtc/xYKi37pybkabckDFlgock
rF/L+Y9tg5VV99bHY3s3k6JhIew4yQgMiIxs2u9PtD8tmyfinQ7I1HaAMJ1b/8FUJCPPrPv4Uynj
uwB4CJGqsr1dbT1H/lWVX8/C0uHJOVOoQ2fFVh0xa/U5PdnEKMESTZXaz39yj07JEr94QXRNvdo3
bVAAF2XQrzhJYYj01/lwv+DYeN8KoAF8jzzqq6G3Kxnxo0jupCd5gWFFpvH+GVNbZibEBDLCDDNK
eIqPcga6os8E62ZPMk1kCKwsz1/KNBWCzv+SZKjlvVS4bCPbQUeuyGSZLG5Wkrf/6s6EFBHvJpg+
qBobHiQiD8Cdqkts24jWK1dbQ8a8ixrM7eKcZs28V42yZ51MQCXiW0qn8XDuwEEWNMrf2MeY0X8v
xDNcK8O+wk+GEdzBlcmFinJj33475ScLv1AYmc/fT+TNHM6W35neb9QoVTuw3xFq16hmHTRWDrvX
VTMox0G3VZfqqa5Fu2zt4wZ5p6fTYEKawdg3RgbyNSb03BTrsFYHJn2vINjzWeURx/mUy3k+sebe
DyUUwDz643aRn5EtGvYa8Iou4MKqG13CCC/Zr8WgGn47qwkTZc5uSA4XAvm15F3i4mzNrFkED09g
pb+lkXMzAKdNTHjddKYZqD4+KK01fq/K+r3CHcys/U8qpRkK0nx7IRQi8wtG7qfPgrN0jrh3lyZF
ouskDmvz1665FPnYqI7cX9UunY/ZtGGnEge0hExWJaiV1xZnBWR6ZBPzKvxxhrWn+MYFuU+GSDcB
nftCBjPrNE/wp2pRPzBbF0avffFTEHFf8ynS6Y+FpU+ovbYNZkgTanSPnSP6bSEi3TYzn1Lsq8OG
d/ze8Km0pPMYHKT5mHeRKBXzSpxEzU51N1IxCgDsJE4qoMUX+xjtHNBvfddpe1UKD5vSp9a/RabN
WcxN1N33Y3zj8p6jzO/Mu4lXC6PyPkneGmTwNjPuBnD+14so+v5H2Tijaqg0XCRARSUiPo3sGZ4P
Bet9lt1ubvt1iYnX5Qc33qcVvt3fhVoTGhi/oDnIPJk6BqCzeHl4urqWDHD3qmjwN0Z5JZ/Q4x6G
FmyWXRl2YEfNxMoA6He3o9DGYKxei2eKrugXy8V2tGJtyyS1RUNnEflW1hr0ekmxDVG8wlTME9ez
64xSi8EnbQ273+asRze8Azn1KlqUV1hI3uBQtM79oEnrs+/cSIEZBRrMJaHApfBGDSr4Bay8tRGS
G2AFbxTGtrHk3BMn2jFdlkpXFktk45buMZl/jRF+bStUraRFiE52Yh7irOaBAIKEQLhJD4u44JGI
iJRfDPwGw3HMOUDMMIztOhAngtfsQY/Cu83JKnYdEAnBuwxndaGSNMqXtJOl0U7HJM2PDE3nbMkc
VUuyVb0RPOGOY14KMiL3X2dCBD3925nAadMOohZ+EMHhXzWTMZNIv6pYiVmSbd7hX2EB9vELyKpl
oY/MwRRsoDPk+r92u3QtJVsJ2TcBXw6EJJ4JlL2LFcTllO9C+bASdr+ZOhRwV6RQX+ccGMSg/V0q
VY0FHi0Pv+I/4T2trI7hFv+0NgTufvJwufgrzSGM9yOkfeKMCiTqBN2CQvxoW+oZMWNu6gYkQDh4
CSn4PTCrxAYb00uwlwdDYBIbFTH3nbT4txFox/fHugtMBuYv0W7UQ09UPIj5tYfYUYcRgZ+m1hEw
eqW9PP6PZO98Bvob5mviBiUIru676Lu6zC57QOIMXJAqquLAMkRM36lcOUodRzmSjBsgrpnmJ/An
PTSu7wymegWa7ml3Yai3A0xr7lg1UaNNlzq+uq80UEn0vNMjuq0Ua+k38Ib1mBrK+NO0SMELD+oH
Fzn2QeGkjgONHvMhbvhpZYEKrlMiY5mPICY20FqzuOiOX0+XFNYjQZ9a/10MFKHzBb0SJUWlwOof
8nQ26/7aiZJZxsgxwm0UZBX6l/whJDCMZgvuq2imWwVBTy5GLw6cZ9GKlJzJJF89ClnZ7+S1sFva
KftsDCcAzjd9CqIvA7vnhEpnSJIym3rIWm+ldEt5XsiHdaDHCec9SI0yEyry0TKG/qxpbWdnrfwB
rxpeZhGAB9i66BcocuzTLW07xeqjMFzAbHn/2RPDFgkpH68lFt9xY9t0bRaSN0vgAozFNHUI5iyT
EtF7nkURUqR3/4aD7qkV5RV5hFCDmKUCbELuwxMdVUZnBjR9l7Jwq26G93VgkqW+s+DR08Z7QsmH
hh7myNbTGEdM5lMh0eaqzwyWv65KBZempRyc15Abt+ipGGUsGxQrtoT/OIC1JpD2IaCkT2m5eaYO
kuf9+fer6eWreahPsqV+li/AYGB/Z9QF+CnXI0AZsdSV+h/8twkMRGMmzv8aZhfhkvcVu8yR9n2o
QITgocbR76w1lLTHqNH3ktCEDyv5ujaEQyPMfvxxpp0Ou+p7M3V7H5c/E+EaH6U4/0TB8W6AoU3M
MiARp6MYH61G7K7PeiGibCVkEnC4lpPRxJlmnvtTQTk0uuvd8W3Z6S7TzSsv5kpTCvMs5eU4MZDM
gp1WL+LkTwAz9kGASvzW9pNxXkmnmLylA4DuELvUcMJgpa0rzAh5ubGYEFnDRMVw+5yb2hs3YnJ2
Nyhsf49zem2LMWQD0fDYenYNpwKRMldQOfRrACTo3EyZJzKkSmx3rKFCaCSbI87y+vXEB9hOmpRs
+1fRaVTwk/J0cI0uuGRDIM0K1aGz4fjwXoNrIFVZCSqWsfFQc7nM7n1BWXJ/yBdOMjYdbm0Pch78
MuiGBaM/LcjEL7TyGNW1W8RCOR8hrxeIvm2c6wjEjwlPLZiKLUGuwAgyXNY1lAdgrrI+Qo59PAmi
N8X0B2SnJU9DIvCTkY7EUtW3wk8h1fQ4CLFy1oKoIaRqv/pRqNw/UvgBu3YYNIKtOyGI92eH7yJf
FamjUSihn2maZWnpDeiZ1e4IzGu5oVMKBkeIoRr+I21BvJosi7TsQVlYXSJUM672oIW8+FcnGDkZ
cu/+Dg0PR1cv81ldwc7IckkypPOx/N487tb+c36IsurB6pFsN1e9gva+PHP9hQbh3JLlfu3JvGN5
9ETuMiFqRcsGYYdlq1nuRObFchGZBP2CtcEFHANlpgjCoEIhxbcMgP2pFWn+Xnw4KIL7QFx6jYzu
mDDB/HJGHw94jiSysIKBW1uhIxe697LTKKRyOgU/HFcgTjQHMGPKKndTMHGeuk4JCZ66n+0o0V2d
qpYK92/pDYA5iJdJCtbe1MRwEDRfSqsT0ivPjnx/4uEJRpxEU9EnXnSwSl1aQFzCvXBy6h1Z9WQc
WokHRPKg7c/6koE0D9JgRYCrzS0Rp2deRtxQQYcpzdNgBMSolPRqDUzktFS+p7qrRHXI35qExWm7
rVt9yHVQPDWqKC6izZGycT/AM6gp1jYGRyZYH6ow4q9gHKfSLUdNMKZdR2NOehUPHu+hICZWeTM9
wj2aNEAtrOuXezu03kN9x6oMiA+Ux2b3LeJ5rFZpz7PNm1H+wT4fE4w9v0G8TcuWA8WBV0de6OAp
1WxTR2PwYndpgW6lJjkMtkmYK9SlH2oSuZuRtuBHDDmzzE9ebduY5W4cn1J9Bh4DoLbu2aptMS0c
QwYzFOvrGoTR+N/JtjV4zTTQwE1SLCtvYjldXb6Jup1QaAAAr4IWtfezV1tu991S12McAFwAvm49
FzaTUvrRLtMK26/+3MPXMdgRBMQHjJrMFrCaqzEbrE4/vVnwsmNR3XxDG/yOFLWvDIA6YWZ76xgK
FJ9ZWt7+D5xohtgqZc2T5KaGOUENmvzn6+I5TKkgXMp79JOMw6WQZ7pHHebIozJqlI2PMIcabbcg
j0NVSSM0iQLxUvn2HVv2YcMGNu2XrMMqYRpnPJWWhUz4H5aVbvp2LX2pRupDcwmeb4pWftiCK2KC
9ABVLaYlfdzaOfIRi+vWMkB1kqNoFhCka3tgIDPtVKNkg1M0GYIH9qhalk1Yklko+7btb/DF0GNn
wN1tfALPv0uxL908mJFo1GCraXjdHcF9ncPSDtB/wT+RtRMq6OGGRnq4sqKheK9vUAl2g7dAdotS
4oFWKNDY15lk+jcxVr0PnVGu/dxUurg5z70cwsoXl03m7p9FM1IjuaZYfnMoVnwrUuwQOGhypAk3
h97iSL/gBusZ8nWQtOeV+5C9ZPqvLpERWIX/xVUAYCFRT5I88k6UEyE7xrheqbehSD3QcKhoYiQd
+QXblqTFQBU5sIOb2vff0tPBDqgSt8sv01JESA0ZKfYwGBBSUaPMIaQgL3aX6yfzfuqfG92jEqoD
6hr6hlNcIITGRPtxCAc6jqVFL9q0Ocv2jDm7eMeqtV1lQLr4kjIwjs/4dACewtFM49UvjWB6ndv/
G/WlLG6+RQLGyGAoABRAiaQ1PwKe5YC9BkqQCkiVIAM/9QKleZCCSbVPouLc/asKN0clH8SNm6UZ
PG58PlLNu4j8+5Xtray3q5VhjmSkf3DYd2WToZW5kIX+UEWKFiyLiYO+ZNBhhE0pez5hrbowBsKw
WBMlh7Tdc2HM6+a/0E1fWNUGsph62iEXkklCMOK/ZGI3KjgujhAOY3VxoLLUDxQAHQEdISAnjO3E
72t2ZNZkwZjKGcfthuEedkuoWMI6Bc2UEcwkgOvkf7dj6vo2hc9px++Sxc6YgOtp3A6u7aLFvxm9
OSeaQwhl/YNFu2kAY+pKvmknnDZI9j/xHYnWZWobjRdT9f7bTewh993h57aCpDw1YU+TTCj9sxjU
pVV7nX+xWHi1lRLk8BtGkwi8gGj/UL/iB07lwqOis5B6lLzAlZUJh7gdmu8emonyHRSyMZggXk8A
Gma21QVzqTtk2vQAyJs9qGVf+qNRR/4wpHFZtILzu1VUYEEVmrU/2wbj5LsGW+vKgNf4970M7QXj
lzGJ6QChp/EyQtnPaxv3Oeuc7M8ab7cbgLJZ8WayVVHYcZJ+SHINUOu1uRzazdJweg8G4jJoE1gA
ZRi17W66QzDVcOcL/GrU4pAAGAt10tAIXE/8m+tVvT7j5ra/agHubrqIFytJLA64nWZCFJF0olAF
0Fl2aYFGymJGBxkpQvB36bFCL9KoVaoDsPRSiL/4hZdwSYdtdXEe+EhNfxycW4f+DUakOxVYJ0ks
mDY5O11HF/n0ENfwfpEAhjrlvOvp0iHqV29y5AuXwrRXOnJpuXXFgKuZjsxwXWwY05eajj7EpHja
mBG125ekwYfADxRHSUruSVdRd5CsNdHvZ+DNKiO370Td5m+XrsJDCfrqnSW1U6l5o4fDlKwosCQ8
65D5lopcTEkGqD5lB12feQHhENtKAG/vaqvDOyluZcdr1JaNH7QdU/jvpA8INudMKYbdDUJG8hIa
suLh7DCsgQSL0E6TZQ/TRqsWn+DB7NLeFGBEk96MUXLR7O7hhmU0XSobgE8CbTA6dTiJ44vQjkDa
G1QhxS8xpxoP4OC8lsQZGrvclCJSoTrP9iwD1jdt3yCKrmQ5gIn6ZxQZqmrbJ+2kpYCCX2nP9jMe
+fkzAWFYZxCcC076PZWJBAtiYz0QxC0TtiT2xs9iRbyDWgjqFSLcQqfFZutgo805DmEu2ttJsq1i
+oq4+4KpG0nik1Rh1Y6e1LswAqVhTgMGaKBc660BcFryTKE8mc1VZdsLTIwxj6JSIFpNcCRz9uYb
N/TrXHsg06ThJqbBi63hk4KxJ/59VDz5ZlIQlPlASQkqqoTE6jgHm1ydVW0W7CNrXgiy4728uT/A
gYSnxykDJxxTL2SqewS1pIueeRkeSsNF6Gc68aABcSlXl3MuFhUL9tqmWMogve/HV3fRdaKkyaha
CXyiU84WpNQtXt1SGouwnX7QeLTbUSSiQsRrOx4TdAmbXz6FxUqBZnIENCq7ZMtVptAPpUYxyl7y
eOaGi5KYRrvrRgDunuujd58rqkhuWk1sMDO6llFO33Mw7jaWtM5Hzcl2FojZ0fNhSDhfGld3EO2N
cY4OEblX8+VvFIbr1yeLXJi5YN/Ya9tf940IWI16nBgMpb0u55H+zOebsNl5w0PRSudP22KkB99u
GQkmsiHAVU/bFzPjgeOKdbWUoTjZ/6knxR4Cw0tHNW3YA1pzWLNmzleXsT0mJxwZuELqn5SE9xUU
S5zlcybFmeM2s6qkOd5TZXI+K4AOSB/VQrSPTP5MjnzRASoWDSCeuCcXXVExh1vhzwGqY6sZoOSz
fjEKDyjU00dtBTAXe59PTL7xsY2ppTadqnBmNHUrYLQvA3W7ySTX0TZHEvHVXmCzbPEJhy7J+RZ1
87wliKjSNzq2PntGbNZqy9jRwrkZRQQVI1TTMMTMdHmYuw7qah29wgqn3zTC7qeaOHtLJLC5TnsD
57+7LRHJM84SxnWpZUh0anSxMmzHyIiWz2KErTtmQmhncF10aaZHQMzsJTml9qYVoXUNHanlgX/W
RmpBR2S6C+fkNo/AAXE2seGleuXHQyFlusgP2rJK0bWAeSMvdO3LQr8Rg74QtK5hsnnbzn7N0Lo/
rB4mbhf0TNtwpD74A3Wb5yhnwKwTPKQNNVLZ/acXpUYsk8NoEoXgofRH3EObgSaT5+KrAT+npeBE
X9F4C28Rc9IvXY6qNzcDCuw0VLPv+JIWKP+Ww/VzBsANBMBFiZHKb3N3Yrok1jn5ZTF1llu+O4Hk
4J2PvbVDu2op6Gta8Pe8hytsIToM3bGc9Ns1rUAwP8mkNc+Mfk6ZrHkNUvxCqQYk/CYs+gW1Ilcq
Q3Kraaeyr8retT28amkmBRfKqQCpJ6Lgg0qrhBqBth0K7DwKRkft33kj40r2GiTNIF1Sp+nDAD29
QnmB3OXbJRGGiukJb03iAKXVjgJOEP/FaGHp1YsCjxCwkW7poNrWYEO0Hp3b+QuoX/tVjucgsuiT
xLs2W9ALUcGFHm434VVQxmWqCdSXIjck3x4f7px+JSSVdYCE6cLLjo4M70UmZC2pKRarPd5xycd5
nCLDh//DCF6SxW9Latb91ORcO6kwsDONVlcoXy1zIUyoN+YPG1mbCdxyK7fRGb4RvpWe4A5XcvA2
UXzdq9mvYpqAgW52qs8YBLr3Yi4zIOcIfDPPh9qokeLxOh07OmvkZeraI2Ek+cZ0gCafl8dGT/rt
JgEx1J1ZNmKcZx0r/W8VJsqEJQQWpdTZm8RXdxC9/2a/PZH+sShk/k+B5oZ5ZydQjc9Q84dvCOQ+
aU5T3wUGC8zlDttN4vVD6sCWaaxed1/f5OTfogEV8itucfeASY/4hoAMevsqzobd+DU9/D504zzN
NKdYrdQVXICg0ofjt3uU3X6RYsYAMOsLd/2FUdM/KUMLPMSmYLHVOxx1NfSdb+mGgzF8DxCtd/iO
TRQTn6LBBSwAE3n/zQwfx1BxvXXubDgdphD5vBfDBnbP65sSW0mUkZKLkmht//llmDvTyjaWQKz7
s1z7E0HzzDqA9cv0SFa+lww2iv5I8MLq/FvGuop+aaCBXpGPCxkme1G7ePE7LZpLEjFRDsKJ9Hxb
hOtEgD2tWWZPMrKK2t6RhzOAmGxrE5h/68GPaBvUixCVjct1vzwA763NZq4XH+LAMhxMdUrHZ8K1
qbvyr5V4LuT/Fjqeu0gGA/3g3LvrtrfUuksTalfiP8BrP1U8Yfhdg7hC/u3stTvWrVKGNxb2slAo
i54GWFiBQYSg6gU3Jdi8TqLstIUVzJDF6sVEuhh8Xdhr8KYkE041eLBRQ9QHtiaHuYh4S7GEmgvD
vhsoMMLupl45opOw7QjHb9aoQUwqm3SK4tSWEXPV9HY3y1h7PZX6S0/14Ssbn79U+QUDNDjq8eth
OBloFYUKqpsmkdyMpIwpuDHnZW8Vi8rVxSDn2LWgtWL9av92ETfQOdDj1kSaHxdIk5n1TQWW6QiY
tYEbXuIdZoKbSQ9L0HloGl6d6BGTBSToFcrAeCNenN5VqT4JODsitjmlqudTfAuH7jTHv4gzY5pf
R/xhpD2kNlPWLmcJ+h/N+aUblweaN1iSrPW/zcFrTAJG2r7LLe8LVwAQwBctWjjPmOOUK5fM/S9X
Br8H8t+lCaOibD3c4FPDW2cyFLFPd93GwaSpBHuxG9M6xukVmebgmAkgpOvJHypqhnjlrmuKsf3j
oiPnh2VnCesK5dLxtjAOd6+woomVpxtLpXPBGaekuppVx7334Wp5rUg6f3yY4O64iqMXmKGv9EaK
qd44cesGXqG+jMrtgJTsTD985ga5M4RXYjCe3Pc+3ktmWkUXsbX8H6wjD45BKhwqo339cxy7oGof
ljQleJPYVzfkWE0wNgJ1nKwx0fpOsw8YS3P9/qLu5FY73FwD9rVA6CwwI0B0ULYvGniux5Rcx4Kk
aXPtFo4MMc0rhZE8LtWDzwIDkNJRWwvp3ECbQ/DHIL1+foul+xyoUe9fga7R6+qSWq1XQSj6Bqi2
bsrUtD/RbORQintsS8QoZ+JrRAwJcdijv3koaOXNd0LYqXsYcmA0BjiAVje0Bo9yq9HdxSPXCjIR
UoJ2ySJKaGP275HNrN2tz8zLt6uFdZIo5MlzKRWrKhVY6fA/jsQchugPaG2TGvldQM4H/sfqUZGq
tSm1gQwEkQ/c1TwUp6U9S7dIHwjirYRfGIubZmgZa3QuNIu0UesgR1RCk3CD7+nEDAw0jVX/C4OX
3zt/vrbJW1IaYabaIxOz7fbYO8jTUWvxPvXwP+cU91gtaWKAH6T2PhO7vi6tSDIxzHCOpnYviQxp
ndDXmKREPeKKXEPq7mmbRFIMzlkwB08Slc3zNQjrwi+ChJ3XTAUpbVlaHXLOY11nwNcsX/4sO/Rk
fd4NSZo0kskYs+/Gbh/meiohAh5sip1xnKcIWc2QuC7Ktj6P2oP18ba1U9hWvBof5JoziWkMDqV0
2Q8ngiY8sQxNTTgZGYwEj6WkxrGdpGrRoqem0TAXSKeqmeTwEDvxvP/dja9TIfdQr9LFnYfR3vms
29SxV5nIntzSHQoclkXo0lTAVjrYgdAtSzmDPKoqmf8eG/m+AcUiZgBMpP9eHwW/CL9WcSlEvJ26
FyLxfoddZk/4lnCdrQUcEoCz53i4ABlgw9g5tXNXEbW27cAHyYw5XfUwrESQLYw+3LjofrquIAQ1
ucHv6phjExtinLsy6xAWS79FkXau1Y5PgRqndfHGdMQ62RsaM3ykR8aNUF+rW8Ji6YKLBhHPXeNg
czon6Z64ahO3mDUVR1OWs/+6ajWOJ4iD/KAmHrNqRRUVSSlRI8tnOiK+LXLG79dmMFsfAklFM81q
kdEXLT9TjnykR9NdjV37OuA211qsfDU0Z3BUEcRy03tnTY20yXlLj7Cfw0Mqwv2LvmG3M+A91c+r
uW02FA5ev9thHDXOeqJnbKGufRBxBSw3gN8Ka7O310NBABrIq3dyO6COv2ZXliWfZUneuR+iK63R
RfZhRBO3KBPeO9oWxBWNEE/2/qkvmxPlIsFlbrY0btW7NUZDSC4Mh5bWEGaV2WqGr7I99LY4qJq0
sjpoLd1CNau+n+o3O/rANC4pk8EDAqlR0LISSix3wkDmrIEAIpAIlDkAMh8/2pIDsiRWL9nYFgCw
Gog/EQJaxeMkEueALl7z44U6lMx0IsIUFXzQuccCkve+xUBGl2ICXnMEHuj/SprG6LKh/TBGZw8y
YShlmxgWE99zwYXZbbWZite81dGEXJoxthN4K1199stEDpRWYnDLMXeLVNcFRWmJU8kjpF82WUMd
WuqcKlG1VfQspgPWA0R9FD/Nql6O6WkViJe5JmThId1lTXU832O9SllyVZw62l1AjLB+3DzYiAoG
ZHRv179iABo8yvocOUMs5Cu/+gzcUpLGeIy7k/D4YLb5J31ts6tsALyphHVGLbESbl20nIALuCr1
W46tvgyuREoRFhlPMCZtzDRu8NQ/cVwvIwrB6y8618tRkXdHHMhJwfbJi0fNPDnwqd9EDJp0z9vp
qZ3xrvsQ6WIy/xon6LW6ZKsT1LJfaA4kGWr5wA7PKk6MLVthIYWQWMhLHp/w3hBu2MLAOClco7HV
MjlrSe332Alc7CzaiT9jVKH7jzWbLZO5hWe6u2TxFa+9q1lAi1WE3HDoK31CAdG0MLDkFSDZG+1q
/7kcjwBB4EQ16rQ0QrfFRPepS5CqssInojMbrlrdoaR5ZDMvnCyvjT9mc2wXPyXwnVhySVNhyXl8
n8gtRXORrxMuMN+zZqfb3cxFrKvx86Y3EGknPncsmbcdqAisHnOrZD53MDr6xaxj4XREx9Oe4DC7
BJv8y4CylwJ3Ki97ZUuLasSN6A0hK63usyIa4oz5wzTQ9dsoQecM1khY0dlr4/ip7bj1GVyjyor6
rwQoMWuJ+6c9hE1kfO6LCq0xK40P1jdQa++hEj6OGkGIbBdrAvj3XteKBzvBLvFknIAfD2fsIO89
aE90gZW9mbzwqc2Q4TX3ksIgCNGMRcn3stk4f8Rao7hmerWf3orS2cKm1+xB4c7XJINGZcQT1itr
MC0Wazm3nBOx4hXUexGdpIxOuN2eoVFAmJx7GMAwkY3+HUPwzyPTMQE0/wDhDaWwI9t3M3ZCXzTl
XQsKMPSkdcstlkyxLe+j6I1enMLeG5eo9MePsvBnihWy51pY6uhDR7wSWM7vbV4mk0yv8dpQbkQs
KCsQ7Bq7yBKG8tuZfp4jp6DU+1qYn+bSyd+8xaNWsjZzD6vwsqGjxTEl2QhwXb0jaql2c3Fdv10x
hC7A3x6EYFkKCBsXvvrARNW1YWEm00KdGWz4DH+4dpzbYnSUGFuhvR1Umt6eX7xM90UgOb13IVok
7mVNgExrY5EtgAKkA5tzk53BhJFR3BEH0wY++7hcB0L4NXjeyldz0NiDlEHYVTRsARTqPbGSZWXW
IdFsp9bU7SSaQIL9FdAAkucfF/X8NvQlTzZ98nZs5DuzzdlOn/28HWCjdYyU4l2J5yxDZ8/wmINV
zoK79aRWgVqw7TDQz1yeHdt/cY2nOl5yW8ba20P5F7RR13bgaErirNv+YHnfDaBsLJH/zBN7bD99
a6XUpXip7/Q3M7PIZV82c8XFgZvbpy6VRx0tsBiR/LouudI/b+o7OJff035I1uqjrpb5B/+/RKSn
Q0fV5kiXqrSp415IcfvWuStPEbiU4fxEdTdlkBi8OpvR+Z7PmfDNcHgzdQYJ9SIy4ORcUTwjxShp
Mp2aL3z4gmh+E2MYi6o7D0wDWhLI+GLDtlFu/0EUGd56b4x7icoiDm39j4Ge4LH+PDnctSvjzNfv
QxM7p+ePkXGK1RtSGmAl9Uzz/LAvENJMIHar0W/Mek1jYVdIUCM+jxiFdzizkjS71W2hdMw3OXFA
yXAajF4DnTDagqYgNKHrFAxxqkY6gC2U0boaeQHpzlHSi+9whGPMg/kNSWptpE0hyA2+KrA1+Hl3
J9lzoSJ5Lo6DuZyw0LDBZuX4XWe4NTiHYG7eXQGlrOnb5pp9xDlpvpFXd8XN+UG86bEKllndeuW4
2yjj0r79DkmPWd11q7VFDcVnKWo1XvUKyG2Fb26MzX6S4IuloGvX/uRAoV9kYAvIoUNP7efXrTqv
41TJCCQB8HDbI9sGQUQWf3Q6DDAF66frB+CovWQLqS/Ew1Q/ed+NBN2GiE8qcv11cALQIi8Ip46T
e5bZ2X+G2mE2CxDaxoor4HXWfUbMWqew3PkPXHtG+2Z66mPudAeD9XNsirfJGZuk5LEVoeqjFMRi
eN0YRbi+y+AAy24YzqBzfD4zuxR38ePQYLL6yKaBPMDeIfdcfWhj4D/0smXcEe7SpmtLDWVtavE7
sMDmlel2AnPBG44iPo6lwNIEy/ed4CQx9tRP4nJqxJtn/3Pkf96jruABuPNBFUxOOmG7ozuJUSEG
xYkrgLIJPCc4ePvaWGoj5OfIlpt49etTQUh1NP8jkzHLUW5X8N/agrgkKfAME4B+IycryTC44kXz
4z45OgMdXzxT2UnWZg5m0Q1PAOBjH3HnP24pcx4aYYl+rDrjvvTpRcTOnJxdZvTp8VGr6Axzbtt0
q0ZZ5yF05Bjc81S8vdxQ8b+f6DytilV+MBaIdQyWxxS2QPnZjJmoDrEvvRi0Uz8UnUP3mRaZRCnS
dQeRMeT2Quu4b4gm1kMhJpzgueLTKDRwoVxllNFl1TUlybXznS/QwhXL6mcq6z6Y5Eng9k8y/Knf
2Lm3uBpAPsW1rriLPxjI17/DpmRSBrfZqHZP1t09VUmAi6a6G/DGmjTi823gn9swJeL9/kt3a5QW
9AiAeLGo5GN5MV8cdugrSRZqRt1ZxWNbNMwtGKZATXwkxJ/7rlla0nL5/FIrBm6Bty9Ale4QV3gN
7HTxm2N+5YBq8m8mgbRW8HBrAZOOMXkjM59/AaEn+ruUATYeq9wVETZQnGLllQ51U+E3w89XKE8a
5W45uUu6G4JDjP66rYgCTFrhSnSmd8yVVkr2d0escJBPTCjXq5LCMIvnnObmFBBkeszOABfOYkLF
cKk9pzSw+AOExvaj6stpuDj7v2w9OIltRNSUiLqi1bcxXsGKjVl6pwTwP48shEaQPdtap78sV4lE
B9Z9qLle1BFXZ+P/HYn9dL3Xmp+M48xT1FXm0tVaCNPn6E5J1sffZYtF+nxl9tGp7ZoKBFuiD7QF
EPYvkvnzkee/UeWJIe7qAY4hNH+Yd12W0e+AKwyMiTc1383cSxti6T182+YwVHB+k1ldnup4n35d
OjA+nB9gqz5zIHi455siAi9AkZXfKpD8Yqpm/H/ct+4+0POzl92poITelUi+AKsXv9hgIlCQjLPj
4OswSqEhVwBUSdFUawckv0xvzVE97OpXLO/RiJklk0iPX5tnEgeJlhum+9m7f44oVcSEJ+NRXmCO
+6O0kfZwvlqQw28wc1KxJf0eScDFxiZcOQgpq/gDQntZs7dVmxl4rfx8bSZgba4CEwr3YAmdgrdC
bYIV8gxepj8b5ckSA5pDCKVHwhBRVHMvX2m9LyBT/BKNFdKZ9oYApc64v/nmGRcq2UbPfr52/N3e
YL2N0WxkxeCGbkk00CXA8hGbNsj2lc3YSsdr34mbjM1qznu+oZO4U9ktLIth5t8F/XgW4Njbnals
8w/8bhkBWvrB6EC7wTucewKysQuqMANsCU6ONTaIWwn6Esye7IZT06288wNpINfrmR6DwC0NZv0T
O2snseGF1seyUbqsFZv+xhQJbYwRMYJA98buUjQFYpD8uKKOweOa4XIyZbvHLlWaPbMStbGbpDl+
rkvJumyXN3VbLEPl4zKtOycbGBkvzmG9Xk3Zp/dNZjk4PqWQ5yjIaGMFGyORDSh5SQG+xq/l42Yq
D2hF80TGAvX+SKrBGvzko6xiCZWLJTwbPlk+yqXjKeQLv20lwCFvflGktVbg+Bu9aUyeWTPaY5Gm
9ixBRbDbi+bHxwdB6zzz05S5yrbWmhXMAyfKsx8hVX+pJ9ipZ23X4aXBXWYJPbrA14M5874lZanr
1PabX4ZZV8iWSl8ON1QXuoRH6j433rAFFGKZl3fbHbs739Mti3EphUZLPfQeOLQtFSoOfFyhs/Ld
GzGp0R1LK/yA71K1pk7ZtNP1zoLWooGoeKEnvb/NxwSxVhXopOzdAPF5z6MybHzESLBli4Tsg0mf
OPVUx7PtXvEiffOh5IFv26wMeBx9z4kVmoG3+bIK5ID28GlZoT/3ssMFZEj/eLWt5WBvkAmX54jg
ZHUQiAMP67JjhOajHjGpYtw8O957StW7lgI4kQEImpsr3aj6bcQJgtMfDgVN9pFGqQW1M/2omkmz
gW/+fHjDPg83cp0nnXMRgCM/7eInodDNHCkunE8d29eB7nTMrccMDVplJ90l35ttWWFj3nSoyE64
eC9ePhrWN1jDOPN9a/QmBtDo5vzW9K+7wIv2FXeloTDcaQSyuVD+/WKBW6m1/pQgBn813bOM+kiD
IFxWx5r/6B782yFr9CZuUuC3ZPvG0w2fHv8vSbF5lS3oKiKe2N5obM5HaMEQWvCN9nFVX0nERSnR
iZUlbBYJuaEU8oigP0T63wk7ux5ywBFt9fe9vYKsrK8L/0kGolPnSjy22yTpida3tSYtVDnWkrxK
W1s6QfLwLS1+4exzXK0hULubFxNOrpe/YdZuMZuOz6S29J4LqRTT0Tpyj8LLZR0nGhwvONWqEMSz
6JHRYPaddnFina9maacH9E1gZ60GoBL2YziOpE+D0Zm7DLJlXqmcG+53OVc3T7hRDdUooKIcVQIj
assBVuBUkhCKIp+t9zjyUUDaGkMaVAaGFrJseSVxV1Bxw0hC4eJ+4Pkx4RMVfYVuTIRk8J4qLdiw
hnC6Ys2wpC837hPPxOb7Lr0wvjPWi4m7vB44QxgK5K/TbqSlvNYKStGvczRLw9IwvbXTJfMKPoEt
FTb3EHOrtN86dV5Yb0Whjt21DKTCqr3CAQFsSexxuO41v96G5marceUHrDadGakYlj8nKEkZU6wC
J8W+/YF+WGbIFU/uB3hNfUwamGGYbv7+F4dOTZqDBjKdfFKKYk4J4iKGcBRPHmAQHxpAkoKwrFKR
0zC2wNONC5oAiVwWOFmDv8BQZzx1KcKV1ZQsOpxGLsxoRreLnShjq27kwXwRUd0jbnbjfeMF1DQK
fncXsMNd5Pwx51NJH18rarzvYJGxlE/tS75TLcH4X8dQp/34ULj+IiIKNuuI5TEqUH/olt8ARsCI
uGK7szwOvCYK0r42gMGrS+yQKOfarHbdEZCQdbHZ7QN8VerHHNZu0XCbT3QJMQdLtg6zxLMSBKcT
mAwAMYH384b5pFrlo66jlp6NJKa/32cSwiXNpy4AHmUXk2iQfak55TXNeZRS/f6l1dNFSoDGR4W7
rDQTGNcgnazWmUIhadwP2jvblH06r1Tg2RL78E6PkBY+PWHWf2B23y0LlwfUEGJdc1OTKVItXru+
TzB7sAYVM+6P/0cDt9pXSgcizC8+va0Bl5sDU6G24mQsOTFzpWGabjs9hQuAbVcH1nSqLDb6vvbo
SsYu6hdLOCuFQfd3MyWFqgTf7Y28drR0gX+d608RfEDlCHivi8FPTRHnyTiPaTLUQogmc4XdD5j5
xDoC8rP09N5l5z9OSWToeEYVetrwZTltmjoOTKPQ0xMzrFTgclZhXfVJ6yFks4ioqsRlSMvs+7rm
u5HDpspQ1XhfH4ROMikefcA/WaC437boTOZHm25PtBIFSKaNbH8H0VcMfkOKbwb6Q/78o+vq7ogX
Fxwjccsci4Gp8XcNp34sT1WKqgCwGQuJMnr4VAXMeQkgcf4r3Rns6vepMr7mxM9QXG5zBlRM3ec+
oft8AniEs7h7NCwaZfjXNnK8qesRRuio4ycFpuQxsj4pI767KeGxyIpBDJG7c7f9SMWvf61MQccw
HF/bJVaWQi3S4aEWNzDCAwccR7yTVY+vMwZKMG4uLcwWmo+IUnn7yfG2skVLz2dRK4Wl+wb2eVqd
/st5ivFp0MS9gqmbsWpeXvgCWSn75NJELsZnGFts6MqYwo/ttigNRDy25aA+3E9JXtyx1KDGxTKI
t2bB62CJQkkRoxnCQ4cwyRevvztNsHp36EYFlN0ouw4a0nnyscmj8bA/BimwoJZNbHjqCp0d/8M/
4X1shNKrTO3yHOzRz9m06F4RqMOEOOInNUG0zz/S0s2gOq1mWDUIKkBo1PkUl76JH2K44WUc+I6d
hMYhvfbHxNi+zM/SzwaBFp0klucFYwexviL+YbVLImvmIllKU3ju1sA1Zsh0E/I/ipPcVBdAspad
OOMrFbjjXLyRYgRcsQvTXw+N7n2Z9p1fvT49it2m2Y74NI4hkJLaPM+H92CrFLCZaP1D3osmuOi7
Aws6UpYFXc6t39yAVhkBH+aMj67AcHKdA5J4tnbsTbGUilaAEt5/DjdouE4Vc/TDsmpIsokMUcK1
8buELOEhZShha95FpGhZTqsyBed9f/lwo+syTI2EKIhQvWM+5XgEpG5LcjI7LkWq1DOHvvgzsPOA
tlqGD1UZ5NziEXo3XlPtdLSpahyjHpNBPBJ2JJXlRa9z7XmpxyxqZSvmkBtErqtWyQ0YffY4SFp7
WXK7sU6zvheGmG5hd5umhEkEBmaYZPQ63B0XaJbbLKyAsOvdJwYml4KAUzXJs3p4SiMLWj+WakOS
Ft9oemV1XXxOz5OKEFlQXWH5MuIlYRmBHU3fnwu4YZcSuZWcC4fgI3F7mu1E+sgHSOa/wGx3WERz
RlFAm1VZ5bhiFsOfrGTTIpYxplo5SspVoV00utHcxDerd4OI2HWuKqabt9Wnxj4Aa46Pg4Xs0dJ8
XevaF2i3fZm9nNoYI6aFjq8/tcnV0xPImuOi6WB+zhpOL5xTq4UNZi29S7NnhrH2CoGyLLt90Gw0
yT1qGUEV00rrBU/qWaxob43esCfFoWElEk8XTejcagQzlVcNIgvvlvDpgq54YV/78tQt4Sb+9t2L
roG13F0PbKlWnBpJ+4H60sF7D6iQM+jtAYKHHsenBfMDxjRHNeavi8dafuJ1Hpp9cWmyovDEtOd3
hZrBfjt3f2FcMo9KvPNB64ybdm8n7bc5y80NcVTh5G1ONwAZTbAL/43hbuLDk933wFG2x6BltUTc
Xef3BAmc8nV4mnVDtZ7vx8rhb7bBbL1MXx2B6K7pSgX9xrn/TpCXXSftFDWxCjWI4ppKHRqz3zaI
kS07Y04tz5jISzfoLCI6h3Rw6vI3178gCLU7WNPKE75Oci0HCkSLpUKTkxyc6ZJrvM5UdLgp0/J5
fZiMxXfc2LLyU5sUaV6yxYiVCYKHKMler2oLLYLN0osjhXq/gGA/SIfK0rfdlS58vnduokEeK5s5
ANMWRntmES1m6KwAYoxVYlLnKChj4ADYUBceFri2n7dIXfOfL7yc2GISuLmFsIkp9ueIF8gRpk7J
xsa6v8Quqt/x4WZhQTP9worI6gNR/3KONW24dWGMYOMw49nzhUlifKAat3cwePX3cluHIZUE9+v0
fZIJ7LB9ifPR8Mfr83gTMtFwF8nH/Xa4IUjqNRYRghluWQwssCzR6OjeFGnwDBeJXZ0yFJm18LpO
ZDl2XnlHSeAKeCj5saFZUD3aUb/TfKNVysguS0MOWF4DVD76hERnYIRHSCG4Ofo6WP09nCnvYD3g
PJ31xHyyqZXAlCd9GeY3JTr64aO+8z7VUwp/Hfw7aNilCnb2njeZ/SycZDYABDrQPs0HDfzD7FWB
ImfDv43ul34JjMtWCdjbOPraL8BJ03GGoLKYK4uB3IhKyO3x0OC+U236E2GqC/AJ2Nk0SMU7EuMB
szixc7apPOEmeKc4r8Uvi7S/oJg4arEDPgGEVJXq+bd5qFjn7obIi9iEzYh6IkNTtN85BHsxcy0d
fiCTgTFeXXywnd3OiS71bSwvNoHVp2DOBsxKraf4vWGxm+Rs1N7HJQmxXAm3vsLNy4Yud0T6u543
OWKUFXgPo5FLfFmQm5L3dVcVttBjkhxiRL54Numkxml7LPWwUXLCqhWXX05jpgvSegnRlNgCDOCU
xxiV+FtAiS9nO3282Lh45v5dsLuGjjevWbALDFz5vQTQFGh/PPtvWVOIMY6tLcwIw5a3y3AnzBez
pwvVWr6u1N1QB6RZxQ3jiXn00XXnSzJxV/TXNP4a/0ai3Nh4ABg/3OPi9jZqtDnbkUj3dNpXdG0b
lE14/5EyrkU+hsq+zznbwK710ZPXrAh7oG7CLE8cTBfI4gu9SfZqb2Yk3s/aWeCFzBbq34lg8tX0
jwaeJEBRsM6UoNrSmnz6PYSPURHkNls/uCQeVS+Hd+JPaiRCBXgWKkOX2fzfcpCbx7NZbTxx4WZX
aSkluvMB97Kkpb0RKcMBJIxe6lgHr1F+GWR+YL2gYrvb1Py2nOn+f68s1itE++mjayQyiV3ddVm5
b7P5CO6lrlz5e78NVf1PpVQqfMfkGNGKoZTRC2WzB8IF+hYgvmlURn93GqP5yXeYWDTJMnU7IAYz
klV9FQvKfBU9HJkjmUG5U5J47d3fN5rpML641qz7JBCVQtIBBm1VEgLiGYfxn0j1MgpFlPEsC44J
AMekjqzVYKa24ot61Rq7JroU7+XZN0R+f+jU1ImRazefeet8rFtbS0e/CUAzPWYrz09sBZNMpZqx
SpVFx/o8xZU42NtzEQ8NKw3b/L9sYdc8FkhcPrRl//8Kt4mPxxPswtOE6McJPtGWCH+AG5zClFV2
qlVCHBD0maw3W+AZ7Pwtmo0wnAjPaSJKqoWuQz160r+No6kPw1pLdOsKxfgUC2dtucNn1biH0kGm
13RLn+Lny6IN3W01e0VYcEDzVtBjy+o8lF3oBY+kr3QRy7mVC49Voefgz0NHJaeFYsTSbZKOXF31
YitR69EOOOjlHnvQqHeNF8lx/iTl3eqJM0TR8apN9VBEbB6mW9eS6QL/ui1JKPUDW3QmAEH8LZOp
kv9UQuUm3w67xvD1W4YRGCTb7quTvoDu2Oc380lVJKFZTIdstPoEZJF5QxVp7M3rtDR5CPUzuZV9
qQAFEp106hyZBrCRjm3JuPXCS52xdr3iAK7F6oXCRH4VIiRtLa8nt0x1BUnpjT2YXDaOI41g1psd
UVKeuI3a3Dooi7rJJGze0jnzc1K7L12qxSBmHigRN5MsN809ft7pL/LnjDlmUB8rCkNIqNK+oD7z
CJx2LuejDFhMRzac6Hep1Llo7x0Wf8k3zncbYj6JNq8PdqCwZdYghp3PHmhOah6FiMWvZSsJmSbJ
/BHFaZFh702VXudtWNKetZtoMBTF9AEhqz6H04jNN6/7sK9UUhkDRjQEWnGYB1CE4JPRUScoJi2I
biNYqHbr+J/Rvjhr8fCXJP205D0iM6xgNRDe6mUpKEHzaII0edg1ysoRFN+HPQtJzQ/4PtJJcSux
/zBYteguzSiqY4C6YiNsFaqAdX5ug6bxbqePW5SxPzsgi3mT8A5SCo7uKSyAvlnqjQJ+mQ4+ld/m
c7Iarq/wcIc3ktbKkQSP8mpq+SlONYtLyIG/7WwGI2utlC59tYq9GQpofOBO+xJCZiPlpVM08yf2
G1PVCPoJlPQ4pyVQ1sRZ52xF6vKNB990L4je9ZoGydth76aDqVBdl3Bu3nQNPqsHqt2Fkw9RSZsA
X4QD5N0dEPPI8HxSHq5tWVl3jmCOYYuBqbItjG4bbld62zkJaK4uiZcduHim6oYijiAmCqzmHuhq
WsLkwXkWU1yNLXk49k1ruY3hvHXxFaZ5YJoRUxFPfE1hTl3mmlA18EQqb8B6KtUGEtXn0f0znd80
yRavrXysDZxTE/j2LxoNSszBZnp+I/GPUPjcD9b+WqgWdav0hAsK54Dt/ePaqLI22z2GqR6FPuwq
H8patzKYE0k3a9QmrE2EAIhYfyTfN/YGZtnFSHrbMjCcKsgAejUfSFqy4Hy67ogENGjmsAkTFIUV
3YOjX9UTTRKn3US9ZPS2DYyxyBTwpWMtt/IAEqlhntaO9OKRfvajzL7pwIksHmDFNW5eu/mVdnvY
TsgNqhRY1ZRFSqGU0dTxRg4GR5qoFKKf8EqQmnPjGzt/XzbpzUjYNbV9rUV/IFZ2pIDStXuJTMTE
5J/hFVTHWRFftksvBdcxBveibKqIX1B/R99yD9Z7VkTx/p7/T/yjSIyjBNz/dxcEEEVEQ/0/FJDO
gdLhHr9buFQWK4R7xzKGnYKu9GDS3DOQVDKYypx10BKT/0+c5IDUY1jwF7+bRDHbA45LfChivkR2
ErQomojm6lOU1YhkTfifkanQAfA3ngSqRE8SzDPfmOKmEJVOse8JfoIH2fbPQn24kjYUxOU5wSy7
HfUUyt16ZOBRidJU1m8tgWDeLTRRxg6NLisqyRm2/eyu/uukEqutkXlDslzB+qIMJ/lKXzKl9LSe
tjvJf21Iz+ZGPmdiqJoddEX4dUzMWFf1Nk+41muPGuj1ty0k/eHyC3R4e95LGgf1ON0cE64AgLEH
m7Yz9VnKrsq1zbJuzcPHAd8uEzcnmY1+gOf7G0CSWhfKWJji0cIs0P0dLtLIqQkldcOmxXTaCqSk
0cHlco9lLJblLcWfbgjGLhFKa7dILfw7rHZNyZsj3gALlZMlRhxEkBQcc/60ZgpJZv579LoMcXxF
3fUYKLZdJ8SXI2AT0JVXjH7xFQk9AdpHOXvXymgYvrSckOOc8NGQIqgoC3CMnNiz5IeETKR9xNUj
vd32ocltAgTg8OKX2EuTqvXDfyr/jWnWNQXUqxERGQHLRhNS97jgXLThJvlwwEoaW9Mas0uv3TYJ
V8L57OXWo/d2xibJTaM6E6/kp8i/tqii9rvu0CWfI+VSpQ5m43bewDekugJteU5S8dFXVbQ/VA/Z
J2jlvwdUCnyEsSmDzCRkyo9nPXz9bLbp2gqs88eeV4uzPeE5ymD5tXZefjDWYTUPMcTlua6S94us
P7CNeh8bedpN6z+j+G9oRNgJtBYXKOJmaL44Wdjr5Gf5nVM/F2LJvTInD5nZNwoEiVg/ONNKs98O
piELsequBVk5C0HjJzUDq/x4jD3PwuHmIy3f16nw6cAREsen4+Z6zTT9RT4J7/UNTv4SIK8sXfPB
zQZD5sDZMBw/DpgvnP2w21XWYW2amtgY3yVKqEF+1+2qizpjz5MtDRmaGHkA6Ly9l5a859zYxqpJ
RjQWNy6dUXRVbxbHyQjT5h6W2ZGEPnIrxzCVVxDANwGDRZSpwS5fDncrJwPVkqNwO1MAxBOVwOvk
Q0HNEiZmU/jvmn6jnti4IqbWYe4GWku2YUVaSf+2OBsZa4d84LtKYxHNbe4yauktnIXy1QsinNZL
hpP3Mly2esL4N4W/PS1M4qVB6fh88P0ccftPEJw+O9PI+lS8DecbYjkSj/rhFpOsOCFRfyvz0kkV
FcZlqB3drfK0Gj9EoRRozMlNArutWuExh/L4K8vkrsC0fWG4XbLmlSdMC/RrnOGQJKL2vn4mhd6G
2C67LdVhm7GKl5lDs3nH//JjkIKOdPnXtLsoHcNPos/q1FTo/DKYQAnppt4D1ZGu0OCLPTuIJcXV
4fU/upo/QrE+wlMISuCPjb2VDTGjF69YtbVmecFFeqbJoIxoR/8jDlJlBW0CUDxtmjXJtSbNT+Gi
3FV+ByJO4fFaEX/y8qHKWMZ0mp7+2JGpaWAJPdSB5fc67ucordcaOd3qpczbOQgot2aZhvlwGTC8
E52DVaB4L0JQfrL4J7RJ+hvzQW0mg3weKmaXthPLPNOWfNQSs+0QD8W/ZUIOPIgiOEczqUIb3xDn
znIVZNdXhab68xmDJttD6Ftumg0R5Hujjohe725TalSRjZgkfMyvJVggOFHq3JjycEWl38Bcuc35
5577e9R4C22JGK4yOW2bey4XOzwy5NlZQpK2JVdyXLeB0bcAbi9Q7WuJpplpLmxKwDyS6bip84Wq
SlbkrRXV4IsYNTswRlLZBXgPUj1WVxXElmRoWQ1MbOQqEWyy7Yn+CWCHrea9gh4qp0eAiPWowUC7
UjLEWFt7aHLEkrxp7ZnzuijvCZVemJCmHWFMMi6Poe4ABipFW+xBHtNZkEYI8DYjChWiJw6eBbvZ
2k8l59Q9g/58ndx3HPzq9+M7BxVboQYDUe/SVW0BRTibRda+peoRquAtmuwgS87iOeuhRV2fP1yh
pnC/Uk3zdgGDqrPtv1QoSdOnDZH5pmY+/6zy7mBttda1cr1H2xp4N989w3LGeGy5bxfFpa/sN5PR
Yo9V6aBT9ICaBRSQUVVVvuQW0MxXEeGAzofFN0BzCBiFgVBqUKmRha8c0iCMtpa/vEVHdHRuC9CF
jnTnissalWVbr9HYjtBh7tHmiuxV1MU8sN6+DQ3lGLuhSYDGDl/EpCN4T+c6qVpqA5NmDdZ+YhES
D7bOhT+P0Am/xNQX05tX4UjVstt7QzDGH7ZqHnB0yWASdOyGm64Zcos32P1vU00arz+NtR2v3YUP
tmK4eZd7UgwhGD4yIsAAlQQiVmqG8Nnqe+ecNNuljXvkZ59+hoA7+z5TU++b4j3D6WMH07mRHFI0
hqu6OyTn6Fpl9qaqRh+m/XFk+oLSDBU6O20ulvleDUidUmjz3wwliAWLnlhmUZzE4SzxiD4cu5uI
O7Zkc4C0Pghcm1YBYEJz0O5CU/nd6GIF4Xwlssh1l3p2TD8dy5od+4MupBf5jOmwX2PlRgdTN8Uk
VrelA6QQ+n0BfFz/1uMam3HTqjpTAI3UlOnH2xrOPrOkhweGKKzudz6mqv4flXXu/VC9rWsiz4Kg
8UEazpPquQlL9Ixxa3akRBN5FqjBh+0YZ+tOuL8PgH1BQs7iCcEYqdvIGtVgIv14hyVHCKHKlwlZ
agVY2jKdf+hHSTFpikNfFOHd9EPMBdn6hqmcXYuVS8vrs07Vz7/EqEVQlz+q2Fg0TaGkmIZE33l9
ySbK4tUeZvxJ9qiC5lLUNm9GjLSxeMTomP4FzfSMQpzXWOQgrPkMCEcfgfFYI3Z5Dv5KTq97HrT8
L9JcyO9ETE+MROrNpmleUnYXHWdR2ZJvRVq+1KayAl1QPpbTB4PHI537BoKdJw+a7EtbBe07dTZ1
72GfIBtnpAr3oFmCcmHB84Toa5TaQNT+CL1iJUbifxKhwaiHCQmovpEzuUeOq3q8xahlnmyS4fM1
RKH/hoYh+0+/ML13XFBQSpXUv51lnXSn1npY2DhPLHUfcyduZrAVhaOOvOcqCT4LwBVqx9XYmZwO
QzXTdDxM7VK3E+YIoCVgp48QxOsoBOsQRfOjkA+avoY6gkyXP/Cfuhxmf6oOQdNVfrX8OwsSBwmC
4PiQuH4KhuGOPKA7bCURjj7cWL1+lT9SVGzKu0KqeVnCoXKs4pXLPjtzFOPpL3DgA5Qw9YdOeN+b
TaWU089vcMudIv+3NFhRmlkSHiDxD4HGylkVPZ9qnQFBHBu/N3s4QqvtLV879hXPF57r2tHnphDt
XYTjvvHKIEs0c835uuJspTdEJWgvtyrQ/TvT+nYcHWhpg+NxR1Y9d5YTUstOyLEVb5gUcSl1Eplb
nookHaX4navPz5rWUSoG0arH+JLumuitp2TqfMqWdi7JsHD+DfDT/cj3BTY5wxAXRhMuDK9BpRqb
Fiw5Xu86O4FenXm0LZsg/8FuRA8fXldNAm4+ID41ztgOl+TvHrZBbdY422haAw26oAnGHCE7konW
VPLPkXsQt0xsKXmmLC9hDkfLCIUo53X0GOYc9K7pwhcO36quzyI+XICaSpBHcllvpL9bn5L05CVj
OShqNdwESqSIAjzrKqVaaTQf1+hWiwhwvNDtCZ3qGQ0RfohDjIPvtSLxRdg7evXuwT5TsgVO96Xl
93PcBygQAl/WL+Hg2tc9FSnZ6DaVmLfnqrmzos02N0PULh3jAr07QTcfJtzXAl81wpc8IjVbORBV
TUQAA1qruSVsthHpKsrTxOpMUvMTIdkgwF7SP7lZ65CewQX23jgQKQmhYnd4PtSEWzjkpANnBHQu
H8BbEvix4wKq80EyUatYWikFJyOZAogTdV3+4/pKND7BvT9ThCwdO9AtCRmabCa8UYwhcclnvYcI
MAm+DR7oPg2Sh1eilqYcU8IPdNwQ5DFfHl9QCzNai4zjGA+ZJXFsTuEiQrsH5YGkq8+JGqPvKul0
biDxs4TWudjQPStvEiKR9ucN3AIvrXxEzaEQ9R96SYLPe/X7WLCLaYd7YvKDRQ5gHb0JbG61jMX/
nt5TaQLIjZUzPYBhApSNhyAFYLW5FVH4mTEUGF0GJ1JXGe/9gSxiNhIPHOpSA2bGWv63urrvbV6m
BmjP4kBz3T43YGDvqf/JaO0Dx2ouqFUFkERL/zxkFDnYhSoPFMv0nv9tRwhge/pi/8DwH2oz+2Yp
UtTBmkAWpHcqp7W+vzpJFAX+eYWlEz9wBHRm2t8DDM642fI2JQcTPizZxMrBGy5asqiClF274ME8
HER0TloM0SzV6n+W5WzuShEv3LjnAxvwxpFaPg4s0p2h1Qey9A8XeK8EvrO479rsNTcOK5DWaEIn
9ABVsYH6fBfN/3pzbpeGRQhJRbQiD+VmmpxPUYD09iS32y5lf973d7CJPKNkrTdSdkDqldQBxpBs
5U0rnRk0v03o4cTXyuwPtf7TFAk3B3XKibQ3hhKxZPjzHA9Iy3Lh7HoZooFGbNC/7hf6cXD2i+iF
/VcWmZ7EpkRz7VtHhls9hSNPPqw8hQr68hRh4L8y15eHKeixiS90W6xX6UIq1pl0RQw4SfupZ4s1
nlNuaUBfVPDuOZ5C22lfgQPOKhAPJE/PKdbR5VfxBmE+s6UP708cPNzxJxRrma++llDZuXJCj5X1
/a9+C77DJqzQjjfKOHD7qgWQiGXE3BPn5iCZLn6D2NU4R163lD3SizlTo/Hu9gOZ6+y48VRU8ylG
Q6/vxaCZvKRuH2yMZywExpFpg1nVqMmf9lcYpS4o7Qp2lf1KYDt7h6i5RKMiYsNFMnuUD3v98E9q
LRImYYo/iYO0XZjhdo+F+Px789n2rq5U8+MSHVmeu3cfAOtlhwwTyEYbLy5MUo5QfK+/LZjNNrvg
TlKqZmFg1kE5J37Im48Kg4uzX8eym1dXm15Sffuahe+EckBwOs62hUBRuDbBx8YerDcZTouTfpME
bnho00QvqH2m0myM8ccochdZcgrn2nL4WDA7MJQVr8u6sbVgX6x4Zeh7qr+px80KAQqyAuucF+mt
bZ57kAuXC5Eagi4z0TP0xs8vJtUIhcHwLEdVcEy0/aoXuN4xGaCcl2pXTUDwqC4KQITfjwkzgjKm
eKKqjMt+HtX9G5DNu1wFrOXly5PPc3xakYKW7wxIn3nuLN2NHsidjgdShEHJydj/p140O8mTimdb
w9HU9VnCBTE7WBAfkumzI7mBKotpeYLSRrVREWzyG5eRpSQPpuZlG3UVnBWb9ZPFamBnzltkhnre
AQPonH9cOwEilbLd4AcmM2ebUqZ57wLNFDKAgVUDXZf6l9d1JCb4aV1VCR2es1mWPpFge1qY+UYz
T4IoYrvu4JuBl0qeWPtCanCyNUOoJmB9Wo3FMVAfElajz8TMEhf7X5+HUouD7Chj1xzpWJgbKr8H
IE6JpdXiFJEbsY7J8rev12jcBV3lqoLS7ZdUNt7Y8mOFSqrypesvxWy+shtvZV4bpKPMsbxVZvwK
1tF2P58JypW9rLpnloRpp5AVY2udVdnIlgOvHrx2Fr10pKDnTgChmg0rzR3G8sF9w54Eb8AD1dtt
IXPjbTlpQvrRy5L/UkkSaNIYLNLDYjkatvaCoCWehTZcrYub9NcimugRfVMBvYtQnvRwkyjutaZH
3uKehgsXCak9c8GPFCNJMAjC1xPnCRqXweqMkdrjX8c14mS26AvijHP6Pm19xj7h+3Crp03Q/GEf
R2z42U50zpDVrTkw1oV5YekrBOkBL0b8LBydboK7U9KOIhEXsNRlQJkmM2sw5xU8kQCUZDplYZVR
ZubKH1h64v07pImiPeBbCAFNVXHEvEbI7vhw/E3/4tfIKdqo/V1I7MFyCpFMMqF17OVuwSWhNBD8
4lfpLTTPWRXcy9l7K+NwLzRoN5GTTgqCbWJvY67kyI2EYiaXHt64jzCp5e86lM59f/wdnjF/m1Wk
HX40H1N7HcGV6Se3VFm1DMoGpvBqfDyy07AJVfuMy8kj4hoPL4FyBR/qj1+vwWFLlqwX/8m12Sfl
5pXRmb84jZf1AWZvLVQmUl3csgQT4ZrWT/Fp59iOuDWoVDzL+SwdTWr3CSH0UMpslbmtVf+7m7ia
7VXERXde3tRSvjXvNrOMOxoOo3tdmDStqmvjLVKSKktLWxLbqaNJQV5UX0WmLdqjiH4IAV0iFdUv
nHPwIRkgdG0PNXvcsbSumyV143z/NSaROKQw1l4aHZM8ZTXG5sEd6KDERDGCUVoayqkvYI56vsya
i0fi2U6H9Rx5wGYtKnhLo7MUYNKC1JOBGJUOoV9zYh6xej8mUW1nzGeM/XR58JbTs8BDu3YlwRg5
vCoR4wft8kUlUAMUnSRsDR+nM4/y/bySfpE3//IJWv6DXD4PVecLYMOYhGIU/SssJInlx/oVyIaI
lmPf32XT9suE+eLhxWx63kfNq1HQrV6cWOZ7or1AeH+Q4RrLb8GvZSF2OJ5RVAfTsXSwJLS/k2Yh
17SGqyiNNsFDhP57pBPAIPRHaReOULgG6tq8omnfOqnl7fVFuOwf6KFcFZ1g9yF5pjh0834zSLGO
HvgpMB4WVmQEusySKi9IX8hmIXYR+T1905e/mKXLr91QgICDg13v4ZK5E1kBq3GlWP2UyLw4cvTY
w6QhIE+HVfsD/GoW6EemT1D/AAnyMOR7emyOMIT23UsIjiWQ2Ej1VYTupDMA6xsGeKzObOUGZ2xX
fdqLrn5LH8popOtXhx3Mn+sdOPjmINmRJlR+SzCZttgcCEctSP3vt0k/d1P6CZshiAoYNMz5zR5U
p9t5jbub9KalYCYIfuax17SjpG11L4EnR4Hr4CysdGviBqaZYamlKJzT9pu3DGiV2DL04C8mRp5z
LH/omnpqgrpW/Vc2Bkd0cBECb4wDXZENjOO0PcJt+vnTM/RG0C/Af+FX1wxgdTMeRWOef/NWLMdU
1Ga+5OZ9NV0XyiUGsDO+lmQkltM3gQOtC/yh7j1mS/vm6UsaavncASDrEbtgMdXWCkcr0v4cRQol
XtbY1sMqYCTqp/kgzVZCfLTWFsPV9qYs5jDGZxGq9c/3fcVT3+KNSqttX/daGkifqxzzDRQoi/I7
/WrEcRWC510mkBPydUAt0O4Himy/D79DpPSifj4MyKoSW0awd7yjA76gmv/upudBZxibIrGCoef5
DI9KunBGjNEXF9utAv6sTOaFLpoAJsLbmy2R41ad90CH1rILufI2BXsYCA1/xMC25KUX/r/oHD/E
q9+YqRduaUVN1qeHeNxue0a8pfT5cl1okldoR+7wDKxhzUY6Sz8bnNdis4gbiysUptvic7pdLxPz
p0ZACrNnKru2ygFEdlUacM1jVpi5U1O5LTFN8ki7/uJVmpuIU718acqc0tHstiCnY39p6fU4DLul
+5of33fmPp8e3Yh15mq1FqAJToSqd+yo+5+HLkXXcjonTe/W2TMuDFCYTy9O697fZstwwBs/37lf
goH8tdF8sy6q3THVnCICxmzbsFZVJQbCUN6/fk9JdxMdc8hukJUEWCyYEvNGzCdPaSb6WVMcT27I
YUgaGy8tHXnhIX8/Qn13U34LXJmfThzi05rbRdoWuAoA4wZDdu25+9JQaLgkk5hs+RwJ9N4AQKpz
fLZ0IW8YrIin/s4uA3l1JmqYvMhkgR0R3p4Xc7hEku4uCAdA5QthqtXgqfjkeKCC725HzCRJvn7V
Ug6YIqmjMKgihA1Yns/wfHO1DM4sqHD6dog5Z8TNe+tno6W8EAB8Ys/nl5cTBdPC6inH+MRlMMmr
8Yy9K/7SY6iymAJ/8GHxpwo5FmWbjxSCu7oZC5J+JlUp2ccMktmK35VNezfGTVnDfZUdYJx8x+ar
1Hi7fKiXiwxP93DQYRdctsI0G3z0eiKavDCJns/Zz+3WAhrOoK1mOXU7+T4Mhy4N6HzbnczMLaqR
5rnibQTELusUVeSdNwk6T9Js0Bnn1+QXg3KOsyDroGABNfh2QeWDcZmGpZqvMxISNQ/p8iPm3XOC
iGU5WqP43L0nEdjQh0mVeCMx+AatYBAZkm4akE7xcpiVWy9GLzZTCnr65BKL+XFjx1YpNyI1h15h
kppBoxUxhzCx91+jhv8CeEV2Sc05T6uLA4GKvmR0Wr7Pch6u8v2bIM90/qPchTVnZ4xXTFFhvmEM
FsxGDy3urhJVZXzfcmGrQTTuT4iIqH1GPVfS7Or52peMVGXqOzNJMrZFVfr7fYfGYaBLyF6vpkJJ
emytSHpHUOsdOI+eTKMRPgt5nzmFEY/zj+v9PUdjU2tV1/kfJYrNPIJ853qeMG0T+BLZpaeOfxZ1
pyW9NmvTH837m9nnablPrng7/z2zMOqV1owau2IypuGvkyau3X271saMuIzWPrSHntnPgRxMwBkg
9DBwcqKkFP1B3apGsnnmEde76J9SwWffxCeV6ifl7kc8NDywsBS9nuULqUIv0hFg/voqdBK4/VWy
ZzPzNbqMStM1cAOFJhcfshxvBiyYYKChQ/aZLFfVUri92J8GKggq8W8J4AMwffWZcsF0BwDyxhEj
rA/jYRAWPXKO9B2AMA1TwqjpcJKSplvSESnGwto9klmkFVzZXUJAYNA8uPxdhEZXvCvAUOmxO5gj
9F+iSbCUg+ZJosUnasTnvvzswRXZ30N5skWlerRVq82PLjLcUzfmC4q/Fjpq9ie1IoF9tLlxPWZq
KWT9UJx6kpznXmARNTovX214B3MAzbgxq7UN2KxPpj4pT6gA9u2YF4gZ8AZ92c51T35Fur5WEQr/
ayQVL2HIMVyfYHF3b8ZPK1xgdK1BvWHZKqdgaykU5xoLdmDjFIPpoCxjH7lI6xLNQnlyGDRr2d1b
u5upsqyCRZtUd0r1Ha4wRmF7rStTNmjXbbFbjEI+yMlSbpc/bpYGOwuJ2gFCDbHZFG8lgnu3eLSy
B2qNY6gsLXH4j3MsIXxabEyyMxeIE/aNQYULrBZAhxFFzWNRM9UhcCewoB5srovY314uJbRj2gzA
o1rq2x7iUcEOiJwcZdRuYIYo4KD2tmlWlUg7B5zGms0PfKwfqfVyxfYP46DLW2IaIqgjUmNTusJF
ivHs5B4wnjBk3TF7BQ/LpUXtf8z1vVxFZdpZNkSQe9K+O5boVlPtvjLcCUGnz22auz8Rlwf6Vql2
JgB+DnBnT/ApKtaGn8w29ly87AOXGdUgMGZIUEkptaShIyzH8QS8hwQ69R2yGXZoom7+VQEeov87
b40hb+95qKH64dhiTJNuE46DnOpCboTohELZlfn3sA9a8+M72TAo3CbbACc/YraP7bcyQiypGaM8
oartPOq1odObLHyFUKAuHb3s6wrg2xTdSc3NbATQ3fb35PS6dNeXeEI23D41wiezHyRi8rTFhtf9
4ozMj6ejPd9/j+qR3hNlL6j7hKbZPTCczY1uo+kblimkEGeUTu82C2v6IZejQMBn6mXzpxi4jSqm
olhLH+gyKO+cmK5VQPp9TuKcRKMlZ21kFiQmKtLzBK1MoLbzMJJ4UWxhBBec3bnhKpfmEsuvhpUX
DjXyFguIdUcc7EQnsCFmF2YyEozrgUDLcsMi5nmvdqqKTQ/jNqkB6+w+i1JpiVRpeDkHY6/xnOJy
zyZtVb9F+5DCtAG9rb/nI21cb+NfKf9qE9a5/7rxXSw/Ym5CMBPLn+scDzaaHgxAOnMaYY776kVv
XYQO8OA6WSxvBNkIDcqy41wb2UjDSW3LvFqf+nGFPXLyk8g1Y7dFFhCQJSeoDlshXBCJoVwFBchr
Mj79l8iOPZf0XHCo11cVxnszhH6IOppxs8crBwW1avdEMUlyCzwtQRBz5f7gkClAnQPZGUTm7JX3
9YZ3t0bw2AB1YPtE9jKAjDoMGa/z+ELxp57Hlza7uGX35KHBJnU7Hr4cLmgFwUbB6C50bH30z7Np
9ufTw5k57Z9QTUIkvy51y9wCZVcEzZav1G20KTd6inlAHZbCRMHlIh/i9TtMoTmFtru+BS304AAv
8YEc4FPHonH7mKaiAkVJMiOu6wBPLRkPLe7RVHXRir568dt26xYwCFXYANu6okMF1QOE1IzXDIqO
OHZsf9TdQP54OX1v9nnX2J8YD6rKRtaBpRwGp+8nsnGxDtogAVilyjGnJuDrj3oAzswAYhNBJmsX
3Y90OTM89zZ8puMMh5N84LxA2vJz3f7CRtwLARt+F8/I/7bipy9FtoxQ8u9MNTqBfY4a2XnvFK5j
7AnHPDIrpP3Uoy+WhULTUCUQWPik2dFUcCoUlqIVAgVy+FnOIPokHeo52FVzsiH1VZmoJDuxrnS7
cT8FMpMpAbRx6rPMiupmqNySR5NiSbpcdV19bNIVe9Bnpty/7oObHUA11DCNpVesVfGY9TTQ/MPW
RE5/PnKxN4+VAlty4qwk+FOoIWU4qTvC0lDAIWFLPLoO9N8YER4QEFRuqZMXd2kKb+o3rnwV6y3I
f76wmAhxAqgK2feYr/k9a/Z/2PcfryiVbB4iueBfZ3gKFiqr3f9+2SQxi8TRW0AzQe+Igv60sCC5
zKnCKSaIYnUvdvnmEfuP3hCF8AHU3XFw0B4Vw8LswltieO17BIp9gKsSEyOJrnn7q2EyNc01Go1h
F6hvvNZ7Bm+bBVo5ubTcEk7jEiT6uwlmGBadPnIWnVJzSCknJs5nID/1YB1ywZSRrM6WQ0BfpY6V
VXNv8uZu3EYWxqDjtl71jqA4RP+y4Ln5cc9d1rstJI6q43u4HmKMb33ASV7KLl4sahNtivrsDpZv
uO5w/60KRcoJ5t2DuSLoheCy++K00+wmFXE5phnPMPShZnzdhWWoOALEPEzK/RiZz6WQhwAtPPPv
kZWZrTIuYtMtFHVw6VczHt7Ipmj7eArdDwMKHH5bu7amWO5faUh2uzEL2x4vx1rBM6Lre1yLKVyN
hhd+vSoWOW0AGhYI9uCIgowLrXAP3k0ixBd5+NFm3iqxE7oaiPr2u2faZfPlnmfy/o+KJV9qME+y
B0NTscYvtIhMm0Yz3g0/gNSa0bn5NCbdpk01ucyyBh0fXP88YmCWkK78o+tpEZUGRHzdkd6txamo
0bep9MciT88NMId75mJiqp+GlALJqALQi9SJQA0rnvMXt6jNRPjCMbJvOZbr1jOPMS4jd44ZDWXv
JgAtUdv9yRAVeGBj2/EX2zN8qY9UWaAjWSLPD+kFrLiJC7txt91e9Brw45uY0CxJAA8ZSAobOqAP
j3b2eDaedf2W8YD7sHZBUfXIJKfidHKEiujRKqA5+5GWnkNi7H8qOoHd1XC0XP+ywQvq9ErRilP3
BIE2hG0AMgxbZWKbW5gD/kUW5pr9rW20wnLb6FgLAIcsABh6IPgQ5r3KbFo012LiMhlq6RlAJ/Pt
OydWX7SLZP3kYYcwDOhda5X0oDj6CqAk16HflM/QKEb9KHvxz/nTe1l8d+JJZFunayVqRgKY4gHO
35MjPU99RwMQowGVKUUpFCjNo0moz8427tnNETGTZEWxOmg49y21Upk1YQnPizO8CeuQzfWCU69D
kuIjkGe/QLIBPdgBM1HUyqqpddGxwSDq8+0MdUcaWeVhTpmtcqxfJeuDKGk5Ga69qYmB91KOJQg9
lFojN42L8QfwUwJXaRRL5FmNUB1ihqbDqtMcGSmGbBwKlt1qzZ3uk9otnuc6hneNM7KC6G1OyHq/
a/nOnC5luYfOZchzN/A2YrsEE/ipXSVX24WU4xKVim9V/GpNhhciJGF4i2sMzJyPKWXS1sfMVDOK
Wln4lm7oQ2tgBO79J1SsC8hOL04Pw1XjVjl7ILd40M2MQVp/DwR7H7w3s/SDJh6Ym7wteXmLsgNf
DYjY1EbFZ8v8P6ILmnF/lzddWVjJEJr+CB9WgAmcWwZEAIXBYTYceXuP3mVcuVJfU6D+6oArMQW8
gdSNeSziZRMJrE4hZfAoatACtXo8JDXJSjm+tlV41FtQXAP6yw5OkaqtKOd3J27JWqj5kOsQDqfl
CbZmGEWWGWfbe8ENpvFQgYx8JD9Jp7RxPHwDOhYey+dOxyQEWp82pvREHHHl+rnuQ6fWt3DG8tVX
WI90DELCp5J9MF/VI294POEWK1EGEOjp4Geqb8zT2rdSLvp9xDlykswrDLYC6sotcZHeZkaCGrrV
DArbWlU8d8TCmgTpWIqK565ihSvcWagSAZ1tsX8Bz8cP1kJtcl3LfsYnpQMvZki0kpjduupBYdOK
NwT1lrdoiNE1xYoh2fzHP0aEDry5YwkUOcHviEXo6YTiY60driEfOnNkYEOPJUx1D9Y3biKrcX9x
JKKnnOnFygrNg3vGXUKDDibwD94Xu8aykrsSELBz/CDzO9M4qi/UDP5bcF4nyQ49MsxVs5SrxwlM
gWhm5EN65GaiQMxs7hnKefAcIoTVItbpng26bl+6+MstQ7bFuiwnYbzmG9sqLImqE1jafsrJB2nx
jIPwEHXotfcEooqu1f3XEoYG+WBIKNuKwnMaJ3gnI8FEtW0lbBtBIR6wQAqUdj3ayR8O4CinbeiA
4gxwfb3bKFu1TJO5UOXHXz8/JALcib2+MmJmh/YlHeyI+Ly6AP6McabQ2NlRlKwPS6EU63NF4m9o
SJjIVqmGiNujbeWNpg3ojc+rVzmJKZmoFoCpWHTJu5DotESzQYuL9EcZ6/bNwdvc97GHcMQm4BHy
/KrHfewEQwLpeH2wQjsvWAWKsXNKY36FIIQsVYfVpQruSmqEzyV0cipizZ63qFAqQCuNknrYpkbX
//wUdI/C+VaTm55I6YSIX1LRd3y4CG2ZkcmgDa2yFy6eES2uIZgHfMD4DXgbDLMB9xyLywdC/Qv/
M9RVsHqri55220QnVM9eDKjFbPCez/5ngrw7GqwB41SR7bAtPJ9/Rx4H4pTHFwJ/iaDr+SMJc6Gq
aU83VXk2u/Vk/mO/1kW7htBioWWWyXts/Xg3N2HT6Mqb4weTMQKHiHz9PKPTluL3UM2qosmJrlVq
QlSIu2KUJD4BxpdhEXieMmBl3GfIMVinmt1XGoy0gOKmxYnhJv8Me5CONUxgwHA4C62UFd6Fwuvu
TCC62N66aR4MnDOc10eaGBYqZYt32QxzEMIkyAVrPW8LqtqUmFmRCrnmfpZQfIiZKiopaexkFvaj
p7tC/G+u44MYzbpb/ovj+Rr4WBq67Qv3jt6BRP+4jvyNMAG6xxX6B64m32tUsU2FO2qK2XDvO9dJ
yMOEjDDXXb+WtOvV8UbOERqZJEE11tIyUTkUIyrcxsEgwCqBoHmc11s1QT50YaIX+3lb+ZzznoDj
LCZ2Et3GU2Q4Q1yWqT1T0SO6Vc6FxAiYHPCRfpeyWx1torxDejrAMsYizAf9KtwCTZWpNDnrlxTu
24tORgmpGXdUei3iKJw/5o0OnwBsjNxh7ioew5jntIWPKaO8WqQZlwDx6mAUfHJpG4PqxMinmom3
/t+OKDnHtQeFPqQ+TucAXygSjwNtbhpOvu1lKOyOma4Dxdi5RDLSb0Gniia7pd6BLS6B8iVhSVoc
kakK8DWsxBDPGfXzGw0QAl1uLnKO3vm7701kzRupwiGn2h6cJqKQGA2fztRn+pRxxJg3+9nakjDz
ZubsRPJzYmKUPc7dsd0zSJW3n4dy/7RpxnOTYjTdQslvf7GsqzctKCZ9qzltYF755rbTn3eWnQ/R
JquShl06c4XsWTA1FWY+bGSqSWb2xhsweWmZ82+mYy+ear7vWRWH2Z2RF63c09cG/4F4FAJgIalB
P1Z21ZTIbfX+yJlcjznnwflMgv3S4flg+/qnxzyMgqCZAU7UQ6OGeEKnNvMEdlhPT5DFYC18O9zU
zo52+iNVxKzNc5gjOgAbfZi9JIefy9VGB+5/kpvDzBdnLoYbI8649CbLGk/PTyGiwNCNYnMcgeip
hF+bSvy2jtpBKb8xFWvs3VjBrzfQBX0qaURJUhis+ngALs7JpzGXIqZx5hSMBKXeTMP7mpfhGlLD
wOkuwUYYT1fcUranJRqf8NcrnIXklAm/8b/c3Wfc/MEy+ZJx1jNrby+nSCTBwHMP29xeYQWlUVEp
zIpgsuwBcWlFTUWsQYksj1lFPjWLZjzfk5Rve2ysREitGMzamLwrDCG+xJPl6mu3mkUSHP7IFyhp
2yubORaM55E2nQ1bG5qStUWZnWHq9pwMCfkWghkkhKb1JdHkTMrz9o4O/yPn+wV00ttsbNLipFGp
1Lp8OdF+pgYqf5SWZ4sm2zKx/8cbekvgmP5d8lNdPV6LMS4PVAMwRAG+uxAJYf3A1oSBG4i4qoTl
mKVJTXjspXGPnvFk2GVvgKeyhPviq6Ucm9P9glOqInxslYuXwCLaazolHa1f5Ubmhu8yKJ/E3tB5
KWgnwzC+mYTul6vxUhJyTjO3sIwK46e5owFkHKqgY+ez0ubtANU9pqimJNMmshvvO3h3rVsO3oRZ
5u+stfxlnZUyjF8FzmSkZGD6mpgVF83xkFk5aQHaL0ekbOy2uKn7eaNhEKlDno8U6Nk7ENlt7u/V
jokYdLTwoA0kZClXAzZCUBHulZVNVgH695wO+jpRKLlzOU0iM3/ejWqpb0dsgAr/Cu22/W9Vbw0V
KRLZjhi2vjJrPNlodr+/Z7CfuSPKf3mabbqRzmqA6lYd15gHp8uuu5M7QaZQF6paJ6dCk5xrPpeN
QE7RcCoBxHU4VMqU7ZD5nyEBO8gLrMn8UPF9mHaJkr2JC2t8Rno5z76AoUMhd8aVqWTTUDiuqnUP
zXLYvXY5uiPRo0AmZklzMd/GYIhm+EuN7ToiJ8YcnDLLq6w1JH0DdxFxyVHrm88yEQs6nbkpqOAA
+OX5C8DoCYkWi8/GVvsloWnn7uP8PraMt+T/WrPLFfLd2KYOPXJtdKUU7MUWbqUnLT4zOdXWFCqw
1kXIQmRJQ5QgNB0OeoqiZ4bcKRxF6R+N2DXK9Vf1CF4msfuqkvITuDvw/cBEAq0//6KOYL+ry7V+
Yx1vCOMgFlwyTnd3Sxma8SQR5ajLGV54uUrafIl+0raHUZiTvZac7RazEjbMLmQK1bvQPkW0BH8f
K0L5koFLspBPIDILLaQDkWUhhW/bsWGc4IvvBL4en/kBTuOd9FCKsIh/tkoPJC9OIzFVv/MGK8S0
jPYNbcrAPJHD0ICqOKouKyjIOvGM4k0Uvd5cF23WglMRFSZIOg2yFHUT1oCamJQvQJ+77EFygVq/
Ex+Z/9LbLd5jftvkZ8YaWlfXl6B0n41RtRN0qG0u1XVlPIbFpfsQ59RlmIOw7Si6/iu8jtSoZdUv
WahCxvn5a7C+JWODq/gxVF3GQhj4HZ/l37ybhSOeMKaya5NsXHz7kFwWRR7lB1IANK/N85F/ZKBQ
IxpyMCb6QmGncYfPkee7DTlPaG+OMFETqy6xj48t9kHCWQZmqHPAsXLcfTwb2lkFSgvcsyDlO9Jm
paN5AOWmGBYXTlZdWcnW1v7PvB8RgOFeg4WtTXyGyIDNJg579sDVfp9aua7ZWb/meArRxWFo6JSi
Xmp/MeGYZQs0jA9H022579oUwAP1i2a2+A/+5/YSfZZdwudYPvKF5Qous41PGaHPzD9L7Xdw1os+
nBFo7grAjPo6XOJ+kyoDZP5t+lJVOz0ZnJ8NFtFEdNgY+myvgAlZl2neSYaZzifWmrk8inungBKO
yo6MkpiBLNr1J3boZmyhriJb1vnN+bFMmyde7Qkh/mHZXYITDZ3MPG/YCkVPkmkOc16UNr21H0ke
cMakHWzaw2nt2X/gPWX7Jbbj2UQv+Isn4MjHkYMp1kKxsJAz0p/8Kqz/4Bj3Masn/uRjEUqGr4fy
ejOklOZueunZz+z1Ptm440Qw4R6BtcjWlGcVcnVckG68bcZQ/Kq1ZRxZGOfnww+9Jren7raRfJWz
NudCAfzfq0ZiQ3nIsQVHDInxVrJTHgIZoHuDA15JsZXCaC9lY6s/GfZK+AbNmcjfH5YT7LEVqRL0
kNkOojgxivOVt06s6ylN2IhbQgiRYZ8WdcgMurMeHqTFS2/i6DaMy4EsUmtXKi/qrA222EVDqryd
xH6BZpqztldw/VAFLkNZ3t33UQg3ATiqP5Tdp9QoSDJRkg8yWDX6SFAv9dfK3BOfoetRxuQxuxA8
7F28rV09Vo4dkueiJxFEapfVtfGf63jlxtEMgA7aJz7T8dGf4MYvfXBdcrr2BC8b882AdMi4I/IQ
nQBcSP/aosUu5/heCn5ymq5/ICLJORNwDxEQ48yTePHjZJjZAu2U4ibfVmXwUethIW8b8z/8M5nG
/VDYxUHf5f92oIawROiaIGkd2K3tmanXkNSDTwRtlKBhb/CgJlwveWHrIlAad5RkUQGuAlGRs2Ay
hP9W6N+MA/R+QS2nIG9OPBlHMY0nI4NweWcgZBzFOqgGVCzrUirSRs13LRxCE3WXV45ebP1vSaaQ
I0n33YcnSmDYSNZCVjyyMAkKrV4fYUDgd6MHk82rP/qc7h24vKMy0SWHfvhZx4hPdH777dnM5X1M
HEFNTRxGC0nJ6GicRzbsQ2Mt/Qg5tkkC+4wDiA3AYIXm0o7XHY2CwRx/Le8jXzsuI2SBlwBUdgSt
7lQQx3i+A+OP7Kw19mBMmKBsRKLndSY9sbr6dGyUdcd7vkNiQFSmtzEMST2e9zDNooV6+yS7iUE1
Rcr5qu+1i1uE71QPGnhk919DJt7pbRwxmonUkENZp/IpuF90AVyTGWVxqQgMzGQmHx1JlKn84Dvi
IGFneER/Z3PdSENJd37xL36o1feGvenJUKyNs6NML7XPzsEvw5nIS0NlmWVxsprusnysaFf90EP0
3fo16mVTgKZpQf/nJ+oTPfMMDdgVK9pcM9ts8prC+w3t1bepcoKFlc4HSS4xKAbeVci6+456nNdn
HohUdjDPFWEodPkxbrwzBrEoNQqncV94XlOKDYM0jCQSjI+TQKY1hGVYwn9vKppKMw4KTS+JBLt/
RFjDGedESOugd8wLPyVrTLEDzxlkLOMDR5unwdDoiA0C0pNB1FvUWZ/1g5R22eFww69NGejKG058
n5Cbgeul9dsS39+xo8MDboBWaAcFqP7K2A0CVJs8myxbpXf2vF5/S7fd25dKmIzAC97hhb2MbyJL
ISZutzQRJH3GCXuUxmcDaAwgUwjIuPv7TdhuV9Qn9K/zyFIQ1KXg3lEHz9gKwQDHmB54G4RE/u5c
/44tFDCgdw8SADXdbC/FoLO7BAP4lA+z9ZT2Ez1RY2s2ksrUlWECTxr5Z+88PSw4xckN3w8ygVqY
ze4rLhCXDe6QD6EejRXmuOsim0T5D3gbuy4dTAzmcn8blP/5GQ5ReVcdTtdGPzFNltfFs53/1T3V
XF0bOJ2g7iO9nI8tu/HsGQKIFCoMsKshnyGi/5IcK7FrQ+pD8oNwRetqmYMuCAUltrF40rrdTCg5
NBCyoUL/LKdehh+ftnKIB5l1jjHpTHYvL0T1Em7Y+oOT3B7u7A2XbLzj2M0pqgGDFsvaF6WfvyLY
bF/3WJOFmBC7o9izIDFGsaAylA9wkYYtFhrrxflwlj6LtsIA/3VpZc9tC4dvRbttA3+q/hLBk8km
mjEcLEBYUJDKwlycKxtk3pT2NWXlzpjbHUKFKANEa9DlGpf+RfMcDwnYNyPs5LyEx41BnZPuDK0M
DkyY5h2QQn1QUrzMZrWm1fE/ZnJpRboDYqeXMc2+zxup9Z/If+GU7AlGXlQtDUPl8wVGRrHuJ8Pw
TvgjdBk5OtSGkQNJIh7TdzHJWi4fVCjvOKvSB9BcqIv3ImaJMAdwh24UVXr4h6yUA2aCP6TuxTsA
ZBIubJDnnL0vz3MZud2Wh+0BNbCt7XThws1f9gOZR3MTgHYJTXqUU9vHRuXwa3IgVEE49k+i6Z0s
GCZgJVvbV+hYN0SuUmx72tQpuut5fjqQQf/2n/9eWppjGaynxF3rmpTK1H0rXW75ptU00SGZeL7B
xo0u99s/ssBUadVPOO0wDRg/JE1NJreliCwcZepcQKEDemFLXIZXP0OkliLZLXK5UtTT3ciOG7bD
TFFipaOR0sIwh3Ql5r00GQ7d08b1pEvD+cIsRd1hBulLd7JTKr+KLLUP6F8vGyPSkia5vjHkW4h5
ttwyoDLWqY2qjsmm66N9yvm3yb9bVbhV0aYaVfILtE/9cr1+CC5AgeRmDUF+YreW+X4Sep53KPxp
zk3CCFV3EJqhg6tybPtxRrGJf+flZTs89Ndgguyi7eykrn4NSFYvovQovA9UopKY2D1mYCyEE9rf
jVHRUCU/aUQM0t6CUAOEn8NeKRY1c4XWI7kTPBwlrN76MKG3ceAR2MBsFcUwQqt31Eo6IxM8ymug
Mf6IAv6Q+MWkRizU1g9SV2b7wawFijpLHCSvodyBsMOKqQeP/V9Sa7ka87tGgcqVZfn+poFZvIvs
SnWHRzbWZ4YhEsdOBjNyoR6od3ox8x+K38BZ4DxggLW/JHkdk9NtosWKubuoMUjOWtRzDgwNTP3/
SIJyCxjRl3Q10celVHUmkFNVc7QPaQ4oiOv63AuocHi37DQQlJex0jClAQPVLhaFF7e6N+hGBO4G
6nIxeeOsySSVrmiByIp+4GREUAL4O8oMKh4AMNMRI2l5nmeA9MjSuYBu30U+tA7AHzDD8qRbydAc
9Z28P8JomPRnw9MqOiE+EWBvab91ed+p4wX/dWqOhiWQ8/JxTSh8lLl/GwsotJ6oeDlGsV2xCih1
CWfavOPMocHt1j3C4J8e62DJOzoUR2n+CLYzj+s9kEIUc/yUWIIAAVVGVWgieB7NZMmt87HqxhXU
fjqrCp5BkD13RlKsiNM6GQwyPF1XcqfT+PAuPcrC34IGlEWRwhpGILF5Ftk6mb/NszQiy/mh9/JJ
VR0iph/wIBXiafS/p9RBVb+7uQMrBQFY2ug+lxokuKx/8s2utiVKAzGq/r7vWUhw7E/dYCh/P8q7
aCzcaJcXkNNLjRLsA6dpc2sLtmcrJwppnPih/xvFXtNLYJ0kIVnztjALARN97PpSDhEiM5EPUJy7
FLHI0u/1b9VGl3u1DEMF+PHfUQcQ8CFkLG1zq/Omb/uqNK7HxH8Gf1RgRPyVSOJXMOJpcDLtBSjn
XRAfJ/8W6l/GlOUDAo/MwooW4EkuV+HQq6ngY/PHAX/ZzyiF89/Ieg6lY43Pb/2F9lfj26RKCql2
KM4WJCCOVih77QhLN/B8C/OXCHbLDcwdsbGX7H67kM2FHbmJvB9m+gQudQJKeY/KG045ySEj4jsv
gLML6rjHcy0IC4b38ad34CUWobiOZVDV63EfKb3P8WlyQWf9g+AnM+A+kqpzXzu6Ulrcu4+QAxJa
teU7nrgNil5jtHwG5xJe5/BlsadnmUCRoaFspC2CVDK1ItCUpj0W0dp9yAoKYlCjLrTlQBaMKg+G
GGFtIV+ErKEbWRgzYuhxCTGl06bHYtK7jDAy7TUNJfskdvDTn7d5M+F62RBY71LWMplJeC+4ZnxI
vTjg9Yr50fwKj/dEkcD5+W51R+mvJd0sHLmyOyYnAmlXs0YJHYFHEmOVUrIQEA41CEd3+aKsCROD
zVdEm+QFr8FgK245Cireno65Z0KPjaLD1ZGtgh74bMULtrKPj8kFenCBHJ8Bb93tOLQtgfDdOxPw
cydReZG/kFHbM3ACYVcXqwy3g0thNdINYjNLwNFU5yCgMEG6aSU7ZsMWvlf3V3FuX+NQMYh1QhXk
WdHP0DzG7daY4vcttUSDuk6oj+ycyoZSUgO28kITdeSYtSPrvKck/ZGRUPTaui0hwLCgOt/As5ey
LWiVjNy1GatHKQLM5u3Z+uc6Vm+egIiLpfHf8FDJrXxf1fNFD0rac7E+osAXs1O5716Cf3AceHdT
CoPsdqsxSLac2fYwnyN/358bq8ct0PM0kOKssRH/8izB94ge4fDj5f+WAnLCaUz9Qwu+tFH33dUR
DFE4I7lvHTeXQHIb/65dQsZ+f0sGSq9clsDAzJsHF+mQNxnx3Zp0w+lrA3ns+dznCaFiFJ8QESzz
e4wM8yr0bQulExiZ5layNzo8IwT8NZGdZcJlR0rj0MW1sPcb0Nn5fn68zDwcC3bKbNeEkIfGlU8u
3FZLGtcQOZ6uo85PPvI8nxg0zqiIggTHmWRC8cndo4pu8brVAtWbkEliEaQN92te4iJFOfRbqHGS
ShuEerz4pzq06gSexdah4NUGYjRRAs8wEyQwjsTCyVT6vHAEkiK3X5dTtGMzC86YhEHHPifZEJYM
Zr4879OwTFBqdzrAzEcMhZgOHtWyN5+xzzja2iV2G0EoiI7E+/2YhuUlPuZkCMfmtYX11ZQVjTDJ
gkamviP0vWf27gS209KT860rdiwOR5ip8cLXLJTtZbRUSY/Ze0Q1soWt2vueJDci87A449dvxDy6
GuBhAlitm+IHDNUc9BzmwRVkd3NqftmQaLujJXVMVKGBBs1n1mzMSFTvVSsz3JaoD2d8akb4z/Cn
jLfUqjmEXkdFZl0DjslrmnxYsptxHlhur63jAiK7H/rhrsPoP0NeizDXP8jWIwVwyCYDWCvdpwLc
bM1qnGfF8U2wn38dZmn6Ftftmc0lSGuk2fcD0S4u8qxF7f7zTPkoN6U8BaTQNMQ6/0HEDlsItY6L
udOdFJoPqekV+LsL2UnI5f3WET8typui4IP4x/dHjzj4JCclez089qbs/WDm5QRk/sSI2XyH9NBW
YBUNbJjIQwahvUB3Hzv9H455wUvGFlFIoBQz72Uz+t6f9ZEIkgtii84ZZh2kY/6DqzpKpub0mOMU
LnrZCuBac8gfN1ScC3orYgl6ydT6pt7ZjxTWSr2lSJkJJRyy+QaPKJST9QpZClC08wv7t6Io9Y7l
+sNYy7Tq1/l6WPyWI7DchplR4UIy5TkU6ycOWg8QnGBCJ40lRTrQ6AhwMeNoGdw0pCsSOf/wjdEa
1i2ri7SiybmbggHdAoQ9xNyQsox36QrznjAzwrnHSSLeOht0P2qu+wXLP2qhSGq7hXL3GYMiJsHE
bEXCPDOnXPiLPs8WXsNG/286RpKJdqpqaLLbs9nlxenC/1KuxYXyVp2NAAf4asVodJKNBfAwsOsg
oZWuiU47ACd1uQQTZLLMBoHkIIVam8YwQYawBlplETnWtZMUwbOuaDY0u2kdjiKgNyBovVgIj3g0
rqKKW0TZjb7fMIK3XbUROUoGUlB5z0ERumVkUc3KfqxtcbrCOv/1+NJVo6PMbIX5noQBKiyDqlFl
QzSL0b51/2IjcOuMahyLSEU7/oYxmpVYLRx0fO5G5+NzyLUcMQ9OSizenMuI2rmxAYaPq+XLmWjN
Xi3VhwsInCmYtEwJukk2TYt7wuu9lKGAuPCvV7tva3qUfkoi3RMAAtz87QwJctn+HPKaWJ9r/ySw
yvgDcBr3Ixs363a2+GZG3uGB0LNvdSbon4AjIPxtXwHNrOdG3iV+4PIu/fSQepdHVcljY2wyWyEE
Ah/mD1HoODfdOn4L9+joefYee1B26bmCpiw3t43dLmNWmztnxO0dwQkbaY6LfLvLi0/e0bVJvwIg
VEu3aR3PDMFpYBWVK8lkNH4d6CmAFUWGbVank/og3opHwwkTfsKvwxKNV/xgLzkZUo7nOPlrJSan
Tc3MzX9gC2tigUX+2D9CF7f3V7hQ5P7Ufv3Tps4dgdehOkj5kbtnJ5QzFV+/ArTSZYPMPBkSBJMi
6UDismMwq+e7FEPDfCVkJUbO9gdShVcCHiHF5LKCTrpU1f4YW2yKpTxq0JgFLjnF3pI9+5z0z8xd
78UypmHddZC7q1+ShLnZJsdp+WrzifSd2JJ2Y5wSgmWa2iAPIG3r2RJll4yYLRbld4MqQJkYGXpV
cxlWqu/KxGK4okL9wdCOQ+p1EJrwQYzTOVVfRjGOT3tMUl1Pkz7cAN5JycZhWrKJmaF8GsXXsZ5U
nW47RIavvUQsHCNNOQcFBBc+n2yAiqAdQQpNjKZiKnOmYn3X0y/aF69H7d8F4DenyaoEQbooM9yQ
ZziSAwg0wB10p4TB3Skkf4TUNKCsgsWe7UnbGZldKvWIroML+6MrRj/1VvrkyNdmXm0t2w5RaW2W
nUG4uo07LAF2Rq8M6KIp+VKB82IKZmjPx1V8lQIpwfn1yAR7+mawSHwmywfRrUiqNg6+/zR/svER
y5B7s2GXCh8Y+XHfGArpG39+HgFnSqNRh8vvQt7XMp4NKw++h5adG0kGBIL1Wd+F4/c2gGUy+AeO
u+RJel/m/aUofVXlXPsD3/HriBuU7UfuyhooSOwZ7LCE1O5XFt2OOrgQHM7RJPFQdhGVDKb239ZL
y+AdQ77dtRD/aSCLaJiw0veHcyhX9OR2V3J5S6ri2FjrAfy/M7/29RO6lNKuQM0UKgPeB6FfnuzS
Bsz7OT38j84afGP0GA3g1D06GotroxpesYBx962o7LKYrH5gB1cf1Ssr5F8YehPts0TU+wgRFn9a
a4zg9EzB6IAgWkhZEehSst7G3b5Q/cwURB6q6xTQe2oVfAdi0OoAhG8cIkBXLgy5vJCZOX1bXarC
W3UHAq59g7+jlqu3bHd2Kq9sx+LxesJD9U3OZFYoYJET0xeXQaZ2EGWsXl+6fC3ZW79J6WqxKse8
Lgl8Bz9CYIi25tmCuEXCZXOK7VXFFlSFk4ZPOjyP6V2is3xvGMAiIuZq/GLe8LJrbgdQrE/Q8Ckc
597kbGJxstqe7TyDlbhskEPeT2c5xk8gslGj+ZrUvq6gZa6X6jONzwooLVBe7l98xSu14t1bM0vj
Bj4JY6OLMQjY+vWGTTTAOfNQQz2MQ3PoTIOolx78Tokkx7N9E5RInLd5+y/8KxfLreE4jcrnvtgu
L8rTemDR+cnoSYbQ4vF3On+c2iJrwZRfTBfei5C5tKx7JhyWJcWH4O+re7MLydbiktsz0ePnGPMe
LGTksgAbQqZUvqwN6nHMG6b8C9mPURbSDhHOO7PIa/TGRzbT7lu5tHCAG3iJ3w1WONn0PSLZrOzt
yysTwSSxxzVQtRJre5XO4d/7tB/FfSup6fh0RJysPYpOBLX5L1tb0B36WVvbxqfZgS5uujBdxl+X
dPD3y344eFoMhWqdl8IjOy9O3U9U0Ira0wTqnHnQj5tcqr/1OP8B8wsQ6PX4YN1OC26gSHk+YVD5
zLwJlLIvusvOXiC4f7S0CaHYjGmB3Hg/mxfL/7gmHSE9ENPotKT0J94oceDtDmZKyRxd3EYJNxxA
3llHVmyCAXPqjNTwPppd0NhIWARHHVG3iP71z2xwNvwQUrwgsLBS1PBOD6+AHhZ9TGhwYpy1zDoZ
8vBJt6b9VOvDq1jLlQg/XJ50+RatZEkwujmQRb9bz/zpHkJ/HDlgAzq+AG6Hp0WQrE2Ta7hTcFjO
zRw0bHqTR08ZVYZFecAEIVR7f4D9UBQgm9hWIaeYSJUMzgqcvyCh8n/FS8c9yUyRGbsSynsU1gp/
vebAAPBZsLdmNJc+9H+PsI+UYe5A0V/k+bKce2DoHgIqFRvbaghnIaRN4OytpbvopYE7bKCZcWKy
lFKsB34OUD09g+oQTUBPLCyqiArvQLWfDSnKkEMunIsi696HzUfl3oQ0q1OiZrJ4yeUH3l2mhh8y
tdpsgWl7I72OTbm1+Mh7kRP0bunxiPQhTFi1FieRyx2CVQnKpK/6Lmy6eNm+Yu6Uyw/Oe0+8NETf
u/GYzLooe/d7R1NExEIIdAmyMV3Zc1t8zAhPOvhp1iHQEMKkfps2mIQGmlf9chhmv8AwOaxNX9hf
BzNSs7CfPGvP9BR/ar/vTXnhPNjannzIKjZOlcMxJdmlUf6ngx6cHQDsp3uci0sB+aDEbUBp9IJm
cleFsqYUnghJiNbDxMg8horb/UB00Bqd8QlMt+P9fKorc/2P5hEkMrr+ieZJArBljc8WvZIFAavm
z6kqq3l8QOxp8e2F6z6FPtGPuSdLDs0Xbk1qyubEgVnt6PqkL4NcWTKDWVCx1WgojuCNFIG+NeKx
evDq8OeO3lR5HzG33PnJ1MA/4nxY6q4dxzAwQt3ywN/qi08sgNVE9xul5o16zNpyDXMvn+Y3VWjO
1qAuQd87XvWomD0l06O9kFxDas6NCW81/a5Ax2OKFubDQwrcwoADJPhuJ9EjAsYikP1HeLSxoPNX
pPo0lutkHAOY8439NYc0W5ncsk4rAxjX3+4gL+8+HFLi7fJOku5vj4BM7uvWWX/a+1wjXDFO8E87
QqYYL6ULjeJ0SCjn/muQUAOMcJl127F+42GXbsSLNWJ0XlqunQb56Ov6dGekCqyCSJFVhr5Yzu04
6t7Ca0jNaZSBSkaNLNt2VzERXBrx9wG15qX6jFnzhYrmduIPbkYqEP6V9WYY3LLfX08HsUUZM8KP
mAS6sxC9HCCMI2laJ8jFjY0Xdqs0SJJZRcU8PfYYHvsZ/8gwiK48jzGNUQlNObPcu2Y/abh6LFZO
PtXrlweuFMv4tm1GHUYPkrNjzPD5ZMYZPWA2JIEERnCahxY08VKnl8Ai6RVc9QYU0HkioTBRiCd5
sSQTAiQjUAf+i5Yk3EQpCKl6qCl0Vb8isEmq0kNDAfRWNr3++zNHR2v58rIKvviHVpZ/CmFh8eMC
a0CnrtIOsPZEwlBOvsLCBwAiZs35/vw66mDOHvkbwUm8KE97SZKlSENK0daAa0k2621Bb3biHZTG
guS4VbIA1d53bwpyofYWKQ4V2u8hAwE50StpSPiurSSsCt8T/wTwAzx2oSjt0N+eJ9dVE2gfwLX1
OShsnPigwO305XUiC5uky2pvZuBdKl08bR204SOhcr1JPC6tSzv/yvRdu6azS8+X+nobKud7uEwI
1uphlhMSErkJAxkcWiazIztgyXJFDJN3zMg12SklTSIUUTAOdve0qG3rr7oE3tx4U4INJVKCDUrw
jjlCUZTt6IO8btMKbwvxhovfNnPyNG5IDRX2Oe+U9sQDy2PmpoMpcOHhS+jjnkQs79AZKtTlIeCD
DUOfhXjeBpymlLXgo6HZF74Jdq9IRieE+5WG7Gi+XwCHSstjL1I9o9ObjIPJtWY/QS50x0lOtEvs
ElRx87wx2apgiPbkDYaJ26tBaazbPQqFK2exmaaIyizoluFx4qORXLZB0c9MFfw1gdpFgjD/GfFN
UTnWynmBrQGg4htbVA7XmFiOnBs612HyPlNJuyqq2GaDf1dkOeFT6R2y2JTnZ843EWZhc2Jl9qXb
3NOdlKWAakuI+OBk0g43+tAYcJxKk7Zkm67t9mkWE10wwCIuU82oHwr4hKXeVVz0Qg20Ebx07XyX
nnd4Fwks4nQJDRtwMq5NsW9CRoAKc8HZYMnGx6xkf06k2eYyfPr9DLMrHieSq8vea6JqLO5I62u2
+wHRzuqam5ixPv6HX9Q/VMbgaT1Ib5uTf0IpAk0qDd9vQ6zazXL9DeARjKP2yND0NzdKKU0wxOCc
Z1wQ8dZQdN48EMjLU/DA2gi0x6faUmdzVEX83RTn20XFHZXias5+dRqpICluzbfd/ssF3qPb8G5U
+QLasBU2ieM+dqtWJCQd2Uvmye8CHjBKGHwt2Y55I19gB5zMiCHGA4Rjtj2YDpR5dXPRJqAJTte2
JIPbjzK9+7YTgay2VSvL819stWB0UzSuUXKU9pl+twsUHaP1lNENADqa/o9J/R3Cnl2UXPV05Chx
UttGgNjBfbNF5UkD5ZidgC3UCxuxqCmoAFp8G7T0GKP6P7tTcaPKZjqpFxwrBQH44oYAGpWDpOEj
bpWnzZJj4XLA2wzMDGghsQdOK/3NKNNRcO7qgYnsHjMQJKOqQ1su8AYyN6az0D4uZSzpOMr8CiNw
L0KmDFLeXE+9k8rp/XCkMW6DdUvrq9acPvWK8vnBarv9UT1KkRf5etcM5Pf/uMSqOhJsHNtPQr9k
RrbWs4zLrtW+h0F+Co14XvVFdLWhd/On5g3zYE+GwWB6krLQOqakp2bBOtYo/2NCK2Yk7GVewcEj
sfXMS20SNPuAQ5LgRUdpLrcDoJ/IpwEb5GN4HjPo9kGxoAlBBDiL6y6V1z3w1pVYG8d+EMy/WOIm
K1XMGbbhl1eqUAxfzjC1360nixyvNGTpgfRFOpYJWzMr4Gii/bczFrAsHObAuUrfIcBY7tp/V7/U
EV+BXk2ZvK0MjS83I3cnmdFpw+dIXJM9Oie7nGNCgtJ963iCJMUHyfRe2Zwsq6yqPJ2EG15anmB1
JfXdaHTiKpZqWPd+E2ROCGdmPzUmyytrjL7YEArv4qZoosjylXJSE98ce9ESHA/2NUZyBrValC3M
aHVMrLw3l3JnPsTHKklgi1TJ7KWKxfkTytpcCVFfNJ/X8KEYIDSUN4O4KVHKsuxqyBIn8ln3PH9y
A0yHPlNZGG21p2t66wllLVR6u2r3a5IjANIprS7oR+taVYhVXSC1U/j3xQ1bf/MwfM1XDiXMwlHy
bcTBG2fotust+mzchtQk2x11VJLzkzKPJ0xfj+SvRNNmrJo5WecsUU4PwGJdvSPZ1Tet5P+xbjpB
eYmjRRI0f7twjJhvqWnYZQgM8UHCukssTH2MpExX3LBIFaNixYfHXQIIqc51oL/9OHDPVmYx73cW
bvLxjVHM3DtYTb0TQAQej6p0k+BZIk4Sc6ZwJ7fZSz/lmdyKYzBq67TvR/NKZjBGz16l8yJv86FX
ZnN86+B/JtoBxYBE6vXadRtWDeaMsNmqE/2Oze5T936Wvi7Gk3GQ+wHzTzZHNxhpZnMrndeXLm/1
tXbwjjFE4LdwSQ/+jWkXZE99d0ffW9CbTkB7fwrX9MKo+H7qSbUyP5C2YexQzEQSouRVdI5yGD74
O+PkrUbjJehTxjKroeppOw9d4SgwuwHggqN76C9jWfQQa/L3YkRo26NJOg4qE+RCsg/D+HUK762a
B+tVnDjU4bO1Xts5iZ7tqJ7SPPTQ1zt+FrnGTeYmaIS25t37w2+Dp5O+JZUKlLoLT7f6ToMKdvem
TCpOG8DOKGakQUqQHdIkXg+geNVszSi7pQ9sZGm9u0Oo+Fe6E4O1I6/QjXKSChFn2uyJK1WNMTDc
Au4ss8dlFiwAhSdBMdNAp7Fh2p5LgcwdGev8XHWt9v/pi1GmL+EKS8yieuVKPDHen/cCLH83Of4N
uDkC4ZD8E4DXIwDYqzCwPAllZEEcjLVbbTY0bJyMiudtC988zKX/t/9QR1A0TDYhMErE2n3Kq/Dy
Rr9eV54DFfK2pdMrsLYRDmSE3qz4ZFuz2wlV4+cjAQMJD3RqcOYrH9P+jAeG7uqQdLlsivJq7PGw
Rj3MFHH86e3cDaDrGWu5+K8kRp2WsdvpJKcxiR3WWAfc6gSUigE3+kqb8t4pl3KXLRc2dzsPDGDD
Hoo2pyzIRZb2GeBGOsp6ek+cBLh7Lh9JJXB0srp+nZ8OjfFFvuvojb6HrXymuoHJavykU8XkDtxV
HSSuNDFJ5mpc/CL792jCVGmr2qm1ERHbNuvw0owslvYIM7kS/GofTHuTYNm9Ij8FhvpZGY12Y3Al
yh1ZkLPb+IOG7bx7xjk6m1SxDuYBHKouwqWM3p/4bAujT0qu+gz291cuqIwRZrtxiQHBgaNK6C/N
f1mMkdKvPwZuJyyvsjMHL+L5eDQr+5bKYVh+OkHQ2a74eo/8LrV5/sA+LbPzAGP51CFcwNPpjVJP
fVk+Zmz4dQqqI6c/0lZUrUyCdsREzyrDjG0/RWvDLN0Q9R0xSO0gTxrM0a0i0VUy168B07HDypbR
GUG/MXbN+YDkRI9+DPxfPaeP4UzfGPhBouVR+NJ+r3z2EpPkzpdsb17qtEGhFTrHkNVsJ1ufAfoR
vPjdNLO3Y2IqJWQSC3FnHruLWtrNZRLiTVxGCgaG+IDbnqQ+v48xUYrQ/iM1TYvGNlbc9QT2WxQO
vfEoO/I/KPSW9TQbF6VQ3RAxaJ8yPyq7RSZHFHu5gTBEUecLi1vT9RBDQZPTONpk01qe5T1F0TgP
/enzacvmSvFskSxSvtMWs12it0UZ5pG0/X8e1Z4KeA/tkBziEwduetA5xyR7BdT183LMG6sZQ7Ub
6ZJar/P5v/1eVW8E49RyhMt/kVDpikad1pio3Tfq+QzQcasjzwnRZiX0ndwu6fDoudIt5XWMTPvQ
dTNlsgVaABpAemCOJ8mOgTyeB0HFViKCuEzoz4TEpNK8GUftbYE1tzuHRqB2/ddvXTEOu5nD3AFx
K7mW2YtUjaz+yHLpJ2J6Mh7q3Ewdwdc6CBjTH1QQKMxEyn1uqRURBuiQIribtuGB8T2YOgWbOspv
gl4Nt4LSKCPfdB5T8KCTZYfoO3nDnbeQfqsEua5dxN5WANf8e3rEOwgBCWa2b2hLGDHbwOoD2A8Y
AOE9dzBSsZjNYHXA4tX5azw+X41ekWOPvNeaHOSCkkalIQeOXixk3FDtCKB+91imFn6cHSDMfGL0
tZ4ZhdjZO+AEFc3hEgobG9rakJTY3HQ+JhJ41Lsgt1RrMhZMv2OOMxTngNMprO2aLlj0mooF4Zhd
8R9erKupEC4KDogZmNUqoRuhLDsbT9lo64GukgfWEOLxVCExkwobp3sIkaBGxO8uP1G+E726xlAG
BzEYMb4UPBb5BWplKAxHvBXOv5aoGChxPCjg/oEGLVGHSftpcf/5uGo26Kih9ennb1fTKSFdk/Ol
arC45UKGSWGYLpn/OXGluorOp5aJra0hybEKC7Pp/OyQnraV5jOAlzvO21FPBHRWsweCIe92F78S
flmBXrgG6HqsvsofVFukP5MWf5igXT2t2NHW7EilkABvtPEW7sEp94COPV/e7OPdJmBpTaYJEkpk
PMnVEZDwSu8vpAQ2bWsR5UBofbslOpyx3bpNSzU3r+ogeE6otv3hs6riyYHATGLmzngy9zstjBHn
kxL1fASLHzMPbd7w6u+HK+EqHQWDFvyWudEXdfCGZR7rpHPeGoL6r1AEji+3jjBULLl311Ru/XxZ
rJ7/09Ya8FRrIsxsYfFOPTzRb1jwd7RhfP1FxfyMN4IelmUIyhyFIfMBKjr9SeHC9YS6A8iQaHko
VFGVmtaThcHcTqiJC/Gd1d1044sU5/0pcgqZ7qOUnU7RqXlBg+MWkdrLRra11BKFPa36Ys7Pr6/H
pcFQGrymplYhJmMnwCwnGUUJ7+fmUT0hiZSeofti3/c4IjXOyNz96oM0EYsw2o19zMz/3H5DCVAa
gSglJ3ZbFIvDeS88OCzqNrnI5A70n3AwuZtDmb0xl5YdUoYF4Ri5LyCpKFybt3jm+oCWZdyUQQOx
E64XSAHUPsbWA8ipLT5W+npLS0p5FckkxKrySXpVBDRhplc8kVOjMNqXcFmU0Uqfg/UIvzVWoWPX
IUIDYOgUSGJwg9V8h7JugJ1JvJrt55+nuMobjKsDQa1JAg8Y1tXrYb9n6dvpHSYAKZW6HLT/L4XN
yURQDzjs+1xdaaJ2VJi689iKaW3s0nGW4+7wYPEqK/bNHsvA4LIEzY3HHkz/+1VGEt2ikXf0hzQC
nMiKwlsBElY0rSir9IkCtkCKQIsfePlYiiQigKpeksVGiQ+QB6Pw+qzRPgMvIzxuzExp6e+IBof3
nLiuu0hUJnCoFhZyM6p2tLjySZKKZvN2tjfbrL1LKWHkM2hHqt7mpMZG+LbgfnSPz5/pHLa8NTga
C13Lh11VkhEQTcJ5FHWoV070wOan6L5kIDReXLPd9nToVMecVGXOlXBoQvgGx/V0+Sl1cxTuqV/K
CF9KgLaruZKXRzNHa3fRQA9Tck6NIctDRWrfTKzcXS/Xqbh4Q49JfnBj4GGKG5Iysv9UUoCHgxsS
fCS9ko48Mt05/gP+qNsCpJR89ZhjBIt8rfvxRClSUotXuFQBalQ9s4efIiuP8AbsZX2Vetze2f7f
0KcZap+EiLc4NYzwzD99Z32FzHUtaG/MDaeRxWomgpAGnQMaizidBKQGYKpttsoSg5vntF4op8Z9
KnY3SpwVZlJ3IRwocxc8Pe1EVOb2a8ftDQ1Iowi33DYIUFZ2i9v3AmjF8qX5OjtKbqpxBxg2h/v3
YA6nARTQtiEbAkQHDRxwKDwf+XlWOEk3VWhry14vW21XAiCl7/Dd4hSh8ql0Y6k5nsK9UyUTrO0Z
qIwAdmNX7jgQc7safiGekLcv6nQbF3tn/g58z96fPBcehc2dp0gdHnwDf+6DbFwrUBChJ/TPY7cq
RIQflDtKcPTA3CvLqyjh8ifgG6K7JBwq9nAhGAv8+35YyjtEkteBRMzt/otEnoiI/CCi5uAfOS/L
m6KhwLFmCqQpBK6UzgcFwHUWhu8z0RpWuzbCzvXc7JZFnwzLuMGbW88i+xgCW6GxCVssmboE7VVA
r0uv3Sp5Ag0JgdwPB96eA8AyA+1Vq1eTdSHiwD/HekPlK1w5xSx3Nrpj3V3G9xXl5+lSEMknwZc6
9LfKGQEipP623Hs0k5nLTwcpC5QRkSjxJLPv98SbHka7rw4mrDozZINWPbZ5bmBgefcieP26hI1E
N9TbXJ7u1gin7gVOFpLplKooSLHbTcwBppH7k1kcg6tQLddu/Z3ThAvs97M/hhV+w6EX9N3Ig7jN
w3N/4RsM0xUGtp8ypT7s2pOObrBDMvDbkVLTKFjKCXh0Ef21xbFN2cmjiJK4FxZzmSys9YXbXK7g
e2y3J3m7qihvEa5j+hcd3Yg2vAhEanVeEjhLbXbt4vgNp30/sv4uYVJg2AUOvx0daMt4k0Zn5oEo
VpLRjpNnDm+e8pmwemv9Tf86o552/O04KTIrh6p7E4E1Qm3n38lUlrI8bX2ShK/E/X69RHHEpLon
KXGsVU//j2Y2pMnzoKLxd+7lJs0DL1NsbjGHXmvQC+vRfThuQWSaUc1VFcyCOONj59SeE+Agqfbp
JymPVtY2N4cIkzKBAlU1TvukGnZbZylbh4CFNaIF+q+ZuEi6zDBCYpgVkUuS2A6hFb/tVg7vGEaF
uIUuIjT28iXInNJm+9QquixpZy8URr7f+jadBvwg2pE4L2eR50nlAtIcndzPbwMFIKAewmPumKMX
CUTB+yWkdnpTaSX3Pjam9qKpI+LpVZfkj3bwVzGgwb1EPe9Gk9T9lJ6elmPpGKO4yP+2lLQ8DzvK
HXhyRM55K2zGBlEIuKfLKxzRh5cODzOkijFQsb6W+OiDZLxFBu1MDaVfuB4qkXTnplVmwRT+/KMj
2srJyYcxsdGEGfo1XL5kYZLTKM7v+IydAGVO4dDxDk/K/Vi7zoNeVatDKw1X8t5NcdhHC4AfkReR
eBhei1A97Wp8BJvVycFoxZ+c2GMGA/cYOQiTZgl+jEGuITg5mghbRPiVEPoK1XRP/qwNOLaBTHHX
8TpHPLstIhxGTJZ1cww9mV3PtV9SuJvjlYo5ZRzfU2LJeXsbYhgd79Zo4NiLB5xUr+sml9fV39jY
aysoMKIEiTFVzJzy7q/C2UBwnQv+r0M+PlkG813Its9oDXrzAxeIWxuY2kcWDqF07wdc57s0+yiL
OKjqRqa+VieYrCLgdv2wZsHsZPkYEWYpem4weBEV9FoYgpmwdNgzMIg3NJxNCBG2KvECzaDwPgrr
RNtoUb3gWFtfBuO0icAetCaOPue7DyhL5KXponr0mWr10i67W1Pmel1SXSzohEJQP8Ktj7AalnDr
Bie+LKFMozzkoy81z+qT7sOY32QrEG3mK5z19Oi0bpEva/3kvC4e2SG0UlSHSzMPZKlrU28WKylW
zLbY3UnL+sYn8CUM9FoO3cId6dmr6kuPpImSKvZdQR9bSRCWtl7XiDmAYIxQLJH5fpoVi9adUJ71
nUkl3iO6OHl41d/kXnXP0r6i7MYhEEAnsIMFVE2b7+dcsp7k5gaLystb0Wj6Di8hfW9f+s4gcQz/
JiClTA8jeeERVe9jCRIm797WG/iAJkK2Im948woT4UQqpqiSA+vI/BUAkHnf7FqgVbV1BNd7N0g5
LC+pEs2Y1ctXk1X3cBvPFkSFcsU2EUP7NLaYorwgtf4PwiXsUoaajAtlDQOvn+N+rQJRL8eA1rJm
WwICAy+N/2y2nfukLaUT68Gv7TKANobhI226MB6/2V66MhYsD1MwMwiYlkN6Q6VsLHbh0TErYzXH
hO1y7MD39aN/x2Qy6wmGzq8OQE/JHEdiNh/HdvAHkl/013ZvTbm+aa5XMFf0E1/OUMYEsqfv/aln
ua+pdIyZbVgdaR+5NmAVd0njP4HGl50NTAANb9hBHIFabPKK2dkviv2AAl6hY9dACfGmz3L4m0zz
I3s0siVGBm2Voa9Edun+B4ITUCMEfOIxNna+Vkvykj321e9VtJ5OEy/PpUjksrF6koAsbtCYUFNX
PbJvtr2Cx0B512y+4F6E5uIOWvaNa7+pomsTfgdC19AYiig13009KbtJ6SCQ2rIzWJ+OCPNdDtIb
t8jVa9qIvpN876OsYrzn9skJL+f4CdvZ1TdYfGjnKNtHPAi1D4d2JFyymTewZES0P3uZmZckJgwu
OvaTiIztK/XFRCpNU/4Q743FPpM1TjCBqciXBOk5YItcXJ4k0UMEwe/Tb5r4tqzPKOBZDU/hLjzx
78VlwuI9gpHb6Kf4K7OL/pY4AROpjgb6SKBcQfRg+mlSKLPB6YICtj7xUmN5W9G5M1cxdNnTB3F7
vKwSq0JdW2uusprx/doXfVM7RF2FgcRy2/OocBpEt7fhF/hyfoolEmi95C51sQhKFURMhFsbve0Z
1p1/Rr59fa3n8lq5SvOkI/FAdXyVwzE64HDWp3veblXZonajL/grViAphOHXfGAZOY3dbQ/iN2+Q
m/kqzTtc8z2Scaal2Y8Hl5b+YLKNpguzGOj5dGcIh8bHey7h8AoXp/Gpb7uvIo0G6XHGrHMAHU2R
4R6SVfcbf9tDMNn+P9fQY7KS1w++vUjyWire/vJe3Zb+yiOlSRX8GTH4OCdWb07Y1S56oTymnx+s
q6GkoJYmhHUhmTCJt4vqHUug4kEOaDGdH9YQwcOt19DxArmFlh1UiNe/3+BaClvyqr0Mq/d31VC8
UVvrV1uJ/Fooy+S91UkR1kBfTSq2wr5ulAZgF37QHaRTaeiyfpiF5dTvDik7dsWtdC/TdCouEro4
ERqmH8gewlUt+mh4IMDQtpeOt0jgbt48pTJ0rGkQXeyBnKKbB3zPtLSXpZdpxljJ0iivcM22G3nE
sBLvXIg/LGB0WgR6z8vYEciB3FoKl2mLWxHXoVqNrVvqt2U4uG9KC/FGzD+26XYBbPV/tJcjOOWO
qDS/7m4ATJi2WbYKHVmpasIF+zhpsP+5y8ym4e/4SkxT0BVhLs48aKz4FeLWlj7q4ckNeP0/NhbN
eJtP/y5kk9rUb26cGzuHM+uuHyRjSM6+l7vuEZyp21dgWCRbm3h2Lv+p+4H2pf/U3C8f5Z3LsyrZ
cIfRQU2n9w0Sn347Xvpu2GZPEDv34xmQ4Vu82YWc4aHIcFZWd+jCSEfmJglNiwUGa3ZiiUJc9c7w
W8gAxooiLfzfI6P+WXCe6u0dg9jbAoZpWwKNtaWIBg+89Sc1imannu0fuTek4dGxZ4nR+E1VZUA/
9lXPUCFQJ/MznSj8CO5b1gsN6HU4UYHRcmjDCW6O/yxpI7CwbuZMWz2bwNQLggvfeTmSLZzllfGI
9LWbEQfFq80sJh3K5Tl160+CWSWp/bhs2gj2QTw7TF1AL/VgqLdMhfVqofhY7s+qH9GPAZae65DN
ulgDJ0PHYXoi8yfpweUtzsHAiXi0X8FvzEuOquzrBJ4f5rL1TjdYbopA1MNFvPy+Qx/cRcUHjJv+
tiji/VsteQW5+5NtYa+vX52DFjf86eycR0mBOvB34IkXb87qJRHF4DQqlStYWcok68LnEInEbJPp
xWoTG3Oflj/73YG/mrNJpOzSGLxiJDpWxfiRi+409a+knV6hK2XwVYEP0LBsMvHJ0ahMGKPfrzV0
Zvmiry1bA1vAyrdmgpYPOtXcRT9+EWqmyI+7GesTbrIrX8XBW7t8u4jXxD+VVnqnsMpgJjOHTYio
FMPsPBJKugIKJnex9+iK39r9UOzcwEoGzvZufOI9pVfw0Ovk7K7W7+EyPciArqyL9XKEMbc5aQvR
b7hYXammpsxLOtkarl3JH/O4jgzAXLj+oMO++HvT7hnnVot5zEVvPpNaGWjJSu9cCm2YTpwuXN12
VttcO43UkKV8VTK15ADJPJQVWxnmtGl2e/De+SAtlJz84GON9sto1Db1E6Uhyu7me01Numqs00sY
beWs19zZ4+IdrgspiAjJec6KI8I8aL3kpSogZXN1nWNtmuwZhUUOJs8pUyieDu9B9tc796GjmzJS
9o4YhC//TIBKK6m5dqOYItdndMSBzdw/TikbYdMsrDhuXi/6KSrIO1urgKJtqL3x3HiAtrbBX0cG
TGQyRMvWOVxpDjGuhZ5+4xIQki5CSscn2zdVQXm8NkGhSxqVa5YXCKMSHTX0k5rdOBHu4tgr1Yll
tResNpvoUVkeC1socLUW9bmWgCV6kwp36wffMSmqmo9VdH/uN3w3mkTdR8EMwytEIcfyMGW1jZ+M
vC6f1+gXbwhleO4oOmvxH7eMu8yfGitC1a8tSXqRi+Ha7hP/46ypkp3K36QKMorRdEvLgcTN6zM0
hD/Ier8GxNE8M4N+fdThJrFGTRd9axfMdA7km4MfRzUAtgI0SBqhBkRboihQH1E2hbWvVvvFLgQl
5QjIbNjyLB/RS7AmUSDXD634dRSCXvB9w2p+zdcHUQCNnl2o59Mqw2BUPtVrLFjVynL8LzYfvcA6
1vE0yTFMGwGRv0aUByHNYps5U0V2F6ULQnDvklGZXJWuYNbG6D+/NxMieN5loTPe/YDDw/YRmutp
JXCqlngsMEK3RFdZGLkiHcjhFtDU2w2ynsLWcag/jGzT91NiJm0CWn+G/vi2oyCYlfX/hjPBMlz8
SItmXn39jq4qdns2dtMxmpSedvfvX13aE4W2mwkvHp7IhEMwPBXOyF9rFChSBwn/UQmUFyhs3d5C
bAyRyIAm2e563lisP6joiKdabaQnnVbClyPltHFUTP09avUrDERIJbMiihMjS8G4Vyek3YD61f16
S0e0MYKDtImJVbmkLsB2xSz7wSLd/7GacNSgC7cShziEEYxT5Cfnx+ftvrbw6sEhW3AzW5c6J+Kg
8BW5tEpxUIPxvd/17w2YQnAwJUGsDaONy1nYhXc2CxjuW3524eV07smrvn0+F2PMeMA5QlysoZhl
VYpt1lRXyFQJpX0FkfRUJhysPEGnjGWn4JEQlnHjc1pDIns5+EwTSS3ids94NZevPg1RiEjgvVjG
jFBybJv6NvK7oRdhzk+CYCLexzkoEcGyXodudfU0iHOoy5w5mJkeE/Gwr/frkcMukCuonJnCRwio
l+7ZipYAAmgfTKY52H82VsHhxCXMLSOfNR//s+kR4Bc8eY2caplFJFeJVG4HykoUYBz7HyE+m4WH
xJT/ICt7Bc4jXE8TuDuaVBMrCRng2V5hiX7GGcTWfSAYGcRLehcgMqxmqNbc68N7HIAyXgHUdgxH
x/cUN7xYaRNspxnS5+ig2fBiD8rNSFFuHc1li9YA3ynT0ANuTpwplDqqg/Vbd860N8hrIanjw8mS
C4TFoJ3a1SGirQirFDb7KWSdEBpfcP5IcJtHtzWw6cNLWIVPp666gL2G7y5i1FIP76xBXYkEjtGd
wHS2Oypd2qYzr1lzqkLOKLKtwMr5sPSGuV8+ujyJX6IkeCTdGqXUoBOjNhMIlPI8rt8dCt4gA8qw
TeGNBZUJnvluv+mw203NRuG2kF0AGk7mPAbHxJQdB7G1vbxGHsE6ZqfXgNvnSi2yqhCoyt75LUxN
PzjOUpCWrWqT0V6d1WqAebyfWDY8hWr55xGjFmOD289yuDMQ6gj2XLruRjL3tLl0hw9S8k0J4qda
rtZT/3xJTxw/wsNpKcJ+OeVlih37JUsNxmduhdLnCxdM/JS806DwNHaE0tTqDMszfi6az75FeRGf
RMPJEcr7RYMeZ7fe205am+VYK3dTdD3YfJm7R/xzDh5a4Oe63cM4/EBT8JGq6BEkKmbJaCjz5lXp
ZbNW9tPRDeBqaMix2i6glEaRDnJP7FmvkSeV9gU930xGRmZdK69gt8aY3b+FRBKEQv1t3ByLdu0p
6WHBvRaoYkOzhhGD3wDU9TrkY79r3HGimHq0iLw6iWbrA8Y72wA5WOMK51nlgWCDpRkP3+bkyCqn
lJmk7GCYfQdUlHQ1pzE2TOPZ7F4kt+h8wTfq89Gaf/2Z0i0Y+j1oOSsgVbe2uaHVEvsycb9h8G0h
peZ6bcrU8NxENJu8AtNmoIWXIppBSkxlvQ78BmVml4okQGzeDRXSBlYGidAEIDerIi40OOhcZiK1
SYIRNn+kNgN3CW8XaMGQPS5WnloZAGRS2Orrh3LhBdrYwxlw2MlktIUvKf7S/ONWmgYK/cTDRSlp
12yF5fU5DeyWmMrfGWczs2m6g0o1KrPfw7ErhtnnktChrY35UXwaKaf2wviCG5/rljCiWC843kaO
ZVJJJssGriYFDW5Hv14ydM332dQw43guWwp4O3h6Ch8quZbNa13d1/C88YrxRsFrd00cO9nE/HfK
eXrlZqtXWQQOuhhK7dxzK6i7BQwCaIpsjV4RAowPmKBVVdBy+it4cD8azkULiASK7z7j517LXrPa
7onQLTOzKS9GKLHGwOhe4VdOPjBpGOTqlw9/0Rnnj+QYq/Ffxo2mpCSGptQ1+a39tekcT3EDSSph
Bggt1iwEVn5oEtEtdCBhGq6bs1p7FDqiglStaebH9s4nTsXxZbelH5fZW2qktcKyIIYUsUMbFp0K
R9p22Kvwuk5wqSijiZ4fy/EcLreJTQ8b/OMyYQ/na9mx7Z2ECPTR2Ajb0z91WJYOLN9F1n4pgEvz
f7qDBP+dQUFcsWpXFtjBRCGd+K1dDyXtIJzYpwtVJvwi4ZH83orpTK296orWWLh/1N1DeNgD0bSs
ImiGbD5tz1yV4ae8MG3TAgE02sF8+YpwrpkGG1V7z46kcOYUjgYy7GtI548o+uPPsUCT0BLH/4aI
D68s7fjYlD2rEdvbYjMyBj/qSKln3r7r63YsjlUzU+9cnhnWarm35/bPKeH7b6glQlScgTlbuvWo
FB9VSIFGGvbi8nMyu5/tWD0/7g5H7jaHGuZP8oSWR77jOoUx8NLD41ObSUMLfE481BM2p9pt3wOo
B+3UKL9SFJfdQ9Aw30Qjro0Vd1/F9PgJD+V7BTP5RvoW73i/qF+ipLeiGBDeidPUo0xP45W+UchV
7pUGKC9fqizRWnpAJiDCDgtGeV+LSxsao6XYhGq89G1+o9yKtrMsLl620arJh2LHBHF2LNzBRrnm
1yXbo4+an+2ma+PKNtjR9wg9Vkq2if94DqVB5s4Z1DgXWoziuhRky43LuRvl34ifa14I8+4C3EGA
u6g2l5DSiOaIHBpEqYVWDXZX5SDlyGglsR+atYUA+6GzwUJtC/6UlqITb8VyLtOHtJfMaqnJs1tV
qFHR9l+GgXcQJSuzO8Lb/bsrKNz7RLuhaj3156Czlq0SuLaOgsx5jhOz36C8Ld9H4yZNydA/r3g7
jir0PlG+svCCLHDz9b6pLHygmGC2mrN3Dwsf3SEyNTf2QkX38uS19dv7WdkBMYQh0v5v01vd50Bb
kY+jfB7RJ71C0PvFFet6ebLsZQ5v2xz3T6AD7ZIgMVpuNEM7j/1QmyNSHa2BeQi09zkDlUyFOgCw
pOKXCZg+FuB+AdhezHvMfiLWbTDFvSZie9WvTZvXXUvXg3ywvKjSu9Dobb7zlOIRTyeAUFBNBKsJ
kpnNgAsXMUfWTdDuYNHyubpT3+A7wLs46XEGpncFtGsGYW6YVrDXDp2eseWNyHYpcOkrq0gswzVE
Hy8rMw0qPs9wkYX/GJumo+hie1UbmRepiY3/3QApQlKHMtmAGVgQiKug5l1UIZxi4crOtyDVhI1E
5/wQav1//qXbur3aG3AOZYkimYg7UMi4q5taMqZVm2NxY1sQH1iAmDn/tSeyRCoBhV70vZWmaYjH
TcaGOxtB4Okh3eSs14mO3VaDnFVElXJLt9x4TzSxYC8nPNqBYVc6+hB+aV5CQuysCxG64qTwKxWb
7pRhJ+eUzPKVUsa5jYDTxUfT+pM0H/Auq7xa4z7bq/+7upJz8FfUF6nu1RiAX4ZMSZD7ghTdWAxz
c5EoUig0NBHvizWm11ejJ/Pqygqqg8KOlkccwRLT1+Y/ABRA3EbZOtCT6YVwhdfIqoTgg6H9V6iQ
7JUJ04wQPEHGUqPQbUDiE3P4MZWBPu/w3VdS/S6eEehQ+f7BgrL88b3CT96/q3T9hHckgt3m3hlt
aIjIiqrtprcho5qw6tM8k/56gru266OUu0UppAxKeDKQUuTrAI3qiXL1+uMHSnxEEKdAKpohb+p2
oKhJjNYZjdwKypPGbnUDkbVx0m1k4RO+WZXfH6v9F9zriUGVpdVM4nO/oCmBaZYtcv0WV224yDhQ
wMT2LfgckbcBWdQQKvrwVLEN5IOqEdoalDyfmTIks1IZbd8iryoBKPhdwCNLYqCLyNAov2dErGih
Dt3eAsemwaoVTapMujnrAzcpfDlUkdYWMYFYTeqsU/33euqgmasTAgQwhcUIN4X5fKNCfPeQgKyT
M1lI8qwZcYTbreQu6nGsJ17aWsowOArr0LkIB2f+FquMKc9AosVF1/VSuHt2k7yiXayt6tl3NsGX
9hAkHPs8RKbRKLcWJWqT+oniWO6QydHZbywzATnqH7giHsmaNJiYKJwUsFURjABFxo2sEnNxSWrR
zLcOER6/ZBirGclZoNU5icNVGAWqpcjf/962G1NylJOYkOHyj2+MdkJDbkdigVuJzKi+7p3MQeH8
mkltMiL1uGnJEPObYE21/GzHq1OMyEedDuGGo9WgHB/Ttwc/9kZonMkpsYwSWDrMFhnto+COz2d9
RdMaIW4Ybf4+fKw+mXIhZ5tKFI9V6hBd3x+gIkEcEtzaWoG8SnoQhTSox+AvdUM2HWZ3cOD0Pwdz
cIVrVrgpC9zTOf3Ivr6jyH3m6c7r59WD+FZh9yDKizXcSnjfr21CZEB490MCO2p1aS0dJSCGOAzM
QTnHBl8fQbkHV6z7EdS9jo0KrSwY95c9zUuGpPE+SRDiOtu9el1LdjQhaZTILuwPpdfRp9TQv2cN
RHNAyXjd82ogxXdM2UW8N6RcaSsHlTehJKtrHUHBfH+prjFwvokWwxxLlcj1pApT5FDtcHC3wcAG
apeDMj6BBB9M/Q7xLOB4Gzra42PawiMKY8w9EQ1iiD+Y9K/1gF5kB0ubr59FNMJWgwxyk75qLzqg
2Mp4b/ev0pLmMJZSFcn6JbpHRQZwfXmv0kRGiG6lgJc23KmRr6gf+SY7AtRr4FIH+bBWVDhcIS5g
qOgHQmlerRJHZqv1N6A1xLHm5G+XKViO6wNZArqi3YPaLyf610qr3P8wLEQanIXwaPt/1ER8/9XV
9lcrxJefDEu2bx9Dol3fcjNJnSu6XpzxmO0sMc2/I8wn5acD+N5O3GctBMXJpTW1HUbSpenk01hz
VTLekEcuBoerQ71AnOf2hDv+hvyyLoHERgt82+P5anAJgZKNjlviVixJ9NnljxYZ15lUFBlPs6q2
JFqBQas8iFp/GO8EECJhOIBdqckqgWi1AeWDf8FsShQ+xTGrnav7RisqPwY1jwsjiQcwVaSb4CUr
obCPolIIVFmTl8OWbBTGGp4Fj4TlosoK0ZGBP62XJXGGGHfkb7PnNRKa0mF3tlXbLNtC6vlgRp3w
9YI4QwxQIVz5eT9a/T5NUFT+b3gs7Sk8cENUe4zwkGd3jro+XCMRX3b3mVte0bW+u7VYIyG+6/E/
mb4wBIpQqT5a0SyN7hHhRtjVNZpS0M156gwYkcUtfilBiQvt/G7IPzF8Hal9wfIkpQyzMOStYJrW
a++TqyYl3/5cfXpDsIOWGeBUNwnqJlq59qX210iZ3NEZ4uUneUvVmugZKscFPY8STtvvf1VKjOJe
HVpse8uARKeFvPxi4xocPtpt7/PjFz/jr8ozaqqaZyy/MfsZs/7RNtr32QKtpm6igP7RqnDpoTSn
cbO7Ln1bWuTVLxcKahZUn7Po0YReIx3PZGhYfGah27raZn8gdd0PenJxulGuwPUpXnkXZnmbG9Sz
RGgXnSFlrnSC604NyMKdX0lDd7C/NWi4z1G8tZ3pdXYuP81cNgPmBZSv7WhDlRjzdtEYBA+/MOiQ
xWwB9StmppSbvY99PFYMqfiIhvq3ix2j1kyl7imvIFg8jPiz2ChBayx4pc8+u8y5JIFjJziL67aS
PwI1CB9OYkfHyszgAAUifbeH0Y0eUR2YQCyfYxBsgSswpLFLLJBkHcdqgTbmQitz0vXa3HAlT+oE
pTiDdC9H3opzerISUq+rK00l4ys4pptL7tknN1Y4+6kp6x0cHwyJJH8RJ6U3HdW2Dk2oSiaZ04ZX
fAPgVd1VD2Cf+f+p6lViAaiSpKYXyat3LHL00ApfYRKyYwNPEJjMD/asleXFpBzqqu8sQEkHYHnB
P3LyOZyOkiG5dD2yKno5gSIo0c13l9Ran+pUYyJBwjsuaLRzjtYcr8ANnuseGLE0yKTg2NUFILYF
6Yyyk0sSthtJXdlalnfL3YWT5wzup3FOafqQncaJ631RIXKD20iMI9R1drDXK5M8vhh1T+Ut2rIG
xETBG10Xd2zFqh328suOGGxCMK/6kAfCjHsfHu/z7VPoAAnXleo0W7JFepRgT2Fm9JdgSDINqQYT
xtRf3IiVyb/o8CWFsfX+04mcAK+v3LTRK8Q1n+DL6v2+oz5jPT+cDItcUxlCg4jyD9EVfAS9EvNf
uNICkeK1CSDJ5pw3M0mPPaDl3bOAxvgkJ5cZ4mBCxHZ+WOkfID3jZifzN3USNo2yQY8uPFk9+Z8X
ckO1/WYwhVWcy+C76tbw9DzWLOGVfkrxq9QZlBUOoJ96/4jrqcEaRAorzZftLpalGSsnX6lgIFOp
+zXczihYEB8GmhnunMwz4b+if+JtNlaRLsLDFDHINWtJMyZMaz9m/BbII50D6Xq32AHaFAD+Pe+3
iCGUHdcTwXyLRZF8Ghm0rIVpUuUcmikqGZjIG++TdcpeJjgtHffdjDkLUSjU1WIBIlmspesRTT+K
klIgyYFWXspm5o5VDzN5h6xTX5C1lvPKd/9g83usyDv6Ys4mvmUfFGZyBVYPczcyC0R06icF6uDQ
apxnLmLgXhFJCogzCxHzQHzCbkHlwGMJzb650Y7QrdyilpHP2m4Ap4lWuLrXXM/QkkpwkX/MbxEL
BfuM+BVld7UxLGCrFkUtW4kAyJnm9+IxHLks36bKeukk/FcRK403A6pQLlTy2M8d4OR1TK2xghNB
EnUPuRrRW8exmnt6nqFEAMKp4Zld1tJJm2rUpRnFZld6I/mn7WZj+MB3WWnPrkYuf2jJKH7gBM9k
xPZ6ACRBfqmR8wJ7KO/GzLXfyWZD4tEzhmSuYb8G/l6WYiej09inam6qZu0SU6B5qaTRCu+rR/kH
zmQrKcKwz41RPlqLFnKHahhkDGB/6b3GedXeNnxxQb4PNT9gh5Ac8LypPuJ6aHQHtPp5nN1CrmX1
foxD0pwR0MVhfXChV8hqcMheEVCQ4+CT1/Urt4XRBcXgtGjsiP7AMMuQngSBJv9DbRb705MSvnll
tOa+SrbHS4ffjDU0GrxE82bnmpAopupoZLQZIX127eCo+UX6Bp0ULK47MrU6RFMJz8Yg9iL5Hfdf
dtPB4HeKbxKqOtQ6SqitVYDj7nrFoBhSb5LM3HS/O6s2hmaCT6j3c/2mqLGJ9jfB92hJgguijm7n
Mz/MZ/2NB69hTmrIesbUosbNVy9AgrF1zak2llqRa8OhYJNnxQHMsrJ6uw/rCUFARKhJTxugJiuo
vgMboIvT5BDAWXseaNJN7fso1v8cOgU5ND9w+8846aRb3/P9xUMI/vSiE6kS766iq7PVRPir2GZq
hXNojywMJ7ANNXyFAcaUAN7OjG121P1b0gVnWFKJvwr6vFHGLutrkWRJtIlys6yQk2YDt3rR5vy2
NVJLoV84S/htwm/vPDsouBq2C2+F4HyMsGeZ0Ms49kU7GYEkroAf8tR29rKWn2m6/Ooxv+23L65I
U7Rio/n6ujZ1NB052H3710Y56QnUrmbWLoHemZHoY7I7BWyi9sGg/9+mysBfMCJ8wfu0441Nnd0N
q0lwphVD2WsjmpmG5vJ1iQJa4z3ewliQzxChD+BXb5E0fESBkO3umMngr8U5xWmK6+dmPtzVduUA
LxVr4ypkfDG4C9ShQj3jcPyFYIhLqggDqEjQjMmWU14TwTKnbA8l1Nva03jpTc2ERU4SSnrADCAA
omtV1BbSzqcH4uGPmWiblQvSfEhqKO0bk//r+oOmKVatVn7PmABTNSp49de8QBmjIrHqxRFxniFT
fp4vMRpxP6VgX/gSe6qmvGTS7fEmsnVtl0b5d8I2OCtYgKlEVGnUl5zwKGPZA4G8JT7xgjraMrzt
mojA549e+5vCoL3rQidgiG0n1rim6BviNoAQ/krCKBZ7uNoS56b9wAAPXpV/07TgewoWCUnz0PpY
mH7qoVDejF3ZQYA22lC7Ub6jV5jeD6TsHuM/EKTeMwNeqfLR5DO6P+jdSRKXY3D7S1/DxHG0YvOd
cMxHZ1d6YDQrI/+cNsXBp3aNnrf/kHt6EVbB2IIyGzzIi+GdVXk1KX5w2fcupAh+8kqTjnvgo2Iv
cNof+Yn+HgXZtcOFoJVyHp6ta29/MbPSpqr0NMBxVrx/ZV6zf48jSI2Kgn16qVl2S86xZfOX9EBs
KJZISSrsZKYNMdwaSZdl2yDqnqpcVi4t+4qpKuRIUg2bag601bwW18wgAbVrKiZJG9+PkVk8K1QV
K2hpPTKQJuQ4Z0GFhKjhFJh8wuOLCwrcCdRf4AAdotzTPOang6OMkb54OX9ApALjkzT32Wvsvnx8
WIvkup5FgXpniT6jqMvVTs4gTCjZV6G/MwgLCqP7WES1glEZleK0VEBgppfQ/PNr3HkTbpR0qosV
B2HviusxW03a7JfSslJpkT4SzFJsdlVrYq5cTUV59WWPCouGqB5Jm7tov0VJR1MwRSXNcHIry/Yp
NLQpvjFES862/t0tQJK2+YAwt35bSv7yuPLuNzex5SnaGYCSCuk83ZPPTJG+37gyhj0E20z0a1E3
VfT3fK4xUA+Wid84tvF1H/eBI2vtEEm+aAeNpQpla1OP+wJ4E2zfL15x2kMIaFSG2W5uRpnIPR/H
XahVUkgrhRWBl5dCf1q+wwufJf8MuX/CLwIh+TdgmN2gRHytrbDQY1+fqkVdFBAx3eRMqYg8H1aV
Nb76cbxfwrrTDjYbUb/1rY8v7zVTO9/QJ2lM7/Igio/lA3UjC0dPd2du14fxMDR5dx0+ulSvl37s
05EHnLMKEiUHfdc0SF17TKDGzyxXRpTY0J5BdOKAUuR3PQwuRr7x57ut8M89uXXv77bgzPVHi0Y3
gMVT2Kw3yf7rKCWMweILQZSczxGxrgTlz6pSRkJ0Wi+KxgzNOAj8zN46pMUEt9+HV4+I4cgykyc7
Bn5JNY7IAoQVGpjvG8goSdCYlDh7GyYd2LqrkANi/Dei5VnSqzqtTBhGfyUjV8s1rj2kKzO8TcpL
TDNX72VTmhQWBgsfYEPQqffHHQ+WAjDwVdfO2EU8S8ZwScTT2RiIrtsycjaG3QBxGmMPfRd6xCki
eWtbh+pdv7Sx5lyhNOOXSKi6v10l4WAE+qji8XL6ecxXP7ROHKvv66Pl7s0KFaSPsEmafMhfxHRh
FyojAvLHCqj+5UUMjNr31WJnPMHSwFRNY5B06Lz7OX9LjKlek1i7YYLTWKxfkrarXPjYkDmscVeu
kQawIyzaI+VXzjJkmI0+wlkY6xoyMa4D0fNfyD623yah29azODK9ojleGEnehmiArawFz8qPHBOr
9hkHkiCqdkamiF0mzMyCtsPI2y//q9G5WUpiKDzbBkKcHdI00glEyyw4podT3wdlEeWQ/KAUQEjV
G21LV0MZ21c9PTRLfYwMKU03KmcaTwbhyoVcOO9ROuttXVLz23BlME3IMHysbRBrNvmYbrKt9vwp
mYk5MbxslrAGUk+qBgSY83c6Z7wniB+vLSTRD6KuWaCIReqUbEg92sDHFv1LoSjZGZkX/znrJm2M
ZZgMrJaO+gp51mGVALN4snE4/W26mjIw+i27qJzcW6AqtXlDtmM+bBoxghlQZjgoBnEWr5BYMpom
S0th+0lR6dIBaUc9Av0WNf8VPyElYTvClt6nFh1+cQJOHyRGBMKfYOZmJNnAdRnTmdT3Vdgd++NO
cGFGdv6uyV9MlCv0flcV5UGc8KbB0xzgGNe3vb2VbEKsL+L5Ny+F3oPpfEnoK4SqO8HZZzgBFZJN
eq0VxWj2iB3VRLDtJ7cVQQpWFML+hWNUjQyinyXyhciVbNOeNob5MfDgPCTv8gq9c8pwjP3OvuR2
bDKHDG5BLUVBdfl3USFl+mTJkvffZKn4bSf09ZbERABSqKgdC396juJ2ce93g/+XQrHlJFrQ+PyX
HYuDPnBDF7tp/h04V2iVtnvft553hAZYqncb2sL2/xzMiu1oIpMt1Uf1uf5w1AjAahOLmO+BLm+f
+j4IqobiYcdsDt8RcPA8hGDdgHwDBSboYmwCgr/0k1kVh1t/T46jDoBlTxicwFOlF7umzNKjJWgg
/LpmdGWkaibYtRnWt92M1wyMwkhHTzPiJw65sTcdmmC52ohZGMnw0t02eFAfNGfJEyE0AaQ5bmXC
pT94m9HEZo2kCaNJFg6ry6QyBUHFyTeaHdN3bIbK1SD5qPtdMnST0RHzi+/r8seL4zazqOzMZNIq
w/IFnkmgRV2TwmL8PH8b2ocrPauSzsx5tJ6rgmNkP6j+CBjSwVrr9ptlbnY9HBejyTV99PRjaBz+
XdSZ3w+DdvXSwY4p7QQnjXzW6srE5Abp/76HGbB6jyng2R6gRNr17yj2gFBKKd3i/weuS1jltO8k
PuuGN9fwe11hos7nlLfUjgDqGFXDACE/Vn/NhBzIiiEPs+88grV8GXLNVo3kDlALLgtLuzd3U9KV
5IbUDNKLXmZCAGmLZ2hytwe+sqSo4CWlMDnDHSTPUSjtiOylaIIR1n4iIXCTHucCj1AHZ1ukm9QO
nHoD+jCRnhKDtG/i8A0vgpPU7rBnnLvFM14ZMK7P2PP3ulYGTeC+RpImy0185EaGrSXBpVb2Sd+c
pEgemtgG4x7tsk0Bv++w1K1nCh8WISvNmI3YWJJgcQ/me1sGGjp0MS4SW8ionxhySixb11QMKrRA
j+W3CFbGABqhfMfkCW6EiITuhdpE+MkaVLMQosmzQ3/2f6Qxp6E6fP48N4+k9SdaqxUYXsNUDZwf
VadmR3oSCI7ZKWWgSyriC3K4oSBOK4tEc+WOkk99qBYd7l7dRWE8/rwGQwLPl/rSEoYaoG351Afg
piZCobr/uE7lRaDLxusJFuoH8LSnnaorB5MLgdsc9/iyOyMjOWyIilMTkT1NL0q2IXRcqAlmBWNl
y6YlIQUBRV+kt8osSMxLBhVtgC7CKojiIsCZdWPNXcp5ltkf6oKI4lzgmXZ5mPU/Q0D16RZrnVBn
ScH9VkJfMDNQt71xY9tS6YW5eH+kjGjUAEJPMbuNupsBEOd+ODi7CmeDPqO3KStTbhjVbEWu2Ij/
VK+dh2QtBn1AKtr7Orz9HBfy1smy7Er/48gSAHjyj5IkaVPP+lPp36IwGkE8g0BN+V8Ruhoc/VLh
xITIv75Z8SrbU1L4JJuaXVfFbJic1zmq+ATS2FlBJ/8SoZz8lvTZ2Bi5ylpWaU3qtMjwS9Lu6R3d
5HqDg2DUq8oEV7cHHLP5w8popozYF39NuABWm49RcnG+rlCbAYPCUkQ1gvUshae8EQjPqn2ggHXU
PStElnYLDYGopYdRJP37P7AbmtcBlB5X9Dmc1rdmlb8ROt8M6EWr0opvofBDdG6aQDYDx2/vYxm+
Qiw/b4KsvraqJeoPS9/8uj1up+K32zwlaO+JrdS/tv/SVeaEZU/kvCVuySlj05/EB26UdK0AeJw2
p5nkH460Ia3oldpfHJ+/6uGgPxsaOIX/kfQgMwfUhmU4hXqGI2RgI1tS1wr5KyZouWCsATUbgPq9
358HNTlP8TxNCfDRBmNaJTeNmO72P1WU2rYZe7gjPSw/i7STMufkEuyokJdUalbIkVNG5Lv6nsfi
ZM8hZvx3B5NSG+DBL/PLQ+fBLLSHNrZm1Jgk1kIVRNqsI3h9rhY+khjhlV3RivfDXB47aaaDKnqJ
Cd1kQyReu1FJIEyEvyhafVE2lSzvAx0a8adztUt3V3WiJVBvyCP/7x59SZAluApdNcf48zcMydvO
CvSugl5QJdWkJb5GCLQQoeqK5GgTC3mtzthV4AYYHAqEKAQX4O6RV+U2r/ut7KePsrGPevWFLK2N
cUbg2ynzx1lGxCFPhe4kHMbOReh31TM9MiXLh3t7aeLoLVBcZOckquiupPwfNhwc2UWb7P+6N5Zs
ONZRnCkWQjSw720xDMUHsYrIbuBwLry4aTpmZ6PKrq1jd0XlhbffGWqQSIhSiOVx8drNaCzJTGrk
JG987kKrd/VTKy7vGRhprAh9JMobnT1g6DIlY3ga2czKX/nK9LIjlpwImPoERXHvj9d9M2akT8bF
ssI3Qd3/kuZEc2XSbmVVcOUKn/WFwv55BMcbuAHGKMwwKBqrTDmSxwTsJMXrZudH+1RhKEcyFe7A
tO+/oJyVYA+2EXDsUp/auXnOMBQo7iF//mDK/9dK0+0XNh2Omtwxfj5ha2iQMReFzTUYOly529FU
bCvM+sMIVrRFLF5D1PFtv3GARgsvTZKixO5EItnTCbZJ+5sBdKwnQKoM7FpENWRuNFiMsofARhm9
9jpXHTiGfCZIQRGdC9SoQ8MVl7p0RPdNnhMEjNzSWhT9Dhd+b0knXzSeYGPT2Bc3VMXS37J4Kct8
f0vA5UWrNjcUhJ0mkbfNMcfchdzzJobCkkHl6ZGq1Cns37SUIOLFUh5zLcgFF+obzj+3WudC4qQY
Xm6+/gqI3SVSYgZJ9oL3yRD+5CsFeLbuMmKLe5VljwuFbwa+XXzp9L2KvGBaYxMgVYU9dwXp0Miz
MDP2roxrXb5weVC81ftjodR/3UIGxkthch8NcHNvtnuOZ7YppAfFpFH1FvYUBDW6Zy2Cgj28sQu9
DlYpyIGdPjgHQi9p68nhNqkCeyPcBMUGCpidyWQh1jKfMleE9hE2589oa8nCn6eNAV+Xar0yk+8F
nvKslbsoNBQYnEP6lt6JcJ5FXkE0hSpLob47qY5iaZQz8bMFKb07y5aNVQjT7z0uEUdqxMtr6f9o
pwp9kvrH6vYRV5YHppLTZWmVTuJepzlrfmZuQ2AntD3X05xkCTGSPr74PPx3U74w4OtNbadOfWJP
iQ31wQhEjmmwXF19X/AMQybo84kkF0Gcsfmi7JNW9FamXRoNQQcsCxokLLHPMGa8nZQvPpzPOXbB
Hgt1pMhX8fUp2LCTwL9152UVjuo17gWnboYQMLU7aYDnayNXtHE4n8oCDjOQbZToIKxReraEf3gf
p/3zJjs+ZOw2uwmg1F5z+p0jBEEprmJ8448Jv+CHRCnVcr5TvFxIWW0v7pQGn8JsaVFpCCuSRLKI
a8eFhXH5CAZw9MgUnAeaJFCE25BdI+vNCcpjsRmrOYCIK641I/pjYHgcjQf0WTkHZ/NzPzZRcxIz
xFVoXDa/HEJYAOLwZMdbPLTXzyP+WnR8N9R5+Sw2yuCiYllGqAUjWTpP7cdQg9UgjfZKjgdNr8j0
WDbVVpK7+PGQbgWSnVezFXFhApCu1ZnEDyLX0sDjeRJmGIZvaAnudY+lZRYnlXiHi4E8wrV0xecu
Kum/MmRilC4DmQrOeCPKgZUGubbgVnA10fJW344N1p97nkFYGQ8BAV17dx8xq7phNFudzvP6oz4l
NZZFlkWRmLUkj/6WBYNGgulxRFyRCTBTbHbJk4aVmFtmLQ4tPuPGl4LyEqbvpQgDxJCSKARJik70
xh4AKbVyrItIEiQ7kNrLvEST4ngjTbA5DP8u0+hWWqTtLgQ1emxHfQBZ5ZhFfx6CCMrTNIVn2YZm
n1aw9TdEAHr8JcX7Ccq5r/rw+58j4CsW/JAmr1S9Rhygvqacd2g/2opm9x57qG9I6scIf65JeG9N
86zGhmL/2tQobi5hLjSxmLpVICSTvMEwDxo2PguIecHNCxLgOxLIfEcvipmpeRi80bFXDOzQsOCa
0FwIAZyTjkhdMahyDa63WnOukKhPRZPeOycDrOPquKaHHhi4V4+0vV5KRq+JEjSN20hjnvfFnCXN
cFNgAH+9CtYkl5dyY20Menwk1Cq/HlahvXgNaz9KfkHEP+GR78dzN5GqwxykJC7700NeTM+DGDJs
xXQ5+Xx1LLej+XFuf/0lncownU/iV4dnwxvBw8v19MB3MdpgcXyMEzqeRIMQi/sUqa1Tr1e1zahT
WgQKpqEGUQxbFpSF1GsBIzAtNhkUF02wON2KpOrNGhIQLjJdIPgyK8tKdrZ+GlAf3x2LpbyB15ML
p+42C5WPYl+GsTnHvhRR0dl2wKqHT1rtErqcUKdGRZUWvSdkyJ7BMV51jFjnpFcYhcPLWxgzXwDM
Hs5vacmoZm7f//pQshaSZXWw09wqntIWnVJKDk0F+93QUNTECsCxWv9TbiE72kW0H9y1Z+IUEmr/
NssYuVqOC6dhLGbwdl4cjyx/6tmDo5B6szlI3hc5ZjJSPZRDWdOJxavrODX+cTt18Ygleos7r86X
O8cIjbawDLqXLc76bRmhzJwBINSp7866pf9pK0HoaQhWt1YbJ/wiivXawL0wmzB8fZUJrQXidY/M
+8qEDEHAhWrsNOa1bgFo+WdfwS+R83i/js4OutevO68AWGRg/GgQVlTNtjmZbd6SkIGqlNewDfBf
Y+6Df6KWIse9i0IUVxYx/Fp6KD4T3ZK441pjryESGQQ4AE8K+6VaW3vQvF6wFNZG2bdFI/dXdRZA
ds5sHeO8DJjAQJKL3/X0mY+bMlGi1tBMX+CEF/8k498jN/2DGYYA3AdcjDCGK9iSKQir3MYWQp7M
MEok3XC6TiOe8sli3l2GJ0JDnPTHpzWjoDeTbYPj6XNkDxlB4QvPVatyf26Lg8DXg6B3brxlZC7v
piBdb7ECKc0JHW97IkbcTviofKM7GkMaUrOw8IzTq5yy6Ya4uvCtlKSSx5s4Ojpkwx6hhmDhW87l
IiaEtxsZQVomZT4tGJKkirmkqEfZloDPGzhEh2KS+ePzDXA5Dy69mn+n7McQkRTTo5jp4SyZdlkZ
fFqW9Ad4F5ezGnt3PMklJ0DPgUAAkF86I7oU7fYCc+vYuThZLECN2nuUew6JSmaHzgmIdpAoAoOW
wC2M5GcTfFybe2Cgbwjz7WBWoMAio/BIJdfO55bW+PAcNHuXRLl58OVtE5xMlcKWx/PSR2zJ9YIN
3N3PDxHsEO2M1nITWIWuo7L0+3FGXF3SITcyE+4ZF2oaI4eHArNsYLLco1MVFb9KCqJX1C0gWthm
W48KFswY3IR0vKv59SGOo2ezHSoER24cEgF4drgFLHLvpw32asI0ki9C/oksLLamjfmYYdrjWiFo
1bddGE6ymici4qdWNo9sGy+Hbp/DijjOfX/5I1J1vCzJJGIcQsl2+se1OA8+ZOmNAEfNJkMsUDBe
WCBkwEnsZQHLzJsPJmh9Mp1Z0N/r/RbEDdE8zsLaJb9qW8/u2RaMzQ/ocmx3nH5XE7W/eQGM3ju+
SO1SubaWAWaDghKJMsXXA+Tx51Mpu0f4G1dx2KgRQ/0/4OXtjsUWPL+S+ciE3ozy0Hhlj2VYJ93D
bM6MraCVfxCxdhOT78JtYN6VeQ/uYnJXhf1DjTt+4ZNwYcS6iJ6joZgd6WgChEoZtoEOultFjCVm
kvPjgRgUDZMLgaaQMHwqusMU/xlvMTMgCEMHh7dO/twija5P8JZy7F8m5jg/QQ0gbuzg46XZyKuJ
+lvZPoKohQAKUJHTYZLDwQm8U0L8t58S0s3DDq4L8DipMieFAPRm8JI1hrljwFHERDMv1t9QRmwP
ZM3X9lvKLzXahDDpEYyjh7pV7bF9ZEWg2KVx8A2qFVymKkFALskz66iPp95R63cvy5LNaqNZ7N6m
MRMpEyYgGc7auY0/aBzj/8uJ/VLDxqS7TXVEW7NfXoXm0KQqZoZIn5FzfMipycVQzsA54VccR52u
ZkZOs+lrRyeyYZJKo83GkUJtYSX6ZcEHQHFv3jOYQgZF4bSNm7aIK0ThhKKSEWPoEmsp+eEZgD3U
WehpVf7v6NcI51mt1bJMiVv1580RcuXRGlN8/3HxLJfSE7YkHREydlkksKbvU+jwIE0+u1TV7lZ4
efWDRGdPMX14dhgnpR2DeEObSmiqDrTcGDIF0rRT2MKDrn2uNurX+VfX0A0461z1OfTKymaKJQ71
gwHPutqvkG3eAGP4joqOmvwK9SCGTz43BYwGHcCDe3cPn2hGzA5cs4w1nOsX3OsE8xoiIKhdK6Jl
5lJN8D1K6Vbzmzph9e2kPk5HnGtQ4iLU4jY1pXmnmSW60KsgwINSYyCeAL2JrRiJYMMQTIoDKq27
dSQ1MF/S/8qbHY8UbqYIVBsDX5xQmTdYDWUcFgHC+/8cHrwhIIn+ZNcQuEUUSDi9wt6qygmV5NYg
JzBiQLPXIQRwFSgg80U5wjjw6qQsX882mc8apu+HfQDKKRK7sJpuDYmt8wIEc2ah90xFoYnQR6tp
uPXkrgfwSyvok+/s0k8T9UDSOy1wKeMdWuhOsfqEyzcbTEyyzvidcxObUAweAic+CGbuRojWn2fT
pSt76lsm+knx8AfiTF9Nommw9hA6mSTB9tUEtXYfIyvIMOqg8mOXrnpozUQ/HXFxfGKQmnbms0c9
w2H1usbXF1FzzDvj7tL+xDmc/qBWtALtEcjW1H6TxxocIxFcGgD/WNT+gY7mUbaprSBumEKiwNGU
tD4OrpcnNie3mtGxBmyBDk/+ncBMGqKAzhDF263qAc8KGlGcC2aT+CTOBGYvxasqdMEQRWMrncTJ
UBvA1+Go9vXibChkGFdVnkqanbaLNHL3maTzeeKSZ9uQ54H6Jq78M+13UKgGc/nnpmMm5XZsq0YO
GVRuwOazb7amIqET1D8MLXl3AIHZZVnnmeRANl2AeMIStn0QnEXjhSxq+MpKMniCUcAwKa3nO+3+
CtwYKqJF2zFgfnOyM3AQO+VgHfwC0yGkTbfXoPz2IZKQwggPozUvMMpLocf85Y+5eRXU3pVIKRR/
Giox6K85TFR7UOo2wZ+yBip7u5G1fT4yxtbNt4AAitOiJ8iSP3m3r2yfsMUxDTguYIavAJmFa0Nc
XKLVIRLGA6EIJmiNGRjuuKHY6pVodoZDHCShzHHVhtB+1FOzw6wqYwMCeZ/BywWFZqEhPkrDiD2h
om4wvDCEtUp8wXbaSME28Dh3xfMxjjgXsVnpjki9k42zBgM8CsaOSynAYaDEHCqsmTp51OQ8Ti8R
HDT9QJUt5iu4EyLzJ7P5Fyr72h2h6tOdIi8H5xVmzVbv+ubMbseGyWoLJ+Vi8VBMEdYdAJwO+PLT
xkGSbn8k+9Ix9cH9+4byI3mKrqLaaaetohsOfQ2uI/xGwhxbuHg0aRfgsjjqA0gW8pxSSGuT0Bh2
qnH0QIdh9/vjOpYOwIBN6SsaWiIpoTvC2tfyi8MX2s/nN5S2G1MCCto+POEOd38VtSuUoAJ8B2WE
ET3nvs/AeEaZwnTtCMJh0doGeNEqzrANoKazcu4Hj2mpWi3yE110sse8lsHwAJKxcYN3bxDfLtYL
9fgyIQ8FfxGhS9S5HNLxYvK2kpuebJU1MG9SzXdqc1KhmYbwTv/v6gaWDMgvFgAVfYecvDMcIRsv
m3SLPVgBHczFwd+easfg6Wt3fptdjWTeBEdKvBhlucLCE5UVa6iagnHRIDNa/i5HeFbVIPkJkPF+
/qvteJxcxclvbQpNKknkRx5krcGPZ0eyTP22GaxFrU6KcxfsEB1VXhrZXYXYgyLEAeFMScY0BJ0D
kbb1ZkbnePbwHKjwSchKRHZTQIqX7xdfdhyPFHoVy4dx0+YVGew0jIiL5VwV8NV5tMjy91R1Sz2m
qr8Z9wVO6KH6P5CoP3XP4s9z0lW2dsK8YdAf93cgO0V5eW2hSm2p64+TGWAqKcol9MZTEoh5atvr
KRD4r9cadIkWsLUBr/ScPSo9y1aAJYIuWqdKndlRpvNElRtHc2NYvNmLZFS9YH6g9HSRB6l/jsuo
FowYk8HhTV5I26fTN7sH0JrEOI+TduXIgSbpl6fvaLayC0yWMEgps/nPO4C8AvgWKRT/HtDy3bSk
2/RGMMTyB5jV4Bua1/hre9Yuy9cLrt6P39hqVvSoWfkXCV0fcOMyjrkotryN00MeBYDPkBSPUhTW
NFrmya5Q/R28EphQ5hHDdroWdoHNRbibghvoSYQu+R1pj99iDtV1d7KZS9Z13VG02xfxO8oKCnQR
sEEu6wgXey93FFY7zKQSyKXlfA+/Yn6Tzc0tEY+bv2CxiKa2vY6rmK0LmFiVJ9gXe6+8Be21qVYL
/P7slS3wSryHc9w95jFU3a4HvHYvFHYJLo/GOTvgKEY3XU8m+fTgz+U4zbKooj3nPrrOMkVr16LW
vlo3tLJKCHJK74bqe/wwSPAHQ1srqutDuVRr43jbDrZV4FaaQSRt3nvl4HjgWpFEJQN6F1AIgKMA
mbtJw28aJKTd2kbh6E4uW5h/P7TECG6dBvew/xAkKJZF0L2VV/qlzHKJpQbd8lJGuKX75Irq4g3Y
Zu4QU22nJv6AVzic4xi+VO+Pc55huoodmdShj1zlJSW5/TnOlhsegYo0zvGD40WlBCZAKkdTebX1
DOgMZnYnNZd1QEY+MwmvXvSQb4Ij6KwgYAcVfy64bcq/35fUjYLsFsdsygN2nhVOakxzalZo1HpV
MTxsgposnneTuVgyn6Rrqma672G7xKcSXUGOSlHs51ChF7wP4ajglYMOiigF0zpJWeIz2AOYeFfC
xnY9VABvTU7/F0e18ZF6M14znf77ASyjyG/LFVfp/coftjFpUGfCqe1oD0LDcHoS1QoEGsg+8n4i
lUabYqFdAERPw8HvpbzgrVz/dtmn+3NDTYpPYOzlx5JWbA1TKVgv9g6vkELMZvd5jw9ZPYEjcmqR
nG9Jeq8dirL2TlNg2JqSmuCG2V2oOWRdEXI5h7jcWs8g48r4snZ/qT1IywiGTQL725jdOfVF2rOd
7/4C2fX2v6LHWTbIuVhYQVuGPKBenmu9w+hwBYosZGFnbecfySj2CkurfZRZIqKsC8y/Ri957fr7
FmtyMILa4BarCMgBSDIK437i5uhGNVvpnRMBkkEKGNeQswSsxuydlRDgU9q2bUtedx6Ocrj/IFXd
2jQmUrOB8jQpG+uToe2OYzO6IFt8uRi4lL2uFnY4KI4SeVVt1g0YAxJwNb/gefHEhBiZEz/LN267
aiRex9HXEamBSFrqDjOEOpA9R9/y8+8HGPx/+jifeUUqU+UEoJ8IfB2SIXYVbKsPsSDELAQlkunk
qKjs09Xv8aZTtJlH6czKVK6aX8apdAGXodlqRq46ZRP/I2Z1aYhbrjwgEbhO/qopZnXRXLLhDLgr
XMpulYZrXSRTkEcpHvqcNUM05R4bpNBKTgft8FSEeMepnMf9DF8mNe8NRBKEfoU2JU0AQyfDYonh
sA4L7v3nCYDVANHkMzXUtrQZXqG6zH+JmBlL8P9h0xWHzPCRu88idn7q9g+ZFDwN3pom73Fwy+CN
jhYrhx4im9mEZOwEsQmwgY4dU2Sd5NtTFH80mvXu1l5RGrFpDc5Z+Ccl6f/dFtfVv8tNG9jhdD8L
bJOFdCcr8YpVUTrLLEinad8WNw00pfGpKV9aWmrrUG/NYNXjBkDcLdaV7d7wBVzNTVPLtALiaYNf
j9Nr0+6ifh6kDMenlU50+qWQ+FZHnRCaQFPBgcL1lBmfrZVq/oHy55nvMaP0YEwGRM+GNjzHtVmQ
qh9L76YTz34WL75fgJt+7NDlu5Y0YiW+nXnSHwntHEAhbcOqwUJ+5N6R84evSfmC3LQnfHwEAx8/
/x0pkJZJMXwNkGCKN7c0ZjBact9FLHXPKcCa4SPeCgTVKReghGEyBQ6sNM689aLqKhpAVpw/JwaC
6ECSDrh9RQlwEvMCiNU9N2JAToCxT6hLgFtU+SKG2FNh1dTbUM2ZYFmIn9rBGcVQnNLYGzCMx8cf
HTWFwUFjr3+kQ1Bj4RATEaFnBQO1Z6jdGBRHgSQS1GFbtvmhIhD+LWiAsySTAkbA/b9syADvaA9R
3FO2+ea3ECUHt/V9w2q0AWul4V0jx1tsrdWpWltMCOrA99XoxyyWfDPg/+kSTBzfTy4dSWzxXQlE
IN3yBo49DH34MQ9dTNARP6LMUfd+lpWrcG1ZCSNaRO9VkIsdtZIaoG3P2V1iBKBvj47Toj0cxtrz
kiQeHyD6NCVw+CKcsZzaau4yTo7dSlAzSBCWgNRtg1Astd7i61+0Ib4RQ5eTFnhSXUvLCxyWI8D2
DSo1KqmM8fAr7mBOlLn36tFiKN3wmSVqQqLVz8m+P4kbzKW0O2taFXjnL36GM6A1bHGaWC/WtxBZ
ZCWSDGB4k8H1QoQZ1NhbB9GQVHKr2TxLOGAl8H9z0qgjqswL3eajFIrNs/bS6FqApSmQsX9p5l5+
9YdepjZB3DJOYKa3UeR1YCdbWTaOL1J/ruGuRC2wvpP9K814aVdG2BYZX2kYfCuvQP+yx6YFprRg
Xk0dNaE6gi2OejZVqwOoQdZMHlPM6axYCZRXs7Y2vcvTSqnkdFaJnETg9ivtEJ9d2ev0mzIdAOml
EgUg50z9L5SodTeZy4rxmwJNMOxraGsmOFaR7n5Db2bYcDOCR/aJwYJaMT0VvzcXEzl9vtYNMyFQ
nPLdSSwFuuuupyKJG+CR1PxgXM5gpgfj219tVPQZKhTyH6wKju9QgSsQgP1EH+IwHeoPzOOFI3Wf
15y8hsdFddrk4o+odVXdw604BWU2+60Ew7PfNoKyjIsQkIRcmIJCSCiipTPEEXkRGr+F04Cktm1l
B/FkVqMG4x5Qxw/OjMh1/viSldBgagvzMGsbWmwpzezrftqHaIUqsY+BgpHG94QEwgg4PjBknMZb
kbV/8XS2JkU621AsthKMVnnAqVHy7MLZV5vO4OSMzR9PrzBDcUPsg6mxAQ2B/xXqy/WC6kKHGlrE
NcaToXdKBTpHvEVvdgR9xUMNDqAJF83TXOxemsD8+/3U+r4dLos9b2i0zxUh2FAqHsHBL7bzNeIO
4Gn5CpEclskgF5phdnQIWbH4ospGY880ceYg4/feC7urJOYHmmfMSFvNzeCGjO+poROyoilP1SNH
BKVMk+/1vptIbei/i1VQ8pbNsZcr+GCkvHiLrJgLq+kXNyyvUe6sDInDGmmQQgB8slkZzKZxRtpE
FIvzAIaWlM2wllrQnOGS3hL6krjXXozP4StZWWH3kE26wbKgvDFhBqqcrdYYWyySa2Zv9XNmshhY
d0LlhNtXSPEHb9Umzbr5sKVjRoositjHvzVZI4GC6u6IH7dfFif7Wuw/vg4XnP24fe9CRCeSiUBK
Xm3KQ40FumP/MvFVQVrrfWB46xcHtSA9gJKpt06p4EPA0/BnxWZO/9EGETe9VCNti08wcwrV7yXQ
mLGbVJhfPd2sKwge9gHsFu6UjFYs0hTIdBUsX0vDy8wr55jI55+aAKd6dZrD8/eK+7mHumWRCaWE
Na5WhkPGgTwutQm09AMgUY5XUu0bBwtVNFvmBHBlIsB5zi3Zo1EE/FA7OJKlzYpb2EBFbt0D5+RK
XZY6YvrHRfLh5tVtGVwuWOWpjZZdWs0hEQhrIEDSDncuKpH5QPcF1E43gaJ7afkB2i1TlWBNYOQ7
cQRLJHjdFltyPJaazO392xMp9ZNm4szvk1MztKVcWX+nzgni6mBJctqR8vCNa9Ok9HDS7b+QBzt9
+EfNKxsGQzSPVZRzv6dVzgpChTa6nYw8GXxP9kKUNMb9Z8nw/2wPEpsaBAkBCDsjN1VjMn/HNUlT
SHJ3RemKhWBrcqYHh33q4VKDA7WkymrEkrGxt2AAjzEMfkPJrgR9RY2vkqiS1d9NinKkG7vqTVLZ
P1jeM3yu8prLIFk1D1OiQsTHu8Zgoaio3Sh9tbG9wtlNfk+fJl0wEOkr4j6hN5/Q2ypJZnANXmI1
/iC/lniBB8M0W0Vim1NJDBGB4QG5uyRgwlVvn4CUz4I4tJHCCwHShE8GUbPaapAdY+w6UtCefIJk
9MaYKoeyLCp/IN7OPtDaS4eMKxv5DHskh7tTLk6CGOqcCMJr4n9lRsiod1qYyqr19mZqXAOi/4wO
KMjsT/Yjy0T1Q6XP2Pp6TqwF0wbhqDtNv9Tgg41gSdWxs98sfbhuW/X6qPv39kIr6RwfazWWZqnR
rEiExPKpUfzDYfV6lsmvUrwQHEbsp7DtYAQm9YlNsFUPrJU8wWdys0B+CnbAz0SVAtHkPd462Ett
h2hQdr7+9ffMyXQYy7/Zou96581SfJqFA1eGP2q6eadx5sKIpm8rlTQkOAfMqdZTEhBWpLGj+pnz
widMCBVpJsJELaeeDjn3/P4+k96Fg58SxG71BC5wfEdp9un/ygVB3lrp+GRAQvZm1NEo/7AYktUn
hCcqpzhQo2bJMhrPmfjoWI4fKGm6Obb1ck/y/q99Um3962Q2KSgzEO88peUIQ0S5zQ7Us68vF8UH
rVWRqnaOjS7PcKt6xFR9jJcAxoSaT+xU4SdioPLfogyCqMQl4DdXmoI2NPKGZfNbHfTyEK408Zvv
9G59HY6umxnG/1f2sdAvrpIwg6mCqQd6kEibM1FZc47+PIu/2WbZ79UgaGDwdFxRiNuJLyGwEiYH
DRrZ+8MPIzT/nNiK21DVc9pF5onm49kS3FdnXLHQCTE7mMoFNzVVVB4Z/W+KT+JxzQQ3N9aO+DRo
WY/dpkg0xBznpgDJJ8F4jR7gJaNy2hiKo+2LZ+4XLzhewcESLA1H8LnpIoTFOrh9wWObXaxXy/VO
TBi8IKe40Mu8krHLFfMa1mFjj6P5Fl5doc8ZbKige3fZ53uLqxVi68ab8ruoSiKuHTEY4fANxvax
HE15df68k4j36x0kGqQHpKHcQ4GIIwTSmUJxg/eVde/0ObIw3IAectXLx1Iigb95fsTVA+AXuH4c
eByGMDRk35OpTS8S4pWB6v2ZeN6AoLU/o++gnyGqrYMHZPW+8VbDA29i5zoYdfYke2kHSGAA8CiQ
L5IFzvjHF+dQhYlZPKP+aNwa8cVzRQNxF/YVEfdzhuJKBoSOY5Y5JBJHgUBnAXLPnmmUMtA8t88a
iTtOhQPq+H4CYE49bTYHrMxCTgKZ5yrSa+l4fk3AEDlpIAKls95GpU4TSLO+BMMfI1Pm8+mF7zXs
jmA3A6WDf6TkH7oU9+TcaytevFvMckDnm8R3nIaci+CbCWmomrv+mqbgVS7haq5+lj5D639msnb/
eGEHzV7bIiZGmfgH20J917JVETLWc6qYXlwwo8bzIW7AodWKjsgj1XnXj+MY/4j3ThgOipntlXbc
bLyL9dW0SbOLD/Kwbu1SiOMS5ucqXU0SPh2VrHRsu/19sdj13+Cd2T16BkmQAz1pUCd90KajkCUe
EX5aIrCnexzFJxfHteD0VCSZhAnqWb39bhF9ToEiQOpNoCMnR5jBXfDUd8wKZWQWAGdW1T27iurw
lJEiIeWwprcmA1aEMFqMP1WYvyHaPE5kIBgYHpBuyGkGrDusT61ce9zJFDAnkp+AUrJJdIGqXS41
nNsDzFSizvTdCj+kZfFM/LOCbJgv3Fh9AqfCEqkJlZarUXjoDI8b4SDVrM+fLUJuncYeoTe8sMAP
b3DwEmVqK6rpweqLojDzqEdwNa6IshmPF1lBB/+HOcla/YX+Dy99TgfIs6pBeNlb3ZmCvNqsFPjJ
raoJSti4eJZQNlJ2ZEYzXoyuGw/DTLacxXUZ6F3oqHfd4sqonlHx9H4C9YizPQuHPnIz7fSt2CBV
Y4wfAGNJ3lV5b07SvG3VL7vBlaoNWalWtAXHo8SMSDDnUu+2Jp/cySwDwG9MkT9i2Elmc8JlGy4D
tLb2ew6KTdX9FtNtJCHv/niHdVAyrUKGEJanoZMTelw1p2PjoeUqu3Efiq6GyEqCI+9W6wjLrk92
1SKY++5L+iZfUQ27kofxTUwWcIO1bK0qnX/hpbNS3XwylhUKhu6tTNYc1OuIrHcJR+s3X6EODpdS
wNbLdBKH6JXfrO6p96+2uE9OcUJ17ox7wUUqiCktMwB8W4M+uHxKfIwdpTndjbiGTYOU/w/j3jFF
x1sxnQ/EBT2ruHw2NQ7+tGGDdA9t4rFCfLwZHpowYceTc6pRJmQg8rDZT5tnmS+r4SIRMfydIabR
cl8ZQyxhP9RSWorWirOv6w5fZDHWwSMlMoaYh/QVJFx+PdakT0AZJoVuSILqsB2ACc0/CHvR66qa
Zki9fzykxG+sIG8sfko5UdXwAd1+dJtaoCeUn6e5i4h87MPgLyJE582a6OlWK6Hz0cGQjso+NJln
TO0gxBY39F81g0MmHmhT8ereUo+hQrp93e2KwTZWjM6Ck+U4LWIuo0m5Jcumdr7VirH3LmrfpUST
DM1cruuvBOhjhGJzWWxuQGfOkYF/YDIJ1RyPdn9nQvupTHo+3Rr3W9Rl2UK9V+s4iv+kogrQVUyg
VchUgbf7oEQenmblmRPnwV+5ar50D28vC4gK5F2G0DJKmbEA3eBWEW6yNxK4mnzEwZi4hc7Vhd90
iGGoRiZ8xKUB6V0DEQPwiSV4QrswAAl/TrBfN3j8vIz4zftfUQKyu7OMN5HTckvM1RtmKMVOceXS
GL988G8uiHNpcr9G0IX5zVpQzxg7qeXzGYAOdeH6jH9r8RlbTSFTMV2KDYQEpf0CQJDRZunS0Cjq
qSeWDqNC+LlNazIIeF+d8rYihlggrkpl55Jd2fZL1Lkipv+uzpgmb8haienIvLBUno0oQxeE+HQo
HhGAWPWreP7KHUVAbjIBawdNFQWTTVPQ8P833cbtOjIHKOxFR4sc6ZdBcMDSxWFYMCHS7snH0J8L
bDyEtyR8TyVwN+8BSLSQKRXcrR18blIwigodPNj40b9KLtvyQfM0I0Cwdvs5BtJtcgbumFXDtfsp
J7fn2Qqm5LXXUsb1usEbRE256Z3OAiYG5hY0T0/6L/iBYI2NLMtqNk8Iz59HR8Xtt1ScCeFuWrHX
QXwNTybYwz0giFO/NlG0LMePCnC111mU0Pkhm+7/iRyN46fJ9PTP5EApJsxgOeusP3ZbtF45N0D/
+6Gtfn1rywXKtQ2nF9jT2ptwugS+gb6FRNgH1UHnKsEL0CwpDKY9vZuZagyrnkluNwCVFfiWDD+q
VA8ylvEAri9HkalaQVG/LXU7c+ohQRvBPURpPQOlZZHAtnhh0J0l/KgceMjvV7G5pKRPHJFS9hHT
EW9h5cahSVup6V6vB6yGvnN8STDMt0vFagJAT6UhCen7aQeuKsSnXwbvU/ravlmqnKl3CKpfsLFd
AJleqE/yQzq8DECTflO0x8lSiILH1+rjsdWCQbo7NKfa3X69PQlW1cNwPUwXnaXcGqyrpO6nkr85
r5bSG0l0s0aTUtZs3kABUNz06JqbPGw9U9SwFVV8aYbtn8S6iZjokgqjLLXIdI1FdW0E1PRc2GFA
udyxtTTOKJzwfELpI1TiFQmF14W03Mdf+f0rwbFgvW3W6vD1rU6dPjUQuV/RtQgzTyG6GhjTFdxj
C6LxNq//l8SYqR/qwNUnQLhAruR1ButtvdfpYQ3SPtrhlD23rnKMSN3mB1JU+T8/JbcD+v7LMOoY
qFUwLKpScpxwPXdJ4eKnFh1/Gpq4nurxUeSkckOOqHc9d9e+tA3ZZOvybnnLBrVssBw07qGkQjAr
Vy6EDIR7A6qSfPq1WHRxMSprb1oVHhXCLqtqSgKNK0vvb7wye94C+15ZAh7R/CIxpeFLO8O5/fhc
qhTiq1tK7BGfFG379qCpHHaNHdQu1ja0hJhg0J0ohhy1Bp+n9kRp1OTxT3AVxnI25q6DMaqTW4QE
r0GpSl0sYYanXwGoHZXSLW9gxoH+Sr81ix+YITJ3yetTxW0WPuLO4WEgwK0EjdYP2f0k/yNks5qe
jKsYD3G/U5zS9lNateKBMC5FdpioIRXUlazhy2K82ymfIk0bKzrO2tm/63k3Pq+W5+Xc1obvLZk6
NgVWO68piGQfyRKP7ubygIZ6gp/ZUcB719PE/k8tJ59eX8AAyGsIYi4dAIN1H4ztkOOj4uEiDkf7
S8ZP9v0bOusCzEdJEp/2eoQE27nC+6fXSC0JrS1tKtNkeooLKwaVst6r5CidMIEFYBrPp03cxrP2
sWiemggZ1Be8MmdFt4vlZeyM/Bu9YSpvZV2Yyv/vnTYR/hMBDq9sZJY9Mk0vev65mFlMeE1BxoPg
2I8pmosC02ITOj4aSTmtMp0gdoeNETxAkDCgP6XQ5qLYdWv06xc4fSa9NuUDHzrihRVkUxwAhdKf
gQyfsvAa5Qd1fSlE0BJV1xGNmQJcY5huVapyqK/zYTNCZHlSLYs8+62BV/lbmRX28BtBLAmvYtJo
mXz+vTUKuEEIKXnyKtM1SBHRZ+YnWCm6VAdp39FonyjJUv/k4vmIcHFu8P2jn8+hgEZwp3kKhr40
RnXdVYK0OV5aU+CmuWG7jbvAyR5X+XKZMymZ/enHPZPDHp43NZLbfhaABdIG9wTTDCdRaL+7UNhE
3+ZNc7v6Nfdo/TaFdHVxlqiNUTmFbyeGetFrQlOw332Yvty0UXqaUwL/m0ocM2hTYvHJNY6ZVogI
YTKLDWEQcEGhWMhBAp1BBAWVjBWloUP7fx0YYmH3twVhtIUz4MKw8qUaAhexVs5YlHrxk385NkNZ
skVFgepPHj8eTZBx+qswhMh3sbVdCLNTi4jYUGd1gm1DGLDUvjpkZalZgB4+7EyYTheIeXXTDUPW
a+JcC11S7b9UoS3WeS2QoCQMeSSh6LZ4fgQcQ7euViTGHEORI47YNxjwFAN+JRyxt6bJhxFqtx2Z
npdE7Bz/B1UnQcD/AAIqMQ8KAU6ytfJQ9qzfOltEgLZcy1EeQvxyLvp1QwnZAk0r37Ic3AnzEvYB
dNMtAJZnE551gMmLeWZjSpvbmKquZK3VJ7G0WRCd4ReyelInTYC9u4S091tcnd9g+pFuUdlp/hrP
+LhV12kIKO2HRo6CKx5pOnwGyk7Y2XGC7O1Apq68+0qUowW+ohAS4mi++bP+eoNMHY4QaWBeJYhS
dEeNgjccD9PFQMTnJ7GTJDUGS0kqyld8V3a0/Dh7PVeuJ2cEqZ+Mg+0cXAffLdNsJcyN88TBDqm9
QJrkpi6kgIiBrazuup7ZdGL7ON6pq5GrbF7b8QGX1AYN3id/S0pjtLBEXoBG3K1tuFsWEzYMnRdU
HypXsVPGaKZ8QVhtslwMqg8+U+kBkbX/simJsOjrUkKkIeDLhSqvKGVFeNp1n/u2Izxx8GbvNs3I
j5J0Oj58XPVOf1cfpqRlwX+Z1zaZHR5Cb/CT5XRFsQN8/hO33r/tN6HIPYEYtP/PALcsu8YW9PXk
AzT+zaqmE8lM+5JBelg1rasMUKzAsuuj7hxnecisixkXZaIeoMDXod3BkUGcXQY4FDGVs6/oHsDi
xHyWLiTax7YXhd1UJ+t14pbEHPKLC4R7NNZT65ulCmZQA8U5MDXnvE7/S8BpZYigWlpd6Yfj6h9a
IElHqzajeSz+ZPEX1omnu2n8kygi8BunbToX4DN1HWStZPXtG0FgiEdKXNPK2AQDN299REnjfKyr
hsi0WD9HdiPKILAWfVYDx9+zOLw0Ls8RCffYOFkndF4FiaPMAHxAujSaoBW2S0AE8Wf2AMr/zd9o
lnj2HyIp/aUx+rpnMQhwvFAH5Z7hd9urwfV8vV+M9g19p8UguUmrc+BGiJliAIGTb4pl2udDxT/3
AjSgvJpwHV2146J8me2DrUFZ4jdxt/hxcH6ept4NbqrvQordapX9BJky9ZFcCutnzLz5Xr5G/6TN
V7TLOziG3rfnwQKzeTlZLgDp3KPGUingVs1XQujJKLmaOXkfNxacFJUWxS6lPC/+njVx8LGqvo5G
YXG7l8/S1/lM8DvmN7TY3kqVE6sIJ8P2ab4upuivy22wX7iqefCEm46KKFP9QzzbnGQtSSFYWihy
HnGpgm+eR2IeTeRG06g3iyWvlpDWjdmDzjdu25cRFZWkY0Zwp22sl2q7sunlV4zu5dtUfaNtSi0d
PlN6O06IWx8gGawq3W/8sjs0a03K3r1KqPCFF8zdtPKGZUN5259tDmNvmkayYp56zhXUeyH3ZERX
dudTwUxKrw20PiJFUuGsuYjSLsv/ww2pK5uqDzwlY1WQy/OIKkppd1Ols303BnsHO5nqmAhf96fk
zQZLgho0fdwAU4yVlXTXcbyL/y/XehTEUUDOKPr+mtcONwCUv9xO41h/UJi00dudaM8ZPXIffYE5
xG968GWt8bBfZSvtJ5OfYXwfYw0p8q4wjZLeQsBlIFi6PuqimvDwAvJsBUv7xXKyud4iodcJV6og
zTlKUzvgyHF4TFOmlkzwKBe0EMder9cG6xXEshZx6wycrycvw5R4s0NODudAtTpO2YNMpVjIlPNJ
4U4rkUmQ/pkNNJvBO2LpiteMOGJ0z4AF+a4NOA9FM9D7Ixj5LXz705ZsW8okxrGg7++M2pmVzMK1
V3vRCWt7Ai03L+3QUZ05UbH2+kTz2soahDbgMQNqBCPjBjKvHXKFY4OABMG05a/1hKxH3fUCjanl
Mh6i5EPhW9lrzc5uOfVfVruNouaovPmovYm/FuQx5BI0MWAtK5bssAodQMDHPRfUkEQfSpkXelVu
bVkOZyFSpAIUVKuKm829NGvovlFGFV1xvuJsn49KdLP+FIdO9Sh4R3ZlZ7woptshv9QcQfRUgxNU
GQVFDThJVwFgzG8i09Rvaa54oixrhYQOwNWyPl54D9SpvN5UpKqsuhIRUpF+jvv4Z1NdnTPE6/J+
eUo45e+a4UOmbwvOiyeqNTjZTAOKMpzlxxPVUdW2Cd0DwDPbjxGXfHisy2Hacq2C9oQPZNoEN1Az
xX0z32wU0T6qDSzogQwR73IEVN2lN2FFOrVYaqQ2U/oOUW6pqKJrvg5BOU6M8p8/ES4KVOaqTgWP
IBk+gRHIj6hWBi00Xmqh7qPLDSjLliyAF6eXBWXKUDvOUqH5AmwqhNbBuULIN3ldaid47AErRnP7
eQvOernCa31FndzanceDYFO8fJ6fPkudq+/KKt089eSQWs9zX3dgzy68tZx6oKW2Hb7FIK9RkvTq
eTi4sFqz8OQCfQ+YCu4Vb9P3cNxgQDv38W1l/WdUkQF7y9xZWHnneaZvcTHnesJKeCpED+IsXCEo
bTTvoQcUMdappk5sb946XeiFDQ21NLOfiJd9tjvJxJ2BG8Grfu8cCT78M35Xp3vHjp0GXAfWa8Jm
X+mOETqh3P4yEE/6Go/YQCZVwcr4ZarWapXJ7Jhhmc17Eie1/sUfhPTy3m0/fnKTYSkdLMnEU895
z6775VL5ix8pGdVsNjKe17vlpPNDJPLm/xeUpFDrPklwhJ1f6uLdJLJhqhA0NEYTQaXvTSZytRJA
n7EVu2g4SFFLKNKOtc9vQ/yrNXgOQo/Alx9iTaRCkBmp80s5EWGIJ3K7Q7tp+A9bEd+xtr6HG+uD
LJnqCaTvbv/I/Uiii9qGCDooLlkgUJnka0z+U4sg3RHSZcsuXhzxx2oCF0FGwF7V7NIyFx2HBE1A
0JCfd5xlErWGKxpzIz24+VUJQpPfZuCL1rV+5teFar1zvFSgHKgzDon/GLOC35m9pZMx1dwWMWge
CgPU8SGefrZGlsvb/938rV6xUi4uu8JersIgdt6ggajq+hE4H7ljdDuS3BM1CwOYvcCI+0S/AFfr
ta0+qGNK/zrMp3bdndL21fKg74S09XzT69ku5CcCw+B4cw3rsa6ynhTQX+FhLJHEbBWuNB1TdV0i
Z3Krem2Jz+GEKnZVJIxSiZXKvPvND91hA4ogMDJ/t8uaoWpvVaWzWdBRl77Sht7DFC5kpda1o2bd
lwM02Pe3omccUz9IbIhqvq5Z94Bclah79VH4SjH0tWuwhF49RVb/mhZ8S4WfYZ9DS+OjFnwBbo2V
Ay+i9NMrF5kr1Bi1pGq7byvX9aBDN/tjIzvYqnBJceV4JnDlwOg6y6jNYMQjJ0kXByEtOoWh8iOc
oq+ZW1FEcywRxopJDmvmPSh+yor4pSPtPPM5x2XXaEaofz/hr4XRzFOezm/PzGdRf7ugkLhs33D2
bLVtLVS8FKpcQN9dj3eDagCiDVX2IZoSK3BUqsDNzahQd4GRBOZsp/chR8D+Iv7FUqDpHxg9nzkc
fMea/4T+JwjfHnoNP3CpLmC9ke1BclMk6Gn2L1EDPp4HC/jpUjJOG8B/1kcP91qK4/JQPpQ5YHOi
P0BqlwbYL+sYlW7ts8mQSgwys6vLYBiRYqjVL6U6PcRETm36Zft+UJAUQ/fJfz+9NqiQvdUJe5Tb
/ZKE7CET39QEd3NKvgA/686EfRTucJJtJV7DEhqjKGF3u8aCck2lC2VUnEPv0E4O1iVJO9T4VhEg
sE0d3O0EnH6vLeELfCM5nXXxpbLO0RJbJONC5m4Ct5eVcM3aKF7iBWPxl/YVh0VMWDTFmJQob1Db
ac5JaCIY6XhnPyLCI0m2GZHEyNcx1YHSP0avw6BndmXFTMUPFkp3sdLwfXfBhyUOmeo8PD9josEr
Dg0JOn1GL2kaHTS+h9VzQpMhflSYGT89vGmAupjYgxdlB6Zgbif3L3h91c+UsG7Ce0Bb9lUI3E7e
xiSPxSIZiyfRw8OVOvt/rXeRi0mSosffKEBlLl8MDmqzvtUPwM0lJSVrBL3Ti1YnZaIZ30cwn040
LSimFfbuVwdg2jvlgw8C7D20XYw88G8RNX4b+6YqrIBzMtQ0OQSDkeTDJlxnsjacwHag2mpEE0mI
jpBR6wHQ/+92oXNoYp2ng5v4N511LxclMTQqHo1WFBVV9cX4gPCwKBdS/nKfBoY674s6vODf9GQu
Hxx3XmJ4Fsls0dlfaiOGv4lpNDDY0OliAiJPl79ZFpU34SsZKoXBA4baV6zXgu0nWf64Wg3VJIqn
Yn6t/J5ojybwFWdGce5ANEMv9z1BaFLe2eDMJMMsJybq0YuKVGoNfMVro3+loFXCgSXTPC9eu70c
WWF2bbcBHVqYDlAGTchV/jW+8sCBGr50qSd1ka5Xw+lZeB1QN72HIkojIgc/KZuuugQz0VRIQxhu
WzNrZ9k2mhk4puViN3UWr2Wh7oSAERviNkj/X87r04snCFQpszxbLnizY3DmyLZk068cOFB6SY6/
JVg1/vop3+7TqVvpGjqMs15yuhcR8MI1VKVd3Z37J3TWAsx+qxHxCk9e29emd546upsMwGRiv7qE
A4q2pYEfY3pso3GCh8aCWzHb6LSBVCdAYiyBTVTMEzGY9gTqhMRj7jsUASQuI0Sqt9glOcbku932
m0UUzU71U+imwUEZhdT9XxXPRQxHfOAlgEWfyerXqrmWO4/CgQSMxKUbWriQmbejpdyQnMTmLuvz
9N7akp0vXtGRMEXBGjpf1PEVOFkIun/3yXAGVvL931Y5fJ7qF/MlOn+GeVM2pRr6EbxMdwuzfJzu
htmtngjH7glVLk2/2ymVnDn9UjCUucI3Bc1Nel198IrGAYkDbPYFAvkxYBq2YxXeiFpwHGa7jz9+
2td/Y/BDD1ouqjdmyavttC9acOLRzygWAgWfwM6HqbiPsA8ln5O16ak5IK/n2v0g8BZWJORdMRZy
NkTsaD9UoF6xcDmoGeq1YcLH18PlBVE6iXddPWEVfV3sr/3oDKQgHA4YG6OfsiNhaqR9szxib1FO
6GBLH9lpKelxE2w4NIf40qQUMxqQhL5NlvfxXKoC+UXms2PVvxR3XB0Yb2jxRd3Ebsez8BN6eJEy
xmwT8XcN9My/bwE5g7bYpUAmnDAtU/7kGDYNHWKkgcrpst2LvrOcNOYpdccs5sjNgWpoCJ/He0PB
20gfCjXQkQyLn/f8h8nXw57vHULNajuPon9AjzHGp6IbNlo7opHlgudpi2HtY/Xc52SxNYJp2Klh
udely+40jSPpDYJYTZqaKSZQwt6/bUkKxZfZ6ih9uAhmeE5Tv/W+f4hN01hvROlfC93vs9Bpf/X4
1NzvsVM4mytq8Hd/h3QXnRtUDSYv9lFYcrX6nFdP5FKA4ckz49OzXLGmD6OeCeXWnW4WioWIxCzv
dKryH/Xe2RgHF/Qf1M89Klba4h7mIdzbOebXsBniI+WtZpobrlxqCVG2RnCrSnhia5RblkgBXc7Y
FZm7y69oGpDbqFtLQJPttWiNtsRODLqa2IeNggs6DOW7aKDRphEaIXlDSg5//sH8pA/wRzPayT6/
dfP1Dcbf5IbUWR1qBcUMEykLxWwb4HGYQ4gAOxH/x7+hvopHhxDZ4T6q1ofaSoIhqe3AQ6HPdo6h
dEOBEfF8Zgji7dyQFTquqCZWi5qXwCIab4bklQu6UmRowqpMpFEQ2JzI74c95lmKuXZsLLkxLl0r
9o2hP+5lUyiyxoHUi8PpcMpFjO00gHlRbKRSwbAGweHVAI+c3lBeztByM3jk1SvaBodVp11stBr2
djxGrhzHbHx2rjC76FOehaPugxiyKGGHsNMFVUWI13n0PmTRgGKnXYrzWCuuaupNYSny4dSxoEX+
+Z2Zol7y5MKe55ymH7TmRVcbu9nAW+G+/QhgZhf5mRxCBx6rm8CONJbao2Pmnv6w0i/AGmVu7ALj
4GmNnzrwbuo8HFNxqXLlIRFCbDp2WS6KMudmR0yGvYGVZc4697yzCvmHXnBof6Y37U4SZrZsTGg/
vPmrgfhkrmJizWCrUa9YzDfhIOysJeFIrzcaRmGXzr34RjRxRu5osvm/WWp5RRC9bFzr3L1hOVNC
A1xV+rKnxu7NY+P8iVi+o9+TdQc0dihbC2q+fVbxYi7csATkX5MnMUVkgfmgaOrlonuWHC/b3+7u
PqFzaJ4NdMTV30JDl9i3KR70GKWqB7ZfoLccuS2qwSbW7JLlikOfVRYJfT4utflIkGmemCDuOjRV
tdTgyS7HUix8ApYrU/XnCy2eFngS/ZHr49XQ8S/4o99mwUg/VfO9bR9smwf20mTF8kAOsFxo77su
ydxvvz4cSkSX5V6vD1K6/gHNtw2LW103PHnQ+F6+kU15YngchshFp9Rf5AI3KKLYFFDG2GBuEPHQ
XLTFL7e5pKCjGbqFqytQUBD75GmU7IExz06H4sfw/MlkM7U2ncsvHL05N4chM0UQdz6vMRGsAoHt
fKQg/ie+NAvEDp3Bsgdb7RUB7E4Ks3d8BuzbawOk0w6xfi47/Ud0D3J/EB96vPNQ7xIAIp/SmJ91
6ncbDHlE+IGWEwYkBpO9mi1M4fE377e3YUZM9E8ThtiqhMNA7nVcZ+EpFKnHEtlIWUir5Qg7jvLE
XXpLSX6/6cMyR4s598gBOgF41+aPqjWc/rKbMG14SvgzlRaeG068VpYep1dSdQL6FjQCwxP89MUc
jXe0t2ZpNIKu58dhsv6qvXgZRDCpnb9wsm9wgSHa3qcOwy7QHPS+qsiv6FhbUfwIA2bMsDCV1TXP
LKgcs/IWXZAim07puW6hLHTuiS+VxfvbTJjHj6ySpie1VVQidZl4dA/rKW3WoCl1hhjIfQhZJ7sT
DVI8CLm8OoWJX8JHcL24gNRfFGd1Vut1Vn011AAIy0f9Mr9xnae3+sMslpS1c82Fyt8gddiaL5st
lCB/NphlavlLK+VF/MaDLUUMYcKjiiRE39pkhGOvRWExyP2BVkUbEmXJganhxre6e9YDd5+lMeOO
cYV9Dw91VbMOujQAhD9sIg6ZlgfJFhZYFC/7NtaSq4DWMvsmE2fjetloMY29H0NzQCfSSO00snJc
ivx9I5JP6sjkkIZUxIbRH67pbWI/UtwxfblBgb7Hj7og99sZBggpCxk2CFaB+JFXd+wHsNqhXisj
K7KV7gHIP2cJpaDgKlewzRpurPj8z1O6P8JbEsKhZByUMiG/PEqxdbFyXnFwotyYw19az38/Wtp1
z3+QNtozBu7fIN7vb8fdjq3BlQy8ilyuxFVWy3Hd8oKYKgMyvLwWBy97f8OuirAh2Kr06eAh80Ae
mUxfCLiIjQm3+hCPQwN32gFkXyJP/PlT10QLSj+O31lhb0XHhdvIdCuGErBXFu8jKDaT1UqIMcNr
EfpVt8sCa3GE0Ze5CvJwzeObyyw4tBGyyJoVG3E5aR4RoivzBpQ5Xpj3GqfNxBBXx4Qdso8ig7l0
4W0qAi6pw4bSkcvCd1Ejbhi9mC0PKt6VRFkWaRmHxDXmKyP4uCCLwJ1u2LpWH+mNMoqgJMPNgb8Q
SCOdgnfc2kZoYJABWD7iZYni0LAKP0kQBm5ENK6fmMn4E9hcUsFeBKdf0EHGWCrPrGDhZleJ1xRK
gq4ncE5u/sF4OTzq0v/lwHffUu7lmo1ftG45jdLdAzpnlR9SKWfJUg0C5UodBdyakmku40+0MVnN
tkYker+L3fz3XEaEaGcw7bBHLnxQF8mOkeST7PHEnmoVxKz3G1m3CHylIr2lqxqNu85bqZUgk2Xg
XfRrw+mmz8fJgO9xokAOHHUFOXcZLpQIrtD30bmKDP0LYiJX+ZBIms0beM0wDx8z264u2Rj2g6eu
S9dDgKWGgPyM2Bl5NDFKNxlfGmexIka1lEYcfGbjU323naiPinVGwyOEslvPl7eAGl/07Qjz4Ai4
pajRbrd9h2V4NhaZnMB10ttnjblHF5APOwzUuFYkiHMXY3H3jtapAGiFeADy3HknYmV6lBUVWL8Q
cHhZDLyOJdeJNqU/Dq04gybV6jR3OnyGsMlonJLEIKqslVvxL+7a5ZD+8UPl1NrixAfpwycmAejb
J//1iQlJvnKNceGad9E8UWSnnr3grLyWpF65Qbg2tWRSK1VYhAti5bOALQhj4InoZnBawT/4oZdM
m/edlZCWyicAI6P+ICMa4Kp9FsQLUuGdwvkS/ikjAkaBqhelRefWeEb/lbjkGYanOYI5LQRBUGJL
WmXfjJv6DYXdbDlBbgkSFcAyNJKOnOQopJPb3Aq4b2uZfK/nXq8+TFVqUqzhkCocSjp3tAEKRT2H
QWCUmuVOmwHPzr7IR73/njO7Has3rB32u4kbf69IXGVpb0L8oPru8wsNbihm4T8WPf0blAn8FacD
pvyByNNTQjY6eLlMsw5kL54E45pjwgcksM9MJk1Sajwxn2CBasPR8KQJe9/5vg+GCnvKEp9MXv8z
9l3mjxnRvSN0Nixa11DCawFGRtAnYK+pbDbb4Z8fYhN8br1vuhLcE1gfmagzjHdQ0Pmv8ZPJ7IVD
HMFVkzS7XmYMBlCH4uVU3zNuUgpK4CXMRv6XjDulqKdE079lkPTDnp2GSPW8LrRGK0qWEbZCXO7Z
vBmk1W4NwBruTJ6LFi2zGXo+NxNg93PxYHycpHeb4L9yrdtZ/uoVcpvVDRoSJO0dOFVq9YZiLlES
HXLWq34D20AD6qRlONXP9RUOgn1pKrKx9Zy031YkqcBxowEXMKZg2MdDgNSYaVWZSTjaiBIPivVW
QyXDxlijb6QwoBQ9hj2w21vJDSB3F+q6lW5T6xDr5SmXi2Odq9w3PUkYIgKdvKazrIVc/kSV60Pv
Y+Y8CL64/gBG3BmERlbUFkPAs4QD66hYaphJbFTfyPfcLmXjFg1tltlD24zER8/2l0McCD5J4m4r
e7aQn7EY//gVBA07Dh/fbf4kotBDX+nE/d+Xqt9YDqcojoJf5IwsZZb6ioctOvOMFaA5NjhYk1qI
xsV2U6vCIf/Ep+UIzAwBgWTspe4d5G/fLQEjOO4W/UVTUjPcggtZQW7DnsBeGAsUndfG4kb/05Z9
9d/XQMInEpTuf5/DQKJbjer4rGrfpZZ/y0QwULRxSGa133puBZ133iivvI/OPnvhFZQNxxykEHAR
yLSvOyTJ9/CMNfOatP0JvO2tXXD5vo84gPCwWMde052eFUnSIRe4vojBC6wEY6k3AXF6Luk8bIj5
46tu7qSxEZGJO24GN7fPu7Yk0GJgrj7dAxOINDJv/y7JL6CVBcP4kD6F0sR5aNkiJngp0kjLTrp1
C/QsLqRYM7eMujAhEi0H4sWJ7XirkRLjll5oCuz+zr6ct74ly7OhnuTNqawBBVrMgJeqJnzhl1Vf
fJY7w14KDQTID7zzJFwoMIgdPBvFvbRAr+9NVidMDVcLzR1CVnQgbL56CCZj/Y35DrgANEXEUtiH
gvgkgszY4J+Yrc3wc1O1smmgX4SBYDxfbP1MyT81hTfm4Job87d9rFy1YuknqudLnPLYOuvvk9Ac
OPSMAeNyUv6az6qp7tom20Zf0GImdqQWp2J+G+H3vp6vhByvQC33GfQt/YdlSn8hv9d3jtHTBsxd
Xj7zTlZW3qkrMJ8mM4eOrpGW5bMEvLYDSoqWht/PSoOlz9300GiUluNeiG9ojITteIEXx3Xs7TbS
UVNL3GfZhAtBzcHczUZVBFh5lBQRIo7DEYCeDZj0SrZMVfN5OMJo2bQpdMdd0+N79wyFBLUSebMX
1/RdiPdKMhZrv8N5ianRKQr+ct2lgso48Y54SIJN2jvU+X2Nmbi9hve3B11P7GxHCL4i7NzhaVBK
22LV8lXWZ/4foIWRxfzNGHTBWTOnqe5uhFk1tXnHymdlwUaVVtmW1evJg5HE0hIJmyZfC4CBiaCe
4ekn8ppmuSI6q/7wCEQi7wlCQC4cQEkBVcYdi8pj9PSiUhBQzqJXJ1u4lcq/Z2kLoSXePmzpvbDH
y4nEqujcCa/i+pvHb809xPtyMicNfTIanKwggv7C+FrVyEdVO2ykp+mxNJuIi2Xed5vPhCL7NUfN
34vU9LEZnvcOXnD860fFTZB0K2sjNYxr1o8X/lbkzqgUp+jw1hHEqChUkZ0Ayi6+NjDLLtPEEz/O
BzbrN6UazwlKpUqRgWAkGV2SpKpSoxGxCa9GTPpRLhTt3DbPcs1Lp6FmFATD47tslomLFcFEvF4d
LH/oIc+WZu3+NbVeGAbrLwz9DZlvdPABlj8xua59+t0CRMclJQAMn7TpNvvpYFLhAVogoO9OksIm
ALGuxulNbwRUV+1b1MPeVxw2kEBZQMH6WzDzhXzd8JQwPJVXBTGHn+dWGnrMCg6rdqECxmbQK0cO
JDyZ8GdAoJnX9UCct/l4S65AhtybCFCa1ATLz3Di7t2hmdiI7TihtsUAA4twF1SxNt2ViOTh1bp8
F2Th8xVbWV/fDCTTeYDkkR3kCp1UzdwY3w9wXGZBLNOmqG4FnXW+Yj5NjBBxFHvmbzA/B/7ngGOL
w8qEyVAkc2/wpBQ1rQoawShz5QH+OlU9rRlxMd4oSYF1E8kCQvfWry7bMJb8ZiD+HLZnu6+8TLdQ
FL3KPpADVM1f/55RSktG6I1t5EPpu4/CXORncG6z1NQcFBqnuVYKt3en+3/KGye1Ze2GpWidSSwY
uhzlewhbXk/uAQsc56m8lbC4TgP/eHUGISaTbXLPzh4I9TNgpEHBrIKcygPNr7VJYBCXIpqCtQk6
f0hPSDDBEdQokznfKemzF4BINnGDxi4yEoTsL/Y0DJYDFxGtOUQ6twkkhBB7gGz4SebBZll6FbFV
lZgv5iwevQfPaM1FDWdtiO8ehkRkAnVhDwMbbBtQiScewdL9J+P6LUkd0k3Yfy9MsGmXUIzvhRjG
8qz2kWLEl6WBDL3lx35cWfqGYPGaQ3Pou0U24ZgoXUjcwr3K41pP2kpFCV9pTkSAk6+nHKtmovzt
ffHU63TdG87v5b1lLCK2ByWdmBXjwOFn56vdD4WBxNy9l5l+R1MlZ28JKR+ksBSHpRVeYRxzH2aP
YKYGddInFtuh6soQSoVjFzQLZlLw3yEhgEsr9IoQZZzHdk7aVUoiH9fOxml04M3YGWksnK6yoS+g
BiiYV/zvsstdnv7/zqvwlgRNxFdNw38Za2Mh4h3bbUJIqFl57ecYCbZcoaEMfSW2d/eUYBcRcUa1
ruItjYQKGQDShmZxQUTyEKJMUts+iKgznh5+iil3nBKcVqyOl3gRF/eRagC57pRmlzHhf3RegKNV
h3Jg5fqS/MBSyyQeQgkqbkgPBVx72yuUoUPApOKQz7ZGcpdVjhPmi5kFr/rdwX/7YVVvoj0va55V
59KrYiqTypAuwSUFdQRPM7uhLeXOy0aKvE9RwLhN7l6DQvUAtyHx1t+S5D1OpzZAAfd8SxeMwRP/
iIIMJYUMtpRo9QPa1dL9qJ4ehzb2DTye6/njmUPG9RX5EMeZXsT5+gsnmeejgxSVhv6xUxbUDsrp
VTu/JCSRjnyZHdssVdjGiLpDXZd49M39nfjh6c/CVGxxVlTCJ+cqpSdjtzsjRSFZaEt0SFZF1grZ
aVi7kktjgZe2l6y3J0ncUL8oZiNp/qF6T8Q/0HmwFHpr5Ji3VVd8f3dZxWuzwS3IOSu03hwf4A9T
oatl3vW0y4BeZEoHlWGkS9Er+XNkWe+nlPUE9JUSu+sOZ9jKBqY4VVTsnzHSQCd86U/CO4t9CH0B
HqPcQIYoqu2sqXAGfziHiHAJ4KJqyiMtm18c0fr9gtOfUrzp1ZQE4/HCFScpYW1ZB0IJBuD2teLv
GZB2lo4Qy98zndiUMXLZRyqjr/KBE4hYzrNt+YzwXXUq3Uw+K/F/zeU+4WRQyS/rFGChCPSCxYw1
SCjiDEZCL8RwaQmdUEo6Yfg2XECX81+pOR9SLvUJEwtx9bahflLxXMhCPyCVcme6D25Ua5K2cspq
Zq00ckiVUXS4iDmnBEDtn0CJjQgNGlYGZO1wLIK+zw/bcv6PUqWN6itH2OZOdCFuwffWO8JOxWQ/
YtL7OaPxMYYFRG8zjOlBz9cQ5LHddJLdkFV+A0h3Ns/q5lGxQCY2U8bu4Wipbor5v3mAwIbmVavm
C/y3w0WH+3b3eco9biD8Z6hS3QTr2KPlIV+lfOn/Oo6SjvuSbV3+SrDo6CABXGdGcHKbS6d1TD7m
KGVpyP6/QzjXPaQe5w/lTflJfJjrHscvy5Hj6wrHtbvMJt7op0pmhD7okOkVjoNNvoQqnG3uYR6W
/C5Hw9xplJR0kVfoMTwqJMNGyYa42vppZYlD1Cyl5r45I6jcQgiHhSNgnMASjUL7CP1+W3BL77kg
NeJMPrpTNH1XNJD+qOv541/0oYvniv+5jerGfMMaBKk0+zhHe5tfxJMYlI6IdnPeEhtjyZ28HBts
GbywaAyKYLj4swV3o8z2KOza8Jd+v8hnB8gQhLBJNd8gYuIWvst65ozi3hreEVWvIUwwIficvCpk
K2N97eXDvuJ221xZslRezLZ4s6H994P05ndVYJvc0OsDfHb13jS0kjYbGNbDZo0w7CJPRIX5OZLb
cl8+soJuiBou+5z7NxUDEnVvlvFJBN4q/V+OXI2M6R9zIkaCCSZoR0sgXyT3Tk1ok3RDd+uzY142
dg/A+FsqY8avomcJVVtF3G7alnnarDyKbK8uFqgflXohOGpMVj10FV1v/TKlGSy0SFpPZ1xjyNyO
KyQukAmq5v3s8CcEL1DbytXRbE9cGyme/vttNFP4RMsT0w7VF9kg530XobA2fAcGW1aIipHa66bw
qfdLwucI1zdcqeJgZRp6BiLMuF2hkSl6K9bblhahUo2ynvrhKqRYGSj+Twu+tsqTlUtJutzwe1vy
3zuHp+c+ciRoOWpeL5Yl7CDYLskcciTHRxZSWEF7QHI6hPbUPYKGEY82LoczJ8nzuL2lpUJJzvjs
IHLnBE5wFT9b7wQ8qXC7Af24a7mi+gktUKyydFwSlRtQUlM9uJo8bwe1pNNZQVEqMjezid/z0sLA
/U7T6bxf103HUGz67TItj9OzlGC/Dv2lnupqPJzjdCzrpNu6YgaUw/VIhs9zZut/5wEuprLKV/r1
4nuWRUDHt3Wkl2wSw0MZV8NHZy8LM7NGhyr17ZKwE6fRVZnyqgV5o0eRZ1F9mDHlAUcCuLvJk4qy
eHuLB3YZWTFjZ+Ht4KAP5TEfLMjm66Ls8y1CBH6Zf6foOURLM8GSU1FSeJkHCDN2wBq3BrpHbx7p
e0hSe1sZ1wgN2qzpbsW/MkicYqeMxwisVQEXm4PXg5muGVYUi+Kywlcgvo6E6Yl4U2ELD+SNgjn/
CCuyU4ozqsoWohCEdNWsfLx81isSHjPIX8qrbNWy884nBdiP/pAFmWXcP0n8WCVYKL/iZrrzYGGT
lSnioHvmyQrDvhNnurRguPXf8+KU2AIceAlk21za6WZeNTEmlYw1ISvKts4RsdNxVHT4e8gLWO6x
fFqORpBRh1WSBOexZcMUfSRjCTpVezmswZCRIDFB/wo+mvS9dbv59OdF0h9ISMQEcjid45+9Qi6e
mj8rg/yBYuW0065wlYwHlg/sPIr184Q5zGNK8JZcM+4N8z1R+Ngyy3Y2oc56D3yv7kmPey3O+R9K
b36sKiXye98gLdq7WiozxlXpw5Kbzpa5cE46MEbGoWlFsblKWCakeqGtG1UVnvvNGA2l54Lh5Eu1
ATZx1ZX2F0WZhv0LSVoUSPAwWEVxJLMQkgFZPOmct2CROye65h9EMx1Q/KeLOSZlkLQVlX7++Kdd
VHbGqMWn38g2O6n/hZohib7OTEzkBDU6a4Duutpkb/Rbf0MhFlbBTSCMup94QBmJ0V//jFrjdtae
SoTYEBxMspgchNpUAZPJFctYnHfL7kTBzB5BFmftaR2hVh5TxoExf/15XDzh+Lzwvi3/NkPnx4b2
CSYe/s6CJgX9r57YBk0U6FpnrovDWwXzX0+q/O3+tYOZhvNzk85JU8YxRMfq+DiXXuE6n80t2+lY
Pvs06lfI4AW8MapZ4l7Ufh3cOshKjYnfQsnJQ42SclxY5ainhjKa1BnHqV31OKGl0eYTJPZcEHY+
nnWU7qDw+zFlO5kQGNO3foqAAlJcm4OwiYoHmh+3Rsydut0ZcDBvMRnIuUnD5v6KLeoI24JAzYge
kDDc0wSbGdeVi0L4vrgAEmO3WDTK9+lWhr35EDo9zcNOsRW0oa617wmFI9n+BMYkjyORFnPHcSrp
O7FVAKYX/yjv34tWFNTwPfynzdLF5MfgylZ0gXnVndcrv8dXTIc9/eDAiA+X5MysroF9/evcs9UV
1TnYU25yIOAzH03rX57eULVMrZ7mZ6IJcayhHe6VPLalXbVN3J+8YvGp5mJ0ZEVfTBSQIgJswGck
7cKJuUT0kvACcgxQf/sbJ5whYfF+y/JhVATrIT20swJW6HtPHHK6o6eJJkqUaDLaJMIK/x/ivi9j
hzdVakQPimANuqfNhsqMZwc17JPmQTLqja0D7WShJtuhoSOze5iqZ66+2EQC/2Wu+1A3L4/sEwhl
b5bS8Pss8vzFFjFFBDpHVy6dS42obXDco8s4fZLRYUuKJ3uLnCFzKJnTxTPhbST124hKfDH/9kOj
nQW6Jk3YLcNmK56yLDxqaXXqGpxsRgYZVyu8alpX3/wlstoiy6kL/MkIhxZhYuVFMsCmfp1mpSaV
ckP0IU3RaT+GGhdlaXVtuF+BZmX0StPfROeUPcgZqi+fOZfAlp9lbBYMid3cPjU8Coe0qx+JMbfZ
YAY+CNWQpBw6rQAzAPURFo9rzKI4z0ULipMrTLC8/bGgaG5TrPL+StymJVopFv6eENwPP0JNVjBc
i6fqPnAlpfQ2cjxSQoPVMUdD6B16lH89vDDyO2McRIqV4wtKtLUGD/Jgd2lLKAKeSb4NumbeaWg3
KmqfPUx+AFSFIDPFdXaaDc6z6PLzGj1b5xZiW6LbKp5PHFkvLcBYPBQ7ZzoU0JdAImsF9l5TDRUG
UMtOIsRX5XVk41cFDexRBoB9mgU0xz1nTOGtQHINl1qc29KG5AVn8fvvbvyhbZkqg4bu7d/26sMN
LZf86+uPyiUjE0Tb4hsCf2gNVQr8XfWbxza+vmjoMm+HiWW4sxCBKrXDT0AltY48JMwBtBSPgQSr
v2FuC6lg7UknBWG+0rqeqpZXO8D8n/re37MrE4zy3Hhu91AOBODiI3oqHRzEAucRyXvmajaGtEXt
haGS+ptlM1wZ9g/1Z1DzgLOekwEeLqK5uzXY4hDpBdkM3Se2Qi7F2HxXXkX/V8PtcgKmJ1Kl7Qkm
Jpxjx0j/n/9QuQ6jULeXFy4KCynkdOOhBLuQ05RClsJ4cGFZn5F2znkOz8IRa2PJuthmoV947j/J
5+O2XaKmBJkAAfmOM2upH4nj5B/+iVELAM7mr1t9wP5ofRMsKZksoCjweRSRXq6JX5drixBDLvqX
w6nFbOJMlbeQ1vc6pNI4ge8vu+KyBS2P2i5AoldFZg19FnbJiT1KzuzGYBH3qVtFmygHLH80iD/2
Deph6SXzwWpn0Y5CEXZxVXkbQX1lNygvr9u59ot/wthMsBtRk+CxQFnM8dZX/EqdofbU6b8LU3pU
2L6PiFRhn6AGWlJcSIQItlO/nU/XfUr4mca9hIZcK2NuZn9yVqG5XDKWxe6WVXzGHhAVhz+/5ZnR
XIlg9NftKuof47BVGHE5TuSQNTg/cSE90EveCZlkYMV6PoT7Sub8Fw4dlT7jkVvOqd024sEYTY1B
bzK8h8/DG0g1IAvsGf1mMiwrK3iFmITg2ggUHLhVtVjkRdTWw6lVi78zkkH/RtLzzAlpXZJy4zZd
FfLWTAD06muLiLO5mYyU7QCJVaY8RO4Pv77nqlfrOZWjWzIhQ87NDo57XEQ90fDhyG4Tsu/xHIrT
K2kkZzGywIJEs884x26aPg479XvTv/PnueAJbfoxGX251POYyuBHPMpT5kObeRLAS596q9jUjXb7
ax5kY4gSH9M3QuGN1874vJJN52tig0HD/fYaejeWJG6w8itU9x1qXlviS9SVNQKeFuJdyICpHoJq
dVX0N69ohO4b0lbVbsGCEt6R1PPxeGNX8PLlPo5mYIvbDgLAfvnXxvjmbLOTMruJqhG+78rOFHBI
jwpNyBwf1Kw0Rby73wgDbHicNDslfAWU4wCLrlfCPxVidV1ErXNuURTjChxez/ILlIwjqUVcVtWH
+8377Swcv9qXCXYe4qpB1b+l4zQZe3hkFwwOMu7oEfvm6Ag/f5horWkGLtFgVVcelB5Qm1zVoQAE
vLZTUWvNPhW+d0ucWNCjKslRwyLS3Y/LoI/FfFRdjHXgwLYHSLd5gTllNIJnS5ukYXj4ugeQ/s7K
qZ27sAF9ErNmsePq4qYoIduV/qF90cxAVo8/EITtNT56s3F7l+Eb2+WBuu/kfuv4T22P0i8XxLhN
8YhgsEpqmj6Wiwgv04RK1hcuMNVaXawgEcvY5boCzYRTGapUb6YqV0PG5EvH6WulRX26FINeEpgS
saFGW5pBeEsFHWsutlPd3RRtOz7prohoOKlSDEQ6NmxTLwNhL7qP0Z2R1sSwf+phPfgJTvmXEHor
oz0qE0S8VVQpsQ+9XvzAlq6A8sTU29dq/p5OoxPQnX90HHKA7XXrV0gB9V+OTrvt+Ak+oUH/KOAf
uQO20tD5seeJj4aKyCzCJJidGf0PUXXl/w5w+/vQ+bz5n6ki5ACbzlGw0GQVLMhIIVj5RMx5NL7b
4qzsfCi5eCZ4snXHRJRqQ+AAIceOZVERAukR5c4EYaXC1ZyKJhATlqQrJw6tQLX7yZmNEx66tI/p
+1KprLXg7WvI9CN5Np2it56XWEIUAH5rdXFhhQd33gIGHa9Dh4plCbP5YQFMSG4vatoXo9V/AHb4
0iJ11c1p8XUDGtZOmxU4A5ma6CG0/63g7VEvG+4CL+V2/nLon/ETZLyNaaRmv3C+iUOtAuphv25K
vDtaSJ2OLonqftBEvjwTWyCLkRm2vsQRSM/OmmzupPyyPTC+k1y0ZdsG7MIEc4fN0a+beu2TXRfe
eLLhhoT0pil93pBRlcPHNI/m1s71BT3X0CwCZBEMC1ZclRI1fOeejMLezFyN64LXD/ZXaVU5l9Wh
62AUsZmqpmspNKFmhPvo/2SOSzwCOKn4+/kBQDotM/ga7zfFGXxWQKYCdlbdzDKEkO1WMpDDZ0ag
H5k8TAsI/+Vtf9HdRj4Zv9DYFjR+jy2TwiQ1xOy5ZV0qVTHqe8zNPYODXhF5lqaM0iGLpJyAPM55
GWXyyLDe/l9CCQQ3BZjoEtxS9gsLmUV3/qFdI8KRfQsPU6uknQD+NZZs3QMYFfFXyah2gb84SllS
88sLfMJGyn1SU0zxFmw2AK1TXHizNIglgLjsWz+k7ZrUdPcAUYNbbsgTiI+qeSvN7Cp8PmPqqtcF
uGI+BYDB0YQ05H5j/YomEB3uQ4WLW5QlKHns8yykSxOY5eM2notRdmynRXfJTUs/HlxrFPtjdLuU
8u5en0sDUlVcRc3F29U2EURcbCIdJHEMA4f5psXrHi4sCQ+6ATiTv/hsuOfa3Gt/R+HVhOPYLZbF
VKrOc7PZIvbhGEykTAogplRFUQ7R7tUZjL2U7Z3OA6tPnlb8IbQtyhMSgzAZEiVfZDeTCvmofBsx
D5TrbkF0LnnCzKHvK/qMC6vK8chL/u90CCuelRQ+EsE//9PxX7gWKURKaaot0b1VeI1gGVUBRlux
d2UdMbKRb8CqhugMPvXvjbgixU2qEqjIwsWBO9kcgDgX4YpwH+flBNxpXMBRnRgEulLUOZ0XJdX4
qoA0deYSdX+Bk/oN9eM3/6OTrkCyOQkdj7s4y3OaPyB+UBje1yyzci4Kw6PrZCZpYyoHHUrdCxNk
o5ZRKtE2OmVw/bCbqhre+cPwI6PjZq54dRyhUK71ipERV5nfk2W/EgObxcFf5pYHgmvEZfkU3cvw
RNrh4sctOMHCh9eLpwyQx9N5aP1nufaJGfXq3dT6ngOtjqiL0yxUvuJWIX64nqb2DdX3FsCN7Tuz
mdvVInzvygSNChIsR4fFzSVgR3bEWGhNDwetpgwnbWASpWw/WYntr8ejvN8Ssi6JxfNQVmOXEXM1
+Tx4P/HCcffoFoaNxKk3iCvKh7kyaAGE8v/80jrsEBPSxiBK4vuETibLFFb3QyW/X4VzzNtvIkPy
fO0AXrj7Pm2EMSwKRZbq05PutzOG8yuVuI6d8pU3KNBojRQKDsx/xIQu5NEjxxRd6/89gURDxoiN
2eVNOdFGhlWYzESP9/+Cv52p4URw+M+RHH8Yl7d7Y519C2eL1OXLsvmrangAGHO6SY4bGdWdaCnM
jEkKvFDhkOY1eTh9l/lYfkLwejxPRK+XHrlWdDdL1RCN3MNZ/kAyv8UzqM82sW+3Sowm/VD3MBKK
gCQ0JWdv9PAaiWr7FyjQJqDmNR2Uu6x0lfe6sCNvK5e0/g02FOFvU8oIlQqYEzcPByCLeXz5dMnN
nyeVB0mGEERTDg8G6A6KlrsM6lvEKtdlyW3p20Oigig68fFHW61AVZtQ/B1pPecRzDhSNlVDViL/
E+X8tZFRqcpjUI8CqnG+QVU/+0wdXDNf/Xn2DFlfsoFhJIdc/MZsuzdIaA31/EkqLqVB0Dgfl1Dj
cfstM4iyCv97I30IeqAMDRjiuIStqp6nFPp/fM5aa6eXtEXRbNrCxMFfSAU9Ib29S8DzjUP1h1U0
pUvT/RoM0mCRQG+w19BPI4+MDTpOf+iz+q30/EpV2nGZyI2bPbsRhSwINDtkSS3CmIuVeOPF3I88
DlLRqr9gT03OC+sYRRKVpdEc1oHCds0UCJehyk5F6vkVOcnvvSUGKkDW+K9haNKlE6R0eW16zb8b
aTEku65sF9/2R9Qx+in+18FGvij1VBkGukguJSn6xodavCwDk5KMaiA4JqRbkcF045r5qBkIbWZv
lbf/uJHE8oxxw/qP5HXBBqiYOcGArZoYf9CDmP+96JlOqo/EPqdNELgTXL/3QPU0lfrdbT+gl4af
ihiwQ+uvLlThE1w2YHPAu4PcaV/VghkTlINdJ2wHXINQaw9/rIi+Fm03eUDp5GBQMbaXb+5BhzQg
7jU/P3IRcRDGKSpJtqdUM3udwtKqyT8F7W+MrC8X647TO45US4FA1waTCLJOouZL1GC2CDnk0kQ+
4H7WKdWeZGCgjAGIQd9K+CwzaQZj1e5uNKYd9drQ+hVi0Jm1sZ0MnUr6DifvOC2NjxfgXa2Xnysj
C2mnOIQNojeXuVzSVudro/hfBV3J3NzuZkSotSmm6yXOBimFVBwnS0XHzKx41AnAeWQRP6u21Iw0
2RgVwAYNCmBo8cv7K017KFH18A+rLljcXz9czgkVPNwDfzYdwjNN4nuG9bgCI6koNjB9V+jG5ioD
bsmK2//2WUHX0EcLG7/Gzb+drLQlNvtmW4Le1LEehHKwh0mWP2tljlaZuyi0otYABkR8oZLXq9PS
/kCdUxKPp1+pQAFhqt9DVnTHoWkK7PPGttDrNXW1s1kW4odqLNg2MKDdGxTb3/5CYoJlppNxwYGL
jGRSn3MzZJdOn+D3Fu3rl6sUlbGW1RyxOsokJpfWZTunGOgmkCo30NtZStVe0YvvTxqdMUUQCdkU
iNkgBsFFaVFcrYNidp4cAsdrtAE/+KSOsP46XA0ZSM51HnuJ2Osox1gJvtIpH3GR2iRLqq65azW3
YsKJOJlNru+Q9j6XbAkJPs+wxwa79H7vpkYmjZRGVwmSXdAp/8N6SqPghH+rpLnqd6FB/eobo1nX
vDOYOVF2pK7MBq+lVO2zy6aaOf0McbLGGByLTyhDJx0urhf2cLl3/XeefeR+xSIMwO8p/AlpaZ6S
AYbjHGtdr6qu2B2uT3VkCz7witlGd1LPmBmd3dzMkltlxmiy2LZz+FUc1FQUHL+fqmgu8vIacz97
81ZbR7fpDxD/mCBRrn7j9bvWuyZloJ3nnXki2agmCdmkBgB6PXw6U8B+nh+k8lDlh3MFmts7tyDk
iHCpx/H22PddCUvmY2aQjk1BSBPAAMVku/72iOcur2nNNjtCGO7ZILV0lkL7HoQ5RdOneRdu613W
STpOoG0ll3bAsLzBKvDnHf5yyuJNVXqYSKvDUbcuRZja8+BYzZh5tfP62Wd/juziTJ3JfLk7eco1
uG8ppgerWwq7PcqCqtHnbu3LLDN83cN3hcfoowZpXReaqBP6K5nf+5Z3su7m/wuxwLgUR6vUE23u
X5h/iUJ/PRTrHRPWAo0snydzg1Lc4P3QoZBBEFAC0P1VAubr2FEsFhMq5fjaXHS8K2c+DFHplFMl
kUdqNlxu20Q1jY3dTw5ViGzN89WKwGiq2YbrSX59zaYMn2tNDWlPeAj3BZUAQEypqhbKL6BoKia9
IGlcc61ecY0fhRFzt5taF1uuqoXOS40wCIaLN/DPHwGPxTDWIU8wBcYrvUQCSy8x3RB0Ox0hVkE9
AAWf7IBENdaKpreh3iSX/WD2n/djYFnkYl+mJS9mETEJQQ9cktXN9h/c66JPRMjBe6A9J67PnMpe
JLz0ifcFGEmrvwM9bxcuhfoSxubo2l5bOzrDZtX4WZ2SsQ81YdOAoiIiUG9Uge14fhsVVdQQIPSL
3/52axpKbpGGz/O2fYhyTyZJzvw1ZDkOiK5b4kciKNVHLdvYu9xhRwduLfHT2GkAa1FTtGte7cNy
UqartF6SFCjac7/UnPm1h9Yv1KaUdD84r87YvhSrXK2aPWxjAkthjN7VtmLpDOYEyJeMGaEQ5f4A
ZOmBpFDMdB1HD7n0InLvzv2ruHkw2b1Q6I7c5LmY0TKu5A7cGl/Y5y59JBrDMuuUnvGyp7qXU9St
sIxp9/NmDsZiclDHQJKPgiSKkAWbrQ4X50GtZX++IvizM9i+mxsxhUmNTQmZ+n/O+GJ046x5ESpW
UbDIHuJDIw3k6vhZ78JAvHlc5Dq+W/2sX4MeidsNg6GDP0805n9yplF6tck2K+wc+ZvGlclI7+/F
UylLT1MhJFZ5f1JwIFAj1R0VgmvV5Pv0bO0l/ELO62Il/fZ+Mb06Q5yTgiCPxA0n8g+7aFlyq8jx
3wHH5J1lpKLSvohcmloe8aIYm0UQazwiA471adzmZvLnpqN0Bj60j5HZm81DlbiTHnbu2rFQextn
Kb6af6kHiuf7V1HsxUWsqOiarz57foSXotZiYZEiZxKz/gk0IjtWahdWjYe9ctdFVibj3RgxRCoD
SVlTg7uoFrU4yjTjZSlqI48rQlH7XtHhoRyIFpZRBf+ReolKd8yNfRvHf7AkbX3tiqBYV9+WtnHx
mLVOuYj3xYKoVNOihzEZ6bMMAwOHEx+RJ6ESpveyg7QpPwuOkxOHqX68B5LeTB7FX7OIvxJ1rhE9
0mMWxHZYCM2h4JK3wewWlc4n+sKPnGKmEJuNGsMX6z5uCJuolzCE2WbgZU4+YyVEuH1PTKeLRkaV
5TxUtGXsmK/iwypF+yhPHNf8NVqy5e1DQ72Imf+K11qwzBbFpTVfUbLDN56A5OyrEZrqgICl9Z5J
fOYLcvVSkY1SkSllPceXYIbfdZi7VpOPIdSf+AROPL6qJwrQqnFSwWsedvxshREODIxvfjkR67/R
dWWgrl7xu6x4qkZPAyMsJ2sv+/uHiUagB03NPvb4GoKajqe9y33b/1zz5pyvChw+SsGHjvVH4OSt
AGt7S0aF8UaYeZOcL8dZ4PncJDuITgcP1l9g0IgfBUwGoke1Yt79bKspVpuV+eXgMicG9yCmdMPM
2zjMONiYjVxAvQIKeCg1IzaqYEXAdSKIwLeT+LcxUMOVeOntMHQVGuAoCng/Wa7cLuJO/QNAH451
l86BZt4J2WDJHd4eLsJD9XDI8Xzetp+tIPhUY6ygJjaOxMYPMW3jQ2m6A4YSqONn1PhYLXtIwBym
M8rjv1xKUhqrPQm0ACSugSbtbvYvMpcI7Qm7Xde22VVFm83ArlqudnjOoWkcMUnZGBEIDdd+dLGR
04SDeftAEyzXtHfmMFmqaK1GIqHTX7KDEe9yDxz5vgNHDj/rXYm57inwcUJ4B9HvRVVh1CAOz1gd
KCG3eroI1lFSH3YFT3ccqeFGqeCs8AxBX0YOHxHn6GuCthYboRTqLtlb4l/XWbAX1LhT/PWe9s4i
Qk/L7St8Se9usOStOhdO/yj5Onxud2OMcxHWb99BVIttKWUbCTq1Jd3LvvKbRj/KOO+uDdqUrWhw
VOKGG/RUHp8jyB+/1SA840s6BW8LFVlGlFLIhS9dTEEXgvQwShO0M4BriUzJ1s4CkeZBMfxyGYgZ
ZwrdFabidhVVkudDDz7a/FmjRdGbdbf68RNp3t+qKhixNbINvleoJxw52wip7IjHc+ttaflVsybW
PSIZSIlIBge4HBzlAh1LDe8E+QuZTblwUH8yWR//K/mePAQRstvLc1P34T0KKD7ySZhmo+gnIbso
fb1nzwZFTylYazpACiwpEJ/8fMj6nco5TrUaUWGuwQJAMD7+Py9jKlzfvWiEWYxQ77HBNz5Qj+sW
gxqodAOehPqski/6T7PF394+MKPzMFYppDyCtnht7y97/POIkzP/ABefBzzqzm6AyZ1grJ59qPfw
auQE/3+saFdnqXV5NkhbEAjLZN47f9sOKWbgLxdBE3iCdNVXOYDSZWRr/z2l18CpjjCCEq/iuGTl
C8SgF2kmqXIBzOP6ekpTqORGo1UsvQiB52aK81hGusCrwexI2zQeO1RasO9kGdHrJTd0+uULZnT5
yu/+1J7/0ChHjZitZ4KBK2PeHE4YsBBbKWUiU9jaCsRq16PJTFUgBoA4i0fTEiXYocDywuUVD5St
1KfAMXJnAAVl62rFx+O0laPISq3Ozm5Sezl/JYxwtqxDRM6/lCCpZY+1FqOe604yEcGJtn3cW6Rd
6tvV0RMVcM0sJeGZz3mk8vMLBaLMM11BtXmbvxD85U9crvs2dAgZeY5M0yRzWwxZ+TrZQGsr+1SI
yoSDtfqU3auiGHtV20OszswAWSE47gY6o49UzMJSvsG/Ygi6z+QM4XacqPzIeTkzm75wQMnIkOmi
sVEubUwMCfz/m/XAlAP0yoLNhxaCD6/ObxYOaC8ny43K+sqGp7w4w14AGaBcIgmv0G9Q22XUCEwv
SiQf4kR/sTaBS85r16mphZV5OWAOzaUUlp63dvzaltk2JIBJB0n/QuE9DtQjxdD2oMU6Rqk6A7Hd
sPjY+Q+XIxvqXE+16hAfBOha6H3fS9p1Ir6SQgWqpsMOXKTYRZL0tjkUSBzKhZUanWrYZZIPwhbN
0xB7W2KgIbpBkGFCqIXahy+3Xk2Z+rh3zU1y9dtVZEOS79kzRZi4y6SgSU5D012bteiMZGztR9sr
ipDqzndYfxGmUCuAIPcaEZEp7j6df9c6+BTTCia9rdrgFk1ctDEyrWuUZXWYN+wI7qsWgensULB1
fG82FYva4Nq0Us7AJtGxDjMV7bdKFCTbj4sycqv15X+0VPX/l4Lzpav3ZiWDR9m5cIkJ//q8zV8x
iJWiKUQ2uyy7Re5wrB74x7tJHai9YCdMTYehhOCHXwaqkWykzRILvmByEiE+G5q2ADUmpdpWRBCk
vrU1IWG7KOxLZbTIkmCTDl7SZLAfcnacDGSKCsuQIoN1JZh/hfx+iC0AyzZEYkoWcdI/QgdPudbA
xOAHZjH+wdsrNKl5ZtPMmnpj94/VlZts8D/8uEnVFQbBQtiau2do8HdXK36z3wCwuvrCWY+V6PoO
2SWEA/yoNBUr3ExqAOG5Xosb14aU+Q1MXITp1HGJOsjAMqoMxXas73UWKw863eiUwywpW4cyQMJ+
ywBvdhtwivv97x5g4nJKpUryd2oQRcFljkAhXdp3hgEe2W7LOmHucs3oOpC+5cKGgXYAsQnrP80C
/dya6wzM3YInA+aUgDASDKusV0i5eWHrp7WXHbaGY6gMKkOEqRHqTRQiCi+DlyUoosnHU94o+p3s
5bb5w6S4GHezgq1YSpinf14z1E5hQgF4wqHqN1P12okLK+Pu5Uvv8WM82t2G2EYE7EZ6+BqBoZ/Z
ji/P0etPa0nUyYKp24wX2/ihPQME3Br0pp8HI/sTdoOEQAUNFdGf7CT7SIAUVeHqjz0hmxfpIPmG
3rsmIJPWNkO3NLmziO2hY3Ecvi7SKo6n2PzDJHKKB7MmMkDg+tBesD4xlI4sTk+j1q/CHt2yNfUq
oghlr9xP6IS37lrGcfY550BRBmkQ1OPchZdPJK/QcsUu+xkorbiXA81IWRj9Aog8EyzVcgPMPa25
r0p27sSIptf5VxBvasLuLAGeIOXxb4XLPGrN0UirKzbvUDslkLb4qh648NY9UgZzyC0yH7se93Zj
ZG0nccwU7BruL6ciLrx8L2PRXwoVcs5Z4IxDVjNQ1FNpenAEP1t6NyFjctPkv5tMsAS2bakOWW50
hzcTEmUGNjpZ2id30pdSTd68Qr9Q7qf1zhZyT5jpJ1P69DdyOEh2jhuL1YKBH1rD4i8kPjxiADgu
9Vjb3mELlnnARXjdrXejandXPYW41TYa6ps7fRHM68f6xV7sQSgl3wZeJqtfC+B3pcAWfuvZzDTC
xRrW/QPeZVgVHh1lzdfI9ubCtOLfeA572MpH5i6gjmXVS2uXOuT8Qq2tx2u3yRJPFhJzWoKbp7eD
4K0E3ibI+wZMuLlrPjlI2qa/UWkiu3Twe+UdxsyIPz5yGtDM9QqBMuq6j6F84d8u2vcFxu86o90M
ayzfCcaQQanxuveaKbdDsqu248Sg++XqohL4UKJ+uY77aq0/9iYC1+YHaLB/lxuBrASK+nSjjdsR
K04iwfcGM7WjNYeUFbCdoOgQ391793K0dsWF++jjoOZOgtvOoJM25r4jPQXJiRVLHtpuzK1M+e6V
6n7Drqaf4mwEeJ66qdK51gkAi6SMDMJ+Q01rljhgdOH0CRd40zPRzPuuVCwsH8dNeblrzZh6UCrw
EFXBp0j1GIp1fH6jT5h0NdK5sNZjBnXPxDnLB1pLFu4zECM8/5a0pRSOJ4pjgC4oUtzfrhcxcozl
KKcWq3+FO4PCBFgq71b89L/Dm8diMkFxo2A80OXe4/JN5zDfG2mdnHkFx5eSerWVNKLOtJGEHDzH
21mu/pDERR6TJ23zjVgtfPswxfswprWECmC87nJdytEi2wF/DEIndmYcgSrE5uEeiAyq93HuZGJo
DPYLkco5oLtVnaZC0x46PRD94IuDmYflNYtgacI2EwFUqF+19Hzbu3PTvjlMdZg8/AlDShuz7Vi2
SfP9/z5rsL+fhFM+CI0TofRR4bYfjz/0xz+2KOknDav969myPXGjfymFZ+KnpqbhAQmC8wQRYF9r
zd4GNCGR3jpuBcjQwq2Ui6CnKF5MK/Ru6SvsiTwoafdAu1y9tAehQQ8pjdbMKaKmur/9zq1mQ+gn
w66xP/J/1Y5LgJoL1ty1HVqBY0uoCdoUo0PSRKa0vmWqEAjraMlZx7uSnCLtoUlx5ugCPdXh57fX
FD40QlxR60ASW0kw/u6cvEMOMUc5Bq2afMIgXXNxWcfY9352ka2v+UocFrlc54dMNiOF3lSrtkxA
ZOnvnGRwrhGbG8y1ERT8sdT1UNPBpbQH0UQVDFQWWDo7usIvFL7ZEGnJzLs3EEFlgTZfJov9fJPD
deFNpX04Aq35+Md1Iu0SKRtDfd8rHQgFvnD9QXSNyGGJ7yf7sLRy2Js2zn0iWNgNlpPnDhCFJOKh
0N0pKTMMVEJoOaQLRe8H8WsoJi8DEjfr5vHhcO+GxlvGX7gGkbHWgPUKs8jJUM0HmHp8sNWs1KLj
mGsbhUCy+7K2hmIDejXkWgKa8BUFZnOGlbxNXM3jIErMBrGrkZFSupMC/+9GDJQVk9fsEzz9EBG6
gwjME2OFhSRHfhGIfD4xDSCu2SlZ7F5GYYQhrWmlfIKOZAyVX3Mx8cJoZwT1cvCXEW3Z9ZPU0VY0
L2hUTmHNFu+Wia7Mj6oFLK5qzYPmZGafqkkQ5t86y7eVifMRwetOHn90HH0UQ+ohR32Ug+VJijln
jDt31Ik+c3Dz1R7gvpA9hTq8cvuxQXspUnuhFB4Rm11AVntaS09Cibxn56mCxW936G9U/+Htxn5c
Rfia0ah6bMrYfJMRJ8mvc+dpwIfpx90fiZxfoUNDIks00zQeh1V4SwBEPOAc2hFLW2i/QiCPQcbV
k4gk25RMzmvpORT3MT4ELg0jyJLHJNNQlr9ufecylMvxOXhcPW7vglMxIdnz3FLJ9eVGwBhWOPDo
UtOH2aQNcbtHC+qAoL9bLd3audTDwGN18a8C3Pn0JOYwCAQiifzOugcjfdOIHSp2m6/vRREmHLXG
WLYgMyMOEGdRqqTcV4LfMcukD2KI2IzaFsyFHmUacXE7qUYQHB1Uo0qNcm9UT2h+dcSQlAOif/VF
mAOtR5MyajjwxIDdHqwhnAly8+EnqkI4zRgFrlWrleHtMpKTsy+Q8c294GPTztOt1jg9xOIvSp0a
fcSnzV38sMPT8lstLt42em/o+hYucidaKcpN1otlG6aLD6I2aJt0Fz5YrKwSEf9zfcXg1fql79T+
JQxgAdo3DKuqC+4jbo7WiOCYPirs1iQ0riyXlG2DHFDk/nj3QjK9oQnqbAjKD39eMOmSf9f8epRI
YYMsQLJIzv+MZdEZFonanbVXgN8V8rIEUE6gfVOP8fcT5foVTWjCEjQmfh1/F40L61/lzS8pk85a
BeYtDR5wNc3/M3lyeaa9JUc+l+sqaxQkss3aY+KAN2+yJ2apiDGSmGzC6I3NXzJtZZRKsnxYFNUG
lnv31GUMLKC6IBslN+0oVo0M+CeZ2+I4gBEnsHMHIvrTQ7qP0jET5FJ8zZTZVmYsH6bakCfdwRT0
pmDnycPRcA4EkgOkeW9zs0IbLqPTtF0r4kavTKaIKv1axIjHVVLrVu/o+FXNLUwJEpGDa/zWaSKg
xWW/eHNrl3CmSabsUc1zD2jUJd0fPEJhLRZ7lI4/tBd8i8AseIjtyGYj6pYb+ivc7y63UppCn6rh
GcFhwK6Xf9HZh5Oq1C8QKy+3PpfY+Er2AHhhiTuRSJPMRd6qs92+S0auVvODvVL3TUa1e3T4P6LL
0HOYc7/WsxWDBIwsIoxIu2tW7vCkDxQ8bI8IXMyp0hr5uYETHBo4AoPh7ybrqNnPKVcgmANTrNXc
qizg5/lIp5C91SoeoxR0adQLLCm1iawIx2NU+NTTVErKwjKMpTFAOCPpAtMOUbZSvHi/K1C1/T55
m9UwpfEq6PxbwusarPk7wptbdB8WUJKGeg3dnQqVshpwmiT9fOzJogBY+i/HmOQniwca2nxvLefx
cD6R8B/+mC/xvkCjp9lMllP2bds/r8EbDY81wqVIlefpcUznY3Hhuw97zYK+q5IRAuV7WQ0C06KH
eOPQ5HvgIw+6ioKk4qZUdQthmUg6KCLFtwknC310uctw7vL2TKV+0wLXam8hGCqenb4LkmDxIipJ
GkkO7oDpDrv1rzBzQpPly2mP4hg+gaGG+LBxbZm7L/xlzM09FkkxxmlSizCtZxWtY788HUyeBsKR
QHl8qCIl2SJ0+O1ucM+/7R13NfaKf3hDv1H3BAyYFa0ERIF+z6vrAp80au5jf064cJxz3p4sBELS
qGehuSTpVhfsWZR4fFDEuEe/1QL1bIG6lauz2hjEBj+gDPn7HwOdamf6PgaV0vKVJGxdLNOpPKUE
ij+xpeNTIJC/xJyBNiSN3kxng7ZWCRpNlIRZUsun6yJkecDg9jEJGPdh38AgBi1YMiHOBFFimcP9
FR8b+S4cFwITc4bKnKzKf9FYDcR4GLfGK4ZBjc9sBeX/5tk2gd4F4SUNtTPX1vQmnoa6WkkdqMj0
YJQtg1K2nQK3j2qVfzO5w95PcDPXjaFKhVXJSmYz+TgTmGwWXbtEbC8XQZriEg4aO7lOz4yboIzs
1IUwXPrQRx4yvtbRwIKXcSvx57r4r+YcSc/jnLT/AZUVl7jMz1CeEYOI89552Kdlxy/RLzSvMD/P
ZJjxHW5538Bv7tfCjHJxbvd4Ln8TZLaDy2tIteVWWccv5VKM38loNhxZB7VGYhnv+GgBfwkLXy/g
cFRo0BksVs6KP2ziMWdKqtSeTU8rpeOeDaU7VWCrlMUAk7XheevQxJk06Zojkt57Otrr6mBWFdSi
an2sAFFNDtpowxATxWjq9/S/1LaqduO7n3VKw/KainmGkhtuHRMKLiAWy2VYhVPj9okK7Hcl297X
3Um+tqUGanMVW3HooExyXb+0gXCIb7ZkLAGt2+q1nGoInLrTZknRII2AI2OzlaIASmnJed3CqnQ+
fVAg8nQsbMwkaTqSgIJHWRx/1zkyt30xXEsIJKoXllSyl+jK1wzWSSVs1B+u9JJccQ5MJ7Q+ZxCa
+T3LlDtEKoA/zSADkigF/zKmJ7+k6LwLQnIJuXKae/IHxaZdGlJr426IMnPOJrt1YL3r6eZomaD2
z/PMUHZuSEXt7nYjQS/LpbGXjD3AleKI9+Ct4pgRB+m27+yw1tJb5RNrI2imrqG3v/LBcHQOKgvZ
K/lWO6ZuQjaWeJo4zjYEczoiIZ3bhsTPN1dhrY13639XPFfvPV3Y6TA7JIWkFMzZuehgRguYo4ZA
mI4XgUp7vmjFn0lSGFlJLfwNTKgEa9kVpSiifFYrfojGPko9xKxR0FXHLbJCbucC/2ZbMBCtlUwe
vIUtNTf4Nf5b3o7dXOXTETl74CzHTFO3xhYE6L9CxQ96upyt3fy+QfF8YSp46OZoeE3NKin7EVUH
asL5lGhxgTPvXFyfMc/N/S2sd9F/XLNisBUp1ZzKIXBDql2fBYpVNr/YsVEldV+M4ROR+mpzxypU
d11d8AKHM1tRkazZPe8YfDH8KIb5LXtysAAZ+b/YYFEk7Mxt9eh+ibv3iSRksG64MNTr9r6i2Qsc
9p1OfbwEo08vvIO+VgWv3nQsVE3ogdLn3EukAa9tspjyb8FqxtSvxeKMU5hDeuVmO/N6Wc6DayrY
rywaqUAc5g+osF/O+Wc38Q4ohKmwousEVjAXt6CRxOhxRUbQvObBLLaoX4G4EbG42oWEVQ9wwAz2
UoSa1G4EOzR34JO9Ct1TxSFVSnB6B8bj4UJdHIG4tSIDgF7mPwzM9iYohtfz7tpJUdZBG5Ii3ijf
kAmaypAQ6/5qzpD4nt4kHXm5hY/yA4x38Kn083PRmoCdtdQY6uIuz4/9N/++bir3zXN3gEteBTxt
mCL4CH/4Lpm7BI1CAVB7n4+9jz/ZyLHyyon9CKPmLdh3/Wn3Omlwlw4Mo1yqq6fXJNmvBZ1zTpHR
8ywn2ZPF2QHzU545P1SSKz4rAjLsm2S7jAh56sYfG3jkc9ZwxOkyhGOcRfv2csJA3haagMFc52HG
SpKmAw0v8cLR/Y5uyGSvFJqo5YyIWnRbLCIZS1q/mXrcD797XAdquUyDvqmonYoRvGsA949ij2hw
4J+nfS33n8aFkS4BimXd/cEAhC4Nj3tjKpsG/kG7Z/JOGOW50h0iHHcWleWe+WXTUxnGY9fbHcMT
i1FRldqpX/nW77ohLAge5oi5wOVQ5Q9CFjWm9SWst1qfU0+4F15gu3E4BWENfaqm+DwXAxiMWLEW
wq7k8sc83HDBXLrZFbgRRhFO/pnE6TcbZkQlkGgRsyPoqnvtrJV023ZL/ujDrNaidF8wN/hNNqQn
kjWVVnTz0W/8aubxkx51eU9/GlxI59i+eahk9RsJOFuAEnz57k22+ouAVY5tiNHHK/voLkopGHbw
ZQqqlBYXYc3rLszIlURqVJEeAKCIhS2XZxH2F6XOL1NqYijg/D67UM7f2p6dInXoNZ1QE7qCitl5
KiOMz7Sb02F1rIj5f+FGLXjL4Z/uGGEevbDFBnXmGHvJa56XZ6JdCoa3XZJ4P1e/BsK5AV8ALTF9
VSbeCr0N9YFgwI3Zakw74XOMQpIh6KUcKCiJfojJBBCyMe30/3pYq58ROhex8qPNqH1u1/2qqghi
gTZ0F81i4tx7x/9XVUQNhvNwsbxRvlTSwNQ1hdGzVcrMHAvBt4IIW4OAwL1eEE9Yr4vMtG0DZ6tJ
wZ7FtSv0ozBwTqYbiYCutHG5prihcvukdQfTKJjdftFMk0hQEa+rQfHWwicZfQ7YaqNtuXqnlROp
KFzIXeJFTxWWUxvFeHW2tH+Fvecn1OrFa751VO8XCAAogAIo0QcxQjww07KOEUa04WZKX5YdfALf
llF+E9YD0lF/d0F4+d26yrUeC8KfHR+xv8KtciZbNHnm1L3UCPdRfkYztc/gwu+XNRaPxlWAlMjo
0b3XYQoFzi3LNdPTL001JoiGTvKIq1JWdTdpbdYVAIxuoeUi4T/AKIp1T4/JPznuSn680eG3WfS4
ig1uVxY40MDKUG7Qc/6P8a5MYZmFmqDWCcgigQOGd6e1pQnmQtUVLdTvwthMIGVmbytvqcKsWX4v
IeLsssQHZBZfHyQTF57EO/edqagIVyMrVOWkxesr4G5QINaERRVr+ZlHFpHWRLS+i4Wabet8h5Pw
++aof0fbaR1cuh7MWqqtrZZeF3F/fUMyyFYNqxJx1aWC2Pah92Cq8TvTNPXEsDUUeQpP4xjCbIPJ
/Ooic96u8h6O/y9cDT1CAhW1/y1HfwctefroLkA1ntJArjNoBvxVkVOjtxaqGCySR26YETSMxXH1
BYTzO4QZq/wppEd0TbvJk6kXRyuc8qIZfJUcd2GmydmMWYOcEu4nfk7l/ITAevn+Yq3MWMFpQSEX
koORw2vPRuACAmdZSOLX8IX441DCpxVqGSaFFjX9y7QEDElcmB7zJSUnq2V4SgjuUAU04RuqafzG
KJTDtVr4y/TfFfZUsudjXmVGpKll+n/77AeA0plKC2ErfcuJtHKgIVU1Ol/iGsUg5E538ifsSKNl
FrpIoH4gsDOKDtnNoPmm1zx4jRRS+UQv9pPxqLWoM23GQiu9H9KXu/a0xdmZpy2nOqyuXLg9RnoV
O+qDB7PLAANx741E5cVzCQsBh/BZ0KOXTVkhOkxaNZ9Q/6FWVxcMJTgb9GMNIUOFt9xOvq5Q7F/9
hD/R5+X1mixP3qLriwyeMoDn14p+rJH1u2WmKa7kZE8gFhhe5hj37af821XKfurRwjFSwCLYmBKE
wqZDethhnb+3L0kZhhs9/1zDqXlIoWdwOHUK5FllUG0VSRvHZSEccOhS6dFrj4u5o8ZLN/2C9Z3X
vl883rl5L9i7NiOE6XhsKXyMhUDD4m/ml9Oh3V+fv+qIOdVMVca3/fKlPOXoTI9Y8HQlGc0MKbYj
NpnRBC1E8IStu7SEmEbq9ijzwrFaw+tcT8D1Ezs5sc46oA59ejH5Z5k1vMHyc8/dYs51YZB61Mq6
fyyiyZXX4SgsCIL8lKBUPuI6Gk8tKKQ3SkqeY5Hibwa2jL/CPkPSEMXDWV8W7FjyrjtuE22Vmlme
D8gvWSXG27SSa7uXYCFuZ/bmrms4usdGMi8J/7tIVF2OWOHgC7Eg630JLv1/vcys5dnjMP2OG7us
buIaR1ooHE9UbRYsp0o7MQwO69ZxCkjXXdtMoh5Vloz2I6ttZE9U6KQSATjZ9EGHqgocoCBtRUFi
mI82P9qBhBg1eEJFXAPRVoMENeNficlZLra50zeNecJYnv7y9Ld5Q6SbKi7lkRsJ08evOyOYbvqT
Em2dxgzXOOWBfTOUw0KORl0war9RFHkHZWyIkuO7UlDhs1Y9G0qXDuLPwcIq3UOAWkE9IWmEu5D7
oyi+8AtAKFdgTpMy4VRmhyawbuZWAwoU+/8xyfQTNCViG5mEef+TAbg3yz3wg4AuZ6eCm5fcvBeU
sOXX+xSGWA5xWFJF5tdPgz0qrlR/djBR1n4GYEoF5U/5JEmYa99bf3E6m+ZCVklzaqD1mcIwXuvH
lD6HRMsZD4LaKDLemq/64tipx73888T3+Ivq+ddc1p/SRNr8EokeAorC4fFPQ8kwmZupKmd6aHcf
9EiWipZJ/Mg2XKA7L0/OLZJ7qjg3BD+1A+c01uiu2ZIjflXQ7yjo5Ikbl0jr/GSreC6QTnkja11H
4gYSIs3Hn0GYzST+Bf4mNhV/7Tepn4WrFtAunCnWRYX4Nh8f8pPe67N2DzNJAnj5KVmaBgWUQUZh
mqsB2swhPOOf6acHjk1bUAHSAhr/9Azj63Zr92MHGPkQ+HKWjP5OsTcPUOGOBQ/uxga2xV1QKaTh
roFEo7atMerjba04VRIOU/Gx1/jI3V8hp4VdRcme3ZZ5EShtVUrTgMsrZqpUTLCrreoj25rIXoQA
uAa/iJE1xryPW0J+YoUjzgFSKNpHo5zXhQgVHfiyWYi48349BXetfrVA6hhOwGZ0v73qiH4vJr/E
W5rDyGBamT2B2/Sr9oc6+S/VfbSG2hrcsyg5KvSPzal9oYIn7EcmL0EO+nFO0MbKYeee9GHRFMBs
+5tMLp3akS85H6BMsgN6m0icB+iVnrqdyrkNmk7/bECM6+lGDbQuM4MtYvOxWd1fudjdrrIasBi+
whSHY7ykYUdb1x+aY9Lcve08Xd6qZKkh95Y8DHLmvvUiFLaohSJfBq+SWV0ACn4a1iGtREPJn+OK
a9tPq2ita6CexZ1ol8DhSNnVBFbKCyUM4d9T23xCMFTbklJ6TZ/YhprmKL47NL7bU/9e7yjQ+g5c
d33c2O7W8Aa6Gp+o9DXhkpirXG5E9dJatNVf7bokCGNM1deoYFBWhjoispllU/X+UVw7nmARgLkm
guUjM07Goq6ipBqhzYlOliB0NPgNqjkzaQGUr3qnat/yFBS7CFIxOUuUdUH2tYF7qdZI2QjIVCpW
oKrpUrVRciD31qBcO+X/nvAI49/HWqWEtBJefc3nKgZE7ltA9S0w5Rd170/VwKESdZN7AmC57wx4
tfxbAoX4utcOy17zPlnqhQosxIctSwp4e113alVeHBkNe219N6uopM5voJ6vTTm49PJtd/qxJhxi
gaJ6Nc3bohE3i3lp556DHC5Sr7Imj5/Sk9rFSYN9gLbYOeYrGlccvfUGLUOP8zyavmLCBi/Nfdsg
33cAiZhvvj47douKSL4/DAXDIu5SbBdobdQSl5zL3PC3NeuZ+0raHGy7kszV+Juzvou7720g2RTa
+IXPw/1ydjFttQgnM8Re8wk9WdVFHLYqgsRbBLJ/TQQ5mEY2Ibg7PgSVaE3XTJfygYDmP/GGJMuJ
tjkNdlFxsWQyfXWH18E3ctY9/kx3/r2dtUCe6wiAljEH4QfHjNyvFDgVS+id2IA9JJ7mgKwpS8Rp
TWJGhAVUFyQPVKIKxbN8RDS8lUZwuauNJzuicpiYzF7jsD+ojV6fRW3ZN+POuWvWCeCZR+yrdod/
P5Cij6oQSPzcvvntOtWxm8Svg4KapHT+Z5hMQpVK8A7+KN5LB4Z5SQnkXptHr4VEGTs8B+AYFUW3
CNE4JVHXOtYKh/Q+cO5phKzNSE3B8X2DCmzi+yWfLTcPFzZCEchQlDdxjk+rNfsbXMtBJiPb1PAy
QTB/7XanqTMCnnvZiRl4kcQ/ABSpch+vA2YQpBjbXqXoEYXt1iGrU58QklTT67Fe+u4/LBC5aIb2
1CjfZ+Ckh+y/UcYl/RCBlERjajkLLMkxghVZBTECh2wf+movdgqZ9JAZoPa5/MCZoCSqAya31yZv
XXz5ProhH/BDI0e1IVmcIbNDH5eQeMHu04Uld+Lso/awjmHpp43V9xk+ONCggTE1CY42mVSmqhvq
469Pz2sHZW6m1NEcsOpJkoZjGbyHKxGXWDAnDArLr7RsYwfhcB2l0ZXeXnQdWJHUKLcVflyOV5QI
Hj2tuuR6hNslCy/Lp5usLRk2sO9Rm6EFxCPzvIsyMngxSMQKtFIm4MyWJZ6A54yEPP/M5RGAFmDS
B576Mvkv8qcO6R6JkcU8THfpHomlOb32VbOoW5HO+XV2ZIHndj+FSV+MkWKMrCQ1k7PepurtNg1f
GSgp1ByStakPQjiQHSvHsLnbgbTPZe6HTGfPpUgN/sLDGEXtBaM9U3aORYwU6JXr3WQtul55McnF
lTVmk/xm4W7ozNe4Ren7rvUWGzO3/pwVQ7VKjLJEUcuQEUR5PIdGQHhaW7k5zhW+UgmMEtyeabWy
iLdbS+x/fM2A4SmSaVBRlcAf7dIwpog66b2qCkc75xHEoPk1T9xfdKhutAvQj+UJYg1PQOQsQlHy
N9DYPKCLrBRSIvoWR3h6vdnaIscOxtBlpM6Bgsvm2088d0DnLRSTvtsbyCxam92XUX8gShQeEu4Q
orGyv7BHWA5di4loNOj2djAJN0QuMtJWny2ZFT2B6krjYVF6LjcuELyx1MPiSVWzBzXmf5XbtTlw
GYtEXASYD46+oMts4Nx0Nfu5CYAGt+4dt44R6pu3OwwUILLW3rWhlYxO3sYuWgUt+saQ7C8tKs/9
3E+Cf0lVlHusSBFI1rJcFKia592ui2FFl0nbFnTxFxY0uV1zlh+UVG5xCMc6SWENpx1SXgvlajmc
J7sbs7M5Ic+h75NtfAxJCyWBJsTahtQKNiPiVXDICG+wIbPVlhfSpbROo9yS+qxvxr5rA+CvNY53
LkZatv8YBvvpkHUqxdZDC5nCYo8C7zmaytBOa6T2euSdiU4se8HVqSWFWsfOlxx4+t341Y/OP9V0
yi+0Rh5YX2/Siun0bHA0RJi1D7omOaI3Khl41skeuBBn8E8Opmn79/dc2PdgRYZ0/WYn4xFTXbGE
DO/vP6ScaGKnueH+29ytbOvF7av6uHnquVFG23t4vOMQYx4648IzHJ9mPxOrczPE4SiQHcJBp0Hl
cAC1iY+G4IMBdze+lnOU9kLYxj0OBriSwf0dU8lP0PzRr9uGVA/Oh8bIEIRy066xpR+Esw2BxFPb
CM/fUVJ0Ubm8e6tgbabuDidKo1NpeQ+peQ24AokrzHzU1p91b5QHz0+m8fs4uuJKbzt5EVJc6hyd
PJrWwx9i6dNfCreQJo08rodM1+6Y+kfX1yuPWigwI0C/e2iUujf5T+WskOm8royu2RQaAxXnoCjj
d/RF0Qs17ntWxipmajILmjsW1s4OWkXposdgZxnExDW1IqXReZ3vQ/r2CtFCZjnXkSk37XmkA19+
DviSzLOloixSWFtlyavv+/yh5Y7K9xxSJqxi7EQZb4KSdkilMnJe3NG3khFSac0ac7ETPrhWl/3C
ofHpQNKkDpPqXcXajUKPXvuj21MZLfmmpMrhwIu7/pVgGSaHPdAq5JGRFhMe5PJJCMGREnM4Kn7j
UGqCKmN7N8n3z7iHjF1nHGk/p5I+HjCqtqreB6KI56qtRNh1dIR8jEl8Rwz+UqHcZLaLfLeO7ivo
MYAQUYnWck3WpRc8aoWC4Gc41xCuOM/TRmLtqvp2hom9wfUm4I4BMsH3t16zSQhHKrdn8beVrLca
HH/wZAPE/Pu0hPdVx7Jn3StgpFqHcLevvPhs+Tb7eOKUmR8GY13Bd9oBPnJbYTdv1FyUtWWjptKe
qM5mFgosphAiRtSEjjLimTtXuRSD5DpF6h4lLThOmfS41zNI4JTue7J52/ZMsHYgw14d8I1S7ZuK
HWZwxvE5U2FqXxeSX8wzriWY52nkiDDUr9fyhpKye5QG55xFIZM/sEVOgYPNjN5QYGQlLn199LP3
C3icDynHBiUA70o73m2bz/mynZ+nHeEj8bMAkmn4mB07CeSLtr+GYTmXmzQTVUmYC+EDMOwQAoxc
H/Jx0LhOaoGrCAvQNjn/UDlF+pOXrCEs+1mvzjiKgEsE1IaLEPbnmRrPXsx/ZqZloMhfjZXf/Fqy
ZZm1UAw/QbghMPD8KIgXkB5+BtXI+wJVbSPGhGk1xSRofepYZXHE1IeNa17C2qC1ja9NAoM50PPo
oY2tVuwsZlXg+0rm7WKEpwa6XKt0rpk5dst50yonlYurr2eGLH7BmZvc9assh9qGUqeV4fGB6z4N
LyAnllIE5+Du54Y/bkWwymO0A9lfYT8Xp9cWFcqvU1/WPWtnsDOWNGhwnzH3oaYtvr8moLQy+mQ4
ah6NqkzzfxLoK6BPj/MavNJcnbsPPAKL8kEq1mXAXd7uz2mlU5ykkQoEhmDltg0Pt/YXG0NOcAWt
LBXbWa/hovjU3eG+n+y8IpgFpl8RF0Qi0Su92aiNgqOdL0GkdG1TQe+7O/aRXRa2IQIKLZFXJRL/
fN9Q02MIuHWmKofLhjSPzDd5hSoBdcQrZHi9/eZPdrSBmodqM9M8V1ESQuBGWa0bzW98aOilEwFL
rzi2fNXdmBFYc2kglRCYgzVyPji637Avhyf/zcNtObZ3ED73LmvY+lh7prFV+TLbuHKSx0hMPimq
65ooDsZ5fQLZt215o8b9KG9iIZwV2+G4+2URQAFMsNhnOYPmpFe5cPKZbQE+XGmCpnrKPpzE5i0Y
CDvkaw7/rOjnEVu8/VXAnFap/v3b2LTomHVLXiRcii12K7SyzxMf2IU2OzLcp5dHK6WcdPa1ntLK
XInNy+tCg0kkrPbnLo4xIyqDlnV3XN86JmgdFMoGfOv4u9PhK7R1IaKiPPKFu88Z2fsQ5DX1YQu5
RJEvcP2ljP/hNq5gTUqaA1M71ZGVVqiyuRVwTyLjIBXJllxoToNwfHaHwMbYQOe+dgJRCcxpbVv0
2g4AWwxlbXPthvumKEbPeBLeitaC0VmSOJA+k3Y/HP/NGjlh2yJyr5c9A5MOa2efMppxoK+c8GKL
TdWXr5/KXeyd9TX5F3LkPrqGssAVJvwtItUhOb+xa1hBwAboJRpGjb/4aGjFhGK9Z576TD7skRfd
HK/p8SfU2ug6xdPKT1/37DlyWldg9ClnuDlz/XMVFIfCazFOeMxbe+YpeU0X7hnrE+TB6YbPfx7a
R9KI7+QzFdgGn4YijxwjG3GwSatXpzha+j04uvWuuzT9qRiV7KYDbJwyazFdTlchL6YTG7KIXfaP
zdZUnQK6R3sdOgdN7qe0f5eTLti/aARSJfZ8knXLte1FPSgggWDzJyONLmqylLBdEQVJq19QbmwR
3fpr1+yHWrxPb/0iG/t9+yTBX7xDeVY0JlY9DRhcQ2rlfVGGRsWZ4Hp5v3bsJsqF/OtORs+MKKaS
QqrYeJZPLei3X3l8KthIjj9U6QrbO5E5K3acid+40oc+ThUd3wXt6lxH+nWHV+rhNjSjrSO5e/Uc
eN6izKWP3Cgq1Beg79nQvUaF5XizG/Lu3vZVZOjK6OSZYwSbUaxbUZbkiJ77gGoRf3n+GLJGKPt9
nH1UVVJzpozP1rqUWgKYgyeodhl6XLg8mn8F0pRiO2blBQr+pCDzxv7uPj75LdcwGdsHdZqS7AKH
r+Z/E4kblIxfJR49JUNIykEZg0Oy4P3MQesLbqNXgdmlCFufCXElEsh/Le3GOSwU5qY2siRaPXFc
ViXmbxy2j8sRY5ge6mVHpJE1yGiP6BS6KIB6+0kLUouPT2KLXYCyvDQDwIPjdd+41r//O/IH0Dk7
TuqjB9zoulVGfqIZvcolg5Mtzfn7yBFWca6enU76tYeZXsFE8Co6aWcgeDdJ10PHqAdMj8NNOfFX
EQBXQ1wQsAJ+mc7NbKNRvjbCxcfuqCLMr2nGbXICbA6zy6hqGYFRnYbwcNyLyt9RTcgrqZJ46tHc
gdHDZEnbrxxIEc7zcYLSBHwX12MBrs/Q3UeljgG2hMvNY7IHYlVa3FukoT1EUGE0hCocGBEODGUa
r8ZV5rcVNd2R2zIn+qBgCe5QVyqyqMvURwUvpiU+m0+taUj/x1TEFKf77cXAEiz61GZwn12k60bY
I4YOlR2fzx96t1MzHRq2Cgp2J2K/mHCqWPUCtxSOQkc3R5+B/R1OaM8wUIdjluwzudTOaqRkFzw5
ybAhl3gHGQVsKBCewADzZN/3OBBvOQL5W0xHYG06h124hOu84M5sJSZQz+6WFnRa3KkjvDrAo7bn
2QGm1tL/vJAhqyiKI31MYY+85CC+AysOib9OhcbgZigUJiHurSJZJ7R2UH9Sq5W+ScpR/CbaJ4VK
yxCx1FIBsluU1eXRlsPPBXh/lKUWKv76PQmrwtBHUDVVCbig7lRuxK7pZbMJw8oxsh6hBFFzXKqD
tpxRMlXFvLXQXE6uOxAKX2w5/3OseGbQKcXAZKiVfiW8iUCWLaRqr+XzuWGbwmET/le36Yr/qdv0
8SdVRrUOJUY1k57a3DvchwKjLDDuQWPfehEFCf+RX/5JfhvImbrNToeV9lS4QleURyPsdWcIWx24
D4Pt+NXSTMYAsbGBUihGzmOAXJZK3Nlz95dj76NJ+By7H9eCIwSxPfeT7qvgl9s5OQmTwCjcnJwY
oYoMTYpHMFjyQRjpx42B5ZhEASy6z/Wkhfc/7QBL2MNNdptIebUATNd4ImVS2MX1jgZu1zMJrDSf
tnTxaN3dYCnLx02X/tkNC/GcJWG8ofQCSfpPana9uXadTdf1xin0GNKrDpNroZ6qIUxt6B3SMh/B
dw7CQw+VmBa5wyDgQ+ZfG5Z2joXHmchKgPrZv3kfutCeauc1SzedUV9Z8T7SFznUApZLV5lBSD4H
8Z4aFtzePLkvfDKreoPNxQpBOR4H/QIIgw+7tEXyk7B7DemQvWYg9o0Yl4cpjhDFpF5t1kpPrIN8
NdGsTmcst6mGrB9nYvzKvteNB0YMBa98H4mR2/6SF5bn7y6EUiFQLR4IzeuTSm3VW7hmbqaZReb9
eyalvtUjy8+v/HlPQVx1qQh6FpmLww4cc27WLJlThKfdyHCGwCqI6gUty1Cn9LW9DDFwlIBtv/rh
MZsidex9VP73pGlhD3I25gspKcKHeOBdXRpYo5TIJX4PnT8iDGVnrUQBClX9iFu/i3qsefDfX6dh
zHRlLNJut/84W4yFX1LxFFieirkAeGZrIxDpwRvUNLL7O1H6XBUeSUR4N3JKr2FPeaLGvLWZLA29
fzjX2QXJnmJAYSe6VLVR/hG5V2vjeqzY17Vg3S+KfkEeU6t/BO9XUwgxFF3qijbbj3tt5mYUa3Qj
k1p0iSgIXcHFUKl+kGB68F6B1jlvHSqty+KMDifkUzVDbpYcj1foV3+Ewa0FHVcmTodg+Bl6HkOy
6rhyw0rsuH8XZn6O35npBZnylrFk8kt3nkd1/JkAG/B5jcW+/I25vDKmGjqZnJZepBl8ncpB+XZg
NvdAqqUMgu3tCtsXtHclOC+DloK+UD+NBR5yCgr3r0Ysc7E+KGzOAnWlBOwIY8PXF45Fnq5Xsvog
8kPrhkKJ4xpmONPOAWh03sVqoLnZiWSWNJlr9eyCpgRyoydLiBOXf3OLgt73oD0UbNf2/Tx9x3jN
WaPrWHZi11JxROHuQemIYPxiOo2698sVGGXI4N7HKYQQY/HzabPj68ppq+1zO0LWnm/9VP7Jd/+0
dLVl/mFSYwkGMH3XDNbptsgPw1igp+uGNu9+RADDp/yGvCpmkeT4Ep/vBOEwmRZdkziggiYhpUPe
9U0eQ1iOrDgm05IViEy0QP5ZhLVo57n2+RB6lkEwxrvVAbOS1FaQeigEfWEdrKGBKgQX0PUbbNO3
tjn+Yoa8uCJXB5dOuaUUKMgiCei5OZRqtpa/y5qZV5hsw0eBTHK23+VIRGgrP/3SwUSAJ6U/Oy+C
ArL3auIbEPlMLjfBJAqDTtwyKiSs+TnA66w/HeuMPSgqYwDpIBajUtO8dv8IKrb6SEnmagILXv1C
jFarUNkA1ow1tfW9vNtevJEx8+eQ9+eM8msCs9vNmCLxeeR/6O9zTbM2+6s3bc6YzzN2AdZRBJfK
8aRdKI/9Ku6C1VKGHpbuqNsd08iR5HQVrkKbjUzdcNapiqXiY/INRpuHJUokvA+onyKaUngZVS7y
V1gICEu2m4PUr9/H6DT3Ll6iOEshwwWwG4uSXd1HE3iAotqNMoYLX9Rm3RBJGPlPijkV0SmotiJe
ptN630IpmKWkzB/QVBBckPBrDJtvx2SrviNBdtgGbwT0tR+/siN/rzxplMNZzKQzkgu8vqVdbzgx
zwt8cI1R4Un/0Qlyj/2msiqr1bvbb/Xl80pw8HT4oF8Uki96RUCqSjIFmOTcJYBUXjiGWj7HgEfu
RgzyWTamduldpFzEzpa8J5TyeVBKC04tkY2redkH+8RjPsj0BVh7jUaR7yc4WKO5U+nGi99dr6Td
LzDH6rbSNuZJVJikVc4l3/eRwNj9KnpUU6cpNQWJkQJtIME2nvnYaAg3XfVI1Nzq8CW0MpUcbQLW
4lXLJVmJMFxLN7UkRSIFZZxbnEq6Zi2tIJKlSN+cKc6czRn4td6yohVm7NHHXGgWShc4L9ktSnee
dw2I6nAS0dtx1GLbRA4K+jYIeEvPlrH++8rstAObEqGp3fxv5mAIBEmoXm/k6AYRNjtohp+SZ+Lf
CNsxQQf7l2EmqnaJ4phv3dgxrlyaVNNfjzbh0ab/KCNE3rmSnMhtuWvy6+BGFPnrY0Ga1+5vqld6
T7hka5pZ5sofyzvvcTumkRAL4O/ioIpwdDiLYkXe9RwdL9ePyXLsZ8HcpKbYL7flYtKjkGd/MMGn
oU/JQnFYEZmyPHmyOSRK+l4A8YfLYVhVO0kQtQQLz57HoDVFM8X6XxxJwoxLhXHRkms7AOFVoBLd
sAA19de4WeuqsYjXagmzfjjSiDvR68aG2XqcWn56r7ySsQTNudwFYTDrCJONJAAaggPXury0QJm4
fo76XDOxWKVbwTCBp6wwrfr0zpHiOZuxiQqGpAD8BhNFKVh1Ov9IXrro+l2B3epceOiJF+92r0fk
5J1YecyT4zJ/hBWbAgUPCU7LDv8b85JyhHz2i/2tW0SzV26q7KKVduDar9PpgKnCO2CGW0z0rMIN
uqHl3BvgSXeQ0gbTMKNinqzifw0gyq/9zROD0YR6lWk7rPF9THTrVDX+nhvVdSoSWWPOV0h8ixbX
YLzFX/wXW3TEONMIJHb5Qd5/Q7PhbPChuwGKH7ue31yLv+SUgo3ERbEa44mCxxMA6yRxWvQvh0hU
a91vDYMryF9jRLDGBCxIabQ+Ce1YVuBcSYrhkbkno7eY/dinUKI/sC1vFJtt/XPHCUa0nqwWW96L
TOC+Gpp2s3EWCxmRNGT+XuMXTcs/qVeeFc1uYA47gynuZonkwcIwaKEQeb8mjKG2tw1J1ls+r3Xh
04WAp4G27ihIUIofwypC6w1c5yOjVed7ojxIWXDyGA2mZqeVER1IFCUzCYIjOpSeNJ0fD1D8YNyK
35xCUwWOmmHeVellKh2nYWGAzVY+eBsMPVtphj9IfT/sGlK8vo07hCZi/DckmmYY7fQy6N3wO57k
Znra6lcSoqvfEkZwSs4Cex4pI4m9xyLW/mTAZhf8w6ZGtDv++Ok1Ucuw6vEBTEMaNoYOFqOWKuts
YWJ4m9NFFxuLkMou5YaPc2uMEIjpjbospccCNVnUbjJie4KMT2aqHRdCIVkBzEnXjVmWFcujeIyi
q/no79ywfIuL2XqWnN3xGWHlGplW5nXjz0gekBn+jnZAS+d9FOMSvIVAWlcdIdGZKEH0W1fBPvWd
O5waDDG/evU/hGWJdeo8lkMvVokXh8e4YFzfFjb3fN8MoSXVaWzHyxGI+IaEYsuTwavBy3j5GtAB
n92A7dSiLPBQMMAu9k6X7yIegFT30fUafGTzuo+GhHj3/VlVyK0dibNGoFxnFo0ZTkQHQ2s1dHpz
zFZ6I7isYqanZVon+MV+r320JdVdiq0gz3K3KNMff7Rscu+4tauXAjvkHEEV31UQSn5HmROO+s4I
vTPCIUxMguEgVPMTtSwbEB1h3pCQYQWNWrQ4wZ0RdQTmydqxVfblthA3p9rD/remt4vH0+dksrFT
VFimtpp4Xy3fBfb3SLB5A6aslUkJBlTxPN7fi+ac7Yz60BkXryz50bSBaWTWH+kDPZ6w1sA3orKX
ZE13XhgvmzNm5QXrHfKEgq9eNy0VmL7ZqyvJmztgRq93q/+I0wYl3ikomNXuw0n1AOqCuRFcoBaF
LQ7zzE/z68Isi7CwheJ+qKuvTAoDVjfHT0amxUUu4W5bynrdjNLfNcV4OZamhbGtaSz49T5+WXUS
JfKGlDYfknF9F5DIwnXwIkgalEcIWGs32SnR52ZYKfrT07ItTGYEpxx7r2woykWxQEWyFTYyuipE
M+UfImVhkmRl4po34OmTjbkMz641hPyUQOcizOOHLgJO8F3PB4Y2qSKTtkTWIxIrFtHEd7Sy69s+
92fIE4HMjo4TXypEpdPNctSwv+hHd3Zrqon8QlTxa2d76c5BOVMaWuh4+AH+ExOyso5CD7oYjyVS
r3S7tQyAJBPVOX8nW7rWaXQmB5xBGAxDn4VEfw/UEXxJCc3Nk1nQhWiFh2+xSFW0PH9QX9uxNJGl
4NXhmOvtJvg+60ymAb+lHDJsOXBnR46wNksDDufLYTqX9Niftp8bsWl5yMjMedBemNkuV4jMpYQB
p8rkHQglaitqMUz4yapiYQAZjpZnYb1zqppxKCKkmKIKIKSd/3+iJEoOPyhjEbyfMYb1guz4ImJq
YjpxEVIQQSyh9Jd5E52XM/uQSQ6zpRSIx/oQtHGIdzq1d4Z6O8n7tI6c6gzpNo1N5a3xolinthr5
PykA1PBFJGXhC1tgsbxYEnONbts6dtjgWzL4q9gJ+xZVcQu3Kb5Wx1b3G54VqvG9kUuvctumBwzl
OENy6sA0eXAr3APZ9sGQvCxtad8pEjPxJu+10xUEdCYQHSyC22aZTSULMQy3cHlvbW5zaagIBrqA
R8Y+wkVKTlsAxxTAyqyhammUOYj0wzd1QAOuqcFf9Iw31X7GWmsb3mI+l6WIXYW3+ZpuoVItAhGI
nantWudUDy+EBcYRi86SxmIApJF/kA83EGW3e9J8JMWMzrYEirvF42Ze61BLpfBH7ZpRmHVl3FGj
EV4zIAuuieiknxQAkd7NiXNCVsgXC2EBKhAfE7wF8HVBubiFUtdHJ8SU8DZu/05tZ1hCsUfkrjLp
oumEnJmpw6sv6ntxDxE5d3JIrMjobABJaQoYykp+uA+YARTgA8uUwcA0TBIDGQlDj3Uz3gPs2Orj
f+XPTNV3hRD7W7NOzX10N/y5sl3LXVecZLlzMgoY0C4Y4EgcOwldmfcYEyRjCS9GKsvnigHJkh6o
Ti+LbbqT3nH7xHkL+zpR97eu9Dtdl8uWUoNlFQx2FJgvOoqUUWzbVQvxYUiFvTDd18ZE9APXLmbd
hUk2N+lArAZ+IDo/vV+rxWDaBLBCj1LXbIvBN9iEWRwnn/D9cBIgi71CQCTYHJeO0XdLi6bypb1P
nvrUqAVc2PVxFsRNq3Vvd4ZHpZQna4696mXNGSRR1KMenEmoMOevOf4CSNa8C393/3AQjY+7pvHC
y0k5RheUQnv308zgOEZVZtUbFLTIHBRzSrETyshJqCiA9qkBG/SLBvrCfAutnmfWtMOfRhDnpv5K
3uXzDbMScNnOharMrk3tASkKtTg60nHLnyn+TmQ8yODdDAZd3lkGzz8/FgBg20cWyumgTqMO0tyz
hrPFyLvjvzZTdcckzFZsYCKdDmvRf72Ls/zj07A4pO0ed9zN646oA6OQ/OzkGsHXJNc7p06W5i2Q
heO8R+X5H76G4PFlgcO8fSjeg6cSOwTQ+i9ITF6lhP+8X8mBjgM4JvFNcLCZLQugieZxcQF9IKNb
K5x7/mvf2y36i3M28v04M1VQbpg8IazWHE+kXxHPugXIKurQN1hSO814Ceb5gft6ll+a7LahhjD3
bw0IEb8rsEnHV+VkrGzltYDle2lx6mmCbJJHh/YmNTTr7UgElCzHedF4DiEIBs7SGM4FBy+JnTye
CHxsPtwuc5UsRBRDF+JyS8EJzxh3cvqHMpf7kBke6R43ZGSCcdKTru+LltkUmACWLpEL4jDnvIYo
iHJlEEJiyDDYxVtbVBdSfQe3JMQbWJKAid8KQJJN9RY4BnyHB54Rygu2oStNQ/r50mCIsSjAEaFu
FLj1VncY8SyBNWNo4m7CuSO2sO19zMwyRywjPnOn4WfStDL56O5OPb7Tnizp2edmEDQb28rjogcs
/O0xoolBBHT5kVwnFI4C+mbRrwwmBJlZLSLDAzjsUaiJv9c4JWjMMgAcqgC+PNgBYYDvm3ycIs0S
XJpXgdGB+AIIy3w7iVmS5WlzQRzqhysWdWDOzhpaintYDuTka8SLYKOBNs+rEY6Q05ImFLbmrCnW
AaebEQ+jZ3W65xlzy6z+GBeafGKlffAIz37PzQYSlwAIentvKt0gFqH0lj81xlkPKhrZbLPqR084
uTT4rVI4yLj4J8hRfoNB5vnRO8YJlK3U3Pj+YF6FVuabebE3SAwa85nr1G/Y75USRwoVD5QXZvzc
q4mE8oRl6YpsT9aXH5NBN6lkLYhxnxusjXPRoky4tzS9pjecPK6p7SERc87aBmtZ/b7WN8CNQ8EE
JwVGj+WPhH69cL+4zx4h8l+NPVpW5M9EyZCK5w5ROoaRUFUWADftKZ/ycDk6xLQQElb8C1CrD7e6
NQM+vtgVD2ih2jJTyNgJdM2DH6MYehV70zoDaamkkcxmeE8cy49RLLWQTee2tW7wrd5ytOVeQ1rg
4ZKZvVETpmnYkKzC36t2fShbyWNll8cgM0pzN+HCICPkpnhr7T+w5V/uTCqfvBPIsuzHwS93ZzmM
teeEunf8AYZWGPqAyi+XLAHkhEzWIcHIhA+OrYqMBXYFwqj66u5+zc2WDb8pN5Y00/ddKdJwtDW5
jTDNGjKsKBMX8HvHYqNoPm6FtowFw+qZCGMwgc3MolHYqWyHt4tcQLzHQxnxyf9iU+rLgdhasvFD
Mt+ELMvo273fVhVK2XlIBb4QcfJC0smgq85r5+H+JjNToXRAWCBOET3IXYuGOCqZXSesfF+hVFFG
mRzp9ueu5hct3AADIkFdhA8C0GNSt3U2py8bulDJ8EzF4WI+zNGpcBJ8tVDb8iuFGon+92CTBkI9
oWuWrCoDnbguN2SqtDZPRA/J2ghsH/1e0/wjqQBm7VC6Ol+vDJC/v782mZAhn2K8zcFfZXZ4ymud
jevjNmbqgv/Jqx1EJDdNorULs/LVipF4ulIVaTFZU56ktVkX4/zGpgi9joA7mYzafPuB0XbVxgPH
AYmyEhQcBxSH3FANQ3aKvfA90WjxGsHrNTuzeLlvB/NhTg7iaSlNFESFGxmWYVFizTrQ3K61xRMM
4Skv3d8LH6alPEwLfi/HvhgZ8tjUNMJ8YaVBwQhwfD2xlouiH2DAxT2+byzrzhiV25qniml+X5EK
SHUeGjqfxjJvMTKLiYOnE5reiAQmM7ZPoRDfUmKGMRrV8C3aVcYlWpPwfkPD6SBjyx49Snq8UEem
suPjtQgBPZBmx6m2ZBYmPjnFiWEiAjImqJhbbanRNOwjTAmcYQZbVM1zAiPJEDoXWrBvTZUVE7Zu
0oUN2m3e/V5CGkFrxPdXqWS/En0AT8d6mgY/DFuizwgs49yjKbNsZlhML69MPwm53YHU2LqPV1uZ
o4Pgw0/6nZEJ/Dak8tY8HHsc0ziiudQhOMW2LEoQp9W7udhJrxohIFP+g8UEmg+oT4kxWOwqD2zh
o3BKKtf+3W2BMNKyV4dMM5j8CrPh9C+jgMAXB8v+Pr2w2abkgiHNVmHQjP448vI/z7ushUxJU3DI
/eLjoS8UxwoBIL4MiRYovxr32/JmKvdC/HqZeyrGib0QfhLYgam0RKzM2ltbLwNrM3B71aXXHPIP
DqshArlU/HVbHXS5RsP3yqJNDVoxNSrWXZ/4xc6YqJ/ZdzipBsr2az2sW1dFVt/9SJlh6w2Rtqyx
wyv/90QMUtnWEIBmzVj8BRILqNVhOGzL1YFg/tEKb/It2BOCkceZnPFPUB6avTcveQAfrc51gRC1
GmPZLA8FT1mb4wtw8qAFS0Ir2JkzOE6qpMay8ABFrHOWOsdw7wbznW/h3KAvX0uPr8Zq3FmMUPUp
oQZGG3WqKELdQ4CqZU8kyO0obDPoZpELR1ABdRQ6cdVENTSNKH2d8jsoBGbDDHK6qgfSnkaJMDzG
GCM67VYiB78xDuzNoYhBk5+46DFrgjMXY0zzR/50EAb+JnZLEGu3t/MRPROA4g0d2XFUUTTmQd9t
WFW0e3Xd0WchGE4kO1dBJEsr8fbL1Ip1QJ038WGHQqHEPVKSE6HZBoOvatQOuaFbEuKPUK0lamnp
rmaLBk715YIblemXMf7soCyF9NVNYfHB7ifnYT0uB52b+9DpGNjR/bQN6IgU4qVn1s/ccMz+PC4Q
HLUMLeUvxLqhmoWketv0iW7+gfYapnCMq3Q/WpPsoseQ2HnmiuWyX3rfB2mKaD8zqPY+4eyUtzC5
eOEchWWZMvy+lBU6SuNbbRToKrTMS1TmyXXFasApdrspOKNB6ZyZDJkUTIeG5D0GZRJT8WGvhdJu
porhRzHpnOdHDY1dqhIUxiqVJyJhZcvKSoC4smsi1NT2qYkPfuyeJzzifo3Fns42k9MsOn/+F9jC
WSnw6s5Qh9W5xSFDjvHlovfBfJaiOHZEwct70BDq/7Id3j8VTQt9RCW2TVzyyOu2vDWS1TspI9gM
/NPpxj4vL7HT9OvcmenlQiTiGpAoZOYDkMXDHSUzEaGwr7sAzUuQCEtDfQNIGkaQ36znwJo5ET0D
zo69o+LLwyHBindh3VNhjUp+y2PsJGlePEo1TRSVPhuuIkUBV7ox0+P9s1bOQQPtHiCK6s09I5FA
CklBOfxt+U/V0IeCIi/WMdINqM4zMe2YG/CeDFcoxDWbTQ3rTAiEPcZWnj42XKNykL65lHbeN7gJ
FOpjqlMTFWvtJpAVM3gRfXITZT9z6hMeqMRi3vGF62oyEQcr1y4vfdEEXaBjPLRrbb3Kf/sIMI0W
ejIosm58J/Y8PNyQ/fasZHZ3bfEz04ZsVA4q41/9wu8DCkOCrXEB1DijWCBpqyqVM8W7nAIWBt0V
4sTCZ3arsnyD1erMvIDelodrEzAXwBcT9E1cbdNBce5Pc5L4VLRvboRKSvPGIKrwezUeCATOjBuh
xxaq9E0Gzp2jt6rQgIUDFcTcYGcE3XIjZCij4vL5wh/uBEfdXMIys6wINEjX28Km0SJKNJ2Kdjx5
mijRXsNsEc2OVIdDtNi9K+9lsxQWwIP9fSFnmJhwxn4wlCzx0KZkYxzWzRlLudZ/RS58aX9z21h4
1Q1bJbpAmCq8L5Sr/Kn6kqyhdLF+QSVoZBvxxeoUfLahJVPmcbYkwB+4kqw+rhNrbCFWVRikh2kV
p52tAsIqaZ/RJYTQA/ZuDlqJ0PccB3bEdPQwcrD85rENXBnkOdBxo9zK2lqIiQXtA5EvpiE6dkd6
bX2urb14jYsia4ns+A8lkQkqSjKNOpAJEaWrO+hDzEEU8T2j3Fy2/yDXMOw0k6yibajf2eaXrqaM
9ecm0d4oZcHRFo3G+EVL2v2wW3cDtpMtNtuRgUzF3WwLeTS770d8F3uLE13z/zjX+4oJuFWDUmg9
TJFZqkyeXLTwUY5bDHnYqNvbTUIcMKtBmm+7EBu/6zrXqJnhzxmFzEPmN86GnM+AGYulT8bmjuQM
sX8Cg9AEMEYJPRq7AKXFBPDLbBjvSTqLnhJyrdwY8Nr08uFJsSHDKMcHO52WSPg0OUycirT1LzPe
tDCl4TUWO3OYtv9jB0DK6nhF8olDbUCm5wBM/uxV6gSDwLkCWmWkge0NY+4qscR7cbYPFNKIM4Ob
tV6TzgTgS5MpZ5Ft9/GH+5BWqhxl83LqII3ygy9O2xHjwcxSL9o5Gf+L/SMTy59QxZn/+z31TkUb
S515QpPAez29EJcHDG/smpWgRHizJ2W1lZus8dcCwNRYsQ5Q2RLQfauJ3XCNa0x1ePvES59P524g
o+Dt1CZ53a40P7KtAhZlo37Wd8Ow5wsmQnA6t73f5WHeK+UsfpPRfqtePrr+K3chIG/ZwzoOBFa/
fSJyIjuAl36mItlQsPeJW/saoGlxleabM/8iogkM5onr2ozgcoQyG0WGQIleEdFU7oPHPqu+HPFC
F3cD0fs/4yW7VvqfXNkBN8hKtLchcR0lQlqQrFwo+k5CvAUIQRsV9cM3T9iymXHyIYofmqohj/7+
nyUIS9n7j+wjiai3L3fhj+bElI8fM3ILryDyiRB79jPU5HmVgvkE0Pl5r9H1O2FqJJD7vqvE4GSB
491SL93JB8LhE5x9bpFzpdN1EAR6kBiFZxvqNQAgAm885OMWbInutERpjDzko0j/hsgiQ7KjeXvO
S/NYJY43WTYrNcXzuZljBNBli3yYHAC32HSAyi6OmjJMTiKoOFsM8GDrKHL3MzjBynm1Ky9mWKQp
4ndrZGh4cAbJ7WL+yqjSU54Ktm+bn7lU1Yzt0CEyD29RO7Ah0OFBXHoc814XPnrAgmtOh6c7cOq4
jjWNhEdzYgyWhsrYWKjbL5h95NwH/Vvq0Yb+eEFytLCa5i+JsLga74nfWjSGWPy+OycPIm1pTLKl
D8ONLB0/auV+Pxy6c3TsG6Lv66jnvKsEOwNa6DVOqjtXzaykCcZVb7U1FC77v432Z1wQ8adT5FPS
Pu02zfH9TJ3dcElQBbDnYRsaJqO961Xxf5nKbMjf7+Z1JW5t5GwYTUh7Dygztm3zMFyGeAOvDTr6
cwlBfsteEqMlI0mPi3WAB68rQ/vbSP/9V11S5pKw3iw7GxqCpKCvIlwx1OAeNPnaeWj3fdTUOhfm
AWzMKib652LMw8X0yTetQrVzouLJ7N1camAk4qrLdg0xiX3SCykNiE8yK7sqFEjKwPjgSH4WoH00
cyHTe5SxJjphs/UuLLnrxgaGv13dNj2AxQ+RkLkMoaTlpMMAYDMCk2sXtr36k5FXcH25Rx2b2+H2
ShWEKqyM5OTNoH3acaakw9+w8MAEJl308euNqHfuWaVVoLJUDC3+XtYAJ4UGIDDUFkg50jZevwtU
KEobf3YUc/quLxA75lKOCCrKv72e8nF/aJfFCVcCUZg4dK09kZLdIC3etfPRJLZn0SWJZ1gTXglH
8yV5qHSLPLuGFUNYatTHXe6w+E15RkPE20SqXIJd94WsP+Z6MotaAzHA6n+W9y2sLDw1x75Qf6Xw
Q4w8hAz0LnzV85MLG7aXiPRa/YKBArm2CKHyo/1CHkVLTWpa7MIHNzNvtrPLidWFDmPu2GCB2aqB
f7mt8WA5fCyPJBdza2JWQhwBvXX3Cv9H+BCY6MhtHBNBFOBfFPxa9N7O+fgnZHpiwta/LUxH3GOb
29Lqbm/1jBF/XeC+me1evmXyO8ctR4vJraGzlVnciIChFNGjhLEPpsPR4df9PkOL1EsecVcpJSTp
qr+tnCcTzx5uZeXEV8jlmUJUMl9I8i0Oitdrw/3HRgsdHDho6TrxL2D3xdaM3ALoradb/5UT/6WQ
bQLEsX+Q7C+SnH/X7+hXRdn/xm/w1U6Y4u2xhOxdBFbFkQhgWJM25WUp60cyjDuigAxN63H+xBv1
byJNcMFLnk6ICgxeHQ64jOlNxQ6BSNuWJWN04voUmwfk1Qhd8YNeoO2HNEMVwkVW1WU83S5aOOsj
Q6yTFd3Q6W5Pju52GulFI/H8uoMWffLTlfCnm9N7kMk8f2WYwTNhpd/DXxDGgpnTBKY8yKOcQKAI
JCdML4OJCS8mCA0PkHqp4SKi6kz3iflFIPOIZHC2wLe2moIr0eEKDEp945VvuB+2iw5tk/MBjIC2
mPDxX5BpDj7yjSz3LRtO/wY62RLJNEPM7VwXlmDg24PdFrvhpX6IXGfFF1GeL4+JhBeMIf5XxVEY
Zq+qdz7hwTlr8t3QPv65+YG9YH6RFf9RHkCxyNzORfEDrigdJtxt8gKI65TqVI2M6SiiX+a+sspx
KfrICWYj+yjB+eIoi5NMRZGIalShvUonkEffXptYcJIG162heG0Gpkwa8c0EQoZpnY8GmFyt5C2n
kjRC8ellHnCjNKSfleYdYpxCAh27C23kUv9REgR8IrT5cJogNCE0WzF5JBWiwCstTKLmJ4SW6RuS
7oEAZH5/jOhhBE082my/app9FM8CWK9dUDTTJbJG2HeCHGpYusbGcWtVas9j0/sgXvBV9VK67uNU
SYaF2OtVOu2kQMPlWnWSC4WaSzPopAbGmPuHZxbPucEspJ26Ejhaiixfg3BtcfJz5HA4/dJ2Arkk
LwEQDPY0p8OIhRIOkNB8zR+lhrPvVqe4pVDZ3VSghEYrYebOkY9kVbzrJD2NEU8hLRuFIJbeT2WP
vIjyLIExqgCt4E7lfNsbzwxkEKVYIzjIb697BUpSfqOK66GYhBP34NIrFn2hdr5gISnSUhM9TLwG
SPOl9nNCtUsOafRh9YrIDm6AqkXdTzHZb4xMNdIM401RNfHdZ+BrDUACqG9mJCcKlSOKgioMWX6u
qDAv0kGo3uQNvQtqoqJrvVNZ0ddBO3rW+DBH3hgwb4nMNlGQc4Qw3qZtuZwNa2Hl1KXc6vflh67D
xkOVzz+irDvzudSzfYYaV5gcqZV4NgaNRZnhB9wIHlfU9/hxn3P5xIacSRuKeBw04zsB4ySrGyaw
aEB7Ov3gnEgR42H6nN5A/ucsOAHu5p2c2HfqSNz7KKhIXE4HQKOwICUU7VIyovP8Pl2+yvH/2HWd
A29swsFTtaNGU6bSj+Q85zh6mN922rxut/fPANwJFyjdCde8tX8zaK2ptFZ/PWd7Xh6hp5ipQ/HS
Ns817TEKZbWFzq1qm599lWtx6ob+MAeDKtEvhbEqsZpMMmmWULS48jqrcLL/6yGQtpjIFD2XJQSd
vqrjs6G6vWmiTzQIlfWgjR1TCYFwELVODWEl5cDbcgyUMxEZNeIDDqgI08v3a79cc+OGAx5k2N4+
xH0WzylKMdTMoXRYQTtzTZDgYrds+DJ9cYFz/01YGPZYIehABVCvP/wLHILu/GO/dDwv2J4nq+Kb
NpnSkXXLY2FoJzR8s7hvN9hiMzDx/cBzMZKvCTdO1NkUOUHvh07VQ5JXAOaeYe0pmLN0tELWYPHW
Dq61lXbYjolacZx0X2z8XXh/fi/QZ8APw2hDDqGImWhrHkHU/SlBq7/OV/xYGkDbiGrUixodT5Vb
vpRmlcyEEvUgrnLrzP371Ki12SaFtV1XCjZ877yG9kix431kJ2GLVpGTUdvlnuWNHbAdBBqhVGiv
YCAdyiEvRjmujRQ53gTGZw6XG1TruB+KVYbKdzAiTzoLFVIbD6+flXQA1erBiYHmZwh2LdUpDetW
ukJFZIdWLdHDyJjGcaTeBzemM1Vi7OG467hbnaYh5ltfWg1mOMxRaXpqYILLZzExUgUNI/ox91pJ
b5fWWsqFFgZqubChwijD7+kMozKYEatcmny0gjfvFCMFa27TzWfTUF05xs9hyD3XxxWqqX8jYnr+
sYlbPF0TELQnQeonJzUYsad6+o24rsMvyA2CXQmy/nvAZdwIoECWEJB3wi8X+BWpreRsLVPgmqPA
9UrlN6IczV+nFnuP+/+KwQ0Jabvq1Nz6KouqB1GoGTRQWXPJ5eQxJ9pV7hEL63GF7WMS4xy/FdE3
yyJck5sKcy4wNn44c4xZaHyCCYYY8d1J1KgbtpQclRnWDNLVI++5cJ3vjZ/ect2YU7leogs6Ndiz
i64ViIQcivfb8Y5Gd4/btirI7DzZP1zMaQz9ydxDm6TWpQd/Zdwdp07rkt8qBobUBl51rERl3Al7
fYTA1hUKVmKChKOF7C2TXGnqoIWiRzjWmH/SC1rqHwFCt4QTsGUjQ9goqnoNh+IMXKdwA9tP35s0
hHraz82uieeW1DgaRlzae3uev6q87I7zXo6AGW/Op86P9cZ50BNlOmSiKVEvqamNu/pNXJC7baom
m7noknuXs8tOewMwlqwJv28LouohRgH245BSVCIn9eqtzSYNV25xbbhz0KBba4ggSJBOkvfiP9gr
nA3XsGF7OuIM+DVHIak6uiXwgXaah1WAYfhpqw4o1bEd7fTmYg4n6hZEfignQUIkvMXIcXLwsOsx
XXzqq0NL9TXPm26N6pBR0nvQ9YIXPzi3E8iYSeYg2GJEt4ks1GQ+ElARVqkwiRQ9wf02pTPHnGZC
KE83TZYujLmUaOisUXA86JzoNiW/Q0u+kAraIjHlgLAG2eTp9FQAAyy74r8+xfFyR3O9BitxAKoc
KFOp+Xvg4dW6x+9gXDci6Jw03BuI8RlxdWabeeQ2Ol/BrvJC2mjMRJLYXemv7qSwKCUrPX5i9EG8
BQl/kfFhqjCxRg0obgDKkIND64ep+jFgNDucMp7LlUMROM+rDPLeDqQwHcn0bTnzacDFaEN1UOKp
U6VU2U04EviAIjMldBbSXzDg3JKExgf8R1/D87PP32cuWYDr1RZVR+KHD/Um8kDBNcDObJ1g7Bim
Uv63OjPPpP4yZO+8q/MqFfFtKP7QF/iP0cv6nTxorZPHhsJkwjQI/kACz14i9ye3wywReFwQIvlZ
UceNO1AdUC3YjfSz2QkU2s7z9siehyRRr3ZzwxKUJGbQOmOSq/MyafLNzx9xTyPDRvIZLoL5RiBs
Y95q24M6ZkJQ5niLn2INCDuKal6wibpauQyFQKWDEmLEy5y+M+qBPoATFNpWlNg8YukccGfTD2hA
t6WkkA6NRGd7oUrTR0O9MUCyYZGg9V3od9ie8Dj4uTflRO/x40Awn8qP3HHmkLG6AnvKxcU0MuAt
zkY5jXuXhmaScknT2VFXautIQq0bVYIDI54ys6RVNdwLTfj6yuEgYA04DIMguMr9kuSZXd0ZOfrV
3spA9W/wvOJVvYMF7CgI6kbc4/miVvSmTgRAncL78nD4hFWqV8Ry/cQmPFzOJWhiZd5yvYYrdFh/
lc43UVYMuq9cDVxFuksqURkbYn1sEPvE5GRWdfbxwTSz55uCxk9yxpZjLOGYpzYy0UVQseV1PkHb
rDauT8YNW5byGa00czw2FmDftohf1GqS8SnUmETWEQ/wfV2SYQhyJDwjp7UFIDaA0/RKcbwlP76U
WP+/jiXelF3BMSZT92MFWdZeXEcoGWNgOtSBxMMLvmQ+TiwLnxBSDDh7TBdPrK3qRjEaMUMBLb6b
on3TRP/GWgJ8C+cPs3yXHcLmWYJLtZZx2xGW4Mc9IT8fO5hQOTSH+zXx58nXAgz7ZTdh5RPNRndV
tbxW4Nx1x2zRZBeNlZz1NTy4R5ncTDiZbhHf+oQteLTsvMMvvfowFzMOMLZ4xXcZUN1VbDkX3IfK
CVFcX5ZDvESFRqyCYBVj5QJiMQUfeU7BBVS1CqnQtDD0RDW++ip2eT3/G+5kfQ+kfXcJacl9M0s0
Mk9wDE/8hjn75jdZCTZxeR3t0+Nhx3YrdwPn8XQjKKBSFgw7oxE9eb+2BXhnJf0N+HXush4gsATC
u7eI1a+INB87NagVhOj0vcaIncHwsUpBTLWxMplTzqUABAzg6lO3jsqeT7D6CgO1q8z/t0+HWp7H
jMZ4LW/4R3NpK+VDcbTtHUAtOU8nNv3NbnZKh2FJR6wYbOcJKfPsk6mna5vVuc8QlgAj8D6WG020
fC+vsOUbsSchjaYNuhfi+V4+TfPyjTo6GTI7lMQduXOu0ZKN4ox1QqM9dwwYWDYpN3imP/VGnycp
wxxJ3qlXXeoplYx5txVbKfJuPsMgrCR5GFnXLdp40g5Zra6eYgW/1Y9JVAVs2puMKSBKmNxdK7Z3
TaXAE0D1h+Bw3G2R0PjWei/R4cXBmQH77GwvTSLHHyOvqS/jmL3sPUezW+ATX6cCM+u8U1/qTsid
gCwlAz/JAV8Da8f64WLrDQFo/HNa5ffACIsrQqkNUR7oc4F93lyPkj0xhOGTnxJby6XNbb3vA8pU
/JN7LuT96utBQngoXcWf4H0OqkKsj403YVvdcddhUFUN28fTxdnUYGVuDCApP0InRe5vYq+8Sohd
rToMuN25YmcpqBkZPuFMIdXKpEjzzRPNxmjpsQ9RDj+Ufka5SXNREgCZYVcUqQjn9X+IPulFljqI
Piw0v2W8wG6bBFDZJdbeOEtEy8kO9BsYYSbj2poINXzXinkxZCMPG5Vb2xSADujKWJdnGWZkceiK
/85z5X81+oso8W7kbcLd0vU+DsOWiH6oCUJvi10CAy8I3XFAVHwkT2hEHKoGZp/TS3ENYcPVNOxe
N1oI32GGqyEsrplUNGp8b9S7JB6Y0hZMjJwg3EYGBK9PCZCe2HPrc1vzbNaL0W9OVb4/KSr586Em
vb+wBGMAKbId76ygh5n4+rY8UpmSAKb0V9ycQVZdt3hOkCP7Wl/oZ6C0EwSIC1XrCg1VE5M6tHI4
h4qQJuxY572+QIwzV3liQzq7Z2Dqw4VBAa5hducy8pRoNd86hRjzq2Ao/kUN4Ohi6i0+kW9O+y5p
SQBXQ/FtUt0pfWFwmicM+iZQPIgeI+3jRoLa7bzeRcF+6aOEFP9LkyX4xNNBa0IbPAaihy49Btw3
vle3wffXbBuqFOcKZZkNCx7s2f87xaov6lbM4SSsYA/aNG+vJ02flNwEeae3n6pb0iSQfT0LiuNo
sylpCVx+8qfvVd76SvwLC2yC/8RgOjHx+c8mr+uOfMqVF1R7OFiDnTJhBr8NktaVstJR5LR5Qn7R
0eikbjO6rTaMGp8n+g8ITA3m6DQ1pYrBiscrEmYlFX4WjcGJOAgRyZsbz1o7rfBMo1k+ECuTrfji
omShogLf1z6Fo9WJD55TyEOirJ8HQkQWt84pN4TKI9MGXSxGtAGmNe6aPDaDOupZa0T7CWRI3EbA
JL+ahd4oCTpwylzHGhfPelt9JeRRowLXxuhnWzNywlkdDv6vPGS7Osip9YlOCbGdz6xQVEAyY3Q2
B6Ze7Sn8I2ZniZiKFiBx8yGnnK+0Ry+otiG83QF+nV6dkjeqgXj8kJhblpTBmM0EofxQETfTaYiO
mtdgV8gAqi5uvFrtysmI5QBTxnOIkEqHtauQXzdarcjuqBQuQtI08O4FGOJIBTU8+LcYEphQU6Kw
6iqgyuOE6CY9HNB6VqZ5vT28T86xDF4NfxL5jUxTvC+5O7aoU8KGYNmfpWvHIAmUP+j8jLBzO7wH
I89HfzlGnRiifkasVa/tGprEB+MOCeAGyKRsqC2Dwjifk5breStETjChO48p/mrsQHWWFVKEzXk9
9b1L6eBkj/G+/A1a0/A78Rf2EEKVQO4B8G+04r0ERixo4uIJBrpuLaRh407eowwFzFEfyduhBByk
t11Jj7nd+MPCrJQuqIy5mkGH0cpXjPcuILXt5aRhCOv+jj+KdQB6QNVqBPNTBMcNZZncaxLbyi2b
y74+coCsh2iB09tbpHMlNrDbGmNo+UBizrweEqUtmCgozQPq2t9Jp09d1epsntumgoi9YX9I2myb
CJlhXh8qQf9ZEHB3rplyKAx5L10n6T9QEsOfFoW2D6adpIlnf/A2dx8DMJifGq3ZXwkU15cVXU5z
co1GyIgew44bbEhgrreQeieo5jbJXrlCkqqZEnocZIj1Ie5xwVzRBOPAeb0J6MEA7wXOUoUbu3s1
iWr+YziIx4n7XuWqjtqzjtoluCnovdRB4zE0Wa/pm1M8H+SqPuujkqVyNl8rrTHC5BN8pbO1Aqhg
27Tkbs3EyS7m+5bOsRYFaFGzVBBzS9rv+BFamPpmvrgjtI+IJRJyWQ4r0QdznIZRcnjBTP7wwkVK
kyGrMO7p9vm3A0bK3sN7ZNTI7R2hunn/o7FDXF92R6t/wmb5mnItRvT9yxP1X5BjySydV6k6kJKr
oIjMdLfXwHBuN9hnwuOZdOeKuPG/VZkzpQCPRvIJ2xJ85aIujQCuOWe6qY0jJNR6uZ/DagkIZBKL
LL9YCGMHaMaD11R6BhddrychWajTEVCjVUM0wRCvhROHKB77qWJKiGhc4vrufEZ1J7W0/2kqQkgZ
I/gl725ODCigKwWkv7mKXpTnDjvNkqY6QvW7T2//jmz5qgxu/2mVvvWi7l/og2VBNypRDrV1TKTH
r3N1yYnF8+64u8YXF78m2Kg7+jkRVQg3/+zIVGvYxeY/buiytN7EXu5UI+j0DUwO9RNKT6pDsuYl
simU8gIEST8qHvOmJ0QC7rTTDOhE1QL17vxUdMHmQYQorRxzvm1yaJNSbDNHKkXJ07q+svNJh67S
nK3b3fT8yhvdpSdRpSOv6nFWK0uqYni1RF4G4iPJbUaOSCeNXNEdV+F1wkDVYWuhiN8ko0RLaC3K
xdxzNuwJ7FYg1sBnfLHFN3ITwYQ+r3WmgZVhBx4au6yfMLTR7I6mU+DE/oxwa5i2HKEt8HlZvGqa
4gUrODrlsAzBn4OhiPeT596JYbH4br4+ZdgJJfUu8EJSFfqc08JMLcQGotYfVvd5PPmDO3SOI1SB
1oHvxxjYzmDaYxhT2olVlXG5rhOnNfWHWSnQb1x1GMDE54cv+4QVdHwYHwUIVgDTPzgHcFhePbfg
feLopmYR09fwzEGQ/sDbyPzOFzgY4Q6MSPuOVffMBq7ySRBICDrA+5jNSySTyChLZGLhGqz0M/5i
7+FsbYurOBqGsW7piHDdRvuukC70PuzWgvuTqUMBvJXaWNcnQspnhBZNS7sFvNikR5PGdpOGq+xA
dqhuRqZZ7TCOSV/KqkeBgeibcrF51dLb7cU2l0nS52LWaRvpF9eeY+A2yHg9Q+/QSuh8Y5Zi9c+v
FRlpUXICIcON/ZjecCafdx5l2PX3SYKA/1NMmHLim3rDFNTzUPaF8c43Fmz0rxGpfNZhuOMsVUCi
0oDtrLFJTWySXJN+JWp3DD3KTRK6Bo6SDW1OIUhFQK2OiAsMld7qFFWXBEo2EXz+Txrvk6LvYhgI
07t/L250h0JoFjZYWRG6NKSUHpnoBEBK6G5N+fbk4z2pXBrFZH0UVgX1mShOaDytA2AJnjg6WvNm
PWTbU1BIUSbdPWbmvO/Jzz3XC1X7H2sSgDIDa7QaRqxfmWdPd5DLWOJIyMiPNkQxfYQzEoMTojsI
U727RsCTIFEJn5hvdH8plG45CcEqlr4u9IVxNG9epXujOWAoQfiuqHJ2rZrM52cWtltcAWyuXd9w
0O/KnQ5CCQTA5yKXx5qvpaGy6qAdUo2KI+xN3uW7SWCpUST7sTxollsLQba7LT8IzU9rNwzc2ZGo
QS7H38NFEzBY+Bg3XDKI0iJkCaEdsjhnFTlljc/qkBxYKwpb6MYNWjvOaEtG/I+j42xWQhGauLVm
OSf0E8zLdGIPIavhXBtKfJWsEI48A122zaqEa/P0SutWNLIHLrxDqUB21syF/irg+I5mTJqOcjkC
sJm3w88sRsgjAydCal+dEP57NMxf4Nw2qAeJ7iTI3XYApV8TzZ/ndxBQqdeoIfj/8hTKPW8Ytf+Z
8MsMhHbDchezjDMA0qVmXgssZsx2ERpkMrrjtsG5cYli/6qxG9S3RZftVflodHW9MwQuBOBvefxD
2rg7+iruAIhb67Gbb+SA19tr5Sk4eypi87TzpQaPQmi3zaJq6HJLuQvepl9aRYcoJ0M6Y6pU5o04
YWhZkYmpuURhVoruvUoin96Aj6cStR+mH6mM1sno5siEK0CdQ4kbXfYprIkfO7xJH7JELm4tHznp
lb3Cb5SBKjg+SPf8WRqgXUB7W8hArWjICSICLDhjMR3SN28AAH5tJieiAg1DzL6UwCrytdiMU7KG
gZ6D7kNu1otIcI/1tTdQTfnefE7EZInIZs/Een+YbiNuZeZDpMUb1+fW6OcJVZuUN3POqK6/a9sJ
y2jSFZi1Hg+jEg9+ZDDYK36cS6j7ZGquOWiDFkQzbqdRw7SVpanDDqSCIl9jvWCEfpnBBlVjV0df
zOalFcKH1u8sRtD9gUPPUOOngEohRkEoeVTP0IBKFdU95KNGE1ZJiGuJq41llJhEXLFCzHqhWs4k
c1go6rBRPxAuZmF726xpG2yavBTvpRc4WxZtgFO3UiyuNKuLaVdUPX2uf0VL0YVSOwndaUAnREvm
jjT8yksSq1yAFX4WFZ1fqvBXBPTyScEBOn5BQhrSPLPiJujniMkDJ8rO0zFjorJ8L6eX61bpLzp6
+0wc9KOM3IYZkVniX8r/Qqlj44tS1mQ+AipPbGjrzm6XV1Sa76IpwdbiAp5+C13+yNh/D8v1y8mq
CWReOJ8OFgu4HdK96+xdA0AjnJEM2rKay6xkWIiI8Q8U+9VxdyWDIvOpozbVTtnxZ5ii13aT/4fz
yITybcjZPvnk3nyC+0ibUx1U5HduqMqdRceUjYqggl3vPgyp+05bS5Urb91V1dpoxFDq8Pw/JqXv
XkbSBgsPOgb8XL8HhiR6UIHY+IZks31s6DXRkq4w1rDhzKsZ/O3fphuchf2pWdF4/PzLvZ+pA3y/
rUEBtt9rbbcjSpC85G6iVS+X8tnK8zYw8cpWlgyNT1NX9CWJUIQpNLo4wR2DHuA/Fa8UK88oHb6z
Bj0h1459v+l+RIaWpLDb2Zu6ZeAoNAp5kyJr9F2QpIz3qxckgiNJvJpt4R7hgTagfksNG+3p+aO0
bhIatc6o5qdZ3wvNwXb9ACoIehBTrm7gMafJfVcMmT4IBpab+Mo77uGXFOm/xr0b8A57Iu/hNOia
RC/VFneWCpXam9KClqvWcSG+sxeGoOaBAVNo/qLEcDtTS+u5kkCTyVgK9i0g67FL38m7g+hvifnT
13ahsXlvvOWg1s2nRcSclmlIJbiEChfERC8Vps0t5vcwKpFSTbUMQORwyO+ItYWOuVRR/xXXxeuX
tGiJcUFzp3qwFQTE2r9W/4LV/4voOKLYIplavByBoFXeLHje8/x/HHkDNRY9I/IMoVR6nXbJw9Iq
o6gvBcsS4eR7Qkagp3SNERoM90UghcHCMOUih0SjVGE7cmvs7xDOyy+jjFLhj5Nf4HdyFs1fv+ZB
Rlwx2uuq1DyFFosimR3uD/4VndrjDCMZfyyn5M6O+IyXcruo4mx46nW7oI3Sqv/w81I8LC2n9uE9
AEu1PhCZ9wCIW26p7Vbye3KrvIkZk4mg2vAPqud+RExhCgTMCkWydegtZG6NaRy1yNc859q/KyZA
O2k64vLNM+1JmGBl04EoqA4/iqAS9rvqE+2Q9Ny/Hzkfabxi2n1HIpciEA7yOWw3yTZVI3p9yg/s
0UzQZGk20B51C6aFlAfRku9rjuoN10mWpsXkVs50fKgYTWHsxlL77b0B07u4mWUDMvpwsbT0vYe2
NWd+LscgFYpNu3nZaoFQDBW63Y30TT68cc9DwZT8o8qwqt9DfQMRDX0wYtBAh3MFP64EUIPhdVWD
eaeWhUOQgf13leT46Qbipq2C4bVNQecdkRR/3nqlQeFPyB+3sRvTwlzDVLC4jeWrsjxeWBiol4N4
bLeVR9X7FFOYDbult8AI6URulhzZpPA/nHTcfTOOo0sgt6N1hihC+0sdw+Q/+/N+ESEb9wys3EU9
8q4WEg55hGhTw4JMKkC2CAD+XdXAgr+CB9B2RmXuQ8NO5EKHwESqp5I5nRFVgYCPXd7k7+0rQfVJ
lMl9u0qnUYl8gsZDEu0bKvg7GFBG6p4AfAK5EkOex0c2g8Ji6wPnbX1ezLegZ0T0o8eTWAd7Txhe
Cpb/CQfKikZq+imv1uv4kDzsWzdXqot/3FStmmgrdH4O586t8CDP86vCOSIuM2zt1AOmz2wvv/XS
GuAXQ7Fq+pRuAHiXXjuvMsPYmGr2UGdtsqFOK07ZXKaKzcuvQ/dMgHQ8s9esvK3syQCTjx8gTXAQ
e5XrkqLxi/I8KNdTjf0H0nyaD5swJ9L3wvCqeLhd3lZH6diegTIKeioN2MUQ8cu2BKfgiVIg0AOM
K1H3rVL+j6MQWYQ/H2PAQI0YW9z1dTrKgG+16wG8HjSXus+TJXSk5exIqWFDPKohFzmo6XWPxcKn
jgcxpkMC9xyDn6RRH/qPVsUDLm+KpYXENo6ErbvhDJRjXrgqJW7a8envej73eSxDFaGwViFFUw+t
/Om7aFoQvsB9jSbcnP1NRO0LrX+lI0T9hEpbmG2PU8Dx7MvXnyMHVQslboWf4klAZhCBgR5o0dfw
POB2N+p2aGMEalpQ5CDdHPIBH5W5SPnO54yNu4oE6URkvhiL2p3y2BzFCitOPvCOlL5eF/FvsWSU
ta8Vph4fQDH+uBl106ZDSv5H5vzuq85oyxcLVcfLVgtuZ/YelGhU59j9CTFk8c1ZGdbiufnXNiaX
83OEwc/l0XhOOmIU0wBxSJMJaW2qLe/WuMwiD7g8z17OyIuMuDrDc2WCgXQa3GauoBBye+4uodp2
h5lq4+6pT7Sm2rNzA38ekVaxsg0u0GhAGsCKU5enZMMNKkVg+FU4FkZRkte4kceKAWZMFmMALLVR
TuMc51d+eIKCbhy2i7iqsJvZH6KGYG2SWwMDKkoA9GlS+yw13USik9kVjp8KNZ+flT8LFNCB3ruW
2dsdL5OHXfdK8j7q2iQOsiUX3UmErsD9TbVCY+WIqHl8yaZfFIUGM1aQvYBICE6bqMBBB6dxWOXY
30Bbos0j5+Vw3WR4xzwyD8ed0Yj3A8f6t6Jd0fUIC8Fr0GHXPZJr9vHnRtLZGsneDLI9RjZ1HngF
gztxSKlCScL1j5AkHadWl1hhoaflI6xnra2qZY/nzCnPeKf58AaYqTkgxsQnTfJRE7/+cC+m2KKb
qzucTSw/wW7qo4iuVPjHwLeW5AOhpRYXhzodSlyx8rJxgar2w55Qr3eJlCN1NBzhtpOmhQmmLK2d
2ilg+ejwB3w3b6HEvdoNTQBvhy4zvUxUzq1X8b0Rt5zkRm1b+C0qvzZy41QhMfzbkf1q0PXrWxXV
xJHsFAGqMJgvjoVXJIAXy0nIPyyx2t5CSuBOdkILmQtOgP3Eb4186Qg2SVlczsMyN9Ophnr/5A3c
TCJS7ZM3HemE1EQXN34m0gmlvkIaysu/21e1UgAKbPa5xOr7aixLWg7+7yZE8mwXUySWaEVEv+PS
KR9y3E0P9v/XfEvS6MK4bRGNUW1CowPO6BBmZ8OqccWTE9KMtnXi4f+Bw/EObjY8YMA2XvnT6yww
M5OUfpQ9jaYJo9tioTvZgwzSqqhXLkXnuokmicM+ts6TE7mTjQ+W2RJWLJ7G2gDR/qQVSTfhPRWe
sgVdOkMCSaqgFatuS/iAugbWQ7I+cqoxalBUeGmcniqjkt70tRBW6MaBAkr++53aAu2p+x/oKTxc
H5DJE/7c17ZqeDbTEtEYGlNjkX5sXTNbm+WBEeW8B+KXnGGbVyeHafnmQGLOwAeEA2Od56zSIkB4
9sk1S1AxZQGvr4+n6+zM7k1d95kVO77Cfe09ouKtU9Y9ztSEMJsRdhm7hx5mkjXL2W/DKqEAc2BQ
/pDCvefTAXMFnq0Ij9ouPyXeuTCrcviA3EBAK118QzyN0uP9lJY+VVISEH0n8wTCyeAYxv0LPiMN
Ugt7U29pBFGZGDH2ZgVbmaNI/0uEmJAWjUKhjT6gv3YWTP4zQ3v/c7+6OiAFJDNR906heyY+J6jL
wXgrPCVyHG43HVacvlDxVbm7ZaTiN6fh7HMIewy/7IACW6H4A3MjszHO45Rl3gjgxy2USxExGdMd
1/K8D/nS6NzqQ9aP5N8tHfHSiqA4QAQsrrcDAXYCvc4sZuE9lhOBSGR+0pj2v7HMvfIPsxzOXSzy
d3AqhpLpnjuWHAKHRM4FwG2gf4rjHKTtALN3wyLrx/pnyD6t2r4E/ekisTB7Mvy5PagH2i7121TK
D8WJo37ZBPvZq4yw2g1jAAO6R3tYU1cEIQ1Qlv8RtScxed0kXYXybSi0NsSwZQKTMFUoW2tNE8Sd
XvqB0T1DozblCsWZlzDTpiQm5Iec8zyIsJnLyMMEitmLGogp4OSsLPcIBivHreO9h2owneZoX82y
g4AyI0i4QQ2CncI3VhwDHQd8pxcZvwqFbZN1ucQplSvZchDXSGjb62JNsOJWK8EEjVlDdNH3+fIa
D0uRpyyVC/SaiyIz0J/E+I/yTkaYVuklD497XCRQC6F8L82dQvDs/Jsv2+KJevDBbuwzv2JT2Tp3
uHD2nz3+jfDwMd0qZ+l4s5/Z20jPsCV76YOG/R+qUGVITJhbnMJvFG+/sWscf92SjCAswtuy1OPC
G587/UxkfEACpgLnAkYZpuJZljXmH0eAVjRiJ4iya89VzBF2zDE52B7p3J0tYgJrYUQyVgy16512
8nTNAaub1j3NiOuBFHUb9LEB3Gz7uIAFKTOORbw/3a1rj9jjBYgyuMBtsyEmaKi7ZYGti6HeYW+j
qRugh5fLJGPgAuT/KQRHzBYnxjzULygU2fwhM/9HzkjnDHeG0OyXHFLkQkVUkN6MKZf4LyZz3/8X
bIwVhtXGrvvFHs7roUdNABAt9JUMOlHsJTsbYFi9wNBKk7h9yiLV+FhAmrJJagtKaPsgygJlzHXy
Mt/O8UxTEoCWet7ybl1ed5yLPic+srRT6DuQu9Q66/PX2D5IqPAGHeVSzYcewQo8Sso82KxQE7Qq
CBSZ7jxhjapQ3tb4LkhYPYhns6fQcCj4oXAgUGx/bXG7kaPXxzw4RngWx5Fk8gmFyVsnAJPTPLNs
tbMHjJiFGXwPZK2/yKbrMpZPwunJLzFEl0m1siOWWaOrVDYmvtf5y54GHAg86AkkPPSkhdMIQOL7
U+FgkXhr9IsAyaj2CwUaGXHpIKTNYZ5tnb14wDbhev61/fq+dcamFs327dPPoPTnEl+3Cvdv6Eni
vQJO+7ZpyWOz/CZFbb/kYEVqs3nFJuT9w1cXZjBrZs/4RjMq5RB7qWHGkU00se4eo9uAHTOcDsBp
AEVAfFCBHAQfvIdG9dtMOdw1hhpVsNTixzZICN0axsrqEm2O96k0ji0rCvlcQzgNbhk/nyuwQqjK
+Zjl0SjseBBvOD7c2yh6V1KvCNsk7E4E3UlhmM6jAc8/xwpJVo7//FF6Zl5Y2RU3OkIvj0UGPj2V
HXbzacg/WguB2lsER8l34uSspYHyMZNZ+ghb02gPIm409gkbIcCw5kH9TLSy9AXEZ9et2A0XRFZD
DOdrw37x5a9t+K37Xcecx64NX+bHGNKZtQZz8nR7nFxx5mZ7YePEWWIBT8668We/Ptl210MfY3FI
Dzxoebv+kQrc7xfggkpM3qBQaj+lVywYB7/j9ObSUAfgC5qXXI9o2xWwUix30Rnalgbgn2toJjkG
tnXBzgX/LuvmpE5oCbXM06agkrbXLNZldjKGTl2+NUN6eEnOxeUP7PrmlUR0431pzSu6WmH3JheT
ykKM5Cge7RukW817e9/ZQztPzy71X6uTvzUVaFU3WWiMXq9MkAIywBkGSOb5HHR298VqnUGhPdnP
LuSeUeEfWLf5wxCuLvizzopedxBAdV3fVAhUlccoNA0NXPvBO6R49/l8S1L/6VDMvnsyHJsyS1TU
7DDO2Ft3vWYRt6Ay1o+/qtQogghoQEkmdIEC3rXFvyOOIfhBBdJar/h2438DDXKN1Y3MxR8schl1
qk5EIboMin8c9EsRMtT7UbGA0LFN+Sz9SCnCaV9c0Oad0qVnSdAmUnRY4mra9mk6yu88kFh4MOwY
AdzifyjF0oFRtkNnXT0YhEVUrMp7w0tHSKzZuk6nU1bzZRMntbL9toAeq9gLUaBn8pJ/hHsGiEbN
J4QTxCyTWiAFfp/TlRhEOwWv/NJQ3/TZuMwt37o0y5TPDjGKjsqD6r4Quxdu6lFBvuw/OnowGOKX
QOV579sYb2uRfl6oIsgbK4KKLGNN/8Eqk76EqXIf6EZB9C9XtaJBuWZ7J/OrUldd1xmoXVj2ioAz
3yM7g11/gK8+eZWDa1mGTtiTjl5oIJpPzSiYYG/lSCmgzXXIqq+9uXBz5UvYpNTNeWounwTv8u6j
Nb2mqzLhBG1RtJ2hVQNP6No/Bi5/MpWpoONmGEKgehegVC6AR3WQHOifb4C/4bapGcaD074i6b77
K1udltlDc4O18zw9yEAl01OnLX7SvsoiAFxvWQdBi6s2Zw7AkxXlTBxiIzqI8f9Pz/nOx2HHGWCd
8kdHviyLtqlNj/hvzpLCuMLl7QBbzNLpesTXvlJbL8hnU3jzkw23XjOOtKAIqIR0rb+16IAizoV/
+jplhbJXjNvBK1NeoiVJi4Ip5nKi46E3It5kNwzxpgoepqahHyMGgANNJdEucKvh7CbX/iPN8brO
trkQqPawdHDHVhvsaEgmjC2y9UjzAzKrwve1jzqc+YeF072t0RQJbMz6BqEOlD22mo72PKl88LtE
HVf9xWPeW2WRfjtICVxkH6HthFuXNIbDeK7x2KWx1BbdzW1EVPxRwWOvpRpFDoVzp3CgydC3pW2j
PmnyoRvXaQtqeeNMcsBALhdkfKE85dc8UznRdM7iHHn53XvoKn+Kac1G1msO5AmnONhOsZIdFjW7
uVfISg8R/JiZTr+PAYi4+ErfAhLhJ5AiZa0nl21qcM2rsHO8yP1u1D/MYPtwqqV203Eputiz/DKX
+jqjLB4fquMGkWA5gDMmE383IAiOe3EJaghCTq025YQ0+xbg22ff2Olxpx2hk3ocr/C1+WpyVKS7
2szke8Dp9J4SscLIWYM963/Dzr3eimRjwmXhOM3ISWmycOhEz3MqCrk4DvrHP5eRpoZrJ7+9s5+1
0GZqz5GIfnt9eNHhfzkA8fHr8bMTUN1ydy49U0LkPjD1rf6Puwlwt/HlBHzebjuS2aatildKnN3t
PaJ6wrI0iyi4rlWwIQpyN2+K26cSrXrn0s60PH2MMBArPyjrLCvkhamf/LPN/+tYkA3HEVImEXz8
Nst1S+B7OFYuIUKOF+91mpd6qsNQZ2KmorKvxKzPIh8XgVpY1pygQC+xCGB7Ig200M5KrWAmhOie
veuZKjgfkjGTBTYVlOUFLP5mtOl0i8nF9ubmVpVRdwV8wXaDrLZB1EEsxpMMZAHQ/s6yhhp+OYmt
hmjK9ZQdoZAlsFNod7f+mt9LUCb/T7lsB+jtYyHqX2B2MLFgfvxyIP1h2G1dipj7u21BHJiGSVov
EzosmJ8YJy7yINdfMagT8ryvC96lnnvHfUJn3S/Bb6NEjST01PbMLC4ndrMl6iZkDgR2lOV7lUAu
goiQ3tiCDgx0kK0F+M5L8S36dcBd0x/tJ6tsV5BviSZ3mjdEhLjJzvjdfh0ViIWWd18Ih3NJ1DOZ
fvyt+4l7aFkhKX9ArGrUfDnywXd9rCh/RZtbSAeZTWcbPMNasibnLYfSo8SpAYaYkRRx6Mmu3ORi
8/XuK1cZDv06udUOHij9oLfO/1DRpVcAw+2XDqRcQlziPwsZtzgBVYXiyx6Ohbp/Miz8OReE3BDt
xBobF300Uh6pmzp1M+9z3SUgeRWJe4azaq33kxkqCI7RYGLgjAO8ATBRcbdeQfDLCygQOEyZV+sq
KhYUuM2Q3lNv6sJ0k1ETvPnGxoBpk03iRq8hQkZdHFuFaGEbuf0M/WIOV99K4dDTjYCnKOKxCWs3
yVc226PvxPhL4G1P8LeliCuYU1dW9Q/2xumV/my0Wf2LtNmVnwvjvXWwviWAUtzKhFHN83BW2PyH
RXue58NE/7K4Ic+ObQ7w2uXVo6VQvL3HlX6Zu6o5EzlD4p9i/+nzBqs2z8rQf609ll8+sJNhGFA5
BavpQ9tnYgJ2aaL2qL8mLa43MnfR5AYzVZ3kxoQPA7lVhJ4W45AB/GCvcGMLf92Wqd1iVd1D3AhT
f9c4miIzQXhLGnwGO/vd4efV8PA9U1WjIfVpdBB4MD20hSOcC4qwdW6+EeLtlrD+sREmtMz6XgxD
mFtMbcVewFq2TOSGZhyRKhDgzM5OD8xVMH1o6kduNlCNgoDiyQVQ9HuhMsTpd6bfxutjGxT+B+PB
B5GhELPPcPReYBwETsiYgoeo8kPvIOhz+O5PUV2h82a1I8B6OyUVfsoJDIrEOv1BKo36Hoe0ckYg
lIP/ENqrf2LbYIkTqo5VRedCjpyQ5MYbBRd13WYrdWoWdl3CU7uxoWtn2zZSocyrwmqvfS57TggC
E/Bl417/LgpFG11XXZx4dh3EqexUKOp5AJbXYcXXg3GSXfP+2X4HQyY+w5cSbKRCX0r6FkPA2ERa
Np/zuRMKiIv6LJcFipSqOAjsDksXXj/iRpHk8nQYhVSzFm2a8x76RDIwbRalsyIScKU8DQN4I2v+
2EiBK9zEj5U9gsXq1sG4CEwjjiOqWvHEMjfbt7omv+nA2X/Qini4ey6fLToBXm+r1FFoyq/PBnop
NLJhFajHLLhxDZPk0BEi/A+/o8oQKiFa+7cVdFA9DxbVqaQjoanYu9GpOXWJTmKhqnr1H1HL01dJ
REPpRpbTlM1xst9RpgabTSMOMmAMl925Afy3bfvWi9RW9YDErBA5ZBnkgYkX/UVlVVACsOcTv8kB
Fvu9p3dH+zF7bf6WeYXnWqb0dtB08O6CbPZ/R3aipkuJ/VzWjJgjbW/rYgvO30wmrGbB9tgIXTQ1
Lfvty+J2yaYB6LbwFAI+ikv0fhZmRgKHs8PRSL1c0iH4JUb+bvwJz0qOY9IAi3wSeXW5XF8vOpWY
zzIaCeHbIg7MNEnS0Q3VbtSSSxL5J4hue1XdnfKNpYnYWbLxVo11oHJqEROGZYgtPDHWur4G8l6V
WkLG8O4fnskC/hzUloY76BLI7F4ASFJlJN6b0g/Rs1rTVPQenr+a+iiuvXF15KjSg5yzRdxLKc2h
Qj5l2LEn+7DOYYDZsZ2FUeXma5j6RoSGmczdmHLI2vd0W2XmLSQxyz1u0LTykwFi9M91bsbIdOcq
Al8+Ht/YJZakpvI1DAfKcaaOh46l8QoDsp2e6A8dTFaQC2/kmgiH8nbjdLzpHbRJPxTtlHYsKDWT
YwbtdNCxLO5T/H8qsiPF+xrHQezLcCutL8paXsX5x8aqIsEfIk1Tvs0Imgy6l9Nf7zBUWueSc+U8
lHBIP9xMwZ9UIAL06GCxvgP+yp7YNENKJF0hE8dD5tJVLQJCdQd4CfnzOdRCwD8h1UgEHqR+h0Yp
3h54P4mrtOPehW3zVrR6VlFrejxvbUyy2fyqpoi3EqHbZobK/9hqfMp06QHtNcI3L+Wr5m0pxOtR
W/nkqPd6SbW5ZbLwtncy8KAZjXyVFru48r8ZCnZbXf2Fiyaz9lNCWOz9dI8WWv0lFZ7H/2OYU6OA
kFFWgoMTY3QIri3l50xfrqIDnarAmCb9famG/BLKvM3MiDFjcG1ex5annSGIYcTPND0DcbiHE8yX
OzOjNHxCdsDTARijXzfvf2F2SfWqYrCd+nkFaihrSGWyjA5IyJ+05kZIqH6ApppvD8/WzSCGjGMl
QDgkf/iI+pFH0bob9PIngfuMjVwonsVHYsxGVLO44XS1R3BrxCXHNzR/Hx/ko5UFOeyy5F7lE8Jz
AfCIoJLEMWr6+GiQduEA55wtQIOA99N4OeFcbJRxYV/ynIwCavzvDEgETJFdDRvT9kZWUQyVM1EX
rfYUnUNmMMjAHhCfyxZo7hVbSZhPFmMapiaAyWJe0jh6rxVnU1xhaEaAXomtzLsvduKR4qyG/CU+
x8c1EGKxTOfwbVstzpu+p4PP96xqfOPZ8TbHAST3Jl+alaxn5V/KcQfgOguTlv/WGzE8e573en38
riRZbsfBjBTh+TJGFP9aLijTQuxrNZPtPjE/xxmpnjw4MR17cfDTv6xFeIpjAUPwPq6VV7surav3
Ydjzha7THsQN+1ZB35nGPudQDrH26d9kpSvNqCqHlFthtyAqlsGYogG7E0jfYPgaWxT8gFFfdvhi
1u8YrhOhWOHk6E00hg9xdcJ7qHVz/d8abP6JgcehE/2bzYGaOOOkNFK75AoG+Hy+TvYjrl6NWz3B
BHzc+Yic4xUbprvWYumwKxEcnLW5BgdgeGe1zq7XokatDpumyP/6K4+atOLrtLz7LGk/3Z7hv3Rg
/mmaDo8RKc+rJzV8bj6dqzMsEnrNhbiyx+kR/H3/oF+bWgCBMznMQ+mXGreFTeBQlqzVT4ADaUri
IskJ52bE17IaVH/wqout9RVCER7laHGbknvzOEyL0E1+vzV1c7wvKZ52z6xGKDofa6NF2fZ+486f
y90gRaS5Lx9iUtJTAvwjIEzgVPb+3kx1g2YUdyexR2UsW9E7IzX5Fn0PHvLbgbyeACbm+dsDGQea
r1XOkZGR7GmMtb2F0B9495NGqiroj+csEJoe7vP1MEWLSkHNkmteKkokbUljwo4ZIgn3n6XBp/y8
ob4Xrk05YkrOc0eNC9683Y3Hf2nyXiGuMUcVAa7QWYwEz0+6plNOg7zBByxJBMGTyTWEAs2Ghr8D
XkjpJbTQWNrywYB07Xm9k69iOzdnmHDa46s9UkoyBWHGyrMQJYGBbqHGdm0w7sNgtpZPaOqAjXNm
qTaeOepMW+tRCR4ywvgjJfJlwV840HXc8xdoBcypVu4uNm/UrMRhISn/BEzF8qCSUY1hHw457RjX
ZUxMi5TGqqHZh29QpYC2y8oHS385h/vAdA340I4i9ipWAf9YEHAd5XZUEjisNOqyTMVLCFdAHlCe
HtIRXQAZmNLfaOekGsoYks77zKRW/OHNHQNgq07gA3kGDIqM48evbBLMsJSKRRrzRaCG4/ouEO2U
rLkLzmqPc9zWxfmmyVsUNQAeeVcka1b3c5sTkzg/x/YZlRf+xvYYdw/qim9DnsFdgWoZimPaPlbA
mkx0/mFmZNQqD9bmm/8wd2s4BXbhWB+SfBzzyhLjYDoMhMGE1W7dkAGkd0FblXYj91sfEE7uTWoT
H7hisj06Dd1i0aUo/K/ssU/4KWHHmq6OtyWZ9Bp81Pl+0w/pAcX7D4q292X/689S63ioRc3vp+66
AnQGyZDy0JReA8LTQ4A9/ttr2qQI9O56bmD5zQGhKuRMe/A33gae0G280ZNw0X9kLF8NT8Wdtled
VxkWVMmlpcqIOut9XqWdfnLRcSAMOfFmtdwEqoh07LsjVJkar4ugD1EZMTDNE+0iGZhygdVC21lJ
PtRQSJZjzYNvGVOX69o6caWzAZs78EVM6CJodTiT3xnrI/SlVIw6FFYBqpDYR4ZMdc3fJODGuLeN
KLzn6RjDQQky9mW4IPsaBPneVcDPf1gftQ8ddpcjnUmUSM21F5swlN7gKDefKZq0LlsENA/NeAcV
GYroH2HKEN5cvZ8/8bsTEyxAFxWg+Q4hdV+sJyuX4JQY0yy0cHKuDofkM5pnINWUpb9f1VQToqbA
jQS6l0+bxi9xCvEr600xB3/W3JxvJLg86Omj4p0l/cLUC0HM5Hr/EyuviAaQDWzx22VEKzuJq74i
Y1U48SNR57tKobIX3jepnmejeVy0el0bK+82xCkPcZhSB6x6bSDNaw1dkEJSlO5lzSOTDmDi0mu9
BLXiEbJtUROgFuAy6hozdfFaeVNIO7ne3+vmdfeRwnCZDwRQmY9XlKZtQzrxBbppfvO6UOLvd5jK
nMDN78as3P9hU+ngefqVbJhdVEhS6ChhIXigjfyeHVx3e982c6mreB6DQRnrOaybTTfUC8LE2WrP
acxSB23N+alZLA5+kcL1Tl3jBic8AzMOD0bIcsZoCbvh6XSYYFWx2nWb5ai5wfrBqdnBnxWBzG1b
TyhFSv0nbdJJ8xGzuNWyWN4c8v6RjLDs3eCiRiI7WyPM2pHGdmLE3NkoF3WhfVjiV0epU/vTGSI9
0MunlD7hH22nWlBt7xHHvrmdA34EC2G9aFyKQXTKj4szkP7z4IkRNTCNpe6Ul4EFxehAvchJw5Ym
k0P6xoFyH94lIFzRnzpUm4wBfCIviST+TX15GcEnUyI6GieexI29xi5L33SA5qzcQhNP4MWsQL++
a+Z/mqYEkRJOWBbPpbYn2qcGkcUb1JTQDNYva0v8EFloLH0+QhOsHbW7El/9bCVqqwBfx1Qxd8Ek
Zul+gIg075unyu6WZkVqF00Rpyktl0KxCDPhkcMIFJ3uPPC6HqI6U4+XX6fLZg+CE1+bH5ZVoDNe
PDnkTeIrHF4MO3Pfwvxvla0AY6w/XtpW3qGu9y19JSZLzs9fz+XVDau36xPGVKirB31JZPRfg91y
9vRlRvkco5O7Jz2Wu8T/6W0m4vJAd0eT57O/cN84/p6npJzScx6wnwLX1mmkX1ptNGtjiCF+M2/3
BkfimH95fSEIAmmzOIbaMnCmXTxmlf3VMm47rkEI76wIEmNekNPRejyql0eLZl1ffN4FWhjXXmiI
Rr4mMYUjmzL8q3H6lbNO2FyXhETZTJcVnCXj4pJ5uw3vYPXuvxCMuYAnr4kmAYvZn+CYHClQZAiS
/3nroEFBpTARlBNNo1+FXGo3utuorUHFEcUDdnUFzg7hq7bd707T0wWqlKHUW3XIzukMQe/TjlWb
WQBCkJJmZMtVTydvKuhcZMZf6n2WN2zf3ndA7Ob2Nsjnk1CERwLKNeoDyx8tNJqZNccXVVDS6Yt1
snB/pOZsZSBnKMlE8uArpLibP7W+bqCEXTPWveHUcVLIjJe2EfWLJ4YoYDUgpEcTpZIjp/aT6kV1
qA/RkyykZMEiPQAmP3POM25JcLfN0vVMevxY3dT+vcDwa/o93jw8Ex0SQtS8u6nd1CRrEQsuztgK
/n540CBoeBtkzb895djczx45YbetYGx3OGRae/wNj8fCgY9OvQkUCD/dRv7Z4WRfhEbGu9Ay9T0j
zq2Iu2uxM+bOQ/lZHEEgYIUC2XBj88c/cSsJ/bsazLk6mL4tk7bi3+LBO0X2k9L2xTbBQVrC+t3R
zVqdtLf6q7w1EwvKoEN8hWl819XedTE4YrhY+1/kcYXhcz82bASXuk8V0E1ko7aiW6UkduWB5xNQ
tS3yumIoCevho8XAtX/2lmpqbWCizyoY7NbJ/ZSAWamFKDFv1f21yme4KdCpsdx3bhnKYxpbJWbs
6cr6XzuPhl8JeAyBNBoR/0X3yrrCGSES+a5Y82+Dqt3PYpaEDQ9sZfhW0ZTC3s0Qx0v1ffGq5jC/
P8uI0aRH1zvAjrsWnS4Sf8yj4ni1v8bE8wa0CA7Q0H2eyPAUqVQ9FV7hKJX7HBBS07DDJajGZH9c
6uJeGoISY9Gj/LFixCBSc8r1uauBtxavicmuoXvJ68BErI4bNiXKyPjrQEzgHJKjrs7yQGiA74Ic
GZOe4u1vfXs5R1lRKh9ff97v1eJxmzmDhZ5vnDqI32HgNbXO+/fqPlzekJY1kUKo8Bd4gfXHGNJ7
upORNUlZbjymH054e8jNgHtXkVx9s4cu7rAI9+PrpakIVFUDMd8uQN2g8WnxrRRpCgiCTE29MgnW
9YEivfwJ1r2VPszKS/gcE6e4MyGrtmxgF6P981ChA+K3zcaJm9vTspvpI3eW1NrKNbrxRCWsRmde
h8UgZtjNce/7QFD6OciwZ8Lty+iarysQhaWr/viGhx9DM61sx4nIuWQhih0FpE2jl/VC0hsU7d13
SoJWMZoQUO7hgTQaODNn7UFJcBcgSBpTQpNqneYZ7zUyM1CwNm2gYN7KvOLz/RTJYPFmO8BBKOX3
jtdqCMULctoj7ebqCmrJDPTCmtp8EjUfIo0fb3UEovD1igz90sFTrjXgOeEf7zFGsWxTccePzqYw
Btndtq1VL4F5fZwvI8Z2G9FdvEmz8Hc9yg4QWw59JRfK6kk9C6c2zc4jSHM4NoQXPLjn3XjgG+Wq
rBGguxvZ+d8Y0VxLkefa/261Hg06Rcrt+BQ5Zj3flEyPYY35WFo7yMGp8ztzEXAqy/mMeJernw4w
+a1PfFM5HCieAUp1ZjrOKBO7lVAKsCoW+0XPHB54xsF+xYub+pqsJHeCmLj7itz+6MXn1ahTqS5M
e6idrwMkiJWa0SXnwkguX6XG+7oQKiQczhyT3hNYDA8WNt0FJrSAeAGxA0dzfvY4U2ub0DIxztY0
iA4ntcR1/RoUbylGmm6qr64hMDWBwwmHXeQoahhVd6aE6uW8MqMnl/ZeDqbtwcklnp+HT7l3/bZj
dZtg3Qw29XGdoNXd2Nva/AHYhtOpm0b4XVHYD9k40l/wrumecZLT9JLaqw0vw6Mdqdl1n0okzyLI
TQTfqfY8aVn1kFeEa/mDuKLsqKDPX4ZlDjLqkjb5rXs1vXZRT+yIm2m5ZZEgDfYZaWZoaTyw0kOc
76juscBHpzuoMmJ8nciiTihI/ebklTyNBE8hRfSi0qQHgniC3eHa6UWuDklRYCLYC2YoJOdYGwiJ
WbCHsFHxg0MPzIz5mswos+28KiC/upU7SIPHrQM/QnFwvJCYM5aEa6sg9ShpZD8KrMZZHSOjrVkU
++Oth8xWk6thRF4a9oTwjSmK6CLoqXFqKFklPFJ10PMIthWFhjljon+nt/b2qJRFtBcKoKhhswBI
Sg5vxJR6BqkZEMk9vJF7kjms6L8+Ok31CDtq0cupPd24ztjQcim8ANoLX9V7LoKImXYg4r/MuUwI
g30hMwwWm01BZscB+hVbFm9C27oz0o8NtzDogHTQT+DzqaCbN0oEc1vezX6cZj4BFdsdPV97Jmk3
nf5fPqvKfGHA2+DVBJ+ybtSBIr5RV94NzS55hOLcjVA8+QxX5UFXNw89D83WzPMe2MvrUDichGOW
skm/MPnfZrAxOY1wYV5kUg4u+6q2z4ExAnxTL4TCCzfBsEc31ftVWseFUWUbJ4Mvpt6s1z93BMHR
f4tvJB95nl+Xmi69uFhCV5Fsfi20HKVKQWRY+e9zL2jsB+JMtLCH6LAO4171hDtlSKatDxRXAd+S
dNPeCobbEQa4wjbYsKyLZxM10u9ZSDkGeuesw1aGwOF2Q6b4ZdwLEuGWlCgv79OqWxM6aNAJ72tU
6x+fGs9/CN4+Yp90m0Glf5ca/0HALFhZoYuL17PaALiil1LYwODHe88ZkfZJ+eFmoajpaaRBNDcj
dAyhOqkdCmCr8wssxKFsiR6JdCfMdo6RaV3bbn55wq+7UHYhdx7tXB7ghsdyy4TIRpxTl9Ij85Pl
x91JlLpseSRqrv4sa48iyJ947VJ4XpvOoeSYYkjc0nULq3OqsCWpR7Coxe5xLLD5Ck7xSvJLR68y
dVLznv2MWVrMO5B8E0ObWfMP3rPJ/61Xr+ugA+eNMB04/m+uWJoauxr9GElbmOuYPFnKbheB+wP7
R/3veBQ3RirQgX61afjLD1pxtWK57+esDLGIDc+DvwykYFJ1wO6VkdGwP08Nc/03MOSCZLKU9VWs
05gW3aBasTCCzzaCsayqg/AoppkX0h7/x+D8k/XXN+RDM/GUBOFW7AATyqeYweWKGqTUapaKP02k
WxNG8s/BMI5o24gpAnIkG1HEG8hjSh7+OqGWYYfxrhHz9+fMGm4Dymu0ttJk1oiC9aiJoy4RDsL7
xL0TClgAj5HiaOqnYPXa2DpPyeNa5bvHCEZKxtabFvTK12mS7avf0UAiEOhSL37ceLHKepk1qGdQ
yUYWhTdYFiB29LrjAQxMUvOFHYIS8vLqPw7gr+7kaj6U7BiX4O+GPglyC/J/FXzI6IFAPGf91u17
1Gh/Ms1JwrpgsoGz4HR2I33To2l4yL5A8s/kw4zLHgyCDlVNzGPnA6IztbWDizoAU3IQgHHxxtKq
WH80JenK1dzesu4W6RwJ7b7BTRnAI6M7OcyhHkcZilqYFyJ87TSBotDfvkE6UZVNZalSGZPUsbQf
9dff1howxM25qM4g+q7zwZlgm02odzlc9eYD+ANeW6mlToRp1jpY5P04viNatAJ/U33EP5sEl87h
Gn3WfdNoWOAsnp3nTyb4tC655kKln3pGQuuqPRfXyqMP5dC0gWEwH8uevmG6gC6K9XRljsr+8Nlu
2nsnJr8tqPQ1+LBmdO3NOlrXlgnFn5VlpeoOJdb+SmEHm5beI6o+9KIrbKGDA+h4CG5nHBOfQJRF
moihZ4ultd3vlIc2hMFIfOZ2wsrI7DnmqYD6EHK2emkXpUdMVTN9AGq+VMugC1wVLE7nczolACRu
k8iXoZBwdW0fd/r3z5O0fw0XQWXo9v04IXaPaajm5E4VPEbas4lac5lqUSeAA9ODZvbbfab2/9rR
XYrDOlZSCbkc/fDiHW5wv8ONPPd7qd94//lwA1uszuvex/SbXHXf4YoVFn1ioNJNmn/x6l8EBp1e
pkxaDsA8i6paaRrgTZTcW+icK1+xXn8lfyuqovyqsFwgfW5roBlBZDaktoeUResqUGqc7Y6zfoM3
Xwrcw+6VNFoXkd1Gnix6fMs6TQrTa4V+1+AGOVoNkkQjA/bFUEf0wDe7/b1zmZkpf5h35K2JMAWS
Qvwb2XT40CCHE7mZj+iQ5hUMlzToVJ48bwskmw2qdpuSpNp26a7BAhDoULcQisWY2v0jwaZg87yj
aotpEuhP0AL2uhPQZOPMwSZ9coccEaJhPD0+P5fZ0S8OaExe9lYbWUwIKO/iX/9sok5AAyMUwcXZ
xnxMlobF3itgoRk/9k7+XjiIsMiKG2/FVw6/mfUd7IjoLCrdIaHNuHSRLBP9wTGJCrsaoUOWMCzM
zxY0oWer7NNRx9hTuFcjhXmlVqq7KHNv8YO9YpXcfAsyPB7jZRri28h9J+BxkkZQZ0G4j1vYju/z
bok1tvrpGtURBbDsM+20ZcZXYWxSGUMFXCBwr5b+Cf1ygcW8VYrwLfuzNFho6NIVBUeQs51amVu6
r7JfJVoJdLSKGAuOrCzBE7rRJyd17v/J3g8lyHdsEWOXkr//B9MUk/IdDJVyEKHcKwKG0gxUwKML
8XoI6ojCmH7bXtUHUd5a2/aZOQOLTv5HljZUQFSZX+THQp4f/uo7pCH2qktD0zy/p2gW5m+oePnQ
u+LhqzfRaPA95TqThiSssgy+4KBNME8/kEdkTVEfMmqxAbjXjKPMIFvD48dD3IvXWeplYHZ5sNGr
+Un/NO/w6j9ObUwk+x3MfPoRRHD9hGZj32j90iJlqEMR0xx5IsMuhg5wCuSuvgjyDl+fE9FuRih+
cAgmarsyyH5er/YOoVhkjvzvWWJoA6B4byHvynh5LBYRWH6Rar57eUAxQYmoERl3H1xUtj4Qnd1X
jikz3X6T5a0tPg57VLfswL5fRHyfveBmW2Db2Rq4rebKsuEdueaeNYU83GwR5YaVG8Wv9LFbRcWT
Didowb/n4OVeY6SIYfGhvVKtlju3H/kDti0OPyBiRlvRFvDbViLzvZhYEPHKVmGq67CTymRORJBw
7QgTYFBoCxoiwmKFogtsgrYG344HO8GUgwcykLgpGLw6P/PRbjmlHcV50AGFBOmN5YzWv0qjxG7n
bRp2I69AcaXKK7xFmlNfVnRKAXAgHCJwV2nIKxrjuz18/IQX8hHfHnBkCkCTYW+BQsDbiqF73ATe
X63wajfz+F2vdvpmsHsbMT9SDTWcT/XiPV2pJIxgUXwotG0tOXbZ0nPntbb4nO99eqNI3cv9YxzI
ivZclvFzewTdsXakShvCUd+mtobuyj05aeVj5ziw0vUm7ZWeVjbaEOdPaU7xiLLNBZW5eLrz/yxF
3F7YtxHWP2uuKiVLcIJmM1hhTZWIPZSqjHv/9YLxzjsQWPhMY60ukVXiPbcXgaUgDmCQ8t7dAzYL
cDO+QmhJ+6UwS4XEsSXRow/wK9o6Fj7gfDY50J6SPVFtFGxIgPdtB0eZWau5AAxJs0fOn9MXDmUj
jppqivra/1V4sqcpqQ78yMQ+bmTrWDVQdxWjc+LcuAEWQqyO7p59mhy1id0xCs82cWVBYqOkBvm5
8yDyzmb0O30Sxi4EKnkzjqx3QNtGLgxqHkL5kt6TsDF59PK0rbRY9sXmf4ByoGsNR3KtTH18iwYx
AqUQCxrq/h8P0Jjgs4qZxAlorm9EAGxoZM0jdDQNI82rt8HlpeAt198RYs+ILri/YFbVavxwC+oJ
0GWnbQia5KzX87rGwn9i+4inyDMt6Q7WJP8DTv36u/4c7nST3zHea19QW5iQ5NIW/Hjjdf2hQoiY
/4SrdRp98F3h5mmWCPHUNn0swiXeZYd5waUaJdApviTIz2YRrJjcSm1QcW7oHp4i9GZHb8J9/ksv
KKpwUNV9a8Uyhb5jTRfMGKaX1ksvSJLu6VewRWDp058jNGrYODHtY2kHdaTIe2fF2tpC3J6x4s18
+LyW+DGuP/f4rRkCT14UQnQjvaH2GlowVDjcER92QjWVeh4oLTBdtZzqHV0BZtLUEnDMrevrjq3V
mLkse1hTUHhfX1ddxwUCZqYH2JQhUlvMmVhJgw0oKLGfh53hoFTpHXENMXXVvG6UCdaQBq/ww7Fs
oFJJzpJT3z+XHlBGA2Rl/tIMkTwSfhbfvHlQALmg03/5q9x1UrG4zKCHCvrbhZT/XAAouYFKMiYh
v9Id6iuB4ZdYth9JYrEK5FbbUnBw4euNyVCR+2AfaRNfHb700Aa5rcaZjIe4NJXNx4Q31OgVR6ZK
wlThFCaEQSDc94Q9nfSDmSoIZObb0On2Z7/PuzMxbZiXDrlJxXGlszOJkW+TH8pI2E4j7xmIpQdB
6pnQcJ7l7GYsXt+6xErIhZd5e3ejTw9LbRNO0QxZU0Bz92XZWL5xqNL4ucZnHu9GORYA2gSA9bA8
DZ2h4dRyGljj/q1rDSBkPV28v+cXmzGxYwG2OgWg4+l3pYUkPZoO99MzW0oUhfqwn3ECYCHkDwEi
brKDqiPYfO+knf+r74APINrk8ancEdWOY5tP6br5DzXBo3qodUCiRBTfj817AIBxeQn0HSfauqZt
V8jMOHACEVgKNtXJLIUlZFRAuaOVqXxRl0w7NZrfcENnpcatTZbf2N0Ywefv6WPGaq6zqpyg0TFN
FlT1+OUbDa7T/5iN28qvf6kBg1HYmroBhspBG7EbzYVipkFvZZwnfrFFL2TtesD9QYZrhacKi3ZL
zETFGckhzbkwUtlFtRgbCSoXihVqXlPFyZ6jxA67qaOq4GyI1rk3VWwaof+emx7kt7S7tVzLdEHW
OY/xoIejs9NpfbEB2aYk7NMjMRSMj/DXyz3dyOoZyvinLMzs0J1fHDAZMJ2WaMC+J0Nd/3ihZx9l
3j36PqcnjJo6+mVY8fiuEU8+oIvZSW9Xp2LnOAUIJgkrypFRsjLRT7vFUfYeJYgrYNaIoadZEqjB
e2jmQB/ETDPo4B7vV0hcKRhce6JjhxUSrXVTpQlZIvSpJl8+GEonz+OBDgerFESrwA/ndHDHqoJU
w009cHzygYHlTFcZcfiEwFQhkV7VS3/2S6MSouvXoDA2baSmcsTh/A07IfSwvpNNGttykme3kfLH
zMBtK8PbYW58TanEdgduSsVKHt8aZ0VRq2j/SSrUMGyRnw70j6E0UxzFXDN/ySIYAb7HHpgupg1I
b7tsrjn/0qZN8DQrZ0Wgfkx1aoCkTkjmJ1xHtLda31vtMxXIxw7Xua+0uKTq0jKcl28Bk0+ZRZt5
txB6Mv8Pc6qhSpIBrAFmSW56xArQrlvKvXcV2ywk/8ty6cdix5MWzgc4+KbXBvbIc/U3xQK3fPi3
G83CC9NmXnU+A+pNu+q8LhHQvG7jNa75QM07MkOmsbaTDYDkaCXCoqxJZk9Nbf2KgKkRSce4OZt7
HqxRNM4IEt5p7GBza/G4YUuN93gKveB7EDgd+iLKf0kwiqVYApKJw5v7pCCiRQKJP3ZLIcopQGDw
G/ssxXceESTZd2DL9a+LQs6F7Xerm34kCQcle07CYAOYSXhJyC2kVymDclrQ/yRHMN402w0NndOd
C4S8nvTzVgMMrKkpWsf25YhHZL+jKQ61aPEfom6h3HpiV7tHO3RWAXNWKxqkVGz2FooiqKQr8ofw
5wdkV/4UEkV0E2GWIctyodntRq64/2YiTjHc2P1Tsfn10A3Cm1joPzut3c/SKEcwI3vU/JYzygNL
67fXep7omTyBY7LnL/8u/hFe2W6dCOCLDPSA3O5IxP4Lzg/VbIWuO4kVdLcVGJ2fRiHbYoCh9YDM
UQ0m2oXcoM9fAt5iMrL1Qx2/by++cOrMCmmiZ6qgPJC2a2W8pYUPAfRViIQaOXgI27oDlMTUOHea
DD9bFdb9utLyRpNXWVxBhmtgAX7vvK8fFl+I/giOSE9y1qRMBPA+RAs4m+ejnBPun3lHe+vNnUc+
eYu7HDS5w+LTh9ggL68r83IGyHpb/UCk6L/lbz9TsvS9mFCHeMay7LOglwBHmgaPZwYLd4oZTZUt
DvlWtYM6pFU9lVSKujWjyiKKhmzYGGPKZdPZXtG9ryl5DwfUh7g1Qe5IZrKYsqcA0ahVDAmiIovB
D1wx8Vw2R+Sd8K8UrvOS+EWyHtUgnceMMDgPFA0fvbqfIys6WanccPXdQqOfGac9KLPWL0eRyqUn
F9k6Wu4/RIQTAORSkNOFB1adMkKGVwziK9IGq7kozJz6uBJ+cHETEurTv1nuQtDnzQKVwWoK9FDk
tvoHoUkE0gzQ8fh7mqIdYUMGiSaY00R7sEuc6XERF81/3QoJuItAqAWOxnrMnSgc9iCURnaolGBb
fP7M/16b1eQilBmeyuEvsTcdFoSw2oqt8UpXDhKep+V0dsSZ+xu1V1VOpssK44/2PgOGgu2Zm9Qc
xUqiqmTMkkBmectCBpcAbQ9JEY83QK7+NPSfD4Ja8ol1hoijqhva6N7bj1NFvN1g/ZGeTTrdJw8F
KXJ9tiOjpRAlHZjTtv6l7yF4G8Piir2NSXFjX2JkoMJXd/55aCGyxSqQlbLcEZYZQULP7c7xG2uX
DiWjxSUi3AsXyNJ6w6NZpnJZDdXqis3MCkRDgqIRvLeQHIb7+3rDV7BNVui7JC7pEA5tqKpag4EM
tC86OM4Kh5PiI8h+MtgC8NIH9OMdiHDaHWzTWPHYaqAytxKWV21toO+A/3ZnIX3F4BSGWV0abXAd
Q5iFSmuBnFBa3LchSJ/L9jv2svr+2Mr98e/EdpJqeHb121pF9KyNPzrRw18qbKxtL2ARtYbapKyL
DAHei76cGo6pblNz02590q2CvHOkkAkilP88QsmMOt07C5XTT9AxCV9r4N5UpQV77HPq2bT2KXG8
eKdIG0wY9BwXfO2CNEHFlJLuGInsujKzYVSBWe2lVlRSpKW9xlHIxCNhFqcky2eJqAeYauX0yJa5
0dCIk40HE80Kd4dHHPRg/Nrjj1jU4DLdoyNGCF3NukimepW/FGkMEYbYK00tABexuqtWtE/7HHsk
41KBHonPYFBpgS2xcsuXGuKpq7QaIFuYyZ6krB6F5DDR5aoQSf5Dl/2OM1gIt5Ntf64l/s+gKAl7
vaATxB3Mpvbc0nFBRo5s3Sx6ugA+wdHkYZqqMghRpDfzplfYk2M+ld8CDX69u24CrM0InrKfzYCh
k8ydygpuxddgPhjzJJQrz+oVPfJfFTZtzvi8iKb1eVawWrV9aaByUIV5SPzuNfNYjWRhqNipVkMx
M4SvgDCVd5Anup6tXMUu3m5uDiOAgI6zgwyp3orT04m/nB5b2XejdjuKtebi+SHKd+pcch/pjZi0
jMwUFyAqz/cLSFjT52zZ9uBPUNcCVof8Q6nNt8QREuuxhFCSvG2zcoo4OCG8YGFBvIh5ELJKfwvm
h4yPshqqOIixSe9sLIgs4ufFXvdGzDlWO1ZniMpcgLJAQ2RdUeY6lKbx5mdreMz9TdLVNM54YQF4
oBPj7LFWM4UmoSv+MTs++0oQ2C4gWvpXfhAocyRaevahF3O0UV9XWNf6baDnPbNnbSx7CdBDcKaC
Y2HOkm2Ts3NRlTmVwzb2SUl+cHF+eXV5+OXB6soDKj6p3AyQZIwCn2yPm+XrLNdqQMUr7C7qFRqb
aLGzY2gvMNNqUJSo74Q79cvGrTKL/TlAILXDtuFK4FCzFzNsR4/tbQt1bvMiUGkZIDov2E2ujwjZ
RcDKPQkHrDTCd0XDbd3kwFc788cHTksM5TUPGOXJTULsW86UGzZGAnh9cRGx5pwGD+hIsjOt3oSS
pY7+GQuk4OgpV8ccgMQOhNSpvHXx2fShP0ovR5iaLfma7ZL1U/EbA07I6iPG470s+/y77FLnQLl/
Y6rRVewPGR6DXDkB6Ztr5Erz52zxpZLFZn0LfNrCJPC3EuJDe14mQaM9KQDUqvo3Dt27WBqZiV8i
JuGe40SBWParQ/nCbhc1p7kivnjmnWOHVxfV7YzSW4Uwky5RWCojSX3dDpBDbVjrbH/Szbef6bi8
+9lYMfV0RX2QLjZQVAJSMF8/Kz9I5DfVgQyh26FjYwr67Bk0OXF/9jbiWeJ/C0UJ0C3kKlI06w+a
JdTNlH+bbcshPS9MHLrJxEPK6nOmH0G/tt0WPDGlEaC04tVaKLprIytfL1JD+dEHjGZWmniJuim2
g81EvLpjRBTkGSz3yAPMN/NRXENI2AO1M62QlG/F1qQ96DaEStunHp+pZKu0yQppF4jqLpQUPJJJ
7StPfXCA6vbhm1vybpTBj1YcIYYM/UyKvXAa0NMRAHr9xtPKYGeU5dvUZ6+QzAoZ5eKn5wKf6g8Y
DPzkjLQwVAUntT70GcqbvNPpRSkYuRtaE3o9TJIFaIefjPF9u+NHtl+aulqvMtrLeO1NKLs1b2D0
ZIBZX74FnW7BC/KRu32JW9/e1W5uph7BPY2lSjrPu780hTQBUMDeYmIgvtoBImGU+u3ZCgSLptX4
1FAh0gI7yky6+pgSIobOhYiWhUDBhHI0RVYKDUP/Ag7O6X7PeYmMv49AWrjnZAa0eLyC/VkHKzGK
4t8iEh5fWjOlbnyjzdDrws/4lj/ccM1Fds0mLgQot0St+pJpGu/9Ui3TFuADZtJO/90xz+GKs7WO
4cEOR/6pV39AMpTpFkvkapyxZLqPX82hhA4vjpORFsKLF2dluz4pQ+pOote+Yu67dozQI8kKyBLl
ZKDLFGaZRaVDaYoZyh7imIRowrogPaZJQyT2csQacY/R5I9fRq1+PYtwGMgBb9X4YksS+rFkS1J7
U8en4XEwPQXw7TjKeXxqoYsa+E1GhJLDcxVAOw8DIUs1rG5rA/G3mICge7ewVPJBq6xr+ReoHapD
os4jAbri+xfKNBqDk1O6k5zq4AROYhqlHxcuWQnEBhPq86mdRo38B5dPuHrpWZapcBqQL75dkWdP
eTkdVUJmpf9OZOQ0Ysos+sK6ED0rb3t72GsVfQf4ZNCRWuBtCvOerzlkF4cLCEovZ+G+K+IFsZs/
BRs+QFADsTlm8OpWaMmHVXwP74m1oVUrbSV3omEbXLT0q6ix36Nep8N9X4bWKehCnDzpvQpQMGaK
zfwEt0muIv59rZi9fhCxgebHvh5lnHGC5oljiIaEuyQJ3kkUCqD/ga/Gl6nVd/EO2PIJ9DlGzLSe
dBA5BzCGmSA3Y860ceLWAk/hfJCmy4dJi41FR1xmaK2kiFg36MFOyEjJ5w0izB5pjrXiFJR7X0ry
+hEo36KVQX81AHTrMqcDR0ZR4vDUDlq4EnRYg2IKsgzSw/CCLqcX6pNaiTlwVi1BkxukHxkYCeFZ
BtamDUDtJbultK19YABG9R8nUBS26C0cEp7FGm+X+Ml0RMB/6JBT4iLc3Dv4uhvdI0pJ4j8PuwT+
OZtYMU+kLVyQ6eLsjsPG+3moB6mh3iGk2hjb3soXqNqJbJYK7hJcAMoY034uMwOGN+bH9EdQD9Bm
03+JmBXdH3SCM2Zxq57b0ebO/kw+GMjvpkqSAgcXk572gpDCPwhA+jedjwhVFm7iwcbrv+TB6hfO
yJ1BmhjZWcKjr54WPdQZY0eS4f0LwWIBliWSJkrijYcNioSixccYNZygiFzAvZ4adtJmFSCAO6t1
ND+MxRRVABmWgvK8fb+ypGoy+yWbW6MVQ9KbWGpR187Ec75OSHfigA+5MHqEaB1KLnD9nJ597/WR
AFNp3ypBnLqDJS5NkmL2bAedlyDpRnQzwEnDTE1F0nrQl03qimHE9tHko9TkgkrXd4thzv5srhwd
sdxkmh7Vus8smVAFWOfFBgjPPsK5OYZ0dTk1J6zU44ru/MZotHCsKnnaP+KjZDTzutjOliEWmhXU
GQuAOopKYuZxEYIoqd2fO+eivf8vqkjpaM2MgMbhe1kzx/Tf6lC5vMjiiHLrUD/gEq2LL5oR1Nwf
0zSvEPWQFvJCHnFllIXApYgBFX3IWeECec/PfT5nrKO1fmB+HIrtjN2IRCjTtFDC5HWx5pZ0GKyw
VAtGwm2lW6lKhGd+UB15jXhEo4DxdCcqrW2KrsfTpTnsaqxM0fLUqVW7q77W+n4ivthmF50GCeNX
+VdTAq9IeDSAaOLqeJsYPw5/AvNjLhv/wYsGWbNDvxbhPbgRY8p2oqhMBP02rCIITT8AUE75AFMl
KsWV0yVvOHhL3dEwiw9agb8F6YAg2wAiwCfHdtVlJkzNu0BpoRrn8CjuNrXB3dXWh4I/EBYNi38G
SXGKQryCmTyCaOBdRoYoeDsV10V+rZioTlUd1F7NJk18u1NBcRUol7aoYWzs7SA+mrBcSXqzP8rJ
kjQUsREA88r2/zkNHzpdNxfdXagQh+qBupd0eUADmV0j6K15TWu1O91nwNCD+wgkex3WgcdoYBbX
gCsgd/lMJVtA6RUyW9VjSqddl3qe1F09lfpwT36lYKci5YN9fUclhPjThax7KQExTSB7KFlTZocc
y/3YnKhaKJVQPi+01qk8jocIndsiqXeL0Q2lqvYCT1e/nrHI7UIZarnnbPwzIbdExgOBQtLGud8E
ZCw90pOWrM0HLgcEzNLfm1IlX6oP66hwLpKYJY646kM/l1YS1w2TJBIY97R6KWFfLDGVfWAEZ+OP
Xafk8d4z/gpsfvRXtHZ/i/H48i92zbUcTUUwQeWUIy0inhlSEoHGbtBr/Pr2ighRgk5mjeaBIsFL
qen7pIZGLR+TJFBsP9242yFXRjcE1UcgBhqfPRRRIjJiaWh9T3exVGo1RLdbUhqhqZwU6PhcBJT8
7lvOg+siZsXO/DsxF3g2JhuILem8Mk4Qr+uLVJ1U2qj3ZYEhNYoQY3TXbXwgLactY5nTDMov/HZK
elLxicedQD+powWTvMz9WLffjHgyRbo13cWLY/B/IBKGWWEkbIK5etHsa2rlw3MfNlccxMkA4Dfh
KOufm9uF4lWYDA6+sqECHN/iQ8QWFh12BzGYO0isLg3AFDlB9JpUZNZWr6lJqF/x+63ysFMLd5SW
BezMrm11TqgZYT2BGjOT3KcBSvgup39fkYiBaYaraAa3zatEx9JQatb/5vYYaFj7+WeTpHDmZbuD
jhQq4z1NrucYXrp5NOaYuR4MzbIkmHvLyyB5UZ29zvpEokeQ8Vf1oN0Ce/4IK+SanLHFwuUESWp5
/mKycTiRD0nTu5mD7wadU2A43cPSdCtQkLKeC0dY1DtUZekZ2tV3wrh77a5VUiACcnAFhpoX41CW
o+CIdrvkcasLGjPaMSlZVRDE4UK3yxrhTcOasY0x7IjgsJEiFcLqrMxDbBXbZ9je67/FhRLgPg8z
pd221SvdHPIrkM6jtj0WEhFyF2hjVfdCBpakqR2YrOC0zAkm2ty79LCFshA3Kd5QDw9SUZgGjz+3
3RZ9CDnE/ywmtDSbMd+Hsz8Bprg2ztt3wyt4x7bC3NyItyilN0OsZY3bN7OKt7/gXEyWKe/hWcu/
zCU09dGCj5c1CFq8gxfAFJvekrPwS/b3VO9ubr+ZhjoFBfesaYb3YxtUH6Kkz6Ql7rwWyKk/7f7T
1eXQePbZa1o334yNe7UanmpQ11A4Bp+y3V52+vdUQRP4s7QeP4RCLR3txnLB/42ZIvCf7Q8vt0qO
EJH6fCY4hOLUSkrZHnJgEU7giU/XkYHs6gzRYpHHkd4lH1W9k73DB05sUpNSOLtepC6JksxyRdoK
w3NPgvhSQmUyJxbzmK4DCOcX7O1yLU3Hwuq8952SuY4cesaf+1kpkH4XAM8n7Agic0IbboLPweds
R/23Ghb1BXP9DWkg8wEpFlS41hoAhFAwTNs/EDvWrM8x1l/VP83UyjKKEC+RfnfBQGqd1yaHTCBD
nYTueBvHYFrWo8+IyYy2eAJDgP9/f5uuclu5ApSbfZcaZ/opa8a7a9YsJjU0p1nI34F0jP32SEZ0
qbswI34dFosjh3F1WOpM/OXxfsQR7DMkwUkHpURObgGtsV7WKSzzQqDaPcUKzZOZZffBvwRJymRc
HA9zz2RqGACPBiF29dmnh97GWlrgq7kVKhfFQFQHy8jY0Mb0AIw6VYarsOnvlY7jRg7l5St2eERf
YGGHryjC4lcR+R5tMPQxddy79GLdC1PEd2gARfZz9ZOZqp5Sp1hiU/4QhpLHPo6NtjUVWsg3jMj+
7mjwubVE0eSp8/R/gT6Kxi13gsFZcnhdu746/MDh8CTqoqrqtL79ZbD7ayi16aLzJ7l8/+fuE2G5
8laYzfFt7ctOEq9VaI9XEjaZ4jiepufR+U8iwIN5D49zIp4FzeGA5b+7fYyrq84wCELICITjzlda
oLDua9z8Gjgdy9jvrZgnDBIGo1KgUIVGDIvIxVcwqOYec5rUTn0kUdqKoBXp1lspQTk9domTC7gp
Ms9BAkOigHrDFCvmHU3CRNqd1rnoBn9I/h1rM0nMqs8FKTpxfhcqgEIx6hNUO2f7tvgsIs2kPzVE
Vw0GsGWuzbhg1sq5Wl1sy9U8dbwDkMPvrVbD2JCkZdj8un77e10hs1D/yRsa9nEIQZ9vZhMFQcuI
pult9QY35/4j4bbye0zS8YgeRknpRjDjid42+W2cs25A4nB4+36DGraUAeSr/Pq0/w/ij5tiSjT3
WoAIEu7dzLSp7JhO2ICdHqofBg7Knd2jLivansWP12HUS3UQhv9rDokipYqHAoH2M3tl+tiQfpAw
qL4iH1/ai43bXsYyJNQQ/TmUahWEXHePfk3nQJMCeaqk16yMEu3z52WMDqBaQ1GKF1vI0QT7imYy
xT9IaP6R7ndS5d4i5YlKvMG9jn3KqffM3AGZadNqL8W/bbcwlxu4tYzhfmgwTcWKPc0RaZFclhJP
5zIwIjvhmzpRgGGSpHmRQW+QS7ItxKYx+xKRlN1PhyAvj47pNvPPUPwy/3xFzDfRfWyUEYp9+4Hc
HwPhgVQD7cTjsBVF3eL9Li8BYw4QPvUpNPmIFangzcnB3e0zTwxMAPpPUCZeUpKXwSkzfgAFiubC
IjrZcKw2xNexj/WkK+zH59H3d86XeQGfwQa41ELV1fayCSNa0RlRegBdblWCDczKPkrRz2uW0qwz
tK9o4c694+MJs9oll291KHq7WpiEQWwlteZCNez9PzMNSoL8G6bNVsC3u3ytr8vnQPYlZ1rsnLsq
YXqmZ/kekTgG3kmSg/Z2i9Ea0qO7PyAdqoIwovF9aG0n+kG6Qy2+UgZzt8rsEmUPwCyC4c72BbIF
LBstxI3jzPjEDnXVJlX4BzXyr+UsXyhM+2AIgAAf9zxj5OJ9Nt2UticpOVZC5hlHRHXJMgu8wHxR
Fze7ucjbrYJ+hJeMxejMtLwphamdjRauaF41humu1MVsQIeh5gHIIFGQHuHeiIqZaVJjA2o8bEJM
9Ak96R7xIyec0Jz5Nasic0LljA7ZSPV90MbGuG0lTtGl7ZUJkMOjVfCJj2R+/nvexdsbdh7r8scn
SRw7sEzAv30pcgaNx7mUosexKt0Jm7llZ2EMq8yxnEVsuymMORJiP3MIKDFuUvsASAD724abVlQo
+ag7e+nw2y3FrB97zvTuB0AP4yRYaAjfCYUfKbiunKpKi416qkX0TDBSGdToSCJBgTjT/LfosGY+
fDqK2HyPv1SmD+zFJi8l3OLTjkGIUr82RxKdqsPA9Esw4zbabBOTZ1FlMl7ofICbwKZZFYSl2mvU
3jUDkQrhn4CiEgD7qa89bsKsSfw2PHDoAEeu8OAUni0Gkjay7zidm0gSSf5BXxkS8mHMt5n53vCf
2lHZz1i5K1TGXL0IaH3m3hHeW88R4vwcxrMJ9qgPaSx5TmJGIvf444lrkmLKORBnv3oPPkDgZbgN
3xFJ/H1HEbj8TZwa3erdLm+n4fDpSsbnnMGvy/At8/XesZ9A+H1RnIDWBn3YPCsTcF55qGh2Ho5R
90pJ74RK2PgD3jFm0dGtCTGOh4jh67UUD2GH2pj/IrVwSAZwjGVQFxgowhqjGzJkJoxGFHcf7Ght
yvailrGSlTlA/hoisOhaCyFuFpucGbkfIrxYFq8B67UZaHiU0LqW/BM4h9sRkAf0aKdQpJFvKPf9
12Vyb7sncKhbQBS4Efq8JvFbqzB8Ck3H72tDj7NEIDICmdkNrpFI1PDt+snkHYia5n8NKsA0+uWh
vBbK6FNDpcNPWgS16cJBBdL0H48VrYuos/xdeU2upFlTXEClRVl23WAr1x92yyGPuG4FWKV34xW6
Y5UG6wIq5zu/14MY1reL6NayhX9oIYQ14TeGyqfJvrB3o6Y0eqmEFiImQzMWfo4RWFkonVbxpwaH
/ylUPBBY9KojjpDXb75z+J22JYa2Ccou2vVqVujqyykDdet1b3560bdThdtIH2aTlToPvyQYK1KQ
nYCM7jvio+29taBPJh4lsmc551ZxAw464SpFgHBNzudfFuhq0l8opr/EBSMdvqJUlO/9NqS47oTI
agF4hKDFTuOiw63HbpvX9aRJIfH1LQBuVAPXf8VlYZ8DO17OVJJ/7mb19blAN6hxS5PHkiKbD8q+
qzBhdUVeFjR8G1SiV/L1n1raZB+6WyUpFJD8uFnIqN2XowxECZAKMi10x/pOcQX/NZe+tEFOe/H8
SFpNWs7kMrUYwS7xgEbYjH4btOfE52IMURCvYSWvn2JjR0woMgJDgHEZzNs1ggnB5mM7yw5fAq8w
0WW8dukRgxd/JNqJEZma0wrguw7okHGVPsDm0zQNm6Af+P/Su7EjSEdufwkhxHEoBsHT4xKEbisA
AKknHbv5771Jaax1//nlKQxK71gDVlR3FPbx+SJS1J1VCB7LNiFTpTJmH5hyDvOe9oIbFJul09BE
gqrjDqL1FPdG5sEc0WNgngNqjtfQpI10nREQlNUf/MTDmioYJHwhwhjf7OPkxHDgQtJZwL51XBbL
PXIh9jzZV413ynXA0cjK0zxNfnF3WOT60vmWY6SFCvuhjuCN93RUX/qsImWDXbxYPRR5vgxtTg0e
DUWg4MOBXCJEllDtLS7yp1bRtsHgt8no8sDrA6Gcxn5kt5+Nv+N2JHGjypTrSQRoT/CKQJC15xIe
R+kI1GYgFRpT9rfZ0MjPjag8ZokdRDSAcFsV7nSsYl0pcJasKYKy8j3U7ppiybaZt+UP5nT7sk8r
iA/N2lwUJ6w1zVc/AeAuGE5XlY+FWg8/76ef9dPdkTJh5IcUdDvm8OB/1tncv2F4by/znCI+8ohL
PAV8OQI8lBu7k9Xa/dTUAQGoF+8HkB2t41jTJg9pz9rL1UeEgeYcdx3OstRWZ03HgKGS/+aw6klG
6tP84mHj+rawIqEHQsMye+1Hf7YhI2Mxu1ZPYmZNAR8lra0oSg+8ut8rKEhFsTVv7Zafitsh8lfT
xfnO5h4M3/UFA2xvqxpwo4TeXh8addMRHtrO9TkU/+AwB+TwuU26t9rXu5FcodcCnhBbgyAtp7Nl
xWgmHrQLZK6+IikhgYY9BqhfBkl9zKf5QmFjDg5nh4vLUVFGtdAxpzGEkQ2dJzM/MTNnGfR5cdQd
PY7Ni4DkfJM5AP79UviCPsMC9ZrbKHCy6IGKSK1+ZpkHrzVV1mgiw84LCkjLZuhLIw5JZCRejz2q
RYay5nVsh5rF3USl4R/gZQi1o+afcu8pS+f+ki3C9MWKBFFUEByKG1yiyxc0wEZjhTWvNWIFPUSz
SEIeksa51xAZAR+KgV7qQ+5XuruT2nGqkdW5WT5sOw/QFDgEB9+ybm4A1T1+qiSGEPDCUOYXnM9h
0NrbzBIQVJFUIV17M75lXIcYMbaveI/wMnyR2V+LZ9bxA3JIChf3o0xtjEOyKc6hIX5uQdsFz9V+
h6EXqodVhJYcVETw5e697Wu5kYBVGF1lJdgjZY0NgXvuUI21TFjnJpKqIgOhVJJ5le3x6Pua9mCp
DgMXGgu316HtzB7BFUb2Qsy77O16+IpgCai/IGC5JGPyiz/L4rvEYbLkt8psxBauD+etOpQav2EO
pQwy2LzMlOVNhGLONq3bytAffivzdpzHVbV/s40zrLDJGOBY8gQgeElSBonBnMIbajPK2kUqqxOS
iitvCUqyweGpzWWh2PIF8I4rfa2b1hHSyva3yVheSWAt2Ykj7VpOwRw2Nq3iALMa/4gOq7zSd3/d
C8RQi6EXQjuEvuW1PT5bl/YlGUc0R0wNuU7Np/qqJ84ZXM/AykbH1Rep/LZ5UW1XMU9sASQQdn5o
A2BSFPTYUYSRZ5TGwcVOX/XMYijYuY5mrqRBooMdDe1JOILyKZ9vySEBiUI7jLp2fBjYtBVmeEpG
YD8d/m1C0Z0209kvogGyvHqX/fmmXlrLeKzzOvunw2nS1kM5aEUc0622CggOiG42u9JVVevjIvyJ
s+BLasW3YQcbzEPBG/lGYh6Qxm8VAHTqTKbEVDEOoXD20NBIo+yCSXqSSByzTC4QP9zS68WkRb2a
SQ/fIGe4n1Q5S474qQuYjyWTL1COSbNu3nkLABzk28pH3h0FFL/4aE0pvvRUny/ScQRCE4fkCRV+
23V1sg+mDiioDHttNaznddInC+2eS4V5ejFplgisCiqagxJLlALv5zNeSrH+To6pjUZMxybJWlFB
h98bG2yv+VP/bIKcW/k5gZ1ZjKZHIcy/UwOrf2oBdhla5Hul3FXmuZh4bwzlmzrq4D+pyzbBNSB2
EKeg3zQNPbmWQLBJkJl+GTWVGV/53ZA6WuLSeDODJD1T5T9QXyRxV8+Wf+SY+uLZwZcpASsHKbDy
KG/0N2KLJFRUR9UOhi9rwvFwCVWWQxgkRajcAchSHuTM8UWpWrZNFEtgMlTOFwZRV2bby6+yp5RS
PqGykGLEjs8694k0wxWgHOVR4Z+iz5uxavlyoq1VmJUX76xrE8nHV1RbFHEJmWcrqVI97UZzO1Vu
RiUBJmossize95aSttOfeB6LrhzkUTsCA7xZqOFJe2oqKBuNif9Z0Ne/vJP78WBI/uv7sl+1HF/6
QFJOvx80oDcnaHZA3zhUEM59FcGXk4Nwtj4UJaBSKRT0BDwIi37dU7SgeK7B83o8e66AfVgAdCPj
+jS1fH8celOMGaZCdhqDqYNL68yK/wqdXdoug0i9LxGrHk48XKYkVvWI26+4+TExeds+BrMbdU+z
Fg7b/s0DXOdA7/eimjYpbQZxPWn7pq5YWmBDcVLftC8+0E6s5cA9gLTF1vE+SMjffJucB02ESJL4
B2MaiH38vWUGBzpnuNQEXS0SZ5GYTtxmdR8zFW6GP5LZe8Q+tV4A3COjQd2CP7PyF1wQU62Y9FIS
1KxXp7jrj/Ug6MAUSZvTci2Hgn+ZY7EEEDfeEuAOq1ljtYuz1hTAe+KiYe6eXZjvAHFrk4OJLAgQ
Ln5d2EC2ByMmiDnXM+VbhDueKwq1SybQCIl5w0d0S+kpErNnr/XU8V8X/cByVY4vT/DXDmhVpay8
WrqJNgJyGSbzx7AtTKloNmP+n2Pok5+dsCUtn/W3zeiyFK1OAUsGKdP0ubAd/4Dx1pqVO3LOImLw
OZT8lDjjWnp1l5+SwPHQTpowu98L+Bywc/PvW3sJeSRktR9myr1/a5zzicqQfS/+rRePebpgJ8rM
1RkZwNsbuQGj0BmoLV86U6i4P4sylsLpgHE2CuOjQsBwBsUyzdoGwks3wilMYXQSRzFcr/lAZxcF
NyGBLJTmAzxmR1VhGreEW+rgrSxIlThIYOZwCxjtGU1aNDABCHux9vUrezJ5MpcUY6GY0t5W1o5V
aefia7quvQs09uSZx0arLAXVyQyN+TeEL9UEvTG0rBNTyw+PqlNgYT3vqE0T8Ct4lsAt/uKQCXVf
itwpDYyIz/+uPDBJ5JogtMqK1Ywer4Y3Dyjno1OP/GaO2X+9BCxfXC8BgJ1nD1Heh5RGjS5Q7mkw
GRNnYf+A+Vf7jgWcqwDxIe3+25SV7022kgApWc7xfabnCMgs+rQbzV27kniUVqep7sBKMTzsE+Tk
FgjjTLjNGkNxWHOoeXmGrXdcj/XhbdAnNxYWJQ+ZkU794M2wD5K2kvwYhqCgnHsOy69UGPlIZj7r
TJARR9qYxM00eCy9KU+036b13vYYT2Dj/bmnaa49lTUuo6igdf3dozVIj6IYsBvXvSvO/7XmGzE+
Fh5c1my0LzVibkbNUz/A13cKGx/4WeelbEHA1jhU6u+sgcrRbC4+j98umM4JoqwxFp9f1CLxvRVs
nqpgBYTd6dZ0Xbsv9hivew15yxOL3lQ4Dl8IUPBUqDtqPSZNlEaX9ptLGhgpkF1R/1p88GcOT6zN
0q6ULowiFJRxW08Z7Qjh3I/C7fCCISEv5+es6Xgffn5y+zHDaOeikqPGCgkUNE9CgzbJTdOO1SFH
hT8CCny2Mf6/QH3QSmt/kHQC3i30Kv3Vfb1u03/JNoZvWHhGg/itBVFrbIaTZwXNzJ5V+YH7pCIT
9rYAzUvYXcUR1/QHSiW0/qCkLY1p1+HOBB10LqR9uYPovr3mDN9jeB9c1nOvsAQjghVsMIBzACJn
yQA/4aeKdfHZo0DErBdvNJgboRLPA+pBi7d1ebiI0IPfWY5uY6dpThSs7b6mEpdupuWdU7l9LAOC
a235+fC4f2AVJIHsOH+bZpl6HDC3hCYlSbaSh/ukvgSL2r6ydTo6K2wAL68QiVO2S0Tq6V8NNyY1
qeMgHnRCQJMW1XLqqOww4wrkflhTsgKVQK4fdKRL/Mc4Vnt8pQkNmYHo+JOlZblm9I/wqp38I0qf
7JLfzjgWulGoJUOSG0PIWRwGsZPXZyzhGkclDjVlM5HzniFqtHYRkDBKB8YDuRUwD0XlaFKUi7LO
6mRy2EvOzQsFnMCkDrqpxqWUwucYNo1Tdi+j8SEcZLHoEG2l7YDYxNXwYu/evhax+LzAYAuUcakF
UKY5R3NG8jEb8eRwKr8u3mNgb3AOzVS+hB6ibxxnzmQH2r/KrRXSo7hhG0KEP8QylBDEaKBszhkL
AUhP1Q2mZCiehZLHOkhIqmgOQdHJkfdkgnyJ69LzfvOIRI/ZjZOMxkXS1RXeQkJUjciV2AH66Inx
IC/h5HNJUdnmdCNPtzy3YJ1QOHTfI0Qzn1tGThwV9KV3NSfz7tYL8UJY4xrleKOiNp8TRZL5I4mD
DSPha6uybSYxYw6Pf9qTOoMmbrUPWOCqcc3hik7ciioRXxyCjOdkjCyUxV4jYF9+jMTLv7NTrfuu
gLY0B7RdvSdxXJ5MJ9uTyK0gS55fuStD+P8/Ck2p/n6qYmm77PXTuSB7YjVSbWJ5PU4BeeB2hEp7
+5tIJ7zgSbzWtVcFsO5g1F7TPb7fzkh6UJK3AODsnvl62zF8R+6fFK9//H+T2mTu1dqeXwumtUnq
8S/XR3+oV8+QjUIDhEpf8dqgOGMMl8uQCDJ5sXo0KVMa8ZLxdq7FwLTkEjinXbkqGxLTHe7lAILX
qAFJPL4L+hU1JkeO9DwsoXdRW39P9zKtpwx9ZviRGudeRCdm09FlOaAsjbaSo2H8xqsePTVimNRZ
+636zIqxhEc+QHG+GiA985PWecqRT/dNXcYozVVqrbeVmcWzSfcg0K63tv822exThHfPmxZGAjW6
86Y3Ro4dKiEk1QS7x1qQlm5eyXATfT6y570c8/8hZFrE2QDzK9SUxVV9yAH+Hq7YyxiZWBCgvqJP
G4rnCqB/112/aQleMj7NAEvue71hdjvpD6Tn2I6RCH9tVYj1YSMs8APJaIEuqv+FbiPMrZKyymFN
ZxY89pY7KoCMWexuoUHgJ84PzGkmf7io3Pq1vGHMnK2mwJfKLUHt2ZNRIOu1pMQpJEMk4KygbnzT
NKbYhXCWRqL4K5/DmBZ/lfThyrvge/1AznFWlID0wDbafBd3lrwAu8qDmZp+avXkEcNOBXB9MDQi
ZD0aC3YscZ9isx2UAjRuXGmA720g2iW1SDjizMWh/lFKOcx9+3+fV6dRHiIvNwgNAS8aHPpTRL7E
m5O/LEM+e3HGntKAnooFUKWv1HRoyC2j7mkMV0kn1xp0k6qd1tcUMH1MVW2bkQAhrLpEsYOvTNcV
FIGB7jq/7R13UWnMj96Aqykn0yeU6QjgwdZ7ClZIZcTG7W1zJ0H+aZNWbMvjwyiz2URh7tlYUme8
j0AaQrT/dzPrPFkOnN2KGb2W6zN8Jy5f3A025L+tizuSRTQlUP5vqJf0jHi0mLleZzR7bgoXDlLC
MRM5EGRUvu7NRviKyXyPPAqFww+XdH11AyxrggmhBk/kGxVUk19qf0R+N/NweZiG8n2sXBjPavl3
HG89N4o9eLyQy1GYlyDJBbR3d4ln2jyvKRYRy9x2zX+htF1NeCZ7/SNkjG2ZRuOL9mP80xA0iD/T
u94zR0yVrF7s1mlbw9gGMU6PbuSKsAhzf9sf7sGWYEq0Mz/f1c+JRrPosFeSjxYwzITs7X9r1gw3
b6KiYvj31CdMTJjVqFMW/a0kl4GFFm9xLb2eVEYnFihbxYhhcikKsoYc7wDNbDWzySVvk7cw477I
USHTd7aMw3kSztuI30Lt5mv12wq34V1a7ykqqiq9J/eMkqEdlhDxy9yh0GpWynWCTNb6iPmZpQUt
H3VU2hqYGJV7AEplaYnEyvtwseFj8282/ygvrhuPuh1e24Gmk1e6af9HDSEbjczF0cjyDgl5FhdY
Vg0vS2I54QEaqR1wQvSO7hR+M8KNGNBJkjiFRWY3QI6rrMtXNGY2a/phhgomsJR/gq4dd7l9xQR9
M4dCNiFlgXuQ5a9ojAyHcBTMjcRMdno1Flr0gg2Xbw1mG7p25gk81uycU/kkLnkQ8vHeuxoQvUqB
+sTcEu5aB03MV2p8x2zx7nNCPUCM73TGwowBG3AMvfBaXZ8OD+/OOCU82PX3fR0vwl07AufP1PO0
7XrLs1lVSP2KmvKM9DDOafQzFLOgfyeoEiZMpsQZYrGfhfXQ+RNVfZjVNp8HdhB7wWgxwo797KK9
z3B/347JokmT7/UIJR+nICQ/ZLTDjUdrN39J8vcBQM9oEndVZlpzN/7FMMJj8/VoyR0ZDWsp4qS2
zNj1XMeCvFab3Kt+Jl33Dfk7h63ifcX0q/8gRizyLSGvm96nP/ku9piOJ4rCVl1HO8v5USn04765
KXZ0hLWuEEaTlp3cgpjF2+eMTKRDk06ubpWdmG9I5Q8Tgc1k/QuWgwrXHTswNaQkOSS2yc15IEWE
gCYscl5Gfj6ibERBZTLojBlFWW6MnI7xiBPyRSI2c0HRgZgDstNNWImMhjBH3K9dww2FHryWmvxO
49wAwDYESXxsvvP/bNRQz78SlllJsi17dOLiYJ/Kyyog5/7zXi2ptQfcEqA7n3NMXvMmfPaIIJ/d
EOxSdXB6o7YvPN+WWIAW1D9u1vtQ021yEnrgS/g/iDHeABvnOFfiZkSdyKIALEH05FpSxF7lZ+6n
OlPHmozG38IaGYntK6JfGXizhRY8GSud/zsWOch3LHCP1TCMi2dgovipFPZgEqzRerNKQ0nHPfjZ
p6LrjHKQq+6GFoT6xbZv30SwzMMuFehyFgb/VVBw5DnOlOavrsW5e+Usnb5yyGg3UQOaB9ayXG5J
3jXTuG/wwCTBJL/74ubP7jf25w4i93PeufKAMPkEgKsJjSxNpXNamViAQreGu0TZnA2hJBu22v8X
kP9qisWB6qIgCqbebrlrTVLp8lKAsQMNuHRKAcZ03KS7vcUJEEgBjURgumZVCu4Kp5icsGEwKV3O
mXrIMbbYN3NQ9hJd3hRjRvEL0BsbV/nBvBceovsEA1pG1pgcXNOrsRyzUGEKI48ZZKL3bChdRhbm
oDDzfQxb8p4NIvyoTwEjfFHuy/trPjfzP7SNsJOILz7EALnh9BmzO/1PsODoQkd3bmPYUBbV44Ru
R2HibCD3yN4NP9QGGgm6MEe6/TOWozAoa1ApFoGPmP0rmIKVdhMDvWwuT6tKkNBgFgys8SPL2Fhj
zgeoLekL64I+IhONK+xSv/69UOxMPGO1BriLHIWf4HYricfcDxyirGBVjceuGAR+8MVb3w6kRYSj
e5DgJayr7Zmg1gi8u9+64tsNM9uySbQhsIJF97whIPJv+xfIAGRduGRsE0n/YVN4XVmO2sD//lUj
jHqHjWXmw3Tqz8DM+Doxm1Inu3OraYAc0LY0JZIc83fhaOCUgVy2oUVaZQHprU8N0BKOwxLf35Uj
8Lfuvl03a5eV+RwBuhfAyaA5TkdIRV1JtRsYljBf/uf3MGDzBjlD58M/glIZCj+ywM4cQfvmjaRO
lRgYassgad5khMZqKj+ELE3kcBNqNfVJezoyTMdVSWj25O2R6jQC43ThsUZvpLczLGoVME3XSATh
yIThBtv5z+40hSaNCQlqpoaZQcn/oANpOXZHk/Xq+9TeGXl7MP78IEU7suYbPjm7o0d4Rdrx0syv
4EXr4M3PF+S1yDv7SRzjfFf2dHlvh2O8SYWyDw6BAsKfpN4+o6B6fnnLZ1MNc8MUyoH9uupY3gML
tIRG5Jiw0Uskqe9KoomfHePUkWm0F+fRHRs7F9+CEUPLKkDcFFe5v33hsTcsnBEa93o30Yki1O3/
1+JSJotcTEqull2zFs+MRGIG2JjpE61oNcHG3Y8pyhKlHZ7FRQDekRGH+nPM7XCyBJikYrbzbGJS
dRFE1Iu+asCx2TA5qa1UCjBX9Aar1+CLKlXsp6w67VzQ6Mw2fePaKdf3fNiQPTV34gwkkU3nU8Wm
bMa+aEXqHa56saJ1fWNGoQqznQgQqyqrKgPf3s49BfWgqe2F+QXYfMhdhQpI8uTFIFqg10XY4GjX
MtyrCPrlgpBj/IGWtFq45SUmsz9J+EIE5Ysb8MLOJ2BQS7OXaBArWQDIX44eDZLKz3g1khpFuTat
rITGiimNGcWZ+kTb2RjzvX/XUN+V3qZ1g2+R43GH84fFfObhHGfxYxLilFrg8MN7EHLxAWSr1OfF
MaIIKmztkPM5p0foUvm/FoM+wNqj6nz5Y2MLHXeTqTTwATg7vs4/ifHMf/fciUq0W8vVXvSndzmT
mG/b1hg64E5WmoUQ7rf5Is6crEa+frZ39mHFxH1aRvv/WbtLyCjJYayM5oL/uyjH0iw/e6mDEv13
zYHIYgd5QcjNNNJAQFWnklwXLNpnTGPeoLxpOhdhH4AHAxAuBWJw8nSeNir+yFLcGJBuJA77Y4y8
4VY1bTP9aM7WalKfMPF53vVmMqyqa4MGW8fgwZIQCCtKBMMub0eccZNX7mdlcvQUWyGiHXVujTvO
G1PLUlPH1AG4cQMBPDjnnv+ziYPp6jmr+34vnK63clqzeu/HQp87Fuco4i+nvwMw0cfkxPBOUPre
np6RwpMYI47Glo5n/nYoJrNH9Blu0Rho0Qg+96cL/pjl55X3UzCRTbU0D8H2W9X8d3M9Cl04wvIU
ufOiqq5KWEkTnqli9rjolWGlbmdjbVQvxLhmAU4TgCJs3IufKhDCn3hzCPiz1da7BaCVrTbZIpe2
aNS288YAtIPoKoQu4TVyPP0Gz+4aFLNO3BhzBMbRD0UgFZHMrzaBE0uQT55+LG6HBcz9oq1dADBO
EdyQV7/uynqkwj6eLkS2/RqXU/5j+Vzyeq8vUjkVhuIT9//PyyqCdBeSNGt10wYbwT/pNCiz5xrx
7xy2C37oGQkyurifyn3NEByEjMdBKgHHuLUQGECBnUQLnyJrw0jowk5NdamrWZYNmwM+MyI1HN1D
KYcZAiUUA0PqgV161pGFUqBuiJIxbJy1vrsfIgB3EI6ooDVKCvUK8T4JMT+DE77btPZlWuhN2HMG
9C3HwxXxivccwi8QWQhxu7JM1Z4Sbi6+cdEtrb+8l/ZmfwXLkYCdJCkpqAEf8RF9drwRIaPH6fsA
sHnOHx0JnJ5e+zN7qhECkONStxpOwBWD49n03JxBAY5/oGbED47GsJJh4R0nUrQbSpniz6186Vwb
Jc3ql9QI1eHvOni7cfKSfJCrniUgmvZkNBlO7+V/7TGNPfh6ifCV6F64gM8lFvy3lFXRSf1pFPRr
Rlm+czX8yf1kubtCrJFWXs9C6PW/OirL9DgyvirACymmT+liVjLDzNshG6wvQWQ1gvc8MqVpto4F
QAKBZOrGuXqgkjG8qeNyCCaD225RCsMCL/IGtpaV8E29Ak+skqnjL5nNvzoYmvD7lUfp0sbRLmxH
RnkiyX2kHvo35c7lmYyMjkvrh7fc9fdVg7jTOFy3//MdQD+p5FsjpqOYgLd2E7Qq50xPBqHn/98q
i4PfDUoak8ZkOZEas0CvyYMzmWNzZ1B+RgO1Clk8DoCGkF3Ue1uLOcRY5mm4MrlDWBK9pm2guhPv
9kWwF/bv+lCtWQG9hmX1qtyCHyVq0PbC3na6vUrxVd+AFUSPmcOUw6jkw5a7eAHFPEHxREZKIARl
XP8GN2hPCsREYn9Btvfz0RPmk1p8N++N3LVJDEC/7gP2/Gqudaq9ZhZB/GfyDAIIADJr5uaBb++0
aq2uEdX+iDvpu907xF236mjIX5hkkOQ7Kqw1lWtO06Sq4j6syvdmQtg1zZhuAb4NxQP61jjUE2Hp
4sPjFKegfsxhN+f8F3ZlPSQgGgzs1ZU8LhLbtVVoxoIRXCzz4ATUJmi4CTedKiPIkWfCie9Jj+nD
ixpqRXvGVs0jPQal9ZDMY0DOpNaUft39S/QBKubmCKvy/+jGETd55GGlKrUKkiklaqgljV7Ob9tq
WMXr4hZV/CIIrnc4TXjL2VmCMWpGLo8wj8DLXhEcq8gxFS3Sf0hOGq8IMDLWftESBWa1deyYp79w
TTQb8h9sKkW31xumqt1zCNkA5DyuYkJIFoS6jQ2uxtFDo5VAHBo7PIIGd4rqa8teNTjudcPkPxh8
W97w9h/gU+pmGN33gnWGzUQ+3KbGCWlZIi/Ygps9Ao0MA5TQgyqmnavyd+R+eG8DBAVwChWnJfLN
FrVA2ybryLoSF5Xi1qgDipCp8Vjytj4aPwPl04GA60ar4XTSYx0TaG/Id4cUsGYV67Ic+iNK2EAJ
0WzKQ6YBE2B40Rxtfe8egKS+f8/UfwhOP6T6eR/52FoI1X8y8ADRDRaxu61KqEuNyiTm6dUaLFxK
ANeV1ZnvdutXoZuoAtlk7aASAkDalqV0ETw+8aVtbD290hk4bjK+zmmTOA6b7O/A875BTePw5mN8
jY396VTrkvYs6+PwiM6+eIUdmZ4I9I8XjlfVSIl2RNOoOHMhDmlIDFs/LlEn4GHeMuAQp6b50qXc
lQr45z5OxB5E0/3FydVyHGmQ5wvAGjQBvm6MKXPTyjIGSOFbsxECqc6H8h2TfgSxmWdBZo6IDMEM
0/7Y79eDNhaFfC59EzlQTMtzDR5EyJh5Zc/3A0f/cRpUdwa0XUKf+NIKA57XP7M5Us4rA+DwXoIZ
92pv9wsX0faDrbN+Kwj83uX0OiQJktUYqQ4ljY4YQk3oybkWF+qiYq4qelV0uqz2q818uCugovZO
S0UH54gDU58ABgKUfyxgFctI04kozjvHou4FxqfyB/7MAQE3cICg1VjRwSRyTQj6uTGuNi7mguEh
Y4TQxfZ05JRAVZK7SofHdfjmrUQ9GfrY1TAanaZVViKGMuJkd877OIXHRl20hVwiAGIyx8gTYnHD
J5FW67dThcwSk0mRZpRqhzSGKYGMQ0MZ+/5jYgyjA1WwlzKKExACDHcboRKpGoSCH9McCwEkVM8V
K6uWG1HDWtz/txMqfwik5kNOFsN5OlU0czN1Hb7QVuoE7MzQgaXDxZri0yfRrIGQOv+WYPYB8F/n
8w/kzHUf5MWCw8KdXooUTRnrMDROJZFrJsvHL/DnOmhlsgAB3gxWWXzObkxdcwBRn+qUoo9KJnhP
maVWHc+X4JZbu4UCx8hOjX9RuOB0d+zPzTmWKvc1U9FiBxqe1OASdDKVIypKStiTaqlMW/4P6uBj
gQ/BDnssFlyeJzOybptl4AD/5909v9tN3rRUrUls01q22ge+Vb0lJ6KFfgQephJELQY9TMoeA1rW
xNt/ouLL/6ru6pC8kn2EvAWcgmnwIJUEoo9gQC/jqwWMpRc53LPQIkdm/mtIInCstBrtu/JmdOQs
8kOWPqdoZL7xDPU9Z+lbul+13gep3EWSdMELMvGBkcPI4qlnuc2AwnszpBrCissZRD3/rY3R+lgB
fsTQs5okJ5MeADarUiqOUeDzO5N5eEQ7BegtzaMwLZCuCl/TZqAKK6Dt1+UY5SjiUBQ55iZ+ifoS
yvDZPccPTiHS0C0aaX1fvBMA8gt+HdfoUFXLTHRUBca1uXhNjFz2mnxUi9mkL9iIhtBbrN0sFyMd
roGhBguhMJ+IFTcCVuTZ1JfFqw9DRVgBRWrfiDeR+vKe06xr4XQHMjNju9/w8qnG90evXpTgb0e/
nc4ioq1suuriVJqju5trdrCUadp9rEhL+28v3YmtV0wDLCejr1cLjwBmF1ouJ4dnAJ3r0Ujol8/v
FhfITv9yOYPjQfNJewJXk5DOAUy6TGGLaMJJYUG0aIxdVAzqytwnw0YUNXnKeBFJUEvpiNbkAEpF
xLWfCR6ppvWErYvrJUpIR32AdqumsZoyWZisl73+0NjqYka5h0zT+ojvAakhYvwkPs5C67PFxGMu
4TJkvvBNcdKoJk84NbnaQ12f1oHmqEErHnXCDASuhBQijv2c9/fVtsostZSihqUVmlsCWrxDOr/H
/qWl157BBINQ9QpcmGMefW650ZwIn57z17IV5H8zUA38/vG75rv2vxCgVEuPA24Uc2BUmQonLF11
q7KzLR0dDvp/bAkXMUD4jLcj1WjWqFnZUh+UPmpqQUmxw4mVtVqpQQcOZ/kFaXCuoZI59wXfWRMw
XvsPYNBHOO/sf/PCipRI6FyBxOpUbV/A8ZUledd55X+BtCgSO9XO9V6OTfD1YdXkeG4ziWQ24+UB
bYi3ra+rWljzc9eARETsM1oKwpf++7QGzJX19o0rQkn/zrhQD23O+GH8IAAyXHkdxKohPn63Ai9T
uVybCQqlx6SQbZZHK+x9NrcbZP2BF01P7rbfbnMvSWeiOjxDoqEAQdMBmHFx6XLDwro0kE+dtFEZ
/XsrtVW8HzpUdoma+cq1qYVF77c4ZqQJylQVgK9sppddxFaMCAIGBqx7WokPd8RV+xmbg+ulShJ+
RmaFrNc6SRX5yfab3ZDpcrJegrRVn9JLxRW+YPOHDvzxUb2xpozqrMyYh9vu/7+lMk+Tg0JdEOQ2
JxemLL2NYvrCjNlwQHov86rZHZTnLYAs14IlQf06By27QY3qV2+f1UgwXN4trklP3uQPjZEsxW1P
sgTxYwCP6Pv8Dh478kBfoxI4VKqB0kH0t5w/Cv95q5+a+UPuRl+y+E5uu1rGpjlU6pyIk1NFVgWz
EdIuEpf73wEM+XPlTF6nH1ZpYgJvHfpuKRjGhQkhLTJrjMTYupQAhO1BpjtWmey8lOcca19f9/if
NdiSht5KEF0RvwC4Oook6slGxoICkkoQNlp3CzonOQAyvjELQhZ3Nkngy4QFjpTudMfMiJu6dWN9
uzjZxDW/xPRm9uBsq/FvETXOXUx3pwcjLqOPT0ZN9Gd6ci4+yBbeUrkI6ze2/OYrRQfZvufU17aa
yRtPG8V0N8Tok9deLFaw+d0v/vLZRF2tAXObKG+OxBzJ0EqwN/xsEXKvMs2pLY8UHAfZ4ZxixZI2
G/zXa7FwtNlxDHde4je2vFh6Tc5n/tP7WXtwO+2MGhW2elsdyYhhnuWM9ld3fh7PMVVt9Os0U3hL
zkJ1N/7TH7qTFhaa2w1T5jLOE9/hnt/bbIvin6xtxqlBdKasV3vGPkmyXXQ0bWtWBgz4/cKu1MfV
dBxeoequhVMJGo/YD3vfSv3lpGKPHL88AmaVsC6TypJn/aHuv4WFwqfyjEcgTUE4r/Mq3JvEUyHt
BeFbbWubj5zETsJPut/tfLNqC0MjcA0FPt/tOZaq5D0bMH1HmaaaDm+OkSJVl7//EStzSiyLHCeC
Rgp3IyMEElGeQ96Tp0s122Bhn3x9vTvpd0mJvFqWgyt6m0R5eumK6aEpGeFf55XvMub6ddKCSnI1
EaEVB5vxDGvZyH+wFIdDcYqR4zcZ9TJ+qU+KwaY/YeuzlE8my9SvjjZb2eDlQKQJDlXFmLAqPiwA
QKnaM+bvjOLf/0WnWJWdO4G70s+O6TOGkboNIOqwUys9erEsGxKxCgMIR0oaqE/Hat0/xrMs4IfK
s0zYs6UO+bRr6n2NgCADXvU5Ft8j7Mancd7wfPRfcmFW6AsM0lCgAcj0gffd5kUUJJsZF3dqYpos
etuYDO4ANC3xNcFgN9QkZQ22v/RqHd3YAxfZ53MgQmCZfgXnViS9N38OcU3mmal/wwLgCqphWNuQ
Sf+MWaKuKSPp8DBHOJprNMpp//clQfUjuSuagHyMjM8bI8LijfME8NN5po1woUPtWuDzJFBjvbhe
hpSWFZqc3IBHbC6MeQ/pC0QN4oCW4pwWhXUtPDJOcxfxvJdsGqb9KEYlYhP3T7T8CKXGwc7Ot+0t
P21L6Vc+a3tAjQiWiIYzqeWLsfOjJl0O8NuGf2C5WZzwiLkXzZfJb78Di5JUlcd0zEqJ/fHDKdYm
xlSQYhZEr5laJ16c6r0WDDcKpcgOfZBltH8o0IMqM5IJYm42D9u/f413E6Xn36/+mBSBZUXc6SIk
K1N4dXo+fc3VgC9cCPdHXNsjgRrWzbHnMWjEeqbuuE94rMNBlw5Uk4rteAuYZKfWkdCBCrBXh1s+
zjjaqMZ60XCzJjBCORP4caBgOzDLihIaiyKuRHrjKkk3/+DAiArt5lpnn7kF9YOuJe9nzN+rA0Th
rFmWtZ3u6a/vlAwM+urZiXNG92Ox1aQ9xZ4RmKVT2AwxDC7S4X8xT/gGU6TpDakXdoziisrSi7Hd
OiR/uqIiG9En05Sr34uiz0nafTZ+r7MOHjnki5uVe8UPG8GyEjQr6LkqgnPl438JnVjuWr1/ORoE
qfb8UiiX9puhH4TTTkfMsWCYS71WU6/X338g3SHP7uQAL4y7ywx2rQxJlFbp5OzW8Wyylij7G0MZ
gA+a01ZNlaeGRqu0drBDmofGrROyFNQ5CylacIBt0zShOufN/BfBg7curxqCohkrxPmy/zAalR4t
yJqtk72jsfF3XM2X924NhbxzN89Uc+itk75LRPt3xG1IHs670EKEP1p+BbUZFB1MNC9IYzKFVFLS
bbkMNgmZnXSyVtFYSqc8A4tORZJTVeVW433JIs/x75vZSfwmfFl6OBJPcD6K5YvddpVHoJFQ4ejB
w6gi0NXPIFeUjVQqRatb5yzd3YLjdH28O48oJsOVvXf+1zdeNIuWCS9pHkNyFeKdlyIDqTRWZHn3
nDfN0a89ZX9hh/96o8XFkn83iBYBDYjQxrK/QSRKZPxUhmBxeUh9tHn4TjFBoVCbTUZDKKmMWF08
Zu1UhZf4RxMrq8w1htGelZnU4wXvOKUWSR//fOe73vu6IxEchu++XpLZjVZf7ITkWaSp1DBFkKsQ
E74kd2Qi+g62kBEcAwJhD8KZ/kCX8XVkayIcPDDW3wKAVrXFFZFwoXfFhzZXgtuzcoIPZD6NRFlv
qFfnHhPBFoj99vwQZkIQV22rVtKClfjMwcZ/LcAMWa6NPCMCG1TL13p43G8sGWjruUurDJi6L9NQ
5/jTs3bOvde1IOZAqBetBb28piP/dLzzOKfBE5Z4DhweJ6SvSH9mTdAOISww5u4C3LZ2h7YlAKil
VpaRxOW7h2cE6FIpE2t8hkVUVKhJOcZ8Z8cLcuhvOSwe8hYWM2qfpQB8XMRZUjYJIg+VuUH16Gqe
g1CrTrINYnAjJ252pC19hUpWKvm1HR9fFhWoTd5QMMSsuTstWyovAAT4epJgNqniY17LRjsdAmto
Wu9RY5Rs37MOEcoGg0Pv/HV8UnBO/YlOIZOMSx5JtLCZm3gSvaM4SVSbHjZf+cfg1XulgI75G1K7
GNtLIazLgVF3a66jQTqTXSUL3dqxKLp+MjHWUrEa3vxtNVg5BRnHnUsh2aryWRwGUumHEkRIVqy2
fSZt5jupC8NPTJ39LgyE2DkD8f5fk3hIlxPj5kEUxp6pqM7j7UWNa4cUXS3hka/9G7QZWOYYy527
fTMVlSZrqGEG4O8cGsGUGs4B0QlqEeSzsEK0cZoEKrHVuG9OuRgnXrjhghIiPkiDao4ATt0TTvbF
O4TsDIbxD3W5KnN4QbDIb4nvNKTPqrSVARSM8qfEtirDkC5ATsY1fhmGui1xYkTm4nD5Lzq7itqP
XxKeoDtPePnzru+NBpMuM3vfrud3gV1fzBmqQ87B7fLkRZxnsixeYRC5u3NQyMMdwiURylz7immo
nogDZLnQP6uevqLMF4UnFecsUVtW6F6eSeyEvzf8of0YrbrXfzNXPrMYTs9rPuHRaI9f5RumKm1E
tooR4Gamq7+079MO9mccd6RaMOmnWI72oTbT2D/0xE8SzekhaHkfl0QmP7PBHxH+cj4+EbI4cBUF
Thm7VERssfu2EmKWACxnUgfw5um8K8ZEBGqH/xRmMsRcKw4AnoKdk8yEwlTOHQe24G6TkFAasS3D
C4EtqLQH1sM0c5z9eVDx+cDBUbKMP2dcJCeSCjBWCost9011+D0cXQmbkNs5xS2YlQB/HQ0HmU4v
xU25SjJrG1KQC2rQNW3c51aAOmDa2ibKUb78eTC0rgH32XvqLJMJP3kXH2OpNDcDrWFTK3+RusWR
/svaFgVjR0CXwbtlSCbYEXVHsUgQ7n+B8qGL+pPZGMxJbvDFp5iKSrNApvI13VhlQ2X4uMtle3te
ON3mKb1hz32BLM0OoG95uc2TDGqiDj8Opob6hVWkpJ8o8snW5CLIF+cyjKHxl6INmHAZgD8RfEJf
Zon/AsNqLtnBFDILup+gy2OsU2P+u2n0DOjcZi7hViKXE3GjLbW5S07Zb/+erRHnc/3nnGvGsX05
wLWd1RpU1K8DN/V+U+XE/NBdhzu5k0d5rhlpHB5/CJh/nJSiDgzRrbp+ua6Em01d3PEkmBNFqFY6
57xg/CR0N36B9AJhoHJgbfioJEVCQGM5cIv1QaFaD0KnYJ3IDJjmpJcM9FjPLYmLjf9jfs9sY1ah
i+7OySdyWZ8LdYqi+6ESMo4OPiKet5r/CJcAUOmwLDwL+Tiufux/YCeTJv3rzNBteQEMzMnqr8l0
VZS8qCkshj2YjU03tg0j6YStNTnFl35wAinfBNAM8sU8kDc2CgNkRkDzg+OU94YG3RxQttR7QuRx
JOqbl6WyJNxhTyR9yyNQtdEFb14FXHgLhoExeE1q9pSGF2Mvc4+dHTePQKfKmyQvSIeuJD3saaAo
8Ps3G30hzZlIIA7+9Xe7APO8iu94ckyKqwwMC8mOcH7KjEX23xOWh49+nma+omg4muFL4a38NE4m
niVJ61Fueli5jIkNDq03gZkXZPfEDbrta478h7FlBb/iNYJaydELLkXMreJ2K39Fnf7AMTFTRMHd
hr42dY+S1lJm+XcV0qFg4U8DxSKgY6vRPHT1+wFgvZPdCN3x75geJrxa3rsODVct7FSDvT6wsqdN
0aH5YuoZd+Wcrj4uHXuCzQLAv35HOrTZJ25IXONijN7uZq/3qA+6ubkHPKaAImIgJPvJNyPVppPl
7kBKslr3/kJBC1sevzNT936QKmYnh6tTEe33rPd/0B5uaUoUx7tPv5GKmPodrPzPW+i/BBk3O6sD
o/YntuZKfxoy68EDOyjAT9wpskFWrPN0ucl3N5fvlZalDoMbawy5E7MhZDAfIg4yRlyY/+23W6Oj
2WioISl/geNTC0Icgm8l2aPEnw4ixhUDKH7om58+HYALg9Eknh5Im8PiaanVq9dOrDH2sR6qI9lU
KSoEYBOr6IXQJIygIgRBZheUhi+49UH5n9BxzgUeHXHeZx6AkqaaryotJkYkJcVWIgHrz14xWzFQ
NFgWcM8CLVYhz/J0fRDYgAMIWwSgc5YWSSzTA24rcIpPC/yAEdH5uJxWY/l3TOX1fyGKNJH3Ke/s
faTqltFX+345v8Iw6AUDDXWr3QuK0cqMcTSu4l//wihQZgmRHtVyYSv3+a8hdjEEmPohVnNkNCHB
KuzGIzs4qjD1J+++V6yJGQ4ik2AVQh7VzWS8xX9do24FT5lyCADL+IAwZEOy7eJpQXxgRvLvJGJG
2SedImPozNMWjpZCiIP928ywopkHmkFoNM2ss4kQEf0EjLryIpDPMz5hne2cORISx7zaIg568sTj
h84wnJNx+f6sVNm8rT3yieVYacoZopHz6sSPC6PtxeGs/zh0TIyrTyRXUU/piaf5Y59j4ITpQxB2
4yXsg6lM1IGVH3T9z/d54Li/qWl1oT0wQKKrJarlQ7ZyAR57R4By5JpGLhn6KwfQTc4YwtphdkYd
gPuoeWSKLmOE5v1MFkpCS/GQI732LyZ3SK6e3Ocv1BWGRGKzyzj0faD47ZCHITaSkXDa5lgW6lid
6yY5KZAKhDyy9SqgU+EqtHsrvQr2qmZMxdQMC8Yl5qH7U7nfSoo8JvjXoqfpclyo0a/Ce55D8Ma8
PNtE2eWziiQAGTDkGzOw9BsUqeWCSbU1k1BO6NzBURq0x9iZN/ExyAW7juRYBsdN4IgxdupeZVoF
kHxlkgsn/6zwtxPYLuoYUF4giiUdsoNXusnEeN/jFidIaJUvL9BuErHI32qIjqPtUT94QhIPqfmh
uDC/yuNnRkAYP1JULikmc3UktIP+NtASqqTG+3Xu4FHbJ8QAhkFnBlsqSgC3UzuUAnpoIp+HPK0H
AdFd1vOSu5vn/qBrkfeEgrY3bkMjE6QXKChbJ7xy4Z31qyoe42jb1b8o6eV6klF7HiiMnpC62oks
HMwRisMSFLnHGbUA1cqvKRAhcO4Hi7HlFNTsRFGc9bd8KDegbLV7fkk2DcWXgsNoGSYFPTWzQUEn
u47275TScwnB57nA/UcRtRRX2shNUMY2CYsq1FVICh2xh/mIYc15dOh65godIxV7KtkVIi/dyCuj
CJMmY7AMthIcmGusVAebf3MWY4R4eznCu2BRicloAxW/YmIp6IhtisOmffnRoHumWAYjIqgoIAfZ
TZD33Hi98WjJFtpKN1Fxxi+RSUrehaYztVuaDa4uNLId50M9n+QlBZB+uJHWpcOqQjvbhWcECesF
nwFzTxUfNw29zg6Wairm49MYZlLQBJQtMb78XICtMPc+iIlzL24wfmEBpUqwpOYvOLgKnMVTESO1
mIdeBLcwhTC1nak7GtprfAiRR9Caia4upRJ1rsb5dy4/UYFH/QBl57OTgfMih9/xgiDLdByLMugT
gEKkPwW0LJBva0Fda0/7wABIL14isVEdEPGZe1CXCM9QtNOOeJnE2yEaS06pNlk+pDoK1Ido5OVV
RPAf8hyKORxiiVuO99WMONQjwQ/BBpBdy1sPIMHkNAtAvTj8ODAOm/R+1CfMLsVs5oealcip8j1d
kdjF8CNVvu/++nCLfOkxB6tWx8dgYqFM72Tl7/WDgSBIMJB+xPjLrkHqNlHUt+NEn6Ij5b5BPVNv
4mC17azuD39sflMIuWNyEpweQYOjiBzSUaHaZfRB5jF5VNiy64hVwLNhmsagw7bSUk66z8ycgEzW
HkRx0CnzXCuUlkpSvonrtSv2abL/oePchQ59QFo+ivBPRsL4KXBRoveqYQd3p0lXE+mhAgBUqmJQ
6ckxEfOoYFeoyq1t4t4Rt0/d+HYveRHrT2lk8yTjQdWfSaHxhhA6cTQvAiK3JthUM/UJNVyaFmwG
IrtFLoGpEhEynzy6aMzue/3KeNKVzFuMunsah59KefGjESmQOvIH6LuaGQ8vXEjg/IAxJrnU0lKe
W1Xo5/GKlwbqEDN45SOy23bIAfghYW4HNyXKmCS6qDvKjcvwmFWW7v7MyOze0LYmJwlj5OyuPuUq
br9dUGyM7RS7iREtTrFnWVeuMioJQ7Qesfxwb+EiCKDtLrgV6filh4GFObyHo/W3VkdhjaNqrbep
rfRiR+wAGZcHzol1jGAxgwpbhsQzU2VEFo8/mwGQJJTI7laUCE6YUZPfSjevX1NWYlvo+EHEHufw
sMwgZVwQKwIcBuUUpQLVbrsAa6dFSbUW/SSmJZFYWln8roywSba8DQ6uaShbrO4sUAnhBpOPNsuC
mSOI2PpWIH+UmBO6F7K0c0nqtw9z5ZrZaLg6MJKefxYhalMLQARxnQTvC2Bl40uEMH7dHPSKK7SK
T/DFKptFlIiz1TntROiG87ZpAnPBh8zKJcraL75cxOvKkTOD/tOidd5A8LGrA1L2LAxFlGWL4C9Q
EcXUKLy0T22+6BgZvPbd+yUlLx2g2eHQ5zvoZjaVS3OSzs5+cuRByiIr5KFh1dkUIVoo4rydXgiV
nc5W9T1Hm+9DfuRm22sbnKlXzNfY6m6gOcuBk0lFege2J8IX/jugYoaCz4jvV5Vh88CMd8b9VozA
yPFhM5sCaUtkxceWddpBZYOvV/BLgERC1N+4vRgSCghVWC4yViOa+SpEW/yNNYEFgMnxJdLN+AvP
Xk/A0/u/JFSvNh7QeJMo9KIJ5ebSovDcC6SmRdEIUdu4Irb6/HOWOCMubMczXLnY7F5x7SITie+F
g7R73Su3seAc2qTdbcGhVYqoYBQnvjgnoqA1eLIT9xIUmlYSyZA+bceU+WF0Hq9vL1BtOSPawbtB
SUUplZslS462tfhQPS+nNFCwBUcsQlwnPnnfsKo+02XaPLQ/Eu3LV0L630M7EmPAxFd12Pwxf/aD
GICJju/Tc11OSn9C56xaM1cAAH9s4K4McxU2LIfxF87bWQzVbp7tskHDQROi0pD0eoQQFcgesYvp
VKxLPsPztqNFBGi7EmWnfD5nJ4ZFTm/22hfR67W/gvLNZ056BFHkXU854n1KOXnGFx5GbPtiNas8
qL8c1q194IY2nT3/XZdyahnhsf9k15WZDMNM23WAQrMcMLv5oh/q0PU1TZxLg24TVRWl1Hgal2hC
B8lFeJo+4yEzlyv9e8Y2PfnWoNfT9QoFMt66Q6oILktZjGsNyppTW4Wl2Xm449gWCf1yS2DWvaOV
iYvR1eI/MUn3cmj0ec794pvRu7VRQYlXeJB6Pd3JBFUQ7HxDf5+9zwtSCo5Q9YI8mnthyaizlqsE
5JkzuN8RmEUPbbd8ZtpBHF6DdMHblfvj7q3eJz+Gf91vWy/DUX4LHkI8luDRauC2G+14FQCqnz7W
YHOv0G4yUKHa6Fo6ySSBpS9fOotkUno2c+FxIavBBWYbOZoge6w9P7r7eY/o5qsCJ3PH+Etd4ol8
rcPv2/8muVOtK+fF26goUg/T3fPk2U/adDLxp/7+dFjj84lPOpoDDmH2/dKbv33Uvxq/4LZ9MKgq
p0MrYHxek86KMmWnPuvXvocu7tXcu8xTNPgkMWDSBxvpuHMbLsCXiceJtYRwt69Wm8sZBL4THMT2
MSdWUj9NklijvKNN5KU/3AXa/j+kE46vufKljZv3bV+ixxvh0MjWdw+Sjh0O+7clwdS7b4aiU4Cs
kc07tiM7AleQt2L5dOLp8vG3tCCTEf6omzOTNdusXkPZALGBkUp4U/rHhMiImM8OMIpUgJIjA1/8
iU3lkToCoHd98G5XIvSiskoAu9IpVhq/ivojg2/0Rzd2aFnmHebNFnMcF9vG99F8lDGu8vv4EcyA
Mf/7iPQqlNAGCZXafmmrstSU4lT1GGeLMEUm2t0nzAM0Fhn0byLIym/Op7kjRInJDgMZuICOOSG8
foEdZO+AZhMhgd8koVMfsI/5pQ6rFpSiFNFU5byDQpzHqlMeRY3HcW3MU6xaXZLe/wtkNzHfK/Al
OuEc9yF8gijqPJY6mXvai3AdJ3lFeJJx3bSZ2t4HUj29AC8FIOyT7cH8VHZT5BZeZ4LyauNheGFu
nPNdXKQZTX4GdprV4X7q15iciig6h96TgXBSUIABP5OdyTbgzsedz2qcgYyLr1Ou4AKTu131bnTc
UJ50wQqseUrDNTDcZS+l8+dxIDccA08J33j7xPf4W00dSF8hcw0lwpiyd2rw0WpOUln61x1h3FpA
NXsa6a/2EOPah5MYnIYqWf4M0Tl5y3Qy572ER26lF52GOvMXgep0S2lHdfmkhDmN9/e4FGapcO8k
6ZaMOtkBslG3pEGak8wMQGDz6fV9ifQ5+oUXDtZsg2p5OUvrfZIkW1OhS/7xqt9bS4MNzLAPVhh9
IiVJOll8df+KgckW9zAA6VwxWxmqdltaDrh4esdW7RicFvOsMCfZd3I33MauG78ynKnZUhlzeIdm
xgUbzG84pt/pVW+3k4fR6Udaf0e0RQKrFlJTm01AungzjJNZhIHHOWaUm/yc8Ea0c/dWdmSgFdC9
TAsbtzel7yY6qd8gvLBTWhflC1g2Ai9eXVGJdmjUD31cd0LcSMuMgggbM/p17uCsLWuSjlYmR3GL
nKd2lC2BL+fOon2G1SLlh+Kke3eAewbwrj7ZeMYORqA8kMBV75LI2GTTMUVVq+iqAMDeZy3+LHDN
vGH68yvv0GpPSqtpBhtzwLe5V8ff1x56k6udw4ARffID9XxbJVhA+PywDede6f9Bs/QSrzLtczuT
GRPCgzw2P/JazgRDsURi9seCPZoysDdxcv201rFRFV9aTBpA0gEPEqwAEAHran3tHbY1Q8w0Nj9j
XxWRnwoA4TRD+cXbfeN+axilgp2kri4H6ydgWghJ1OoOQUDJDX2aIBmXQasbbn400YCmtgizlnfn
rLfVUrwYE11BOUcFgu6Lz2Man+FJwNCeWVGJqOA2odgeaVnAvhBKMUdKeVmu0ydada5n0JRUGa1X
535xD4zOzbei7ommA2gU058pKAN1OfO/2IJ6s21C+tRNoIJlpOm2QwOMYQvZNqnOFySVajBHaHKE
AX1+87RclMn7WwZkEyn0AHmB9BPL01D7pc5LQW6JZiUMKW4s4O6Ksr7VJlxBmC+qZzxS+b5nHF1f
BhZmpGk7UqonSqGM1goMfF8pzj3S61FwTygoByA1NChqsDP91y7t0/3IbnVpkBRhRoJrIZTLhjLz
bK5jK2ax2gxhakAWkWMzQTARwZIQZL6J8BdXfFpOAzj7QrUDhiidH9Hmb/UGjcvJXYySCqlO/DXN
zlSWZLFd+OP34GRBaJyeLwYn7TuDdgOLJ2eQIv3Aj8c2tA7cr8uKIJs6CktRZe0frk777cmtRilq
3lMuJdOvXSm83W8UC4aV9E7KgzET0IvNCg7c0UGbsOfZTfta67FgD6UfPjD+5FE0uZdXR5jBoQj/
+CD17vsmGQqmcuihMETuz3IOjW8caklAYc6H4V1UEG8Kiza97HtWtT53PE8pFc8VSy1eFoYjMedS
JcBvp+yePvtVuE8W7a+TIrNtvAZIkvlejkVWBd3qrgdwQs5i7ZUTo7EgoIxXnniHGzsOz9wqz3TJ
vIqnA+0NafZWQFphwNjvMRq0Glbk8bSJI0Q5c2mM8QJYjmJBLSAM1bGj6muA4eltNgRon7ORlSTC
Mkuks2P38cw/0A4wiH8WDT0Od0lYrG1Y60Z3a84P/G+0yMXjxGgfM+deUPjRe0sUDt+HRloYhxNl
Xx6DAhDISmKzfanMOqY6YBmgGp5GvCVyUBZUA5b0Ligxj35GZYz8XqTiVY2rpvRX2fDTEThjjocB
EEPsuX4LfDxHG6PlyI/ixmDBVt2dqLQ658XeZOSCZx1GC53XrwKHsAiWoSEwHpzNPrOmVZCoM16f
DPe12HbeXQfrXt+PmnxZ2UHAW/pm0gMZ5U2XVF1wCoqFUR7zCW2yASPRCXQUhB7MwRMTDaaHrEKz
feVZOjBbGr454JtczhMw7+AG89R7oHyeoB6IyoNVnKm659BlyXWclsXJjljp24SKjURbyUc0/3Ck
oBDm0uhhGovOYPJN7uhH9pOuQVav8ZLGTyvkp8rHJ7s9A0jhcg/iNIYrxJmwOgBQaoZD84OdRd1E
lbA3PchlpSPHHYPi02QZFyWm2HOYal0/Og6wwo4lKW74o4VJt+fVK6PqOIL6QMaDfj7FXdudhM/C
B13IYbRtxNgfattjGn4czV0epzsYHFwgV7UqpDkWoqbfnHG7QPguxIXyExPty9bj4Lkol/DAZiua
HFYOOVA8uAFMMsRVnviWZdPh9tmUN3QjI4GfsKL7FDykAlb5V9dth25cZPoUBCagHAakx1YFfpaF
XErB52onW2lS8FYrOknyq2R6I0DYka+kAZwtK7BKZE8XbyW1Iepo4YJ6yiT5N7elKVUhzPqE1i26
htqzbU2aML+lyqwPiLuNRJMvg3eoqr3gy9+Y8GbC3EW/OJtVH0H0FDnbkVZtYLcg/D9fAViW31yf
g2ssuk/GoAeLeApTFfjE+R3qgJpVyqR6VxZW1cnG2Ip8DIAsh4HuOR+C2upHWcngu4gdrsvLYiTh
tzYjMXp11De+f7wWkV8x/CNVCWEygUtylm8RNTM9PP8j/ZobHd1D2Q9vsH6pWAh+wbfIS0ke1cr+
CkMDGdFl1UCMuG0oSNyMKIGDyLmztO4ghnexSsf8EDbEVbVPhVj4ukoqLYY8EYazxsZaYU/R/ey9
V5rMwAyYsnGUHUnUj3VQGJdXjxZWdje96Uax4BvWjU/bEVSNi7ujql28DECedot8KUkpGu2hIPt0
aCvrONjcxFefeUckCJyraUg33yBo5PxMmlMUWP4MP4K2AVtIBlvptHdGYtMdNS9/hcKRYCf9PQRU
TYxXfRTc+syZMbJyRJOEVe4rJKOEdD33ygixBSAm/nAJ+Wr+L5y2jj1UUi/+DXV7J4NaAUBm3Fbh
1XDKHbRJJpgKeWfZs+UEDx2UYZoFKuRAPUW3Fw3xUys60Y7QU7P2wqtohr9CqOmKwqL/PY8HgW70
YX/LQ7jeV2Xe+PWezmK9T0EyCxcZdu1EPLS5ZaNwcFBakjh9RyQACuuuBZZd6BOuWPwk3/rBpV8K
8aw7jCujiw5TCvUYU7e56YUGalQM6crIPCYWbkt9aVZCFaHTCkC6UrLoRd9NwGUkGJAPqmWg1CZU
tVPX5B+8XVzeh9pinQfN/YgTzpeVS3hzW7fRFcuK7TCQIP3JxUlZR40kMmH2pzJAihG53bq52o04
hAHuiCOEhSm892D23M2AAou+sNsK34W738+17SWdYyotMcwgybx1h0irFb/PkdY8/NKQLY8t5+Yn
JRDepq/XOXD/Vk3ac/TDapyRf0cl5XwnhrCMA2Zrvtfm7WetgHvfbBiHWN6k+wjOi2FMX8Fw1L1G
Hdu+odjLoQgUii+EmCOt88IWoqYmOwbWc5apBb5ekLVKwk2UIWLLRPbNqMBhmu37vU4vThi7Ohhr
WSNBL7o54MAAIxXb9xO9UntFl06JqeItgKdiP98E91XqhLLDNpDucDCbT9NZtvzPyVBhVg5nRwQJ
8jiSaMr88SDJB32KYWlyUxc4iWlTptnCazBxDstBCj4nfLpKSBa5j2lfFlC8Bkxr2sJH7T/4XwPN
oyTjmIfpJnFk+cwvS9WdxRfLIy6p/WoqOodl3X0RlnCMlPx/DNy41h5/GoS1qZ0psc2aLWNBMN8Z
D6PlqiSrS48VJPfJ2e1kF9vlvXge2rhRw7lLZBSGdXxR6E/ug34TttfCU0EiCf6Q8uwvKish83Ga
DCuM7BULeeamCpoUXdkCOW7z79zqILMzgyRqUpLusah2qALYX7RRMPyZJAAUseMMO30ug5NNy2Rt
9fG4xtqPpy45lbSsy/RGQf/CnSscFgM7faHy8Y5564SNtvMJ51QFDgw7piMfHmVqdIwIKFtCK7u5
VB1cp4BlOSxmYX3/flZT+VDeITs1CmR/gni0/Eg5gxKBui/d2QeqoT7SfrlYjUnWDXzvz8sZMvSV
YEFvy/86V2itAvPV+80dowKGXu0/3TeBOqUgXfkp7btV8SVw+24Vwte/Uj4cqmaaDRnVJbTNxSEc
Z2wjIxZ5u4aONGSCFvqAjK+9L218QlL2w6C1HUUvfTnhjvlDzDJTc+PGR6pvImqk5//4x3XYNO8U
oQJuplnhAp4x41Ua6HLAV0JEtF/+7AiIYssZSmCtd4r8j3WpdcZ8rU3heQsl+e4dWLogFUtLCnsj
4YVvT7a0DnmCBX9DoJTgygfxOO145Wt1tgWWpKbgPeo3Cm2/kZ3a2wkmfvoZJ0k+or/BDhxOnFzK
8KgfK8vwjuQqyPvWUQQeqVNcQvHgSZziyGrMSgj4AzBK5J+oo4duHn69SwZAKPaRKid3TyertpDW
4kunkBYmvOCLlyQfW4qcs1Nt+TGwmWSlX+kCam0oxpCDblEAzov49ix8XkJu4G9lLyBn1eyL3XlA
C95unysj+UmK0J562BaZ4fA5gzelvb3If5PZwXxl/9cOloeuYC/9WNvhH0OhMyROAMAiYD2LHcny
+Q+gQYwxdXmTqcSizl2bBmMPmg8SpjCg2G4BDaKDwmYKO4FcQwnKUJsac41ubDqmsIs9KHmgXAqb
FGx0nSoC/2ao2DXHt4+6WJpQyjOFtgSqrad5bIm0u8P6RFgFU8CfzSy0sJzFq8G3pNZPqw6u5opS
OK4Kgf1+EwWeQae3qAUZ00/z1MmqHdnLmg94aJxTwRvWLTnfTkn4gcMfAwBjGL+NaXiIKIpaH7jo
RLpRboS1ozUi7V9vxFtyzBV+t7SuTsjJHyBcuD0YmmVFyL8zxSXvikCo1r0aOPbFuu2OOrxRSz6g
UhjEimhqNQCYV/RXaeE9xmsH4EhIk+vYWcchuB83tvWfhaVBtap/oF3cIwN7H9gYITlwcKNyE+tT
KyNTAA563ASnmiH24bSoFIpT+A1JAUshOOqJ2f0KEXbVqZm3qmMzau7p5TWzx+/fzPu+aT81DAdN
L1XQarinG517BTjIAKYIe6fY7YGC+4FN/LOdc6PG1eBt6gnzYpz1YN+IDLwDyGxezLzCvObwUnCH
XlfNBHyQQvT4Ude/ht9h5KTa4yw1rf8PImmivgxRv0AhrrIl+LPuPRA+iTLSc3lQBDeWX9SyYooU
7QkkdGE1DV3xTvqTW/ShJpfbgnjbtutC4nbcJ+iAeAuOSYA8L0Kp3eUlYyZUc0OSNd8zN/Qz1G13
tbmqCt/mZxHyzl/nhxfomsoZxy4wnE0etU90Sno4Pb4HG17cCGtPOr6RoPfoiJo8bOCCXlQ5nR5f
ECX7piojVPpptPfdu7pC2h/taGmHogLs/atzQvrd8qvu6HeZIe0H2Lu3EPX4wLEOQ3oRBWOICm8S
G6/hq/UN1mFsWIYsw3pXmgOCLiync/d18y9knW2WoXKntsBcxTH4MNHmCWQUbl6itzd044ShFni3
PPmKKKzt31nlbRc8Dg1dOjuXOHxGsT/ErBD0L2RLINUUUcfn/meaTFkXGikQLw41Fl/Hal/+WWiR
S5A5RpVQM3ZfvJA7Kw9yGozV9yOvkNvy++SVIZb0DIRYkBZFLzgmyjNqYDpFDdpDcf0DQGU56FIp
3bJS/yQZmABrFt+HbJhwnqJWXqimXBeKUMwvk6qQzaPYpBbBNmy2WyePdq8eOFa7jBvDSV4/dumF
AcHU8OaS8z6lI8E7zfPcXG5MY/b5EUDHEh/G12hzSm5wbOimb1zaCF3T4kaDEZPEDO5GW+leM6KG
2UcCtEV+NFVhZ5Nyl4dQu+Makp7xoEUsTvcj+yvlnmM7vCnauP3FSMDTaU3SDpxintBXuQE5ndOd
w7WNje0Orr+oqfQyDBTPjUJhmdf4CfECAKBhs5h/nFxJ7LVgnKqieSNB6Knfdcj51Vlfj/gwSLt9
tann0f23hxeIC0bbDECX8GRWcO7Rvr8uOtuALLbgth7tYur76A7PP1p/T6B2IR5kZmVzAB76D5mb
1i4+CWW1NJRT8yXRgp+EiTci2acQ06SpPdoPd2L/7eglIfGuK3Fn6WLIu9A+ZEhqB+K9Z8MmZjJS
rZiJ7DBbgz42SQpsFYz96TLWL65CnRRFcvVjoayqfmYMI/t5KqnIx5/GuWOJqakHy6ShYnTknhHh
fkHWIrXXnZ5lcs3Wjat7HJWD2zh+59geprj1E9BmUFpBrK1FPAeXpUMsQ3jZGhSkbUIJmYe4DkPP
mV99qev9pQ+qxUEBIWR/lishXWcoyoC72D3NCKuPUj3l+HVxPwY8Da+EdkKW+0acqDDWJdErLKOT
mNLZTVE6rgtY5WvTDbgT77DQkqHEhxWfPmZFBLD8mb5h/RS8g57IxRpmQzlSiDAWc3wsSDDgkBSN
BOnpIp42qH8L0mEBorJ+2dZbzUuLWwZefpgjAo+b1aMVO/irdY+OHjPPtTyyT4ecI5wdXcs14Ijm
yaAbXZIo+0PC3hio95ASHRnodCwGhGTE+akomoeomiuY0WHwON8kCSVwQNgW8v+MNYRobE9m8wyH
oyljVQQ6i/sYZigxfVlb1PqxgJcxdh73FvIk5gsxmsWJo12smTbm+ECCqFHkGsfrsMFNbn0PJm2F
4Q/KljG6T/l468m4MYK6mnj2L9W597C/qF/jr80RGMQNArjyNAVtyEhsaabbb5wBa6aPsz0rPVWO
5FR8DWcnGXRAUBZF0DctKil+rR92kti6e1pft0JQjMAjJM8XG+SmnFOli/C+G0V1p9xYv1kq/UcD
d/PsHSj9u8Du9mSU19h7MpgI5Vz4yvye7e4M16eVNKmBhcov+pIa3xuecsSDF581sxzRut+bnC0J
DRJuDIkwVxqdzeuDBYU1+BotY/8VJBEeZsCvuXsoocmBxBTbwWtC2w0AWwNRA+hEdB5iVNjn0I+E
2l//lBw78NHun3pIw1A9Ule8KWjR2ZQlNeeGuF7bMUuZIVxb/AcOZnt6HkTFbqLfmCTamIUltknx
PCmxEDDNXuMRGEdunR8+bHjNvgmOStezU+8vQfvZLugxUkymLhge9hwFdCbFtV81V+ac3kQekBVd
v7988I0I/LNiECuuaD1ToVxInUhVUBGh0kvxy/pCCQKeyeqHLAbqQx9zWZsz3yhkEUNCel53P9Eg
istANNg9cCpPo1ahbP9sFgm+GJnR7vBKvVwovtoM4TBclxhkAD8YT/3ZwN5XfxGjwm+fSfG4U+bo
CwQ430aplVabQlZyNyuuHc2EfHS4chNbU6B/bFD7cJLgcwZbKnp1u+StalpMwuySI/3//LUxksJb
00E1KsNfBvmEd7UmidPAknShxmA1N1cxpYQtvTboaVm8Lk04fusf8GECKObzhilc3VDq2t5D4MLd
RsOML6EePmxr3lfxWGI2PGG8kpW3jikuV/Rhc1QZADzlymdk2qFFMGtrKHA9s9s51ULFFddn4mk+
BpMMj4DyIDA8ovGOtsqNyMPPrpcWLLCdzsgxs3+m4AIp/LcjrNwHkbRcww5L53YR+vAwaore+eU7
FiVd4VNfn62CHHAhyAmqRXJlwuCOX7UYOSeU7t12XYPQugL1tBFlvMsOrx4gfzJJo6p0uAspqD9E
51CGQ+KgHsyleSs6yUEVlaUjdp2RDefFy9/l88pZfBFfTZ3FqJt/9+7h3v9MX7tarf1EVAsoaIOw
NosOyoBsInt0X2ml/dejMmzOquTXJQa2IBMmro57H9gGWY0qJ21fHUccgu188Z6KhHS0ke4z+GG4
y3oUi7m6JCK+745pjaQ3pPe0BfN5TjhJxDpXI554SuZmeUP9xtVkXsceC07z8s8h+qbYgoF8zuSb
5uyVp/Nppulj0fQPhrAuUMQPyjVW7+FLanU9hLk2Zs0gfahB8nNFc+6jNluAzwiNfSypZ9LhUvoo
fXAZdnAZJ3FY0Q8iZMmTYCec8uWL7L7shlsyaJgiT0IVkeStaCyAxJy7qI63y+8ij4X7foOjsvnM
YHfFH3cxe42OxMaW40IcCip3ffb5FhO4+Pcm9wbXsDFyyJ2hF9irohBPatWmnRBLa7aIvnsqqKhY
erXO7syMRcV32NyZA2V4Pym3d9PvvmATCy22F+vdjBtPyBdTBq/NcmWOCEbmlXATszcsDYTpExt3
ao7ngMX7jyDIhWWvgIAjNBh9Ieu/OFtGiU7cFXMLJd3owFOqsiCbSEHe4xexu+N0OvfaJ0uP4ecy
uSxabZj5+K0vkaHae0wyZPkFaQA1FIiPwVXJ4McMm5wj6ucfRnzvjQEPYn3XG72d+lEd+iCuaZZD
lgAltqCNXDfSyl30n0vZ76Jm2R20e98O7H32LgvLIfl15RtLZo66LfV8ZTPbDOruqeFoy28cXPH3
dUU0aoyq4gMcgWM2ClfC3Blg0qe8f0QfSzeBarwsIWNaUA6Y6tIuY856ceXTs7MZufSUmyBIuu9O
qVmihCVy2n+lyciq9nU6vbo/suo1AaYn39wNvVV2LbS1ePXtDrmSfpbCo6LTOcj9lYAsfVtlkR42
NpgNTkEm90bB1Reim94j8e5NaOH3huqp5UQcf69ap3FA580KYEWs0+jZ0jeQNkmfVvk11IeIZ67s
M6N1coi6y4MrA9SvSd961m4IJWI2HtHAKYID7jg51OjFtJA2AgWFDVygXKgTgUdQiG2PmdqSz19h
pM4zSpLuN6PdCx3ANvLTFQ/T/NWDD68lKWDvjEFNQ0fIhhLZh/LrFsX9tKrXQJA6y3D1KLKaT99R
Bx1E75AWtUPqzevBVndbIxW8fsQaBrE9pRGsLGDQjRKlkl+OlJ3dSxEu2mXWNPPSy1fM119Gfbpl
2xzNUoF+fRaGlOvkkuH57XlHyAJityj1dkXVqLNF8ziES1/RX6YYS0wIJ+X52I5UN94iVR+COpl0
I8K/X1p7kY//QvrCHtBeCQssQNjj7Dhu76BUhQyg4C2uHJF1s/OX8Epd16tShJ4bul7sJs22BXCM
Jfg97SlL/nYWWnOkEbw90e2cojT8qNXkrqVtR4YSXrt1yNutqhsLkz3+qnOKh/a64OVrPBqZiwJn
aH/X9z8Qu31cdm9XfLWIwxLYho5fOCshGqMrkMl0sFfHBqYMcddKLG8cgzXFQ5JiOkgxksDbIz6Z
1Ie3sBn4SyX9NyDdPIxhG2SnKGV9LrnTpXKOl2WRhtC2h65FBcGyNV1yd7YT+HqEZXfMGJ6/pxN3
aBxNz0m9Rb3MMoKHvqolbrsoPe/EMgxfxQP15pEPUmEle5s2b4sJB/I2sDtUpCiUwq5RFWd2Vkir
W0N6nOA5y/al1JkyUeqoA2wT09O+x5CVvioSTwReN0ZVQqNJK7JLa03ixSljHu8LSN9gRTQsM/qn
/R3j4gDtjEFltXEr1OPMyscN/1whJvpG7pRQH1FSf3FUU9YNbrK4Xc78QojOlfO4DpAKgvkLz/SD
Nqba+n06Qu9qHmN2MzdQvbpNYhrVx9aaps+BaLw9v/ne1Iz7C2xidx27waQuLpYlDGHKMYUSoKai
1kv1VpvKsDmcNuMDCVbGibExzP0NMGlfyWgJ7Zp27hcdJNhFH5ZXPQKX9LhXL5P1QZLGgWje5RCv
50qHp17TpIG4hqPxbRdMR1zQ4y0qc4AOD3UJf2MFcqAFswE8ib/PlwT1ky7riguL8/gdrNM37Vma
oxAXYefG5+0TjZLbdw/k/DX+Tunrh5M29a93qxBDq1P3MCJMK1Rwi3ztAeZjxHrN0eu33jwYGiGh
2udUEwlmleq7ia6p9xqs3ps83WcTc+A43YSnjBjbDZyS5QrDJMc/8oSL5iZUohiIzbkwP/6rOhy6
w59Z2okQUYZI8xKxYSxG4VaB2XabUQh8S4eCWq2wA8xSwHLxqNqCGhfJBBVhSGXpoDTPG0CsUQzE
v2+j1EMP4c9DFFS1Iy2vfwZrq3DLcgezdofHIQZahBFiaRY7D9ADJ1zpPMIfJTqhHTWmPu69f2t6
5M/yWCFHEWRbJtgVRAumrNL/Kc5mIROmROg2ZyIXD3OO0YAh7xOLXKCUp/TuGyEuxK8ZHtaCt0II
4PywCfMZ22Q+illFc/gzqpi0F9e5c/hsUv7hu91KvsWMofrAsi5LI1/+wACEjmHelnVsde+44/hI
vaXa3Pj03gYjyKckXGurySsc6xBZpl4rUJkJiKHjg/ZqgGMv1bIsHQbj661bQSTF0Fa6dEP5AhZN
fPzLACL2AcgPxVey12gfOaQgYHX1k8t2ne5mtzaaDM41fiEuZBZYmcsLOnVYtz5hILnDgAtN2p3J
bm5z55AaMncK6jMAb1ZnDUTEkyYjD/2DowuwGfluqJbWS/aSVseBGTaOYhmoFh6vo+Ys7SG9VqnL
m8WFKabeipddvcvQArGrqC+xWn+eHhq1zpr8gds42JqjXDsC8ZKT97zhLNHbu5IyyyhzgbkXGZOY
dZpNeR6deNfQLvVKGvbjKPLJyHzAolgas3MzUqaynaJ+G69SB984obrMrnw2ZtnMTno0zbsHm2tP
j1S1Ez9F/HtOpMQRa5m0LI7/ncZQM3K++ndaQD4Jlt1rEPGN1eB2/I41Gy0Guyvl86aU4mhfxboS
RGpP4OmKDDkveFFmhgD+avQeEIIuXci7qTDZjZGYeaSAFXNyELZMsa6ybIK0yFkYLSvbFQB3zUzY
tzKEqdmLmHAxf+vzo+jFtOuWaI0sWnN5kkcz4Q6YxBmBNjsfPPbjj+H637t+cdOhiKvThKWekCj/
ft43wTxvsnm+02SRuRdHORBu8Iv4MicpBeKCVoQAEmspy5XOh+l718omuhdPlolnU3K6Y/5ZTrOl
ARYZOOgBrlaIJXqyBCeZHymRbH1QFoHi7rf73/Rkylx9yxs3K6ulT4sRRRrEULNin6vEmaUIB+UF
KXB+FRP92/C4Wc1SEi8a+D7t44WEmdM0jKZcHbhtO2R/07fPHv5hNCQFzGQzJy8GdyIOhU+IfS8g
oSVh3oPqtYyieJhoquWNSeDBWF8rITbbf3QhDmVoqDeZMQLCNA2fHPlJpFxu95YuDyJmrOYSHYEK
9P6Md4sWS5FVSuHWu8p4VQzioyMz0RS3lyOYkzMKBoyZYmVQH/Vj8JMy4F5eN9mBOsJM3QnYUrzX
6LJzN5nIqE1OiOTm88Jq6bXT9skPBZDfKoGlvoVToWzjbLNKRexa4UuDjGOCTcbR+Ho4eH3Dz1rc
wQZ4Z3VbtKQNz2sAX7fsB++a4omvNhyVSKcoqPreH7Q548izPjCGgejuarWRnIkWDlaec9WrUsB2
teHtypa4lhpBLKVTmVrnoSnj/0Z7hsUBvDys3OuqEKueK1I5ofOTBQq0uaC7ZJlW4GtAPGaLRACT
viBnJmzEvCeYYwVt2Pxy+9uUUjcyiS0ncu5EtWYngsBLZLtTXpA/D6j4zqL6otNBatTx+VYTKos7
b01SiKu9bk7DbUzgjKIvDoe/UxLTt7L4garotOA0yxLcjg/QZ/24BSAkI7WepoFgujy3PKM18rgT
PP90bkpKkcXcztKyywIT5GikXSbpyQEyjtKHBOSRyRNSW5g2kQmo2M0NEvsWVgqAKx0ZojTBhakg
gJ5FkVSs8Kl/WfBQtr8MssUGHYsXNn0geezz1lHThB+TbhUfL6FL31SuIChahYugr3yvuee3/JaV
lJwXPco7F3DUhlnZPP6lasiOJC1ljEx3v7EHZ8135k9cAyEBp8OfkHowJIs18KuWvBaLrgZ+wAWE
aPnLuVazuhOma37+sTsRSUotEDSYYuHwSuj3QnVyZuFjRoSxZLROXib/YwmrLrsvPlATrl+Mz64o
D0ArcqTowSERQPyUFAOTvaVKlBMYO8hoCPArP3+SDQKqh7C5W9CeDO9fjxa8dcPFF8oVM1BzgybU
gpNkZLqffSOKqHr6z0aAq9fUPLeaEidu0cZpYeHkThslZnltjGEW7v3YZrEWpgSr5y37CPXi08nM
4rR9wsFYtAsz5JB9Re5Bq0G9yEFRDBMkAS5Y/c004AC3Q4NpeOMNnlcmaxbdXgFbKbVcvwYdTozF
CxeuL7m3siau6fJi56BezqmDOFblpg9y1baLICRIxo3xCJzvPK7B6hqLvIDI2BYBre9ydeGy14l1
JDBq+LLr/pUcGi3t+2G7rhdLParQGoyuIE50ePIQYIcaILGwwlStOqlV9L41JGgLDtqnxDSO8/OG
shWlqQ4LqVJf3/uB0LhmzzaMTupouCg73maektzD72AH8t+rCjH6NZRBXeumpdBBQ5aiAe6BzizY
Y1U5OTK//SUxOVz3mFtnG3MNLOcyWAvD79+f+SXikDMsWkeSGiTYT51OI5qzedgTJQEjIeNjYNgp
Bl+KQmHD4Ge0cvJpAVpth7sC/ud7zUNFf0+W/Lbqfc5Xoe+dGM/zTRjDRO7YuurecLNaVfg492+w
rk53xb1z8gsPpaITmbcZm3dz7qSfm60A10AQGH2zuhRkaJa1ERQ71GNqD7HkaVApwIES/x/RkOME
KrGWLsDf6DhOGJIvAj+YwX0x5HYspzDyvCDITWI4+B4WLZwUHB/649F+xhmkVnIADqcbYotvjKyU
mmCabiA4WDxwhT5ZVcorgcDlgcgJr/mgPDVJzyDT21BpHZhYa7UcYKI+5LV4ehyXtWA+hw43O4pA
lrT5WwiBoW3ebyuMMHzgnniQB0DF//J4tlt3gsI4KNH4/IRcsMY0yGG+s5ggriPQjaaceAyjgTUr
wm4zRgQtNJtqGu8/yRpF1InRUE3Qu5Xk0j+9nf5jJojvCJHO+LbSiPzUo5aSd0he09rgZyixRrVk
Br9cLKqdn7Ob5S+WlIk3F4iVrm+oW6Ri2M+7hxnOYxxRZB8/gfW+AKOxGTRbyk5FPhELmqNZL0Pa
1XggUsHuI4bdOXbepqwtOvQu5Gnu2nwKqfW3b9DJdyFyzkZPwRVZaSls/6HQpTe80gA9AXTn7cXM
wyAECKtWlxErtm9XogK5Is/SKNtuylm8ViukbxB62oaIeMM5c6Gkg3ZlkH0TnFAcH/6KZ9PwctIj
3UHBdCE+mvY4c7ISaMM3gBcDFona8xbQL+mBqL7amnG6dDpX8cWlOA2u6zvRVWCugD6U08yZ8uPP
kw+hh3Y/ZtIbR7Td7Erp7VBlhECTsmE4dxnM3nHofuKGeQ7GQcUZn6VzBglNcZSdOmhTcGgKyNhN
a8UZlOQTCL8gHH37/SKIldfQcAirDV1WFqtBz0tO34tpbTrDELKb4pp0HF3vwQKCK6i91MtjsWN6
M/0G2pdX2KeyZNWEiprnBEBqfnr87p/OfLLxjxI8xx125KdvKwQrECJDUfoVMflcp3FooMaDlsUs
Im9oqYbwDQA5GGK/u++QqwF4KBWjk9PFN/aQ3ewvQS+Px2Fl4xOFbFtiiO6phUWaMDq7m7BVeaEs
ca5/vzsv8w0yOhySYsTVl2C3dNQzaLhwwbbJMUog0jdHp6aKLlNBV1X9yMHcnpx91G1Q82jkvuz7
7qfuSwKe1NDWsD79y5qP1GBfeVQgzqluLME7FesWGXZCdIGFP4LLQHy4l2SGwLp3kq8yGuSx6EBO
QSW6N3LRQjNOX2Am/nopG4Sa++s69PFdn+KWOeGvEgGhsuyAXWDJuui4CGrrTmRfrILsOm1/5wWc
Hexjv3570sU0Eo0iDHszTspEYN76R9N97eIWXM+1ltrJaBYT5hY8mriesZkr049kMykFuCPNJnYe
qKF+o+HchMHcKfPKxafbgddmkjcggN+5/p9ApbcU8+shgkPdbD9rHRe3j1NgmUMZqgpL4HVXKwi0
VyMDbbLhtAYgPNusUri81zR1dXfmYlthW/QqqI/FtaokSByAUMv2MUuBGWE1rwXLpnWIuBZ6SC3m
R0oUvuBW/7M8Ap/jWxXgOIp1XTMEQqTU5MVAYA2Ot7G1AF5/29jwvVsUC83yOvsHfjIbNsJzNbl/
48RAbmFNs3FGqAixCTzUGbAt3ccmkcnP9lUhqSasbvjBub636eSDTjewco90WHPEAFaPhqKXhW73
iSmCQtRBPDx/1zGFOMuDDYg7XYUcQepe4gpDD5rF0EOVU6d2m7RD4UGOCqQCpSmmU1Ytjfh74wbI
k02jWQJfyD+YkxEetMjw3uXMIvoLq9uCqn8om1CFkJmJ0+L+D14mCDxmTtm8DjnvHvTX4W6SwVrd
C2miiu541Gl+btV65ENreuH7BM089TKYm5E0Rf1Sc36uOax48S22YDnHyiVqtdU/xnA5irr0HHxD
OF7tMAnax9pq2on3tZwW0PN+ZfGaE0bnAtInKBH/8NC8pS+X31uoZqKuVHnuDuapVgR5woeH3/38
9LHvVLeiMXwSFesBS/3aF+uT24Rfcw3nYiBAP3oBSIhSBbmKhluTEFp4kPObcHmm35mSv9elGuAi
trYlX/crAIRiOsjUTH2lmt4eNEJn8rnEqsJ4/d6SjeUsZnw2t7StLq1+adFbS0uoYL59uBQZoHR0
QIEiufShpYuLx0qoInJyu1BuNw8a4KUotMcUC1eiOYDfGdSzuR/6RMiMl4Hu7roJqdsk03JKmTPh
g+zcuGGeelygts8ZUQ5/1vE/j5Rg46WgLVcUZeExWCkm7c1fZY2vs8fR0NgSN1mYqIHUxEcOea+y
zWjIR6GS42ZpdKVwfA6zBjPfQTGn/JBVnIsKv7jgBgdbhwzdD/3fJ0xlXMa28dvJkJdCTWFVkA9P
hrtyyRqxpdKIQ/qC84QpsUB8c24jqVf0H+egUOXnzIzT/f8qRE3pz+Vg/JATT5diQp9M4MX+x+uU
B8JQziXOO9x3hBj/87IJP4OAIR8nan7tDAHveR6g2j9p75wjdKOBplfM95aqhyxUFF1IpVVzWo1u
zVutuqtF9tE6P+9rwdleWc4Dsgi+w736Kq4l2z/tbprarpd4l66tFLs0DqyVxhJxAtJ/A4g8vJhb
n5yzDuqQveYd8vqYqlnDkO5eAl7Eiv8FF0BmoLX+0HXdmjCf6A41OUgVc44rvjhTBxZe5EB2sT76
Vgu4MC2QW9YFhddMLkl0gLm9/i5B4nPdV/1w1Cylvw70j321C9+TPUp3/lgWi+rm++p5cb1CkqS/
haj7qecG293NSwUxoYWQx5tQ31lxGUENhm6WK08umEtRTFfrr9fKIloQbaH57HWCSchBpbfYTVk2
ur6eS4vacwKp+SQqojxWdZw05EW7zZZYZSWjwOdSEle4hGwnYM3uyXhaF0H2wT0nLovslm0zzq3b
P2gSzKKT8lEmwzhWUgNXdSMmzUj9yc138iqcTQGvcR8LfvqNmbCWPO8E7rKeu2q+HMRPnk7uZCoy
1Si2uEVjBrkYRta76oGAaKiITa5eHUTHCU6WOdgTpEjVpiCaN75+4no7/cJHnKXXeBFJ7H44ff/Z
fddNVN6WMGInYNeXf7ecdTEUo7teV0MvxsEwYeZIYQdIFBZk9dKY9WPTXZQXXoEiCZ6sHeXYuFHp
bUm1W5uctYsXQvYhqZjm6BdRgNxamwaqHLQbxpNr585DyWc8GIuU4Cnh88CCCQic9JKDvNToUiOD
CTTe3z3Mor5GQ+8eIo0IYtjV8/qS29M6IO3DYiTON8ZA2kYU/wo/eAwYufvIYsAQO0RzZRAzrs3I
ZSdyBf7P9lm0TBlunf7IJcRag77hrbZ0ygseDMyfXBOyp5H9AyE2msLYshxkUZMiTxhnark5Oquv
cTAQsQTKicRtAPbAlVreUSa9Lywej4Au8CxrqJ6lz23gpy9Iav1wlIyIxFIwxa26IX3TlyUoWTx6
tTae2MurjRZYOO0HkyuPAzT6/k2tqUH/zz3d77XP+tTVQ5rom3EMfqWN5VC0UcHfmedq5phRYB+E
Imw9yf23lseZId8siNUan3eTnPy1Z79RjwggOBdd5U35cHAfRzRACVOhvOFIfxedsXU55TMBAdRn
6ktrD+UFye9FyIT5aYBAGJSqu1+fQCZ1dys6Q257nj/C2AUnU+MRKwL47rd+NfUPm38ndMMoAJRu
Iu+uNVwU/zfhfGGkJnOuD30/mFot4GYz8MpbvwBkEH49HzG/MS0ReWsMoqzLRipksekGYhz7K9rM
GDWhks497/XKmrpaJcUwOHZXPlolhBd94sJCd3YFRXSUGDvNdW/ls5FM10W85x8dQFR9I2j2Zr1o
p609l+gAR8L4dZ8oj1rJ1+DgSiSkZuwaQ1xGvtuQ+9zfug+3FCu3lPA2OJiR6DXtCM2lgg9v7B4r
Hvw9uRy22yPPDrCqkvTyRQB7Vwx57ilCmN0MTKtrrlcBsQS0+yml58M5Ke1cNk+0Cv+ma3Cunl/W
1tAYmKyIQDe6m5EIDLMgqQ94WN+Z4u2IfPHQBfeREeJrsVSVV0fpXgdOVMVhoM3p3xCmVhZNqhuJ
QY9FIm/g8hZrol+O95Uk+BY53ZhMV/XYuFRZDwsbvg+gR2lQo3CKbApiKs+t87El3Xom5PeQShlQ
sGMyh3AVE4U3aAUJ+Ryfhts/vBOBQpdh3OU+HAinzPMxZnZ8FZuj3/n3FHYMyshRcbCbOWnc9Epa
I85czrqdgOCKx+K+xEyXNcjRCeGZ3Ubbz79Oc0VE77Aw2R1rOlIuIqh7I492YQVb9xQNnkXINVze
Kb5OezdTun8Y/wRhYzSMkAiluW+wWWkBw6/FNSUtgTi4LKozPk1wJBO/t7TUVCVK0vZzPjyzBLnD
k6MabDWh8yw44BJiBFdQ66HvZetnzFWbSuIbB/p9ZyBlu6ot9+VIhWr0F3RZFtJL5T2bVKhjuGW6
WHXT6QZwSS6k7d3gdmYasoj7EAnFNcIv/6cZc/K/58D681bn3A33XO1izqkSsrO+x8oYnP7EH4A4
xNUjOzlogHB898cgV8tjG332QkhaUdX764wLrxt7gia76n3rUdtShlU1E/9YpqkaTCyt07Mf3Qqp
dJ/UMAuXQd1ziYECiXo2ee/sWBGM5mDQQgG4dSLPzn5M0s41YiusEU316AJ5QQ/Pks66mmYxLRR0
8+iDrqvxYe6AlVYCHM+qqBsGjKKS4aTdY5HoijkwMUysQGeHeLfZIr8aHP7XSyY1mFsoQb5aOqzg
cMshIOkQ/jSKqp8BVWXMkpf7bKv0S1sZaR5paDTT5B1xK2e0xc2cvkMfiVt8AX4bOHTbl3qbLVa2
HK7XhFr1wqvJPRL8OPNYRIrehbXbPcSxllz+9OCUL8Tl43K4bPw395mL0vgVamSkLpPmSXRRgahc
MHj65OjaZsQsSFUefiWnQu3DClB3W8IiPxO4T7TUB5YMbWsbG1YS7bxViFqknYv56jT5DIeQXBsM
1QgsAFgX3EiQuVKaFNVuhoKiV8LEfA/P5EXmUGgyPVVSyzmsIrBPXcPeMjZV5GUgO86xk72s6K8t
wlZVc2RnWgYhSI/w2F82sxS4oP85lAGmx4Wrzvfh+IV18e/moQOU2KXsj97qi9FfIaFa/36L9j/J
pgS8AykeVtoY8bI6HShrBDI15sf820GbOsNxxKxR/E5p32UoQ2ZSdAkhd94mAN85AtM9KH4p+na3
l7CaOZcSctcTFyXI15PP07Bbv6QtXH5FAj7mNdMGoiBi39AOemx1BRXkyOIqPfFHPb/pnLNqUA4F
u15UjGJpkR6GTM9gOLJYubzAjIF0Fd18FlQN4UPrz/6bDnwrljIqVIHBjFO1CyCO8XhAIZaEqn/C
AJ5BnDZajo3puaV9xndKD6PWK4Pj8UP4v+Iqumqzeamemj+EvEXfO3CS1sUeve0xgNnqZZtqL76y
+ibhgvoJBimaNhx/t6TDWugNN3WH5CK8UOHLczyBHJPQNi0bT8l8oXWYxq+YJuDTnFZX/spKFXBa
qaX5Au10aWPiSunjmtOgWrZGazfiXbjUrVYPIQseLk2OI17QkPnjVSwccNmR/mgUFBMwF6b07bCk
SEDPS/L/AlcMwL5pxKKU69IKuBfW6TV+TJ38CZBaPV8bsPamizzmH8DdkcP1IrfvtiO14GC+K6m6
nN/I+36eoFDP/He42NnSMfnqj/SPo+ZgCOtKV7qyoPy9PSesz9+KC7wnkzrosDUF4vDYDYBMpHl1
D4VbX/nTpWyZepwqATEHu2GXRPWvysj0185IIiRW4GTi5tnIt5F2rwgI33EBqwr6uG7ifTFvEYVv
rtZ9Ulw89GUsKAq+8x8SQI2vAm6Ya+Bl/+qK3JXYRkJeOU8jnGoc/IiXSKQliehfjdxgFNj9An+x
F1YoEhJ15gUC8Z5WhRU94rlc8zqWNnwRG0lTIHWvZ2u9LqTekaKEYVK7euQ1OrQJqjC3xAOrWRZk
EoUM9sHQ4WNN9hTZs6kvJV7CG6pB0Oo8KeYjyf62Bd/OWgjTglFw+nH29l0d+fe0mwCrxR5CxuRr
8EfT/McjlI9P4o42t8Rb66StUqEgjePUuZUC5GayaCejeTrfqxqw4IeB/Sky78Gr/12P1W5mYJj6
8nhxhkdOMHZG1tgEZGVI86fia7sVdKC0rWXp1HYzJoDlwoY3/3FC1P+QT/SCOjY6I1JtBlONSanb
yICzmZevWtYHBQExjMA38z8DNEh+WKEijQuOivUxxZ98TgWEAXOERYw7vreoLVzeH/372wjjepOZ
iywTE4QrD/wpU5SATzB4+cx5cyUn9ln6MMUYAeQd8V9rkip5OY5PG75HHbdLxxJEfJKwRY1B4RNC
l+SZ8j3+0hWfg5+MYwEF7i0NUBioqd/vUmhWdi+FjbLVUJtHCXYc1qxHq2itHGHsSEz6lfkb9Daz
uIAy9qh9vbmh8kO4g1VNAwUmXxtiZfSQALK1wjp52o3321L5/NeDr4tU24gCYpi9jmVehYeRW49d
tCP53lxfqVk/pBENk5QuW2MnUz6PYOXy/rFBprduYx3Vf4p7yrHSYbSk+/WoMlUkTjWftNfUwwHW
31PO69C9HT9xnEOVJcOOWoe5t0UXMjmzotqJ7+W32RF/tsqL1sy5aVINpsOKd1Hgkkc5B+FRSgb4
OzKjKALQheBOWjQFkxBHGAVbUeWXki7aoe3n0RBhFIajqC77EB1vJRU4AXvwkHlevgycM4jbiKBW
9v4VT/cVBtqKvfPy9/HyNAfykZSN3FgLmzHgjX9C4gja/PQsVcxbZuVo3X3JkkqnYNa26Lc8Ik9t
e8wEPFZ0wy/rX+VEQiO3n4K5Vd5KCXb/O1cPN4pvsPTDTfXVAgN74fetjpXJO/ClFq1fCCk7b8EY
ck3uvbFEKKevqhc1fQ/WCuZ/JspGBhLzrVVacL+7V3gE7b5D025+J529iNkzu2W1czh+Edr6coqw
us2YOhGnlBceQEQC30lLsc0yWC39srMdtl0MRLiWfC6ZF4KC+tgXh+pK+1y1kuibn45p6XS0ftZ3
UlLmoc7K7kDcZHvyk1aa0VtuUqXqL4QhtT8a/6Zeae1I3G+Jy85rjGaYwEyyXv4fyM6lQyYiOKRC
qULCb68fH8PdYZGKctBO1FnEw/1y2gYe3496eSGnZkRnvyz0szhlbvcVvu0zWl07nhdpQQZEnRiP
Xv2opwktlQ6ybXw4xBfSjCDf72Lmmxw9NiP0mwGYkeeJ+CraIaVJG4M115FB24Ap6bSZeV8g6VPk
alAg3JDxjnAQzs9aCb6aYZIa/wQT2kzItTthtHtMCUKiHWPPpZ71KWEQ4ecu2M4HEiTeQ1rdfmgM
zzXbclvLXe34ode+gFMHFCFa/Rwf4A4R24t//Knn9MxlOMh95LKpCJ9X5H3Yu99C0E0+unLzfxS/
7QmC/hIRAjR1Rs2FIB0dLONfwM3kyaRmq7sfDDKSXabJz9rQFhiphGjrwSfcLw8zYpnmbAAO2Z18
D+5QpJmDd7X1dpcjscseQcLO1ri8OX9Cr2pKBCuddBLRe2x/fLjNApri6lmlMfMFg/1G4muoNHeo
D/RYZ11KMNhk2SzxX7LEtW5CPsG1ffrJX8qu7vrk0ZWIm4T76p7LOHHSEks2hVwn/RqDQT/ffk8v
oLXVHI60lelEgTarmQDxT8xYq/WGzh68hu3fsG8mW4rkZSIRX3SII0o50/FehBi7s4rgDZRs3vgl
+6BUtjvU+KltsuVZwPztG0vDeg+oCuld2Z7hSbnYxxDIRVhIQCbiSsmNLI5Hqtvws8piNX5mTLP9
CEvOxwsxiOrFBMTIPy31e+94QOlHNKMB3lBBvUYQu7p4N58ZnOELnbrijpjkEVmQSHuuB2LraW1o
JSE3OdhlO77HImbgFflR9aDvAILZzih8/z07IKkjIM3XFFxWxb7MhYrFgUobOngUf1aH+t0RW3r8
AVkrqY06c+eHOFYFUsQF3+OsdclRvzZT4wpfcdEceNQoHU7XH1UZM4CaRfpP0PVCpBOobnMcEokD
/4jwD+s3Kg+59t49CW+yS91ms3q+UbJ655Q4aMWCKq1kuhvhjQ9N6jY1yEIkvwekNvast4/64t5i
hdnDbXbagkQAe123W03lqZgnPgH57WmZpT4qqjeCn3N9CIDjgywkNdavBGW5X7ySdQy5gDjgaUnT
eR0k+SB/fO35XxmSPXnpHBInNXlsx1kUUiRNGKB8xFEaXkgKY12lfYu9tJrpt1RSxcoqQ71HYlJJ
gMDbxmixclhOL9KD2t5mzWkQBoS3+s4mnU71FVzL49BgElaZYG90R8T8xfhw6dATkO8g+67bJAwr
bcAEdKqjPuWjMVMcZ7gOJaDTuil1lYO8rfSAMwqDPuyc5Npp1D6dCMcT9zMOZa5Cb+IcLW6OO5lL
CGldk8C+1KJXgrN2xDq4P80wGpXpLlqZ4nGUosfzFogPTswUEwLh9VecVQlmR+6V+LJGmT1HB7GM
63rDTEc/CL3Xsf1eE7bqnw4P38c9RkDEuFSOHFu+94lok5h+WkXAZpFUzNU6uzk1puaDNGkN+ill
ayzFbQKhElR2kdUZtx7lOjMfvq9LRbkRDQNHx8fnz/GOsIn8TIUEM4y1mKOvFbfJ8u+mNbRpthTo
XoXNjwstealG79y7HEQ6ALa08TKg7lY9Cvf68FZSAUFvZO6KYA6KWUaDowhkOLVBBjrd0xVSNJzE
Vv+fG/QDF567gsrwKRxDRj+jdLYkRndP+bzdZXlFD+HA7Vzb60iv7r6P3Jjsb69klr1mfEDF0k+c
GW1S5ei4vr+WmWSGCssGxyV42iuN61PKIddvR4wb+kbEDWHMbMPRe8ZpRNOVfyQOp0CSNhn19Hvv
W369gMVJ+TvKBoKmuzLpXsKL+XFvPGYqoolMfF0J+v2LJtSjkm2TUzNqn/6ttI5vuY7p3hlOL8h3
cTh68jQQMkXO2PnQgJ9NNjhOerovW2J0LZxxfoLV43raqQC2GYvOhW/IhNmgpN6uTAdfZVqhJ6UV
LgnU0KiS5YvsZF5e6TfvuOfp2SPv052Ukiyb2SJhG7Qytycr6qOS63/tnThFiemOP8O8+a5zBrED
Wleq9z1g5ZmRyLH1cUHKCD9GLXG+txta8FfebxmS2vNLwvk2VX2Lhj0WpEFrSh6YnqchBBi7vACl
1DoWJC2R8gmGCL6rsOBHkFzVEzzaFnslyKgj5Y3R7FlSgpMK7Gb2PVr0x9a0QB8nRxsYQgujWT+T
pFI3BR1EeLUZV5ngNZB07dj3RlxGlpALRhLtbDMobSXzRJLFpK0/PrVf3EuRlkR16GBeljTJXGm9
HpIMvfkKpCaH4qfzST2X2xGJSuIPgAPAUUwa/WeC4IJygdygKEaSSuPkeU6Hw3Jn6VnhKQ2nkaFQ
G7BJKgerMcQTNcppb79U2AmS7Jz2JVdVMphnj49/z1i05mbJ0YCyEX/YbmPR2Dp4fY1TJvNCGanN
gFkeiHCwlwe18zxSjr+e0/f6nCd7RMNit0fqbI+ZDe057LeE0RRog29D8u+nubK1KYtb0n6dUxur
vKVnk0cHpYxNmE/cyshHQDASkaKbRvylPJycQZIBjXG9UPKboTVyiP6YUaeg2zWX17kvOZkS1SXX
D08twCFV5is6lDOMFjq6MQY3keGQY33tYYuwKrCJ2Vqe6yO85GOdKdwEXlNtTYrxD33W8sObIHGm
Ml9xSk87xFHjRDdu1zuy+wCRNmUHoz+qwJAMW3cGQ0KZmlT/vTiMZMySwc+XZ8HfLGHjFq0+Y+bY
lP8rczuQRr7froJfZQkkjqu3mxOylUHd4YBTv9s9n87GWHe2eaE5zgKP6dKdS62TNwyMwJgrQt0V
AfDosA7NjtWr4OOeR+dYh5V5cOxdFIQF0rqv9ba65yyWgj0RRREQ4eoU5jgcLbSAxCnEg52JzbHm
aRxBbkCDyuGTLbmG0yZ24OAAVoEALL005epI8B6eAYaGhlcrdCBnWReFtZFXSFwn4mrIwQujsoaO
zJjitiNLIDeaHcGrf7+s8Z7n5dWy+511zEvgsCnuOpIypccIVCmSiy82t2FAqk+DXIhodP060HI5
lqu9gEHB7cutAvAXXjNC5+x7izspPq9X1JgOyxhciIYp7VW/Cibb7TFv1w+/ZrOfwXqK0zibYBuJ
llFKABQUR8bU9j9EeFOhDIsE9fhlVEc3T0cFNhvKVEgFBN1+nBU+FNgAGD1xnfkMuEZ0WWL99K5v
kRdAYksCGS3gras9mWY8YN8R6zWNHus7Ux8X4nJMv1zHp2hw9eD3SZzHzlFynP8xx1DE9GmJzeVR
wuLiI0VFcx4PtBF4O2doM9fIGXEz/EpQDs1P2m/NwbPqRxz5ib2yMjzdPTVR3cMOuMqb7Cjr41lO
UjQNxclXUNa/knuKx+rKq6bkwVCsA3YEPtCYSwuuanGrxfmOBGhtPCcY2EI84qBCTQ//fdt3h9tB
ed8trhrtuinGJXuje0+sw12SkDTVQ4d1uVY7DeuYWi1S+XBMF8VtJ9yeu1GVSyMZ+IG8YSWwjvMH
qN//k+Ld4T2w0rbEKKubdMPtxApT5ffKo05/vaEHUT1kiiChSit2iaOmUXnFYGLYep0rXNbvTTxO
PVzO3KIzJ2WWHv+Jc/v/rkHXKNCDC766rRooE01DcMmuFeGNdOHCp0ZOSg1JqsQ6Kb+XLKmNkupA
KmjOqfxfs7TRsSFrdzfah4k7zXZZLSkycFYRy9sXSIyRf/hmGtfUdVQTQTy+qLmZSX/GBPCu7EIh
yynnXyM8SiyvGlaZE7k5S3lD7J2WidgVLC0TDolSjYDRje7TUMtWYG9VHD8lTR6sUFaiRvvUOHTU
YO+8/wLGI+CAOiYCkqE87tzw2JKLq5EO/CJGxtCaqprkxyePnDd199c+Tl+eWECM1Be4506qtSli
MdHgbSC7mjJ5piXOBy62H8GvOKKYq3afhOE/2Jdvh2O9e8RE8cS7+RF2DjHkdl79eVXXIcQHupR3
Z45DWgENvdhW6GZ5o349WwJ/9oNVnMcNf4piXnSKR2iUPEFXkKkl2sr1Er2bIQvxfemHCJe/gDKS
flODjq2zKfXfox2uu7q49L0ek3/JiNfGtSU0n3WIaHHkhAXThS1Ag8uuN31veQ0bZmMtNgMQ+I9i
WAaxA99SVU7ulht23tRg9CGKHHE/Poi5uUYHJASMwq6/LvzsTcrZqiGV1C3WE1Rn/g2VDnh5lRCl
audBA5zeawRcKigoQE2bYnfIZ2Ns62cByPlNlEHwDHOf/7vKRDCCtsaEV37LkX4DTM/daDjx/7El
k8wKglU/kaya76aqU3PRYeOrp/DYa2PwHQXJmEgIRUy063emcyZJdnJsWn2MqP7D+groouVO+JYq
WUC2GELiT9lKFGKJhgjtKBCyYIr3AaEStWVXC7n0KbAOcA9VQVpVwIb58PH4EzRQaM/jMZEvqZEN
1vBTstS7cDpD6ciKH2xVAq6Wr6fFUpugZEgu4VsNZ0mbKBipHa+7V0/tlSGbnBE/k7kJYBasqpFn
bJZ0KbUL8pkOrorRbAxE/PI9uCiaOwFibwT33AwRdupjdYE0/58TbKbyp9rtj/9qX1klBMqiHGOV
chLcbCFjatiC4ry89UHFSZCCPxcrtSWrncJ5yorkJOMgpOW7r5cka8WHmWJsKD32DVb/ZRCT+790
p4HtZkXFB4d0FSeY4YQ3RUeY4wJ/7qAzikEj/JGUIUGV4u0fWlf6XmNRw6NaeWQyofVJ457ZD2Hb
y5BwTCvAvNssCELlQhD/DnwGrv73F0Odk3k1eeD0DiubDrARxCpTuM2OHeD8LGfMQhd1+VG/C0jg
gzJPITcVTfxwstZ5NFuIfTxQy6uQ6L3KtXtUl/HiZRRkcdK5ESUoWqyNw01o7cL8mn/G5g4VyYzw
o2EzZmeawp4fZIRJqk8KMg/HyWQae6W6DTnM/EK150CnEg8OrHDbil1X01moXbgnk+UbwMnuJ/hS
6ut3uXqMfRfoK5Ln0b2cDPX8tbdqovbaz5p+s7MUaq0cg+Aw9hywFhL7tCPKUn6JkV4ma3Tfig7N
vjf8zuRBhES99dPSePtfUynKm+V5uhXCH9dp7VK4wSkb6wr02iDd8MWn3VU8+Jwz/KZuPPYFeDUd
lmJuAXNI4W2QQgGWU/zjIAqOVcAWk4JjYeBcFQoRBy51jCo47KRXHFgYPwpp+2BJAb0mx7dHcX1F
LOoToHHkWaOvGpqhPsso76pnokRwm72e5DB9RgKn7100e6uPaNfdfWguBN8vK9lK2/pk0QvbSz0A
MIqQHYZojbYQaONkkF3iAlT7+A3oY070SYI/ni578nV+vhUnZp8nsyLmxejG4ZINzeYPi8BXyJl2
2rk/lrfqgmc5/F9TC/SMOs3nj2lH27V+7u/36Kq6zjiqVTayue/Tfs5yNPSnXx/U/bK48P4ZwH6P
iKorgq2T0N2eNe+coylBc3OpzOqmuO8Uh8bA2i8fzHcznSybOcAgxcrHCy9v8eHO07bPzZ98X5Dy
4mNOjltL6kw8DNLxeuUK8m9M/Q7oTt+KdYTwSdZa2XvFcJn9JcVAdRMlbsy1U6Uf3Q30hGhclJJK
VLZdX3lqPKuHuNeW2ggtc5hKjwdFQfGo0ZWyUwj63p5Jw1ieNkbl4SaP4CDUBadHSlxTbApCFh92
EaseogWhRRQkIYAar33FJMRvT9QBOQhVZ2WOkqkTw9YSNIoiXBtNu9nmMD+NB/suDgE0Gm9NnZji
+cQP0isJq6UVUlN504sMUvz2hxm1ZHEKFifzd0tkn1kK0qXzPGanSGUPS0TWPUSIyknFCdeuAQCT
6mkYJ90HX6qPr72yUOuqXOTOF6iKITwQ/zXD7Bc1Es3BMjoSz94lUuS6lxzOP1/czr5IBLdCv0S8
Kj9aID8iJH9+5x+ckHZKIwGDBkKRJqAs0kZZWLLfVaFRt4EMokfS3z/N82kgsY9HCJiXXBlY20AR
tCK+7kWRgb+DmGFGtIgvz6dt97YBlXw3rEKpbnh1DaIlMv1JsmD39U1t+MG3OyLMClQL66KFmIHu
OHJMCYz8AEbRisXahoivMePLSNRBPgSCBVtGYSjKALrENCc7ikKPJ4m2VoxwXPHIgrz2BPXumIUy
74o6PygE/goibLJLvYMIDRz55Lz8SNcdEC/f81pnZ3Wk4znN9n2DGknJrZet24dTIHPX+pTuLbuQ
hnDw2ROpoNTMQ5hA2wLnXEevuvA4Ug6iX1qw+R+1tSlqOmnGSqWZ4NTDewO3D8/BhLg0dp9j1t3F
a5paCXN/CNN5R9pKIrX/aH5Xwi+hmIZEtAvGSy9nCz03V4S+Eabm6z+2vtxeK7wTBDmIy1EmqLeN
JNal4l75XJUYoKNrSB3DZgjAbe6n2q2i86qVPAiuTpAJtO5Vqs1X3lmO0kfQNYJvnxEbNRGtt9oO
WE2RVOxmR/Z4ZbQGyPAGEXvAlQxbl+Zhh0NRy/FWUwWJDaWvTSNWX9PIz2sc2XT7Mw4QeBPAIzIL
XJ4G3kTj4mpsI6JNRduIlLbYj8jMCTmJ2HxeXRuNsshWYf7bL4rW3ySY73oJhm/VJIJ0K8h3qdt2
eYWBzFgIGjRJ2/dOUl7XeuoQR1yveWDo67lweYiPChT86hXFYi4QVkGPs3lbLJ3wqpibtKc+X7lX
nmdtl3tbTGVYd66gfNtZfQgBrkHGGzzmg8cJ2cOjKE3jVKbkGRIpj2riXbmxbjoSHRabnk3x279x
jNaOIBE5XkEVlLFLNKWpWzrA71aZZcXgEpP94bmGT89woUSltczv2aiWDpBPHSN1hUsrRY1iV5+l
rp0tbkkDjYWH8IRxSYPS6qB3T/VmLtMu9zXSPnk+SE+3L94VQczcDSraC16dTHi+wrXmzOwjdazX
r4G10VK26kYBcTY2SY+TdJpOwBze3skq0JATmjS6DJOnXogEX0mwaVFSO7O+eMVqEH+zMPQiAiRd
X1UGB7LO4vIfKmhPih/Wdjdr6squEVP/Xu0i8QkNiR5CwtQ+81Oqj55UjH0mA5AESsgt97ZwZRSM
LwjPA4zpo2RxeQ2Cy3+eX/sSkDCO8Ph1l+10Aoe9qvhNDTJEsh1Ph776OCPPz9r+wVylbgIcaPtm
w33OXFRJqKfLQTZzTA1SRrVDN+IIMdoqv14ZvZsEu4TVyL7YzBXzFvTMASXjuh4FiEXzfVkA9Kv6
u1j4MYpuxXCoHB+C4I/gxqRUWdl8tznwJeFtrxqM+YwpHQUGcD6lzK5q2ZcDvZtKhqDyYTT2+BY0
t/G3qCflWnK/dtXxnJMfa0Ade7T+Crcc4Ovz4AvM2p8/t7JjK5Rrh2RFWaFvJO7sKYHxnKwCiFPm
dJ6iHNWvnr1tcJ3QjWIpTQgwc+Q8brP4/TEwPv9f5ZStjeTgs7Dx/VYNwPrU1dQ3kY4C77Y1QUqi
W2Bxaka0f51IAQgGJmNl6eJFmn9F/fYWiVgEASbQUsZxvuXWGGjE6eugH3r+YJ7LIDjzWWQvtoPA
hMOdkvolsA8hvYiM0BSIZXPkywd+EHFPyNulGQLY1d4ebfn9z3bkBxZwApNsV0RCWs6GiXe09ACo
pDstEUusKahr+SSJgmF3VtVFxt94jxVmwMIqSmBe8jDYMmnc9kHjJjJJ1aMY2P/RFK4h3YJy/XFi
Rx+H5xXjsqpaH2L0Kz5iIuLgudg5A0C2raD+HZWkiUkxr4gzT5kNKX83ygP69RqRO0NaMiVUcXVe
n9a6GqmxI5XBy21BWCP4ggQqWV1Iq+WSICbJdnhQluDzVKyR80SpdiDumsbnODgduzs+O9QRK3iX
VebjSG2OKkZCqGcyXGh/Gm6XhNktDLvpa7WGM/g1D3w7faUW2ER0Cl+F8fXFR7ea8B5KAQXmFgSP
dqsjT+BBdXP/wb8UzNBt3taG/0mfMJaWGfZU9Hn4eT5A7kDYz7mqtL5UUJiceS4qOP1hL1XPykPB
UGdAL6rMSwqjWBtMGUaXgF01QNKSmluyH5dV4DIwqayce6kvsRP1phwBPhTtBxwfImvN4POcYvpT
bHgJaEtncwDyp1YlJsNXfwWbpoPFTjskUHuxQWKwfP6fVJuXjfadqs/8b/ql+m1Z9c9m3rTatV1K
vAJaE1GYwjgGfvnZtoUAdkTfy9PSjLjBdkK1P//ReP6heJ80lrH/xJdrctfk/iFsPUjrtSF+pALq
tkszgXSG7Zzt3zYE/rGsdB86iZb1jMMhTDA9Ua63W/x+2nv38KD3jK1rfNyiNK0Kqy0zfn5Uxo1g
59L854GSTq7ODxpLUweewPLeoiNVADJAq8Sasu2+ffbuPvoWyirAAwM7rD+GeZRSf1lXc23b8CE3
vEXJGqtw+2uC6i0c3/O3ykz3ihst+QmVQdNY5gSYg1BhwtVqnRB05zX19YOzfeYAziAwoVj1Epxn
/YPfkwHOvvVBQMr2tvxtGXiXGk2idpuR/nUw9mRzJxuYO+0fGBuHeALpRPaVVdP7XvdHmF9atIUI
itsvRpqFl+M9XpK2GEiDN+qBD0nGR0F1PYS79bEAXcuGSfYD7Xm/Hu3TFlUWMV6r1pOOVmU8tB7c
Oo9IpgAd0sE88O9aHJLfuYFGCp58dEZTppWgm7Ip7i8T5tIQFU8WukiL6w4XJ/yjncuF6ioAwJaE
9blY+EOebJIoN3VDnsk6TBQZTJ+GpBgsnYGNPzF6hg8tYiXeKJ7gdh6G+K0b0F76hrl1MDgNQZz6
1yuEuJgE3m9evaDdQkgs5ebSfb8Iur0pRuRnpjfNwu3wbxOaBdDOP/Wk2uywrjhwChAZ2ZP7hnDY
N1BBRYwbFemzlAvtH9hEtpWqNjz/tw14nWZ0RYrvpiPfjdG/wEJDNYmEZuWjxd+qbgSxr4Oy5iZH
53zYiW1uCkxAp/GJsM2Hd66QyIRFtSUZIvZ8RnfycvEfAq3oy9BfYFJeS445R9uN6GQo3ja1JKV/
GmiihC7+ysXuOUJNIr90GtZkt1e8Cy8xYWhr55fwV+8MQ2M4hQNfX8QG17fshUMxNP7nnqaBLao6
nAUrs3HHcQPMvozzHq+YngYASqEG7INzXKlNgDfgV8SU2TSXG9rDpPWtCJ4Rog2HFCFhDa4TrHSL
KBJksBUcxhzqp0q266B7BjWbOfF95cTqUMixdeZNvuWSmH/hpwyQVNay8vJVAZg8OywtX/5WV+mO
Xtux6/r2i/WemwJEQl8HNBjpoLioRQcYRaOtQTK5RfH99BrfAYyYUJ+6bA6zaskJKHYwuud5Qbtx
w0caMQD//NXYiqxFEscDG1zCT1vuF6I12flAJjeHaF25E3/HGKrpWL7I9roW+MpiFBvxAHN8X/2/
kZSlIQx3qYwpt6drrsjjlN5KEDD3LD+7R7VKMcBq2DC8/4+aIiROlM9PRa832oooy2fCkeFaQ0uE
lfB3fmAtSD0vKGGlm2gKAEfoyFKik4hXD03Q9ZLWvqQrUmHBMt/y68bnBJpHs8ws3h7RVdyM98JY
0Trm6pePJK06jivRLyoad2iy/PMlwyYvorMFFNDlDzhEzb4UIzDQyNvdXFqgUk9ufIiPvA/wb+0V
XRMNgXPTvuM5yQYGFwx7VIedhuXrNvGoSAomc3wt4XEhB/F6kteiw/I+zg8QiV5YNyC3o2KmSIfF
rIIBUeowKOCmKi0Cq4IpBpehDFVpnU/1+svhx6nKa8L46Qn/lrTPgo2D0M5WhqB7zg08B3Bl+BBA
H03WrG6axorAQwvK3SM1ATpRfUncceXckXFNUA66SOalz+Tc6SPaKfOhc61pjyjDnjCUja+m4P0O
b62sTkZ9QKrsQVTUPYYRVikPTtbc7ovu/J4fCGLjcExlG/0n+zgQ3cJTYxFc+1c+4d8EqroXFKsJ
/6qXSu6/fMk4GZjCUAGK4FIs9CFvlYlzttNnUAUymAUy77G8YuRLN8xnskwayoWgjNibwyZaNVEd
AlGXsxReTPUwbhUgVKB5fUSWR5Gc0u1kwtDMmdQmZmnVkQAx7D4euvEIm7oUwqGTPeH2HMQ1rQUk
xYeru3T1/Ajmm4MAu1CYRlXmgLnrRgKfDOUHemiIGJ+/iUn1vSEcUPetNx68E3bqwzhLXBgKyxsl
yQxYCvJCRuHeEpCo8Sv4y4oAApLfPcKoSyem3okkaZEuvmz4GG2V+iSmNOr/ADWNBnKDiFlt9hB0
BUweVvWVIYt/CRHSNyj5ro7otOltliVHS6BtAJ3ghwnIM63VrTWwEXDPAf9DWlsOiHcQxr7k7csO
y//UokhLKO00Au24R3PWt6AG7/8DWCR1fAdVtPt/l0JEitzvwOPUAtbbjT/rk8B3GphGF3Ibyduo
3WKIJkJjXkpWU2OH7gndU/uaiucz3Sr6RFZ0kIcdhlKEK/xiI9MT3icY4iI8XWWnesJd05a2bNXy
RN3ydcGgDUm4i7/GRhqSVxFIAPV26kipju3MiYhhbayDEX7Wc0q2dramFZ8mgl/eR7LKGQGnA82a
1BczMtktAtBmoNwHj9LCz8fzbsZ7rlAkRRGbHCbZPJUfU7hjtkojnjR6Zkde03/Vkaecr+DKPQzO
KjCK7A4eGh18UxhR7qMBGrljE8XISQ8mejZOV4dj8bUVNoCingJkc8qpN175QOVgY5eRwAX/X+zl
CL/1qVJ+TJ4vpzQaHf/bTFvQFmJ4161uL9fDwNYnqm/bhKtpvN1ccngJB5HYXcrAHYPzxhQNFH4K
aYOQ9TNfhKFd+rXOb+JvBa5fb4bAMlrEJy0sGwX+Crerh38zN4pFITuk7hzsS8Wtav4CjjehA37w
alNAXxH5uQ0fGli7c9lu+mW90c7Onh6i5XMK5exs+ymkYAaL6Mu0SM4kLY+msT8tHazYK7YC3JaX
da81vOk6IL8/cRPX0kw7z9uKl3T557kopdnYtdbDUtvDRjerxB1rMFzEVW6zP5KwsBR330X6QJ71
h9huDSO/SrxwNYEZiYjXxn8aV/CLjKBx4KJz7PMLlTfGFENBmr0+bqwjE6fEThIw7CelY8uNvRPD
Lhfl+2dh/Bsv0tlb7ealY2FgyXJZwOaIltkNR/4wImmqZmKHorRyv7hp8uAdjbbcPSu7ScdRXDcv
gznpsUREBKxtwSmAy6pgzJNeZZlKkVVrPRgi5ZVPpVLA7Nz7rtWhtVkSFyeYG/c9594AHAJydHpH
r05w8jEdc+lFEfQB8NoIoOc3BsEYMCLt2aGav+17mwYclT8Ist8RReZuLgMMjj48Ww0/k6ZD9Tz6
aP1xinYetQhjrjPuI6IlQWf1zSalf0KVwq8N8XS2/DnG8Np5vCHUgVkTMUIUC1buWqFmWe6eSK4h
+MhILHCGG9q/DPn+/eBRyug4mqM/sktGdVa5RlU0CFJsqwnhe+ZOlLNX/xwOS538ahzHGD3iFuuT
QO64tdeZGNN/LddCmS4oY5YejtsH2vamx2kW3KUhqsLjluBc+nTvcVCRFJ7nlKGQDgNpwDsZBChr
Skke5B5AMEimFx3A84Xt+Q+yTpoh4dvXCkh2q09FPvjRgSElsBVgV1vWyrjTVTvwHZO47hGIz901
TuY4QqZDHgWvcTFG9Z7V4DtB7vPd5hSagpesQfQ9dPUsyOdbRsp6imxskokwg+iwAb9nqXmPBCQe
zNZcIk42rlzAtqdCoUqBfi6e8fjk5TFBlsRhqA7C1mbg4mPTyjP2ww/6Gaj2uv0U5N+j4+mb94OP
UxPs1uraUYYARANIPjKnptdoASqlgPipBK/MYa2J6MpFw40m71pxS1e8kH87hRRJnIq0XKp2EBlz
BHltImH6j6a2uoF2fpHPXJw6ad/alK2CsvnfK85ok8oQP9fkJMVHq62o+oXpouakbonqo+IAsRFr
4tDaBp6WV8+o1qXZdcFOzvuM4XGpiJBBjh5CO6TuPO/QhlBxBtGEUKfyTo+B9AQxWNdR+Ha4+rqA
G0cE6JxH7sy1DVVqZjsLxg0LumZKPsdsK54+eq5qaV45DbLreTp0Zab8xAFfY1uBQlS4H8nZsNZQ
RoU3EM5Y9sEtz0cfQDQty2wbQRetdnBRcCzsvLeMmi/cxGM+DQHps5wt0VWgoldw+B5Yk2qy1cLw
ESrQfViliIbJNRX47ggwJldHNA1Oz8KHxYQ5h7M2UX3OA2kAgty4Nwd3yXEgD/77yUDK0m+FEI/q
SHDNDrSmf6NVJN6zNcjeApKrMgM6vDnEprYVRHcYadnX/10EgTBR4g/iBFv64XjWbmsiAohKrJbJ
n7FAKZbTYsajshVzBxg6RNHUhHOijVWD3mlorwK52EzHkHnqxGaHQ+NgiuI7093zD+QoT3+5zWse
gwwKwnFCoS+ymo0wpQoGsozQnM9e//bl2jWXX1hDjXH5wwoL+gWtKt6GAMQjWNFEMTj0sn17jrzI
9CBGqD10LbjLMHrdIBYA7lTeihWe2THUkvbnxG+5HLXytq6fcrpNif0X7sndGwwwo19hECZFgO6N
tENYGvSrC0FwIKgDQaw9x7ZbO52bNZSqdIDERvY1FgrgEirenh1GnY3ZAL37NhXkaP3hmhWUJ1i2
n3SEeLK2HjWkUKONcCZOrN+DGpSfj+0rfs6j/PAfo6LMtqL6GbX3fqhHhPs0p14LhGGtGiFcXeRB
eqDAkHqXPaD8dnOc02GNy7BCBjZTvlC7X8wR8xYCIeVHQ4G6XqGFg4GDLxwGtQpn1D2Bw/HoS9Lj
NsQxq8HT9Tqr8wD4z7IwB1Y2JrJ5RUWb74qGv7FFj7PwPV3rPxHMZRuMRkVNdIXnuln+woqeczeb
ynp5HEBpH5gTpcK0Mb38WW6xcckS9WiOQIU1kCJOfc/cui7VJS5TbPwTfMHCQR6LI/XCV74S9QFz
DANW95nVNrbUMDTYZaUZ+6m/KGfEKXomvJEYFgRU1p2dR5oEfcJkit7DuchWIoEIQ718KFUOjyZZ
Aqk65DrTvQ6w84Kxss5+ro8Ac09ooHbTSIai96B8wNWssrhRq7cOFMV0Gy/f6DAUgiqTsLFAu+bZ
IOHN27sB+SD4+ToEDa7uGjM6EwAR1mcp6jgNasastm4wXL5fWdZOzaNSzaqkAevP02XleOIT1vse
eN3ZDu0WpyHUxkV6NtlMYxNPFm9xQ7FacGPyKOL2j3Eb3HpX9yp4ikSYDjT91tMB1IVXKM+ABpSQ
jmy9QmLlX3XEATFC9dv4loEp/B+iyo/C9xPLbCpVINcxSP3IckhMXUEVjm/IK+f9HCyDJCXjFmDS
UNyhowJW4Rg9HcpCxZg6lvyR9VxWDr7qX8G9Vl7HNv0US/qGEIN7tpwkk7jL59jSou471ucqCgPt
bo5m1PA8YvGw5rIVTBkKLeQJQatOhV5X0jZv9/x4BhxHollBpKA0cT1y6aCHBZ4i0s7xQO9upHdZ
fKDnNM/QOx2FpnDfOtPakcle/QwpxUsmgNZAkBMFkokVKOuypxeFyYFBr2G2qdJRrJGh+mg+hW7a
lB07OalgnjHHZR8jNZJSA7pwO6l7FQQ/915seII93tiWi6jbWhoyu0QWlvNLVCdQAkRrzOLqrTtg
KD3RgmWNyTdsk/Fa7EL+P9mBfByqpEIVeEXj1InGBUUynZAb9Orwm0od5lYPT1WpC0wkk8XEhM/Q
azLRhDxoHoVQ+KOCPYqmkAB5nMGq4miiMd4MNiD14ROySCmXi4VydNED+Uh0MY+p+7mcLp0TeRkS
XQJDgoUBo37INA32/vqebrg0q8hKqCAok1zgcBS/yf3eSKD4GIRf/rHxWqlPwil2e8lBUnXZ6e9m
f2K9MclU6GQ9mRwlI553KhCCHLrCVdHLUC0Mc10zP2LcGR4Kmip5ugJEXyNy/wwlY3YgYtVUbQKp
M3pkkBOYP5frFERedbcZ/K3YJkk8eu/4fJQyAdfr9P83tvllJSI/hVsvuSnmCS3f5Iy9esqMaHEb
fJzXtbShW2ruSORquGFcmQFGapQN1gn6D4HV5+DESgWAPqus2Nf1gNB19DgQmSenh8ZlQrOzeI2w
+ke/a2yYuOUSmbdc1Qsurbkvlt4DvDU1HsKafDcx5abY6qKffQjFD6ebbaJtSJRarqioM8YuU2lI
7ED4b4ezRzLc2b5btgJH/FldULiMVGycwycQ7+CFC4e5DkRH+k658lZ2gnciHVeIdxqoJkhGBokf
kg0fttc7KVqw2FIAONOBIcLPPklppy3/TVyZWTIa7eWiH5vmyT9h7VV08bgWcWf0+tdY6YRGtCbd
Zt8PbNupPAyxd4S0TxfvahrjQj0+6oevAF3yQhpee7GYf53gTBzrBQpt1DIuhlnECqoT+EQJm1py
1hKOnesZ/519x2SfoFEW/u5e+1ixJOHDbCOf2HWYiyR715AKUkg2tEnJ/Jf5ICKItPcvpnhk6Pbv
7XiJWCe/9/CEQSAK+1rOflb2KEgbXqnE4xAB0F2i6RKRbniaWpa4hEtD2Pa4uB9SiIlS4YpX0dBY
VqkZ+nRjGBGDNYA6AkNeXwkJ5MQM3uTUvi/+S41dlywpKVPJJ+9KBKKesjw3WG3z+ogpWrGSh0io
6QwhtxGKosmLbp/TaOCPN9098ABoXcUaRhMZBEB2s88+t5qpXIqP7athaCZ7eRHBWmdDjtOz9poN
t1QCzX/NKMXuboNrkeAAj1H5X8ck7SIZwyBdHlM+kXpZ+5wY40x+xM8INclpZ441sASKhdmqPKgt
ROLBNZ87OrnYYr9k0Yq9OHwdXWU2R8r5hBrwLwq2IOjSP0VsnyeBh7a1kojl4ahmTmFC0A0jGfHd
sPxLAWuyss3DZ1+UVMrWiItvACtTJdt9wOno161CJfu/1gl7t9j8PCJY4moUPCsogyteuNsUBGzu
MuBqc6bbMkplUoEd2Jg2bf6HPhp5vPzSxWSYbEtYJ916jBM7KFZAy3Pax8C7PHn1/wHTpP7UtmfT
HFegfrCsrf2nrkFqcJLrjmj4jaLgbC81v7k2u4bb/sp2Uo7MlRLIu8+lxoEZeIzXVZPyLmWzNHif
B3XkqUGwSexdcVCICnE93nhg8D3YlrnBR98lBf3FKz+oHv/DxqHL1Cs4Dhn/0TV+sqfzsBIJHIO8
O6scqOAl/t24EQM4QoqntrYbaaHGJIIrIAZURjNp2oHUpCKrnmYVrmS39t9Fd1oCRyji1IQtMGGC
4HmTl7IdnQGlIDJYAa+68HftApxlZ+o3bVrvWwtIOzsFHcaSx0kY+hymy2Xz11TnDFWw/BasumjP
tyc19O4pOc3oC2VomerS1mqzXQOMub1b+5Dd9RqKedNlCgbnlfk+2fdjWG9/6FGgWkMtirLScokN
FaZ4Gz6IqmSnAEJCB3e+A7LK8NOSg/WDLKW3SDLRPVURsmbWgzDitUjQBTJKIr+skG3hg206CPNe
CEcH5zYPYQqjSuwFuKYtyqPVBTR5ZWglOZb9JTACSzmD6rRTGdmRx8f/ODFwqujTMo/0H9oWneBo
RBvMggIWMM9ndbhHGu8pvHfgk+omRZD9JT/UQunM9g+xKuKWUzweXR2nA91MRPQePUv75k1HrtpH
PxwsQCYtjC1n16mptxmE18GGGVvTdjDCK4b153GraHPfQDFna7QFiDm1Wj8YakPOxFxgYdfyj7tU
6S5NSi9OJMpaU5xdfidf5EuW5gfneUvTNtYLf4fLYoKfB7HH7YRVnmiU3bM+yAEaQQj0gXOpTyBQ
qjtPu39Y2Nsipmc28ymS8XBxndQIlXI7CnyZY6H/NHNvUyPT36s/rr3XiXLXM05qN9bkIFl/co9A
KIpPA2redt+pshA9oRux5nhoG6NScrAutsu8Rb4Sg4fAx2QjoMOG8VPChGdth0U0FCMEie1m9r0w
yLHj4buq2dYfGyMEqnwr7RdDyFVndHZGB5fOnmLZBBr7tN/dN7bOF8qtfRiZbBnsB9Qu8GubMxMe
YPgZqe8kDaC9Zs4WGQRTx6QbvsG6oE5cq9qx1E3M/aVIXqTreyNOwQCtW0tVddNzuHds/gX8cr7J
QEpO8asoLnQVPmDn+IXf1PNaWjUAb6IyVvukDmgBxkrJJcCqgycfCJLJHgV2DumGeoTjij72kHCS
rwgRJRs0OgH6+oPzOiX9xr35kKgac6dFl0qDswbS1YIF8gJrFKmyApV/przVgmGM7DJXmX1VsbuO
QAADbGLpgCjOvFXiDL8p6Yof9LEGu3W/VzjIcd5uzzF0eOU5LZVUBVTdIaOHJ3JprbIcwxasicbX
4aAbW8nL/mj/K/jAgtIwFtUx6z4b2YYjPd0fCwE8XG8jEyptTaH8UWfHfqUCQtgXdcgmj+EDpVRF
mi18nV9GQ5XnaTMTtPP1ggBvdXknuq4TZawp3x7jTXgQdWB91D2ahiRI2h7P46MtNdeRuiPmMa/Z
MFvOrDR/rsFwgNL9cav2koQThuIr2uo70/C/Zhl54B44qJ7ewGKIclf1T8+4aU5oxYOWFgSOU6lX
w+tid9NkNR8XMhYz8EKZrGZocZP3qlb4aowxHqd76Qa48k0z9HYsAMqetDCQ22TAjR9pDKcFOAZO
+n1xDDNlXvZ1wBBFGA3gCIsihh7t9QvItIxHYgZun0Uc2otWnzjuCFmOdxBua5Gew4Tv/YAOcO7A
3utAme6wCeoIfT/OYIf+Ncho7g2K8mQaeLWUNpv4Ld/9MiXBJx9EtzduhGr6xWtqRaA+dCW6xBFi
SYqCirrlBy53LbrprM3RUrGWumU1i7tU+rDDyeeAGaRmMQfolaf5WA8IK2xqreD9y+m2xQQxdKpx
+CiAJrwHGbNIauVJOKOK8zUImyuT18xH+ydI7U8zcqmfTxAZjKedENDCrbHBoTUgrfu+evwLlby4
XANuNRlbaJKHPkCwIgxofm0FhAfii0kZ8FusuDJ8x7i+gHKsJZsJlxNdBrxUZ1EbMK4jCFAQBFP8
3qCa/FVHTcew8D/qvmiOFtiuMHctXpVypZ/qZZ6k+lTnf2bqpE+TLOlA50ZsecMsfaBBCFX8l5Yz
K2ZnkJ1IRDiFEiXAYTGooT4Xhh82p4fsas4tC7xOZdj/ZRLofqKWcQuIm+kSMciULSjyVf+ibf4l
gjgpxMI6cg8dKBkzJMxflgL8dHuQn9T3TbqDlxW0KGxJjqhtmZ2rGKkRGALCXIALSQcbfXqoRcwe
y/nMA0kWMwUMkO5GhJczpvXpyojrQQlkz8UQgk2UALVPMS1RixIHWaQXIJeGa10aK517Ep4cO0iF
3VhfRhQ/EUgpa512zH4/YtwTFs6CpI4VBnbG8i6cioKqKNmd35V4T/ZeBB1Hpy7iX1bRBeE0s0iQ
YQ0NLikMfe/LT7isQwxFy2JdJXQTps4b5qfTx2hHehlq0wfQUoonY0qydbDMHeC+FDQWKapXcihW
XrDzeFSG0Skv9AXR7EPcYaFMPnbB53VxceQ+bUeJ8Sj9lxXrQRL4/i81SuGBgneQ1KwJnu9VAMq8
qv8/x/ujrwlLVnU+DFy0Cttw99f/N95jrc2YWvvsumooA8yvpfFiTwnJ3+lMD0x9yxaCcAixzQYt
N8r93RAzUCgsNFJWBZG+AuZBDDp32k62dRCs795ed+ttYm3gq0pR22NFyuNxJ0R+DW/5hoKBZtIv
UCyUryr/jcqbhLoTHQoDJLaY/uFVyNxh9cCeddEERllRK4t9BTL8O90tkSe9s7uIfb3I/y84m2wX
ilP3oP8+B3ZOOQW7VmjAhfgyVlqXUUouEjeihZVUqqn4FQYhLz3JPp5oSLEU5ybeOc8Y3ttNuUmE
jBGXvMXQNYeug5zdXznPI5YsuzqXkJ6OdBexyfdmFGgN75Sjem+qpjwRcZzH+mkxZpPGiB1KHZrU
BCPipQmLtBLe3nhgy3LF8yQCCyP7igHGL4m7YJBZeyP75V4b592aWo9ulrkA6f1ewVYRFYF8b/47
KA7c4nG3NEWD1fACYmc0EMmsB+r5tW7Cvd+MAWDqYvfCaGRumVgPBT4B0WUzTD50olq7oEHUmN7s
A56ot+PIlMWn9TBOqqldxo43EPD5AQgzR+vJVV9qn6TXdw0myq82XmpBYb9NWtl0sIUulNkkd5TF
HVD+4+KTneQdjc6hwgqDSp02YXpbPfiPjHpOg8XL7G2YYfMexX/TMfDxqtDGpIbP8G0Mfujf3YEy
x2nZD7kuOZ2Rxd0ZBF/heZvdxTmOYkZPWfmXwpE47nnZ/yHK5rM7r7YgOq/nFrEHt58JO3lCllnD
xxwjCdyM+BBJRp1qmb19t10bEXMQ3LvB0ir91FMOa0ToSh4+WtfpPVzikVbV/V6mCsH0ejS+blgY
sbxMFCiGO28oKdvlHuUPqmIeh4/krwLYZK4VyJsG2zuWXrpeFNtzqMcm55olT/NUcaryKyXOiI5O
uPICoOd6Wzb3QhZNbXpz+8mn3fwzSX3s3X88FlLOKJZy9C+zYfWoDIh2VbsdJ21bwHQW5D2Lalpx
UAHb6xYAUrZHggfrbDLrf6AQDguk0sqM1GYognNJXi1nfCdyL866vhpPVJ/Nt1+VdK1OfqkOVuq+
NK5iWnhFw2KITJCXWqEhPJQeLjCKb3U9/cmpnLPCFdJ3la/FYI5yN6W6gmNhZC7Oh0vsgPz59bPJ
skl1vGmXjd6MGerl0h/GRjwgRyhxMU+4KZthHP0661+kdoxENVsuISef05ax0/A2w4E9NDkW7c5B
E++0ShqI6pgrFGuZHAUPB25f9Um9eCRGXqMeVrYBOlibyXrClOCouWosuXUbkLV+sF1+QV17canU
ZHyz0SL5r3CPykiIOiP216+hXH2TMayle6ibeG0HKJRHwPp/2Ztdp50kh1SJgs1+vfYMR9ABUeAu
wh+Kwra9jy3AURLlrZ9oSTjTkQYRSqp96hgErTkVUIDFy/As/GSfUtDzUq50DOf69jcRBVYZ32Zh
B+MvA3aSyKAw6av6gYc/Q5uTXkudnOau7g4q8rOrwKRMUyqLkbuADLNEbLdaDbC4/1Eahpo2Ld1w
tmJmuS1qMjVQmTYWOk7RW5oPT+wlULCZMLPO9Ny63kd8g+uviDfxBWgi7KDgiS5dAMXY3+L1Kl6A
PvjXn14T8/oEwOfabrEzWNmdqvt9Zvc8x0afru7RnfGHJ0X60v91DDvCJm/cYt2aa3XTYcpRS0Xu
X1nux6sRRJkcdcLeJ7w5rugj+pldEpT7FFElEbhXqgri3MCRaLCcHVwNInWAUiMkrhL1z0PMCQpk
pDVJuj7CH7yGR3bG5MbUOdpkEi/DNatlWuqD+CIJ6V8yDerEo5G+I5KOIyHfp6PReGPQaOAc8Bj9
+s+IQ2LwL/wgem7MQr9yGB8vcgxlR0c5v3KJ00lIw7MT+VhdLtIe0R4pXPxGVWjoE3VbAt4hnf5e
lApWay2+sQDQ6sC4OzEBNDb2gV3muCNRwQ2lemAr45xS++ullcZxK7Q/dGBUwxzGk4IJW4QkZsqR
JuCh+RKMcgDI8XNZtvKSsUBIcoRH5g5JSfHwRHeRTxLPWrFtHgYLwkZOhOnO5Z6zvD22jvNMZsmq
U8l3lYwBhcX3RhefUQpXl0ebKgUZSfB6PkbhkPEEik+Xh8zKmLHbn++edcmn5ZVHPatPsatumBf5
/bqWlWubQKEKfJ6hcA7VnXyz/HeTONXsbw333x+5pUEzeIoAD/L1CiXRZ2T2IfWtzmnsJ2sGAzuf
92shbmklP9ZRlanX6iswdwGUfBLMiGWCV58ou2lJt9ixfOuuRkbfsGcyNI133YQmCIbwZpzw/XTm
gDcXSz4zP1GvzcaYbfBEk7PjcfYjb+CH5d46n9YIv1smG+RmZtpzImAEWSVsQEKQQCNwDVDBXU1V
opFdCPdw3pF5/2e+Xb9kThF85B9DNugtIbJL24pHRIRz7onMKwulfZmT32/w9P4SEw8EzZxeBZwW
Rfyguk08SjDzls5fYYR3U3dwNVeaY2OP0Tr6giWXkys+K+MIh1ckda3VYp84HZ4p34ZX+SkKc0n8
qcCrk910Yuo2lmxaKcmn72OnYgcdIll4enTtLZ56YVp9uUqQ2jhNYghjZj+cfLjQA3/uhRKo0T9D
uiKN/oIDmjLZmEBDqGCBjOCJRbhEPdfgRI6/GzXhUrba9SNrcqVf41Ia2Sq35ROxbjXnFa4Fa58a
iqt9vDLDfboPqWwPDqGQm5/mz9/BgBwmoQs5uOc/9tmaLyMi41SPBbT3tSxigONeVONaCth1g6JM
Zys4+BLiWgxFpZnRzQ20g5Gnyp4qiBpc5AADTuBrOz+nwox49FJKp9PVTIsfmapUyga3rgWVmCqG
1XbQHyppJi6xHlaCdHfXTrTu7K0+tCnMc0umCH5q6IR4OPsTfTRIIb+7p5zUfyUaJXxzRE77dXCB
Rw2TADYXLnrNapVdpPGVLrDKlPQDw+aMixxU5kYqqO2V26vFfleBRTTHd6NMKvjRz0lXy5kT5aCK
Xd3Nvzci5N9S/8Lt2MpBAH08Kqx3K+br7qP64Q0yckylc76DLvguGn8KbluS5x1Muvo4uYBkvGa+
AO5qtCFkKkKUpOGMJJGAOZgTmEAcRGINB86vIBiR7b+nlrvBHNxkg6kZOzz3NP1PmnCv84ebOfAC
uGD9WAqxqG4rSVxmsUyB7NF5GajWGHlFE5O7Qz7pv4/RG3iQPRCBd1d2yPrhLqWZuCJbaP92YeoC
3OBc6hPuyOelm2p3isu6as2sGNNvKIvpMxuQRFEBNtET2IlNxsyFUiZ3jEPAyUet7Ezq6pxmHuW9
bgvdPNwTdDwduzGLb4Xw2/TUFDPBpEAg6mq4+x2vUeZ+PG6LtDvWgXHEoptu+9R2mbsqVeI6G83S
uJyH/iZVfFhW1KoKbo3b39dJKEyPd2fgE0EeM8uCLUwDLYceLU4EZOC9/HEQUE/h6NG2lQcCns4T
abBK6Pgj92fTuCa9QUVkKU3iiwMPb81a/Y02klH2c4uTduYMca8KuTkCSSh1SMWNXVSVefWSktmu
U9V2XpQaRBFaayUJfzdBgIK5vymSIcmHpj6iupjvuXPRjLpIJhPmvtSIAISJTSvPeTMwnO1mrn0/
07trsDeheNkURGRrc+kTgIcgOqFZc3uXa1MIUPxcpsNRqNGDAisv2toIz6+r4N1+QzHVVz3doBXc
UlqSRiGA8hfX9jpfNIQcfsPGQBVZBHg7rus3Ze+qdX9+NpVCXvtKEJgQFmhjh5QztNNrT60JpF9f
YB0Hw5TtIcReuGjj6W8E8sRn4qpdIn0vI5ar7HlSWlUwq6N9oPeGlL+c84YsyECuU5KSj+Eu3F4N
pPzERkfo+xYGja+eXh0Hn+1qIJVqzTHCW94E0wdcmqjvxYvCTDyo4XjMQMO1dMlsoY7pdutrRfax
NAaJc/2BlUS/GM8HfYhrucBmajTjOVd59dasETspZ+mU3IZcqi4gZUIWN3t1tr3dIYORAkTjO5im
SipWpsH3Q+pdtLQhL3tL8/5c9RXiju9jgUzdrkiEyjbJFW+Ud3BuE5tX0zLVrhKb6FaZ6AK7GQHU
x1YOxI33C3JrfxDTpAgUI3h/+2CkvhuDXy/gWgSKIw3IajUG2nZF8g/7QoA5/aoZ+39BCX1nDLrN
sb61eKmkTGtvOThblbjgfMI7iAh48YldtXX6FND02L+b2vgVfg9O+AktOzFqwu0afjxvDbHukfBj
7M0AWbTD7eF30c1K0TssENDt4TixdQ2fBcluCr/VW/h3UlPuLTCVymWH6dNKRcpc8rM9sVjdUjtZ
AeQVh0GEs0urIUNQmMZPljmM3niCLaG4yiuN3QTadiYsYiY+vHO594e7xIaDVCK6KhZkMfI7H/hX
62MvvAJta+regIuHAv4R7QdvM1C8NSQEZLwixWp1+ESNGf7IihLQhjfP6/mwIdpTIWwjpcE7bbFw
Cu4Q7zoafkz0ykAAdJ7jE+5GIy+8fGEfyfG+pRsfpfOdFj5FAuXUPcOYs8v69wN6J8qZUXzOCTR7
Y5gdeFWhKmm+opQn5XhiIGmlmGVK366xHt76LfIkd0SDW6//vKOf9XMA3Yrjif4c5TP9Nv74+66H
h/tSiY30J1GXaPakYnNTQjapaAPln9ZDsqaUsJ1XKGOVjD6lsXSIrKTQdMb9FnqgEIus0fSoGkgE
+RDDX3xBIgQ7i1gl5qX4siSMlwrowwGMaKo94XFIpBxZNrwWwRaYgS/MFvajXN7TSY0xIWbDfR17
iEAhEUf+YYYLD/xU4mxTFYhJuVafCn8fwJmYzJoI7J1tl5P+Ir+tw+EvaFS/2JVe/yNBlWI7apF+
5c4g/D0pJBM2GO0oZyhAYCUpY1lfe/ShsQV9EWTPC9xuMHZL++nacgvUqCKDs5zUftMOxV7xgmyy
onCkXiND1d584F2kEMSMN+w/FDEZjkHyNpD2+FRRzJgnxUUyJ5u1q/JOjRXUonB9MI84lkhL/j1E
y9XD81Np+HEDtkJDjNyg+DIOQF32uKAJ2/AT0mAJrbzFPuxUeMwshQySF2JYwOO5mHEuaXs7hyi9
abbmiRFaP6/qspgh1+9ddJGx+Qce5/V1HiL2obxAxON6pL5lxCLB54KSje8tUSD2X/yd6Gd/z8Dp
nhfQVBZu35xaJOL+YpePPhevJRXwF7P68ia8tpMCSxWtJiEg5TR2NW4j9v9IgPOoELLSdiGs8Awl
DwonD/raJYtHY8J6+fU8KvPXSZMwuFNS3RpKBjgx4xQn5oxXqzVHCR13Bs4Qr4S0X9q/tFl9xXJp
OdM4ev9gnfO2kGzA8NnUymdX5BCcI4E1f76QAdtWQD+Hw27atryfs9oI05GOuMTT+npZ1MDPR+8i
rW2htvcu6oQvUR4YbQ4fRKu7a5i4m+LoD7WXHh5KUXFkhKsfPixwgh69nQrFNsB7CW9pxnqgRPUe
+R8ASl048ns7b22S4OI/NZcmDlyeGh+htdWVlHpRr1m8G1eYQtTFX8W+QomLeU108H9sQneiFliu
KCgWegRMPGgpR4kf5128d4EUAAus6TZHClNmRh5sNTzja+9T5phpDraI4ysHXC+AlNHuLrdZkXiQ
5kxoe1RDla9ZX9TyyCZTCbwWmqlZ8fs0UMrf4R6PE/OiHYun+Cf3oAooU5LLdG2LXeLukf09uAwu
jbsVlHZ2LVItk+ZxPFg48DYLVhVXi6lvHZn03P2/oMIG3P1+6iPvLFwnMaRPR9Ar+H3pwM+3Q7zB
bufzw8Or1fftVLXvrA3UGMpOfM/i4vcSYf7ImhdXKGmmQb+jCEMUL3LH5lJ+swmtinm0/kDeGscs
/p57H6d2ln5tPEixZairtwJLb3BaB5KxqbcrXJbPydIHtseiMXM0gE5BHw/Bmkv9YNqiJvzLj/zm
HUv0kjtjiSRqkUyauN6FYv/eTuQOmhDjW2RFf7byTkQh6N3JtrPqGwFSZwbOtQ2dx+pCqYYApHRp
cAXC3AyVYos3eXBprZ+W+aEbHLeDSinRQF/NZf41bcdPJxK77M7wNYA1wmc8f6WA/yhzA+1nSiNP
77ezATBiwV6L3bfDH+RCuaynvOtTIr/3lZgMUDj4XDh7i86v7YavKF0S3JX5YyExwRMh3yg7nsSv
eJa0nGpgmNsyiFR0dOglcQUI7jDTaoczODx0X8dnmr1mTu91e5mMOa1AAFyyMWur9wW3QGLPLtZW
Upwg0RQssZftMVVeqXHneisOqVI9sSyJRjbr0D07iyKIoJIhWYuwyNyGZmUMYqg84gDs1WKoqbGp
9IE+z9BT34CrrfncRPm5OXVD11YKn+Lh30ULVs3Bs7hfCSTV7vx6ur9o39dbDq0gDDKgwlZfwvVT
xsND6Nnz3c45NgphzfT1P/bF54AXVrwGgpAKxfaKCLdrzxO7iqN81nquleAd64FhgxqoE/OM86qj
z2wR16erz5EdtUj74UfyCMHthY82xDZI8tB20TTTxTyQXvagnYqHqokuyRB8vvz6A42/LEjTguei
oURM9MdqyA7iU3Cloyl7LqD8Mwyy2woak/Ahhki0rMiNNU7PwOjndatiDTa90CuamGyAR7qIlGJE
gaCOhIx7h5ANZDV6d8GD0E7eeESMH8nxzXNhADfHtLd0SmAvREOqhhReIonVSAW1WG5gLtzvnHfB
DREHAoNffnU5NFxWxQsKHDjDIKinOrnDomzFrErMfHuC4vG/wJ9Ihvm5abi73JnrL6kM4uvCsDYI
xjuADZ4F94w9cU+3372UymYKyaQcNSAoiW8JLj28Y38pgPsKBJP+fWZOhi0+6eN0FmHX1TDCgvvO
ckbok6nSHW9ZWLrkpV04/PTihaUdu+7Qvsk+w4bW+N7ii7KcGAmBXJoLRrIuaL/TjrbVTRth9cd3
Dvitr/IDPaY+rT1Rfft8ag2Qb2iyKo5bDssuaPtJn7W4UeTwdfiFIoJgwvIwqzlQrsFiTlOgO/ja
sNBpX8ysx3WgEe2Vhous0B0CZDt6D4PqBclGDjTVE1yA/Urwc7l2ISCKWQbCnmEjfqD7GIuXFHKE
htPQOTFRq/izA/DcZTSQ1yp68a6OR/w6zrg9hzZcmUKlknpN5tL3qVTQIZuDhNZGfC+BTNC0ivan
mwT5WagFJ41TzQY1shd/21jmTClRa8PNxC0vSklvfqss6EinuIMaJ+LQDAr76+2jJVBroSPPZ94g
w+LbfP76CWpILl8xzzQz7k758kxNbpG7sOHYgzSaAp0v/NW4EA2ifFmva+wVwb/s25BxAVSU3wEA
W/kJlnM9y896WBb8SH8mt6ibt3lqaq/8tKOQdibL9q1IR/Wmqgm6S+pf8ixcjfMefNMAxIOmdrhb
P21ED7P5WqWzLddEsumM/H8SWYBVyhbjEldW8SkwW9lfCvoKuJE0pw1+c0Byyq8vsInSHQcgvdE5
cYQDQLgZGC/NvKgnW9ytGs4gwKdUhnqKcd9206HnGPqvQKEtWX93QzXHC4DiXqRy3zayROc3DwoF
EtqdYvqB+z8+SU3t0g1oSF43RYrZkhYCHbIG2Tjl+WSkBDEjU/YentYxgaNOwQq1uKwA3U/AUpF2
xi0eF+ZkrDTvE7mVBMnaeHurn7ypkVq8ml1z7zDZEGhuTOOYdlzefiUR9OrDOClEUyE8Y9jHAQY/
psPSAV3TgWa0AdJszKzxai3apUDlUFJzsqcSx0xNVU31tPCMi0mp5oth3Y0WvXPHzhhEpx6ETDBE
wky1UNVVhkRw0/eRBt/xoDNplU83Z6aLocNqPMC0LEvfV7AV8XBgzOLbKAlQmIOCWrewrsfdROsd
8ezdqRp4DRskFBPrt4drVbv8ZZ19MhPm573Koj7yHOEB6i0EB/T/j7ZXvC/f7EAiH09JvQ7FVKTr
xAAuaUQUBo2XaTU9zMCJH5nHB5wkYunxHL41Cs+bSzqqg36LtGf6GC2ETX0tZ+x8UUCdnayumjrN
G8YlRhcKE3GrjKrNjyaQ6cLC+bul7KB62Doz+vK1JT5X33Q7VMyIiBS39xQC3QUr+VZf8IVoRApw
6lJbwMhP5lJeFy+4bndDhFe/JNuXS5u5oYRqNYIzMuWGcq0lE0FvCZ68Gf0/uO/L9t12okNnSBg0
vHpiML7yRHZW9qMhstZWqkjq1eBmOgVOCaVlc+/Oszyce7DIVdXJjjSE1o7BOPkSaHzwf1aNQ3iV
rJEFzo5VqO6AurpRnSOULuuK+EnutIf/4Gp8NMwMnbW4TBQrN66jUInoSy0biAosT8WpvhezE5q+
P7DLedSTh6N9qh+j0iwMtwskRQM+shyeKMxHru7j9kMuFFJOGVe5lltFJBT4aj358siRjjXo1giY
Wy6wr7gCOLhImNFuikd10jF5wyWze4tsmeXxD9/8sr1lGDPKxZsIOyBlq1lj8uFREVXEYZq6OhWZ
SLG64axsXuap17XLr9vdmBM5q5QBLbPovNSfiGgg3eJfTqcO0+izdrrVLwfCwcPzJlhTqCz12A8c
D1Wu0VUory01iVjqyAwqcU+yoEQ4NWYFi7l7hFOXPBQv3RzEQfdBgslIJVjapaYBzdr0WMvwJRnX
zcUH41QELXPDIUVaQr4fYig6rYWgVY+WcZUv7hLqUc9pUAHZ1eHZoVedZBCssMOWRh/kzkNAMfvb
eCD9I6gxoBgtuxcYEGrXMCzNSD0wVHYR4C3dj1kMhzqceULE+W4JOv+oo9lAIgMyQ+J9xLAcMgSJ
kMLWBRPQCnuy4oOa4Ey+0VRkRyEvVZCtRbPKcf6dODsVHm3TuCApq1X63UkC64n+ai1cTcz5jUgf
zhArGxsXgE8lXKEnKnyfKeFGhmUkMGAq1US4I+MDyrGYCONJypxXDzBk2aqunj2pBWDA9lGujMiB
fvdMuAtp6gacLPmRIWX6kJcEz4SIga1K8/Yv6St9WIFChwM33//lzg0PILF/xNeR4ZzK+Die/reP
gTSAwM87Lw/nc4sL5Sh32UXskO1gUAswgXVLpFmU2MjglM0WzMtyhYhoN76/IawSWh0gdvGxrY3c
+/NVWhBW9QGGyhUVDRBUlzsIZzkcyQgl6ePVuPCunq+E9BNbQeRAeIyZCIaki9J5k86E/sCVH3+a
Ymk0o56dRjwYU+sVyDWYaoXBcwLONaMoRSDg4XObg9dA8Pa9Gqj6UbmU1EGS1q3oPEmWnVpp9/oj
sETq/j69Al8XszgyYfxdHXLTAOzi/jAEeOsH+YgamWUJPfqKtUvxE97goxln92mBbduHw5bEWhGZ
cMNneWladnj2OHqN0TAv+m5qTPkjcQphuXL8aLKcGtCTcSkPKj8PowRdQnVex6X7Udu+IMvU3sWl
YzgMCXUx2r6rD+WdSg38bDRycIMD/dVJRUub0EPNabSYBRTSQqg/n34B5pp03xKptIOIwcY4P5De
pkvQkvBmUQmdEb4zYDzJLcsguubmHtkRXf4wVCdaUHu74TS5i2Lvn4/sbVT1GhYes5FYrN1P49RP
Mco5W4wvIxipeH3Lym1YVGibE9LTo3Y5ioexf5D2cVwo9IVESn3tqwhTq6UWw56cjuaFBr5dp5oe
kWcqozbIU6CcaX3F4HuhyhnKHIy4Lfc6G1hSlMvyh3C3hE4472liym0Z0+QGUCH3Mf+NnnrwPY1A
i4FX3AL6E+f4V/wvwiHBA+SwUGtFYdmhHZ/SaufZLPOw7XjHZkCQbH/SdLDsBRIeWIKmuVUKMFME
CPzG3v+qvD+GDKllrzLbC7au3YO36gCKHcAH6X+TPiJh0Zx57VuhyhP1yzfD9dj39Pkf0pBmCf+f
7DZMm1kYKyMM7qss3JqdTcS3F176wESpdLsLbC8MPP9YZT5JeJQnpD07rrtcZhMX1KdW3WXR1EqD
A5xCYs+mwGW6X3vneaZnBvwN5gCMh/90+eaqzGJ94oN+xYDg4na1Uja1voSeBwDewtyAGM8uVsZe
hCzhObeo+Sa8eKAU/98SvAIo3KOTYU+KBj6p+zd/yasL07lN7COHnpS9HaIHPG4tk13r9/g4AEz5
6N2ahLzulSvTC5qWnHFFfFn9aucIICUV9p3Gy1yo1rgDekVg1B6t10mRC5I8A5OwF9ZESn2vSWnq
EeD4ieYbkr696VNy989/PVVvjjtPR/Jd7FgGvwiyEPwCYgtc7xUf/aaJfGirAs6jot3IjEULVG07
BfbE0guIuN+D5rOTR2gFCJfDLUVLq0/L63uPUPcYabxfuk3BBC0pWNPXTYVCLekGHX7AUGbuhG+u
QLFsc7GkUZQdkM6Srk+8PuuYFGZ5nKcmBReEbYNhR2Qd7gPY+iRxV79b7FyA0dQF1lEmYsLJF5p0
qf7+vVu1rxnboc+JXPw3WuqDgiS4JX2jEkEiAZSnDSDb+k49KbN45OrVCduNhTKHBBXmOqziZe6D
zxAWg1bT40SuHLSIi7/qX8OKAQ/3Z3STEZhICjLJSRjeOynTD/FLU0/oSw3LHY/8J2pwoRkgK8+O
tinVsFm23cYfmfjIy7XJlhbAriavhGwW0TYcOttcUKcM/4XtUuNJ69mRAlb6BOD3dpRt7auyFYuZ
Xzpyni4kcsM9lPZ4ODFJHsUVUiHak7WQO1upxPJ07C2o4xs2KzM/ISk+UVccdWAyTB4IilCs5x+r
+cWgqTT54qO7fwOEEOvtoPLcXWJLxy1lQyWxG7GbUPXUfJQEauJcDnAKXpWM24hm54G8qn/XHGKu
IgUVpm3OB+6wQuGs6X3ngO+oJc73bDPIarDBeoaHbMuFgXpLnVTHvj0uORmhHxM0N+7/znN5TKZ9
MRoIPuq9if4M8yucHsQ1lmHEK9g7Ou5prp/DzbLGwjAF2ay7+XmViMcgHu0OamFvmp87KT6DSmWK
7MHG1h1sMbh4E/ajaFf3Vpr+RVe0BBddpZTvlj+tPB27LNEx23eFSVFljwPlqwzUdOOJtUp39yTT
3hOJMv5sABONk7nxCubQah6k+eFuQ3NZNHMvcIraKcyQUY4+UJlXUvjOpj27M6UerHIl7NrCVl0x
qvmM+zYGA7K+ukwV3IF5G+ln7r8vkI9Sdp3PK6a8PlwLubkg+77No597qT4r0K+hMvJKumbAUH8S
mwLDcs1Cp5cP7fwlJaOc6dZXjwWhJGxR/eNVyzIIhQedfrdTg8amLJQjoqYjKPQtWXdHKs8DBdt4
LEX+JwqnfQUvfiGdbSVe9RFJy5W/3vV1OJE+lrqkbvfck+WA9NpuHzWDhh8upQnmS0vpBQWi9au8
ny/kpkr+/4XDEmaK5ETTRAvKw3pa1Ijk22OORtxn1HL8otnBf4gUs6bb15Nl2hC0afhXbdFxwigF
XTo9y+Z9R8sv5dHwM7NnMmypPOYKkyp9BvwZU4NwCi6PumxyaEvGJEfz/K2kgjVJe4zMlRShUdAa
3wAEInvtar6y1saszsgqOXf8iZEuwre1YdodiikCGHo2lwjC8h181LlkHWutCLJCB/eQSnqLj6Vd
uIlN0kZNKQ7H335cACAWDWf8CDWx3HAaAhxaE2DxAFAW57ylbrX6KUnaUHEhHVoJXnwHzzqC6vLg
uLUCoi5aSXEfZBMgn0LmwdGHN2KJGqX+trkcI5jA15vEyyFf0LcTjNcMQ1k2q14ZVgb4ybuOKs6Z
k1Amdeab/OdTm8DvQNvMvOX5uVtONFC/3bTY9eN1Os5scAwL4x3XxuBTTzzf4nI8SzPzUKjbUGDJ
ufLQWF+oFlQZZNwNfIp8pHIQbepL8ATdO+lQw3Ew3qciD71LLSOxOCX6oH6Q2FqgrquGdZpYivyK
bPnqSijVmd3mf8neB0QcSQmJEwbD68L9YJNG8to8ZXRQHHRcXXKPE5M3Bd1hm5VXmFdOPZtK8GkD
B73CrC/M6KV+8Xfc5/mC0b8pNVe4k2AlJJEKf0Rtl6zHgkOJ1y0pFXE15CNeZnYOTViGfxaVGpns
qITX0rGI83sHejgtx7gsJCRRCUsjXqFmoBOR7TBqolyn9b6n/2cdhhdlc2OFytJOa2jcLPb6khah
i7V1awXqwgADgYu8ThWiYOLlhwrVDjWMQGdzCOAQVhOV5iKVH10pu/wSC+vUIqCt7+h5dVFL1bvF
EcluzqAeBEW3edg0t/t78KoGMdfQCCMIRWGiAtGCf8+TK+vwcZAS2ExLIKBG37Busp88s2W/9kTi
tK4mSTRE5NxrkKTgrK/bYtcBp6MKa/get3NFHyRv6Mbki1VhwFkv7UC0YGaAEVKyX7aL0YlEHQrd
2B935neEtgkJwNtU5f2Fx/Gnankpsu+z6lckpP3jPsZgD01PgXfLwN9PHMC+lp0M+8C+jNYBBJJH
QHp8yLM5xk7mJiKiUWGiQE+aSXWLrUXoVBVG/zsGAkUMRH2PrQH4Daza3DLefBfDCXeQOGKjoaP4
NWG4v33EDFtbcA5B6vuOqeWLLIMcj/+LTkDbcN2B9Dj+YEFL9tqmFdpA3pbda3+ulVUSD/hJ/QiB
Yx/beStjt+/+G1hQdB+9LgBhQcDD2wmJKAyYwiFZB3yiE9PbZuTGwcPFsakoISyWp+CvRmAbiR0a
mAyxrZqIKedmT/tQD0xEB0vNNkgsUbuDPanTZotfbEi1dTMOZzs00dbYZf2RKF5Ud5Un42cTGPhA
nHZgIUCkjvpcfHbIh5LNSFQzi4x70mqOurFIxBYJSSRsb360v93Q6MNm12E7cb5Aeq8XhSpr0USH
qndRDbHFTWs+d4TBjM9+9k7V8rlNR5xSgACaANEST9Y000J9fyQ4hzByw29bWj6wUvJdELgA6b14
oqbbc8Qpuia1MVT+rgqNRDLFtE4Egb98+SGJV1szB60+xFFadgU6jeBGvcyIveJejT0bdtYHAA3V
0sxgVCTk9keu7GLFulkvw5MHpwrJ7rH9b8mhr+xEArveNqqsExtbjRtv+mqL7GjjfRELJGeEODaj
V7S4C35fS28L0FRapkrfMNvFP/gc/cQ3Po1GHzisdIqSRx9WC53QIdygmMVL8IoR0dK7E7GCvpGv
vZajo+PhTAL0IujBQ1hF9SavR5vWAmoBbcukVh2vUoSdo6lbuj9mxS3iIhPFdNbxOxb4qM/c09pP
F3gI3MXaYD3NvbwscNg8kViGw/LgmLbwviwdSJIl+Rr5qXYcakrjqUZ6NWSqyF5bSLdrYbyAI/mD
/N25er8xsHtHGvSsld2m6qFIWR6Sx/gFgqQqv5Kc+VkyUJooFeGc2PhsHoghu+EBIi0bJ8nWKaJl
iqC2tp+SJyJ1yXMEnFWkFraJojiLW9Pk9z8PGb6wHAg1a5A/w0aRYeorjXNnueZ9yOZA3zNJnjNp
ZpVlMrcMTgzSCX86yDsJjqBjeiAB/IxigEMBkL6c2sZbATpS5tFYmP8ZkOnlhbq4LNwWCkulIvEv
nbmIonYegA/gvHrXEpHH02PvmBdkXXOwQNKFSZhBXJCMb/GTiKoF3tQvDOM33DTzZ5dVTFG4y5Xd
+PEXTqmYNr8jiZ2mqKs5ycczHHuKd3TnzS7nVTFesB9RmtwlowVmqEmtcAq8UrHmixvO4NwusCE5
95wiF6dtwjB8FU/r40t7zDN8dTeg8ghVOxqEIt0J4cKXyTccbiON1Y7pOkH32M8ycu8BjTIDMT5v
5i/xA+oKtpPphtPaxXzBzjocbctsPqGd8B8r64PEGUlncA4PYuLpR1fD9EsJAe0AAnx+xyCU+ec1
tyFn2e5YcszOFQ2wxSACxKEjpvrJq2/arBbdOKzCQH2xO+RWzkjtauNKjOwwebr7xgJlOh2zshLP
Y2XrqZzvllMFV6ucg8LKRWwdQ0Y+m0WhY6WHpYvsdQs3q7L01mQJhZ0/I6Wr16Gsa4kzSSWvmR3n
7tPG07LLMFKfAf56t8GssuCkqBWBnptP28xmCS3VgpfAADRCW95aIV4S7tmJwxoIAQdeCeiUUtQa
sPAQY1MDfy6Z/5FT30k4dmZ/k41b5pXUpMromirhiDPdzRPQUlAYP5ePzNv5aci3efKGo6z1OLZC
sYduPMDrtvs2T0jQgVCAbYwE6/sXxrkVNH6cP9qNOLi9YP/Z6HS4lrc5Scd0vhickq7o+D97jNRO
2ZHYFjdlK7wz8c2h746Im/Hkjd6CYh/8k0JO2iyYZvpFBBIy+QAWeOr6FHaU6z/lQVERhifcSXxR
Bx+7kfpIKU+e3QetAYrxd9H3ZFOlSytbuhLLn1munS2gqEJ9MS8QEHS6EzQZugiTiC3ym9IDupfG
b3xOnVf+GkzZSS0UC+bcJqkkEmikmMKSyD56EdGAskRAIYu8zyQoU41v8jvliM6Xl8kXE4omnwdL
A/lHPCeUloukuEt1imJkTWFa2+1FxlF94aUK1UVI8AcavdyvAuZlnA7LW3bP3iiBan2aOqkSfQh4
ANZBSC6h4nxMEg61YXUYppjn5mgODlpoMzsdoBvMX1Grt2EJKqKWy6X/NumX1ixKD6xsKsg8C5T1
dbfvshbpLz62bV1UO9pnlChJ5yonszvlNfjfhxspOzh6+BP/+eVnKhZKasEuBFUvnYheX58amL0C
kiCMNQbi9Yo3OlE77wRkfWubGtofsLbn99GhPnqaPnacusmJoNM837/O9GwdPynsGtQuBnPfCmMR
x0uM81tYd5dwglWhQDx+RTR/MhafggyMAixwFgBNmzhpeOxwm+GmHtRmRShsfkccr6yy7WqjCqxH
0391MXIEGE3wsVum7HcC5/K4ZBgk3h24ebFyb0l9xq6nzvh6rdtxiW60GyWkemaen4hmGZloX4A7
uhIGmO7DuFi6NG2SBBR1nL7Ml2CXLCVlzALAgwV04wy9OcLq1xyMjCKLAkLJJ0aO/ZdV8RDTkV6q
SrKR81lMzkoiMv0dgffDx6zSsPG/PuZjRs+weKtvJtc0pjju6r8ZwdCc+MxzZpWESrGc2gXTrPjL
0twsBjHon7qPvvMfSNir9rqCb4VoLoEKQZ807TzQisUmZwdsEhJ1kS+FurcirswQ28NsiKwklUHV
w9rp7hBaBtYicrYIqx4XFDNXqNJfr7oFJWGFpFuSUU3xJSzm+SSM3rrViWHBAVHRGaV6IwTHS1Ry
cfXaE6jq5fhh6vUCaK2cQhbIrsOY2XSMVM3i1wxj5b6K9Re6rtoFm8Qjr5V9YMMCnqtzazu9P9qy
RhPLax8giktEt9D3SWTpUCZgPR7jtei7hFgSiJ9QSQ8DMWMiwSKAso+aY9YhHwhKj1IApVfIfXip
8usZ5xB6cZop8BfCv6D2KaZkt/w8O1lqzwncV03hIr+cI/CCylvtWFpnt1knaz/hzyqxSB7UcdQy
hpZQl9CdIb7uhegrhx7jLKLuqXmBjNgmL4QevwzXWmV6weZApLEkYIiP0EXn48iETUaNzTHjLezW
Q/gLPnDQ9KcbGZSRDorMi+aC+GqOoph1NaMxi6OmA1aYG9+4g12bNl9TTprzx6PdcxrvgmmU6hQI
X8JFrt0Z8+x4FgmmLWLPihn1v9H1spYV1/tr4ADignx9q+Yw+my8jWV0Zp+0TOkDY+mO97ckKEmP
isgkiMDFpaj3sHi3SMl0jFxKsCbFnkiccOo2jnxyzaikxo6/xFgYj4oiMiQdKJJtSnY76K0bYjFz
k8BNRlBuH97faht488JszJQW9XqTB34osPZ1y6pk3AylL7Q8eawwpbhlCq82aMULZZhKm7PFHNvB
0+DlBND0+nMrmSA+rFPmboY8tGYDRmnBNlm8ww76x1O9gokJ1dWW9WmzovAFsNk5yspXPvbC6maG
yy4D/FGNiUcA8qg6v3LF4l9Hra0FWm1UrmPeVyzUznRyptqPJq1jfhQelWc/fi8yOiuDEbdxr231
LX4zQwITr2Puq+4IILUEQ8hMepImeN6zDZW+gLdVbwawCYnOTuPcCPYsIk4vGc8wvKS2MnauxhHZ
lwnZ+DJMgqejkqVOe19DgburEIunc7UEMDk4GrvRbtHILwEYP8oqy1Hff/NZBKPgn2mf8izrNWlE
MKcrgT3XJTMc3MItyhiEEQyVHGBcivrHAStyxUb8GxC+lHyOY3CRDg8yBqeWas4VKynO4mwvzKtT
uP6MHvXElkROdzfbjK7fs0R5qKPdhGlISZqDb6OD3csDZXFLUsomktmQya9t0nWeIPm4OB0vc6Tx
owuK1z8W5cvq9mSCBCq5ViXm2MSnw7JqYLW7w9YPtTRMQGZgjhGHGQPvO0Sn+SwgYYDUWmGWNBzH
nlPz76WvOi543nTEaz2SE26N2B2ZeUA03f/+e83Z33KPbsEo7wzmw6i461garE9kzyql/5Xz7cPU
P8VsK/Iwsizt9n6OPeYKQ6GnQLNHdOlxXkRcWzrBp93wqvm/H7ikFyOScV+L8aK3aGwzb/uvzTiI
kwTlprOsh27zfe0e8bW6lV6EHNbfA09LXQDWOjzNwBb/h3XDiItdSzWj37T78shlvoyJRx3xaru0
MS8MFg5ZSDomytccDEJi759vZSzFctULYMtrNQ205yXBgbGeYm09dUThitRj47N2b2gFuGyn9Efg
YeekrB+ohWugkoHmbCdMUNONYP80+0W8ImNdiiqzkp3paeAioFSS1T8ZwT0mretFmrUKyANlRpH9
lEwolLqeqZK5dNIzZPP8s7GiYWtt03c0Hwi9s9gzRYN1LGoqZxGLzFPraVDQgwxUSbJesq/Jn+4K
ORphQ5Hpi9irQSdUBFSIDjb0buHx9d2fZE+Fgqa7d6XrP6Vvh78Zs6i82AxEZWeH3H0KUS2pfV92
/yET16nSTPO7ccOUjYRqEBIhwXDx16tHApEKVeEXKGRYiPis5hmU2EJ1aj+6OSlFdkCJsA8dFHXW
bv85bTQRpqbTLeOQVd5HEHxVxBP8t8Hq5aajk0xQK5bZnHOi2H8Vg1Gk54IXr579+IyJU1yYSLBS
uwIf43FhmmKQ1dhjSVA5jQWIjrzrapYklj2dy20WbjasQXIF6U45GrZ7Xsc3+9wvi2atyAJ0vEbn
ryAjVcumhSt3eh7ThJDjeyEW2j+7zte1h3kjQCEhGLPtFqpMwy2vePNo9J9I2RLxgzspW9T/WkqV
dMYPyaB4lHTJI2ZWKPV10J8dYUysI1t1CPozGmXhR8KU3wzSQx47xq1d3NfIvEHMFN6N+yp9gKQ1
nzSXxRYKbT7AEDMHexXR7kHyPGeP/7PjKz5tRct7XxNM2DfD90EJukDFBHzEZJ6I1vhVOeteabsT
WpBaknkHiWnu1zKiSc8CwStbYP9bgGKyhPe4utTVwi27ncpjOX4wXITmf4r91DBsXricYx4w9d8d
YSoEm+emHVKQqyrAZxOfijSd6utBriTFs24pnUR1kFC/fSXyjl/9EnGRJcoUe6gjOJTFA/Dz6l+K
tlhpHwicH0ihOdAMKHWOUke72TUBFhjIy85GFYS9atPjDXdpf9jGU0DnBoYTsflhdz/GdSj7rH2l
/nT3PcnEODMPQ4BytiumOLckcndS5k7HJ7nUubfvol37nh/KlcDkITZbFQdCCqN5QzT+HmV/NYS/
R5LhBrcTIC2JZTABJ+aKRm9PfVatRsTKt8rxmv7T/rJtrbeovCUsxLF6eWenU1/HM7CWOXugvHjD
e77ulEgNSunqMIcA3AKNC/0mwBH0T4nvlJQowlKTPnmy7i+4uHqVk2o0lxAM1n5rKn8xwlmRmpJA
Iv5rZB39HKB6djm+rW8rt2kcocy01b55Ioi2KX11sxegZ81lIInLqXlyI4beIJyQDKZm/4jSC2BD
ejuMVKSAItvophTRNc8zjXTew5rMP/kqMcsxTTrQswIu2ggHMcL3kFPN5tcX/+x0dKrMU2Y3Do1u
QIoqEj15c+OXFGvzy0xN2Qc3ye0oTmyuWtheiIIsLr11UoMO48WE1qfRISpgB5v1r1FAk+yskZGU
hQYR3uqnRSHPnJoJfrsKKwybTFEDzYpiUChRSv0L070aZYIzsaqpYhZj9Z9Q97LX1oYnHhjTEmUl
WBvLTDBKpdWrlC3/wpqd0KDSvj3dMXXqqtT0k+25KdvH5ia56ymVxoXNEy+9W91+QTOkAsGdXUVk
3ZoxnWc4J/S3x3g6kSL7HkEBV5PpoZi0ZBzdi8qrnF9ScCCcmD3brcDWMLnYMHTS3dfguSQD6Ja3
ed80FWaFoAYbhdENa9vCxsdRxvsw6j9P9TcKwj9NWHb7PWxuOGxKW+MnV3B97jaew4KrStu39FlG
ho09txDc6cc2q960u7mNYR0VtfshijeseXYvBnQmxdm+4G+Z936E2QA4nSg9lEbxKT5PqwaO46NM
VPMfxPyMs4ghG2OlAgfwzGHceGGfqfItVzDmoZ1KTmv2YI6Loyb5ODv3YrSqDMcnqqyILT4KjcON
/T5rydVbSwzFK02AbNxZQLP9gozSrkBtv0OESXsmhAtWMvKb3ULKsrbgQ5pZcJH8E9EUQmK2AZad
TlQYWR8poGjBxaspCOFYUfvyaGdjEEl0CgkPMSnHfkAuFIHHJMDHPa/Vnrz3oWohkTIKFrYtqPPW
LX0wUAN0FnglIbeNha1AgWrXBhiPyECrl668AiKWLGV78JGmyNzb9+3Fy9kR6F3+EPKnnhGuqiHM
d++IwSFRA82HGrwoH8YGIzcfI4acuwr0D2gYtHzFH/OPHbN4zlO0rJ2jXCwQhB1oV8OJzblVA7VW
87qZyOt39DhUiHke5fUKZ93ET1own/aOU5BNbGtI7434Ie68nOnZd7yql1Y0Ry4LRmrM4OEiP8ms
FNHlf9dqLTyqXxFvd4aHtRyuzx7uhtDCkU093vexvYl8Rpd7bf1XBoq9dk3XcEQ9gQ3y5C69JHGO
R8EO+b0Yp8AL7ttSkaUWVK2GnCiMbgpc+ywncX4o2wa9AntS5lVsItJxw0af6jOttcFeGkjQovcM
EL24EHiq6iyUrcqINfLBMvv/7XKrGNvNtiHBMnnKZgFoM49ml9OSFO1/Eij19pfuzA/4taQq4m/k
y4TQsub25zZDm7TJUokybXU1TTjJamemt1kR53fui4BcfiTUe+CQJbq/5uZI5zQO3/9hLS9bhMUW
Zm0lrRcSq5oYQl/pY5++JIeNlt/+zRziJZxxCHg9AuzgQFOA8AfzTVZC2LMpo9hWVVfzfmg/aTEN
z3kqUVS1HcT2bQH34DvOKMZTT2j+CXjq+ORpje2WETqpeVp9EWk/J8CY/bH7w4e3VPvgYNozAw9S
9PuyjPay+JhvswJtJ4zUpMg6OBOrfvx2d5OEDbJZW1/H9JPBxeUxudBcyyWowbEGaRUPaGpvpgQ1
WLG7RNQX04tRD6PC1RPrUZAMGvgpU0Z5x9t5XNKPjKv/nVlT0RDaJojUhV9kPCgylLiSo+2jDx/P
MljGB5i/hljP/7dq/eVaJUoMTkbEFyUFOpKz1mkfpzMkWrDjzH4Ze0/maXA07f9dJlbpFm+CwPKr
NmY6F8xBOxVqZgsYc5EjFV4q4ltEHqAMTnFbnpKzef7+S8KN0PCfZB3KOpVqV3KejRtIWmEd/7xU
/jSpNcrSGE31QP0kcToDn4shHNIDmw8qoDP0MZH53s2orr3O+LD/evWG/0pOSRCWXD5jSW6MIYL9
8QoLFo0xDcscPHTLtga0JnWhfPmjKa02aV9/U1YQWgxgVPfMDW11/fhR76mg/hYwSmVYTqXW+nNY
YJ6el9oiRDlqajyeKiK+qj/Hp1nKaijqYBqiEhEq6oc4D0pHICWlEEi7WfI6jR2p0g1VDnJFN93J
J4mow9G8hPDMAl5jSQHP9EICeGu6Ttv3L4fXrkGEEGQevxfcyaPl5Sw1BYLkp+919/8YZzFWY6oT
25GYNHRAzipu6/BjEgP1T1i6I7Fmn5T9f6eKFGIiq1Xj1efNumqnyeMbAqy2eD11MXamKfxvN9qF
lwlcuGSGIklMhTgrOyxsITM7ipnZpaIrMxsH8BHRFOUIQ5IAtCzkUogOTf0xNhUYIWlUl1bGvYxh
Wq6c5P/sZ0FyBOMf9o+wT4YPG457SdxSOg5V3yR1U/pYBony60Mn8Kr9VxqCj9oyMCyK2xILzjVL
qjow9TnNVzCdvlAuVH0EXLB2gHDRFJ3UHy5aa/Q2guDY4ee23sC89d6xduRvREtH5zCKjfhk3p8P
wZ7hjl8ab77AQZfX8+e4bq6Tdc6vpzJ66K5zijFWvwRRFFvEpVWsXmdavD7/I/ZhH9fuQ8iP7E+X
0r4x6s3W745oFUTrYdJKQp8OxkDY+ZBrkBmfYYPzMjJSsF+q2dsKncuXAOv61C68nBKzHz8X1tz2
xqGbb3EhJvsqOqGWz2OjIY+ZC8Jv51m+hi+LnTt2JH9h3dCt1cSkORbvy67y5cdpUIx3YrHKU9or
0mrkUfeSYoCMsSROhPO1UMHsta6gbs50wk6rouMM7mpP7hiX1lHz/b0lRXHmHaqMkTooeQiFc1Cc
6bIpErNx+XPOVffvV+mg9tDes4OIVqqTDfNlPdF34KRN7K9QbLuyuQNl6yxJwhd4kvy4ya0sUqFZ
rfR2+dqe1+gUKLfdla0wJ4QaXq0bow/Ds4/xI/hMynnWfbG0bdR1m+r37uzGpM+C8nEbonocDAsB
NH/iKCNENCiXAbqV5+OleB/M7qXv1qp4Xb38GGUfc+HrEcfPJUJziaXagITMvAduvvnUUZoxAPLH
RgCPhzw872Na3OrdMeN5yT3yujV9Fwrha4hcZZ91+SfDPlnIduh6v7Ud5rJ3TQgKg1Q5ENWmrQJh
oSpKSv9zgubwkOkCjYBoHNAsZPCPqvNu/Y1Mv2Wq1bHsVuSINldYMIqkFAUGFPKarINgxetyP4tI
Dsojp4c+TPF7I6KK50cUWhvO2lj+TLCHyk1qbnheuqOAw6sHpd8EHjdB1qhKfP7tTztOxazJ17hY
QoaanCl4SujVQvSTU//G8XLnXecn5WllgOW5nisqI8awdOiWILj/kLVtHDn+cAMZNDA4rBPXIpkR
kxltX1uY8MFZJLaPuxnNhFzMfxO1r42O7vn4nxiu6+ePO23jV7+Rqi7alovyQ9r+GbyHcUriybsi
b4B5899h+sB18WakxMx181Jhf3yAMehOsRLhO8dtlhJTj6SDP8bLGUjdGV55NFWonDARt8fpBVEW
yo3/qgWQXWZtcJTodqwSumIPI98NTUMF4qD42XsVyyzh8KJr4R1fot/vH8qw6XR94cNlEwaUJArF
JKzeN9Fx2T45/J221sK3pZrnvS/vNa733pI7yW5CnnqNqqdvnSr1+Gn/Yys3FV2hRbGgYhkGpq1J
iezu8tt7joaZKp0tiYP6Wi2gFQR70a95lG84HjwWy1EBDjVDzl7tnOQpl8wzs8+AuswSA6mJH0re
I+5zqUIjQPMgXM5mnE1ejGoyIr/mV+s0wZEIQSuXL5YV+Bgal7pu1/uHTVraqxo1HtGPD4E8vptt
GKUARQmYhzr8FrtjZ0iBuhhvzhtZw2NBafXNo55LoKIlvLI6HXwbT6SRvN7ehB9E+itfBNvoKPuX
tzCOxLnlE6E0JMhhHzXKE9okVmNn2eTA2n5VXlfJEfzz+67cw2UdL3M/2hpj7Wc2vadXyPx7BLmG
xJLxBJ9UKlmkVYdNZya0BpY3cPdObUhZJy4YKL/NY7CLqk3TvSl9lrBqZDYmRts1U9aQQPunZqQV
dUyMz5pG/YH3YEfxsYdtBnWC1XmlJRFZXFj+lyHSuT5FVwNaixdmexfzOwWbeUjwRKjqKW9LetMH
IquTjy8l4MFA/FJpvWjCkHNNlzkKc8r3ghfcE6LW6zoQFIXpLys4qV15nXcs/5cYkffTBU+gce4y
P4fDnjmNamdmCHyhm+89OXclnG/8ArXvtDp3inJPdC0+Rr+YjDqOWrcWgrtbVCgEwJRxknN9X0OE
qNQVeiq6iJs+Rq8etxBuhHclvq7KYwXilIPYzFoZ/JPJ2M904QjzCLAnn240ikgyHYHpCvy5ZPuS
ytgsWjkA/PEWRMXNb4FCd4vLCWZnNqHzLTmmWUJeqkVARsuHcOGTNucguoecje+NVsNyXnNMgU3q
0KKfqm2SooUHglNjD16qidhpxtbT8RXpBvDQqe1sqTDrIBLolpNe64lh+Hdek4NwM081puCcZ6uv
XFh/kYT8CwIt5PgbqWlPrskSAOnk/foFMFjtWXYsu3T+KeCoXAeswafHnYYm/9jctWUqw45nrDpq
QlyLAe1wUs3i4S7snHw5wNjJ4ynji2fWl4fvbX9wBjoiSf0gaR7HG+3g/BcExJJFzbYVt39yH8VC
yDoZTdCyb7TwVsex+EjP9foiH06L2qvvhb3sGPFrI3ZP5U5Lgg4Z6+8jRCuXJm0vS4i7EctJiXBt
JBpZCVhRbig5EZTrGzkxv8MFLLq0+Z0ZrAUniG3GybqOaGvDqTMZoKHzPzHNLg4qZEqJyVQCBQj3
3nfN/8Ch9Y4f4FppXE4UPJKxLrlqBDnl94ayQO2zRS+kL6NAyDM8HsxrszkAynxZbgthrOi5q6zj
iAhTZodfy8cgBLW4OCajw+W2Is86Tt4D0Cz8MrlSayxqlbI3PgvnHl93N9JZoaL5Kigr+OJR3Nvn
7N19mb7zfqM3OGpMPwLpxrewqvkvkBP/l5fHzovGEgZqRptjrL9njLbC1iijX3Yjx40Fsli8wXuT
a4yZHslr9FSuLwOt3lBd4OusL0fDed0vD+7zn8Lme2ZXXZwJSgb6xAE/6PO44ql4gHZkXZqs6zZx
bSZvji2jAmNEpIx4bY9e8PGcPbyvMORLaLeWzqA4tAMlRBjyvdtW00Fhhr9HmA4IuiRABKwz9K6E
X3WALxuPomx5orUzA6euF5K/CeKYjuOFmb3ZDbyiqYQ4FoiSNUmetoJEW6iIzm9UZ1kmYWGPu4E1
e5lc0fv5hv+bvyp3Kw52p2sjK+2kc6j7Zt4R5gBe8Gz7C/1mcakTddWfwxWxl2T+w8LmnUhQqk9s
DE731tBvdY8KKwiz9zqb8oB7WvGOdp0jAIPmDlwx2dB57fry+KKQHeLLHZq7js749lyiCM7cBwwe
+LrKb9s78rIUNCKb6jx3jGZ08t8Y5XlzfE75t2HHPiO15j+G7i8LDP03R6Xupj+0q/Z5zRWj1cwS
cnEGEYmxmwLShwlqUtbyY0uvT7IBileEPTW/pj9nG11QPa1dcXrfNDr9rGh4Cy4mr74vwEzOH3iY
ffTphJ/0qnhbrB781cE68nmg9UehRMtv3n+KWeZwFW5QTaY4TPn9e7UGZ5tzUDbqQP/N1h/dXUdx
hJSNEd3worromERLAFB0g1zmDgDJMvvlltUjV3WVAv+C0P5Hunlz0EukL0Z7wLnHK1zS/shxFHp0
DS1Rnc3q20h3s4upxKY1y0j39ZMYg5zcZI6oZbUI+npOTsd/fOmAcIkiJs3E2qL0Dxwl2y32wF9I
p9ak7rVmTXIoaUGYSPw1xQww1XkcMAbgQmBjVR9gMiJ6Hpca6/TkqdiEI8cwKYVI0HUVtJEN3YHB
cb9uMaVeZ/UoZDksA79z9r7dFzd2kHOECjo0uzRuxqYA1A4OwwksCccVACMw2jTDvkhXrsml1Cr6
oG9176Sze4XJDzK13sd0280ITRp7NRKOjtTt3987F1jaENaccIUt0kxixJASj8QTubmHxI1c1QGV
TH6DVyIP5cCdyfI8nZhmiCsmgPLZXzXCZxIk84Yc7vo+ax/xR+K/WPtKJTEVYLgbDsbDsxFX6jqx
wuPb0Mxxk1quRpm4aCfhO61OpNI/1/EXRPNyNWzT7HAWKFE5ovzE6WAt0VXIy/KGWPS7zTIAXZfF
uJD5h0S2knPW3HNwY4jSbOYUaUVLrikB2pBIbvskFh7PU5q20IWgwo5NlbB8J8fGZy/rBZaA8VwX
zs5FA5Q7gy52cQNB/tRrOfSLI9QXCxr9NiuuJ1is++IH2D4iwbk/2m1KkKHbERMa0gsYtrGsRa7M
dBO5pTqLiFwvDHVI6VsYBx3jCVPupLMGvgZx68NkSBXKyjNqam9+A+BcZopdrZ+lWl6wdYL+IHFz
OSbDUPx2nK5b8TfPC7nJ/ShQs3sHxGWJXrOJvGJ4IEfOXLH3uBTbkEv12xdaQp6HI0vV/moM+PJk
oUTTVncG3k2+wJmpo+pNMCxo5F1Fo+YlZ9uIP/9kJKp0sQsGPs+SR0tRazSUQuTDnfMGw0sed/Sk
ShnMMHsdKks4gyzVCOUYCzykc3ZSDVZZPATK8ZmlQABcVMJ1AKzt3OuKjD/+lWgPbnQ7284+Dx2M
8RYt2tAcNeADwKv8X82ERvFpKaItQ7UhBKgg141o6sPHzrt3e/QwzsMO1FDbHc/SoNK9RIfs/Xsx
AUbCwIHYIcTMAU6SIV2cgCdzw+WdAAcx+wXxcd1tpoee3H2H8ywE7tZTGDs+eh1sBB5QMMJ2ZerG
FrlJ/esGpWr/M8ZiD2nH3ED8S8W5W33mXX5qSuF6GEjDa/6dLxO34c2Bnbr0DlMcL6j7QFRZpUKK
GU3tj0rTj7HGVU3oGuTcuWE+nwDxclh2NLMPprAcokGiYGb/004FiKSmixfP+Kl1h62Ev35a+7Ft
bPV8Qzi1oatYr+hYjzrwvI+4SwLcABTbnRetor0DiTnqIUamMRJwT16Nn5O4HhRL7A1jY8T/yp26
BQeu06efsOjo/2NJDB65nWWE5qM8XqsnQ93rBHJ0Kz8GYQd0/H+O7QVYcQKKk1xKI+set3oX90wY
UQO61EVSCEd84iLfEVESyhKicwKCr9elOqqdMhWIpwFN/7iRkF2CGtCjgxU3PtRXoGD7m23oVfL5
SFkxat41UrioRZYHct68n/ZPCX+RShcniaiXBJi9PyProgYzJEu7G46vdWW+FC4rJiftEj6nLWxW
PzqqbX/MkBbxZ9yfLJ/ppo2yCiwZaVcpFjc18iXoZjUMMrLDdgZfNnjdLVLbrlSyrTGyhcXodOcc
pddsAd8rIn0LXxdeWYlMvDNDPx/xIGTPlPQ39l0y4Cv84wzyLkDTiC3dTZXQGgdPQuwEEh3SyJh4
WRNn08wThbmZJIka1Hm1uaO7onjhnnHHGh/sjh/VsuOd5si3l9RTkhfUcfDDyKODfAgg0rKxsQBr
zeziH3mWHsonSnb7zMPuXlbrWRtPbff9ECPO9BbGMokLCT97QnZ22hnRqArVtOtx1WrlsHdAn5y2
5fxKVnUecvv9rYtPxI6mKut4EPLgk/Scnr0b4G7EU4A6AskKyWAFhhgOkSoj5GruAKL4q9ey0kE3
0x/gcw9wXy+hGctpfaH0t8b5WaEwc9JPi35Tdfd1DyAv23davw3C5oEbaETK8PEjhPgneMdSrAVC
ztvXLtuz34EmvNM4ui4vAuJJU9JvMML5OW1v+r7xbIMQk50Vg4zfLU1WLRgoZNxDTAaiEeTO4Zkt
6XurU71vqZ/J3tIgZqiQsyQ3KooY/sXfQ4jYddd5SpX+osn4P+oj60pUma8IJzjfnv1sg45xTtK2
eD1HEObEOCyGvVhMAi+ieSLw7quZJkj5WZWNV75K+RSoXdDcjQ2DzKLsb1BLVpzjmgtMDdBrSeV/
ilPuyb3rxwl7ljd1Y7/2/C1RD2HEwb9y7KKtcgP9/sghm+Lo8DFcwwjglzpJpwJoKVydddQydD8r
wOXMjxSV9tSrBvdgIQ09QgO5Nw+ECvlAuBxQRK+WW8ZQMZPsayXhzosM61QiflOdrAPDIP2N9NgI
Mmrok5aJ0+Lz0A4iGgruUgcGFmjd4ttoRlRU9OBc4/qXdOd6j9MwuuHn+2tgFdtPZtiNq0SeBIWF
UBVqIUleR/Jhv5C2bmDyI+jDMVSf90xCrvHRYx0nmceQVZZDgeSU9JTUVZC6/MZ1A8ezb6LMfGWW
Bs7n1Q3UpbGeZPN0qSqaMw1McU238F3jp6qum60pkg9jUK2r/xdmCaDkwqngofZJ4WIGRiQ4VeZx
s6rVFkL8RhRgLJoWRQmTifiMUb/AEcS8jOVwl2NPj5x7ps0fERQ6+krQv7mVuOhFBku0DNaoynws
hQmsq+K9abQGDfBT9N+kjFzi0J6AgClZso8EPX1jtiKmoxi39XNAvOKyhd13pxe4NE6e1xJG1+sD
z1w4DM4PEhxhPHPQZrlxsf7StRbJHvh7UQyyyIC6mc14OFLt6+w/xH8AmQAAkhz/CRthHV+21SUI
Oz52MRsM4W5D7p3D9MN3X1n7RwNNiGayZlD/FBvdIcAm2girs5i39H9HfRPfsT9iNtwObWEAFhMD
7O/LX9nmAYJYwWBGVgOh/BWqD9n15C6E9zU0C2AUyXPszgYFGLKrX2DC8gUd8lbxzDgST2AsXQDx
tQLmsaXHB5NY5uGnFtkdMLL06fCBQMZfAyreqX/qFU9Ka35uR0VDXeApSKW5+EFNkareqIgQekf7
HhMblSdDVPfEcJlgu83s5OyggHfrKLeH3cP8lzLUP044oqjwdGtT2UaOG/4mc02lF5ADDnRQr+Kv
bYNJo6ytMgPU3sH+i7QrKX/2fz8HcgTzcH1TZp9gTwqIdACF7GvP5QQ+wNf5X9QUFdvUEnewzI8X
t0KGhF+LAIzdqfLzzsUvBlGp6wg7OF51sQu5CiBQtKSoO7nltVriYKiHK0Ru94cK5dFMy/1IkbhG
8uA8vrgprqZq2TwakNj8tYdPrwtqZUz7KAQDIo+YDxN7wAvOH2QvlotwwTzmeaRNsKx8AEK4TkK7
GZ7cu0Z8ZkmGVzUqaA6BpuNDMbMEcqgdpHDpaaccUskUk0htNiaX+4l+8klaGFgzBhhA7fr5w+D/
Uhac4SrQqL61gviwLboWyMiK7v9JEYMGpzWKO8YFB6pbNvBftPII+qFoME7MLtekxdVPUUzMJkmH
uAMrSnn95j17Vtc0ty60jnHadTXcNCX9IP6FGke3tGg1Jjgf5GHSxf4v+oM5PBx3YJVKzogafeUw
bNvxpTXLNdrhlPnUBbMXu27yMNILRLi8uNwjfNgDSyejpZsBEENcSoEPlApEKC1QDqLg45zjttp1
1Rp3MTU9U2M5ZrdqPcsO8fIjcEJ9oVEQt6OuC7uWye/VbWtmoAGuS3l/zg6D3X3OsGWXPqvaURuA
ve2iF6wwfAwaqXkle1s9aJheU4V2PN/CA9fVLCEfzyQ3R+aIQdEKfjrRf/y8fFt+JTL8t+umZ0qq
NZKLqIdk0PTb+j8I7oC047zLQxTmkdZqzY1ogN1PFA5ljCneQ84I6wiZ3wYdzdKlJYbuWKPtSnr/
mAEa04PGi3jXt5j7xiQ7XK2K5R1ZFmx7BLP8l8C/ZaJ1F75blOSHo0HjsJa6lfgiEElWGKvYCLMV
LrB3vsMWBa6jkyHYoquRn4dbui1t705qpjsMypWyI/26/jEEwPEFAOjLk7biVM72o3ZwlRH7B3br
j+cS/SbLAiz/kOZ0YhZkcwEtEAhbNSluevd2Cj8nZLxfmzIeIgegdnsigao6A5+jedVWyMIiHr77
yCjWR5Wc7aRjf6BkZNtvgVbNlAHW+9IuaWyw3LpuPrLrT5Z1ex9yvsXVzITK0apIEtwJgpectGsq
dV10fSCqBd4ITMpIJpfBoNCpenCO/JaZMV822Ea7ysmdw4fXaoBSFBVMec5ccw0vwQ0pRSleQMwH
b1WtSRINtM+Q5+hlGfnU0faOYtwQTayKYrIe0T0jwvTbTEBgu7y6FguQcRyogP/YbVm6aGj3BIzW
DR9ZC9o6n/X5+LwnhbZKkehHZlA7M1OAXNnCSlfhLombkqgnMo8gdMUyk8moVV/EZ5W2SifZVO6+
HRZ0i0wtqM0dKDKO99y4MVinEA0duZhR3URKYLtCrDRdebm2dZCmrcMwifZh0F7p+aTOhDu8gDGg
xn0qYM/ECUB/FSy69x8XX4Zk78mMhQHphyecFgRBqov1A6zdfKq1maAWE/IOczGbxHQiElxmPo5l
3kU3rm5nEHyUbZqF0+jNcKJQ6zLNfdbGF71l18u8wBP9ON9t0MWcLCG72JMLz4ZYYiHV75NoNYsK
rKJBW6tZ+HdBPDTVtrPupK/mLjPiq5H5QV2LiKLKm62o3uoMJibXsqAKaKUXDAVPJK/QLFWDmABH
wrwm9bNLt9f0sDixiM+SEQeQqZDePC6dLIwz+bHAP3rkLkO9oyI4Hk7KE6oXknw8Q/eBbl4KOgNC
9Y52GZotuDMsjbSY2aEvm4YDwbPQd2mmJkTq4V6LgIoiUnrtkbxq+5vnTIsWdbKPMFvpfen6fB3A
oYN0eUTR/1whON+yqj4euA8lSbUKMiJzx8aoEt1ZF8m+OCdg0OxGXIruDMIwVcFYUaqnGsxfVoLH
salD0tr49+KVAwkyOG3eas5C1eMbDJ6RnCNw/6Z5A2Ygc5siqua1v/bUFZWyVk7wUah9b5xppTkb
A3WVgGN5Z4Gjk7SzhaXWO97EOSYEi5RbcQDkhs2ucOJON4zzoV9jfKQUUzLC3S7EiP69+7qfww9v
ZHHfatglKgYbDWY9nAiuTjA8qLp0yWY6qIZhLgn1uTmK6zg3wZdg9hvc3pSC+hr4Zn7tInGSHUAx
x9gF6kKA5Xs9Ep3UeAItnkK9z9biB8YEMVd9XCpH3bgtrqY2HC2n5YstJOnBzuc2mCEVBWgLQpdh
7uPC8xsvYWXrcdpbzNaOfpMnJfJxkuJhOQ3nmGjAV2qsJoqSjs8XYjIUf9Jbl2Vu8HqDyhIrdTqk
kcNAvpgbxVfEz/xNJlifrYQlY2+zJ8BasdZ/yrjBVufLm65FtFTXXYbSuz1h/kaAHR4iWkjk565e
fVuqsIzrgtV6SZpjxENCqgCrBf359d7gsZUxvhz4dyFkFr9a6nPrQGdp4ndHH8qBZLet7ZYJ2Ch0
d4vB4+qutzZ5RjNFtJRjmRb4ynMQ3JdgBmFUxBUbzqzoFVnabm4Uxmdt9+PBbo6fw+st+zr02SQC
ksQgViNBwzpmuM+ju223TlAeh0PMXiHkIa6g1+T30dPzHLLl8o/ZQ7uG5BCLtBSUO7AkRd1bPYuE
aPYWHEdcBLQC47VFkxfpzOy/jr9i1ILTlJDSu8tTmvTi3eCvq3XNwJGxpLEQguW6V13JGwe9BikA
A9bVPY9r7P+j8RFLBOZ9GyxOt8wKnehZeIXJLkZc7mWYR5zfpdq3+VbFqmYhLIJBwcZm5JzQDKNs
4xKKtLnNujmP9G6QNBse0+E41tqyXrTIJmzjHoefPg8W5tnstQKQew3nAAos+iBO+p9f7713nKgl
vovlV3jugZCVpF/GxamLpA1HMFEdbMg9/tUq/7eHX1IK44zyAdIWSIxcfIYK6ReHod/FbG36M2hH
C8o5CxZFQvdr8/emelGus8WvS+CyIaDi3XjbmRyrBkpRAjSFVq2YT9cdBUxrP6F3kzWegGMzBhqw
PD9NdY/045OVWHjmlbc0hrZ9oWyyujD26/2MXd6jJjTuFnPx1n3M/IdnxR+qBoJzUmlRgEDCRysd
skEey1W7xz6rTjCc2f+2lhU9Muki/KbitT4ADHXmL0ZN9MlSa+8HbhSoGpalwVg9NoRSf40m5JVd
itPESVe5U07HCYOytGhHZl1/M8rf17oD17d+xYanoyJX6LVzGmL/aYOoI3UDVjw0Amm05Ub9KVH9
ZWgc1tfmKOPmIBNHdV4nNahnjMgqN+jhCQvWw4RpEy1U4F7VTnoLrG9CwG8O8bw1QcoEBr1+Nj1J
gqNXA9A79ZetMbCLin7kciGFtnqMURp/qyNmfHukrGNGnHuKxIJ+VzHt7AhcVE4ODyTo2bxZEyOp
5SDNpChD4e7fznFsT5B5lJSPFN/0XE4Ve6AEcxxOt88OaGYR8aUafrbUJ4rc1lGOPGcCr1VGDU48
G2VaQqfRqgIuEocjABL2sKBOSflypUpiyBW0R3ePGIzDcBKYqj8lwedXI+itJx15zPq7cFRbrbb6
ecBpwcnt4O3PAXnRztYMxtty4qKEHvraxoi5H0ekYZAeiWg/3Q74cp826AqriiNNsSZ2etsnuKEe
sIb+pt5aZMHwBLKZEt9iJJol6zN0beI+RJQK7HnBJZnqi0MNT2HMUcdNDiUdF+r+HKrsh94/z69B
UIwYiPZ79PdUNGwWQyOzBAQJacrq71klswSJgurgjMJ4tl5KH2397Uod8s0/HGMehlgqA7ndoafz
xJ1m3A0hXoULqsbf6pYJqtYoo8DasEF8EFwkm9iu4eYndRUPfjKGD1sv5jSLVvbdTx9ltCiLMdEj
sn6I+BLHR2lNihycLRoVY438RKGMdU5s61hkp3F7cE/Fc6xv35jMoD5AvXTWTnasI4DXAgrZwQDF
5Ol9pK013r6qnxH1phvs/eAy4iXb6GC1rYws4nJUuwtMBTpDsUMtSNVe+duixCH8kvjBrduyblNW
IUR0L5VKG63z1omKjcQOF9X6E1mlvu2WbKya3hj26xgoHwd+V+auG65eu/7XhvWC9CER0DrgtgRL
mzy1I0qiqNiCjueB2YgFxQabAoEGzbzkfqZ6DmQLcyW6uMFiIhNVWm60K2IJ/M+rDNId9V23UyHM
GzxE75ZzcNPjbqvmdwJrULZrituhjEFV9gfR0mk1cX/Ri2z0ftmiD/1Nz0l7ZMDS4/cr3cYOkxST
jjLXt1PXpzrwRgg5YnXs8/1go353T3F0BiS1HSz0KGyP2jBZeMkuZ3m5KUbWbc/C7Ru660axJGOI
46nMKn/75h3lr8+7GfjgSpx7Azg3PAp8w0yv2Gg9brbsF+42LQ/MG6DHn/LtRiIRnsJ6iPhVFiGA
Iw35A5Yz4G084/wwftVXZLM75G7hpoJzCISlME1YXNWLnFf6d1NKWy2jLbn0rzQ3U/OwaTwsVG+0
dIucdCEjiGct5okPDpSHy9oMnmBtaI0UzVRIX4mlvq4B2v/Ae7VmqleMc0L/kD9RKPvLjapUBwfa
p5ZaKO5ni1FzV/zSM7gI2oO2uI8e9Ixju++sG2dwGIFSid4fDRR1pROwwz7vV+S55tZSGVXdApK6
WblT0qWn89xXqbVkJRE5N82+orU1eG4BP9raiMq7hzUMhfY0IOHbSbuN5GpniisdGUlHi/Gl39La
nMj+nFcou1BVIYmHxWKMqgxo5vycS5dcW593oIqWNQLonvRHfrg/fPa3Io2aG9Bxj92nEKZ8vZbX
grP+EdXftoMlyUVwp9xnPw9HtcrxGgBq7EHxuRgnGLcQL9ykUNe3qE/CaLk6qLYMpcd3NSRFajUp
ogdxNrOg97hMFp7adWndN1z/6258GNEQerhTWJaVZ5HIEBJliU+t5AkBAYtJVbgtB/1WB0hT+j83
zEtNBbRQII96E7yloJC/I+SBralFKByhzdJMBBJmbh6Q1FdUVzT5U4lp9Gj6jAVCvTQjZJm6fwHE
BZHOBubZqkB9t15zvH0zzMpzw0TTufLrkubdfE1XJr8W8aFki3qYKOwi1cxmFTV/8+uBZnDuMZrf
okb6jXmqT3CmJrgKoX357cxfV2wWbR/w8quRqVl/kqNsQSVKUSZtl+MjHKoz5+sNRadNjZc+r4oW
yCQArU+h3fsg1YA+F1inlyvaGnWcdZ8LLZ8MMfN7Ko0Z/OSw6R+hSNwbA4vxlXlBF/N9qQga2df6
s6ld+MDa95+q1LQjnFnJptS9iGaj+NTtfisiDYez/cHMEdNDPx7Fc258jsqXmiTmZwZRySOjiCip
Ws9YIB6HP/FzLdW+/hxHm247ZrWef27oDcjk0AlpA2KRI47y7pNFtMOrxfgK1ROfOTPFJrq9bEOc
ZLiE4hcwttYhbvRIZCnlEGGvg5M2i9uGQCod9PUsTqgR7uYvBrgYrqD7zSMZCCimvfHHZNdksyr6
wA9FpuhhF68gPO/uFwNWaJL9INW5qrJbYvew+15D7Q9jQM1HjsBvzpbQdknuM0RvehItizem2wJj
ceBWZSW5tHJFY79ddLTGiG9jTMQMftx9P+AyVsx8ImCjjCTCPfGoaHJ3+R0XywrIz8Z0Fj+qdcHs
Q++jrm9jSu5rgakxdLWJE7095NFVBHsfrCYAIkNUyrp3PSbw0A8NuloMkSXYiaYMUDtiAe5q2R45
idTmBcPEDKLHDV/YuObE8EE6S/QNNtcmNBH15J5wde3ji77UjnsjbW/VYDD5GMic100KCKGoqL96
R6gT85fgBDiTz0FRTweFecm0xDKxl6DMeCNDQAHNId3kuAOxlT+Bp7bL23Fkpp+s70IXVL/JBXwY
TvVt2LT7PI6V8TP8BPu6aWkjAVdmwgDljX5Pqt56NHPrpjbahM3vWzo2oX7Yb1ngNWVANkg6L8b7
CFCnG1mq2Bx7tq45RZ+tSBAl83qILGQpOmbTa2Fkv4EUuarI8WnS/Ar+hiSlEze+gTACkyWqdn0V
lKJ++qxSEdSg+9w83q5mxVZZfOJPXrdb9Dx6l73hOFQBO0KZf68nP3Hdx5Fba9IIz+q4VqJyNJUW
wDUDu7PkBZ5+PHjH09cv9v8KeWN7/DRROJFgWr16ta28/LVBt5kyXOROE94C3Lx9EgFLurTyJTLB
5/s7SlbLVtJ/fWk+mrNvYUlnstPC+ue3DIgtUdG9pZhZ8NOAch0/68c7q6R8DNAUkdJn3Mv6Yh7X
j7LA1V+D5oPsG6XtS5rb1tJ4UgIHoUKLM1gQgwLiqXx5rb4uCMbKrdvJ+VgR3zWLdsRIpaqwJqBN
yBX0hHOuFkOVkGC0SDsdYdZJtFDkgpUR7Cy987DOdNG46WASYK0dovzF1aVeB/JGNg4tnYZEYp/o
gsO70cNJRmem+P6UBNrIa7SXhGtG03DT1oBCNuQMPnKtwg4NnkUMe0DYCo5Ap8wMAv9Kd3JFe7fI
ku33cTnBCM6C8eHcOjhJrv945uV/1ZgPuYH85QpIGq68tmmIbW4ifI9XL9fZtUb38RGqfS/zuPAR
wRqbpC/nAhItW2TwYxqA6P7f1nm+OJ6Jk5aBn68fdMS5JrBfo+jdoVeSuFJiuQ1/qbstKPOX3zHx
cqMTVujgr8DS/Crp9OO/uKUFL+98l71Boox8oRwIANaTiyCDeNh6jmCWelIwN8UR2ma0PQh1x5bx
vp6xi88LQkX3XRumOz1NnfhQFB4eu0KKT6Gk1Ti+0eltLls1own5x5C5ChoCmmgKfUNV9Pj3Ysuy
CrGSLADrb5yFfHJMgx4XRaq3J1M5pnOwHpeeiPnzzpjvOs9arFa9yvVD/C9NGK1SvB8YcIISp0Ym
gUfkFxZO46Vci/O58fTTThj1lPprjY9BB9dCFPgOZyFnHU0w/N02ie2iWtcOhG598WIQyaYt8NXU
NqeCCB0Oqd1UU6J2+7HeOgWTC4/1jnnvHfLEfbsrvMBnuOOT+9iU6BgXKjSfEcv7rISYST6Zy/ym
793Jr+VMfM5o6TzEYcOovwxpjptj/9fTEqdYzPMEeFAyP3j7WFJIlLy7G9PZ2vzZjb60yDpt0gde
VoL7BjaiMIsciCc5QJPB3R0kaHmgnpK7+GglsU8SBDR1XZNWWn0lhymQbe6WysVTkvvQlhpsLa9/
GbQcXEOkDR6oEUtG8POGn6IAZejQa52i1G9B7/q1CDTj8HStiar9L+P00N6RrRYEAIrIslyB3scm
iTm5Rb5p6Ewin43/D2W+AlzZL42Qpj5h9DeWcwWBZEpA6keEnnMeD+t+BBdA0Y0yY8Gol7rKX828
qmaudZ2N7CHbcFqXdyq15ZqiTnxtRsTPI1V/Jrr+WtGcCFoL6C1nBzgvwebLn5VcwOpDz8hoz6ju
r+slIVrBZRU8lmPASMeYtjm/FgjcGJC5Gx5G4nrVxr0sJhUj5JqxP27zCGdPCCzDUZ0ttStneCRn
VbT6RzpU9QEe6B8p3VDOysO5on2+4fPnqPA1w64iIrxp5wuI2IEWQsSpV1mh16MoQHiy9DHa6oe4
UYjAqWCSI7JC1AsrMJ0I6a3a0KDfzT495JLHKq4aD6I65Tgc7Ic34rnREqQx6saoMo9eSA70CXxL
99ABLSDufwhgFhmmF0UNaoFfpifyEMYp8/S58KJ2p8xkOfHiguMTl9CkU0SyA4mf+xY+d6G0XjUN
ExikmBSHc3xIeooom36bCOAjZ+VNJN6LmipAYPaBgV6HoWSQSOzjbjE2yGCKBfXfGPdlIzlqJasD
5zSyqFkYjHgsNuwnFGCPozf+5KkuZ3HbRSBX0hZ+/lF3vYp+ojyQPl904bnU/6nvCSmU1mmmi4aD
uRxyWjXTwtJCeLvMZ/Zy6EPUF78FHLnUlYkBrGkdbunVo3/8VCzu1A+rb6Rp2dOWotTLSQr3ytw5
4HFNvD2WM9aNvj5QLFaWdT5C2+EpPyqIAu3hQvfWDauzL76wxfG/QYWvtF87e3bUli5K4DZPdyfJ
m0zlDyfPXkiHi1zH5D9geQcASg0Rtcto5VYMfcS9U4qAdxdBIH99pIDj0fEpNFnWz7C0eXhu/2l5
ig8oaAdwxZ8Y1YcCkXsmDGt7BquQzNWOdGEnnUHWvT2FZGmfPGs/PeTbSCwNppw5SxWZuCz3F0Md
O0/CoQUmWJ3qFrzQDkZvyUG5s6zMH9nfKSnVaDyREl4pkIz7dVgNYs0rijg9ypYkrO2DpLEI+qQc
bYvrpYn4e4dgD7lQgw+1ZH/ec7YIQEeanxl5YXEGrV5GTaHA88H3zMr95o2juOKtZLlIUIx9JwPr
mL8FSkqx0Hrzh2yyAu5D8GUDMd6GM570k9zJLeR8Bcp4zIGNWyuNnfluPUfMFlMGAP24tpg9xHys
VvmVzOf1KnGw/bR58JFzUGg+CRG4G48BHgmvgcn4BkpnR3RbyFktD5lBWu3goBH+KaRTWezkO8B0
entgjWa0Wz8dCM4IcTwKl1CkSOvRmn/3OTKbKAT0nuKnLnPiaUOBe/nOmhMLcGGGcZy77SJ5qFly
cFQjwX2HxzBqvnyJsnYTEapdXtkQpGHlYrB9N+CnZFL1dSkoZPXD3rjt5QXUKxk/zdnD8owXbiG7
hwR9yAIfh+sxP36RJ5VdiFYDo+uYI3n/YVgJcq0G7WkGCpuobyBzQZlwpftmOygdp8HZc6QUCP2t
PKrFzrCmJKCgAQbIDtxd8+w9i8vnopzOWokf++ZBPKl8bVG6KmumqHKq089YL3bjFJr6xoK1xr7n
25phbQ7oexJq73KpQ4pXX8zGDug2fAnZUUBGnBrYBP+ftZXBc1bCV2BUi7tfxTLMJvwn709keFgi
Ykmz6z/R1AOaYszrV0O4RTIqm6/HPM3ePNGEe/lgyRe0lqCVSsbSFRPk3aRFF/frrHxxjn906iAj
BQ9M/JD1t+viQgz1lvP4DAQVdkjH3EPcF5E+rq7vNJib7uP7NwlkDxfspBo5eiCfH/hLnX04cKZM
Xc0xHDNfx+icEYhlBfvsSVYabAyAGUHplVAdyVoDnGrmdwdZ/+LtKr83i2f7P9JPwXTF2WOGgrVV
SCHt2FovE9Winjg9f7h0cZr4EK5Oj22sDr8mybCISI5/niLUqiMvUkhHf5O/CvhxPP9FT0Imle6n
3vd0S1KDQqlxJnm+7jIB71rV4bzOupvGku25aB1u+jLdItkhWcNayZtbZLpS+aphXWaOjL1zOOPI
cC9mPlLr6hcLCSAcYyOxQQVAH/4CmJFmijLI8wDxwac41GGCzRIOvg7Rv18NAW2vuYjyNg66M3nB
5r2WF4oAwbDc4eAUQG2E17oQQAiZWeyA0ryRfRP8Qyi4OHOjMKID9oIUm1G9WL9bRdvoaCUMWWza
eARh6Lpz+i3ipMiAeVXaGK5DkMgUa0fI7+MEofjz9dCRc7lhelPFUAqvW8k7T8BnCrdH//qnlO3m
12hw5z2hG4SZP7YDfch1Oz8sCTZOCE3NvBkPeX9b2SLQXEC05zd8hvhPobSV4eC914sAUu93PyMD
CxOdS6nNgkniYXC48SoclSDPu+GN9EUFOpTKtxvJDVTJg8aJhhSQN/pqB0sa7jCWD+a62BadR7b2
AAryYTHl/nehOk16ZSTfof4wCdc7KvZHqXi3edgjDAcE8GAzycPTgavcDmNq3WRCGwvCazxP8I1y
enyGh5x4b7ezy3ORgxf6q7m0FHAHchPTy5AEcZ3ITOmrmOLOgzjhpDBNJcQwRPyjB+4NbamxL0+k
Tz2eX46zyYnv70+IBN1h+SiTkDN6fplwtUzlGFne3piDP/o7wzXmyCEioZyZP9IlmR7PGr54QY+M
S63sRB41Cc65lGL7M6Dua7fSQoWDuvUZLrLUqgd3B1XqRQoaxCv9uwaOeq86KEHJO/kp70n52soe
YzvlfUgAUA3DUyu1Vq+SLlRy7i+ROu2EEM1Z/udnh8vuGWaoIpYwdINyhil9tRR7tDvzWI4oQvi+
+i/8UnMXhncVvkqFOUxSCnCIJdLHw3zH58D207pRQoTiYhPV4IgxMi3LqQatiNzP1D0PWIhwhNAx
hOYLvl1Eqc+UxvdTiO4Nz/PFR3RTnLr5DcbDqfVvsVHk+G5CKJmVxq5Sqy23boLcW6M2u+zU0d4e
Al1H6yytl8cthpGe035/llXscsix9R1VlkLS1Oe5vlFgbJVpi99ei1Pqk+a93ZhJLdo0Sb9xWcvv
2q6lzpFxz2f/EuaLw9i6O0AlXdAHgn9a2NExwff03/L/0XHdrPgH8mX8Wolvg1+//jyYnG3pySdy
09h6GfvhrC0PhRP0qfQLckLx1OufB38U8XW9s/5sIWsPii0kEjolyeksIaK+cjODzgwouHNZdxQE
wtT1kx6OGlHpTNcENSuGeY4BfD780UHnk62wG38+zM8pQVIwaW1R4M0of15Cuvu6+15KgvaZKJYF
/lzZ/MOvan0hpxmgsXIY5Pzylsd3t3ulo6TXC6bExLw0vKrE+Av3gqjsM6RwYWyfD+jZ0SL5f6Mx
/BxHZYv5Bccxc5we59kCtBbnGywoCUv7i40Cs6ZrXgTFvkIB2Ny7bHNW0QPQNwS3WIjnkLfi17Hg
8+eyMeobRZFMz04rCMwoQODy0y6RrJqtJ2RV6+NyAme33Q6rbvSyjyOd4jTwnloOe/NPGDBO2FBw
M+ufhA+vsP5XHkOx1nxmROUF6Fpme/pcumyJVovXcm3atWiimz5Urjyrjusgr2gY4+L+Q2cbamJV
5561TCJpvQL5IDWBIRMVZIzCWXj9gp6P1nJQa+ehZ5ei/0HH0MlEf3Kx+2nNoVltIgBS6+JH/hpd
S8isUl8KWVsLfRMPtm3mYvwHR5lnhk9+FkjvqEtE5QHAR3tpcIitbTvAFzOvvkMvaoJieyLFBaZm
j1KHVL0oNy5o6V3UovPEqe3RUDpXZ8OBYvjQB3oSTA5rYNsbNrRiRMs7D1qdBQfxHi+miRTWql3l
7d7AMz0W2PGh/CRznSMZJ/R8QA0f73Tu+ZRretRCie43y9HCzaswcg2JFvz2f3KyvR0XDPEkhjxI
xpAPqy9agNYclCCmDsbWhoooKMFwehYEQVOyVMWBhbP++jqyW/Acq111HSaLBmPy4DBA1Mq9jOJ/
1M38NQ4JbyLbWmeIryd7jB7wizZ3DwbnlNQmdZpE+f5AMsUswHgO62ddPK0TlgBPEBhM0hgrQRJK
ktFPTcIccyAEIABa/Wi7A3rpzAZNM0CqQbSOwO1Yq5Wl7MJwRTrJxyXH/1pOH8NrMZDFPIJf5iaQ
rFbwO754HAan2qrtcJW3ww2v9AHubB+Sopn/RQFE86FggBOaMEbs7ZfwoLC6KEK4qAbW+OzR39BW
ruQAklX1kfAmibRLVD7GS5SPmrQ4xtrv/1z0taMQskjWcY4GBjN3C/n39mZ+Yql+03aG6L6f3fD6
jQxKiZpwn6rNbvGSvYCICVNci6mKfbCj+kyWQxxjgwgXZCoImINTXJB9cGuzr5mqo4PrGVzCOO2y
mCDV0xmH2c62cfMxdnCAPOhuyMNYIDO8EU2NwLAnEiHalMthEgSfFYUV/McLhJX6lubh28BDol5w
cbqBpdm1aiC3fISbdV4brcEw5Ye5b243vGFfMm01k8mO5UNBXgLUiiEOf32x0BGUeuKjNNDWBqwb
T+EJRPLQ8wBbLt1YXvtGffiM/DMlpav8Byepb1edayGLTSSfKEilZShngUad1+vL8phpLpJHYB41
v/JPhEFbJYHeWQmhdPm4/8B1IckuaI6n1maeNC1RrnY4vfe56+PXIyOtUOiAiln29RE1l4rGfZ4R
ac0AAQHBRc20j8xB0/b6NBLfVkdXt5GKkWE3jWOPVUDug6UrUYLAc0deUUTP0LRi2beIs2EZNpP+
geRc62Co03Do5CxAvg/NeIebQLoQ20qoaQ0ROc3maOTYPqWKAzqnz2WPzeTrigb8W2ZgXE1pLrTC
2ODf63PgvFIo5AXg4HPDirFLKkYbgNvSFevZN2qoLvzODrplrrsX+Na7Qh6mZFdrsod6viwvc/cU
zSbc9aH3DtopuKTxtfNr2vVi6kLJjhxCnn7nJ3F+YUWZMq/4scXBxLpHUI0UJbOVVvmiwXaA2NkN
kaLTgP/u/MaHppeSmlo+18d9FPZ5kTZMidZnyYS4NpKdgxaABTMua63c+P63Y+DdOCbMkbCm0xVt
0MXLYhgwp/uBC294f3rc3d8osNIL9XB0NTJasTnzLOkD1NWATpyKOwBKMXeX6aV8ZdhpHwEQyzMv
VA9ewbbFnZBBIQL33Y3UDDxOtE6J/Zo313SlX9IbdZY4uV8Lwae58b3h6/Ed0+ASNFGg9aOmMnNz
Lz/DD48LGotRY+gDHwkt8vYdjkJQCQQPoc4gi2+AbaCEcAFGnYFH8DDArfdPVSdMFar4Rm5dZjzg
ki+YTKYs/HbH5lrjP/zHIElW6AVLahWHG83UopNLhkSLoFCwN4i3qSwN6mxMEjqDyYb6+pbXoJfw
4bMIcnMAwlX+XmZszHDoWDh0eKZ08SwLEEiICFiYeldxclxfYPzR+PAvmyoh3m0bCjCVNlZSm3Ju
crhDB9T0Kcw1704/pelmeJvnFfempEOiq65gkpgkL8stOMdVsjjWrM/HznRKHCiw+DIZ7x8Y/e0L
czx+G9yj6xT9te1uI5LqyW4Ln3nnzf+64poZ9KaP9RHtitZM5UmtfWQuYsSjMEdzxoJ7njZDkawR
PwKywx46uSlivA2uoCaBNjxyeAP5cabr2KiEj79Z81pvNllvo74dOblByasfwNxRSZwOkk9ITkAE
0Ti5ZChFtd5NoIEZqmQUF+aYJap4kooHKLjFEwY2XEr+QyDpTpYbbgQ0RhqOL/W9kDvZ2p7tqmCM
8l86o9kfKcMSOp/+e+PguJgQYd1Z/9MOJ3Z9S+EGk9oorlsY5VRxsb9+BGAEjDTFfCdOBhbT4NiX
jEI7rpXvbJb0NbLOKgUMsDk31bCy+lS32v9UZ5hTcUphIHA+s/wuNRtuFc3dSm6DSkq/xW119VuU
7X43zFK1qDKGe0LzBk03PEsZBbNfJH8D8rEkDPM/OK5yIo/hmbpI98kejmXcESHj69Xlcna+dtAN
nwo5c3KTJTFrz54KCVMLyiGK5GzzU9oCxd40AjebJxMw1FjNQJ7s5QY7d/vifFaQy8vrVXx++65O
GLjCkfPsEFC2u7n5b8PBMDs1e3rEXPNXNYwyeonauO4zdRSBDLOcYQ1NsX/Bmsf7mAPaq1GTIhvZ
Vy+PYK+wJ3UGcRssRcnVHVBbJtoth0dNfmOAkJmHp1LLkpnV5h2Rq1SESRVLuNnJWoue/NSjFgL0
sFl0P4rtmJIPe6FDhnkOkn5vaa5/F+1mE9jd0Jlx/EikektDNwUAhbIarE2+VVlCrgXEqRr7Gd8q
81M4aoWrOlLpceZqr0i7rOzN2REl4tRzi0ctIJIO7YfWxD/0XiASINuhzDgzqMHZ9bp/FR2Q+0rO
PMpyDHcGcL4M6FWhX1vfeSSMnME5jd4NOttIWcafP7NbDAIrmJ4Xc+W79QVWDdJErvU1c1TAqOZY
AtAbyZ1PQiuoZ2garm1kkjU/AgQy1q8Cj0aFY7/nOJwKz1ftlz/V0zCG0bSKtzrlWWSeJBEC4hcR
oR4w6FZqXihRoWXLGOYcaP0/EZk+tH1Gf/ppfquVAYh9gtwUIUSwrKMgOfyOVpWyngeK3706Lru/
/3F5gVACRP4zn30Bz7mWC9KS5hwElMU5aOK0zSLO2F+9rapwLnHZON+/GxM57re1uf8cCn61rlss
g4wD4RFmnjzUADPmi6i4gs1zRbzZEwKwh3u09hkahQDzGCt8UsNHcGUFKFVd9NYMM/SfACEaDAc1
gqWtRLp0Jzwr9ys/2DXIsc+/cUJ8uiBOWYuWdcleO0bS1T29UPhW+9UjoowdVtfDYOcm10Ba0Xf/
VDWWrr63i3crwAEm/z1TpBT1vhJa5jhw4r6u16tJw63anmGPM2BHkUyvpofoE+Qw/Q0q9XeGIpBk
Ri0K7EsGu5sK9TZ01drW8Kr345wAcNwqd/ghu35ZQzZ5tZfwWtR4uL4Ljsk3tkhlsBn5W8oQH2YF
PFsMPaGXOP2HN9XDknutR+rMD2791r+IeDswwwqJefmwRmp5isad/uVz6JOo9oYu2omUSLNy12KD
8yij2x+sZxa06Gt0j0IxnROunWsqyXQbheCfTL682uviWyp52RhmUowWbUjvDS2isVZDOZsqfvFe
Z1hjfzXtX/qgtzIsIC6RQRn7z0c73hGpqiYdQf/rbV9/dDKJaiCCaIV7NTXYbN2OIrqm0y5tNkaJ
P7vwoEGQ3qBXHJmaQb/whdTkxpiEArnCCB66ynhocyxuEf+nOWE4TlAX6NsxJgh2t7/JO4cLdMFf
CIIm+DAC1Toldc1sxx9x0tFYf0On5YXv70+oh6UicC3v6R/ZlK2mlp6iHBUmcdZ23MsHbwQphQYq
2AeYobyiIxVn7LdpX9vrj6hD+T6a4547fa7PEKMnTc1uGsauQKphzwnJ0FhzTxT1Zk+W9lfe/UWT
tiPS+AX0tsEqY0VaQZ3HZv2er+Iu3k5NfGO+qsHrpec3xYIniO5dfNJo7O7hkjaV5MvuUCXvkbv1
9+QwwKSRenDFV8LKFWqQNNdbHIRCE/uUPR4dcRyWHpu1fTxZYgaCOoXkfXSslMYAmMGEugJIJGUh
C7jL/DbKYk1tld9bUUmHTUPB8+ucWuSY+AlFByz4hsjrURqhY6NqIaFr6hGBWReYxjZYxLN0Hzl8
7S68RuON0k5aPm7E9/S35kqfoc7GN8Indyz1IBM8MSKDLby+dkndGhHNczANg+Cuavgyj8Cz+S+c
ho27LWuOIc8MJD1nhY/rNAPvUQD/cJt99fy6X066jrW9CBAffbm+KReYH0xET0rKJoyPDj/D1+Hz
9jlkriuhbJ3+5WinSAcUfGyK7xHHZeMDabmw3EdAvgylspUPZheMjDLqaZjNW9z1HrlNi5FNn2XO
IJx65SEir/z4RWd72BdvfbGrLdEqze12tba3M0JXcCHwcIpuaWAAokDz2C4FfknyeSkKRR0AdL5b
qxuyg5olkSf/UCcjpUP3io82byXiuqG4XBUMo3sOKzMxGLnaviCfOhUig6p7gY+UBaP7w6h5YtOH
5gWzcpAwZ0k+HvAmcHVC1ITJFvc8fOgeCsilJ4X+swsNOhaGYJnPHOpm4+YsvpspHEFWJwceseFa
72+5znEf0nFdkrRNLV39834eYfJGEx3SnfYrlODTjCFpwjqP2cH4dDpOFU1cdbmxzT8sZtCdeCXE
c/H5JYeXhz2Ik0KjS3a+LK1+VW2yMaNbnIb1lF/VdsMJA4CSNUmRYDd8oHd87sxRdXLRo5RFqEGr
y6oyN5riPHxheMTHBezRRmGByLgVbwXcFvLpbcKyck4GEVkuwvr4ZRpjWEqJOPgbm6mtO4RS1bul
zykGpTR8VQnBSsL0LIIyxTG+T2ssnsqxs1vMqBvN9T+2FEvWTCIuUCln2uS0gSTV5QOZhzv9b+J1
vg9Y+wGdAqxwpeWPNIahvafciNzvNJXeu1TlNfx4JXtW9E6cpC8RWYgyCnh6TaVef9uk+QkzbB1q
63GcPpK39Y3eIwNlbTNlHNOq8zYFWndHqQV6OXtGt9E2Ks+INS6EBMrvXk8qHK44s5wspGHf0Jhz
qAk2TLLfamm68jdPvQTTlWrQafTbp6YJB4af5Q1thkdul6JMXxDvqSkgf//StttCHpbE/TXyF4sF
yBytSDfh3ojNxQn0UgdBdzyyZQehOYtOdP9wbd035RXYrrWxAdOE7Pmkp+FCQ1d6+ETfYlo3cA5X
0MNBaJj10tgfRxDYFGiTDbeWyaFdNcblv+9uAO/pi1YG5+gDNUZroK01BNsBp90rf/wd/vddkEEa
OaNFnMaKGaZx0k9qU/fnhAsm50Hatn5gi+Ofbb1IiXCmg8Zy3BNcmmOa8EKi93FoSo4+0Km48QOM
Tjapo3JeCEf9/IJmShVRBfyvfZi1PgJDPsTs4BFRjlN5cXvZdw61s3n3woDk2ZRZTnDqsw6idNdA
mXEy/8Ehl6OYQfgr6mJeVjV9mLGiA0nEc/yx0t0+tamDdAPLyjvIuBKcObLcPT759fWf1RADcYMp
MoLCtDJYMEqInP7yrjjO15B2WuSMLtzSUTl1C523RK59+Yb2Q0+lfThk2RzlQJ+bJNQ0hHvTBXas
MHqOkbAL+fTzvzJ2RimUN0cQIhFrJYzpUpxWf8CjUTKnVqQuVRdLRxvaGEIgarP6+Z0NnwlMopHx
CzF0RhCmBwPdq75oCtsFHEcG5PECMD30vHDTfchYMcTkVbpEdJGtQdSmN0a7AUbmFRwnt7BF3wcm
9rmmoVOmFimmIGu+Z120MrdhtYTw7GGLQTde4r/ER0jPDdQxQekPeOyWcRfR+8Ss4TSn8501ym2K
/qUElodDzIhEfVfC1wpj/4iHD1kF0A9eWFIWKkwjKIJ+YQKz9n2XuIpwDqtq4x+S8cyALt3WMxN/
xFlClFYfAsMTemtJYTGddlG8t0dzU+Jvd1LG8GeUQz8lmmvVFBwbFuHGXZXJng41sR2rHa5zM8gn
kduT2lNUCaIMvoeAKrVGj1ukARp/YBJW68xNPZYwdIk/C6bD0wgfCay31b41fZeTVtDiO7Nickw1
BY28snJzilXhpEHw//jomeGjXFaIomit6co3jkNtsdLxypRS39k2rmAEP++4kE2E6n1onsY/L7+t
7WXM1kV9JiQLwemiI9ojTbCjt6VTMkZwM6L64hFYfSfRoh0MmOfvt6KSUZ6k+Z1ETBOrWhkkr1Ap
T8Hv07Y0qR7V7JOarPGpvavcyCXZU0UJNTneLUtDleL/NejvgpXww5vylkIu/xkih3Y+rMGEKqgG
Nja1OKUa9ngEudnlb8W6tauhQ5bw7pnAO0PLzp3Ka1mBvLboLSrmhrZvs2kcrWY+I69Sa1FRx+kF
silqSUfsniFVCCtBpy0WOhU23cUIr+V79hPaHgtVydmCL4AmJn5GMlsY9cgnoMNcKgiUDxtVahfc
CwBabyPSa/H2BV3+EyQK+l7d0ZMSia7eTqvXKqF5EBJlQLozyPDgGrFyDAh3xRx9jIfERaXZ8RGD
DrywGHJeiBduwHaYR5o3+d/y1jXQvW79vnzLg4T6Bbbkro7ATqiiLeFq4EKg2+tuU7cb9APwwZxJ
Du0qYNQqQUgtbw5JbsziRm06GmKEUkGKR3PQtxiQ+gHljbisSMOh6wrP0JFpQu0/jlIyeSKRSeG7
A0/Np35v8GvsBE8zW8+rvgHJf/LTHG3qXfMXI3JpVj2U+QjHM1QbfXmaEz0uahBocuP5Ce/GOag3
tXL1xJdXk4wFYbUiy9746/aZzUYdLCiMlVPC7KLOu4elzdYQetKVibaN7+dqWhCQrM1wiIetqgaW
ZnS5Ps9lj2kLy1klkO02tJBVz1+TQym8+lGnoOCoxFcHdc1/hSxk7Qe5rRJ2Vk+MxLQfGb7D6Zxg
gwV4UZchfI6t8TedWAKBXZVgB39qqasCXfQD8EXB0LfGcUBzJ7hoesWlaAAUcBjYYOE23QsAf4qL
BuNW+Ik2FFSK3wAS83kSw2ElFdZthMqoE7ZFvhF6pEf118uU0lZkLdGkS+m1e1WoCuywUPOT4jrB
O7bV9lmMmstaR4wCfkLFraNJSzfeOgH8r4mJNztznVy7deeRH8y1RbwBYMU6kdaeZX8x3hK4nKVm
tHeM6Xkd9Ka0zNskJRpYnDUqqw2878GXtDLB8zaJx5tINXEToUSm1ZvadwrGb/p9l6/xY/JmvPs5
rSbRRbr3vuvJ+9ZxNW0WH+Wj6rOq2vmSbkzTIE2DqwEkn2Gm4w9tKL13+F3eYAsKVEBrsQ/KzP7y
28PRTbAouiOiFPSOoSeOxYxVYkhzMjgoau0YQVXhUwNxHKAOcF9UR7wRQD3dCsEeeCqBn78Jyksf
pGp4FbtlAI1z5DFL0s/7EmwN6n8+JvGWQVb3/dNmic168z2pEDfv1L8ekoC8BprR0CuCxOO5AwBH
cFo3noi2iy8BSsot2HJw/zhxTxe/dbOVgQ4JqslnSNwQbMekZXtx5XqoA9q1tobRH0i1q5F6b/Uu
9U+NnMAgoQgh3UKJa0auNVjvDAq9WOaQS1C07Q5wVyW8dzAb0OlQHLX3UZ6MSckaNlhbzj+1N0IJ
kxGo+Lr2vYI8WEVAE8vhthONv1ogbPMtCQi3j8PgZXx4GHm0jA2P+rz/U4h2/3JpNm4m3i9HqV+s
jMyLNwwfewSTGdnKkNpSvl0I807LSay2ui4BhWFBzGfn833ID1eOAFTp7aqMR4tW8ABtPI4X+wiX
0mD2bxJlyKZxKSMSVcsIvl6bk+dymq1DqA/KooK09FHx1unKmch3K2xJSWC5OcbwSLVNlk68Mvbv
Acrp+P6MQICbRdPQKnSYG0bF/9q6A8WKn/1ZKDjQHUf7TuyALWOoKAJQro/RD58VT1NxG/b18m+j
OcpphcFXepRidRXkIJ6pL6RbBw+55Q6CaudAdmoYlSjG1ygzHDDrTtEWjrzPemMYrLpKuV7zvNZx
2e6bVVFxo3zcEKP0O3AXC+i2X0sDy2KF7OPMOzXwjcdrbW20sjajmuxDivI311Dz9YBabQUV3wUd
7j/WTWGdag9NiEd0ipoq9/ooozMqDMib4WlRSfSUSqHJghV/adluynzTiklffQpGD0Be0SvI05pu
KmmSkCyXQXimgPnQ+ywUuZ9l7kJxRUnZNQW1MN7/3agtCPRJfRZqFjVDFOW8Nn5DPRT018n04qaX
D3LS5w4DIMeZ57tuTLpzdTQaf/NXegXYUXnCtHKABlz756Tm/sxWJ8s1uISrEQ4V2FNE5GfAmZ1A
vqSu7DwrPPg6ob/+kRXWZ9xbiReSH1b5kH40S1cVCujL/zlolDCUwE0+VF2/SMTUh6R6+9CDsrYN
ekK5fmaVY8X8093DVJ5M0q5CQREe4TrwmuO8H83r2M8c1NMK8QGu53da5yvb33CYHDgjT5klJEvg
BVQ66Apbic9JjXRYdiMKFLlizYht0HjrrGYwgv3ppwnsOTv9BxRrviNWg7nRwse5OOLF37PqE5kN
/XzHdbRw9Q4GhEo59Gbq5Kr/dZacCoFHN0dSqbDRVT4Y87baxNR72ZcUlg/hOq85WX5WvGyNUr22
k1Z/bpC8qhVIlXWUHcHMoAV0Cengr0JLcc4Y8GCIxJYSBWNSdw5dLwLhHf8wKUSz0pGa+3aTEsAN
Txgl9tK5WQ8KH+yAdez8myLfENWzXIPHh8htsXaKb8jpSmXIbheh7UuUgGlb+jfvxIHHwLFUKaIl
ai+/QTzSgCYtMOU86QKAoE0Wb/v/3bXjchgPp2MWbcMz48ubB7TgKXrE7691TMCzJjyOklcJrBXz
wZdugZFRrCddtJap0veuis8GjmYST+5tArj35S7D2RdQCEJIGaWcsv4OESVSdmjrKT4waDD2mAwU
cn6baQXxYGbNVIQv2AXX9mOnBuEZaqHHmSjKDy+V3rooqBKbe+fZk01CAuQ5LpM3lY7We0EMPlgi
w4RafHWhGM0wWJkWnbWWehYTZOFvZz4h5XsHJ1fA/s3bgQ41IPhW8/NA6GCmQmZaEwUnWQFX5D1w
rt1mwtOgTckqp+zcG1UEwokMzEEzIM/kt2mY2XkzSN5OI0E3NC1dDdw2/3Zst4MqqChH5e12WtRq
aCNSzCktWbvWCQaK0080cdyfnduHLmHBS7YK71Trp5tIaVhFyjx1IAZA6IP/1NKmgKHL9wJf4/R9
tZHNU3OXXxJKeOCNSfvTAfsY0L19pCMgs8LGLERYQwLl3I2mTcx/0bUP9tN5yVXWUj+9eK096uoo
D7VxR2zIMCAIOz+rFOoma4FglvrcaTNRyWodNYsZtbfY/lYlE/SxcnfvTiTeBOB/X+1gUapdRcUS
5NDwDUoSVzAVfx6oqgEgfwar1bcm9bV9+u8kKeAUknuEE/KSRp+dQEprRmd2AukYfTBno45iBreX
LPRCeWEva6PRc5k/4xmZC8OFxaiYSgrO5QXSgBECdj2PmCfHrm3S46+fLdsnI57Dh6jg2MaZeKKQ
u6FRNBSwb/ojRH9MXRh7SozpCyi2irnzX2HjxnN71kjaug8CvAhOyBsksqZ7EN4FAOjcyDheNqib
Bn5wSXco3P8RKqO79FeiSbOBfLOZBplWW5i6AGbazSkEuqh/PhEhCjiCvvTOjCLl1mXCjcideviF
tyXfH0Ngzh81uZC/zPSfRK5xp0rmWWYJyD0eovGszRVbIB78Gq8dS+TRhCNs26qGDeZZCWMTT+j+
AIuyzaMWtLl/8t7APafruzRUBrP9CdbXXKKn+vC05UszRYViIs/S7COYRB8sROCMTY1XXNRpWvd4
W93tgmEc2Mwk+AVm0rApydRAeFHIds/BthmfYOKNlWKnat9pBxD4JgvliM3r1ktlnCeyeNDbtncS
AJ8sJS2AnWe4NsWZvBYrb0e694wkBr+Rk/mk0xlradMgOCmxaTDYFDGcNS7/UCWIt7ucTHc9lMRY
LrMh9++SbX1ElVU/i2t6bi9rF4VAfcK1pjleu2aWW5r7GSaZIiExtQVo0FNEpd3bLUaK3pelgB8A
Ed1TBjVShjS1FmrbzJNgTScN8gFrTinkm0Lmn2C0r+0Ja1ftZuy7h1NnfieV2VD6TLpxvchTqVMi
9Tdp6Q9ng3IjAqtuobAYM4DXF6FGpDu4sd03hQSciNmRxYBQQZCxrLteGFnEVD0VgFv8Lkwqbtwv
wMvJoWAE54qnw/hJ2n9laoQbeSTVglhwCHmzLxPz+4pR6UZskFM6J2Mi1skYm1ca7G8BxV7YCccC
AmSSyGMhrswpY8eqCKR8j9Z7zjuQazSSeZ7+ac2E2I88BkdylTv5UIclHAHqDQOdnX11IOHnEiAy
udoYUBHabSRZzgwrDaXAlGgHrqu2b+jdL1yuCM0t+awHFK5GaViODK+sRdj+V91SsiGx0wKu3of7
6U34YnqR+c/6bGhJHZtame0J5iCZ3U9FBVo82vJbXNgBKS9tTxy29ty9xFJ9kyYjsgwy3MXt4KWr
4DSFIk3uOEnIri0LbN0OaHzxFCz5QRmDuXA7plIo6yxvg5VaZCx0bBU56Ez8H2bzesKYyVdX5HeV
s9/iY5vYe0z2xMKn4vGyts2swBsY5h4nv5FuO/JsvHo+/ITB58BYoVeCv6yxk9EkKkp3kzAdCvul
nURFT0l7wdThAUUTZcCOUqR/dmMH75llGZ56Hzq3tdONEh42UzKOvJ2ScbwUDbETTlAvBOwxMb+6
Bk1/lZ5oOvSIvpx8kPZC4aovROQ2eHWA/sjr66ekdEdg/RPItta+P8Lpl8G55qp4sOXNUl66V92t
NHQf5xaBDq9tZLT/tyZdJE8wU/GIY93e6NEdcu7nyEfNoIB56G/jRdDfSkocNuyLK8xvKIph5ajn
ttYBfj+f8cW9L9f/RgtB5yZJWASTxsjSXyC6d42JHT06/dh8J/KD7cmzWyW/waB5ied0+RW3IYzZ
LPe/ysVTvO+g/NznX/qjJ6fz1Sy8iSBZ1fGh3CxQ+U91Y+UXVzF4qFnxIecn4BzhR4SZi99oSfBZ
bm/vr4aMRvcTu4jbmrRgp8Ft5PAQRlbjfgwto65aeDx+16oPw/hmBhZfXzLVNZjtKXZnE3jyRx+/
WBWo+P5Y47pUCjtmwu++w9InpC0TwFQVXfETgcOO67UuxDRWiVv69pD2oJiCBx9SAxnPebnuptLa
EP8m0ClDv1sZUztCVtmht6O3zxuxnvr4JrbxYUTd9IM+KY1g+MSo7G07Y0yT4A4qOivZi5eQGsRs
t4QLVXrLe+66SZS2K0f7kEYH1om6zT/j4mdkFASVgmhOB7ttre5d+hH9ENfTr7IK0n7q4OrWpRf1
zG4nYtOTnaTsTpfQFEk3QJm/OFDciroTK162Z5iwMc/9Q3fPW9nWl9KNw1vAXDr8UYJRf4qMlv0h
6bWRb/dNswaHfNSQ/EZXGDx2tA3Ate2IEyOm8s68MyaJ1KfySatVkPW8yAeXqyuIGEfHwAZ9/VQ8
z5VgU+EPUO7qwLUwikIjBL/bDa0WzswB4FS1QhDcQTXrUPS3XnOr1KuoRvnCNK8hh2tXJq/d5OZ9
7RFUdjSltKgI3kGWMQBwhkbWpXQq+t8bB0WyTAv2M8kHyJRSFxyQGgMzePlhJgM0LRM2PgNX3FlB
PW6d+J8aksAH3dG2yBCuqZb9Nrj5YO7lWz3IqgENRGSH26dQ69B0DhXePynrT16ytLIQDeuJP2PV
PO5eafVvZOwkhO3enDFByNjkJn86IyzhdlSk1SPXjBqp3q2gVJZ9Nw4Pyv6OWUuAjKX5iQaX78qG
+4jICluB5NN3pPFVf7OSKv5SkrN0tRidFj+wDpYA6xaDdHkpsEs0UbI8+aXuz6XzuYrN5CxSZJqm
Ps/dV1E7lV7NywOaxF5rw5HQ9dpNuU607V3joMZFV60m78plzItufzZKSZRD/eow0DYRQOpblnD5
zw1KYuCn0wU11ejcSm6ac+iwwJLZJ9IFRzgSDocvL0ST0B34QkFIgQy9jPQwT1xvbXdg0Q3/dzoZ
t9bN/U4+C505id0D8sKvXdy2gyTCPyfjez1fZY9JA10CdA4dBjRc3Aj0cgoEVB6RdXjPnTTo6HT/
SyzwYtdBQiz1Sh0rFQyPWwi/2NSJiNB/9HtP3umKR9Mytvg8TwaYNiKi5pmBbaPSgPsFtkaON4u2
yNyV4IIZKJtfuioVISp/Lj/fFUF0fTXhuWW6LJ8FUEXxCT7DiEN65YViLAJ6exD26x3xRnjEteiJ
rQNOeV4RbdQ4vkc0UM6ji5H89k52oM+6nFtPebYE0+2r8UqeJJ5hw0qbVubOBJcxC5DmmWHXyaS0
uMVELuPg5JGFV1YlyePG7hByvf4LTMqBQmldlgtV4p4u6AMGxN4xMzx11MMXAWSFzyvNdAVqQwEn
VL1evjq5B5C84apSGxbZ1cwoytXfTsUvxEpAC7lJUv1dJleFIrMnLv5Vuyx59zBjGuqbHo3u34WL
HTuHjGNG8MuVenk0ZV201hixFdX1rI1ANJq/f1227gDwRvQquMh4JwxKx67suF32TXNb3BVqfks2
g5Wuq/8cflbwa2EWqRVP9DakQw58w9CB3Ol7ScoXWyZsYbkcNWkFsf6hkKDDsPz8dgh9TQogSXbF
akDZzlOp/F/cusdolTDsFLjyqLDPaQimb+3QBwEy/Qylko6NnPr5F11G8fPDp8qLp1ABM6DVXO74
LJielIHUyzsrpxDv6TI5kxt7kxADONw63SUDrGGLposj1WWE8iCiz8LU8B9I/MgtARaETwB+rBQ7
fG8mFx6tMBvaw9GBW+r1X2NUPYw0GUQRKK8qyh+Wk9z8zIPsxhufmryYM5ASXV50W8TR3tokJltV
u+M1JXoyc0aMkXgCoj6N68Cciw3cr6zqlPbynzYFHdz+8MEZkzOXv2J3op3jomAuWcqqX0jxDL5h
cv4zZ9idit/AU9V70zgIlYq99Klk+adXJWtb5rjfS5EB74T6m1WWBsapQJfRg6f9SAsIO8punciz
/afY5zJq4aw6qw4y++Xuoba5QPYKOF1ly0TjTd5mwZvVt+wyjpScqoWhA/9F4oDY2+v71+PEx0uo
3cCqjGa2+vB3KkueV/pY7JZXERaPTP2r/v0qTaphdNeh9tD0zvS68G4VPvyKqm9qPuOmMhyMApte
OhASb17v3G0od2x+eGYNIbDNaZ9Quj4gmueSjtsv0g0ieKdMYHs/ZS+p8bbWkPLJmHV+daCCfKUx
1Xhk8p6kW/GJWLVLsf5eiSmfa1LVnIJhZFuz0rj/Qlv9cpbNIbexnFfwe2yCGB95V5ksFUze2uNA
IBlSxAC46zEjLZVcuxJg/5skEEbqMpHoaZU2UFOMA23zpKpNlANjr5ut9CE+jcub358exu1IhRHR
9GYYizPfSdEkAC1m2UvxBZH4L+Z/uBCEySTPhkFHeaQOEAvIj6Zj4Pt1X1mFh5CpbmI8wcyd5nmB
IsEaAXL45Pe5VWIZV/Izh5cyhZ271fCuD6uCG0rbrQXOPNewsAF6Cjbq59jf8TVt1D8bnWXQwafh
mNahdFl9An5QW/l3uXoYmiSbJHpILzvIm6hgT5u67CFKcGmstjMjqtEi7xvZXBB+/+o0a1cA5BVk
+9moCb5vT2fy/b3SBqg4QhyWfzp//AFt0+3khX60p5ZYCn9UlQrR5EznBvKZN6dI3gkmx1/NeshU
jiqud5P6P4fILCFiecNA5XFtHgBO+hJ09w1JowQV1JdwG+HNKNYu1Lth+gPgAxGluQzvzj8nqraG
4AXuAheBbrFvsSTpuAFXg/abMsYMA0c20wI9wFG9EL1AtM5g7ZFy3JY7r7+81H0F6ayYxqgVt9kB
UCDSOF1lFMRlnMp7v40+DdvQyH22g158Gm6MABbBK/vqxoZrBWZz7RxCM7sHA9qxM1TVTuUhixuG
FZdwA7Ze+8wDWe/syCK/lcmJbES0G/ZD+77F+QCKoF4kFLWPdyc3EKZebtD942XDAo7hpvgLQbJi
pePPl19dIOrUTb2a+z/7UPt2FpJqFpbidpFabvhuL9JU1wDTbanrCy90RyF7Bw1Fyne/emudJtkC
y2bHxWeKF0NloVWAOCAQxJKk682dVGRg4jt9p9pDyHtNQwfHI7Lww5kllhLYjhn7fumzM+z98KkI
Le2trem/2fFUpfYP5T5gKAyL+STUlV3FihQMGUHxuunhOXW01t7sW25wtSCkCkS+/HYSX3SX+9CE
GJ1gi5Xj432f1txZD68VgKNX+Raw+wWQ6/FMiZ3kaGZSGM4U1vmV4CEVWowrXPfDgWFbqXEwjxmj
Qyn60oESAirTAcAvMtmBV3RYOyfUsWx33FhLWG8i/yK7nuDVRmZvFM2b4KorxlSV5Po4U2Z1eo9M
w3GfzAI5TYIp6JhVXLaE4HcVTDNWTCBLHod4cABmT5DEKePiyO/na7dIq71/qEbwMy2Cz4FX9GL9
cJCEf6qO8rH1zvFt/kzBtpllzMi5d/KbheIxJru+zwpKAmECqe0vf0ppan57+EgQQEsFNtTuU1cu
IE0+WEYXLKg5Bc/eQ34b8u63+I6s3lvgdaJuL8jNXwgVsszpkqIZn52qhlv1teZ0SzynQSbfWpek
rDph3N5ZA7jk3WMvUU+5V0qjDpdet35BQ/NycEjgA1ZxC04k4EP+HVSrPIOYpTbWtTPA8rmnO+An
pn96RhdTl0R9S6G/HHkjao7Pfh7HAPiOYo/CaP8mk3RovC1+xOY4w5ZhP7shMaM8UoBiOHIZztJC
g2D0Wz9kOxEoFZBgI2fyBKsP4wLDd7eJFaMIttTgq3ag55FtaSvZuIj9YFYYNGZl+UPvLhzUaw9a
ziKNGo65BgYGlnOtaLp9bQKnVZjcxn/t8Ql/mUNn2O2FG9K0XtS+6XELN7hUC93os2T4wKpI/YIb
HjRpqXENHzvDuPTVi4XmdI+DFUfhkpNeK5WjaGadmcOWEv3EPJRwlbb8XsT45tDJSisFDyvqTABg
Yd9cJdUnZonPqYjcsYzLUJOlXQvq6ffXROYboJK4UfpnLF0L+vU1gcrRSvwqC/EhjJNiuamZT7UB
iwJtVkzpnG7/urAZo53Xv/b94HoZKeqrOdQS81e/g4G837f8tg4PLXkSu1T5zQtHnhpTteJ3x6Rc
To7Own4lXmLVHuGw6aCUARRHK0VdyZGmdu1NKLvA4ue1seVp27jnCvp7vYe2821r57f2e0Yaj08/
R/I+fLwApHox+TVq38wbSVUpctIE7H0khRz6FuULmv1+OOzgRP+9uTQbzJ9jxHBP3lJWvcGffkWP
9WmihBQurnbQTk7rAMOhUYd2d3D53Pr89Eqqw+OmIuifhe45zFTekAc0DR+NPagk29v1dARK5oCm
Uy07nHeq512vh2ocwXBzYD3y0d36+8KZ5xJg7/z5MAg9vc1LKQb8oRv0wMvH/34MLsRkyHU2rHWs
sSI74FkGhybWg4fvcEH1C4tpejCAaLuyRR+ZhQXo+4GJTE78KUMxD2kGPpNK9Z9cTIdIi09qMmSp
gTEdJkdR8voTnPCdZO4LjVV4+DNZb/Ehv28NXZtIjYOsqsb0q1OoaRmkYfbRpiWRy3kPnGrKOGWS
v3o3T+SAlojqf2yas2066IpoQ9Xtek4UoerlGAuB5e4ysPqGfhI0Aa/POaLiQJeISIU/VfaUgkiQ
IaF9Cs8Wo7LF46JFxZL5ISPwl36aTCoJPPh8w0ub9MkUIzOiFg53nQETeW83nwOZxYVa8KUZBlWX
zd91wALd64xQ7dhjE4zd3wOZq9236P+vDK5x3ugtGIHLjUyqMVvR8uNzYoX6+LnsYQwlY0RMaMGA
K2nGs0fQ5Hm+2b2hz4g/FfhfJ5re2eD7ZN9i6wn73p6mtAz+ptER+ggnICHvmnK+RXBcJEaqRjwd
mA+NFLQ5tSzLbw1AXrEH8JVWYBkMLNaiB2TldLkgF5Tef74ro4LcIpv0FDX5OtnUA/sRFgKcSvAV
oKNRKgx2h5oZsf+hIwC18aebUADKg4M7G90O0M46tm46kbS/CluI3Q7L+BgWxeErCQA+xr3IEiL3
jiyzj/2x4pq919d4kIdjekk4YzbivNkAYVYq1yJEXib5lJtpxKproZ5oYIIIjx0JFsPxBUnt3x64
NFhdEdQHmX2sJE1LsGx8TN+7GiFXAoN1m5Pa+sSiKmiIB6axXnjx3wgkn0k8hvUvJWelBVSLeQPH
AX1O9NLqAliabsVTpk/+DTfqXkEvlkjzyoQElGzFC+OmcAR6ajxtT4oWTdR40WDUg6oO7ciXQxOJ
cHPig6KHmJbT77t9OHiD+LtUJ8r4iXnvR4EL8RQCf8T311WbxfblDXVu8PrmB7pOzZoFj5WybGOl
ppku/DhHT7YFKOS7W4FfvBCOOzG5G2jHeg/hO5bWnxKpsxoVhW+5a1rOF+wJHaFPinDryHXQOYvL
jXfB1J6ZtBilawL/fmBOEMjKTZV4pFyRCLcnA1W099CigcHoYmFbCe3y5XMaA4P5djhAL6/3Lu1E
nAG630vtRP8wNTAmBVbHEFq1hoj9LpXwxnWlALVPi3vdNtFRYrcGcSolK/f96pwfB7zbi5Kq+Qdw
IQbfSPtIhZYgKet1CseqAZ1UxkWuoH4pXeXDB2SI0YxupOGWhzW/IS0O1G0E/rBgns2Q/Y/QeSq5
7cpecPjkIdsoNEHII1VN6+h/TEguEbyCbZCoYtaqV9HtEFFsdexI1OhNUfhSSwTmaqJegAn3m3ZC
L7ydu9rL3e2/eZmm3D3/9eFG5RAD+UuwTNncFLqey24hgEOHwTezLfZ7wi9Tv8cbphRSXPTH4XHz
j4Wy84i08+H1MNRBo9zI6XBOx8BzyzsGfQhqOl7O/03YVnj+QPWnEu+nn9i155I3zj2STMbtX6On
dmQVnXG5169983mmjeR7Dbe1MhBuHgDHQcuIppRrejZOFecE59vXJRiturJSGQGe/DzolIbAM9yB
kVZBtXl7B2hUQuSFSlb8+XZ0F/dPB1v0m+ydRb8aZDD8PyHjkRQca0c5iAwRNC90AJVOeW3J5GTT
3ZZ7V4VOvxUX7CuWPZ/TvgkME9mo2QREAdiZnYx4T3XszEtOeBQqr8OV/k78+/rzL+RKeG7LwfeB
7jYyK8mgusAyblVUgRVZ2ZDetnuXczNkyxD87E2Vmm5uutfDC1rHz6B6aRUPg+yJrDCtxVyMuGgq
BeWACt31tHcmrZ5hlzoEH7QdkyF3L3TQYZqd62xJDp40QhdAHViucDusmokvRTbNYgJLE9CtSh8o
CU9ceOuyBJETMOYuGbmtjYyA5Ma2GWxJhPwlJypD7h1+HxV0HFB+p5/6YoiFIHTl/s3QKDzAIE3+
X7yI+6J32HBSLXItQ6Htv430KCjfWRNdfQRLyW84XJDfBfAzreuNzLt7aMXG9KB0F3yb4Ksv1Py0
fF8LXrh71UxLmJqqqrxdWilPeY9vLpv6TKjNWeMKNbZVPDQ3O980hv144oLLLbMrZmy939lnsxmX
TkkJgoWiEl1KCzZTpqhUzb7hg8abzlt8I/HCFRWTbFmxefF5CHjTC4xCIpz9YgJ4qEdMpiOZ/y/e
W+yJNN+2VzKa5TnM1b3xStzHJ7FafXEtoKQ5xU/EOG7LJPGbXNWulgDeTAYRg36nyY8o8rHPRogJ
P1553QaCy6UMz02pKRpIhi3B/rF6dS2TEiH8DY/CjIC+aBAIhCtHoTSiFDWQnR/R4kwb3YNMKrXh
JeFruUeTArW7g7p80W4Ymy5xbvpRfbnPZXbDK+YGJu5CN5BEEudDFE/0OByrI3jKIri3/JtduQSc
MWGpl+ZQHPN9UZZeSf27A1FuzzGKwFVp3bsfugdDYo/IVutxtcppoo+CAsih3YkvQZsx1ZHBs6nh
FxgzQ625lOxZqLobgUZJiIDfcOuO/HoJjXqkxz8nyu2XQBJkjPnCyHE623KGH4fENlA++z1sv/xd
GklGNSepLUiWy8AHNxjcHBxSWkQ8TEoe19hNzxlfIPCHDFvgUtWoq7KpxpPVZ9zKwR/gWfncKlnF
GW9jUnvjhHdGo5pmZJe5WZEJF0775U5EYIm+aYaqlpBzd3ytC+nbBapsCt+MTOpWwJOEK8eCBO67
/V/19eQJWE8W2vfQdZ5XyPQD5vU+eGWEUW5MHyuReALuflSW8sCAWXtndjJksUh0oaH1QKWHFrNu
PlJG52OT8X6eFNem8zVrZaloD9/ENCe+yyQkkZ6ip+Cu1nWNApenDOjsz+4yzk5H+9SEb1TEC8u0
WBSx+AyyHO+hGbBVP80JC1CKpYsKNx1EfjV1auWsD3jqFYfMVzpQtfr4CSvP1oudOjb0gF0/9jSg
xNpbYYAvTOiJMALMM2Qk3uruN5qIssaCj/uigiuGvwZ/wexusYZAO9259GoilrbmqjUHeMmt8+69
nkAQ77rG5+gwi2TkoIqe5zc3paDLmTO7ynb3ogcDHFEe/74xYwIvHvpDLDhLRfvLMDMeWrCzLAM2
AqhAcMnLHVOrqC8x9afBI7G/ymAMPIrN81uBzSgPzQ5C4vTnOaUTdLtJdI5krxajxOWVavAylEmq
Dk+QQTE/oO8VtBt0hfb3dqSEU99H1njL7EUQOehnyzKKxS0HbkDW6Ll5v/ieB2c4EWswWbljG/iA
yhLHx251nQYHbsRi6nUOpvPq4DenBBQxmH9POEe/Nyb7l/gZ9M/c+jeY+rD5Q9V9CO2jKQl/Xm5S
rsfIMEY3khMBGamR/apulBWNdhEj8LjELYSeUsEpahqyNqhvFrHisiG7fYZr71s/J970Iiak+i+3
5mBV51yIj9TfA8otl+5A+WaQHRRQgbydRMmMc2s4JLjv7/Um7bj6EcFTLZf0o6HfI0q9D4Plw6JO
hLc4nxalWOfQX6BKfEqufpImBKPJriC7YS0R2Z+k0xTWEYrvywGe2Xugt7yJjc53lvxqBRuLh/a7
TTt1FV2TGa5zE1bCj8+qT62qbninE4gYAw77GGhKo47omUWSto2oLq39/mldOI2dVToqvyNCGi/3
kUHIlGJeG6FcWBQHdSIpDjWOaX+dHONoXueo5zWydjFHBQSLwdEX3kg3s5RFy6Vte+vRxbennkt4
wGR5XuiVg2tuM3res+C+ut9AO1h7qeKZsxk3FdcR9H3XAn7TQMpYVUoBhleihddY/aUEY6M1U+vK
kQRjhK7Cbl36t2OChMTCvLOUR+WeYyl1mzoAF52EJ1Zv/Y5KKI1ZxmrQADHi2qMU4Mx/0SewjQ37
vy23RsZaeUg7Ryqx32rwjEEDRswSXkjtCBhNnNo7/tHkETMwXv7H1HwgdQZm61zz1sR3KLMi0Xv+
fVdytl2EATiNFgT7V/IKkqUFkU/g7NXfPEuZPSCHBg2uToGtYE2z5ERhUbaRBzf6/oB4Edt9RC/P
8ryQs+mpvphPE/3tgJWVtXQStQSBfU1E5PsDpcEMH454qua9f6tAxtP+wCF/BCSCb2Rskk06obXd
CpeXnETaTm3UEYZS4v8LAmw2PbOGFep/5N8ZOSYNqObc+A2xtJsiYawMD7MlBeKitUJ26HTerWg1
O+WNtdlWNh9YdH7DlRQgaft7MwX4NAqvbkddVFVVcShdAsWR/ibh16tNvlqtO7HIwdCdXpGI/4TS
D5YPSn2NIYVDD5MH8MoyThXhg4pLiunZqLqkqzgsIma5eMWRwpL18uzFsiUYsTcDw6ri0PYsnjWZ
vRJm69YCQSw1Lo1mJI/nKsK+esz3bZKGgdZai9jUydJw+xGW1FQ8+cL5c1WFQ+k2W95/ivoEFz8/
pG5jzfxzayB/soxBhNlE3KOjHvv5WYr+kXgkeWjfteTft+2YxXZy3gTNXFc71mu5bH3Coootagy/
3Q6WSeVe+jVxsA7raaesMn9XVchxonna2wy8AnqXeFtUOMGWhyL8ok6DfPcz/VHfEj9h7o8mORMF
X+ica22VukO5LhrE71luM5tfs/7ZhRTA2b/OuZ3F9f3DC7qCQvCSsw9oXS/i5rP2t7v5YZCZs+sk
ER2rXGtdDTUu+7UBwrjrXIClnL3yvUL4u5D0SEhctSHoIdCauuSLkgEr4wh/2g5Ak8GGcOXLtLTa
INMHzK42qlIo8aXdDRAfou8xEvtoWfybf0tx4qZrcBj/HuNEWynVAWgH1aEnTMrnC/mcTyxxzcnK
1z0/Bjtd61bWgMhGnzmAHWxDtvzTEwPOd44eFchDSUMjS9kZNyEXgyMmBATXbPOrE3ot7UOdFsWx
Un0nEz3Rr6lX2sVIKy2tKDABLkS9WBmejTQvoK0e2CmYiHYpNo2rVts1YAMeN+Od0kpDallBpZYe
EjhJAfBzOT4bGNe9LbGzjpqUsmTwkirq4xPlV+HaNEgpNPHenfbIlX8DWJe/8mv1cdJR2ugvKSXy
Lo4JhGDNJM3oOCukuZBzb0Q83kZrun8kLqml6wpm/l3oHxZXRmerOP/4newuvfSG10tjuZZrmsGF
OxasyED2filenQ9tYEcT7bUbS1IgTgvZnOQZmo+ytwhrrgLE3+o10WdFPZfPu/EPUL82RGqi08Tg
FDBsLeXMg5fhwi/qBAwt/TL6czaE/CtTG5vVvz8FGQovztF5Rsd8mmDLnFTEBSHIU7AAx4FIs5lE
bUAFQY4VLNiSNXcApfhOGx8E+nvu8SJ759D+fVyb97Kvwfe5R9SrdBpA/axk2rmzYk5+CoZ1bPoD
oI0Uui2J1IezSsfSqpunxKwtsp/fiX7bs4o39QiscIAwGhGhcKKYx6e+PUDeOKIJXsDqqcdQiED3
LXG0duyH4tKR3oHWL7lnlIR5+0K4kWIZeaNoS42fD3Q/ULzajzRrj9mRFmI+C6CBnLEZOUxV6sQC
o/uAnXeORrTjve0eSVbg/8KbocVNSzxL9E3pdFtzxx89mzaeKP+7DVSjDQYmz8sRlKZAvXd1t9NI
odbJfJSZramfaY9+3+IOo3CVUzRDaYabZjVaHjsFuyfmX1a9skYSja4EnHfme9N0h27wpQIUASdl
sic3C/YwE9FFu5BcX5ViarZ2haVtjfwW113C3okjej/vJiqF8hHEZA/deSr3cyXfg/CxSPh3gpJM
prCouOe4U6x9Tu0bwhCCXDhp9RqO+pp2LGzx3LQc5y+E2KKlxxttodUedIO/z8Y2mDJj5efz0Z19
iivP6W1eMr4dJAfz+0qtQqQ1q+gTyuCt7XBB916QmhHVPvj+xOm/1FqgEGWYGeK2qC5NCqG90iyV
M5Xp9eZt3I+J3frjVQpxD+YFogvOrq/n5TgZ6frlmuxU4O59s7aAW82PUO7/p0ef9JB1WUBX3852
5UaL/INwy2/2NCRKIg3EkR6uZ4/bmH889vNLu0HbKA9/h1pqlWZcF+//tCo4+q/2NViL3Y40SvTC
SVq3mrDyexTxjYvMyvr9eOJ/VO4vbHXSqAOQ+vpR77OnoCneMIrWvbEZu9hTU+1uJJ95EsTWzLa4
031SA2iTKghQJsi3kDs3IsYjoc7dHdvJIl2sLhjmX48PQncWxbiIS+JAzyYxf3Ry9Sv0h5WgEi4w
E0ZWZHFvtrw8l5OitTYCgoeW0EesJiP3nHCsEAvrSiRfH+MSywbRoZXfyfFaEtph3riAebWh8xq3
2KhTORhl9VRIqHOIVzvNR2Erw6IO1T4AhrJwgU4hArKNkOg5fwe5nbmwsuuYlA6FmidG/d8LDEQ7
jU1/3BRoFRnFG2cPQ19NpzrjZL5mxQ5d/nmM43tuSeJ+ow2LnVC7AJEm8ncVkszlt8OxIvebQMcF
TUIvo9SuUMC4p3t9lSQOWc84eotAwW1rIW8jX6Ql/HAifkdJKCNOKhsOzaEfZiFqeiNICZYs1sBR
W5qW+D+VESn2Z9aaR52d5b+c947CuWZu1HN7f8J5zrZjxmW1anU0IThrwTQ2nS8lileW4wclIK9l
LfSwERJQQ1FGMKBrWpborfat9wDJjgm9DwFU51lrcjsAje8hqm89k92W+Mn5NRjVwlWJELvx0DAr
7Ub2S8Bvh56yi7+yYopJy39OBSeZxHqqT8UIaupRWT4/GY8Cujy95nCVQA9wdg/ymvmZMGYfNjQo
u0LPO1tdP0ABNCt04WHnjhyiXysA+4I7SWkEfn1YxKX3NJdH2pWq3K2dYqnpH+dMOdW+uQSOWGU1
R3ZVIr6aHvGPHyXMcfZ09GBZZZcL1JGRPRMHegfMytOQRwfSN6FNOZMudwniw4vaQ5flWoTE4dTp
N0wDL6jEqa/Zs8DDqIdj1WRQ/0X31gQey1Gx9USB0Hfix2C5bPIJLXockuvBvmPb2OxhxMVOJsY6
UkVPiMK35aJxwwiLiYLvATBqWFKbQ4f7hSvWX9tUVRZhMUMv0H5gzOT/9f6rPqtIkaNnjQy3NSoh
u8A5ZSIgcIaVibtLWcjAoA72lOIDHSLNWzPH1deW/m3bL5hlFWV1iFS4ge+l0NsxR139H68sApPl
oSQqX03WVx4sZ1xTkkv15EVHIiVG9AlBtNwCMD2fnaMRBJnb1QTFAxdAcLGQpn+EgAKEEk51oFDB
DL92REoJtUIZJMSVW+BcJ3YM0vOvHqCzKHe4ShVzhhVstUdOHJ14pcrh0W0leGlRLkbTTriUSdNa
0oz+dPsARC1gjUu4zwoqq5neq2kZojQ824VAAgWfDYDGHOPKAUCzqhYO+wfAo/sempfCzL179/vg
/BNedr72VXl735iv0bog8UDzdVYqvcFYsJBZODwdDjzE8qsI5C54Ky/FkTdKpXTt+RNeeW2jpGbY
jk83CoB0wBgsOIqaFHi6eisvr09qWjlmHpLf1MywnayRNt+n52n2VgI0lMFqP9zBe3oDI1axoQbw
wRgksN8b85aUwoHpCQHgCIQAVADo5SLlToxZLx682OjFIRG8JeOHtQCzPii0aO67zIn4voecQITA
mgwXhkkmiwgj0pNgSh7ECzOGZ71x/CT9WVWUhdQTRpHs9LNw0+blfVbDknAkXXTRSmllkf0LOMxx
NnTdtsn3mp2zWKLVb2rrP/QAJONEs1oeCMXjdt7rSe/r/+4pnMdZrazcZVin32nwFlNf9ncEQ48J
p1fROONlT+tIthbLz7SE4oEsKVgoL4jMDM+2HuL1AnuQF5U5mxNCaSMH82urAWGfk36v+hvGNL4d
ZOevBa7n6JU2ZUJQ+Rij8Wgl2GGKac9faT0u6xnXU4pblIULIP2vaHvZUy6JiaSkH7553IKmsU8G
HdrptEeuMqfW+GvWsFYhuXAau4GThcs1Vvb6TllVUARkpfQGhRkpcZP3zF2gDLURZVjmtaEmME1J
e31uXxdIUt21aSWZaMDSMlvPRBPJ6oX1Dc2HzOszoVQW1NSYydKu+ZGi7gIcid27kut8RqOgvE/+
88MW7Lq3GlOksJTQY2+c3Cv7vl6Q3gDAE91wxza4rFuZrdxL6FR363f4w3kIYjp4g94GlZa3WBlH
2KbUrjSFGS9bo/mPQK983GZ67ByghTqm/PabeYmz64fzrE03Bb2BgXTYxxUZ9yLwDj5Xp/mS4osj
CscW42934+6M3flIxL13Fs1EeCSfvmMFX6tfBgGiR/nHPuG0154tqlumXmJ3AmjZHc4ix7xN5Kjn
t9fpcj33mvxMdMG+giopx7AKd+P4/cOyd1hWXles+f5IjjfJ1SCHvoS5Rbs+P5Sn25ck/JmYJZG1
4umD5S2vc+Tkf75rG721toQoVPP4+/EX28MUxYZNsgQIY6YvYFLM09fAbcDoPaZ27qj0fqD47rGU
dQY2SRNnOBpbNp2JjVeKDsy4g3FR8md568pvWBp4l+uP3QILMVlJSveViMMopWKsBmLxWO4HiyAE
lJXLbAtWOjclp1nGyglAEzwqE/zsOfpplex9LJBIbC9mfE5WTuBx1yKU4Z6suto7nMicPesBvEkW
xlVEsRTo5JJlCGIrYFjgKChSjPgUuSiTqiSuZyCdV0qyrlyPMU4CAzFw2mt1oAHnYuR6kzHWFx3Y
TUZXN9Jb2MRltlQWy2CxiYeziA9q/UxOw/QmQy+7775EaANC7rFUTtpMcKLn+Q2hKaxexWzGQ36o
QfEUbjbx8hzTLjck5dLYJ3m1HDyk2DBdknEIcEtL32yJrL5rLxxC0kbVflKqUMcFosO+WLeSozHJ
vsJxOw+DdGhUdh6LL/RLI+jXRxBrk4hm/QfJU3Zt1d98Td7CYm0tlshGBo0/pxT+1wuHuqbiFzfS
I53RYpC0v72/b8XjSCjLCGxsARAO1Etwa2wwuQi9l8JtUHbqGyzJMeP3NP9oYixC+6XFmyelLeZg
VOWEcw+UEGm/Zg1kjO2aEwbkD8NHLB6lxrNLuTePpKud2uYHc+a4Yvjl5NciECEem6IvOZdsqeG3
xPHw7SCQYj6hNx9SdUULTXaM8virTOOp+4M/LRAIDgVmwmtAtxXI6776vYDIm3A7lD9TEH9PBC/Q
mb9ZjXCVaIdSZx39O4P3vE/zsxKDeDeDJLBBVpesjqB3gx3eqh/Tv5letfhb7WD9Ec3Da47fYW/5
ldq/IUrG2jKFatmup4H6qPE3I6gZVITvbMDqV3gVqToX+bODRAO5hjZ/o/3i5kY5O3Br3VXssYA7
rfI57H/bdzcJVJpubub0q3Jc8l7Ar0V0IJyMoM6cTmv064e1phSkfw8+xFq0DAELhkX8Dyo37C/d
BwXhD+pV7va3OnvSMpBKB1hKWPnfiQYIZxot/rzR+b6/MlKXYBi7vYEwCGrCW9mxYozBV9eYZFtj
DdS82xp2PLjDtUHYT75NyhiA0Xp+GidMe/JA2qARIovHW7x1DaP4tLxszUqO2ztP++QO4sBNW/1w
Q5jFF36JSLSt/FP8yhprq40HqiP0B+9yvUnjNKz/5y9BvBeANFIb4byo1wtqdvS82YUJRA4/wmO8
b11lPY6n02pSqSb9MXMV3In+t8grj091rTH5KnIlPW39l1wG28LZj6U4GOhepqxRKNb36qeW5Cel
uU73fWycFfFx02o7zS+lzvvSRKovdtj1xJ70bUZDR9bIceABV4Sljt7/bei0yKsanGyE04xDatL2
j+S3Tx5Wn48nS9CmL6y3tA+8ia2GRnKykbUaYFBPxw0t9x6YChhMQGbVnLThsJkjQ/+vTV7YcYSi
T7USCA43wX2/5G+f3NDc21koNQlv5velkjyDySXSW+BubKIFVC2CN0+FxZrqGJQf1tRFsh2IKRKf
/VtDno5XCEIrww8YzX/KKHny7vD1KryFGTwhI9BkjozsCdsQp1iS8WDZ1z5jptAjEl/hJWnNhGnz
S8sn6vneBYA4HbpyQQ84yoYrJqAPSUhGyWiDck9UmvQu1j8zU2fiZN2Ho/tbGZ13LGqfCfurzhbU
dGNCD+hFBkY6LS+1wxlgEWVNHsdEg/7mwRtGngC7hcdOufWxn3sEeQWGc00vYi1qmRFp253ZIGK6
L7MMRkBe6mJ6JeDpjycbYNg0lOK8uHD4K6jvQ5RZzseLDVZ6h5S1xsd1mFRp8wkGIrDvoZ7Bt3pl
5r2YvL4x8gUx/Np3v4bqyQhKBgoCTzxjnpHfX+9Dzl/y9vhvWd7hN9kEe1FVvlzKUpDusoDTdh42
NKfrrRfdiNI+L3m5K++H41Qc3Eh+xBh/JaRsVdm0ofjFF7KUxjXt06OIRyCmkRV0+062i2ws7Iac
ALd7w/eiIo8dYl7uJEc5RG8jGmIMbaEWeeaSye2pAk4m+SxBnRNPBpfYdJyN0C222Zkz35pnuVc1
U/lSCBDezeq1N1YjO0YJNauZysF5/+gxrdus9mHnv6LahGAxqxe9yPr73Y5si1tCLgg33YSPEMjp
3Mx4O4EbGidac09EW21X1M/TBzww70UztQRobmLcgzzp5i5WRpj+yDewYPlNzioGAohWcW8/h/LT
yZD1Z8auncED300pVSe8TfkbOeYPj7ZvFtKo1GbNIQIXAxfMaiuHCf+F/HRLePDt3bVpP+dd7Huf
2j5xKkl/fEoV7gwavy2Cg59YvmkUycNLYReVzsDjOW3N/HxX4VnU6hUR15MSuC4IGmOC0Nc8AuEv
51AlvEHLXfRZRWHJFJ1uD2dDiurJiwH+y0Rqe9gU/hc+f+/1TVaBvAa+7Rr1P2DKC+TSzj8He1wF
+xjJWaVMjmfhaYyWd9EcZfXhSjf+3rqoGViOBuHOXo51XZT8l5XLuAWIyc+Nqw8nC0eKQYkqGnfz
gM2olCCU12AbogJeK/U1UccnlguXibBfm2wnD46KubSKOEOV5TKurNKKb6q09zYtt+0UV/3rZMTS
T1b3RPrxpyV4oYUaqdxQakfYoPEo45dbnBvemLHSWKyjalZcLoCc8rYV6NTYq9hOALCFwwiHtxp9
4K1LUfniq8G4hB3VzRIFKYwPASLcPYBjg06az9PkMFd07N3tEePCMcIUF6l+tOitJpHFBQaey8bD
9drGTKEgFxmItqYkxUj907vO7qx7A0eYtKzacXq0dceDYHe3vjH4ttNFMQ2pRIy5i62NnLXxeUlF
U5dTMXuT/hFIGZ7a2OAGjV6TcaiHwXpadeCcXn2iUsI4hd0T9+X9O1uWtOHhx560WUjoXb6UfDoG
NWryqv+93f2a3FQ5szPOX7ViNK7olBTgox6PPnha/jYpiIE0EB9nD5b6O3R1d68jNzx0TY8kcMBU
IXu82tawKK9qWlA7eMtgqWOBvrjyo6t4Kdi30VoxTHQOQ9Ltk6pQ9ZURAHE8GdFzxz/YZODFINRU
o+fNO52GBeFeJa2R8F+KqN96TOevT7h4+tzTxR21MOROjqOnva0fxFg6ucllOjBgWYmndKLiBLVx
lqhoIfaiv6HEPjMtsX8zRpnwNVw9tCvMXJWY+pvsrARkGrpNZj0aj9s4Kdsztv8ll9EnfRtt9t6n
no/KF8CVhrxDSdUyuseTjHgqwwiKOyyidC9JdMkIsCxgaf5nR+DkG6EZVr8k6k+I7kYHCKSWQCmw
Yf3/ukr4Z474jmw5Lozlc/fRsKdIRLD1Efu+KoYyCm54xm0eZi7ptgRjYG4U+0aMfmn85PUMRvVO
Jewbj3VTJvOISV7And4quxmGNxrZGVCQYGs+fk6omu1t3GjwFGx5acD6JqUUx7tUqeuJmZ/rMcAS
8IC3Fl1Sprtqqlzul0sqzGHsCsT5rSCXGY2uMUscKnYxie7La1jUxF2SsPmuT6MDg34HASf3tegU
+nNEwcGi2G6v4WkYk0XeYf4andMydBX8lzxa5f0VWpGF1hqKnbuygGQUcQNU0uJRWtNvRn/fX2Yk
YWFm9jiGi86tpmqtdtvwi2qomODkiaRJFBiOOcOtdIwNY/EDROFG64pV8mxuyfBiYU6intpUBVl8
g+jGGXEo0m/vflxV3JKHJOpNzhgPeqWWpqgDBs14rYaXZbNKWOs7Upq6tkqX+joNSQjzjCXlJYaJ
EiUOjazFE/c224pSjzVik1Ldnx8Me9ROCVUu0L+y/m+D03zv2EA7WxQzemftz+88SN5rNK+ce5Es
fW+mj3p+zXiSc0e3+kR6GjvSCb7KpoVpbmxMUny1E/PNXee2cQ2h1odnn8oj4aG7ITeCPl5pL9ab
k6atL6oJfXXBCtPNBYx/LR9UsX+lKbgSPRWQAKbDgJazXrNiSZZ10ZMoQyOwAIKngjetFOUZ6Xpe
Qblw2Z3x1nwuLqt9u8bISoOZePUNiWaiSgO3+RM4bdFXneGXspUJaHhT0XYrbWI8bVY3G2Po+b5A
tx8QVF7Zyif9NK3MLJpzpVAEIvloh543UY0R7g0et6KlrZ2J8qFrCfmeqjMbZUv9OPr/OmAdCKVC
3o/48qPjYyqsnXA8dqgx26NkuWrrCzNtq7q7ldxpPRx+GFvO7MnO+sGyBVfYJozaUdf3g6O6DnJ8
z8046kXsbi969ppzC9I8NBdVN53FceX45yzMrD4qrK25oWX0B/dXqX4qPCz7NSF9t/IeDc+D1BHj
WD77TtPaqEDOMU29C0uQIG2SPF9Tj7bMh9i0aiMmQBaojmM4503DJFVezRNMlpy+LOTADtFE4Crx
F9ubILoljn3HxY7Bba2yQGEuthMJV6APgrECFN9xvPbSXYpYwZcbdiXEeHrq1PFaAvyaTn49rZS+
Ph8bBXkRP3LOcY4a7Mbr1l0j0XieOjLvnbIIklRTDixAKvMn1YTBist6DGueTVmxB6xTWu4fCJ+P
A3qIecdt6pn5CuYahboXOzFwCvvn13UnU2B3TB0Y/T/4L9olGJAsVak0WxVpH0+G9QQZpI8vZr6W
0UXRCKUEHPjLPCNxlQPNKzyj65yrWjXD//s0eWmO7CnPWPFFxNOgtCqFL1rbv/boAHrlud4T4lco
1BjYyTVLZfSnQVDeQ74hkWQn1SyAaZ5y/uKVeXGSIqw0jtJiC8DPftfdA4IgVxtK/61i3d2riy1j
zP/1TwLK5m2kjF/b7UoJNlCbP/UhYmMmtTIGCWb9pw26cv1vGRhdXUJXRAwtpUoXF0fbR1IvpJxR
m4xHMeKZ8hzhcu/xeHiGs8I8JTZfrDtafSwYqhlWD6eUihsQLqrfZq1wP6EtLDwASaq0sL9QyFvI
PBdDXW2fYeFxHzkt9eW4EoAZZ1koWqRKxFC9Cz83qM0TfVI9nFhhrXfIFj5A9lHKvbpabU+uQGsO
hfo69fSu3vYQXYcBgiEeavSKKElhzZjWrDIAc5VFyMjsanyEQ3MVvoTpg6pz7/I/l64HQ+dcnnxD
6FCLHb7hY5dX3zWRDeUwuwgCzdktX2Hig3zWxiz5owOLODsFPdN5Z1HXXm24weAJKtJ3IAVLZOhe
+uMzkanI5/y2uLFR5d5MMkcWK9zO7snFX+kb/PHPBV9dD5qVw9SAsub3kYvxzyQi2eU1GsWdpmdd
MLNKfW4+E1qulUE/2cVQSwR01M692GDW/2Q7wP4S0VIaHGoSpFFXubBtfd755wNsIn9CRa1yvxr7
ggZhsp0iK/dmR3ABaTnOndHW4AHePn3lOv3q7xByHNlUqfQjf0a0cWWJZJq5dCvAvaiVbKKmPIvq
jLMsta+KBoSv1bDsd01tvptr8zvfpxSD1aPsNcHpCPzpkBlHfJ9d+KhCeIX/jMBmS0PgH7n4zvrb
3BqaBtmSJgqgMMKoVqU9/bN5MSl9x8ccMUs20s9GxpYATzr5QKs/JLn4gH8EcrFRgBrAT81XMgis
fG+qRkViQDVj2Y+Ci0fQ4Bqi5WzR6Axm4/99jw9+rae1LeLAgZfUfJwI50SiVDe8i0GHZuJys9Ca
bpesVHuEyus/t1auTyKZK2HlWliM2fTEZZUtWxMX/pP49TQrqMnoYcnfip4HKWOUEmL6Wx1GpyAj
jvJwZPYSjspKqIhTzi0amTjp8BecY9rtFKgPX8PTECH723YVGKUryVBxv+rdWDkUHWpPvxw9NWuo
BGmjFWufAT7bX79x9wZoSgjJaIPpMnv+XcSt34KYcIPakXPoIXMavRtTsT1cMrZGf2gfKTP9IISF
jEjUPIdjBPVM5fD8n2zOwFhnU1T03EZMTcuBzQnTdEPMmSfXxodiPRSEK94mkTYDgNJCO9E1CkdU
AOFwM+fDkVj8bqDA/Rjmmd8IxiAlPKe5KVzYmMUEf75BD5f0h2FLBybWDQm3NbXnsv/7DEn+izGA
viy9fYDxUzaritc3IXO1SCQLCCvlGulPraOsTmEHV4L9m4AJXQiykSy0BEp6F88D7+Yoi5XOrsy7
k9Ma1NP6rdQRhsV7kA8+4ehR1CxvLZo1mgDPEoH4/j4b+Hemb1BG/22tqEKo0syFF+ar9USbQAXT
DUZqDPwci1gaE1pi2phQGurbL66ualIjaTkBh4bNOtUdhkuQDWssyVMO+4C63+lG881ABilKP29B
iY8zZdyQNQF6a+4o1Ky+bqSZ4oVZItw9oCap8l8YW+eVZnDEVQOWNvYDND3hPIu4v6gslANg0Ld0
ghF1B5mg7DfapUABAVrp+x3/sU0GX82vNXFqjrLhwCAt0Dknpk1JrGAP/t95gg+Sv3tdqURbxN8d
umHvQjLwGUHAiYwJtdnDiFoyMqJCfNcVa0yPX2Bs6vwnCM3liTLkGZksOghh5ucWIU12azfY1RF7
B3NXJwEbp3D1YmdKsaJpOxj1jDure/fS+ntk//w4ii8pMCbLFeHqqdQsm59DB4gonBpH+8K97GXI
04vhHY2rVKCCo7CdqGbYE2O7Samwd6txkV6WWdbf8xjlMH/DWragnFhInQsJriyAPVofK7NCdxXI
MEKDCzjSz4Wf7tgoctZyz1FSkAdcilvroglUuchjPJYcUm6HSKfiGK65HS0naMKHj/GS/lFBiSYG
6VYWnw+l1PZfOQZVOAjwLCoSomBtYNyITnslS0lrVVzaExGRSE6mcYqcC7iJqWag/fuda5/n/cuM
0/MJYGNObpk1aBPfmHxeIhrLXTk57XqbAbs0jiiHoQKX1ZvSbS5ucPokzZL6nw/bbYenPLyNI57r
VsuwLEbSlfkwln9i0NlQiMoYuHbVkWXOoigXA1sAtIj+jo6oNcB1jeEM40wdGKzk01ot7HTkNz69
GfiOXyaqwl52TEwkaDbxlUmoN+e+6G1sdoMwwxg3azveeNGx80+CTZzB3QzDx4YiDGiN9DI1doic
wUAcP3y1Uw264r2jvhbQs4IBje+soN/qDJNzR3XfDhSBJf9JzUAJwcAFKfT/WiRigLjdcVOxLo7s
nkZM8e5S6wnyoZYDCDCG8+vmWrBmjO19STBzFCXS3SrA7sAqVu+KmKisPgRofQY4sdCV27klwIxd
GiJjl5KkXj+tVhDCIode6GNN4t3wmy1Ffd4azp6YyNsjvYds0F4NOxQ71H6DCXX941O+j++m4UCe
yRRYIgrwbVERKuQpSc8ffwz46FJwjpg7AjPXMWGfdPrJjCNB2eQ5mqNrBceem32A1jLFN626+LFD
sGpMRVFXu6dEqTpgpR+h/oIYfmauBcFhL5imAw6jrdLgvWJ67SMlPCzvZ+scvKpq08PodGWwR6rB
EjRa4K6MOsgyTfO31JX65jVGeVcST7Xnvr9KAIW/IA2si3OEPG+GEvMH/xe3Le+QK0OAPPwO1Pfy
rSIqeXruZE8On0wVpDeZV89JlbIKIHAC7JJdfhR+CPtwZivswb1da5ammMi6RxERnCq0FBpInwwx
+nHKMiINmG/29sA417/Ux4VCCTG6JPk9AHRvcrCu6I0IlBb7bG62v3MyY//OSkn+vOSu0ZRvUjET
qxp3XjS9dcEnnK4Mliz6rzL70xApxiRtszsTPTvM7K0ySyp0QOM45vQBsndNmQCv8TFaLQcmTKcj
bqDbf9xTJMhgX+byF+YPhmUyxpzuEuaAPEgdJt0O9a9PTCowk5emHcEGQ5eDwffizTNkL4hhih0d
QrZyEtM10c6LGich2zdP+6kVZcnO2XHRAV9nZv1xTI/wCTUStKMfrqI0D8Gqa42VLWqVuGhXWJU+
1x4xpmrkTNYgijFYvhzpIi05vHo8mwpC7hEaf63pdh9hVlVFvjvYZHrPRi7riCZGTOreSNFQqyS7
RCiMy8wthedgs0AVJVQEQOmQxe2w7VnsENZxDwV8WcgdzpM96oyaV8AgncxsI3h7tMerulpP86SN
DMIyHTNwlPpqBHriXtKvoMeSpZvgnDfvb74feonua/OlBfCLnNjlXBFUT2q8m2wwc+kXUNB4DhUg
6966+o5p0e6NsZihZA8Iq/oVzlfmC4MSsgHEkv+t+pxW6QVk34md3S3TgLpiAuECWbCvpvxQt+mE
6ZrSgPs76187nu8QXJAVY1I3u6QHlPxkyMR8kYkRrYDwk7kMZpR3OtK8aME58gu5paV6YJQ52dlt
q3qpcBx13JuX7QdFzL7yC35tAmkyomZWnB6VvXwHjn2KogJqXDsDbFDsL9IbhKJyb6yLey9nG/ic
iZ/Cmz8CmZBtbozDdcO5uJs57oNBOPKlgoN46Se3A+noj+8ANZXNKg3rgF8jbTlzamUvyL9SpzZr
KDdQQ8nbBYk0zOe+3OqTBUl8YdW2rjOZ3rC+M5wADbv4FMAhbC/YoQv8ZBPkvCVVl2a+8mOLgZOI
YE/VRmcBpEXH+1yh1OybcbHngfw8CPejxpHxyBD7cjysnFrNpWWX6Hkig0txjTlb3VRNQ0BPCruL
r/DPyZSJjMKzFJ14A4HdmH37yb+Z2yRJS1WrnyIFIjfUj+UhXz/RGMeaq55cpwH+K6sgacCkWp7T
qHqSyiBeykR14ce8AueyfDvf0/wbHuie4J8RtiLKMKFBqmNssaDmVPRSPGm0xq7cT2A0s7jORbmS
nUttBli2t6MWI0w3kHBQYReBeMWqBelfJjIbHsgdVK5DweTOAMC2YGOWE6FWFNTS3vSKkVJ58Irx
vKmldfaQU3jNG7fqQapfgJAyZOBgZSMF+ZwKbXWXQztteOQrRIWrb968k+u69hoOWGwWmLJjAMhi
RylY7ezNYBlpaEmf5FYDhGMV37+p0c7I0Xw8BqhBFNbPagjg1mkjqhjA8J7xee6tAXjR84cVRPHA
oKwDgkkiybVju27WDVVraPtA60NRhTxxqSY4m00UwgGBJwJzwgsTulp2YeeMy45DT0/VpVyVgI3d
k1kL/vZwCVBIE4F6qNwvKgoykbqJjOUtduJSW/jfGNY1AV2AuqJlIq9LFOty+uGRz8beEa8cx+fW
yPjdyody6r3rbU9a+3Jpt50r+ruhKektkfPrnqU3NbIs61MALFj13mxZVUK9w+pMXracB+5kKUQZ
IkaAj6+K7BFyeUW9rRGEoWl2jBnWlPecAEFL7oMC5pMe9rMbjQFKab6vhuxtbNAieaEjG3lUPFJd
U3b3gbi1FsVe+CfDmJhRTZKm+C/kboTaB/bEiAU7L432EZSECtGiTafsBM1HJ3ZjIf4hoeey2Xu3
oFbFGG/rj6/J+aQ99LHFa1hE0/8/K4EixBxJIzJeOs7OnVbBmwSbLfANkmMR1r13VKBdptrA/7+L
XDeDKPQzNcOCf2aMxsFR71LUctsOz+nNcyfevAVDrrmvgwW3rbtQDFn+vN9Da2OKcnvVt7+1ADxz
wFdPVWgzmDdZJpZvS4kRR/RZzJ5lUT66IT9pbMNa0+GZ1gknYfKKBNiv3jg7En/bhQrdDaA/3LYX
geZkxPQ3W0Vj/2J4DGy66I+t9vp5azRYc2WqG6+W6nJBE0cXqkCcbcqvLmeXOOS8DmTUqpBZL+/A
UIV67Sw4SfDsjpOWcYBUPUI+CUvfDa636pwwh0VazOQ9wNhkG7Lo2gXqWHuNvKZSIb5JhNisqduY
e0m1laDq/0/9op5k2OGQwZBo6JxMMFUW3t4XobBVGWLtsMPsXUTl05DQy9j6A3E6LsCA0jNJF7gK
tLPuDUw8/KvJvfsaA+qR49X6TxFq+4VciQUVTmYB4VMtrFZkZlKOalztuz0RUsMSlO1HgTZnItWO
c6KgcLQ+bkXnruzbTMd7QVDC0JEkZUBIYYqyDI95RAa5ZKJZBRULJ9SkfD7y8QulwHg1G9uXwd3q
ol7oh1RQx+67eyEhs+6YJmsrZdjsmtUY478Lr9IMy8VBZOBTcXoRfTusb20KhOhbqRRZ8Aqr/mS/
XU3gh2xRqaT7P3ETSBzfWlQw7YR34KE5rbkXIu9+cKRdHut840C1fYj7ahkSmpKUoi7hOZJY34gX
YDi3LJdhKmGQ48cHFz592oFk5zc9fgObmCOUci/GjUVU5SiWZVk0tUbZgH/CORcgJ1h5QB8G9Xss
mG9Dv8eqD0Xvzu70Fi53SSwMrxpz1+PPtgC+zvME+j2cluIQtsRDxkpDaQioY9LdlwoAFpS4t18z
cmaS+sBbt9UidcCfbRgbI6JGVvGAkWD8tNbS6AVAA4cvI5TkYGAKLkBMV4XZpauwnIbNlgGmCqsI
lffD/5BlUF65PD7x1tMLY16ODibRC6+AGcw6kaPaW4gKLTV5VlQonITr2JVLt47XXSMPHyh/uSt8
t+yzY11yBx7RBi4tmUglweQeSyl9etDYVjDHakt7cwKmVv87PnktyW83FPgTJvj7+7+MMc603BiL
13Ad3czs8QCZyE4RnCwI/dmM2tXd3QgkNbExScnwOeLTbm4u0+q8+++20KeGtygXhoKYK2bOiBNB
jYHRA8GAjGDvj3LzwBX1vmHI1OW6HmuGZ4x5QwrYaultmniTdjhYtRc0oCOYcbjQ9YwO2Xk6Wy8s
M2l6zdLqmQQPMViNOPrJPl7x755sVNnTDsOLScFhnacX4CLyj+gMWZW7Xvhx5xBXvRhfZn4CbpNr
wB/a8WQz+jpmAvPf0x5bV1ewJbNYZchHCcky5qRw0iWAe7EOdANvwZoHdyvTBDmWLXKfTMMsx4Ou
h7rFobm9N0c8grSi/LH1OgkQSLYhHWLsz/EP38pC4BmID2hPWcz046xwrAU85xldCtIJo5mSFw2k
/s17OStHztZ+lR92FwLQ17o7VBrtApVnqDQgPYg3jq8Ma2wVfrZg5tZkuKe2uQs/wwgrtbGo9fm/
O8ozFRF/QeuWF0vQB9THfaPbZa022wUzIDZAWsQCDSGomS2JEPk9DSMGEQ1OOajZ34CQ6k4SPJNb
8lN3Pm99dOwO+2L6h50Eq61l8cvGjOYkNe6dtDlNVI8garFyHyqlV8pyvn5kafvfndvUK4nRRpqG
+aiS1HkDKd8KAP9iDCBTZt+XZrvjlpQHFQzs+6XrF+A/IGz+LNKGMRTZVtFU7lBoyQawqRVM4dRt
G0dwAiQQ75nOwtA2IdQVV7sOT3pivDlQnsYPQInDyet0h+psvrIAASKlVQVVzwOyaAOBmN3xDbJR
biyFJj+tkeKvXMxlCg4WJ71Ixb+WWdWrzergmeZz3HERk5b+giru2RqgLgM2CyPKTJBrHnlWHMCl
qeDHcqyUPglAVhgTGPT7/bAoJ7BICkxnmN8Lg/eIjUsXHixwzxCBcL5uOT2AgQJQkLUR8Ew9vZ5j
B8yxdEGdHC+pA9Ssi7EwqcNsb1e/ctmV5Vs80ojooAWpzygVhImrNhGhJN0FGRf6UFd7HA7Pps3P
ItSjjYwG9RBNVe6EogQ0VEz9Nsxu/L8GRdF0kaBITk2BQXnds361KHU8epXVrMpl+Ij9eaCas6vi
p9kIThguiDIjKzELis4PF9r6RxVSJfnMzl1G0CKl1PRP8hqNBScMZ6VLTxhlt0i4Ulc9CyV4sc0t
8wXZn2XsYYRfg2FTjsM8ESsejjocb8g/ugifcgnsyimmzMlXXtAo045d0xC3P/qKT0w5snp6pVF+
RQdMSeXdB+PQP7Qcifc8RdsoLBw/7FqEaMKo6XNoqSXlA++9WcOJM6wZETLE/5XZSEW3TS2Dc+26
2BJMTjbDGgWRNAVnNGUXGMe7zXkv/wrRDHRX8z9fK/0VwvjqJ+f4Ut6CNLxx2wzLPa9sgIPRKlIy
DKfxkRIcKZgt9DYlGFxwqxAVc1lTh+5Xe1pgdhAQq9B62SQwZz0kYcJbyq/AyMJSKDQQzV0UQmno
9KYl5bLy8DqQCvUvljqgwModY9m0IsAt3TU4aW7n/A73R/70v3DezCh4dIZmL4guaPHlE6JeOCLD
zp3NBVFz4srGVM+Dz3RqCocCBupNSFOI1anIFqSHhA6mRa/doOtVDBVpUhBVfK3fU06oVWpgVXrU
2Ev3A2LXIhaeeo/PBbH8+Uvo1+4c5yF0hl4G8uFFmzQDguFFpWgr/8TfuobFdCct210r1lLRtXRt
GnCee81ppzlMVRATs9S+WnHP8/5LGFph7OdoeGxlw6vqN/xZNxWT15bib4WWUf0KnxfAG19S2Tyt
kVOx2JbFxcDv/XFt0BYSFx+Yya8SMXxneCdIkYmOJLd3B333apKN8H854f9LF0bwsZ3cTlDJPhD+
//cOFczo/GXRLFoPkXV3nQy1EFASBN3v7VIEc1MA9L4HSkQ2o5QjVyUgFWZQRlNuQ3JYouYsrsIa
1iX/u8AaqSPRedcIh3n1Gz2CsaT5SkR5NSE4/1u/Cin3+6atRewtEHqW1qEkCqdwuEOi8qOWo3GE
Rszizk5A64PdJMbx7mqu/A8Tju1HdO8WjNmnbK0DQkA/orQPbmYULNc2Inkky1Qn/kZTziAPPvJF
5OzuRpIDcR+gfw4x+J+n/oHQylZRBx7inoYLOT8JCggSBW7xiSdhMZ3Wo8fd0z2vycYRQ18b74gQ
jjkyubek1a0n4Y61bFYDnesMafMtIpDSBcpwXfPrdksYyLAg4PHeifpit6z48Cgi2PVL/4z8wFor
15lE3xh3lXah83AZ0QJEDWCh0MAT/C1HcfiIH1vdviVr3wRY2XJpaF7djC7TamodtMYLSiTxvHhe
SwaWx1ws6O9gx8mH1FUrnEWCquKVJ+cb8g+QIJ2mvU5wf1XpxaxmUzna23tVZILlDe9cSr/+UNiS
nQD6knzFqZELzHLvMjIZRFytJZIg+nOoATYC8zQm0zZ+etwnq7WqAlvPvpjj1qNk0/4a4xvP5bHt
+b3bxS43SRuBq1VVEYrbF2Vo8pSljD1ate+QdqapDFSRaHTl4jVBJPgUa1vw/jwTb5DrIgJ4VFg6
jz0KNs9Q7ZIBvdZwy0AU/N2BLIbgUViYbdbfi3P8F/VxwHeb56DDpCxbvANdFAHE81OkNiah/tjb
HD8BzGH1BUMcwY6ZQZVL0b5sBh61MVlPLVJMpd8NSE88NAgM+HpGqzuNT+mAajjzxqkVcIJ7fm3w
3q12zjyC0c0OBnDWiGFx7wm1UGOmXe/QMe3VkMLMo8+6HC+3zkknMitXVb+M83OS/Qu+VzmeD5Rq
T8U6mxU/LHXm+gcudabndvP1b1uLUNm8BfXNpNht7VrZ90m+ZshQxOQDsbFvVZMO8UbL3+oJyL1Q
IIKxl5sTCb5KU2H158VvYLIOjgbEpwzFdo6VZhi0iYQRITo4vSGC8mlX10TjhEueeR+cyZ4L6pKi
WZ4PAmFLR77uPJL6UIaGlbGEFG+yJcXZy8mDfZlAy1+/ZYk0CuCu17ISW0g0wVt/9TstGjZSrmeq
4IJwM6ia0hWTGSV0HsnZu63Hwr9GB7pc3FTSQliLdISve/1k2V5sijP3n0aBYkMdsjQuZffbKl7L
ClCznqamDJz5g+ZeVmUDI6gfjDVRLrh7r8lsygK1+RaNyzee3CS/Uuihar9cPuh0f6H9a5kvLnKP
FOQ41/+ELjjGArjX4SvEZV7j7DRuxajnarDcO8kf4y7ZPl0vHr7eA7haFsXk8WxSmDlq85k6agrk
wtFVYO1v8Lt8vWs2IeTPUmXR/19lxLYkK0AndDohIEfy0N7UutyphBoFblHRLsS5dWs4jMzByCJf
XxtvgcOtFnE9sL12Bipf0QqInNmyMSDTl0QlzzUdvwZ5851jZ79BJ4ACEGTZ+K+QxhJuKXG6Kpu5
ISWNRzncPH7GVCx6P5IVpGokyAH0sHVOcB0zWpKL/I94oHxv/8cP+U3XVsqgEpVFkOh0p9ac4JGj
wjayhCDSlNeRMXPJLLJ69cDCtLozThQ6CVXzHZhfc1Dqo/B7nd6LHV2q4KrorFoHwiXnEBP/lOau
hlAbFBs6ql6xb2Xl7Rs3NZ/P134CGqY2DNwgPU4JimCx2/3LvlPx4bhoZk5aVtY66L5gKNpBsPx2
Ej0RITEhvE8zRlNUAVDNAAd2TqLEajud2xUSEzXDrnHq9IvJfIw2tQJ+ctHqzR5nAX49Dl8oeegQ
tJLLlTUdfLS42EImVBvO9pQtWZph7z8hKwLGC545ZATQfJytJkr1WubEl7NMDi5DwfjeEfGmOMJT
v7guVfDBgMEyC2wm99j0CjAQfaGd/4l4F144RWG/A8ZSD2b3Iva718fFzGtGMDY3NPygRPKjWA2h
QOohvErEYWKCzFjvGAfuThrYp8cw9TdxzQh9dJWekHU+78+yXSxDQAlTV9Y8CzdNghgFY/HTopeZ
3WRQTpUxTiUSEgioSXAT5N+khU+pulMANArBsPu8q8CVUKshiuahLqH0EdYMOLaG3D2LgSXZcHeJ
s/CB5LhX8HpWfOHf2w5LPCKJ6H248TPwVtFD4utKdDFskDQimc1QTOsPCuSDsaipw3k5bgGB7vk7
MKZzlfLyJs5COkKviv8+4K7AriwKvM0lhj13q4N9S/y7Eq3zIGLy1M19C5ZssNisBeX1d19XCbgm
1omoaO/CE4O/8EqPQ4xA0S2+Phnjn3JaxVUKiZkOeyz1p98sLhqrrSRJXots8RZQ+R/Vk+P8x0Vb
kDK9Dkc5wTByU5dtSmuTObvrtAOyT3CSS7pu+dnf6f6vbGNyeStEXSLUubBDLYodperDrFaZKi0r
NeqT1WQPSylc1feTJ5u50uDDqYToR4U/zpNJCJxTBzN6NnFu3mlmWKrjKe3PUqOeERLWuJLmPYch
pAelsD6Nui5gWIKKHRSlvwFe4KVE+BPtloQM5/xtMsJMZ+N9kYg9r4ARv3gJsaFjAztQTaeOzm6O
Ly7TUg7ISxWdB/zy95icEHQfzU91tPDxhMVGnqqiOoZfTZvJL5dNzH7pBXUrAN1SRogYcVjx8PeF
aFAnN9NDi/HgCeyENoJu73lj8lVN74pS5f3NE7pRyrbgngiKke42rw9ijMJPe0gjojI8xME2MkvJ
zCw7bTcFD37q0scEFoD3EqPgAhvQPieQytuUT/QSOrjsgXEFjnxnNrNPRpN1i2FGi9Z4vC0yqGUE
7AJHyJFov4bNQPpFuu85J+j+4b3bH2wNZuV33ugUolSEuwasG4rPOAM4NcoaQ3kA/ObycJLSXPQd
5sNcLkIZIJOtuRB8VLkSagET3DPqAzw5ZaKWJ7Dltlvh6A6o1SohxTOOQlFlD8HE5ayLymK+6+fl
pv4GOCPR7+TZFA7O0k3sPOPeauNilCd5liCaDq9BwaLp4FWdBe6W3L8PvTIRMb7WO//cw6M4GCJF
AHTbH1EMiFOfz5ahbh8q02kq9v4JaEdCEUIwBQEjHjJhp8C4BP4siQlDwthV4CcpnLjF/cy3RPdy
gWW8AiGRUV2KRTkJL20mgcyprOKhO4Mczv7ammu0LIjcAf43ir23yAwkr5SoH4jAr7mfGDKmSkus
PwjuaK2J88jqTncjJP+ozJPSpUAWwGvlzx2UsYlpfgqJ57XhIrER0DnlX/UtX6+v0IV+XhHL9F4B
2JkdP/i7FXxgrcUDiO1qQ0+hOYydtBp53ZpfkOu9unmA67jw/OOSawHDdKmK6mCUK8dsYh8D7tVX
cnGIoC/7AGAO0V3O8nO1JH9pITCxRuuAXJ/6732z35bjfnM5As3WUntfLJ9YQVve3BIFeN8//qf7
tZMlm/USnc+WnONdW0gDanQlbaQnntT5ThypDsxSh1RRWO/xRMgX94NQoRAc9bqvme/To2GKVFQC
6vgTNiDWjVx2WAZgyoMubd6CgmU217Jx1IatL3sSaZEXybLUZWqrTz23H7rMggCJCnRZjOzrIxMo
Cf8ZlZkk5MoQn9OWaBiwSjVQsWDm2pUbWktLzgyp7J1n3yeLeFe2G+tP3KZeg3tNyBdoxt8nTBWi
ECOf9r2ZaYxyuTRo6tTtgVBB0L0mZ3NUIC0KSGJj8ORdMV6BxPIu/LUihltYa6/WfOCXslO17nOF
T4HQXZ/pa58DF1IEBM5ci6yw7ecErDqLejPpFYg0qb7yEE6dkmu2q2KAqHd7cahWFkHvauk2/ifc
YQe/Dfo1CIImJWdFV32Yg7Xk6HXof8MW6GqXdBT9Um1QZvzRhQ3SOnZQi6coMSKZSpLUfAaFLdGT
76fNvcwmYHw2m4b/ds3AT+7bJamu1VqTLttTjaZDICuMaMxQwc69jWKMMUzto60g9d2q64/qBfjf
SbnYS9C73wE2djTscNsUCgOkwTl6DCzNAeQGLOulG6NSijDTw8O/CjrGzzNqQ04aoliDP6qiJid1
MXhzic01kCscEyfV/f5B1D8cuG6K1i+fzLcexLmwOCe7gJtHcUuVjBoLg2wfapRmGGkT/3U0f3Lp
Qe8FdE24yGgSVvnEmLKfHs7PtLR3FU4CRw5uzTd2oJDVxhiSBKicdHbWA1Ymz0zTTgMDLt9FG0SH
FBbFYSiymxz8P61SJhKKInc4CWnhZAg9dfkXaW7a28ysgQJ5kvUHymTAqsHfMbgnQPRh7+c8yvlE
uvPmjWAjFhrgN9MzoGQ84oD2Dx4O2nout5HOgE8g7PFPlajCAGzhl942ujYJxhee5+Lr8Z/ZFTHm
gVYLCtdstJEo5thFIiVqgIFWTdwaGhh51Ib6On+O4N6H3yJZvF4ASjx4wmaIK4ArbpN/nZQBVVHs
T3EVykLBglIL1HTw+6iRrE+T9zWlVp3PfU+ZZw3wyUreRDpH/Stk4o5ll9W9LJLO+Rtl5atfZvpJ
FqzKd6wLM7q6JSDFRw4C8Kf1MlpO8AY/8hf1d2UKVw0WXvNmt1EDzcW6z5rCrTFFmicxMDlTInUQ
nPKR5iGvSCCe5vDDB8Pekefo5ZkWCdRbNChqm/CW1omZlJFEFiRcNxa+EvgTs1LMIlpnUXmXilfm
ZWoTxGd0DsYoOqTco3bYJsXJDS9w1hyAPXxFFSUjlqkboKZOe7Gybn6fwt8RC7JJ59wRpYNu1K6O
DUPAt4Bzqh1PTp2Dhwa0Z+mAsWNLvrJ/IhKQXcQIuVNzq3N3rYyVr2muvhFwKmyluFMflaUm9cSz
uFsw65dmI5oD9SmBn5Rge6OfLFPIJcgXnmoBSm373se5ZjQEKBrmY/0uOP+E5pTwK4fozGLHqVgh
MPGYX1Qp3ahuqSaOdYa1gDpmTXgOqm1PyBStOw0ATjBlMuHH+DuJUuQgIZcxc5aD9XTgn62FyCAi
cysf1nDe6AGOfwKNUXSvZeGMkYGifSZbpHMCBBlKf8orXgal2JIR+iuvDmaIcTJxPBSopZ8qyLGL
GuEFb0ZZkAqa1FcPqmRK3eylogA4mIkhuOyYczKTGOMOw+jE+uToIoDxvjnSSV8M0qHDQs1keNMS
lk+Dp6O1GQt5jmUeDWG3SLyUQ405pxA1tqWDzg8LcC3KkvqslXs+k8/z6j/XgLlvEYoAV0ZgpN+H
GItXp9p3sCfYc7yrm4pKic4OGDNYxHNMfuybYvUnV7PvbV6FI38NdsumRV4aar9m9jFxynedhHKv
EF0hFsu28sH5+Ng9PUDAwlmJkoW76Mcg+Hnt3YgDJUqpypBuffdR+1x8+QKDmqgyrPVAwbiQvKFj
e1As6Ux3I/RNY56p5tfytX+oAF9tU/S3ZLxVyKzWaGw/b5eeTr7fCLLqXyR+CpfzgQsZoxpngKVf
Rl0U5iLDOK4KH73/oMcmdbjjYkZmYJnGbKkVIJhmn8XRLf7CjDIn7k+KT3NJVxR1XuhRH9jAHIoc
W0vy2jv4CGwZJ5CQZMDRQU3KEhUnnkpQ41ywjlMypys1gyXASduqBk+EAw4BtEvwL+Y80qZaizUs
rU0utSBLmrz7B5DK348o2m2vZGvkVPGPQ6zZDP3d9c7jOOlye/8U41mqm3A6/EFY4CgAg0ELnmRt
R28oEGH0StHlLwO8kvkXFgS7EtJwdaHx0/r6tONgTQIIxTD0eE2dopqRJp/837jOHJPtCJ1HsDfV
75dWzgNLFsLgxMnMcg9aoJ9RH7aw7j0lqai/nohb/4nN3JUpegMpNBMVc5eqlwLC8ME5emaexuzg
0S3U9MdypeF8Gcanr6RWdwn/8V201Cre201HSV57hDWHieocmy4LlL8a1P66c2i+qbawi4IHYaDO
mVq6zPpiaNUYfuJ/b7v9RumQUHyzGYTcbr3n4WUS1t3rAdwhGH1jK5NmTLu+C+97NIzrpE6G6ZD+
7CplGl76BZDLv5QddGiNSrgIel7TL3tigq6aD3Dl7wvPXVPmgVhu4iwGjy7veSP55fWKxtxwUGAD
o8082uK8un7TCEyw5JpTJM9wZJjj3V+hTd1db1kUXWcvewHcpuu4tehGGNlAX5fKdqi/ZLVKxN6m
QgwAf21vYpLqQmp57vunYIwS3LdLodmDiTLEVcFYw3V5Ni/5YgVZtLxi6RDRqXq8jVR3kmEwlRE2
sWbY/jVHQ5VO8FdKvhitDg5x4tCPsKectaKTYw/ctBt0lrvL8ed5QsCicZooXtR4IhTfFmg0oyFZ
AXEdOhoIlQbL/Svsfpm/hFAoYOvFPpBidKal/fz7YGgl1crXz6mVbpIxKoh+f8d02lSxQlDVMMMT
eaeSbSN0M/gPmUCp+G1ZZ63fiRdRUf9rb1ytk9UPl+swwqfrriIWnUO489UtpDcaPjv07OM9Ne0W
Z46jxMKY2FSe2U14quUu317iWtgr5CGRiS5BlPoHASotJTvPYFQFx8gmdJed57u/HeUZff9z5Tta
5TSfa1DjvMo2pPZQNjFnvycPQ6DD+Wnao3WXs88L2ItioT+/DTrJ+2KPlj1akYwY7wpbUxC+XAXi
CNUYcgMlSdWwcks3PuSDpM6ZisJ5jgib4ApDVbz6haJWUVOumdpmKUaSYIlqHHy8xRBTsjVl/765
XEmT3MM31bBT9UUdoIDVYql0Knp3KDqCJ7jQTWxE7AMAdd0adPd40bkj7R1Buy0/cwpka0c1FJFk
xHzVDR3OUzhBT5gHC03Kb05sOgZ17EsnWb3kvKSTFMTvrWUlyd5alwOSedvzcPYgx1IONW43Xl/y
dH7lHaVbpfSo7gZC7Nq4rEuwzPxz0uCiUctAjyc5nG+ypaEeKjBTLD9zAzWU1WEduUa680IYbEwB
OTJQBoQPahLCZet5ej2INgBOW3WEG8R03g9SBlq8/wKqwDTm3WEsktxo1mNIMe8TCJh1B5kksQ7N
p0Ex85IKU2i7rOzN55SrLkBZOSWyBGL653i/lANTO7IBqDmMGDFwyjXIuG59c/Jp99QoAtQZ7r9n
FBxwHkH0b+rXFlmhcd1w0hldZZ4//qGshyzgM48g+7W+/6DD7HdOgYtI6Su/WDqIgSmNyyZBJkZ0
+yPnWCtYLilPpBN034G3jjrZbnEcHUJn6MZ+QFnCIUjVSMzS21kTyKdXkyQqX8vZ5/rk1rafqgS/
1PeVBJl54XVUZs5Oa0gsjg7Oy95VyRJ7tOiQI8P3kIXo50fk4qYoBqO5M7FNIGhju6DPqxDWzIUl
Pr/xt4Inr0M/9AGa4Zyw+3OKu9rQIba+wGbtIo4UAjmTmolaQGNpo/ehjUXNDWSwhyRebnfPDCpQ
sDm8d82WmRe8rCYoJwUdj6AyNPl7z7SYhWh6OjXcPoB9XXCOm+0FH+nJQwHoPWABO4BDHDCT1Rql
nphlE39Jn3+QMXfwPAsKIU1dRZfW2g22HI5+dJ/W+h4GeNEqgn6ZWjyMe8RxzuDO1rCote8NQmi7
escmY2gSSCYSx2Wi3lYjWut3oJitwYJVfewpkkgiMe5DoaEb0wjzFAts4KVOVC1+bj+WpzNz5aL+
fSUO8xrarPF9q5wiHGd61nP6tS0BLt7R2I/yQOd9zwkRFLLnBhZi2SZxuil6iFvNnxO4ZUXCqLEd
CSRvvaCdwAk1D2vnrowf0oVSBBi4YFZu2KWhe9654uB6uje5+gBysUd9Ub1sNQ/vivejGuegW9br
/uB4bfTR9nx0GZqekDYM9kPhcDyejg5vJoIxUWbHW96aHG4npaaAWHR50lgi/18VQ6gbG4Jn2waT
ntBEhEUMAc8RapBP+1PQSMuIpWb01hsdVHphad9N0PrcFPHEhfMcRh9+/xKRfuC8xvdslV/+zrih
l5gp37Ix5+YhpuMYXTOvn4s5nGI5zTzr4Y/Kkk/45edXm9aaFW05E6ZhQSyo5Q6j09I7KXb3o7NJ
D5IBTrz5zoRmtkjpUQ4KJ6M4kjE0epzjp/0aiqrdPtAt5LkMvV/WJIHFFYQ3c8jUbJWF7D7Et1KR
iVozG7iW/QD2LvojUZfOcuZRloID9O/DEKBKyYNy85R2qbVVhyqffAsfBaBOzIWQRtQzitLwi9KY
UQAbV6aH49w0Gu0F3eP548XgRbhbXERfy850QY3yqo9emgtJk75nCLHd6BHAVls82oMqSdQjCmOX
bctiggzshuZrQEQc4S6MXKKAmEoQ2L2vWKqUnA03Ag+zCxx12z9M3amXgLbvh4mI3ulmAabM1Tqb
VLYP195hd8SaPZdegzBKQ0fB2dyP7oPc8z4kdZ2xCAgubUKr0ODbTLsR5I2BXFTuoeWUj84cDpvS
kjHdk5lydeZViBXqykDTnhYc9iL4iZT2BO+B5yStcvAM17FsDagGAJGeQaqk0YeBe3c2KqXXvmq1
GMjl7F6bRretkIdxtKAW7PbPqUvyw6PAFXtHu8SQUfJSDzDlGyPyzUQ2kF7W7pESoR1p+clk3xuw
g1PtrWr3daw+r6ZWKSqLgLRkKpfvZd1X0xzPnubwNkrIJRrHjvgTJIBjZOQKFKm2zPzYT38q196N
vpbqjYk2SXmLT4ycU95+rDcykibgHFQjD9BEapRzHys36WeNkRB2rne6q6E3p1BNQYXnLqCLryuK
Knh8YlVbNjFsKWDtgZqJodV84djiWV3Rgqam20TDgV3v++u5TSlxOAoOmgIe8kdcjMuirhkZXjLk
vXPMt00+dKj/eYIT8EkhM6Ov49zsFSzsM0v+/VPdyzA6qd/x7rv+EGJTDuOlyw6k4Fv3/1Aimwqz
CdDPcnuYgf5wQiYQfdzvHrxetAv2mL0eHXBN4kAAzrDbNzZhuWs5nmTqMr7MVnD32g0ifBlxhzjb
HRSyPCbAIvSwgcE93Zldrpdc7RMsmaGx5rzGGifK7WFTP/z09cxgjy3L7G2PcVblTgsBmDgrWnak
4LbOlYZy6K4TidwGrGCOfS1PYmIERRGonmTLqq9+KKRBLcJHtXG9SR4gtHlXKAn4oxdFXdIFJCuU
RJWgeSOKm55ub7llzL7YrdvHgX+Beuf+QnV5KCBc+eN4CL5wieUKD1y/ap1ogRYddyPDdHOzc/pf
op3oifTsZuNmKtvChC7uOrq7pk0fsDCG8XKHSv3Vn5Zhq4SSjEThH2R0eLwyfp5GEC+DkyF36A+C
eLPaC2JPbjF2hKLWD4moUZPunfRWF8GNIStfQSkdu8vvhjH83zav4BSaNdczN/NUSIUW4EB/ljgt
DnmkTMwR+hku68Zv1jNMiFtVFi14LYqFcfjsVIDJbw4ol/peKkZtgJhxOHotcmQY2gVEWHIuxqqu
CEsucZ4/4zYhujIEWcB/1x/7rdWPU43c/Exp11tmY8rbwv+ACdHhVbRIDg5sSmWjgX9cO+ISxM+L
NG72jUEXQvQpNdJ8e69k+2+qKt5pzs8Irfo2M1xspxH8Z0owhfGnw0yA+pp6+/IwWqYJcyuTmaFw
wsK22nLzzE1qBtgBOMDv66M7GVqwLT47x2P1pnomxK9LE+v2CQObV2/MMw1AfGz40/XnynFJI4pF
2uy6hAig+4K6L7T+pAgmFrrmRpEt6zEhF1pb1JZNy1DeFDUShv559xRkVff7xMcgpEMSUlP+coFX
ta47SAahmPKYwgyuU+cJt+Rhzj8g4XJCF+CWEEH93VNpzLhdSAu/oSKljIr+ENIjmYkW4hWoh7oQ
qngbYWEXwjQ3pSxgKOuWjgZR7gBucdYXFAThJx8G/VA0J4ti7aeg+LVlDfh08fdXuvln0IJZRN0z
9H8ZJPjVMrcM4gAFzFC+TnO4XOoYyPy8ysFx0fgUyrqAvfDCk+zTphh8BgN5Li3HC1kBurgGGW/d
Qo91CBDxFTkSRyxP2aVyeaAj3q6TFzZ+T6My0QXasTic7GAuT5qWPUm+v5H+6mNqnMEJ/eA11hSQ
3rYu8wLuMD5tR6Zs7Pop9vDi6hsxK6/qIk1U9EZ8m6FdeoV9lH+2znG4OzoIfvx5DbriqJ8JgJyh
mxP/2gWkgr9IqAX4ndHVQtCdRGk6grMkE6T5VSz8Ja4zbU5IbwbYOArCJPVX/O8KRxhzUIpVBQxC
NkKu2cTKcqngM1EWzrQzrwnQVwHY8Ri08c8BMNVKV8BpuuMCC4d6+z4XwPloaSW9ktIClU1YLZet
spk0f8mNQK/5Ncg2Yq1pnwz+WxhXhBFOqme74YsjGHwl1KZ5cyoKg4pLQ1K3PZhXWq41I3HUF3Gm
9z5I97BFPmyEYsKE82BHI0VSafxSctHYHjBAv4L4zJ2azPeLdKeBy1PbR9qAb7iLUaSd5I4+BX3I
eSf75z3JvOgjzKI+CvrxNsUX14Qx48URouz7+lDFqdHhfZ9upbYvKZ0LMJBA+wWlyvilw3xBX9Wb
fKkH5Zu8bLy5/wLKM9NKJ1qFjX2c6e8RMDNkc1YM3cASt6KfYan0p6iGu73D3Cs7k6J1xBy3fX7q
xJ1d826eSFPpXEm3j1U6/cL0xgsj3wVPXBH5trrCp52EBoqVSaDEYHo8WnVK0l6kUyVLspcCy4R4
x1AVzMenHzz7VvjZgCKHVqeL3gZIhvoIjxkuXBL3Z4yo5+vDp7x80g5dIunu+bAdEkR76MPnxOQh
2GVWYEk2C8ACv0L9fnMlaR8jbc6Kdwm27Gv4PEo7p1joCg6eHk/IEPXxcRnP20Lzr0aqnJHrJzDG
L1awq1NGPV57Vvq1PJ+dgUvYay2Nd98d5jMAMgxy3bHP2pqH85PhpXD+MhaE+SoAcLdd59dxsAXw
TGyZqgFy+t/sfa3VW7eqH9bvEqXLh+Wwcrh3j9gpwr17Nq+RFL1ifU/4SpY/V7vV3pF3XKTRETIO
h6jbOhDnUdfIMMqkddReHOx6hA6xJTVMiKEADrmoYvQ26shD4YYuF0+uTXtsAwpiycPcOxhQdvzj
HSkvbWfyKXVUvfBrPkXuihniLvkiWbaxLYvVnKqrFAprg1wx+MbsAZPdyFO2A0Ehdf07BcUMbmP2
5Ga1NFno7Ak+F33aOTc2JZCyTPfmEhGzYL2RzCCh/9mGBkvCKLDhFjn5NleWzmGAcpLCecJ7VHNz
2e4F2u1lG880CoNL+4E7bSmen9MiaL6T0G3b2pntp5KC3FDMISJPQ3oZhy2sxPh2S9BkKG98wl4V
YCXMG2L/MUj0dEnON3tvAyaQO2A0sb6tIuklsAhLj00hrVggIHkuI277Q4BOd9wzyBtOg4CvFoeV
zNWZcRwjbHGVFFvJ096a3NwcOgGf7hPbvAl/iaaoL58a4HitPI3HuLiYIvTFSmEEt5OnAYhpPXIe
JZfL4t2Dl0hLu2jx02CXf87CutkwrjY2hRj99iE/jBcB4qlhyFAE7xguzsZtj4KzpfvUo8qPZVYj
mGVz1BPxKx4WgsCD64xzmNT4e/tuvW1qXDvqjPSEaxh/MBVCkVdrTf6jbOR2OMvJnquwYdYBP598
3xb1e1PZlGD6uAbQUInkzv8oP9fYdPqHkSOpdMESdNsHq8kD2GhnYEgJ0SsKbQbv5SEtDchmGYTn
V3Iu2NuERuI2jvJkKHbArN9CmRD1MjOPafofSklstdB5Qm1sbhV1FiFMnHyUQESGY2RseU7lbts9
1URyhgtBOUNOrHgZ1Lx3YZ9Kw9+tYWPovg3RoIVd+jFSerEGNwBsxqkHVU1/oBc9V1/wGdqeXmde
LZPcsTzCm48fBqKA8o6GW+5R4mb/YYf0InJD6PLCsP4q6orykrfsaCJkNXPDKB4jhYncT//z7Q3v
IPyPNthhjuffdnjStrtvBny7072vBCR2vnTcJgPnz2wNKTWFUdLCFsjCQ9xDh1JESZAE+VyG525t
AkX4TJ4ZR0fD1u9KY/4xvBoNfHLia0OSTsA/kWFIaW57twxn66POFeYgnlzjIdjGpBjoC/eL/7YR
zDCQkTxEkk86Q2ujrbdVlNhsFSgjXlW1xjDFxhtkLQyZtHGVQNEPXhJfjQD1/cNJJBlVr10SvVOy
CIbhVxP4kQAyzlh5KyoqH9ahOeuInuPWROx65gu9DMNHMMVLFpibmZ2zvpwCiFlOKxl/kPur4NKm
ybJPLtG7QSubN+Hi7fqSfKxbBJpyxOzDmeth1CUgoGeu8Y6d+IoywYQL9xUoATEbxsxxt5XmzRJJ
xDyM7sp59j8fycyDaOTzbdq8jmOehg5Q6tKCpj+AmfRaLFmauCQq55M3c9AZLDiv8BrF80axjU+x
8J4y7BoQEqWZ6wAWXBsATtT0Nfe30ODcBGSfXFMKlVz+ZLqQJNtwRkIcqLmEnsGfUGKSbglXV3Xl
liEWE4qmAl/5s7gKweql2dXTKErVeWqpR0i0XHbHSqMmLmhALB/JUvMTKvN4DHWQ/Q/hVGRytYQq
BKOCaEd+5SLcDNwloRtyPMy57ysTGX7ocBshyLB9j20etu4aUoe9eyjPvHC7vNbSLUdJEBhwJPCA
cFN0Rwtxm0lRUZqjPIxBCLLFt+OLgPOLvDmus96mAfob0zoJO7pBNLYK96E3q0EcB7TapchwkA+z
xqbpFqFHnl0TP1Kgvv7/R9nSuXKGor0l6AnXiBO2nEODKcVmQ+d+WPF/o5ekvRcKWGKbaJ8Az+AX
iEbLrL82Ss8s9L6QfdBa2DfAn6n6Nl4GEwByQA3CQjNUusGT2zvqYSqMQsLZHggo55V8danmd2N7
RFVBCuIt5a+f/2ldFtcA7KonLC95IL9MeUWqQQTNTy/6yVhKNSexzaQAD7rOVn0j9XCg2D41CM9y
7c2TIG6RdoiKuwTcCXVieSNrUhj4doKuqTtIRHko8iA3aGEQYX6AoiaaZp4ol6NXpp0++WjA1dF7
Tp/eU4F0TbNicF6IwJpbDb5VosK8stZgWOvaB1UHUiS1rZs1TGlg16uDLWudDLVM5oOJr1eiXwAT
CBDP4wZtZCq+YKtvh6vgN5qQ9I99c8HERCnMwwsVLqNDPovFzJl61Ivk5u7gMlvjhkpKsiOBA2jS
1pRp8j7QuMB/8r6kjDWM8TA+XezX+5wfhuAFKtB3tltCaW2pGffJqtZYsazacAV8RyPtwuUOjQt1
w3lF8uMPMWH2Vtt+/Vldek7IgdlnE/qllZuCl365fLPbNE2WLKHd3mWVFPaSYZ/KppZTGnyujEX/
gGp9f95CGe2FYxFtzySYe/khasLAxDjbd46IVz8H9G14T8YOm63L/bXsBqBo/JzkvgTjmZuxFXuX
av06hweINpzLdpaBbEwmCLaepj6iu72qvLjSfym2GsvNsXSKotVy08NZy7PDtNMtv11IAly6uE77
ArvgayDSVPGBvNk98svgUHxCosSLw6othmY1lR6ko6BzUbk8iKw8pjE9B+San/UUSfSZZhtCtJ4D
fESu+ye/tJ7GUYYsL1yn16uYkhHK6fmLdlSv6KZhcCZhUqz+liK1HHtF3NsW5hPKGgJavhpeHnie
nLh+6BuM9H5PWCQ6zy5S87CW9FCRFspf2cHidFWVVpfDPDDRQ6a9CQLXgcpTyuEDo6t+2LyU2KUc
JULiDT8vIy9DmR92MWVNJ59eAvJVO5DtULyD7LIl13xIDHW/+73qQ9v9owIYlnfQirICwPIdR8kf
U2XVFGAhMNBs+5pbpc9PZbBhcP88h/YT0mE7aq889mfV5Ccn37AO4CrW6fCjirvOcfWRakKsZIbA
XOSyRrQeqhaLSgAfKlMaAu3C5dswOpMGJzfHLT2BOnIqKfEMREwiDlZkYY5idDV0G7pW2AzZXbEE
9PprUsVywGRyV6jVi6sIHuCNaeOf8PiEyMxFDD3OiJG13lFkjpDMUznvlGZRGqbXqw28d91MzKY3
87Bl1W8Acbm/28og2ewBx6LdBly6h8KFBD+AlBw246s0i1+0zs4wkij6jmy/caMIDjAQzaUo7viV
BHRf+7bMk/Ge6uO2vhoIH2dvx3MyCt2AFAIBVvlZJel1gWTgO3zP1t7yZh78Gg3QrBcCCiL7jr7H
Dbj+l5+uUKetnGDXZQX6UWGYrr5yx0nXJiXLoF1BLiF29hGXIf5XEDukg1POde6n8OOsw+x9MhHC
NQtskk5fCWX87HK/7div08hwiJ+r3pbYQ0qst+fn9LpUhG/yx4xpW3Ge8Yc6I0nxGSZ6Sss72PlR
+gcQTiXxM02MzO2dSNmnzpcf5SkQKeU3SjFayQFF0h45MYUdcz+dvCTFhqrYpcBNyfCY6KGpq+XJ
bdubhxBqZQIK3HCj8sR0isoEUag3a3Fw5RK4i3G9IOZbwQlFt/fu1gdQG4iGyGfiR1i1RJoPcSg7
Mu4HlWuUMMHR+BebnLc8XK3iuZ+DJU4sXchY+EkgCCimU1JlvaFFJMmnJoiui7hNG76F2etBpbbv
UhbJ7aDuhFXQQ20VYA8Fr5PC62Oz3IGpNVIPAgWGuF9NVQACAZDWYmVdh015pB9Q8/icU5qrZnD9
281PeSx5P7LHNfhV+VUbQw+qTaOCe3+T0rd1ZNT/auNN64xKOmxO1nIeMyOeW+uE5Oampz5HwGYS
P34B2uL0vah1hIYaFFpeLwAN1h1/UcTEoIlfci77S5GgCtGh1eHUt9Ixmz+Nuc5wi+x0+B3SRsoz
ZpEIKOo+19OyFtAr3Z3+fld6KqaPlQ0PIK6caNlwXEhWFplAriKVSstIFM+WyDzgvI6PtSvwPxjc
+IbMe695ML3mKmtZ1gTCYgl2i7LIOwZN5wTm6zRPZWmz+/znhhKV/R9inS7KZjhrVhBj+GqEM5dz
ZWEOFOvAArAOKoeyFfaVqP8oJb0cnO6AbDGkSrzLkQpGVyt3mwREGD/CrtbjyhqdsmYuvQ/CdrAv
4hWKbhh+QFfpSbHjZetHgXpLp4oeCc7E/LJzymC6OojNB7/E0ByFpaim2o/K32SrMIav1sDkwmf+
6Og7UOBmDZSYV8TkAeV+zVjeK15xDmeQBGp4ROs0SBt7yqBjHmt+1//+xdvdeK74mThIFOTLvolt
+qttxRntolmCkI8q9M1JlcKrUHfBXaVFg+6xbMGOWILyqNsy61LfHa6+5cPJZHyR6ooBFzOOI2AE
ytl7XQ28f6oPpHdNbsBrTemngJP7WAR/JmKgfZd9Thf2d6NqNEcTCquIfQlsgI66Exc+AWTXCnwt
EX6/aff/yXgkBUjve4iYv4+HOq2NJ5PntWe1NdrsnfqfG2m7z0W6tkpZdDWbte51h/RiSSRQPOi7
aLBUUJbMeBy0gklQhB9Dbz9l0ldfn+wmKgjkk8M9PAsK8BYf0yxZGXQvAGAKmigPA0zIpFQ9bgah
m7azLiHdVwWfR6NBaujS1tw/eRX3P6kR51V65i6uSKbkqJ3GitSXKEOasKxVludrelRlNZ6JAbJh
Fr9/FBrk5BFZVb6NNoJtleiP2uv1w1nmxwx1JNdNG5jTlDdN5ufS3F51SwcWQ9tSkcNyJmpQub06
i/j2uugGZrDBJnDMpycbXfMmsEUTn5sE3o8fRJowCaraXwaEpI3pdPrvQ7EnqxoOOpmRhkmBr4+5
R3049vK2u9Q/wZPdscZqpDrSBtk5xAORmeHOR5t51qiNaYt8Y/X75YlDQgKkAmEd2Y+K5vYO5qGf
Zyb4V0GH2gvpluW6GJyAraOzJcBt+lXLDzeGzSHcnYxCoNVYugXWM9pp+9L14JLtqM/eBBRbdc5P
JIv0D2fvpx/J+mQg+T+f0uBVtBTn8fNRiP+R7aOZ3KUod5n7wS1kdbYdUUx9630XZGIE6oPWHrWV
+oNK4N4cZAp/Pirgx1dB8Gh2ofIR+1w7X7ckvUsLldIivzSnjrUrBPLxG4o18poORXs3WCun+owt
jPS6WjAYRRRs7EK99Ef+wyRuhAq0IzDN2g2wH+wvL9GTIrHK8JNUINQ3fxaQlJlAycBYZOPHQ/z9
lhbzfXqzNG6prWd3LAw9NCAg0nY5PDj0ZmAjvsM4mAxA3x/pD2PfiMYNE2CYmeBpbbjWWdIneyzU
hTtQz5MN/+SXhXqGCM7VEBQ5xqtEw9r7kVRCcPYzC5CBNIcOSjE7pBrul1Tbaj1tS0p2T6WQqzpL
ZO9O+2gXvD38lWk2DS4WnC3k3jdy3X8Wfhes1Z0TlQYdDhDBZ1LVJZOqqFtjEYE8fcatSimWPKQR
k6Gb0STqULOc9UuAVkRY0VFgkgCOa/4JMpHGJT6FuTlj+H4KblQhtrUBi0B8OuTDs1Ih5QBoNPT2
Q6EAYroNy6i07I+eqRLSf5jMp9eVsOStIGBLnIDuWsyTAI854iut0glbzsq1E6mqGSewrxjSURs/
MsDDZkIyJWvu3PEHm9qn2YZkHehi80XdIvXQcyZM2oaNJva12tVd5+dHD1w2YVBKmHBvfmNdWTpf
548kuKsjauIKoEYs4bCFXyEdfD1jpGnJun3ZmmeQVx+4o3FeELP4Sxpcp+UtNxWsvhs69gxQA+nU
AMv9u5VwXIZCGY9PU6QMCAGbUonzbg+oF07qC+x+83UgHgaa6SUauD0qZa4qpvpv/Wy11FvY6+OO
aOmsI0qxQh25I0JPeDf0IZv/3p41ZN+QN3XQOX/B+Q2kj8wihyIHHbvg61rvmN0b1HY+Uwl5Lz8a
KarHA8Z2gvCaZplSpI6iTOBnE24JO5tdaftPlVw/o8+AW2Go+s9x5gmL7MatcAw03U5hsA68Jyy4
Yq+kUufB7TPtx0OZyUVnjm1GehDZtJHPfNP0ugqpGgVy/61uTAhsprRyurNJK/RE6u5xjwEDnNw+
RR8RIL35KkUGkYGpZytSTc18nNiFYHdfRan4xQcIkl/X+cwJp1ZQPRupZhpE0LXcyH9UVt9h0y8Y
2MBW0TwzmsWujsUMSycaAXHhM84kQPMLToOYagMp3wkAjhig/cLYpQ6OgAdPJ3nF2xxGyEiEumFP
bYreH+2GTo8/t+ijzDDXU13C+MF2TbNiy2coCCffTUERPO1ePOOaQYkUwEcH7V4/G0vWHbfiLmQB
ZK9dqRMBMb46GEg9sylx4g+Iy410naz0DTasy86vEY2e0zyccet+BCauB29CtSzLsbFFQSzVgdAv
qHF/UlL2Z9BgS7QvX7H2exG7w11AvSVSijt0vr/K42EsGBlkdgFq7NCYIJCJ0jK4gIq5r1Zw+qun
KGhHzvpkKeze48xQAtc0qMH5UePRoG7OSyRW4rF+6WYYztqQGWw7eIFkYOWAj+WMgWpsp++2JXXp
GyeIqCyvmOFGnVmUSzXPPemaihCgc4sGQS1O9vPKRMdxm4z5kuJ+SSj4c4w2zdepuQbRTDCDRelu
efDFw5hwrYLAvjNoEvUGvzy9v9hBuORG4q7DMoWQlVdRCnAispXEYzEGQvoKgkDhpbjQFQxYFYIv
GtFUasnNCNVaFaLTXgx8sqst05z1QoRPX3r6lNsRvksNjLOIB7styQvtF2is1xIwjd/Sq23S8meU
VWZUSCpbHG7jtxjIfBWgFsuOUNwP7k8SwUHwDHx4vtCIMitQp1tJena5zKQtES1XNGDEbfrQmLC0
AYgmIJKFoRURCihjY6D4QZJoa2IkmK/dG7oPL+0d/qcf10rmHMJks/rodgWqjvYiDsfrTO3ejXkm
QA8h9OpzJqt8Y+IlGEuHces5+buGLodZCTguhKQzgLWf4LDXtsLrVRmKUj4t4G3mVGobG/0Npen1
I7VoBtDvgDdCMUF428UOQNhKhajTDv9TuMls4z3kKFlXYPfU87xKzj+rv+vYlZl9aKTuXXFj0L/h
ecua8jRHdriwDrzqUGCeEFtO9PKEHPY7La//a4hHyT3O1XcthZX4UpQ8bFPIHh4xweJqI9oqQA/4
fUOrGl0dgUEPdELs3n4GV0ASGn1AkGu90Ur5M3aVbgou/+gi3vrHB5A1sc2bm3n/dJgYKyCaIQPp
zF1YEfPgkOzCTfw/HkAcvf7aegI0dMA9YWmIoBlO5F2bDtOWm/Yxme6kn1ibQuHHkWc3viCTQqVE
LxivIAPWgFQSw57xbmngchIQiqG9dl9i2yCyrrq6TsOHCZ4GY3/k9WBP8kMKdvX+CErbcjvS3hdq
V7s94yx/V4Hy7+cL2RtS5faWwAox9Y1rStATlB6a8viS1Pd6iMaskuybjh01LUMWVgOttXwNZZgu
eKnFK5YgH68pS0dMe65qKOY+Zq53EiISBreSR9RyyEdENX1hDUeDQA8rbcPfLHMMq76LrVsxozC7
WVUMQq2DQ2fgaWthTwTGjbGWr1ETL4Flerupq/Cv0l0nHxexoEI2AsB9f2mTjlr8n5rGD82nK24M
aiuPzJd36314KVMghdhkUj13ulHzQsYi6A1Kcj6WCLTm9H3f1fekDXdrUgehApPvTjeJkokXVi68
WpCA9I6g0yBFGGerP5tztmjRqMWPZ3iXvrNiIYTEz+1+ktZ8r3yY1sn4henZ3Ap8/s0N4tVLKq8s
wUxzqsP8SFNarQFT0MX5qf3bWCHrPBag3ax5iSU6FwglOUfDJ9IzAkPgm+c5WQxak3bkN2JspL8S
tIdAaL5KxH3ljISNxP2aQQwcIgXzZIxyjOYTmRA0oZEO+dlvEblQ59UihM2qLpe0UAj4pPVbDzUb
zNdn0eCETTQXVaswbfHxoCQXIgYte2ClA/pHDW2zky77Ie6K/Xwm+yNfNPky9lLUtDuRgf0y/+KY
7gRKwEtof2Z824yZH3dFNF7+0qBV5OTS7P4TOH+SnJe1ZCTeTNmS5ImHi+IGpLRuqQbOWQEapHh1
4WvcUuimyRLReFNsT9ZAj0FuroLANgP+nSCOoHpArJ0aUhDCIiv4HVjNRIpzbmQ+RLQaqUOhB20X
Mk8G+rcXCGXS531Lvp1ZanJhnhlIw7EgnP+8ZGTT1rz3DaWwlem7dUaDf0CE+tjJ3tSH2rzqMnT7
yFbTQGOJ+18w0oOg0LenNtkiqz3nQSnzxj499g5W9ilqMqTaBYRUPpNMHHqPJNg/g9UaJPgE+trB
pry9gPJ6W7ZJzmvSWQTKh7TTCOaHS+ZzV2OeiWsoKLcQvifhqx0gg02ZX0GaHiZcVNJqI0mRZN/q
mauVE4Saxw0wUj8iatdXvCrUF2pUUcPy98j5XBkvdIT6naeuw2tOb6kpvL8lVq4o3OVNnn/6yWs0
73yuh1Tuer2NakQfD/dd3tAmxYHd0eeEAjW5DoBgQDZ2YBz721ZDaaG7Ii5Tb92YLKg6U46wgYm0
Pnad9BXVPdBXAFFh6UtXuSCWeE3ZfjoV+5A214Jw+wO4NKhwfMpeyqp+FnzfkhuVQFOVxaCPMA56
VoDhj+3sSQwCFmToqJ3J60DZ8iwAGPr5P5izlfNjsa3IlAqnU+KMU7FcLuAlWQLgy/7gi5fm+CpL
QUU05BLX339I/fSr2nzDeU96Od+FpjGCcmhggU4Pxpv+vMUpbuDVdxSKxI4mKj9v1UbsvFFoZDah
E+ont0gpg9vPAe5sraiDXR7DMDNQB9lMmaoaAwBGbjtgwP/xgY+9qmS56Fk/v2DJRD1VfvtTWiDR
v3IFtdSeo1KR4lxeqXyKjXqQ+oCFZNJe9EIjqUVLmTBPKj8sPaxWRr30N5QhnXOT+khKK0Q3VeLb
EoGnPKRAjbh8NjUaNR4Im72l3bRJSLmtCwiShg4ddPUSEY2r7s/X3AleYWaDyiTEQ5H1wi747zwD
SYKjZOZtuIs/EJ10fb2B3i76B/GPK7BWIPEPDq2SDlUZNayuBEYY72FnWTg56iBcTE4SaYoN+QiX
iTqG4L/dM0MnogOTIvBaj/gXl7G4I5hqbcxY+ostJ09kGbnReVHb5dMMIal3K9B4WQqhbTEtuU5Q
r8RbUtX4JkCXfBzeHVVX8e1QlpdcI6AP7sqIUZ0DSmzzEgHqOm9dsZZGzZRIF8EniKm0t83Y+RPy
xEauxssKyC+qZmnmUQle0lOYLheMNOXcci/OWcxUKR6RdVd1NMX9tZf5GryH2qgCBUzvarpRwkaS
rmheRCj6H6RhZ96rI5hhY+wboxOzzYxU7gGuXgXWvsCPTy/k6lcbGuIdIXzoI3O++LX81RnC06U2
m9o/c4aqZpjCkfEeLel2kASOQlCoEN2hBaRmyVK7TEUWrs2CHvZHjeMVthKl28GROOSMczHFwL+T
4MqIsQKsHmqystoYyTDNQDf7LqG2lPmJgvHvAQyyC8xvt4AfLU/xQjKD8cD58VoXFRyEUpJQXnZn
scTAhSF+5TOVY1MK382PndK+Qin1t72JqxO/PUWJIXn6c6owtBLtNBrc8HBFnk0awtQFKo20boRA
+c9lhMPzNxx3ORRBjhGtAdr2b9tkqHRjO7WItPY5quRQWaU9BnEU44BniQ1fNebN2Um2gKwflY0d
3VlunBoMof9O9UiUbv+l0m4MUxJNj29oXkl/MgLxEqh7yH1jiATNn5iXkqc3vwjOoQW1pwZF445l
fnZeMrnldUVe/o/f+VA1URKpjDtow9Vc0j/mkHbr+6s9VHyDOopNpudK4e+ZrnHgBzetL0dhNFli
h+LCSP9H+uqmd6mGb1Tv8jIoAKmbcdn2RQIeIDae25kwQB+Uo4Z5MrgAERKI5V6PT/fHzds9JUv/
WjHjxM70R9nV3KSUiIvbSlExeBWWonE4CekamHrFNqX8PSva2hQAtaXd2tMBwOcPU23372Pd5a+Z
YImTt/gsIbQiMNL6Dhz4uDU5kv+Vuz04n2nBeeC8dH+0c+I3XKi+LBFSniNtdL1y0l60vgLRn+U5
0ke7LUWP/PYXeO7gfB10IDWAj27amAx/K2XkdmaxoR4Zu1Wkc91e7iIj1+trB6llb+1om2Uuz3Qm
NtSP4nTYsNh7l4sV2LnXBlAHiILSvucL1JDS8btdb8kfyUda/vfFUTlXcTVcbRNuTRXkuoQBZU40
BfOPrxJ+CIK0vQ2C+zUeuvR9t0uDDMEe+9VsX8zBkuNozBYhR0uqLkMbpfE284wS/ad6WxX/vXq5
3LbNYmwykEDAGsE4hrNOYf2ntmYdyykcT5sYbJy7fUKaFuVW6ZUxXXbo+lSskLTpirizV7BOcSsF
jYzyTSasADDvIula+HaoQCYY25LGPbHfLvWeSMYHLH3WORwnfR+cWwkfb0GbiU7bOAlI1Jve1PyC
ZSbVDxdNIr+uxVU++EFFIwCT+7UuK53P8TTYG4LIDfu8UZLykKOw/AZQhOcurg09ld3gAXjVy0It
3joTiDZ3N9SzyY6+kNOAFUp6bVpjuVs8qMibpblJUV0UrADyPXTQrTQKe/ORikKcCvyaNCjhrToE
ccaDqcu5RWUnVJSCtm/BC90O39DfojEdGE0B3z1IVwIqa1buTdHil5X0BKcuzvkmib7qtvs3aG+s
oklWXoWRHQqDfEdsF8vxEXeHGE9P6CNAIoj5cCsNkKXbZTw9ppfeGvRMXkpJWqswGTZO8V6293j4
hI/PHyAEXxpFcf044458A03OuzbAeyzdjw95GGLZ4+f1/tjqUDxj/Av4Ty60PKiQ3cDM7jB7dYmU
LWZs8UAsxwufCGvvLo2UFYu+sT9Xr2n6eR0BdeGmUw48qj8ZrxS/zo5sSovULgMcxIGKmk5WkUbb
EAk0vR76whVn1K5gGe3/FKfPJjMFD+BG19nUZ1Q11mCa//JMbYHPqGCX+OYlQ3MP1AY3s+8JaUqW
HHd+g8qCMhP8ZUb1el9NgeT/jY/L8tf1ymIWvoG/qC+d2lBo5TDmd7rCBTqzSZFpLuA68pq2bqQu
AyYCqtqImJWq1RlvPCRxalKM/w+7A4cKvWdkLsu+7uAUpbZCwB8F8wpFfqhi/W7id4ch8ntrErxh
3TCISzzwMV8IG19KHrNedbFbRsjRVylqaZ9MTPYGbFMxx07s3EiZHpruse8BKXFTOQt4LSLzNnPH
1D5CAJYyk6gMbq4llfIixrUf6doZvuSy9gqM42axDz5sg/LSFVfE5fE7qd521BQhqkerkLHGqq/z
jR3G7DduqSTcOIyAWRfHj25hdcCU7kETpPKLr7iUxqHkfQZ2XiNn+Iy9VjK9LWHXcFY0fbr09+ZE
IIqg8sufjV5APNS3AN04h3cLTI4I3NYMivI6OLDtNsGUN26oIvuE8fz6shiqrJW7vkG+vw+93Mkm
U/aVIowb2drpv6E+llEfbTMNavVHgdj+xTa0HOtTd7CtxDjq1sZi4i6JmY1oovdj+DF3LOgdDr9P
Q2BiPYG+KO8b3DXHnkJ775K53SXQLcXh0pDO92R0YSbDYsPHuHcpOgfj7RlcljgmRaQ8hXFRGQG7
QUdZxMqWswjCxLVFwk8VhtR/OrhNAM3scI36jTNmdIpJdTd1PQnYkikBYet6+HDpRdV8YWy2x0ES
TwFAFyos6vLVhqltaixFYOzVPIWJooo4X76SmDQdhjPUaKoLrHUSoafGXMPn0cqWCMR/gcA9ydjx
p1JMMaJV8fRUQABfb0nUFo9ngyMwy0GUmnegRlojfbs5yy8kaqtlB79dYVy9pG2UIrvbV6Faom39
GhHVjS0LRWUI6zf01MJkKKu1rqOqJZ1lVQgOcMmouxzI9+ZsaEDsACDVUrIIO7L4WTn8m77UalRa
f5N+ADZZu5R0DGlAeoyf2+gTToSaomaKOFnwMamSl7VOfzyMgUsgEcK3bvDDWnpwDtTPcu9ii21I
xVkQLujKmDSiZ6ztXydShbTBs580mLhfLWXWBB2cd+kfjENO4MClNBUkuNhnNFIFDZTMIfPnESXn
jmj1oTrM06s7aJBQptyBKxfnovNbfGGnBKaSldGkvivFdskOKeYj3uLC0NwbtzTdAjHkSAAZE75E
itMgZUzaQMCsVu2iycc7xegVPCSWxFfTMfchHjFWesvO6ifb/5z6D+DrYWZIVRzbbURIEBD2IZul
cI1YIeMEKUuTsb8aQYELNfA8rUYbKcPTUM0LLFfwfL3sQCoeh52q/Dpii9U0vdHNjW7GuRHt5Ghm
jM8oEw+K/43ewjQfVKc6FQQtutujhi50FdQ0ot6/Av94/30dCM5ljXg2uawPOMoulZ12M6Fqqi96
MQYJSb9qxzWB0ecEdrmx/iPE2kUBD+GhxLinUE1xqKMPz7/chUpEeekjgbIPG5FY1XvlyLk3KJwy
3TUE3nCKad1SK0Z/7nqoT8SvvcIDiuZEY6X5MlI9TOcqEVOIjCqb9xdy8bqE7JoqZ74yJsCOD3dg
sNtqUiNWW5LXcrALy7URjyNSiGpDBegn3mnPgBdAIuUtfQ2Wp0v3/S1vuOqzaDjtqmwE4O/TFaG2
jr2Dyp0k1e3H333k5XyWMi8PRpTbttj8ilkKlNlx51x4TU59f/2YMougnfZDEoUjuGnz5Yz4zx0y
QzaoiNQQWUH5oQidgAagZ82dEYx/NtGwygyazXZvzabyWiDjDEJLkSG27tLCjxBtNYVAJPp8Pu8p
4vSItmcct7NNJVsssezgFiarImhv5LYlRpeo0oC5EzXcQ6l/AoqzpdsdVyNc+TZqo8q19+/WWgtt
+29+HdaKoc8A3lIDxxynoW5A75zWByIvKylrSDzIsSNR7vGJSx0Cis6ZhlWfv119mMN8AkwIlum4
pyV+1jl9eDurr6D3ysdhd9wzPbchkiAST3EYICR8DZtAuHZqk5Wxp3dNW+24y25LZwDXDYrwNvi1
yCAM1rlBOi+SV5Oo9+Q8aqU8SiklLehIRYaGajTebBndgz25HUECL5Nesbs23+ZvZNjd+Eh2NXqK
GoUJ8P2rIZF7fwkiA1bEFbXctrEHb3dA8dhoD6qHWI3vpsy2GN0YDGLxXDXwVudHmXm0WZ5WOp1p
Jj/uz7UxT0uzjldQIch+8aedWydS+SxO1bWta9slkTDGCktJcAckc12yH7rrk86R5/pZU4b1lEgk
jPkegoAtac2l8PDd1QuUz2Ux/dIpaKB8xeT+tsBIkFoyyAjyKrpjfFbZUBqtVL1QW718HRLnwEW5
Prg/d5X81OE4OW1VCklJ5b+5fYuS2lQPO8Z9govrTMdJVpM8CmW4eTg+R9kVAFpDFn1Dr27bOxFh
u/EP8jPY7BFOEo6MnxQp91TH5udJ5SwkqVCRfz8Sg4fnEQi/Vl/2aFmIS1LWN8yb7FTbVsVSTQYv
5YpI6iuy/AJdZOgRIrBe7EpHtA2pG7uYal3GETwQtvzGS4/EyOzItVZqIiFwCbWkkwvHzPcuuHXT
s9HQgaIB5/98kBOYlQUf6lLXU6D6cbbDVjTmP12+em+aZcK1MXh5+4JBE5TAQr9M/JytzCTHrCj9
Q4VafcF+waYdvu4ZeoVPqrRzRSP595ZnIADgFCVfJTyNsmI8L/HcW3Dt3qkS28pBXXyOCUIG1uGK
XHSSxBBz0K3f5CnKVDVJ4KQoUH9Qs5B0+AVjTM0EdZ2PlUQCKMgA6DiJBAD6sPv9cInWN/+DnpDE
wNH1/jVAbX6+mmETzFRxba5xF3Mt2aNYSn+q6YhQ6xVRaWATxx9w4jGXgJx26BJyqQTJnkqQduwk
o4DMBZHZgRGxsd5VxN4FFZ1H6bwK5SfwRDBAFZo3mNDS4Lukd4Nknxur2nxiUukODZAvcgDgBr/L
2pfbGODOYqQAq0jmXsZDKIcB/cV+o7N0vGPHh2rs627e4wKhXS1B3kcr+OldD5OwKHc3SBVj/cD/
I3K5ozMxMPX5G9eZOaMVLrya8ENWirbBAxzkxk35wgeAEHcdUIefXrrNtWxDDGEkC3jRDwgsx3U6
dsOdGDeltw9mqIIjYuYuvyqsFD49voqh2+e7GzHaBpATT+7D97HiwVwgaP4jCkh6V9hrWdi1y9u0
WS9rsrtj/J58E1j5vBvnyaBK6EaG5rN9pd5C1iIV0TqcHofdeMe+1d2Gul56kAKjNDSrnynsw/IA
58g+uYRbqyLZHpfJglaSnLDplxZdTn7ex28EoL68TVsHSQJ5/RKC8pI6njX65SwE0CExd9nvlcw2
jKcyo6A3TrURnKDAmyZGzLZe3Pi8IHUJizRdkTE+DACOC8vX2JN4iF3583EdQN/nSN9QuT6cnaf4
7UP4Uih5+HvmWPtrIuR33Mc/Rm32coYCTPzvZHZ2s1qsCmctCkd6zxMlGVMjW9h0/Yg0tSJYTnc9
6RZqB2A+xO7slKe1JEHR3Xap5L/blHN5UuMScN9d4C9zkke0mBjWaEEpQF9XRPQ+Ijc9ZTvmYj6F
6sEA6yR38sS7Q73OZG2uCb51NoZ8/pv0ynGEHdOg+18txonlRqhdwZbXfqRraelvU16E9iLYUBys
NSXAjocR3ev2gG7eU+a/264gM8+OebeWUI07Vjg07WNpi5tDlw6ElT/MfRPV6aBTPtrHX/DRKq4Y
pXjTi9h4a3/hD2FbfzsP2POwxhmXOlbPbN8hiD+WlH0UpMK02FtMvfw8dvceTT5pcCTpzOls5vIP
NOXkjARbPpVdX1W9mGWuTVWx+eC6sZofoTHvVoq1xy99G9GKvbaXPb53T5ge8YMFcMg0S8LkYLXq
c0HPy2nFaeGEat6rGsaXgL3YBSUgERq2ORyhUYKr6fR2g6rp4w82a8sIz+cCfTIniciL60QvOur8
YuoDq20ZxaUIuPRYj45GX+E2PqpdNf80jTu/mEEB8Ck3wvea3iyZC7836LPjN4Ovh+MyPFGX6zNJ
88Qk0LrYUwCuzF0PA8EbGvfKK0tWW/ogd+ZqB+B/M3Z59xo8lv2xuA83rrSJSrW8RW8TcjafeuTX
AZOkc0VkORRctgoexNkP3VIBsVl6H8MlDUoUX708f8GxfZL65AdgcDtl47UPOl9Eli9mVTTlX+me
iWT130E6kKtY5r9HxlOudobisHqZBhFQjkC6kio0PLCQHAEIClUUW410jGi4olF0rUy4me7Ka79h
8pfVTRfBFQXulnKgavKWldjyLIzwM9A9LUDC6zxqXkWvZIfhUlfu3sxrdx9OG7nevYpsVpcJjWhM
pqyoLa4tvnsa8dHGanKVvJHMG0mu+wMbzhcbClDuZEY4ccHXaymZS0ogLsUYN7Iwvbv1yvgWhSf8
+/WH4She4bzEdHsYLLUiVJGLUVj4tA+KsSb5mucmk2UBuGZWRCnPemblbAvvNGL6xpSyZhby/mCF
kU2b4JNDNRXI4ihyj/cTyALQgG1sNLrwsXRFxtcZZe+QaeYX07CWE3CPIwLD23JmDq692IPoSdNm
+B0YvwpcMi5pyz7QlixYTF0Vsa1fjZkUhDQiG7Nmsv20/T++otiYlbGQy6o2acU1eyWAP8ZxCIIA
WFMfjyKGfeoOzTS7egcnnzOv6oRPr7tyhd9P/mhAWj0v+eNkZh/2R0tALqr0QF7zJQVzmdO3G0SK
XPYyKj4E8DHFcXLdQmoIB1YUHns7NBIHTy1V6ILd6DCccOL5ZeKxeqQF79ZBzIOEGriUQYo3kY7a
O98sAjWXKZ1XUFN+c6VCrIrJV1bL70aClMQo4ar8exC2sTcTf4NSfYwujWMwG9PSyCIhtzSqehrv
woSgyY9UP9BXo3VEcKJR90lKJjoUfO5aKfe/1rLmMvtx0bjqcU5lf0Yo1UaGpabhyxAA+zW7xhIt
Y7OGbTjG38o4zFFe9Ky55sSxXrPFFqhMwey2P8nJV5iSq2/tBxPBl4GBoVW1/Fm9BccPqQv+dkyt
i1tycDC23BBF/zWIR50e0kcaMKrfGf9wuj0Xpnpff6nmWxjIQTW0aaTgRe1MyAnRE1Ae96n5g8kD
DWHbsskdWslOr833/4HahpULRd5UgjEc2plScx1QyL2qze3g4AIV+zPGO3P8bitsnvIZqNE2M3vl
opkCTLeHeaVzTFq0kkmHbk4jn7vwlFFNokp7FAofLgpUrt7MovOGTowfY65QT8ZiU22Qn5N+88W8
x+kUUNThJi8Qf7STyXGQeFJcS2lQfMWjTvX8e2JVGzQsPOJIcGXS50QLeZMPzAqpNQC6no7IZ0n2
AdZxCgW6zuR+1anoG1fKhLncdOlkqL6SJAC51IUZnvbrRGqY5QEKcImyKwG40L5qmtBJQRrD5n4I
Xd8r1XgBnlXj4DyGsuvgT/yvrpdkIDHg2O89QhlRu69gLRFtGEnoelvnzSBZT5t7THQkeFEYcQYp
RJCset65L1Gwoi7QILR+9uVZfgrDVC1WZmGXA0V9Gym1sO7EUOfHrsy6yy9lKpeOEGaq9+h1UA+D
Xo+qvKDa7E0hpI5u8M6GPuwvwmVlg7iIXJvRS4AhymYv6mzPZKCJte/69L146Ij19P+kbHtofswE
YGN+0qpT0LVjOSxlmruaP4W03fCY+MTKLdMM6BduzFoldPbOfigSe1igT9qrCn0SAB5rS8cGFIG6
NEDZwflscmBKlxQFbwgE/0QY5tQMJV0XSk/127BOiQqtCvt9USbmLyTxfonyDCGujKwl3NhbH7f8
elWyL100BN6PCJYdRJvuv0EiTLSQw0AnW4IZZBCqBJKkP4E8BeEL9MT3YJxJQOk2Nh9ShQ2XzL4p
ysM1vZKUeqNvYsv9gpNFhKGuEEaOU45/E4vtikiDvBL6H4uLughBXyOm8iw/dMa/MmyL5+XB1YTD
nHduZUJv898jTO9xZS8oIJ8JcOLXoq4ZZAPHa8oBtOcoaMceHfxSUMLgRUDE/PamtoCBn//6v3OY
hDPbGIy1EODCpefBhlIApYyydEGasqwO2sCmDHJj1EEehKeT7c2tzPoosdzhUR2/qq5rgNn1bLZV
Gs1Et4CJZ3C+nDoe99OfiZECm/+RtoGt+oLiHpNEIoCW5hCf6q1YOmw3tO3Z1F5fr6TkgiI/7VzB
2z3E4MIOvWMf6paF1Cnjja4eMZwKzR+QKU6iGnnMw8R2ybPkst8LeccYMxvKcnVZ1zzpRP3vYQ5M
BOt5nQCCTDJenctn6SCvU4B5ggDAj5uyvNiAroxPEjxAvpoXlXuYbOFe8LKO7FP+kK2I/Gzi6ED0
ytgDFYUSj6XVDkvWCO1XXEXrYO7yqNwwtceT01KZgz6+oZfcSdMpLLlj/bDVlaHVKA/jW05JGEXl
5e0tYOaaYcJTt/h+IFzO9sGlBYFuOQURShQc8iZD8wkZIt02biwA9xwGzBq2rx1MiUd1JU72iIHY
AkJKxlT2gsvidZQM2VKfGmXgJMLVWH/rMsbuGjYrIZHylt5IUlwQTwY+gsbbDbaqX0Nc75sfxW84
X7hWhtg13Vpdzk4SdV4K9hyBg5jNeHVHv6uBe+hTcNQDZ7iSHdlhhhT57MVFFOXsa7sAXkk32yoI
TYF2ndYA20R8RrwIG0xaWrg5RAH+U5HOxMqQyzHvdsfhBNooB5o5e8cPfoBqvC+Q9my4W0QMNOth
Ymokg9feDGrkw5lu7vJQsmrNHSdhfXY+Tktsjnrk1t4+o+OS31NAyYe95EOKuvmarOshn1HFI1GN
QOiwbCchtZHBHe0hrSaNHAOymz2CmokdKl7qavfaSzCMMbYS3+wdXHyK8nCvyXbDGJqp/CLBuNSE
uXCrRybvHHtzcDOsJKPnTEibLiuA3qWMBJQhTQJqCCCrScbvXw+BNQWmFaK1cnl9uFz9rUrATuDr
H7IyVvqSG+fjjh28CuWsMhaQR6p4NQS2hBHZVAl8rAe56uWlkaL2U9Jb31h6+Tr3JkU5DCZHZNvy
avx1WgoFdUjDQJzzf49xaPznVe++1QSjF2UNa77UbTqwOhS87r/qJZRGub4wliSXVK5dhaKTZZWC
ReSl6rEvwaQKpro46IlhY8PvDxV4z15WDnch41lc16aaAFu6YVWkq7vpOhxOTBgW4TXT1jKrGT0N
tjuH8bqAAarhmKMnoHlfBELuBkZ+9lHYBeMkCw/KAZSbmtxAsV6cZJQq84N6OJ3d2ltgS8OnAGnt
KMg/MMe/6rX9GU3s4Tc4dfCj44xHqZB/9pGV0E1TWcVEdznQMfic6Ub+TBrsutcserne/nfBa5Kp
y9EemAFs0qd6BIN7cSBhv3l7nCNIhNamoEaBr2QsdQYDDroj60uXISCH2aqMlJs6mgnnSxc6+q7E
e2d8MUMOlDkjyTBdwC7IfrSsCiMxKVlZmt7iaaAuhp9leswTJ0yVJ1Vs7dkpt5DsJ2gyVD1/65lm
lJMHdQuV769sc6fo8qVEVHGsJO8qvcFnfsEjlsvdC3DJIQc0JsqHDTWQov5zymW7rxQl5RlEGLhy
4Ctba8RyqneObr0pl2S8cvcQEOmUFsJJI8vLsYXA6OjrX1+vRoV8OAPJNU0myYG6cw9UtWk1lDjA
ohHsACGO9Anv+t1xtZBV88V7iCgFBz5dJKkMbTRgXxSlszVMu7a3EHwZjl+mlKVLEjAVLztyFxIk
P2yM1HXI8hGzqulsw/1V+p85TR0v5KstX/suqsI40Ev0gRII+FSIT5RwClGatitxYE8w1uIQtaYh
94eVq3UtLDyjql6eyFo0j60/h56pxuixwc1AL4EoRpi+CD8hkw1/ni56woLIuZx/hlmdvsODm9Us
utwMsu35YjAdSvUZSTf1kqVRbJPaWEqxS3JHINhfLtfLebttGFbC8dablKQmyDQKVJsXYMErfbea
/S/EAKx+5TZyVRc9626hi+h88yCO4XDSpOyvtUOtlNwIOXtHtdvWDOyGXEmBAZpUUr8I2Pvskdq0
2Tau3nq6IgbvFN71t+VoUrY3NKyroFHLmTlNwLchcY/XhABAZH4na6+7CQ4HAyrZnwRiLtxC1G9n
yH02rRQtM3SCACfZluCvFAYNeZaED3Y9PK+p9e9Lbf3d0uAe+0uTPR1uW+cDkos71BbPr7Yl29Wb
9VSV+3RBqrXCag46/KsifBGy2fz6rM7ps9omAv3Gmfgx2DqPmmg9DsEsThlYZ4gu9UMxcH44MqnC
haFjymEMhZb7m+YZuVaSuAmZVjWWIqx32UbEFRSI9Su/ojJFPrWV1aofwkDgnEA1S62yPbs5Zggo
FseCtCHqgaUZOZJaXpNAdJvDv0jBQmfPxbFwrPItbg0ZLa0sXmTP52SRhyxm44kOxl273lIPjMlP
A1Vs4sDv1KcyEnUh7jpYsX8/1Tui86OGuixAozgMVVSiIppbjeTRMWcnest4Xt5ROZozRnv5g5Ma
zblRQNAbC9T5BISF1a4MsMiDhUZkBYLwBrD8yIvluosRkBWDyh6Zp17n2TJh96MKwBQXZXwgjipi
v2+hKgZjcMnHfH6cNLfLI3uF+l11FYasIcujMJg6AirqRiyydS4Qc7LwalR5NMM+HISqYP9uh2ND
+QgfmbHoWlE6l1oat1IXF3jg+h1qltKP1RJVqBnXW+86clQsW5ZTujHkK2tP/hz0pWDxoDx0XxEO
42Tk4l03BK7GacOU1UdJGfHvn4EzIE6zEQAuMvHcVC0y/rSck/vkEX9OA6prL0FXAtbvAzR4W955
XCNMX0ckV9a+JoUjnoRz2JcoNr3Ip8T4ef9AQ3zud+6rW8L5ve3L1SU7Zm7Rn2URjPQk7iOiFt7F
EjQ4TVeLLT0g7WEljw1wiAbkVpFO6Ss1E/Do+6Fg23BYSoi0oa/6ryOYdSxdDZ5sJFOwWss6Z7d/
81E3XMW9A8C7JInkdfpWhLnrVD3x7RP3qK8Wog2s1cpE6IeWZpiCzABz2IlYxqPkE/YKX30qqqUY
g91fp7zBYFIkX5g2DOmfzfBoTtxx0Xks+3u/znNO8DjzxMl9M/wqXPGdcLqyassll26kHQghwbQS
1TwxqEmHEwfsGjQgF6om3niuka2HJofz7ztLTxGwpFGAME3CUpmm4AuMuhrY9JCNg6tvICuRfnAO
OmOVLidtGjByqrh0W5YR+EBfI9M1nMN6OQmgkW8wKlDevlJCLRUDP2pu3hlbgGmUY4LvWvOdQW85
Xx9qgKwwIT8Nx72GQDpBvx7CZFNOalWOSxLozkCa2JhNaXX1FaS5EKX7ymOaSsLLOInKGSDRGv8F
CfGyeQZ/jqvzvqKztc1cRoQ2uAXD3Rbz71biZuGIOkv4doTpVScvaqF7aHHbwgTcOwapcEj7H356
rJkublpy6f8dcFoQ8uAWKxBsIDb4qO/ieirK+ENrMoon/aegML6Viz5sRVghaeiWA+qNaIMmqrO1
wUi2L+H2T3b5kfm6iQFcnSX3RBNLaAR412WLujAZeA0eh/BDGzwyewuBe7Um/K6RyNj4IazivH0K
vPxXlsCx0sPdAOxwQUbLmcrxY+uVvLGn/cawzSGr7Bh9hP8iWeU53xfAWpzYGGUHAeFDJq/WGRJu
X0fsiYM1+j3UkpHNeAJ02kbWQVcTqGVRUaxZ3Um10kmzWIUD3ti3Ma8D5kgrfG0yq9cVo+x7nvnz
RNiJhK2RN9UiFzoBUNDsxhjaIRh2z1kcMoXYyGxPwDd29Yr49zvkm8dzlUwKN4KZuh3FR98qGyd6
TNVA2gtVGsvuQETwUqhtdgn0YjLaIkhOHOc96gQXDbzeFSk0AOwVwO0vBJdQ5Of9Qkdg/yJtMSc8
uZ+TdFjDp5iPXjuGxhSNMfWeCvkYvJmTC0cLXENmq6naxZN42aDD8uL7Ptk3iYpVrbKVE+39M4qO
4xxylTZ5nnvSfUM38SqRfplMmmf/3UwHbjPuRWnVD2gRtAnICBjK7sCZM7c+8Cf7m5DhfngkVc1/
/u5mDh/S7M08CY954EI/3ZhV4B4rADs6H62YTslQX8Rho4arkvzJ0hDHOE7wQxI92oy/EG6D8vj0
esYkshpXL+svOoF4sYNMnWUjofoxz2wHJj/frcn+/gclpr4V86GQYAjbiBjs1+WtsglAdf1ZDMpQ
+zH6nUF0D6VkH/TR7fVyV8m4NZrJmz4arTbUio5wizUe7yJrxS5iFbBzcMHxgJFF9+o+X8HIPFyI
7NuV0CEOKcUub7hIUWXkmwGGGyod3NTSGBaHRFgUYqpr5Kq9Yiocyd0UmGVFiKz++a+Q5MUopOF1
vLacTg+qyiNAGMKGk7FZtjK2/n3EjffEZSgZOztKPz8zcHDdEUxqN9b49Ofkeu9JFw/lgpCNy2Og
NTdI+gZ1fp35Nwt+KvXyfc/8M2Nonv6IDRiyzdgN1Op8R814FK44FM6TQghaanEkluUIWfcOhF8P
OZgjDteeZH3PVJ5Cuk/OO2ouI0nO1UjwYsmrtxReHkBDDS1Vx64RF7mFeeAhC0gjVf6DRlRsp8xA
PhnmoAM35TRsJoNI4LkwXjrXMfcqhiQHpHfOIPHNt7GTG46IvgvY8vwHPdBfJiX+Nix+8zA292Rx
DHOFETLqnORD947hmw5jC0WTrlgqMsIH6fIyoKJvt9DouHcJoEUkE7JxG+EN88VM1srxmuvSO/P7
gubpARARkySoFCWIAZHeMFvXw8ChZU75PYXUNZEANmks//ypNtfCAORaeZ/D840qe/Ig05MSytdQ
3+ZGw942zE6dgT9Z+F5Uuf7l7izfIqiaQpwexETFvsyn2/aEN9D1Pr9nawr7N1xs+hQoSIJCAxS5
Gi/BlJyigw+8QJ75ttOw+Mzz2V9Z8CamkFA6pTMEmC8HYESvD8vKzPbS8YUkaTvEzwzPhZvgl0w8
pTq98DlGrJIgKZR8IlcjSQFjhOnkTmIoM5eMQN1LmbPyho+0Psodq/wgAmsBkdbO0pDqP70MeHDZ
94XAaKRCKWLB43nmyVkSCIPqZdHZKEVP32VkpLyTpg90BOnx6Uikb+RNInSIHI8xD99aZ5p5Vuws
c7Gi0XExjcbdL9tFtRRxVW0GlZFiiKfM9nqcfHg86Yi84zeQOlwpio4osoKDaaVD9wxAtt57otnZ
XxzN7DSoj3aiCCz6qfOsRjV3a+jNJmGVxkucZkIQJ/IqkIV1wIt9jqtpx8Q8EsSLpaFc9qeECjRd
nAXNpdS+ct3a/p5rJM7S48nxNSOWDGjUNie5vyTnGItxCTSxE/VzcLLwpyrquyY2NcGqp2JdYxXw
9W7nugw+p0zwkIiXNGi4SeT/8Ashp5TZean2hzRxrmAVVYCgMRs+Cl5hkzcznrBG3BpmH8vUWPxi
x8ECIIeLuWEV32NWxSfxQMBhrJLbsHJmM1sI+QDkiun5fzLE4fMmKTTmI4vSv4UgcnuqXuy5m+v7
G6whhsuzPN0ULb62N7SWklt7xe3rvRV+0iLqheUAfh7dEetNvPJWk/HJvDdl8rRFeN6HdDwX3YjF
Af1vVn3LfEy0+RoUrd0IaBdBHJJwsnh8LMl7niXKKrpV06AAfmnTgjhMS13hAVjG3n4bdGhMb5ch
RaHLRQ2mv70TFMr17e3WZI2hXeaL189MllYhJm2bCJv+I1T0Zrj3HE7tFicVZ8oNjrIUcgVU8nZX
Z1nzAd39KdShppBjVcahj5RbiTZvS1+m9QBgyn21zUG5iozdYbm/yesETLvrRwz5vcL+0eeBcwEU
WWi8dnCseYqFPNcfSxxerWNBMx9hrnewrmU7+vbzs8cDqcN+cxaw0SzreMHTaPwjuG2AJZatBJTO
ECKqR12GKvSJtGErh025t26edWSDaB8rjhN5lyIlqSLalrolY6FWnQDoNYb5HNyvCsemoMrFRvzu
qgaUH8p72DnQNkhRsVCb1oHkpNJMNj196O+2jMkE6RGQaeqeuVABUxS/xC8pmM++8z+HIkHlqDTh
hQ7/YyW/Gzy1ANIpVVjq5SCBm02tB0r1vjdRsvT51coxJIyUyupZCyxNPoKlAvO9J0amNgze3iJI
/rXRNeKcQRFQblCqIWFLuBbJQ0/A5hQSS+PzTq2hA6RNki7KkPA0NIzBNe38sdYJC5yzU4zIKfmm
nrILEpicnA73e3zgC0WsH0s1ShbhwvzKnZasafP5i0wep7E3dSrv9fwgP9oPvjUyh8SSne25LC67
bj0Ko9CTIuV4JNzCnHjZ45tA68e121DIHXqUK+rjoTZ4/2GHtq2zgqi2Vjrgvu4OWpCfv/CR2nYE
8hu0gu3CgsJOffMBUYfJF226zKAahSWznrnYoGuzhDP7scN1O/PxqCMPUx+GjtjLUpbeCEnXCd0q
03iFJ6FemfOF6RMfkCdHmQdH02YgsDRK0PMNY10Pcs8VRCVHY8vbv9MPgZJE5HEZ2eB5pVG8HuCS
aJteoxwbVVH9gkJ6nPVYIsFe0JT2YnUasU7M615WIKrtLeXIergSJLwlslvpfzlsHFOFYZzeWFEP
M5fw2/tdCOCKF/rxG2FlaOYbdWN+k9jewkuavVMT9jc3Ww0zshVL/ym5Vb/gJhd7P/iDsrc7foMx
IcdYbZdrdk5/io/6EZfi8py6G1n/yCShnlcb+EwKmhveCjUPCrigF8HAICtKj4uvnbpnO0KHHlP2
mdSA0Rb7eCuYQVKbTj/3lCdH6H08lugaayVjktU8/DzNvwbbZVPyXFGmPd30dikMMcno3cggPKXt
WT//dHZflhkoSs5fx1S1CTkm9RDEfxFY7c2WVUPYlMR3n5mMmbSAOedhMi0JaZ7e81a9qB69mq/N
uQdIbpqUH1lOw+9pjoZJebI7sBDAfR3vAdlMOiIz/7K5lMd2Fxr3mEsZSLGW6Ciq/oqJvhrOmDj5
GtUpMIeVWXpYZhz/m+eMOBWwfS2vdetjOq124NaB2/LnE0X0oH/jc+o9lp7mFYcAfnEJf7vNkz/p
XsoUrF53H4CIcHG/R82M45IBO0TIHUpMxXOvItvbk2SpumXbwNQeAkkwi4aXuZD1ZUFfGd00rRKn
uBeHgj9YSMgzExjsGxYE+svsMmHqIiJAgoAENROI4vO3ndJKB/Q61crOgHK6iXjEmFnUb7GG8OgL
RowElM0aoI4rweYDa3gOqF7tLpXkwkxmO6rpzq2/6zRzz4eZQGHJuMHzjU1HBqFz0Hz64tBl7jBO
wtHaarTiMz/UvaH1oKZOwsTNEgVcWmNh3rHjkd9FnH0jRzdjHE0U1Bq9WNj5iYatNmIouS9CEMdt
YPborgmeSw/ycTeEirCoBytp2i64n4iTGo4w1cl4e6ATo5UKFP3uWn6mnoz9Jo5/O6ngKcLe8Fov
GtrBwfpsMQSb2svKoEA78uBs/w7MiAGa6d4AL/m/wnthh0U0OuizWS2mW33ZJyh4qOViTQCOzqVf
lhgAzGFgNUeplYdWzEHDkEDJmsYq298DWsYyj+8BPn8p68JiCDR+re2GSY6rqflo+JPCOTqVQD0n
PbrQVS+Ak1TPdz2HMd5m4oN3+U5W7+/njSEKyyyVdv41QRzIXam/9BrR70VAhQ2Yn4UH/knzkIzm
wqi0eV0cVmGcPt3OTS8ypNi+6fiwOBrJTDHpSIKe4eZ9IoxbuccL6vupchJePEY+o0uY50OJgSay
NBoWLKtYNy5of0N5ydd8S1T7vNcov2QoVKqjRCrEwe2+Edx9P9WSAxfOE3z4Ue8wr177cWWmCI1g
nh0nwRo7OrJxB9ctVjFSllAHc0Zwl5GwRveHFQauCikN+EqtbUNFqHv/IxjX2W05JlZ4Rw4zIcVb
lAxgAgFVBXzahpH5lbzjQFeQBr6nnWAWLgw775kyxlMLqj9JG6brDK4vYlGHEXJTJZB76mCYRG7m
NA/QCsEmlsGPSPEKdlk0/7xdlHa2ZtwzscCt2AN0QgytTPCuCgKCP5Fxu8NGFwH1uEuO1m+L07yH
zz/VoYRhvjh3O4H2UkQxoVkQUo6tRGK7VYOa9LGYc6xYwbz/xhnZE2p5ihkudj2d0wW4/F68FQH/
UFgpZtU/FhxZx0UTruEvgzkauxF6DpzRu/EhwikByInV31TxQoA/wXNuzfNO5pBJyRZ8OqE81Brx
5gHDmsBs+Qgx+xaa47GKCCeQXctD1+ynFob7FXvzP0WJTb3/e/gKmv+NoVz8cBp+r6Fna8m9K8y2
gdm6AXkB/GcX29tTgThM2tSn2XfCCG08JX85hZai1ECRJozYNlEXgHdBsNWzsYXhK/ddYMlmtQoB
A11M8f5w7DP/cG6QOnqWCEvm53C25t4UdhreeZbXCpGmTNe46vFzM2I/JxBPKXraAfPEF3D57N/2
HqN5fdWvlxytaiZtO83BPsJ1N+Px1WquyqNpx1Ie61raEmZmwvZwiBehBWDjixLpS5DFKSMmVSJC
5DnxpznoTk1mM1Hv02c3vbSS4oE5sAo70+jmKntOvbkNh52H9lA/cc4KN4jnhFJIs1284Bv+uO0P
zbpOO7gwoMkVBoYVsH/mMhbjj0JmQNGsdh3Dc2u1irRmiCSob8yONCzdtUQXOZoPX6bebmQCSBNs
1HhdzxqRYoC5z7GD3tycbx084aSvF778vnzXhp4KHfH9DzLbqUaaI8INxTk+s1bbs0n+FIIIl0i7
pxW8zTPitmgswEYiN0jTOiIkO2PbT2Yva8sWzQUhHniZHLgyTUUZAXzHWhzGrJPBtDqUTEgy/0Mc
LLNWb36T+1OnujtMMToWZk6hZYZSglMGubMGv71BdWb3CnF5hwcikZStyOq1HBPPld+lOVGNduQ/
Bjaf3i2P6vIcqdj8hKMyMYDz2HEkGj6mJ550PEnD+eTbBafnsDOipZb5ha6eaZjHdWEPtgmBWrDO
tD+U3BqzDfuJBEoE+tkbkX7nArSAK+7UJFJ7VAewY1ohBHUiBI0P+rez/TZ8svXFaxs1Lj4brfU8
S4TC6ZEvEzoYFOpIrpGQfihyn2pmPYpjcMTLdforF/S63I6xSh5b7m4jK9Vrr+6FtSVQ+ID1JnQi
pgeOb/LotRirtOmm/7tQQJpOXedD//GqAL7cFxuqQ44BEjdD8Ysa30k0+DGmqbkQMqSVc4Yaee+X
iMvy4zLyhUw6zFpaiT8BUUW4nzx6X8oyvR6uPwdF7ir7KpPCiTI7KyXa2IDGQxoiz6NYeI0uvB2q
CEzjWls+HdK/IxDvvu+9A1NJQyGVBQP+A9D0Gnxq7rAtWY7xBEk76475K2rvQgYdTWXwg6janefe
MT1I+GYlXsYxbiZliJbFT3sfB4/0zCNO8ly0i62Qigb55Qn9hQP2sl+tNxm0C5BDFNoUDg+VsWga
30v48A48wsN1t3hRlOuSM5Zp8VBcPX0GZS0ALwVRzskkLydjnSIiWF1HWvrbrNfZ231Q0It0k0Q6
0Rsi5q/8RA5Xn5f15hMTMFA7JfBYSk0rUBgkAMIJwFPmUe5O8LQ53IbUhgyM2If1mo4S/6CrbznB
5eEFRaGBkUmSghdA73ZA9AcSS5uyV+I9AjR5qK1iNvCiR71isjYEPGjMcaKDydOqcgfrgfRB1oR/
qC6jzLgipuCNacuSmIjgPAshXM+26YZZYI5lzUc7q+vagAn84EtA8MAs9+4VMPtsTENZOePNpbHw
gtBkQWcg0OoFYk/DmBxXZWvdcL3Expibzvm64GX/g25WSwgprE0kvTf/uQXQcksY2hOn6m/VW8Ti
fQEG+jS07x0LKfCgMQ426RGJ3TfWtbTUNKZ+HB1kgoAM5TsYL1H1Olt57vnv3R/4vaJ0AdvlsvSH
m7H0Q893xM4rXmnJvUOLFoIWubnuk8kUeQpAyYcDWd2c/+0FbIZX00b+JL+8F76jWU0IABdKGoZv
SDoEH3IBXPlxPcMGNuzgSXYmiAaiaUWg7kNIsNLPb+1qyUcajJh5EcC6CF8H53kQ+HvTAd6Ztzw1
hL/wEg3EXIsMdTKP284jbNLptYP/Wkxav9NjcnnR6cb4ZrL/cdm4WO1WQ9Eh0rPZW58dkEu23USX
Ao+16ez+SqemwUGpSEtEPkKptp2+tD7lzxlEIfoBKJaLCmrN232xoUpdpgziRRufLXQdgNyidL2N
VD9reW5EB5dwj6FfFbADJU2uxid68wv8thRcOxol/qPJeHaR3ttKnwgulDkl6+zsxkDKJF3P1BIX
jJzr7ADnOrARiqOMtEfeortTcTp8e6gSzXiY7AE9oz6xyAzP22pQSTic5NiMbIzkDJvm37rvjF3x
Vt5dsGbBqDh3D+ysNKzhSl8CrCeWBV/IbZ9+WouHIPsYKNavVwV+eH+PLJzeSXJLfm46xlysEQ6h
s7Z5c1nn1+oO2wrZSs6ZTXP95KwPm8F0tsXvuT2uSlf+vjJ91veCaMo4DiNEhlAjG2WSPW7E1hRC
DvUeEqRhtJMi4Atdw+GRAks2gYUch+O4Xvl9+Qe58J2p4dmuJy2JyH8KcYP+LKOtqekJXyV0MQ99
oyFH4xbHwA53IzK7kQB+dTGKVgVo2OYdQRZKfXuCi4VGj9hKnxoOcx7w4mSjxyIboFC+BbYGJZuE
PG09fK/Xol0FK7w+nWUuTIHLjoWx1LZbb7wGW/tIAeGtSjYL1U+hwr6rxz1TC7ieii33ap8/qpLp
uz/AMCECmD4uC9NAYQbaABmc8F3I1hXUmIvyF6TTRBtYv8xNgxr5EQ3Xq4agwYDB4oaNk+sdj4XA
JROXKN+2Uak9itZ9I/Wys+uq43nqxIe3MzzLPyCvmb25aE0m9ep8u+o5mkpNnAIV+ar/+bjRqN6b
pchENKIVrnJ4WuVO8hsgpmqJkVsleRNb+5uf5qUpURWU9q9yHfts4OKpm2hcW5q8HuQbrMLrhMKU
88wkHDz91M4c4JY7ZyuwNWBBLMo1n2kSZjsYS7qwtc+W8q6oVw6W/67hjRnFkleXMTHcxS//qRS/
XNJyqzkXV/TOYWhUm4D91jlUQ+3hj+vRhHVqNToH8eF2IPcZjVOtpAEv1Nd9m9T2XMNhnP//pyuV
YInrvFIngKPSLbXcuhBHqkAPmmpr25i77VEDbWwrVXx+4a84YkybFz27hp9fjxg3N5GwC+yGcIqR
XG6VNoUdInEK1lgLnW8LRr8hcVqTJ4pY6miOJ8kXUTNmbEIseeFO8kVpZr92tNIByrruAhZG6ecg
G/3SN/kIL7uXMpo4KQur2m1IsuVRsVv5nJaM20amBp6szvF/T6FKgr9B8NPBDUFd3Khn68t3sWPJ
gfn4yJykqVOK/FjMCKg6HAwDAeHKh8a9GJ9+68p2Kmdz+AovQVJrE9zJRVboUckGFCU9bIgrscwQ
aE3W8GNRnoyCGWjpFmQKz0Bq0DshQG/PmEyyf209liUrAKEFz7iG8pxqSrTvrgJWf8hWDRKODWra
oA7gxbv7NYAcRQZ7D//5LnBrQUi9QFytowqlEeBmIaXzE+bL262kqLt4ZeFhDeuL3zwho4+LAtCW
7/z48ysxKWU0SGxXKkUPiT08/+OJ98sWRVsqz8eforvFP8bDHkCZYQhbfmMnSI9zton1XsZXleiv
cSt8UHpb82o//sWm1b5jIzN+h4JErFbRorGN0An2w0o4NTM0COYxIC6w0wNaUTYHnrS8l/sf2ugc
VJH+dKLAwrSkfKR+/3yQKqfSI2Ioi7CdwTylA9SEbYZlcZ2RDodtJOvw/3S1G8gWr3D1Nlz/SdpG
5iQqbAJ9mz+YqwDbn0IsB5Rpy/DjsSee+pt49dvHKcxCHpoWKtPFjmlp8scgHdtGedt7qPeh677w
j0swHNzKysIfDtJ4HNmLgg2dXijrmC2J6Qtb7Mpek5+SYD0gZs/vK52Xq0GA1UbS0XtiuR5NqILV
RPfBP0p5LaX/mkEDPp2qG/LmAbHzRje3TO9ALgeYFmnHXUiMTJsG1X3M8fo5IeUfLh6vbZAae2cV
jtazZkDpityq+mGyW41UV3lT2aLAl7rTNt9METBEQs//q2EjfA6k/y3Y5avl3VrtT1CUi12wwzJh
LFAro/080ww7QufskETOTu5e3GMH24MywGp4hISTmv0UnNM2aYDfYXj+zRflztT6DtE/oRv+pFLr
62mt6UTJaF1a8NBG7dfkAFyM6c1IWospFPQKyTQkiGIkepegWeGmUH6tDEt9/kn/qneJBDoUFI/h
rWRbIymoXX9T2G9KxgX/eIPDxvRzbGVX1lFy1lrEYzQcopT+tCg1frRyz0pNTsh7D0yjdLdF1/dy
FHZrQART9HybVhwm5jqBP8E2t4v6WEOKlN6pYcLZaOmzrxBSUQgRmfDMNB21mlsqjvsH+GNcVxF4
A8esOjQP/xiw6uKQOu8cyjkyOOxzP9cIWzItmI8CcZibZPlCQICBbr1iUzcc+keMzXXkk2Xj1xxZ
Q+yqOdutoahfjfPrGRFeCMap+nmXES1CELlJntZcsMMEp8+2SLzxOh39laYAd2uHVB9KmkJuprCF
FRfrjnujvRnzURk1HN9xcIlm/m3t+U2qv4Gq7APqRL2tKnEKDUZB6zGy5L7id47/iN30OuO9tvDG
NAgJvC/yauBkxHfOAFypShTTtPEGZPFx7CYSqbpxk7yGlq0Wk8W2YDY5Iwpc3v/fRpYyl5FCwtmM
XBhxThHP4/VpoLWUBWwW32p0+AjM5vFFnSW89+QKFl+BmZWYkp6TkuQeWAZBlJqyMyofZvFOEvwR
ZuuY44ZOmJ5Dg2dutg6sRgcBSbJX68Jyn6Prjy2n6vUxi/VW+6f6mmpivmhKmaC+Dcl7BZuN4JPc
d9XEqTfFgRamqwwV/WlflHQg3oi/GFKIb/QoU2VURs1GTa4b/zXVUZn3QD5iqH4lh0ZVEXcaVNvK
XxcnHGCN2be60XnUAmAkI+sbcxqjdq5c/0am9lIzQpitD/DGL5FmC2KxIHeH+WQcHMauCE1U6dL2
IiFndO/BUV61xxChz/7IcG5NHE1HmAoRTLraiN6efVH2IYa9x+ri0ZQEmK1dmPe0hts7qQMAn1+M
8hzc0qlPLtbIBqOCvnc9vrnRuO7tsM/s+elYbMCbyptNptr/U0/qUXEIiKlKIBhw9PePqLO+ZV5G
TrSMpRQYzOYPkI4sv215AETc+NBWrYDk6nw5x6AI750nGPxdmhbxA7+9NsYRJMtjU/lblepm4oJH
GuJkkVGFNbK8AxxyodYCnHgG/H1R+nMXVNnf45HYn517WCybiIEkyLMIw3jub68fHPHqaPKdMByK
W0iVoGvs0YCePSoPGzgMprcRzXhCz0x13dXG5mz/ErH49oLtnm7kwwOFFrnv73lG72/IbDtKTGop
qEKOIzueFaKb/6uILp0Cifi/Ci2wvQnrRGvcKBIR0msAFtnJRjdcPcSYJ/QaC1ucK+t45jwG/YRU
oQwF6Jfih0y/GETc36hZEL028xEt/UnwdciqwW+Az7qnZtN8YpzjYiWpX01bqt4oV8+kUQldnmYf
bPNwMzxImu2cfosJBrXKie4S/J90cQnqcbkKTq2Ao8RQox67+M2C9Z3sYdhUkJHgOEuZfO8Ysyhk
TzNZ6+R1WOzfvMc/zM8cxivl+m90IDxE/V4Kk79shj74vk1lcxO9y8GStUUuqNXaXKsvAm2H3UEQ
IB/1eno6rWtkk1d/XTgVbJeMqC5v5tKaVei9kPTvTV5+yk04FMiB0bODnocBje2jVXdhcvNbHKpm
mPmrg8EYl48/RNRN7LhVKlW1mJ03QNtL3lU+12qtvzhkzXF1hczVFdnUHtbnZAdpwY4BtsKieyM2
Afe4H6q2StLqWhT5KjWvwE1/pozbGTGgZ3xzs4d2oiPKM5tVlj5OICaYx0JoG/0w8MgAw0ATxOB0
8lyanpFBLxUWRKjF/sNFsqtQGPoN7QjEwHD4D+R9Q4HNKtRzCbnGVCbxVyH2cHsqYbdGc1Nj8zLG
K3VnHxtjVc4dt33Ys+fdV8DItK5BbfGVf5GchEdAMkbHjwEhjD2cp2rb+jPKS7W17ONkfe7YoC8u
k+HOpcGH1Auq4D3arVmGjJFqV2+PyP8fcFT2oYc+AIFoK1HCPH7+JY8wpzhPBx3T6dyw7cPB1CFH
XIlINMBIlYZ1LulxXDGNh8WZ/9CtF9F1QuWgeDT92+cujl6SVN+u2MWdyin12QGuYGdgU3/LdArg
aUPQbYaUc2ewZv4il8jKQ/a2Xf3a++tpHYS2NfbybTYyaBOpq9qKmHaopZob0z3Dm6Pzb8Wsegms
9GFSYk7FfVRC2ZfcUTsz8ggkiNFdRMz4g+Kqg+gFp8GlKMZYOQwPdi0GeVz44q8T9tJMhGY6Q4HH
hiXbuffkzbV5+53CUBQYHGTZbkXKPqzYzUGtUDf9xKFFMmMZdmsTnb7qZdu19ov+2A+yBol2wia4
C7mgroU3soafKmImYjQNR8PA+CXBvpZA9WotstA6Mudw36a2mEKn+PrtroLZi5YtCEhSoC8AnzdD
I4ONuutopC5DzXwTk04xtReRiHlIe8QGHstVqnxxOhlSD3n59aohkUBofg2pCHyb3IaDIwb38TTu
EoX0/Ff8+ss2OFai07ujV1Pe3Yp9rDufp409dW6gDd8wSG8Kmp90zI6Fm3lHTxX+svpFHvbrTdU3
8aHAfX4njy7/FHaT+kJIYFg0ctSaWamu9UitQXR1dh4765FA8CSAfLadZuRm6c9gCdv4LUFu0+jS
OKGtWprK/4Q66xQzKtB7VsMyXs8xdbFNqC6fURMhPfNSm8BLkOtIS36vYyc42X8JB7m2pVk6cSsk
BKLbBSLytIDxWPuxIvAezENoAmvML+oMrImgQJSeGy0H5XJgb6sin8MykTmltHSweemTh00UdDCE
JIOzd+eUMvFUV/D5gZr9XIGeTfXtUQBkVmgMtCcSM24rvpacbxJFxHKWuhKBLxuYVfarjZ9lv1pf
O7bCHi2WmuZ8f46EJgsIzSjdAJdG+0X1wl6MW67ZZ1FondcROKYc8FNwIWDWf+wQ6/TmpKBKgrAn
SS4QQnqTDq9q71v5bP22W2YS6fQB75bqJ56Q2ZjvNfgwIYPp1gmkWiTpVB5cLxalImmrCxWemjZh
LoX+t3KafYLORN28+8B4zLAsrs/+JVnnHGaLaMLZAKgJNkIXyN4RPAcgGx8lNSxT9bNV6sPnXotc
8nQod9I8MlupwEntfD9SKxrW8Z8QOrmopisDdv12QMdz+asAsLNH7OwIBC6aV01fFMlauk9UVQD3
0yKht9QduIh6eOs25Lwb4Dlrdjyd3m53Inj6MFalXnF+D6ViellomSPGiGpFRhaW/ByqDHH3xuqm
K5Ruq7W1uzMVb0DBmVLMviGsq92n4yRD4qTaL9fRuPekV+TRRCfeL7HJFvnHYFn9SC9LchJPrgh5
g8Wx9+On28tIOgJIFeKQGeT3AT1Rf8XBqhEGFpyBjGRE0loLruWTF5jM/hy2kBRaTOHbBRhiId7Y
xXu2pWgEXD3GxdnqcaGwAPCcaDQSJYEy8S8UXlelbytlHSFCrxVJNpPVQV2xU5f5UTbFJDlkQgQy
7Yx8R+h/jNwuwmyRTAPAMA0rvtHG7LFxI0rJ6pWo9Bb9Shrx+2dDdzZqCWugW2yh9y0WT0n4rH+J
iZg61o9qDOE+6qQk9QSvIb7wvYijlS0cF/KGt22/KuMJmi4CYMMDjhOFLAB3BPrPOlQn+o8ZAjMn
N3v6b67ggNHoslrGMKwAP0Bcf9ynUAreylYBV89O7AythRFgS8TsEwWwg6TNkZOknq79Vet+/yna
sdoJ3M8e331qX+IQz1wRwXOs9WNh8/mtigXQX6fAsgbr8nok3lKki+HV3qA6SmJZ1WUBncS88YXM
PYbAXLQoi2cIhd4vVQDtnwD1QeEyuUymWLz7/MYHpszsoc2yd6cdrxu6BlElT2eisr5vqs9l/DDC
B8lQJJLnux6azomtORny+d5j+rD6rmo+0VAOfKGZW7Hw9/eJfW1P2J3+g3wNkJqMPxWXEV60P6xD
ta7eK86vHy+H9ODclO95+I0xsD7uuMxwPi5qsRRVbPF6khX4bajuKPsocxIakPa3nXG1owf0n2yi
qjnb7ZJerx5YRrI2eSHDAQz5HN8tmpdbBUpL1Hm3zf0D+NF6t6BkaPbv/wrOn3Zf4tpqQl8fBAaN
lcrHMrTpS2tzfiYjLqu8X3qGqGNfBlDjzIusSPqZ8DSt43BtQ7rqDhqpRtdOXkrvwxqe870QhaHm
IPEl+w096+kpzag6y/E7FevSINHltqH+2tOu6f+x47ig5HFCnG2Vl7wJFMdZtyxg9qk3OLWuBSNk
hI+x9EF4O0tKcV1ILNVyJqfZ8zz/Gv4Fv76fH4I6yPgMwQXKtvSyqRv/uRt17PemWiHAHO92Dr2+
uVxG6PZhD2Fka4i+5j9Bd7EexkxNSaSev2NzRhm/KbcOK6yEJ54iGWk6BCqcJAXLVn5Ri/ZbZbuZ
DwDJ06tN0BVEK6BrddYOD8WxDgJCgkUWjP4vQUIwUayt+tqaMUfP+zLC+KZZRRpDke9qQuYgS+Sn
uQvpw2dhMBJVv8bjX43r3pRKjNk5RHTG5jTq3xw511S6rdx6NLI0w44XfFAUofu8hBa9gJqGdX6o
QxyU2JQMT8LrOT/L6QCC2NhyUYVpVg9CxdDrGgTNHZVFPeHIxVXcW7aqgJZneD4thp6s67pVSqDz
6MoD/9eVR85k8ayofTycadO10ayamGd7r+OoA0SiUvThz95ERZgTjXlW3tO5CZX+urpCJou8xdpz
cXFkBD/2W92f1wri7ZwQwcd/kVAvm+ClAiHbEifbWc7UYYVAEaciZkfofnF2PdUhIDreVg9CwouD
7zjmcOC+ffRxIRDmHJvXUxzZsleNaMtcFJblGYH/EurQrKDEe55rg14iim+9O3C+udAsgZLqjR1M
BkFi1XOEkQ+i0qbLHwhulbeITHgqXrEkHt431feJgn2xqDrzcgzWsUy0gKjIZhkaeJ4Yf3ImyWKe
l3Q46nEQ1cL9h4R2yWca+Wh8KRVrqkDApS0L4f5OsvsfhtYesTsNY5dnQr6AMUZATXnaFC308ZHg
v6ZkDR4c9o6uPdq7NMN2KaHQBa53cYbcG5J/Gf8VylyZsPQv5mwzpq6CjTwww2JbN2Rr/ehcSFxv
RmngCJi7byNI61HAftvrrA5/7rHzk58qlXGY+Uzo98BmPnhYASvxXvRSJuj5Bx95C7R9n1PUzCdi
1QmdZGWGo5CGzpdw78qQ9XL28QtaBcRDZC9K9H3aFeZl6FY2ooKa723JKEdr3MYGrucn1DYXTvwO
qUGRxKeXgwZN03osluQK4uVe0T9yl67DG63mgTtjO5VzxnoIJSCqGzeBVuUtlG0bCyTP0cdvgkN/
Lxxh06yAHU4u+358VSOiF8buPFunj6b3v2z6Dd76TatSnQVje+ZtQnT8ED4vUsBpyPYlH8SsoB0J
zAqJXFly6tmdbD4I0l2YZrwhrtEAKtzfsAbiBpJa11nQ56fEmNxrfC6nF1RrtPsuYRBDrVwtYcJ0
ePY6lcyHeDQcRlWzMIexVeJnKrPN6CBf99lB4gh6CZs+dgGdG7ugyjwczh4Z09GQT6ZCmW51L+fy
60l/UWSqindkymyIjdQ6WnByaZiRTLN5XSkZbJeUHOhz6pwLi0ijTqv1lETqc953arI3WUHEyew2
tpO5oTyBBtmednLIEUngHgl+uV8anA/s+Qm2+rwStjf6arBStZawN3krWKzdRoccrCU1Xh1ThPj7
ogDNrTTX+ZJkxJBVtrsUYHcF5NI2bwwd3m8eDwoAKaZ+lSoonHsKWAYm8WqmT0xGIwnOHayzHaN3
b38MH5IJ0H/wWIYAeMrRlXDsG2gA1ifbtcKS6KevPFM+wca8zSmQrfHQdFxVsH6lpEloO1VTOeNc
q5+SQoRPmH9Jt5B1/kg0iCGBC1ppmi+Zxtt+0EYGdHXqJc6uHc7PWhpo9BdJtGvGvlWU+iQ+L+Y8
Ap2yDaaFHssBfuPjQgVPoNLTW1TOvFy4KxICSX5Dt6t+pd+YSZ4ThSsqyhUK+wWaoVP02Wpd3Pvb
aK2EvLahtV3ytUMXUl55JSRtZF8rf2Trufpqg2QqO8Yn9lKRepalX/bpHqwVGKNSFkhYKv2rXbns
bpYxvIi9QQzud7dhlhVjIYEit+BnKvz8HBe9Rc92ASOrYjHH0jrf5/66Pie2y8SIfZexKc8Mdv1y
1mpC0E7hysFikQOs7FKlZ+vIMRRfnvOYlWJ3d/ZSL8hLmYz0q53as2bmc18V27zfstftkYpR3WiL
+YpAR57ac/z0gFyDtAMUchkRrmtb2oR7VrpE6GFY/9UX3C4T28GDNJdafFGUcHTmpl6QAnE9ufus
jqthGU4Q3U9vfy4Go/IQv6bl1Agj+pBRSi/EocmeyVmQvPGaZ1y6r2nuL3Wn+Wc15/MJaD50aj7Q
9/bBRbw8XVfG+/Xjrhpl5X2lpOzriqxrwzzavpxyUWGu7mwRn/leTYDR52acE6MHxlnW8e5l6vlG
01lMjKYvv2AFbPMgIYgxFNepK30tXl99KnyShTpe4qp2ZBURZcma/1pXk4jtOVBWFF9Z0tCKb1xy
fajQkKyKGCfi8drdHCqFT6cHsz5jj5hY2m1ic+5UEhjM9V/ynB1fzfc0zSPswxoY8RalRJ5oeV8B
6G80KDUiIrDgsU6JoWI/J+BqMZFWXeCsPLizDuyBpvRvITzBpwRSHPLMRoJEGsQ7GIZHZxYf8v72
HIrDo3byHIbqS2smznzD6t8yELkfFZl5FpUmqw+GJ6kGoL1PULLD11bB1gitMYB/KEY860lV35gx
52aRhIeyU32C0i8zqCIxVA57GoUSfeSgqFka14D+oU3grpfIpJ1Drbru5mZyIkDKDJ0rEwZr0SXH
zUsSmpqt4weYfwNiRAuQPCLlzqcSaV0WO4iK27SMYe4ggLsK+cweL/ByZamiswrvokl/xFBD06Hz
KleHe/VTvAw/sGxIrkoLTmxe6cfE+JSYHh0ZFndpr3KXB+VaXBtHsBgPEkf4Boz089uXUDavG+4V
Z8+Tv1fUo7SCi0fTZNEi6f44pC9dJIxVqLoTS3o26YDxaAQ0WZCmXbQDucGHW3Rf4FsF0cu/sNJ8
FYJoTG4VAlbicE2W993TAq7zlgA3HQgM+VLLxHKHVwhxVv+0Rwui4+cTA1kRHIU7dXKKHcf9ql2w
4Wc80RhJq3oC0HTJh1dlPXt9ayREpewOOupbqMTiJcS9LwRCBJNyIBCboaq545fz/aw1v7rcWI4k
WFJHKCGH13Z98yO0h5VnxpJcPhmnLGhe++DlnWYimg+QN/5RI1qZRuXkYbOjXaMhCVM9is+S0fmr
xoCY3gT1eZJVRj6GsI3rPZR+Xonp/INi2zhyAp4kh6oKySUAl+z0z4cUE20+l+T4wWf+5f1RsXYF
5GxDkEe/aL7ebU49SHWqvsY2Qbc6tNyPftjdapOcpTI3D0IXCQY1jYfDTnEUUZvk7Ne8MnHq58xd
ltNKLHNLP3wLy5m59Umw+L+CuBpOTE6Lui6GW/WP1OxVgrnAZy59TSLMfYhKK+KYoDPmaPN/IfhM
grVL+fLwlhUFKlAD/Tzu8ujuqRRNERh2Xdo4IVjAH46k/CSKul5cF8tUwB3TnzdgPalqcIq4gSk+
JVzyDxBHTrl7QJWYxjTrB6pgebXSvtBgQUoCTDYn0P/upagpF52VqYq/mF16lagkh2RTdHD90+h/
+9O7yH8pHWKqNHjJ9n+U4lrAtl1JHhChlKxo4MVS9y96icaNjo2FfYiJVhDHfXLGtHXtk3LGdO7O
SMF7yA2/r4AN7pO/XPk2hXOZq0RZD15DOna2qXIUvWgpXV1F2WjoITKc+7jKV26FTZ6RulNvCLyg
49XrGJpez+15rChvWqPSdoq7NCKuwAWHVRHY6f+fNshzYLieYxFVz0M08w4mPQKxpnUf6ljYH3vF
2gYHKIJ9MyO6GIzDxKVjKjtznplcV+GllvF3n+tdWH0zbE7M6Yk9lGjurcsYXrUcA9vmN7vBDtxs
9XHZ8lOThOVGa6Cz+SCdGVje/jX5hs40YjSh7wetJQGFFq9RqVW0fDme3aTJ/9FQPdJCXCMP2xbX
js/G3aufWns1S+HBUQGW7MbJT3qlaVUL7eemD4qgU3OkCSO83VKzjx3OLp7xxwwmaMJXNCvYy0ez
KNfCtaxJeyuczJ1vZTFLhu4HV7yWMAeHjaHBanDnTtnlE1TvegKs6db8bAj8FcCAGZADRmes+vE4
VyCWhZY7dPe9Dy6BU7AMpO7hWCVM7ODgtV2I4M1jepDCsWcuB5u34Kop7IsShci/YdCPZeFikqJ/
RFdIwIqI1FM8NCUsXCgNPmgBqpUQ8Dpn1nkxchB4JJsEcU3vwty7AiC8b2QkJ3O0BbKWTIi/lj1g
b64LAetcU64Zh3PDm7mGfZv7zHq2wv/7zBhA4dhUZVb0xlihx9ESeSSVtfj28KuAFD9NdEmrl7j7
KSEqFHzXQGC/3V1okiac6NQzFOT8LaZyg1L9wpMFvXtUt9BnDYxJUNZlicdhcyl+Ct9+qMP8ryn1
y/+u1Cb7qmhEOBY0uhWZ/Pt9Camftk80g1YkBOGpqyoX4l1uLnSLUeS0jg1LIc789G4D3r+tRkKG
dr6idVt+x0UBOAd7WWUtumqY+OuT3U41DJKANubTzUkydHhGRYg35ewFRuZFLZ8QxqGK3jsM1B2H
c4jbVZ2Ca74TXXQUQHXRAWPyNFlNB7hCwXmqHfQeo8lXEZIH7oMLNIVTs2NQK2+rE/qUyQuq0Y2G
GPGfSmJ6VtZagqh81ar7Deoh4ZPZSUATMxmblDyoLYVXVPDW/XJgRvKfLT5bh0STTL8ByR/vI/34
ePmmGR3T3wI7VTMBx0Wh3W+AB6B9j0BFlnqwWfRcQgXhuEturLCJL4dkHIVCO+6bWtlCIMn1ZBcj
frW2w9c685jHYvRhZleYURwm7VOxHofHh0dJH6dBcFjN7dhKBCf/7P2rqM89gaPwbdpkA4tBNLNt
M1vPM3lZDX58EO5BIn+8mUieZECX0jFeWteWgp7WWm/Ttfp7TqyMWqWzAqmDgzw7NFCShok0guIV
UoNOxZ5mpQpDtiZi1HTWsrv2YB1yMFWXsCvn9EOz4d9PPHAXBXFlFRGXzT/Hl4HxUTCJ3z8J0LdR
c6bb8S2jKL+siubNw3tC2lgsW/oODsr+BuyS1xaxwNVN+qfoAzAMddgj3J4er4vx0WtWxNQ7gCDW
bjCcYZkhH1jRuDAHuam5uUf42E6s5v0k9l5RSyYf5Hf9qiwQgRigyLK9IexalVxIXW0aWdDmrbJR
A6nNmLeEVI/Osj1ClwGGc6vlRB1N9T3gkt76cdNtvIcFWSFvw6JT3KoaQVy+mxuhIUcSDeRJT+R8
uEYHddn6r0XMhiZjYTqYfwNdTaqZC3H6cAU6GH/rIa6/FNlgjje8afZwcj1hItVhbJ0G64nzKeTX
xfRtuAOKa7YDQXK2WfWgf5nOPkL98EDMdKu1QxR0Dpw6OUisKDwlcQpS2933oQMJLyquThOYnalI
x9uCbhSzU8n3hQCSj6KDeFKxGwH7rflgMWF3TlTFQ6PmOLnC3zvVCyz+69Y+8qmlmWCX7PHiHz8b
0br8dQ4dNTxfC/3UF3yKV5Q7kHWmHdDHdU2Y5TBVn8R65FYZfLEEhR4x/XnRex2G6myWo9r2odbT
XQD9wm1gGRq6RiC7H+CdDhsEmKnSWGYavjP+wFW3RaWdT2O7qCnElkcGW5shsWio4kBdTGpT4u5G
VoruN0zGIXY456MUPwpQkvVWVpikrqrgRrV0YbOxTYXebNSrjsBWBcRTBIwvky6Nabjg8Grq+lLI
Uv+CFEDJ6SwinFUg3wQeeNxOJKXGUi6xF7X5pkM8zl+vIfPvTEEdwxqJ/y12PG4RkQm06h4w9MlH
Zd3St+k+s5FMC8SuaJGm9cjWLwNWFtFc9aI79SnHFJpQCgCrhpjJMSEhzagJDTKjBWK7al+pwJpO
OWjPCsamZOgDA4mbTG943nKWOdqDhVbkwYyCr90k+Hp4mv3SB+BJNZhM4vYGR/dt1JGT9Jwz6Onh
ywMqBINCu0mV7KeeJbn1BmQ+UnUS0VRZXlO07I0IsN3WOa8qb7iW6AO/BaRvFWWdvATSe4Xo7z9h
UYmnTlcMbhEz6lJNOaSIXvdUyk4Guf0oy0kHGWSX/39DJO5I4aHKrc0Gv+lQO+FmVeu1GzvpLF4G
5KLVbFtOGyayxfCSN7pXrOxVpvn0VQbWAlLAqvnEymA5Q+Eft8820EisCZgyN24Vgot6eSdy4DvI
QyF9aXhqNWAI4XjTLG+v9/Nnou2L6QFCwRfJmWDjvKj9Zux3BJpkLIDx8DGsAiZX0ipyWylUtl2S
qgtGpYNZ7KMcKLv0galMEuvblNdPFkbRnGRNlk/FTAynCYUPaCieMMv0d8sN52Yywcj8jeeTy0v2
zb6qRXiS1LfbllUl11Rc02RpY0k8veLdH4OQMhp0/cGyJztva/IPuIWIDf+C1JIW+Fl9AiX7wAqQ
5Ml2jjjQZ8axjwPpgzlyu9V/o15/lvM8tEqZSeAQmpxrP0ONxy8sg5XS6igpZbReBiJOaCFpdjMT
y0q7FKT/yA+Z7N6p1KgnAsjvYPBSdb1qwnUctghCdygIuwFUdzE+h8bNyUMeYqAFsIC0Ax9aSFJM
Ri53xHiXx+uMWc98Kh3bMogpsocL4YsX4lZiqnm6DWS3bGsqeGPKVol1bKDpqb3ohaVyWr/6Wx92
GOqUAj57Oi1NkSfKjmPkHaZn7Cw4nIRVc2cg9OIxVMKk3WTEKekcwWAhBmm1DsGZkB57z2CO84Oo
jlbpblO9exwhXO3AszgwAqmvPM/XCUqjNneFveuz+RoR+GWCFURTtuFpuiWkcQWKv9YHYl0R6t5G
wLVR+/shm02ev/Zi1diBXAoKuqY7uCJKskJN41NoRaqFTaiNTGiTFUWlWiz9gWk8iSoaGyeVY6Um
+MHylRl9cmvtt9p+6ZR/T1DEaZrHuLIvdjDhdsVFbpcImPoZfv0r5IeKJJThoW4jqjRwdaGOhCgP
2zVuaJugH0qjDzU8AWZmUq0H3oKMFLE08dl7Nbl7o/Gu+1H3QMLKt8TspHqezuDpJiWagjv1LOAo
rdAgoZmBkK67dwB3AUS7YSZFqri1Ka7eCUHbcN5niXlfEjgEcWhMcNLgXd1fwNJVgjOqoaF+/kMP
1vHVyP1zT/t7LNTwwPqFzLtty9dlA3wyXvejs9Sya1Fhjz/LWiy2YLbKLKUUfIgIhT56jbLgQB7H
7wmrOihVtq9Im8NhkQA8ZVzB2UpZjJcpItLYcIAJrz+DGmS4yWBUSz7HV/VkPXv8I3SSTRU4WSbW
MkP3J+vlEqQKIEfv/aUrzksyqF0FYNujbvxCFQt38BATFrC5Mju4tcc0tzSQCVrATt7cw8RxETGz
KWM4ieRf5E+to9p/xUnwbVtLOzzXTb8eFDbdzZEtxa75D6QOgcHhjgmoByAKBHCjyCZHcF4vbMC5
KZdfOxFKJCuoIORuKMqtXx6PQQnjZ/i7GeTojMSUfGkk0GE2VvJ4Kj2DN6/dFAMIAJTUo4/+wbPT
vyzRU/ek1pmrL5K/+cEyhF2b5Htppez0Niel8Hgi7ZUIErUpOlNJTWlAoKhDtOOgCs8lVViskVjw
L3pry3YpRB/A8QvjWcBXz3hxUGjkEwNhEouOsmxunjH8D49FKhSCmNO/QUdtkbrHnZ9uJGodtN0d
zq0iA5ObDN7XXPSqwxqzLdhlNMQEEHIr3kHx6G4ZcIqguq1XOmc9RcjBaAIRnq3oVxUrz2E5fnqi
+j/whdcrSl6aa42KjmbNu2LxJZVD4nOdxizeUuF5JpnRY7CEKWgaFJBNMDeOZS3s41/VMPDq7leG
Iu41h7nHmHIRiIOi4dZ7fMVuYeTyjVY5wHA1yT+IAWyGuRAsXg7IoGNVKzw+uzYZFyUzUSSWj2Rl
duw4/HzLonU0/lQWTxf9If3g2zhIgnXYE8ouWMY3qWg09k7hhCl1tU8bbvzjOf3imsTaHw4VUpJG
h5XEDchdILmCXwPzfrTvEHa5zUN+VqDd4OpaEb6izV0D6iSIs4JBaHe/OGiB+nZLOYd2qpkPKaOY
VymWbruArbfHVzB1uQ8acPAJZYA0zHTrX1RnGBKsVkDTisq2+1GtkcTXPT2KMykAVyYjI5ijw04L
Ym/CiCmQ7YWhM0tpOJzJ5lymWpQIY6pvaXak3WQmRnxXRBLT5wbg3erYc1tNHRgPY95g7Uid+rhf
BdqYZReoujlw3ZBwJSkcAFuOZGaCdFShrTU0rYUBVMxvzRJgEnlwJkquzm+kBZ/LtvcjrNvQZkgk
owlIzkP9SkpSRKxN9o0JQsjRUbuQS7RLxB9prV6J2RQIl1DzWDrP95FCpbM/9Bla6fa5sWA3/4aB
YJ9wKxXBDkH0bLwYVUyEC8zoWNY9KQUQICnhz+aKp3JbO7wzvr80Nv4TzMbhkZu+XwmZRMAZD8/+
UjOb2Po+IT0/V7/pZ1PuhMMmfI7/A3fdovF/g+PlGnuyLi3A3/9shN7VrhcHyNM1R7Qzdu6pDZCH
aMfWim7acq/n4siPTe+nc9t13J5kCzGhDHPh5DNC/yF+W48WSlSxtTE892Gl8r+yFkyI8QXNXxTP
D+mVBFoSeeEtRiOZTDEohIREojuslCnzo0QgKQOJtILWlSWzdKwWyapK+danUBJFRnxkv6hicC0+
Qa2SMvlqZRceF25gsGlSTu3vP2f/JUCslvKPsYZGKK0YD24jK2Ra1Ol6kZLq65J33GctMM1rlaJj
mfBpWxX4nfRsWX9gyqWKz0v1mGZTyT2rVxr2rsMDlFtisFik7fc2V8dUB1USOZA4xv/USt8TP6tQ
3RQw1DDVUBuZTPvm6IMzpwWIcEH2iJYoqSh+X9MCC64DYONv1/ROLLZU4rnK9vi+NOKtaLSa7Zx7
k8LGZNNbhYgZqoOrgWwuhORzcD/YwIQd77ex5cq8ssH9Us4fC+5iDoYcNoj9thgrqv//NC6T5P2C
6ph+OsVPr4PFxO2oWyzqZ4zcm6NC5Tx7LscHIyq8R2Cmem1ZqbtrqHpCRFopbRfPJin6YE2/yIsg
AYZ1KihFX222vGHbnO1dHoAeAJBvR25O5Rf3H5Vn1CMqFzGrka/GJDwc1YngqCQUV7qChfiOhMay
rP0t1U5BDFeT4ML5gwpXhQ+aQRjL3aXQUwjy85+U1yLTWuHxGinNL4p+KHVf6KLzNKoVaDW7b2A/
glspnmlrZnssu5kAYAdoFUtr7he22kwfpVO7PFUbJLk5YUvFs2emE5PoXFxXIOEeQaUVs4lE2Bho
ryB/yA7dfxiSye7nKikNkinqWHlKst5nMxUOhiZzfiLtCvCMvXPsxLJT7yan329oG8eeQQYBAVI4
p9Ch+cFHqNbelSkKVjGOcW5TDINOT81WP9giXRjUbjy5YX8t9ISzpRcpzdIqnjarZPPyrYLAXcOn
57Nn/ZVV6/WyHFqOmZjgjXxLetmofzwRxc0GFYG4zAPeFyakHZ6GWEanC9wCfy/Gl93EJeN6dtLE
wFHakdT+zbit8kuq8kd1tJruu9yJz+DRuqhivm0CF+Ww8Cmc3y4Ypa9Hpp0j5e7EaQyBrB7BVv/I
APRA5RuqXnlzYBhf3QGJgPboGs4R45q9mononZrUZvPsa4XLfhk+SPbvn1JdC8WyTVK3ZHJAzzuZ
bZ4L+Pzf8cYzShq7F3vnQTD5ZIzNLK8dxTulPilgWXH9fGRQeY77kEtl9DzaprrXgTCTd6mOg3+3
gz479v/NgGgVfTgLbx5oa/1Y4i1UEcxL1TkU6ZZ5Xh3VweHArzqxjg95MEMh2+DChUbPePpoYBu8
dqNyN1KKN5Zzyw63LvTemN9IkNA/uIHIfFH/jWwAocNE2wkO/03L6xGU+nqqYmPJgqsTqAN9NZNI
Pe9tYcEiwYIJGVBWvRDrrGv5ZXIfV1wtJ97hiI3NwxnAfNevlG9YklsF8ww/SIVn5aiLjLufFOd/
Ot74GbixKO3QPJATlZnfddyCyL7kKWweRkdm2VeYjHZA76kMoPgGIKuh/BxeAXSB07jy4tmmR+Nb
+rYBwt9O/SkipjYOZuGYz9wMhkU0r0td6GVMn+VFz/RwgAvdr0fkaLbpLBOh01eOf+SPtuPNPi/U
7Iou1Qf5AesN33/OaAh7A1jxPGz2NBD4XSeDG05m0gvFZY72amrZpdsA2CBUurFhzZVOH8taLXd4
Xk/hhKBks+OJtdbictJhnWj4FXGwPn7QE16W3gDrJWN9d5wXhUcuW5yGBt8VOS/BG3p9FS14eHMw
Y2qTcoOd7SzrtgV56i8kBhIbXVBA9HLMsJQE3bKGysVctlEVFk2t2ALkljrtqqctJhmI49nRUYak
dgUkullP3BPADv46Dzcwk+srAKxTbKorTvEpaHVrhaz6MfeSMWqIBVAV64s/1Ns23SIK6Wtak5as
5j3sFnG1BXqDzLgKRhHWL4v4yGNn9QKKCc4FYM9lfpmxFxTnu0yqysUTNQGao3XmxYZalDCtwbVA
iGzA1GiwswAEK2OmXGwizbH4rCXYKi0+XS6u96CzhEaJe8K4vciEk5lg9tsX9NSi4u/FQ8/Uzg5d
eech6fLj0MeWxoDnYIUQTWpdypYkULu9EA9R98fX8o01c0B2Z766sD7Q7SR96Ru7+Uo93HiBFfYR
fXLPrCb1qO4tTTmKMIpUscE+MDbk0rB35as4fJ057Vu6/P8vOaiLWE4MV9HBBYIufZ128IPIPRkb
lZ/T8ne+s5cZ3DmMeu1121bd9u+QXIVJhshIRgn/bjnl48AQg4GlkWcgbbfSnqjKKl3r2SPbwz2u
xnAgjLPJyjmn8aRT9B0vM7uN79G7xg2CoW2D9mHgtxJl2vNWwb4YytNQAofQHxs/CcP780a78cZd
xdd6menP/bEVs+Gi0Nanr3SHzuP8susP17R1TZre24QkfS/JBC4Bxgkr6ne7jsd9ZFpvPjE66hqN
0cp/GNOwwnx4ZAojbfqiQ+ZBidnZZBV+UexLX/rJRaUGtlAX1+J5Ls7mmVZLhXTUi29Oq5FCIGHf
mTALSgJJ/GzxOiIz3TuhxBGlej/ICH+Gb7M/vGA+3S0kJZ4rzpx5zkOty8hZeadfAfvhDxXpeVYy
01YqPOhFsmSKo+VHvEN8vgwu+OHWzHLJkbhIFQKlOCkmQOTKJOlaADZ3F69leXrMi7Rfja+VnsR+
fpRadUSXp21NR6BK/WBbpkWbfAVLzNsINZEtGq02bHDvn3NrcbyKF4wt0g5O4aEtWNDIFXAZoYBH
RbST/4C8wEKkxQGZwOhLPy6hJyNq0/AP8oE7k3QeY4JhN3zmH77yZj5UKEXP9ggYpycHKZHWLCkX
LNO8vkDR16xzO2P394le0el2GgNwz//QAxiWPUYz7QD1GJqvBDJyco3r7Fezg3rQINPQphMosJtB
uPTTevqB1FADK4WTuUHuyTQkxkZljspdQ8Rnffs0TWtkvqgF0EHEfH5S0/rYx3znZ77Wc6oJig37
wfBU3tFmWD1LXeueR7ShFoVOn05fX65xLLBSO5k7yvVPmBot8ysDlfdTMoCMUuM218mSGLD9ZOM0
n2WCeQzwtKWIg9K3m23P8EPqtlmM6eXwqU3xG9EOWaqdmpo9v3v8oE6fPSaKAtyas9qfGtnyLW63
I16ky9bcYXWOQiew6VFkig24hTEJH9j0/I08Y83LmSrlmV0TcZ3ejJtZm47SVJyl87sH0kJYWcZJ
uFFVKlT51yHHUFU5WD+5oiGWo4uF6wZDgfVMoFdkzw/0NX9aVlfRmNt5kDQaPeWiYeFLxUdkHQDg
biTJzQGF3GAu6KV9t/5cUXQHW9cg2lcvzNevteBW/k3nDfnYdh6gVuKREgQ2tFnKH24LgmI5uWoa
u3UltiQaQEtHqnMHU12I1w4U09wLeKyYZDWWrMRw2wC5hB4UuI6Gu5NooECIMxaektccThu0TACI
0szC8ylmoCs9U+pLF+mCXTVHbrNvW0YFsVmuIeBKZuGK7lC/q5tJAdHxxOU8n867u6Tcqqcs8t9i
UHRzyAOzwF9bZyOeQ5oSBEgZ8M1XN8gYi9sRRbNo6cW7ajS5lOXEQBSxDdkSt+DZzSjtGhFasSVF
D/cCO2b8ZBFo+mhPI4RHh7iyTgYbKfXdzKrNxrTCxlM9ELuPrWgi4Lge//Ul0ZdjTJSC6wTleUZX
sBATpnJCCMRnnyRSZRI8vQvCDqp+s1LI3erlUhJEdJ3908aN6hH1f4CrpFD7UdXDEVlQtSa86BIE
BboGZpnL3sTDrVRuE4Mc5j5/aWcbDWi1pY6axAtDnlCwq5hthlgcxKQH9EoGfzf6klwgd1IjNztU
ekwdzoVMvC5y297Or0sy87/P0ldJUtRql3sEuvTIiTS0fIqVSD6LUDnJsTeb9qJu8HG7HIPaDUlO
YAt4AKEpfr6ELAv7J5r94wPWQtPuh4YjdHCKS5oO3tWmDvx7wcK9HHFF3blImujAnuqEfotOyLqH
m9nXFJNQbQ/x97MYqT9XXM/wasOf1Kl7RKlygwvL4B3V2V8Ze0I4xHE3D7qrayb6rvRAW/YXqZtn
JwBkDFZUTSo4LApQf6+11JFVmpuy4gKZ5z3TJ7vGodoTMDRAtWUTTNlACtAajcdwSOA7JyJ1SnSB
KySpQjuubZY3egjgwZ71JEz5S7NsWqBy8vVvm2PEtLxUX+5oGV9bxV5XvFe1N5rU6Mq3Cpj2l+ri
c+TbXTZ+ph6By1/Vfzt7IgD8jBIYEqzkGDd5FxTBrc91+0muAkpHE9xlqCAH5OTEEzkBzpGa2Ec7
h86BMMDyeMQRJ/g53qpUKJeqQBnBWqMBYg2kfCe15QXqXLxgO93yKkPyQkPLwgLvQuWqXsjIPpa+
D805SVWNBbo58xCS4I6qNMrBT2rOqW6+epGfm/PCV0ylv7NhuAlz6q9EzEyZfaChX3C1Q2V6aSqP
Jg85nMAMJoQZT8t0EMAQVi7txpiSpBnPk/5PVshQfmJ3+d9jnrBdY121xLSK2dDdgcNWC8XIz72X
EUdLqB1BczlRYOcgKG6O2aq1yVhcxefkI3EmKxj6Ufg8B6Vv4ytVfq0WVeqSS43zd2TN8yW6VlKV
wqUgyIanf39jFQSTMzbnfJewvVLe7BKqpy5ZN5BuZwA+Pm149bgt5pOKSDUE9mpkhC1CghfFwiEC
WEV6YIWligWrXPkKstqxaHRxcgFVutOH/7Qz4gzZMw1kkFSL6eJXBZ2iDYvKSySsM4/N0Wd/VpuD
h1FCmCIPSon+7OVcuNcP/+7Dq/lqdvzPfjlVs6JFIrzgkK1iBx+Vq5XhrOeTbh/uxi6OE0FoBQbm
2yIgG0bb2+rbDfUymC0Pw2EN2BkFamxTa514VSy1ULdfqPwJ2SzZ8hqPm4LeLSsbGqbjEWJiix9E
9tSSSZbeh+5OORV+WZtM/AlJchus/reA3Y2VxjumqB6JzdEI6Fp7+7QjFY4vi0P0Hfz2siRbFAUK
yMB94cpjPJ3EpZlvoarnGyQlNP9PMRAZ0NN3v9MsI2KZvHTbLPdEtkkOAdWIpybS/VevAQzBOlc7
NtxGmFgPxqxjIuZ9pWtVfHqZoL9fH7SCfcHt1lI6lLQAHCvNDoisW0JE/nSZknwDwTffJJNtChP5
WKVg4a+daG3Pw4zSw9zGKU7oezcjhqIQ9NjzcKpjojAxCY3pLtURkZUx5Jgk2ZZns8RAN8bFtRWX
APgBIpC2i98EYDWyrLn81bBn9tZUUH4k0jk3jdp2I77oWZmQGAU4cisCusUsBDPbmP34DnMM54l7
i2O3Q5chNY8bsizCA9g8OUKqJrtFiEa3TIq7FhsN4DNuPOuf9PUgcwvaa7xvghUt8SswoF1dFGEo
U0s1X1F3CoJzjhUPH+rZ8byOnqhrFWzi/EuuR7eaIcIl5udi7ly1Auu8pPrAqCD0dbXjMtROQhit
biQdrDUDO40Lx9qjhOG0rerAOuRPDP/DVS8X4qF0fapSMvjKSOuRmh8KxA4DNJ3JyEx74wSc3E2b
lmH557ca5JkK/vwW/tl50YMEsOinHLDexXiWU3nxxNyc4ooCIlXjtfGVLatYwfqpOiDnsm4LFLMp
He+48h/vIEMIgZpkwE1qcGq9EGVxJysoNGjR7GoQxUH2khmgMw5+KEHbQUOiN2ZQBfEOmF/dPXNi
Dnu0U0cgI0Xv1QjgCa1c+OvzmKeuU7hTEXX0HfBvha2XbbSgThcVHm3W9vvnuafWAS7lhKQrHau0
NW3SvclcjWnYBzIADzyq4zFSEHrfgi54yoOA63/mSy7kkgaPbOy4A8VDmrnYsN7Tlx2y9wKX/mGW
P1caiEHg/oiUR3NB1Gi2cW1V9VBFlWD2XI701humAKMibaC+gDeJytRz9gUre3FkFUahQoCrHKav
XX0sxbWIcOiB70gqCg2+Ncdw6ioJxlRj/jpe3JcFf4myEEMl5L7ypmW6S+7rkR23J9KxbBvBhlnU
k3kS0tAgrV+O3yDLWl52soJAoahe8vQXI02jJ6nrRorKZYY9TItiguZ3xooilVBbYVYMzBpjH4vt
b/QOo6Zl5zCN1OI9vwEEbST/Mx8MyXEhdDG8pF1/dXUZN7B2J1LCIqs70f+PMFHUEbrkG0nP8ScX
EzzHsT226sNaYePt+DeLyliEN7PeWQYwP/Pk6HV3EaRpyqI+UOhNoLZfJrw4A02C8M7R+UKkC0ph
hVI2IcHFhfwr4mzOVmHvoK1orXEHSIyLN3Y1gOTBGwFLEox8UZenPlgUOwbabvYDzxLtCO2vgO99
HwQQURyBREWFmfwoS2JArXrd6T5FoDoVwrWkp3TmpQkbP48kw/B1in+8RxS6opcLXH7OwH4kw0Se
CQ+al8TlPA9H6UrJO5dZhm71XlqS71mQeaLk+C6l0MQ7WWVZyHC8dPR8skModIzTNsZPMh/FYUh8
EDMuavC75tnKcmIQQWUKtHdVRkLFj9shFVowP7UDR4lCmdj/mJBNtftpf5TdtUTIR+OJCqYd5jN+
J1jhir2fHT+BBxjNdGR2p/yF4IusJvzeCJvt1QL9WKiZXICfmTaUUx+V3Jl+6UToh2YNQGT3DvtC
yy1qIfKetv1GHjmwu7N0wiY13y5EDTDck1sADQqphzazN320XMyVAms3UQZAatBzzLVykMFigy9T
nPV4z3B/UNIiFtybCs6/uBDsMBm5gbEUKbg9XlGJwKqnrgWiVANr3A8CRRcEc8kDLwEy6/RCZSQN
q1ZCOfYt0itZ5dpLZzNU68WVjsZPwKhVQ52xF0Dg0tw7un7+u1D1ilOBQ0aJcIefEBM3sHwAzu6S
znn21gG0kSi+IW+tB+14SYGkyj5+hmkP0Wqj/u2ZKdPn3UAAQkt5DvGZnR02Jx25eId/F0x1xE9W
lRLAX0VXXzc5l9AOeYwmOtQsUl9HPABv5xAMczzfxyPU9M6DmwbcTiXuqCIfbcWZfg8VUEwn3zyZ
A0wmO3NA7MzBb86N8laz9CPa6/yXUy52eyNkYx5I//kzFqcTU5RNTaH4OqhvEdCxY+coIQa1fLz/
6oW+LFtv3ncbkZoO630VGJAZ2SrhIAQ5pB+IihJlnhmIfJzGZdLmkqhHZxWIhPgkkRi/sxYzFurP
Ub8WYfwfbDzRapIfsz6ZW27hswf+PN5k7yx1jL2/NnKFwAyaKCB10pUN/zL0FSPKwSaRZwYVnoyJ
MnORoxF4i0o0ZUDWD8N+hgRSKKa37Uc00QG1LEhDU4qNbDzaldFrI9U8N9rhFps9TghqHlBmYpVX
PIpHDKBd9v7GqZPnJ3N7olMAYlwxeTDt6lKboxMjjOQXmKmi2PjLrp9ZGI+DdJMIXzu//BY4RjHY
YLbbIf7FhoeL24BHqBPNB54V7i+Sjxve0frAKuwn5wt4Ko194w8D2WrtbrDZ4qT9I//r7+bInrIA
jBgFbh0xCe3MnTnoUNYYP7Ynsgtm+hHHk/1JHzb59pDcK09IvyjEkCb48lRByy8s1nYNF8buZw9y
01B+7Fnu9KCBRKDIeJzRpA6lOjDdM+KnaouoxNxfcrZL/R8bFpNyvRmlelgvm0iiFDUfKNbbuRTH
D2aB6dbraiEuti7BqwcQXnbb9+qU9pPQ8V4JbqRdEKqqo8Sx2FeyeqUWh3UNzij+mUxvGmD+d9cF
Q3cu244SniZNXZVSHjTewqNbBmEpT14iE6/9quxRN5gSpQuE968ZMes02WLEfvkNSYjkhsHK/PnA
/flOJS1wjvockd9GFrnaguXoN63nCKcbMzxh1kS3IRnzOEMdn3ZWJ5q7NWFu3SnxtRtaagRRuDyR
PDF6bvNIALpFyl8nLLZ6N6rFcs9uve634Fi96AyHJIvNPPLntZgk8Plcs4+O5tR20FJIdbwUsyZe
NybrZoobo9QuUPpn85q5/XwD7srtp+a8JmJgNEMWd1AIOLZevYKh9X68aXvUY1x/gV05NeAXddvS
tOEBMrwjEsmEVEJHw/iIgvO761r236zESGiQno5/ROuK5UJCa9hDIGDfzePYvhMmmBFClpbSZRkt
auhq/Sv4Sw+8xyx3CVbTjD3AD8ac4A3IXN/OSb3DY9MZanWzImyKIoXRFVv/LNWTDrdVYO1d8nB4
KgelLls978rytbajkKTGFnaWur+hOG8CpQFlpS/GCyAz4vAakBxYo9qSbetINB7HHkHJe4ySNLlB
8ils9wqSnYbrkACMgCP+VTXLdxrzfW+Vhe9eoWns6oJdEuL6+6zJBX/4/uAA2eNxr2QSG3DIyuej
5yGOyhuniGjQkXuhtMzv3Kh1k36g6zl955r/mHKLUo0YHAdan8JsptywNxxSvqytyXOoT5E8dO5g
GIRhEhkYqotrnHQagsmDCmSRA+dp8jnWDcKFM3XOMRU8auegiM9dOZDZCzT8FhL4RtGMGZ2puU5N
gcrzxN0pVUfR8DUmUJ1h8cts+1QjhudlppHoWAkbrEYiMiOOKY/tBgbX0ts2LBAgv6YdteyZMv0q
DDS1CC3n+KVrRVEDuMvfIDzgY/jTyOekhVD6UI47KAnBlJ4nThsMV9qziGb51lIl99vV2IhvSfI1
GzxfXN79YRZC/vkElmoFTs7wJ/ohs82IARn6NDRtKZy7cBdjD7yLuEIsPheDfFWXVw7HEaNGUHX1
VUJ21v9SQh90giiFeSqkDqFUyymMZZo3Qo9F1H2g5L06LqB3Vt7WbbZyQCeQNM4pHLI0jdyooalK
iYGVhBRijBlS3k9gq6B8rpRTjgGl7voERrm+5nxo/y1g0pIdZL+hJPT86PM69rMVNl1gFk/KUj0J
Kb62vh47vROoGBO/t/sK8uyHFhxeMSwzdhY9IncLAoOSh+NNR2rygxwwomV0Vpdir+M6mqEFay1i
wypZ/Tqui5RBJ5tuAytfSzwPzxwVih7nYejZqNAMrOUtkqg18+k7iqIJF/AsCRxLier9zUZy1UMH
FsxCzHNAnlHRJ++35CtIlwtgIN5+lKOAwY8ZGjhUCBkybAukG/gIzDorN0UOcJv3rWWIKznPfRyK
iRNtM2NYWfyJg4fFjaiNAkKsXaRs7JmOvkSMhZvnoJ5BNl92kmu8AHIUNqCWkIBtW5Ko6rFNDajG
rVF2UnYSCEUbJmIumz/AkhcsqezZZi2V8N5cZME82yGvP6qZlo0xO/WPZuY/g/Qb7W3IRY2l454F
wr+Suxx8p1urPp3jobSGlk3BJbmpuqOVD6wqqJ7Z19mA/wa2NXqa7v7kSdO7pYFrCh3VBxVV4caF
TcnvEycsPSCaQTgqQtnB8dlRhrZWmFKqz6XzH/bPyNORfV1yBTn9JpEGy2qaBVRzlBhwKZF90w8r
rqPSDN77CvurNyaC58anjK4nOU94dHo9DXDmwRdmOsmOCulU1WISHggmNXTkP8mNbjVxWkNikoQI
BlSfE+V8UBPNKKzdzY0Eyg9LtRXTRzWAgSTj4/ZBFCRAdgbalom7OFwD6UJdjjm2aReR+O3TuQjJ
7E7TemIg+TRl0K6qW3YjxtLN94VIym2ouQQWYKyy9S7uXSqs6E/CSH4WPdUGFmA9+qjGeVJuKKsz
kGNdW7G8o812GhCiQT9OmJEdgxwCI3FWzyHBkuIG59Rfmlvv6TJjablLssMMS2Fuu7zMBS0u4x8Q
UVQi2Nv4Aa6cnXTpdLtftYHvf+qwKm2mmlzcMMDGnhJMaEGJv/nhKLTFYhd307RpahJogY8/LpCM
HZdm8w63Bfmmhv8B9AAR03F6dOZBYa0YgV31VzfoZ5FmcJFeSh1zV2fFu7DIcl9RJ0Q8nfVv1ep9
/q8y2LgejEJBRM0QX/Eh6M4uau9WUalsd173lXaFB3s966EruonddEZsOkJ6LoJDR6PDrgsKUkVu
sSiXM2bzqCjpDg1y8FBHPRCLkFJ1yh2Nt6L+PRX4CS9P+QhXHvZctVK9j3CwZiEsoozv8fBHlZag
K7YHFt2NVYdSusqGhSnbWH2t0y0Uy4pNWX8vjlrZRsKPc69RJkg7FbSXwFhFGneEQZ0sfxl84LqK
/9UxJhayD04iuhD1PUEXLzCGLvGViV93QSLPaCy6tpN1pwdV5a1V9lmT8pBPyrM3Wc52jRLYNaxa
l0ZOaFzeALDIOZOUIrAmyC8Hc/1iKosRkDRQSYgGFZxpL3VHvks7QGpXGMtad3wCglK598BfhMzO
OxZQ4GqbJmMKmkVLSm2YuGPlNm1voLZ6DKfinlnTp47j/K2qOqWfE9DsY9FmrZ41JP1hZE1aTghh
y8EgEb/wUc5agKJCxHkeoOo3MkG21tdBUo5PkuPTaospASvSHI9MM33c2FsliE01mhBne4C3QkyR
3ALfiVR0ZXb/HNvIYmHvEbSuFNTelYdyLIK0F03a+CfvJv6BOxrGVSLECReQf+ygf8XW0qOcLRKT
pMHom1TLnbT5SRZXTaySVrGHgQon12aKkalvRRKX05rR5NRgOhc5ab6G6m3/+5dCaM9hHBLToftq
fB3R8CoTLrao/c5845K6a0y1OQAS6ZubrPhJayB6Cf3UrwDWHsMJPbA5QA4j7F4pTwCEwj7hmvQy
uqWjTujqtucmoDD7A6KT30MG0ITyPPuX4R6PfVkPkz+WAEXJIYjV9fl6hXc/PkfMHM8LdaSfzr3J
vvHWY5BchZftMC0f72bMXYcwjTioNREeQOEdNBFwJIk1C6Hygo9DD8SvQrefGDxGUXNsXFqfy29K
r1At8h0mz525YKk7lXwC7Cpg5ZaBNMLyPiGP2vpcMw8wyJ9u8RaFEocP5D5QrQuhlM7s6T+5O4Ui
bQfpo309p9XdeItGk/SWggpE4Fo3pKL8To76OTs2YIrifItJwY6sctzRV0YJy7S4aRBG6aF0UYPV
RiKBlqSB1YDy42StLiFfNd7gvksXjP9ZQDxVCb+BYhcp0d0YwSEmKIrHqtL6geeCOomoJl+qR+y/
+0gF67Wepf5sv93K2qtZQFyStnd7vrJ95HGOlnwoQU/C2/KighKMu1PZt20XunpRJRXvIggGXXmI
GiFIG+JlR05XGi9p7bXzM5hjDfAxpIBTB849uxHhtvZQAk4T9zIowrR4OTFAllwXXP0BmWIlJwME
+oEbYNv3QOFb8zrBhJzHluqLbleNYDxNVieehgQ6iPDY1AGt4ZZOo/aTW4dSpfdcuXgk/S6IEG9o
YJA61eJGgB7951YFElmRoDstp2K9W+L/P2R7VY6uqubml2B3SJB0F6X8G8aRUfsIvKGR44zqXo1T
AMJapOIPXxcFAnNBjHTvvNpiHqOqrxwonX723NPjLPvtRTqrWFTolnzU0Fne6n73VclFO0/FBjZa
wVCCrz9bVii17IEjW0zwXa7gAokf9HXeJdEj8To/o02uvscu3Cl7GOZNND4cwKEtAnnZCo3+FSK6
fr18FbRrLjrWnIRpYd2yeuy+FqNH0IgVoLBfv/idD+2zt/I5uZuzLs6+todcUh8COGyWdmo51ri7
38+EPkHxVOpJIcEavtclylaUywPeR+JIbtoHmdFRozZFSy08y9dflkzicYQxCpYDJSSkUKBCJQNU
zuCwxvOsSK/lG/yFCT7Uo33YStBGyIy+fg+oLuHxttetQyFSECEf25NdheGUIH39H5KK/P0rcbKE
kDrcK9iR5jWmJePsA3BCVgqCjBUanJtKl8dcmLziyIyyvcHEGRHPT+88ECq2GT/+jVtjFj3NUVDz
XRwO3ScqzVIme5M9H8VvtBa9a8wbqeccqG+bZtuWiGEUAXnsOUGaowpxV/K+iJrZMLDC8E3XO6Rp
gJ9d3Q9YNMdyetLzBOarL2qqlL3U0KhhuCZOAyNOpqJtcTqEWYDxInGi4oih13du5/6+rE7pnXpe
YUfA2JfPgtXH3bLNgRuURQmt2wjuFbfGOWeQhuL8hMdWEeKgKu4kMMJjyVYz2ZIOHXUKZKTvfmIP
Fmr52bLu4qo+z6w3YUm84oQfyMi965+qloXd7g0osXdSaLCwiBEsioB5ylnf4te6APkgIeRtT27H
iYDVocR1spMoIG8Q8NYXZMX3MpPrsbzbjPHXZgk5Fvmh16cLS5hRhboZCrbgF+Dp6pSoQO3a3twk
AsF4E4ryZzbVuHHYR/QH9D3sthevqMYi5JD1Han38M2ZXXLIdg5C/QYorj7fWe1ND6qEQENxqViR
HfuED+Z3ak8IhLxtDGzGv1IJPJbfiA/IMICXDhGDhrdzNGH6AsvfIO9xuoI0mlVaqrOiWtoPVnSZ
pAp1rQ34S01TN1veGVFinZvmHrktOXTnG7p/CwH61YfPd5RgoF/kHbNOqpJWYApEMLLotiwgA+nJ
gtYW+Y6tRu3TJeGMxOYbEhJiVSzxWZ6ie/8ZdkRdiOsaE/chIK6LKTJlyo96CCJFSwl2eWKx5FXi
9G+Rpuc9jsdwYEhRC2DpBkCe02R8RXyUMT8GOZeINLhDTcY7KvfxAwfmEi12PRzXbacgLcbZVWnI
f9WE3Mli3xKeJChNREs4L31kb8he0hnOVwe7YcQOjn5p1/cbHUkDs/uGrIrnrhlg6aZWb45POfN8
VsxuZAUFTGjC08XjAPnzPEk/HqgRiBFexxoMJExnXBPkCw95imKprNSM7oEA4AF4BymB4mc782+s
ise21lZDXV9VyT9gVnmlCHptiztnQgV6echpyzTrlnewbKqcanYzMTKfL1uh8P83zcY6uwHS4AAX
4BYjj076ZrvwHrnmDuUEVBzFyxEBmQ+11SC7jEuBqieQxXr+XjCNvCqVJQZFxm8tVPetcSMDKR0L
nywJ44acDqM7KpKMLm7jlVjYFNXDwyEHO8feWjfbu8D3/DO+4sAWRvIQF/1jKil6s3yosKvr1wvR
cfrtgy+o23LuYfJLs9t3ron4a4lLapUd0nrN+nmwkAe+ZxofXFKcti4b/lJknrULo9B7k2gKzBkP
pUWFcoPPTWquQJQT9pWlcP9rAgMXUcR9sj7PO5PNtGsZWriCmPaWtCgJF6iHWVKWS2sMBLnqHZpJ
voKZuKFWtxT3kBueY4R2NrkSGAR819fVnCOGUa0c098vMccj2tL19OjBiF1H6qEsFqGGVfBTiRc1
K9pANW7mxZa16rpgO9UqW5+vUFOt404Ssc4pijDdzo6LoljHw3B2VawSV3oHKnNWr7FQIxyiAL20
/oEaciY7pzvgrYVbscNteoMK2AVExccJ4eZBBu62JRMIGdLO0p5jd9p0OvFYIRZaGzpS3J8eeZSh
ypLTNyNNz7ChovV5MRWW+5vMFjbpt3MGE5Jwjb7o//RfSQTKvvbQFKsYeb/V5jK+9B/aJ3nA0MZk
QW0vzGBfzPwDkru1zlFt7G75flZwbwtreT2U8yMDfVyIf66sD1hQT9Lk9OJ97N11QZKoAo0O5ifQ
fqq+OWuWv0o6aUq7Lwsy4sVv9L7jLfm+7T/1OZ+0PLWW30HiTftjMxtYwLlAXO9ZKcKtmO/hrvy+
4oAQH1b6mXKOZhxeku8cc+TK8zxJ5wk+NiMEKcrrKTO8pXpoO2f/nT/UpoA+a+I2T68pnZHh5nzo
Ob9qfOZ+LltFNROD+AmI5lgajH8JIVYRHVYwFRnGSAx2gFAJJTlNlVwArpaOkWvXVQW4WuedIHqR
RmR579uIcFEAhgEg6zv2e1f4HLRurBE/E2TX7106LBA31Ru7c287qmzu+JAGLqZBF4hTzvJ6aaVQ
0y5DlIb8NdtKrsy+ZSmxXbVDSqLxz6kC2eg0NplMnKP19A9JsoqXxXyMj2VeZJsWPk7Q1L/q4OaT
ewvnfVkvhN4QABbffa7wxmq+aIzt3PWQFsyX3j2H+cJLTWCQXYzH6p0KX0Jl+Nmo9aijGRMWJMvz
BUdM9c5p7bLzYK7z23XDbug9REqUbdh0yV1aCBTF3NM1AmvswPVYzUYnB+Wrg24OP1gySj8VmcLI
K+RH/Gupe6hCQWKVqo31ZizvDZcE5MpJn9uj1SX4AkMsLNaKM+n/cF7heIJ9vacKlzn1E1u+Ydea
3aDhuWDwiXF1AKfd4S18Sl/Pf1ZDpibBQCa+VQhquYGZXMZlcauEKlSBM8tvhmJ3CH+6U8D6+4QB
iL+FuofvDdNMMqNy8k/KAfY6DydtHK/s3tr9kf5EHOQSZYKwxP0tZa87bIfTQgUvwlWVYHDmHM9x
qCRbm+XhQHeE+dMoG7FsmJd8dXhO89gkZ4W/LJBAO/awZU0OqdfkFZ93Ou7UVWHEQx/vWtSMVnuk
iwVhoCAXkpBkpJjI/Xqznd8vkiFz2hotj0X5N0rRKSTFlPotvEPW8rNO4eoRjP5QjS9vVD9bhopn
1l3+6LhT6qE+JZIuUDQixcKbEkXsFZatw0b5T4UEaaQkF4Nsv0uiJAWEwR0B6S26onuPg2lRH1nH
LSJ2pFAhjxBFQjWQoGs/REUP5u/NjK3gMz7m37szeJC79U+MmlYICNhmKy8IkLzcx93CJMRzIQ3I
3eo6jWq5M50VaF3Ku4pPJseGCorV7LE8HUZ4roNh+fbsbZC7eRQCuyQQAkcKNC/MTFFq2+5PSAvO
W8oo/NP8oZwLqfw9b6S+pAve8TQ4HP8F5kUIW4NhcwZArNMgSMeU1yf9eCI5aBcuh+eHBe0YnGyG
+u1jDJhAbiua/8+QZOPZV+L7y6xAtT6PX697ZZ2+rKs4KB2I/kav3c77G0zgVHw4fQCG8qRF2SXQ
ZG2ak6Z4eakDdmwtq3ne/6jakX/2oMUIFE9b2GMvVu0NZt8xRvkJo4IVVaqJk4QwFabsOBuFj1v2
vW874v7BVXq/vGW3p5Sty6Aa1YOJ90pRfowgSkQWcucp/hhY5kChtawcaAYO0R+42CdLcV0s6rC+
kI8cJlUdnUx3PGHJKErqDYP2k1+oZOPjlOA5keqRMwH+PLsrbKYKqQtFxvtg/C3+b1NLAIHCeG77
uic9cBD8ohkiD6KM2fSNI6cGWL+KtuZwQQ0pqPsZU/In2JhFv60rR/KVupk6MWw0tT7eq101uxn7
C6CE10l4/xmg2yebD1mTDr4IKammIJ6ixLQV5AIrk8UKn2DDIRopdm7o8/iK7BvoRrMUltycMNey
icB7BGGNakBxKu23PpujxkRyuWLGZyHMs1tA6gi9hsATKAsznKnPS8O/ysO8kOCevU51PGXPujho
+eTatzbuRPnsua+5WPPydRyNY2exJ/0WiFhuAdxBe/0i8zPsGDXJni3duuR5AvGxIm1/GX86wDi/
KANuhK4cg/Hg3uLfTDlzxsIQf+bDWGP0kwdOGBW1fMgIJMTCqeO3++UIjc+CdVXV3gHVAd5Ek9cR
s9n9fZ5Zm1lzs6a5PBOiVaxirgsM9Is/1csvwc5Kejjb4OkD0BTaxfb4NEHBiiXcXL6CH4zLzPNK
tTajCpacvBtBGvp3w4Ip2MnjH4ZVFRzk9nnBPQVPFl3L1509uLu3VQb5CZqbVQ690eHnCOHnZo2Y
fkv97BTBgrPSkVn0FxDWWAypdzLJRmZXh4OxeGGYpa82+/Bso2F3Rx4F/frPFK+n/ynZUWXQY/2U
AjB1/3yZ4Opn9HdFvgOD41pX+vCPMhRNED9hwmX72yRa4rT94fmrLvvJEuKSramkJH2DcYEBmp2p
Rc8wujaHxcW4/JBRWzmtPDUlZ6MMHJT6PClq3Ji59FM8SkjZMigFxnhAwB6IYmFxdLhS9spWYDk7
4zKCakOH9lfnEATvHEyH72kvpXesWlIIUiULtTt04kSM6iGObIo0R8JsNaqshLM37iX3PHr1Bs0g
iXF6QgYnO1ckeIt2DW+aNtA6c1SewXwMa/mjh5pTw6jbXgVn7T8Fv6lta9BdR334Z8IuZH4vMfOf
0HaaD40Wco4M3EtLPSpgx6Z6U+XjsQuVoXFvoQk+MW/OaYZlpNfzMQ5OOkhXe6ew445R7TCUEB+G
FNuK1+1N1oZlgV9tp0rBxsjvQDuKZYvKrJho5Ip2nlz76BBmk5dkH1ySFX2NVPjqQQ4eo2J8WsHh
6HGsyPy9z2SH20gDyzasQg9vNX57sMi+cVU8qe8oA75WWuARmlLtqiB4xFB3XTkpTqav2Kf8pBEI
PWbV/z1s9TnL5i+7Z8WZuDsZLC/Qu3X4y1mjCsKUG3qWvaFW3ScevTUVMSC7JL3JBQ5s+gH4lUEh
e5fb+fAbwsN5EcQplN0CGfq8PqF/L7f61/bHhZE/rEGKfd3dC8M99FsXFh3ofJn59s2FVXVvlZYm
MFqv0sy05VI+7beKawduVTkWicwJlGefaX6rEl3hspBrnhRpsIcazoWMyig01RwJ8YDmM5NehnXA
zJVhf82aAgRdblxWYgcjEHr6UNRj/IUfN+Hdg5WcuWucxC9gW5t2h687HrFC5bgMiE/zsH9Th6Ff
Y8d38HwxidCXfnK+HPjq6XmoeztA9rkVw+KIB8x4z31efd/qEiyA4KTxcRUGq2JR/rmbUmL6vbhH
G6J98/S4udizZD4TNwDObdEciCmEO10ApJKUZIG7fXRArHknUC4sVKGvnD3cYf1Xd5FVJ9SjtR9k
81kzVUV1ERWKEdJaQMTEfKhFqfO9A5VjOO78yshDfsj8GU+7hZv0p9HMRJH4DcYzvQo3jupE2BiH
fCoo4YTcaEoHWYi20Eh9coFFVdCh2kcnHBMoWqBZYqibJ2nNQ8nDjJOP+eOKOWnC+22ns/gEM4NN
rlM4jA19vZccBjfvHDHwjeeRmqjtAOo1zB6zxvsTeNj7wgHXl/P3257YnND2pGRnf1wefinHOa0X
y3R5mitqNjkcBhFhrzYZuFyR/l3KErEPJhNOxzTZrOb5PAQJCM78KhKRwih8VQRkqvIRmxmycrW1
BrbRUxNqzDb3tuF0MPd0PUWUQMRrl+0D+rkSsYMfl31QXSRCNejJMIt7k1tTRBv2KEiua+duvYL5
JtceazXBUviEsbOb9H/SeWi7fqruM3CnZnCWRaNCJtgolfIL+hbp4NllUKlOWu5y+b4cOWJmg/Kt
mF6CUOwOaoQTGJhlJ9Kw8JlpEAPwqQ46paWCLe2KBSUUsbajxwt0TwRQ1vaoqZOEgVWqPBelKIcc
cg7x5F70wohQ4U/WfrXQFbySS+zdO6WKL/FWituWkYT9hLY56z7GZYkoU/i1DZo14fDuzfHtMhom
rx2VlWhBIJzj2xnXrngzQcecP4Io4uS7hvu6r2aEyXbyh70E+Nuc3C1ZN2e0/3WSOoAES/TG8qSm
exON4gNLZ9l5irm4vsedfV7unwqYY6zjqEkNv4V6g7oIxm5fJrpHIomOK35Y3ib9bcLfkN7QfoxR
CrpY+XPg5g4Pr2wsFVOAf11ntREnawOIhBc1u/jPwusm/846vSdR/Cx/+BbnLKCwaqCNRmhRos7d
HggCfLeHk71QnbI6Pblr3LqA8pycHxAbIaPGEmiJd6+tvyCTQO1MYsgfFrHvDTJwuGpM0kF/YXhi
TWt3bHVi0rwiLh3qfWcuYkGmS2koLzMAev+tRv180NnUoVqILCFgsy2CkF7z4GJ6Whxlh9ccfRzB
eh5PwmeR02jRSo10+JR4W+BLwgvYoJgYd0DMKm0M6lXTdDzzs540WZvjJngNwWBWdZBlhRWNCi4p
vN6P2/1pZi3gvpceKvJC9R8cB2OT5rCWqT6NGUuhwh0G6MSBGFgDeqGQsK46jEkXXTlTmL+nZhzD
uo+UV15qZHUFYd7ofGRu7tkaQNF7ly8MMm2eWkQDboiLTTNQsd0U+AeHd6sxuVVX7oxNU3gQwSHM
o6u4F3wtwZrjKsuKwolByvX2KtDtoIPz4wcNWtj5CQTzBwAnuTh7WXWDv4kOChiNNuKKx2SAjDjf
LHk+5mJn3d6FPm5ygrOIXJEDPqDHr7UwheE8TKpZ/hyhEIc2Cesd7FkLLtvmr+HODV1mTfndgYox
5sFUqluUMfQGuzEv0ReKUxyo+4UObsIe8KIO9Mc3qEeq4dr6nE6Q5y98qtyzNFS8/yL42+ateCcW
Nu3UoquEFFoEdgo8/U4CfP/OTEwazoW9vF9C94pdn0jjE7UQbKzkAA/21+WMrh1gbQv7ewGZrXqG
cdBtMrx5h33ggxPjKU8gyZqm5OsZxXzWfnZPwHr9X6Jr1tZBCvPXV7b1YAaUaAyVBPg3e63nrWnC
pqNY4z1NBAu+Z3HA0vVX9p6cS2LmWZ/FRefA1y57pNcXMHP6sMIRzm20iUATShdExtwYm6uieDj9
c9DvPDqRAuBVuN0tS2TkGT1V/1o/n0YUu+x4+zLxrYHYy22nDRhrVDkqF/Iy1YHBNUCgwf8LinV/
k0j5oI2SRbVRYUKgbJHRNRpa5AOdRYHmBjNYegovwzdrjRsbcaMlIbXwtq95fowv7G1ZTN9LdK4C
49h9AvGQrIAKx30qBnJGx+bkjAS46rR8hqWhxA7zHNQa3lhl4YvOUgSvV9mwHTINKt5dfZ9F32nD
Ilcf0o9lPbQX5Gs7vqQVoaRDT/2261/6/GT11FiobjeqD3EHCbRknxgGdLJ2E/hyyI5xyb5WWx0f
jmPizoUTIMSFv+TleHx23wocl6aW2bPRy657jCRwjGZARdU2623FhC0migi1Mc/c40lEH4zSKtdR
irad55pbW54tAgIS752MhErR910FIbdGS6wytOBIqhVGQ0nBog7t4SWr3cVPOq0xJ03l7/7oYG29
sY57LeUvXuGeLaEPF0JuERdSdTXt0Q0JPxQfIz4JZq3SF6cOt2WA8reuFP4eMUx40APe/vpqgwuK
Ry9eSxFYOjNQUEzrO7Emb0u+suEM9FwAH5c4gCWQrGI2PClK0EV9sZaGaFJoTLp87uGiI9/uTTal
nlTQyRF1CRYfjP/OnZcJ7nG8BKYf2juHj8fnpNfQam3JG3l/NH1IODTJKQzJxlD7oNpI4Bdj13JA
Sfdw2/z50+BP1T1YbOIq0XH4hLX3A1VUbVTR1aMrpGDTvoGwjUPllHDwvlEuZ4UYPX/EMbYovfMT
aKMrTQnS7pIxG3Ep+5cc1zR+mkD7EqBaF1+1D1LeRPIRe6nILaGvT1Tt2/87PVsTxNm3BF6Hxpg/
761dgGo+bTq0piqKz4vFChtxBBM28AjEvJGigV1lvuIjS2pkiQwU5CCnInrU32ym2jn8aaYl5+Es
TVYAxPepcd4CJlJcXfmA/IxElXYZMjx2IS8DXTEiRws4P/2Ps9PY8Y0uBQ+F3FLaR65/YYDl8Jrq
HR3cNhsnt0NCWKSPQfjbat7pclSrjPjnBMxBEzMXLQoACT62C80NFfzI4+aaiB892LAa7lzDFcmJ
mu/M/78Z5WyfVx5XY1YMjWtD1txtIz4XMgIy4YmiWT6zG0KgYdgg+gGAsppbl49ix9qyhzuTAjRm
tx+A7tVDUSspxegbAQ/sHJodsk5IJt6subWnRNZVmhva1fCEx/kFpRGTwp/xfu40BkXtPyeKPvP7
vEGVARWnXg3k2V8Fnkl9x0okZ4vO0kG3jsjoP1GBFezVvXlnzQaNPZQd/nsbRa5q4X8tf0jVYmqO
Q7WY+ys4lYmaQKsU4STLM0RCUBGhvrp/2GmyABGTyejPAoMhIX42yET2cqjL5yEXJHqq4Hs1QY8L
E/LOwMTpPEeBa976Pli/I75a4Jl7aq/Dd542GLA3nVu7hg8yyXxII2XpHmnPNoUO54pmtqAmGJNF
QeqfjnX5nW/SPL4dgdvYVJbOBrSoQYZHxOiTL8/zjrNicYqM3PLeOmz1AbgtSnE3S9XTQ0xDhEPO
9ntZVpBdH338i8b7A1OBdPBtdh30VmzQ/39m8mdJUHmPAAvozWFBK+ft+gVEX35XTkwTagxClV/G
sMK3fFpw6la1+8CKm85FiNu8ycBlP6jA9dXVUFrtiB5w3cbznHXHDKGCap9klQEun2qN1k31aRLY
8sjdpKrTOW5qGmGcU04Z+svMuYUerOy9L2YhK7pSngSNFwr5lOBJ8c9yPGiVkpRWyGNp9TlwnRAk
KpZKXP+bslOeVMAnWqR2yyx7f5zU7z21mq0MGWfzwazaq+/dzzmrC/TKDd+018DFDxdhj1XPsiZo
TKQeiakIFdHKBG9lqFuRD/FmtrkCgwFg0c9IzO69ULawP9/KrdARs4sdBk1yp59QROYxDW2eqPt+
8hrbkvficoEtjKEVR9wPR57RSlTtUC2/vjE7EWL3Ew32vmR0gFyrcekG5IgtQ+gNA5NsCCKpHqtE
dG05G/n85REs737/idMzjncchxqphPajlm1Kq6L67JbBAvsRfj0KehpebSSjlXR735wLQc6Vt7+R
Nn/37qiHhzDKwXUuJ4bzCAc4bS2/H0Ksc0crn0RCKHlrDXQ+e3A7NpRhci3meKB2H2erLRSCGHrS
EaoG2dbE1OuRi9ONbPl48mzjxXueJCKB+nG9A3bq2tnzm867XHqIyNzqJRW6/ejd4kxeOW5G5t6h
0UUtm2TIIUScD4Cj240LvwNTggRrl60IkLECAe+BcUMxOwhjcIq3PNm56SvJ+gNCGFoFZ99o0iJj
qr1TLxLFG45UaGKFOceD/lNpJMiZ5ufMSeSHmLU7N0K/RYwn7keNU4NXqR/J9S1TDtYXX33QWdG0
XBkk+nnBYze9o7dY0PZ/PWG+LoZ03vzwrackzV+I/1ZVtSASJ1lB3737y2zXEDz+Lnp0+glSyx6D
jP92d/WgsMSEu9wwoJOHXiJO8tDiQFvTh1gyuFkd99l+2kvXCppwixnWS3UUXvBqptEOztSeCqo+
aGQY4CoHZiXhfUfRPXIYwiW4Q0jz44AP5YhZfiOG/ALujQmXc139H4u3/QjWi09yAZGfhCD3+9lE
Z9bRS16hPKBnsGN8q5gbX2xY3BWD7lSDONtHcCiTht0GZMSHIsizhWUKuhdXXaJUyjoUmbKCQ57i
x0q/0LkC12tOLt7z7U1nsGqoSCiJE/t2UWl/WzoabrmUYa7w0VaejiquF8vV3XO4IyMFqr0ohfh8
K7GRyWutRG9eyevxrN78XY0ttrS2HYmdDA4gzhp+ulfbY0UVVT0m4286tcKbF8zSIqP4Isbad/5E
IZIldOcdnSooBQYySOswrC14K1VAGfICgkW84r96sDfqC2iMbF2sNkvkQGE8ZuCcGQin7cM6yTHA
fcI3sySR5WOBIDBQjLksEUdeQnWyf/cM5GX0o4bjTzUsGEeEtwfLm35vyNu+HF72FYQFKI57Bbp2
+PayoSoU+eC0MIPpMdeqdk/M36GWNilofNDVoOvKR+YNxS8k12w4RMomOraHsLLNKkdTCXQO7byk
mEugq90w/vS7mIyedEmSrZ7AGeNjwBT7f2atVb/CJapRZD/UVwIvLZPdiwmTkY+Q+7RQXvsoDnWh
s8yyopwNNmXAGVOeMKxsc7+lz1b85KFPAFp5EFQVAWT1YaQazewsi+TMySTrBXQdSfTCHS8AZlFU
bzkC2iW23O/Z0iZ53t903EuS7HBja4Y53KQpMAJLLDSxVutc/HMdsp7syluM4afEHOeRfMD/2mm2
oM9ks6kpNlGnRM5dM1xr+vLLi7HztJsgdr4U32qS2M+uOoxpgGVayQS6KDPpUrZLEFed7hKziQtk
NWS9jBaTkOTCS0LEOjVLgCBICTMMPUbu7iDJVoDGPczAUpMncApQ0UPOl0js4qIuBKGDpXo1/nsX
rReC4bqnQAdndGt0znhxN8LgB60ryfQgsTJxx42XJ7cKgB2CLqSC9Ufv/e2hjxyYpVqt4slF4xvQ
R+vs1cy5VbtdY7hzLmPukgtglR5G4X+PtVOXkz5UBujaJ/K0f43iVq+ebPls46QqlZ7T1QRa2TUm
sRJ9+dydbdCT3WGkm1sKG1WaPkavo72/s2ifWfcXW89ZooizLE6J4ShYO29aqcPEtBLJsOf/WX99
4HYWrZ/MF74w3pYuhHDtjgFnry2ZY9JMUl6u9dJcBPq1S569+SGWBeUvMskOXUAZDIXWEYe2T8zl
ZnI6C+MeL/enflg9K1dKYegEMbrBi5j/ZQomEtaQziuF/hRXo/vgmllWqadzHrgj9d1pqv6rvSAr
DpfpyhllN52RWK2QCqUP4r6zCkgUwCnTi7yeooQ1ljnr4LMTrrbQ7oc4iuNagL3pxYSyHUhTI96N
gGzaCusIiNirsv7XOFdJ+Ylh4xGbhHAQMEfQxyMXndF2aNm1Elt3ZDW/kg3nTeuzPw057nogsNzX
COugAnAbQblf0jXueovTb7Uh2BGwvA36ySJEDZdA4r2u8KQB/u1+ZX8xdoShrNy9+7VR5qIgpx3+
iagRK6LQdK1EicmK91ez1s1v/s3szcei5+Lz/cOKSFGVuPDC2eKfI3n2jJwPaMzIwZqByTpRhc78
fyj95w3gD72pHJUDyyXtpjfCAdSxVQ++3AkV31wxBR3pG8RWpYBJtfI6gDPpg5h86dP54jhxfbBX
VsrsKNPqlra1XpSqowuym+jMavIgaS+zD+NjrH+O1X5AvR6s8gpcQaCh3uTfpw7rTQ0D27AMiBph
4+dp/0PxWxG1bhmYmEve1njTUpN370USLlVwU3ela9iVlpbmt3L2H8oqCdYO9dcbiq7ggpvipY4x
8K2XKc7r5vYLGOUQde991IRsdzQXcD+mwjvWnqFLJOswBvc+81n9e4PnViJzfEPBKPWdYCDWQIEq
l2aY/w+vhOd9f0IQprsVYTwWSRVPeZSAeCDcFak472UpOqhg7VIUU61fPlws6fgBmhwNADZeuoym
/2KyciN4eACVHDre3JoVdV00rDb/RNMCm5aR07OzOeLQZsf2aAimsHqSdsN82v4AVPnwABnKdg9P
D24pbcHPRVH7YLwRCizsGvWovn5OUtFKoSKrQYIo54H7z1eCIokx4Q94cMOJAnpraOf4XoHEye2v
BLCTgNLPlZJ7ku81w/eUBmSrBHHhqggyUlrKf49/Fr8X9A/05tJFRo03BugG9SBiAqFd3FgMRgOL
KeQnkOQ2FctodxMdtUMcbxPxG78GoB0GZuTgD9k/p0NhsMgpPiWDT4riizzipnf+A2e261bUDwnv
qv/KuFerYCsMXIFmmlwHCKmrYa66Ps5NaGOwAONskE6aGQkTOdEFFxX5Or85P2zudnyTVa5CuuRO
OLqHtTLi/SjmRTUwxcRRmB6uGsqCGqYdKIC7BNIKsBiixzHf2GEl6FJovVmcg2CRDXaVj2+Lrit8
N+00FzGtIbhaH56oPDqBBxQfS6ie3cM7Ge9gCmpDhWAz7g/d14XKn55/l81a7VaTK+im2MVPkLrm
TeKQDWocmzFPMi0Aa8H2Xm+o+nWsPWzWpDooy7ApDdDvfhJ2cnTjP1U2dQnUR1+FwRZgsv4Uk7ki
lrQpf3Jgh1Ee2dks9wPHpl93no8rETLChsIt3d2UtahRiFd7kOg/RlQsdgxjFMYEeVU8Hr3fHEjZ
E/vbrI83TSfANuuMA37C2HRkgIX1+aqqKW73UwSWrftmIfLvwrlXJtY9x2228rKCqBlzcK2YXxLf
+jNDZzpNwoWUaktCWSYTVsZGq+V2rJwhgVtP5/F/k9zKVAJOK6x+3z4SEjiA3SmJbbrs1qjwS42H
sHlT79fQyuiTKCSC952v67HGuUe5SoGTTRvufkrwL9qnjfc9NkBUjmm4AngUWewEFiODSpyEtzIR
89E99Ok5839yH8oskGjfqWcnioV8ZB3/s4z9SN8FlL+4z3UiAyFaJ4PVeaFIY33TOUgCKWVuaxCZ
CBBBalEkT2Qmcycfp6R0mah1foY91A3xU/FjVnv1xaISIz0DCQcAjZrgTKLXEQQWpyLYo38HmOmA
mPV+HHBL1Du7WzQyLtFLxBntb968x+/+YrDD/1X9/hqL3pSAfSqnM0XDpGaZL4hrpcQFOLpyRUI/
hrkMKiKtFeatRIg9QCbYejiH0gHXqd0lYIdHFZVMJ0Xo6BjXclzM1jmsHEhm+FGmBW4AcVhX0EQU
pbYvli/Fe13cvwtgqN8O21pW0TeYIjBl4UzJD3P7jpuwlz+zEsckZV3uYNVwyw/Hne8mxLr238Pl
9GgpO4A2Bn4B9MmRRgYxr1t7AGiyX8yLNmT00s0UBzgfqZ/6FGpxFmFBQiT451uHGCuCZWz2AP1N
Vy5EMYu5uX1aCNG9ksLp6BidbYWj/pu7RM0RM8oID+9gI3sCBTCHYZxxRmGK37gNiJ8OiGLXh+vF
tUbfIyXqFQZaOa4IorY3cngteuwTf/NjCnzjg6YKh3feOky66E2cKSYXxBhkapxlKc0W1mnojlFi
Yaa7c6WbEzxrC0FhccS+NDIGJmJIFFnxLAeoIQNbVhuJCvHiIM9EUkxSbbx1WrEUSGGG9zDAEc6n
IdWwHfwbXmihgRXLvDT5HId5WLwYR6O6YA7OLPL9ybn3lECCr4GDSbZY7Oa/ByhpCFgP+mzJtpwG
qX7l29TeANtcPitXUV3rZUgTqC1Clz1fipQ8TgN8TIOYT+oCyxNloIF+TTKKoZbQ0SZGmSsYqi+K
pjnHHaXFTJECwrNK9Z0Zda0hVFg0Ry+3hKLp6UuB/ehPRHjIjnA/Im5kcNB3ip1v62zqGNVGx1X5
BWMPnrrgjdumVgVxzpYPTyTSxJOYXz2Qa2JnOmeu9ViKzgrxX034R6NBxZqsWexl/VNpuEMDvQeS
20FlU8ifK6qUv2tOHrwejJ5NeZBolaOnKwR1XkXB1BZvR6oILCcOlTvAL6okoAEcxDuPB986UQJq
UIZVDtfv5MwgzemrGEYyAOnAqRnnOGu09W851l/kVdSxAV8uzwSV6nr+iHt2ROHAxJUFJiHiJlmr
WIAjYk9NXcgsrE5BGeDiqd8hMZZRSrPyo67X1Y3Tijsse5Q7oH6Vyra8XqogN1aAR9UlM5Wks09L
Vssea8iZNvaft7sLfimaPA9+p7xURMCBDe2aOwJoSMjIKoG7CG1fxjgF+2goQHf+AVn40xdnoATH
V3tKuVuG62cxAcKkyFiMrllBGsmiUY+IoH6U/13SO4HdCc9E7ntDqBjpA9uvkYLml1P9NPY4dV9D
UicETFsKODJ6H7uPpLFr00jJl9xjsrsS/T5vd5jwof3z3tuozAc7/ZquYPHLHygwq7VxrCInOMUL
vgLs5GxdpPE9VYRptiC1haJLdnVRTK0B40HoBbqfLu//KWk3KLFEg5NiL3T57Ef0rPh7Huni2Khk
EiIcvGURdAXM3Abou4GInxFygRl+B9BRYD9KGS7udFiif7dtAihKWug8xZgka3qdAwS9N8xuDr3D
zBqRy3yc3JCYxg0t/Uu29YLWuDGs/B0Jx1Al0uLPmQuygSBbygxuIE2zJU/K4C5D1i6bW1ZIKBIs
+DYNcnfFcgSGHYPFJnqDQ/jdpVhV9gQoX6YvPmlW9O9V8hTesLkUplkHm0ntfvYT8DblFC3/4Fo8
jtNlsHDdT4ZEYYQK6gdDPwAhfYVvaCJeYbIliUU2VOB0QD8NyeJyTXBooT/dKRAlglbuwJKQq5iC
p58jdgPpVLDHAtODweEThNSdk3EOotmlb0EDtOcLUNh++rT5ht/XI5ifCb/gEDkUCAOFOFiAmxmy
yZHWqVYeSR4ENpo67Uj1XPwsGDcpoTeScBSuBlGaIwJbBMHQbkszJR+qQyUM3arVnfCkeUVopWzt
kjI2dyoVvOawpmkgwVqaiL0194vBLfhAk399+fcSkYO+hY/e2edhozAn52xqG62RneDpqpiy2wRO
kNQ6t/aLHbrtz1YFs4IqAb9CQG2JTutBgh1z4m6rHLb94GYiM1iYd8JX/dUbDvfuJLUxtdOoAOBm
D6Dpr+A+7QZSORPbe6UufUfG7+JfvyXSsvFFM3D/ULGflOlPsgU0avxWQe1dFPq3vvhA63SdB+5M
8cS/hh+TChXDqLzd7dxq3jl/RG48ms+OzaD1NSLhMhFZgBonxFt6vl/nttLjMzSVnNwDdZZJAFg7
Ib8TM13ltu8tMuTqFtm0Zg8jk3xuZubNWiBk/cH/VTVX9cZddxpinbAQQNzTRDR91xZDg6xu6rm8
H3NodnLARx8oIIjXlAeBKxKaD8IVA0PBXQpyj6XNVyys/1LvpIsofHaszUglJ5QDsNAFYLWwvNIG
9VSXTikCpmPsuSpytn0F6xIkIhFA6TzxLTq71MmltOTC61B9ilz3lduv01B+L5CxIGuNn6+YsaZC
g4aWrfmklc4OuN9wSwyXHTnfLhCfGTN8I1Fq/HW0f6N5PJim8JWN0XZ1+Gp7/Qb/KoFPxhcXvqh1
m5c/SS3XR/e82RWytBFVTajzLEnzrXVuFX15WzqXQZVSF7Me5UOo0ilS6SNGT1lofRSkHA+ggE+c
tFNx7D3b/k4omKY/eUyc2ZBN0roT+MSIWSIiFyn5EuvD4+1pGLF+0OKzJSfRxCN1YGMRtuuBv/IZ
WbEd8Ernd0ZHWiAEuyThRUV0bnYsH9fAWo4n0qJQ1bCVHdhnZBnceWgIqUfccPINrh/ePBkXI9V3
OZTSGrlyyBHig0OOncqlqU19eSqqQGV8zNyqAo9vupey3y5g94CeB2wGgaSERO58VA4BMs0cT3fA
/Rkzhg6vUYCgrM0iI1agVo/+aSysKzi/jy8zGxTIGz5v3ajwmdhqhNZtLxJL0gJeXlTlD4QtcbHZ
GJsgX7YkGHbmhA7neTcdx3A9osF34neUZKXYqcNqBPR5UnMu8J2TyUYa5VDd6MLEQyodkN+K6RUW
qkkQ2usjMuQLZS+la3KxweIvi2aLlpo3VRkgxapGT5ZwP0w7odUh0swA7yo1vaYrIRX45LDDrh7/
s+7z3cmR+mBjT/j3R3OpI2PEP13WbU9D8pua4nbmMFrWAMCVYzgKEWwjRnj3CYVyU7pRAuYTOgMY
iopFkjy+cI1nIBsQyLwU+Ujv6H5u+UWITOsznkfq7iroRAtl7eDBheMWayERdOJm//jqrws4Rf07
PdWiKJtJy97FsmaU19Q7VSyhe2ikWM75weUvITHPKp+GQeykhUb8HJWlDukzhj2vcsLhasS8ctYn
nQVmDF22S3iOmgIeJMoDis1fRCiRJWtFoxnwDjICpRgQeJ9hWl44et+X62UF4uBNPKHS69pxLDJ/
KItke48UElS0ds9O8OTGtbJjyWuiMre1hcSKXdZC5Aa1/usjnNvg64gyPha5av/Zr3U7jkta7hFf
qp56G5hsaVqZ6V7v0pxOJbg6xvh4Vrlw4vturnYiRNB1eRrHk/TwTO7vJTSIG+ovW3mS8FcXpYX6
3WDAswc8bgmnXt/mb7rWttnMaZX7CfhDeJHJZKkdOpzz+m5+ph2sPanR21M5jy2nab6jboC9CMxi
fdq04kSCo4i22Ud1y+dUuD2xLcNW6tOx+/w+gZGDiy5Wt1HdmsG/0a4zHo5gt/PAvqD676UeQ3vr
odrime9VcvXe25gnImEi5hHfIkVtzJUqkj/TGLjhrv5EKLs4EHVE53/8zLwdVRnzqz9qBwvgbs5M
CcAo5VJCSsKZGAtUzQ5tx3KiEtgquzhyajn2SPQXijkSKMy/tnW+9l+zhFo9T8dZ+KgeywuW1uqF
S21byPdabNKhaoLRw2PAWr+vk62xDhgZ5CHMuXALEKyrzzWkBub5cIX9MgXqz5k9j6WOOOUzqQLR
kgYJgvoM4X7bJQoKCZg5SvBCqIdycCZPFH9D8ezTurOqJ22m22WzWkV1AUXQvTTxKcU4GqMHq2w7
l1gsk3sL8C7tsw7JgScKnLWg2aZKgG1slT5lAyyqeqf/HjLWA3mDcSHjvJ8cbncbjVoxMTrgkJME
SfiuAeFYAUoEZCNKI6EXtZohL4MPsWYQW+pFoiruoCxYIOM2hgV1fDin11nY8gyojXyRS0qAE4q8
WaqeclETMH57oIPxF3VKR5A2r5kM0xKZTmUZ5Dh2r33FUJhgNJjcZaahevXSpp2aFSNeiuRf616t
LO8qdNgGTPL4yeop0a8x4WN9y6x8SDu/JYo4Iejj9oPpPSqRnrEvN9SuYBMdUL9fgl1SEDqd/L4C
8vwEJCuFLr0OpqkN7zkUDXO7baozON6ktPc3WeaKtUtQiH4niqZjyPu5i4eZq825ThT1XYGRv9Gp
3MUUL1Rn+soG9Mh5G4w4ZkhxXvGi+jCD7CWQqunyLtZrZbe8OBSwtS2OY5yPRfM7+uShLd3RgkaJ
bnLEy6yDsvgL6aDdezsf2A0rlG+4YicXRKjjgWtEhff0vLBKCE3Sd06CHsqTBlyw98aIieUSZ0ti
7K28lCm+eDgX1hXLG0IN62UtHUGlI0VQqhulVMyo2MvPGyD78Y6cfxDN9YwWYbZZycGUFAptqToE
3/B4LMMHiVNB5XxEBLiUkHjOdRPzCl5nfdn8YjnBpssJlGO1iLnqdAmQQYxSdIg67TXUbrcb9BsQ
XBQQsCXYs5AAs/rdyPv3xe6P3hoKvD+dnczaWYliTi0NqQrNqoi8K2Mag9PYxVE2S7mXGFoEs01I
ty3r+CbqXsPQpDDmLrCg/lwIekQ+zlHb7/1dnCKvs5kpjxQ7km82dOVcYyf7q1gqmahwXBdLe+o3
1tH/Z3FIDciQcV/wVV2vH2JGXwqbw4AeaMzQgVTGcdpJdfTtDSSJSTP1c0xnz6RYR2Ffv4owQK8/
8Q2DSt3p7Pn4X1iCqlQLx1TAMMcZSCLiBIMSIU/82CnxfcCXRyzUUFIhRSG/+uwIpreC5sGisCwx
Djl2dRl0P1wD/8Hd6ibA6Ermq7kLwamm4OhaBXpFNB8Rli1e38tDoR1JQsavx3x2J5F8Koi9Gzdd
KC0lPsJjXNRsC1kC2WhPAttFwkGNG6SacbVEv121Wz9ar+i5O28eCodackDIP7W+EgRmDBbazPOo
9/pxBqEk/I5kzrjZny/4dgozvUT0gX6dAjeZ4et0cWxho1DRG7WUiTQIXO+oewWqlIpBOpIVgUU/
0LwhVKwIMtn8p0Fbn7bDAGxJO9TMXu+5yH1fjAEwsQyXqotHalFXIzmXBX0j73ScZx+O4BfjrX12
f/UGJc4eHKmN0h6/oCUJDpVRRCmiUwCU7G0IfbqDvxF/oHwEhpG/xKdyvlVAe0/SpgJPLX2WJbFD
W0EtZyJ93A1oCyIAwakIJ34xBuJmbIAZo1KNpR0O7DphKgJHdoO1TQGWZnJU+oblrPfMp7vA7XC/
bQZqhLeZtWn56izWxChOF9lEz2We6VprVJTBb52SL1N/46/sYeDe1a8lXx2qhCcfGUe97Tn4PVTe
iZhyukj88ZFS2GtZtUM11lJxKkJGEqsUz+585vCBx5eat4U+FocfBbIYDITQNA9oJkhobwQB5qPA
b9EXP8lgFjeeM9d0L0VcgzMEmZo8JLJpomcmFM9gMmvRUPdY/PJy/fQ5OxlARrkrtQYPgYG788sa
deyCZNhTEH0FDhfBmmQ5yclXuNyUmMvMYJtr/cHAFZM7o2n+EFiFjL+An2jp3qPs1/w3iYYuLzDX
hdu/ZEYzFYv/AJHCU99AAa+y+o4/4HpqIWGsUokw6sdss7Bu+E9MSkwbQA81+y+uSV4k3BOv4+Hv
STLM+3gL4tEhbd25uwnys2CPcFV85k9DpCO9hN6i0VWdxtLdte1jdtr14WyFtBM9vUP9ikVU3HQ8
Tw/ZdFVGtYoMYD9lR5RLDfir87pGDcI9EOcdiY8TP1wajAoQ4ii4/oM0ERhS5QSfur+WCwRmOmhL
fahdrfB6M92gTKilCOTTk9RDwGyU94EY710hqmK1zkyBDjv8M0EVNv1A9/qtoHeeqxR/jsPCSEFj
us2YcQh1ZhFctCoowzfxFA5am9yvjN13PBwbKPKcsqysVrlY2JYpFCofYoAMAl7AmxHbtpuqqB8t
LiqtJe+6mKKM7nEPKMTA0vP7APJZZLbf73RA+7V3ucwIXpp1K4pAAbnAv9Arjq7EBa8FEUML3Ppq
DsnbTEbJa/7VAi8DwiJExFovIoTh8m5MMmMBFGzC+19Nr7Zs5bBofMIsku91Ur5tjkaJD/nNREaU
bRUh0evbQzxDpI2GPdLaGCke6EUVlB4jl3lvTcTWjG1kQpQhoMgyFZ/B7wayrtIJV8LqoXklhRg0
oqobUhALhseTzkMAtUo89mgAt1ra5xcVq1gNxesMh1AnAHg8yKIEaMZTkI78bWiJbDKWqeaD1RET
yX4TQIDp5h59Wj9r0YQ7EExRnBWqlmhuRPIua1vaDNYUarQJQprfl+RyaESIFKPD9VB2piG6LC/y
6qOWm6gsY8oN+kaJ1lBURMq368eRoYQR/X7a6O3GA1xH5YrsNdsWyE0qeg55/XVrRK6URbe3KH8f
DfWlMMYmSJvf4oEG/M3COaXFs0KLE/IkRDOFwoeiSH+V5mbh+oI+yRzC0Rk6K69dnqXyfjqNmovf
zWDNSh6dp5fO9Rw49wBf3jz5wryaRLGV5YS4OGWGYlpD9sucvUe6l0xOdrFNmFiD1M/8HS1KjGWD
myBhmpsuzyfbdoNfUmTwXrBQqt96ecqfqgLrR508KvQhPJ7X602pXgdFsXp/bktSTQq/bnPUdhrQ
wBzinM7K8na1ILXLGXWvhXuJqHemZOt7AY37Lw1XV8gadBAL7XNMBLGbzAZmTt2Z2N3cbNgQLknQ
cTrpz79qHM+9lodEzx57j/goVmpUkEdWEoIWMqWIVs9hHN1YAbvcDtxkFP/OphTO33DKKpUPWOc7
pmAEjsx5ixBYhQ3hJGATMhwq0OL7+khU1LV3VvE4EcDoAXJYGSZztUEZB7SIRTYUG9yrL38Xr7wG
QwxsmEwn7nFTaULa6Z98U3BJu6l1dqXYqcxQPd89++LIjeGl+zcSo8FbvEoLNJMdPEjsWkTW6hSA
5OHeRpQ/om5JeZV4RXFlf0aiOr5HEaRNEIvnzYLz3R46p2iA+ei9S3DOP+PRDmTcs/qYE4QsBgYu
01ewb4uDiXLkzuuI+sER8Fc7XsYrqOpnp2qokDS6gJ5zMBnA2aiT9MxpIviIGdxg9jluqfkL9hf0
J9LRceI1W1J9zV5ococz9u0KH4pKWnpCVt2Sjvy1uuGo0SzHatmBuEMJjsG6/BRvNHYVFQGnX1Hq
oKG9rSnm3Rz2rekUb4n/LE4e7Ho1vqmBLrtQqm+V+9UN+KnWlzb1zGF80CGpc/Kalkwb9e0KMyP8
nwhDX3hFJEniTOr/kEmgQZSnNsWkh7Zl+EGZl3XcCHkkN7U1o+CE4XQpNtpNXuno1tqz9N3hZDJ3
uiWrkQtDrNYmkm+wM0P8GamGczgvrr7K4/bT5yG4W/b7hbT04xfv15XQ6BDdqIomG+tQJNknssrJ
5YNWZV5MqJFmqp3G6WfXlNj/E6t+hiUcIN8coIFka6iySdKXWUhrOKvCwAIrIXLvvjsII8dbKeMk
ZVtVE+f3UTLw6Mgy+ylSt9FW87eCiN8hmx0wEnDmhv4k4lKRtQ98McOBOykmNT8bCKd5/9xiGPwS
sCCMn+nuvJk6l1CQ4iYjQbcwwtvVl9pg/j032aRDoxdSLR3oJTfu1lp+9rhrwjoHsZcVw2rOsHIQ
DHfRkPXag3tK6eXqFjIuC/nvlfW06Ost88qKHFCW+2a1U3zv8Hmdm3d8wCnrQmaDGCH5P9PxOAu5
zHU9YT0AFL+7Gq7bOJdw4XysTSCMJg/bAxOY1E0QPmneu5n+CCbGbQxcrcg4+uPUSaXN/iz/TLcV
P+1Ok9kl9ao9/0cXGBp2y10IQG1otn1to7XcLlXVR8qaaXm3/4Bv7tNazuj+b9MrODwaKZcGmmPp
3mGPLn0+/e+glEzfvVa0cZLX9L3/9Iw61ZggLRwD9UpxE173uVTXTxOAuIj2Qio3qvkMHm2Z6gRt
KlRg3fkS12o2XPXtV4jochA/wwr1XG8zSejUy66RgXMOS93gtJLy9fUQQBZd04FE/3IAhVFp3YQH
7o5kAjRA2DqlHHy672AcbhUHvHZtqa4W0Ga7UXLIhuBB6NAXuTNcBtuoGXGsN1ukd/7XDIZydmyy
ZXeEbfYYz11VqX0lfpPbuT8WrtlT25pocUL7YLb/XQfLl/2BiDXTN6FAvDZF7jmgC/hKnTuCavoQ
YE9NtOQM6izybuasIC++RiaAyLEclG3tsmhGR8O4ma3ujhbC02ak6++iML/prabHOLICTp+r4bFW
9NeDdeGX0D5AQIQIDqXdyIJ5g3QBvOMqrvlJIIY6GlDcJgmSCXVHDDliuVbmq/2VICyD6TOKeQUa
84+ufNAfAjLfOWwIVALm/yzzVxDiW5IZBJtLbxhoqqz4Iz/FYwe/DBu0zoK80IUfLWUa+tAtRvOE
puQ1dT5sa5bAPEqOwvFvVZjFTJ1vUtqL8owGaGOp0hWuXT7Khea+lmsSCQMbYINKRvmY1tWTzp1F
EOwTmFOjhP1wJCRPXvRYBhLEjulNAUr36qhet7QZVib8rsFZ/yZ9FOqM2k5wTw9aXjVhuebGnSzN
D9bEFK/M8vmiFOCGUZtEjjUzIomi5kdm+Gwmoh4eMQe1Yb7pRUFhoKW2LeRsnQMpx0CDvCpU504Z
/plLRBtwXk6w5WEQZ3u67IR3yqMrO+sjoIYXtCq2xCP6zDgBMKqHketfPSFNBumTGmJTEbWo1M9v
LQq3GrKFF8yURf43ZPazFxkwLQRtad3c40VNJLmrwNI7SalU0rf1PyyTm9Fh0Wm+xBW/4c0+aBsV
qK+1R/aRM+g5yAZq7quQ19R/Vhz8D3AZSSl/O7DOLrOQzJjOd3F2EDDZyR/0+KxT0GYyLRc6WVcp
HBmBwUH9IcAl2roB4uI//uBZBWwIDR2FFPCb2zgUfpju62na4l8o2JCCcsVy+PHPW+0PzuaFiEkX
tqfE41Lhwi5aReq/h0UzUXVyofepHYlDUTF8S2XYzF+H8L7eRZ0C0zIBsASFbg/ZMts9hLT6OdFG
nwpikmOYWS6MA94TR2tH902e9mID2QYTv0xfgYwCVZPth4e+H2Zh0Q7axZKFzTO2qRVWgajZpYwh
T3SCayHXigS3qOCMFmAnFTPEvZ33EP/ipwBamJENMCxAIgXNLSBBbXDVh7q3FhmqdshbRJFB8hJp
hvkmkPImZeD73cK5FLJsd5T7+kKnCZizwp7ap3R4cV79+4bpddFtBPSb6YGRlngban7h8puxXvs2
Jh++jFLnSaSagGb0ZCOfQTVCHO7ji8lb+zhRAxre9WceF/899L60fZAw+jhzaHEnIdG4xrNaesaY
RjhlTfBXXgoKzzEvLxi/KdlAGcjCfXrL+pfNxw8oNOTAmaWDJDsiR7Qex1cv0uqoUz3xlOxZfJyJ
VplyoKuGmTJZAgbRv2i5UV9H+8fjL5T7GeL7GTnOnYSlRv6n+PKCzQW2cE3oUMX2OD8yiJvie8Yf
oJA1yl5gb9LoCR3YjUhdNwMMZBq0vZoRRdBMl5CnthSyI/+wscC6ch9Bn+zCV1fSUImLATvOSREe
VmBOZEV+o7RW3TYhWNzGfgBJseL+NTjnJ7Z2CsOb7dB+m9sf6lnts+oQvGg92/NXN1PEXQN44Tcb
NSNe866EGoOBam5TBnXTv9uskM+MoLwIOPGeU+5OTTMCx7LlvxPmhEa8QQ9d9m0hlve/A1wT/j6n
EaNtj51FUl76vd2zKC6g1NNWKi/oNtoRhwY/3G0npcwwGDpYshxtY0y0sj8n0aH6pV7kVrNf+323
cur6D7us/XILAxx3L+4BKx7aY+GIr9XH/qmS7A645y8yEJpYrILynuYjK3wxut+ZhhRLK83mWaIP
BhULWqPhp0ltfwCBDJrpq4uppgMR7r1y4baeDM1xcfNLzm6vl6F5IKuBPy7pfYxNEj/51ecDQnez
w9qqAjra+aTzw5tmPZxDPGp/DoOwncTpS1fKWq5BYWteRG8siot65hmC/3TPLF3jFqz+2jSq0WTK
0PLLqJtDqyHxJuBT+6Y3La4/LRo/1M8DU3lhChfllRVW+UvX/Fe4b3QYpeWpR6rrNW1A1hMPe9ga
UHtHUxctoiD3kaNATT9/jyiOk2pGUBcL+1tPUxhR6LNqCamocPmWeTu1gIOsamCfqYOngW2DK5Tj
0j6zVhebwHUXUSl8ukvrKG6zWxJYDPs85brRnqy0/MvdeQuHysTwYOleHgW4VA4M5x/22rGmV2pd
GDiEOCYSAxYvRmH99LH9kqUel4QNMb4rB9FL20l6ahrjzf6i2r0UnmIvv43r8Ph6vGFQhVirM186
19o5TSJ5eFacfXkj46fYb8fab1s/bhvBSNUfHz+GhgFrMBCG9w2i6M/BEc02N2Gg+bpaI29R0BgP
LsiStAJ452SomP097tv8hPbNeWr2MGIut8ofG11lvprXds2NcmXrhTLAwfXKtvMKtpoCUWBR8D6I
MiD+aoNXr3NRj1mTk8VWQrKhASlOmXbKa+ehnJ/38FQgG83A6XNVkd58y/7mjBLF0EAJ0H/0mBxt
bIP/YSwlm8PKhZxbbBt/ZKoAHVlpNyYr+GUtv/n9Xjdp1ViltLdshws7aiPRlKIwHtD3ZgIb44dF
/ahwI0VDpuFZXCtuNd0htlZf2vObT+d1wffW61gGCLExioCDaIbsU3eQ/TtUWExtr4xvMxV539dc
1ZnMY5hVEo4itC+ycYgNP+X8fKNc5N2AsXZ74kw8Z6DnAZA6A89VN4MCLZSdBVmqml3iboBr5UKB
bYpgkxzYwoGTiU44Wfncl288uls2U8bMfv09j2gzmGS+ow6tSXnHHDngZd6MtTZX9C12rsKiAZIc
f2QNixa6QOcQA6JQKvGxDJflSM59gULqOpBlZTsIQuCfGMXZ+1v078kT1uUhDLXz7OeqbipeOTys
gw7NV/Jk852lK9Y4ie2ecO/YO4rxb7BAIb8MckCgr/UINcdxeDI6851D2TX3aRtE4n0mWTi7EquU
5BwaylGZJh3w2Gjyliq/yc4e6qjq2q/iGDYAyaaTQOQQ+SUp1B9Ozb77/samItO1fSRQsHKeVi49
P6zfPC+BFelpSQfnVzZg2cq0w8y6iQHxst8IzUkIl4MImExkKuWH6JtCdY/Dw+Uzk8xG1iuDZ3f+
tXCQrS8CVQTTu929NuUm3oEPXMzYei3qT9qCU8T+aLQO15+1oy53JzyTYAshvoi0nZGXibX56TmS
z00fLbZW7bnUtV4DGIBTLpJbEYh1Buf5p4EWFcPOFPFp7byaJOxTSaOtB3NxAZF1cdCp0uIk6XnN
8YYuWoIHXbD8SNlC97TNXEsmnKofRgvmQkTCS0FVn8FXCdWynoBEEx11rfVYznzSXSRouOYI8rPH
OSObYZ+Y6TXbBjFYXOE2CMdtI/J4xgxb7wU7zr8+vD/2GzdcqOAKr3x4Argb9swAAIxQbjygHofn
4n4VOA/adG+xXp9vcy1Y8KaUu3Ub1OsGCo41avSIRySZqEzApkDyLF0q2r6r7yYfO+PUizhhb7Cn
jnMD6V4fF5/7LfC/AcrS+wsorpisR6XfWOodQXLnUVZlxX9dZlL9aEg3ByGrJZgkV7+KHML2luiO
IQk1sICSSWFKJMaKJnVGC/F2kQOd5/IeoVLUz6BwJvRUT9YJmeXaTsk6PTdQP7/WAIkg/a+tH4ee
LjNrTCHTYpO+T0RceaW7csGEBpuXUrm4DxnRbiWTf6g4HbYlGgfiyJiwJgeABlPQRPJhznfqWVTp
j2Ah+Ct4dW11vrsUMTNAWj8TaF6pWVujFqRhWSxV5IZNEVMF2n5F+zKJBF0axXhciyVlcUCf8rxX
JnMWifUMfksJE/rM7TeCa2PJm/IyX+bk4exSn/9w+u4G00FF84ZB3GhFxVW2o4TxMbHAOQsG1DLV
3eK3aDNUVe915QhvXDmk9pe4RXVo6GcUfAU1BJ0NDGi9fU0MXLRPJoNHsYMiKcfm0TsN0eH0ZIYu
ZGJrCl3uevsfW5+5qOIJem1HU7W9tCkRaK/hUkV33QbH2E0IIS1Nl8juZqJl+7a6w5UHQeVW7Xyi
68T250P0X7+N+BtN5VF9gucsgMrpv9ULOiFpptsRG+3dv5zTeGgyBWm/wNCL8IPn6jmwq99COXoH
/RU4zLNYxLhOy8g9ifqZmlwoNgI38IiDDXi0IGidIq+VTd9mwnllbFdYsRHSCmOqSqWmReypB3/b
JkrnNfrrfUUpZkwg6wtGroKxohcdXtYt9bm4ZnX6NdXl2Swl7I/jCbeeNowwKwAbXn6dEfKFou2C
oX8gDh0Mj3EOy9+jvK0LTqgcQVWD7qqUViOcHN3wi1G6D1Zx45c02hI3jI9WefPkIr6IaQclo4pe
292v35FNsOR9YLu9iVHONtxzKSfdjajLz/MamDIgyQr91t91zsZs/sNFFFsc8vO6x6Lfm8xuChdl
rwuzZMo5azDiGr35aM2ISvGGJvKKIxXJNLbDOpYA/uRCma//yCZAzeosY1MthMc5JEnXgIzuQL4z
LftVcxmU7oLXCwadwhJzQov2FL/iKziVJuE9jmHsa5i7RiCd/e8SrO5ZvAPSCH4IeHkFTeX1MPMN
G83iqM3VarXgJL2h/YfH2oU5bfZOyALL0M8RvcStrb+LRnTZizkmeFVadQsaeZyDnKMWfCOheB8r
7T+DiUPcxqno1xkAlaflqu4OgjwvOXxYIo2NZVU/85xO6c8xtLqJXouUqhsQ9V9uGg4a2MOfgGwt
BxlchaapaPgs7sdc35ojrpYpbbIcIFnGrIznUS/pf7uW+N5ukLZHtq0tvpbQKSiE+pAoyX/wwNox
f+zNBHG6YJCSVZRuG3jHV6odBHudRyrQc9n3wq4/5wq4VbVTp/XRzK6u0UYVsKaDV41elE836Prf
DRWBGACjvq+XW7uKjyR1dkS+Hy/QHZ0Zmx3nsVdRiuKkGcQrXxIOhHXbuuY/+66GRKEyhduhGN7k
rSWni0HMiPScxu1MrvkQDl3z+Zkcq0Jre0OnbKBXZfb1FUNHcZrOxscVFoxXO0Oz2WHEfQrZGezU
muYDp9NxE7xrOCKhO1/9ocdhLB95YQ64w/SIp9/X84FRgftorviy0a6b1Q95PhL39nPnbg6vWUsf
xWyPUJfcU+pKzDqHs9F5X6b4J5oqFk9PGLG1CbUDWeyT0HiIsQcJBhQxYkN6nFAD53S8n8y2cK0m
ni2wRLK6ayYR0BNh6NGqpVXtEKo6/cNkpkIke4E+yBMZOYDm0rqedinKWcKMnJzEQJSL0LbHU1pl
PfncvhVBKjEV9SOsxAqlJOJ8YmkNUYcdUOf9+/DgeCK9l1sqP9+t9GKbxmXhHDF7MKD4KxicBSTq
Ci+D4N63L40CdUUaOzdZw4sQ+MLSSq7Qgndi6zwR7wdLgUrrWYxpsPu4V32DweytKwvU1ZlE87bv
YuGLNI157Brq+Oy3BwZOUIWIHUQEvOT4uO94bjIDm6lwEiyWltjmodro1fC7UuuPA1+J37J72Frz
NDPWy1A7cs7HBpEGrDDuqnhLfgHmpClFxMnFc7xMddFkmO7ewo/JGCaHrpg89Twzw2lQmTMHcnlb
xdkVsZjtSsQz9sXhc3ex8lDbJMNbk+E/EegiX7sG3jd7ybEAWQFxvrKa2Hb908cQo9v80aH2GGbx
1hug65uSBsMsMdcG4gMy3MkzPeJEWaEEDuNg6OCkxabnshUwP6jePAPatWdc+iZSEwUzdqJ/B0p0
jFWhBfNqGYCPAWs4/FOs5tkQH/mUZ9NMps9vvjG67KgdOfT6ThNhZa9xXwq6uTisVk0omEv/3aYJ
cQX+DjSPba7vKVxbbmOpew/GviZcqBg4MIxcIIg/2UbhdANH87Lo9qI759CnMMlloisGOZS2t2Ky
pmKS/i5HjW4vhpVk7VrmgPZxLqqLirwM/OxwB6zyPIU8xOnGLNQQJC3xs6HEtLIcwtuZX62XY+DH
LToomoyaR7ue66f40Xwqtj9O/KTy1W3UsJQdya1dzG00/e4IxWcVBcqnO7K07viNww+mw4/bJP/3
Wj6IWT6hp3YXUsJ0ZMaxfFOkKNy+RfyW8+znFIhgBHYVu1dhUWX0V3C78aTi2+zv5vRuxn5qdJh4
XxrYP+l2JN8b1THgdU9v3kU4oW4vZO+/xaY6Rm/98m3h5V6/ouTFQGaUSZmeuMh+Q87ZyGxNBbmW
/0Ng/vW+SX3ZKy3SAqWeSw2jnOe/rGoA5i5THBHd7/SbbBhMOgHAhjkis+vi3Mk5XyjD4L9x1i88
PMLUf56q6eKz0XSjpUT6769A9GwwZcTEZ8CubdYF/afpWLT8hvYyrRXBSxNBIp8qmBULwrdlVYJF
BIpQEuVIWhtpvYjd/yQbNa25gaS7Qrm4p5gP2zTJ3b+v4dvmxicTsCzX9Uevd+ZP8CIKE+UhDMO0
+L7T76jQ/gGP1Y84FMMgQwoUsZyrQV+wcNqdDNXuYZSlk98w/ipQs4fWTO2L+lspmHzRI5DW0et+
QJeY4VcMkdygmdybuIo4Nad/6JUG66WECMm7s2ggZT0/fhoLo1XQr5xVzcBKTSBF4XrjNpkqbSdP
vd7NvpvAR1YTUYQmItoFoW4U8tBu+tS60P7a1OyBsJB10qt/M6TesTBNil1krd+o4OqBGXYn/ptC
nkcLb4mll+xJGxKnSeDfvfBnIrF5UyV9tDc/busuJnmneiNQMR3BRJr3dAcen9KQ5XWuLGUEBJAf
5dOSqE9tqTT6IoRr+5pCHldLbydepr/X+Jh3RlzZk65pg4Kd+Qn5QRO9ZRX7Q8hzayDULzQRlOjI
QdYUc7FZzkdm7RjWnX1/7qTIZYcu/AdOc0VYilg2oeazDO/rA/nD2a5LydsL76jdeyU+tMpLhOfh
z/q9VOaXqtHBXyNpgl+vCZDjR62dbvUl3yKV4p878HfTuj69J1lC1LXDM//j5FKX2m457d6iVdxE
eTjIVK30oC0ddryRPHeEDLrFN91kvRB7On+DbDMNU1FX7ck46/YZSCbIplFpYeZnQpZhRgnxbq+x
57hsAHGCkaCXyixceIhUCXjiiFtXg4EW+XURPKrTln3Y+paQvK9Y2ozfCf+o6tBWV3jfflcYH8Ag
5BeJfJZ7HlR28BqrCiD6/t+PyDTrfpJwiO9kUn9sdifZSmKLyq79kQu0ncG1f4j58/jOqsx/d3Ff
B9iuZWG10I4ozDNkUzX+eyi7P6EGbBB/BlTp6zr/JdSnr4ZqYmiTKh7fI8g7HvG3gPYytRLnwUbT
oWkNupZ1jU7k0jw23sntNGThf8+J57EXofgJsauACA5qUwSjva/TPOBFaRSeeCTzE673ROt67T3K
HH9Y4B4z4E+wE8e7mAKqurwsZDimfpiMMpdWYXfU+DpqNFX8I89+zwofAVplkKp3bAeb+yrmgqBq
G9BoaCLLbxZ+jLTJmGbKf7OjoSKxAxHExiVZNUC5hxUcHEzTn+mQNhHWx/pgFHravMR5Fp7RBEHi
Z+SnOAWxo5z+c5xP225rsr1KNFnI4lr0+4A2gr+vUh6uI0GdxcVjheGqe5w3LRF0YW2y2KTwaAR8
QaqGUcNY3mYDJqZpDoaKFdrnaEnT8HJECY+Cfxm4SkPxPbJ08U3++WRyX16Co6Q/nFYdizSGqWww
VzBSlx2AGuNRSNTxM25Ks3peEz2VY/eZWpq3N6BxCbECV+4frtogSHRAvLwAuE2ReARh/VxIdjFs
3eXc9xfbY7hD5HAbvvfZvPeqXRiVgFjGAIoZbeGbosasjWP1+ZXIji/V3sxM34LA2tdsx0jlapO7
nN3rIEMKXLxiKNaP922FTiyTPyV/oNXB3yIBLCv57iDSEteb13QAAgukWBYOl5fDG8PjjvHcXGyH
P7wdg0n5R5zdYHcJTV2Ksrx8IlNhbRvON3j3QK17BQ+ehCAfjZhrxpWCoHgWwZhSfcC/4odu1Im4
+zywe8cXYE0Z2m7aGOvccEmqsHy5EwhQQLjChrmqZdnErbPRUQhbocTrmbd2yG4Ue9fOd4U+1kvr
Z0dlOiS1P29NOs18vKkBXeo/n78GkBjo/ZA8G8rGONpZPlsF1CwRsHHMntG5SvZQ92Dc1h99GX3h
mPyV3K6/rYAMM+B0zYNJsfV06HbXkAdU4BOpFpGOB5B7ebNALMpxCeuV8FpPh2stL6JxWnL9N/Yu
pI1DHdFT5dsXo9IUGR4WMxMXszgdL1RARmXT0cBRPHoJNK7HZpCgHagBNRHSvRcTXGPZhfCThV3N
uWdsLL82s96mMhkEPXetlhRCLGhEmsHayl0+fVAS1SmXpvi0bRVfhb3OLQCq9SFoW3/SNfUUFg45
jLzCzwwecXusOme/TjC51PVDLqUkOjhgWFMgXugGcK1/91lFnf6qCOWosRKZ+HhZHp1t8t4mvn7e
A6JiE8a+lSiuICY5oW2G0ZWg9dITN0zhqYRMPikKiRvLRp/TIyyt1sjREGktduTvR1eujQwT3V7Z
uSPY/cLyqnjMrJssl28etzyvTNJ+KGNEVzPaAuOd9TbZ1Gr0F9q8RhznOa81vz16A8a6zbB76Tlv
lX0aXsPlA+g/vFP9p1XF0v0dhKPcxDpjDF+VRgbVDBWo0IF2kzgaMVIIo+qxWz8ENXM4MQR6+RVS
d9NICBDabNZujbHV8bR6p4K6kzhpBbFLnBZYOW50sRSuxesvBE3wPMA+tdDuxsQI45r8xhrnPTkv
RPdrRUz7o5at6gwnbxjIqH3+W81bIT5X2bTZ5r5yZpukDjvtrzVYNG9o6nXSZvz+pPSLqN9Yii5V
VcdEzYHxUdplBO2MjGwaE5a2k9ZMxwEJDSMzhk+09/qazyopts+cwoJOvrIOBU7Ukiz5ErNOmHTu
QbJ8kzOjfBcMBqb5Fiw5sQVAIQAaF4VWssFkFeJFUz8DO5CEX9jcp1TKtywliBxVlXvC0DQtXymS
UmMZN9fRqqXZEAsCmAsR46SDOGotTrk/045qcqT6f8CR1UlFPJV9JVmtKwsfSJqXC/C1QH1ISuUQ
k+W9CfeEMy52AaXjZZ8GTC1w0Xrwl/cGfZbJq6jZaKQGtjg/T7vFjqypd9JBEjrpdPFALLg1QTJm
08V6JQLInx6XsT0qlqDVXHi5GDWhXAPrBdW75OV2KPD7FWvy6S3+PUg0Lsf7BtstQyongsmpgiRN
i9n65R0POc26tInupKajWymyeZ9ATgB5rANPMfNxNJSrJoMQYrFdjJtGE0o6ZPMSKkf6JUB4M2SU
LlpVixRXSk+Wl/2QZ9k9BV+hv33C6z/Jes7XaWh4h6m2GUhHVNuYVA2zyVv0B+ubuIOZsGdj0/SD
vE0qGLxuD3A1V87vaqJEtnHJUTa2Bp5LAHnxvHGftrQ1JP12J8ly0Ea8RZnm2dOWT9p7JyRc+cq4
bQ/h9hO1QEwPrKWzfKbtbTwbQsnkQEs4qD+GVswRA7y59/3kWeehiztzDlEpAkBdmI220Xb7cAmh
jsCvvHjLqGjnYE7OZINOok3d1dQY3t4diPegeB1ZcEL9Q95mDb4LbXcTaY8MUusaX9ok8Dya95T/
ZWk5uztNI2EhVqYph9WQrnYAmw0553NC/tmVJkgX+1d4udoEujTFAPqpbMpimZRQdN28uZXQE0zl
6A0z1B0x4pGpXYoIwrYaUcW0SMOnwyrmD4rG1madN1+s/j4y0dREySX43amJfFpQ9kyZUS8nNmZx
Dqixf13AvtChplkRpuXSfTk6TNd3Wzm8uda85AfsDEIY6jvz4vGX4FIY+q2R9u1MvQTbEw9cJNfF
98sVOmVd/51tXqLXeeP7dqMYR5riCLLB7CPxoGa4S9y5ShURvp/9CeNCXX3Y00KIwnAl/e6qn3cC
EePbWhHEPsxjHk8HPcxgLvQ2zkrt2y4PWQwD+gg8olxcS3zfGMYtN3FYpd8UCfxbvBwA6gxk3uvt
277bcSH3EriNBqdc/dMvMb13dxgYMapxsElx0BYIbYiof9IA9UjLSwwHVTe+VUX3KF2muzDViGVI
ddXe3dLQqwm6aACknHPYEGHAEPoNoDyT53kgydwxuJgJZ4Bw03DnOhsOckgdEg1ElUf4WKq1ue20
JqCd5kDJKyfRIIYij6NqCWODtTg0jJMfE2/GLhSP82e/T65sd4l8ILQXV8MbkatswKaRsUlpdsgG
CEpW8pYoewGMARhyk6JlwfryWTtvUxn6GVjS4qdExBIRANQAcJE0oLHjXzPy5pcxPCR3eyQygDVN
BoyZNgKaGCFdRIKCiT5EM21z62fcXnAUF1W8SmwU8bYalFe3hGP4Ojl2GNERabPbVCiOTgP6dfdZ
+bv1vp+8j+abQ1iRcQXgZCgXofGCqH9r4X2MZoATPa2lvCRucSztB32fBpvvyK2gqBGeOvRCRA46
8QjMfyVx0I5dDYR7vvDLs5bc8Gg5syoBlinjmihC+P0Y1g1GjQiH/AQ2L1DnNxK2aV1DER37m2UO
2NVTJNqiAqssujZp3+87FLZsoQuvrAv8+BppR+UAElTgtZH19Qx+oZWsMypwQe0F9w35D4TJV92u
o36pQZRNOAKwvneYuzpTiLwwzJe4QddJqMYFPD8pc1YUhl5jmJO+EYp3dctvj01RhKDVfwcHljn6
GBYwghdR1edypvof3UyWYJHtj8hJzdb9eU0OJXwUqLBKkjGbSdv+43fLrjX/RPureGQP0cbZAE5x
wjcYbv8qJTWm+amVrMRiPjYul64/KwtSutdznIRW4HVswauaqqWw+jx1ZIQNYdLNhegcOdYEvWcA
ITsBiUWwPm3vXpZXGACfTILLpDJSKgnmsUqlmBFZjP+d63WgousN20bZgv3RT01vnwvho3OVNckf
Vftty1Hwut165nX4gt+hWWUUC57Kg5rNfZ5GZv4c6Pa3XppE4wwL0QXf05RAQ26kVq50mdctbVae
HMOYWwcMho5Zd+oF80m7H1UiLLYCrMoSCLWAVkWIqPs21T/odF7qg4a5yqqfEfPK043CixQp4ItB
qjb/9pf4cgoPtYB9shUFQVQP6/t/3jgFEh/RdISUkuJC4OCv79yf/71b5F58irN7bAlbqG4p4WNt
0tSGPT5olxaN4oninKR0fd2q8xTcJpo166fIkg0eilavrrnGM09pbrPM2eAn3mz2wlB6END7lLPP
GZpJU52KzpX3hitJDsCrRa8fw/sVNpQMjObikeVNDm1JCc0r6Ojllot2C0dpKbIkiukDMUx6s2XG
f45pEdJx1QT1SdCo/zHC4d4VMb/Q8BYxbF2RoEn+sKfaW6tU2BAcZrPQytC0uYvk4zsaDi/wmHZY
6/+sCwmKi75yV88hcWcBj8Habyvr22ddlK5fkqdTMHq0vMYBS/3H7di6xwQ/Yz83bBFu1EXuGTK4
WmtSEl9GlgB2cRwxy1bJLmjNGnid4c4hDcPgHrSGc/TOmkvXp1+UfxJp7k7UgK7yrDxC8vnEGY0O
XgdEECT7g4NNUgkTkZ8J8YcQ5hfvnmYHwDBQWtwhMTh3cp08JPYpUc/27Pk2o8J2BLoXslifKvTF
BWQA6zbwASDbgrWjFPIn/H4AuydbOBF22fN0LrlyM0bXwDT5rhJoQWH8UBHXWCJ7in6t7PeABs/1
eNPVqQLMCriSLim4QIeyVMuf/8cjOzRDRJv2xRuOETAluLRHInXO6aV5KaPDidq/1iPwqzNdgjKt
2i4vGXe3cc1teQt3qSgEROc4WrlakKBnc0di7sTtwR4p1HqQoUUowPRFmLnB716ej4G7dGJtuu2P
G28eAH6Cr03zir/Eqcx4yLPjNOLPVdpBXlaXf5Od0BbGdlp9DqdYcJrUhdSPuOpRmGn8zXiLiJLN
IMWoD5m8G5dD1q0zlMKL7D3ffvG3A1z7ZpAhA/UWT4Sry8OQEJn7hUftld77yTzc7fA8jyJ5hJMX
i1tPJAkdqui2rUuZsdzhoCcrb1fZmC6FlZ4g0A62uDayD51gucssQsXPPTqb337D1vS7+FYPqa68
TNNAtLkg7mADUH25AFGuk5BxnR6Fxhpfpg8zj/exkkhWsxTDvfBM8Z35lA3MKynLBaETgsh67fJ6
0gp2POteezU09JyKLZfh6APXqqP3w5g7WAeuwqoN+AW8HUP7BFrtyHcTAcMJlUhn6sjZgoe78ARp
nbK5OyY3yLsxmkKP5AcmBhdcEripAlG8b9Wx83QvvUQcNMZvpk34uGPsAQsTW9lDGcDarkoJj05U
gu7trrUEJfs4BValFhjM6OzXwzPGbnx1UcpNixU/ZcwrYO1y6RHKjRpUwEtcSIUVN6mZsfZKPM1a
3/+rQ5+W0ReWF+s4zVI/OqO0YTA9OZ7DR8pmNwl6Cd0ZZh8ftXfxu5WwUy6Egz7cHgP3s1+CfDJ+
D4l57JOWxLfV7Mb+Gfjn9q9mj7DVfhhDgBeiF4iTpr4PxUZuZ1n/hnsMZWuOOUIsPCQ2feDKw27y
+W55KrAaryh/JCPEW5MGd+Xl5tBz29Dr18rh8kj9TabzfC8DmvMjbFL+PepuQP48ZgzQ6gKEdxyb
pHVrzTwx6+08YRoIftjmpesHYy7ZeJws0Z9AcXbwkBsgrmVLu1qNV6dnzps1RwTwPX9TZmof5JeS
ZOHXUQJSsswenll5udn0hG8pYoeXSjw2DUd+fL7xpZMniXubMrZ+I5QiSvS9SeepDZ5VVXXqoUnR
OcGNvMhRn+w4/mUgHjccXR8HYTavs3p8oZJ6yEUaokV9eyfBTn03aL1RcapZZDfN+4quhT4tECcp
q44a8X+GtYmLpGDo48m+6B4U/I6Qv1xVJXhyog5N4Z5IOd4vJnLKhJXMDyRL+ECRq2CLbsi9kuka
C+XFEguvFCZTBpB0oN8l0n7XpkMg/+XfmHgKj1zi6qvTDPEaut8mbT5wq2SfpLZGATGMn8c2/cby
7R/VaOBjr4RqKhxfniLqYlq6B0u95+8QJ0V5P1xkUaFuNreg4IskPmpw2lZ7JDuDu/QjRyIBprtE
j/Kjgc7g8zbLpPL+5sF2/YIa0knfUZ+gPnxjk5kGS8DUxXMx39zr4FasalB5dc4ImTKHqy6Y/MB3
D9wh4d9PTyRdoR02RnlnZgwyi04pgIYxpghhQlQUi7K2KznIhxghuAc621vZ3oVYHCwkX3cTd0g7
kUqAuAT8uB2wiPefOTtMm74rtlhMaSE0+J9w214Udz88wpQDur0eHWF/m6Hlki5npMQLSVh3/sl4
1W7fEP7ywNzcJ5M2isiSBBWUEgNkogryLEgWECy5u73WVJUydzQKT8w654uufh+fuuBfFVZ+uDr6
KWJrNIPkhB61WaFHueodsoo9IVeY5pDwMQHeGUV3hQZdQnGWaZh5s3n0JK0vDmWil/9jxIbxnHvO
wr7r4uGlCdjdb2TrCmITfg3GPKXrWoCsBP+Vt5hnyyFH60QhlaqAyJormShO7y179ihTjX/GblXl
jM0i8QfnZoB2T83ypUJQTJyjAMU7IZyBI4ZAqVgEsDVMx48Fk2eXFMhBGXhbHXbAScpFE4OhpG58
d+xvjV0vuW/s5X/k5dgPna1JVSQP6HBQ+Zjs6MOybScbQl/3BHigVtsQttFTIIMcIuuJ7QXy2jDi
URwu5C1CntDYZWy/yqztDvGGY91q8rP90zHalNeF8tqRBT8BnQuup1EdX9qbgCeWRGUEPNDB2eUB
+gSkI66Aahkq5ECibj2FZlHjwbZmkg7kfgd72N5Sgf29azpzD9n7haZ0KeSly+SI7x557FabAlFi
g6tNeqJew/U+0kfcTJZF41mJIESWaohYOyxzjhzejkHXCrDMeg7Mn4NPeVJecp+auQ4QC3TJQlu8
suRsJQ2QRbmjIt4WkBFZXsJQ/X1g4HIA7zeftqD8D1o9nr+1Y5yeUEvavqr5fu2JCobfuHclbdq7
IExXm82Xw38N4QYDCAx3ldTJKeKG9tlYVa7RuGJF/DrZFczRpvrKAwmsETEBdxsGz+x4h/BiIc2P
50LPMG8u0xN9IKb/LpBNJv3bzrdWFuDBXpg4T6zRq7yHVP1MyrCgFH9PBHoLmO0OnrbG55e/GTA5
oFcctTmJXy2oB064AtuDgxEArGlPHeEQhSOkllzt0NbZKI9QjZwNj9Ymp2GEcJqcuX/oCINs8Olr
nzjqOes75imTcm/1SyyUXqH9UWe4R62dRXKfbSg8u/KBhtUm1TBqnRXLqx9zdRUi4PE6Y5c/X+dV
cn4qDpmP02aBXygWiPMsuMLr05+igcjyu4QVC1XUqCaaGFx61XLOez8+qEfH0hCu+cpnMTlkGICS
+Wdyg4RiZjehJ9Dt3MctGlFDk3rRRma4YBi/ZNLo2mdyTqNQXZd5DtYlNW6R92yDH5MZahQHrq+k
9VHSKd3N0nwb/7v3lmHsY/jYTjMZ7J1rOuwZnXUIyhUJzPz6jAi60qxdb5XEF4WGOmC8VShZEC9O
qLCdsXDPWWQaBxKyp1gmNsKgdYPoCFD7guCaFcYdYYf03wj/iFSFdvZ8E6Q7ei32349p1bwCMuud
GugkJTPceuHkdC5PIqCFwIiUS8PSb/8rw+7nBgMhuBKi96wQaw7WYegANZh1BZlw3Y0/nTH9h1B2
5pVHdj3HSi+E5JstYwzPemt2jmRgEFGqZ1OGdDhuT7TRz+3XsXQ77i9dmNJzl6ldtNLMdaewN7aY
JXR2LruNGOwH399D5Vbi4UHpYX+mItwkf/APwhcDc+4HNJtuzhrjaDCmcPfxRcglW8yuGZJP8FyJ
YO6nbsZPFSCIbEdjNZ4UqJINFnNmdhByuYNjfsXFoChpDv5EZg3WGEf1XS9h4G0RF7m5NI8v9Rd8
gVujbvh9R9FgQLUYpfIHq8tXzuSVxtxoHJEJc0tPLh80qDKq3TwK8OlLBu//iCcWpqjibJ/4iPTD
E3fHnhGiYdZaSb8u1QmSpk2vyzEyULzlpwRXg6eqAhjbM+AORGDo8d7AX4rKdpXKkB/xqG0QAPNL
RCeDc86ifWOeYOXPgZ1gUE6Mjo52a922SBHpMYx2901bFsadAMdvzy0c8FXrqMQ4zRRoZoSX3M2x
ZOLstPed2IQBrGc6xheR5yUCX6mRqjf/RG3yBdZ4Q7uaMCylZQ/aW1Cb69LCq4GlOoGPbNHPVt7M
JmFy4jDl1psjRVRLHRLh75zbQHAUYWgJ9zeEwaMrF3s/st9lJ+/q974wExQBG3fdROYA8Zl60Cc2
mVvFcCpjVuVu+JKjiIwC2Aat8Bu5qJjz/uj+RqVreuvFiR6M8NVbCxpl5KaD9f878+o3q92BNskE
LPKefOMPNyuPaH5ee6JYdfjXTT15R0xyvgrnxIkk888vScPBGIZiT6wOUm7LekNJXlY6gGXVdWqD
edjReVhF6EmXNpm2rzxdm+YDqiDiGCFwt1xFdrPtxWz+ukKgvXJE5xOZXAuhG150f3nyniZtCmbx
WQZNhowOFWw3L2n7mFCyPCZcG8SPuwIBo/2+PzT82B0pXoVY4NwwDOxdREQ0cF0rXGP+DzVl08Av
TQX8nGkLBIkZ5kGfuKc4kzcvOjRUp1H0zE5WUkwH5ftj8mtx3NEl6KwnKe1SC5PUBKLomxzynB8D
2lUSSRalTX9flkkyoyqppmsII2pEtNRxmL8KitqynPnWgs96xk9lHIhiuT6e5zNwwJ8A3aLcPj5R
gzyZjm6ez/93nEYRWOEwzfOvHEVyg50HtpS5aO0HAodS/UgsV8FiWB65fuPOtWdbNuyclpdB3Flm
7G4WzhAJNG/I1ghASWxuhRwuwGjU+AWniQ3odLpKsZuxCcwz4VK8It9IYnpDuq3+7jBFF8eDp4dV
zm8om0MTzD4FXYQEOhz7waYEvTlqvJ7XF/WAm0bdkT2Rla4arOG6z8/eFMadjIsC5AgVS6qHb88z
I9UnPuBIlQjYJjGnaby+hloih6KmFuHvIAkt3ssJfSq0H0+esAa5Qe8+cxeQjODZyZU5lfMV18uf
A2CI3OkmeS+/ZVS5qruT/UehN5KoWBZt6NwmQvEW/sEhMN8m927uGZJd607THWfAgIveD7Y5Wjit
aFZV+bd8AFWTEZvoAE5QMcF12M1CohwxGY5YLlnXdtMhmSLPpH01XGdCzbxNvU5jJDXJmkyDEMMZ
Lft6Em8rl/ivhk+Pf00Pu3kCXs7Nj8fy34SoIf64eIp26+6ae+V6dq6Pbka4gegNRJQatwhajO0m
q3TSqRGGeRmqOtdbr9xtBnSKECkPdf/E0CoqXSrFcKigKxh4yheH3b5Urg4zN6LRE1Ci/xR1jGDf
YjuA8h+w9qo8ajXaHnqHuu+tlsOz9LLscdzwIbfF1J5kk06QAJKzcemBOA+f7DYQwfkLsXQuQlqm
DFQ/8pQxxqAR1gDuZxS3rTMTlTQK1ipTtNksKDz3d7OIy2/m0l4oaHNbOgD02pVjaEQjlyQ1dcrp
DO7hjBnYDS83PscSqLVKK8b/V/fgGsrsHAnbS5WeP2oZJ8FhA2QwwQIv8Q9FgkSF/EaXDTDoFqmm
fYo/iD9ouq+SXLVuFflKPULRC9oeWhobxoL2k5Naqy3VKak3d5USnC+tyGUPjzntgC9fNvwFZuQN
p0JulS2kWmCYJsaixslCq3Oqb3zikSJ7V/HjJB1dYgnTO4W7cmaRHVAWENgFh+15/26JDJY4Pto+
DzlnHWyPNaD+zlFR6Q8mdt5wA2i/5IfYE08c4IYfO+E0WZdk2eryRbf1wgsrPHqhbQeoXjrSJKTm
mtrICsHv70QgypsF0CfzKUTPiXn0IQZGnU5mFZDH9mO+OZD0qRERunqD+TtOPoNjxqbaUrwSQe4A
rkeLVxTZgeeJAQUbFjd5XatwE8wVG+DH60EgZpw245X16SGoKaUnlfTDPf+cYBUJaEZuHqqF2p4W
WpYNNSc7FG//OQMLcM8PA04YgceH+qcD4u4o6xqLGebDtZIoyCm7y5w+laKM8YFLIZIx2cusvw6v
smUs1FX8yJon4W11Px1yryUDcZEQMIEL3RxE02o1mmq/ml0l6pkxTvX7uIX9bP45hOAqcKH5ymNx
qCeAcfF5C4QyNHcdzopqD7WqT09jsPKkRxslJo8tO1sBCK4xEtBqqitqHt5GdvJ0gND0EBmGDn1f
kWIaz4Ssmi06iHSph4QQCOO4HVGeolceK9V2a3SLX39cfpw9hSo3DUzTg4K8HzUSTRh+cUFRoqXj
D8JVHsgsrvUDD/bv2tLL4hPnGOYnwezNiRc931jFIhPYdyx+v47jmpG4oWyO/2wDqEd7YmLhPFSN
IDh1WDjzCEOoLELbMwWr7eJrxzl2xf1RpWiQss2WuDfVh/dznbktdbViHWoI7hPuhwDF5e8FUwTS
aZd+vVogV++A2ouRLEcbtMYYg2s5EMs+hkzhL6UpMV/xVgd9LX6DLoQAZxNd9E5hOsBnRT49FpVh
I/HaaA9hKYNh+NCCRMAqSNukheQx+KdnbUvQDbHbmYx5dq5iGCfsJWPfNpCfGmrpM+CqHlEmcBO5
IImavCmpbJSTX9LUquFPnD+5LP/jenEfibJpZgf2NmVB2y2ur1nKrcPTDX3OGFGIqI8bsl2IUOdy
bh0R9g4Ehk/TUvXbVEsGqfIoisCuIGmFkubYtKtzoi4042rrD0e2SYTWiXF2eYynCYU/HCQ7Gpdh
P/5uevuM+rPFAbCa7WmegfcIqzt8CnNBQTXc8OFnX5UML1ZD8PkjjRvm0/xtIkJ6yWGpfpq/zchV
hQNNbD6vZme+5ac7sruaGmSauUm4MU3uVS18cboOXUPqlKof8fXY8dIiwANZhsOT33zQKuQ0QdTx
2dPwwDJmCrFmA82kAz0YG+s5dv5VPGJEwYsZvgWWGh0M8tCl584ttnGKCwzGWEKNhrs5WQXlK0XQ
Un6T77DOx363aSXW80TUPfFdcD2U3zqXde5hi41PFtE3AAUnO2PQ0OOseCKm9oO6Nk20e/QP4l92
/UiCgNTZROCroqrDvdhz40CtgVSsuq3r96eFDvBh+6c8qS+R2z/thRaOD+mxDR6sbWQFr7h56Th5
CA17cDPm673UACfH0ZNacy0++AmX+EPHVEmX1G9T5rlPGEmK2B6Edk+jZJdhMqP2qwRNzMkWLbP0
UKWKEl1PRo3rSuAQERda/x4uzA0GxHHhigRcSnrQX/pswnVCsuO09Q8atErcuS+pzhtHzUCeXkwQ
OxJy4fx88FV6aZybIrmCeex0H27p1AWas7fFBn+HF+TGi808SzuOSM/vu9arIbsF2uNQYl0J1V7e
bNDhw5752PrKfxRxkOGH8e3b9x40fcDNvb33LYKY81g+OgL6b+nfiu3a+S57V2q2UBae0Z0/s/1t
1x/1xsiJ0r3TmFm+ippSWrugQL+cveejVnrHTM9SnK1r1GyxnjzR/mIg+2uyFLVJPnGd4rh8jbuj
LDFOFZMNczeJgK4LlXZ/jasQ54r46YMX/UaFZPSJRBxAF3FMC/UYPjSh4s04zfMuL6/U3nH+6JmU
/gEaUPQh87eisGFk1ufP97fB4rU8+t0kxiLQIzpint5gzr5tBBBhIL6XGNDqmCP2E01Lr+0PptZk
7ZcFJr+svBLkQ9uUZ+cMUA3mMMHIutYvo2ZoGNFJ8kWDdJI7hRZVkXOcasIV9jRsn/xUx3fjadZG
hLuvmXALiwOU/7SdZ5QIt13Sp+wJoLWB68Qar21gouinF84sb933qQcqtnEbCJDhmruM5uUxXMbe
4HiPOtVc0qc6Lbb7b76zbQgAe5il2lZuLbcY4K9cEexbkMKDz/7RTCU9IbQy7SI89WWM8LhDCZ8j
Ko03aK/0YkSM7MYH3yT6QkSWKVNFC4r5ebs8n0zeJJ3A/RJct2pR1QucOkJ8hfyi3HDJb1N8s58F
d035H3G4sFDg3HaR9IjJZttV1DOJuGv3WONuoUcni7gaVNKV7YmVLvebP+/ZHmvAQRXJLyMcQF8D
Qck9rVTB/9WIqVoAa7fKasHQfeoRb0YiQVEniTQqnT/EGZrk2GNqYJBSZmPiYP4TUnYGc2bHOAMm
RLRNfHtz0nplTx4Ky2S7RUpFjrl8IayWt5UN5B43U3ldkHsx33Qgp/pNGeTrRDRdREMPZARSZnqT
XqPyZcH/V2yTJ/BXHWjw2OzTD1v3RDvo2ijVAjmbWZUGtTLo0r9cNenDW3rGhJc7uJwkarSCUQ7x
vWS8WEc4C6uuPanYSgwwYFFoVRRze0SkdplcmVd90VeKr5tTahX5+OKg9saaj89L7JVyHGnpaT43
UQ3xewu3ELC2wNGNXJMJ+ZAIztGHYq4Da8guaFse38Gs1JLiAJ4aVcw05cZ1LnqoL1LbtQIf16OG
7TqNcvjD8inY6P+n5DbyQ6j6UH/8WZysT69bnG+gv/LgZFi2lDGEjuDFolD24xIAy9YmmXgG7zCu
R5NibXmw8MYPF7pj0b0oZAh1wwcpPIXPy08839AkfkJZsufZSAbVutFW8Zb7z58D5THLkEBB/+B8
moaFlY+nVGiJGocdIZuhLAZNuCOWHuXTJUW/VzbS1/2+0f3yjPwPuh+Y2C2WYoheg3uXu8GkJ2mm
+sofR3+fj8KMpti+bf8lkc4iGnaPRwId3dFSdAv6udTBVHlujTSDhh1rd/9d9GHV4+wM63V6R0N2
2AYUTTZU1JJdpCM07O2jLYWIpjAwf5Yuu8OWGAlk3bYnrfJljFNQnS/GvCu/WS+NDLsq0y//h3S5
KijieC/kpBOLi/l2KUknFnLtAzd0KBgIkcOeVh55mdf9NgaPQmLmpNXtr3LIYKxl314W+kPY+M/4
frLTV5KaD0wdc1tfHswVirhONI2ngi4pXTzuAZVqqqD2opUfpz4c5pfAarBByzg2R7puFc03t6AZ
YzxfjFPoMHVBdtiFLGr/C2137seHt9vikG4Zmve8JQQaqEBn2xnDJI59NFiwD+vF3bVEUUNGwZii
58rebaWX7lx9oKjytw9KJLrbdasFoiFpu96u1IRABNDGiJTJO+rHMjfE+9biW3oE9yWM/kFRNM0a
M7VvPpBzZSj6a8dvEhjt/+WubhMZL+QCUPGG9eOXwgvqJfYAfQrtgpLTlmwFvxA+mUBleC41oS6v
X1Bxt6KLuJNvEoL889AcovCnT/g+A8aEERZKvfIZjtN/PRK2T/5nJkl1PHEKJS9X6WFhg/M3W+rA
MKckA2fmy6jZXQ3+bmXHX5u5h/U83sUjRsLZsy0oS36jb8Qk2aGLxcRgNPYa70MtfemMgeIQeAtI
wZL7JK/6gUK7KrvXuZ/fVARHaVEwMKQfprBOIpzZazNJqMzwbDibJZgMc/l8COTye6KzCKKffXj6
Icps/VdKG1HkTHbEdAFf9NTn20XWh9hZRlTzGs+Pg0l5I9qMLjdTfxr+lNoKffOU8xafBZd4lvCv
upu5utcSC+Fu3QGKSp3pUjFsb4pXi6lTxkDH/GshvXeP3eyCP7mcKxOYGHvSus01CxjLplMk4m4q
KWHEB+FXpfvpFCMcabzeWli/HLWYS2AQrR3OHTrJ95/jlMmfZ+gN4BoqlCfVVAjgVeznSUSq52ou
UJFsb8dyKyrNntL++rT7WVAzi73pQ4NUJn6kspJb0YpLVGRPZql5p6B062/IS4dIzIAQUj1dePmq
hBlqh/XeMKDkajcElhBVEWjKhSyqUKPWATWiUkUOMdS8LvicpMaFMd4XtUvinyMOhMUT6FaqYvTM
f54AqQbdM6Shu6GgINlpsSie9WOTne8JXhXaxrPMbG1NXp7DOrCPqywHjVTlnmRIm+NlwR2Wc6rZ
nt6bfl8AkXlOVXx55TzFKAvsQuOvJNQN7S5I6eEvs2gvC5y78ozRIqANwZe6rG0VJOcRWSHTA6Lg
9KiBAMVaJS81J34s3hPFZqhfLCHXvCbb2Z12VE7d6QMilpLFH4UoUm4bh/7ZlEqeQX55gd9oy4Iq
C4kLLj8O+X6Bfs8LKbmjpuOG7mdBtry64G50ompj4Ao5qNbMKvEbjOcuu9gtD9cE4LYFqF2qBzSg
W5vH1rE6A1lcEfDYiYRtxcM9avX9InSYx8D29QAkGBBmr8mT7Dx/jZyt3oU7emWm/KbeJsR7HoN/
Kg5wPk1Q4P8lFz5Zg2eEJLHY2MmEfcaKxNCtlRPxCqkhdkyFxOf/VBfsIH2v9KepHPY2wkXAu4xR
m4Hu/QYS9hD+bCKTDAhQQyXraP2mbvCwjnpGBtzdOdPXrfTAX+UiFQD79ciePMfadK+WgdqDlOHZ
IJRJvsuaAKnja5Fk1hvCb8ybhd6HP82yR89IZE5+cZclEMyw+oiFYjcNrTKkJpLmJfqywrns4Bd7
ZiBBSximI7EBggd+4G9aTLuAL5WVYJHJkwsvBpgQ1b0hw+ooDfpyJzZG7myhWmBRYVaGg69Eq9j5
VEQuMTEFu/858WJYJrP8k5MdQuvDca+EoO1RpKrfXnbPOCBUxww5Xh6Kep8MNdWLhpcD3SByZaSa
YbUOAAn7e4FZSCzKfWAaawu3ABbm2pSJOu0lJXQhPGfJz4peFL7WXuR99lmms/3Iw83EZmsK6cLc
bvjkCtlSyAS72cb0MYnX4F+ctcoCH+3niKLpPkXvAfpunIAv8rhbczD5mVzpNr8SPERMGNJHHoEv
84TRAmOMLyijOlAR45PlP7DWUeJ5HVdHOreSz5yPAGvgyMkJwY0rFB6vv2zUjMa+0z0V9mqhJSC2
rQR3AQ+smH/J/9Kor8c41OOylieF3GZrx63cTD1lW3Gq/jiij0HvyMicC2rZdqFi0I4BgTeqtXZV
NZy92NCUIQgiScOlgCHs/LUXpPqx3rQeY9HWkbDWMLwfQdMIxEdO6IOsTSkCfCDR94GQX+APmUHm
trGmiHNAhw+BRUk7Mk+r9TFfnGfbW1odxDuAisxwr67Lo/+LczYBKu0T52o9wRkclowxRdbMtR8N
aAvVIDRf3Yp8Wnf8QokxWQM5HSPVjQM5m5mThIKNL+lyyHWlyVv8Zuz3E9Qv7EerZujJ4e1sMi2j
r4fXlmEuq4S9ckI3eKUx2+AqC7ip/UeNrItdQggWX5qTRf1fL3hbdvruekDSeP6Pztpx8ADTMZ56
edOp6CZ9bJsiBGMDEDzLxDR25cMDQDqo1uN1L5fnWWooP0qZ86xn8NeZwYsNtJGjg0w+irTxfeqW
VAdtBnR1olWLaL4f+UZS1661omRPGWBvODhZeVVIWPf94UifPR8GPq0Gx6u4gNkrGqpkFK7LWLpY
gzL7zjySlUJ6uWxnQ9rCHX9hpGrDv5blA0h4rh4DJVyQvNUiuHL6ZTA6pJO55wqKp3RTXWvUx9wc
X3JEbR60FCyapWgEzUDRh2PfdBOvY86sw9lGHcbLpsBsdtS0P/SH+Bk6iglApATDwbRRLuJabKlY
s+y9gsnYArEK2Cs87x/qJ5u9V5YU6FPlDSD8v8BiTjZguSrDLYNnPek/pHzRcj55RGC+LcFgoAXZ
/nbytyfqFwn5DgAlRd8RxlYJEUDddRjAuz/xYgtLUdbNg/hEWul901O23FqR30yZtxjWoPCIXPPO
TjnnCa3XqU4wAMw3fgm8OJUa21iUjHKLnmvP9f2nihZ60xkWsvsPwnAmuwLxM07h6+hn6SpiLPlL
eqL+0jITSH5clZSpaGm5Zmpr/Lv9j/BuhlVvKg1XxNagZVomO3HBbLFmyhszt5JMPCqCybBgqOJ9
86Awi6wN9rOXzcjGjjb8KWdL4LpDN2Gk4S6u0Puhu82x8xS8Y9zaPCSNPYoabDw2A8yLvns93C+v
/m0k44pXz/77Iww6sP6Y9y4DvVpluGzIWGvVbTgQS+eW2oRb+wXADcmXjPQ+Xf131vxmqFS2OBC3
eoLlJCUtOcYzMWs6qJx6ij/ENG4YqtoYsJ/A4U0hbaFXOZHQoGVLVHMvFQofrjvYfa1WOjCnG/wX
xjnQkQAgWjHgFBR9NGjjT1P9erE5S0vLhY/qOJaEUlQX/iUISQ2aHJ8f1xhQsJ9WFQTbfpz2gipr
BcFLKpznlruIfDdEHajdDJkQOACWOZtNdLamqJlD4O76ARlJEAuWKdloRYmghrUP3Aj0eM83TQfS
PDaMc+LAmmBWmVhsoMZF6rva1LfZXadSuzrFvHHV59Vou9KRD3P8Bmtwc5ikUzCPgpw5BOlRpxap
sYpdB/10kq8UcoGdB9SlwAe7NMM6LCuK23lUlu3Zpb2js+/7MNon4vQ5BvJczq7Kh+67jX4WOY5C
3LJNOaTp9kympdRrA58BVXCr3NmaNDOvoCRkuzBtFM2+YTjHktUFgd4M3TD5posAm5Rwyp9jNCqv
IiReoT7dEO2k4mXsY81XqvNpIFhrX7lngKKmJ03HA0xRMFiMI73ogC0f87kERmSf47YWOxD+ECS+
ccmTKj1xiZLW72o5Q4Ro13+NXqw00Ig/aWTfsjAdQqE7jFqa+3RBVa2PIyyTmxXxJtoxL8w7rBIc
+Ak6VTPQj3Z7l8STi3gzs1kYIe0qPphtWGzrm9pz/3QaSa6z7nyqJKIeFEWQPx1ctKyl/csZvpwS
RA1puPBqXtCSxWbfGv+EBNajpcdDsoQft4RXx0xnpv0Yfi0e1lgncMKIzMOR2WP0KYGDXt7shPN6
Okl/sgUr7iTniHJ2VUUHeO/vzQTXgMLOf1rVV2rURoFIS+8NvkcIw26FMLNlJrfh1OSlrexntLge
sHCiHzcf4ym3xtSJUzIWjQgqEAoTxzvKNjYMe34kNffvzGRxYuwUEVGgsDZe/AEmoHk59d/moomd
cgHFoZbfVFCCF4DOtT6LSAXXT97s7yNXq6DD3kNGzJYDYXUyK9/8cr91dqmO8NJEGJxuR78l4Q7u
tNQ9Cu8/4v6Si1j1z0SpR/NFIaPGAOd1qik6Kclc52Ln4MlRMEf7ANx5xPIrO7PSeCKYqSVz6HQg
lRfuKTo8/GwRLCLF4xX1vJrUkjYkeQAa1WQMR1CggSw5cneWsjOLaWrSq4t+bSUjUkGsxz49talw
6QIbTF/V5KAAuo4JM0IlVS+3uSrVI55hKPnDU82bs2Vyduxg7Wg5bV6BpNLm4sXeYy/SqTmZT4XG
yVA126Ro8nsuVKIl32OOlhZMzFmSi2MrPpiy+7C3QD/BZYMJ2eNjemKiJF34EFosv50Z8LqRAqCa
eCEB2hxgPYQcXZiVmJt03zFi0l5z6/dRLk+GLQP5ugUmvF2bRaEbV1jFCyaq6yvRJbL0K2JLXCpA
C4E+0LM71qfp4GqDekWY0NddsMl9H941YESxtAwyIP3+k4P5mmu16dEw/ZAwNKU0Wy2AG4wNCspN
NJgPlfxIhKlcYtXqe83vtYtBBbAFU94+n8DBN/QXDuRbOSgLEwbJOwGHlvjLS52SIz8LFdkvYeA4
rJ+6I08joKZmqHGIHzu/EwbrhepAAbJw2CsyyAEVg7hdinSfLMkJoCPKaTwVQrfSuS1LJpVFgXLm
j1wgSoYJyVulPeio4UCdrIVakD8eZ/p1AgKmutd2T5lFdwHWvj1bni6GgBQG8J/qWrwRvcITtDPk
L9cs2hIEb37YPHtEzv95dcI9gLmilkuq//UAjDu+Q4TIp4ZZd/oehumHTeMeKUwIZgTwBxFfQ0cD
ZkL1lyL7L52YYxyb+ZpPMx2Td8GGIIxmGNuA3NR90aOpzOXIcYRI/XJ8D8+zbcSaisDyzmc+/16T
61QK8YNf3UVxQWH9QUITFMNndtqNyAckMbND7PtGhalDabCxS5f31L08yGzINks9q/R6ocF0DDq2
NcuqaeCHIqCBY/KwU08w/IOuP0aD/uKAhGNelLmIfmLHaU+AgbDmRrlIoDPz/kxDGb7G4nHl+y7T
XCNY8Dxjn9/94lmRkMljf6iU8UhiFUZSazQAND3l+zKxRG/C8YddspO74aIO/4eyem+OjEjX8CjD
iUfE/u9oRj9LxS7VNXh6emVHmCxPOItrpTJZB+JlID+Y1b7VQGJWehMmqHgV7nOFQbkmMJ7DpAIS
+OdYuXcNbtpxXBhK4DzbG+TKLc9YadS7X+qldnRjykeJUN8jKhfF3eq4SV1axhg4KmJqKjhDvBBK
+3Aa8UAkzd2HFYR4aBbV9bYk4sLC07UZcyqdCy1ysx2cxEiJjOetAndzTLTP1ufJgYmGE/uncj2m
kC/DfYkVUFS3MKx5RujKJFj4L/CUzwkeJygyVFZkFSP9XXnLsnaLmOyRu/HlhuyNWB7GDcXQpiB9
vyVIkUsBur4q7g/bpIdcK2rz/SHH2x00GOZehZvMxq0wA/GD7tw+knI8GX1aTHuEGNDumB5SgasQ
IDoL2yiOphr1wtRoBfGu3kF5m9jZtUyL9Y1iswCxwAuzNXUG7DB1DYlE5hTWQyovvaed82BNiA1y
EjoqWzTCJd+u0Zxk70Y+U+hktRadST37P+PxPyNLs1kgtvjHXyVmnvovSjZ+meAacPFNUcoh4YJ2
j5CsdAobH1cEwZwWWUXu1WGKCoCD60xHW5iQki8XbylnZvVAe3jnvUuYwyPo0GJSu0FoqnGcbYWK
1llFBODtZBL+s0KEqIK1mgZIjHKmx0PsGrQ14ODafNy62X43KBD1uehBDt+s0A1aoikbP2ZInHep
T/RI53HiNCq4u6PfutH74Klw8sYd1wHAmp6IehwesAL02niUDxh2fNIYxx78htA7jIKFuBC3+QZJ
nvPsntsSUZ3+RzEaOiCtLmy3EmY705VTpP9Drma21mfoX4jn40+gDFcijOm5JhfTnJzfFfctNGcz
4jPW8W6r7SG7Jo7tX7dTCmMMGxknTUKjzea7E2JHbgug4Nhdlf0XJb3ZqWcUiVh7tcPv1ilnLB5e
9gNlVWxHLI808lD9s5RUalJlpHqg4TZJLZ7focZ30PmW2EjUqJuHKw7+iRr3t37wQSk+vcHnaUl3
UBwBye4PTHSV0xNjIPgWX3bklmGPWf2KGAq3F7Nj/e4Ivp0kRJVbf2vmhA/UBX/JfzEg9H1ltWPR
G/VRZg38SwgWX9jVlBvoj0a2C4FUKZkvesiTPrISAxoKxceVYggendeAvr6MaH7WA+RPrIGpofbK
anuBoH8tbCgdoVQcm4nZiO9iHyEmSyNwykqQebRwS489f/5iGCdiSMaxNLFVAl059EkX1FXGeC5E
c4xezbT1a8DUDpIuiEhd81mHvKSfrSAnG8tepURTwGrrbGyIjH4PLoPitQ5c4Wzm1pzJApaqV2E3
BTXlVF3DKoVDvObmrAacRiTOKE/fdCX33rRJMqm+BsZ8Kmv6vyzJYQQGLkT0M0tgndmRmfgJmGEl
+VF+sdn/DSNcMGVHiHXIrZ1j9jmRZInG+2AQKTRE7L3QthDm18ON3LyQ007blMN20Sz9p9WRgNk2
5ZUplIAo3WOAr/1masUT4suOnB1OthS0VjCa0O2gXhfLkBk4i7mfEDseVySHGfx5KX/r4KXIw/rX
26yI/Fs53u9CXs9h+wEuRL+qaGWx1mGR/N4KwzeT4qTncm/tKmgbdV8y95/4YqKMR3B0nauC2Xd+
eC6xjnbCRAWtZjyvQeBRlXDCzaAF9w5mA2QGHE1cq/BRGVxEAQs/xVnrGRxbLUhxY1hFZumnFuah
nOxdRN1enXllRAioIvMCATjZcbRrt2KZYPSE7KcRVnrjXn3c5ZjcnyPBIqzFjHxy6SWkZBDjUi09
cA53+PA4DChjWxgfs13vIop+t87EliIA9GXtFnHGZl7t+UXWkY/jcr1yEnq95aLsrjP2X35PooNY
tzHgrtrOrJGdG1D1Ydhv2pkXCP3zWhbUAdI2FI58AcX7aJ0A17MdS6CmWhXI8QX5/OSzHP0s9PrS
zlBtgfdlKmKupBBYAyuKMoXJueqprYdMMFw+VbGIkQIVU+/j3jWbL8mMPIo33mS+jX+Cal5n+ef8
yTN3EI/Cz6OxLt4v/ZtjQvNR0F5bPvSsID59l6a4OVmcGB//jaipu1okAtDuq++xU7E4XbM0lCK5
Ff6inBhaxg8frsEoFhMGkrkqW9YjoOfhwa21Iz07AU+yUcdeIQfmu+FxobWolqMR0d2ibdkFn3v3
J+Vmjl3SEBH91Uhi4BgdlvQj6KaDOfQVJbJ1ul5eySDECkoMZAACAENbIkNOqyoOG2kaN8dD57lJ
dK44amvJgPTCNlIVIAcvkcNiabxEmE4O6iovROUjngXcEpGjxLHbWfWWGUmYd9Qyq3lJm/l6M2bZ
QqbwNXcCeXLEPfLr6s6kETSRKGtRZBFEtbEegkoNaoLiZ+2TnVvw2y9ZcWxpqyZl9cMeqmPia7RY
ilzjcz7T23pFPbKV9N3WEXqOwTLQkEqmUBFuoC3Ef+z6Ruz6CSzHJsJyoC2EOUuLqJ5khZs7y5WP
9So31ZcsyJBP6tpfyyeknchBE9AGyrjHzPbv2V/hqUzaSSiDHl8d4IPQjiU3hANdSrvYsen669Q/
zmTYgS9jhhy85NomKVpfnPCUSiJ0NkCKOxo8qPXi5UjQ0mM+uY/7x7PNVKBWnzLw7NWiOWz/b48n
dcIHdLq7LqKsHtZL6pSDUNpOIVPQs8UvjqskHOAICrdZ4rvVcyVZzzwzJwi9t8K/tDhVVs6RddyQ
ih8EJr5A6fW+3jxvoldecZtDoz2gK/jFNxWZc9QehuGCMAgOxK8YMq9C7JaUXtHdmgqH3OO/m4cO
+OWyzl7EYyiRIWTDZgVlR5PvXUgmkQ2fJQORBCwsgHOE/CLtRMCk3HCb8+JbsoV8S9a0SrTjFrUT
TQFIy0bs0E0+F81y5WmXkp2/CH51cp3PhbVszmePgqEvIPZ64spxdmorvAflBDISd985LyGMk+Es
0CoqUixoov7NiO8XO6K3zIglDFBlRLp/R5Tt99DxRL78Lx4uLBnfZDbzDmd/sJwZe3co1YNf/5sL
8YUVpd3gcfH5q/BWHYQ/9yUc9AwCg7ItTxG44od/PnOzqWmq3JZrhUkfjT35ez3k0dkWBBxSqzjC
HI0hG9ypA5DO858OCiySoU/hxre/+yjrMavNzGwyokmStiJ8fusRwKr+k72dMGscLMOaLYmEma0o
Q3rpM/6p52A94gk5D23fBatzVbhbyjf4KTZ3YNKiURi2GM7nj/MzL6B8GE7oa2ar+1so0DfM6JSR
JXGaD5SjSwlE3hdxqzNm4O+dlAfs6JiRsN8tX3UCdofeJDjHlU/7NaTiwIhHl8KVX9vkyS5SOq0c
iq9ZZ/kuKukl6j8mf9Al1FwZE/BQYB75ujGYSdf4REkhPzbr90VJTAOrbyJZn/aGcJTHJfdBqKDu
CA3jmUxno0kIoP9OKhOME07t3XoC97botKqyRo5ddrMnNXnqNUgdVDpBrv2dMKI3er9izG4V5nbr
XYqtRWcCWRjkuhPa7OW63dbRl0kVGeMud0oSB6p7k0rg6StK68UJXOhoHivT2/id3TRYNllp3rC2
o4X9N6a0VRDgZaHGEVFGNmzE3Tfpxnu3/v4fJillNnq6Ld1olFAW7JwDSJ8eQe0VXiy46+XzrZ1M
E30en51BYW2QXG4EtG7pV3aZAhTeLzZSUd4tmLpPyTkf/LpnBN8qPmBTt3OM+elbSSXdLiLB2cFY
mjWmg4VIVmUZPsULDCTGO2/yyp9gwAVSu/JU1jnHSZj0JJUKiZa0BkdSFRuZHbQwetaEDKQLSH6J
d801WPpGhZ0mbtxX8t3J8kYG4RI7kfANrqLvFbMCoRQysX8fHzIKpqQuTE4v+guU/gtSUc6dq6Ma
jwGxo4qz7XMZQcZg5g8AGJXz28fA2X+3V4k7gxizsomI0M42lYmw86HR3KzkMmRpnV7g2ry6bTwp
s+Lc8VLyYsySzlXNWyo43yr39I2Dl9JpMiaUdO3rBjqURnXaA5pvYQzXwK2XugEVEB1esZZGvFBs
pFKDMxQ1JTmoSz2obFLF8LqPwRv5yitwHFm6O9N1Baw4TLpmUTiwyWdXySf0w/8Yi9t2gRToQO6Q
Q8+vuNB2ubAsGNDPJetxzTCJoRWNUlFgajk5Iyt9tsw6An8IlMgEjkVbC5XT/oazbTxVIYNf0Vjt
KLMFMsbCLdJXJQ2jYMYYLdz/onbN1r9ep63+opXX0OzUeXHubuyJCPShOAjuGaEuepRKJZ3v2U02
9tXHP5EWuWyIKUSudWJK2YIw31Dl9nC7sMcBurLQL0wumwTPb8pJkpkYYcNVR+PseAgsvuaYQwQD
azaLYYGhdboAPzWGSK7ZII+5iI3y9hzK8rglmjj/c2pWXCRruMaKOd5RvjBgYa2A6LR7Wv5BkH8W
I/EN0YcMOqR7NpeG8TSLLfx4RTS3I+EcH8LEH8aRSBDWJEmYNf3CPNFq3kUF6hIPcXnYsm6YYWyM
NxjI2NC7DlzXRuvlaFL6PeUlpzlwD0h84K9W1Gq6B4aGkd5U95MPM/LJqomoedSfzjvF2YvUR6Lf
0j7oij+cIIhOd0V8HRt2Q/W6vGOZEdI3OfMNCaoQDuiwh4DihzYpQryhlbAlV/VBy2p5h/9ve3Gd
eNnzt+JhPR6oktdmEw==
`protect end_protected

