

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HZg7J1eicTLULECaPz6ctaw8y1kpWgApgtfn3Q+zYY0GMZZHrstjvvtt0rjShEIyHEmHswkTon9F
uInqopAFVg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
L2/HzTdtpI+DDWwQZLtw6a20VAniDvlrZ5k0iYB4G3h22Zth0ONh9GaVxdnh5RvsADtDStl24FLn
89acqSnMq2//5lAdWAp/jsSUiUTqUuq3s51XcviRecb87oOU+8iTczHYM6EqTAd3Utr3aKQ7HiMo
3WL0mQVpCBOpCQUD6jI=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OUJeS1bwtebGQThLvBFH3PwBsgx/p0nU2VJ+e9SC+Hrio/pbJwz4o2xpS2Z63xJ7QN7VhCBN12gu
ZFY5Ng2Sgl6wTkLeA9Vhfi5uJY35hY1D9sWB0j7MhUUJxRIFWIWs+H/FElpBvWn/H5UtcrDSuhP2
nLymA6ruYrGfx7a8Iq4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AkdqgHhBI+1kEGsbiaO9eH2SWpUOBQkGBwaPxgDJYtBsJdOF2T3rxHzMH8aRRo4rOV4wq7F5qDYZ
2bRKyZlKyXwxOIrgHQ/aFSyCdbfrrJedXNOvayf3bMLKWGvmkeKTZFG4ie8bYq1NlzxjEK5tXh5u
do6EoDDl64fqmvjtPSKx4xrYKjkfDGC1J+lF3Ws5x3iNXrNkIqRirBHfL2nwSIIbCGtaZ+SRJZcG
6fOBaI5sglgjVMndkM1UDvQGQg1m7SekmV1gNbuTjfVG4yDcoHwJCq9TChQTCfG05c2xR2kyrVm4
vPlYfKMD9L7sptBiihT7k+285Lhb3gyxkn+LZA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kU/KxTFv88aIggtPFaqaw71mguuPJV+CvKI8SqHLyiEfFwnEl2rRaQjfKPPKVY+a9ar3+m1VrJZq
XyAytb5FrHwHwKJ8PWa7bc9KeMqYCg0WQyqVAR20oTRysvr0JW9ZU5xcZQIfn1WQOAidCGjGERXk
D8J1Mok2babDuVuQ1k1BLyAGty6ATMVk3dUAR5LIplcmY2dcgXHhvtTjcDGgu02ufeeeQgDtYdEr
XxPaZ/IuZu3RKlqS+LyaN7GLtQ1sl1FVJL4oxiYEefZ24cov5R/2KmrDI47bvcitqcxarcKhbIwt
EegxbadS43xqD9JDNFUAaaCu542z6SRuS0zC4g==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
k6DApHKykfoAVe03+cLJSaTvIyV2mgyg0ee9r8sDTCqvO5kwFuomMl0B0cjUO/4j7+8GeD0YVUGW
M2t6DJMbIxuNlNctJRXzSjxwlBu2lOTLqWCd5V9OOHutCH8JEU8ndSXTE8ecj8B3ICDoE/uYntN5
p9eeS5YN3Awwuuf7vpsiQrcsy5iqvO8GW2b0InrBhe5m2bb+CK00dsnS6RTA0bU4RH+b9zcISWyN
JJFEeDryWX5A5kyBX+Em8sHpW9ssoOlBZUuAR6sGhqbdC9endcp3vkYasFpW89RPhQcAE2DOJVLu
qXK6y8bpxJSgUq7bdln2TJUwnHb0mgJEbAKlHg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 114672)
`protect data_block
pxeBj+oH7HiLAFExL0g5WEZ4yLpBBupIX6FuMPMN7xUnxPzKscv02hePml+mZYHSmjhtVjLYt5AJ
1Q4hXSuwKYKijAgPSbuYwPq/zhSG8u7mr1qvTw4aK0pEHtQgihRK0o0/dl3wSBPnI3kEa3dgPJcq
vwyZx9DauAE9fhrO3m3PRo/RTVa4zIx4CIgtbEC0R5OJ2DIW2ZqErHyRhwRsajz76TbOxtuc5rXi
5otPzAn7y3puXmbT+xv0QjkS514dt2ReHxc/Qz9FfPUBrbIAxoniiYInxOzAqVhIwpSWxcORPUyG
T9G609YgdbNdWMw6poF+i04JJqUBoU0sZ5VfuPePAEmpR4HDQA9mrOrBpT/s79DNiLK11D7Z1kYw
RO6z9Ver3yoltbm3vVGe4tH022kocnocLHRBI/kAupEmUbXLjP0/T9IWnLsrEn+B0V2m7iDDiFlJ
gDa1WATYB45nUK75k89lD1p3rTl/i73Rb69CpxWx3cm9GCteRZ02Yl/qx1dSx7nryfuyIuATfR8K
WEMxZBeIdZFmWEkVhcg0Jjy4qbYHJwaK4KiMtLfVw0RtwOM/y9p4H8Vk1S6VQ6w1TpVjXl4SF+is
PrOFV6nKjKm3wEUDFbF8a5gs5f+eRg3dUqhwi02b8Coh9n8uTognJUAsLHzaSACw50RnB2fR2U5q
dy+9EWL6/hOeyJH2vRanG8XTSFHr2yHGAUrEL5J6PzZjM7jc69E4skouSJT3aC6pVH8h8O5yB0Oq
3pMAoaSXoy6NFrd01B8T5IVWOUxPBqoqpZ0a1qUOtojAxpDwSy4lR9QFja+36NVlQOivwTlpHNjx
h9QngTwFv/D6U+ayhciUsF4n+9qZsZ550+/VLlDPv0MB0y3/5DoEJS8tK6GEvQjQPUAnkJcV0bOi
HyZgaRiGvvDSUxbXK6x41iY0RfjzGNFW2ybkq458IjjmzGHF9rlJ3WTAshLejtgivw+SzBoE6uyM
rivNraVl1UVtPg5a9ysAVtakWEq3baaQ/6zF+Q9gGgP35V2VI4h0AuqGhvYMCMQG7xNKIiM6kTS8
1uYW4nhyCxDolIV8mxaSBLe7J5xhvF6muO/tOV9SguVtHNZa4DfLlaD+KF3Ga1aI8XkaQPeYgLkv
Z/AKVek/COjDOiTc6jlKvWePrDSSaRMfEuRgiF9MpWNed5FR0PORpWs8hXRBwboKV/8rBjYwOI52
3dZPGk9WidhrR5nYqEtFMufxE2T7arW5q6VHZ1dobQtzXLLwJQhmS1utIeprABwH+bujLuRFnlk8
2Vio/5W3wRT2VClS1wEwDDabJp8sRyciMA+urmjXVzxlU5u81Om4XWvvGlSC/KPx54nuUsxmNvFo
nIlvqBIsDrdi4Q3sq6ba+/3Q8P5skxEgE8xS+FcuKzP8Xrft+4ryb/T8FCXAVJti8m0iQ5i5AqlP
oeUtFwYThW7JB+2uiFDS7IZtY0Cq8PNgeenwqrvy9iVk5lyzJIA9guXvY9934YJ4TkVo5WHLKIfO
42sNkRMqUwR3/sB+GYFDGh5kuds78Ir9NeqReDIH3WkVuzOukgTtYdcCMfm7pJicarbBLyLwVqde
iIJiKKF0+WtQNArCU7tKCSY+sDEZ4nEYwi2HdKHFwcs1caGnyU/JbfwUK/STWp4rMAW5mZHAnCMl
inKUsjU7bE55TgEELO36HvdqOVnvGRUAT9+9nM5GLaUV3kO17ZIZ0CVCFJVgcT2YRp829QO05LhA
I3ccsGX/OwtvShyQaMQEWuEm0Tu7AXVUxsLRcwl+MXezJ/zVB25YKhnxBv6ZabAov+Neyx92QeV6
kHsK6DUMziczzpogAAUi/wTpTWm3DYz9/7QhVjs/b3ulsvgINrFUgfVwH94GaK8/0jbAw4dWe9cd
KF+oGijsZG1sxOwXGqRyRMO1PGbMDpfCZlkaLoaeoAr2SHAtaCa4SmNtECiJ9DPwj1PgN+ceg+ZY
C8tdzgLu5fs9gBDuIURXBsRFpSs+hCvDQsExrGhK1tP0BDsDrvg+Nri5Oa2+cVHuohyvyi8feT3J
wydESxokcdFip6Oi8xK8Q9BZfaU+OpsckxdcDxZMk4Feumov79wYGGB57aYUj7OynPVOkEFOMMBe
I/RB7UhExJewWXAcBqGDbkpVzbsfelHsgbNtMj+PYZ6m0QSsjTyOMDqSL+06ipDY5gW5Cq8UQBcw
0CUctANV7wm67Ojs18bqVx0exHdV3jCGYGvYyFSVAO24Ig4abTKqorxGwcvblt1P+yD8XR2h5isK
g+4dQ9D2LFJrPfy7uWMN2nVvtJs6DNwHe02Ihf7Mmar7hyBaYoCupN90oQWuTKQHtUorKYqxTO3K
NaXQ0EN84GLHo14CHWx7V3IZqQyZlTIjs0kXA7v7uM7uKxzynOH9Va9115oPLfI4rpajq9PVyhxa
XRHUw3E63m+VUXUNluAQkg/RTvmu1yp01P5d8AFXvdoBxuk+DKBtO1lnGf1lGoI/hBTZvGYK5onA
QqYgQSRkgreCPEKkIFA2/TnjKve9QpQ6AO0igMqi13PaYLGLwBSmHTkLuBZEuFPcDpXwp9DvLNeN
F1p0C/xd5QTK2vzS6YTL4b+q+CSuVacY5m4EYuoBgjamyhG1FQsQxJsYlUBhwhonvxPPDEZXkikF
p9bxryn51pXFr1aXMy45P1Fu4e3G9gHHm1xAMNOyOmGFr1/pcLUMYf3LSu4WC+EiRz5o49Ch8UNi
Ifh8Ep+Keiio/7gC13BR6dndnod+YQqSzwkaSIinviEfAmCKjtC/TbyFWdbW5bJUYGQbFGe/yon6
L46zq21qXmNqnOhR5n1VpGnFt7nZf7mbaF9/zhujuvN81QqZLzoCQyK9NT4ucUIumIMOvtSe/M4Y
oiI3x02nF3ty7hUUIRem39nZBz1gpOre4UxhGBjISjCokC+KR4WVp+SFbqOUrDSv+vbL+h72905/
lXyZPVk03Bx01T82AFQM6Pmyh1/E7cU0CgIGzZLTrSr77n4WJznr/5+Jnnr5p+emD44Tj95RGysd
A2IJ9dyI7TvLgh4H7ig68AjKT85f9vDyyBuVhGlTJu+Edlf0Vu/WZ7I13X8NCMLDRCJWdQ0kYagO
t2xjE+G4usfGHcvkgLvXc36hbWAp2cl+0hKijmLrjFPz5PkEthGCcNGM9qrO2h3wIyc0cKA/VkAf
QizMEG6m3ekjjIa0/+fWeTsEigOpMWP+pVf6qDsT6S/sgBlbrPOLAOrDXut6iLu+gfmhlpQ4Xc+3
iMQwySjBFJ7FHFDQPl9Bvcl6sD2OJLRjarP62p7NeJrFjddpUoHEfhiDinmuaeu7iKq2lvkPSRGZ
laN5L/a2VFC/i0G8TnSDunlODzWXA+J5ArNdceay42OG6sgi7f2TCxasJgUgFISH6sCpHQ8o+m+V
AifYH//EH6oNxcFQ1z4c6vTfXqyumaQ3WYWmeW5CDRKZQD8DE0skQ+FbtTsX7WqxGhW8FSyFcK1Z
BWRNKY8I1+poDl4Djb+4smGZebF8upyRTB0CJ7U0yOVr+c0gHuymh+nzQvbnTxzE3Ld9KMaN+Hvz
gE+7Af31kg+iRRtlP5Dx82jCbZY6KUehWfaCjKazvzzMBNKgQjDAMDVL9xCXRGQ2YXehqhZz5SWJ
RVJz6Z2sQNsO80NaHBo9GDAoC2mUksCbJEwsrVj5fa+rcTwI6rwqG/sRhQVZKpFnk66yJQ/7d4V1
VC0F2ww0kjidd1u/k7NXyhPRKusPmIHV40Zs/kqo09TkQ560Y7RIBG+tOoKw5++DTO5RT3/MzZga
h6nRHydg5IYb286nO5HSbAG5fWZ0+vTFYEOwlLD3mUWyKR7/cQeUgUqKN4T7VLlxYXQkxwwfB+NG
pRaORMgaX45VrMC+VOz5TF4vmmal0FEAniTQBYaLkc6Zh+FMPbp3FjXLKx2811L69ggBgFqNtL/1
Po0ZEViO9iuj9B3id1Xabh60YSeWh0XKZFe36KhMQHuGbTGt6SuH44mju2qcEFANIsLoo4IdkFXx
dFgOz6G79Njd+CYLqbokYwhKXQxCo81nDlMLPeyOolry4nSkdgDbkgxmq85oiRcYZa5nkesV0Gmg
BWdN0wXOuYmSYYcTBEPOEHP752vu8BgRp5MUzqzd9zuyYe0HbN29tcK/ROWDsCnhXNCnXGZQTFvV
aEgLGfmQsUuYeLriJAzM8+QJtRqmFVSJH9HZ1ljcKjM8eNJH03MMzpR3/gigXAdkooHdqNeE7U8w
YdWDCHPOQ4Uh9x/ZvH8rMqk2l2vUVflqYPMQpa+40+KP7ds2ibJWjkfN+33Crz+FSb2hAWCkUPcC
jUheQ1rZaRIiRLl4KL0NgQBvd9lQBHMzxq2cV3RF06CdRyakUtHI4vD7HpNbLuJDqTOngocp9hJZ
oZ/UXIFWbief7Ig/gqs9EX0O1ie8nwNkRc+kmWgff4TFO452EkZ9Djtj2aRMx8Pys5knljQqMyjV
R/At/M4uoonp7wjW3Ah7rqssSCes9OUA/AwASJnaj6Mb5Y6T/a6l79KU0mIyxoGiVXczdDY1NA43
196zpinnRwU6SFzhhIfBPg7EI4C5pH8mnZqWv9cMgPvZukOmV4GwJJzI0kDdozEi44UXTlqeCveY
tMxr2RABkrT6y2G8Kwvc+4eNtZNyOXyJ5XNraJIsBLJpWOrx+9rTczai0dPlq/jeTX+LQBhw2BDF
S2h/2An3EgFpkEmmC8gel0e0LJITNQKo5pO8Ege6pv2szaYNLGoWX/tS/+iUi0UFZfsA88U0Ixck
9N0eMFwiFWDypW7BxXFWwEVn5zcSOBcSCAAeZI+LWRFN+9HPEmpps02VwhHgDBV2eoSrqyMDg/ef
myTFWnOKNMQbMVV50BBei91DOy1v7VDYYluyyHwrA4FjQm4tNbZyxAoRDjWOYaVHZocHvuI8tkJp
/nzfXEzaDGE2NyQ8ivC2naZKd80Rmsvf1cIXUo4wo22CPyp3eqPbI3X4CmkLTc/gKpuQHyg+cUWy
pprAFPqwnpTrDhXUssBcehxqUyzjZuaLe4I5g92oi//UatoU4KiaQtHB9yT+ntt12n+30P3bnVHA
16p0qN8+PUL8LXMnmWpNzKnWYBz95N97uGfeibkgc3FazmwlrEVIu6nJTtbopLBoyoU/GNWPIRfq
w8x6URZKmS5ri+1F8uTYze5pXu3j8oQZrSZ07dn4CQZtKtVLBnOgD9tOFVOKhuaX15kIk2rrYz3L
f+1YoSEUzTmZyzjEuJdxe0HBo7qk0mZoZzUad7+J8U871drddDsXn39IOkp/bmMHtrxKVW1hqQ6M
tOMYAQXhG3v5du2I1GJ3+lRl2NegkxEla4KNSCKKc3QDt9TvAbZ250cBRm6IOV1xLG1DLt6lZ6K2
WxgqLWnuFpcO1ddiaxxvlNpWZi/EdDuzhoOQcun7Hps173NbdpJ1AnkI8KbTkMz18AgyayLuGq3D
bxiGyzRYA9vBViEMV+03HMseIja7XyQkQO2ToZ4hrBpJQloa9LhWfNHpTOk1hhEkz677y3GoUKsK
iLTtNz0OPSyz1J2ziCIWGfSfylDCkTRSjQLhnyvy51arhlkQCCZMsSVZfakFZh9ZHPi8/vdYkjjQ
YydzI+nVkYzSVvt4vnH5sY8zS/yk5PB3rJUDVF/P7bivhVCO4QYZWtdf4LN9pzwWwTm48zJHBSah
IhaBkz5NpC5SgJW5TCd//WG5F2XJwwI+gYNOdIlxFgfGU/B71wHdvUIROuhLmJN4pLmpnMT9MhOx
mZ2HpcdsX/GR64GxzwrrJLAu7CbTZnN5SKaM/h990Agmw2/bm0AcfrU7gPPgX8GN6MSffkBcWjZf
cIIM6ZIP+0ZiTGibeXR5e0EzVEW/X9HeXDh87axzvDhJ6PqHsyUblEotBq9tGRUXvYgUqHDksJQQ
qWc4mkcxYvdmmsGBDl03FsB/5R1acHqRJp3mGHU7nRZLqMubFwr0EV6l0pU4ZCGKwnjS0MEoSlwS
NhzD41NaFtQzzqIrBqg9Ss8mVhtehT8BdqcgxQHmNXdG5a1RE7jryG34dUHpHham1aDTqTxef6hr
sGNIcTb09YlxtSHyyEiJce254YReRFz08XStNAuUU1W1EcDIkfszous7Udc3ocnvxF40buWUPTX2
ZpApDnIVt6VvG6tfmZRgGZW7iM7TH34iKECa82fHoSwsejnNbWOm+g8bVKzDcrqhB4ylhPzvBrmD
lVz5UPGP7m7iWNbSf50KINgEdnPMKbtn+8VqB45SMvuJvnH3R6C13J3h/ITHNX0uFh/Y31KPtdwb
EXcsjZwfD9Qse5p5kZHSI1K0wBj1R8L/6l5Z8sQ5huMp/wils1yTZkgmRv7+LHHhnxoSDgmSI66y
LXH0cr606R63hF1pOv5zHEFcIknMM6IFUB/D+RqVAAT/KwU8t+PBS9EpFAFrNnoLrzUUSUTHFLuj
SbElpe7z2RJX5tMjtmAAAmDrI27zGjJVr3VA5bdx1+vZdXNEZUex5Wqr+Ab6bDPLlUoYo2YKZKIN
9mLmUvArR3zlST6r2ZuREhAnIWaYS1Rgja4iQcZTBpo9vh23j4SamsII0iTRtvDdUPrJAhYGYA4O
e7lHRBG+GZtwgg5bLFB3ahnFyuwncxciMs7IdOeOlL/Gyallxi+CLjtar+fxT10mZ7Xlwn6zjJeZ
NAvGzf3P4b3sCFConWCH5Z4XzOEnFfSfMcjBAHxrB8hmcwLl2lQofmeFrgOngt2Ob7SFQVUZcOZ1
VH+nGCsqbS8rRtFk7VGRtgunVbakze61VBHikn3DfgKan4G5cm7xvRfkJJn3lI8+G23OT6Aq7lXU
lw9S5nxD9EcokfzX8qwQv5xn33Ebxc9DaPgbfERbxgaYEoQ4yNwIHWjoFNQtqYd/nDiG44ZzZkLr
oQTQSKnJZHDMVhtI6Vmc010gHxjFLjL0jpHummFNwBnoCLaAr2yoqlXjfWjlBwL2paVZSClsuwYS
FaitqJsnMkaxpLrScqb07ra06qkKYEawzjNlmDG99oyYhf3iIpQwtU6sP4uhW0geh8LsiBiGXV/q
Acv65/KJtpxqcdiMsKr3eaB6q0Tk0wRTqWnus+Irl63Ott1m+tL1UnELtcZKJfQ6zfbJzNhhAGkO
+gR2LUmh3p1Y8vlSBozQgxbYLX/Dvk7nSbXa6wtuKVz1GQ3x98vJBJpCBPc4PDi8B/vhotaFlQaT
PEMYQThkQxrsuA0bJCklr1fIlGhgCnWXXr0KFhEZA7fLNf31iy4i1jj8e59ZXDHb8munFEpK++w+
+WliQcxVcPVLZJ9kog+iBcA3aMj3EtkLQPQpc3aq9Mx87aiMnV8Jk6VJluJ1B9bihiI2NlHOpkvy
3q7jlmaYgb4itsVg+AhEl8QXABIybc6EZNU/HPGXMR3W8Pfce85vXWwRMZhIqrXxGqRpBOMfuTwA
4FIoUNCaD+5GYbIuFwHJqK38den6OMEhE/VduS9+w8uG96mo3Too6oFO03O9vu/SFackdWaxtZhi
sgazkzVSCAeSZO+frXpQGBjuTDcNzRzwpb78iSO6d8C7EcJaLg/pn7Jk5nRCamwSSlsIO/g/GqsU
84Fsg6MrKYqNIgiXilf4djk6K44cMFzM7dTaK6C5M3VlzMbqccQBkV2Mmsm8MFdoYN5P1weUZJnS
EEgp9sscYVOc6pj6fWT0BM7tUCVk+/9g1+iIBX/Emo3yhJyvlSAr0nfQvkK08LB4hjtOWYBCRMHo
qiI9ASzVNAtpOx2wPiADFWx++YRO6vg7EvSyY+0sZDCKY9AxFDPjqJtqpSfT6LVkkAHmeBIZO1d4
WRAKdnPgVTBQvvKKNyG2x1CzMUnGPs/74u+yNpYUT3Gigbmiuzq2gwR6N9egTe8QsFojEOmpjvq9
PslcA0G4yUF6W+Q4w9OjIbHRjifTR6qx6K091LbwPRrTOYgoVz8pT3zsE3P8yonLlNTfvCDG0lcL
hLHBmp6usKqFSlm/seXhiGO7U8fGjEy92AsSFkfRZ+R8LzfYRH5dJzW2BhJQuC/LVWk+SfkImach
EP6lBggC03HDSzLClL9Q6QWaMl7u+dYzMkijvCvHQ0XmkB2It8nsZQYUU/gaaIHrM/2mVIP+nmgf
2fD8s09QZ72+Gpo/18VMdHUmoNmpvy6lqA/dqH05URkSMOTAJynRp/G6BgAQRXfjp+ZrJ9ZjxDT7
4oonh+MXnJQd4So26IpISlD1T/uOKcc7Z6COhQuSvMGwK7JlcdcNcPS2DnmPMWnw8ZIS+pVxDFya
WSVD52bVAjvkZsq5tbpNhxrvTP73MOJc2RWNiwCCXrLt6+1GNgfHwFspYr1+Emg9hcL+x3O9jz21
TrcB4LJaW9Ky1wleUDPf4R7BAxxneTa5UwlKlzdFqQcDMcOQ2RYGiUAng19H5XPewChBdvekI0j+
vSXp8zbXa2yaih0XEM7lzRzsiajV/Kgm3msw5X6/F/Z7kvrc3mZI9EM8UNB03CJ2hLOdzmEayc5v
T+BYGzWL+08bj2OjfAPpETxcqU+D3Gej74kh9DTVTELmCJbVg+oGzfiCMVyXpEsW5dzhIdP56oSZ
LCIBdhBi101ibDVLZUWWV+wJ9pICH6HYg4OE4mJJcejNDlGBti4adO6Om5G+tnau1njJfOIx70s2
4vQvw1mAy2i9B8hE9xGKyw2cbg15Dr5d8pBrHETyapabE+9swasAgGUSCOCiAAWssyuhEWQJ+B/F
eQyVBg04j8VPacXHSoMzhKrJ/EJDBlyao/UkSsoID/A4uVFHywHeE3JHojbwjQXJ1hMo5EDZFEaV
wh032XKMC9jICbwZSX2Hv1+S8lvc24pJXazdtW62PJKnsnkSuR1lTU5tXaB0sa5FSZGzMTVGfATv
7y2j8RGAbGYDT6ahwFqoL3IWEfQKE14VdB0UhdVTWrpkYEPUDhv8K+ZquEmNBmCHg/cYJRcOJ0YW
+YyZa/gR/7ppujXwGnrZK90d8DjKUufZz+pF6qE5qb/noo4pqB8UU06/zeV4jTS5HN0RJq9mgsUU
qKDy7u2YqD/0rxqpCPI8QkCGF7PuMiHu0szNOKn0cEsRh24n3HkKcOdPYFQjbxJKAVWhwsd6/G3C
VBEhRHXyn2JHQ20+xnfssmhbXfMrIzegcig1uM8j2/r/9q0NA2NeUPqEngC3ge4Qg+YcJQGmmdhH
Ie98bgHzfgnyXwdyG/UJYINd8bouS/1kSdd3weolHryJvIKGC6ZWabrNX4A6dakA2OKbYJ7/4n5u
Gbq5IzP17BzHuZptZJVivH/DOgVmDMdUta31W1beU5lPIL8cQA/+Eer5MCg+Jm2Tlqk8FSUmbRQR
ZID295+Au5j11dFVQwAKFrVzs0OdcbejqfumN/V3/qqfp65L48EV8sp1gz/dqSnv9ZWrCk6Gz5zs
crTwbLQxJLVyPA8nMI+8zJWnQmVAeDb+xTAbw5AeTTtExjQSk16KWtHadqsyR7/SgKEbKEAZLHqF
petiKammL69UT1It0GjpcBaELBlKC9EJVo2586tky67txgza6y3TkrICBzJoN6M925K/8jjQ2xnN
Z7W4iD6QYBvtpzpbDj2W+0iaZxhkCvF9HPx53ESv3Hbj3nUt18Q3njm5g4FxxHosVxdiy/B3jgg1
SG+uT7p/Q5uI3c43oV5XdO8s2JAAwEpiTmJWoPY68vYD1itGa3qWaBXcsSMMyhsWVBukAoxwF23/
zNeCyUFPvCfnUDzcf+eGwQoRxRWBuLbJH989Y0/iU1hgVVSvhDiw9u8Ob4eAAGJjNG3xjvkLIklC
wg0jqZbdW60hMBrp4/DWI2/3RIwAGQuQuiuybxJOhAjPjB+JJZ9ISl1AZTfFrnmsuAKtPQ/KyKxh
ZpLGuk35EVNCFt1T/kJUOwYK9g0/5ssj1pJj0ctDHNxo+d9hgpMJdM/E98kdASnOEsntf3WLFD5w
yQHkVDa7hMmLnZZHHNqsMtS41TtF7nVJgu7SWsLvtKTA3asPpu+SGf8lHmqNt1AV5gq79G8xQpn8
eIpoA2PI1HJxATmKruAOQECNgEIBQhivRKQUB21NvMWiKy8HN/jWkzAPloGDk9cBFHgoikM/Q4kS
8N1YOvtHd8EZ0oHXeOeY7NBQzU4FzLrx48rfLHwaAsJoPUJcsAi7CPNEj1FwRd9Lg9S9hzL02NdP
KetNBil/ZGvstnSRqoRpbjyIwZ9cG2NxAL4v6LhwS9t1fN4UPkXquRGh6jlkz7qobrbHs9Z76mS1
94gOAg7xs3FDd/Fss8Pu589/VkEYFk/xT8gAe5XmrHrB+daF+WR9t0sA417GHFgscmrjT3JqPw85
7JzrJtYXb/4kDMsovT3xbMqgDeqjDK3Q8IH4NTFHFL1wTl6iRwQqgH/zXsfmZBp7Fhuv82YVA3/U
9oMuUTYIT5lqvWx2xGkW+gld1GmCkzFPgo2XjvZV5cb7aoAC9yWgI7s9ZtDmV3c5HdLJlz1ZmpQl
juklg+UsxzlW/jGJUkwyTws2yVzorKKPGRCkEXXL8VjCWBr5YckOO81X6wN4Tc8k8ANeA0Jh8L4g
QZQa19PeLcEsndivtdT/12QWeVEqQy1vK97vQha3chVk1/RAWq0KFZPFcrB4cRAT9NzwbuDeHC3Z
4XxvlPasX7fieoAt5CfqQqSVQeRTt/inxMBxqmYIzu3vhJ4eyRr8cND6J0EHe24ImpqlSCZc7WYc
i86OME/IVAhHGUfY2gnwOlheAW4yWS6/RWk9BtRKFLv/xi6DVOm6iMP5Cw1ylwLutjf3cTPLZ+6B
DuEqpjlNGk6cAd0X5vD3ox0nEzeQZPSHU3swr/ipVlI6/tJnfzPl+HjH5Cyox2sK020WA20fW9Af
O8wb3ODDc/8F4CbjRXyJ+qCvLVVLIDhSZwlc96XMuTA5SzTAGqCtSI8mSk1MdhVtsDlusRnLcAkN
e0sefPyv6x7dAWQ46+dDDFodzD6i66DMPc+1v/N9SXBbH1JUHROajrzOCBCR5amSoViNlY97wjnZ
wLnMSxEYwiTX8wk3XWmjIbcKLX+Ya5+qPS0Z2hCeur6xRIq/tZlkyL1OmdSImnvSaDJ/mxMXWCym
EAfQoCc3CZhSV66k00NeFIqLkRbwCWR/k1V3v7s1mVrWj5uTVeWG3DIc/R0dHkkSJ1oxrLEPQcqU
kMT5UyWNbLa70aAKNJoKFIiUXpTsH0ETh8RL9SmQX8a8EJcsWmsFLMfZTxrTlJCDcZZ/PMM38nxn
A9Gg8U8I6Ufoe8EH+mIVa12ZjLV47kR2+5wzalLQmK1lqg30NPAjjnZd1rrHjoEApPkN9Kjuxp6b
aHVqce7XS7ASMJ6UZHqQrp2agBUlvtme3QMXkqhhyA+R30mZZ2oWCnnV1iUl2YY1bTfcYy0KLOJm
iBDeDrQEEjGEFAss6DRc5i5q6sgAA6Z0XrqLCITkRTyJJqFMukZhZ+Wx24qzHk7aJWYphdDg96Bu
lVCGfNLRs4H30rTo8R+uay6wr+SHVfoAErTvLenqP7L9W+9PPmXC/hejQTu9gE3eCXSvJd4iL64Z
P3CcCBurzOP+Uu6VK1grNjxXD4KTBm7zFPhuyps4M+4grAWVjCqe8TtH6JejXdLrGRT17n7jhITn
jm1CgEA8YyNWwEF0DgOl0klDrcqZsqvw0h+E+ABva/iul2bo8Jac28SFVAvYmvLoD1aODx9EaVSi
Bmm49ptLiTFd8/yjf6ofxVk03VU/pRatPW/eJLq8eNPq9C0/wBINaMjW/5+YYLy+6cq9mWm1PFD5
c9Gr1BotYYRfQg+eFGSzMkjrx/fN7WwHiFIbdT1mpy1t9oFD2Yc/P2jorcRIqSrJbknljx3a77Ys
VsottpgKu6P5bhr0907sBAzd2jPYvIdvQGd6KInuvgD9PR9cds/Dm941w5IMagEV/oyuVanOG4ar
iPC8lDwG3dRnEOLupYi6pWLlhRx0hDUQhntrka4xWia/VcmXGTiThwzDg95JssngDln40V2OE+dB
68low1CBD/n+UwPT9zbrdjUbPzl1+GpfrLu5mbtuJOpoWNUkklwjcr8wbapR+33FFDfZ4qJfhf2t
B0D+ft08hAcOV8YuxHfa6mhswFlGlYEEoIq05l2/XqCBrY11F3x7D/DO+3fkMrw+pEj/SWFFjVzY
PAgLRkrUNEqlp/bK8ZNhqD+64e/W6ZPq8RZpt4mK05mCZujrG3e4LaC0qGlS1SuDxFl2Bz4uP9nN
pdFe4dvYeE4J509QIiedh03kHfgZdYb7bajnCC8BNMtzR89dIc0t4V3tp8x9lV0Hr0tMxV2Y82fS
qFaou+y03UYRc17N+mPylXOS3J7tF08KlDYe2qD0YemyPOUUd2ZdAoSh4LIelZxy8/wC40TJF1Sk
02YYFo7o7fWTKQxlabxjgEMFeb3GgqhK3aTEBNnT91Azh7Xjc+rM3AEZN+ivYR/n7EDFL6aT8gOF
uRifrDw1lXooxRwnbMvbkc6Br/sAFpp1c/io31mqtX8xuf2z9lypBXBNAIK9ua5nnMiuGg8mQwak
StfBhBsIDWd3AWEH/nHuBYrTwuzEXjXSyBiaq3m6vHgzLvtXQv/05dGEZ6P8j1K2737qitBoTCs4
k174VOO+V+erl36DzaogDVflBwSpV9N+oHcSVdPXkcQWTv+fy4Aty9HTV979MapLk4rwQodwWJw6
/TaRSLjWnUqJEEl9DLCxn09n/3bVqUOuXXnKCYEx0UttrIdar/kloSt0WnRAI7+UQtlZKKQZFDw8
b+srVN+1B4/snLphKJ+Z5moOR4LpLczQMEGTA7FpyJZMxzrqn0YM4JGtmvPqcUdIWp+fDojXe0GT
UPcf7t5H+IpISqhsQvDx70owQ4YkiMRNdCzwaEl4x6hU3kAQAIGXCNL55aDZ4seRD3Lejn7ygf5E
Rma5eSTpbUc6GHZMukgZNEEOjGEvN8TW8BZDMYtfDG+sR84JG5wCMiB63REoLfIhXWu83BBdJ4Zi
VFTaAy0onaAM6VXjctA7A2tWSG8IK6lyjhP8A65zt0YslJQNYm0mWigi4/t1ixA/pxL8LQMh1IWR
5GHftIsVnskHc+PqvdeGv7iaa/KTSDhnas++RdIQcET43qUoi8A8+istuz4FJzGVP3v/sODFqTR8
veg7jnRIupzRKqUwnj8GMFtpyzaMekHXxABN3u5HnWtAU/l7p5amHm8QRRwJN4bAATDNz6Dmvl+H
NL/mc30tpSz93M5oa+EJ7GLgf8AW6e7j/dOtoFrc5U8HERa8DR/xRhri0YwleahYB5Dnb7tlLyJy
XXrFVZblKKTmkKTDrVqTa2FMr0fXUEs7pFRQvgtSb1e7jn1uPGhSUFZa2/Z3Rlwe2XCMzHjtLj5x
bYQOyKebaBh3DI/bQkhpT7D0oewCO2GKYanlJWZ6yIfjUvSpAUw73J3QMWlmfi66h+iwEq7hZBy2
Bx9qE4RmPQY5AEP9JzD2hg8WkYKLi1sU0+1lOE3PYMC4y0VdabALY0aVBNRFkN9nBvISnb5M2Gav
6jvCsovFQX4JIwsmlOLZ5QyndcF8cfwBsarSW7eIS7La7B5bGSGz29pqLUBPUWJK3Y+ZcoI+Y1AA
0dF7Re2bpNVfP07DaE8UXRiumE9ouWQ61jgWyBxWwYZlYmaRQ5QNPWpQ7Zp2o/cSxdP1XQpso7vL
PmmD/q0cXnxgP0Eb2o47QN7fHVp5fsvq+uoUqdwsvj7mcrxWQGL2BLy+06g2WFyMtMPOzRFr/5zv
KShD6sDetj1PZXYa7vdbmhwfzG2ZkJ964M3gv17fbB8cdqUcpHgHc898O8pfhCrksecV8ZjYojfz
H4Y2fRSaoZhBir2cfU+LJxOPWNszqtU0tjLMXG2LUPYTi4YLSklolmHGIotqcRy0SWmgfag1+cHd
CiYoCwrN/6R2mzRtd3etvfgXJ6fS29d/vcX0kqLBFZjpID0nOTb+uRY6MoLFJEqaHgpdul4ea3NJ
2LHCthX0uudlqArOcceotuHDgEGBw5Mk/jYoFMsjhLezHaBx4KpkAXYrmldYLIz+YbY0DME8xhi6
C3wRIBDERmoPAsLdDMjH9JGwt2PCaJMX6a2QPWDHeWRjYGGPv2Ez1kDiJZoloHVgwphpZr47ocaR
H5cNI18kfiKn4MqRahzO15dq8A8K09yFUxxQhedOwpiya5HLLvu+VAnkR94xbERvfE2xYYgzmSvj
tOFiQnTNEUw8M6NNCkkRKm2rzkZiZ0je+dg8GsxlGJSJYa0JxGbyKl3OJ4w2XDjLVXzadWG0x0C2
DJtGjZB2e3RqoCNmN6KBl78g0rKApXMGqisTw3eQYqXu/zV0Tk7yuyHvrGb/j7D3wV5DFHQa/Ss/
bjGUIuTafm3PHeWk1uIMJ7qVV7H/MrVF1hXJ92cHaKLzmL4o5zAQxZ340YwIcu1wTh4Gu42ww5G4
5EmBhzdXCiiqr7pFS5je4M/MG9mAVg0PFP13tYLydPDulWEiiXUXQWXhHhMcRbuEFmnjEpHYP6xy
K5iT6kC1TBFCu+iQWeGMK8/OOhFM2obQ5J6sV01mdp2InIv6nTT7ziZFJFvYUh98XG9VEIypZzmV
tpje6uzA6W1W006dvx8uNYdJ+jIEeEzcEE9UXHaQn6K7+02vaMDaF+ASRPghY7O/0kjuvKM7x6/n
F9YebgWkkPEUpoWJVGtRVE6kT3xDrvTlAb2ZFp2aQ0y5O669/FELf8QPzvnFBiIe5+BKSbLc9qTL
5PyKIO7/ef6G4DFMycqLRvbSddmgIxuj+k5PocO90X71GZUIPYVGcJy4Gs3K367sj0CTVpnZq4FA
9eqxY5AL5uVIeSRAKtxCKmofeqBesFF6cceIsvNH9DDafj3Sv8CkL1yEjh+7BTbWNRxFTNzEWUqQ
8/RZC7KE6VgiChrSq1kaYtgS+dI6OIlPRIvyW1VZcdyVqxvdvsdq3zP1xjdr1giwOBRLW/VL16xZ
GrGN4KU4BnsDDe65l8/8zDIfAuwpdb71P1FLcK+ba2O81GCgK2BjUqmW4KnW5P+TC9mtD6f7Uw5h
Pe2F3wHZ7PAa8HAlet0iG0VTcSIfeabcneGVaoaQwWPnlLbIywfnsug5HXQXYvmYuZs9tQhMf/PZ
8q5eNgXkIyhI44q8shQJ5k6opwooGAKAaShRgjdBWsMwDiP/b5djoQKA43KGu0Z1MEUi8EonzAi1
TY8pHRS7E0/W/nLcryTNzb0jOrjK378i0eJIcAKmANwksglj2C7atdA8G90/NPOAHtRWOn5qKxBQ
K08LA3TvbNWdje58rXLgEyOeN8PR2rUUvrDCVNyAyeRyMPDd8+6k5FESiSifgOz4VlB5ZDSgOX80
jXTWEnonUZAV1z5JPbxFpiPAduA9OqdzXYEXIQD+ves3JONdtwboo+0FBNsvhrl6pLRDAZkLL/vl
MU0GCrouo60ZyV8BREPueKmUHC1CMf8pQe2+ncxDuAUQmOpBhIpApUaLQASqhSWR6/3TQksqGmmQ
CU/anhpaGUwO7kQeCBlK310BC892Xyy7IY0/JDLK011b5ijZYG41Wmy6eXcCHg0SQJs2SrqNj/g+
zY7Jjeh95X0CfssA+1j0EbJTY/ILhx8OdpqPLYLP6seJf1WcDidDkmzbezuhIjRtjZpkSpPHBjZG
tEXcHL/1BxUw8SpAdgqr8Ot66E2xNnkxvpoZ1dtmoMzCVJJ+kLBzSzn7UbgPFYnazqIuZxk1ZCOM
xcmvWw/39M46Pnj6UphZK7iXoIqqG4I/L5Rg+Q5+/3vKGnfAPUr5DJ/5md94psoizDm7G/LzaZvm
ek4qQLGLTY9zypk8kBiFXbE69AGEenZjQkeeOfyfJTMRF+KlsunugcrBzPwodxgbbeBs2ftOqjzD
OsY/Odud2oc3z9ZysoU030FnaSb5QTweUlb6V9AyyHoHCSz7DLRfcXB2cCxRgqrfwswsL3dx7/E8
6o5i0tlmabkabJTh9dX4TAJ2CGKbGiTU8Yypoy/7GIPIbD2zrgm3PfDbp1y3pzBN63UfAUI9Nlw6
K2y/QBxL1uXM6PqIY+9zkCvTFOdbeLK/2aWWKjTmIoG868Pe6k368igkVy3qMSpbgMyYir+qxRvU
MkR0CljTeX83vzkafP7H+tvDVUIv22n0e7RtdH85pkGb2pR24GrgFKdzPYBmafBUcdUbp7kuexX7
fEUmJVKtiHITKRbo1NTWPO1NL35Q0ZeXqLPMgCJWlzXLcAkuWMG7IyXqOediyHxepntZpmeXGsAT
9YKjWs5v8mTnkET02JW0/cPzsrCfHL/GmpkC9RyIH+9vpXTd/aqSl/xP7/IuRrOoa+LnEInald4e
sDzF46jxd13+fLEgbeJKRlTgnFJVKo8RayG4eif65Pse6Vb47WlblVVTZAVPu7ae5GU+jYS60z2j
dpICsnFZuIlH97ggO6uGR5cJkMJsfSRcxM61EfMcWJ0aH3LmILkD/dYVyInNdvnglb9bbWZ7PFrJ
W3su8R/YVUHwE3vqgO0XErJdbvq29YlbFgPLaEwtH7OTrCBpsg18lzMIsbg/NmrW3A6ko9++G+Tf
8oJO3eQms064CWoarc2Sx5hGERyhTYHM8stsXkuZim2G3bkn+GEB6aeUCsngUdCBKV4+BzMhh1hp
3xX0hQsQzmEep6gpO9SwBrXGTQq62V9fNw4xryGvaAoZuzfbhvqjiitW0AY2dUU5yi/LMiIYjay3
O6EQTd345fL++dXEolrULSd6IBiF5PtyaHIzJpMYI2M7pzxbRYZXT6OZcsqKEZ4TItyIQFPLZb9h
haJh5ygn2PvHsG/xAP0Y0miQ9N6bGNJHQptvgnZnLSbVlFLqHSFhUlQyxk6RQ0T6Xsczdb2dLDcK
vOrSNSuv716IBJiEldZn24JLd/a7ZdgoaQI5NLswiHQVkEqlTchZEB8pAoVfa3gmR3hesr0r5A0S
v58u5IYtWpjHux9XKdOKNk5sRwSOaKvnol/7gMbwz5N0J+IKOWp3ZrokgIDygZeoq7sO9AwKQuH+
O9Cc7flQKoeHscTJkOHvtStTtpcZ80wk5EdWu5qGZTPpmaZinZ/gJW97HZwgoOitE0pYyF07MM5f
c3wOwuj+wPM4PP3qFVSuuy8VxwPd8twNWe+xcxrq20LDn/F0PZ05gmmTqpfTYOfWZXeJBFDj7XCL
RzCGScAxkCe4LUWwRJzpPMwXEt3BE3M+998eSQKKXMaQkVwcpOj96zgg4/GbwSrIODowhfmKmJvO
GGXDUnFhJg55gVs02WMenHxCm9H68CNxnMhQIdx9MhtoQxWuAUReJixMsvCtyj8Jbh+aMO7C7P2B
9ulPI8jjSCaYIBMeNJMnSpk/pjCHefTILW0AGyCukl/4DDIQDWY0s34FMeRKOZnGnIALEmIU/nAw
1sjXooUi8V5cintweRUzMXRGBiNW0A5yG1mYoNCN2QqhLsk4H64Vfqys9h4i/Swprs7jpaEOSO5p
aHk+gfiqA/zTYxhU5PdbM00CcF2Up6z1/xAvTl7c2OWHS64nifrQ/3pnLPrO8ZqlpLzV3/y3Twzh
/lNcnYlx0Tl4b+Quc8KKYhuqmZqiLV1pXkkhxN3mt2lTqJP/m3JOhJYgAZ2QXtkmrUqb3blt7BXw
FRNPH9IqGcO3TnCbO4fKnev18qh/9ZyEWkxsbRtlbRijortmkQoBSBPrUYonIiSkAtsZULIejytx
sDf+aNgVhogCe5FyLYiSvYxRwb9uqP0DXSrCRl6KVxBiUe5mP3vfekqpjNU3frNoXCNUIO0Ti4Xc
D0SwrKHVER7oM40DOWgZnXZZ87MurPzVJF9dX7lSFTMwRQ38OTZkwA534IxEN1R5XAwr0ajVo8zi
AB6KnD71xB9NLEa3x2Qnj6mf1iOKCQTGlR/ATqYU2eFNYERJQP0Qjr2aYpa6nDFuolTST1keiljP
Fb4RrWDA/fWbGsBOfzzUml7yB0moTkEn6Bm/Ogl+k20hLjHC8NGYye853PpbJK+Y0Krva/Ww7QCC
nF84il9skOW0AKT8P22HCiseNBtP2d6MzzH4az6dZ+YzpmvqY4lQ0gcRx0EoOaJdFqFlL45MH2WS
hMKZoTHxQZFNW1YB9Ub8v6FoysFfpTlq0clY6lAsQ4XMY7F8MDMZy6qHOaLUf3zjAsc1eDteGvkK
bxxsDRflZ9yPCYvkYOhzOYixCVuVb6ryQEBJ16dablezpkEE4L9GyGWbaPPE06lrLH+LR5wyli4E
ieWbwv6z4EfmP/Rw/XACURSma5RMcWmRb9F0oRg+9APXHP5AmsObA2UGJQRx9O3AOtwgfTfDx5RK
MfqobX5nGy342mnnSQiQ+KvWRpppJhSVEk1Y+FhNuiD5L6mfsgosSRKKhdHC0jATuElbl1dN03t6
+z8Yeet8YnI0/rqBry49f3rQRPcdkd7yWY4bdbJlC54T1+TVmLvN7ZQUpwPyVXBpx89+iiMvQnLH
g79Kv/N6xWtLKEGjO4y2CwsGMtyok8vCgupcwnAyNygVtXL78X9FTkLa6nSzWC7v0TYN++UZLvlM
jdicV944F+lNT879camrtALM7JURVMqymAcqRoAIo8iLm+QiyPSMZbnd5PN+S1WOrMtoVNno2vR3
NHd8FMVkIPhn78c3hFoKDe/bGWtAPCLvFmtmlMNdPvdxnCIjxTRzH6D2d8REFY3zgfmNsDQV0829
Cuvh0mAHD8w+uJX6tA2wT9fwmHx0fBCBnry/uXakCBeFfCLLJ3X1uOFUgJIGJ2S4gqLONsbJ3oHl
LFrlh1r5oLlX8JE7QcBEUIoNPP2J3ICO8IAfNVq5XyNakzfVtaW1g4/NrANEg+FFixfaOpNR/vay
cC07T2eOqB5KynKjCxCrt/thqN4E4FSTGaoGKrw6BS4o/Ixn3MnDvc9F57n2J+wz8LVq9fOoI3JL
Wq3lNXNXnyWlQi/0HkrLq13+dbd5v/mCmx+RgbECwvwxJa40jTRItR19+o7bGMo+o9Pe6R1CBtrB
DDbF750QZpIscFBUN7qKvIpKkvow6Inpe3kVBWaBriKz4ZWTzMMkZFPp7elUc9u6NNxqG1MA2tU8
UmfoMqHG/bu2Ns3S2aRhg4PAC1nwAQn3aItHT6NGE1LWaiDOpIGWP01fTrZGk3Jp9VHKQSoGf+z5
J92xOz79PwY9/ejrovN53zbCTtuye/wQWd6Wv7s/cYXVFvPiTivqsQr/y4iInPzkNPXjvZdykktG
GTO9M5fjD1TrOi7cZ1f5Oxvl/uCBZVjMmdIrTaBdUlG5MWhLvoXQgFl75JGDxs/11uZFe3rzAGfE
ClDTskid38MnISLIgmnwK5wYNOZ9+NXNDEUnBZCUiD7xSgB3hN+RW8UzPlz8oCVjyxAvFcIXO/6v
MyWdZzasVF8Bo1lOyUVEo6vyu4ujLChMk1UDMF7dEDzq7VBnZTYwVAFC2QWsczKO5Y4vK8gb0fgX
8i6zP8QnBHWhSdYKBlDdn5wT+WDUhX4RyyRL0gDK+kjMZkMPpbiC/crWgN5PeIuvKATTWkmWgxF1
kVcH0L/0hnbkxEoGHFdWDZIf8sY6OumoJj2igl2YCTVCgPYQGQvgnJeKmAKCyp6GlH67sLe+yQE9
M+f/CJjA9zQOCrYk3q2BndoEqNamuVvGNr/T4B4X44yoLdo8/KMr1RsYXcotsZktYz3phs3lLFfv
V6WWpLIuM2PKE9cX6wQmrZ0FT2p0vnkmiMMDoq07Sl7tf8gF6W5GdfxKGIyV/y80Stw1Pu48Rmun
CXy/URrkGMEKNK8SKqFAqP7ELlnBx6TYyOehHwpzOCJXfv4xB46+fDvPQ064TXsLW2sOxjACQ7CL
+CrABzhvhv5jBbXnonGUQXL2YCjM29yyEFMh8HPVtGcj4hUVczQFbh4dqmUG4586T87/u3zTVvw1
MfL2jbAggkPJLL/VDbCNoiyjaDiizVMPp4JmGIF9KTwdNebPSh36OLQSvAw/u7IzKZpb/nFDopkM
yuIp3UpDG6ArSksv87gTQKQz4VYQpBktn+gFW/508Avyamy4O17PEmVPNc8JHg7uHuRDpBXS+NGz
IgrXYGqgIgGxLX2TN+dwGj7J7vpayUvui8TUblQhchft+aGMZbJ7MBUIWBCRMtrNeF5QlxV4c8Pg
svXFnhLjeRNR06y6/lyg/ZkxWJIMVD62k70RQYo32feAYs/z6y7PXjzF0oEVfT68hRSg/MUq0ugV
TYVSIX4w2PHI8SPlBC4MyNejC1h1P6J1jxnfvFmuZ61iwTGVFZheqL3AXPgGHPdZDPlz4pnltGCS
I/GgI84CJ0Fj+mFTRL54cD+5dzP1MrM5nGieFyz6gfPKi6Zwa1t427o7HIi8V4Kt+sLzOtc/xPOi
UIzYGNhPOXZgQfkDMhcoLQ7ew9OJ0vdq5V/7up0O41q/xd2xu8GbTt2ZXBVDrWY20oPX5l3nR8z3
sZM3/nnDjwlOw0RtqV9KaxXy4/p0udxPnMCf1wrZYdobCRcgz+2vRrFjD1iz6SB8w0FvyGC+v8yK
im9fPyvh1a20usuwT+Q9qnRtFOdHbElZdvGGZZbD6XxOmIYmV7mgN28Too1INCx3bTA6Ho7hR2Lb
qpoMV3vD/+e4u4n9vvsLJ2VBLiP/8ia9W8sGo1190anZuTd8zgvHi4WPhFvwRoLv0XnhFxYpvK+I
+HCv5P1qecJRyOxK+GLfzCedbGh78caHN3UY6Jhw7xna1QSVZVhIS4db51DSVBJL+iakqieOcyRw
ujTNhozG+89OZDzJN/QxdnYwJPPRZynElMDbGGU6e/uE0VVOL0mq8gFyel8ufUZZHyEq6ctexQE+
g/xzhSg/dMu7cfF7N0sRJF5bpFkXzPVe8kDIee6vKWxn9Vj+v67gK+X54NWlnnFAZWi+MnOznodW
kecVHy1KS/BUUHY+CZuguDPLUjs5WaeJuWqpnta/RoICrRHay34duAACTzEMB+gNDeYKtBkPEKP/
kT1DR3kQmTJWUgDsk12kSjNVKUVsh4+oWAD1bPkSC3D+PMJU1K+g8aISiXyvMaW9BGG/l8WsMyQ3
445tNRI3q5wOvnQxcufF1/Hx5x5b9yoG3RGoIyd5oVug2JVxn8uJgY3P7kJG22vJzeG9562cwJmG
eQxf1Y7Ytv84V12VW/E60pFRs/255t4qfN8VYJj3cKtI4HrKBc8VVRlkHK7UjyroQ/jLfQQxhzjY
40nKiOVszGzLF3UMQ/9KNmjDiXoviJrdw0HtuJH9Yjp6WwQsfeBlafG9Si/sq8yIndPHcFqGwz9E
di5xgnAKTM0NZKqPrbWo45M38/Cjrkd84Ou5jDXx11dYv2mcXwsZSdhN9EeG7l3RTBKRwwhG8Cil
LqxMMJmyqNo4jheNOa02FYuJ1JpjYPyPbWn3oi1+y7Zc4Uqj0HfKosxiCECZTLD/pPrpIJ3zqQr5
mhC/HfZknEUQnuPItYTecpN0k/0oZ1EZWH1Gje7Yj85pzs4TjvIxbotJdcdwhrvt1DiOte5oAwWd
X1rpbTBisFs/aQBH1mITDewLyB1M9/W06Othuu/dEoJ5rQuxWI+urI3ezZkdua8ObX7kXcJ9wfqU
tU2yMupKnY8+E5Hn+m1iACYr+bsmlgVHhPiYQ6xTW07FmM9rofxhCQspX98X9xNTYvFRt9FvjmVM
+2iW2jXWGmO/rxvID4BJCqmjJr8TdcMYfT2LKcRGwRg+H9OkIrXC8JmITGSHDzTN8gTrb9GJi9Jw
lAizAf/Bdiu6VfGE80LA1pKhqoSTKrOrywv2908CMAMnqxlekYJTTHneiV0wgEiucpEpGXXZDYfG
DOabT3Bo5Yq+wDjgMZH7jfQIjHO8sctNXDGeuIDbjvXesAWuIE5vjHFqyv083lNfG7vTWwNbUonW
eVvb2eqd8sa7oI7aXfO6wMkx6IZKQHu0MqpiqG8l2L4saVbKvbiZIMnbvJvIWcwQ15+sMQKzyYqh
VsOwvs4plDceLHrVzFbrpXQM1XvO8W/s61AZmybhGXEh3bxrzEytANZTtsK5JSRao2w7/hrZ6K2L
hNfnFdVDEWk6cy0hSCUbNpOj57QFauPNzO98GAfLP3/CZ0PhDreQm1/AdYwocWW657+LantwP+rb
Qz4Un0blvcm+K46ezQMmk2CgpmR8q7w3r974vX/Q2Xi1Ruq4Rsa7xMQ06Q1o32li18CXy5JQIHph
puboLY58XmwKV8BkicpAOTJ56yWHQVsdcpd/DoeZwv1yrsVZYGUEL3knjdvjR7DkgUEK5ISSRibt
ZUEn/TIa5SWBYmsf1AkBPLmHG48SYrnYfb/3hEL0rYFBgWowAUvgdO8Ek7N3xt6bnttBZfHd4Gc/
a1y8e3ecYT1dMFI+IkAS2o7L1sMsrb+UwS/Z8QhgN7Wc8N57qiqirZAyK1nKsaM7k3k+UGTHvfl0
4z5ZPnhJcHdtLG7kyg4hzBClXxpU2XFhQESV52/4m22febD2aV3EnD/gx+dvpm9nhL/EwQ5D35Bf
5mGhhkQ+MUhkrYfPHwZU3Oi75RG2lxyxqnPQ81ULsDjTR9SKcTU2NSxL8Es5pzn4LkYWOc/1tuod
mt3zBUqK/XB08kyWER6JV1G/Rg4Bg9YBkYVU32EIZx7Ma4jX5uKaeDDfKTB48O9KcVXnLRQa+jFf
oopuyV9Uo+Duh15mrOeS8zhPmlxw8go/3ninAny3+JpmxLE3EHbeMtg/ZvxcEYxq01Lxobg7lKPJ
HrM6+79lheKU+t7bj0ZSnj5HBTDwbplbugU8hb+iLcXr1HiVnwn/5+r6uFJ72gpFTGfiMeyeQU6z
y48v7kfthM2P8jU0zW0g75P5PebImhSaTn4lGMaZRbz/of/BSMDnhQFjC927rlpZ84elEw4pgakI
MgB3yd3FmUldXAywsg3bzNAS1xMOKr5YZrqlkotCy18l/KU/nFIamdlg/CF7E9vzX9aL4GEaD++k
FKbqwclow1VUbFfNs5ycyqskw6g1Eqgw+lBlHSH0ZLgpNHWe20+O4/dMhwluLeaGm3vQlOsmPAus
mz6QOfxji05dAWQt9/uCedG/ESM5dGWnL2Vgx2h7Gv63lZiWrUeJmKv8frA/kM+6AzfZdxbVNDpT
LdOYAnNZOqywn4V8LwprxC/Zq8u9/Nwh4jfAkj3FWbu5ag73xkHS7odzEM+db8vRFpMPQeSDkl7x
0QvODGxehvW7I1QL4CZ2yfjp2hCeKPDZ+JePBddU+p7+DQyzJeDsBNiB0J16ZXefwzFO89iVooes
oVdrTgijJpMr5RFROXbEzlHRUebWh0MzndBtrxOGyAUNLJXtryAHQioQ5S4OA7Uv1MJeT3XQKbeC
aewwmHMCu0v4cG7lFtXaSbH9fwi5VUBMlh3TLWHX/BhLDyh0DANWSvtkOIqCEFzBy2iS51Al52ZY
2t6txve++5GmudejCnjxU95h3xn7m6cxeBlG2vvMghlNXRuScP97rhDbfgGep0kT0eJjO7WR52/H
1vhFchl+/irKlTo8DYUqj4SlNS4t3LtLljtOC8PkWlnam33tWIw5xC3wO1fwJ/wzpbrAy+Gvt/bc
QX1WUl77n4JEPCVOOV1P0WDkscHURxKVMiGnZcoXJb55C7dL2Bh/C5NJvaudiaxQKkKLgTnlH8c7
A0/1gDtJzSt9JLS0b3WzDbB8nkTCbjAwDxYlyirTJUpQLRGTsZ5jy08WJs9ZM1YXfKKJnClknsvs
Sa2Seai5Fiw1QDQs0+v+J493yw2FBrOCno+/g7AoaqsYXqNoiGekY0rDzI6nTWDCumB9Rgz3lGQa
T1EBg6Am5FzcvbGh01/qVe47tlcZQgQgL2rvMbpCFwyvLUW0JM9Dz8q/8kEQAWJ8EZ07UEMiKtnP
BiNj2JqDbiStbAStcVGhharDi4fDcoiCvThfGCRAhW3X8guTkeS3irOy/aetrgzXyl061rLhwvkV
hrUz3nllBSft2X315o/e/Y1lhojQjaGvclHlfHoXczFl3dCJZzkmGPbgHhfynxTv+iXEXy8CQMu8
UnbvccEIe4Q+R5I8HfbdS0XojzHAQCy0AF1PNRYADf3+3d8r7hb808MjFWFjsolVXLYCPmytCDv2
7NMhkcWuKZbIjG9zHIXHpBQEq5QfufWGbuWhja1Xjp6FJlRLncnrl6Oe0Sk7cBHt5jzV1g8AmfdY
KNzqhVzkJFYWGJy6VRXeqlRFYIQZ4SEBR3jQwfa/a4PbZ+hz/qKbAbeI/Igb1WQ0IrHUUieAYJ0y
7ixX43WtHpjGSj+Ct07/iGOPbjq65sCj6XEELlnxjG/1ccCEc7ZE+qPsv5R2dlMR2ITt00KUOrJ6
3FM1Xp5H5x+zDh4hLTBbQGFsdww0PyGn4sFdAkylqvTeCwmreLM9AWADoCVkhbmvU5ieOwUOqnD2
UyYweZImS0k15Na350Y9heKhzXSEJoDZ9TkxFYFIqNWXF7hJRUwQ8KzDB0f5qMG+rqla2O7lVL8i
MuLxqqyB04vYyUwwAPzSz9s5Y3WxxCKj32qeUwAP4bAUxmHhoygFqmYi0bMW8CduBp/33bXVQTZW
Rh0JjyV+Zqjz7ig/eJk5QGhaf+Gloa9TD4vFMH64hsVJILqhZPpn0iH0mdjKZHY17Rs4XO705W/i
Bpa5OFVylQhLelCGIvlB7FFSeWG+gLh/Cvs3a47R8wVK1imBs6QaUBKP2DWQMLBJrLg/jUY5hCIy
6ZaB1PQ8Mzf/SSR7DyFhu1PWCca6MIJcsce7v7+NmTY+EnsCFI87FDOScV5rSzPhKb/ZoDCU52hG
FUg/CBjiLkizs5uC2+/p87lA92XWHS/mqDo9Of9BW1/EVYuWDbLyVS84f3gN/ZUVmeDWfJXt8WIr
N6Ev+0kxt7xFGqiO9/NMmXBt9hQ+yJ10e+nNYVLrwE6uWm4rXPclt50IHy8N7Fg0FhaCmF/rC8Co
LV0TVNrIAl3Lp8hOFKMV7sDiOzuFRk6CaCwqAMiItSoAlC81s8WVetkdExygN2POZGZeCR9XLxQ1
793SbQHoxBwHF6XhBp6EuJJVPxI88zOsSvtblMrJA+aEb5LL/mr4z6CxGzqoExFu0HC5R6Y7VPNv
eM/Gggg6MuSP+Ix+LlUd0O9txXRy2necW+TWWvxP6dI7ZBf4JJC7Z92kFBvxfGcG8xLFw2DSPXID
uGWtSX5ULRhXMREKHiZ+hDGr7NbqISYAJ80Esrijzx/OKA/vAWWbJWBWn5i7SodiFYJE2iXNiGRC
7jfS3BZ3bpt7u3fdKv+01KVOgUBjmD9zjqxHFcU7AwWqZdEE7j9OtNgb2OnH2+6Pcdyo1BGn/mRu
oyvdAl9osEKW2IuE91PByolzx27+W1yGeGu4FQH3HymKnRadhaHP8sUPpx12NVrAwO472K4yQob6
reUfhP+eJF0oOWGFAHcHXJMrCA29WBIm8qjr0UUxrqafzg9OKTLt5sEaWooOiCUX5XBBPUuyyEIp
s2TYROp9f6BknoPr23tZoxpu2V2dP8mqhli92GXTMdUq/2MgHua54D9nSER9PxvZDirtNDj2c78+
rN8IjayTfnpxdWRNErJUbav5EjIC8vAfvZeCdVc80TxHrnLOq2d0zzWwgprvKz8oKJHhancNrbOf
nStBK2ipgOE7jWeTY3LUXyS5HfsOiY8g0ArPIqJ9FoZqqilJSlLuBzRvff30TO+TI0vMIWfrMSNU
YgeS8F+42A1ZAq6UW6DOxR+QYDlztnbz2VvqWK61m9uZ9w7qfXSvGVveivGqEahPAH2dY9aDYLhy
b+ow/HfxK58ffxNdv4TM33QbRjcwBBN0BITwrwO3nukcNBNhW8Oi7952oPaTCuQBvLgZ72JnsMfz
uHOrbvsDdhIgIa+MgjmQeTmHGLePTEWhxDJQFpIGCWT6k7164b/uDgDBysXln74cJJ7DFOg8qgiU
I+c/JO6M/1KCIyvtniNEJ5+uMaGOLOYbOO5jFKZYD74EkkinsCPhfHitVW19EACKkt4VPPGETlZL
/cGKTYYGK0AR3NCpVoHz+PQIl8CjqQdytjxhI13iq+4VxJEzif0YTeu1ee3FunJgrXG97hvFyCy7
OasSDTAbQbHFVUU2By+WC8nFmcB/dvoKRo0UlSfHMM/SCJPpQxBHL3bJb90AkhUmwHq9Jg5lPTq7
hSmy4uXDImbdit8LkUW9C6tpL5S3Xm+kXBSRcSz0wSfJ+rfpCNbSMZkTKBaE5q1tbChVHMzvE7wQ
4SEjRNmSVaNsg+1cnURLp2u3c/MvsSyB6zd7hCpb7HVcdt2YmJ2CBg2MROFXQb9EH6Mima7kgiY0
9ZxELibE5+8G9idM4LFz6TQyRxooZdiCxIM9WcFgROz6JI0MVNxismwwgo25hk02QkEsRwRN+Pjr
INUD3n971S7aMWRjQRM++ZMa8HlRoHcd9Bm8l8GJin51KNfDJrVGXcVjO8lmPaiwhrRjhhZnHhpg
/WeUKz46CoQNYXJe0kDhHAFeo6/5g15OrgYvBu2sa2ricjLUCvqoRIxUHVPx0lnirhYfl97ojAzF
fZA8sCv9Mnx2ufJY7+oCfLzAiCXGya2sSehHopAcEV9Flmcvye4anWdp98qm9Uyz6j8DlkvXDfO+
vSI53IjzAPa2Va7KUdmkDVocIllk8QpY8m1ktifSLybjMElpb21tTxaoELmzWbLG6RtkEjDqjI+3
f52msNKKX+gHjyIhv/yZ2a6gCnTJSs+/C3D6FrSFxoPVAvtgn5oaF2Mh24krkTBknNuwlEDxOHyQ
hK5DHNDJr4gQ1rNXMh0IWv8KYedFssGDXiM9VFSh7JB37743cDa8X5Dg4yDrbNqoNVEMjBURg+3T
TRADCoAIY6G+oi7P03GzwNms6lSNanktvr20xE495wgDPNDyLRi0JRWIskdSf2R7EsKFExwsnCXF
WWExGDxrj8rFRaHwAKJfY76Dnf+xFEvi3wRuNBIp1wdnU9YDNnK4zRw/lhSb46/S05+GXLBbzfRY
QNX0KCKmnL8+BXkmM+3pgif+9jBzPBZ81OCgCFfCemuBSdXIfpvBgD+xYpTBp/TXeUUf/fHg7Bre
s9z9PGok3vlq0DECbl+y6cgZkHIoLXHh4z6ZHQhZ60RzsO0SSQk+QEoAi4SPn5a3hvhjAG/EuARy
sA91cKc1kKjaWitXXy9ScetC2KRVFpwndzAzkwK0wPAoOu8cxVCJdEdUOXLh3SX6HSUn6FWLRH1h
NNEl8CIVd/MsUX0ua/NAmaO/S891rMZ1pWgzUL4HRRhx2wG605Evvw4phUM3Mni1a2krPt4+/ycn
sXPBXGOw6Jb64P4s53bHPoK+2Dof4a5f3UiRFzUzXKy6QeI4WTENnX+wgxdafw5zs03eBoluB51g
EvFuxVqaBX/yisRLFpjaLNkg+Xg4rotyOQ6DDZcjN2ZDIoNxbIiATmqAzda6W+uWdHoiXQwibZC1
n9me4tGr2oYV+Tf/CrFL4tJr76a4yEy5OWD00BwAuCj6L4ESgVLwU2J9lAY+XZdZsS6t++xr/7a+
irqboLix7CPUPUBp6t++hlxtsHB54J8TgBUfiwr3DSf0CddOg/Zy7gZsezzG3ryHVenH2hIvYb1E
PfFIoD+Dj/pOhKX5gJTc2TCvhEXPsPu1PL+QFfirViR/pBtYxfmoAe5PiZJOl2+kH7EWeHljYtLN
kIKL1N1jERXUcfDXR2kloHexASH7XhyoS6qJQImH44laBYEGVWfavWFe5jdaRo5DA5+fJHNRY+rN
JjN1SbBLkcVVOQY0p091oPVBSjYy0pHeyf7/lP9pDmJOYT0uLpMAqDAW4R3y7z1kMpgppbU2Omi6
sPKc+jFJENAY9NNb1noCfTRbn0wG40dYdHWibCD0HmMAdKY5TLxogPIB+dNaP3nyq2+RGUvMV/nD
0M0ggjjp4vAECo7XL2rZsTJrGFbapwZOmaNJCnUVevirhFhC1tE7qgqpb3ONZvdImpRDuQ1Tlpvz
88EDoMKHMWxxYZ3XY7Ssj5gLw2dEcCMJA3plSARd2vzjehBbppcIVC5NITN6m92mzFMjD6eU2uxS
vRq8ThvKhCyBMz+y/6Kvi8oXbZi1OH/murK/bzYfRkZsw6AMksj0wRwp9fyo1RMzJ4JFRYvDNcqm
IeXRUxF+mOyVFMi0glk0ahOlySSwkrv/XA2yPn+h169Q2ixy3GOoTpCtOemAlBD9E/sj7/fCRGK1
GbNHu6C1+28w8GJECXXDj/opldt2l1PlPLy143l+mqNCC6JUOZiAQkpBZsRLV6daMPZzc6Io4Zy2
GubCOM8Hh9DlAOQNlsrNkH6N+gn5NH8xHuskkb/jJ5lAOSZp/UjQAAEooNSsX6ucbuBqP5IIVR9T
OWIjOMMIeZ68YJpLQCNcgebwK9yUye+N9uSTZa/muTtq/IJeeh99V9r4jVnt/ErC7Mq1/LUf8NmY
JXfNnE5LB0wzvxwM2lI/HBcMsuPib0VtgAH801n2g2Zf7F5l42luMl6AEgtvYV5UGC8XxPHr8MFN
nOYLVcgIWv+8qDjJcioD6WLAAS4DKFVzt2GXF9uYL698h3v7NK/h5VhGMIuliIgx7YNpSekhiwid
l6UNL6LgnfslA+87NZMJ1J9uF6kys4G2ITQa/7AQQpNBsrSKYuMSP4vHSRZYxPgO7Qi7c2TyFZvm
pv25GVmM1mbQtYHVen1N1hAaiToxo2GABSdTUcdvLnT4akLucbSlt73FA0gwxQVF3XuetKzFl18c
RSQzm957zdVtevfWMo3YXYtkg7QW9P54Z2mmD6ucK7Ca+mrRuYlX9c0aFilpce6rm3M6wW3g06Gk
mLNRDfRCD2LlZQYf4ISEoGoS+XXDdekzzaHefxjAXnTZ+dbNY3HdrkbWMjWEScPkfdT76aU/Dezm
t016FfTubgcp73tMKjvdjCc8LpiwQ9TViNBH6izZa37EERu42TiTPw42tdCd3J8S++DJ+pWwX6Gi
wc3aehwRWxGcc4aOHu0g4n+buWELjLJmDU1nDL/meUfQYo3t3B2pZEjVrasgpi78buL9WKYV4wzZ
0DC47Ck50ZSQyrzIuxZPHlz6mZ3wPiR2xsP/woTXh++j2uA6vRvjR5Tqyjy7DgFKZDL2siahrNp/
seje+37o7bUAHy54RJSFiKJlcQ49+ucQFWqUuzNjb+RLsd3ars0YEVXkogZl2/yhzYIDt2etzMdd
CwR09iPDotyAsCX5l4lGZl1YJkONQ8gGJnEfqTWd9lK5TVPzSxusR7y58FuYupLOrlPPz5G0HOPM
Yv1uGs+2f8cVp2O0oimRerNnQG8TJleKZzkQikKRm6fEShV9LNBEisoN3eLdKDaUhWpXb6PQWOyh
GPq5Jbt5/bh9ynd+h0tk8tdscIfiDo0KpWm5DC9ErH7U5y67C3ulxo8zxJP8LO0nmlOHGZce+V4W
Zfy47qq7NwZOe0CcbCJvLh/qlYjCLv+bYXKbaw0jLs0/oquoas8fbm8hGZwfXqQ2hX37kvjdMYyy
RmKXYVqy/yteMRcMD113fsHHm8G7M5mRSnl6zLW0/f2D6moqUwb134TxbLP/t9M73vdDow/82OW1
dMfKnEGsh2clxDqmsKxYGiZ96USEjXav6NLI/wlSMggTPIDhOElt4huwwUFV1SxlhYO+rATf86Bo
2OY5S8XSEUW8+6z/YBYvImeLSGZiNYjN62azmi2dZBqyLG0U7jTtSdJD+LoKhU8J0X2jCKGYfyt0
RkeCTMfZgkXS704CEbdlIXJdMlz9D400ySkc5zpISGGzuU9v6SXGj5beSHbmrFG6z1MTxU0QB3bV
q0dQG23EWb8/dAerE+D0N5BpASXp6s2vqyYSdC5gtIvACozTAAsi95JPxwo/vM4igWC48ybPd/8R
zM8gx5szFPDXCNx25Q5Skpseb/T1iRImh7z/QQtNl6cvs8N3nx8JlC8+9C5G7224i+XA78IqsrWo
OqPluG+HnuUCLq6CfqeO1aJ3jbnBjDu07eu9KUHMUh303Wl+tzDlXm5bRoG8Ki7T1ZDMs2dOW/C7
rtt00cQk+fCK/KuUSkUy9tbrmzp1lrihWDIUaPCtbqhQpWhvF54TrsAhzxHVUfI8C3MH43+U7Lia
8Qtlv4Bot8g/LRLM1niSUDDfkn0LihnMOzTZVFhIQqDZ+92Ro88cUprpvkFLUJJy9pYIybBo9AWL
k9SzeyDMr5uTwKAIBkPnP+C/llu+gcQCXHgse0Rc1Aqjb0GYlVmaFoy3Il/TJ+OtgIwJ9UpMfE2B
PgRpDijruEEmyjaNWWRQZ1PBjvKh4tcJfCjdRTYAQa0ozPoR9Ho/d/EcvhnqyswEI1mFETM83pit
bNIB14nORMYXNVIOGtJCABbg201BMrDyuv3+2gJv1qTlg/abJEH15biLYnRJOk3CpBidt59PwTK1
u2yobKSOilvu0QepEPaQvBYQm665OwgihXcAchGcdEqklVFEQ7pi6XPqQ7FMCzHa2dQQxPOA+6v8
eF/uu1dzywjnPoZXnnBbCBa713yGM6OYMHEdrEdWTZyMmjYUc0dSMv1640lc2Yg6lINul2AMu0YX
ZPqHsJ80zgcDMFn7vyiKnff/yMYh9DN5emm105BYbyyysIB2Zyb4fPmfP3MM3QHvoBNgj3ZtwMaF
eNaoYUUGE25M+wk7i3JKCI8pSYg30K89LsvQD6hYYV+7bDyeSHiSPhGrvbIATIj2pUX04K8CPMKK
jIy2ArqnWrfYnEnDcuuuCK7qVt4ssto2WbR1JytHtjdPffZcvq8C5EJgkaWtBi4GJxm0Dpw2Z1p6
F4M+8qhSZr6FAhLHCO3zdFKTa5jd5mLz1ZLHOQwaPQyOcdJXrIJjz7tbu+4VFbCQxZmVn3iA+a7b
6lPhf/qSD9Kc+bGcJ/1eiEltRr+9BaR9UddtdatL6oBOk7FDqWiPufvA3dfZkS15A99BlPLd6OcQ
nhtd5LT/pEYKx6n5k8o2hijOX/ent6AKqa8tXUE0zshHHzF72YQepdvrxjO5aCv0aYv9RmwTX/vC
Bbvef/qUwyerqRTnpP0ZIencXzksjCsbTIQItswA9vUug/qAXqntK00wKJ+8GDzlWHOfLBUqib+8
UF0NLN5E7fRIMubH/1Rnkp2qXOamQ5c6KD+ydHOTL1FXVl7DUcOCs4vZZ0BOwWB265wYh19LFpiO
daMAYFfkRt/yLha2+mpxu1VousVNKTBiEMIOskvr7PksDYJdC1T0OTzvoaURZQLTqVe2XrhOsy2D
32kQ50R5o3VGqkpc8t7cXAnxm0J9/CcKbveFEszcxScgcpYI8902PEOudgpP4JZscT4urRWUXYQV
MPyil8Dh+fxUHunknk3zn+7VEmSrilzcQ/PTMoMQ6E5Lfm5QrtGI7iMVPzWAXULgmnihLHk44sQS
iXH44ip8UfeBtGGSz5It5dcNePEzRxjy4A/4weojMc2Ww7xW/c1hlcA2URsKLZVPvtu4dmefyP0U
RzDD7fhccdpDtan6xUbeh6rXjT90KL65FJbT+Q8vnJSf5e3znPxqpcqiNLspGverWCvZshBBobZZ
9dOeBpyp8ZwoOR8jDvwmAMl2JBijyEYpNrI2LWE/bI6yRwwcVznvZYeE4srbS0rSwgKia2jiR1Qt
AI6W4Bc0oqnAnKVn6Qzm3EkUw0AISyB3iRJBpGS1208IGwOVte4k7sWDMwiJZyE+oHTRburtAXf7
0FOcefE4F6Gx8t3gCY4fwa4ekT4Sp3MZ2aots5Grp0sPwJzzCFMNozIhwRVLSlDhlU7JdH943Npm
85Gg7i03b8IJvEbqPdIjJe5VgzLRVXIF5GZNce4WrWkY84DdssoGSlt1aAUsAZVf+ApVpQ+tqaS/
CL/rQDTrrqL5PSSJtp+Px8QXVUsWFlbIA1nDIMMcKOKo+ZRVl/5KEuDw1VJURrjOEe+jLzg926+F
iB4r+j/akvmjYNKopU9beJAodnYJc8tXQMlC47B8v6Ak1/QI9tNt8bWDde8ufBkojSGLP0W/px6p
uB1O3mOZyZDD7sYWybaxeVoU5dt9vJ5oMpN90p7PV6LzQ5RDfexwjOEILViPTzco510anFwLa5Fp
yEmpPpYVFb4XaG/drfkBZVGlfK8hagpVyIffxf+6TRqGt6wKoVzn7cc2QGxUpNqIqX0ErA2lanek
zuf0fRBOzA5JYQq+mFjJXRAmLJzNZxhprBxysjVs9Fl5dVXEaR9/7BCXhRZhal+A1wS/boK+nVPZ
oeTB0FwexhqtFn1FTM/tu4QenUZc6cG1gtdv0UdJT7sOc87NDu5FR2VzjzNFW8c5PQyFZTTEupQN
w01isBrJ/+3wfT/cmUWRPwSugoWnT86OBHhenk9XlJJoERePAQJXGLKTVu3EEMFK0bgG/139/fDw
dLd9XCPRsDBLcyPiYuR4MeU0DnfNrSWjXztJ+JuP/Q1wGm+ozx6bJcUIPKgtzZRfektv3M5ukuWZ
1mYXfVqK/5zISFaFf/D4i2TJ/Y9nkqcSX0a9iPhRbb6SeLCMWCywFLMEAUV/Xo1sAcjAL1bYzfby
QmTGr9+xTPrf9RG2dcVr9XJZGcebG13J6ltWaOTH0BZXpf6l3jSSDOgGIU+I8Al1gFl6HnArkxfE
Fl24LAAfFocrMmiDx3Ztl02kQDA+AA0jP7WuhmcSJft2wyXT5njIlBsT7a70SvD2trXse6rSwWlr
mzp4WzRYl4aQgNyVk50TNDYFyuKleBkUN1ob5E403SC49yblBgzNte8D0ov33kqrmTpAfhRX5E7X
Zrx5bNzuXvnOeUdu0Ur67LGm5NZwgRfzW2r9Is38wAVs/ap7Zyw+IW7/y1Pi98gIcbFJf+etNyMe
Y+0EF4SmX7ciYTbbTrYvRl+wtCIrihMVcwTJljYwTQ7m251362HtbvueM3DEIpNYrrD4NRg6Q4+0
hCxeryOgElpeX+i7+cPHrUjZ4wTWedL/SMlmLTkEE1NOhb+Z2VKTHc65uWKREf7EM2aoODR+WqRQ
su3X0Elz7FatGq+Pw6up8DHSMHIyUIw3DQWZeSfptm6scFgZyXU4m/pIxrEO9p6l89jw8vLQNO/K
mtdyUeji2W7mozlBM5lfjRd0i6+4xMdDKOXsE5ffQLZ4b07nvYgGLJfrBXMmONzcLrzMuaP1H8Mq
CCatgEu+kEp1+YXqF9Ke5RPnGbJLspLW7gmWhOBOGHAee/7aw3dVhp3lgTRL5te5VqppoIso1mCm
lgyDXgW+U7hV8xy4GV7HSy+mRhjDp9G4ePtJyljS12l3TAZTm2n/995figNk3PAMazFTVtY/x43m
6MalqjgnQhabZLuIQD4fGdd3ATM21VDbcXf5WbTp0G9EobbNc9TRK/za1zgHmcM7kBaygdgpHVaD
Ilpms4Phflx88tgSv2z47SsoWXMKGgru1k94F+zMdaxiUDx66/lUeQH5NrbpH4ecMjPwxXcWFjh5
UbratunVrLNRKPKvrh3JwN2wBioQQHv/h3GEU0QMaAhaNJAmOKOAxxhzxbTZmk/qhNtLI9QKuucB
jStgPpY55N7byPA3RPRr0BNPoL2l38ZV5poJM13JWJmTk97xNtjt92XWg7HkK8h4QqIVAhMX1tDg
Q5O6vJpekfkzyBo1NrI2sECPNGAASw9cGecgBmfuEuqF0WGsQb/R0H/NvI+i4etDJET8ehrwg8ov
nki/NFq72G47GGnPxGv0czHlLxqaIFPprUkDnDOGfBBwYccI0Rr13atgSmUCUyNKkwdGwVM9ONFp
i2lAvX3idJiK58Ru5+5BpoomVkaqDpp0hqKh9BCbHLva60QCvtcvIm1LiNmYviFm56/TPgFVl/GH
Ij8IFK6g/fl8lZsMqP/4BVc3L88OUAAE8ndR94qsr3JSuPgLN+AGHg1JsnA7YMY91kLSNGyX6to/
nxdYmJfFpHWDaR6eLkg+QObZXxPIFEj2hKEX2s1C+RCD+hhqjGv2p5fntQioMC8ZYzqG5RF2g/Ix
uGskyyj/qJo/HjxmteYJUqXvIu4eBgA8x6eVcKORo512kjZsDtkX/QDoWZoYApBKgmezJHo4wbZU
Dk6CwSljC+kyPOykzsmZU78dds2IV+yxMrbzb0hd4g9UKLHT1HsoD9kWyar5ixpL7mxhoTNux2Jn
MJjVLvXRYJRSmrV6sNqehITRhBLg+NdLaIJa0tSQdf732GWjkYPWT1nP35Yat7kwIXkEMuU2KFc6
OW/BajLA2PqpLOCAKCw6dt9zDw9RJxQLnW5zUVzJGnuZp1AzVb+DJ6ax/f63bpEjdAiB2feExOji
uTDzvOqC/QXB4FCOLWh5tf6ji3bQG3zCcq7BG5Wuep75e9bLKBXbm4WPF41+NtdQr9OpyP8onhIE
xUuGJzrzJ3LrR0sjrd13NzpNnQecXJ1QLRweJPA9M0i3cB3vvSl3nhBVkCthMvmJ+18rl/JLSF3K
AV/8snIz79/RSGeLZEfXiMDMWXLu7E3oU+YHNDdR32HWPayCJaf9JjFl8yQmp7B4OBPjn15aM/Y4
kBSsWDjZiQpCKiIMJUi/68+EBSj7xsoY653Alzp2TO0LbDyj7mocAQ4rsGiW3t7lx6iXp+j3rglH
QYMRQr5qahZhspgjC4hAXYspDHewSS98YVfGzIHFwa6Af7+OiKAOr9zm/kWb0PTRJKsUY2I04GIH
wm6DSiQ3WmVdN3FcmgpS67fi1qR3jfcKIMLox5Pv6e8+1RsSI97zsYh/LnP8F/3elLThbqQ1PkzO
8UrqkaAG/iaNI8eLS+huW9f60iT4b6FZq9RC0X95qUubIYhQ0IHkDelGIkvwgZT+1m41k8ogld2W
poIfG5hgrdVdA3I6RMDaVrPA9dEjnY1GkYXNb91JFXPzfZksxNHRnCf6gmgIrhJj8FYSyawKoYGn
eWf7lIl+cDIPk2kYdfYK+xRwtyagxUmw11mhJ9JS+nt0ue2dfh/b3KMWDLth+3up0LyXj+2RaPIs
mDRKwdDWvTUku2pOBezqtg2OwrmBlmahQJrEw9+x1R24ziQGtnc3NirN3HQbk3hlI/FY7kPTJL1B
Kk9BVYFnL0qN+F/T1eHgl6GmE9e7wW1CRAkm28ZOmsnMmNxnSzZ/YaHlcxUMgVaCNc/Qr+rUuVX2
dB84N7SJKhTeCEDKlwd3APnRPwFf/me4xLCOq5um6ChErl0o6iEHG0qZun+fTPKtGWKsD5KDbIok
Gg67AKVoepzpHJxlR08JrOLAWya9kfbc8eqyPrDFLS0h3/ycsd/pQAiNheS80CzupebRNIKkNIOC
g37FtVKdeikmFXHp2spKMSoK/XXKCJZNuxymPeGsCW7K//7EEjMz+qt4maxcIW5Ouuts0YEcYsqE
AB0CxHctvzoyfwH19CLn28RA1Mj1OtWB6X+fsWEEC6laG1YCejrKHJeUt1InguGhiWEnutMtb4Pk
dLLWQSCgUlpu4xFZ+0UWZrJl0h2GabsnYggKxu4FK0mCwcITbsLwkeEGfXc8zuZlQk2g8lOY4E5B
PaL1C3lFv6/wK2nzUyrSWIj5hI69F6CX9EQjsCiTFN37kFnfQMJRYK2iyK6aAl1BHwnN5Oq+wE8p
pkCf2avJ2AHap2uM9aQPjVnVszwob9UJoLwxC9ampX7q71JYvK/l4UurnTP/9fdPognNS2NcULl9
h5bs+YCdYJN80imfhB3jmVPzHOcQJLK++l3XFhHwBM6orQcMk3uPyCZEz/qN1kFr/NjHdW8KmCqS
zi4tbcdODjmMs4anDwPyHDw9dxzuNjvXzaMeS25JIBFOZQYpOEvRpgokVJQs8OBM79sFTsRLbSeh
pW73eS98TIyoJXDnfU8HaWQYeGXalEhs927U194ohMwTbRo3+6+uZrCSalyeMJ6gSaDC4Nr2CLRl
WrcWLdNbcIE15kShJ4CGceKbYFIqytcWSievhg8QhRN1+o5+kmjXQ2fadNdB1pXUc6HPz90c/iO0
bqVKjxmSTJnF2D6OKrakU2Ompb3szHLIyXlSNS9pvlzSo9uRV4h2c8zR6r1m75C9wIbexANiDUaY
NlCx5JWNxROg/EDA390iW/YIJ/CEVUPS+zitsh16SaEjoC2E75OkBKh4w3fzXqEccJZh+cQhDyAi
rQShYdzRY/XE1tWMm+FV1Jq7l9rcrlnZ3sX0ZGIHGfeX7gLp9jN+ih0Ni+/fr+nZZRKU2iGWciFo
OrBQsESGk/NfIwv89gl3q0ZGgCgC6G5TQQyWfu12GUI/cXlN/s9fvdiXS6zoy0avafdZB9XWvfx5
g+ysn7YqdprK1FZUsRQGqBYsexlAcmfaSulrZ0rkfkwTJcD/fidywMAB+Cbdiih0+yNsu09lCR6s
uIz5wwtKM/bNvKIL7yA7xkdWMTxvNkXZpxu+9pZ8jEqkmdGo0cpcmWDClNPL/ZKdXY2C1Xsw+Y0A
qHYzQsA4fUEp5tME7HL6j+1rRCOaHbNZyoB/n1teny5jKeWu1nIsJksF6rXiCgjWysFBHCAK66U1
6QHAASEFl8meb2AjkP0E9nLSX7lJYmCK6qQ+N3RXLQC3KpN6dfamOtkDEltDqHuam8Mb3LFc3c6i
v0Kz2dhG02lQjkuo6fLGHpHO6kFKDhCPDPgUJeaHXiyJPum03mcQ5g7ufdsmYBEEHb1egvBty0gw
4TLo2YCIFlwuGtaN4DjZnUpGzgCVIbpcbVCCnS7xHnW3qVEJKroSsmP8hqNxADApL3864Zbs50v9
PiD5rRfb+8+XiOTYvWOctYxAS2uc7qe7PZMbMrLaY6t7AUw9/gEk0tE3Tlm+7Ekd+qxAQbxUW+ih
/wVFQ/+ueW/z0BrqDFfI7lRCOPvhgs3cOwqv3H2wiieX0127ZKfgka4u/gUohKWieRuiGmnBd8GG
Be3aOozSNRtzN8b3Jk/IX6XubUa1yKNodq6qG84+/oQoDb/+mI5imKowhFGpVrC6Uh6CoAJ/FyLS
nNc+Bx8tqy5IDDq1O9idkN8m1JPPRr66AKKw4xGYfTeam989PAy2RUifBayha7AgX45KQgKdkisE
JSsnifUfZ//julpuWB1qbaeObkwOFjaos5GfGg6ufYge5sHppKzxV9gN+cigCCtwVAafNPVJZd4O
5LqfPdtvQkhJCch/krgta2/pAqRbuLlRr8YDNPUriu0/r6AC0j5hMb1ZSTVhRVWhwWpxG/tiRAxb
yH5kUZmUNhy2dBIDLYvP1HzMbWteTlDAyF3TqMS5nt1/yG+zIBpEPqWlfeq/Ytx2X6iC8N3NPjRJ
kfc3DCjxhz8R7pb+HLcLACqs+7Lqx3Nhsdd7cP1BbWOX2PKIh6Dvd0P0vZdMFTqSoH8G9C1sKWKd
+wxCjFimHr36tRrbdl/iTNitXU65VvX1eDuRmUrmGa+dPPjX1FUXnankKxV/C5annJxZ/wJChPsG
HGwTrLJ0ZtXI4UW7K2Fq/25yYr2G9d2fXj4Rg7pn94Mix5lFMBjT5vli0a+F0euzcmskYmcieoN6
RyUNXFi0PGxzYJmPnNhFKqnrtJ4DGKtngQlCXPQZK3PKaP7FwFPmVzGLKLiVng5+Q6W/jw0G2tgB
ljbbdOD/DdkhFFvPlUwQDlix7qXRoqTgbnIJU/kpqEkIfGSOTqeBL0Nc5uuW8WcIXzZYrdaWX3jL
qcqLjrENkRR128ji4ro15giGFM7bvAcAPomvHyzIxVokaOMCljdQHT6Z9LG3kDadoLTYQZcBJyc7
Uc6UgKTjXiwD5obyLi4UaT7wLg8V8daKsNdCRLU2Kgt6LHFBP0/NQAsFtisDHuak1S0kkYHbMGtu
/RVPYJ+rKUz6Eh3WbXXl6dxvz1opBKTPDmj6KG4qYx6cm6095gwjGGk0sN7eK5VkBQiGrEQL4nSc
/oPXMIUBLXvS5wV0yqCyCe8aun/0L26G7LjP4nFbA56hVA9rfOUgLW5fMXxX3dW9ZdJsUeahUmAN
shdoL9cYgI7uS+09jU/IP0tdU88DEz4rzVLOgKUbowsZsdW7ULg9Ym0LUm8B7V3jBwQtO/1xn8JZ
VI5O1IuNcNMStygxCNIfJEJLjbJAjcX0upRUTP73fEJAVf4pcDgWA+A1f9uIqAMRhRrdJ4sHtKng
l8NE+aqE6pivPtX513qOeRhYeGNDS6sv20G8LpyyG3TLxn03uVb4il6qBL+5P5EfKFIceottVp47
bV6rK70ciEnJsKbtBVffPCEk8v/JsjWawZk0YtDkUbhsW7l5W1IxQas06y9JiVYrdVAG/lHdpzZ8
y6dfRGmUMp6NQ+gczsTWQEhHf21hDj7cPkZuQ5Rnm/ETxh55bRupTkOCyhWpOOnTgzYbnPuzaThk
AfHs8Ru1KwLF/ND7B79rN4zTa1AqxvqjATOxdSzjyjRkAfDj2XuNmex19p3KR4b7PibPjgqeV2uU
Sk9h5GAltf+w+g5apeC92QfOTehJMwbw1zMYlSxctAutHtMtYfVT0ZPWvZqym59KtuAYRtV6bQY5
RpOrUBO1kMZMrmH2OKBkF/zrmtCeXge1Dw0yf7noE5Bz0CC4hUtr7aaMSffUMzpmFoBPpiOVszLO
Th9Xex9ppwmINvw3gUoCPtp2tGDdMApUP53mZLP/E7x9tGM4T55WpihDyyFpmrlk9oV1gGlnU97o
UZpsgNA9fvunsiZksC8frbFK3N6m/sOebKCyIf7/tjViFWaL/mF6attYccxHZeoR25HZtQSE27Ft
laK2jIA7CCCB+OCOvTtAwfggW/rJo3yRxqH4ROvd+FzYD+G+2Fvqpe02hvXCFv+8iCcRLyXz7JOx
mu0r2lv3ZOXQoBcZKSc6aWRomgZSDEtnHDMbM3SMXBnZVrTCq4d/FNd9j9PYBLh6EkFqO1VCbxNX
v84/D113lvj7Mra0PqjUooB6bgkIwVq3eixCw1DhcejlhNd7WDpZO0TlDW/mG4Db/3Kr9lw91ITO
QLLLj7Dw5gPSdgErJP3X2A7Nh/ZtX+piuWN6dahKk5AUnSvSGt44qQxRBKC38tjxDfQOXZ/7rMbp
vTOHSzQskzVpIohWkSVgnzDe9qm9oHq0wexjsmW7/oyB00oHSdo9mVKoeALWKjHyttl8/095zdxs
hXRsSe8XIpGrhrOX6Gf65PdWm3byKkzRhS5nslPNzXI2TjMnrI/mEVQKX0n/jMaAS3WtWPI+CMqV
vnX5983y3FQvqCb5dyg7hW7A6eDr6YVp61NDQXO0DW1hqhQGT1q40/wZ51dMmAwMi1YPWpZowSZP
XvzREttqLjtrv0KJhLgMUjlMHF6E4rz7AgBuj3IiFDMsgczeQbXPEs/J3YEVLc8LnRxE0+Iyb+LO
lMeqD/MwOwnpReRk2CAsQjQU27xtJ0JhBAxYcECdNAmy30mYqjk39IA/0+g3JdScRgG4+ooGyffx
kQAJI0NI+hTT5Ll19cG+WHUV8QVuQ9gGcm8Boh7twcFAUHBS/XfhsJamiBN/c96HaqqqnEik6G59
bEeUmI+MFzdP/DcwG9aV6Smpa9AEXMfFc6h5zx1Qz+0hlqQd3KiwCZ7c7/OfYC4us2Yq8ARjR5F0
8UoWQmk/leShkkH4USGr/8UUUUH92FfhkKYdXeffqsc3TQPPpQ74OSIloE/77pycveCs5t9azcQC
5m/XGC+Ovvl/2mv1swhDqO4GQ5sDttroiwLpaYODUH42LrjtAQr90a0OiSZsifF7aLtWa+1Zm2nY
+IufveIGWvpWn+eI9OhCsphglu5IWuvJ3jBnfw6XhNDfG0NcKCyl+cvZ/wo6y0zM6rfkd2Do2Viw
BkPztOdKL4BJlhkz9RanOh56omlvT3dCyQGk9R/dRz/fx7dYGOYMfDhHvBoCkHVBMtcmOh7C7LKa
xrgWNTuRDJCAoADQQ8U7gLcBopM0XU4hzsU+YFUK7xN11rZIMcSkJzJhAniC+Bfemn7bpNAkXqg9
rMelympTpFOa8PI4lcjryslVkXqotqO33zxCnamq0yUfU3dDIaW1skliEIjxPlrQ/VFJSbf19jgx
OiDQdvDqXDwhEnwzuMr4ZwToQsAB6SMM1dMX5gXLX2JWiFkB6OKfxxI8iEvndGrFd/UWbK5Dn7cf
ked/TrsUTFeZk3fsk8lRKJYN5/WUZTXGl1l8xSdLiRPHWgxpQTmXJzgSeW43e402CqfKnh3agh2e
g7VJs2jNhmcoXB86zJPcc1KY2lpB5axZCXXWmspTz6MpytLG7v4ZjUx58aCN9YR/DAn5vV6DwPyC
PRhLR6Ztlxz4MFts5ElHSmCNLsWMqJsDDRkwz0zcjEB7pAOZZ+/xJ6tUTNqEGxjO+hPslYjfXn/W
NHd6ASN+qHXovLRRRKLhU57N/GPqKxCoq/XaXlwnNIHVLV02lvwnn/w/heF8iqS4gaxDv/iMvZOX
sMQUK38MxWacknRVWmFOwSZtSjQgTPUfFEEfqY0tyOX22pao8pCqx9Xc8kwqB5oGBDI2EUVhTga1
7sNypuSIXGtxUnBC77QlJa8udA1MpB816h5iL2ALD5rmYjHf1b7xEMbDQjEbHJ0Zri1mlJkz8aF8
1t8Jj1TmVJKkcnFmHcQ9tHtf/uZlzn9Pl1MIhZ3WMZvZMMT7PmTppdxUXe6cdE28VsuKjDKdr/6G
R+W8R6mKFYfTIrH4EC4Jw5yzp5LRpde6P+A9AvzhgHBriCTUPFVh+SLMjJR+QRnJmked4/hEbCe+
II1c2XBl/HqDQh3C+k1Ahwwvuh9b/WOg0Uno5p3jUts8AkU19/a6qbP4UN1dN2sZNX1IVywiGidw
XQu36VjWN3NnqoMZ0lDWwsA8Gqmn0PsvBGuil9RTbbRCkqEZGbuQihMZswCNQa/LqfiwKnm9Obl1
LxhxAneUfGwc27ChhkhpooYqsrQ9jTWcPgO6tyeLFaf/s2R3XoyAL+jB9IZN70FWZps1L1secvTy
cZmi0ps1ljG9OG6wpaWqfpPYad6pKRNwd3KVIRjCNdC6DZvx7tcd3WmlqyjgB7yit9JGM+U6G5Lp
k7Lk8J/J5ydvHZQZgpj6q4MeRNFoHXjF7n8COHf7/UQqOQbdNxh6Hf8dJluW5nyFvwRRjUsZiw0u
IzivyCM10s1CR7xXe36ZPBOFKV1QoUz8kQwU0GVhOBDB8LKJjR+9JTj1noUwqe6G4p6krJJLy7Po
qUbymb11gWlt1hzP220dZcC5U89Q9cX19kQEsuQ2mmFvNIQnjLqLp/ZB7NOL6k86CLYpJ05eGj0w
Wv3+WqI6zOsRJ/P4xHn6/9H7anKkuxHzJ5/2kzA/aHPxiERxLzuf3aypl9Wv5t1Jag58QsJjkire
UFAfuI6gFbxh1UBkumyS405EUWf3sk9PC3uDg+frx3FycG6JxYlNqfg3r4zDKsWVCkLYZRAYIoxr
8ViYp0xXMl0bHh7RXTi6WleJZEBKxEWmZWUzrqP3eXnJOX19bN2+/4aTHySQRnfp4aeG/Lb2Rf6M
5Rfi8G/4bE8ty93g5xDKXmCFh4ZuZwMB+mmk/Fd943c9qfZkfoV25aOaTgHtp0rPh5ebGm05DIrm
2DvcZ8Dw3vxqp/nbc9YZ886VjeNTDx677xoQuNIbH6UDJFT4eiIEaMOKbbnupcRtPh8OPPeFikDd
Sn/UXir6FvpN98GJ9LViC81gE89ztyUrBogQZLM05b73/9jBAkz09GCSFoF2dYAAFQtSRbavkKAw
D8oD4pWAN3Pm4Q5w6gUugaHIa+7+1kUcUj0TSY6MuOKeCcTxS6pJb5shEnBgCDU1C7Ejz/UedOw1
GlF653Re5qgN/hEAfhN3hTdugiRfOiPwRCfJ3nQDkIcvYCDLySxN9LtG+lOn0GURsi0e0OGK/PN1
suweUIDN9gQUQJ/5G74ddsTeNmTt4HjlZKh5jNdClTJG/eOmZ2onbcKbaCb3Fop/JejSWB7uxWaW
C5RZIIyV0nLlZUMUIeNNVKlU3aCdIzDgx5KpS3uVBGhKYuFOPmLFVt0IRQCrJxFMGJ1AwVEGlh+c
x8onLSkuABAxPZgeVpH6mpFvl7ahxlwLgaY26ca9msowSuxSgJtICooHNGwErsI+q4WCKDLKg4Yn
MNmKtSJvdqr5ptCTtv/JtRD0XAyosdbbWrchhaUOcw+nwC0pW6OrqpvZJkCLYOnDCHgpjVrpTyXZ
gTQ8TfXpYofN6Ocdy7thLmCNf+z9fPaIaBuYcNua3ghgeYsj1yUngRZKDqM57Mx+pLvjHZtpblpf
24I2F/1bpL2Tjm4SSDKI4BlqALzI5mjWneDOYQqF9Z3W5EbYlFGYEF69Yck0FHQrRSNKVvksLl9n
3PqLXrsAtz4tn+v5HJ/Q5dBSxR06g5gfx8KOUrAKwAf7hNL3Qi5jEEh4Snw67w/e2OF2TfTdskjA
0bviIsXjl59TIqDTTW+xCarHa5QfEXlLYygLTT1exQ5UntKkhPfZYngWdJUFxPe/e7rJh+Hnjuxr
ORhgy4ALo4kLNDV5fYLyPi6TXUbjSIiy7jKXtQLKiyXv6LZj4e27iskICaXqzPmUhtJyR6wumC7Z
Vd6L/CubQlXo7RFoMGnoeyQSGrApkhLHcB7InacI5VucRC/vOqYgSrwWhTlIH8AOLNA6RNluqlsr
xe3XC8plELJUH/GDssiyW8nsWGwWcqDgH0kx6f85waE7LDZEYt6lMUl7Mbs1PRhfAk3JXgWfFEnA
P2lZ8Df00M/sAqAVSRGWp7tQt+YQabweydsl4TUBv4GtYvr4YJ9xox5tm5LjZGywC4l7BWej1yD3
AlwNc/IjWQfVkuibn/FWtgtV0kO/gFNoD8LEyTRjQg5x6TxSWjaEIG8UFL0Q+w1kWYdsNZH+iwmx
82CsKcnYeaLsXhp45dDVpVvoAxUr8wlSqur1CNoMxdUFrr3MTSBnLPNxVtAm9XPEuo5qPPTs7bHy
6SHyZNuI/0dktsYo3yWBvmjwEXjmH2hWZVrs7vpqTFb0vLRIMPpww6MSAtJh6U6i33GHlYYAqQAN
q4Kd17IaFnUO/7znrE+HcfI7wUATXe8qU+7ps3ern0aZhbDj7DCMYWBRlSCo1WtSJ7AjRaz4NXPR
mAlAQwuGc+dknfgYV4BYKq0QfZ9OBSflz6bvkh+hieTJKxnk3QKhUxP1lHdQIzvXpyoDOMXuF6Z+
ktjxA/YiQ2VF13w/Nf9jilro2VDj7eb0ovPLE0vhOaa+NfSTf+jUkf7cmdiPkFKC0ZhjP0RmcWEN
+f+VoWHdLl5er9sul4zOt9tf3zwPrztTgdfI/p/lWE1lpcMTTHp6kMMYPh+OHXaaj01NASyQz2o1
c1WTf6YWoRLUqYfqdEhh6lw51LUIU7GhekXSIXKkSskpRS5kN3LG+9RY5OdM+mMhBZcdPtyVmt7j
ZBCloLETWppGFbmKQGPT1YJiK7q/UmQSWM9/EtpQ0qVYJNzOYRgSaD+SIvxnjx8lv0vkz2fudKT0
fkLhN4jvsU11WUr1wEbW5XWZyXvRnXENy3aGGnPBi6gSr9/2OnTXgalnmP9feqnf3PQ8576LxpE8
XYidybednLbktjvTwwNGRSBCjjQ1cqhk4pFG2iqkoYpphHsl2Sp26NjbTJDufBYMWtWfLWxTHx8D
+GckpvFTWlG8shblhLAeNUj1CqKYHweRPYak3/6pYnn3Z9APwIWorbeW6qJ/tNqrYsAdbgyA1zXw
4ldX1P0HYM4mmQRt7eRFnvSVm5ShzlfPd4ME2ZfX/QwJsBOs1cSiBVaa9wbNTeYoK+wZydWk9pup
p9G8Xngj+kgeE9EWcM83XF/A+7lauQAohp/mOFoyBL7eo/3mvt4XNHVpvzAXWMqEEIHh48PJkUb/
iwU3jx8g1G+PBxaaxQjru7ebSfzn25gjTDgF7L6w9kUhM+JbtQGdj7UdtIYPzmkPbHROJdY0ZpHB
1Pa6X+dV5CU9KIkV8/YiYThELG+FDsuPBzaen2Uyclhe4GX2M++gWxvIQjdqlVuSyQjrUthKlZGh
EiCOj4l8toHi4dN+t1ulvjHkia2A2T/IQvNLP9YDYfe/4NuJdIDV8R7kshEutUF/Q5+W3C3QSegC
ExPA5BSabBO/vhd8ePKDRh9ASvyyxvEkgHuG7z3jY9ZLOn1aWEuyp/lq3GAJ7zGISkD8XtHUzyWb
CCkz8vKKJ1tcAQtAeit6dnW4xr1G0Cs0Q6Pbxxx5A66uSsaaGYtizTzI/OyjP0O6+nq1kTJHQwZ8
JoQ+yeLKzTD/WEJmcfR55NlGJT9AJE1f7lbKf/012+MK6DFL1jwqu7O16C8wFkJjB+NbDDQWOtyk
bx4an9a/LbQXX0zfwltSlOtkw57VVjc79Uh/F9pEcnmvNqfWzMZIZXpyT0BEmBimRDxyIeF3LVi8
blTnkbOhcJo3LTBKrtnG7IGyw9mpo7y2Q8cmsTj7n4XDJJgIjuJlP5yikLS67qU0szPZgVbBOzQk
4t4mykD5wdmWp29Jj1uVC1W02wdrWk100UZ5NZgHT7TjYFz/ZFjkF5CdTum7Z/hB9x2UihTdAteZ
p8Wd1OY8+nMzAOBgdOo6hSyrsABchD+QhnWndyTUyCLiabCf3bfnMhawX8sVdJI4hyxrhS1HvRwf
OpR/H6bJ1FhXojMt45GAn9Uw7T0oBW+qM/cBiFnq8+KQ8dTNYL1E+2jTj8JNWSk7Pa1VyCuX6y7u
BVBICKyUJtW9ohRd3x8/svjtUy6JYqVuInk8GGIaZvihTGdnUGtUq5rwWDmX/+EG+OkgPhJtJFFg
PBOYmYRio44W1t/dkq1m2Z3sCY7HFw6GgEfsuQa7KXCb6qIMVPMrJmSNHN3cMMdaMuo5zpxeAYwX
kCozJ1Kz8LwhABs3LSmXimmRwhIysQbmcwhp0xu5zSPM94Us8KJ3L2pPnC94YOGWkkDdP1JdcRAw
wzCzXNRuwvDY04BQUDrfq1o2HhMeV/vp3E88eB0hVLURet5qRS4I7UXqg0TxzNW6FLu6iDLozjkv
Ggsk9y9XeJ4AsoOVFVVKJ5rA/ha5pM9QsCS67H1uZXft09gI23EnJpDeSfCgBEaiB6DKe2EEWo0Y
uaoVfdkRMIe+qtGQr+7s8vBuKo+ylkmuoynuBqOidsSAjIOp7dUavY/y2UNfnKd6pzLl90JYe8mC
dIXSnHgr8HD7OkHHRMLd6I3ugZEJI51ZjnBw2Jp5asH/7NlgQPY6z0qHzR05K8CkDEUoOovridpX
TIoRsnLoPnqTTjm0tnXhnFdBRgYnuyDK3Azd03P0ZQkKPARHDT4QljgxEP/u/Sx7IHE/MFXoOS0b
b/dvHLc/+vybxdiuWVOxSodMeoSQg8YxuBq24YqK4AxYNfVCHYjlIHkToHfyr6juQjC1T1otoiso
VyRat2IIF9dRI7oNBhYCiT0VJ4hp3wIw3j0zbEB3MbY/2RwV1LeC82L6UxwPPlPUb7XKUw79Yqka
2Vez0uk6XN2qXgDZR5uFpFsUKI79Z+ehX8QS26J80M4EojSxmym4s6ej6Ar3JlQZ/YMqE5u6rCLv
/Izhz/ZMuBOfeD76VooggAt/OykIOSkz1DZUzYywHT1ShtjFQaXlyPHcYejUheMDebJ3esDNyzwG
BpYpH6t8bQ/Pu/NiAEkt5K12+A3dLvE99rJ3e+F4FVGL46YHIJbvrSkp9FFElw4ZgMq0wUNYGFsb
uSWif9DhcPViHKymtK9s+yv9I9QBiE08JVH3J+T4ts8Mn/yEGp2eOawOOg6lHlLJqzhMEIFUgDaS
sfC7RGbYilONclmhwpPYhbmZpWWenhVY0b+aiKxFf8+TUwMVO/b2mpYjr9DdVUhv4J2O3qYzVWlk
ABkfbfEz6xpTwC8xdBd6Zs1dd4DbltMVbpSHJdSeoj5TadN0EevRjSxvhE7TDTXGaNzUEGDJ8akM
+H1sL7nTn1tGK/x9P7+wasSmaju3VBCIMP+WiWUhiXhS4ajr1GnACDApnwKDPA0I71RkmqD8t5U/
5x7RcVUjV7dqUjUHznHHVu2P2/7FYiHBnfHVcuncd363zZ1TfKEI8BOFojO+kV4rjqDduCXYEFml
2sOk2RkSm+hx/PqTBEjXJv0LZCKJ+0xHnfQwkcPy0SRz/xxntRVVrmqFsN3BUx1zS3oie5n3KBbT
IcZlSGhOVZDqK+wTNKVgf+sA0vKei3xfw49C0kSD6s2c+kxZSdDdNzxkFa3ZlmjPXb6GoJtWUkUU
R4vnj8Hu3uRoFWcFPM3i07a8AaC0kF6o3JKr+HxT4Mu6/5KGMPdzi7+8ZlGN8XNBZFjFtaFyP3WG
8F9jdP9lpnNKdIcr55m0ecqxtffIVHRsJoiAScU5EP82hOSM8XlMAgA12KoWYE5sWxWVRVZgw2DS
i1+5Syhotu66LGsQ6y3l+nMW+AtTZJ8Ns4oEJSVF3T3UYV++8WolyiG2HPMDOCXgUdk+1WmOXyuI
iknSzH6obTPe0BipMYbZoADd2/kwutNsivx4LLFBczA3hdLmnYsc33voqdwO3qO2s/jD5b1AVlkW
e2Z2VUUD2GFDdWxjuGW4aYD07VMHLE5d26t4G+cJnfrrypq+PUvBxWNEYCHLSIwr9GlTg7Szhm1f
GqbmVp3K7dZeY52lxVRE+NSTKiPgWVBUAzOE7Jqk95uuhzE0Jzy2PoUp5GOt8n7D0p/xvi7/Unjc
O92vaA4UJz5tDdiNyicI0Bo7rRMF9639I4AkiBcsyLn9oCCZfhw/axUFswJ0Z9g4MXCMtcIj/Ccp
DPYlTV08p1SUw3uKzXb+qyAnE4xuD5NqX7PFGPrGd9p7hBjhqmIZ2d64eHqu2g2xrbGovAgPvn9B
9DrGMcAPQ1u4RmFVbVzxyrA9uAfZwb9s9g2wTGrVdjAZ/SPaKR/MperGxEQBdhzQTflwSSpRZuZq
SKrgpGixJH6XmjFMNqObNSw8UKf28jWM36E7gDCC6U6uZwb2tc+nyeGWRTY24GWadgeXtxxiysie
jHGo3S4kutGTDRv3ZIh+3DL9E86SipeetXYlc930XctcG1nz7UYxQPaaC+0EU2z6mCLMnZUEJggM
cS8sj5/Z2UgHwLOXDdg9d2vDJ4o59dutgOVgTedCISPdcQXRYWG9ftJoT1GfmpQzLNGVEBazHo6w
d8yukfI2WoRtzD2f1PzDgztRSU6bQj9nx063F8dlHMNmeF/zrXZyUbcMagHuCOamkK861n/4C6fG
k+4FCrzbXnq6SrvsDkT9hMKzun+aXDuq7H7nj2qW3Qbe5Fmhkwe2y5anRmZOm181dH9M0q+LoY2U
PADs2sGwFT0Iy4PfcadRujov1Tx4+ktXGnnZXBfTqt0CEGaSooFrfLMSxhRyDVk7CKdIA/1rPWTb
0gK03LZhLcAuFTQroBwXS9cClI3zXgBCErzFYQw3vl4+9lkO/tCXPaYIaEr03gUrjUIGK3sge7LS
6lo+dd5IB3FKtGE/P2mls2pV3R1xbVzr5uSovFEwgufclKURhK2XcY/em71V5npXCsxf8y9aF97x
J9yWjHLDCyRibDmxuRp4swCFshbhFzhkkuNimKiHu2nRRok12QHtZm8sGba0Hm/kd+muzdL7TYOR
DVnLRxPdBleGrETy2ZUhWl9yxQUbvuOd8Xw1eT6u8XhTmRyGwiA0iaEdhtERwsrfdiz7AjQr4Ynt
3bbigVMZ90znSAsjTX3QMfFWSjp38FuDxTfD/tzaiLUWlmyuymH0t6irRaZJpOS24BuuqGP99eAj
TLPl28StAMX1zwe0J5LtmkZCYbRIlDltpFQqsKd+deRLn2HwKxSPaJvft7jWkxp7iA/sIy7VJChR
YzJ+GTWybnBooH01h9r2M1sHA30lXlhlP6vy+mk+zDbL+1cJsQgc44Fs0iZUOoZxHPezP70cE0O/
wPV7p1yusYBL0JfDR4HnwVlRdY90MMSntQjtDBcNxo/fV9L/DePf8xH3C69eXOIkyQ283JGPJqc8
JDY0RgRlB7T+L6yaotgrYz7tju0PbKjQRMQ5VKAxZDHg+h3kP4zYUe4zphjMM5CA9WcEXREc9Yu7
4/dvJrXgt0cJRWCvZvS9Gn82ngz+sLes5RDkoDC7ecuddfvnJmIRA5gzPqNhC5qxMBcJm3XoWmvW
7jX61Vxa36aj8lfezH1a5dvvvjm9ZEeIn8c+vUnO2i+AXKnbe/bHgN1R0UlWeO/vgdEE2JZUcvWs
QnzeLTmJEI40uH+bpSPdgNKTgygyAyRZs7k5qSQNb49pNjF0B2F/Pbxfgsax2+QtGi7QtfjCpm7k
DfDebbGsGdtzKxPn4rBKv87HbFEU2JAGtbwvYovi/3HO8dY1cLBqCLd7bfj7/h3Xs+DsJZTRAxG+
5AxYcNu1MDBmnh+9lZUcrBbaAD7bSEakel2STHmkwpIwUqqk0abER4xwucR+FdN9j6OAUA4FU8w3
YnxVLcQioEvNY35jpH5LytDWZ7KnkV0tboOsgjatPifMwiqMTzAD8zWGdM2Fw31Id3MY1ptTgeS0
UCKwHOta6cLEwI0zlGXvJvqRS+FIZsBPfXtTfeuAV3vICmyppn4gZQW847jPH6XVcwbX+Ad0SNkT
7INMInCpMQNOeg1bl3A0BMqDb+B0upwm+CiUn3VxCgrbIuwoA0RhD4cJt/OpWfdLYw1qp5b3H0fk
ZYU/NRO5FLOwXGZvK6sAtHY9/KrcIlm982u3XWc5etp6KvmRma/O4YVPtDYyPgyZgRO+9K6otpVG
0kD1w0GMx12FPrSkA+wlkMn285MMvDJEaeUAxSI7/oAHV9oHV1ijKk2JbjuGTVftCVMHQyFP0Dwu
vmPZKBQudQKK5jJcwVKwNSpZ47x4cfmQhlT+VmnHFNtwKm/WLh+xJH5iso7BFGn2dWQty3EylbH0
X+oqMfz/ExadE/qveGhFI1V7tNN8Nqz/Za6kagb3yi7NjMfIxp9WiY2RtH5w/NvbGGpbAmkVtk4C
3ygIkHfXO8PkBocw6HK1FtjyRlteVP9Qj//IA/NxyDIFf+hRFUrzlmvaT3xmNQ+wRIG8poPU2s6d
rtcMpkMDFGVeEdLTBJNGD77FdoGuSzAlohm4HBk9FSCCHkMS3POou9jtEuhlb183GdX/32/svwtw
qCeSh26vJUsU1zbCClRr+O9qbdBcE6wLzzOzRmbim95wCZTjT8DpN2LIqoGNIxd/VuNmQLG8WDg6
XAEPFac9FQPYkK4vb95Sb+3ALuum+hejOGyBYo/FHKG0nv2e86SHYBJkpzxMbEisu2zfyYX0wtTA
+AWJe4nABvFQtLAlS+rT4ucc8ezD1ipRy4WYrfS5TlCXIZehI0SDVCLEiaGx7FeFHMwz/v5CpoiY
pXrFXk/vAU3MaIHxrcEvkBdBwAedXRQt6IvwP44iTG9aFbl3V+yTSzNJV8cRPMx6IBfJJUahPEkl
PGEN4j4udl0HF9IsVkxbgcWsOZQbe9/ICOhHMrjI7itwJnT+cBjGE+Cn5MYJxO/RQ4wSu9URLY91
wJhJYjzAJsnq7+5e9ymcy5RB5jt8CgXCPhAU/syVOlkI600XwraydRFza2wplzg+hrko/1Akf8Ee
z4blozX0bzqPdPRitIgavKNHup93TcvEF1XS5D10edjY73xJURVh7sCZrWXjMWHrKvS5lE2AbFhL
6MO5xuCLjAS4TuRJetvWqG+F1rYe8/oSk6R3hAhhfjImrY6c4Dg6RXZEgXh1PGM4xHZTSOwN8N34
ZHsNr6kwPbqpfaDM2iup7qXUZLNSRErTokvJysv5zXfCsVU7NUmFqaE89MhgBC+Itvus5sbFrYOG
qTkGK1HVV1YGnrDy4p7i/lj9J0W3TcPmNtVC167Q3P/0B5DXqnBNEWqcnlhgFZFV5ovaVpV63t93
Rraa11rxZSRNxjHxeCIvo3xYapQWlfr3jKIszeRB1JbQVkxXydBP6VIP4Lg3xzRKVvb/GJ8rp3b2
yuHnRs3WvvOtZrU6YsHVrY+0WqCFNg6yb5ttj00nN56FBQm1oXJToHGwa2G1wPfMpuGp5hUOx1aC
J1QOxSfscVszbHBkdGWPDwf0fAsdGnUjzYL54IXQNDcJcb040VVBdFdtW8m/tq2N46A3UpeRsRlm
Bn8nbfaqRSHfB21LoQynwM+nL9wrETkWd+if0nIf11CabRrvHo10U8iUeqyWJsl2m88MlV782kB3
WhqTKm7ayvUY1xM7TtE4Kn536F4ZDDdDzTj1RQKjVLYv3lHKm0GXBWMGSA1GZrcdW62N9IXnroFk
mrsWyRN5qzc67OjrTAPwN10IQon49M3yGgG7z3Pf+Znk8vZBtQdUN1HpTzwr1jWHb9RakTK6YWzw
BF7XIBlJ/LeDj4uC0UJNnAXHGjOgRLo7dzoQof+BvZoOnnHHd6ijoVuxlqVC0f1n8gd+plLNyOIJ
ObOscet5wm1S7Nx1fM0eZoaobjYaH32wM7CmCg8CeZmxB1kvefRB5tedsujddkqyG/uvsk1wmFer
AlMBUiIjVFMrIDIkdK3mWpAn33tC8G88sR4AbesV4u3W1pofqwiCVRYdL3UB0gdCuaPIkfNSJqoF
j8rttks75quUJpSIyR6APiYzFfC9oRrn0LWZPabNPPgYlVgwx3xYyk15+N2gx+7FlPStNFwEIUIa
cWCMureeW8ho7o2bwNvKMJPeAI9rl7TbUaESwfoImCoEpWzNikcw8j10xvgkjWHlVmlyhnmD9cfm
BJMX4XJp/0wE68KiUc3vgk01fFH1kKPOHkdUz+osn0+WJWO3zpSQWkI4xSEAxQ32x4zcyeoBMVPQ
OP4VhnOKLydBTXsUwtOTTEjGcBojoCOMaaHkd3KicaEgkuPJjlL4vrwDS60r/ApyE0dROV0Tp2Y1
FYf8UFK+6EetRkou2Oo6tNkOIeqPJMluINnUdwH94zsgWHLWqEbaCVQMPyyP4fchTWxCRkhFaqAW
4//fOOX9CTea4jtuOKCq9jukNZQ0fYhcsfP2Sg7kqRw2eelUBZgMd6JWJ5ZaBcZlNfy5XeMGSsRX
y1V83I5CpL5+lrxYEq5ShL2leYOjOEF0Pxxx4UstU86B11Enu5xoXnVbpU8K8125/PCyBhYx94fP
pcAodBfF52NUoUdp1djm8hDYXLPjC70GV+luCYr1bGGpJgZXz9Ofr62WkeJLSuKEi1VsE6B2WzGB
MvFOIN1/VTMbCxY1nOFazNQk0Yu1FbW9id0hVsymTGFJPFytxLpFGOfVlofe6S8pXTN6NNqZFgfF
J985iI7jyeVhyodD2pAMV/2iAq2mSNsubfnR/yIfY9NaGInaQ6cuUhpYN7mB+uG+WNNLhu/LR5nc
/lilaKv1y6BaH+PuPIfO9ZwEZnC/TTDKaMPXhtbH2ZGp2CIF/Y52Z+3w2EJBG2tRdc/RjbWOmF5+
pbdNyj3vwXbaVU3xectPPqfJxOnVWCBH4N4Vt8mC95xaVSApwz3w8ZJPOGcaQo0AvpbllsXgdlea
kRaJI9xrmN/HZWuUO7yjO7InVfZhh0Iioo7TZpnnrUxmmRGNd/TotCgqH7LEWGFumncso74mnhml
CgLYU2fYhRYqSzBAHqI7DOKAN5obPoSf8k5Ioic+cdgxp3+jUKHwk2Xp6ijVrxtlwkpINtpvNat9
mDLtNjPF2fk48sq0soB/awHlTEY/a2+EkauOod6nLY41B6isdiVEipS5lwBdASf9+4NLZ3YERgbC
Vtp+a7qT8/SLsZDACbo4F2E+mm5u2x7aZbzAR+DJncBs9TLsXKw++6MBfcWIVgvOp3UYrKtJLWrY
CKfY5qLM+Os1grtwxGAoApTK8VeAGLwrXo9io4usWPZhnon289bWtDKrTf1hZaxc1s82XFV4neXg
v/7rBGcB2fLTx6kik4/48YU/gJSt3rAtZEVkqV3n0ZCkJYMzdeleazX23O2aHNGcXGMIg1ioPWyK
dc94woy7rx4RaSJwVd4GjS/Z+NPCaGlnQw3JPpm5rz9kAiFsJxlPc+VWJkkBTVC/eVvQTe9IQwcA
lBGrZx15k9AR86q/puz+MdABbB1+JSKpCOJuYQ4yV9PriqNGoend0GfF6pfnFOe9A3Wegsnu0T5n
Zl6d1AZtPanfdzY/98sjXQO3/BR0B2cSGYkjY6GVJ7JkwD/W08HjrfH+Krz2HlUZERh/SMLTEODH
Tfo30DBYM9CQ2M/cwFF1TaE0nCbCXKJkQX0Tm+WX5pfDQYM0uSZQyoFQaVbeYO31Vy5lxi/YMKRn
Vb9Hk2V2t7yqchC5AQuMXyp++7iScTrxnaobUFgFTTIJ2Nx44nvX5xD+MXyK5vaGzcQvLAoKPuW2
cmEQRV3zRJFhSImvdOOi38rOu6fK3ot1D2Ubqz5P/WtNlj56ublFZ3kMphM8Bfd+gY18DtXyP1i9
P4tjdvwCPFSXsPw60fSh+yd+VfWJfM3/BcGcdbP4B6GP/Mpfu38fE/Cgjep1dLJkWg2Pp00c1i9O
aVQlHqV5eK1NpZ3/1LUY2qGiI/0cHBZasT7ffhXaD6+RU00kCFCl6GkuEi7Z9C/RLV6Hzu5M/8hP
dDbi82xttjQMkCJ4wueFDqWaagSXK7fU60Pgb1AYybCM7TW62Zo5UYxLDq8DLr5edEAA2sWNaODf
biPQ3+YAFeHq8+Pq+Y8F1j8E6K5nLq2NhtS0yaewatRIdIO2+0TX6Y1NXT2dSe0DmLnIRCCdY3lk
MuVucGFqrfmcxvW18rDphCpHP2Ku+Z6jgoYTIDxC62APks4Pb3nWnf5IpFKfoCsQcks6YIUHYBIT
nO2hKHEiTZizIh8eL+nXl5UIPIRlIpKdiaApc+dFClkrvyxlCZKHvPXkgIQtLyyclB5D/AMDnesn
+DboBRoh9+ZMWNwKUbkLcyfg2wnWQhpoemcNUn5qxJKaalHqVRJ1QvNhzcbYUnfvSnE7foZaO/j0
WFGRlx7JGX5uF9fhAx5RC5onXiZpRYw92vQtturiep/bcKWBrVy5HrKckBf1YNTmyA1VxacqhJxz
T45JxutvFc6b6acRcQvGdpoOWuIHFqlnNd4Mvg7wMMs0AKqqAIkA0HVqEnaBEpbM25pBjnru8U2K
E/EOPOOc3LlHUIq7jYnBtvtuVVqHcZQWR0Qv+ms5Kto+wbzeo/qOzPovRo3VXOchGyaSomJ/b5lD
kaE/D3bTxm9Vi1LcSDuTntX5Oj2ElOX0qCL8I5TnjuIIt9HVNAnsXlbW0fDBMs5Mp/nPyOX9Npv4
2IKLMHJN8JNgsFk+x7yxICJg8zG18dfQPe2LLkCQgLKXxM1MaGc8AwIqddWBL3zyd5Ne8Pg2cX1b
uNtltPYBwgfHfH9jfFVidmCyGUZgURpqm6MecJM8MdiRIs8nbNQ3D9SkySlo7eVADMBPZbz3rzna
HZ0GHL/ZOjFiMdd466q0GMd7WxVnUD3bXoZLWYGmPcqP1DLBlG0Hn+iKlElbsf5YMaxbDnQ2Jynr
wrmtHUb2yiovu3bI9bjlYivcOu+8KBzumU7440tFjdSDYKUjTUNa+VsBaWPCtIKsSMHW1TAhiALk
407pCMmM7+p0Yp8rQoR4w3rdpj6UBWcNXehTuOgq01DwQqG9p+JdbgObRSf+lemJ0lyOfQTtdSs7
F7IkHM9uV7JZjq5+8nDqSfkUkADu2m4tpVfOBK2GCkJFEokPRYaruF1053VfUr+52X6PpY/nylIU
1fOW0kXocBJrTYIfhQrwwXecO76KfQFESiHqfKhepTnAnA8uDsNwzgg7Lia3lFuQusfWb2m/dFQR
06eSjBoq9HVeDa3Kp2D9eISifNO2ALu/nG7bAdtJhS+Xr3lE2Vqi2IBD6iMrD1q4+AujWeofdxk/
ck9qUWe4N0RSZEVnTZ3bCmzUhClPoUSc250WTiwUpmGql2SaGzf0Jr0BNgQgp0T5KglZoGhKAHYO
CRcAuYxOFekueF5nFYcbhoD8j7rMfMCUzzTw/TJ3AVlBWawE47SJCwJGjdi/7Z5olHQem47q+P7o
oC7pme8Oz79txHz3+klQWxC3RXhokfYGvtj/9H5XAVOIwjZcfB3u5lJc5fvMUiShDJf2v8o/ZP7T
Kp7hIoyATY9neWNcJ+f91c1aHJmIjBUuJVnvuWd4Hu5PNojcC070J9Lv4DsLK+bxZBFnKIG25e6n
q0iovD2SOG+ySf8q/RZQFWamwpo/ZM9bRcZFAnrCcYgOwupQk1XPQ+FLgizM3EKPYuL62GbDkwiW
PNoxbZtGz282ArcDz7M7c2UHRDyz1hJdGtktiJ3yToiPmHH3AkyY9Nch3DGF5E4P7iKChs5Xr4hy
0JfZIxV8sLp9uJzh3NOmE1yRC90I5YcUe2VTMinUBe30DUe1lMkeY+DR+LPQ2KEciwtXK7NgkzQ5
pSdQYxqGB9qaNBI4ZROXLDv3ZvM6FXnwrYoAHYVyGhV6f0cyl7mQXv0PNlNLWWH6U7tOO+di2gBv
Bo4misaYD6UPH+wVwGoFfpIzhqXbCRGwRsE5Rc40nYFM5Z/MzEP02qsQoNfJ2y17Ehsm2Str8UN0
frlzJYLZHN6Lvs0M+rcxE3WJ/hMVX1slzDN/S/dEcWE1MxzYZeD48xpBk4POwOyX0ZwgKaPALgdb
uBvyioKm6x830IU/OSphfOMpMPbS7WzpKQ71KBETY0HeyCEopm+sCxCQer2/48QmqqaXwEVPG4fL
LjpUnuFVJxLEv/x32XdRU3QiOVkUya50r+VhS6GgDjZjwPbhuMOBKguhK9CE+6m7dDJMAQzLALJu
mPKZfYAeiT1IbpQjXFJTz3XiBxFsjZGRH9JcNRQhRnXVBr4o5wvCBel3oBmfkNlEkU9Dls+J54Ap
ecH1jNf16/V+inLvJET4cZlApwhgZHD7UUg2/Q3VsOpxil7fCm7qBnixXMX973XIGsrX1uNY5sKe
QzIy74T9gJrHqGaRyTuGyhX3p6TJBc1OrY5yhEnZEZ9ZEms2NbNWZ78uvm1e7vz9oLIceNSdUgkd
eJpXNNG4o6uiz7FvY+Wpu2c/alaPwUXzf1uXR8rTagTsmCwpXjKE2a3yU/Pm0s5uSpuRINSq1Kjn
4V4gfw9RHQp1aTf8fPsgx9vaYuUv5goC4KE9Lquj/z6A8IjF/f8hTOgzlOHUhKo6GDRG0YeeGed4
ZKbzT13y47vq6VPVOgVX5nk5iKXJSa3PwsNbRrQtl9HlHfQSUh6OhSBBsI8AbvPAXRxepPWHaNT4
cGAA2w42/FnX3USzylKctz9F9vVw31We63rHfAA3myBczju1kyjIuIDs/RmeAM9pf4zu0UpFjshn
mXAQWBSCaI4WDas9216w4i6VR+4TVtLAtNH1Hj9XP17dsuOwnWPJjcWQ83Pos+ag6fdLZwKSB0KB
2lI7bf6cC3IeV9zqpMPfpTB/CzDMkzhuDuMT2T78LEBdKcW6ZbajqjXIZg8DHOyi8Z9td2Jc/UY4
HDunl9ZqZ7QdVCCGTfOHIV6YbNBN7UQm67XnWUPsVZ3uVmHBnF1XEOcuRVZ9bG+AUJcsacbpK+0l
FRj+5Vhwi2iWSAx6igG9LzY0nnVo0/g1rioPjugbNxdgZDc2RHGd+gtoXCIx7VX5tdTEhvdVCdB8
J2Lv+PeSRAPZ4AVjra/GGnN4bZM4OK2Hd92urBgRUh1j1/WnXu8edFc+Gx7kgaEj3YD8+z3XhqCs
gwOvjVRQ67+9paMTSB1wyAUr2UCcgz1c6/JHlzq58v8YkjjTRVUPbOQOB4tmdz3fUyj0oxLMLZYZ
9k+3zsyPkd960NQUfPSzTngxy0vp3NTCKjynZ6tuzb55OCJp+t5x7IuN7i3oLbY4J6i9n8WUSIYR
17yTvr6EFarMnJbqJ+n+9k/gSOIoii7y9Y1pwncf6hZxJiMqNNmd8iysSTRHi0mbcwR2rXiYvh1o
TnyLtn78CnpA2s/+q3ZwFxF+NSy3LxyQrkaoPRYabzCXzn7TilZeIRdhV6Veh2MUpwEhlnlAwIcT
JCRWpy6+pzF13slYnocIh/YriHLojLtoHl/21a/J7lFSTNJIjaq5g0PoOLnsgsxYALYyAnRgK2cD
bEK4Qus6e0UZOQbZtiaXU6ODoDl+esgrlYyykspsrJIlJggyqHOlxAMknMzIcsyBr7XQMiuDzg7a
91cL7hlCmkSBc4NmQcRWJ5jbd6yZGvM/ItxxVbYd8LMhqdIuF8CL0GLesy06Xz2ZLUOVCNT8vZLb
GXWLDKSkJNBGauUjHXWZCc3QPCUwAmm7NzTZjRLIet8kv1p8aL+Ixd5BDbblcm5TNeTBPbwmgCq/
Td0VDU3vB5wrAV6EEWOdQ7jBCTiFTDO0hh4hjf2HYj00DTFaniYvb43yC4RihTA4GgYR9H1xm+u8
dnyLNrWml4pZwm5T3srEwEES2m1fhjGQDjGmhx0uGQVAKbj6Ff5WRbz8zQX/yVrA94+GwLtmgmKp
bsOBfLTWDcdRt6EVNGyyCz5f5PWhxR4Jd2jhH98PIhS+ey2Qs95ANbAWUqXjug8cKvHxk74NAQps
j1NxVBbAIMoFbt7vD/MdFrnm7KrVksDxRPGk1AmUehOvHj4GT4n23jTWLE5hao8r0nGNVRm1eqFQ
oewpKkIPepQBYAYR2yrPSlVXtQGSNJDqxWN+oOCwxojEBDRyn7s9FmQ0EoPsoCCyuCuy1konQNDC
XvtUsvNyGbmKFAJIV1FIIxoHYjNMOcVI+PsTiSEQVbwh8MzmJjR5o+4R/HfcbC/yPv3fabIqq4ca
5IlAtjz/biyjuk8MffGw4Lplyxft13dIbNsGlMsiljrIFof9F5Z+/h2jD5BB/U/RpKhLTCG7nnCk
XSY0dwcUaQjye/eHj+fA53++569J35hbpG0wzEK4xvNw1moiTHxOElAHpbro5D0tKDHqzou8hu6U
+RUHKDWMkk+gOCuEnVT/p01Bibt3eLIvu3pk18cFoHvj996DymVWky4uJZzdE78OVf4nQhVLWrei
cCBzHE8XE/4rKuLcXCYdHefq91cJRgzZ8IHm7Kz16LLkUb8ftM5V/F+Xm86k55NJInPBMc306bw/
GFwC4+IzmDxx8LrPA9gV2TcFzQNHZs2ggLgLvP12ywCqe9KNS1qfRj3OeIt/A4p4Msxhf5wYntRl
ZCvSNtZWyEnYENvP+RZa4D32KL+CvTR+Cil1sHkW4vNEztZLippK9KdPkzKxX/AYsFe50MnOeaTE
1QLmvNdQbguw5shE+yfVZCmpHwVpAWU5qwDIv1oqoqrNhCyS6IHP5+OS83rJm9fz9qn18oVEgLsK
T3mAzaZ/JONdiuLu/CUHG8XE2BfxW309RoK958m96Abv87HSEAa78o4p8TP3cExAxKua18nQdlkq
YnLepiomOs6ibi8zNR6bDlqRiZ7HSb/h90Xjv86A/bbfhUWKHbUlG4Y/iG74wFoOvwli/4+OYGr1
8hQrVDw2wrvwSaOEKVNJNxz2p3n2NyZ0V1h5cFbrxOYKAHQYJ6fBFxiNO0pvIplsEHo+dArq09jk
HrdN3xeo5w6Xk1mb3X2Yy05hbStzdrHuHQHsUoSVA6qbuZwmLjnilWQC40PD21qYydiI1ONLdNwO
YgshvGNrdCyqH7s/9t7gsK/yRn5ywtLPdq9S4eLqS2gnvV2CyzdgScVtrSMjbq8Q314UO+wvrySb
VMCSTucVxwiAtEPlkpzLCmdCvMBif6fuVN8n/RL0kP8yPQrmdycnQLnD2yQI/rQP2WbQW4hdjsEn
/OTimvDjKwUQPji4EfyIwG4wo31437t0BjNHNZZDDlJneBefUr8yfpyVo26uUMIAq6TaSvaZM3Sz
tq7/n54HUZUC4NsDXRC0fbC1VZZjxxK8LQ+vgTShu3/91nr8s8AKvRQFGgndwkGAvonqJsreoyPu
hZmGBO74xgsYUD+6W17YHTWGadt9Q+AeX9e6/reDa1JBuozmkBV9UKHvEgudsHqnM6ZJGfmn9tor
8fAWeYctbwwPCx0nhcTJqoETVRFSJFgG74KjstHXlMk5LoiHF8MNfQhdLiqvSjtez8xciV0+N7y1
v8gomZJpb8WIt65Y8Gf0+h3Zy8RDO4SIiDyq9h1pbSh4B0V+DNTWOzS1XR4AC5kII3p0iOQ9sJVG
GAnwCY6bxj5JcTWu1GsOxXWFH9wX1AwlXpPjtMxwHrd2PwAWXAW7CODMJsGvqmBqNilfCk3TmZmd
e2AbZJSgxBGjBXrif6IktCTAcB238m1jZJ64xCv3ybATQ1BMaqI3EHR0aSKF17HQW3FphmkS66r4
AGILK8b+CgtEJVlDz56Bu6Ei/j488U16fwOyraG1N42R5xMDzE2+gH9tHUBdpUX5Dqo/woxqelq0
8xDNfIZyG2NyCBruaMsTgiWtKzPrdR9y8GBq4+y5dTGMEcRSTSVsoXhGqYZ9YouJsGknN+2E3NBN
6d8ZASGL60CCuaXjGpG1kS72ij3I99rBiWIbITEw0s3qz12oxj6ShVEOzFK/7f0jV0lbShhwCB15
j3WAhkPvYvRBmIZpPNozlz2mPpLUgNdohF3XP/pYrHln1Ekffb8rQh51pXFLbVupu4Ef5/Z0qIh1
A3sFt36a0LYO7jfGIUSTbs8EcMJRpzg9zIdxSqHa1McwH+owicurMBODID2wEeNPr90an1nYqlOc
M8VKwh8bJUt8IYGgahO0p15RY587lBwsXDkK5kI9dt2k9hcKH+F7WhRPOf0rvjSBq7EfvBmyk3ed
m8MiM2TV+4TnOUUf71/Gn8T6AN/6e5WaH+/5JiMN1Neg7+H1G5Tw/CjVAHHT4YSHS3xJl8mvt9Hz
B4TGUTd7oIEw6kW1Bk4WNUS7+etRHfumO5R3vvFHDT2hB9IDBhpi9HN9/14Uh9fzMfSwvttGd+Ve
SqfF7hMbjMKBVS6gi7+P4qDJeFjQJEV1WTcp0NNPkBkCSIryhjjWUnL41P6QcPNW++7vcVxcDauA
21CPVTvrELpOKKaSuO57LsVhhu2cBSpH11jlEHqMqpwNLJQQGs5oyjqneUhcsL/CENdmFZsrREDX
3dRSeA5BK4rBYLWIYMZX441QCrLflTU+ZwUUyAhgPekyaQbA7sfL6hbd4AHrMKKBVP8UsXUx+SGv
npGIFC0cudbIkQAhSzJXuqNkc0MrLSo4REtf9qxMxweEQuL+sIGy5w8FTdg9KjBGl2P3ivHB/Sg4
UUTJqDmZQx+KdZGfbq7ajoz/okA9Hy/bPQL57D6mURUBau7UKPT66j0hx676s/9OmiXvgHTkhyeE
L8FeZTCyhRLnudMEDOH1PHqOWZ/aX7F4L2KDuBHbHpTUJGODzDVIvfoBC2fXlcDWi58tM0ItSvmx
+oh1R6LsuOjqO1K32HeqAmNYEvsf7iNJWFlKjgloHPW8j2/JoMDqBXqGaDQQgVtE9t+Ikw0YwKWa
rfJARgkAcXEIp91JhuLm+ApD1JwyvNni24hCYzi4QF9rM7SbEpTtuCJl2rkf4otdTSFIZyf8TB3t
XbVrzmrxuHdG4poMg3yWESQ/+0yZRV+CbOzwIsZGMr4q2NsQkJrPbHKeDknO6uiQUu+D2j6ayg+m
8ppp/kHoClU5Ngdq5gH8xyE2czU7MYkaL0Aqak60gCD4noUUbs3vzPofe5C93TfKJ/D4gTExS0AW
3ief38FIHlOzY9lVsXiWQ87ets19SH0Ekqs4wQXEbSOD8L0GVBPfz51oh6ZmWFltedkUPD6YtSsX
pcDYUG9OkH8yuyOtQUPxQNXkhn+2cBVqP/CA2WFcqhzxcaBZNiYN+wM71+XEO43i2se9TL+03cm6
/lXiyvIdSiJQqt1jApOLxnon+SrMLfAJ68dzIMWCDzYsc3+GnwYVd+D2lI256gyAjw/AdoEf5h6z
hYwh60UFqJRmrBBqTDmrIc2YVH2buocWsR2JNC4SlxezZzG2LfYCibQQ2LHJ8nKAQ6AmTADebV2m
h6lDmxyuz+o7wVnrb4zvaAofCEH9win4VwcgqwS8sFJx9+egekuHPEHZUsnTcPL4BKr0cHYvj15A
dlu3pDiwb8Ib83qVYklbiR0PP+2ndQo4wAL2iJZoZlIfw2YwKMff3ix2A6+jfN9L/4wXdRt2NP8h
yy4+lYsIxgqP46OZPDSIIOqR/e9LgyCQnPiVd2t0w6Cp+JavO/8S4CL2kypEtNdUYt6w19r+PBTq
2B2ktjk8j3Xu9/THZoo47DP+/nU7AQfPdcdDxG+bPq7HQqBAdpnJsvt6EBJWr6GD9PR+0zOB9Wcr
df70AIV6AWu1VdpwAl8yo43omCk3MFyJSgdcCBs/aHWt3wq5nLjowZHw3mtlI+DJ15OZ8tTNCRGn
rUtd24OproXDrDKXGhjgJEHPTd9aholrscw8Q86McElUbOaL/fdbp4ajl9NBVLGwGVqd4zVfHK/+
tf9Zj89s8mmPWcebSVwBuBxfHGqjlyXbMtOMKT5GTxh2PygaSXJGcmpHOXmolgAobAxNl60M2AwN
wDCE3+PUF3/4BkO0onTuNyWVPU3G5ULon9ZHqUygoJiG9FDZZp2ifYhPCjMMww6K8hGYuySxg27T
FeONcdvz1BILcVBkrrm5XNp1G02S2aIKpCCMCx/MyDEPqdfPYItIF8ud0KTmy69H0dBEncBR5OcU
boBamPTmdKjQlSHJ79+YQ5i/4Xs7wnzet/u0zeDwUI6sE6MF2Hfgfemg3mDqhlqZyEvhw9xP0mcu
sKkkuvNbuvn+hQ+ohOA9wJdk0pwUdPPNWfjXTg/BQdIgNs/q9Cq8PZiq4G6bPgoDK9tIgh3VFKbB
TQGvoitG5krdXYm47FUDKVKxWQGbL0VYRUoI83QgzG404srDEfVfFRQ+5YkPIn7t5AhWxaC342ss
36gIpsBMCNuqck2I3IjR9l10U03DW4yBadKd+0Q/KCrJ7Vh3bcSlt1X/VWCU8DVsrnHWfS3e+HK2
En2Y9HlZ57Iprxc7xN6bztJRGTl+UqYBK/Mwc9NPGFL6s8p/NS/xCNhznHGrjtwfeuDlC76R9h9Y
TDXb164tvcGzlWjdgcHiNr+l8EeaZCfOkxKWSe0LwxnFr020gCOTqwdo/KUON+wRALwg1NX8M3Dg
cXAufnMa9d6oEUkn7BUeWyO8qWbrSNj6nJqex67rLj+5S61QPgpXLOgsTRc3k/mX8wbNmRTtTLUg
rZf51thkRKCCxKMpmsISoKKfDWjYXB/wkc9FFJWCdHk5PzzZIhLfziPBzaYemsSsUl7Tt0bZce64
DM9Yzd7CfsTqYxlTIlU5cJCjD36wL/LRMi+K7xc5KLwJgvlYOb/q2ZK2WYJKd/AN/qvdD6rnclDu
cXTlZfDtD7LDHCtnqMX1zDqGRvs4lzvHQ3GvJZ0jHE+fbwcyreGPSC2LnDYUWDkcUEwcK/PpTmOE
qX9PGSsFrqpIs90nLdAuqnxjUvSyBbF8NKGgtgkiXM5ecVIia6ssq0MPuyInGi0BmLPEQsSbDcpL
z7MfzRcVDTrvZtCBLpvBIbX5wmMECKX/FMn1iWYH6tWuZmYcA0zomy105y5IEASgnLSBSj15jnal
lucxMsxKONFe39Wc8BOtHoXX8JepTuLzEw7ORH7JVLC2BbFDRYQnTjwO0MHo72RdDpZ7JZwnZAfj
CqLxU5LvnuBYluzhrh8hohU21Td5TYTAmjqNqKv/CanraVBVbCn5v7R8t3ISPin4Y5x6w1vwmqsn
Nxn0clWore3mLeCjItKcgszec7wuOnQxGRYnffVt7ehwnSL5Xryto/MwySH20hByT5aS78+GBnd1
pmIcnhnm/oS+M/qJh+BfwsKbqJ6ODCWHAwMkp3KVIRX1nq5DNlcp3JCy8gj6Nl9X0V/Cz7Vqt4rl
NsBL8laEju4uWph+QC2ew7/X4ET3z6g0gaT/9qZAPYj92J/pYHS21lqktCQq2GzYYUcVE5+U0l6m
7KNmgpeyPGvSodY8QuGc7yrEyquGXBfERMe84XcPELSpZhLNJ/qFDkX2x0C5UmIIzeQEx/irs2jg
b+AuPG0NskYN8+1jaxov5oXPOz++5P5+9IYqvW0nt/f9ZECFAt/hjmhQdyv18RMldgNM70bb/9oX
uZjprRKizeUTeN3Rc5Mck2ns2HzxUt+ZGpqbGL7YHcNfwblwPKxJyB/vrxWn7z2Mts2VUlhXP5Vk
1QIHCSciqryM79kLGlM7JQ+h4CwDbCBh4hbnXh1Rmpgjn3gxu8iqluaWbl93E0OtArofzaMtAjot
0lvoe85NZYT4rR9la9mbTwZWXWXD/5utRSsTHPiBsHZ889AFVYABxBEMqGf68BRYq75IrJ+40Eou
OhK7ZZ+MvYA3ZglYtB6RhPJZcpQoxn++g3LN7uO2EqcedadPpCGJhs6ZZ5vDJpDZZlrm/H9ydfna
VuLoSscdNa4xIuA2c2NjZalljEsIoxLCj8+o1SPgiXE4x1VQ++zcKpU8reLSfadtWtnTAl842olJ
0vUdnUSpTuXXxFFQUSNZ+BrUWKYhdz86E8FjR2IzCxxKKo0Jlyhs4kuepGvKCKabqKOfqvOeTz4T
O98N2SnxioAyA+m8Nv3OmexBmswgvZgnv0hkUj4q3hs+Y48lgKonU2EKALwPd167nCu+s5yQqyWW
EKiCOnfZdwcXpxBgTaKdPljHn1ypKfFBzzs1L825qXihRrd6ityJuATITA30DRjOwltapOe3KK0I
ZO9mDqTu6+Yb0HrIFBkzSSTA9uew2F+dMsLceaN73P7FJEF093lhrdGbSUrYfYuMU9s/soypD/dj
fzRgCKC9eSmcEEW7eBRQ62rk+olmqywuCS7O5vsQjtRNVvrkhdugZpNCaHHIR5SQgzrqV6u56fdM
JZg2m9GdGdnegrF+Hf00X87Bw7fmPzqwXh4Ld3HENwXlls7Wax++57FrKkNAs1wU4KMF1IiRdE/1
PSk5ZPeKldfPIIqT1wxgHNdrnDDdVGa6wUE1F0P6a1PfYz3Re4SS9h5cH6XGEmh6xQfbO9XKNdnJ
mOyZUSeY1Hx19AACuPZsOWMP1ygnDiDRuukJ03GWuFC8h9DM/Cdzk/n0qR05Rm+KJ2kAS74VgZf1
4LbUNkgqFYhSBExZwi6UnKh+Yi9dAHCZV+5B3+sQNOWFBtIR2l7xeLf9w9bDpmWLqbzHRBKb3uT5
4fvPwV0wBa9R7pXwsmZv89Jal18ZPmvGgwwUqwXNDbdzCz1A1jEGRjaJNATACpDFX1SMpPgnDRZM
FoBI6m+arOgyApHWH6ZvsnAdhFK9oMVlIr6OXitN/KfKxkiLPx4As8Y5f/yA6zlOQGV1Ph/viwaD
N5q0G2ves1sQZpZc+2g/FSvQXFfj8hp2GovU9ifAafMhBiBNCV7aMT+cRF0gXWW+nBP5MGQDHV+K
lBlMymHpqYO9h8cepMFvsGAVb65/t7aSO2s/+wzRlNil60133Wr+PDdcGVQ0oOhggiMHN18Ln5Ex
GxclSHLnvntjd7JVsGMoGryCNnjgUvLnKVYyQE/5o37fJnyvY9TqGgnYOtBR+tqplKhrl7Z5mSDD
lF7JupqHFVarWFqDx3XnlAHKScpvrnX4WfwWSf2UU2AsYw/YJqI95QMmcyz4uW1FhTCdv40e5spB
iejF9sMCNoxT17MfWwgA74InMNkL5io5QCLewzIFeZf5RldGAeftKX+XnoDjS8hPx3Bzs6XmypnC
iyFCxDZQDaZVzc/GucUmwFWSHXIZE108NClhKmOLNYhL6r2UBSV4ZXDtvFW/JghF7qyYLih0/Dhs
g6udusj3AFP5G9SkK8bmB9Ia7+oEb7dGxGWFEkB/x1NbSm2DSOP4sXQNmydSv5ZWzbM7jttPoqHR
mTfVW8Eu8utvBQnuXrlRcy4cuiNz3giQSpN+mM3iGJb6OKhBYi16XWoRtlKQoRDpaYvrAZMbuXkZ
+xn1Iylwlup8Z9LLV1iAoUv9dCcK3qJsQe+IAw4FuvppsXzt87gxk3BavrOVVEs4cAsxvuojSE0N
DB2wHbO3TXHioSSA5TM7zh+opUhpbe1WTy9neorurHbnLKRknq3AarOL1OGS8U/9Va6dxPQic1f4
31zqk8mbze7ykoAwvuO5XB+MLKPEsdf+5s/IT/QDwbm/iXcXqEozZHSJWC/6nggGFxzrzSBZVMmO
G8V92DgzNbxeSQNCiaYmayxD4HJNdTNIIehBN4OjBy/LQGKvVe1HQf4yZQKPDsInknCCQ1CsLEMO
FCdCh7sUh5OD4CvP9B3dEFkYX7hmsAwarSi1gQmOEDg+xxlnLZmG3FAugnHzrOtvZRYewwobPdpE
0BrW1YuUs7oXyHswfj/qDiTHwwcYp8fkIngMS1Z6nhjSKf95hASLP/NwYCjeJIlgGvZ5za6BqBV2
SrRcpJc/mQh0Dw0AJr4++ys6v04Xdi6jHz3po1Nqe+j+wGkuEEvUMnXx4BcwQxeBO4aO637fvkxb
kJEWq+Tb+ecg0wn391hagAnxCNr5Hj99qt6F2jrnaJR/hJ2hRHXcfcNiRAvNFcuUWL0Wni4k4ZjW
+4Z6NrSdS1HIXpqNqpo10fCDKhW75s4xHP/mZu3QL8SJb8oYtmvmEd5uy8fsVI7oBkno/fp0cHID
+4EwDQisKG8dZe0nFsSbQKrt2kGZWjkPjR1spItT1Zqb8acUgSbfi0F4x4BkGpsIR4/y1mqMJBpP
f8cerLg1UuvlzLmeItmf7UpsjxhXem9jZ2YXquTkJkJIQUFgsv/E5nn2er6v354Ij7Loe6WJSMLL
kh5aZgZVyGNYQorBsUdYxH9+i64YOEBaKtWiwP6Qhb1Eex+BA/CgGJff7KadU14RX8RjKWbtznYw
xDpjY931szZGM2lnicRJ8P043Kdc4n+W5fI05i7ZXs9aNtrdxQ4jqsCfR2HIAeZ7sNw+6Vst6xbF
dKVbMoRa1KDEavDbpT7D+tYIhuJzGsd4i11fi1DK82Ste1UvBov6HlQmifRTJ7gAuKYTCqTas9Xy
RAJRfY5XdxpIQszCBuoh9o1lii0+gspQ7nPgVEfnJZU0Zn+TiqtknUpUsiHhltJ/iPeZAeR9GZbw
jHrOvUD62jdSQ7D6ejJyK2OB+z4LtjWpj/lsXE5KfAgmeTlZmtKV7cP6O1Vzo1tf+xxTUYvbs9Sq
/YyN4FJNhyN34wigjcEOVKnYuu4rXvFRe4ggpcBIoA8YxV8Szhto61L0L5HKXazgewUn4uWgMQLE
7hfvbRI6c+AiKXsnuJ1G+vEbgCZ/+LcJNPb4GjWT05V15OKOtgWzUjpXbvazn96sJRHUQBv++6ds
8gagN3c1m6ZpoRs2xsEzYWVTwuIq1zFu+7NFuTQ987VzCIs9Fkz0G/9E+kxu67Vn1jsIC+SYb6ud
ZDhs4u0CUxQexaPNcqKM8Qg8oS1fqZlns9KMc72v8fFk7M2wWjiY3wMrVeHN8b218efvRgn0kgI2
XJach6LSvr7C/J7qv+hbWdaQH9Pz6fFYCfRCV7FUf9yXA3PYYm+zFJD4auMlx4l8qkL8IcVI9x6U
RT2IYhEUDxDonU4AMNY0koH+1E22AO0ksUkeKKns3txuZKaJ/07nrjVa1rNkvzuKHe/OXPu8w8ms
YT4XLLJt34VJ470TJlrxzI6LeDcoqyZKZiZMAmmNsn71mLhma8cKnj4jLkW1prZTipadc51BPKM+
lAxYFNIO+LiAncE3IQcqexfyoGU6vTgPD6VyKC5PVDn+Oq0/QNY1jDNzViCmcrOjUybEoW/ZQOgp
cHXbJM0aJRGDPCKlNiVYAYe5DtpMoqxVi/1114i0UNrgWog8J3MjPwpFMpSWYZOUw1ui0s68uRt5
cLcdmtcPhmgWhB6+5B1Bjc1Q4rg9avZH6nRbpkDoEoyBDr+fQV+XCRI2jpPFrukXtB8udW4x3kOS
MgBvsp7LRPKUgcV0sSnSxSyo6HOmctjLMvPoP3jafU/AgE488pVISHwPIhqV2NdyigSS8w1q6UBn
MwCR/q5iFI5T1S2xG6ZpdwB3WgNX+V7PECYaXRnsB+ZlD5kCInuxt/LXktm5in22dEW6HrpSUK+R
9TnLlfSFxPUK+F2+4Oxb3y2YunE2UyZTSHXayJVQ0qb9s14Oo3IYs3aKAuzzCZImYoAuEv6ZHqeX
0xFp+rU3Kb9JNZai9SrQSNGRZuQpOK/2q+FRq+yONE9A5DPKwh5C2KXDaLlLqGZblEUTsFzPDlvU
iTcPlz+0o0TtaveFoUbM2IynBNxzYfbuVDG/sMcK4lDbZSZ+USHWmCVqDabVF1MYI7yrm6jbABMB
sL74rlIAmbTahivItVNjI0H9wA1d9XeClILYJH1SznCfu11qYurEQyUv7+MkbxW9sIlHo1nsNRSo
Qfw55ELOdjw3I2lRQz5M7U/ybmzpx6Ss3rO7o8RabtGGTSZa/tXyJyTsh1PkF1HnuS+Sll3hBLse
rtbhwfTF0jPeOxkRXSjxD7uRdnGjYpUPv0bhu3/9gRQ/bOf4+R+W43e5rrcoajKdQu8wmFk1CaSH
K+6AZYSkv6d5BLNcQvzPblEs8o0r0DY3HoZ/+N6EBRd02CA22z1LtV7pZZ+H571tELVDHEKqmrLJ
KPpkq3cNGf7NY+n+SFVQspYW22miDzUBgXsCwkB72y/qMaOgWftukVGnpCR6D+z70GhqG7rs/svY
RxdaOygQO+Yh8FEa7/MZu1MAmKJJiQhot4vfZU4aSHeE4rt5XjVua/PWhDgqQiUxcFmkVQC63IKD
l9i3ppelBz/yxbjlyqj1aPWxhZ/kyvNGBP1eYhQa4ksM0gt7lQlTwMztG29S2jPIfqFopl9/epQq
VS/eB4RS+YJmNftc1mT+YIEmt1i1K+S7IggD7d39+60nX2pnnp+3t/S9stFIsOZe7cbn2kr3HB1I
CxZ4nh650FKBVuG9f+L5E2f6J5KTG+Th4OoL0/tGhlcrDGlLvlv6lr//6Yj0Kt2JmgMYJ2e8mi/P
nYtd02MAuqaSuXJ494oby3PAIxEDbb7ugjKExa1Zy2A2hKJIc2/l73rxdUkemWTq+WWivrVLLQuX
B3RQ13Z+JnSl7nuZMTqy1Gg8m33U/Zj/Zglv5tgJK/IPu8t2wpWOW0g5ogsOLyleMjkfGffFJaeE
IM6fX7HV0gX5NxSowH4VKjZ/dESpbhHhylnVYQDvkLgn2s50K7Y0XtVh1nQZudeLmrPCFsVLcVVC
lCCnJIT8T3WFqGBd6YtvGCN5AE3U8bo+6ycfdQN0J65y/KtgwROoz9Ao4ilaThovHE+oXobjx+g6
KgZY9dH5X5XsnY7/2gVYyq1V2n5QQ+2x42u1+8fWS5GE4EicjvSomiD1OpJStHFF0oBDk7nMGAUx
alIRP14PPYNqA124NAA4NPNtvWc/uq9jZ0D2hGMZqsNyfY/9aht87tSe3H1+g7g1pbrb7dCZNBNT
KY7uHmzV9lxp3qPNO+Y5ZsOt3rYa5SGfGL2hMKuwEppgYB9iHiKYno7GisqR2jAL9oIGWh0kTu0M
WWYvaN3vtKn7wn6TX9T9Aq0ja9KQ5QzIUvrqD7ume0RJJikrsLxh/j7kF74J5hkvaIVp4CMKfIDM
jFk3vk11bbNUaDfWk5z0LKSftJzJl3Fw8wwdV7RhyktvGJcWRdN5cp0mK/6ENF+0vVDyJyyZfXEm
HJNQIZpbmY10ruqN/MpAJGUBHmuYK6l/yUoK+Nf/AYtkzRUpvLLuHG6QatjP6wGDP+oUFJWRYZO3
AYouSZhyMqdCoRdU/IhXoyGXuLl/Bx2hrromy1QN4uw8TLkgIt7fFSwsonaNtBCpmQ3T1r1VaJts
vzdHsz3ou5WZydKWeLr4nSfFYXr5wdk+qk4bpzapjyulWhN4nuJT1iefROqWIknORZFxzcPgXUOc
f3tAobmaxrDPKHWaf2C16L05FuCbC/I4J5JhpXfl0a1Z9fukRXlZay6aBqC3yADXZ4TQxXBdGo9O
+y78+AA8N7/HtLqVnMUg1u1p6dx9Cry9IBE/v1iJiLCf+FCmpt3I36NSveEVSizNr0bfY0ZOb0Kw
QsrFjoUMdm1l/t7OLF9Gj/6PQKPXDkgI+mLZHZ9R26iJ7YmQhFQb7HIqj8Yamna5SF5FBpa0wb+3
2FLiOJDCYzdY+gcw99ygyM2iYcxlaiUK5FqWO63DC5U229G6bMj+2RgC8mYs/zs78APNKkD/18Lo
bRaK0vJO/fKYvXCYoUU6soxpb64sLXxP+VUv2hZW+TeLWc0+hRR25xHbpt4KXalQ1bAvDn6ITEHn
yyrn1c/TAYiW7e3oA9rBMiMuMhWLFJeLMv2LWX+3t//Bo3tbfgLUY9JH9PgSLH8Nm2k0U6TW+ILL
WtHZM0wkhbZZyxdOogBjrFPj+JNv3yBOnuUUq+cUakorqAO9fxk2ha1PDKWA1esbcxY74IEQVMZH
uIf9EIv/jrQl9Z9n9GTTrRcSOiwKf4EdRXKT9j88dBTslNejs9BEB7jqqOyFMdRSV6FrdVIs4XSu
XxUGmbvUwBdJnsHv2Ykv4aOm/eVZ0jv5NQha/VX1K1lL1Hez8ASNPnOveNFOzUIJ6RutTjxyr9Ay
SdH9cyL7IQNvypQQHYbnNHU+XiYYDErzJEXtDbPxlZ/9sMF1eNubG9Wl6zLjbrh5iQKdx+naMWLn
+6tplCCawAGqMT320AZtBQSYQvAqV57lzYqtoWeZiWH7RtttuSRt10yFAOXNGkTtDE/yYkN2ShQb
rc2dtpwZwngP535LnU+TEK9U/ekofLqcv2abOcf9Qco4cJMUttOds8f8WskFEqO9/xmBSOGNk2Bc
/LQgoUxgKG7jBnJ3cfIiQDzbTO8a7CDrAdN0by4Kw5U6jO4YgtkpRhc/jmDnH4fYxDMAj2azyTjn
w0hjQQS+K1czdq+6r2EvQiy+O2RNluMSXZKBNiqywou7JwcVuLRTbnqEkPU1K6CnRGYvWcMv4fi4
McUQZVoEL8MLXZBmozDtj5zDEY1tOAz7fy3WUyZPIuWpcCq8adnuU470IWzV3bca3ECqVgg84Pw9
fzOGSY2DyMP6MIqf+BvmLMMZTkGXV7R4Y0YK0jk0Y/SJid38Z+A0kqMwA6Yobo4hGEOVMZm5PsH9
zZSxDDlw+OmEZ3YdSWxSgwVf66jlIusULFNNKJA/QW0cBm1gyTNCN95UnfLZR5xFvvnQ0hD/tLh5
JQzZW7yxGapCDgnEYpbEoN5flmqo1uL8BFRldOT3uUSoRtoETe6aGoeUteAwW+Ni7pqEpo+IKRx8
NsA+q+8JZ4GaFyr3LSHr1DotY0o7odUYwVJtgFg7if4VInrLJRYk16gA+9GyU0Jmki43+0zKFVFg
eI5DIm1/8EGd7o5REHb6AjRGP6AsD+IZedA63wFOdYfCFXxaefm2HsyoRSs5vulNkmUiZnq3KvKJ
AZCDpHYwdWofn3fa67m0WW5DKQimuQM2OGpGSqokGA34U+5/xgNh7fMURXtev+Zu0knwwkh8dWVd
7JsDHo0i0NKuXbQmYkBB28FTpEEkPLAdswiIsilvK/rIo98iF13iHSt+T3ya9YpgG2v8+kjoyj4R
uDnsOo3A94282O53QgwaqI955YL5vfhSSXqgL8d+Kw6pxNH+Y0MriTRr6vSIel8lzv+Zs8pFmCv0
5Ay35ccsdCQnhZukEbSUUrlULMOEa4BKArEqbHhGM8B/7G6OisSU+BK2eRw59enntLCN6lo2hIiW
tQzUn6mZBkgRWJHTBXEpDvQtWnHSVlDMzZ6S4sUPVep1PYR3ZYK0lgqWRUYwWO92M868fCC6Tu7z
z5auVDLFvv0Y1pyPIFwds6YyrWUknWlf4nQ0RzzbTGGgmBwq0pG4HEXqcpRWyqapMN9EVHp8eqQP
zLgUpH113OwOft1WDHDDmdg/AoQIHxtC6lfZWranQUJH+1AV+hwpW+1uDhoaEpVH1mf6JiWcGsKi
PXxD5Mnq2ph2A3MtJpNb99Gwg3i210srql+LkLjFntONSL7JbeE8zl7mR/OrHbgVUHNimcoRFQi3
KfjO4SKE2ENN0hzERtXN9X0e3MiuKQylGYX73Al7JdiIcnseRt+4AYAMswwk9GhXnMM9OLWnf1+F
dNPpKhK7QyvL+0hzSBlsND4ROF8H92xCtaZ5QyKziEVAgjeLWEscMduXwz9+mjkUsT/BhLEvcpY1
q/1l7Yr8R+tgXERwqM/EG6btIorEKtvFNvBlk0m9unza2UfPypSeZ6RYm0WK0u/AueYNpcXlnawe
5Q3V5djPyVUazgV4Dfq0kkyL1nI17LgHf53JCnJmo3MSUZiqSx2cNUsIrHElMShlxCoeLABZTvlK
kP4qtrScdVV3OSb/DW4GLckuCQ6oovbU7VELR0q+cQqrK4QxFg2VfTfy3jpfYD9x/8ZhdNoMR9mH
rowCQWfTWtICjXr8jq2WiISpT4VGyx3mQZovwu5Eq2BpbpDdTmmT3rqHJbLaXXcJDQfbiVnVn2Ue
M4ehwDE538kQ4glZOeDCUjNKtLnPI8fVd3wgiMd1G788WdBj+YvsLd0ck+DJmmLt8FVUFEXQiMQk
Ipb+dMYnp3tQBrpB/C+D2mUqdh0InjUHn7gI0KqClAc34QA7kQXoixQ5gQ+9VsG2JjBxkdcp4fTy
uUhO/xJjeKXe9TVhb4O7mSVPfvkUqQxwhUN5fYEvU7td2IR7blW9Uo5zPBzkL7q0sneFoVxwIqfB
9bBOb9yOb4vvsKfKJDO1w12C34xSVq7rGWtmMrNgPmopQwg0dA7jys6o4LIlv8PIiWw1/PZgFdjU
lsMPv3Dr00bYe6oPx9WiRr+jKQaEruYcEm9XfP7DhdmO92TTJeoxbvxXeCyTxoiyFdYcLDL7mCIS
tT0LMXMVcET0mlwhw0hnix9nIQnIu0a97kvzn/65m3oki6zEIP37wdcfk77Bc8nnUySdDt0sEVyP
7gwO+o2OcQM+Eas9++7B3drcAnEEh6Ixr71nOkidHBtXVVqzzK1EvaEOzil1p89NzwTizSqhiARk
/Cs6Q3vnn5pPBJYgANRJnvib7AGrB33+yKnh6sGnQjoYBzm9S/oLfc4qE5t9DqpjnBRoRwQwl0s9
fFrAvMWxZGezUFjDoan9lOBAghgpJ2AFBBjViUhaX03+yitVu1QEqtnM0A55hVYYabHIjIxpxJ93
p5EITCK2Buo1TBibrvPKvi8V43OuA2BU0HSQc7KvMw1zoknk3ZERM2u36K1/970ZqmCTrpInUx5Y
NxbZyWSly/HTqJ8YUM2/OHDYQROQIib5MezeR+Rx9cm0132iT7gcfMFAMam8MRVPeGpxE0flKqzR
BmlCQeraVneozpeBcxDGua2PF4SiUbqHpssKYD2lZPHKQ93vvh1L08oCKUtUMZzQ0MqFBvbuu64R
p8JM207Lezr2s399h+iH6Op3WuxKh6oEBuIxdjvZBPN9DrBlS2uYoNH7UNJuEf1f2Q9hoaTGaN7l
qqfHsTZAG5A0icHPfH38kyw/N3Whly4ZxJaTAms79O6rBjuvXYMaLRkcMF2jTy4ObjF50RxjwNN8
mE1eamRpxDu1K2KjiV+rHOsB8zAkjPjeYRGLxXZkH6Hdj+/T3cqvqoXoda4rG1/tCcdLX8AG1y9M
d2RLyMZH/ClnmkV2+Oe2k13HvJPw8rJ19v/kgL6F9eeuuOy+67CNnKNvnC9vkWSNmM+Sz6sSl0B8
FidiRkLp81SOStxy6ESpm+GfaWHMppLyR19BltKybImW2BBoVZc5Wn8cr5WR6iAWK6cIu++HMf9H
nd49ujh28FB4ffhzWRg64Jjwwwr/E9sL7t762fF3Fr1BawaP0V/MYSbe01mVvHnjsleE5YpNYVE3
KudBKsokxYUZk1rCg1lgrW1meLyMSNhnIUaURi7ahCN/ncg6JgC7h8cawwIny5/X9S3KSVq3qAlH
kRQH1DGM48qTVl5s2ZruMutK4krs3vdsxxbU41R1nIrYZzZZT7mLpYbWJQgkArb6AVD0iO0nM/yt
OuITQfiI/bHyO5P0YQyynHb5SAGTR5NeFMNYySYS5VjI/2HCnlT/Ik9GNfPlFQjyEpYaFH1saFYc
KWiIi9fYMlk5IccwBTJFfltVrfLGt/VfAT799u+bfCSQBRgaZaxbatqrCAoE7/H0/2hgQB+RJbHW
btXKNjkkJ6CWXC4e7Y/X/n7MCDoftZhr/YtT/1fZiIZtPF7GiWdXzPmQmOHEiVwGIf540XACq8Ec
D3HcqPk+Gh/Y1BwnvhnaFu72gl0T0JwTPF/t+vSIlw3IRDGCXMKadza3Xa9Z8NdEwM7K7aNzWu+M
gLR+BIoZURJDYaK65VWed8qG5mZmHsPyJfkbbWX4AufBluzTcofYitjgrgqkvlFiKlUFGex9PZN3
dr890ylSIdjbz9PY6Fj2RSVCbSYNMzYF/RDLgi0JmjlFUCMO6H1g/PXUH8qC4Bu/q+iEOfot/ugx
eIJ4EYSSeRrwmDGcjDobl0y+3Eue7X+YnashNG04hKrSbqlvqhF1EqaSEE9KLIrZ24SBYOxMF5yZ
85BJN48xcnMWj4wUi6Xrb3mQtCHylckIpmZZGHU5XB4aSj2UOqBWliS7n7hqq/bTP19aQtm9hnfJ
jE1MUSaIXAryCQ+YfLyXJVGjMr/C7d40ynpxt6aqKLFYRzOhLI0WFO9EXec/8EA2MVAitpY2OQ5Q
RH0S3h7kbipm84gCpDUZprRThoffexm6okvYx7PsfdCZQE541/kZB3JCxrFBguKxcBo+sVb8vilr
tkNoOcz/999SlDKSKwBToRuuGGTzLxKJ7y9R6PSyT6ukOap/30ytiBd8PDqYzWv489kUuIAohqDG
ll7K7F5z01SzH9W/VAyoZeydj0BU+Xk5NvIvI9ktOAsc+FjhKfcsgHDWlElJauFDBI9AwM11X+oN
2vD05zwDzccy8HKPbvF/IhO1xc8fqOpwtbm9nq5E5ELL3e3exy9N8eALS+qM9/mxQ7ZRd/ozL9lb
iDiB0dRLU3gYqjj4IDXQ81rBHTqUMOZkMc4zO/cuHS1jCbrwjaOq+fOKzVZs7rDLljIu2Pazq7Kq
bfYjKbhrBZ4vtE5c1bh+NXPZ5lL9D1WFFZha69M+w7HIuel/LCNHmXBCRTd1mkscyoXb7kXGbtak
JTP/vr0fTyi/TcZ9WHx+1xwvcCHpoKOj9Mu6zoy0OYlVg1dB5jfjwAR8kJecmZ+NzXVLu9l6qf/3
UPs57VHxW3q8jUc5t5cOqSTwk1UKIu1xHg1UevNkxrMrlOM23b83RVFKrpCHvfcoVfW8NZXykSGK
AZbchOg42YaCTb8u4YW9Y9j8oqIBLyVBdsfLKP+d03vwSQX+hTibg5Y0xgv3MuhJRPkbelkMZ1+d
KxMfJW5vP5fykqUNiYxen2WDLhUx1ohRTjMrZcXY4ojYbfA9/VmiXbP5kn2yb9IRjtAy63mfC0CO
LiAFS3jsn9PBtnRpk8PYg+yx4XSUfnUwXEDmK6YPjkFUbjfA5zHMlCGwsYDcHxS7xZGMcvVjUga9
pEO5FxJeCQ0CyIdiMcLmlu9EplyLFVdttxWc7nqhQSO+jKn7wuLOnFtdb1HPtSGfwV+zItqSgGnP
ApI/unlYSFV87+Iuvrs4e+MN1pfshm0zrUyl614v9ggkiAxS4z+WFw/vH9mCIkoiZO43/+m7l2Dq
avB7yytHUwQkJ3tonECKZV51ubWlokglhjZuCOVQzGk63WTGR3kRMUw/qHL3f5EScUcFHTYH8IAr
jAIAIAbRhA+Q+jch/ILk0Eo7NeOp0+YzJS6m1zeUgDOLIIFEJtacRcK6TMExc4r1sh5Ez4WtZYir
QXSep7hR8Mnku4b22TFP97bM15yeZO391wCeL68zZih9yGwr/D+ju5VM7Lfsi55MT8fzlG+MOUkv
lx73Ck0X9BqKGJXKWoCn4lUazmZNAJg4OmpILldpM8mX3JLwoKWnutava0s0BsCO/ohyJ0OzwEYT
4Cug+g3lxeaa5PkumxcbWqp/H6FkKlaVIUNMvsoI5AnIsFVbFr6HZ5sR8myFdzzxFfVdVErzKxxL
M33BfnwLgxz5/YKD1who2qqkPIMliIrlfoaEqkNW5seUCFK5beeJ7GpqHZk7ff7mQ4+zmwh4kSWf
6W56DoVSUpAw9zhjrlV5xpCMpjgtBUhm22QJqJPDkYN4qoLkVvkc8AdYd2ob+RQcmrdrVk6wxZLC
+QgisjOmwO9xM5r3VGzVn0Kywlv1j5DQGwxsYruRDd8rleY5kZVJ6IaN/r/Iyh9rj8RH4eZB8fYn
+1PVn4C5s0mPfMPg4YzqGZXi2yF8D1TWVEyw4sxzlheMwxMtuOWtw6f6ZgZNIr5NCmIHmf5kOHYP
nPpvn3/JJ50ZRsDOkP9ZvdaD+7IpxT9igi8ohDoUw/JCAGCAgs5Av6d1czfF7Qdzr/sRIAQ+HFsj
Qte/lYYoHpDNIEWoOzlXoNRoN0HY2jxTQxNqoKwEvVG+a0nbFgOzt5Am0GAoYC11RgQvTGcEXrLp
mtjO2Q2dBFyssdtcc5dcx0ngOrHc2Nb4O4T4II9YveGvH5z951GoXpiUKM2lNIehOctcD/dpT3iy
hOxeenZX/cLUUatefIH4R7E7JO05xqvZzBqN+MtDzXMqMl4nFvAbLeU/JlzVeX0ljxr312MXhqCF
6708T8eMA6YVEnTBQVRm4Wmfe3LtvTngf71uZ0i+cCvf98O44rlYCkkb/laPgSq5FvSPxnRRa9IH
ys4NXiIOXt2tfbN/oN4J6HBF9RUaePbiT4BOysxe6MmvXOm1iipjKtpDgG1ZO9BbGWaODvRHJkaD
TD4Cnj5fM2zXUOP0tmBxSrbrbdsM9UAHdWKKsRGnfKPHAiepX5Ig4UQFbvQ+a+Ys5D6QwEajP9ma
7GS9iHagSNR/saWGZiyizKYx1zxWwj/5FHU9TmQMr5zHl4McKcfqW7MAaS3ri37m2K7K6HchF7c7
7vyN5NQyZQXm+7P3fLTSBniTfTGiiFVvaD/TD0GTaUCSNnuq1eoR57MrS+KJ5SAqlBtvkvnMjjN8
mxgu351WecPubUVjeUGcuWE4/nHxNe6+zdSMJcOGJRNV8k1tCs8Df6GQQOYjByySUipu45IOTIFY
q+PLia1SJtHHaJXmjTn7LmAQz6y6W173X6e0HjYZHWOZF+WUkrOzLlF0gnMlFRRgsrpOR/5VNN0w
uZA5/aL4BcAXBcZqvlqoYI1w9pR1afKvVqF1Ppq8TPGnUYXr/BjayBkmnupHxniLVA4a2PfIH2Fd
fSsqvqmZ1Qo2AcWhFGnNXt1iMAKRQCnyNk5bzVwPA28esIrLWoWgf/18EdpkYKwYehJU2PmhXxaX
1ofr5V9InYaIPqMkGlw6lNFxNCcuUC0SwcfB5IaQtaTxevoDuFbx9K4lUcB/te9D6kvToiL7BTID
XPQQqhdijDJnQdhC16NagUO3sUwlbQxEH8RPajEL9xZU/0WZ8bKdDp3bbqd0CUusNeuYEI9dqv+8
5mafII5wvzC2opTUCOfJr7wBlLRY79WZf6Hc02DhmNUcRNJrOeETLgg33P6YRLagZdNaZGU2gtY6
rttRl/p4QUPgWFBncHp8f6UgtZaJcuufnCk6gyhmnVgcpgsP9UpjEzc/kc15ulXcIyqbQjK69CHm
it1YomOex7yK1XGH8cnXJ81ukcGonOO7QmCYykmenUYidGocA7FstJybQBnVxTuYCeXILdFCKxjg
pfT8vq4mlpgQHKZlFwQwCzeK+YoifdAcDjRe36TPs3t9ADdr8qCi2h9YBxu2rMGWZie+uV1EhW2d
/GxfBdFaZMUW44Lnbtns+gtTY601JlZqsx8WL2gaZI1zdyWuq9b959hol0DstJdZ17wQLi7x2hkr
EExNCGXUlkPR0kC5DdBX2bxYmYemxyIDBv0RllvizJt/zPqqhmh51+hTAJ8vyV1udwjHaX7ySqQF
es4od0gy3BEU2XqnuadJQU38JlPPV2DjZh2V3IbxXSQlaIhoRm7dpTBfYVRhddTaPfmGCNYEG93L
3+husEFKtKPee+7yKpGmWWDBiGXTz2pUuLQNtlGL7ubzeXEgEZmZnJhGTfY4ArupIiq0CvFRTx5Y
vylZnVttEzunaRMdZ4GZhUrWCKigoZZeg2+4J+aErBo3FqK8M0Rf0DVLiWqMenZz5GeVB+wSS+FX
S+lqeCMnm/UkWEPoyfx6uTOtQTCunBPLfiuwg2Q23hhU4nEY33c8Tke9OA4lLmPzPmhm/4sCP6/4
BTf7J5AOqwvG1102yJRWqubhRp5/KLECksUn/ccX4aVKob1a8tuLbm1YlBnZTN7B1xkWnefz4YM4
iQE0Fft5yaKVJ1J/dvhttRlk/tGVcXgZ4Nlfo8CuSYokBHITur5lpnD8+YZ0/IUKFZIm89IuEa6t
9H3+e3Ixetmz5Y7C7cqqCB89/5orLVPRqm3TbJ1Fs7IXZrqCBTHQeVD0SD6iwml4RmUI+cc8oK7f
HsRSxWhWBJ7Utv8DylB4LuinwBeZLeunnl9rnqPmtm2C5E0Jd3RE49GYxf1QcMWlyYPchP9GXUFp
sDjAYT43fQvqRsP1MkSWU/zfZfKlGab5+046xL2mLROhK/anw89+g5qxwz0hleJmNCXRpEdEF6Yg
UFhrPCoMUF0gdioV7u1v9NsQcgo3CwPOWsCM5Sg1l5Pi4C4/O9YVbym0bjI1mz+dQu124Hu/XlGe
Bryeo/K6sME26hmB23UyzvTtzk21n+s4Hv2LggW7j41L7q/yfAQfGAtX9U7c4ycpOoCLHCZQctEc
M3qWyZxqz/eOK0vdTKEtCQWkEI8N6b2X5VbRSOsiuiaTVmKWptLmDVfdZmK+43wf1nUt1WTdIISX
ZrQrv5orrdfEcGvn9iXYWul+HqoqYZ7djWrmJbEU3QPADDD4lMej9JDZ1SnmHkh60NvxAKEZlYtZ
5pltPu4LPVj8bZ80WpxN1sb7KbMG07z5ppOy/8wks+iPlC+3pl4X6eCfwE6bCuWgXcS8PfMHTwXd
/AAlbAH9lHeTC8z0b65vfxeCq/a/FKWOC0doAmuv/7TaRhMYm3CHLQ878O8g4kOVasnUC+2rahB8
zNQ1h4MYuyO+7joHmpyEUfYsrHqf6CqdVXwdrobYtMZ8IPP/+I+VeUeY0Kyr3vWEXPP8Kvq4Mv1H
WoIw2e7KyJm8dhs1PWZqIYFS+pBE/CY7lXiNhAR8pZMooBhQCAPWwuCUj3+rPPw8jSgSOUdAGuT6
dVStbINsomLULXXzgU89H62xF9KjDTUuWsQ2dC05uBICrtGZTvHKkeYQ6rNQL7gg5WRjNkHCfCJA
OtbI3chpOynElRCsAa52ee5asLIt4igT75MGwxoIEtClP/qk2RjJop7PZ1yluzqiuveeh29k6JjA
HufLuqt1VV+uxbuXR/deNFvgSTD/WrXxsPDD/H5TtM3ksAfxvB0TzkxN27Dxsy+s6Ij07icOJcYj
nLrt+EUZdrIJ5GQ45xKlslAfuPp0n3u5n+i/+jFZUvbi4y8c+TqHJfcEfxhQ8LfOPTavO2sT88tH
OpJRus8z3g0f+XgceGMQ//gWtFDmqrddnpetGVq7WF9siZUMh0T8/OSEj4aJcgg8rrkZ31kOVcZZ
F1DANMyGHyWDPKECv4pHlTEOJQhztGOxBPgqVGSOJRJW1CFwzqW+lJ6dhsF9blG3kZKKgY4ZdxI0
KCVSBHOjniDSX/5XV/6ZY+Nmm/xHh1of6KRnrreHQOlSVtcpoNIPx8WilkZ1bq0cRiUyUpTFdRze
3IV37hA8DbepYHLMb+dj3EZvyeEHXrXAlZqNubpO5bUrd07DhmHH4ZDJQZXLUpMsdo0NjOYdHyoN
ZQ4bs7b9/JF4mjR+3jgnVBQRk4271gwJ+ClHKSrhRvwbXz3Lbql62UgbhiCgG/KHrTV8V6xQ2yn9
Pvn402120+CI61iy2RhXuBHtWt+vbojXGGU5VnwZgCfLUz7TDJEkJ/SLL3klp5nkenVdMS+K8lg9
r0N0v+D/R2iS/DFnw2HvY0KKM6JO/YbsIQWgJm9kPxaSgKzZF1rxpR4mEZr1xZHUFtB2zN1MpqtE
aJHViS11823RB7vKsSzyZT1cCFj8V9k8kuf0mVcGqV5hVTFe2Ll7L0iYusy4bIX8TPfzOFjeqFd5
LzMYFBCidtBISCqHPPlXHpr5Fy3aOehD1I4o/zAoYK4Zc2Ej6iMj1l4jotkgjrpeQ/8BjH0/Xoug
zY/s3KmkM4WRCU0RswPqGeiRy+osB6n0cBwGW1A0z7/h5FIvT5B3HZKcAoxSVaj6BHRoA5w98icq
lwq1e35QKGdP7Ho9R/GGxPqIRynLxEAz/SSF9JqLKIBG+CU1rd0QDx0LF2UNJM18cWyD7p3029bF
Lfoq3tntK+LGdFY3eeXxvui2UPrsCLSR0Hk8d+uhLCQsSvtW0XI02eumAkRXC55e9muZei6D6UgY
mDWG2tYaRSGnpazm5vKwqQwxujCw+fP7KruW/2SpDmpANjw4lDKz8+n4Rnhxw0x7d2XowrWjQnxz
SO6KHfy0otk7crkIISXkMYdRlVlu8xCDJhXzS/1eetXyDkFst5xbE4X58jGMkwEHFeGk/tAlCAJI
j/PRPews1KbMyLF1Dcsx4yTYOkToDjltpaH6lkrJCF0jmVk5TGrcFr9H3LEB8NoRnI+g0ZWhCb+C
ok1QDmmrtypfNU0pTwtbTJhqo7mOhqRN7nDBcZXaAYDB/v2Bvz7HCAylFi3sfzy+Q+27AsbAWCgl
hi6Ns66aZxPeagUFiY50tj7CfoR+mOTQFx71TIJBqMW8nFT3Fa6bZJtxZg+cJrUai6PtKmXlvNp/
9p7Au+ZyKCH68ZPMwrqCgsv9MrxJp0JMWspnsxrTuBGvSi8JJLCtktmiJIWBEB6Qf9NdUx04V1iI
nmGf3Th7AHEx42GtJoRw7GBnuXCzbpDEh627ZSfxfU/p3aYzqQBnwRM0tLGiVUguBrtXVTwKwDDU
Mq9MHyJDWofHuYq5axrzxCFpqzQF/G0v23D7/v2m4DTA1D0nk4JYJHFlwjOrYr/H+Z7bGrsb0360
aq0w75S4vcDB6bi/05pwqQxUOFsTf91Oi0ryk+bxBo+ZdO3hyIHuhlCUsMaVTC/WQXL+4ZdyB85F
UmR1C7Tvj1gpUFK3r8bdQly0Gc1zGqVo7L3hAX0SQyLFHY2MkAqDs5ebqakf9DHQ9tGhlArn0fOf
PqGeYU2bBzAOgr2tEGs8O2bFq282+lFWwOCMAhzWWjvLaBILZKbTORJytNJhujNxucuVnr2SGwlX
i7rdfiGHqzN8AvIvc0W/V0JI5qKnZIRmMkhPBMtYiyBYyFiGg+KEfk7dr1kMRLR4YguMmgM1ERL0
ZswjJZaUff1FDkBLjHp31BcjRA+YU+bFMrVgwtXff6PTL7jWeaEgDKKi8kmcjDnYxsoqYiJx5Za5
M7Cw1Jy2GQyb56zWXk1gC5iFnSG9T2BfQzMLOrnf4jbbODkOYaWifPyimKV+S2913gnjaU8Z8PEQ
cc+8wQwsy3KpT2yGn9AfLy0ZLnzjjLjoy5fyeSZ+M4DfdBaDSjq6HVltmTL/TH5E6383EMzdVSqB
ZfWSuiu21JaGaAGjmAqQtpV/CiK4uhKjaO7CXRnTfd6/0nEQeWfzrkBQX+2URY7dPOgtMP0FtDcM
lVzK5+CeGppt3obAI2oFIPeKpGKVH8avNyb7e8mLv7S5V+uuQjGd28stdT1sN5u4Adze0EMhvehU
HUak/0PEFg2qDLjHT3725ew3Zwfu4pAMvHETMBCIzjMvN3ZGyiCj3WO7opC6gbiv6J+8LTWyOOlR
5ZoJV6mdrjHOuA9AEHZCnlIcGydHenLKnaf+o8KMiGND9f475L659u+itnwr9s9xlszZKzejjyQr
Gdha8XJsY7Saktl80lfmjjl55rxUWQqoMBCwgb0j7Rf1wArMEuCbye5gxrcuDAOAxEFyS/Tw/Ohr
xOwcIXuDYb4vh4pX87WfEgD2T89LamRRVG4FGHAaXUKc+iJ9WZlQV7WsJ1iIHMfR27MmBoGOvbtW
rGDCgcORiDo/ARqiemZSRO9qfcukhqA7zJyt/7AumWkFa37UrpNf9fPrIcq6eMP9qXwCXMwVifIt
VRFHJxolL2Y07totRVT8du1hQfUYnRuqs7SlUNp/rO9pcQxQ0t/PVyfgOmWFYk3ftfMIKcn53EE2
KG4KaseiY3LVzwGBP/JNC1CNeEQ6NOY34yRRdjBEq+KUgB0g9fGmptZRAAug397q3DvsfAT0LxlD
xReUhyCpDlrZX9kn7wdTJoJ00RKtj14kZIUPYQlKi/bjOFOkiXZUo/3PIMWvJtiY31IhHt7nk5kn
zk+NWRaFhMSpEWXFDyx5fo0Q48v9Weu1gm8uLApzx/Jff8lKoigE5JId+GrH1J7BE9ZlU9jSPXfS
lcvEoiSX2KJkru06vcSXyPyOvNu2Q6STGW/eLMv637SWGbTNHoPLfohSXg2J6Ju/QoS6f7EbfDwe
ShiJWZF66GMyxTdAfmRvsH7txNBZDLcR/3iDe/4RFp/m2kjVasFdWWUUunVEdrpgyKbQ+b16WTWi
8FZ6nbsJ6fWHzNBGkypnbbsFZYoUkgYZ3+fS8PtPuq6c8Bhpei2IfGyMTj5FNk9Fe0XlJ20VEKoD
mWLoX12/jcfcRVrKyqs754/19bUVdnAzTTsnSqPV02ExeEJA5Br09zh10WsGQnRM77pTAdKTWOvn
HaI/HbFfbOL1ndH9MNr5EVzmNzApyhpkWVfqImKFhJZSNUPWiBTTCfug+5ZPdhvYwHz7RZT/SRnr
p9fDWfj0Aj3Y2f4p7KBL30n67IihrUxBl72KVVIntM2KjWW1ZQ35H71JQDggZP4li08a4gpSgA0b
be4/itwCA+ZRSi81ckWvqATUZWXllMvG+UVd7pDYN5MuBhs5MzeF2Or4UM9SzSlbgKxqaAGH6Evu
GltPdLadiBAmwBIyyU0SKaWO8D0u+srSocwqc/MmH6o+UkOCVKaiFVjaSxgqz2U5rG19v4qUP0LW
m1uhvOzaJqU3zDa4a5keTOTfu0mdqlHXRkwW7tRlcsy1AcLLkgRmkqbHCglOP6XdoIDTs4vv6yNe
EnVuSi9N1KrqFi2KOC1kt3t5ToqKmuBLCsMTOI9F6IS1ZOYgbsOMYMZx824S+w1eAKDhL9eWW3z5
msdrLnQRPSgqTG3OZ0eozKuRs0FG/tSwvuSEtUdUueejETi7Aj4ddA+KQVyiJwohVs0HZBwZNr3x
lZHJ32zMIw+y9oifbAj2KpJ4wUDl2j74ThIE2JFvQNs8s27k8bqWKE89aMzbqZD5Ev1Sf3axw5cx
hSxiaqEzoxX8z5O8EJeUF8+2hvxPYOFLjQpJ1+lMSy8uGn+raAy+XwZJVD1njoZTQuWz1eQDJIAK
T5hou3Mw+z6MScfmOg9exNlkU9wW2OUPRUQcMPHFyfD4n9z+ET6nL00heifdVeW/5KCVqh/2kFFJ
4V+UWSI3/3h9jZqS4S9pUN3KBOdBpYMJ2nPGTrtBgtgWzulmtebyO6iWTDUUwaTSBd7CYpdHJH9f
puJfufl/mJAs+4//wjvUvBsM62cSZORpkYJ5mzr6Iq3s9bt6P1XuLLMNjhMBZtyaT32ZqdVaXK3U
Y3Ubaq1DhcQj6OL9HusDLF2FPCKt2L4l2xFvoCJCzBkGtzbvckkB2AALkpw4Kcc7Yuzs/99PR0St
BzpC8CEA1hxHOB7WRkq3ia72642OxxFGDLmaCwojtQC0u+1MRCi7HBrMWBhixs3l9cvPzLbKQIYZ
udX8cIbQUlBhD+v4pq6gzrH5jqON1IbnaxmRhyX1mcveuRItwJdfYBTK7dCrCR7foBEofYn4d/++
qXy16iESjr46B2/Ld0ypatxifvG4R+2g8Zq3hcUTU30K6mHVSX0IhFEW5lceNOlGg1mqOFuY2Ay7
eev3ZsfxbzPjUTxP8EZoprPUSwfzts2CKmrTiJFsHXY4blPlcTPjOt0OqysOOnxYrGthxC5S3eSp
6cNT7kuVYSB4zx87HPMTtOnFwFqdv1c3/khxQN2TKpcHYcMTePcaryqOgW2Ol5zH5z0dNveVdqa5
3VaXXTearQfuAJMhMzUaBuR1Nsi2C3G5GdcXq7X4dPVKLGtbChr/9Ed3kVZN/pxrIKMbKx2xPAu5
0quzu3Dr+t7UobuRm9aRACq/4dfnyxWC9qCXwJ557fvWRHKh2WZxq8oyj+vrs1mDeZXmnTOgB/S3
XFOnGBiWQUPDqKBokW0LUwybIumQrChRIGGGbrc+d1Eg8pCWZBDKfCrWBhejG6Rx8PkfecH17CQT
2xFlZazvPjDWgmQolQj9b2dZhFSAC+S+C0RwkMoonC7F/fKkt7OzJaYg7NHfSat8Vy8ooo5HhgPN
D2Yoa20VVW85ifACTtZE7gZ1AmAcaXu70gpq5ynlZSH2rJhAte2Nn1be9KeMZDRi9plXTKXON2JF
apMO1MI+lM4xyyFYxlEZFwnHBs1DRgfD9S5Oz2xMhNjtK697SujWm6EQH+kzIfUV6uSwqtfTteo2
BGY/M+lQxeIvFFhBqWmYaFAWKnxBPiXlEDp4S+iYFAa+ewScvRa7RQ5SLEcxHm6DW2YZv9eEKlek
DiwbFO8zGD+oVtIfPayN02+hYIdTL0npHaSh5rbfX33efrROXotD3rySYVJ5iNtefNSkpK2bOpot
u5DJPRCnYxbVEXmf5kV97knaakdlIP5ls47CHV4v2puTGnOm9P4nuRo5sZ820JvCznwT2wF7ANfK
GoyvRc6HbHe8YKv/AsNGjJoXwyRp3A21KKsKzOMX+DKi0mZsv/ElBeHlbx4pcQy3FQxwyD9Hns1b
zDaK/H0pWjJ9Say3YYkSdOi2viPW4w7wuGU/YRxz49bISm/QdrATjwZmFyivWKRhA2R/gNOZhwgr
hDRYqpLN74y0yYeeVWfolbSJ0JMxIOTgJYsvCECnfVPULwew+GQusUUcuUXP7Zb47xXA+nZ12fx8
sqMRPmdfWpCWv475rIjLc0s13nLKHQnqj8UnPj3qCDq9O/dyUT57MFoF871VoqMMK23gOfY7v/Ka
AmRO8D2Yed+Z6PtKVEDJA154OgS0rm99i9e26yhQYnlRodUm4Q5HJMuYUIwCIF6d82o4sSXT34ie
PTjGXInnXTxNTgwQ1ShN0ao4CC8z5ocYzUs1955IRcU/KcSS3SZ9HyncT6bq7cU4hFY/Ejnlqw4y
xinnzho6AGWxASm/cG4VlaRMTco5iLi72GHOqPKs6RuU5MES0ISRv4rTldN21BVxNP+xA9H8Rb62
CSxuOeSDUvMUHRwGF2x660PlL3HLqI1iwt7OP4Lnc1FRyci2sCjFf2hrY1PdY4SXvhYibCEb9bHP
IeUqEz49t7xbk11oLBMkqSFoGCx1JXTmCKLszGdfQM3KCc6flkc5+m+AGQi/B4k5slaty3hBx4Ux
9XXdO3SlsQduiXm9EAq+5m9Sk2hrabiosVoBWS0wXATKkCCYda9rT3a6M7Kyvx9hu5VydRFSRA2i
CxKfX0R/e79mhGVeVlbisp0MydL5NqV9vYSHGCN0YHtvsuDmXtK3AfGkQc3XUcA9Nnh9mWdR12w/
7mjKN/USKmKqcfC+LwDZNdn6sBbvmdHQUWI56WMVoqHY+PjAhCRXmOBcvo4XFdeDtB2QN0VOfOX6
jrPvfVMLaOkOSVUSgFk0fylzrD6rHqtjkOP9qJLiocdzeq6hW8A1BYTjkz2a5HBhaOg6YsmKN229
s76uWS7ZWtmK0endqMXg4iSU//kTJbkp6TtAc5Hlwl2HjQqSlqJ5sqmi3YqbyGHBzaq+gIy/yOTI
m+V5I27x7qh60ypEVHB6Zeq6u3ACik5vEBzhmpE5Gy+HXFuIW2GbzvnDHV8w2Iu/y57t6x7Y+3KV
GWfJUg/DVWuo9KNTK5axzIn+SFNWrVGwkDEN9v0qSzUguhB95eUrg32E4HW1Ly0CzeGUaTfhT+qL
iiDBjxz3UrFctJMQiOlosv3jjghxoU/YYD4EWXQs6b8fQg7/X6HQC0IGC3B8njNfKfsrh4tm7o+B
nOR7eVercCULUkpSokDQrLECOpHQCVlUPeBEAa4j4gl85XrFwTFPH5s27Ueo82u+jIogK8UY/nzF
SYxswS2i5s1DBwc0VINWqSi9qDu/VUQTm+hj5bONN1w6n+Ro2d5Q1a/Dq8o3kyg6vlyCDfrczTzn
PI3v31EYfYrRdV6bmfuIGRAfcWK0V+qiFOQtweV9b2CcHAIqDZ8QSZsBPh3k2u3e9VTrqqOGkbFH
gEabAa8FYT+x4jHZ84WNILKgZp4PTHFV8SxAx5IfD0dbk8D1eFqfAlrshLkUHsbFT3a88bVZaGhN
sZr3Rb8QQdQSj1VShni/Hj1UVSILSVJFn1bp7X0nCu9vMqZOPRYgLoA4dKC79YtRnUGeA7dYiMQ3
k29DsiH9J+mn2FuhP6hKZ2iWNhYWV62Zw9megyuMuz74K2wFGJumcf634uDtP8dzI7TScC2p6nDv
wwmGonI8S3mCetWYy0dyhRjwbGuACr3+oqHO/59Oizyf8t59RzBkDsXLgo0PiIeYdEb/E4udbeKv
kEfeTF16sN9+0VFEiIYbDRVwEcRInbKA4vLHMDzMAKyptXhmpP3EAoYjU9eRL0tf9pB9ckZtFQQw
ieRr1AIW9uVb25ROFhMCekq5n3FQfK30yZHj58+e0z/Owekai5KBvsGOIo+FxxW1KJTYYD+ynLyS
mkSUVi+e+6nW+kAitl9nMxavxoXxR+WWId0oFFa4TyNhLV/hjUcIbOSBPO/To3UcEzmtWIhQPKXN
hi3mTbSVJf4SoK81ziym1PL89BoGOMDeWCRPBIVRJ4AafflUNgirQlahGnmysZhHzKqaQQSta5/M
Yo455UdI/SginSWvi3ZBlCgkVQ8xWqh4jRfuhUmScKgxEclLqNEAzyvJZvKVdkOZhBtxOSEouMgo
WPOsRX2Sq3xkf8y8expoC750AVYC200a6UOun5t9witaJDcpnqUYVm33z/im7cF/OlwkNCSnota/
04Q/zeIxIPYK7HlPJLCit1OmJITR/bq9tUjRJw2/sSJw4B+K571vtgidRvkeWAh6sSCYRclOSbRD
oRATf6dcfLSX0aL67RQFK42009/r99F8yXPCElRayDeiPX4ih+pNUT8Q7UK75PhigVXVfBFSuDod
ypecGzd0JObbErY2dJ91htAxHH9pwAYiA02iqVXOyAGm1AAa2qX17ZA4gB95+SU4FiujCQkuKYIs
sL013whPOgNTjqmApt8jYtI58wnGJ6UwQL2aZjGZYef+wMIRb8ec2+LxETSqZD3sMi6rx+Aup7fB
AhtKdIS7UTjpaJs13qL0SLwUpMWNvtx1iUTCDHs0pb8mJN441aoUleGddJERr+0eU4tgydkT+5Zb
pk41hAeVcVTdei7NdtDFOx6nzhSMeA+uJDyLfP8slLLpRgWdIIjVNnQSE1ZFq7DnL1Jf8LWdXqcW
aSOOGVKgFo6OWHyqKVRe0XBVQ3+frFEc+yOUKZntZtvPlcG3J00Lc5hQbKhb8WQNhrnInA6R/ycQ
W9sG2y+hURrTYZPOfVazWcGmfhWkTIOYD9qtnNeGTI05l0yQRRwSMrqRbwXwAEf2DYdIdl+e7uT7
qL969s90GdH7nscaocGhdqbLNyyekss0MpGkuvhOVZpS3LGiyFlFeIaSmHioGXsF3vsAk3EndgWU
eD75z0BtbJCkGOxUVop4Ly89nnOZZuKhJHNGrnvuGoH9Jzzctz2PAFpgioaT6P2qNTd9jKAbFWj3
p0CNkphovD3YKrf0F24xNb2bzMOJwxkoJ9AOZOzAqbf73GAAorYWQDeitmAN1UY1m5Gv0b3PHyG5
ywfZNF/2GWY1HC+dcEBWNTbqr2T2zFvA+4wVRU5N0hVpiliUHJu3Zdl2b/XG35H8D4qWm5rS9Mei
YLNPokw555ooa0S5LAtgoZyGrfJhC/Ta8QZVAVvyiVi00ZVsD/ZE9oRXDbbrMu7CR1hSW6b6RdQP
i9dLtTjuFCNN/Ynm89Pej5Ks+j8hQSbiqXkbROo3gbFtxypZYFleYnY8K97/nktlgDHhGnsVTvrq
zoVUKEmrXoen1p2eNNW/er8SlfEZ/P4QXHMZ9Wt+dXG7SXkKisSWp75BRYiy0JAevbZ8hQl07ClF
JaCliomgvqaEkKWdKQ++YLjVztHl29GcsZS7vJPtl1pLiW98Axi3pWnzetkULP55nGdglBWSH4Pg
8yT1xpL72O/ZpAQ6dJV36oJRiDb/zWZBZ+zi8h86SShMx5j1a9IFrHdrWJOxcKiuk9DcK0hzZYhT
0MkcGIvJQbznWyij/vFxzs2dM7We9WyKaKgw75qjRWyvmS1yC5vbtgYcFjhxMuUa5vqQmgVgz8IZ
dXJv47O7UHGneRWG/bliIjHngBxwNwDBVmiSj5ra3NCgELFVW9HdgZGfFlPIuPtyZfAfnpQHOioE
TwuTM9kBUO08gCiRmbeYBiq9s0BvH9pPZJSaqHcSoviNYFA883b1+08RF8uEYWomVjRI6IkDBiqU
3fs7sbNUXTtHE2g6svVEbeJ+GrZorSjPWz4I6omScHtKQ63KEYwlf6k3J7K02EXNakZqbgtb1oFz
6DnVmxkF2ZyDH4Eo52o/lFA6W38lMLc0mJeVC7dmQycivEta66tNGMJ0YouQFlx14Wt3uiWgd2BE
D+A3SmUZsTkrNE0u6lRmeVlnERfxBs/7K67tkr2Jc3QaWx0Ze7WsMmGJ7Y9dr1aaJss54xMgh/w0
+v+scnnfCjscws/wSwgIYeWo0tLEc/1u9wRuzd+2EguH/POcSD8Oj/VCMJ4vhWv68Ag5pkivsdcn
JNi9fh2+I2O5ZLUeq1x+B2fr/2Te+pKJEIbGENJMfwH82LvlqKwe7bF0k6XZhGiHwINzUrrzmWS9
povjrMX4jQBseCIxEeYsLmdKT19nfm6SHzvWhvTWjrv5VSTHaLWeQwO88cFkx+ENqjVtTgdpaekq
SAjHeO4SLHIo/sSkSQ7o8HepQWsux7LqsFfK+LNgjcNUYd7l9NGKreRS1Ian0mVDlZMTv3I2lI3h
8MbkmM28ascX9wz/VNcJETVkTZi/3DCl+R5JEx9FU6FfOS6X/ibqfwoy2e/hUvmhkw55WRA48je8
JmsHJy+vwXj1IcSKal9NjyJNoBS9cFOSvlXpv/WTKw3SuBh0GbWu3w/lYxekIFPUcTFS5Ybu9quA
ydHaP0utZgRNxe5IRaDb+vIeXnj6suhJ+bFUFdJjVkiS9Jzws39DdzP2WLGWhSZ0Tih5GVPLalV5
aZd5fip70ooswzQWE7YlS/6O4YDwRFxUTj7Rfk8wBGHAqtOglLP6PSUiICPOhX7S+tpnpG8L9fex
Y9kyIp4x6civpylL8aHmE20E40Oc4rOPbLs0V6TvIIxVLZ7JKwCV8bGPyJn9Hs8r9cZHv174JbUP
PuPyLJ+szr/ckUzFmPEBCxFY/iaJcMOAX/lq83SEVFjuelRC2X67OmuacSBX/W7lSPwp5GCmJItt
+bjR+rBE2oH07MFl9dAMuL4AqCVzeVz8Ha3NAr9phC3HMuY75S7gF1LlEcDZdz8eL6TKK26w4cjH
/zazB7vOVtcKn/ROgDNIG1+ZQUuRVJT8USTtb+v+kcRfYLf8wtLts8cMDFODQ4NJ4EQVkv1Jqwjk
tslqiIgJ0zhvbEHvtpBAQH0nUso4eVZpZ3N3sm1rEJKh6IP4DLlhft7gh1bsF5H3dgy+D+ZAqMKg
nDJ4Xkxl6CIaRp/kVAy0xYJ7rDPHYbt1djAZk7jzntHi9dFFr5DaejFzZYHnCqouuaZtd0z5syGG
jLgczqFOd0+VRP2G7/Skw+NUR4mcn2HF7qoDFL5bmndIR6j1OFyYaWXNwxRULRKLYrWxm6A423KG
iJhm2PGC0uCrjc9XOAEKe9vT4h0e2f5kVHZteoA4NWpNL7xX75+m402qXeCDz9qjpGRLRpOIBYD2
4yARdfEUITPLbLG3RR0Usio4Ne4HqIPBhWm5zR4O0zqjA8P+EYVpl6fn9rvUbQDIshD9WvoNi0g6
bqwroDA+lRzc7A+f9ZvDyYi1yK0HkGv0FC1XB1P1u3A91NOEOsDMOe1Vyy6rq2O66H/OK7Rz7kg8
NIFYsdrMuG74MBS/7NTkvlWSBNDbXSSb+zoOQu04y79m7WuULl/d059XEDk8O1KmOEF+W+NQiOf+
ojMTEfj1Ho4OZjvQJN5Gw4nPGD/CmcTVBcdMpUiVucouFBp0x+ixJMzNQnsp2EABAWPcS3jsjDfY
607J0AXTaCyqA7Xbs5gV+tGL6hl/N5U11mzKKmTZ+MTnKojxfq1vJmKg3hlJxX1vsGfThZcqp4UC
IAKpGI4JKDMUwm6mP9/TKbRXlgMJCaVy1HhwxpDMKVlBEmlYBhaBSCYAH7FLKshRft+HuPBHAKor
8firUDCCafjibbQ2kmDzB25lKdW0QRBhXjlz9agCgf5RYvW+YnoIPsZB0k1DlHM421OBtl8O9V1+
99hq4GzqJYG6rDacV6qxRp2DEevPIXBtV8NHPaEg19iSrWSUUWo7NIGW/zQz2dFBGZeNNBwK0ZRk
MHFeuJLwtJ8bmpE/SO+WcTNUtVH/OZxbxN6PKiCbGFN/bi5x21ZRzKkP8RjH/Gmdqc116KZ5nsXa
XpOmv7wPJLiLTBzvrSrzwekXOCXhDdrfhQ7158JWa2WeeqmrRpC27EeZGp+qcMnWu+Iqad1D2zpb
neX2DmMlg1INr//ovh3DFAT9GNbxgWSb+GYV254xoZJrVSknZPnptfpmJA9j1AIH4WkwGSPzB3kD
TJJa/HAW3ZLBblnUSpodvYDsUW99FkBuqD6ak0wvaPUcvQdb7Q1fCC+C9jNpS//CxaBKj9xoUVvV
y+t5Cwr7Zjd/k1Z2o0ckq5G2leUyjXEAiTNKf2dtwYESFyDbVsWJhIl5krrxSAbbhs7fsAwKu0xQ
H2qdjpjErPNm7dTryDZfZU3Yxw/8XQoeZJ6X/aoE6GPYw2StFb3UqaGrfbHJsdHw5yTrOjuv94Ip
9TCNRq78VdN87ciPLPXigssBjpoiBjsSKK+1icFggx+lVV6feqyvvbDx0A0+X3QGnJl8BFbvmSQA
NqPo2YLVJatgbYXhZx7PQxXcGPKsF8vo1da1wm2ObwVMgu5nlBLBj/2dZrCMtyo9qwOyT5l3NVcn
UldfJry4STJS4uhj2IfjxS8Wzy1ncNSJr4LNkhB8NpSrj6evsX0AlPSwG6L7AQqf3fpEdW6vny4n
R5UefCCllx1i/7V/Mc6HFD7XBL1VrMqLn64iirSlOMgFSkTzr6ImFR5hmuAZNmwLSVeFYPOxqiHC
1NBNdKha6h+HZfferKT/LNRMtZmlFqtTMGgN0/Iu+XIOumk7VT0GwXsIENoX2XepWQ9ut/uREdZ8
bc5HSCeMe3RsSD1Xm30/+nkH1ASSP23NMYaJ8PpjCC5kR52bykMHRrXN2lGbKrddbv35nT6UwYes
9CrU3QmNtTzeIrjqKnS9hsMVt1lgu0OM/+T1neLf1o7k4JD8tLr3cOkT+kQyH++v0cpTv4lKN5bf
5XiTb1J9Z3sBw0chCTRpFlKw/i8uwzlXoAPX0mj+u7G5nm8Pm2Z5eg4T8PiW8aqNo9g6t26eZID4
I6Bcl8+hGECavPeoSpHbZSuU0ZTIR5VSzYl1vwO+kwneWLi+ZTFOAD1qU1DQcK7TghAuC90ps8LR
TA6l40SPks+L/aibLULcaviKG+kCtekwaA03EvgJjWTpHePcW+jE+XmblAvUHaXMuwm7uagHlvCd
neVvKXIqK0yW9pMGdNo33B5wRlRMSsPDZ/RsnkjZvwphGyi6qoz57KGIVaaHSEnGfDG3YgnHwMEp
KWYO6h44SVquJtBKmDtiu+EIcGZ/j+4gDVi8YdKawhhEgxn5npLXFzXBg3ZyH3CqNby4iaFVEHHQ
H0S3ypLDgY7p3scMos6myCXUaGhUx3b5hf7BqMa4/R6yFxWPSHE9ghoYisxohYHYA9lJEQCALi+V
v7tmT5XUh8d/N23SErm/dvD/WAyW+1jOseMo7y4JvSjbOVIW3bPZ1zmBZyMIELPhHFh8YBnPLayg
jpa8Zup5R6CN7PasI6Af+a5eKBS7z0dNfeHSBAKKeBqqZ4/PEu5njXfp1qagVHXMqtoBJtAihV1m
eMXi4MhDjV3Y8i/2aqdTS/4/7Gd4aBbGbXZjfeFHFz1Dy+LCFQPumOodkDAmKCYSdiCTGkmwPQBa
RXTy4ijBfo4ynSLByPYJfPTEhLOVEwZ/PhM7R8y5KLnIo4lVDfabYsQIQe9G0aKiGsl8/TgzkdMc
9++Dsm83/s6wwwbdFBuBzI2d9sUz/QZmPiTD8MfaJFOzFjoDzWmBBGPlBHdeHeIAEH+XHRcTdAKL
ogEUKSiH2cf5I9M7+B9fLQBtstX4unJASyrCDitEPX1OPuSCSledJ2TF9130WDubfSqw3o9v/Jq+
HuBuYJwlnE9w29mQIfg7OfO0n6AcWgPCxWc/c3y3b0AOQJZQk5HNFEc9n4WKV4AdjdFNrmOYZfMl
Y/Wky9zbW4ZRePtKR0wxtP7JXgzvZMlhiGwerKjQ+WJAUpkGCkE/0x2WBJ4Eb6l3wXyiDF/DuFJX
GZyMNvJvZhPILdGCyyGGW2XRv03pCKc5xh0OhQDH3ztJtJ4J+GBxVQEqMbua9y6vA3j4mU7LdhZD
6u2MLbdH9dnRd8tucxGuuUCGzrQgaqfzqGFPJeVUtTjrs8a4zbrHd8DYNplQsu3WcGI/OGpPbCsK
rQfdeq99fEC7tHEs3IxJ+ERXktmBwdqzZYWLY2YG8zJ1ZjdTgBJiW41X2uoOyxkmpd+lza3n78Nw
2n7jMl1aEg1UZFYxqtf1Pntga4x3smrW1FjJ5Cwk4czuctoSiB9TDDuaoSg8XejeDjaxHzEqhkUt
5gPyUVILyke2jNIhQEpgsFTv9Llb6bDNSPRwg8ueXmCnY2HRYr+fUcVwG9xDGHNTnEN8Uu75vo2m
uBI3dDya9njPikpcgxHgzZqHqh7F2COg/sKZI/8XrAAPUENiqOpGT6U2oETATw2eyjcYyZBgqryy
Bmel6qCSnhYoO/dgOZEYXVmi9Pth7QwXKZuXhvZmx7MV96fIYJBuwX2iH1u4368dFYh31s4Fx8uO
CnXk0v5/BnK9do5WpKC+EEnO/SIK+3bJilBzp3cD9qZEwMtJWF45AwpyEh5IahpfgV3bCkZKQ8M8
ZcNastvOM9EwW9HhEnBptYuWSKVvoz32SfgMnW+DkcEQfZAXFaztOhZ1iIHGWK7LwcXrnHZMb5T9
eigXWXA7kYUPxjKqO5rYOUdYf/Y6QYIZxLuxtJ6hdYdj/PV9H41hd0WoB5TsY6++pixeQdR1knor
baI1tMK1EW2Nn3qK7pCxg2wpODKmAYGHMirLa+kQNARnaSg5iSoIienSA59mBEePYnvS0QPb3ZAO
Q7aQDQCRlaQhrbO9jfQ7ez8emVE68bfE0uREsz3QEr7hFPs8oAUbVoLGb4yZulqm+TxCszk51t47
mQ1C8j+uOYfLZph1BuQMzOvFNtUCZXJe6rPn5lKAoEumX6ufjPo9gg1QfGg5ISTLJkKoDC3nNEkM
OSOOm1gKN/W73PUS6Qt5YZcEU3HYHLRuJxP2YviZVOlc7iGsgOr578ywHNMnKYWGj5TV/IOjhnWs
0pN20vO4KlgL9MOyQJPzioH8BdjB56/Gx9ie76MW+nG7pmqPHUJRislse9ihflFvliokpHW4qZgM
sPjSqTglnAw34d5a0u4/0AEr8/vBXfZRQqtJbVlksDYI7H3tmatQcjregPjJmI9KEALaF7YVm8Lw
nCOFvXz50joADNRv2FBQEZVK4ye9zkoRCg1etOJOEUIG+YV0eiN9NtESQMvcTDhMtfNYwHrlZ8b/
jFlga34H+UiXhyIwbMMXkaO+wr72+Npwt8+tfo53N/X440BdsQFP8v77U75xdvm+Lgi7NEbLqdgI
GwMj94KyMGdyqU0PxB+/eMg3f37XoR0AQp9NyKo74MEjbOvkJS9CqnTIEsCx9CaWF2TGb9ZUwdK4
yDoq7mwJvIgst5dMcvMx6JMFXZuSaE1e1WIFKvCCH6t4gwgukaRcTv+v4QzqQypfoOBlN5ebacd3
kldQkMRms1ZZ4R0DtvePWYAXTsIBRX/Ns4WYAtkF3cxqcks7RVwunLbrB+UR253i2QsUbE5N9PPl
YeNDJtrrUbtjsiHZccpky8rKv4ZCsp8jOQ0l4OoX+A1ECUUUd3aCxhkdL0Ms8cGNUUPxcyTcl+KE
WGAnCoiGXuRLkzrXyUizilALMeuZ/O3+i0o/xgn44AGgnDMzfR7yzI9pigAHCUuE0s9YpIWSaYQu
XpIaDJpgIUpZEbFdoQn7RsqzGaxLm6UuQcVE6cqXSj62NQoU+c+iZ9+j80OL2/MRQCRfsTIypjH8
+pvsKbKbn2Rgi0QhFduVvE4ZsTq9yYPLKhWgmHCyhwWaByXDHNGPDRFAW0KxqkHS8pJPOA81+MH2
ogqFktYe/uDcVleotpyv5xxGM5Ujdz6nlwvC7aAIeVb5iWqNBG4YdGNhjUbE+HOI9BW6QU23NAdJ
d365mtkZSfCwa50rQphNf8GFi6zjH1E+AO0m1LZBNuqGhCNEnjun4tbbBK02+xR/kliQ+KlOtaYb
cmOwSQ0osQR1Wol8TC0pFdFMD+EE7r83Azknc1ws4NQ8yymzZm7DI9Vq2+HBTWBtwx2l6OtPSYRK
vLEBbRK7KkLHoEzhSdORSQ7V6U2lyqePpn0cZv3mpqAuuWEuvJ/cY+u67WS+oCnm0TljzFj1IsIQ
ic9c5MDUV3SeAnaWPh5MK2XLbq56OmKRC+maBGAV28+B6VzXhbnKL7dPtBl+BnI3oeBmPW5g38ll
l5CHY6ihTdzMR8t8Rui0+DmUZzG0xS4RrKgaaOO0rEz69ndR0Z1X2lSe4vxIsyJpMXq+iPthvi+S
ltW5haU06/5wgBqubbGEVYAzu8GFKIaT2VWvjdrhfgR4L0HDycqlwUe2ngSYx+LfmbkQKhBSPzIV
rnbxHw3WBuBa7DPY9wolwQAU/TJFcRAs8wt23ziza8ABou5TXz3myLcAvK1AZcSHSkLycIHSbY5q
4529kMsqUoF7AZIselRF2wyNOvRQTTKVixEYRcyHQr5J/de7nnTnUZGgmyH/FYfrKUz/PL67X4q+
ZDQieuCfyxiFAGLyzUrm4wg9ZKhhnX85kQKPo6a1VU3JCwIl2yUEObsDJ/2kaqrFpsTqrdgpmZjO
AGXITyFVXaJHzFsXJ7fKazHNoyAMFumA9XugS96qbT5GnhlBhNYzcIigW0/XHiVIx4hGoBqPS5lp
XByK6nIqQCm93FtG9lSwLOR998Pdz5Qgf3q8FoFjkXywRhmHbiEke9V9c4/grxAuiCiXUISF8imT
+HDjfzH1QfYb0c/YIpevNI7V55z0TbQ2YffmoURD0DA91ba6yQXzSJYreYMKupzPfrBy1NSKZMZo
D5NHqZePLdINGxPVCNbJY9ByGvtQUiB0vQXZPu4yfTPcDhrOMMI8EiS7L2qS16P+gSWG7xaE6SVB
XfhdHfqjreX0Yx4ob7MN1gE7qNImr3A4OqdmbYOpkKiiW3suYqkLUm6FEmrl3d5em5ggKPWdoSej
gD8FnV4N0iAppK88+/yTQlpSgQ9/NMIj6y73wfVJi/r0bahqRu3KIEzhpOecAxsDr9CFdj8ZaJdp
EAeTF2P7FlZltl2Nd+6jFRN2XIv6aQz6BSVpK+hNdI6i12SoPpcZAOeXGZNx98igAYbv6ck+Ad8Q
GIIhkAVSfyzgyFKqbo2nkX1ovZcLYkn+axbLPHe42ZGpsLTMruOhO+S0OY5WQs2EA16hvItkKVO0
rRFPnfkzm1YKTHbyPPXA73qT+svdOjvk8FOUIXgKA+zvz7X63xPsc0FeFMsxmEV0aA6LE7ZtAOzn
EZC8BE1dFV6O51ST9oB0gVZrKbby6pAuJq69k+kY74sE+G5CQ3Rxj78PvxbfWND2wrbR3unQJXfS
MV0cJwBCVTLAXcnrr3moJjUs00gh4SjU4v4zEYEllCyzJy0hg/Hp2ISj9Bt7M4olyRwSF+hE9o9g
1zOB98V+0SUPesw30jqMGg5+ROrVMFLxGVto7ptSz1EIou6MvcMeiq3vy2kAK1j2XKuHrvNbF0QP
zPMx5bjS/DfyMoo0kB2WqI38Ja2Ed5Uwc6/YtzMBGpDimJXHni3UGstLF67zp7uaL+jklMCuS2Pz
qKyRGPySE2rsSDqS1/TDkC74W+PMXJdw/L44gCLeR3yDkXVEi3Yw3pRT20qjHoKSQdiBRywU64m3
JAr5JFIV+eFSPMbRfaQ/RUh3Xeqe+7pxEHn26TomxtOBtId4y1f3AnS0rxvsRw9FW1KECGk4WrHr
ABdxKUGFJmOVdiuiEC4h0gC87QNFRxF/sOWhuocoYZGbBf6hhYcVQ4Gi0ggghCSsEtj0UpQExVxq
fH9lLnAJ73itiToH8GLKim1rwlrMRC97WPnFpD8ZeW5haHeTeu+IWmyVUQK0MMmkUv6NmzUJ0SGO
hcibIPDaZydFB1uVaT72YFk6X270+7rOWXpzWU75+QNs94BNe3msdIwdHC3BsRkpmmgAndzvD5Kj
0o/i8+oZJr3zai6ZLnfLAkjAAUHHIrUTtoymAwmx8nUIRpq/hosdmDdBp5Gguv/I9ccOmSjpQBrI
euRE3Mqsa5+3DUQZYWHj/A4SW/UiK4eZgxMNXhFV7ZuNYDaoTdO1CzwB7JllEPix0+GLtZQWKc8M
OoRtwfIRyXZ4l2aZfpiLWlWXt35+S4VxWGChcG4uIrvhjYGafe6UwO7uDaGyfdysSRwpKto3TYRa
FylyHUvO2rC9wytcrA/WBa/ufvtXKZoIqA16xhqE/AmriVkLXgRPl9osNks3bIF06naVvJ80A6K3
5DNnWRn7MVGgLiglEYYI79FYxtYCNG0faeh4xVGDjrSsoiOilnqLHmt3tOvsbkVhSk4Nq2NL45ng
g0JOoGgNOG50m7C4IsufUJFSTWsrPsWhysZaS6t2c9m2aa5RYkqqOlwitzp4yP1Zo9Bm+khfanfC
Kfz8ypMe5dp2Qz2TTLaS2rTh807dxtDI1Hdquvzk759gat05LE2N8NX44NRSKDpiMxqY6mHciCNI
WbX1UadQORdwnieaKc4jycAKfa9Rja8cQTpr78mKlkyMJ2NQty0YXfVGrc4VZzREjY7vq2tpPCyc
PhzGxXKIaHOXwZ0En+J8sTUYDyiHlg+I/Re1A2oJVVPhEJFyZfBGq2+hr5RDJ1ErmZLIpykfW9Iy
TnJoCqUIASfpPOh5E9UYCzwsADvevpyzelsR8fMbtOxohkj3ARJqz1p48il9dYKKVfvEtgYO19vo
0dJ8VWEC8JoExDzAw0HRdulZVKJw+G6O/Lv7+Mm7Boj4ArQ6TCHn2iD0VhLmlmakS6CfYruEwPdP
0m6ln7FhvHaQbFMCDiAwf6vxQL92WOHE/I6Y+qZJS85iXqEP3L4bZB384PHe+bLHsoYQOf7EUjxB
cxapVBVvgISWp7IqFcKytA/4wL1a7un9ldNm6vTrG4JTpzjjUsy+cRK0sF6ALdqLnVimTaVz1MM/
viDzBlbl6YuZxyrNousqPpzKsHdLV8+Hx1xPC2Mii1r7raE905FH4UfQAEueBUAb83oA+Qjb8Hr8
Rs1x+caJMDsIB0cffDBkpEi2Hw8rRuJtgy46jebKcZ61idc7lk2FK/7bps/Tlr7wLMTOh3UmnlLf
+dc8gYx38wLuuuBVlhQVbUDE5hIXP6GUGOs0quPc4DO+bpvgI7x7Y4PvAp7OY9EpeBbhRfr+cTHL
XCtLmRFaTjcnD2sqvwIFLpfolYyExNrNVxUvEMEaszl2vupYkn0Ynlc5oTKjeZK9spRatdIuP5Uh
PsQojtHZryfQLjhKeHC1TQO1lBarXhZVrKz25RuEVOvaGd8vxPBiyxtQKWxVC6G+UoRrW7OcvNQh
9if37jtYesrMYNZNHWIMbN1vgJ/tHVAWRxApxwqQuWfOAvlDzE6BwPqZiz+Ud15ZvWfQt8xmxKfK
i+th8j6l32fzO9JDtr5ATDj3YheED0svsbAQZ6yhHeu0Z6ll5BH3XlT6nsyxNaYGH7XQcWq5iljL
o2uZMGUdmM6ALfFnBWNapRPaM9hiJy8BCSQmWruZzNPcLxnvRGMRHDXskTnc1i/Hs8SmsSUegH/9
HYkXZC7McSIhG+ivEH0UNtAm/UHVMpwosDl4sdAoZ0VX/iPhdJ/GKMKthY1APR+AWIgdYvQgebgl
DaKgmqBj5CWa1FwyP8NwQHSmN9BYIu3mHFhA0kp8B7RangdH911LG3xbWOhVWsftbsB3X9Dow6tG
RiYqcPcyDRKUv9XRE1qZXYm7mkbstyO0hXOJQ7Kuz72H1CaTp+QMUbuq/jXgVIxuekYToitZ1IzM
nPuN5hepJ/lpqbBERjF49+JbXq7e40WLq2I9KWqJIP3YkTuy2+dIO8qb/3OYbtDUnz/60Gr0uWol
szwHgRIjBulYRW6RLg/rRcqMXdOrtKRd4NST2J8VBowh0FcxnFzy+fYIO9FwkpRCR8taaDszzIft
UHrMGCOByiYRR1OHmhIPMxpMrB+TmsjWstoCmuasvh4d/T7v5P2E8bn6a6B75AFBMZ0NzDPFy551
mzjNVzGpBc6AVyyx29dxSSLn7jGB/ecaAm2ZaTuoLM05n7vECBW6ZcpqTGY+gJPnDAIshKjh5TYI
9ldktWL3PoSefCcLi0y68wTqPKIDzQghE+Xn11iBZJ93A9bEouN4VOfS9ec596Up14NPPdmhyBCY
KYK6kBSTg9WHEAyWw1UaW4lHcT3jvemN1i6eCTmXGVb8oLgy/MBbXLWYgjzPCHRxCPmXN6OJfHDh
aZQ4bjnZRyagBwTW2cx0k74T69AfSaNiksDcC3TrIyWsEgT89ni3ioQr0lX7grRpMRtPFotGQQEB
Q+0O2dhBVbgOD60RNyRoFAspN+WsJedRYleCCiI9BQoL5qy+idZK32LiH55yFkqwUOyAeJ8IiJM2
W6njf2iEMhdLE5qp5QCwk/b/Brv0z0+C0IPyMQ2iBDMJd+4NY2duNK+Xgems3nzkqAXnhoOwVmS/
K7LsXhOs6tyWBAJ0YiCqSWoqkhCrDI6IM3U+8zcuP1VPjfSAvCr0ktYUjbWGASJr2ooebNFym6iW
7DstgUTd3942IHJkAtOHZ7C8vumoQ3zyZ2KOu3x2Ge6qwcEhA8nYVZr5Fl9JLvSGxpRJD9eLCPJe
1WJIUmSn6UvgBbNoaHspwj7lIW6qWoYdmgUwlus6onloiPxVt+lLeoRCL8UiyptIOADazt8echsZ
ZUqSRAkNuvfMmyAt7DvBh6DFOfkxZxy2ZjxmE3NRKKzBZgb7Z5t86lQjM9QgqDwmCUkOPujTTFqy
8f5TTrm8/Gn05AyA3hUhLwL2QefnC+9jmL0lDyKd6iUezKlTXFp9iHEdJDnx351K7IiCienEnqW5
ZmJVgPZtfdGtIrLZv1sShxXdv6kSxrWhGNnUeXfmhSXcEqN/3ZXJ/bVCV+LbsasZsmdWkoiyDaM2
FD/jneELUne4JFDNAYW1hRHR6yosWDIYO+0iZNUbCn/erUTSgYNg4cFRWYyguXUOhV4kfNdjhocc
cNFWcWHzRTC+d4PEeyBH4jJgkwFDfPTIeYgHqbnrg1HHMUrHqCBDT08LEx3dhLfX7tfYw5rQ2pyy
lMjmhAC0JnK8+38se20HDIkphoTiBKML6JGxVIkoUaZCTnsP5N+Oo7NzyKig++cqkKrZx1cADdXp
feL5qmBjO2n8/+SLasLfZFZ4sjXbXFcLTQzUFHfH6SZqh1cYMXTgWDSkR0FXmWYmkWDhZ4NB2r1L
l4jI7Rfn/Mag6c/THW0POTM8GdSfBk7Zb+ZCU1cDjC+kdZEKOCqo6z66xEot4lqQphN7SVdHAwZc
UxqfwNjQBA0uv+p0Ug9+Rf3knoTEPDJiQ18SjG5rZlserNDyD4qlj+gXhk2tHEDD4vH+IG8a48xM
bjM/lniWbEWTIXVcFTt8UIRK1mb/OkemQPya7PZo2saCceZU2X5mtA3QJTtQuGmnEgt/nV9VjjQr
BWoBT6zNGwkyjtF5edQks2idKgJyYRSMO9KaqkeBQE4X1idYnb6DrGraCd/VRwZ7WzUUCMQDMqPE
Z6Z2AqUDzwgMaHkOprzo1KUWaRz4NS1KEEXVHaeKo+TUVYKy1V0hWkSO7qaL8CMq93IsxoVkdfEt
IW4I4WNoYuqujlyrpNLiem77STLBMj1p0foGgNEPSfl4DZlZ4OOfNU1BGSqVQ0EQQP7z6NFhqlD4
RtE6DOybJ+UKx9M878TICkVyrOuJ91LpAw5upax4C4EiX0lnNQmS+tux93b0lqbfxgUG56nes7Mb
a5BZkUymEZS4WoCREVt+d93rqAzT5HcF5gOvZo7tCefz5u7nN6fM+IhVUdIs/QLlcprEev6KIvKO
37SNiMmAmoBUfFpuVNFbMrmrJS+YLgcaytT2+U8Hu+JMDIX8FEz6O9Wo6QrB8Q1LB64yLb2MLVgu
Zo8Kr/f4+vUexsaWbCv/71HHfqU99I1t2Ib3t7jE7YYcwdUqvpIstl2dz9TnVpaVSTIH1oUH3EVC
wQ9350mggab59vci5zVYn/uLHnC5tQXTSHyFgUH5flV2IbIEqWygW6iCbOmUch/Ff/l92WDhpvJG
86Cspr52TeIB/I41D6ljASOvuonwqUklDq7oJRBj4SG8bDiOtZ6qOJGeRiwurEm+0xht5HWkv41m
gc9fNDCRl4/wt3mD5lSL/TydwcX7+p0qytiAsq6Ipr8nVoz4bOzVGS3O0ffgwtxE/U2YAeQ4Klty
WcKpLrWIla5FM+cIeex79J7JqUB9tbQ9lZmdj2RZbn3MvxcLJU+zV12iy9aoTK9KvW1jLMCvABqC
NUs96EkEQDx9QpKHYABq70t1KmdrIP5lkY5+A1sSSkTqgBkSm/MpLQdDkGCbiVePp5qAo4EJ5gMw
aCgmVlTZRiqTlgYy/9bpkpdQed7jVD4+17KfC4v6W8VlrLsFpdf67ll1dNCGdQn9zbbMUv8yite9
i0dRZ7wLTxXj7IwogH88UBvV/THHG/5IStvHhG9MkhQpO41IldokGXKq1dLkMGJQO5esVa9PCgCY
5BWa15KFLfwmQ6R2CLRlDNep0ta2uemCp5eCs/ucYs8kYE0/W4QcAZq9YJ6OwFlIefVCPFs/oy3F
nRm2pmvXQWMEYvKH4sJxJ+C8INH85yvS/RoG76X+tEyWLs0uDGVBAEJyO0FPqbel5fBl776q1J5P
kOH72zMKvM/Huut2njqhOdvogc8nV8P2gkvnuzg1jjzBj0/XmXNe/7jXA+C+2wRqcYGiRKOjfaly
JRPUUWqaBfiP/QGPkNOCHE1wK/9xl5NeFJuT1kZ6vmMRS7Gf4fOdGAWDWOpK5zKikuNRfuY0CniJ
a9kblR3W91XBB4IS8902xBZ74J7ugK0dt0o5fDcAR8EA3JwZ2sG7i2+d1ujq0vIT5RvSBEwsMp5K
MP/WRXe3IHPHeu1/yKtzn5FWtqhE+mG4WDHmQaeC4cJslMj/8qjVmWThd/usZRqgkQ7ORJCbksZC
yo+6Ln5JLaSTNAcEZvY0Dt562OmWZesWooag5f7503X1UPBSsGXFhnJn9HT0+rXaRLKv9GkALIzt
N4VIxuF1TV/hBoQIpFnvhaY3sacDGynN9e3UlCpGIbnhK5Uhj0cAyvuDSBeruwQN8crWDLVHgqOf
TXaSgh/YUzPEb6fwpw7P0a+yCoIN9vugpqdYQt4JYL9W6d6wXNLkrgQioAGA2ZB30IzYHMDthrsO
LFCXOf3SchbBhSe04rvc3n/onC9hH9RYbB4YPjgLBZUx7u1gUwkIJTEDxG5nj7VphcwLpLgnUO/q
zJXdVXEhKXgsycDq9geVUdyXxyJpBy1/8WVkEw3Nvr0QSyjJUCvY2wFLuOxAesGXWp28z3OkYi3M
GifVZdICo+ExzyGpwXSpfeY5U/cVURbEwHqKW1UNJRU+6Cj5NMHb9ksWdo9pwQYM/LTDtII/VcV0
ztvH1V6DEzUWJiAe3UjJYjNdFZXdSqBsW6cyZ/FUAih33UQsOzwdBgqqMuxr+8WyCphs7VZbnVdz
q1hU92YgLVnnxtEv88Nkww8pYnsCBNkW0dX7/UKcl/20RyZdjYgBPJB/yYHNEh+Iz8jyoDPa+prs
MzSHii/uF2NBwVtrDH55yaBBYbWyM2DgP01dkAvseRP+5ITgGoAG+P6Z8dgL9RtZSHsZqi3JrX/A
Sgw63bmAjXGFzoXrEEhJBiBawtoz21BurQ/zFM2xUNsmjrjjv2qLsVLJzhJuPudqYrMkNv1uNbx9
ZkxSdegQwEEEKAfT9E2uKpSpLiTG0DVJey/ghNHC6+HzRM0OmJYD419a8PHLpCmUxwZm26Fwbv+f
4Z2LRA6bXFMGENCJbB/TZRDPBNzImmu0lN1hS3l4FffhCRpTGQaIzDaJNbHk8nxSiKm4lD3Y11HJ
A6Kic2YEStRoimW28yzM9wQHXCbAtiNbrB8INQtwrWDRF4JXhFzpRYUiBkzUs4GugFi9hsiRBypc
9kWOoAwCrQA0QyNNxM9py+DFlhfM0z4GSSD4KxA7xzr1N1/d42d56R35QJcuYBA0CzeeeoQmfFKf
r3F9nbKTref/PGSOuVSHrC8gi/GOIKa1VsPQ3xTErS7NX88OeARdvjwpVXoot4sTbm30ZAEgsaRM
DfugQwd2Gkam7NivmyTsRMSI/2Y6Sb6RQVRk1BctTy1iaZb7u/t1mo1kJufK+DnEEN+MCY9CMQfR
eq1RWidWza6vaeGK+4UZ68rysMkCjn+joTspffRlfLJOIIUUbECYEVxoEnttyAKo8e+8oj5J84fc
FLJ7T44FNfbuPsDQqL43yWBcjwqhQJpCBKh1ghc82nKbCyzvpYQ8NFpIG4W6LKno2P55iDKYWKA8
bLN5IlEEP6VTCH0VYUmVXsX1JSFPMdPkaVHSOjOwzLivHQxJlmTpcR93CQlNeton8Co9rSFSazMh
W5+ST2EtW3be5f4pRNf9t9N3ENH7bIRLijhavScs3IvNFyVUBBB4S7oTkaebqPMSag6ff7tuisIa
dfMWRfWWGHzWmA4FXnFaMDkenoYlnCTfjHubUeaX4mZ6nsMRy3JNNRlgrw6dXvNv0z+hqDk8nZO0
pq357gMmjYzed79892OAlrRIdQUozU/vRICdW7Z+4QZRkJAVNC5jtDA+79/HsjI+YBVPWjdMvy5O
N34cT+Z/0FFEfTVOG2uoQf7zeKm+5048x4YdmfVO2oveW5ZzxlsdMcz813x1tzTx4mqg957JWtIL
Nbp47rax2/43v5jIAN3C+inefrRvbwsse/lzBwXMg83XMwHwcQn5xeYOu9EFWHT0pNRVC2pRncS0
oG993o62NKHj0KktfmxDqn4TuU686xWEryJ6m9udGdO+KR1uBt2FhQ4OnRaqlVm6iXbhNj15s2oQ
Q9EbsWBQ7AMx+GspoNA6C4cXywAnJalJxj8vZw3NW61kicv4S7kYTz/0ccVdGYLe5uBHv0Qm5J7s
vtLBPOE/QkKp3eu2qkIARCDmq4wqZdrZ7Drk83Evpvl79lVHehKCniTBkgZSQK+/P71rs2oxdy6O
ueVkOnY75eRtO79VqVtoBt4AKYy5c26mEuBI3auhRqcLyf0PAO2NnLj9qzaHP7VZRAzHqZoVVdeH
gJLLziD+ZZNMQh+QRDsd/HJzdi1+l7HFc8iVdV6Ez6t37F7n4q3/Sr5L0+XcgWEhCy7OWvpcAPQS
YmXCbVQEkdR1huPc7U73MaAG5P82o3QR2pVR8uiqidAzjbmeIBMKGX999iHpwlhF9x3uyXyte/b4
2NyzhQ1c0HdGtT79Tu94Ji9/Q3SroPNNakf70n3K37EliSVymwlSaBhRMFDAPtm8NcEuBFOoYqdx
lvlldzqu9q2hm4oDP5ozTLeoie7if5noNJG9bC6waxD2qVE93h9gSjKYDInMBQWhXN1Xbb6pulAY
Dj5Rp7jndr4uDOaouZpj1eQzOd9seO2qluJkfnwiEPk+RoJ8WHfxBOxyfCjZ+kGYTcF67ekMoC9u
R0HFYC4yJ4ZcBrlU3c3Th/V3yRTCCjOLPgWsGEWovhNOolTeB/WCQ5G/DyicTKXd+Yfro7PLY3uI
x14/FZfXQZUXqpi3LzaEsZ15Et8EMHrOaAnGxx820RYwV/Kr4z00/O6fI80aoS+xUbtDM/0YZO50
pFkOhy9iZTSfH1Y8xeZuceQqKKgn7CPRshRQ5FD7fYfr2uMPY0cTbyEDPC8iaryOIOGIJjKej5Xs
jyyuF1HFNwLeI/qrMfRXtU+oBK9TxgB2QCLf6lKT/nOCoge8btAcGH90TkS9dD7G6UvL3ti9Pv+g
9Qm1WBE+rvqp9ulPqDB2wgJt7B9RjRpC0TNVlTZqkuE8XCoM4GO9XGeNQmQ0s+YpLlRlcRHKFbht
3LBwRP0JMgzPowSBR/a9c3ooxr3/TE0YM8BnipnQm/F0UtFPTh84LPsy9UAla+2TTWYjArqNKtfl
wVhcd2i/Bi0OJ8yHbkg8pI+kKO3i5gjc/BgxPe3kRB12wrrPf9xJf0o1QDvzywMZZu6M/UWBmJqp
rHQNm9BmCn7vcYBOOT1Mk4oAgakLz+fuLrIERqtf6KQz5IiQFVXvBODmDfmRCz020StmKn0h49Qw
jYbPcsolkYy48pfXJPhkjoQ8mqszmbDGLLKkdYdsTxj8pi3FBJKTIug4hN5COwLsD3Hfv+Lr0n1W
4oMpUkQL+HAIIFWXzlGDWXuSAz+2CYv/A/aT+q+eAre67WmVCZ58LZ7HMyaCtgvZPMAbHQbff8oZ
w6X7FhzC5LqYYfbZDbzbrtsPnzftqLsm+61WisxeQXtVbx0aqHrpq3/fsR5kdqpzz3fYK+c/Nspn
lmE/UqLp9871vUvxCsBUxhSCa00MnjN6C7tQcvdwnRVNE+JwZ2Oa/ewwY4aZy3uLNz4WNhO64HQu
+2gFQb5l9GkzqbEr8yRpw3v6ao+rQ5H3Tjgv2t2GfoSHkpj5J3uroN+qpDnh5agq5ZNYWs1JL/PB
pxlYvXG2FoJykLSu9r3zPdiopRaXRdVPB6aXgcaSjpbEmcpU+Jj8Gwc/BeGcH+O9lFQQrShODVqp
551devwDV4ZtgNkNQwdHURuf7OKU0zxL9pPI0hrwBUcQlbXdaRbB6VQ0X7avm/KqXVnd4VNO0kqV
J4Nfb1/42ZwQfim/xIolCSyub6DWBROsrnDCUJCmF6O3TzxpZvollXmjvF8L8/bQdte+pE4ZgTox
ri71rZlNClNTvAa8J9yiyx8v2F+9SE/WdFj4pj4ih0DXZBgTRqouDu1Y59maiD4l5uQgl8WIUiiC
RDJiU+qn1K/a3q6IqFJhz+Z5yVnYvrmmUZ9rz3pjIbY5L70CgRkzlUkEN6TlJIn7Q7nbKgupiNKu
hWfxQ1iL/9FXZolO7SFgmlWBdvDirnDXbMuNsaDPOsCSwc8tNsTEHlaxtEVlM4gS/Kcthd2M/DKI
b11g6kKJx+k6aecZgP7yetZeMlm7U0ZFIm8yWjAaZJegHZN1EZyqsb49wLGNfGNglsdtykXg3Giz
twW9RtEADTa+cSWWME6vzA7uOy90yiKZMoN7Hj0fen5QE02SaxB5oLNBye50+uAgUIlEIXKe8W8U
8f08TjHMCj2svwmYlZ08JuK3vLWLKeb9TkMTKomiBDMZ2RePV4P497nNbNZIwYizH6Yc2YP4gUQM
Fzxw2l2TiEX8o1DSWtQLY4Dvm/bCm+0o398XZjvMj6DSULSzdAvvO8h3AeK5n7kraORO6npetRya
TU+Gw7cGT5c94v2uQBeKk9SKzvt9FMDHI5QU317Ak46wcDa0qXKaDnvBox587cB32sMfgNrFkEAw
8HNWPcV8wUwfsT0puSdlJBV69DbpMswu9UEtXu56F8hODca7XSrc+dzvSBxyKGg0Gxc15aFLr43T
QK0D708fmo8Mhld+3p8FFjRTimBh4E+swptd0m2oDtbv0fFxCU7pv+hrGY5Cx20+8CRyoteub64Q
KN/dmAk6z0azZQUWzh3+Jmwg69hXmnp/IFRr6gw2vBuYp4oCozsW8EhnGrY/jYPk87SY6yVzDQlW
yGmCfVCWeM8sN1fqc8RyZm2Hw1n//Oj8J9zUeg4wQzTEUJTHSa3dODiJdSSavvVfAsjSrfVpb0QM
aipjDHaydRFi/wLDDDtsB2MWWMx2pjhcjr5ZCYnsXiDlPNDLG6i3XijzyW+GYFYRtehey/EcPMQS
OMUYq4D3LcMKKAeGICcj2dbVZr3x3FGPrcioFWZ056Myh7RxOiZT7dMr5qai/J1Gw3uuBaVBcwpS
A81sj9xSPYCvJSvtLuEmI5Hx1dY4oloj/1yOpeQ14wr/Fcda4w02uynwpycDBcxfMh4X/URg6dNb
RFhqy6HONLDsvGJ77kqmFXKbFpR9gVpRX9HCoSNYS7BC5Q/bMcV2AzDxK/MQTodz0uVXxxWwreJW
EwilXOVMRvD+xKBpsUVCHBKoUdFqaQEfxP/Wo7X5Mj9+5OCE6QQ7fLPG5l4wO9UfSTZgJNhzv0VP
I+3tCzfDxwgB3g0wO78qSCN7z56ctr9k1B5IaddluQRmcD0iJNaLfrQNHKK1+sWmvOU5qR4GYQY9
UXytBzRY8SoMyUaNjCdC1vg6gZ5Mmf2CWrtn0lGnPvTqdv4GhV2e/VYm89sWCCFmjoTPYtu7d6ox
gP/FoWTlLsKYequx1X9mvcdvZ7xZQTBs7MVjeVnFDFLJUbX1xHojjn+69XXJF8/VvJnx2G26um0C
LwHUO6JwWlnNJQuYK87LLxtyIu+OOMMbZznSxAKgvcSD1a9SqoJBK58JOLmv5C00y2bGVURDt2fI
dZVDtNU7A09MEyyKu1qPnmfhwdpQpkrWuSh+6261uT+gtCTrKcxUoo69/I6r+6jsP1sIIgKgpi3q
TdALKg1RHMSndB0LVA0SS8xDbQHJOhWhF33RXRRpGtKUlCFQEY/35WeOBuHCmPNc3cdE4GN2tuuM
TcUR3a5kizC/QkXJSPtnqjiIKZ2NYXaQXGlySmuBb8jD/FJaEjy+3uK28JvDS9x4hnxOC/K4GsrW
FOF62BekMb9J3WqdGM+mLLOtNa18bSkf+dmjz8ReT2W7xd3tHgFoV0wOLboctuBnk/ISVIKO+ytQ
TzwdU3eRG0LOuLBy2n5SASGT/f4dDHvMrDrWdWRe0JwA5xFucj2aCrvCFz50nwn9Ba63so0gYcY1
nAY6XdwvECgEyToScTJTRbB+PbnaTWriheEiWBUPF+3DXFh40d+EsLSRMbhTBQyU0WE0lNRnhvSf
oKh0VyJmZun5TscSZbu/ZwDeTSnoRIKJse2cgVhm6N/mA1za6zqS1Wnj2a7LT2oqqUgoEot5szit
h64DgzyvB8RMg9WaaGQ/4aibsRsjg1HYAWLuA+5pyOVU0P/NGpY5iYBGqBxWtQboQOfTbVfjf6e+
1tBpGiniNC0JGY53vBLEvFxdrFHJjoAjumQUDn1duCQzn++eySux4y3KY3ds6VdmN9kD2gJoU9Rq
W7J7KFtO6oX1NGS5OuiaiwAS3hM/adagEmK7J3fyKVEqhwzjQMcMT4K7Vicnkx+ggFXa/DaoblNq
9W1vsBYM7MTjRFrbDT1zt8I+pk4oqPek3lA7Vu2rL1W3wDl+DkVcgvgoMisVxn0WEC62BYbiTTtC
UJgRc9lIA30V1rIFEAsyqk/1kYzpOGP/HuhjB1gODgzms1j878wlNuBgcbj9LtmqNQJIutUBvh2Q
o7Lhj6TD7D67Ep4Hmypy15CEBY/qj1WhOHjp8+kqrX9e5/e9+9axr+9e1Of8KebQlfYeyxp+3GQX
3wLEmxJlBMzUm5OvhjWzgpBK4HCPxJ7F8n/1l74bsDcfTtwtSb8rtDTIqpsNY1IrwzyZvZzJz8Iu
f9pXaDtHnfG/q+xKzrEAC26oeBPYCcaLm6ZET+8IllNglAmzjAn/i2mPZHyFGhmLBmt7p8GkXECw
iBgduXsDzoWrybJauyHZHrvd8ULeLILU9yGQP4XYcZyR7UFAFrz6HijLlNcUYjYUCTHQwFsJjbcz
iFkFI7YCBykvy7kXVd5O7qFTg+8ic+1JHWFWBdq5oSw5IqhfmOT2oFcn8yjMYKQ+To0XYwoRyRNz
w7tXVVYLUL65kMApnAGbwW8JoiJNMayNW6cVl23tcYcd40tiDxFcMbUlOAZnp+rypTowwrm986pT
z03BYH2TPz1v8TTY3n8mD8Im3Ab759OsvcRjn2ITrgxCesl7lW5yl15ihRHs8iflkJqthbRHLiKj
mNbfrF33EQAunw2REE1AWm+gTqogcCNOZaDHT4RULut9d8HJ7AE7JxTPqNCkDG/+o9RzgpeWmYS4
5/rFfohPa3fCUHuar+BV78vnCKWTOb/+FqZ4idK8P+xTJ8biHA/BUCBD7gSOnLmh9BqjBDvtkoh1
8w1xZmIXjKRONLjaNEw/fetJpUPjnirlKfdaKjGeXvZ2XQPU6M+HksodhM84UZmUjBUooPsWRPU+
aD479vwNpIYF7SwglNkaYYBb47OUA2wxg/3EsSJygZcH6c8hbdKsRx/3RjOMeu8jt2bjthKyADxa
nIppdo1eJ07A+yXwCD5uJ/g/47uOTeygQ/UBYNY/x27o6WEj0px2PG4zYCdt1lBjbcoM11MBFTvZ
v9IUBonQ7Jh7+zx32uKdfbZun1CDid/IA4y7UBdRJsm0fs97DDORBSumf4lfTBkoGkoW4f8c+EQg
39N073/rG/trxtd/Xcf7sP1dfJbvGkrlhFF3jo9lVpiBdPGAvuygBHpCwFwfHqrrTCsUVuvUrFAS
SlyP39h5Ef4o7UAwGq0fyP1A/NKE2wx1XphctNY/qiym8aIcIjOvXszoX5sKHeD9x+PcOR86cRV/
zLnl4nc4k+2pFZx2haIbag5k6ju88XoI1WQCoGJRs0teGvBfBlZWGizcy9Pbv8R3Qzrz4rAE0c+X
t03o76Kks+tS608ap3ZGAQRGbsQHqwDEvWuqSXm9+FiqmC8L3G6NWSRhcwGpdvJ0NonSO3j2gDjV
I/+rA8jhrh6aJWRIetBWdOR/WZPzsclCiYSoKuU6x8EZcjbIHWxv2PM7/QlytPwpJzqZ+nNqRO8Y
x9lLTkyYeoFgjGF5GtEKn0Jhpdz7a2sZI+dQ8VMIDGZ463zggdPiRiHiKlL3qknbChejM2F7OHOs
1ltuXosv+7wyiG3j1Qp+5KP01RSTU7SRPsvEcdIGgifqxqjy2dKERE3gpesZ5xKlh1J1kUjguRLg
e6EAW/stNituxR1dXx9BnH0+KqXH0e7aEYVi3BjiBrS9VEruQc+uk14re5qi/pgn1JP6IW2hGDno
S/7Se7otlKifIPpqowJDU1SN3Gl9kHtMbz67RIdwWj3NigFjASF2/oc86e1SlBvrD7WyAmYkKAo/
joAQ7efsUZgxSyXwlCARw60NkzGkytZBuLE9RCv7eAjrXFmk5612URqRw1xTvr3z4Faj5BBl/66C
6M0vMK/5D1KSxkHbVD0LeEOFVD5ba5SbWzBZYxiC4tn6JIhnaZIHAZRTP3QzAqz/HdStIZk5Ggz8
UDSiGj4uB6nQIAjuBIXHDKVuPtX4xqPbRktlvmjsy8KI1YMdp1jDld1wzT2e/a6xs6cqHjybhfy4
bM3d+GTCRiFCQeqQYU+DHaf4yTvHnz/YCUPk0Ew2ou3tf2XeLV+wfrI+5/Y/mkM6cS5KJ5yEc5DP
LaP7syPGOtndbBKley8ZaQzeJrAK4MhoynGovOMtmIDynIjS4n9Q65868ml8xLuSD/FHMYjG4cr/
5Dxq6NlsYPTJZIIp3GXWoxws7CmHOQ4iJfMXxrknqgpDro3wwijJg3E83VLxEa8OMySWeLhhrnaC
mfKj1TmQe0XjIX/jD3RM5iLDd4MyFWtQlNjxwUVWqTO7L6a3E/juTRDqPvR6IKdbhNr8TOdj2scI
DzbQ/ilehJCFAc9JBJS11nkvXWgp8ltmnVC6Nkx9fWti6eNFI/I0QS5FOoIysWSMArtJNRwFE+cw
OYMOAlwDgcCcXJzSjtOQbI8wY1m+gYEEKcH/e/LjPD0IlK6M0vtHmaS/GATb2qskbSATlhiXhK8J
6td+MhaLW/RXQIcUDuMVHP3LMlNn7b7iN5OUx18cGeZ2i0UySW5zEdxiSh12x87XJh4rE9Ezdh1+
sUcCJgiVvyKncFNxNC6VZFY8CXK6BeL4SjuycoQqQ+jnBwk0snhFn26KW6kI/UoQGgh9iVaNEMEK
51N36uZsZg0u2QHQgdZIeW5TmuP+q7/rTzDTzjnQnRvf6e5Fntluq/dxyiMVfM2EF3cilFU9lU8l
ueqdJflJ7fzwVqXtSnDjAW61PoVRUWPuH9UNSMpYaCW6WfvxPRBKUEZ7clXkxXCZ3LxdtSP/OQRh
OvyjPkDYzHFeUz5ZdJ1Ipvw+s/oDB0m2l8HXjz3yqFEW8DTa22rDt3WXqa8Cq06OcscEqk0vRFPP
IwLLfx942EaSCWu01cHaldrVP6F5lwI4zQGecdTjmy7NZVKMgiucvv5AwrjUyi5QxLix9LiLdF1P
Wio9cJbot7usDOuGWlAxqyHa0myg5slHgYxwD7owmaKBjrktDlTiz/lKwi0FfHiDUcO5QGAniGKo
HZ83klyGg9HlArV0IfXkKHPauFnX8AgHkHvlpw4F+3EGG6Mv7WxGrtUaW8H1WPOfLyQIH1P1fhUD
I7ey8haR4oh/B436+dtSLaLsJEVw0J4TZwSioifqvgBeDs88GmviMxBYxL1P/9jDaZINRF2g/qRA
9nSNHgAFDhlxcGpLG/PibJVT5JYMqd6/XJ217AFOW6Hjv9fMqyULPYMHx7CYF4Aye3HBBjHKdiY7
YszvbnxupLTtFVZmbxuqkHWXw+UY++5UVGc14nEETvGKB6/ilUBnBZc5izlZCPNwTHFawPz9KlzR
ZlFeDnMFGUANbZlfHrPtZcuwiK97ic22qmX8VVEi39vj7LJQWOJRjr8eobjFWzWuHJnqU59H8daX
+U0ChkmaU+REJ6chRpNSuMxxh5pTefeCSjhCwZhzN3o5DoHaS1pJ/lroAVG3kHo5fB5lssM8YwJc
JLb3LXjEtZUkDZpJ5LMnsk4BnguN81jrK98Nn/6PrZfjIlm4kS7reHSyobskdTtLHWyHrhdjYXgu
v4+wTM0NKzhOOGPJmuUCcWEh7jjx/yMh4IN1vB+U27Cmvhw4GLyww/z/nhWeQzqATgtFSrXq2vZ5
nV4guVNXaDrcU3I3EbUouSl1mbnkKuCvHyBzLyNBiPHuab06xpjLH4kTy0o7xjdmg53p0e2uAsFR
zh8lKYva2mJ3K+TI2VbIVTXalenpXN/CoLNXU5mhoUmazD6aHXt63Sh/Ns+IC9yR4UsUUFqHYPWa
bk6uTd46//xW2SIMg+gPhS3G/BvuwF/3IfvF4Rao6p7HOsz4CkMB7IbcDNIHrn7xH9AedlMvwoWY
oV74hn2b3bSloTfJXyc5uoP1v/MOcBKpcVejHbABUVA34gAuW2kvGiZ24yX+NbLevB1JRTj9wSTY
oItfTn8Gdik/9p0rZxl/5Svb4qstY4V6hVqe/R2qCDo2HTN3vQ2f3Er8u3+/Po5Q8Y73PpzGnntc
bAMbZxBHl1euvffYvQCA7+sUKq+3sErk3JNHIWoz8Ks4iBdk4gn33cRYn73WLW9+6DxTx8A7rPMs
AjtxZ7sNl+Ydrsmh1a6A/ICSvgI/KPlXtu8C4DvZD24D6+OT8stYFfeMVaMeQz8BBQT6idHHmY1t
0kRDj8PtXxt5E4VrbQC93W2D7guR4FcVh9vGqoPaA2NhweSMcmvgq2ZLdDBX4eBoevfu0tIEIz84
42XZ07OXJuA3rZZeroVEq3D9Y8wmJqSxXPLOC2n9oCmppmxm1T2gFKvYJISWLip9M+PmK0nwEyzG
wQLxW8xRuBVDzdBxcCyBLvwqPd3FUDdbhvYyrlqONkZJsc3nft80Qsjmtnx6HWO3PgsHzDQp1nv+
oms/G84DrDfZkSgWoLeEULCy7DbnaFv02l29OWaqHtJnPPx50039jWPAGDl823spdR3gfr5pPnBb
HjZOnqeXfR4VAHMdWpXIkrKvVcAjChrprdWZ0RwdpEnxktFSfdK3t+FRsjAAEZuXabnqF9vUOqxu
KMivkFYWnf1E4A2Li1VnpGvlIopBErWN362/xAIA+Nr37+UqQElocDVmuDdOsMasEAXVVf+PcDX0
kryFoQLLy7LhNhb5gyAj1/Clm+pN8SHHsaFN9ChSon+fbHe2aI/6NrgKVpkoeELGa2h/L0fvCazR
iMsTSxs6ZlDV76edINQDdUJe2dOTPdttkYrboVJbRApe819zPIYuoFzmR9MWv6HTlmjOVcapfG/O
p3f9UONeNAuGGuteF+HabWHbm7/W8JUdyHjDG73q7u2VcLtFUCcjuX77PT7stYmWt2gtKhYTGcCL
gPQwPUxYu4TfjYe7aW/YkKhT73TBrQZ7p98DauRIw6LBeEkUlLMKnZD1/EXU2ckt0998cUGY3htw
BhP3l2Ei0OpNuVhqyk2JfUKlmQKf8S0iLSqK82+XRJpD3Aej8nrZJ4wHX79WebSBcjv52wuGZAoK
/0781nLKCjnB6txLzbeQu7ykfCmQhDiPzGwypExLkkyqEuKOgx3Jqj0PVRJld6X79IB5F8GXgbIn
J0zcsq14NvTWAAtJMTmdWhrPoGZJ1JFGTOPxwEoyX1TOxITnmkk5jrxPU69WzUHfeul6ccm3v7IP
nhVR4jayY1mDQx0Tuy+Wc4QwjvQOmC9EYtLAOO4qXvpNJP/8QNaMJFGTtKfPGmVLlgaKXHY3w/Pn
aXzh9gRtVJbws5ABxSIY6KQm8LlYiKkuVnpaXmrC0txB/UejaQ0bxh/GM2d/FD55HsTZ9Ftf0pkP
Q4PL9+LGBMFmq17Rb8Yp1bzS2DT2NSwV8mmVQJaeKvxcIQ3+6Dhe+Kfzyg+wqUz2eW5+qjIhcZIF
LjPzKQfZ+0UoJu0JtILv12pZKMz6vuBUFwE2LEZkTd55jh0OiE7LOgR+/7SxZkETZp3KITLmPgdm
w4jXV7DH6omHWrTGbPsNFMRtf6B8vhi0DMROAJte6WjBepUHejxf6NdAfzxJPZvH7MDsQRo2pKts
sjpWdzaXVt6yr+jER2u6zOZvf3lkwdZ3YjbrcbxTKg7asvh2b9G3CWnLCY+CdZzA3GvYo0GWZPmi
CsEidR5K3/azo2s2ylYAIGrdKjPCoLzadyLuCwcI4bcLvdErNgcbJiIO+iOlsLvproLLC2Cpurcd
315BmHMYQhUyjIFSwiJGwYwZ5KuDuWATxqARrQbyraBvTWtDrMbwX/h108nsp1FDGzv73VyYRyMt
rdGCVPUY+ZyV8EzBJ23rvZ6wop6B3NQuefHmI4sKeM8DfRun2eIIFypY5ffvOw76bZlA7Ez+AAVg
zO0p9wpTVWETDdESxMEXF6J4o4GL4LLjq4udhwXZf+Gpooomo4O4upz1m3ZH9TuiGvHJkcIH/LrI
kaqUS4i5y2ib2ynyNWrOME58tuPNdPFoHuDHYPHSEh+ZM22QisOFpZXlwE/pZld80PUoS+WjWknm
sLo+gfs9N9SuD4EsVEA1acBS9gbNFnhJFLXRNyD8DQxm4CjWsgAmKKdpBGCAQrV9BUQCl6xAKBvg
G8vg4HS2Uu6qd83NeBIw9rlznqDHXlyfCG/MmWh0ReqzCmC7Kf6MRbvVP6rkdHmbv9ZBGc+h5vTl
HOFpIJ6nhbr9bSzhi8WWn0NuEfua4P8EQ6O8WWM1HU8Su3eF+USk1D84imRNzg8p6hl8IUbIgCd/
HwhmYzIl5ccK8rLW2/npnpWRn/mK0uDqfwXzczaLMNr3h/Onh9yM89UhqMWbncC/tw2x2TE7kJG0
xDwVY9HhmuSa68pRuSVgu7/SCAz1wflgqBLuRuMOs+ZOpoN7jXYA5Md465qZ5TwHPJK9pBX5e0hT
xpkAxlJcfveCZOQc942zCHA6p7/tUlnJxN2WfwHdwrBVgjyXLi7Wl3x7OJeoTl1JCmlrcINmk02p
3p+njuOd0i6n1aOV6G1LPrxFNwKfW2gY/fHSyb5VwEVVcdRG8vH3h9UHMZvxBDwQLTuBmvfrcRxE
TBEbNDTM+dbbEQqOCAOfid7n1vET/YWcg2qz8L1TIs99rwkN1gfTGCUla3XBdxiV6cPqzb9TC11P
lCQZ7KnnJG0PUw/oJPmrzRfvawoAAV+65iBBEcU9Ku1uwwb3juJADmjxuEeC9QCdkMV1rVGHVdOJ
epJg9ODDBHFF1xrCsR0oFxzYZkON3EKUNH6nURtO/uJEKojDdMoNYtMVVjmxV+MZqUl7HYxFoTlM
kjXRHUrdyHYgdh3ya4ZFJOxJTfRLp5TpiHKhiRJz2iZ2egn6vrMQAj3lZLinZoutSHNgATK/I9bW
Yq0hryCg1cagr4Ak59sxfHv8yTIa7HPTPXjNR5boFPFNpEWdiWVPJ7aRXYjsbnpkxQpvJ0ci8VGh
e53t0bSmh2vk4V9VGPtSnPP1nZx4uIRzLBNbZKSZ2dYynxHKSlXXq2wKdt4t9QAP1ZohACdYOA2s
1GQkIFpdaM0BtS/34OSMiByJ0YtOmCjKqmh/32HcCm7ZwIN4IFxhp52b+klow8EP/pg/5eBVjDin
J7EzyNRxE0ecvgHydonWwy2vTv+1R/dD8WeOc/PmSEt6PV7u94MN5eUpdRPTuwjBWjy2xsYzWRvx
VcH/Fe/qAWQK/+5xljQgdDbQ7mIORIMwYaoRAVeII880uq7yxv1BzYznga2CCLnpcBCpwlsbB/0e
bIcUZE86fWs2JvmDP6l7nm4qcTjTGZksqyMahCAJ1xoro2PuSKT3+nWncliKJsOOUYJ45HEpva5y
sWQEN7ykemHizKjR6QQy6CVctiTOrM2gLL2ul91lUY79yzNPWJc5W97cMWEpLvG1lzSGdXJpEQHY
rleB3ThkIVhuQiZ/1lhvZCLpMh4dnMlz/LUbJpk7GRCeqJ8WrS9WRuTZqstQQSGDWqhBXXvveQN/
NuMKD7mECe4qXtX1+NMrXNiM4sAVjcjPmV/ikfVvunoRGHpY64eZIIgt62HUwURC25XHy3gAy7hl
Ih5BZuPPpjzcKhHfTn6Ts8Irds0B/yoZJNDGHGPyiTCw2PgGoyCXGlFjL5vy/HIDXvJ2U1CM5Zjk
wsFq3VjPqGhZOi323VGfe5XVAtwza0BMnYhVT7y7R0wr2R3GkXV2R5uuHe1eKFl8CzGVJkmh0HTc
R4Z2LXNSW4RWUQplMFKp8T7S1EqHqW/qc7K/GrZ1dZ4zUhsGdPME6Oo2BJuj83XAIN8az8xcyrh9
+SKSQhAoYUNMfpmBGA1tCGWSXzCk9EjdlTQXbulERu9dAyQWut4C4OgVpfuDAPJoXnxO9tA0dX0r
splm3DmDmHkhUkQ3vGCQgSA7p1K+RFNZiPRW2/Jp4yQIRlbd94rUFnrn/HA4Nsvw1HywpSPe38YS
TSFlhsD2TibfOQ5iC71CdavuOGniM2kYWahimtD8ca6GyrWyRWj3q++v+53VYd8MehJHvzqAQZgW
aAgkUoUjvEYbg673vSVX0nIMQNGvlAb3zT2wov8E/UjttpbHUSIGxRoc8aXTXiC5S/uVQQHa61zt
yEPfMf3EH/yQde+rZlMWf9/Y2EW1dErMpVThSdKK+xp7LGgeM4g5YhKgFpuPHzMlIwB4f/sbh1+b
voOipnLBjc4HLoOD27C7bEuHTw9hohCP1QpqyEHIidU9ISnAMa5g+Pzt87nTOD5mOWZ9QNYePumi
7EmlTkLlebKNkQUFLgEfHwpn1aN1o54MY+0qbG/hhhB+7f4B5wJuJKs3zjDwsy6xbwJmO/5wOOAs
3G2le4WQbTSpbdRfe8kTlUxYUU5nr8xSSq1BOqnHFTAy9t1UJdzkyPj/8w4pJg8ZQjfReyi/Zz6D
YsrTOR3JXdo1uYYg7Gw+OyBdDuzhfku4jeg3Daonv1cXbJBv9WGT2PQd3n8XjTmjim+u45edeM8e
2M4PdECurp202mknI9StM4klLSeu2QeyI75EsZ+/3WXfCuMEGKcnsgKQNKos40I+UW/2+13N+i3K
9WhHzEtng/1sNlhJi89Pu+AhL4nlOzQGxKXLPskAiPckLnsaryHfE4mjm+VSjOtT+ieF9KKfpQ9P
Aro4fUsU0Y/T0hTvFhR7xEhq2PDLNyTINOsWrhjUyYDRcFdbw5/Cm/gEItLJE8CvzEsApVz3ZhQz
FXAXer/QkvHX9iKYJnr0FW0/3fGTyOt8FR6RRugEWIbUREDKT555EapYw04L/7BCgKggRVdxOPOs
VCfaxhQWs8b5gnpcy3n+D8C5rL7oOQlJsQPlOi69pwiCCjRd2TQwHXy43aTf+K1iI1WdDGiGZxBk
PCKv4u/a+fX/5k6dWNhvVWm7n6Vo3an7XoDcQv47uhAR9CP05J/JsBfa7PopwramZhFhknYI+HE5
V4X5ue+/EKIneSxr1E+qbnBt1vVoVketscsTkxm+HzsCSSmBVZ72KGJs7YMqbueiOR8WUeiBTAy0
YZkwtuefI51SjFjyV6T/Eup5CxyIcDUUZ7S4gJBaXzMKGNsRdXNmRIsITvCGyRI/8w2KESPFOoeq
vf8Z4air2iyuqJRGFgo0/7C3j3X9TVtXeMNjKzXLp/pU9ys+3Bp3t8VeDdRL+fPwtHIVy6pxkdtO
hS3duHTLccxEoHK41vanMHeRSd2iqllt5djueS7HRbK2ahFFuUxQ7CcDSiB4dYYCT6TOs1Uw9+nB
jWo8joYecIHJHz66eYD3FI18Cu+5Ss1jEvu+HEVL7XQxa1XRxu/PAudYuknyTz0f8QqEKlxU9h18
xNdkAqjOz43tGLhQwGTZWc/USWxF+itUwaTl3KwUisERDXwi351Y4QqRN6oD8P24Uxu9TYOs32IX
6ZpGM3345B7kqTArNvzugqAe5rruKN73lwSoKgOm59E6T2xHmG3W06eCMWof7Hns2MeVt9xqlJQ5
OQMXF0MSHhCpeaIcXaMVwyF5uC9iOQu9Nn1gO2BjrVFuwqaneFs/Ly1TZ3M4tkex+8LyfGkQ9nhN
OfE5zOf9BWsoNfioQTWECrLwCC4Qf1n0g6k10BD8Ij4f8DXTp2BWuuwhdI9Msm075v6Tkw04jblA
9tUCoHdEUAwVq1P4Wkdjxd6Wn8jYknzIqjDdbYFw9TQt3FzbOOXfgdPJK1QLvTAprhIq7Pn54lTS
13ym49CUDy6Ld4lw2jAQIJp8KMVzzKGUkJl4w9YR2JthhInVzT6sAGnPMldAngFAPwr0wmXncP2x
Jzr6akT/ALuv3D5366+jluCJOMdFhh4wht44iG+MY6E8DYkNdTY+4rEPh2xCCOtJrj/A/eGHq/+O
p6SPZU5wR8FSle5mrTVwaWK5oCNYzRYnp7A7XdIe6Cit4iVDp2JwFPN49vRZ2xy926yi0ymPjwco
luoU2gqUA0OVMYWBhTPGyQdN9tkywGJBT0ZDl1Z18gBAuA2i1wrGdqLdPU20nW9qv0LsLNgDE1Np
5IUZjKMPUD52S7NKs+dvugQHNqBLnL+stnFWVSLaKx4q+fp+9Px/cddMq9GSNkWJ+sm7lXzZRc+2
DptWZCKjqYsCejYbW0+S/6BXA/Zcv6z5U1cuY2SBIKFK5kybZI2fjNPxbM7om1fruGjYbxffRJLZ
NEU2iEJUjR1wWw0dKGiWBcsAg5c/ssfEnxJmiWGtI5fYP+SI579/JBpGhiic+sQHNA+k1tWK/DLx
xJH74pwBq5+YO6ktPhQTheAa+XNkUMEw7TiX5FpdDpiV9vEQAWReaYkEFiBbWBxENlfwZczn9k7D
XtotpewIvX8rzZFTiWVJn6djhKT7XSWyYAKrmsTC+zi4fycCub14K+ST4y4QaSa5trGJm4DKEjlf
ejuq3u1dQHRo+EPB5P6fe4dyQz40OwLR28mcMrdDGp9mKjUO9y+bH1OMkI06ojMJPVv2YFWPsZ+R
HGsVCytHqCPD/XKea5mjgDkL5x9nYJx+AYcLfcGmgcjs3CjlS7i9uEA7iijgdTbBq5NXSRFPnDIL
Pq1DhX9f1IbogxlNfPkpiJgPJFyaIcQkfknfRl9MzvETB67MqaM8eGOsJF0vODU/VeuwC98NIzAQ
hH9fij3WTuUViHGGmCqnFPMF/0fGRxDbDQlYmMCkQX4Til0g/w2mt/zo7FbFmUSyZymvDzYV6+hM
28agedjmLbWBDEVRSZ+UvVNtNVTnIR65REHjziZKf7clisR3b7CVPrmzkUKoLcss2rm2DFpYJrbL
uf6WoCUXgOw2NEl9Y4jxWW4IbQnkFSHiDt1FspCIMMgYU6w7248+CkbTdoXf5kMig3/no/6KDF3x
VJLJjAIV9WnTUGAE3BGybbqvj2brl07KrNQ/5LFf7EzOKDi0IzxS1YsKXaqMbB0MzhyxDvR3M/oJ
X8Vp9ttaf5FxpvBmPq81yxDaCKi9EAZOIVCYb/+MxB3Q2tnSu6b5b5g8uO6SR0M9VJDlqH9tlhvc
EZJJ+yqajC/z9YLnmxz2yq2hjTyEKRxJDP9nzZnfduU4E4zrjDNNEHc21utGtU/lQ0/8C6waG2w2
2KYsRpm8k/rQzLdcG9nUXxzrugvYPiOh1PD0D4k6DEOif2TPOEV+jjLk9VqUtgE7wBlL6+k8o6kX
2zxKaafJwf/G1iOml73Z1i20S3K6xrjrPbGRqFoSGTF1yDrfIieTANYmLoftKwmVrFIARVq7GzbG
z1Vt71TVFzqhG5F7xafJg+OphdrrD6saDZMpcvHBH9f3jvuj79soP3ptgQ3WwuZyGz7VRG+SUFjR
bQVtCeOUSJ3dNALpS9hupZvMF6vgD+pEQKVduW2AFQ6UItL/Kvoh9qfbtaos9KNZpdify0GO515D
HXABeqYXoDXu8ARx1K2FOqVp33Vx9OLrJiIVTtu90Y1SFVtk48To4ZJZhQDLJEeGrzEwX8qRcfEP
DNaymHOI7sJv7S8iZNrJLgCMnaxzI60Q/ussXvoLMcgZUW2HtixOiI+RBwkoe6zEZhv9EPp41FF2
7UlKsPVWXJ/bE8Zu6jBaAhlNh/3Pv5iwkyuDk92O6ODVVbqLVadqEdx6B+C2wrnSp24sLx5NRjK9
7CJ0ujVs7YV6jD7BV73QWvNArbd7T9Z7O40krLV9pJa9qYR56cer141vK/Ut3xc7toQOgeSOM+a1
vMPXDsCh/QlB6bV3qihD3jEu0lSLcQV1IWxgzC4R/RnQueqO+MmmdnJY0jCA1Ihx75k1LHLrP/5p
soxZnb7/fSb9TGbm+nxgvzTGzfuqpfaIk9xzvaOfXJZQusQlW3hcmyyws84xXeSWWjZer4qSwyBa
1ANuzto/sSwA3mlu4ftP6+GzAX/oOvPZKpAyOHqwa7s3zEYtr6BKU7ARR4QTMSpVvM90w+XKvLWU
Qh1nnBnkR7Q67SRGSc05Iy91HLb3r6SOaYG9/i8ZWKNZTB1YsclhsbrC3LppplWkwtcIuGNpmNne
7c21TvdhuKG9FolLpqO1B6/L+zsHfoykpz99xzbFp6O8/hD4FXbY4GJbSN1EyHlLbbs/CFVtPYz1
LorYvbTax04nFwnDU/w88TVGjhHJ7Ij5hN4Q2hyMzTfwyyGdnZ80X76fpyJ/7lr0Zp8dF04TKt8A
YExqhsKcJe4lBxt9qYftPHUJwf8NBDeHQPgKXfsXnMQuxnhGrNgxsZRyGau50HS6LX+B/y8EpZQk
nyzo4oOGoHncJ1k3VumudEDzaqd9hMSjFNE079NhRW+eJoJ85JK5EjdBUPer/UL4fAJDeiiDA19E
Url1mx2eQ6xqH7wbQZ8eEAVxRgCDK6lDbbpoZo3xGvVu2aG62dnA7k3I9msapKWzUtvlYVaBhbrn
dx3WRgavDBPfpWGVESN6q2WLbkFvv/3kuTKqxyRerwelUTz3AVFioKWS2LITSB9vLTylKPBcWjJE
yAzM7ZWwL4Bd0vHwrhYQ1vcpd6JvE+hroQ/bQ4rHCLTiblN4LGjmltT6T/ZBb56+8FHBo/wBHP4P
hv5Vvmf80a9klxfrLIAodXoqDTDlH6fPDVnmSfhH1Lp0sicirCZWB7SuQWSF1t/n2brC07Ec0v8T
0cqqIdB2QULuESbJyIr0IRlCSLM/3aY3xiSzSgHJ3OXK/FbI+MBcX/U21vmayvzeDlnR7/01+kfI
34G1yl7yXNWV/XX8gsWjLW1dKOKXjXlC1GUyF0og/ImgFKSKxj/hIzOhb5SbDqFolZ7I+9BbF6l4
vBbNHOhdF6YHStzEs3zQyl6kIHDvyTwMEZGZzLRqFeVuY9s5COX0Ee1sBRX/Em3kB+qPlLQRe376
hmq+myyQDpe6g7groU28oMoB2vmn6PEdedE1+dIyjQ1D1KIqJHiJHkl5rB/dpNesfAOuE1bqSn3l
faLriuOg0xHAPAD6pEq3+MkyhdPHYW89Kq7SKmXwHzJ0eiX3I+ZG2bibyTxpEPzg3FX9TharsHyG
i/KQ4yg5WT+i3yWzNmpnkISF75UJQnsxhHWGmVH1srAj5WHiW9HzTC6DAl68CXuvkQWgDWZ2gdGI
Y8gvKfM+GSwt3r324xhaI2mGzSScLmvDJ9KebGKOupn3KdeoZ9NX1JFyx+AQYTScDK0aG+6iE1D8
sC4/9RyocpErCbGIld+TkQ1VM222eTENtlSALn0u7/qhdnaOGBbNDFraaYEIbuAfaqbJRa2XwgN3
+UqRTwCt4jidtqJYq6JAKxwLQbioWVFef5tZaxyBfoa6mD6HCJFPUlVbMLMB9VEwEsiQKcPo/UpJ
Pb1I8DTWpAgILKPTyRd7CR+CoKlGvLudSZhOwlNwQBIoFilYGWOjVWPsoVODr9o/GWon+z1o5Vrb
rT9CYlcVjhdPTMTRexe4m0HM4misjNK84EGR4TDcnjfjSjs5zGKqIFDYj39gIhm2xNqO58WxtHZH
pqCxAf5cXlbHUosd3Dh7cNqGGo2xv2uPGYM86z3JtANBG9xWrH5CR1dCpLtzF7JBln3nNHpHYor+
LpUI57Om4fjoOD0QJubC1Vnkjv0rCM67fxe9GoJsPHa5eWBUFIVYiLlseu3abkekUc5jBgrEUsJI
0oXBM3GtqvfEZ9XhIes2PSPjzgHqWEAU7i7CRu8eXhK63A+VBKHW1wPBO4D1g5E8goPypQ+SIIbz
aLXfHG75NqJM/xYIFRI/hmhFCaUL9PP4lhDqE9yJZDRRzDYzvMQ9gLc8HUfea05qBBz8IG1Mza5r
EAktp6SIsF6Ej5izJcwmeysH6xJ2Wq10josHW3QvRPwOwzAraBP8ERBjd74fFna2DLAWlv4JQ0i1
vuRUjSE24JMNvAAvz8SvB3EpCqTZ9D9TcYzFbgXBJk6WqLLbeiEKv7YL9LjrbTjVKiTWeljTlncq
esMvohnISuGABowmyBk/esInZzjQtkLTfLbt+uhEtciOj6Y7NMd8/hWy1VB8yYYxU9kYGj9gyINW
FDA5ZDI1fONpMMrDy4/dnLiT6jCfoM1KavI1KEBg8TrT2jWW2P+sk4fPU1KLZCNJ2+lsvwb8oQfO
KtPl2+Sp0L3yeauqj2zGSjvAj9bSgiBIe4bRsgLcjh80J3u+cEV2lqVjO0zArUFC3olXNknRXNk6
CuzWU6XvS650SrxV0Cjg+IW6xoCZ8QIlGawUeZRqzS1EUcaHHsNXOv3Z+Kr5WAW6kZXrEXqsr9Tk
nDXfHrit1W412st814X1E61vQ71RKmDXNVnETOA27D6b36zObiBSJ60rWTw+XJZ26q06DhotP+h1
UjupBUbO6vBPmgwq91Ef9mnnqfG9We2mHc2GNUceHvjZmfQjW6vWyN7612hb1g0bIpgLgryAnlEY
AZ3stQFGtuPv6Jhp1m9X1jPjnwfjLSWDOJkDioBZ7vUZ8hsLy7UeuoeGNtlMY1017M8RtIxBs9XK
ZrlBLtE4dmlbJtsYdxe/eaWIm0mQYchAu7BugOyeKFAuG7+mNlawXpxnMIfQsRGa1cELCsdgJl+W
G9oBChH3fSWCSsfKnMxNai158gWlqZtA76IvfI2uzSOkQ7V7N5SsXAo6dnxydAMp8UQaJkMxL5hd
46sfoFHpuMB7B5NHNtX+j0YAV/zomD4Uld6QT3kraluiz5mnTuaGlREZOCyNSffdJNlgftesFhHr
x6vd0iL6hPxEcrqILO8kU1LCn7pXdckmiXvDoxagOEGPwtAXKmZwR+XipNI09V2j1DnUMSsN5Dwc
f96qmiW9ENo1HKAF725L9N8QdDOGJZ3no1rb3T+3+3bafsLlXA1Q4680qOW4eEB8t6TSPJfEvwZ1
JtdoqgJPg886qqZQK/0WCJEBpfiZJLlg38xZXU6dXQRwyzkkiZP2n8HVubM4eBJk8EaYRVoQVK8B
0rU+MfS74zHNja8Z0UucLRUAHC+Rn64UVLhL0hV/wwMcoM/TrB+fKBIuylPPARAfsk71L77LG+0j
iDBkg/wItzJ/KWFts4YvOuvYhPmTrXlE7FGCp/EWHcSFPx7gdqqyJqIO9sNcQVMjl4AQbVjowN22
2qfZYUs2FdceFf/uTyIeWlhiJU7OCQQy2QYsU6sdEyC+/f812zbdzIUByiTq7miNEEaVvrc++Jjg
JAHKfzOyXR+bvuwgO8FM93nn0jjeyrXkBh+Jnsnl0H7awtwq8/G3/8NC7LmHeek3pErBNbv8l5l5
A4JFbO/45xBGZZJFbRIoMOhoxr0GWvUjbfnnifTJsYuV8aIFBzKihVCj6MiNV97BjoDEHYZ3mUd9
sE8sJkVnbyNrhNYG9Kd47sTJm8EvBcFfHvucKVqlHl/9vjU0LYqgxxOlhtIiOsJ0E7xL9ELuk9jy
alh6LbWwBdMG4ovEuZWAIYWN8qePcgxUQBceFXYq+oIuTq1PYRMWkcp3PMJK56zxF1LXlvVyhdVW
JrYuoHSsp4JWd0WbU3Ni+7NW3BYYFo0lLCDHepFEQt4QU9Ag3bM7LfYk/6QjZO4BBZ3Pmn0Df7Mt
BLlQsb6vA01ZRM9jIjD4ajoEbbMCpo6oPl9XtEWJFg39C3HcmbfvRxgcW8lxFgZJLlWgxyB2ZSGd
Je7SeMFx2IsGtaJ6MqV1lOt8Q3VoqUevw0wQuBhwkZ+89zplxbDHBX1vHoMQrAbEA4sYuFcuUdzb
hWjtQVKb0MgbQax7ly2FmtsFWa2kQ0kwERpvatz4gOuQcdj3VZqmD9RsuNvIaECDKEi0ZG7iWOWH
k/3wf9SYBJD0TgY2VpK6Bogl4dkSektyvu7KpmPQhbpXNrle7MzfEgDn866tp6oPswImo4Mq48Cb
iU6vEKotbCkZiWkr1zoazckZal5a6zQiyhbHxKkJzN/JW0PZCPaF1edC8/oQkuinbM2+ppNLxlYQ
rQ+6+2q63nKHk2ghm3pCK0zYv+umYLVC5GafvUeIx23WKdaRwZMEjBu5ilrxCnFT3gc/nJy6/+QN
T1PNIFPmwrBQGpTUbIPM4RQWlIXpI4Kb6D4XN3Hnkqq+iglxDLePohJC6+seMO52YBDA/y95jc3t
AbmggxyK8ETJsg60rS+iEUgZnymEndk4zzF08BXpSUGkP09j4EAJdLQ9ehH0pvDb4YKAWHdUqIK7
5rYchOYSJpzfJFST0dR7cVZBrrvs2p6NILWlyoJTofjvhM2BSRgkE36c26CBoC7/cttC8cyvEQID
EuVGDQJKwSxXKQEpQDoI+TM8MZsJ6kCT1W2P5XxeVNrFni3a6F8h2fxuF8O+GOK0qS46bYgJYLUA
KuycH2Y+UrKXUWc49WADo3P2aQ7vxDmN9KmCO4+V9Jfa0dfGXgEA3+qN0IuIEoyukWLpwWJEOX36
XzI5pUqRXbQ4j9y0lELwG7u4jZhccCZMwUBEKWZghCpFNYTRrMnK7doMIl3arCW+GE0GQVeMl0aE
gji3pvOtZPlDOdT7mJv71xsxB/Iejxg0aP45QjIpDirrGnK25ePZgNKzEsJsoE8V/pzkld27fQzT
pyRjJfRPIQ8pOR6nCplrown3fiscVVwV1QFz4mYpv/5a/YcTh0CVBpOZqG4uQy52LuxYXtVUkBit
DFC4YhkS0anJO3Z0ERVkANGy7bIUAIWJVOunIwr6J4PUm5Kpy9ZY6+eSrPNL42rB71Kz1wnQRxjx
14EYIC5oVmDAhgZ3D6qjM++PnTQZgsCpqNx0ZiZNnWnGo16+SPiS0p5aCpVG0jw04ahKQq5FCA9G
1l8hVAgAryxEuUqG5Gyi4KQrFITCnBB2eP87XDuSPPiEQxjmsFcugcom44rz07wDbp6gHZNUtGYZ
eniez+R+duONmAEORhYGwfrz5yY6Cnedp86FX3cgnf29NbeZXCXd59oQTyPbI/B6WFpyapQOsEAr
RUb9OPU1qlVpIpOis2ZlUVdiHBxbIdou5SZo/oDpUlrS/1hKI2ZJ/wwyXBSao7Gi14iV8V0FnLi1
dQktTZvbgdb6ilRv10jO0GPDteSdotnt2zu7QeNaZp0Zx1juIzK+Vq+lzUKWGc4d1Mz8jF0nIu3c
eSwf/B0Yx1YKt/KYBdjSW0oiefZFzpB1rAJFKNf+bZsBlNdsuEQsy7GFFC7Z7VcrEDUvYJBpReHE
+SCOMp0BX4775YfEWcefEiaIs//7RicARoCCF3xvraBWCAyRXaOdEKDjO3kQL/EAgDBngeEG0CUU
zKLA4NTLx9rz/+IsJ2U2+VZVsJEZIWKcZFdJ6jAunrhVyyGfPKAURUc6jgrYE9M5mI6SkC/A03bg
GYQKPxrRQIIogUuVthLkLG6KIUKs51E5leM4Vko0mvv80OzvZEeAEMGhdWLBWEENi/G25j061swA
ZV8eDbH5oJMnSIk+3U6ALOJpKLKq3inQcmVUKq/C2hNgGlLapCNpN2UGVSAAmSafhzpm6X8kiqTs
JqHIi4Fy9Xd02Yfpeeygki5e+nUIAwiMUW4inCkiyTfDhLPOBt3HYobET6o19hcdfxfuUVyhskJv
+zhicoIxMaPJM+m2IsLS3in7R7IgO16IQZ9iVxGtYrzstR3n4ihJ284Y9MBUNUWkVJIbCTyyNtF2
IdhLpq5Ei8KpN51CdlHkYbCcAfDzNttzlHYhk4yj3kMo0M6FeKzXh3iYk3Ff3n4e1Dyph2g0/hL+
DCaQN4Q2yqNIDBfDopfjGna1BwgAEgreXsTgYIRYgi7A/ZYvS4vEue7raSOU1BH8VX90dqtpTHY0
LfNMnxurTp15hNAMCxZwrijfK1MXUO3ph/7Fe31R9dvKdOlntHtIZ6sesX1AaaeN9p1iPeGJ3FZA
FWkHYIKPiCs8Pr755ym5k00iyYNhr00vOtyAOP03ZHPs7wjkxeQ/c0kfAbTPdRfHMME2JDIfDRcn
K74WaOJnlSYfwdfrpsj5N7tb3fYA7wi4kZDV41j74bnIed4GMZNeKRkF0ae1Ef6GUgLZ4dw+29uQ
j6DP9HTlEnnaALgTKC9MQYXAa8U4HmItxk9uvQhW2Z9DFBPzyuRN2Mo98AeO9guNo9w8fv/TDy2F
PEXK3Wl7rSvgto3JC3mnP+GgQYfWTUEvcwIdxOj+PocestK+sk7Ph3EjIsGESfSvtun2kD0gqclg
M9hnRp32TiKkT+M7y5CNNzgPdfYEm7+NDnP2SAkGa6NVmJo+jhs2gpnTIXgvwA6r5X8CgON2zCzf
fCFiDKTGFT5OLh8Qy2PNvwu3QG13pwLh8vgw2TELuxTRKEgJrPZCIzgVwggemUxnrgMuFjCrvEaP
PQyuMCSaTZD7Xm+exzFJ+gTlMAN9wl4ivorFdaTmL4+O7W/RVzqTat0k8H2F+V35Uo5zrcjUz6YD
M+BuPgAKCet0TnhNRg5Q9eDOvr2BFtTk707VQ0DfbBqLJikC6XiCD34Y3+7nBNZ13/My+E6OQ3P/
MmkRO0bWeZzjmPZfae6K6sdSohbOPh6qkeQy8s/Nn/mrSRKDI6IitgDRp2NpJHo8fLbv2lqd/ERn
0VOjoTIUEkUibGbCZaFmCAqvqkKdzbL/3qUwjjiVUjbsJZ3eMlAnZIAonymcHDsfs7UJfM2qidpl
7pBuQT5QsAwAtNgZT1T0xRcfQPKibkCVHIBfpAXEZpKrcy6njP87kCImOmKvKvSfzTiYfPcpUW5P
UoOOTsB95ea7DByaMuFEKtFJUO1edKoaYtNGfMn7MCR7b6gMzzYjQJQ87EmMHaYwVYMr0ryEcY0L
D0vrhM6PiY4VjZEqv/eK5A83KxMqwTwxkhEvPTFjtOsH+VVt0tiM1Kfr2dS9xPUMepRGprrMMnTz
TxAIO0DOs67FskIHMC884xxxoZ2d5uZVQezJIAKigFfaiqxnO5nBRYcqmfRujljMMZcaL7X+57vP
xyMi2aWI3pMKsFZaEINA1+ehGAMjieMDCFJ9jagW2VtfEwpaOkqgu9+YCvGhk+dYONMm3h8muluv
xAoqJ8SVIH3njPUtpd4QU6z1Zqrho+RMl+C/mp/kEH8Ob8hMUljpMBF11qOwdcwkn8+hLLjXKpJv
ucWH5ZG7WLcba0l3jAQts5Gau4D7vF3FBBXe5e56d/Js7sJ/nlanQX10mUe+uh1C2BA1UaI5XgrK
Wd6/o3DFela3FRv1UEiLgmFFx+JUvEbHjpr5use1HKA+5t+3gwesYxBo0L1PSel0kHIvEyOYIRpB
rxftVO2n4aUrxLyftiewUdBqvPkeQYNc72aKEn3j4c61Ia73QVRi3rvBov5ju1d/epgnpay9Z0Lb
XjwwcLjAnqYAsHwAQhsgpkVwx2UFaE26IGJoQwKQOISZ4wAKk0wwPR5eCaa0k2xRwfiKj1H1QW7L
08DC76SDEEQMUimkSz9IBaQYWA34UkyeRnsxjlKWwqNTTfwJ9gk95OqeM92ynj+eWZlQsW0m/9SN
LYrNvhuwFyBXNAVvWn7zTrQM8//iD8aZZNEYziW9oQKO8UQ8gIBoKZwi/1lAQJ6Rd+1h9PkM13HV
qfdDMF7Flogi2TFSpPc5RS5S9n9FkHcIWLxS2SDT3F6hDbV2v5bd2FZujDDjkqdlxrqXz5dTBU5I
Ws+TkXja9T8/3+F/kGaUSLUOXCdWcDnzv0nmVzoP3QvDafGwlHcGtgmGt2STg73As30wT7LR8HuW
ZttyFLFeDeYeg4Q3wYee1278D9PgTmQuSTMMyjOdJ/8almRS2hPL4+Y6iqLnBoeJv0LHewIQj1e+
TGctAnutnKUKBH+fG4w7kAHEcVoIVvlaXwvyHlbNZ+UoKbjuhfsQowK8r/8wQNnzUineAMg5mV7L
MPBWuJxdaO3gy3Q4lioTyY++9itPZichoUQGVgPUo/hgI3srn2WOAZpNOg8fQIz29gh4/sw85h6o
V1SkMCNrIRbw/+EfWx8VQwzUrTcERs+vBdyUugIRdKi6RNpiszd94ac+7mwc37mUzNYGscU6SNNM
ovWLZKyrfvMrHuYTJyyAdTlTxHFkp/WPe5se6/vOLDKtxf5pZ09UrTymSZqNWKxvIXR6WMnq6vi9
4VBNKvd791v8EGg4IT3tt8gc+cO2VxffkBSy2ZIi46BeFeyywztbFecrCNz8eZ3RtMP2TtXNVe0U
Cdxue/0vx6FvXRAjcUPvlyRTMvPkSc4GScFoyEtBjeHdcOPLC3n+B6ogUN5Wt4gWLDGHXuF21XA5
foRCIycInXdyW+VIN3aMHHJwa0vduVTEy7Hm7D+B6tb3Bc2KW7pJgMxA2SMPTldWVfmF/mZPlhNf
eTsraccqTsEIjIcKr3V1OXLKbc2RkY5pObbExrWHWQMF8Z5L7QNTkUj998PNX2rvNPcgNDNrbXhI
skRzZBxqnmYMt8HPoI7t3Sx9cloNrSjlHfnQy1Ee6KF9JoiK7LhQTbTH/4lrCjNlx6aKX/v4t/pY
cArgmMdQWWKlUXfnJ3ef/pv0yxN/YTv6OscXNfk7d7ABTRi+tu1aP0JW4qOOX69ZVBimq5BCQK1v
nMalPt3seIgWIAv3LPioLiNGYJouvt0shA9DuiyMaaxvrZ7whsm01hHqcoVAow5EhrNDD1PYi4qM
8poBOMo0004LjYtRME6uXt5TI+kSIHQ7lpa7SWWqeIRWDtLjPxh2/BVmj+h9DTO/ymFmnXPKNFiM
bQUZeoYfF0eF5s64qhEoeWq3YyPOLWYo/4MEMdf74o6YvcaYKSq4OekgYri7bTEyX3a1TTQGxGZP
xEjMsup6mUs9MoaPzrnvIuX44WMDHDTY37e4WRIiby7yerT2pBtDak3cfDAIgINMPGsFovENwO3+
Du56XTj8iQsGl/8dWhxSDNybzan1Nc3GQJS0G2/2T9Ip3feDaMwVdZCZwTC/xgfXYCs0DQJ/q/+8
7OJfcUEoSRUr0DXSZOXL2juvgPb3aNEhk+MPZDKEOdZPkskTebizG38KccOWZfLcgSHh6ytYFKl3
8vqEhLjSWho6QAcktBUNn5boj3IGWGdDSH1msMtgBd+3Lj/u6km+ReH6lrc6HA2b1qhVN26L8Fel
1wvRnNIcdhnvwWGt7xMeIWGn5syw1NN+lc6+MP16XlDl7WYUK68k19gm1HeFnB/poeQe++BVERJ2
OcChNUOsRnApxhQJ+6omDBg4bRQd6fdZDrhRZDoHmLYsN5agekUdCoSUKJokdBCrp7oFC8QKhabF
trXW3kGYu0yVNq7qH0tsO3VeApJOgDOBq5SZDsyFoOfe5JSx5q6Fxc1MfSPaOISKkL9pYron3yWV
k2IaUb94jHs18tKbXR6eOsQdJSZBXDZNwNQN3JgIIeRUl/PnGiU3XM9FbP5EuUD1znEDA3ydjMRX
VWEC9WYwUQUyav+xrt8O+P6mYdXf3Kp0I0FrXTglTWbFWK/l0W8LrNYDcii8pdNNZ2hGs/tArlsG
FgtI/z9F1IxPhC/ISyKKe2dTYBiRa+fTXZaFHayU46m3nGEn14iOeckooYh1VYAK9/u27RJV7395
XyQ3eLSUWRR6bYxZArbUUdbj3qpuXItrcRUjtAsbYh9kd80Vuzr0arP8Q1nv+9tbUPkjSGcO3fOU
lLUCOHpvr9KbuSzXywc1gQ75dqCjfYXNbHbUqoDdlWv3jpFjSrVJAYaK0ms7k9HSCRMksz11RBaq
dyTVqrzOnMjmYGZGlp9lZReaPOfxCTI2F9Wc2fUKSDl3PJHW5OMitP9IoZIF+AS+Rf9yYDNQEYu9
skxohJiLC7qxLyER7wImMH06KF8HbRmcWnfXDckbwRGCd3SDI8viUNfjNroXxbcwQa0Bu4gcKiaP
yeBb3+1N1zhPXdDv4ey0L3adx3VvtRchxLaBl2CwR7besNal1S9EsyP26utegVI3+ax1f8/cn0Id
+gfBKwdlCoZQXy146qv39oIjzwDaqn10/vvtxobomFErEZ527JVsW/NWLo2++VGECURIZMB7frEQ
X1HDf735MF5IU/fyktPXoQxD/MQ4gTSC6RYQez2Jvz2FOeW+hZ09KgxlrYPdnTLhRljLjVtTUabl
dg8yAwW2hFmJKa+Yk/9exmpYUocK9NF8uZDhxn2H7UHOd7HCZ0Z9cNO+OppARvAr5WHOyPqBJt/2
D44V4uBAwmsOwmUl2GRPPq7IWRrhPaqj7dfVdVRYbDszgOe6Fx2NNwW8Hz7z+YaexiqlbUhaZGZz
AxtUK4uqigG/8cZ8PADOfpys1ob6Pt3u2iU0Z13fj3R5WVEmk3vgiqDdKy/jV16w60od+DJeC+Jo
Y8hfwCJezxv3GObxCtYafabUAlnxvxHXikWInfzITrVn6mnY1ncx0Mn2/RNvGPeVqul3HykQ26IK
nnNFHUSBx0LF8efGdgd6sK4FcYWEeItSQbwj8KagUsFL0KLgTYSg3oNyU+9SzmToLBqAyN0WSl6l
QFBCJDZERpTFcMfV39Um6gk/HTIGr1RnTqlsP36YbTl1UTC+7vxaGYKR8+76wajyMRLhp+lOHwQf
97KMQLPN7mPlEeJYt7o8VB78tg0PuAQVtCY+SwSJ03DSAp53XzuWt16zlrOONqtA1wavOLAid6yM
ajyJpakQks2vEMYgtEoGuD3nBkAsG6LwerR5v+sbq/YRS5obNUwWz/+dscfwi3qmMl1/sYQJykO1
yAt0CXMHNpr7GagJ9abd+XbD+F35k/c0YXtP2yZmfdSycYu59Q09+GF1U8KzIqXjAsJ5ZY7ingig
6veH3ST36p3K24vQM9451i2Pu1Gt4patBPkSM0PQFiLgmyZFt2jqNdFlAL60Gl0GelvPW++N63Z9
0DCYb+1PaY/IAjBlfO8GMSPYQBix7CA3bwnm/amFAbWA0xm1qsI8JRQcxCHY8nWBuZnE3HX8fDNu
cm5CshgCwwgbS/kkdxbd53kxgUZ1XJ7u/wqPb8RnDS8kzxSSb5VX3r2nek9+eFjR+47iP7ap53zP
43C39hbxTchZaxmACUF4IOfhOMhoNfD/lGn5Jql/b0cZDzStVNPPZibn9PSi8bRxoZwn5AE7pO1k
XWj2grcAC2jEPW8zlkR4s1pqSd8GRlxSadz4fYZWC5MFfE8rTX4KuKheaLTGsLbdUEvUniC5fDqH
S4AE2TpBJcJTgQaULZTexBV5zOY/41oE14VrDne5ap8df4a8T7VY2Ec6Cly5cKBw0MOrT0lniJSz
we9AUeOW5LdWV4/Hw1swRXGBDJ4owQli8E3bYWN4hwpAQWsp6YjVBKNNZmL0qTtp6ZtkskrReGHl
hgGRfldaibwWcQAQi4X/EWGyoSfDIKHajYVieNBtf25fxibwLqx6aHYYBm+1ueTkjCw96zTNo6gb
wE8wVIzT5y7UIAlmatC3GGxr81ABY71dfMII5WJtdec6nfOmiP5MyZ3ogQH9NzOwXo7KKS2MC9Xy
V1cVobqpWIUUqn2CyQSz9AVeAo53lXg/UghumzpassAQQqVTuK4q1e4iB9397Vr+aKcUVwLiQ7O3
2lePgT4c1vss2zIJuhEsokMkxHy1AA8On41ok0APe73nu+JECVyeQjctMC8Wt6g1SvNLgjKHjZ0f
ALNDx+KzY3+/IQT4g+JPotrP+1tmdaAXGvKqAdRvptG2qfYoNY2mDIPe/awufP57G89kqouU2lAv
O/TtOUDkZZWSGYJfKubUF/lUskSxX9jMYHZT0+KBd3nuwyc0o9Lt8f7rL5VSEj7R8k2tMPEftrrt
B6APnJzypNiY2WQLdqI//Ak7SQFmmeZbKx/Ng049blgcXuT5B3y+B1eLCgUb4VN7YEUQCOzzvovl
zxVFLJM0p/x3nzs6aqt2uLidG6f13aYEvSDS7Xf9900/IandS3CxDGCzSOKh2M6wFupS12xNZ4sk
VIeqn2pbiF3k8MY4nluK/Wb80IH4ui0fzR1LlIkJLHUAMAefcXV7VkxpnFT8pcEIAeHp1c77vM2b
6fDWizLrDyJCOdDSdfybMgEu+CswQkfW4dxSKaRpE7I0m0IO1DhJBmbk/suhgK/IymZrVH76SEMa
6UFWpJ1uArGsr44G/Vdz8W2CQ1DtbV5Vj412e9BBFmCkyJcbqiSnrQEk52e0VMddKMnNkOCRCbPh
/67jaU+YSpEX8bFGdCB1E+v7Ntnd41qkhq+JdePF+kCuDvXJJMesR1zeJLwyF6eZdJgpSqkQpMgQ
0UNirT/2sRN5qdUhbL1l0PbVdl+i0UonrK9gn+qNZsDTVY/ryqRT4tKuROp02IbnQHsjIvXhfQYv
co0HIPRNbbz0V9jLFEQWfoLLfKxaVnTbWZf+aYONmIL6+Jow4Tj2CrPomslNr8ebQAdxnDqtanDF
5Cv9ZM1pHQnw0NjZK3RUCmHzdQzrXNZEOIuffvuRZvAfQA7+5n/VVxG2dlAUYRKbkGISL+k0HJnu
EoY15qsyXak2bRqULAhhYDUlxGyoAwGr7YH5J0EwEyQE9piDk67j53ICSAzgxpALx6H85hzH3+sj
WZQ0PPXs9Gmn4EeBHonbPfUJZaVeY/yLWrxfu+Fft+A+OMov1Qa0mLbEtLuVe280E5IH4U7w7H2z
ve3vSJjQDikwHZ8DBBfFRCIBVa+gZ30c9ElUmyYROB4kV0viRRfBxeFEQpPhlpweoTbtfPeTdXTX
tTkxAJ9+SyVQ+Ugpsvh8zaTwEgKM0Th/trgZU4VlUV730pSLU9CdeByYxa3mcZvSf4NHgy/JPEaA
KAuzTwzhO/+h8b5GtQ2nkjiK3pQnPwIor14qGjkiMyZ1nYNbtF6soP8HnCaRDNqxNZaWYM9ZEdzK
5O5WgDx8mGMvjB1xUDwSIr2AP3jEFch4kYfdWDndw1LRgqRmyQqPDfnVGwYG/iYI8YGFDCA+z5Jb
1jmkd7/tz0vLjc4WvxWvKVQAx9s8oSZ0Qu33fVk0EGQ+iKAW+b4uRrB7W+oF0Eo2biyzWTKD2wiV
X8v3CTCQGQp8PwdcRPzMuekIn5JQS5nXBUkMcuOlLJXETeZBhG3ew8daV9VHWy05W+nWD449Zgnf
gBq6A2ZTXmSxHJVRv6ny1mj8ilN7/bELuAHqFtLJeCAXANSozlPkg8ZgriSotTXA97h4BpyEnZda
jQI/UJbkoj46SiDLERORR6jrOvtlvRboxpospHDkgKyi8WlpRADUW8qcRjjCK2tKIx3SlXPW4WHR
3erS6K9GWOjyllC6NFEd3/hcYFl/x2urj0QGoyJIu5oShr3Xs4hCdY0/qt3daXFrsICP/spa4x3F
RTqfrgbOpX2SVpFq69F/ZDJFsYmSk8TDZe42TWLX9nBJmZjJCnYMp8K8MYJ3YU80qP26JUstrGap
xtzKREfkdWKrh3iuA93SUSgz3cUVzsM5kqp0BuDSBg83xZ1sZT8qqJJd5aksT7tCWdjSmiV+A0wR
elFYi8NNgaf1Boo5ydc98BxTwbGmC8bCAzQKKNMOqy1347otLn+VHp9UbCSZ91xrYhz196gAkQKk
V7Z9ppnH4PRtpHowe811RTy9x7jfSRuRwaipkeLwOpIDAmT3/MJOMrhnOkVLGyL/W+4iYBEaig1m
lU/xGPiaXCqFkV+02S1qeowzHMy9k147PdA7EdYJIEnq/zTHij039S0YgT2j0LBuSZgh93Z4WEY6
WC8V4MpNYWpUGSKM+YBByIDfB2q4h6Q1gjGRyxVcz+6qn6Si5fD/X9F9czuvpr7Z6bNrIBoxvV4+
UUDEZtAm9HW0UM4mOj+2LsQ83buHPBDtB3NJk+k/osyLqat32qetpCjcPd1Ck8Vnh2O+RlVi+HVn
9bZKV8akhf1CS8HLTDBWNmQyBwX9JaMA0hcIxlwBBwgOupM9wkHlQiY4e0U0fS9rT9CqqOu0vTOL
B/0XJTVd+GUn2yaugJkE9vEY/zeb/1Zv5zzTOhz0becm6Dp+9ShazH9LFTubASO99GwiZP52PLfa
6RLLvn64nh/lCRznPkTZzbbUjW+sWFLYtcLfsFthj5PLAWZbsrYFUvMxTaY3CAy0KSQkUKzhUnxR
0y3G+3lo7pysRuzFbd4p0Zrauyq/qIml/KCyIZ4Bc+lw44dUkOqansytfia/UZJxsumZcBTgnBVj
ZOaIvHqginNNG7ZNin2V4z1HFH8qAqlHrVmEk/rCYK1wTz8dRRCszn5/NUpXFfQRf0tRpNyqaiT9
0potdQieVU9OCnmc6/DhHPaBOSi8HLdFL7nv+S0PQKeCS/cHcPvaUo4sO76BKRQjS9mJP10Pwkga
k9tOGc6mg7zFAg2i3WPtdvIb4fyjspfGRFJfP9CeQNrqwrIHQVHVYGPjAF1KPxlPfxd255UIi3c1
vPovf3dSYA+/pvRRUTaKEMmgI95KKpJyY5q3Sl0p5myaKehbsuclCUxht8VbKnmrd/e2mOj4ki1T
PFdfIDVgfeHSFerlr5N0ljfrOdt7qhjER36tpYm5JLAFZUoKeV2LrpQn3OPYBr/fzuT10jvYXus/
rAnXpo21ajF08JKUZUVuNVaINWT9ElPirfv0uBEZ/GY6idqK7zS7YgXkBYM6pmY3XiTCCQs7mIoz
QtkjnhjA3LwkJRvAqknptrL0nKk6uxHn9FdBeIGdIaeUM+CLB/1xhZDApNq+GD5ciNHhMuBDfrep
/vEsXTQWKCZX3Fa1dql5RuZVnzTLlAKtei+ZY1oPgkhNMuQFZ1ETkn2dxyVzuh/250ohkgVET0lA
sOkJu35D1l+z4177B2OfvTOUD4D+OMkbN9cWCViKL3CPwOpeUk/v8Q1f7sZueYoeqBH9hkSbttKK
C9JRfV1KJis+eRl/+WULOLIMWU75mbn7cODkett9TN2qGadfM9XRvEFw+g/7e7LlLC0tSl3L2xIN
dHeGQXvDeMnto36Gm4bVmZNvVGaD0f8Q1d75nlpVswGPEyS6pwlWJFDlJKdBKqtuhBCE52UMro2V
QUhzRgZHTSlxc8IQxqfeHWqCP6jQOhrNYv6wYSE10438lw2unetP2Jx1SklUhuxiQyKSELCBf5gB
nATSSW/vlj8Z9UQM9cFkU5DiCB+lG5NOVDBKr6ZDBjiwG+ipvMqPs2p+9vrn4x316VD2qEMuNbBK
El2H6K8aOsXGKfB7YpAaDL2Ct+2J/Vl1MUKxh+xEE21sbB/xqdBZPSC/bH7B9JVy9r8bMXuQhqtf
DhlpOijeg+bG/VQpEed1pdZHTFtkHzq87cis53/xTB3AzrB4rMMiNesmD82GIeeq7C0pwyHSrmO7
NVTQ5vaBWIGwgngpR1amMJmjnsC2rVODDnTlN5smhg5jbTaifrLIx4R0wXH4/brLU2wD/KYRJdCY
L4JLh7CwASgQdqGqvW8IwPttrByWMjjWrqT/wsLw3cZiky+wrwM+ydfmSiUwE71XTGC0CzUE7MmK
Rn8ppwVf2rmI4d2nN4QbD+NL8PkMZ80/jw7RdK7cB8zBIWkqeIh8KNLgfmftC1ikpmR8HGZE4ASC
7Ygz5d8FKrGGSWjW9maShzeFRNJZAXJf4WMINlyNb2tQYKGhjcFMn2YK1FP8oxtMrnp68DU3Ln5f
tOIU7dVAtR0N/ADVyfkXb7HEkniGzvprglj80zQ4zkgNnid2h+vBilitqdhRQSG3NlW8sACMwfoo
rnbIBUvKcf3TALzBqDm/MM0kYRJGIcYfsbirEjHJd02NSnYbRMJdvZfZlgLzi/Y8iVblyKN+H10V
Il8QW5aagRL51Tzjin6clrk52+pMfZCve2FWw+n1FITbbvgOYO1lElCK8A1Se04EFq/1gF2FUC/l
/rL3uufcDgoU+fzoleUyp71f/oqeW91qDDCNBka8vWRSZajjbUXh14pmO/c88QnyefHMkk+QeUBm
lLqI7ZLU2+dGAACf0ZwW0YA70KxO1XLeFJYURHDIpF/mAeXxRY99fTQR0TpcYPu9yXYE7PYd2uPf
eIDkAdV0aHYHNFYfDxTGzmBvTlGcsOaenSu65Rz1BHQVgexxvD+90pTPz9fR/jKaw8MGCQQ1al4b
9Wu9MU9VVGOo0z51fKQqRDdN6Zn64uYOitAn14uNLbEWj5eS4LqOOs3iEa3JEgZe1WwUU41/7k6y
sYqnyGjqkoYB61DtULIYVBU/SS0zAQtueoUF2xZ6kcFumcPlzKvgn4G2gvC9Z2FxC4wo+OprTqDE
ZlpqFVfdZ+IF8c5K5kl+WLT9h0XZyRsxPwXA3IKVUpfEW6p6eMr0TIvOEfoC5Ww+o/14hYiqzRDU
fhn43ClAmMGDd2EPKaSozv+HObKQxN4DrX2dALtCPXOApQu7J4tyuX/L2jDDpgmSsRBlHXCMfm2O
gNM0Nzhc/7RnI9Lv4UmerLBp/uNfF0f8IPMYMqNyxJJhVM/u0S37VVBuPZgk4P8sCX2mm9fwB1m6
8rjPjGO0Of4FXR6dzA/I/dmCNj1uQhnW/gFmCl+XCaScMkUHOOuNOh+LOTejhtFgkKzrAbGt/jLy
ASuT9024XGIymfrMC0EoobpFCWf+75F+ahxmwsOrkam6f7HrKJuAWyuzG4nLbWn98gS5s5cEUKCm
rSplUkwsoPxTZxvB1EErDBSJAdZAzixKDj0aBi4ZpDmT3hnI4+7dOvVnI091Vj5w7UXBeu36G/2F
RarA2IoreH781PMUdLmYywJ+Y1ACbxy3D77YACwG/KuR+ujIJUgPIe03d03BKJSnnCJy62Qbb5t5
LaKq//dtF7YfLQPH2pz7idAb6CPgYtgV5RtrGmQeAQgD3bgvGStxFBUXuWf9yZorQunq3PF9+4cI
uSg1TOwmH2g7TCyhjIRd9C83lek6AALghMJJmpy4oivWzEUeCm41j68KE5QTenYBj6/iDP8Us8+V
A5VdX6unJGC6OBPXDE84WcdbXOU44Uy18xODpB1/l1hzSiJ6uo6Ic+kUVoMmb7NUcYB2+QFtR+jV
4d4+bwp5LPwg2IgGijGqZ6dr8fEqloVH/c36whsnFXxKTiXJAxNXWiBzmmKz5cDdxmGVvX+dUquk
VvE9y+FyqXmof6ymuad6OcIfCUI+HWB8NH1u9D3UF3khBkXXHn97koHPdlLgvUmLgNiByB38UHIV
wshjgRhqktwmettCcnN8Itp9vmRnxT8zYRft9SUIgMgICMTO5Ea/ZtkP0yn6/bxopkjS3pcDraFR
9FyNv0+gF+JO3hZPnVpgwIUp1D3bHfW9HuUdeIfUwIJGTW5+BWt3FuwbomAkEfxEglvtLEnpWvA7
E3DrfLeOykFwAXQn9iG5CPp2uhJ8NeEHLlhJqdt7k4MUYY9poIxI0VtBL1TozhOwWRhL1rLShm00
u4HfGa/asKsLjWA4o4XCva7o2EPvIsEP2DDwtjGMHiKqzymyBIMH7ISdC8PqDGTySPcteCb6VnWC
ld980gurThbdDUpYjShQ0gqzqd+AwIQwi6IGckRdYLTxyXVMqvSiThCRTIGYH2tot6aBySFDVPRs
fNBwqVF5yBUhFMjZIN9cFYp9rogd2007xpB80cj7dDStlPScbrw4WL0y7dYZfDe0fcXQo3Wlm8JL
y3SWDFdHoVjGPRiFsdII2/ev075RzJn6z/0Qm29XF3G07RKhtudFgsiA6Wm0W0yBXSjKT1ggoV0Z
OTCtRHGqcp4FH4NKXRsKJOc/beJvNr+2i8RXcsoVpYCM80y85gRTAyawHP2NgOjesZm5+U6ue3+N
5xn0Za5PqzSL3YuQfPvCfLidqN96D/7uUDdz0Ry5bU/SpYQ7BbEYaZ9rXKqsBQUJDz31wWmGww2U
QZ/RVFKjqn/po+VTrTe6idmqh6RUlzjyWsBYgI7scRaMU6mu9wqdWcahG/ITCMkTJXSOIibp4/QE
gZu9xY3hIE5ZghNSoNOs7W5TklDOaJXA8rraiia7PXQsEUW3yejBqXxJCSSxxMjHQXXWNbtmS5R+
V84Yajak44M2ogDCUXXK3L/kG0q/4PUg+ooPlmpv1RsND0Xcknm/Y72KJXqAysB8X73GLNXaYcDq
abubnoOLMh2KiNdHgvoOMeOgcg8MDSYAs3YpEW9AgVVIrkez9Nv9FKcD6tQJBUbWe+k3tSShHqJ1
tMaderw53jfAqW2hmOgJO7ozuiEXratUts23kLRl4fQtPczGZt+UxAos3AyyMPu6EZ4uLys0lC1l
6rfY0eA/AgZYIn1jaT4Xo4Op1osmWSBp/NCFMVPQjQDfkGm4tiQ5ebgXQ9y/Q3TzhYO0cAPTglDG
jIhxzFnEtqSPexyguS8nw8Nt/imUIbIipUp0D4IkhiYBvdXymS/Acw+53COdGFtiMDJqdzcFRj9n
P6dfae6yH28Bg6Xd3XM8ZWr0+BOJy9oBHrEOQbh9Nu5hImTQoaFZB+3dd0A40e1wa9gpSu6ZlMz7
r6JbFdMhK9nw+VX4cdAMffFDSSOe79AusVPF8zbRkUMT40nfQ7Zuwch0Cc9qxFLHkdcw7Uhz387W
CEoKT459YoAf0VMJdvXbCup2GMM9k3OYS9gcxOAvx8ea0PqfbyjzxgQX/jTLlrVxHl2rcRO4boD/
MuRdeKh00cRn+teQiLo0PDdW9IJ9f0XEBDUEZNqTYA65idpmGnKogYXkwUJfe4F6uKKdyKmNJ2/3
7drHqCwt+gUfChw5qfNDZHV7chlZKIvQZ4dZvH0PLqC90P/tbAj8mHeobA6YzkeiS+Jfy629O0HI
zFWAe5jJxPxfBkA9GjnXh40Hc/x4GG0KBjV152gTF6njQkariDHab84+Bg901f/kUS6MKUBxu+3F
0JDgrvd4TOJx9XXkA/JWUyfVCEZZs4CG6Ofz3mqUmTSJCxzOV84GqPmwyg+ObETMTieoMwwSeyVd
vJg3jIsFopNG7VI0AP9lZN+pEr7Mm00xm3nhxjqA7Vsfui24BM0tR2/8vwhge2Lo3neglr+3ioRO
/kr1X+m3m19uowilPXsyjCAS2n2IsKS7lwEYr5qosF0tY2u8ZSHLE7ZnmOfeIRGiUSz9bU2h318H
j4l+IJHypT6s3jnwKjujZJ+WDFxrlM7mxOJ3ZsRNFJ1LSKgCiIXmEXPJBF+hsvNL3OvsGBiVaMyd
I+GzyaoHmm9lcoku7H8AeVQul20AKzqYSurQ6s9BLNnOpa6CgzTrPkkY3IVAnt2f0Ujc96Y+dyDf
N/jWgmgmIH7d2Gr97OdELTfa3NO9WqjoDs2wNEczyWbKHu/UodvWDpzSw8RuuH0aMeCUv+2sPFPZ
G4bXgaKJaZmRSK9RAIPGyVzUdQx981+fQ+dVLURlEBV9H8RJwIbzPeSRHGsjhaKt2wIchaX5v8cL
AeV1vGz3tU60uLwXULVZETKKKLt+Q67TTqInrjfAXere7KJj4yn1gKho+dY4j6RDRqMLzpnRqTBf
w6s/KeaUSSyWUwLntxwGTFJP2qpa+kip6FUNlc9wjbmtdntJRHiPobTPVXFTLBSvZWO6C3WN1RSP
YGbFmHZQTM9i9xFIuxOfnZrJ2QF4E258F97MYSYYJJb0W+8vU4uoBs6seci5Vs4+vDFZ0W0Zc+cC
heNmfSOkMoNiJO34zUWJpM6+UE/9bhDYFQ6UDJVCG6EWkbnJiO9p32tl01T7sQQnQjydnovvQU3T
HWWG8celPJjrlfBxYTRRjjCW/x66sNcuwFpN1ftNNHxRbFKvYNrBKTbUPHNDAuORVgfdX3F0zR8y
aKXNRrI9tclysrQ/lp7SvQItaNKI65pc4SACrRkZUdHCWZ2inkyD6P8o0gsmhPM6BfJ9GuBWihBR
Dcq3DW6QtxZODYc1kmd+Pg7lIsNLPJUzI6H5J86sNp02IqhqlbPpAxH32IB3W3qPIaOQ8hBlgLlz
9nh0qUfCM87YpJpOLGo68ywr6R4yCN+mZarbZ94mATyzw2f40LYkOkjll3P++1ivQiISFbwRFTkb
TikvrgVKodkDedfKteWwNKs6aehPhQ/nHfNZ6/ksg9uVR1tQK1k8ZIras07CZYAiTvVnMWcZeneu
468lSUpKqW/P5yHl/LU50s+1vxCCoqD744dJ03N4fETmdEKBe0Dy0royG8Bwz5Umy7FvBt+QpNuS
otCjNa/UGYZH/PWBNNlnQWofmDRWIO5txTd1es4zKlzO03bEtQgRhYELOTi+3Av1XMB09dNlN2Lt
mNwBOw3TyhhfM1UTs5rLwYexiaHO+LM+ph4mbCdie6uU0c3dyoCMeMVL8wSWpVqjT9trIfvFe9gr
7GhN5J/rBjLL35DTYGfBhsbhHJuePgB+mZoAdiaSed0Ni/RF2JOA57buxlNjo+8IhRftBSN8iJ3W
Whr3pq80mBgH/Tb7RSph7iZjyTITekggts01gqATND+ETOMWr+G0n2kkSbla6JV8bWpbTGwMLrkk
3vq5XL2Q8rvGHBG8G+BZRK7TiGmKQ9nsXvlLrvWB2yOJBcqR51NAgehrA4O37E1Z0DSE0MT88Yrc
QwtACFeqySSDdMyoKgi3Z1TCB4kjs5proyMnQb4t+cdg2NJzfNUjUWXcJ4HrIoS2AnSe6uUVudN9
wJhIxQsoRIyyeCRvDHhmpduJXvXvvTo5I8/Ko5uGK+AK3YvkiN4utdgunc9M1O1OguKRYF6s7suE
ZNb9yvrgUVObUtOQFMTyO78VIn3UMkLC3DDkXhcJnGj4VpHqmOGhhWOvOG4sE2UvI5RnXdbxJ5cY
CbkzONygGwpmxQ7xDpou+pragXHjvvOsNLkzOoiD+PNgzyGFt/R7TvEnUDIasevUq2LLKAsiN/i3
FveKdKcYwlTXQaxAs19/kxXhkrIFYTHXDsIYnfsmJ7WX+RPFX1O49gYkJoIB8WVGwsHEamNIsXzb
v37XEChnjRcMZFiRTBTS8nALfcW63IKk5h497nVrHZrhYdatdJOo1HtpV7YkxRUaXs7i7QWOnIBp
av6//s//HB0nI/kYLfoxogGkRvdVef5b2EO9sis8IDptBNQC17bbA7DBuTKJNqDCyXzHeRL4v8hT
Xyitw1YvqkzTOAImfRsXdX2vupPqlFkSw+5IYrZAfYduSXsUEn0L0x2FB78rh0hcUoRymMOS/aMb
hBPPnKwDUcfjDYf5xf+/NT3ZQxOyrI7hoy2V+j8Tvo3VU/rGO7FYYhw37TENkBCRYdYd5LfWC2Hm
9SMjnJjT9OXLOfjGzuBlCHAL8oEIRZLsD5Z+oZDKu+TfPmnae0343qOE6DbNre9pBzJKcdri7UC7
LKYgeE81i0NyGrp40rvhA+IAQxhA4NkXlbXkyqFJ2VgnpkCCh0CRPcv0ZLJcow474QR1BHnCehUe
nFXOvLStGUXvGzKfP9/nYHmZ+8vsDKJhlawSZAEJz5LKJFlvuIl6vgTWv5tLdI3yxSd3Kh0tQnrk
0QWX8zAk472GqPbC3uQpvjapIZ9JG1SJO3CdU9TgomUUOv1b5Ek1qubdwev1lAGZ2zR90C7TNBvz
EtLrAh4o1ROt6Zkue5cB2IKt8jXTlEyRWlfm4ogVU4RiRmhcgTNBdzdzkCja8F5pd3rqnZmLyVXx
sDsfEz4VVjVdUJyOSImRKRqLBnVUNs7f0KshxGDRS8/WjjUoyo50zWkXWC9V4X1JaAqYyl+wYl5R
rgpPxVDJzPdaV8CwY0yySJOY8lR/qmGO8U/CrHU0x3cN8GpNJ9AjoxrAzq/vG6PR0DoHFPXArwVq
GE1zYvi3be9lgeruzBb+/DyyTy3wx0E0y6hwGByB68uQDdqe/vu8HG3tQVkuCHsqT83xs/POncE6
pDZVbjEqoqdSUrxTv6P0TT9RYN8Oqe8BjPa+PZ7vj4zOUGtIWSTJazDP7FPy079w7L8CVbchSKaH
bLMGjCAwjFLbdSgQJRePIONLtesQs+XqATVUQgJx/s+VisA7ylqOpesPo9cA8VucFGHxhzUQfAPO
g/WfJSCGsb4GYd5JbFxamMRU88k9okaGTNPDrSx3adV4a755SIy8CsoPlWuewTyoSw7gPclm+bQ1
q3ERW0G+avj+ZzRWUoVORvk2zg0g6BHp8Gnwg/U709luEIxXPk0Ayxr0seEM49IsDMWQsSWKchfU
Ys/eowa6eroSMkARkcrc7XpuE15MklB/Y9HCdNcXsWXy3SmTGIpL9mkq9y+eBsqYizZnapLofMz6
H/7RNqFSuiamtMod7Gas3PmCcQrJjGpFSePavgRlq4X2PdMykMXCVOgYZoLz/i1KferWZuX7Lft9
qPasBHx2Z4Asf/LCjDKHnE2oHq8levLa+8lchadDcZiVMlYReQGxnjMAQJt21/xXwrVg145AXhCZ
Hu272EPEhJgAqDVJQgP1LEs1BNQzLmb/omjYtGIVJOw2MOJmi0LE7y20pNLExhb9ZkVNxg2vDjAC
nvQseKjAa+DmiHqK4IRRCpfkLXEq9wyvysWVLPXgRQZMCa6QudGjzjWdmyVhAKKvoZ5EWoo+26BZ
L1/4Wa96fJZbcwoJreRb1mvr66ClTnaHuVTm7LlE/wbzxZArs7q5ChZZH9NmNYt3CKZ3eycvJRE+
6osr9k3yYIN2Pt0lATD839yawM7iuFZPfpDdoegPgkbR3nk8dq/MhsAmvzMbeN4zMHpKJU3kG9Ew
xCsdUdFMiJlJS+ZQoQ/34u49Gngop7VkBXg0heFFGDRNJaKiJTGgrKqnz1ERd9AdeI1XRAvltBf8
DeZ3PD9QglG30fRwaWVKZ0AkgQ+GoXFFXU8DuAi+ZBMjBrVFf0Ar1B7RHn4zDyqR3buZ01xl7Orz
KRSUf4GjjPjQxH4vG4GVorUo/JKq50P1oRkXwU5HPdxxrX0Zt+gf8CaJncyWhqqxxHhsMWdV8oH2
vn12iuSul3v7NHZ4qm8ADph3JN9uLutDtX/csLD7pcuaioDfEq3PU73UIJdWzM/qerJJhir2HPCB
qgJS4GA30Nu14zK+YWEPq2hd42jAP45C9D6+PEWKuAqPWz7rAqsCD7B+Hb+yzDzUp79c3z8KxGqJ
3fFX216Qe4EB3vimqbz/bcFzV9S33E6RyFioBFNJ/LwLRTHwW62Hos7IaZeDCj1Qsg46G8BbT78n
HDKm6SeEtIUCQBRbPjBAlEZV6LJNtHresWK5w0McI4zE/3q/kRmFqWvvF2jebBpZf54R+9h2Q/LW
o2mexQqW23Giwf7MQ0gLmeAHeWQ2H3x490bbLMRQoFfM5OcNftkK9cejHtsyzVt74Kb4t+xCeKCH
O+MzU+rTVyRTrph6B96bvqtAY1oOw8ti8WwKzYxrXK5qZpPhx9efOU220279fYjL2VpnBZXgpZ5Y
reZ/8ZTJD1iA24sa1yqTrorVKd+0lS25hm99q+PstGHz0ohCKCB6YY6mY6wkSdiNHriWGHsjFv++
iMkE7C22puCiWio1ExR54vPfp8jGh4FZ53/aqAWM6dbJW6Ei4ojsqOCYE/OtLOmS5fSqey11jQo+
c0xKqwmF4dJWwFGCePDZbrTa452Z0jt/U7y6SP/IMxRUAwAHszkrPRgbCX4t1PsXahGBtbgwMJgr
FXsecunSDgWtevaPVjLZoEjmoCxk0xsA9V09M+XlQLNq2T8AmDN9E1ReqdnHjHJaOwOScD4BT/Fa
RyJvpQbnyNmKt75yIGVNNRXc2B6MhYBN1ghRfS7tVcLIakq2UHejKTK417YvhggUhNU8MYJ9V6IQ
iRXEF+ur5/9H0UU/pRsM275LCWOEsZIHb1qJZ+Rn6r7FoyJlx7bQV34QCCEb6FmZc4IakyFoh9ry
MLlfdCbS+bjo+0Y0S15gMv4vBhRmYJxRDQCgQzjY9562ZR0RkGJ0Iz2qf2qPyrzAjXKvu/j0kYhX
cJeSKEK46VNl5O6KrTMq4jaXVp6mbTfgYKqMUPZ86VUcaHL8c/r3j2s2AYHoBREwl7S1KnWerN41
mLjOR4nzAmPrjvrXO2/D0609aUqko0DVzlbv3bFKz9+gLvft4gL/cu++iRz5DWTAMjPzIiFCtJCM
eBJjOvMvMOQsthVYcOayAn/PORze+SJBArBp/0f8DGIWqVJTs5GGm1rYnwoA4FXsO9eqZcFCuCNY
HRb/CXGnocyt+S/Q6vwpCH/EzlTqQfStegB0yWxR4G8bGZVlNht4VYcj7sABZBaPjjs3tKxDOJTS
lQ/VRoK4SfgPyTxkai6ikhZMK8jLfz6+2s38h4ozCDIoZxv5QsPgC1wCLzYCX11FN9F6/IJCKNh2
FQ8vEkleDCYPTnsHBg3Us4dQ6efw/BrH79cEgtN3LF7+JIgrme5IeO+oLF+RpdgxpDgXLR3uaXRL
MCMpP9K8XeQTs1I35vszAvqsOp+xoUp3D4LLjNbEBQPQfRwiLJcMYOyobGUcyuXPT8qDtmdJAtpK
GEslbhnw7VLxlikXddd9QOKZ9QWFZDrj+llFVghjmIbvNA/H0f8DnUfdF7u07OXadW8/Pb9DZqi7
ERU4tCBIb1G4Wo/9Ns5rW5aRHHFwbKUgcXoEAAseYhDT+PXZ9izthCYx1tLDVw02n7MT28wvz7im
6I31UL5hZFQfd/xo0zjRad6GGHyEuEy/u4GrRhi9NOEbg42IcAYFRX33SQ2waMo1VRCfDK5Zm8cJ
uX1sO8IXVnQbpcS7y8vqDWF9rOL0LTOGOoWPbuhbH5twC6Di5K87kzaqRzrHt0nHkwNr5LVmI9rv
MCKo+xzEXa4uuFVepHNrJ8/eOzYdJf3plkTE6LGC2O0KkgVF04mvJndyXmE7hCOuIOGzlicQPFIt
P4F0uJsZjOPqAS1WOM3BahqreLyQG5TbIBriIcEyqnzo5PAmDz9C0XP6FhoenvccdVfL2AFHMAye
l6w2TgMJ05/gwzKu5RMcKM4kJtH74btmFU1dmdYtfEZy2NWc/0ZfCkKrw+2ELMXaD6DMqhsFS33j
OTiauhRuKeraLv8J0lw5SMhThQKMa4BcDeQjp3IzbU9y1gKsA46GTQWpS/+ZqHXNsq/bHi8XSdCo
1+ebuqQ2TvcmiKPnuy9KLYDWgUZNZ7HeKweeGJM/iliSbYW3xejqVttQqMvBmk4VCwZLIccNmrne
8pZq+E/XrqWDDvipTAksFum5Nqj1igpyUdD+JkP1IHg0QFejEFqQq7sYqqe+gYFHaxyKFwwKogm+
NY4ifLBgr85qxnDCtlIggTVMD0Xntnu3KOITo5At9+2VY4dYr0Z0wAgkDuiTaDOLDDKDasVPv7lW
jFQUGrr60Pwcbd557KY9qJemlASW2OfgenH4GVZYD2tbWzKLXYH3QIEqxEKsAXMMLvpOcKQBlYB7
50HBePr1TAmTDX1PuUOaC7WbtP2HDa7naPzk/7sDPoV5EL+rcpVtAIpXYEvzUaeOv9ZFaiHCj05T
p3k+iE2D/2nsRZ7L7kwDlY9V7fCTa2GP6fhEsz8oK+kEmM5Ywn8haQ0auLezbfxT1PswR4Mcr5hS
achWEWOG9KodZByByNTNMV9WKGaphgxSRypWnAXgddUSvLnzdH2vsoZgcx2b4EC3uNOcP8nbvUTR
JBFcdS9TDs/c0Ue45WLxzC7tcW/j3XVFFjYomPsqMmdbeZD4uGqh4C0VnfgFa8GET6kVxryAam5E
PyXi0KjEz1259pcYCOV4K15IsHGXUxjnXs5qU4SS71Pm5ewNsrgYnxEjdwe2gAxEU8yyUGcJdS5a
qI76kA4Wo65U74/NBpb+qd5rMqvse4qwMuxtfutIKWowxbUebl1bw6BYi96eCC25MuGIWDqoaSh3
emNpWfNjrmIXvaFe31oPk+bi6samukxlmoJ8K1MH0WSd5aVq5HPSEOphziztuRR9TfPBbDgNBhfK
GfMp1gB5RtI5bixSb4CUgAR06lcsms97saiBseh80+ScAmIvmwU/QNpadgK+3w05wHS+tDqGY2xx
aeRyRndRO3IPoQxmxVrYgeDXxWIpsaZbimqSgIMDh91U59Z10cK0G9TwIbPEFDmCN4SFszMKB00T
nrVHRK7pjjzF6QBtiImnTrVJR9Wm2JxvpvWHV41sjdJJ/0DP4NTUlK9FbwO8Gh687YYFKUe/mGCV
NCeHsoK3/5zmBweb0H6AsBMb3qkyxrvgTE8rKkNpkOGrioib8FQMxyfHFqHh14IC2aBEl7mUiMl0
a7990lunbZ0buTw2nnsMXdWX6kMw8ZjL0z4JvB4pR2NYrkQ0JlbHmWAqJfGJTvtS7HmwRbpPDK1g
OnrBJ8R/ncvCbGw/gLZcxSrzo56UQS7bNttW4j3//zW8qdaun8TD7+w4PHT84nSDYmLyOYV1UwfF
CGR6FOVDKsog153lwTj44sEzdoaXO4t98e8nExLFJ6y6VXy3zQ6i/vlQnPMKsrLt33sOeHx5mdwx
XOGGuHDglbtUmspyf90xWHMomDXIgDN/qa/cidy4HC5i9CKAW55bqN4O2mfvH/8D1Ov4lu2eFGNM
3ruFjViGZM6Rq1qsBfoxvhjSNtJtGojIypmIu0PgfolQqYJ/tYb5y3wFAzu1WP1HZU8WCmPTLON+
s5DzlKyF6A7A1nBoRLNvdMnF+SdJVGNe+1qoa9fmqcxZUSQXBBeAWGSZ3h/dsscbgtxX5El5IEkE
/+MG5TXNl7MFtNZ/s9zh5dIE4xhDSYxc6+kPl/awwulb6CGt370MilcL0Y0yxT/AioZO8rfB0TMU
gcbA7yOUOhiEQJdX8+Z8uln+BHtdCtsAuILGXOxvnr5wg4hR6lRVmkSp1Bu/m5epCIJc9ZCAhJWr
dLIa1tYdS1uMR7+XNwYq62VWs9gOG+ww+JF1lQ3qNZ33xW3Ii803p7+eqXV9mF8NFLavcW2tjfmw
5KUfOGZhRhDpJN4Cj9qYR7gvP5c5/HPusAdC4gA01ye9wWQEwWh+zkY7tAHhrlz+ZKEKeUTwB+aY
7MembshTqcZP4h3Ml+T13aNFQMnH3nwmUDJXSHSBAWUYFoeTROEX906po3rVp1cQIO+e2EW9flbA
qeZffoUcMEM+6ZRqU5G91wzTuAk1F8cqxSwlRLMHujuFtVLT/ikTtxg5xUm1pFE6kGywvJ5jN+p/
T8UegV0spZFNaCGUz26EBClAHiiGJLy21ulJzqxSLDsXDBcvXItFjUpJj1MDGI0Omx7XjCqQ1QtG
ZJ+czcnTSAGb5TAHc0+3eG97qLzzVyRZextYl9smVbrPr0TxQMEiitOJ4XIJ9mwAcUMmTRwJsIVD
TAVXbYJ0oagRg7H8UVvUe6ciI3CyGbQnTfgBIYxF7ONcMaoLccP4RCl873ZOhxWLIx801317CjyY
PQySZ324Fwm4QXyjRnvtqiTQPJgeq93GuufSguGTnc/+kRfiXSlma8RX39S5JjOWos8p4nMlyWiW
AGVJtZE2OqtMjvaSmQChGCJQimAjOZnsDI6cyF0iS9SHdvs83NCp4PZvbbJYkx1W9zWBt1IuLUQh
rXSiJRS1WhwG9/Z58GSF8XUo2p2sXqTGJfqXEFmV7lNHUny5Teo+61YIV8CCjtwYLqOPaaNrYUgd
KNJUb7pYFZ+HOxi+gLUwmdXfPr5Vr1FIGuLAIxVcQEeZHMVxDd4+fVXlPex/YiOho4olG8s+EBMy
EGaqt+vBXFOILo2X8vNKtNKs9YklcGKbzU3ME7N+OBa5qcJkFIZvlS0TjNCQXmgtw12G8rbShDcP
Va2NGLDA0L/DGXory5DX9YYcGOGZHVN3t21jfiSwRcAe07Kig7MIDSutAT5O6uh5FKCPQdLyOv1D
14zHhTOSLJnkHzvWk8BNvtV0j0e+lhbmtXbStbiEmIeXyFcwcGVI/j0H1+Gw1REo81DJlV33WcbW
dlY9habw7l5M+NaAsohwpmH1B/dBSGpHA/ti81zp+QTMJyAVxZai6y5CYqw25496d1kjf88pqGO7
9s+XUI55daGSW+MRWqzAFMq21NnfcC+EdqB86t5rDPlOLcPVfVWslMa+lD+pEJZi9pwz6Jedctxx
JdyiGWkAAX9ZuUeT1gOLqfsBnZNt84W59FUJn6w3uKKcW5QxLwQMQQYjTvvEIideuoA8LDaw/OZS
sqztp96+KVf1harkbcPXNnkQyEvGuZTw5n8PeSLI2Z7dVubFnrUNCePfijz5u4tMguxqOKN56K9x
t16o3bj9FO3kN7OOs6/icMThmEOqx3t+fbe+vjwwB+vI/4H89P3uhqCyhc1wbnpl9vn5lrMA2+iw
5KZZEzSXV+oVWsVNcrg3Ojrwhuhe9GDfdjscq/9cdAInpxuCUIuUu6rhk6scXKdA19nXq4yNJqzR
uH71M9n3cwa4OuIi9SHlNQn4rVLGeJwqrnAdMa+f3vjRFHCNcdlaKkgRPDZr+OTj/SWmWCRV5yx1
FfqSlKsqq5xYfhVfUF+8JRM20+eXe8kFAAi1hQYkqysRnCjyMaaPrjQCYuzvbnrdl0QcQSo6doEw
Tmyv0OkUo0H+i4U8p1qWfK4eFoaNGTj1ka6XVvwPAj/dqYxG1JyeTsgZ4WtamsKT0ADWPRZ/vIoi
NIe9Vbq+NgO6+6IRTNpEdFpkxDZYADAxa33zjsGpAbsIVI7xcx4h1YtTxhOXV8h+iZr+x2gWWChi
PkxRcxLr0WFcQ6u8ZYoQKatAigELiIkW+qUrz9ftjdBwDk9rNnJG4OFsUCI2P5OoJUA4NSZw9E62
+RK02ipNQVnYj0w5UVMcKoN3LSzwnCWgDtovdWOATZIz4IGutw2TnY6gW+s3hFnH4sz5GN1lbJ0r
mfQeQ+X/w7tiN4ELpHDfAm3s/5sdWa6zDXB3NcoSx6v82Y2+E+/ElUprcnxqsrQOVdjv0MuAaIZ/
TgE2zWJG6Sq7OhUE+/Vvo5ReKSOmt2h/0PjDaav+cTGgRCIydUkzrZgFsVQK9kZBvc7U/S5GAiQp
mIFu5HqnzQLrCXMYZG9E5grIyhoAJHIu5OlZ9firE8HYpdPQ//VS7fLcC083iXnGC0rlPpHQvlYL
NYQf6z31gpgmil8GLMHdYVxAMOTUYCQ71Z2A603pY8eT/ciwY4+lwywGsepKektwXLE+DuMYLrBV
9UHt9ukwUTQcAEqCBNSkyz6haJEAdhrnwmibllpC/tykTltw7GyCOi7s+Yy+Jtos0qcltIb/CEzy
7INg7CQ9zp/orqjqpuB5s4chEKdRjduLAR5UZXxEafml9ewq/dtQwukDHtT039Ciq2tD24XhRPqz
+cB0Gu6nA08xqdWO/w8U7GcKt7GmA9C70UJUuo3hmvSK8vdIX80g0mgEanRYgZZy6ano5AZDp53l
g7yW9vsKuNlkeFdM3u9RLG/Pmub1RbnGB04g6VCtbCiTwgvtwks8XoDfd/uKH08udZR3A+MQeKSX
Ny56j/3sNhCY256E2eFUkc0YfV/ztmmaYXbnIhkseE/ncIjXz3q20w6JlF2UrDjY8RdOjE+M1j2O
bGdqHOedUkP6Rvsd/lSkhFtaBgsF64xbNEfFIEr8dCRaRdwMCatywEQOGUdB/HcPd+goI/SnMRDO
vRzBDatFfdCL+j60To3h/RkL4fFGtse+jOORp7ETOhGAKTtyEJ+0VJ0GSarNshwmUiY9XwM3caFt
kUd+mWZz/Xc0m2t8htfKSZp+VeAn1PN83NPltHhggyqbNooqNt+p6G9kQ669MWAS7IydNjceTN4c
5megOVWe1pgZJZWekvl4fsr6Bk59odYyRejJY43GokNks7vyfFparunbtkVRj9Jatj4x6GlDuPwj
sgtYx4RhyxkS5TA2VZhWyU6JfZ9NuV6DxIccjtwps7HjCb4/5mYgcTUQt467KMf3CX8pvKeejpgx
C0kjgc+U5KAC1T+AiiZUJCXTD/3wVbZBTia9zMhO+EfxJy/A7IKbNC/fByA6ti2CQHewiUQHHQY/
ezhpd2A71BqHw2INcYUdxGM8XVYk1Bj7FockYwISFDv3MQcO8+C8OWvcrrDyH7CzC+dzWJSJZY8y
yoaneKuXt0bGAuWxYJ8jMPd51kuZFLh4cdCcdVOYSwWUIdWMcUjd8c+V136HSq2ZFmHrGNeyoMDJ
8J7MUik+rfQ4EFuzGF75VfKuIa6fHdPtaIegFhvCOXsQf2HEOLMJk+4QKqZB5fN1CW4+br4k0f8G
UPxPUgoPm+/NbUezdes3LLJV0130O2+DXHqYgWBdgLRqPGDDPKbudlXx7Eomlcr+Hn8nj0Fqr7OF
6i0YiOzW12gSEmod1Q482TqS/sU3A5lxPcx43ODVtu43ccUE25DdVNFGTO3TrM95pFRg5Ds8ZnXk
fWz50+puLua2uLePsD2HrSrXelJCsmVpMNBZS54zMZcCp9r2+gx4NsK99XbI90oTSYHUzZwTpfZb
7SXE6vqnDyKkd3dIxYB2spLauMPszH109WR6zTzLMDfsZO1OAs5oje7oU9abQTgrF5oUiC/VlMIn
vvpv5moLbRcJRDS2WILEHq1AVns6wDRPKjHxScr1qKzfkicBLQNJyYATt/YXF4B2rlOti4ln7Uq2
YWHX7pwq86lOJyfCIMC3XdxNIrehj9ED4+hEdz9lu0zsEw5KjT03JHanuRYwHUalN/BHXrKyFp8e
I5SVj3TbJe/LUKcHf/NMVi/5tDgUzUQk5YWbeTvyvjBPGIaL7nyUZ6YvBKKamiNpNEqBCozgZ7Ip
u9CvXwh+MeQEhr+dXSIuj3ZpyxjFI1zifxtQ++uK9Pgzs/5z1pVrsGgDzN1NI/tFgXgTPdUxUiDx
8vJbSMt8TJ6Pv78wX8KTeL2qxNCLRp47u5ILXjfXij1odniRfDozNkTt8rQH1Q7Q9SFpq0pjzAYG
4dJEI+KF4mgwYPpFhoDY85DIhzgis/FE03Lnr5J7AIkK7o/QUAQqfr8dmn9dVzGbQPIfwsSkfij7
iy1ll5u3OLtndUoPvu7dsF06ntN29vZwW9UH/gZf2eQNRmrdAkoenfXk0MNguUnPGMSRgsE0UuVO
bR4cRsUMHvETRy3+SQP8p6opXEHQZydGKCm7OeVd88YKor22o7xvcFzsW8A+FEirXgG3RD4+C9Ld
V2FyjJ6AOjyg8d6fCZdwOXb5+dWwFuQwT0DIpSFtYtL4by/p1SXO9di6GIK3tTHEIVKebLRV7HQi
eN7ZAANX0pNr6MaFd7K1uF3sb+zMR2Q4BSHvQ6PHuXkrD7tbDnU2JS7h9ICZV7lsKgGdq41JLvEw
16ZaBzCCGlMgJRiJWtnZxF6GLGmNqF/9VVnp6T3h0y1/XHNvql5y2BGkZveXJ1TuDdW13oJxs0DD
1n8x67gHmR+g71gfqliH8VxAm9FiwY04lix3ZZ91ql2TeORBfUKSbKQMjG0lgATVxQF+0H4sVCER
nPu/iOx/FnesEIR6AupwQ4ypSepcXJ+MXm/ZYx4Pkp2iyR9ufcubFGVlAjYzTp6iJjRVr6d/ms5s
U84ImYeRT/Zr9z4naRVMOC3wh0pU4RQ+7ixUOsFPPEjOn9SuPCUZSl1dkSjGz6IL/WkOwoViidFm
oDjgrl6mlRsjc/BH0AUom2WEw26H/pjrKE46H+gU12Z+fZcjtJvwa9OZPROsNbadJ1oXRb+tAHNG
ELuXjHI2AGQqeGlzLD+P/JLeI6DaTa5QUZSZxEIoIWLGW3QkTx4NvmLQKN2b72kICshjdxngPnJP
U/GzS7VnwHwRTLa9arIFPJb8J8VHz2S+1xmO09vzYOpb9rel6o4oqsIgOLWPu99fbqlHFJKjXcZK
rqwoNpwDtIOFNPbKi3gXMER2qqG8KOFTT4PNi8AYR/xpj0Ms8CphrIbDBlLM4TH4+6Lktcjzt838
VCHM+4Xjo+80Ea2zQLCFnsVJ33cQvAdwuw7+O71UOSnLRn+gaOiF3oEBTnWaX9iU3l+SveC3AhMB
WeOy7HI9JyQDQqELGuCZqGuBowgtYvg0CtdYv8zj/NwW+d/aW43+i0qMNGbZnjYlhKwrpgVlLDOl
AYpK42F2XwN1ffH6CppVkA6wx+YRZDgZ8WskKEMgwStrSIId//U8JROGaKTLy2K9mL3qErqDFNXQ
9WE74WftVx95jHuBQe2XPezgA7fTdA+4nWBYlew6j4wXFgSOgV2sUc51yWyqsKbPnPQAFKEgB/r8
V6HmLdIfhFhJKEvRoocJDqgrFPGlIACwLo5REc0/UT7/9fk8lBzY4bYrPVcljn45eqZwp64e/bjb
/9ROyj7HuaOrexIuF/o3qJOM39CheUxrLQaEEA42++F3Cx1ZEeIyiYeZDQESB19OXPEsHLZ6euEo
DEXvbwBVw9hLRmfCqJWUDa78pScEN+YV6Rp41t4GA3aqo2JSAaNloFWsJXnb+fNlfMo8W5VI9e2x
z6lhqVaeMgfDqC0BwwT9q1/9cMwCGIKKX2l4TfbU29kyqRESrq+aDK9mlrv/CIbl6pphVt7CHumZ
Rorsutr9+5AVdqcuhI9ADJSxW4hoBdxxb1Non54q+MiwwbXiz4uXd1Qvf6YaONd6P8iUndkcVQBo
xRRu4n67hEzn+M0YCEAmWnaoY9Zf3uoI/IMx4Idhtngy9/pqSRiP1QuRoVIrmdJ+H0L26hH6eLoh
5PskGTkBsQ4a3sj6/Sw1HrYg/qzQjPqr4eU/Fo3CJxNir12770DWCOeBEwAD6Pu9X7vPWnY1K8m1
VJUiiFpC1pxdSUvfjQyv6G/oLUhs/i4OAxBd8L4NyeZbb6H18kGfes8updoTDk4r7PikLisYopol
SqZ+bgXIUUTcGNVfP36M/n3vOewJaZz/GKvJfxPBa+u9v2oCo2aN8EzTroWJhHZxOashDcNCLqA9
IWHlm56UmoQVt05ODtHJ1oWHsw3+9etabj6wsb0pZNChPkThx631xroIzT1EWLUW3eOGGBhSgwRt
Db3WnDl672xxmcQX2Ahaf+3/vH8T4DU6FyQ0BO/zWS+/gGIeWYePw01RowYi72Z3ml6JnMgJRQyr
jey1g5yy+mqRBC+PCVlyttWZ2u6WepSFA2Z07MiTVspiPfbr3J9LonxhR8Fo4hNG2P/l++0WfXVX
5zYuW/MpZKZ9WEXEy0amd0YSFkLFffHG37CqsdOsImEh7tqAystu8juHtrXkWF0IiucjcoOhuG5K
efwWhJ+OdscY/uJ7uLmbYDA98sVCzBv3Y7dRnaAsbNVxyi9MF+gvsjOhHI5HCVPE55RrUCr2+v1R
u+FXn7zci0lkdTDtZvG17u4BQgOpORHhRIRanMytqk2QTheJSvTwWCx25s7FN88Nm0d2WVqVTqfE
90ZERb0ZJYi60A1d5zP0HQH2hpNellHmgwuRF1YH+qqdi/HdcyT14IqV8xMnofIE42L8ZZYl2c8u
enTPutsHufltqFvVUm/lGr11NsULADgLB72ZEVf849iCW1IIn+ZRAIZed8iwMa7z+MgmxpAkr+Xp
E1cNoLx03o3JA6CNI5KPgvy+ETaDYi/fkm4AwHxNydOK99ogWBQF0t0u41euAZHSYejlriiuSMac
aoZIO2gNPZJtkMIHrT/ZiAUbOC3qqYm0Umbe0lA2o6lwUnpn53RBdkPYhWK48IuWFkHUzY43ODrZ
KgfnqM5PvzH6Ig7K/YZvS8zNkOjy2hoxK7NNPCWmaPAo0rPy+U+hXdWxJv1DqNvA9awpi8PgCcQ9
maEGwIZ9R1HE4aX5UgPsmquBUZzWZKwdHAV/asfjVHjQRrBH8r2WINMxOvU2AUUILlg98X559dqb
BVYHvQamopErgj/iaMIZoKcU4eZ9WIhqt/aWuOtMJZ0084XfChcZPjzerZ3qlzCh5HeFFCxpX2Vt
T09348cQNJO86cEH4WK97SJMgJI/WQs7FkvR3TWhbyuutvUPSKqLf+OpNTGHD/r5Wrfl4U/1r/Pg
+Ys0gFYe9gsk0rN5QQZCoDjE1CD0UHpZ3uSojl1K9nwYtE+N61pm4PjV2VBidFzZ84uI9H8b3jgS
WA+z5y/djUBS8DBYc1TOPnixg0RECVZt2QB4nxPf1vms2jmOXLV5nURCqWo8A/oTQeaqdZra+AsW
B6EHXn6Iy5PLZ/nuXNVPj7mrew9LWVYYns8zJ2uA1lnpuPWJlcxVOrsGo/4phgUwXL6f/1n9TKLY
y1XHHZry0z2APJ1RSx58V5YdwgtRr06kB+/luvaaSJaexmlq2W9TmW77ICZkykJfr0tSiFRlUTcg
6BmdmW/uBiN+9VwZHv0ZzbjupyzzkBDDab5xoa2BpZJhA6e8FnMEZGCAI4BvwIyDazCg+XqhYK75
Xxlu0FkX2FQ74curJ9MbxvnuxZmB2ytLQO+pdXOcDO+u2UedJH6o1eMmvc7NPdvIdvbmWumFoT52
L62MR+49lSHGzp4l8au3hLVi+BJ+69OKqtKg4I9rgJHsbkIP12jTd6hISmywBSh5haDROA9m/g/Z
VRbqChqDg+aqbtJP/selQYPkYUtwayXPCY8mw62hyvPIG4gd8mf1GsXW9FdXLTpUzp7Cf5JKUXi5
V4YXNqrKWT/Wpbqtv00+hD5aRuzYusCJINC9AZd9vehuV1tVrUSPlFf+ZduBSbmhv0ioBdCHok4U
XjvYuglaKryIIqlCQFnXiWtKH9PBGkHJ0POjlrvt4F7QMPLySP4uQNGx9jo8X9XWKElkBYUhBzVC
QJrArjhYGIviUl7PXKQN/igrc8gzaGm6Hod1P3JEJXDRIL3sQsh+siRDcPTKTBLutzUfh4wJqoZM
0ABdFAiuQ8H8tzZ7cXNPtvWAkXyXKqj9AG41ciBjI5+R0ZRc2djqYlMbs/3OGcy2JP/OKs7Ug0hR
KYzpOqg6Cl4Mbc6OswSO9it+9wP41NPrYkno88QmgJkUyn3SQ+Trx5mNlrEhhaLoL1iqtHyQBTzJ
pMfxwVbjkzFPGGr63ntH+cKNZT/BmgzI8bqOTzOkHCNbT8Kg6JABH0n33xlz2iraEH0EHdYC/PW0
h4iXP/JV+g8I8FU/iGzEN1lc/EnlmxI7Jrg5DeFzTrZ5cp1dh1SWSV3E2/tmxTgVnFV1aBBfghtg
iLZKKCBbwzBRk0fsWU5R4kbHnk0mdQlMvblUkrftZT8MNasn4KcnhlWWxSbxlcGdQSC6pxESTidB
19S1nbXwaDKrm+MRT7mVJjljAKasf265ZGmt0viRis/COqmKivHdsIDfJCNgjlDH6zv2QsZWUa6W
WlJJVKOzg597EtKAzJqfhHct0IF7BUKXdVUBjCR+JpD54Jei4noABmgRnH0LaHVLbZE67GyMn9uO
PZPp2qKk8HowQ3Uiw6d8Y+AElry+3nabWx14L1OPwb+zq5bfAK7FMt2gwXSwQKZ2RvAvb3ofyv72
H6kmDUj+GyUVcxwkdR2iRc3/P/abw2nla08dfpLE0HOtj6/dN6c2S60BsiXYy2Osslwg4SQCwtzG
QISOOsp+8cUJVKvZiRluowayu6UfKyUAXS/Ns/mf6sXabaBTpI2TGTpeVFverLCX3532hvEdhC+C
E3anISFPV4Wl1jHevT/Cq2HJlURdshF00WXd4THM75QQojPvtfOQ7rLg72xd+HyUGOy6Y17ki9Fr
7Dr18HjHtCcTSw3zZ+uUAaSlmaWqZgd28/009o8kncyOYYFKbdVhMs+jyPjR
`protect end_protected

