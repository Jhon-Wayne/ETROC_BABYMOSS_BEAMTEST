

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EErsftIDJVF0m0AzARUB1bTNfa1D65PKFzXVCO3IcVnfdNzarCrieLdbzQivIMAadZGQICQFGhS1
QckM881Qig==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oVVLyVCgNzQviLS1eG+3q0tFr/JK9RCUE5+xAA69a5PzCR+NN1kdZCFY3Hih5lupWCZCqlSR2yxj
T/gFuX/P5PwLJG5+6QmvoI5i4SAxY/rHrl8XM8Kicu6z19CTYp1SPiJ9834l0f0lOlXlTmn836kA
Wgmrcs24F99177fCyOw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kW4owDNqb8AMzEcxlafWfz8koQuLn9mxd/TVVOMuiv8YQ3rvx8K/DGu+WboW7BU9KyEVtBG1MjQH
gJKixZB+7AY25kT/0NwJhM5YyjG4KdEl5DSZuDhsBJip1w/5m+kP4N5/vcsnGSfB2gcc5U+hEZN2
tOLv961hH8596MgBAeOrfvnWa5SH9SROtve5GcJIcP2+J4rtDHR6wFKwG2xp/9kU818nQ53uY3x/
7USyyE73h57I6tiR1+FD47Z14CKQGy+J0+yoYnuxOAdrlqmEtQAPiwIuHmV0R7zwgIucScma6/i1
zxERzOQ0UeBZqrcJuNAcQN3PnQ03sEWGfc4Qwg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iAL6wKTA9iQaAsMi/04OqmErqGG219F3T4DtEhjCOkAVV5xns/q62D9v80Yu9LkL7GOPStNaimH0
0fLZZNbLN9aXY+LXsOjLmXKIRD1NJHFD/6y4EmfJhRxv4wTaSxMi35TYjtTPOpBQ9f3kiGqvET6q
oTK12b3zP6bRyeM2ZbhHWjG88vLFxPuV0/g08KIWxnwsizoJce9xWIbPH46yn/atycdYeI6hNlt4
AsWLZjzzPTaNgwoNSmXe6Z/iHwOsFgDluZ4wunNLVxH5Ru3KpxGf9jGPoEfbj76tqe2kxC3Whmb2
TOD3EfgrtAPEX3iiwhkJ68FGwrBXobVCgJLrLQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AYk0GVXSV/oBWSOxjuGlD2oLlqIfBX5t16vozwXg1+siZJZSMUHEbzptzgNoTGyAuDaMihDY3BLO
EtrWbX/36HzF6OYvwf5POdt/VXMiD/WmbkoqBGEm8hBrg/s//Xc8uwTP0aCjxNObZuBko/Q25mgQ
30NgIumW8FqCkhPd5zaKXjVEqWRkZbVy3s9drUMCg7SmsRWiURkSk2U7gJHgxqNeqEvn/U3HMsD5
przVbreKAnJv/RzsnAueSJ7se+zz3ea7TcdOm8FG4lJPtFHb6jvhIcFQ6qftny2xQ/73EGrSBx8k
emkzKeZp3UgSKQV+dZEMJkjg6+hPhExCSG3ddw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Z2aYnMPHx9JY2YhtHwU80KMSOWZwPC6TzLQf1GQQ4Vnr361DuLoPMu0MbOnkBR90QGDH/qF7P5Cr
Ly2yiYO0/eJzmgzCpSyJ27rzee68zFBRRDPmlOAN8FHZvnbWm8t3N4kjdk2vzG0NcvKGeDmWVBg8
WX1YKAu49GjIv50pk7s=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZhLzhPI8pgMrQMSYddC1+njODiKwQHec1wBB4U5W8/l4gRoB3jhisEMfFb5EoL+ePeazVA8YvpBO
fy15vYUdxOsCKx+vVBouvB0iJLQJ7MJ2yB0Atezf8W/dnulTtecMT4xYThtmLmUoLpjc/XY+sv5+
kYuBtkUrJcr6xJNsQtV8JIkAU/9rh0McphkltAYVfKvFQQ4iPL6Vn52nStdWLo/EzZRGxkA2w3hx
RxGGI0fCa662AzFgfo3+9jW4FVA/MfRfrEnMa/qSzvX29NQHmhsMx87TbESpFUhf8rcOf4pNxnvZ
Kz+Rm+SekS5sOFDAnkaGJ2fOU9v6YhYC3w3/eA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
zgFw5JI6UUvwBouz+903b+zCQVAqCLP+cWXE6KoMLY26n43iueLvEr9YpeXyk4vKOq2NtbGH/zDs
iliOzbPfIBfZXNscyaklCZaa2EGwF33MjBNZZ1A/rtCCbDyk4+xk5elKdXnlg9OCS/dcnPWTj/TL
j7uBEClOzu6naIrLfbKtkNvg2xF/HGDbzomKgvgq8ln7M8hwBHzSuCTJoNORQuxMa2WrbHKqPGiK
qlh1oEPYtQ9Ywbv1BKZNxhU2V/sPYhD0JQxZTG1zCLTnOaQWyjVARg2Ptcm+B3HkC/FfLKE66UjM
nj2tINsjs8kGS4dCqIdM7G6p3nZJo06EwZLxeHgFcESmaTVsRnpNfCBfp33LtDjcCCC7aQbCQ7cp
xYCnugYh2H3hz7i8CZf/EWIh+KTw3eGRFodsNmLbOKD9/mHDbkysj2s1saG7hVw46IzRr3Ex5J2C
K7TkPz3na84zO79V9OMuC+qseZyIkjdt0mAqwb106libYhFgp/eB0R2psvw7Ue0DEG2gjdbLdl9e
WRR1YhYjWVGIZbUmi0/lfr9RL7SaH7V+b42TeEeShfxyr/yfqfLBnoR7vYtJw5t+Se/O3WsEawMp
sHkJFgpKkpilR70sMzf4YLJfDvBjJrGAthPAjZfB113Zv7qs4kMbQPXc460ZWa5beBCNrz9rrkCD
v3f4wsF4r4+o5pEEgs0UPSQvR46MBG58BRsRkHdI3nU3uLubEU9C+U1MVHsdrpdY3HRI/wcPvuey
Epg5uV3YqguQIo8YDSchHXfbaUyrIVgQaMNlJ6yTIc8QKBLC/HPNFK94G80N83wqcP1GU+V8SM6t
ZhiWLbRBwvFwLpu/REa/TDAR8AEaHrD86CM6vLCKGEiwlFrBAW3GYurAFUjrlF8BKkV66KnQ/eo6
nnRrKzH5XhEDoz/7+XxgOrVqQx1vt7ShsCJTt3KJRedTNhxQZPvatEYA2xxdlouRLeI6q9VUZkj/
TyUt9obCaWMtfxkYOK8qSZmYnTvmWPL3GU9Zf714GIHUxUbzZI88JZniJd6UEu+Sc50RojxOWj5q
LlOu3oRTRUDzom6rQxDq+XMnKY4yfAWmDDa8sbdIr86nOfS4l2AkQACVIpGbzYzJiXzI2TXdU2BN
dwDMPXMg4LziasAGc6QJGBbhmbRHOIrhTusizzUfbBSSeOSBLJxGiVKmJHgCS6c3zIW9OTZ9r/2z
HEAezFENSC04nk1WELrNgRRniwcC8Mu04M2CC3OLX31ZRr6sPn2NUV8jKmWT7TkuiMukPRfAY9++
Z6KNg5DxgauAnTjpp1XfHRIUmnI1l6kWeOvja4XZFQE7FIsYnwHkEWGZh3hRp3CqCiNEAtSBwaoE
WGTfVChoMKhhLnRUd/7qddFh8E9YeMN9EJFkFvm9n5lAQsQ4B8ovoA/BoyXl0dxhj+5zFsEj5cNH
zi7m7ewgGgdZcqQSL8cLT1TilGQ/cTs84mEd+7QdwQoruiDJTSwh5vTQg8vmhsubL1FVZdHFSJgY
XKNQSeJm8zNMysZoKX9cOIQlI9C5r/WFDHRk2hp9SFNAaHiXDfFcF9CWjjxij61x8UR+qBFTpDHq
dBlfT0ixJDfIWGhMf9gSfsonJtlDERax7s8rpOfRmdGJ/pLr9B6U5KxgjD0PatLMNH1fF40ck+We
wpzDwnaDX1xfbq5ojNtm4D71Ki+h36OQgIKYBuXkzlSQ3Lx6WkFP5/D1VGq2D10n/HbjxF4jeqWj
6w0LrI4av62FQehUgn9XjEvwr1EibxiogbhVhJQQSAZR224PE45o9D0AuoFi5pU/dnfSzGxNhFbd
kK5n8Vc/kshH8WGqiRqp2sxDDGT++3FU/TuL4y98Tj8H1hZ1HeXNpCF3Jm+IxaLzsKkCHoEiSPjy
O2orh894oPf7ejwMFVoB7pmGiq5mWxMHrEPmsqY44bbIhr1aZp/Q0AWAZXKCnHG5ZJQe1n3kv/NU
K1FPt278O9+pFcG308s480LPu2mNixVk+4Zb7HCf99HPzfjFAMT8eBZiVyqN3Wzxguv6tbshlgom
bXyH5uCkwUKonF/SOpahtfafv3osi8+pjrQfSFA5SAjeyNytPHST5mYnf/KeRWTzaXzyeQMufxzV
dEo1i48i+DXW6enRMggScM/nC87+LXPomXW/yWw33DDAxGiefYkpLOJgTADM8Qs6tmHLSHUxnP/c
0V8gpXb79okoabaj5BoZ5NY9HLlqnwyhewLL6ug9G/GkVeXLIPeV7avk0V30JTtKdoNM9BaUeMZG
5mlVJBaL4Nlx3r7DT3isyEXparLQdC6rVjq2xINitH08nWl0mTGIQlQoGY8X3PoP+Tbrw5ry92+C
KjnHlV4fle6c0e9jwq0h33Mgjmdztr8b2tspYYI6W5WQ8SMq2bvX8kAYa9f16A9I66tH7caH2kJR
GAClYtSzZNjsSri1e1Qr1THd6mQlgmBM4YPXOT9bg180lZDEvaveEB/OLRBf4QfD8uJ2CvKf8MAk
Na+7sen3nxTH3Znhos6uGlvckEEDWXNeMdoQiZVNNyPXUB6mTjOzvtMDiCFbrCxAtTM1Pra/0RsQ
ZDur0SF9eFOz9mItfB6gb2URGFtM8rZqXp8iSpUcRygMbdsxbToaxASNniHNUUF9Nl3LcDTBwS0F
hFMeW8sq4ehMK0dYvQdLRcspx0fl0XC6N1mZhxtkUP7APzAZ4MhEv9HQFSEKCNr5IuastTrV4lqQ
jg7TFYiyJwTbIxVIxwmg+3AhUDFSbwAJp5V703HOHMqIpUsUKeBV+VNV4qsUF4YdUKSOsmJdSfiL
opQo5h5TLsQgA3c1Dq/5SPS+7lEcjpRdDBZuFVZOMXqWvFRuwx+TvEoiHc1DWQMX9oc0s5mPOo/1
st+uGVgqxD902UJ+lyAdsN+yedkYbzBJtnwi4Ed+E6nzZf/NTvkLC4aOH4WDhhrwac+ZYNuk5+Pm
5pM0HfUJWOogMWmuD4P2gyEx+n/a4Gv1j0hwfJ1AXQlqz/OTZGb6gdKBKbFHL7TsHDeJx0liR++M
t/xuM649UuTKjXPXqR+980Q3eK571SHGlvDmCYeM8mpUuKLpwQ1gSM2P0dcl6K3RxX31/67v82ys
Hi5hnnfI0JveBE3Ud32Qm5NgRipnV3vtad/6CjPzjTLyi9oUAfoGNsLRe41FfyoxLuI9RwakX9mG
bH8cwJzQWqE7lQ5Hx2JKWGNItUN3lhKAE55EaYyZcclA0BZFIWBm/c869+dKimVWZMJfSkvM9KIT
AcnuqkNogNYihSsaGLN9SQOtNZxSjtAcOU+m/xV4bg53/wd0rdoUh545ZrAF/jVU9e01IGJpCmi/
Eqmd+WL8waxLYpYYgu8a+JEFrrGnCiFoFfCET6I+6GppLkUUNRwYIz4AfWr5AfKOH+Zfr2cTw7h4
xxbRVlmO6yr7XjEFLX4fcLvtthRaYtimn4FhIOVEf26Y/OYpWhkgxzGiqp86pk30nzmsaIGFrBu8
CLlBZ3crF9jf890ML0UEvbOVx8qXX8ViqlGa90ph5N99UQ6HPTI5BdTmPNayCVxHK4imaJEtzWsB
dThzP5VXNicC5svVVgw4/RyBUzTzzwRGNfqF5TB49RfEFLQ9pOwf//B1cKbaOcjHtqxCvLof6s98
qBbKaNbFn8t3rSarpo4+xf3BQrPnuWQ3ErMk/TVWmIu91zS1khaeX+F5Ddc24Xb5HXucAd4mlF6m
Y+vanC5AUMRaAShkVMPncJQWW7UNxcGVyP6vyhy/pIlKNEBYZSIwcWkgDtAWY2OUfjJo50OMglfq
9N6cZwTpkNR33jqnbGdhaR0p/vJjDH1BOshjpo1feWgHGkwriqIFVq14GChrUqpH2yQLov3NsVnH
PLSfcN+KQ4KMRqX0ibmIaj3nhnT9f1xA1bBa/t3tEoheqWrxF7q5c8uh1Fe6SIok/AyG4k90JHXK
9GlIHEOrbHrdJcWGqSmeTYGSbE846XmcYqW5MbitWbsj6dQ4L2QosGDdb27v9Pk4ASXyFtxu4xya
MekQWswToaeh4bxYL+dTGTbC+42YDfysL1wbnBNkZcVXOWW7u+GpWVkZCqzvdUT0yX+vfZfFCqMn
sVGICYVgnmVScM3+CqHJebDBlq8YgaWDR8TwZj5XTYRKJfLU90caeX3NsedFfHJbXGEATV1WuwQG
Z484N7G0oultLCFzsNQWlqAWMyzeQahHOUpls56H6TPqXr+EYz8Rb8K1HKASfw7/PRwVtDTJ6o89
yZgTX8W67XW4R0PyzhbSNqbXom/VGjsCeSBdEXR2/7iQqMdimVqP+NfukM6+rrH3P+iuV1Lr/WFF
Co0tJxmQlsKB8DSP1IwhqX7zyc7HQNNzEMCF055KLv9mqZ0llCr277FCr8YYf4NF0jHofzzghz0K
qIuvmvJ2p1OFo4PZh/qDBR6Az+tbwG4JX32bCCDvRY1tn0App7fq6yHnZOjGvcezQ+A3FdsSB2AN
BqY3xZqsF7DqK/tZpaxaTyAp1OFNGH1hNDY7AceWMrCSCbrkBpkzLc79/L4ptHqfyLfNKeGNydfX
ThwvcvWMnAp+j/ig0tTR3JNfT0pxU9DctQh7O+k/Ggwxd7nur43IhXry258cmQunSLCAbXsgZ1zR
yN5SdM7R0SKUsvXtJIdmmyJvJpCj4/aHTQd8NrR/PZAh58BewFJoTiRbtsf+y7Ge7CFg8c+A+eus
98fhIZ5suxQTqW9AhU2c/aGLKdSsVwXXbW0KnNQZg22kiAJLU1jHaKLGfoQ87W259dP86yoq83/L
IqRxGjIU4l8XR4kcAUH6YWm0WVTFoOZ8BB8guhbsN6wTn7+hfrecv956BNE73et0yEyMqaJLrDFW
Z82KmWA6hfebPnEtJ82cgy8/gMboI+qLzL/b1bOGigVTX456TddWfGptTT4B4KO9kaViADgtjGt+
St5FnTLjsJjR5jhc8wxS32YZe7tI5DOTdSFrsjHaa6I2yxDlRcqIYTmuxIeGXmV9te7oz9HMWrcr
m8Y+BMy0AyblFalrjej+7G23l3+rJWtwcxrok09QK8gdDz2kbv9sSR1NfZgU8qhYuLZIsHQDacSM
A7yspjw/r2Q7/ZnZc5Qr3zgYaKI508n19Z+v172QfGHHsR2BCMZrvEo0zjj6DurMz0aOVCWFVjja
i1rr8VpNVCEPZYwoTbTRpq6ux/TIbXEUIfz0SR9mkE/14Vj0WS1ibqrvHmeaMe/ZcNzeJqlt49De
k/f07tr6uloGuADrv0Jgpq2QW+zIOxsClye5f7W3jSPqqxhwKciJDenTJiMuPf7dCXR8pjvUo4Mq
eMAdfWNa8x6d0ZlmeIrDhtE5G+yY6MlJjcqCEY6ZTrBlKKThqsqLgzMnhlH23qmUVAGcBe4PF5ce
/aZQIEjdsX/gaAhWF6H85GLRnw0nc0CrELqcqi1WqcJvAtSZACyhVzZssrP0xbfnMnwjniUTJjeV
SD952fyaW5mtWgnYq6tG3htHZ4NPX/F+uUsNDOcMixcd3Xzolhmrh8QplteJYm78bKYTupCbNXWW
U6/zwMRtT1Xxsw9UKzjiigDY77v5p4m4Z8WERh2NGB9P3f5n529TZeuo/BLdrEJdeZBgnXhxhLIN
hTIuxNsxUEvQ2Lwp1GZR8lqZsvRdvwRbp91ubVJVeHfDtg3dUyMosUQcJvjOvSdN/vdwuQCzhj+w
AiYY9eJDfzUh0tJqaMF4No5QTCRGZDYl0LqqrgOxGVxsP7I4zD4AVxzHVXsRKtK/aSWMw9EIvNMD
4RRywcU8xQ7hIJaTC4hUFXZ54JnJvL0iEV29ehYWb7IP6gelaZKfjkv5QqYHxz62/nfIAunI/tJS
yVfgEng/aFWc2QgmHCrFZp8vsjs6Gldt0VXkeKNJMcaM0AWtstqMi12Aa/OZSQy32l76EnFafhpP
U8gyLQrTypW5+zLos312oRoJjJ4uNf4lvLNgfYlO1fhNQa/2oTfijBCNfT+S+TF8Jj64yC0sjeiL
kTnh+j1vSQ/Cb2OLbxfKZkqvmomjox+n3iNsaz7f23Rmnzo7goJUgTmPLejRP1UqsAzDFrWoKNYF
eazkBl5hrctT3h+QaSXaGFDL0v4RxJ36v7DDImlHmMtf2k7Z9k+SAnvdyP4ZL0Dric7cSlFBnapD
1lRvATGR0j/i6HkUHYSCP9J5LFuQ0lmu4kzGPWOA5q+lV//jYXPxNwImaKPmpH7Ek/UdIB9UoWzu
dEsyhfqmMvWFNDtrRszWQOX8RFfUAXMF8tHcoj3iqbjyfZ+pepAwiUDqk2673XNAh4eLoT7YxtJm
UfTbqC44Ja7V4SwvIgQux0pyMmgcyMv9slAFIghkBMF3WiAcIWTlEq0euVNgAQmdfRSEZ+p5IZ93
mFGAAG5SHiYptJZN2bpGSfGlhDbhFGOKs//kI5/SEIWYdO0xKJkH279uxAdxI5e33cHJRe864EHz
zfVpkgLus5QE0WL9xP82n0l1ZccfRfggvGyy8CdVR+7Ap7S+Afz5UvGf9KGoOO6dYYV7ouoPQ1Y/
mShfOB/6Wnm9ApRLrB6OHafdLOm1Kw+4V/Z64bO+C28EPAdj3REysWnGgYRu1ZjFNxXaldAbppWJ
9TloCxG1eMm3kxAubrMpv6M18lAUSL+1qBUNXwushUQjJx6LXjGzlbUsMj9ZOR9DMOGqA3lGyxCv
9ILDSa2VDd3NIzkdauk7KHj2Th/kU7rsBRsaBvZTN6SEm2WlTMyafjA1N8hLPMzRsUuk5c9zZ5HU
h8qR3heWbREZydHpc10xscpHftVjRgWPCdOCUEJiFLKgmhJDKdQ4EPqnqEP/h90z/UK1fISF+d5J
xdyms2J152Y1qXI6uqeKuXdd+kw5EoZInppV21QRJ1sSGJca0LlOYCeBSUIX8L6xiCNaj45hK+EM
CL0a0gN/c3iH8sAgfdP3WBSW24U6p9nZpb45L9sxNVUpe+J/D/3a/ZQCMaMfyC2H9JwDFqZkx2/o
kLhR61EYn1R7vIDwqxmoplhTWN0ikwSZexP3RmMO+GG8jc2QpCwm6ZRlYhqfoe0d+3vETMdngYak
gqzoaJXpAQ07p/hu+kxZYxCWEngz24ldCTwdMGaDoBDQ7B5/JRkJxj4bQ8MywBf1/S8TUceknmGz
+zmvx9amFF+HPqJtSQsno9gEeIvMkBhclBf2c+WqFIGgZnINxSo0fWfd7kxu7Q6kt2pTIlgsuIa4
y2kThdkVuk/1wlSQNxL9Up3GarmPVbdMB5OGz1YQfuNoikmrZ90xWIQVYaon3XI4nwUlrrr1ZRN2
gKmt5pUuwwZBKZ5kPR5gyX3PiAqOpQAhG1GBJLNbpH/KJY2nc/vBwdLJ03q/oTF68rOdC16CyGAj
mTENfnJvcOBPazqjGV8gk+tR3ubDiWW8Dz6eXS/dmJ79ismCXu6wrY9nYDUC8MhenRgYy+l2IfgE
H4msNVQ3cmFNdzk3VmHHZQQDshFZauuxX0eXErLSGMad3JnSOu4asDbEf0n+MK6s6NMkL/46ed3W
tHHvGo1payG8xMbv1eoLMWvmCDL5Re91ib0ZEdS8hEk4CmfnvovL+gameWSMR9lzDcW+hqiyvCUG
BqCmGU94fxIPQbW2s6V26BFlr7vjdqYp1oe2WB7U/4AcwHFKd5S5bACRz5LjAJF8F/HSpxN4ZLGS
Iaqlc56eQMYtyVis1JCdxR4IFy7suRqarXyVfLm3qJl+I+yG49CnC27Dyo3f60Kxn1T64oNfvwCA
6Gz1zH+AHA0mvDg5ukmWQ2An02k7EOgSjXJgYFQAtYhNRavnEDnTK66ZjSfU4WFWZaPcrki0s9MX
C1sDy55SE6Xt6p76DqqhEMAAqBoV1frUF8nvap/ztf/gW3rfusddVaNHlI3b04IqQG7W+awW11S0
Kt+CP7QjbK2a5lXxNlfJjNzZKNH7ymlFtXGi04WcyjCGL927gy7Cj+QWGx+4eil+EG2QcvhpmC3J
e7TiCvha8tYxDmBHv+QYHs1tWBJPMA2alPvlmctTzGuSr6G0dxf2Ca7aC5mMah+K7u8vP+qIlplL
02Po5+8j5cUxenhf/5WLwQRgRV3MA5ej9io94dFJosl8312v9kYy8jszs+zbypFhkoAKpV5bauv+
B9CQ/yFV7Vh3Z5yKVuwmkRQQApyUNGTJWoj3oQUBERuYusjSCEv9Tf8l1vjNE4qKfkDPHPzzZrwp
Q0yd6ELHDpL7ne/IYhJBb2l483OsGHWJ6+e9czyuauZBxTYLKTu7aRW1IlAwu7Ah33ixHh2VRp2n
5RzjxWCNEZamhE5mBnDZnaQ+VhuINaDSaRkw0acUdWRhubVHd7M+0Vl+pVX7E7ct1OnvE1Dpbg4l
fhPgrxFifpzFmGfD2iL1ucCRnSPBWn9OI1Ybqqu3sA4q3mlU75bLVu0kEKkWagMqYc//4221WQOb
v49pprfU80+PZFpAul73jWFI2x9RH7SeCVaaBduCPqnAd+I1pcco4+Ww2x515GV7cSNCAgeG3lbS
rVdfryO6j4824tbbIYmgUAavMEffxMUdMKXadViqb+IM9YLPWwOvhdTM+SbeWSrRAUPpOuXvZR0n
Ihsvk0uBNnAYW0yr4wJoptg9Dt56R+vmrcn1ctUF3AJKoksA45bhHy8dYN9O5rKxRRvuYgjpn3um
mZ515QMljllLnZGolpquLMCeVtGG65VApsNV6yLcfV88oekG6MMyvdDNLuXhmhQ1N1KlS/2jyG1v
PLSfNH7kT2eQMk56Zen0GxvU60zLzMPuqBitNQuwmjZyKwYbicBvhPRILFKRvDdLw6ZOU32NIg3J
TyTnXLqJ6PP+iXYuqxGkQlgfzwdmppMcs3tXSCopiVHV3WEfBQ6dokLHUDjd7UQJIgiAK2HmnOrq
IxqxqksQsYwbiSJ9B7hlcChhfRPbFwKVCZTf5MhxJfTG9maJkDEnZVzcMydbC+9pvn+9JW7iIpPQ
mEd+ZL2aj1ju/ascI6OLlKZhqRE8W946T9uMqXxYqMu7btt35QsvzQro7n1CA6L7CzO4YsvKhvnJ
Clk6u6iVfCuH6vPRAu5u50WYqPvxMvRjtVBSz373YZbSLlV8W6XHewwV8E6DYixwN2Ee/P/nK5WU
gtoOmRpmDaiKVG35oIl2bLOTfEqGckrVhXtqHAR63pyJGdLh91A96CvamAWUFJeuUizkqi+kGa1a
KKQapqmXDKr+6XNN8bn9w8TNnbwT2a1I8ORuV0ypfxf6SsqkpDsKgS3nETJxhJcPFz49WbysllnC
cCnQvB5eYV1AIAoqpAOs96JX4bxMnSwxesVaMOhdWTl/jDsyvNsyku7jpV21JMevIuTq6/jHtf+t
ugJbuF34+sBT2M1eMz2Wlwozn9QJRAfHRGb3xksqog6Pyk29z3sGW4od6hDGsUBZ32by/vqXQRLE
SqQfrPCy8BztwkWYOf0fBudQLzJCrLNQStn+7kOOBejIjKb0/NPVG1vmEIAHOII+0MBc1r1CrKsg
hEdM181t2OAdMIggGclAKuDJNKV1h2z9ZH4Ip4exYFNtL9GD4GDRMF5qZMg+4DS9FJvxpDxaPkYH
tJDLoM2Q6+tOuLy94pV+Al02MtQVYWJ+opg2s3ynKY09Dj1uRrQTW+e0QWKGP8AAdAB8BhvST+6E
AwAc+BnFkq4iq3Ctt2W/IfhU1+zK1N+8nRdjiarCyUszrYJ1FiWkaEjn+OoWS13xS21lLPlZNagw
JfaR4tSL8zKQy4FdAEyiyWSPEBzoupet0Kp5Bj3vOU7yuh+uH6rtt2i3aRWITjoT7/lbC9+S9nlg
6iqpocnnxq7BGH6d9Btk4nLocVrafY3jF4yQHE2oihFgJyIk0Zz/3Jq70u/tOO9VFgfZ/ceDRn8+
IrwwGgKq3I49lbAaOEMVlfl3I4QkS0yr2rDYoxR97vOZ69WdnwTVqISj8g53YtwblB11vTHGxjOJ
iVjOjTonhposbuBH/zusB5zxapwV/FGGdC6/VkCiLkfklLJP9psRasLDVYVfB3E4igBodB+FKMDI
sf4+WR+80+YLrjxr5wDfq6mI0FOwAK6MJtcvFQ2dxjVSf2UrERFV7G117e/QVruejHXpzppSYZ65
FGfV8sVyAbgQOLOUIS4o9EqlzTLA+bC+55WmzdRxBhSXubg5gvUm17bRqjSNqNgXDJhqcYzsKApF
ut6MiiAV7aNDaSbQgsxo/yxNDo38VZcVBkC4ibJOqYmPFFbHZiBcDzy6ZUzs0l/9/GcoAfe8vP3O
19Cg7hT9J7E6hXXfcxLNM6MhLqNyrYjF7O+UAAhsB3wgEH3X7tAk+AgmNQRcag5I00kELX7Sq19l
/f4g26rv+yG5JqwzDqnv6undSYxgsqPhhiN65adWpy/f/eqh7f3YMaobZ3VqujR1C2M1lqVrXOAQ
2UkHefFirkf5n/IW+NGqxJQOMMFp4RL47HVDdqYRdDaDcRN3Iw/RbP2XYBD87axfOrFMRXG5xvUG
g+iRTWzLtgb9DrFE/BYp3KNLd9nqHNcVrGSDappSFZrz2d83zjejQPVfnVK2shcubcqsH/oRucSG
miIJO8EPrE2W1P82/MNQHkYUp/LmYTedyyaC0UyqAsRKLi1mjTpNA8TQ3KUVIg/rLGGAwTCLeGAT
PSPHdfvIFeZ12SpFv+r4bJkeuEsfc062abP4UnOxscr5clEnXXjV7BcAj3oTe2IVB7KkJNN5jhal
yivjVD9gaLPZj3obPZalg6y3z3nRqq+YtQK6atTpDJICF+9IwWS7wyGt95w4QiB7pbFL+3C5MpAl
bQtXxfUkj05fF9XgChfASWv0f+f+b/RmBolgGWpXllyeXejiw35uA6NMcOLt5ghzrkhiR/EC5qaD
xUDGke6tsEz3k8YhIgYzo6pThY4XUypcnpsjkQBgQC18/dR5rFQ+ha6UuiPGdKSH3QwmW2HkoRZ9
JXBmFfYSE1awk7CxaBhgP91u4/VICIK7rIIE0sj01mpmGUAlzn48GedKMb840EXag5vOkUhwXybU
jNRd5ofcuvOaB/BtLXhgdZTng+7I3bKdnSXqOPB246eaFwFAmT/wYaC97TJ/FFJG+b2gj7elmErf
sLJNe0u80sKulR3ahoL8RyXuWdSaT/1hSEGef5S0Lul3p+m4jW2os1Xwf6RGntOKzTDDDWuaj7Lb
Vra6FI7r7r/DNd+JOYdroHzuqTldsiyHsAVWSv6dRvofYuaCxDUl+XX0OCDUkk7hYxnqDKqpthbs
gt/IMvk9iZYzawq97KbPRnb7VER2bB7NHEe13yI17QFz6vcOzdcD6ghQk9c6SDuTn2Vg6oZbB0EH
32ITpg2b4tAqYkThuX7FL40zJriUdvGq+Im2nWFHhsZktPSKBYaUN8reFSKLAQLcfqH/tLxGWkPT
bbDJpwuMf9WVwpOgiuaMh9Bz1eUmqo3p6jr+AYei+NAMsODhKSgBKzySJ3/+57iPJZ2AYq1csyKZ
2ZzjfY0npbnFtCPmZ2PkFC6Cbbq+h1qvkzHNz+tE7scpuNl4aPXN66PRzbZ5rkSPBuY2A7ayGDK6
5CpqgeWjB0wHqggtASd1PQjdv8lJVeQLmzNJr6zr5Fb4Y2dcJeo1ukLolEoPaoxZE0+5EiL/2UAA
WzV16q7xL6GuDb8rhRy4MYzT2vhfCMRcjkG9kYEcNUWrD03oTMR/sJ7tE0kYkq9AoWf3/eY9BRMe
3uJO11yAPmYG38jaFHMACCs7vzT/CEc0H0YcjACpN01mUlon+PS+QYsqCTuZ9KJaenDzfhCrGapp
bHnxLIqE5UbpYrzSu/RkeuyFKR/LuFKE5HyVRScfJnzHODfB5jjA1siHWqs2gwhwQG2BSxDVqFkk
EyQwF3BoHk3k3bUSBhphgYya5t9JMML6fUMfVAjV3XyGfnnV3oglW/CiBj3PyUJTc3LoY4Nktlcq
Ou9hW8EwVd3LTo9ls/dB2I8Ky/wQ+HtUR4ItU8BH+pwM7k5KggNAYzcpIBBgGzeRrATsjpCODo7d
1f4myObgINt1rbMbAQSDw+9xIZ0HifaN8Adj1/gtNI0O9qiXpZO2yy3phtX4zizq+VPf6UIBj0AQ
5471mAZYo1WrwBoAjut5e1sfX+XgE9n3Z8Z3PyaHDgEDkT+t37fKj4Y77jyrS5bMyfj1EGllYKU7
V1cyWXqIcGXYk7+Zg5jEWWFmEMV91e/uJ3m3L74abUoWZt5+t7G1pVAcpOcK5wpn+GPwKUFQ/UvO
w3NOm19PMN9PeSQ1/vcFAueENAV3hDMqjKKymrQ7Yz2nOE1vuE4yIhx5VF5uxl92JAquRt1nwDzs
a8l/OnMk+Hx4G54M68wHBvk6O7jc+/MLqWVwobXqHRDkakjKeDrILMF8qP5Cq8hTrmPCxAW9Nmdn
NP12H5oheh8mwTxwofzPjvk2vdGwVZPsjjyZ/LRpJxIahO9r5oqVne1eTsVJYC/4BteVXMrxU7GN
cGpmo8o1gUMeatNjRfTsz7kVCF6qMEB/1ctvpmPJXBujc3Texla0M8/EBkdhzk9/odjjt/5wzEhl
fHr7n3YqUghXSWXCW+NRKVQwhxdEOa9/mNenrE7rkuEmvROX/s3+Mp0K4tphA0SdASdR35uKJ++H
wJ6I/mbdRvADkADxtVt35Z5pBQv+08uKEpa6E/XGWNvKOv0KJuogwhhQTXNeQvrgYRTxolRayo6l
DNoc1ML0GGk5bu1PgswrRdirjwMFLk5saehSQhXe44BG54NlhoDx7BqIUIuEY2XZEcp66gYpLcYq
A97kgLRl7L30S4MIL/5dWHAZPwviuf7THTgn5/crYpsdht6Maf4czM1vPRwIMTrf41c0DqPsbyaH
ZigaRSrZkDFJr2MHPcbC+tdOnH7dr2PMP1/SLH+W8eo3RCB7j+cfi133vV1zZ17PmKpxOrjQxA8P
paRHLq3d3N8JmAw99bMEIjFrCM8cdq7mQioaqr52Wg5sAbnmg3vBDNfN+YpPfPvUNJrdSqSQL/H8
kXAEfRfCL7rG96KygrtzzMMD6WDQX30Zp42KG4IP/Ngydwex9TP0s3pB8l9iNgwUhVkXpTfqC/Jo
JDxgbxW8gP6chDGIMuhnP0iWZzb++H+qNgNmyldc4lNKAJQTeYJE6giWMIAPGNDbumEZdu4eSaGI
J7iFqYoQzmB4/yzMG/Xkxoxcg2pFm41B22F3yrtyjepZGL5NJCYqdRN7Ych/zFGfTNps8WS1VuoF
rJymbQWPaw1B6V/2S/Qk7xyOawgfOWhnFzw026iXEcjpvG1Mzrh5j8Cl2qrWJB6zjikjQQKAfs0X
6TXPoVPS+Q8Y0JmLExU73CUZT4gm5DsQ7wIoxTCcSzFGxRCUddoKUw89en8BJYG8bVniwGyJIxbw
6dZ8T6RFVXbgXQG2saVS3BGHSw4kAvAWWNKyCXyyTyxOk+SQFnVK9Upz7GkLmArpwg9eIaw5PDkl
ysPwlCExZL9mEdAts2lExyMKfQpRDo7WTGvTP2LlFp80lGZ0CigWpsP4+34EcdcZMgBFGbV5eQQt
bkFSZXenkLM3FLS59XB26h9RVnubvqxrpt+SULosVDARoI9OfK7mxcpFNcYI4PzXMQ07BIFEFeLG
TrRXgI6Zw9DyG6yqqRS6IAtC0C7vbtTtXZf9xkKFqvmi9YnYM4GW1Pj3d4VwRxUTXI1fpVpnYOxp
0ZvpWGudfSTDicWIc5H+ocV5Ixlyaj65mnA0scybL435Oow3xrK8bZf8dIinl8tG3XlS14RbQvO2
JKQ6DODNCPujnCBgUWlymENVKwNEmY5O40Z7o2q9InpNlw6q+FDXLqLaQRqW8Ks+hOAw3ldbmDGz
E3t2hKMCQCFbyUoyT2md1+8u8UGyShcQkomKH6w2BWHpw5Ho9rp2M8TeTtuqXZ2OlCffJDZKigjc
+7D3TrUhWfSrgB31psyAusg6ZsRDCJplgn7GbmCoZ2HrlIcwFeM86sbVo7F+H6zxU6vG7tDA7Yiv
mPvLfs9hpeP9c0lEgpLMTyo3Fdulp+XMW1e8NwfgGSFn1Sy0WIwBDhVaKE3eN/JRVXdEBwJ230kz
a/Bp5QObKce5KBL8tpyN9QxrOLufKVhzl/JVd+Fy97j8kvC/xrawM3E+nmaYSKEM9oBfcLKNBBrz
Ra6u0QyDI0OPHQd6fZxkUwut7QZ9HJsPhe8d6/Aveu3BdS/nhDGuCOQa36nm/QeWoc2uji+g11Bx
q1CZddUY5MUY+GjGfP7Gvj4AnIN/TLKoBP0Y9oK0L/gvtDuidRdHi6ZyWRhK4dYInCwp7ne15cuc
LBh+kVoncW6CC7il++g06xUOhFCSv9iUMPN4gM3GRcj05WBJ9wwTTGpCqBbyDbAI5BYzm68rOlkm
33jl91qH1ww5ionAtQQp9vSKK0s9rLRZ8tRCu8rAw6M5EB9l4Q3RMxZbDmThGdGuFGouzOiBV3+f
Hyn+08O4kZKe3JKo32RFuwc99bGd7KJUOhVMw1zEPrFFvj8HQk54OkU2ggiPmfgwK93FqoR/SSOJ
Bvkt/dY6k3YsPbGexZ85oCAuNU1T54Ux5MvbGviJsVr5eg2Jro8sZXErd5ZeKCqwXVqDPHpzJC/R
kka+HlUrETDv+veO51+J7+BKZuAea7w7iz2XUfzDZSk+mTJDBmD4lC7SlLJfIRi/24paiKGCJDK3
3wSjQJpdUOabZIfBW9j0wXZeG6YSq6t/jZIGaV6PIqg45wL6jASdc3783q3e7hu4ec4bZ1bQA2lA
uDkoH6fULqhVHa9zA62NoN5HDvHFAJsxnxZXv9+hBsoLyR48aAUl4+YM7tlNoQXvCgCNhG2Nqjar
G7a5JFEuEU0tCfX4uJU1FxAlymNkeH5vKSBKpCY2i6t/ILmA1HBPZIoYggLfLkQkpGyeD1yEAjCI
LqYa4I80a+qTqV8TG4x/5ufRLhnkHgd2kNqUenCLDJEfGA7Lsiiy+q8K+ebOSLqdACNq0fNxvG/h
HLpJGUez30/WfmAokLQl9B0emZ52m17JcHOzTASM4YpC/3h7YWUHUrCax5M+tlOXyJJXvDj1he3f
yF2bSs2qoH4NngV/V5362u8x4HsJc/wBjyRTO6gi/o9rDkfJeQL/9QHH125k03ZHZGj33xqml31j
k8hpVQjAjtMUdmkErizTK6O9K+fmVSoee+MI8Ut1x+bxu2J6PjtFddCDfxPIGh59vVtyoWjArdlV
CAFazpn5ASdfB3RK/SbmYuqYDoZJaR+N/x5OIrpuDI9p2LWw/6QAuA8cvrwLjp1LqgrDfq/573ky
jAJbDxnm0YvcFbh/FBD2aRL+mIXj4vt3Zpdkjz5ufDHB0SDe0iq6vwrZCQgf3cj+7RRfRRz9D+sv
80Gn6TBzDWMMiz53KIAldfzdVh6gOdy8Eo7xWpaeRnJ0Mbu0hRvJxEc7PzEjI7ngycrmj08dE6Fz
a+t+AUzguu/4tPYyQ9QoDqEn1u99isIHrq561ECC8wYQbKivJbq5jT2Tw0vvhC9D76G86as448Jn
0byUhPvs2lz+N2DRstDMXrRIU67Ol/VCW3AGMSK5h5zVlw+xYYyBQ9/05CH+8Z8N7CipfXenbwyN
QKseOhZBVWt2gWMfZQ/d/OWJw08ZKCsT7MVU+bXU5fs0ZYEkKpDk2i/NcA0vrDpYfkfULTXLdD1c
uFN5J2wnuwv2vUMwkOj3F20m4sBSt2zwmQaScU7Clguclwn931vOl2nWWWX8GejSacrTXAH6jOrV
nBR97vJzoWhZraJMHCtPWU66xyb/RosZQjpDwOnJ2Se65dNSv+l6jYKYadXi5ISPGsozJ0gr94Ry
trQADNFIYKPCNOWlTHct9PnsIEH5p/o9lt2Fjh+4hEy/lDyT1X8k0oFD/K0TTj6yqTd6NaAdryhL
13Gx4JW/4cKKu48+ozjOnLR2ZPxW+oWtrDPwOWlvh+mhJlSvV9j+l7V8DHDgobPI4347OwHLT/Kf
E7uM6M7NyXfVWZo0QsrQVpEph0Z6MTQZSD0RR71uDPuvizsTj9ae3DyI1iZmkeM0kYie9dTsQEcZ
514nYNkvE92nxFiffwwS/vqm9nm9zXUuGGOZcppeOiwwVqsqitDl7UVhY/xUWIyOlVobmOc4qu/h
BfBgUAEm57Tqs+t/zEqKZdd3GHvyX0Zs4yjYbIm3J5hxWMaAczcyBLTYSOxm7JNMfNwxM+OjqSBy
YGfI6YF+dBxzLK4vl2j9/mS2zq54EkedjQDmLFpvHPpMwsU9IAokEZvXLMlzemUXzn6mAu5khpTb
0z3zS6UAylRLd2pEJeuesfB/+qq+ZVtYWM3ihzERQm4XWiOGPyNdoVcddy4NYSF/JC7PGanv61ax
ipL8XzH2WYtJJBeFDk4iCstwZChs6PTTjMA5JD+9kUJ5xrgGh/QQYwQAQ51ERvld703bdzJJNqtO
Y3K1Q+C+V2SSut/2avdO/QU2WVfxqoA6XXOyGjth0hLqijxFEU87rLgZQLtKteWO6eCaLa3E+arY
01JN+8W5/Qr0Q53zX4lehb9bx5IfRFA13AWoOZ8sxsYpMk/LdTTncsk3BNR/EfDk03FJXIGNay28
70cCeIZAa+GURewsClp1P/NIVTPBD+X8STsKpChpy9m5OH6UtIkdj35UHNg2klbEfuuE2iSAT5OB
QbT3o6QC/s3PaDBfX0wB9e7Cw8wrkyd3x6On4hpTFMln2es6B36z6ZVHVAvuCnNoa6U66wMeApdt
5WYioDiweCaxtuienOE6lkFI3w7A+9fnY7ZsLYZKeu2Oi7UtoNpqIBwfun2nNRUs0j7lzJbUbj12
Gj5X4z+jzHYAerBd16jF9BE9kZZQXXiI4YzVZGyQ2nugnLq7uyLwxrwgu5CpcX+2QGi25ZH50ZpQ
IvDjJvRczT5DpllCgg0YIimX/A2JhbfE8+nownt6YFv5CMbLL4osdSuJpXm+7UlXhhMzWK2VzVFv
rO83Z8NLodNXsujOiF83nEaFEFWPx82ArUykD8Jpn+78glI7BkR9wusBKmPuOGffAjNWIo0fj+Ar
WG4NB5rF6fi/oobPO8n0HI0w7mFSlwI+/+5e7D/x7XWRj7FVIOWn18MLgTz9HjsvCkQ+JH/UqF+Z
cZIoQa/ojT7NcbH/0dD9MvanN0gDQLXdEktyh1+dFnaXXyep+Bk/fMKnH1c1s7GcYj9bv+IoPpwL
0azaHQ7MyRR8m/+lIif4hH3nQwzdDf1gKaWTotsPFfeo9UofBz2IjJNVryFzb83QtNRkNQx3vLl/
2UBQyK5IkG4YMk802upynmiYkyxxstMPMIUbsrvi9RGkVf6XOgJmwfbCcaMq6tX2jY657ZaaCnPq
XGeWw16I+7Uo5jQB8n8u0sl9c3sT6OIadJzgonwGIbLL3vN21aY0VvACYNGdb84POoWM0SucAhjB
5xs0i2eQ4bJHrhyh+hEpp2rJY1t6dV3K89/Op2tQfpF/gFK6h2jyLLqbXECrqCENwQ2HROkqWsua
/eYOv4dkWnsHPKFZ4WnO9gy6eRrBoLH2Y2FwtF/tMlulGPQzMeZGGUqCbfCW4YL3uIzqsFMqzMQ3
Ndd84RQlwsVy91ln4aLh/xEM2TQykYdzq89GkwipCr/67cQZBHEYNxU3WBwp6kLi4LV17ywJQMts
hkILnRMYDxuQTDA5I0bGyxszyFJ48Iu6TbgjtECEPaYvjFGEpiSAifMQZD+vO0tB0s/SQV4fmimF
Q7N/XbaKbo4/3T2sxs146itXy6qsqAW1FlGUMym4dTwyUB9UUxXQp+uFZK9qFACOYkDtoOyDmT7S
n1yAbURQMq3u+9euUa2iZ6ImJOv7qYseKf9y1IZax1xLBsSSKiJJFzmuER30mCngXZUXy/8yn57v
FZgTelmHbevBYqMj3CNi90QAD4k3i0Vi7A+NP7AeuegGa6ft8mWB2P82u2O6PLC/jLTWw2PH/TnN
j9ES7HGTXVVkcBYBQdyovXhlteY5bmMVhpR0YdcIFPYmOFd9cmP21jTuubSDyye+v1OjWiONSIE7
I5xIG+vv0cTYwBT7tQx8B0u9Ml9Xb9uxsIjX0+6bpjP0UcjSzuuaNRr0x7dTbg2USHI8gBH2xB5T
DvzfY1t/R5X9PfESR5q4YvNTB3jFFoC0JC5AVflfmuLP4m7Sa879W546J4qi23f0rjdnf7LvSOA8
TMMHbOoni2mzZrjCGSzvGl6uU1qYIzDi2Hus28AYAS+2Y9JWZAieNQRMFvnIMAO82u8xXSjZ58GG
A5EVjaic5s88a9zdmtNUN5ZlOm9apkBOnQrI7tbDwimYdZ1V7BfR2o/HGAMbCXzZ4Dxfbe2NV6Xm
Eqhngr+ynqvzrpyWraC4rLrjmS3NkhRZWWwnaCAPnkWTQm3a1agrWKRCoQibEyM+y9qLqIpMyYOH
MRmfp5ZgWeWJFFaPmGaH7t/RDpZzhbAv4+mCM60aUBOikHYsXs4OsVlsO/UuIvudWROANBR3AKy1
37CAVjX8AcUkmXBxiuYFHjAMb/apVDCAPNBlQ2+Dgx5BLyQwtq4S3wvJaadgInnI2I2yxiRM1/FB
CZc+00w8lbAS1YYWGhvq6ssr3BxCIiR1Q6eCuFWdoTcUqYUzX2t4ESDZiW4lECbD7VbXb130DuRI
dM2DkPdEV0/8Jv2bLxjdo/FDVTCxeQcoeBq7KNm3naLw/SUv1H8MeZzgCNoJYeLTqFOjEkK1E+9N
uvEeXfVI/gDP15MoiR3SSAoTxtSTTY+xLToC0TX5pnQWl9IkutG8RIT+YVJMOIGZQs5I3Qa+eWym
jX6CUpuu5kNdMwM8Iv+juT5V0iFyXOd/nFzZkadnNyMdQDVTKRDZ6FWcIjOQKGYf9cEheyPg7TeB
wzDeiSSZX0ksRibgQrLvFAS6nxzRgKlbjJagdQH7I1cWQDfUEZcHKbBG7uqGGHCymsg3FNZv0Xlh
M6YfnhXmyL8cuM5o33+ylzjHFC3zZK/aWoFx/L57cnLS5xkv9iQiWWq1SaIZTkqNtlfPDreQXHYj
ZpS2TPDIvclImZiOC8A1Ibjv9fVMveaztpspztp2LGrLp3bGURkXcmSQuWjRs1oo06ptXxDd2jfe
7/s4pHwMoylv9A7kbmJjAM6UUffEHuBj5Ja97WCFVd0fQC4f4Okztzm+v8FHEsicNnBr6Q9Equyw
L/MLEDOjL29hGQdO5whO6g5QUTu2A4eIhdHXrQd0+7sNxqd77esBsA0RyYRP+PD2rUSGcBxMhiMl
HRDkDs7pipFf2JYcXkYcYTgydhU4Ai1Rd2cJ2h3E/Ds4Az7yxt+Ay7szIPipCZtfC4WUftUBQ6xf
Zj9eiQNBUgBcJmNg6UbbUwL/8WATMR6kgGX7P23RARNzliicDjp63807HTZPgA+DCm1ynsNcJNeG
a6A9DJ4TLjiBN2cUcze5bjfMb/9tQHX+1kjmWQlJHvxifyM9QBCj6VfSq8fkhNUpMciU551WL2Gv
mjZcSJklpVny4p3nXbcVwPWyH+GQvck3kfghJyfx4A0HownRKvnlaba3QYR4o2x4f/iLsL64brNq
KGyG/YU59hafI7fpQSt4oNqxJ83dMQHWY2/MxR7jN+B3GcnT261dq0AmvgXiRSaSfOsrf6hbLSs8
VCUDZqTSAWRAANBZZleEnJh6rBroC1QnsyhhnKNuAW+eLoe1gZlp6tN3qkhlBY3vVxQFvjXXyyS1
mILq/BtcDjX4crk0EMN0WeT+ih9Opq57UZoRR77awTUTWe+qceE4g9FzPGfpKSZ9WhhYkeAOOPCi
YQYuphn3z8DtsiaySB1QMzdMAIRYGs1JGT4F61dCdTX9KAqyaEBKiD8NfqX+VH/HA0yG+nIRCAeO
9l/T+PApUhAcWfAnVsyjTk9uE8SauJYvUgtgY5hJknW8Bg1Epp2VtrZxYH2z82Ma9zv/lPNu7vju
hAlXQY5M3AXL/rydOxpK1+AgwF7u0/NfTRoNGB9vA136NhDHtw+PrQi37H+zF3QBD+evAo/O0v0e
F+4pNK9lFH+1iq4z4x1q+iGv9D060jTfUT3IjtmvDa5igXquv+LKaDXBo3ffdbw1frW24O+NHMTD
Y6R1LtWQvipDuhxJHQQRIaSmLSFM8V90iOhawfeE/6OzBYFvedO8Yxf+LWy95CGnqRyjOgrMvful
2C2o8EDxqd9cvs1EbXVykyaUU+CJiTw2SfYlJmsjRKSBHw+RvOGFRDuyCcm37HBZo/RdRW1pNQX1
OrIvDY8R3PKSilvEWM6Vu0r7xuBmr+/ojCTFJXC62NwIXpUJpRbZxRwaLIjmq/xP7Uc8ffPICviO
CHbMcbAbJYYkBbKUxdfM4tDpEqFbMkIziVJoHrL1wLxqd+AHzkClFN7zeBpEW5spfF1Nh5+N28Be
Fvq+7CX/zjhrANh6hYvflD17mdeCfG54BErQJSLMiT50IxnxwHIl3CdZZPsLCaR4it/VyvpfOPlX
nsA0pnrsrgn6X1zrEILBAZepr1iRqlj16olf/Rtq2FbNgV6ljAUPxUL4VI+KY9Mx9gtV/0C2Lq1k
XcbmpOVYiY/X8GmypcCSSpt5QwvkQHqP7t+b5oPlQb+S6oznT/rKSSrl/yF+lUbFbg1aoHrhkKO5
jEAd6YK4C2R7uuT6Kg0bAtm5lUT0UmJqoGNcctjjwll7sTNkMASF7pqCoRf/0Rg6thW5eEV4GGLs
UxRznWxMYkuUetfS3CHnibCJYv1zEq6431x4A3UCR0dDduWoNkAyNKtvZ02dkYEJ8zHq8rzpgPe5
2pvvTNtDGmRJBt6PKCuEGXc6B4JqF/d0U2QAguvLCxDFxtoTJa76KQv3gVYK3KrmHlIFmAUs+SLS
prLmDbgZyisylvCjZoJsJ4OW+Ylgez8fTt464J43Hzh1888XtJaF/ocVH04GbdPpjVBM8h4hxQ9n
/yGsSrCVTaMlopMGkvRFNJ/C3r8UoZ/UC8CkxhSnkfM5x5voPvvXzX/xMUwhfR9HQKsm6sFZxV4e
+9KBfk6NE4birZ99/1cngYT0qMF3pdmGHMxilgy/2i2koU54Hug2MvNeJogxdDCW6n8+c3eLltCc
z464j3hlozxad6J6JFa+ez/xC/I5czi2ttGHeokEt0asUtCfpABj8iQRgtel+qB9AO2VwHl0UK1U
8KTMH6sl88wSdN2kvORe2aHx4FXYSW28Gjjfl1jvOVsmk+RbH4aMAYi/lQEm8pRHOxMclj8ZHkL9
mC5hxRppzMn1z3oidICU0LmGzbwo9EqaABSPgF0Iod8Cn8dIe2oyOZZB5P1faOG/SwpYBikgefhm
InpKnrq7kN+np8sAU4kdwMctsHYtHbZBe1AiPomdXihcQNnChAEIVDYYu3/6ZP1A2MX7lYr+WQzX
QzYzV3rSBDPvBmCHyFh2ohlZ/XHmhWPQfL4Dfmgyvvo/Kse/P3JK1YR1q+9eCYpiODVJ+24Mu09t
bQyxaSiFeUNbsovP+NV5KBtSRiYGxK87uLGblhZziJ5zN8GbjhTGqkGH+UA1nrHbuPk7QCGoMOIP
JoNhdVu+zQmY0UDoNkHU6908aCb+j3v6O+hKb5kJ3AnA97x1kHrCOKyt/OnWwhhmFT97hg5T4h3F
ZcHO1Wk+Yzavj5v9FdpnT3qCaszeCAaKhxxUgxfwiQFPl4s5AJ98lq80w6+fx4GP3PrFrsu6B7eE
oyFnXZPiVGIyycmBeF7D3719rp0x4Yfr3vl6gNf6fRTMUTOlp6tJIbEKIz+TU/hGgqXdPDJy5JIY
ykzXq58c2Xz8PSBC8+3jzYCRkqsLvIIfzQ6Lm5RuhAbUek423rI/fCkj2wyR7kKn5xw4i/7H5z8x
Q7oIjcM4SOHsj6arztGAojoXgbckWcxZCv47ggD69ROBQUoayqXldQU1FypOXr+RcaJDfKwf2XHf
bGtYz6ahWnd4eTmmNMRP0938F+QBRwt6+k34OSwm2MGGnyKIWBcjeAdkmuvB3qJBkIdntOlL1jjj
SX2MlJz2N/NmmDxmLgACEZ9HXi03rXyWfeTB3yxJ3HEokbQZO8r4vuxHILF3fjeqHMT0C2F/QHn2
ONdaqWxp/FBPEb1qwChNM3JCxnD2W2lhk+XUdfMjq5YwsCE8Ep5H5qguv/uBBDApbkor7MJ66MtN
R5rhxDjBxItF2A9/HM4xqsfwQKrHZpmpoQa8zsqElAJ2ThzAX/U6pMD6YuPKo2VNZHRVrqTxQeqn
w0i5LMjxi3LNk0FKToOLGnShdH1ZENXcwbgVrqltX/ffkP+VGZVvliW0THS+il9orrS1NSjPPTCp
9Lp7x9JUwlC5ne3ZKNgfTSdp8XsZ+uOo/5iCa6oqNcUM4KHO/d2qgAKUydR1GZE8z+n9oN+rzKib
kyElitAi3UJ7YqkKRXF66qhgM6fyE2BH7xaURQ98aF8XxOE4ueFU0OJuYiKM0c4VGIxts/SjzxsZ
bbprFzxv9FAaxm9NeiNe+lHQ99s5y0LM/3l7nULSJwmRNcNMQluXNsC+K1mCXYxVqbGlj8ktNP3w
537qvKcCL827caj872T+xw8EYgoTZgZujcsh3CUCLnLzAPs2462nP4jWtgFUw3VcezuBSd3kUR4p
Nqda3J7vJadwuDo5WbhhbvvbWqPd8fdVarPIjDmc/ZTdoflaVgrIpzuNyEjb77BQ5ppO9rxmYgnI
rs71qxGVnEwLelFdXP90J9rLB3RA+1HQvzKCoDaHT5vIgHtVaIL6BkC11/5bRfbncxyfxaqW3dYk
CC0ldclCZSViP4R5hTuqVF/GGb2KG2F/uDMfzN4iG8119GwWDyXBCZqMins/HK6/YO0IXxT9TVsp
jYzmAW9/ctJpT7amP1NAib9Ff+yVDBRqr8zCyFoaFUNqYOy8YFIifI4jrvSwlFd6OuZHdRYj7xg6
jMnnlm6pP0Bl8v193q6pc7cYgecxP8beFSNh8jNT4NUnS6yo6yKBtUC6MXzMLPOC5vGrEvPVGqmT
E2pVdPCJvr+hrrER3SxM7YcW2sgaWSPrYOEg0bFrIbDXxXADtVmXI1PVavHtsYEJqPpP8fUFzNo3
Q7lNQmiiY94aI7P0ifl43hr+WQILMknrggDTC5vRLR0CkP5XfnFLOaYsfF8OCC0R1ObTjGHleBPy
wxOQlmkIdfKtKp+fbTMy4/TwxNIGfjcEmGA0Ld+xrVjHo28KPNqaldPqtRHRhjEF8qTs/bO3yCF3
qb9Efxg6UzvC5KICvmLtoT3xk/7hb3S6WvjAmHmTBMgrRk+4zRgelvKxxKrk2qv/LRUDxMcD68uC
s0GnuHpbRm6IudIyqyMhgJVebXqOvpsXTSmfdmKuCI9AzoHZU8o4Wvt3Jp0yPz4cpB/0kD9SdR8z
qIB0AEgB8C2/aFTpXXELiQqsPHknEyMt5VwsQI2QT0nvpAYFPst/YwdsiBsqK+n5oQEEcdzNJMJ1
roPzPMpWZzfLtb3QvCHSjoP1BT6zZaF1bcyToq2vVNnXdAp6b2n4dy3zdAbLwy4JNLeU6si1IZar
7SK72D5AboUWPiuzS12x9EczgbD0YhT/6elr/IqeUt7tpxq1jVS99YkZ0Z6MLEIr9Xq+vFEL+4Sr
WfWm4lpbSRzz/znqbTYsVl9ByS9iojB1LovDuxp0IYkUbHzRBsQM9PUNxfwnDkC90e3W4G3Puv9r
gnySld8CsHLpD6QUN+aIuXRPseua8Q4KYzh6RT6fDbKubuJIEji+dn///3tzCF2voWLmnCgAAJwe
+NxpM518KdzP+F9t2U6ME7asP6eUJLHIctrav2YVepSUQqSTx/23gD3L1ZgGtCJru1jv6HZvBLDW
ceyV4zGBD1ykSQjYvRurDxWBAUB0ugKp5i+zynVAAcNbKjUY63dTMSnObqlZEc1BXaUBW93bIMNk
JAT6DXD0ifj82AlhC15XLoQncoHY1JnJYA6GKFxooa7KIN9fgsY27RCdF9vNAJA5+TtcbXg81ijC
fz9iKK009P1sEcXC9tuuSUllX8mqb6SxiQ9yVHeiyNrAVqxkBrWh+h5KqVBgr5QsslCEjVVIUWyG
J3kNIqlteHdXhsM8L+eCf5C+6BewRBFVjy2FUmjxH/CiklapsVVmpil0e+ATGfCJ4alZ5nXTt4Se
uyU6Qp1CJP8x7q82ZEWDOSj+cP8TSUlb0z4yoMNV5pvZu/tJ6rXzH6Ac1a7UwfB7bWYqkNd4B2Gh
Og18p1dxXeZn/KC/iyv66hx2zOhvGQvJxqjjwm8po/EyoLH8oH59Icfn1pxHVuSewjEQtKMFnLQk
QkR6lBnnAdt4JYoreTXduVa2BayaWFxEUhujP7bHdJVHGTTztfR5y43YB+aN/lNkUHNAw3rLXd5b
jCreZmCEmA7k1ccS4rSa64yYsQ9pnEVLCYtcA0Jp3jqFzhitdn/kDhLiNOfTA4sD47KsWrjEJVQw
KI9gb0MFXqWqDRT8HdiL0Q5j6iXREIU5DojapddOKiaiBm4/om8B+YXU2GHAeAXsgyOdF5rkIkzQ
paeNKSTZeLyvb2aRQ6Ut5wDGFiPFyuVA9AS46CETxqjAKYI9DNgpA/iQaY3qtWNc011bjJ2LKGuK
occ2moxo/xGPnsWePhcadzeW/MOUqfBcU2r6JJqUqZeIWraERf+tvKN73PlcgGeQZ8s8vE8zJd3N
mxPa9fwMTXlSBMfg4aOwgrt+HUtMNz457CdwzhucA39mLXfJyAbCVfP4NTlcULuPVz7dq4myjl1g
FeG+URRDQXuZI/qaPF/BtpOb2LYa9jKBWJurZZOiP0F6qDC3LwVh+nlsBeWKCpxPQO8brTbwpuBU
uzctAaRUkHgP+bbtFyCxKTjvD9q7jbS8Y6dRoOQHlX2324hNTsksWnI7wd0tFuCzdbDB8QzjlWAM
gg9rQ+foW2kcO6CExP+dYh4aPI8luY1lpSxFSzzuBYcDD+H33Axt1jlP5C+/7lDL3qyyzPkaBRMg
scgITjqlwnnvwcX490H8sWqiKA2ZlOnuyDZtrhmXc8nUtgvWpTxE6v8QrKYJlXVCzx1zoOfkzG14
emooFL9dxFxKCrJmMqZEhRNnb/EM7ikwUOcuiUnYgDn1ma9pm/BqjDKG1Zu01f649ntYhdvHe1o4
Qi28V3PtGHzQCrW9qqmRseCCO71Sgp0hVwcWELzM7teaBNQLZtushDzQbB0UUhLjW7FJOtzDxhpp
6dX2SrNCTz4gyFaklfCH8fbZSoeUdh0jFcSTnB9NQMBMX1UShirVlef8ubCSiNrdGPrq43LwDJlv
tO7tpiLuzEDFGlhlwndQzUsZHFats2+ncwx9sN1orr3tcjEc3bdhJBS2bTI/QWUSs2pBhw0GMQ8Z
5uC8QjuRo/5YWrSxp4+RMjcqlNPBxX+quYAjNDsBANkp0NzeRuVLDIhtFG3lzroa1NxoHWUepaxU
Ud/sGHhy+MKza4u5QZxu1wt/0/gCq/W2zKr0uvQ6TAt6R6sZheN5DftEHwv8OPgU0C9jGMGmwlBV
mLKtk9onr5JT1BiEMCGgl4adyod7r62clDXbHLRXzlZv8vnKOV9ctls8HyBp5YolMAT/cLW+aWwI
GE8A8sNADxabnvjHFafqB+eoyXRlz1rPEeawOJb1J2ixq7c6a3AW6dSHfvhOrogLBaxLddYffyc4
/5UU3cyW3cT2ylmk/WhGRYGcZ9a+KpBQQdSFHDiEHWi9mzaqaLkB1rLcSn3wjnADUEumVw4FwaPa
7Prsatgw63L2Skj52rWpQbeuAaFuavNto28ubK1QDtyyqkQtlMy/QxrbAC9R+ffFc88urjY1Ws4e
+b9+Ff3RkIGFy6YvvjmIMuNV+oSgTdCMxmlwsorq0t/3WxeYwREgJirK/DAu7Ot7h898czaDNYEI
J79qU7rl/10bik188w97DHiV6OdYNgTyBXjniRD4TtCdkXzwxY5AWqU6fAhYTUZAitIuq0jFWecA
dVwkvvWW1CyrNbVFi9w+IN4cWN7YDR95kDfco1q8jQUssLh1dET1ilFdDZ8jXRsrwuJcwTArc+CT
pPdWo9au8AFvucJX1FqgMx5pgAZwVAF1BD09uMFx9HxdYMuSP6V3FMfe4hy/FcTi5h5Kq6QHdZ8B
ch9WEhobj+UUqNMVpjHXYM5ytiy0C6S5h6+4VUs2lICwxCoeEK3lA9wYrku3sYevJBZPtWla9yS0
0g1VhdIR+stqA2xToib38NCKnz2li2tgHw8w+VEbrZUNKNNhHd34bCObaNIWcME7X8hdvpmj23Uu
QLUry/seo9nE6mxssUXS2/5/Nb/4N2EBdh2psZdVS2t5BQh+o0XnEMdhS/Uy4Fpahhu5Pqbo38Xz
eZAtKXqWoxdvx83D2qbM32bfNMa6P/K0bhk9+oHTSegBstw7vsvEWqTVhfb3mZDDBDCoxOr4uuor
5Pg0DrIx1cy00CyKxeF2xDF8kwIYpVEvSrrpdfRQisrgCoZQT2M2lThVto1mREKB6q6AsUYjgFAQ
P4jKQvnJjM+NYXqW1iINawgTqUvT6QhcUpHxBlkmVD/bYIzF/5SImqFaGdEYTol08awtKm6cb1ja
RaKmbvAwOptX0cT+aA5tcxbiZH7dCGFuLuu2DjMluRvSrECMICjpl2xonkh1yCXo/YvD5v/13OSc
SMrG3VS3u4vkv+Ky5RUtQ0YdBOKfYWYdyocx3NJV60WHaiqnPd2s54OStIbvNaeW40cmZdOFquDQ
Bc4xItDNnesvnMFEMHW2fMvxnXl428PJJx8c8wP4t1RKJpPmEufOBO/k4hX5oes70LbV7KvP9Ae6
uivApp6HMmeMq+bGjoRZZ1jgkuZ/bDYmnKEkfchhvleA1V0c9+6oC5Tqor7q9wL/OpPOWca7A9Iy
ZwHpTHAGtdPcKIq1K1mMy4mMWIIMCQS4VG2DiDKxndZJBdkUmHsOovFq2/XVQXG30GZKJ8j9/Ked
GJhk+lb/RXNQntZJC1rM/9Em3VP64Rr/HJB2rdrUQLX95e7yKA32IKpv6VE6wcQny1uyA3iGw9Ul
daKx65Ei3nEBxcRsSbVg+aKMBqBrASYwBJhRfbkvVPjIydj1REBW35pR5SGFnFzYb8Uw6zc+pkdS
o/LGhe31KiI7I0mpxyh0BarTgcw2VUu+xcVIRMt6Py4aGdW1WmcsiDK2q3SN3BcMd+pCrqJ1q54F
x7i8wEO7wZkvmp2IUXiDZWN9fARyS8DdOfbZpypwJMGfTiaBupV3J0f2ZMxjj3xybOKpQgTf59ZU
GioRX+eiCle+gJ1QnmKNaOrDiIaK6EnJv+7i3nTlpCp+Vq+3p6o3Nm4ciQKXX/Qb+4369PaFUmyT
v6eVEheTKBT1c1Yyb30sel5ZHZceJ+Xa+AQDv7ZyCvDT73TOL5MunYU3/0ByTXet9PF5akvATpGT
qS6bM72HmH7hzdFI9v1x8ofxehDD4H+pT/dFKjlfHwGcrrC1i1z9AvGrHrsYU/V1AO6O7yJYyEFH
VaWL8xEMNe1WqEGNUiusTIG7wBZ2u/RieT6iAjlZyqyBCPQbilPeR1BNOb+eb+KHn/cAv6HtRtrW
NHR9tOww5t7UtoFTDaVTYGQZM5m4WPGFTuvB5qbPmYR2WWWHIAf6gPSPokMiEYckBoc2e+/rkeO1
BQcuMWRwNmASJ7Wnd/lSXq470+PvJt9oSIhhr30Zlkle1cyImBreKRUGZ6vQnhhV94w1JPFIpeB2
xxAXuVERT1VM5pfp26AK1ShQWkH5PxQnNOOOu4DuY/5J88laia5sgK7zA3C+wmCCj6yOGLt6kwlV
/0eymFjcwh7X5ZDvC1iDGPkd+qTb2dv8roWWSKMyxjeMLyaykWgtRBO24fxjTriZJ/vOpJg9BgDS
VUCDGpoy05CHlNL4OShQNA86u6oxcuXhhcrUdfaQQ5YjMeaxHO24DkpfEz6t+p56buvl/25bd/rv
3o1lzgUuk8LodYePyZSJN8ClPQxlWC4NpjxmOzXKGdMqLL9BfmfgjbC1qGateN4ChjEZGRMd9qW7
UUJKwwoaaDD5zTWw+6pmZ/KxxA2doM56n/NhJL1Ag58eXlapNV9uK7Xbdwe8S909uv8OiIHkNGSO
NiX04wE9LZYM3ALDdwASNX4AgzqYjofnZNisqd/bKbX2mAnSDSoJxHe83EFaekKZOUXJKGsCHMKC
HBXQcOIZG3XTRzVdyOmoAaqlz8kBXyLzVHe+NH+c8EYY9hCYcBM9ESri64qJQK2TRz6IbJNsAXMT
ldsSnauL0IXC9J/I9fPF97jVUuVT+rBp7exa8zbT6MOwuw5xcZdMFmbGOh7uOzK3ZWuNy/sAl4mF
4a+zHsKg4sD+eSJ3zD+UXYjvjoFSneHGjJOUXqvsWq/zJthqBHJaL7RmoTS9LXh4h/o3OSxMHpYm
m5GmL1IeWcwZ7u+MI00FCQdA8ZTpz36n5MInGRD4YPeteypzu1gk0ShoftRxPT8wiZMxbyN7+JWY
rVuK14w7e3vd83T7aERincgMe87Y+7TP1MLVdLYiXBuc+U5GBwU2obYFTkLKnE9Ph/5Nk32PCrkB
ARnr0IZNuJvOuA4vEfjsmqIXNSRDzIP3L3c00/PlSVDv5YBpt/Z0T47H4n2A6jccO5sDD62RK+X4
6nCuhDP92dWivNvbW8CUYIwFYmx2+pBAfdTOw7RtY7uDK/CX6a0GZdvxRlo/m+imImmTyx7d87Od
Sr1sav137QVyLC3T/2tWV8HXfWVKKANrxayLh3AQDaOOWMWx9qy8qp1YpXC+KiSttWa9Ty4ycErc
UcYeoYoqwJB6ZDVaoXloz3e4Fo050dyxnHLddfXV9nvbQypWybfA4yiOH7EFW5/xkgsnmGJGEuZI
wyL+72l1LsitkPgmxSyWim4mnobsdcTbGSToZxVWKjMz69hbXYKXgMymEGvwIugoJKAJZ7YbugQW
LPQgmXbbeEdHTKtcghQ2Eq7b85EtfQ9bO8KKKmlNpWeK5FEeBZ4+JteSvZGpGoCmP6iXY6b5X44U
r+HqnYORIRXKN2kEiInhaLyqa6+yephmp9PTLLehFAvbW/obGKh3HcTnjRyxjlsNc0XQjSpLqxVX
gKcuYUEH/J3NWU/g9niHyC4LVOcA26PDeWz/cItAAaG9HiI7fMiAAaRwbVFOvAqV32dBNlViantY
93zhRCG546A3FLikIAAw+GMQQZTDHEfIHimIQPT5GWvtXqe83PWiUhjtTce1aeZvnN3KGK9plBOE
GONophtbLTXLFBhLuIXX1utbsihPrShzjBI1RmMFtRIeEdpwLPe8b9hb0Zx/N5dlw45vjmUSmw+2
Igokp2FP8v/LYVJORM3PtBkZzG/9xwFqq+/GuwHxrvKZwPrIbftNF8q6SOkad9E0I+xVRvvJjx9K
bGbOzEEo23yyqVteEmr9Wmx8vcw/lkneVreiTcQ8AbF3x/JIYEDX5WC/oZakVuWIBSfVTlmZDb/9
/QLjuk+YrpKg6qT4v4QMMT8N1a3kogr41BCOzjXU1i2tieB+Vsm/ZpDu+/eQbhyWnwuKIu39d/ZW
d5C4NjPLJmWeMXBwtOTecC9nFZ9KMyGmcoHrrt12JM6cF2Sp7flwORXHEg2bjx2dECYF1YS5WuwH
sQhNssUs4TY02eqwJqy8pXZ34Cn7W/+KZX3OMSsiz0eyZ/3YZQ9uozs97PJhgRkDgokGzm4McAXY
jutpzXebw+7caaRJrhlfeQSzCIccZEV1mGs3VnC3v4s+lgP9Ga932Q9wsyLqQv4L1cICkf3kxkBn
mwbgkaJkoiQK+Wrv1W8W+o8Fu7FKTddJP7yl5tqsyV+Iw0FxYBfMH+BLwlxzSZEs2E3ImB8xnKh5
JeE1cS+SNMcCH6YJYyGMJF65ErHtxcriobOoliW3Lh+jbdoEbpfEPww1sVEf2/tEFSOckMboZI8I
GNHUGsXZJawIHRTD72bdXlarZVBOf4AesjdbXGd0I+cfqx+120By4dJ8NMbs23Mk+hst9qTB1lzG
44393dviUY8WBDQ1Qfma9SasczaaIKZ526S7UZ0g/W4CwfrFvvz+LgrDG705mZmkwppUHdJin57I
q/rsF3DFGkx5esYxdvECYYfI4usD5cyywK24LNve+HGTDbKIPibBJI2XRXynTAspXrCTzOC7+m6x
67xDQrD73U9kLwuhGieuDCTCy6zFGVas6759gb8QiVP+3a1CfWu0xUzHWYJT0qGUFTopG4NV0hwu
ORo7pc24LBrWpaSkHr4W01W/AF6s59soygzF6A+8RTk8JeZF3gpQkyrqVFTZ4ee2ugL8cXooDz2m
ELMeBK6hvoObBQtF5r7RJXBDwg2pJ6E2MK1QiHh/G5szKMYHHrfizRRGdmkYZCj/6lItird84sVs
A8rJEVA6D7OVhcVUMOaCaj/eZc1ZQO1U4PRMaxg8bMHast5r4xOF2YtQjXM3z7VSfKNp5WQ+dFpY
vNA0YxeqZFmFjBVzCLgzShzxNWqeVUEqF+KDFx4w1kSVjyzRe2v1gpgjCs/cYh8VlkLQ5d7t8Qe0
LgDLPL5JuOxlD/Dzdl6ZUguty6oDf2r68bBHIJz3vKJszgu6BcNkz0fsOkgqS6J/Xy2KkwUrfFq8
V1Qlv5Qrw1vBINpIg+gmHKEF5g1/ZZHsCvPBoKhsqCxv7Xl6+Tw8PuK+Hu9kgHjuvCa9b2pDGKFA
zt9mfMoqM0V4sMBYXz7z70ySG8EmK++zNKuz8bjZeydUNjqKtMH79ce0z1JRcUn9GbbuOSoIYY8L
O1ALg+HJ5EHbbiDnjCgWcEUyDd+m1/cv9gjCFvoMOrP3L/Gw5PyaKQBF7nibZbPePwcq4nCgBaBT
Ys8HNNkUBvBtIihaCsHinimgprP29YC75e0+BXz7wGk8uTBOOG/fJ+jtepfxd0Gd3X0oNxkOpDjP
ITwd5yKTI4aExj/ocK+P0M1xd3ED6m6+xiEh4X3IzJ/kK5HW93NeFThaDj9KOVmtLSU20MT2QeYw
nneE3CdvO5oNPFcPVZmVZT9YZGbDqQObWwrkLBInva4s31cYC3komSe/3/Y2GYxJqEC9E8pCQJi7
cfwaxcGxwyGvUaVbckmdP+2V4XomJRgnOvfYNU9UJWN8929iW/7P/W9E6oQxoPpCIPjvN8enqLyX
R1mr18oJPvSCrtgsvl00T3OoNCOSKKio7lbPi4s52auApX4LK4n9ki22aZcXWwxOfVYNXOAk2fTd
xzwyazdiwfG7QkLhoL836wPEDljIF7XKGBXa3ZGZswAt8lsmMyWGulhvmAH0tdKvX0/rwcGtzd4o
KAG39LNSLz65VCR4JpopIhbO+Fx1Qv//yISxqHpYAuEhbZwdiKuU2A1iEqHuO5/Ye5+IxrsVjOMy
lVxbbT8o40VjmBYOQxNDVxE5ylcCCyMx1ciA6Uni2WV1x6y/dbrO555DUqR6C+tzKQ3GUTLrfAha
zmMIV+KUoNPLHesYAL+xb6GC3NIldWCVxoy0B+wEZRQPQnOINxE090QppqmG6a4QljV57HZ9zvwB
DzZ4aGaesUVorGzM/CRwhp1dIaWLv1eZINI/8GPY80a7MbuJAW3/aqafxJQcAKsbWQhBV/NK16MY
ESIk3fugMsPM5CX5nNTNFTHflC3gG22FAtn+A3aQnDEIBMvsTjM8h8+hpx0bvaMLw/g8TEaYezpj
NuptbW7A97lCx7iyg6iLT0TBL79r5y7T03F5LMGteGExv5H1HqP0XYwUh+eSESip1Ffpc5bmL1wS
QAnJzNOpXlf8MgDPkL9AP8jIGB7Md0vL3y/VL828MZzWReZyXoNw9lT7+YyPpxiD6hTZszZlH2ql
KteWCa+R3vv/ZLV1KRimYDQ27RLXNMeC9l2ROITGXj+XQUSl8LFYNJehib+Hh8DExIk+GkEcezYm
T+wRLZ3h+Z30TYmL1WVwSZK+rPamJ+FbTld4+Hf7AUuvAaY7Jr4Gs0EvxjFsGG+BdGev9a1FzHPE
hTG1N3mP9qr0JOwD9j3jDY+EemwUN5Aktei+mM9AAl8wgpAsfhXyWUFbu7URDdnOzWDvHhNojABO
zNYXHBijSksKk6t3c4tEDLOWaBSTOb8jfh6h5u2adF3Ty5nXfA/awM8PdEOfMz5WpHgjCeupLPXj
pKJ8P4/+FqvRncm8amRsMJMFzY+rgJeVHHfPWH9BXZOZiCVKPgcEtvy4oOX6THUfVN2l4B/t3mPB
BMAwexmuOcV8j/5HEKmmg5HazwtnmBSbIYCDWkjze/J9kulkIwcKgcFQZjVEDVb4zoi8gCgnr88X
BZckABuAHdOjVGYnCzvPQgwdK0Vksv54ctmj6POcrGOeDBtu+P8kSxYfiwhIGssypOMDU+Dye+Rq
fsiF8nR21zsYYHP59zQgynAiMyBHtDUPf97mE276FFPEuFyBkifCz/ooa0eUS8ybHr9Yp989MpYk
+gfdgRHA5TSeuKQUNFVDarStsh0iLJ2QUB1MUPeA7VtE2Js9a7Hutud/VXGorEEzAUf9EocUUPQG
dIS+bzk7pOJ5+Iv+UHAuojCj/ukDiklKA9VqEVzgXOdeUBsW0PKRtZM+06HAcm8S7AwsIih1P3IM
V+nboPflwU0Ultk/hO3V6Z2xfcAA5Xc6g4uvedyvujML4bY9qe93nJk5TxmlXV8t9ARL5eouzHvW
VO2/5sZqLO0WkW152MwDpulzJKXtc7skgCh+4ybVzvWB6N48DrMTdp8gXy7vhJZF77HPgxQz6iUj
duh+gzd4MipJ8GukBqVqSSEuM5M49sOqJjudiIODbtnX8QqVLqydLSQXMwVjRgZ6+NAEQPB8YM/W
MdGL5Hs9BisuSbr5SuzgVHW4tBgSj+R2e/1Cr2t7djC6fg46yJGk6Jjbfi3nfC1/9nD4LF3bA0ur
AluzRwKEknlpduogyXJc3mVu4e7yyYuqNdg3I1kej9/vcwYVy6ysZSn6PblTh6ylmte2/XJfO+B+
ifNEryoWPW8OjmzAUIStQ+Pkbt8+na2SgfqfhJRnidNZ2veu58Glrpnxh/VYz1n9srbwf0jB7sOK
Bv1WJxX8+n1gi6C45HewQCs3kM68Kte/yuuGecAElPWTujiO+Qy0LB4a1nq6kWb0HbivCfhX0juO
oSwwvsD/LZUsv8yY3gk92ZsXOB7WpdLo5mr/0/fu0WemiepwRt7Uyv+VShhiMFY3wbtH14TCQvU1
LBucge3jp1bX4/QYQxsWMQziXcsaZsTKc0wEMRA3V3WCHGioidPkt9Ey0YdiJ6WfpVU7eQkH3UE1
duPDUcnMZqn4ril7cnnMNOlqFFuMst9FDRKDo56kmgL31y9owfXKHqLRWXhFbA8PUIXuwH426gxD
hp7/fNl/zriHWLVBXtxjVL/HJPNAn02IVkt68kjPvb3iQPui0SB/y7l6455Zj9KM/y4zpod/5caO
D91EK5z1YNtxjBNafjpfX1i2dFKdgQU0x2RgNyNQu4O2NwJXTK389Z81yWEvABhuJnaxWmjf+E29
5rTIf0AXBm7WBBDrCqglGrZa8eEXJxnAUN94PTBf+8X5zz7ILuxJcjClSPuUbP9i6xTZpNu1Jpkv
I0EAnx4hQk1vZVI6DAgtodNFKjCDpH9G3F45MdK0pyAi1pZ5IsvoC/0x1SU9LzrmBmRLCmz2R5/Z
fqaFpBBpUX0YEhVofhYdYHuJjC8VK7NATk2ZM8FFaEBWvEFS+dR/H1hyjlZl5cfaaF+RYxVnJ4i3
97YP4UFfr7+//G7gWTx/wrioSw66JAX5KA/OsWtyMR2s3xRcdlgsaPOrUAaF/W4dwxYcAgwv8qkB
dV7BmG8fP9gZMdwSNLHS5fWPaPjW0pqhpOQf1duYL0nR5xzNIwoTMV2VAB53EhIYeuCtGqTv8AvU
rcBxHKMkJI5rRgjKhlE9h6MgDtvqbw3M7wZcLewecKaOmp2uWRe/gN7m2NCvpQCi39ib8UQru4be
DarsN8sodkCcdLrD2z6NO16fYbrvQNfPwukMXMOUIdmCYKQD/fJ1OIMLGZuex0jYGCzOxbjxWUe4
H3m6ox8nQLNqReTg7xe8IDi/zSM/eQDhrGYvE/1ersMYa/1h1Nx4TZRhDaMCrrwrbythfcpnIt/I
wiJiczANDHIQI5dsY1JA1weJpn9FvLkrusIRVarm3GosL+kPesB2zSgZbFDc5+XSVfP8xvF/1fST
hwE6f1Yn25yG3RXplu+pybksORvgCRVsgqE7KQ+xMSXJh3QD1XbJN0IDJBlFE7aCrFihleHX3QWK
WejmI9NI4SZ18UcrgXHFPFeIGgAZpoqOYZiwrrRRjPNS8fdie/LpgxTrBkTDHXbEVTFCDcFJBz1k
N5oNHWNQEkvrr4qjhJbyOgHACxJNvblvOsdQolpYKZusmTAX+zr4ciAeaSXK/2Pp8WsqjgvSVnff
sd0msEjLiDu5PVlKXCY4PUyj11/sQOLnwLyQtQCnC/oSfbSvnsglVHYyXLnPIpyxMjJeozmg01cU
TS6BskL36LyZVmYYdsFaRDgM8uSTBJMW3EPVmT5v1sjNFPcvo13YEXdfCWVspOm3baf919VTi3IQ
kq0qn5kaFV2V9nRmmHy+e9il/qhcf3B67Vs5kHBq+M2nFYXAmTVL9bczcOrGsIYiQ8lQO0JpKjq0
Mz5D+z/4xhoa0kFgL+13F2PE1x78sCC8Jbn58nZSCRcFYzQxNZkCjv/HV170E24U9gb3BDzdQSyq
KKmHwo5oVR4skk+swSkTbVhQG/ZzYZAYkObkF2xFrkWcJZ8qgGiLlAcFhrJDuI7s7Z/w2jRL3Y2V
tolTcu4uFYbFfTZWk+x53vrv+ETRtSVaTa65Tv2uDNX3OMyaNXOkAvhw+joCHUCAS2x4YRIFCt20
h0u+D+RjiLv+VsmRsVCHSbI3Bt1BjIHbZ/AoRA9EHnCk72mW01lsk6QS5aT3PsoazZIsgQpbOlq7
SuOlkpzmQyvJ3YF/YTNF0Brcho0TnhV/lOCdibYlSOiu98g5qDInUJN5rl7CqNdOL3qSMMke/GqO
lIDU+8luSH665ZkD8EBTlUsTv4pVS1d3lzeY6vaAsFnRFPFJaUhB8qxWcirM4iRXQ28PpuLZoSML
KSr6Ag1JZAV0wO6jO96jccU/drEm10OOjWZf352Cl5HmVtUPXNAxJGTAOC6LKbMgSlTNBx3WxOEj
UHc67xDD6qiDOiNJDThCD6pR6TAH8SDPQT81mccZMyxdSQ+/1FsKwsS/55/zXGhK1ZF65zQptIyD
WZzcX4DzFcuOln6EJ0q1/3lJtxHLk76IWpYuM3PxbGbnBqW0Fe1iDqCeSAbMAHMsdiVadvdwb3oc
pKDU2GpAtv2/1kZKV7lVIu4eigNQfzL7xKKdr26bM9CYU4VhKVG/ERVTJoU8DnbMKDAGNs0wxcw1
a2IyyZ0Zy5587qwzXCwUXNxbw2yz9izy6fPBf935qQPOHmuVlugvt2MCkYHZKSEwp50DytKIHlSP
lseEAjfkNd1G68dmYuqVZp1CPhe1VhzvjZRraQ8ai/A1euVmc/WcEuInDudDy1QBoOoLoWbdiZ4i
PRCCzykYpV0Jmu5KmhbdRwR8UKpQQKoxsHxjY3ak3TXsvqPNOxuU1okjskAjfUk6x6hXne5gBgIX
LbdWLFE6YxkVcKhbdKNZ29HsUN+0bj4gtpo7G/gZ77eVB3ll7nbyoBIKGBlCqubiTM+DVSRrKEbC
ahKceDTJ5Ll6CLjvSFsHB8cB9g/dtQR5blF9LUXpUPwLiemsMiL+FyWLUZLw1/SG56+4Faq8Zvc4
5kLLxW51MHkG8m3bRjqVzi3DrlCHGKBMFI0R4NLO8iJEyidqELf8mZM2SQ3YhdkiIRb2quIX3rTV
Y6XYnB1dp3EROWdjeanFJw+bhfyk02127oVJA8fDxTncvwIIsLMahuAzA6Qy2r3A0Mm55PrqIsuV
VNESmpsH4IdQUpe+mCb2cc3o9eDFKRBD4CDGvbDWerx5dZz68XI+n08W9geqO7hyHlyWc5XSEj1S
MTvwSsFSova/NtoDIf7cHSRD6gFIrCIHGdVLzB0s9EYzxsRJhuFjYjkdkmVJrrDCZ4Y9/cnzbMLF
UIcli9VLwKRTI1usYekMWbb/K9kivwlbW8w7hLlYPQ6Sa/H74BgvOpQDJdwXYaOTNF+J8hBbjBtW
LcW9a/aSxo+TSldGBjwL8YUqgnQZ93dtl2aD6F4qqrqpA51TPMEAku9gxCtj0TIU54wHCCDLEbBW
UeIj6ckOwkLt3bvW3vqbQr62euFwjzxZ46ewiMzjY8rgu+qPCvsUlZP5ImSaN00mCPO6LwbX6tqF
naQCbeRk5wZq3sOeYvOQIKgRJmuNLkQOIm96e8C42GzJu52cEigNzj1kcsaMP11Cv8iijlBvRkXq
wPDdM09i9tqlLsQvFzNTZMArIyZ1ZBCX/gBqhovEHPPXDvtIoLUpVUIS6CQyAGAOiUiJBZNWQrwp
VgFO1Jty/8xDL9wRBt2xv4MLqA3yYkFjHwoAQKF3HOpENr+ylMz7CS3NP9gbybaF6+SaQCxK6tAJ
LTanrmVn7eTp5YOELICLIdol3HPiFOXWTvOa8I+ACzigHwrQO7AAh8Vsj/KLdHbg7DQBguiJxsRH
wTA2ixkx2kVwkwOPaJ/cEDGN9XEfqw3WfIdpsXK2QnEWNclzMfnrZmY/JmkfQPhr8yju+WarKvgj
pId6OHkyRonylajyJyecmRbV+RnAn17YC5eWgZZZjkUQnO4hH8Bky2rOup27LApWqbWvROApiHGv
fxLo9BZIY88ZqxUtkqmeyCzzB7s2eQGWMML5q0ht3NNP1+k6Du1COTcuS0R6uY7vmFk5nNIBvq9l
dQbGOiWxFNH8jV70Ch97v19RtFF8ng0QCxt8fNztLCiFD6FGjRF6wyjw22IWneE/w3RU+uU4KRxp
4YHo6lRMr/wk+rLBz0dTFufh9VF5bynCP39ikRBuesI/l8YMvnDVQ/aNQmD6zPFbsMqLEhgP1xau
aMXP+bHMemnwJedesobjG7/nPP0dBz6mtwD/ZeQh3PycL9SMrF4i5KaD9FwFU496HPksF2tcQGnj
/lO3hPwg28rgSLTbI4i5R/dY3smZKBvL3cwcKhFb2mIB4M15lM5xL4Mq2Dg1x7MLKPu7SUDZ0kHW
p/dzwcK64cLaHEH4F+WxTfJzqBRAiA/U9ZZgDnV7Dt5w7PFCxIuU/fcEcwV1CSMf66nNJyfprw3R
sFWmRv23CDCP8wtfpQJPgLf4+WVK5deQpPseYDU2k54mRNosgzKiFzLxzFwnS3F87mgWOZ5HKK4j
w+0j4DonnTj+e7PPDv1jdig9z0ASt14RArh6HAlucwRiwo7Zu1M1sD1HV5Hq7Hrrz7hBhF2b6DN1
b1HLWid9003+wVrwkJL+epVNz4VpxytpdraiQW9pf4CFgiK8Q3sPSppfLLnqw+8o1PKqai+bqm9Q
HpuHpCHG8+oNvsGi312jNgCeQgZ4DGQlqSy968cMx5z+wyt0nWtOXIev3gztwaKGHj29rWZDwAaq
0wGT0ajOgCh+glIvvtm31CjWj4nHqE7umsUuM4xyKheVVf3ZSsySyJbTjG05lGD1/lmRo8bbDQRi
hGlVpDrqudF8cHGfLg4TQJ5fq05/2Pd87KqYrcomI05rJtAJsn++su6SsZWvHKOhGtoGcYccY+HG
ETN80CVxyrAjWqz8hydR4XO+wZS85FjdIm6BVY5QA/kxN3xP7LgrIwNjxnDxRcZ0580s2ilxzfsU
EN4iHbtylTxqhEAF+gGxoF5LcCtL8iXSjS7iEfQboLhUD19dbhxvrdRiWhgrTJ7vilpMDfa4L2t5
V0IGDAuOipwnRWjqfA/0MwRxUHOAqrs0Wr2eDt+92v17uvulH+8cW46l3IgMmFRydMNrBXxHtEFh
TgGzaa+HsbDngIu3hkORD8Xpq7R3awNb+jy74YpRJuqx/1bWlymVgxKOAVs0C0xJuxpjJ2NRy+es
AoeIpioqlTAsoW8YYp3HfudPU0d7nB+hYlRKogWxW1EvBcahNwa/Wz5izx1BrDHoP8O/NRVqDH+P
gjxS4qP8lFMg9tzzX1yLH5VaTUJdlQUXDEWpHPsr63NkeGSazFlHW32tbvDX7Z/8IabL5pCSFpwt
QZhszc+hTCSdLK1lUbLQxzacmYyWxEcq3j12r6pyBZTFzC4uK3rInUg4St5tXgATXVPm0TjO6jZO
+TP9KzwSx5fLWi2LAM8hEnBMw7VdC1Ij24dfwjQhVMK6llv1aasnLld7Asb6k9b+1RoVsBxxIj2/
AVAUXu5u3hfmItjwe+PdXN9T6EMupDAcOc3idVV3KVZmN2ARH8UQXiPPVda58xsPca6f57LXxsd8
gDRZ05U4PdCJBlpMKqmA5UdWWV5npSFH5YgocSkZEYGO82+OgD/wr0ZdNqT4C/co04M6dZ3RP6vy
4f0vQHAIaT/PM9LflzxrXQwsCXKibeoISGQ8wqolpaf29z5ONU/lferH42LbOCcgyor/j/667M93
j5fJ89PficoAbOXKjwtaMfHkLbMTDfWWlNfSB/+o746sMT5kE9YRIfZKowp+2vajaBwU6o6P1h27
zeqn5sINrmmBW1K+27zqlK1NGHRy2e/bSx7OUCx/IPj4aL14WANcHRxPdQIjeujUUXYodZeT+iNC
lQuftzEgPIUuRsOUTWxisg7yM4V41k0mzqGyPfJMByBNlLEGPkTXZAzIokFoIzQbvsc1jnJ4AzRh
aunZN5t5ANEc5EFRdPx3nc/ebN/OB9pjMQVZxmm2VqjAgmZW4XRKMcTYy5aQOvt1rCqxo2BTYNv3
WPftb0+/JKy849pyOfFje6F78ZSR/NJmDFnFSYc4N/4zVq55VHzFmUOje8UelHY2XYwRPE1GdUFG
zFMXprygMdp2+ShaSpdwSuIqmPORuE0BL41ZmJ1G2tjeABqHDA0qqZDxQtyb1IxT9Be6iTUWXBsT
mYJO6mkyz/XxIuQI8RVO1fxec+Ab3x/gbd9AdXUPBOi5Il8UXWc+qQLOSHtTb+8Ela1r6SEFuAEz
Ht7iE2aR4LcM//GlNN3PP0jf7j9jXDJ3mjowetXpefUsW/2ExbHx+xd0lQHNeXBVe2bmATxffwFt
ntl3jg27yZLWbQc5f24/okJS1wOhoYVoOkqhzCg2FhW93q8keLJhvMmVSys8PbhP+VC9i000RYQa
GK1P54eyore/BkIt2ShhTHAALgotTP5Iox8onal97w+4f2rvgJ8N3zwUbYFLFEIvmtaxct6S4pPH
hP0ITDoNqq4ImAqsorwNh9NqKPSLMkWA8y/bmBYnhVLurE6cgGbmjh9r7n/FzmMHA9QuUfPteSx6
EILLVzTmXtguQDyPdiIhzlS2rK8TXLJ+9X2MuuCwEe36njqX0hKsQSdVoCm/arX4U+I1SgFqtGkO
sjZ7WCoYahGqxQ4/eB9j0f6XT5RR1rt392u6eYUhy9kewCA4+AQqEGYIvj83fLrpLj+vSXakt37E
LLBstoeVjebku/Th309r+gGVQz7yQc331Y6Tcfuk0yGMGyTDoOjbTgBEqOjMEAYaXKU1Wul1Whck
xXQA2dksp+CBuPbniHgEqA2fDbvVapHIXQpXSFKmoDy0O3s+R922jNxPjAYPB+pb0UDnidpdVKyB
6lLwEpzrLdCjR7I3MKoNTnRJBP8oKUKrYDRYjbPE53WFWD7c3MlrtZQGEe1sa9x/Wuj1kg94Di88
rttbY8SwtT1w8NyEwWkfEoqpdZh73ZghqKqqqMB/IFvBZKro41Zu+MPrCb45RNd70mY/QsSxOp0w
dpQ5kfbjrWIrnhC75BbNPdMZT1NYdMt2aP0c2LeZaEih50nzaNxkTtaoc5LnpD/uQRhuFOnwsFxN
HIlJRw0kWa35ZL5iXBIhwyrsofjzscrX5BE9G3zSZ3dJuEledqGEtPr2LNgroFaEFilEBlVnjLCX
dXOF0UdV/w0Tx78sSo8lODTMg/l0HY/3qt3IXcO+zxKAjemmEpJPrKqbs7XimIsJrspyOYIA2wTK
UsRLap2MdN71pdlaiKm7GUtf5BqZF1Qb1NJW2EqHUItLGMCpDY9IrBbP+vEk2c72Egz6Hcsvx2eW
BuWHO96Kqi1NxfU2YnfxwHsslw4UtkW8pbaHD+Ex1lMtSoXva9HYQH/mXu7j20DElTyBO96Kmi/Z
sLW8XWYz55E5sG9jv4V34VB5N7KB/o7WVFfzUlAkBFozkTjRLJN8o87AjhGk5IH9RHEwsX9vgnAl
tIB6LercDN2dMOGwrNy8deVToHJnT303Tcqco7cT0z+frRri6YKVpsTD3fNoX9A/K6W/udzY0miY
5ypevbm3uN5K8bs6OEBBkL7pedvPBh4NihmjMnyNHHz+iIXEgVkcLyaHlkt+eUtDAz9NJnjHTMCx
+Rsl4PqI8v9AC/sRFJjDZ4BKeCQxDxZcjHfJDVTiBLURv7NVSfenLaAN+w+gdDSeAOLRR4qR40s4
gzef703ZmTUHnipKlGZ8A+7CRP37r7lzn0V94Kc/RQnOa5kQKXzjRdGBT4e1AcDbkfcdnO5097Jd
V9HXga6a6R8Wf1vQfo6Ig9Ge8GaIrM5/DzMhthEd+3XWIdxmQ7IumB25W5nf9CvNz4xOcX8RjVtK
dQYoWiW4i+tHBOQBiUuMO5S7QLxLZRDbV66NYeH/Th2LczO3N+ExioCh8WPPShGdcJbAt2E07uhC
yER5e6pNB1Vvd0CRd8IyzdOQ8LcWFqj3F1DK1n9rig5mRvcVY8UylAim9KaOt1tny9J9jIDWhahu
sg8Ce2ZIaVQKZXxMyyeFmkhzSq70Bpe0/n5PujnZ4XEjvzuNZodDAvbSka03SnF60zGvZi3AMDut
5OjHty1G2ygn8jVW4S/440TcgPzOIsfOZqehOeRteljHFqLMs1I//GeRy9Q/euMsvFgghSHr0xwV
EFPzOiOYXDqe3Me3sIQAQi5bSzmjl9kLbI/4RkN7qwlDe+/J3arrtldYwQ5nrypaJ2qth1o+eqak
LFZTloYd/23tDoYHtjVxVxny2EmWnqZqO1qGw36jH7sd4vByvOAo9cocNjrMi/UX7HxLQuI2DNQ2
W2ujKF6Z6GKHiONmCkKd+Ytd7DNHKiDYm5WB8zugfsRTGKJOhNpJtSQh7QWQwn1s21yOI+QBzKHz
UQpdGVfFye62SSMcwbBSfx5KTwUPlF42kAJgi+DcCcVSn0tMaBtMy/YZ+cYQ/7NqwDGWAdk0HIb0
cbfTMNgU8vcaVzO+eGHpkOaXw3ulhmtg+agzleyu7LngHnoxRnEqhIxz6VYpvzaIMZX0A7buT+Gd
5zWb7YOlVyLXHijrAt39CEngNHHPe3STbIEO/ZUjnnVZiHXYRmCmoRi4ucxym3Viw3c3W5imhiKb
xy6slapNxlF+ckKpI6Pm2yVkj+rjAcSj6+gooif3IIUeebkihTpLqRR6udoTbbdFvrXTfw4wKGD4
Bv4JY4kN4O8eLtnRuV7ocs6yrpfbPt0NSbGdJgFE31YfX6P9MEyX2njFHPtDfLw73rR4fmYZDjlf
dgj8HKMX3/nPDIe3zTyLgXvNctxeSRgjPDHK4zSTV988ZCdAf1p0xFP0hngdT8a7325TCQCCp/pS
QHxYXkGZa3gzLhA8AbwacCAMo7QuCvZeJyFD0UXgD/MMrwuzjKwOpXLONxJ/HoDFWE8RMdgDp5+W
+zPEm3lJVjzxh+VYdSB6vz8Ev/4dhD7JhkWrdpEtg27G671E4kPvncZvQes9916OB4LpnFASzIN6
0U8qGZSPOG4Qz94PUQkAdTDrhDxJeJjMyIk7QrK+HfqZingBXR1enUr9cweva90BD+66b3WAoIon
a4aepHe8KZs0+r6uYI5ZQTi4o0Y1cxbXXCk+JqTonc7D/tZF3DQ7YGp9Y10YUA/V+RA4D7uWzCC+
WRdEPsmZxZnJNvXOxQL7XjDrAI4zfKoWEKQWGtkzbFnqIbUofc6LGq7qQ2tFkT93Y8o4lLltsuwJ
HzpN3aIIrkxUUbuQ26xG60DMYZsDQlcAq07pf8kP0tJFJfecRzmCYU/NPv3lU3lOeyIE/ZluOjZX
ZokEtPQf1IZ41hjOSYBfik9iSVp7Kh3u8beB0cJnJA1tqetiG87uqVZP+c6SVj1QG2y2LhR72bX3
j295WhYNXmoZ1jAF4sZS9evBh2OQ3sjRoZdqJl55N01Q1PJ0y0V/iTUNu/gl2Ig13bRnrzQlaLV5
X5JsMgm3aolxGa3TwJtuiVaOthX1uqpY9QTlINB6KbvREdL7H71Nc0qA5H09xQs2z2bExG/wh7sM
p7DDD6q6Te89h+t/pFI9LjZE4UfXjFhOgMncGduYWus4mkdwb9o2ueq5SNg1wLOn4ROO1p141fpJ
X2giROvq6sHhST8HsHjftHnAN0TEUNG2znuTBmMlNRHRSrkcbLHw3a7vS9TzuWGM4nbuICFdG3zB
36uXJQJZiAMTfe1PwFq2NReUomAhRfC3inG9S69O+SjHcxkcXwHO5fcyGCiWPz9P3LIhtX2lA143
5xJXdkDsz6AI/K4Y9v9G7pI0gvKxN12Fef/sSIkaT9YZw5bsV7lLLUV+aUDgjS2lzNSGBPE/MwPm
RLJ4HJquzigAip3ZOTH3vg34BVrxx3BTnHjChfEhgTeE+Fd/HhSIUC+g3a4osWBUSCvPr0O74Ee/
Cv5/YwFU3NBhSKNmkgQQW7wXN5I/HmyRxN8c6JGu8MkG7nFUSj/qVr7nuPjB8ol6q3ZjKN88pr9y
eHdxsknvnYuGJhNJPF2yGtSVIsk1ZivV73y0hbFl9jAuNtj7wXHWPQdMafOJ5NNNXXk6ZbmQFQ2P
FuqHoD9C4h2zE8fbxefyrQbSOi2vdo8SmvUmYZRdGrSl6ngHyn7iBSpK08oubXH2UQicyvhneJui
OfiX6yVLybc9o0ASa6yytHWpS21mhQgiD09rIPsNNeYPEAUChIfB7xAAMGtygGX+iVwWPIoPfgfO
lQk6J1fH0irP13uoLC1p8v3azQGOyM5hyCT3H1NIpbDladXaZ+wGm+FHtxOxHul5zVKL0myQ3YRk
O99JfgOjg/qCwme6NnMh3H2POI29dY3dcg6DEuFmD/YUjUQXCd8sxU3pHBWlOpVVvf989ilDdzCh
aHc/hcMdybXQbAN4q5hSBZaBLR1/4I/n7wIS+ikUh0Y77RXYWhn9cVxm+h51N6KULiSKCFbERKJi
cfKRBf3fKzdiptRSyQT8G2YJx3fDwzim8NObt85fJsLIgQJjl66x9Y8wjlqt8uqRuQhkopeZJqF+
8TGZUc1AjAX9Ucjo15RzlDPaWv1jVqizR+aAYG13Jts4GSWW2k6xn7iWju+0gLI6i1oN0WaxC3/d
L6p9mg5T3BH3kTSaTI7WfjrLbvUCgmFDx6WXCu99pF0bi/zbfWFHTUWZm8iSj2ODrVHL4irU+lt9
XnL5bR1qqpXZrNMPIn3qFnmCwF1a+egKquvw8+NZYmRXKi8OgUwMd61KB4beuBFC2QMSyR1+jeyg
ikTpG1mlSwVxzUJMwPqcdCVC4Mdcdisop+oy6oX7YeFCFs/Q4IjuXnXpzx8s0y9IErzFWfeQstzC
qoGilq9R680h/IiB0fD7+NYSZI0KFwGlmhYIAEc5LqcNf7W6iRO8WycJhldvkfy+lZfgyaEZiuUV
vhv6s8jTuZoSLxFbirwT8NRBnmKem2GXd/JU0ICKelfVohKearqLKiL+Jp5wu7wyTlZLleQFYdQD
wf+bATVgGDJ4AcSpHvGRk/Qv/DT4+0BgRE5M+672QSUjX22ZibWZxJCodgExzn2VxeoUQuBAmSUz
7gM8izGlkyf+whPMhuWAzwfyiqwGK/BprlgVS/JQcfUV8AVF+MYCnyTMHT1xC3HNCfnmx7jho06L
hBgmI5qy/9sfnCbpqsdQ+QnOaAiaHcUj80FZkp7EBS5NnwXuCp5lYlwk8QQBHnv6zfZsbRxpdnya
CMsAyl297w6NfldfAca/4rtU4NwpOmypB0dHU+qMZP6c5Tkk4ojVbXiVB8C4rSIKw89gE1FaXhCr
jsOWZ+wmSye9Cf9mVyHU+XYC54a9uUdbEdnoUx9/4GsIGJnx+hporjlJjhtHcmJTixbsQ0qjM2lS
kJue+hn+qWi/MQP3fv+7ExaWMHHFnmE/izrmR1BsKd691CwnHhq3rMPvfhxIOPMxpGcL43tpszja
xz14sgLexNjU/pDBcu7J+tse4C7+P4ymv9Avn8zqz5ZdqvhkT8f4M2kcAsyVr7a01W5hJUoRAOfs
JorHf/hPwE/zfg22o9TFVinQgVSfvDhCo0SAe/QSHWhHZdtRNSwvgTt3Z6IWglzE2gTf2rxSgA/+
ExO0yNPOk8ILoYcGr/TsyjFm2EXaqfkVhXh2pNd9GgVv17YY4h83oU3dsyEoyJe7vrIrgWih6L+J
I4VZlQZhABegicmWF4CQZf39MqBakhUvrAf3sIb1aMzdcPa2PHsv70ThN6/fnZjijQBw5+RR/kqO
xpDaxn6eht8oUB5rqIZ+GM+iAiCxpKZD8c5tSlTqNFMs3SUCbSaLYoVRqPsfoNmDKnA/iEJWbu14
sYJQjRqNMQH56MDgFnuxScgJ+fNAmUVn44KwIBOJ7W8YTOULZG9SQZ0/cvU+aVXMikbBpwo/3BsD
nhX8TPpAtsN81NX+pLVf4pYO271ZCEnajdzg5peKRt6ScJuwbzx3cKgeHtA3BMNXBR6srZb5/6nd
3yAtscRtxfdiCJ/SEW6TBPxo6XzP/4WDsZz/DQNli80ldk8/icyJzl+buWiEbN22LlnCc6maxP/m
b89kIww9G/MbfvLU1FrC5W4/f2JKNW/vgsbbvTlpFSpMT2PgyGRvUlNogpVutBozUB6DYIYh7Rpf
1GRqEWGo27EmGKbTYvuClrmY2BFP+ao59vfFHCXEiaMcE9sa9lQwIZzQ7De7tta9Ck3fTtJpREBc
G408OjE7zJzDPHDLjfLF5edWBsPqebbU6yhOYMIpysNXRe3/tb6Gk3TK2s2aHzdfCTcyVE0R6pGL
uufubK2aXOQvJymPaWNl8LfCE4M3PZ5OL1M/4eAllWYovgVra2uHgXqDJ6Qvz4CXDkKdWfjt2ibC
gxZmih2gAXrOIBRpqyIq2geoWrZLeCcdtO29TFvA0zYAGaiDmHSExZMxfT3X8NtYqj7/KPqh2vX+
PcYa866DQZimgSGmc8tVHy+LvoaY3ndY+VdJvV5MpHCxscnegAubWhw0TzNSHS/RZV20MCeJYiKt
cWSD2oWjIgMcuMmE5sIMKOqxVdGnzIAX+baYfOKFfIZslXF5zeRIavY4Nwwh4Ou3IgMM3DJYcmsY
mdGOLxMF8IKQCVWnpwGAjRlgKdQHeL1/y23xpfUAnSH5VH1jzhWrsmufCPkxNGsmnFfK5o538nCX
D4dEehikdmSI619CQ46PRYQuhuko19xLFampMo+9gOSW80kkCkUdiSSHiMM1spodTtGytp/OaPyy
KB1mi27p5fHaLZ56GvH2P08ik8Fdaf1Trn7iUR6P0l/osQdyvIh/xEFPrjerb8epOk3ZDvzp9Blj
9x40vBRcFWlwn5Jj6HCBp+mfQF/5Ol+3GxjlXPgr93OpRHmsgG7pdInkZN0iAckK6jLQSW4PF5qL
l/x001SOl3tdCCfEzxeL+fH/x/VoxLe5+QEQIK5nlMA2V15C+5yTLToQ5pheIpF1niG1iVFW7Ry+
ZxW43WWTQTaP7dkRvd1kjL1q9iBSw3CTZ2zvT2vi8HeLDKn0+YVNBqno5D7L6dO6rak5Hbve1vpw
6Pu7r9Oc5GCFWk7asPpRI7NvvYDSMEWgu7cBidRhcBu85dUs683Oo+rKOODM22ShpngdoHNKzm2t
4WmYr0mVH9gaViZnqjRDKfo1PCxnM6fyTS6qr6D5sD7rHQ1wtz6+nWlXCppcO0Rj73s7riDOb++a
SzcoI99BGRbNzSY6b4vuZQVnmlK+teOlzl/bAqsaQR5Zoockz57Yg4HMp6K7PH9WB6baWMeBuK3a
65h2RwxPQqu8NAR0oW0cEEfkPGVG6M3OFI9/q9jpgcBS1Sx5YCH8mEcBjeKCngHuXVqjGv/5T5IN
BGuCLzvkIo882unHPtj05x2+/vBmutdo2V1fjIcWvRH2X8VeVRvbUegjDH8x6I1M0e7X+FsZsH7h
aZy7h0EKgZ0sR+++HRd8sU6p5YN3XSlG8B9FDgIHwRToNo8wZRw3geHDX+ZNS9pwd+0Be61T/UBS
mV/U6YlI9UEPOnCgsiyfjx2IC7wOGmukvfAvIl996Pe0oUM94Yb2hpYING+JmhSxKNMO5wzowcbp
yB6wltSDoB23lnr2JOUXhTUCkQcYAo0bev1LXuSd2nIlJ7baClGp1rUPKPwzWXdAnpnYoN3lQerk
MW97XnzrIinfOx5a202RPBZzSopFa40SMtQfBOR/Gpqacn5jYUr4KLKYrw94p3WwhwDCOjyOiS3t
CSMomN2mYXpj1wC+bq1VWPHVc+C5qDUI4CCzEed4zAm+0DnoP3sQ0bP0vchxRn3V8LrUTfPNt/yM
0m6pu2wcMHGA5KjHFBAWSB9jFMdyM2cUvgZBjlpMujtbKv566UoKC+aIkINhNPuQX8SABwlklk6g
uJtBgy3348pnD0SjsZoFmDV9soIAGiYe9TnfK4+Dd5TTInxm+IhDXmRNbx5tVmJenvNu03R3zpHt
HQDL3FfT+MOG6wuaRP2ChUTUb0SzkFRVxrP+7F+ouxJK2tt76Yvm/iHBDU5rz1fQPkqhA1hFt5r8
txNLu6gqZn6DWfhYPAUld02T/D5F+z3W0fuAHLX0iYqWUrqK95AeSdf8ASB2WBapu1RpL2VIFhnG
wuHopNi/4ihmHasOnGse74b451wIE53Q43buS/tDXgNv62tjYzoHecj3inJRhav/MqFU9i02xxmC
5ZHHgVcLqXOh8aIdpqktlIUBHkppm+oTfexfPFo5tP+0hwb2nCilxxBDf1NQ7pWjiI4fqnSxiPtD
5MwJb94l2r3cDhyaJ78fGIcRAiEP92w2k4VnkJ8dkvMSnqg04567MRUcaGQw954ESl8AjRqvAvog
zMpBqO3QJjKADYtaIhw1kZkYReJ1+F6dXlQm++qWS+cKx8SjFaBioNz403XbQZ0WxOizba/882Ud
77NZ4CAOy/83uy8HQrMl7yt2HdCWFS2gsgq4xhROcI8pezEtn+fips2B0rUBE8sVORQcuQpANBYL
yqWiQVZR5pFxIgfASVGas8ffvUsLQuRbHIZt+bwmjKUhYXbYuGlwRWN5wXmvFzHmKjolgZ2RmoUb
0l4HGLRkqLsxQHNg6mxzLMySD0CaKDM4anevnzQErMVmSk5uv3voUnUUKA5AYxlFh/o0195aAUcR
tImucb0rbm7oXaLohR5MrRvgblvyttY09rvKnB2xk8zJYYsAKSj4cXufa1cOw4QNXD8fkF0ViUTx
Xrrfh1W4YgMcy20PScFUJyAGZ6ytwp9r7Wa8oQyt8WW0YoN+N/bVHxgOHYkQBkcsVpA0b1/7flPf
fd/ufCl749SHpSyZRmn5D8SwwvtYjsFlgbBiLVPfq50PEno9Y5lq76yEVu5Eap0QR4xRWKrzX0/L
as72aqO0NpsksEuJi9j0pbkRFNT+loiGpHif4HC2SAZY/EEEE5aOJUzxnODimIaaKllkL3Li38j6
WUcr0CEGPPRWAH+dZlHrC63vke3PHqgZ8wZbTXbct/TgWqMsmdo9r6DlkfHDudVFXmtfid2NAxfW
tF/Hpw4I1N+eiczaZr9KIEcofCmLZYCewnNjhbbfHS47TQkDPL6TAbMGm2QtJL6wNxg/2kfvG0p5
8Fds2xOBuEE7bpn11vKw8sAVmS5LCnHngUYbByH53qqOYNbxi23XpAR76cLp+UjgrxEpAu09b62C
BbyzhtJrjovqORdPBnodRQx/SOBT8fOsTUU9KzMJ6qdlNBSISbAL5NszRIReYKJZyXxQbgU3Z+Mg
oixkIzNdBIkF3b+bfimnr/q2WIfmytnjrb3HSgOKzX5Pf7InTBcOKITHerRlVfrNPC++OG3V7u+v
ArYPGUXs/wwTPl8PaGzX1Oo+pX4lPShImq/bsk7KWuQfirNvPONcrXw479U/xiHjTe+411uXq+iF
NVJO04xLI3c755p/3yYHz4Uc7gCJj9Z9MK9zS1qK6eHQ5bxnTueuQObO99+yF9GQcwP7MDt8bnda
IKX9GSB75m/lpyC/8lNjtHrXSQqutCcmMA+8xsfiHmpG9O53G9Ertksfez/RIF+k7LZZzhh8Ynvk
6Mvd3h5TtjwUMayEg3+QhyOC9oT6FE2YmQXeKrNmDywA2Sc/v16yoKiOZT2gbIKsLH9E/pFzuiVz
ZNVQhKe+8CQs/63XWhm70dZeH79l4IPxhzgO1Ylo7L4nqZU+Rpbj9sy8tO05CiFd8DfyvckDdIZw
0rqB5hyf49d1ZAcK0ZCWD5WSM0hgC6NtuFJIQ04olbWoJnE0B/Ko4ECHXsh0Ui434uXZZWWNPSkn
CE4dfqCKmdqTaT67bICsT5pwCFlWS3geL7JR211n99sGI7TOj1FOpGi3dI8rp1sWRcR2pxwZHTCJ
ygPk3BaJ/6ghbLU8qh8dte9bCVE9vt2fqhHeI/uSxs7xU0TIU6/mTH+95nayFOfjhYPD/6i1jJvT
Gb+JegNcAjOXvyh40OA7AedMYGOMLVjcGKR1EkYf76sclJZ2Hcn8n52f3femVQuUXhASl1bHrhas
l2vRixroSANZaNJssWhn1AE9Y7Dr37xoFk9QsUsGbiT17gsABccykWp8tT3H+kCBOJkdWwJNU0DC
FRt8RJK6tPtlAhou/fbjCgknfzg3RURLHESP5zqQTGurVnrDfc+gqS6RnVQJ+uCmWj10rlv+FmSQ
148lZCL5qfuaxICW2K0CkbGxpOIlVuxsMZwCdUM6NwoPuf4zutAzRJ18re/Bxtak6PdJUyxST1aI
crv8E8mAY4tfDSPNnvwz5vavEQsh7rBPq74Zui4jtxoz6r3RNe+7wVzrFtiTtgyjiMvIL9BRbPY4
ShQikB72FnHsxEnsbcZDTlsKguxzqHI58DXB//8A0rfPl5QZ15rwjZNYBAqXZMd1Xz993MhYQXqu
IXvfyg+UKn3wXXnOhm1jUQD72ZGee9fkUjqXhSkc7X6wirr5ws2C3V2IRRYg0Nd+JO2OuhobQ+Q0
nS4+6j5U6RXzPDvUslXJGa4lwjkhV/+d88c0Pwa4yDiGG7V4jLYGjDcmEM+PXc6XP5YV0TRI4JmU
lmX4gJIpsTfjS3I+Ld9WnmR3FrUKnxVsRsrRNn+TzvTSytsco+8QegSJOjpgHLmyHSLjHVZiyop2
WIdhjfIQd8rX6B5th9GkBvV+Vs3c9+zW3kCXCMYmWVQI9FY3VzmFsERG+bUdni4VIIOyh6ZGGSWF
CwVxBu5r8wWc69v+VscLnBYLKMpJEPNImLjg/ZnCUZ8AKkl97kOEHvzanXOPMG+WFri0EHgqEgsN
6poNxL34BuGKDFkdYv3m+B3ueQnMNMt3SOMl3GOx93F+KfRykHCDnHCf2ElghpQvs5AJiud6ScyI
MjyP8+hd85ucHZSySpAVv7V66EVE+oMjrXr4JA7mj/W1nr/oDwDS1Cnw4E5lpd15n97WupYsNFuH
UbZwdk1H1TzvAInZE5tXTzgyEG4yEttJsWyXqwSiolQwIct6laEM+1oGiLQ9OwwUMYF5VAFkeHPr
czP2tcDgjNlCdIy7dVzyRPkJzXlEPzxZS3tN/cupqJHmSJ5pKCrv1qttWgi6+ZPRwf+W68aELl52
k9euoyPRGe29CmEWaSYjiJH5mHtFy+qwgNecMhmwXAQNnOfxNdXpx6L8TNy/6dKBc0f+xDs+Y0qX
sJ3L4gNIQ4A5068kHwQSfm4WbVIViWhtk9WKKTxwuc/IoXMLnP7Vu5wcaoKV52YWrSp5P8tETDLB
Sz7+81xERnsusU6djX3uwhrlSnUok6qamJEt91TTXywT0jPnVTtpPvSuQ1il6RMgO106PnsrEXSG
umCl/lct1QK4PQzSz5qESA5Bq8UcZtrl97sq1zovF0UsiYw4/mNLEQJxwJKi9h9Wp2k2X8vIcYrO
d5+9pMlCOo8iq/c56853/py5m2sIt9ZpPnKD8ikNdZxIfnpf8VTMT9yvG/XGhH5DdIvvhhNr5LVu
pks3HDlhJgQhIjpxkHz4dWDaW+KKzA1viAfwcZtsJb66UEUeJkEojWxMWfyFnx4q5Rrg+wz1veam
oShHf5AuwFhvbpPlDTmlAwZsC9n5gJ1K1/ZtCT1s1tYk/AwN3Sjp1C+v+u8tkMA5VdHOyEW2x0aH
9dhuaIylHQh9nwFoY670udLLjayyawI4jXGdxFaR7oxC4+Xc9dnPTOD65ag41e1N4ExlOc25SS2I
DVn0dCVhulLiyLAT/MUbOO3KJDgON7ObWuPyiQhlNSP9th18EUe0J4GIIlMItmuBSnM/Ixz8lkXH
kHOmcOMAUi5Rb2CFLRAb0p34DVLQGD7t8OeylpJmQXM8box+WoDviJCfluoDGyMAqvpjv5xJdg4n
QYiagUADWP2CMjyBqbvkW9HFzKHvJF8lF+EpYdQChswIj7fTaLAJZQIijCAfw17Qo1iRB+Ze+L5C
t7fGkmNkfH7rxj7WXGI8/SLwvqWCrfnnR1SX87cCWpR1t9sM89yVGrdoOxA6qDZAKdlorFy6hnt9
ydUfuEvXYCdyzXyz9ckKxC42LJTGElxxVRcgJ4SHA5+pPjUgkyzZhOD30cBJhgUPDK5Gj7YPoYbL
sHEhkhKblQxI2l3gnU8cfFGw7sXrsRpQW+iqLPZ0PmWbIP2j7CvZoElFwTRzfiX4mwkr8DHghLB2
xp6QPJpC8E1/DK8TDIiXKHOKMinIffYuIFUF5oyfsyDOJ3JFFG5milFJiHX0YONkPodV5+/QsDP1
EsOm3rYb3Q4cDvFSwj8Gxdwpj6IPcMhxhlFO8EPu3Okrj8dGaXcoamkM5ttmIdUk8SayW5dC/iD1
K01xRKJpA66qLY4lMj5oGumWe+/SmRqV9gwvRmwnFa3WMD2yMTpdZ6mF64XDr7e46pEjZaJBeRPo
U9lHvFVTJuLwbYRnQCA7QEv8amFjHEdO1YeNT8tMeaEF3xZZOMwuvXjoNK+xNC9TOSQ6ghoeR0hb
/GRJjvX6U7pVzbgdiR+3Vgfo9p1+u+PrCnJCLeVl8zV6pgayBlX30gbvVRFpJhAye3f14ES4GR+T
F0/1CM+GDR9eWFQMw185mt7r22UMXqGMG97DulQZnSRKVCP3dkiSBIjRscNMnmr3qYGdzonuIv9+
g9rSGrldApad2XLwmIdaGHr3CdC7VYFboItZ4TH4JpbeCZ5sdt7qBg82amJLkyZkZbI0AdNSC5W6
+9zW2kRYFzO4hLWOFqLIeL7kzxZoYjNIqX+NITGCi03Qo6h48VRXwScMbPNyhtTlp3USceyS9FQY
WGaE/X1AM+FGSWDRMedpb2lwMrKQIOdu5tahHuXn4qM4GGl6vLkinORXUKKGlScurcOtIlevhBZZ
1qufW9ZhP8gOqha1JdR596tjZqPQv9qbUWF120sypA/HIGaVR/72CgHGvGBgJIdAXUC8Of8vEgGh
86sLeliAEn0218mREKpxhHJwIcxidQh8GANattl8bnpirjEbkM7klGwlM6Bb9ubuf464Var+nLFp
gqHE8Fj7JOQ0MDjVg1Ydf8hTcCEmrM0jtiELDLeNfHRUepOKGRzHSAXE9Wm/detnH0Ii7w8ASt94
0lNdh7tMpHcibQAjqiJRY4udEhqfF5CGbNoY3MZ6bF3xFBSVPYi8tOKQUFvPYyQrro+ruWju4Cth
FXlti8b6hiGpEwcqB+8LswgneGcmuVv/mCnArXsT25BLvqtOg0miUA6b7fPFBGD4tyYJebpKnfDP
rwYjHcf4URuJuV31Xk9cc81v/oLRJ8DqYvZea/Hy6XeH52ZpgH/qqEOAyVXGn/qS//iK7TPa77Ru
3ryXMBuebuNcEab0UrAWo9GXD/ILx8PXuYHLg8CXwhBIq+JuoKM1bkbp73rGMhBaLF8tlO5bNxBw
Q8Gx/VI2EtniWT90RR0qLYagyKF/fnnzLgJ++f8KYv9XGOYqOxgpyxQwjXQLwJD3DUGFOeE0ADKh
rBpt7J7+F2ivxPH8JpyLWCTRVEx8ehg0CEBUtr360CwqElal5oj83aOdNfz0+iLJK5rM5gLQEh2C
YsUGfcYOibqoIeRwdPWqV5IR3u9eLNqIbbSKltdWwPlrtRdHRKCYh0rHVawOMAIe0oTDB24jQi4/
Xh043KEM/QtvvN4Snxgycg2yMU41c4CqD5iurqOoffCUrRzi3Bwu/paBKrENSRpVEgMgh/+/eZ6h
4J343PVGvhwVyNaClvYQNbEiad6t9K+ctqxuyBYOKAjmICAsUbR9y4Q/IRmzO+7Dl7YzwiOe6+bR
RfSltoccHc8aAX4lNOJsDXwBfPgzvG72SeaI0alQMFHdMcAQ3NSq/eFo/AN/LQBcX2a0gKIXuo7c
YWuY0ayImGuW5ZYwYLizCM7AKWINVmQCha6NGZh3PnTxTheSDAnA//EvAvnkxSNgZduxeRej05O4
Zz3rtJS9QuuCuAOelvdD3/DdBVSLX2vZPGENAIhMwIWX451vhD1uHgHkJtSVMKrwOJGan8I2FZ07
+U7FnDhCn/Hi1uJsNo95wz6T0C+TL0Z2RJUgKzeDPOJ+1g5owFjPCANf6G/R60hft3OU22n1k5r9
0KaMEsa6xS+yz/EAq/2hMFwoXrQBHkllA8OM6K65bxO1KoEW+Dqh91fa4dNLWzDQXuplPO7hhcF8
k1UykJdbae1Pzc6ofuPgUoU9YQVIlrsEiw95vIw8cAuErckzUHrvg+W0PM7XuT5LVfLtu2hyfahx
pMQ28LBlyqpSTE++29iEY52HQwc6sXmyFJlBJjTjapkaiqpwHXwqODOxuNFl2//b4kLUymZneDkg
+JpgKLoSbIwxTscbMHDLOh4w73QlSUKjYJm0PIUiWXSqBjdDjnpTpcJN0YwkKjjEgnLsRwa64m0C
my0lezaTmOAZoPa0T88gLlNpLC8vzioZ47XhYEbJGpRRfiD9YUUr3ywGttWWb16haAPmfwwG82/b
bB/bwq/XgKpQxNpyTS55hfERfAuu0rhaQQAI24+jL5CagK+rxTr/PP0OOK/Sf7alrHNwTQKPs0Ww
zSZ5/NCx3nGfu3ub1V7PDmLLySaoiuj0laFEK0DiXbjdVwzzbk5nQAPeXWtIdLIqvblJK2fhgA87
JQVD+IoSPa25h+tj/By3WZjjX4hduw0qCBwhCbV52OPzlaeSfElsRt0qd2+VnQX/lipgRHd2gKgD
h0B15pIAgw2hGR7+A4xNd1unaM1WarVlzYhmCWNZpQif7+jITqBxNv4OcjgQyye5mAYIXWzSAGlA
hrGO3Mzm8vUVoZQEEDPFCcUnROeqb9vPeCvUj59kBovy7RI/snGaEMhx6cZkNt4gH+3WwQg5+qwd
IlW2Tz9l00ia0UGv1bZ9/LKPJHtIKph+fPA7WT3uxmN8TP9CE4wc960ZnY3UFj5MZYVPvafrWbjp
TXcKxDIB9dqxdegJ+xtSuFUDjK8Qo2Q0RH+xoffE0jxq2XXNRIdrtmCOmdjA6vG3+xlt6lMCcfy+
a9oG7PBuo7ar/SzffqAwxCmTTGIw+VTgdieN3g8MpIjiMxlZpWhfEKvt5fD300oauu3f+NAiQOvh
LFusps72au+Kt/ydJW5XTR8GjjWCurLylcFWhcjJZXm7NeHx1fYYuagZBxEZsjR5kaAkrEjxJ7Oz
psggQDc3rgX/Ch3WuYdd2neCoS1x6v3eO3Q23rbsWetJOGDH7R9j8zikw5h2QicEg5UljUCXhwG0
c3hAk2hQosfUWwvi6PzTNL4IGq9hXsxLUYV9cweRXLw8DavN0DSP4gsqlEj9Y0y5GRnhXbIVFkTq
uAiTlpmfR/CBMxO9JtPAJsVhlgtAWCH6/2tH3M4FX1MWkDfb1FZMWgUUJecT9bujtB9/JhDRpks5
M00yo0vF1tXZjfQseuFmTXkE1t7xhPrfq0QpchXJRqnZ3HZ9ObXwil6jlBYek4bCbpkYXYmWrns4
avp5kAy5aV7OLw+6v2KYWSpnIZErooGPxoWR51nPik5YBS1CUoEjjffwB1hqFPM4ue57i5A8mpME
V6b/7iiKFnhVeZJsIC3HxbTkX+24irtg1RKHSXz0H67QEbh44/Q6POue7Ob+P6GSVCbMg1+qL+IH
IGcdkIGFhKo4WeDvQNzR+hyviEYum2v/fD499g0whqEkOglujfYyQysmxgGcQA2bUuaT/xI0j3dv
hnnPqxlmHFjF8vHF+94Ewp9nFD9QKElG6wYGVlPF6LwWV5/68LnjdjCTOGXiccAhR4xf8vO9EBEA
ihJ4DMgnNuBpWzfIPOHPL+P1Cobcbi2Kdctel2EmBAprrndIyIDQ6GpQf7TQc6UgHPgUb8Zz8WbI
CYsc0KUbIFeIoPukiRrw4SWaxjLduTAt3AsNIiAJqBAUDuJ6heEynq3gBROTAcOXCRs0fzeJ/cGQ
byDAeClpnEdCW3q77EqetNOiKgM0FvG77lRZ9niGWp+l+RvM35om1SoA+IQiVXfDIheGN26avOUs
l+tTrp6hthGQy/tWhG02z0oTxQ/qzguYMxH7TmwjENIrJ7IN4k/DnSnDDj+6ERB+VazUZ8gS73LU
6ktCWJG9xIGldZfZvIp+7X/jL09yltChGG3VCsos5R5dlpIIJcjKvUh3yf+SbHlT9xOCZkaSesVP
m++6pPmaJvtnPflLM8wNKE9y9KjasCnzEM1/ndYSRBoC1d3VhN8X9yVxoyNDNSDsI6LA/ukMzkXg
90Qq6r8SJEsjYvzSra2T8vwLnjuevMQqjFydOfpD5jHWcHyU8KYifT1L0e/9Pz5pi8aUNyRemzM6
i85hx2YFmdCCdjuGdi2agaJSB6Eu3m3BnKVL9vz3VQqvNejn3LBSQeDxcZf+20a/tkT6gnnsR6Hv
nculhKqek3qE723nafP5lf10pXYwwkvQ85++u1KxW4ofxD9YlSJzu/SUqFO+1TQMr2IbNSCP7jyL
k3Zx/ocs7ISY+VnaYYazFQ0mRNqJPhEvm3RqhchaOM/JxX/ZqM/if2DuxvkE8OvNgUl2CkoEgjwu
lKAK/FUHVaI6srt+BapWAWetIDXPi5ksld+8YycQXhNo7P2cgKlJM18pljQ2tLes/ZUtZxMdnQip
43hKF6V+tSzQOEdBjrZKwtPeNq7MAWk6F/mWz16KcVQmO9E9Fw0Hcoq8bQ2zE8AQAwxl8jGe9yV8
59GXE5vmApfZTtlurmp6SZ48eLGvIexu76XZWjvaBzWas5uFrUVw4310Cc6dt+77klKkrM55JY/H
SH5ziGpSLDDP34ShOTNfzQ6GNBMQjzqBTkfMLN1Bty1ckIoKeM0QQqOy+P1mx042XccFvrroy1B0
IHPjeUsratLecmwbreUhN02wHcnTtyOd2uIdPLK5wD5bwpyWH0JLDwg/kpJoCkImuoCa+p+QPr7F
PXelSPfXlsiIrEm4oH0gb8Q3TJyDCvy3f6bQkqPH/FeljJFmPWaF3RTXiIz1nYCiRKQghnej721F
Fzn9LN6EkRzEmLnGm/BlOZOLvaniW2tI4epuhBUFgPtrMLD4uO6KngOXTIYqoWMw6fh/JvKXaPxL
OmIA9RTI3WoASsi6/HrCNa1NW3MEyG+7uCO6LAyzlCvcELYYTy3IG5/woZHGaKZxgQFjJsKMnWl1
PPxfWqHN7YkDDjwPMXw5J6YlkfghnkiUAQEmCx0S8lWPDGLnuWsJNwKkPVhxAXoXtmU4gYb9tw45
G1MwPgQU5VcEnBx7ajZcvw1LYQlgAnicvFcK0A2Cz+49LsMuCNrfn04X01mykJTi1twRZeSNlFUO
sr9io2M3vHvPjES9eLfMRWfINoxoLtpwvEK0HVMZ2Xmb+T0OBLp3NpnDy2+mABcIYezqAiOSbEOa
kGjRrdYTlKfhX+mtqYQmH2f0xJrk356SdvQTBHZElwgMpR9AwrNc8Nk1oQtBNw2Cx5lLXvOA5qIQ
ySbzFd3ymyR6GkWVd3A8i5dpHOGpZ+kT428djQkWYYj/1qjY1pVygovdmIuwFYbmjGfzL44zV+rz
Uh+3t4elMUIIN3n1aSmS9p4QAtd08YOF6Bz6eeCK09kj3c6Mb+szWb82HRB5W6sXJWlMcbwsY7Hc
E7mvhPAPjDyvroCGSVH6DzXjY07fQ6c1h20NBS5H/ELmbYmRmH2IKLBBr2CZHYOBOxT/AFNCQsTW
xDz8BCXB0qzq/Gwro1AUxKmEpXfgoC6NznzighcBrpgGuV7QnVrHAx3oZhdcs40N1eaooCoGAKzh
LdWa1VcHz5i/2Cg+jws38YAwhbC3OGE3laLpRv46jEMB46Fm+kGxPv+W/2vqV6uH3Ayd5tPn7vvA
zvkeX//TbcgjLAFETmXyEKa++j2HTW5YQtkS5uZW/Ne4VXduGtsG2Mu8/L6sk8vglnlBSeMldH5t
/ZPU7sxegJq4l819bl1CmEosGmMZVINxg3DeWE9DSu3GkDTfdxR67zTyVSZFOBAidqTyHdSm5v3m
zLCkA9adHok2CnO6w3IEpxHv+qSEEg20s40b68oTWX0Vf8maTHgkShPFP2PBGz2WoO3V/NX2mAgE
oKXM1zgaa97g3W0rtA+UV5Ndzx5y/u/x96cZavSAGzOtEJ6lguSVLyjjrXQdqdj4kvxNIqrpJ49W
xh6xt6HGHBs2wzYuz4btFzfuu7X7/rC9AFACTQVYyT9lKfNxgSg35f7mwMwOUwHN6rofCfivj7fJ
e85sUITrs69xE0/+jgfxRDj60TP9WHk9MukCqYMYDQ7hrrYE6MY7ILGwbOkNaekn15EQfV9MianA
OMbUaNMv5XLG1LoPmvOATDMjWli9hs2hwARoADsEeF84sW49pZQn9dR+nCgFJQTNgZIp6u9FJKEc
HUzfsx6SBzZdSednF9hURTwYLHzD4aIIYoiPN9q+1FfFljJteBMdpRYNSnyrbBxBeJ0K93N52Epi
lWRrivqSDzT473Z3ujAD1pVG1gqPkxjBeYmmJLtQA5gAKPEMH3u9GZbmYjjNzxOjOZeK4qYudPrj
ZRQSUueGkrjgaXJhhifFFsVF5OP8Ksw8/A1VKRjYekP4c+FWnS88jKamdnlKCwdP4tBziEql1yaP
JWRA4wEj2/p+Loy0Xys2h/R7lA0s+0+PJMMzWTfZny+fvBS7Hs87mqlo/zl55tHusSDxTqqc8JHU
Tyw4BdHDA3Ek5DqaxYRrnl0nPfybb7piXEo2rFWaQntsBKHRxYBFSycmOPnSfwBMJfk/tfk4XClr
pGGSpT6W3MBz/lVbbnRbLINOeeXahwqC3Ea8L0NWsc/LBBGPsdEJYmX+7SJ48JCocibXNDaVwVj0
okAF3mLeLswUXZNkG/2ADLb+QdfAzLtmLkraPzW3Kl17GWZiPUjRkvZPMlTMOUOn06zV/NjZgIAE
6skgZXfL08Fwt4qSJgC6MkV4UGssCytOWm+kUTAupcLcQ1CzL7eF4myXHrePyzpmfuTSAH3AbJ0E
s9WQcZjJ7nBWXUM4roEnfQbsxT2SE1hRwI9AjRD5j1+JPgWtdU2kqFl+ctbxZWJcmEB16IBKNdpW
Ni1nbwlaQa3aiBpmiJM7ACl29Sm7xx/AQ+mwMEqc8Z/bjHOYD/fHVOdlRzq98FEUx5PilwFjTj5w
Fp8rzV8Qb89CsgH6jm0ZDZ4hCoEgAoBy1i3Whz0znMenG9X5kQI1tr+q7o8zLqNtZ9Ilqora+7ye
w8cZJb6cdEQc14DawpjQ7CW/v61OVfEjfSuGeMzKRTfmNh7OABGqYXgT3Z1FHh8m97TllfT41TVb
C/j/h6LSXZOZYg7oRDnW/93JJuXVrjYz5U3Cc8n9AEqIi7E5s3rLPdaYQxvc6ZKeX5d9qnjH8JPU
EqtdIGbFcr3qHv4IX51PJEiZLs5otfU3N7K5emKAn1I/lavLTgTPi5kYfOnx6OXJ3wkDqHYuKD3f
qRoyQbZ1LUsQRYQKltK2Tce8P8KH3Mnr5ndu+3MqIHAQfG7qfBrnspvNHEPnKVD6Rr/vXqqz1PK7
kz0QlqkEvO6Kkev2axMtLtHZ8NaG11HY6Vb6sxyN1WrodQs4jvV2ty09CeKS1ZKl8E4C+8IhmAjt
r9nXNZTBF/jXCSQKbnlJVIENn/nToC12SshKnRMTTOWYkI35pati+MjSlTVg+Qr/H12K4nDyqgum
mvutqmHugOPoyOTDFcu5Eq6CQONKaorkEHZmmq0Yio0qzJZKIpfAxui1mA2ASi5DTyfP9MOiXxeI
HufSXMvcLK/kh37aqGw1F5is5eLKDPqpJU6vTzhPgViJntTzb+krlHvrvCjEmV47tlGufEpntVr9
OpJ+BTnIJz6IXzFZZReC5avYjZ2Mfpenk8MPbulTunWCEtGjfqVVJyFUxRhpHOBbdjqconSGj+nY
VEC+8zK3d4Y6BViEJNiq242HzxXNR8EvJu798ecinauhfP7vMG88ux4Vz0IVMc0u71K4upIcYl76
UtpEiRjsL8R9MAT6N8vsJ9EsDdRdUzYBkPsOOzxCJpb0WBxSXQYPjy4BfTwUoVPyAGSLw7qGJvvZ
zqzf5jgFGV8o0QOdaqcnn/As7mIX2bJegW2au3KcFgrn1c4fsb4mKXNBCZ3P7jglwkyOEE2IArW/
wXOV8NiD3mQYzSqaGP6S0r860faAp2YY7i4+LhslsPa0WBt0WcYElEIeITkPMN9ABKWmPqz9HVgk
joRuyfz7GQ/DJ7qfHcn36rWIp+Vztd2aTI8IlRnSbMk5lJw7hBRHTqpuOSogbG3JeQCgfFwSkb+3
WNH+CdJQl9odiu+tjobCMXV8HrznXR59viVE18T1JycXryeEtSJQW6tFl4BFYRXkkH7JRrmcdYBz
+SYBz+qVl5LT3mMcv0QgRhvnBbaeWAgwk2eRkb2B94bAwhMLijsVDDCNPTJtbhzNyHk9vJs8y+H+
aiiQhrPb6MaFndzGfpxeYkgpzwS+82Mznxbj7CwoxNJ93xkSqrOgSpkUjIjXlKBethRLF5E06JoD
t8cBclsGD6zEpOH5gjpsaG8UZREcm+Hmx/1ISjIVH1Nwq4H6BhkH/NxDF2FQow0ws+D48DdITOSj
JTMsnw7UqzFr0FVYA10INZC3/dfP3iF83y4Z/Clgkpfl5Ya/kGfcRLcCclBWsxBu8FFBH4LC8sg1
PbSv63ouGBmhuxGqZaGO/ok18/gN/D58mC2GJ3jANOJx/vLII2Sb1Re0yMhT6C6UVQVs4n0BHTR+
iU1JX2fwlM3OwNvuoMbxDd4io7oMeEoSkOyaapwFp5AxfoIqTMmXEYKUxcgeermiOG787OEECMEC
CCKyK2I8JX9FyZnnQzlT5AC1pw/saVXl7FeCFQPlDgDtz/2X4uMa33M/7hKM/fAS7SoIBNG/Enon
/gVoJlscPLBOXCBAeutAY3Tnudoyh4uRMEcxg7L+ArDwM6Yj8vPRTsi4WGySwrIhGFIzITbz42ni
7xtQ5l87RbQ841Y2TGjgTgwX/wsqXq3nMuhG4snjE8sBNRT9N4eWnp/4zk2XfjZEl5DPP2OLeOGE
Zxg26O5Yp6bdN9IJ3OUhKUxAQtKqyEh+RACpSdrUL+7YimbXQzE1kKQCNtkPz9KespH7putSyUVH
Z9eqyuKtlatv0DBz2gQvSw5x/Y3Pp7gx/dr+s01dkqhG1UU+ctlMAuAOewoR6c9f1jY5spdN7548
Sq87GpOP4S3/cGuGdTEeoaHhtWlKP0YLjxDUkvs9EQ+vqyajMbyKwDTbOPjZoF35+NXZx0MYBNhR
yge1KEnnN1bNgRWNcMMjC7LjcGBNbAtUvZtvkBAt9laLnbmM7F/UT9vHgc5q5IF8D7ni7m8VAX3h
282Nxb0uUkjh2PmQoag7itSM3NLDn6zWyXpXnAK9i09VCMZYMbZLGYT/cxu+y0GglLEsdac2HOjD
zSE+hyhD2rvygDP64Ll1ov1mPpG/R4LZLrvdcBo8mEKj+Y7TgqRCy2WT1IXm+mblRULx7SXhRuCE
T36Mb7uJD711HGsuCuh2hDtzccHUA2IjQTI6xa6Tk2LC+0HZBhowZwzkv4NV6wOMTup5s0oQ6Ci6
RyxYWqzNGbvHabTDcDCBo8+ypI/IC1KbhFaj1uVSAxkNiY96gcan2fDiN+AM0McQhHhLVYKNRFUO
bdf/kmxWXuOyJTT543D7fkpHYUNof4M2nyrfJSkNEn400TdRCgGZNfCF55bNMgkZkvORZ0u1L1I1
PV9Z2z/cz6cZEGL0/InXQrIMCaTj8BBCNFYkqC6LaDwoWbQitQrn8X5g4GZl6Zs6JrvxlOcbZk5s
PB0P/Cu0/avw7QtirXvyTwqs9HAbrUCPDx0cppwZ/OKdUyQfMH6mK2ko5cg0Prz2FnO4KN8xL+vk
3j5OpSal5p9TKbMlNFVCdFJrRewmB9lj8pzZ1Pxj95PWft9ckUSnSuD4S+LwCqtC/W4OSrnSuqPa
QwLCg6AC8FLDbYXDmIWdmjRiDzI1niOZ6qTAuVKfL6hYMtzBZj1b+y76w8De3BgqcsGRsZJdoSk2
wj64Mm1hV52Cz95GSwGOnRkNNhkhbeWeQt121OHTds3/u6Y55fVA1BIpvcZ8noyV4gVd5PIQJvly
9Qbx9IDf9KQht2CF8P7rWtXrQgOGsTIanKd81//6yxxogpIt7ZW3cpVQja2gCM/0zePqTGEoKnJ0
jWS1/UqcBi8wlCT2FqsFpNKiYFi64aJ8afhCS7eT4TMFTrWQbN7zU0euH+oBbUisDqwl6Z5b/9Cg
gW6ZAyt2WfXcQBKztrZHTWCy1DQGtbPPSbYTPPdgiPkEZ8YaAPF1pSt3fa5bFz5ZPxO4yqIvh1pm
rSjUwkvH1KW/F7loaiQBn+rECVP+V5wbSaXkp/iRFAsQLU8p4aGAfSMmlOvjhEO1cB5ijWkVxEma
i/b/SHmnRPI36zgNVi3nUyfUm/CQxMFNXatlXrCcYJe++hPekK5W0KY8Cb5Z+bbv1Nrz+M7ZNptD
r6T3rnHNjxqFg0CQedPoxZMIbFj6aFBQdZfCzqFgQdRix+ssGbu9auLR71RCgCj2AC2T+nqSz6jA
cuKZs7cjLzE9vUTGH47VosZ86n3Vd0MsocMcmLn4Jr8G1BULlNnVV+NuiTDQ2Frh7vZ64/8FmE/F
Z4sB1Deukae/P752erH20/AUX2n+sGl11G5RiRoYpGw29boADHvmVi3GCtjv2nfBziDYkLwoF+xQ
SjZpJUTOAOO2h8L/ZTj1npQdlflq/M8LUwQfGqhNSnUz/jcLUUv4plVzLsytWjCLxfr9/0EKsJoZ
D0q4BoOrZS4y/+H6GCOggXIAqpMYD+RSTPVJSIHx0kbHmEq3W6iRIBzOrCBEekeP3FW7gW0UzaCB
LOkvMfSErVuJZi3zeq4qA7dU9S/5aIEczrY7k0kgEJkn8fhGTwek1yrtWvE3Ip2IIDoDnx81dJoQ
Lm8Y4cNjUzffIEmqiKtJ4neEtGRJ5qdmcczDOd+ZkC8sg7ymzA7WDHOdp/dQZbDPz/+Tjit6egBi
sggXl1BA0NPAFbZv7zphHRM/c0uyrSAzx4bT6BvDl0NAK/KBCs/NQlJ4TcVGCl0KYP4hZtGj6Uf6
HItJNZb05WMfvH8Zlm8ExTmbFeZHyBcZ4pW733hVqtYqp3Na3onegFXg74y4t+tN1mqz+3/YCrvJ
OMxbxH+YatEAE5YPlQUf2/W2YL8/5tspRSxCIbhp7IUiDVUYYZ3Kdu4gKTmmBjK5qI42aJLORMBS
J9JUt5joNfaHiiGLaG8MEE6tr8N5o9vghE5cUXF2PRwbIScR5fAvjc91VlunjKriu0nPRbRQaJ0m
SkOoLQcztCeZYADVu0z0qrYnR1FjQFTYXoTpPrN/xyiAtsrUWrxUn7lY7Bu2g0RDHT05xm014Mp1
EzzvkfvBrTb9BF3I3EXJNU0yOzWZxUKhrcvO0XPCqo0mNtYm/iqxz4V1fSU7q151ZWBd5O28Yh1l
EiONqA8kGd5+MogNQFaTQGOEo1lNip5BIDUDqEqpcF5L5skT9iBRA0NWsCmDfYvkSj8Jh95CmtaX
tVGzNesbzIiWtLcCo2YFtLfhg0aMH4nt/5zbo28GuWa8Is4f36uV5ei9nw7e043bpK+CI6vEEu39
NVNVjti3W68W2LVZW2lOZvAzQ6biyXU9fPcK+UZJd1rL03PlqGTdgYKxCU026PEwb14z73II6TQ+
NTb7JjQ9BmfrMZ+YOC1ZX2BI0NaDItqGRyuWLOdSJAzd1ICHk0fzhV2XJaOQvQYwLAO+QV4r0XgJ
uZna6K3Ex+F1X7QMy1b73TgkfB/cwrA7QTMPdTzOyzBRkF1Q4WPJx8ngHUQ94+AJpqHERAovc6Bh
2v0UlqtgbwM3trI7C3VPxe5nlJ+9xV4fZSf8nT7ZnanG5uNirpB+Oq337jn3LZ0id7IAvU7rUHUA
5KBBDmXByTBWSsCNMA8KdyUoJFTEgyW097NZe7bRZOndumOEAU+jamngu1hHDswiq9dWo9XoP3+t
Y+PFQBXBU3cB6Sr9Uc92zdlI2LTYoqXAE52sZT5J3WeZFn5t33MR8exhMTK9lzhT0tWIBXKAX/04
Ndye/+wP4BaBilaQPotEPJ45uQtLeJnC515x0FLPtuCcX48Bso823LuQISPBXRKuHECV/yZuXb9t
BnslJxMuX/baMyR2vACZWdt3zNwPAFQg/gOHFG71Zp9lELVBeBXMAa/72LClMt8QcXUqlvkZdjkg
rZZrjRQ423fH1j+jYeFTnjXq/GAgpxSjSFZ5vuUZyCssAOLFgXpdIK5TdYzoTM1bvyThKwzAgT7+
tr8pi39em16ZbQZ3M0k7M3w2J/seYhDvQoZNihhkfcDXo+wIKzpc/v1FkriM20BcZ1muyye/ax0H
BGvsb2jkmK51Jl6/nbwdoQGGrvJ3hFHIP/uuCDgfauLFZZllVr0pwkS+J1IQvG758xG6HqvO/W9c
KycYJiy4u8+FSnH8UehKhQvXFrgHjcZLoZ2N/7aC8oOkubO4sCUq6pt/ynCWZYgJlrip0odXjxq7
xMlk4PQdZUuUpxUGkpHd5KOlZ6hsyt8zOf4VPPme4kWO9mY7ZiZMiCJo+zY4Bj4DlFG/xpUxqpR2
Rdc5eWsr1ndT3KA4SmZsFY2OQM4XpNy/NhCuOZrk7VXIxB02ChfvFVWtpA3F8abrFHvSLlQIHKBS
tXfsho6CSwq+wC9Qx6Y+iesMLyeGPFQiTmLI2RPZY4exIACF6pwCPDIrp2ZsG3C2Xi3lMwUHE8dh
omC3PiLWZKYc1EPqU02qP2UawzgQ/Yc+mMvxd0rKPQpgmCOfxTC8cKuJ4ix8lnXg0r7M2yaUCFJA
mU21PHZE4LMMh3FJ85bV3l3uQI7Spa5XRJfygRyJvbjtqs1dkZI1ac/jvvHG0TqYGPP2evUBm/to
z0AzNGMA67M2SrUPygwbthrLxW9MTn5Yqh6s+XZJCwm1p4seVDgU8Ay9+eSzaRF71pBGGzpB6ERi
owMd+vFl8mty43CCo+cycTELlr5G+OX/q+F/uk8MMkkOGX3pU5fHo5AUH9Mb84OXLcWuj+BJcrjO
LInEh7eXNsxw2ha7jIdZ9HjhfJxq16QkuHAbvlDgtW0wvsrO5wP3Zq7/yXh1ugl9SjupHeZl38vt
u4Zn72TPJ8W7uY1vHx/tMIkvnLUt2F5uJvHdHajRry6J7vLbOh8y7VPEi+4DeDt1L2QVjkKZnhx8
+8VUXbM/cDOVL7ntuRJ+7E37gdNTXqsfvmvmw+o3DcafX4CmYJnzwnphsv80f1RsUZvtd71A6LeV
i2wYeJY2fwP0CM1Kt926sdt+f4A9Qah01tN0cjfUE+eMjwNNb2UsDh/9jyxp9uMj+lD+p7f1CSQ7
NZHJBXvV5uzRpauNs8C6zIzAEKlFemD45MnhvW/4IY848NAry4Zzim+msi3R8/OsXL9xXDC+smRd
HQYuuftTxm5ZzZUmusZ540KO177Rt3mGd4YIhSzeYZNwfZzTlGQJY5sZXTQFftbIp+mbTOCMIeXb
1x3ZHI/vkrSS0OxTsPiUydmi8WK5bPN6EZvnMp7hdLHRTEqYDJaHMwxvEgFGEsRYus7xc0B1C8zy
P8tF8lwvxLovLot8ucOXnyJubtxGVAc0KTqCso2Ttl3WuM5iVz6C/TEOyllt5Pki8pu24qj8XqG5
z9mpoBX1A1mDGm7b15J6keWKaGHd/02NJLI+Ei8hKf7zQM+sGdIZu9V7YdEksb06jc0QvPEunGqp
ZwsKjSBk929/ybA8wL5eDgEsjW7sEYpVp4X6rysVHnYsylZlkp6EFcjJ89VyUHfxVBitYwIhxHhf
39gXDMpYfldafoDfPTa2qD0ea5/hB4asIDO9Ln5RvcTuH5vtt8Hcz0fvL/dLoP+jwqT9g6pbi84K
P1Pz2aZ2DmZjX9vMq222jrwJ01XBBOzubCaEBhHRg59SjV8xEEveQDqu7X/YZhhh1wLpEUy5Q5Yy
dY6uNL7dk3HzWSGvyWOvKAW+KYof5XIbV2aDanekKch5I4eaoO/kF777tRDb3xrs0oImvPl9OBgI
iDuYkXdJF6dTYlil0T7ANr50HhHi/9Zg1CfQSfmuy0c7A+A7MYPqSd6LEmhHCiz+K7QcHlKlYUq0
xue9+qLnP3Wd5sNiuIosh+1GcjAsICbwUAR3y6DO10fzMlSEJEYCzy0pWVXoOUanboi2UJeT/1Wb
wBitARSz26mbNK0QyzyLcoqA/8dfOqmJZ0+D80w+8HDGCD0jURNqOOj7kWs21/2QNhbG72NkWE0h
PkZXpjWSqfs5ZZWmYpL35Y+hmTXAIPfdr1n1lj4GJeNQqP0qJdR+arTlhcn2pkMD299ik5b7A5Zb
yKB87LlOmYyzGtwh787336S8vd0lzvkW2N/muj2zy2q8+YcyOdx3slsCfBek0CGt52VP/dTtCrUb
RMM5FcXl4jkNxcCfQyyg8FRVdBI0iQ2UZd7qGaQ3439z/Qaythkq+mdoeKb2m70toh/1zIbVCTE0
hZUP49Q/DRswOkY8btG43sKuEccRthMFPkAo+OH3vokmMV7YpWC2RIp8DFsRDKG49/kzTPTFySUe
MG3l0Qp+oqPwqx1XS3dwpo1rr17+DdLN3F4rlfZ3yle9HPTFsA8KlhUJsuQMjbRlwmEQa58SZ6R8
RMRx5T6MKqbgasf8PLDwQLSZu12COszBRVkWNRMwAV1JCSDb6NAdjG/NeBoyYsiGLaUP+GM7gNHS
0L0wteh/r+d6TxnB+YeASoceJGXYaGsJHlcEZT/zoLytI5jBlgU+qN+dfuRBDrhtCRIchTxL5j8W
fZxa3cAXGUPZITaSeaBhaChOkXaALaRJZ2yJHnhCem8KPjN8AwyPTef/lR0kIlTPro+hpHTD8RtN
vyM82kuIKZpiEW454Ramsm2oD3kFFXL+2lmN6cSoHFULW77CJsv2y0FVEgwDkUj3Qy7QinPxHnLp
urZMMXCE8b1vOP8StMcGYyJkg2oln6glMwl7ItTeTwJqBTGI9r4vO9J8q1Ic03Pk6Ov5BZH4tci+
aVR/BPNGURl820rkIQ8dOoajGeRXHGOC3MiniZTp7VJucaxXMZjr9FcoIsiWb4JNNLc6+qK9Oizm
R+4KHk3Qr9U6jj6DanAQtNjM7RcVAvhSEUfAjROZvuFBxCqknxINL1tnqSoTku806HkQy+5JZeNF
dRpYccThAey1HGhp+R4HO7JR4EbaNcvhVOIoXN4MGocEFCRPmz3fqjj+vIuvO2xe66efbmiSDWXO
qeSALI78ZPv3zfkBsTSgS+hk9IBiQ8ftUj2twgvMkPIPj5QML9tMh6aLITwKa2hB0l8o++SlWelB
Om53TZbQiDZ3tiQ7BtiO70inz8KmLmeIbmzCqZgWrl4hLSlNc1A3L5ZtHkNuWwz9saZXJ2hb260P
fSFWBZ7xmckIOgdw4cy6+tdMdzf84ZcC0oj69eM8kIJeX762zLTM8GIQeXGHe17/umbfsy++PPKC
6hKO6lmTvZOkOmYbmmEm6cK/q5aKuej7JQ4ntnMb/CfqUroLWyuLbr7w72i92SMQa9t4dAeFugk3
zeIjF/Km6vsYjA0lrK1HgyKesWxzgUT6trMfHneaWaLr4f1/ldSjHEGB4gM0hD83yl8R0tt4ywnb
ADU7HXUGopds2PuDQlyiZm1iNsgzBYqNmmeEDrf8TXkNH0kia8Vva11Jwvc2AXbTpKRWz1kNvNNP
ZTnnxmDBklsCWXsQ46fRLuN/EWT+LBUE/tM4nR7c+QbF6d1YWhBXr/6EaL9dzGeoyIDGN2WjC3ij
4Qj7wT52qCiZ0HDXpm4pEw+/V2BN3/koy9aU+HI5M+bRKpP0zJci6gmtpl7XmfeKR6YSu2DTpqWE
S5zvIO1QNBuWu+cewl24aJPKHZ8lGXze7lLdRvx9vxxWd+78oLDoQf4a/33qnAFhpf4OFwwFyeBM
ywKEK2u/hcDHNT74ecl0TnUuIZfFLt8YSoxLgdLji7r1YlzSH0Su/BaIRsPz94TLJZfvn/w+tcNG
fH9V/CrHvoKm8uhamQ7N1z3Ood6X/kuQBCdBD7hhpJwhSMhfUH+95nJe92cqxerJkjKkRcRe5zD7
ApfANzvY1WXsAXr4HzPZugm7X66fwHRziqf8ERtLeXMWJLNVsQE1WnDu+Kx5C/A5gYTfe1Nwv2ps
cs2oHvlgkjJSvFvVds1z0KZ7Wu2LxHdvzHGJM/S9+SdrmoB5Q4T0XW6Cb/QPloxv+sWiMRmR8eYc
8lWtg3vUzF/tMjeMYL8y16cSVBTI/DVEXqt1I4UtBaZ6rL1jznS/P/BN8/6MZYxikIYVnipsVzEq
sW9Uf2qb/e8H3R5TpNpojD5sDJft7gr6yAxoTrm9eDFSVMzIbOLuGhjekRHTVzAXvpAKmojTR6kz
oLjw8m3xRLvfMC7uaHToKdJVAd1QJ9yme7gIGWQqjv8fAW/yE2R5FNmNFBA3yQB+4gLXQLdvg0aZ
EZ9ln2IBeSeYT1KUcl3NODumGURYupmulgP1EcKFV0jl8KKOZymOMXnZB94wAj9PNejM6t2fjb4U
Ttcep7aA8W/+nsxwV1rq6va0JYEY8Fmhwv+6K+fE7yFfM1PsXuN4ofnrF/j0N0kP9j0hngFXTHsR
wytdQhL6g/D0bPfultgXA7yCjA2wqopkfIppp/I9u5mSNTYugBDkBgRRFNMnQljBrYAzyWxkhBc3
FjersHImiTSpBsZcPLTFf47I07OZlToECg3tyfmgDEOx1/dg0t93EYVKviUA/eJdhBQg+/+HVun2
1LcNMk3Zad4HR57GtcWl4AWHsIDMkzL4QcwJbB1bJgEQJJzKMSr+8YzlkEX7A1aqhCP+5Iv3qrO0
TLv/JzGNQ8TK1lDdTqJNvGJ4zLFC38X8CP33Th3DI0J9rEsFt4lVzZJxq2mSNqcyou4HACsw5gVP
CNxESgSNXJ/pTM+J/7jHtPlcsfi2NqUksJri4mggUqTw4GvQ3w0VEHLc4sV32rD003BzbM9Ez+qr
OzZM/7vivRr2e0ImfKAp0+SUBJphuoOuJWNgVT0PzDXKNiIUzakLwT1HNQCSM8C8Y3fd2kVdOL38
cWF4FY5lgaMi3SbOjBuyX1GiWd5cWnFtPl1TOqK7mHRkZynt996xFyndkCQuDNnWtUlYNvGkH989
sOoXxXrj9dJkI6/1QJRXKrtuoYpCMiDOjlxOZDch9GYsFrc3iSiU390l/7feeS/64JklYJ8fHvoy
qSTcX9dmqTd4/BloroARQnv/B8tLt+vYIkrOTQlhYg4vAlH20MAK6cBxWP+/5W6KfrTSGd2UvyiN
n0V4L5N4D3Sd7kzZDSQLuSIO5nXN1mT6nAzI7P/9q5FL1GHf+hMT5v+W7uriLz+zQEpBXIsmTIGm
6nDYXtsh1pULszz5FG71g1I5p3fvB0RltDQ+JP1hgggoBLc6BJwnmCN/rhOByRuzgSUikvC7JZfj
GY0/YjTtTkLOZqjmB63ZDZQClogsAxwKbzJY1tHvb10D0DCoiuAHDgNZK6eIh8Mpne4CrW1Dcy7+
NbHpJ4K48Zg/DsfuTLq82rl/NAjm0e2294+aL5M/X45vmIIRMdIz4bLhA0IdM+lHw3CuCnfajAU7
JxwMU7qxo+0/UZLNAEp3a2re7I8yerePneUmiq772m9cKrQLt9wVgYpYaP4PHs1jyEp4JbplXzAi
zrUpw77dcvIAOcKw0NVL9F07WS7oOcxKkVlQDNe/aEj+FdYmt9PoFMZiV6aOzuf4bkWFF3rT6wnj
i7UppoFsZIW0tmOQQIsujra8VEhBAhDekH2zmp3eTPn8IrQ1ryyeaEbK9frhrMyBzy82KmSCckAe
AeEoEhIU5Xp94TBemB5Ge3FHFx+hzqRfGWZVPEFi+XA8/ZH53vII5hpF8n087wxny3PhkqFiRzv/
ZFUEAUv7SXJdfF9MuUF08zECdTNpHb/4+NCPpEoZfKaUvCWlywxdFqiXZ0lBsKbTcjasP5JFzvga
QBSuGA2ZxsV4fBVobrFop4SxiKHkF84RYYKeglKcIgL72GrZb9/75GFTKxqJ7DBI8gOXNNK/dxqn
q5/PtC7FOx7x+IMJJZiAMX3lhNF0jTHB2QO+obg017F7xCzBWx9bXdBs/Ymmx/Ly+rg7wQxDyaaj
aqgEs2PV6PG4zZnDYwQzy/AxZNMYzf7EwZRsW4YBPB7pckOJW97DZW6hm0SV1zptqHOyMPt23Jz/
GdrJt2wzAvnhceZyk8x1OZNODCnx/j7uuGA9T9+5ztJRHLfui1McqDwPIYBs6QFEw/p2p6KK7Cof
zYEN4sySwLwlgYC5N8wu8jCALzKC5COFoXWq40RFDV59XvcE+1OnytIXLtSI3bsbB+ZoUQFmsWa5
E2KirEqR9+3SZ2pN9907akcdw4HN5BkHdQdwwzOfkpXMnU1BkCg0ks5SIi0rTlqoQcXMyPjdFIl7
6TDzRlCpJmOXMz3CMru92bCANxX5PVTA+NUZiDBqCu2xVgP+SEFE+crCiqr4Ciq5mrR+GOcv7r1k
ckYq5U2r49pnyaBSQf3B1SrCrKTrj1kkisfzEYyoYWu5fNDMxcC0V8gjdGpnRIAwL55VfKY3DdPN
/cJ1fw9W+9lNRhAwUDWrRJ36bFlXnVfSk8nos4VFF0qpAdVVDVwB31r6lST9RdZd7FlhDhFW+pYa
Zd5/rRwKZpFEMd7KAqbqTseI5OjsLAW+G3wKcOHJRCMgskqEc8otP881qwJczbFjCbgZZeoiJK//
UTv3RBK0aSl19sEqFB3uJyNGm8PLojabY3H2VNih3fqzoslBPPug8gDd0ZGCTcR9HGSEj6xBsCZU
jZT+N1bXcE+oBaaaJR0MM1bP79PnoNh7og44G78ByrT9Bt47ho+LkHMwjFWG8+gcjqJRLONCC4P4
LnEiaT4ryZXoVKj9QDyqO0LvNWOKxDWb/qtDFWT2X/XgtDvua9kfCcIlWXu6UlblExu4+hhi7Yc9
10YZQFRb/LvbQ4ulLL5ZPQLfG6lipe3Jubr8Nw+YQef1cVyUIM6RyuteucchfR0XQ02cj2z4WAs7
Bl5QmnRl3E5AXCQCjMrs2QBcts0JpYYt/EDyOOYQcY4nNOuqN+aM6NhH90m6RoT8dNkrk6HmrHFD
V8Ztwws+rEYyMe52Jv2iRDrBXfc4c+I0620V1hTnn9meFQwtKiQT2Lnk9q+QvnclE0M51JJtJyP1
bbUbCQOt5Nuvh4bh8URDrzt2RCHxLIU9SCfRZRqMyj+UxvHdoycbF5MW/P8Mnua28Jy9k/qxH9Yh
3uBS53BhQRVaij0EnHsTJTF4E/BadYuQR76/UcGidI9ZqSgHunKm0tASfP+Ny0vnqJRa2pHOCvD2
XpV9eXcZetS36+d0vezHhLxL1fGIr4gHFGzA3dEh7Fq2BKBckpc07bsxzM64/z5xT5DH13jwJIGh
RLmVId6cvnkFFG7riajjy0b/hfCq6HN9MYAXBT1uT3jgPn3RDLvGUzQCwtjLgKjKEeN/BqKGDeLS
4xMKnqx7Lp+zYwiEJxsaWosEa0qEij9ggudPyvu8j/DCRVnsq1CSXu9hOsnwGgazoe4xjLpJ88Wm
Bx6VC3Hht3R4ESnQV7vC7OpgH1f9dr7yBKLUulMQ/SuYxCbAH0q355XOONS3Z/0LJx+PEp/EwMCr
hW6e+KDKauU+96vao9weauXPRUz7dkAocs5u75FGSDUxVhFoFzbEhilXqTQ07+xB5ma6zSQq/zpM
4iAAs1wls7oV3H5iyl2Jdrd0wGuEGOp1T89rKoRyt0ZJPSXTZqEDJhGyfzZAIXMWCyXBGZMeOyj2
ozyk6JcciYddLtaMDNl3PqExovsDiPDV5WHxm9XBn0zikNgbsFhVgPNjg360hYC/YLT+n+spZz5Q
sXFWQ8JvfWdJldtCb20QrzanAkl6pMiBHbqIaDCrdvwG1aVCKvfQPZvccUOU+60fNGAQWizx5bH6
za3ZT4OC3EiM/0yiuOpKTVXsllfObJXRehk682rh/UKnEL3hK8LSFVP7/l+HPJOXla5uYDVqYmak
XlIRK8lSmKzkskFjfSYks7l7jLzpuFipaqKsFAcsxDAsZrXQeu3u7wbFCgHG7NRm76biTE/BjW9I
RT5DNQkDJ4IfQPFl75jlSSngJ/o6xFSJ/INHLBG+BTxtPRdeZqflPWXPrUx/lazpaXspdqOfUmlO
Mgjjwtqvc6YmkF7GOaeFkhxi3lTxGJGGf2kRcgWyBLXR0xTJQ840ou7imH6edZpeXhFdMotg8X6c
pPKX4osbHDiHV7CtQtwzOulV+IzOCBNDsmTUFYhispAQ/2o+Pufk7hov3aSaoEEk5Walr+ZSoK1x
ve5FFwOI4gDYMAwybYxrm1ldMo9nT4OsIwQ4oPGI57/QdiuQ3bL3zWfnajAuRI2/tuoLMvWAi+nU
5dYSGyWeHyJel1cXgwDeR3yQxvi8pafwRjoOq4DzFPeNRtge/QyK8UvZoZBVFNOQ+FYmdouWS3aW
JYXq3yBpf5Boe3JmyyAwvursLLfC7DLwulg3N/pUvnCxTl/DJzKIKaEl+kcCYBNt5NytS6c31Jyf
4FfjT7AM+ptfrH0hPsFUIGf2mTeALYcAky96SKk1Fy2GMxOX1DJPUo1Y/RwtwSYEqSWw4nMuQBvB
RWwjuCaN58HXj1/7JpnPCHwebFfPe3HCJW6vWsIpqenVA7U/Pj4HkVwMbN9rwH6iUOMmErXOxA+m
hP/OvlEswMtNApaTuUiAfKnbal/9zcK7z53tHXde5KPsl0st4vMB8mwYbfzyp6FQA+feeQG8/MU7
cUEsGsGVf9Q8W4TwEZqAfxg6/47ihu/SpReWds3LLI2rxQwriF/QYFphgiykLhJBE71C1VC8uuej
gyvVF1zPOy2Ot/Q5MnPb9C+QkwRlGj3VDDN7T4Xw0HHJAKXW8DoeUzoZ87MdXr4Fq8vSgEWTi4HP
ND6VAgVNsOIlR/oLzXN2SFdNVBr9GHfSaeqTyYX2EeTWEc51+l6d5g31kgjKrqVgVGHT1x93bPgE
58S+dUHPAWkdUPniY8GMAnhdQ2U8Dt5fE/fpAN5nBeWTqrc/F33BcAXUlTE5+kngULXgC3CA5+XP
NdVTkIDkuPlWdSRoEh45ydhGWBN7iwofoCl9Kfe5R/wlskLDz+nC4XHP68AD+azn7hbBUNRfAG1L
3Ud74fyOR5xJuwjFz/6ge0Tc7gmeSfGgzQnQk/SR5J36EIx7PR/OY9H6QOmjzJZrH7RjoJgiaLCN
esLnTTQXEydNYmJHVhcVbJ63xH14hxbxlwUaH6l8pNyf5b+CzPdxgXwXjZ+3KwWirTf6/wPyE7/d
YtC4aOwseQY4+yOjEi7NtXFSQ7tbe61DxIaW2/OXv1nYQpnz56W9AdemfOnS/X2F/cQLFoAAKtTJ
37cjHIWtFwLXRjxt1pXohm6Ofb9r0uOw7qURcuLSxByaYAvUwVD7or2s11KO543ITnlbPHG7OaJ8
nn7PVAU/zgxU5aTeKPYIRuGfY5yZyniZVhQ9h/wb/cadYs6TNvz5N4jvt/9c6avLN4UVkMZK34Ol
0e+F6D6e2eSwdHdvk1CqOFcvzbpYokfMJXOHwdmFiV6QqecLAC2p5sSEcAWj16CK4aF8cKyb+Kh1
ueMpgSilP8pLl8Z/OzdaBZJVgP7CO4uis7zFP7eb1uaMgBCV/5JoMZYfKbDKW7aZXeqwq23kP2KM
IQUZrRiigKhJ/xMP5aBYMBYZ0Uu9bPr+EniNA7QBCrOFfanqs+ekby7QkipJwnyH3F4pM9+QnQ+v
cfEd9CGoqutAMMjk/uBihNY+qLFllIkWCMJK/cYsLorye4QlVxD2pUUDOlnAqnBo6bvQNMOBnKXM
npjNcPAySnANoX/9s1yHZC4m3QoILbo2Q6vPKkwWvqAc6B+83P0LDF7S3rHau0ejMhvg625UjcGm
3tnnPcpHTYdtSTKWlDDu6SFU1iBLi+K39aUtxDHlF7WGY0ziJiP5GoCEXlK0poRlGpxLTsZTCjr1
hC8M7v0bhraQqDJTFdxaUjLi9zN6C1Oj8deHfMz1o3McvTQtGdy0rA0H+G8iTBRp4UU0qa11Q7Gc
Gg8EFCnSFqzQHLn2NpBsp4UYbIiXporNxi2QEVgJRTBbtR0Hc3m1M+vveUo6YcScxio3Wo8N8qJ8
iBcShSXOBOxV6qk/O36I1lPi5jCBN9T/EMjF2UwimFZH6WzgeRVqxIM4iEhhyqlcIANSkJ3nSujj
k2Oldttb49GFjjwVDPJo1YrKbNsk0ytD3traKTmKWykAMqwoQ0/dW366zUVQ4qgiKu2+BC1kPS3a
ndI7nJwsD6uqNeLbZaPzK2a/rEdO+VAt2PY1SAt96i6+kG3EjLe/ke7geJCOuKuy92zUjzgKHW7K
tIEKIxifZ9A8r6KnrK+JrBYLH8ON86bDBFgtvV+ogmtD5nLq7x/4NjHPwvCidgM7T9GEnpJOegc5
3GrkfmS8ZwBtnbdtNOg5itVNQDK1M8OYM1e2AYQZDbiYd4FYMFhPGaNqcitOel25tmnf9MIfIm5P
NHEgULcnmLWkOSbJVda8ETk8JSO/N94bH+6dUMZwM1IX4A0w9SNDHxDJjDj2l7/3rKYBnMUyCkIQ
g8rGc8q/1hYGaiylGQkJtOtquJmKj43viZFtU7ZEwBcNnUzCktBJ4lmBzzCUZAuUt75zHNluV+7G
c1jj/daFx2hYN83O+117LMmIXybrPbTTEQf6FDPUw5OoapIytEhSdJQH/GFZ9J18zGRZanCieyK/
rla7e0F4wNWyow1CDABU+9wFUBTsUaADSlpubFWSd4SDQqP6pO6uL8XXSAcvOSaoApw6jlcOVeOV
eY0kye/5L0imGrzAX8IaIygNthbwrdesHTGY8t1IOk93dk4a/Kix6CB/HCzN8SlJ4DyzzZUuueH/
ULHVwcXq+P3ciQev4K2+b663jdm/X/GmiolUT6GdXhrY3aVERlOD1LFFmrx/ydYvUZiTR27vyPk9
sfTcHWm7+2rPgf7niIVCL3ZXrOXUw8uwWEzZnxGJYA2gBR1dosPXtVAgBvb5i86DDnLx5r5M6hbR
RfzKjQ1JxnsAwxgBBhoJawWwTTb5WLhHAIK6wM4npFp7jbl7DqMG2vehvtKd/repe5Y3Q8OqRRw/
CIgEyPe/DEEP0CEI82JH6NRrvGtuL27C/skVNDp1oGGy3urJ7eT/c15k11LE+xc83VfCCYSz8ayC
TgELZws5tx6HcH1A63oX063BIvb5StDq3o93UBZAg+yZ9PLJpe0sNfoy55lkFESxsLgYmSqWRUU9
2AKm68KNlFAmMbnxgg4duhEWlleNoXJgz1gXNymkyAKV1NUVBJvHNVq1v2WYHd25DwB3dGdgfKpi
8q8OZHfJxeNKXJz+V9WKxwWJdn52OxUioR8dkYcUvqbrh4EuqvuFjgUDYY8N9PlOcdH4iu2NdM1F
DsYAvxVFBGtnIEpiZ2L43jNA4DSQdraxXqBRYMAuNF5VBOAw6xybIh03oEDSpgxztkHTJzV76OFB
TofzqvD8Lvv7LFDLOb77VOL8CfUncaMUcNqYwFdWlu0d2db3mztxZCDFxBc0seSCIvVrKS9n/01y
GDv+jpBctDWRoNoOONjmYSbnBkwCdfBO9xtNEfBE3tObr67xim8GI/+hxjz90QtJGP0eidM6aUSb
wM7ZnCe/mFansae9lqqYZlrsoPyQ/UMuG2DYloJxKtbN9z4sF9Fq0MfKLV2oDgBqVPJEVUIr0lyz
VzBn1ttoGhymiI5F6l28A7yohsrs3jQO/5H022aXhcHwZOIsWSV8rDinJpv8IeJNvdMM7AFpkzS6
Ki/cAIW4MyyoEz/r+51GS5V8AxjWxR57B5UcGbBiwj40k3kKC/jAr4AcxcunYKK2s+rJz/AbB4DO
4ZDIGOy3O4e2mV18Gp9rjdWatU7KdCvosiLvgUoWVj+qUJQybdJHgh+QVz4jxd+6QAmooFYw+qT7
tai5FecfJGQcrfStOlSx8x89yMSyCPRpJDnRe9SJFCqkknn4K+MZcwO/vRirEQEoYJmKPRjgKH9R
KeHPdFf3mluivzzFIiZfsrHQhfX8Ot6e1TmCmyjKevCXQPpG4TLAGfKaVeB2p9lCI3slX6e0YA8p
UkDtKXRhUkRi41Smb10PNY008W4weNN6IU+BStUzn6oNSna5cORtU9sQBx3CYejW2ON6mMYAZQbf
KPy7AdJiLhX2spCgZwDhKp6ZInD2PeuejNEfO45ztMSyctvQiyhEFt9FwVsoMA/mneIc790KCLvP
mXyRst2vDhPbn9rBHXU7jOSlFvlcNLasYcd4ViwKfR5RtxzAegjW1G2BFYiwfzRwXke26hqV6+YZ
oS4PttlJXgKqFM2XpyRbet6N8Gy2DAKT9cbQv52SSveDcr8rJA2EcSVZ2LPeoudizHGWoawvSsYn
lkcmdErSe/vPO6CSro0uOXnNPbfhbW0UwqMIa6tAkG5ajiI+XhbnS9ZBx1HcvKhJ3Hr9WAfXu660
t6Lu555BHczB3BNj2IeylXdKqG0oDcl1ueBTFdWA9J94+aprm51Ui5/VAIDmvKMst3928m4cg3/f
M40+OtA/Xd/YyGfS3GWSmPZykq/VwJnjxj1s3ZfiadNfLc1GjBBAoM0EA0ww3/KEw1WiqrsvqeZO
P2xQA4X58a+LMmEBDounqerMAvvnfhRKo56YNeFvTku/MLL2xkMNUuQ/kIfWR2fhGr7DPTNWLnIW
faZREOjMxmGZja6WV4JxKRlAr7B08SE9p+/z+HcEizkPAks9aHp+wj3sfcxtxQH3J8DXye1G+9Ew
XNKPzI4v3tJYNx3QnMYfsVZh3SjCMz+RvQYrHOSMnUSe71h7nJDjBTtIGQSbAKKzgFrKf9RGrkZF
qpGUJJSYhvEF+OyS6jsQFb7peff25TUlS1VSPQb6ZoLyXehpKB0wvwinrRRztNkosyMFov2sNrYh
XQ4ZybyQkIVbtkZnOM5G/Oz0foRCbJluYcU4rYoFPCO6wG+LAhDMVE45+opPE/0WCkP+mFnlpCwm
bp5EgyjQOUOodda3yWxzSjiFXKcyaxj9Qp6J/6/rm6GOEJB3CXRESHTdb37BfKAiqcwQG02NlfbW
5p1zL1TEuk9nOGMeiUu3IUws6gjnzw/LrtUBcsIdNceVnN5PUFM5P9m2iI+s6bR9iL8YUR7ygE8/
kI2Qe9TmWOlgd+wqwkrRY72bEObvOzKpII6jb57OdzZuaH1nL0ZnbBl7zl2g0FXSu/Q/Vbvaii4X
Coo4WVeVYBqCu/XflOTaJw5BXcpCnEo7O/iJc111L8Zi2LBYv8L9h+y7lAMsO8R1SSpJyz8/HB0O
o6gQSeWZTLM/KDlmFqY1zjaYYQRuiORKLLQ3L3CzbAaLYnbk7dx8bwifN0W3KciQiEjbENaQQJxn
kw5GPtkTTjQeRuDWtUnfIdbrw0q7uS7UU4ZCcCa/jeR4JvPGkFVtjNaRRfM3v2zESMjq09d9q6Xu
C3NlHIGv2z3zqgPtoMFot45t0LU0v/ZPRtLOLGLHHF+VUuVGh7ZR9uUrGGQ8QqMYQRmJe4XJhLGV
0qMsAhV2GuXPR6WflqW9pycpLsYDFsaWLrJfdVKmiWuDILtBvRByuWWdG8/4x6MTDKNY3s+luyZY
ho179o4h5+tBFDco0e09aM8DtHGrvAiMhzSd8474JVwfkp3uHeaAPFWkAMhKJPQph7lzv0E+FXdD
SRkwtq56L/ejW5WbrbPXbnRh+vNqzlY2cImepGYEhJ37wHnwPA5WespCFLQxDsbjvLU9y/bksMpG
RqZ9QteQ6mujhJ6zdivsTX3UED38e+8+yXfvaiXcO9V+/H3aIBMJhNXOvS4AalhPq2dm8k3q3NTK
6/g69Qy6M5EFEF78gp97igKV5gpNA9V/DCvqghm0W1/21D4sw4yX8X5hpdoPfgT/q42BDJVHvSL/
3R30a7B7HJgo5hAp36a4s33oZTMZiAbTafQFjgihTYeEGpRY5hh/V7nExdkCDNd0fZqaXdtqUNIS
JZUiau77O21KIJDZf5Cku+o0frSxcIj1VTTcCLV4G/+K2fwPpt/rKkecyNQJIdN+IqJNhHt0UWVo
YQk6NEnMcA9k4Uqaqr5ej1G4Ar+/sf5lJs9f873/xrOBDISBYZ64kG2DJGRvulMzzCMoYkmeQ6n3
tp0ZKZ/56YZhf9PAmIVjpbcIv8w/f+rVBhkIfZPjEHcuLx68rEAS/0u1xFBhsg4VELrTtm6yEN+x
lT3e8ihvw8bKpUyfay/hsfHJCsU0OccDr7HYgYFXsFk/iAr/EyHpQewrBAaT5/LZ+zE65EOVljRg
dl0Z0WHtZJCHak4b0Nq6FTa0aCSedYFShLMp4ygyQV4CyUwyQGYGMD60XJTrnUuUg0ZCeqNfppw7
w58U5lM9XFxqInN+W3NffiEXUvZM4npYLrrgKGtE8yVev/cyuQtBuZ5px++Mvc/KohindfMeSJIm
I4szY95cgkuqLcVxJhPNpd8d3vdY9aitzx+fT862Yu5BvHv5syo69uW1cmQL/0ZIoWkqro1KL4fq
S9Uim9P80JQnHi2dJvAuUknu3MUc+IcV2QQcQx25Nx1o6sUbDGTjMuPpevRx2cVCFS+c+AGMUkKO
ycpaMEVudoiP8Puiw/nx5Mdv5OTwD+MLHVoiWgOhHvrBfgQuhzjwQvvkOrsc6h9wY6ckt3The+rl
DXR/laxjdXQEx4p6HeBP9qVKNs9cC5DL23+kaXCg6SdnZbSH3H8aFd/F5+SkCoPuagcJnZf/bIfv
l8b6zbGPRB/n6dwGd/9Kb1bMB932b+zzF8Y2nKTvtJWGAz1Df+1hwC+3PE6mHfWML9xfsKFthcX0
8tlQSAe5Dow6SemDmKZyA1de0c3k44RgkdtkIsbYD2f+F1PgjHWShfwxqWIvdyPYSaTgO/VxTFEO
jlIQd97R3y8cTyi2OM8rlaODCmxuqpPUhdlTedEPWd81rtP8S3l42a9aqjudSCP8sFXFweCKjz5o
sqaRBAHizdgii59hlBMM/x8YSC0qkhE5VqdgkYtFqrzDkzK7/xUIu3bn0kB90M1B6a9LR970EXgY
OonN4AWkW44Zb9XlTSTTWOvLWXvRBwzTQMEDFNleL/GcXMR/AfF5/YBRW8AvtBfzIKxo4jP+7y5M
PeqaXwZYYfXTA6jb3011xvxHO/xZ6jpe0Uplt9g+Blj1AOyQPzM1nb7mgJfhjE59BX/8JNdZh+2W
ivWQes0VI2s+ZWyU99XZ8HHcZA8/FPnJTnVy46Au5LRRAMejRPRVa4vkdxf8It+TBg01H3U2pFxW
XEfxyhns3LgpngezrZ8RcEBUtbShvUoar3e24wizTgetU2ecKgUzSwuaHy3yTVaihZVn2DPDMW4O
KenPV8MQcECBjvyeJbD2+ic8s9oNBvJkAoKsSM69XyP4Wk8Iaa6RI9kV4esmVsZ0Fk3zAFeD6RG1
8iBw5HhXnF4RCC7rNGWr0QT736wWnhL8V2y7gn2KYZ0Qq+kzD59tLcLj1KbUg1fpxaznjS5zN1NM
KHTaNvc6kj7fvl1RWAVacXxEyY7+Sa4qAz1sZ5MQ0UPs468s0oAOaLal9sQUJu4JltDddKsxmMIP
3XcAk6sJw9uQrn7hpfB71ELdiZtsgWOkOyjYpHapbUAocPVte3KCkhdw3pprxOAXLKzeEPAjIzEx
EGuVWGQA8KmPisLc0bTy8iuxM4/HM6Sz3EJ9+Y/MHNLXsKBXczffxhhNUgs/gnrl2Mw+30h4cb18
aqIXgB2n/2fCR8O+ezGlxKVsUl0P+3x3DjVff6OllEqkRJi4EAkwt2/z6zOmL+DD9ZwLZwzSAsHP
WTr0kdPvKji5bvQPy7TTNHbI2LFgmNGP0BaFhuf1SMv4f8AvEPSWlUVv5YiVJgHyUrgH9Tupccyw
7og+X/PejSY5JJc9iqEpz5kyuDV2vpG9lhUWDn944MZK5eDUmwEKeX1Q0zYUD/AJeGPHeK5WVuUd
rRRZEZBKQpq2lNjvQAvHCWb2YilscuXI4O0HAVxMCwckm3BcbaPMiLEVdy/6KSXbGBjSmTFQJWTC
xkxqQyS1Y2HGl6ksmttCoOgOm39RiVaVd5S17Q7D/x+nOCaYFKorphKmiRifMuLSz2T9Ja9uGOPy
Q9k8ogT5p6f4z9+9PRdtlAIVZBSZfG03HVWl81jcMHNIx7DG/pxSWnl2TQe0SbZwf3RUyOpOOEYj
ovLOj6BWE74z1clJffT1euJcBLUTX4/fYBKPNCI916yCLsV53nRzn6jvoifC5nseDlNL+fngoKH6
C6HtUjepEc519L5M+GQWkOqj3+MrRtn2weA/QCGfpU1Com+O4sBTKrR9SeVTu9VGQ3mYQgSTWIe3
c6jexJ+xW1TnBdfIj4U0tsaxyR/P/gssKS9xJmZRjDQFMYsTgyr7vivTlVU4HhQ1I0Aiwugwqe3A
0WdMPt6GX/tYEMa5PLZvwtkKcFfPTkNIYXwF4xerpC7SaQjgQ7Qm6QfTT51Jj1T3XZf80jrcivY0
4z9OqmXxmhcSyjr63COKcKeDpmyjmZHkrXOh6SZKxxgBxHStbaSu2wJXjRDYKL1DdYS8GVk7S95Y
a0aJIFiLwk5h9u3/SKDjTrqu2u2EepB9qDbZgXxB/f0Ug9WHGe2mmzhJubw2dtP94gpN2izCmdQh
SKZFU//2Nys2rgUUXi0tFRrvQseSpP8HuopPhNN5KR+fWXw4utiU4MwcTV9vhyMdTySzggfVOGcn
8J/R5kJwFnapAib4yKa883ZLc6j7gOKATDhkab/uKWrCTkabGzbmlmZcXrIR2JRTrg+fakV0Hg0R
aDHsFc6IvVqMdQGJsnRKhSzhZUVM+RXLxa2BT2l56+Ev4QV+0cD1JpSNwyEBr5RkKmXhSRENbWzN
dUu0JFMiDwJWESikVucIzuAHTSDWJy1nVRlK8EWhabpx8Gg31BB2fmOHivZTqDcTlRLg3ecBPVFo
WNtqpf/nzltl3r8wxUD5AYaKxvKw2h2yAyQ+XjNnpo5r7RsL80eIDGao/uLd90i+RExSdgsyw+Ym
YU9OLLzRUgigMOsyjK28+ZY7OPK9pnY4L4r9c6He49W3SqlvOsVfMw5IvHO8RZgx/1TtdzvhqQbi
x8XNQZKeAy4c0YE3Uo/nwwm96Al0qJ6ExnE2hLhlGXJdlWY25y/ikc2L5Ja22LN2plEed1JoRAif
kfjAm4s/oShq7dbCiVxSL277qUdXpg89Ws5xNWxd2zW3d45uvhg3oCNMkBDetezkyybwnj4tSqR+
4G5QQhwrnIrXyb+G0lDo+J+gcApLHsWnzsonM4W1zoP34Hqe9zgeFrW9KJu6nysiBDcn+uMLAgWj
aCv7sHk9aOHnpVpelhLBJWa9D1MX2MICsg1MAVAi1sE/nBgALp2eGuWEHtuRcigoTAqs1a+j4XLs
MN8OnVV27xvOCSm/tNaPzGI+GG23Vkd4lZlEFFjIf6D2roEJTravIoPEMqYU9/qHDdmWdUJmyKFp
Hid/5Sd2hcFCdpuVc0TciFoW53j/xGqivcDaG8TVIFyKdrUJzNJWKOJBOMEcONCTEDkawj28ws4I
stCYvrdX6lVTE3eQKVLRbGbMDK//TV2OQgQEEbhzzjBHDuPv/BKb87qbjirs5I3DBfHk8mtWE+V7
xXg8IlkLmfNUI5N8MqvgZmZtHlzAR+gg2dkasTQSLyR7DL4zYWt1om/ZEc/NRGrJaNIexSvtgmNw
hkDZNs/r4pr/IiWxhjhT/qMASwjWCEIftDgxr/DCudZG56Uq3JDCf5/iA02tK8lLP3gp0wsRWtaR
EA2isQqU1h6074YkPb8LZRIioA1V8YrZ+I/v59L08je+U8QdEyoN366/dw1tqSKLfkSajUaph7FD
2/3sGL7/CPK3DhbjXzRUtyA5s/jZr2tLAstfe+WAcHbJB1UxKpKAeVyjyKSyxrPqz5XGTKtWrwRf
c0LmRVuNUthwB9yf/z3V73QPgnxADjT7NfAiLtMh+SpEx0doI+G0b/b6lt8zfP1NJ8aDVQgT4q3f
a+TIYBNzeibGxGxacMff7xtXKdOYtGL/4gSDaWO5qnJJHHCd1Uasx9wnAfpPlYJpHM5LjQ6uEN6k
Poay+dUlnOop2nZHjHbmA+YU93PSQEugztCmRQ5DOxNiYDtnnmEPYC2+IgI0DOz/cfuZIDhO52DX
AXbzFxq2Ly3EAwtIJYWk6BjJf/4ujS9cAPA4xVmMiT4jBwhIJLzwrJI4jKUhUbkkC+zhLHuPRUgQ
ehDhBL6xsAtZhPV2dyC8IWUkmsgyJi0V7yoX+aEAouO7UCztE3O46S6oOuhjdR0PAOAstzWOLU0S
f1gbSNcH6qtVBFdyeZSYKgD6R7Ue96QlI0VH+hIOMuWBdysJrPSHPJeCkUE/qUOlNveiSyOpfySF
SI7ipvy7oJxxfrvvE+bcO9x2qYeLxb5E7aRRra2sU5cLcy1UsGV0YqlfddsbNrbOD9GCfpoF0IiP
ZAGKrv1QVTSYoCLIRxcCAld+fErbdYKclkTWFmZZ3HskjGfc/Z5c7wxkAtSLgks3hhgL6zO3h8Yb
m6SnwxfLfxb0U8Ib23NQ8ilGrP0bl0a4Ls2g5x9I6Aew/MYUCOYUjYDYTC2hBqsXB9ZcazG/qXMn
2PWiJJgP8pmwE3OfdW4Ko6Jr4GIExv9t8bRSM/asYqHEKifUonCMjvX2n3Y0m1WJLru4ln/Xg/BO
nJ93Mbs4xATG/qeDxGXiTPBxPEc5WRtsyHaaBhFtJ46/dbg8R1IDQPDFGKINsUlwPceIl8PiYFeY
rajhtT+A8iOwc495q+IG32KiCY+x8zh4qbzfHSXHms3O1eRZzKfDrWdVDPxEXUt3qGGzieZ+nBPr
Yl9bpkVXeetOIzQo7twBbhmv4q5dIcIFqCCHxccb+Qf1PuX3qhMYeSuBeMIza4P+l5MNIT+nKcbt
mXIQH1/L722cvlhWxKFwUK3UxbTO0PjZ3u12bnEgiHuMflI9bD8tM86uyVwidR0PXd934v6eOmay
Dd5EG4PuHfjRdpHC9oB7aObvV1u+C40yYY3/25BOK7dy6y95vsaXeFhmfk5V0d5LEfXqdkFY2fgQ
yD9qApBNMldezZnBPgqL8yb93qXJwcEdcQ0AlDbzP6/CBRsMA11WxC83jhQFCvgcVBFJvrdnw9cC
Tm4a2PajyKXUKqe/PkNf2t5cpX/J6f+gDW85OAPgz641M8N0kAwzzMelMz/g90Y7yxESlxrYUyQo
1Fa7D5CkpHCPg/QH+/LKY+sVUu4l55O9OOF4o73KoiFeyqrTPhSGl+icSf+yD0Dj1RWk4kzab5dT
MiTvqeQFtSDvwIVKvMywVgRruTo9OWZcgsePiPVBzq1fzMNb1Ur/MWu4zhpwbkmqyUa8dtOlGPgE
9KHayivIEdf+FlZXTfi21OjaM7WqzpUZkiT1ahZQyKELavTWW1xOmc6ZHlNvb6DOzX6UCpP6zhnn
FI9XtmVpNJYUWjdUWQJH7fxmGf8AP39QV01mtm9VyqXnQknaG8oFtMXaJQQiX+ridzeUU+GzRG81
tXmmnpI5q3AGJXAj1A4GNsdBsqeYOPcsMjhfM13UwtKKnyUWLMS/Gj0NawK8w16UOokMiuofTQ6L
us92mQpb7ErBej0jAqeHwdnt1Etmp8LdUrSHCyhruDkomEiTICIkDSl58gl+0rWhASf+/mwFs4Nv
oV7rjy3ZVMSOLuWPwzcAwkTKOKelt7hZ6i4pqkNfjKJ3kptRQfHcC5R0yPu6Lb2C/B2Dk2WMf5Th
FNEcaLHAmHX4wBdG0L/3V77D6kj4XNDbH7M9YO0Bda4U6Nx56Y9CIeKpslX3T9OlDyK+yag1iuJL
r8Xcve1OBRzr9U6btr6Iaawsv7mECL662lLF8ew2zr1jyxFI0GvfVNA+TgADmUPHmlghDt/5kGJg
mRfexLDQMQjzY68frLRVW6vL8wd40YKEM3eoQg8qi7fLEWYj+iZjhcYz/JxiUiws/4f12tgge0he
noH9JpnfPQ2uaNs4RJaFs0uPb1CDUBmtZbqx1rY3g31pO2gV4lGYGf3DOxC/sNQee7oA7q9/Jd52
gUgPRMIgA6MkAVYwLdJqvY060EVxTP/hAFdybItwNO0S8CYaQ9eEJEE6kob9OuMljZvEkV7gqeI9
4nFAqVYwvL5VofI5XG+MpFIUilYrEgW7RMxuBUPupkFbVa4zmGppBDMlrYuVe5eN3b0c34k2M55A
OFqyRVbOIJlRbSGG3cKgNyKmW768gK6IB9CJ0RyITMBo9bQjZdE9j9ZbFd1qYKJCZ6XAhUwCLq6F
IE6Vop+zawlm8n5VzTJps92KvYdM6uYKmq88m/WZ6RY9AN2aUD4KOy0qxlrWH0+qEf/WMYtNMJ59
tPaGWmts/5ivcfJJ0dT/Ohh6w9+4po8wGz+XEARYVycSOno+sFHBDcaxV+F9V26HZyUWa9pe6uAp
8DSP9UmD1FwazLoSNghM86xQ/qUh9KKmClQ0pbtjrzc+Ik8mGAlJMfRXoItCISLsUjpswBWZiKLm
EASVltlp3fTjRisS1W/xvVoBuZw5sMZhEFCd3zhay08CZMPGUtWJMFERA9Tc2RcnMJbvfsve5JNU
e33doNYctbOFs5SApzor44J0LyBqxP+MRo89qaSqHzicdjXZwklVsYiR8YXw7K+x61xznX71QR9p
sxRYXgjPDhWb0HA2AWtFaboYUPLjAC7jTlzLNW5toEgvOiaj2Mo5N+rPv2EuXe3VZV4NUqps1Qbu
CttnCVPYSZCQ/d31x5or5rUJuzaLpP3F6GPiK492XBfu4iHSCiZxWeAr4OCPGyIIfVGcCN5MEGrI
2LZHkyjydDJCFvAIDiq9iU+R3CgTHMxMI7ZmlwOPwB/hrdTaWO0N3BRc57gV7Gc6rbOPasHMBefq
SCMRCKTLbmwpw2KMUyEppSyMSJTxpr+w1PK81HSuxKA+5YckH0KEY8pz5EEu92x135aZUh4ZVRkv
QpFbnoSQPDvtbMqeor3r4/pcbz40imn8V9aIZbq9oZ/bWARWq2DJCZma9clXc+i2+bRB+G3SlZ2P
E/TFctt+2445BTyOdhWkW8R/KHXhdv7Gv6KuEDD9B1CbJ4WHevrW87uSgnxvHzMXbJo67228lppT
jJoeO0qgdkXJc4wduLUVyAm8hAliIhzlA0cqoV3ltpOsZxATkKNTbDFPF4TvcUkQ/i5yRt744zXL
AeIq5TM/k0In0mf8XBrJW3J55H2md6zUdfFco6aY4xxVAHyPSGt7kDRPCbsDLdpk4NjdfQOZLtiu
8ack/cvOnTCigwYT78swUTDDvMmh7QBDpfYdT0clTzMGXR5/1rPGzak6csavH5yUNYIjLpR3Rwi3
rckeTDZni4QavowH7u3eymOTggrgKl2S6K1/uy63soeM1T7bdGof1BTPhEyZ/9JxIGbV5eJz3Yn5
pwuC0SL8asiXF9qeuuIaJHRAD+VebSrwe3/EmNQDapuUy4AZHwqX08SkG8we2xftoHmiN2ukwf45
e+te2WdOYl+lfbxbLL1vVPhIb+dBR4U2pE4wtWdvxopNyR2cMysd9zGeobXb+ff0FR3oMEbD8zAQ
lu3kKdY2Fwq3o5giNIFaPHmWnXmWsQev/0cxkc82gh3b1B+4iK+GBD8PJ69/KTRAhF+pM2D/SODJ
5wnuMzxgqxiI7LZLk9j1mHgth6PYRecKVJfLxFmqBCp9eWVm6EAR2MVDuh1AH9/NR/bG95gniNX/
Ru+lKA1kQT2VgLMMFaeAssMM86k+55IQtG/TJvhdiIoKL27rSuGrpUafWdDFAJoUuN419X4gpODZ
1gL0XQjwiwDSi/jdUnIvGP2DIRy0+KWZQ/jddEUD8ncxbptIxgIQNtar/878bl2YCa7fBuyUwjj1
biyvpnQAPpow6bzXF5muSWh81l5ZE5P3xplAz6XGwGP9YrxlDW3tfNyChg3A0xZydwNnzTRxvnsj
bHi/4zHGPbex/qa0Ri7ZnXepjtzBnepot9FXwcPnciXPCTj0CBzKOhoOYhdKQKCl8bzFkD4By6Zz
ax9o7RNDuNS144c75yISKcnQZ8Cii621Sd20EYMvKunb5A9gx8qkJIl/lv22+FOyhtJheflKbSsD
trBeWavckBEgGVgufTQYGC/Cki6yyUkMcMb8meLonVNqhiLMOf30YQBTU65NxNoK5L+M1dwdEfNS
V6JhMxg4+C42loYAt+TzE3M9Kbnn9rMm3ykH4uUGjA0QrpLLOLr17RsqvtFpkZpmjMoBCua1BLSb
JRqNs5yKSuYIUvOqFxEAMdamj87KPZpD8tmZuwyps+gQuiWA/kfy5oFxBKP7ZsQeZIcdip7j3mO3
F6x8pqapVDwjsKh1ZDIXbEVqpCpkhx51nFdWbrfGEFsFwRvYJXnl2EaIIY1hnzZzz3WoFxoB2oIj
2q2LIMRRJ7+UxB+PhpeYHozxOkNYnAccwnqXNS1euVoMBncF2SqIuoCDifa/TKZuwnryejlYlj55
Uvsn5BifKjUFdAVYJhAvFb14/B4oB8dm4lPohspAalVqmFr4jrQ4y012gffyZYakr/yOq8PlHuCg
oDKv6kHY25U/PEP7gk3L7O3PmEZfyfi/+c0/+kmsg5Z/uarJvW5UKj/q9LK3O0+66H1WqnSnDPZ6
aEwa3+UFEkkbnZcMAISdqF1AjK4hpXCoCCdqth3uf3+Q6ws/JenNHnYO83LTHOvuaILT9vHRu6IB
Te8l3+WNMnzteMOeZSGfPfEOR4GkZWF7CAKiKRSfrbpfM+4hu2zqIch3wbTV053aFWKvklODI6r1
V7SgNtSIWVbgWPUOqE6nwhPmL/s8neLx4CZByYtFJQ5ZL9U5E5GVpi10hOPmcoX84Xe8jhifTfAL
fVXVxIZYCQmhGY0+FDFrbCOOPZ0AUmBs64qrPQGyg9nxCMZUlpvSbI96xMLN/wnuPgEBj3L5KIsd
RzI5fCKinyveEjeAt9n1C02YPR4dHuGWNTe24q+dP+IRm+/KdG8u/MRCsVD+tkPwTCAUheetk+23
zBM2Sk3E3ecl15DXw9G5lXRlsAtkt7HUhGGaaKTayuJZ77DznsdNTl4oc14a3oJm/dU78quhDFK3
OBGJCOsg8h6VszDe4xWD/assuXt1Zn0RFqI1YvN/qcXw9cF8arPIpNnEFdKyu/3bWUN5aAwhm3j4
EshXQy6NQF8rEwy+AFBeYHQcmOl1bTp7WX4EXDuBynBr6zkyxrRyw2wKx3tfimOEKv7hGXvrXbvk
0bNsCmqSY2GEQhftpuWpLf/kp+bp9XbMZLbaDxirAlx6hdXwdG7qWyLUzbhafRk1sMy5U1mRUzs1
MfHVGyLrsM0ZJ05RWORvSmw6x6J44Q35MNJ8U+LNGdsf+pxfn/VOHR/EjinkvJVsyQ4DHeXI9OyU
Ki3f4lVidF4E1WofNizaMnhL0kfCybRYtdOHqiTPQSIPcoZ7vlNMb9X5ZcgEOTxkKlPdZ5OJ5NAP
T9P0zi/Oe8wTcHZwTo1zxAcl/Db65GlonKXG5AjfvQtfKJurPmcHSmz1RWJLN9FXr1zbxo8WigTV
sR743TNyH2Xn8ZIPEtnmghlgtugbG0hEaSLZKkvwv3HXbvuo0M7alfwVwWZLp91up9ILCkeCIBhq
5PIdIYB47EyQ3XFSiFXgDpZQx52eYfgdy2JTJhArTM7ibJoF0R46HC7JZ+K2jYAMEKutaVZifWVn
lyUQoXtA3e5WXQBee78aaVZggzM0JtvkF/jIj5W/58+6yCnVrKPUtOmlgzGS7xe+twnwKd88soW7
h/AZL9Q4637ify5Twpadzkv/Q4HeWBlAx5zmzCvqg1wbwCCEyrLnS1HvyMv0ps8RrM+78aSMIMQy
QoQ/lWrKyTzcPUzxJO5N0Pwd2bIVEOqxCLHNwQvDB05z6yF9pFJC5b6bXIyOAIoxLhS+xgp6jRk5
GiSdo9hK7b0gY9iaOJAth6WdTdNsl1KTsHmftlYo66g5Udxd+0lfNJeBIrpLdrvnit+AhqzW2Kgl
vS96l8Pho+NL6x7PKP3/FX7NvijnZI69z17ZhwEUD3fpveilNUt7iV415SFhxw40xQZG1Rp1MHia
wuhO1yBZaRQ+sb+39NTv+9OMocDraqHj19yjAp//TuKrtaCzvEUfzDEzARNu/BX1eJcwjNi83+ro
OYF1QnsCh3q7f8mwiQfdjb8bxfm1FWl3lagu/dGkZFReixjMHZUZODHkG+R/CMs5ezq+0nopGZ1Q
B9X+Wm5eKHXPhB2HcgtMHZJ+iZwLykerXPGQX+fHkezc9AdZ3grnHH9XKBUzfcZXhhcRTvlrc5wP
jDw9pqacRpgBkv0e+BEVl6wGuxOW/p5vwBMQQ5F14AAJl11BpLnb2KO5uuRDmj/fJY+wH43U3WPn
F86boNSVWsfggw+yhfj3+njnr8mzn+6Yf86nWunGhuynXqu/SpQ/SmJ0zEmTmH2nf3jx8Jq7xqMu
xIGOzNcN5hGBFfMBLZfGZ5EnZCuOwhvsf30tlzPqVh+862tHDR4n0mgLFK7BKF5dyGEB3oxNrhZ1
/RiovdiEgoHdEtA/uenF+ecNJZT+CzLwLhfz2OWv0Avnxt6D/Sgw02Nl9FDZqRx4z5Qme7gUmEDF
Hkxwh+b8XFq0EoTB3wDeLsPGUiUPI2vXwQKv+412TGHjSTHCwGwPT0Oaw1OqW/TK1vYsj5n1m7tF
Sd0M2basvJR7qZh6QcivEG0S/1c2wlXlPzTeOKql6Yidw28fzTkKvb+P4RlMwTjjdUAAwNtXjFH2
s4rhtwgCO6WyhbEk87raIjsb+T9G4gt3bdN/5lkt+44I9Ukq3DHk6i7xXvxVr+1s+Uctu74NDcgF
1jjbipFFLyAR6Cy3gbuf0yXHZuBTBggimQgXK3FstvuG3dGcSoyYNKn+soKKouWNYFhSLcHOeagm
exgW4+KrtJoSDyX+FufocoDtN0sXkOhmz1M6o2UZpXFUZ9nA0uKZUh6DRr0+ggKEJ+jgmIQ+PHMH
gdl5wGOAnUi0WKbyUPChoFgU135JDRpemQm9GeG3IvvZPNiNLyVHNO8yTWIqjm6zt/Aikexv6Aic
8e88LnfeEhW1Eu7EviYDm6wXatsI03jUsPfYzLCC0lFMEy3B/uio+f2rfnzy6+gML21IwtQZrqKu
GENX+glYhiZ0k9qI270JAvhQ/MQPFoWFr6BnYonYhaEwk4BAtMkCiUaCFuLwCw8xfYjvLP6kO+1P
lo+NCjqR9JhKRjij1TJCjAWx+7TybSXEJehsVJM0DiUbcTVVhcNJyDSqJtsSTCQSbiyL3Ev//zng
hQaO7ZAJN0n4EjF8f+A7fE76F4SfygLpM3/LB4kEJyNjGQ1COKxY3PBN0V9z8wZH2wE9pykCdiie
Q521lPMdew88CPHOZ61CoSYv4mfpPyuQB25w9ZGSSpRxlQMZiMmetwyP07rCgHfXyjVZAds3nRtj
ujR6yRnsayz6fAyZL/snKVNip6nwwEmn7l1/jQgEo4215EwWmu9DbzfTQur8H35ghr/dJ4WyoepO
xCeyrj8QEPNXE8Eh+VPrR58ntRHq4/n+rWVNN2VXv8nJ6FrW/5p+ElgcVqkk4aXybP2Pwc73VW5B
gjALSmArPyYKt24bGkhchlJciE88fQKKQoHGcqgVSnB+3b9btiZ82+yzma/hXf6Rw9Le3jWQpMQ6
pWTMSSYuCJE50gOa31tYBhXnkw0C12dBHrj240l0pzTXsq8xMXMDRB4LhLaBgFNHN4DGm48uQjW7
WzTP6txuPW/J61HJL70MANZxN4UXJP+dCwwrtNAPikMzv+46vhTz5m3HwO9UzppnUqKZivc+EhRI
hC9NprUIOPVRFhsaqiz0Go/03EUz7ldorRNm3X0YQUCoDFv8X9EV+ttmHSLnc2NR0iN1X7U60k1c
X7o2uSH8K+C8HgA2Pd8P/elsb8+nY9sDxzAl1c/b2PAcJ1ziiBTJVzZILCDR1Cf3xVsUDdvqMOkP
tNb5O85fQbRdS8POfIepfBjLsfskA69XQtEYWtVie3OrERwlh/OsMmGsG3lZI5X/7hr0hNwXri7g
6Umc0/2iiBSaIUl2zLIV+tMz3GDXhZjL7+nVplWTtkA/ROxSShi/nIy758N77P5iYLe/tUlHrsEL
epI7wyOUKcnXWWKdZAGiLNCuobDxUBHaJGRyVDta5Y8/cikKwNT66i48p+85PjMziS4svxIZ2yda
YLdHW88vmmLTqfL2+f8/VGYf9mMfaeaDVVuKRVQ2okw/1GWnyeMz082nttGaGv7ldmP1+JoJCuaf
EIqfy3+F5PmYGb8oGEi4VRI8rk2Ri3lkPnU5pBoU+h6c0ke9POZOVI4hf1fzqOZXgG9dpdiWo5XX
8ZtneRn8dJXCjYI6ra4HVp5XTHICYVcBQ7yiFkRVQXFqdYQK64ujPEshuw6gF8b29zGKBeH2klE6
4gIoCpBvf0in8tS9k7zHTXXMM7uPpQEvwUvr9Ajt3U+yn8TeaJ06RgU6MX6RpjV+GrMcNhPbJvfM
fF65DVwDxIvCdd/4rnpJ0ZEsmBZdwrvBRAHWLlCXoyBMFva3Rh6yEdTAOHIWKOO13Xesv0V8M8IS
Fi4wc9Fj7PyVfxh3LduMK82guQOdBQgw3hRV4OtbVgOhaYPnAqCiPf7SN2WQxT1WSxQ+ovvubzAb
6dAuWNGvxNPF4BK7q3RrJM0y4AIQn0JEW+S7MNrVjCCOxPr2Xb7PnsywbC2Z4TSs9prg0jNtNYR5
C8c587qjaO/lf/FVWLS+CBgBu3ueMRNx7DbbdJmc6c0A/pkecMsn528sfbXkJz1vY200S3hltPfV
j2sexn24ClzZhdb+9m2kJVjRAv6iXDkOXtzF8ZV5Fn8bdqalq5IKIjV+hxxZ5Q7jUy7XUiNYxdrA
8LbpaB4pqSx5I5nROcxkRCCp5mvJxIk9rpXEbbh/LrA8g8oYEWEIrpKP0qjcOcLmFtq4TY9EeIU/
0cWelNhL2KKD9dojueHxqjZLXN0bcG8HGEIeqHoUoiwl4UGuSfy69rhlkm5TJe6L34AHtV9Gr3sS
wQSO2osprsZObqwuFtG5OKfgBLxKv04VhaI8E9wKj93cPUAQSLti2HcsaRpsLCmuTqi+R/gGakTs
UQPU2wpMwJRJrMlUeixMgs0EQp0yCY2wHknAdzXG/sZ7SqdJCMLlLdrwAConolM0guUFbgViYpM1
hFU6IdeZfdXs31Ub9pEVjMLDbMhcZy7XTWtYkRV9lCCTgUKus0El0WXOnppy7Q7jY/YHoqTtHght
TxO0WhIuV/RBR6h6LN/X37JDOqZ3ohFc7MtsKbDiXx1o1LdWpzs3ADjgXOj6x610189loQs3/j9v
5ANaFXSj9kmpffNb/yKLqqDAUuPRLXW0YZ3qpYpq6AeY0I1z4fcaNhyjHR0jA83zWP3yGPqN0kJH
QyITWDfO6/d40tG9NxCCcXzpUZnU+CIeiFmwOK28K9r3+mQlRGHO9N8zl0xNgAb18lvhrkyEKiCB
QFH9oFsmIpANb6vwisUoNeZHGy4gIyeWMxYU2ZHEEamHTy3x86kwwqUZgQpKDDxZaqfNns3zFzpo
n/8x8pFnYpW8gLn64Nom1RTSbiRguwNqZNeyEPkcOIkgRMlgiZHzDbMe7FrAhhbVUZd3OR5jqkaJ
X8muf1VYMAJEOPZF3I316WnviPYoVaVKldI53Keir4KzF1y+hGQ/j6KfjREYcJe71NRulWg9mfPM
PiI+7l5KGkmH7FvO1j+Nex4U9oIVWVKf4cclRlTKwd0g6EiPWSZwizc+PO24Xy77Bm9zNWj9RLCq
lkVR/jN+QCxqD7S8YDYE+IP7Kyrnjox9bIHfFxgY0IsNoKaSTj6+fFwACdVRKQvKCgMJed1CsY2G
8aemhdNA+2tqjpiBfz5KhuAM/vENUZliIYRjFticwktfMKn4Wl0t1XUv71BHJO8wWXDh7Ub3jJRt
OiVk266lGD4zEVXMLQ1y+GtfypgoOOk9Y3quKKmkYxq32TssU3wWoPXXZQ9rLXZ2Na1D/5Ttpt/X
x/MSDOiMmtXUgBz5evaWlfLBTdCclekdtR6XVAr+N9ySAeU0IP07dzP5o5P62ww7TpBqqqmW3DQP
yE53g4d5cHpYpQyGoUsHHF7ZVJ2/Qixd3Ql7GrRlFHvwVVHXXQyhpPJ95L752Wtu2eZByh+FZsrI
QmPbuV7ImZZrxcimNXv2yPqazBKhcplBTgdxh4cQrMuh7n8QzsM8QGuUEioIq9/2cd/zohroYvNr
wYc6nlz1qhWOZdnb2UXaYuPVdiGapQfs6z1mANwGtYSQzmsPNBEkmXz13JaIKFDNq/1YHL7XisyY
3t4wUsbQ4BsxgDYKjRrd0A8lP2O6QJvS9TlK3K7Nsg81lKZu2Eud0lrM/iMTb88faDjXsLEA8f2/
1FFYdXkPgX07U98oBxWB6shBCyq1SCzVEnckCYZ6Yq8CY95PpieNv9bM+BXs9BkqWserUwEUSko7
M5nSFdllTis2IcTIO2msHJXgnSBFSDUUUq7EqE1tXls1KheucMNg3cgLcohk1PHsr2KdgaY/ibT1
Z7TBlXJ6uR75ynWf495V9ZzhGQRl/zR2cBY6v4ZNOORqQXrgXCoJ9MYhJFs+12KpCa+ltJbGRplW
zc3x0AZgOqhxTysraljjBK/ThdUpZRnA3JWczKbFlJuhcfRlCtmvxFT2uKkoMOT1MG+4DG7YBNfA
WJUC+rW2fnNw4hhsyPrBKNrz2MpUJ1e2KAx2ioTLGJ8+bW7m09jS1bL+LwXl3FDiKszRcQhNLdxO
7MMQGwzrng1jTJvQiNficiysU/0LeFcDKhNzx2dwyyqdSq/j+cS7wtntoErmQVrbLnAZaBJmyyL+
auTJbpfxsceM+ZU71flCCPLq2Qc1l99++cAyDlIklQGMsMoSLBep0sW1rn/KvweHyYkPHpJLHyeL
tDcg3CBC/g5fDncE8OMBFQlKXFYc5WuAqNdqaF9fq8hlWoc9vms9zKUf3TIvdHnnqAtxNm9phIU/
ZjebcJNXajY4RtOOiyxIDJ6IXiTjTLDabJBdcInC+cQM834nf8FnhxAperEY7dAG2n8fgzklKtO6
CxkjbyLmnuKMVhOqQOeMS9sOJnc+i2E2usC8M72XkWcdrmA2+MGQUaFu77Hy6OLR1eujokojBQ6Q
amhWH3FcdHC84sOYGuyxpaP/9GmToPS/NIOGkB4rBy164TFrtXSCFGEmPlCrEKn+U8CSmwduuG8R
WbJXhDyuml2sWsE6KAf5O3Mv3P6/6zP67LoJDQK0oL692e1SALBSV3uVqw8XykeomxB74/zv0VYD
X9XyqM1g1xrGoIoDEUlwq8PFyBpFPN3v+my+pmmiqQ/bmD4M6SrAvBO3eDefEQZBqRqFS8dR1OVK
oNkGxDbpv/ZE8v6aNP3RLoCBXZ67dOv05cs593YaB+h7x6KLJZKcu6kbwYMjBLhGHH/OMFRTTwgQ
PIiNAHwmkQvMzP99M2YSOvD8DP1JmNI0HWsZVZR4AIm78WgQ4aXyVCX/4c0g31MtYW6AvTZOtotu
F9CxN24zP9YtwLxTVBhUxQT4yHG0L78uInlWhyCtm+hqvf6CSq+V8M0vM+cphVgX3CJBgnbtjfVg
sAkNzBg49ed3xuXpuJIDpMQGb46GnLKBVVYXGqJFWh6TpRUEr1rzAfXVNjWI5JJN3d3fBSNSMGml
ERz84u0isAAJmBFNT/LFKgo+dTeZyzwWLmY332Qos2T/ymtsbyIJlU7U9EtUSNHaidha3Q9d2zlt
TUNELJNGNjcnc5yPZam/AgmfZdb2zVFLKuxkyrxuRnU+clGJXtj8AnWmWNiHmJyXZ64Q8dmT3EYZ
z/cAKgIOuKYtJpuz1IfnuoI5MbT9H4ht0BoEiw3JxAtucM/jfQH6xo6cXUFgvrhzVq+b0SMSDnVo
D+nbZJ27bqYcNi0E3iK0PUZQ04LlMw7aS8BMc2B6ClvowfpAbqZji6L49AA18YV5mUaVkcPLQJgU
hMl6gceFa8KGCKYynhYRmFSOv/4khy9todj/gpAPCHzIWxk/dF6ZJFnepIr1zamXNNXNO72XfSHZ
3MLJ0iDDdsxvgONQT9Vo8pY0rkUtLucKMOrG63Fsnb7PRVQVSL0J5u2Z7XQ2xZSza+uQimFq1BW2
/hbLCD1KPyhZgNZXItA7qD1XWA9qrYzbRWTMeP5EhCY21CE5bk4M7Kky/eZAuaomp4vGeZF0Svzt
SL9be8x7zuozgrUYvggvlanViNXjHAtM4cs7B8lA2Eq154mTyz190dyOibrKr6VQUcwRBZ83UVnt
CNw9P6ZZ9r8smwNxTLdaLVyvTkUPgJFibV9PvB5ZTYlVll5IRSPpsN47UGVwZeWSN5y6irNFdzJA
23h2Zcm4puvfbCNx3MXvoWEKqL9iKSgbz3cOE5hjnSIYopNgI6LAbV5d5ScygPPzR3YdJwYwQ06J
GwlZgQ0YIY5kUZrBQOqTs58dkt2pukc8S8zyi6iCEFldMW61K9W0LkJxBfEr1ZW7sIWEeChAW1Bl
iU0WZfuj11G4w+pgq05IfzAqKVq67oF5dQg1pYAhn7xDg4ZUbLWIA3nApaWwtiNyM9LAWVpqzRu3
f/dchZU3CiDYb60EV9mgkpa2QoetxxY2CaKH10blbgpamL4jvilSwU3HVhSkO66MtKxmkUqg6jf8
stf32dH47HPAZ98s7WYpzvIlOLeqkD3IZfPv/cKCqmJ5AB7tlZ4/pwCO5qG6VKZOA5STM5a1w0w8
nUvUDWuKbUwT9s8FwBWJj1CsefLyliIoLO/AioswVwSnxxnkT4j7a5NLh5TRxmxWtWjUeliCCygJ
KlZONJfH6XJkI3TE7fz11MGdp/VID+yHWAZF28D6KyJFyy9533HX0Q40/4LVGB+F1uh+AdWrTs7w
a15PPhJFHDixJ98sUpZ747EDEMHSN4fgxcJAyDzM+eXSeGT+37A/YDK3hkuVbqxQqRlEdd39uUBe
9umMBv5kG/EJALSQC5Y+I/VjpVWmEJ1LGuERZ33mTELJxuE6zgqMgt9n5kYWJwJuVgwqCwTVDmbH
5AqiiKsr/vGJF7xvthLeQEfe/LU6b36E2PHbCuuFCN025vc7Xn/1FHlcXnsIMtVIbHPCVnsvZgsH
FZePfriLUoMNIIdMqCkp0CAMz6WleBlu6182OkuAKRhnsyCpl7I8ha6PhWCAj+exYTrAJnlzy2nt
25NliLjN7tkaq5wWw8jID1sgyiLD0fJ+5aotMSYcF0RgF5kq2iQgLvbH4MSQtVQceHo02yFsRGAh
ND8Eul9TVQaACwXBG43evrL5ZLx252lBoRF7B8v158PuHqR3FLbySezpEKNYAzdAAl+P8fUexyHC
LCcz74CD1IKZ3ywuqReFOEYJrZmFUxf8oSx04vDXXLAgsmO0TfGWPbrLaUp0as4OCfzvdpaOM84L
Qrn8hVqHWDSD2RNVVjCeojm+RHeFQpCWbSsPdp6t+IRpL8VGkyzoTQA58qTIvgzlMd47trk7U4FR
UarRysnPNkCFOQWvD0tZ7fWYb0OicCT8P+Tym4PSwud7OhEqZZUj831qdhgpoxsIof5Y+Ujral0y
t7DpuS6ibFwanRiyrwZ5dFp2e3KK2HBSxy8WPPac5uCnVW0FdoXEUmHXQjGCDydUW/KvAjt/zO4u
273Ip1W/oame8UeSNQwo9hX7FakuTCV3dghpQKEaKOsk5KFQGlnRWMnvFercRceXBZJiWvTVF9jI
HyPg5lpfsHFHaxyIe1m8OEI7xg6r43ncapBroXm3KmFCeWC2RMQuACpXiZQQQLgyGrgmHAlFGn+L
JWzC1c/aI5ctGwzRSzgjQ89t1FduBmjX40kmgMxnkwIJlK32nlOP55Gy+8jSFg5yo2b0SCj1Rhix
uNVUfqGu4jZDPiY4hWjpAIZpnipsxbPjEe27aqgqOKvDZL+sGaCLSqqw6FyHbyBghiov3FsywKCH
NK6HN5nL+qd+8DTWd5OvSy1fDlf9U57M41dMFsrPkf+7PegZ3BgJL5e6x1HLwiGyR2Nl6ZeJHH9h
cMvU1Uv1hEbFYrkqgM5sWbqeaOUorG7kHDkHXdVwU9czKJlAfgokkG+majsU0QI8yftNsru1npK3
IZRpBgrqmdwnsHCDz8GnJHxDfyfwqD3oLxqgK+GaA9VnOIqW+peYCWBLNzKlyFw6vS1VZEbl/BLy
r+HLQb/pJ6tbQ9/RCDUH3eAM0ZC61WMF0WlLtB6IGJz/bTgwYKq+QGSO9tX0bu5JFLZnSqp4Pxxr
FFp9gZ9Uw+nXulF+ADH4hgWUP1WeA0rWJtp2h8i5fT7PwwO/DC0/xbp3MpyjxnOlNBpZFzyBEbwy
Ggd217t8usQVzmbZWMP7R3qDoL4+I8XgkElCsad5RlSiXfte1MQjrGd4cbfGCpmXt7CnwvNVfj5u
ecNmczcobGzzx35GJ7UWPI2xHaT4xoj5Dm7N+w4xhV+OsLBZwuvGBOaBYPCa5t6LoFde/vSZjyVZ
WjaMsMjuJTtzWA1pQYj2lOZbhqHw4cjsolXupSvVPBtzjgIKFrif4E0P9nqS/wcQpL4c4svo+OvK
2Mrixk3OxLUZZVyR1NjJ91pmYP2Wys2yn6HqtBFyLd3V4ZR8qQijm59/dfo+hqXdk6TbyzHsu2w7
jtQ+sXcc7h7HPVem9VzW2SBZupOg9NRsjCuUfQ9+ORp57WtVf0WG0L5BeiCu4jDF5kC5D/y7FD7O
WIZ9da8xknhsx1XDGIW+lBCLndQtji26PGjmiuG1ZPDz544OntIpWrGXau0ziq6upzBc3BJxPQf6
IKkyN3nmRl3xaxnuY0QLRD3N7ALbwxX2g7J/IlOAo5UCcGk8+dKUB/ibxLtxFHH11enxbcCpZEsE
Jmod5GLyh7FBL+2Uu5PqVAXYfNiU25tOGaHxal4O0OEkdS/7YmguYqLdUtv2TpmMSDmRT5JuwpHr
b4Ehx/xAShx9BgFU4LJmJLbkJsxDSW9Hf3jleNiW8nobOh6gPzmHVqc1n8tTAAP6m0Uoa6zDSTF8
RaBr0hhGn5RaeqX4FwyZcwE+iLZ2aIRVvQMGubnGU9N0Ll/NPCCg7ztr1AlfX7dFUTDfNYtr8W7S
tsWlD68IEqx7g07VKFj6ylFyNOh/RWNlz8e1oEyku0GNG850my0z8wij06oHRQq2JCewh2w/7LzY
eoQGPD3tfPUjK7oR/liIcGARdCU4rAI7PU/9flubjJn+feLHjxcFkfbKbsWVJa8pZhiYl+pmZZI0
tyQsOgYTjz5AVyAo7rtYcMOZibbaq2J5QMWYygeTZtWlp7j6g34PrSKgOnSSxOPd3SLcBLm1LvxE
WrjUgzbA3yato1YB+LLuVNkXCupsl8i3EeorYVjv9FH5Xasce6cSJHMN8iGwhcnPCaepW+E9BJ9a
GO6IoqXcaKAaMiL5+3omn371RQVG7fde6sBgbzDqJWuPmTHZ0tBkW5pXg6yvv/PI2jwvfCh3fQBF
lDXN7xF1ptNmj/I/DWoJ2zKWOu3g2aMOnV5GAOmceDYY8QeBd3w+k9Sw5UBwqAk1NkpW/131dwIo
iVxN83d92gL1kX+N2SUe6YAfbDdchpl607CQEOg0BJf23eA7EEPPn8UMx866RF+OaXyr+LmGU4P9
qqXU3XLOZWmbRJcB7CKwOdRV0GWE4iXeIIUvm/VobugrV319TzD3fQYTrq6g1FahnDFUwKngBGZi
tRk/HTwvueo2oQVBYq7osYfw2vXNeI9eAQlHLSW0JAzJsu9W48kdkklhxU8ZxKLDNi7/aA1rPu6e
WK4Ki2B+HqVb/voQUQWau22bs6wP17FenEOGTMGUV8GK5Le8Q5St8J2q8ziwnq+oFQwI4LduqHEG
W62EI+enZKNQcOe/a/kQ5KEYjLIqNY4dS3Hp//FR0dXZ9ii+rZI9Z3zQzcmy0nZHkAIuH5iy/i4P
5NeUDblSykf2pcbzOKGi3pD71sniZKCnntuNUZ+D7izFKUif8kyHhBh9wX12UHM6Ei+i8QuATXMo
pjzG5Gh0yF6PVAuSMwk0UuZNojOYMwjBPO+gvZH5oRgmB6/nKsD/QNqNRDyvcOp3Zxsac9Dmlktu
0X+dgRCA1OeGeGLlSXsqfdSxla7Gekd7U5YzCoeFMZltCGzILj++QN/0LIf3np8mosUHWuq3qxBJ
4dQUXlnQnSi6Al6kilIORIqxQtjGBAWO3IVEa9im+ndSyXcKCSCu3VtrfnAfG2VpUcf+0iA1HfLI
Cw7ddl2hUqtNMWtHpD3Sqd7Hk/fsgnrYdn8UxfODqTRt741FMkhiwvIe0sAJl0gm2hUUFqnnTj2R
aXdZgmmzUjwiUowA5huykJIZDbTvTZpmzlZ/RLWee/uG/kCyB3yTbA+ZjV6wcDqrG9KHySApNB5M
ErQgF/EakBsgRNh5mAqMOHsNTzx02VE623c4vtBmfYcHCHcRGGDRyr50ICib9uXuQwGOY+iNTkLa
/yIQz7C4PcxzOAyPHqXBsKCw7iXGffiACpbezN/HE4NvvL+L8FQFBi/VM7MfMqRU4e0bpkc0bRmj
40jDe7Mvl42QXS92MzLtLC81NVYgYGcSYLdBeqBmHiO5mYzZVNfofjxgi/oq/1cIemcMwkUysjip
7d1hFcHe87bWa/sij1yh7vTqhjTxQIT4A/NU2o+3QZrcWnm2/YUyL0WcC1pvdYUYdm0juB5FbyvO
j0XnNnPeY6pETa1IrbgIZTAbbRUMZjMicevB+dE0OgpBKB21YRWqdqCf5jL7ojth32PTJzEWhUV0
fIvmLeQK8fTuphluhE5CzWbul24tYPlHC74cUB4L0eaPKawk3f6s5Yepi1FoReGyu2Xmim8UGVCd
DPgywMlX+oPnJoq0EeipdHSG6gp8gTkVz8Y1tnIZ4e93idAd/dLFhjBGWmC8aIuNVOyyRd0p24lh
bwpjHmeoqokecHhmqLcXUEXwe+RozAjiRbrsMSLN7bC623a73AWMoVLQsJGrZmVBFTiWX8IvwLix
WbDOEfaect4LoS9v9XUXh2G8C5EtSFfddiPgw43U/yXB9i7Oqj2U7fWj15R96+DdutdqTk/03i8U
8J/ZurdekO3PkUXo9v9jVmPxPfrGfnIJkGieQXrbl7TRp2+mPrHiuxMMvPPRqA2woBaHo6fEaWAt
bGoqEjz8F8IHyzIwzXKJOXrdMSilRe/6P1sBQbNDRB+W9f93812SlSoJ4GCGx5BV/yCXqewP+GKb
aya9ed4FpUccI46kDCkJ18TnyF9DEsvW9kozJBJ5ii1zw/waA0/wq5LZvV3nG6/mbJCj+/Iz0eEi
hsPMQ+0KQ0LUype8OElQ5MSh7n87GGhq0quTEiz+TFoBn8c9P3CTr84hLMP/sepBQaBxn8Q7vPp/
CQZeKdHOS7EViHqs9ZAJf3i+TsqsIjotmSpwR67U4bus6wIXcZW87Lpgu+SEsjuNMLj95hAe/ePi
apTCsyCdb/ehoTjrAMdLgjK4dujtqFOJdQejWx1BkkWbxFiX3uSZlbA92PK65WsuMdu+drAdwL+N
gPKYNq94WP0+aOnV0o4gZviXcwHIpw3zQfSCDzz5rhxGozzoL/k55bKOPOR2Qa2IRomIRSkop9j8
T2VjWlVTmf1zoGphyQpj6kGSpOBntYx4m+FzGO6RENTP++mjlRgp1BIZilINcpLA2Agi1Nd4xAr3
zrYUvFeEMQqVC8Pm+2Qv9aSeUpllx7PkMzP/gzGnG2C7EuUqN50Ukr724fa9trj0vTJYq1w+rvfM
gFqXjaPVL6h2eCyhk3lLSxCa9vitfcgS7qfOr6haHCzxFp8x7t6ONyvd0BGikUfPgnGA4AUtfg0m
SzwRU9AKyioqDEUaxuoGWO0+tOoXKlIVjSGIiM1xnR7a2nd8BjSXfuSxMeZeeSTv+79tRv6YvRHj
T0kVqVmAP09qG4hzN+NKgHx+hImXiWkUkToh2yPx/T7AtpRiAuFajD+oj5Ey2tQ29CLqUbZOCc5b
2UwaJBoYWiKLlreFVKMx+SQj2PvPpu446wALTZoHMJOLkND+pEx82h2OYgjw5Ym3PXr8+6yKrgJi
Fju4jEJ2t41DS/3iSXfkfW7zNabgekJPg/KGsyJH/3PYQ8KW2kAA4A5a0ihAebBjPTQj/Xn9BbLk
k7WFJrZ/oq1lXcFeg14KFIUXpQMTmryb94iphfg5K5OsFyBe68M+DmRwz3m2cb6FcWtCnr+Gwcr8
pTUQ5/P72DSUXUp2Arp+nUkQOABvdhksJSV2svUzrwZkzjZGahmiy3aUJziM2g2W/dlEKI5w70WE
00nfRC0JJoKkTBLyOsV9ncMzbG4+S5DPzZwbBLBcTY8d9BoZWe6qw7QJXHExEZEKbHgrJYV8WTMj
di900hLJ77jTEzvqyBo7WVHjWgsxIz9MD9ATW0Y0OPG0a6BSLCZ0RZrmZkuKoqskMjGJjayqp7x5
W5Sv3yT2uAlwFNzgXmd60uQew81TX2Brcnk07sKuu5o36tLaJUFAq6Qx3sB2/oYZFtiJuMyM152I
WTe/u8diGNddge6Zhz0skZAU4MConh+paFlMMnQBUSNLdStcOaMAFjYXjVxZqCNy4fjD4sNgjRKN
/jT4ak3cPemmmpOUGcdyiSQ+iZ7uLZbQ85jGMTmII+wfvRfRWbzUzJet/4h8iXBKksizlHZacnam
OD02sro0rrg/da6DobDB3jpfziViRGoyPxxfmkqswjUHNHJwQF681g9FPQlVIzLaU9DbGaCqfHC3
yT2X7qv7Ncb0cMhRGGwn3CAY4n6p8wB5VplbzPTOBB/Uj4GsIDqvhE9bFx8Vp+xIB3rU3/89vh+b
X/2vb1ayPKY+4AcClS0/9NSzyPg3Sa0m59DPfji6M/YfUNw37CbeIsc5WWVmfJjlO+pkgsHFQp/w
RUrdjo/2amI7MFt01M6C+WBUW1Y8S8ozceXWUgNAQ1o5kxZb0dLSKtrJJkiWu0DQm8iNiAtjbXw5
bvbwuTsbv41TE9eqisxdJHbmYujLkli1X4KtB1pUARcX19SVuyLdvR5HTJxWu/lJIE+BJzP0zC/z
Bedr8EBoRzhneHq4XxuRoEBanUobvubCkN/Eacvdhq5/+uQfqlt+UQhvVU082EI+dXqOVO/7kok+
MLbNAGwgcPVXkYsMmALNBIV7tMx8SdNQH4adFjpsvA29pwiIJiIsttZtnp6JwuTu5ZYzYVDQ6Dh2
3rL8+s+SoYOP83/WUfhOr67uydfSpoqGY+oeUrnEhG63YCnkSm3lq7nI9qq0B41j6qV6aRq+58Et
yuYBUnvyQR8vJoCmxKUBlww1QXbMegRMOZZR2/BuM26KtvOmpxV/z1U6I2WWE+6xk2IYyQFzQPZ1
0PmBHhmUt8y9aFrYJIVQHB+33XSY7ATkIsXaE/5XSwdZouRdESvjn7mEKyyHZWw3xD3ZOhsJ1tTl
2OGD5fHNUAdIyKQOuEXDr8dEkYZ1kBPDg5ns61V+twOrhKsbZu9yRWZNrt0MkzIw+x77toWOnDTd
VrP5Ux4jfOXnc9DTiaJBO+DEuZGRA5TfRiK2+hfOh2cCO0vezvDtst5brou7nUSNbQfuzl+EvFax
YW/p+XngZX8sMo/caglsMg8xK36UPpvYHpQdMl81izAtPvAOywxfzn3yWlFuioJinui0Xi4Lzlid
YYf5jg3FnvSJofUD1Z3fc56rt4AyrX59NgpwbYNAH+fdjJUM943t6tAbWT+KZbPMK1uLjwqxsUd+
XU+IJDWWCJq4DU0kCg8fNfrVowWSaAVT05kQhTYfEU2CY18q7oFHpKJ3/bwva+Ti/zO9irNkP9Md
1oHI2/gD3tz6kNWtXMhTCKgBT3s/dYA+oz/7RVlVyn4xFprQEWKY7nAoYWcWnaTuTjwav9wp+acW
3EFnd4Nlo6xRcnEt9SHXMaTL6VWcfZrx0F3z3em+oiV/jwLd+0dYxbdZ6PnMZbuMW2xx1cq3kf+T
P1H9wYCjMenE+4P7sBWKldSUxiAGUejy3EF3GFhihREJQbFPcXMXDfN/eqAUTaxJdeevd5qIX8Og
kRAmonJQdWlg8DYHzfqSNFBg0OJIzCZxpxEiDPvUUyH5DmiLdphoYaa+m1jOR/YoIx9K6j/RI6r5
7SHFk/KLpb1bRiStFwSw/I/WIdiDkCjwR/1zOYH/q3pyagq8bEGgJjIFrC+bf67w4jcu3TqRc1WN
Pym8rgNPfCzbQ/7bXvj1c7P8IPe8WVfo9YUsjPRPNmelOrMBCEiWXqKfbPY14ay6BS4lZRdrfWeZ
5C+z8bo2enhzoAvDzOCTGGEMnN4dXINAJI9Mkk8vjwKxMaM8NaBlVuPxQZyisDe2JQmqibNPRBis
tyROhyomdEfyT/zeLslRA+YWUFky9ohdPYiSbc13Mnyo3jn9kmn99klhDc8BMuI8lg10FrMezjkG
qgvlijrMdJHdsvQFkUvNPgqaVKGg5enC17KqUOYq0blS2976s9Oy62qZ6JWRDnesk04xRJZ90dN+
n90y51KfBNSZp/g9QN0HYsHdseY/5I62UKruN7Vyrxd8HlAnMA4ljFph1ScZ+RbXL5Nmv3b7dvA8
LexWN3VBUUxvHeDf2WvIj1dCi5ENizA1eUA+txzzpj7i+KX+LEOEN+QK6ifKaIz2FIW07UfDllaO
Z7eKhIOOuTNa8vn1n9PZM1zVndKkM+/iAHhYgS2mW4IgPiK4ErLMpunljDAyzYcc7oG1VG/ny7aT
P0WalugvbSyc28C2Lw28ssvrYY6tInGcq1veFhBrLl6LAhVsOQ4K/Md+jCpwnc2vulEw3d+1Kgrc
3pj6GVlwMVBGBPeHwkIhU2z5nDWl0QA4Fj/GEULX02UCN6r9STwmOjrIF6XunubwUTiLsNVfUZFG
28jDaWMRy2EhenXGbwVeV4XHN87s5taU5gXcDcSdQc5j9l4U/ChbeHpIl28bU/GXR0Nj4CRJBqKm
dEC8WdPvCtnC7DXKvpmr8xHrgBJy2bZZgu40ffnbJaCY3S0/tRy09+E5ycrc/XTjgRRnnFl4+2jh
m9oNeiSUp9LDaM7/8E4dVeHKhMQRlWYj94ijIcPP/EqSv0XMCztKTShFPZJl2iQcWOMC8w6HuhYw
Y7FxZOp7HO8gbsn2m0fimkYEUr5xvtI/p/atEeixWMiUEjVsX3Z5O013ZEqyMfJL6CAKbLk0QtlQ
vFXdUV+4Vn9whqAnolXd3YLXu35N/I8CCvi2ErCnlGI9AtoEfLl8A3K4J6I35oCTUWImidr5iVo/
EdCp0LggXAAc6KVzbeEW9KsLpy2uL8XB36xLxkmV/TAb1BT9qzC+b9XF/qFLIpDTyXwLfN0HM16I
Bss4rrZ7XIB3uhW9VeKrMnl8MUvK/8VUTVv+YAPfmKd0/V7idzuF7yNtPvP9zqBJbB56yqvfywSs
98bnrPNaJMpj2YRM/AbkXI/aTWceCZvj30JWNBCCmXEhJBTROOeGdvtpQ3Bkc7aDd1P/fhZjzSze
tv8odwrHuglin3pxY4L6d+sUbU5lujGebSVq56KWw41RAnPAGoah6sIqqgf8upvZGeXMIRgRfjZD
dneoJ9MbvMhkBTrAexNTOT88CdtGBIzwBukrGVF4cw+kMBaJc4yAwS0pjsk9s457tccryx9faZ0H
zRGlasOXk5x4Vonm1rZ8S9cORb1LriWWHUypD9kIbg6ZcWB9XZ2KDWDSDnTKHY0az1p1HJbtBV2T
wmbMb9e4qY80oU9Dow4CEh4Hy4u/icURexO2CSPOkPcjRwuZVaSpUDiUtW7PBGUKpK1n9vN6NNfU
qWYuBH9sjC59sJpSqLAPXAvPi7Hu/Bbz2+1u3i2EPSj4oUD9uvflqH/HdMy07xI1ScHcIFb7qU3W
W1S1nukDMcKBNDzfcNiOdXrr5aS+XUyEisV/QZ0KLPx9ohA4lqaELMC5gyduf9FV8NNTV/zhh8uK
hKVfEbSXxQ7VyoyZhB3XiA1AXMUmSK2uQTp7vuI/cPDvZlG5mAujJ4RjagxSXEF7nZ4sU3ra/lvC
A17ud5AlB9GMhMrP7ZCMGb8wov5E4f0UQ7vDaxdSu0hJdkjuaOLTWYwR/vyKTVen5xsgEkDLrCkb
w5OYCVNIkpTfgRraaW5UB7ByjyCBuyE2u47aS7qEaBW7nTKZQhkRcEWjjNq5QrC2PArrbqU2STx8
50b9wC6rLut7LCWqPGL70SetvS8uuxldmF2169w9f3ahnb/CQAmY+uqn/Au1feM3dNIWLQLYytHu
ejWiGhUS0iLxYi0YSJ+e8qewGeUOXyCLLe0r7oQfgyiUcSZfGgWH2MtltvwGDNIGst8qctYHOKx5
XoSmzWYupqK9gA7JVExFxB8ArN3WdagHkh6P53e1Dy3je/tUSrgtCgJeh+YX6LZosYwdbqgIRXgN
8yOWh6C/NLsA2SeC7hXcY2W5MO5EP1enb2Hmtdo9JQO2GPXuYhAD0KW+sa8b8gBMj78iN4CjqquA
oDGi16/pSgQwVthv/addNpMBuJ8y+IGAVCg3Gwbu6w6Kyv1MWxgn77JAc3zDh4kAjTKIhgCUUNPy
FU5KAIu068bXBobLkJ9LnZF3Ei1kHS1CB55i9/9x82iZxwEYKYEOql3sLLEvQoHpwBUfBd9SGUQ6
qWTeLQjrfLNqjZ2uvZYtEsY54Qsxq4Xgh4StXJvd6HTSaMdeEJ+NN3AyXRHWAjnYhdKMp/qYTAPt
cWJfHFEm9WYBN4ZcEm6B3UEUkRuiOGXyi/pMBhauSBzs71QOyZ9M15bJ3d0s76sKC8dRbXH03Gd2
7b/oJBq/+6BOjMqwjchVgVPBpK/LKQuqIa46Tya549Zyx8DTRJQx3WIg9pfz2Aga8NGlKeMnh+ZM
z324fXm3vjM00/d911oDpeNNCDaw59ap8Au7Wcto5b1GYoHC3t+Rl4vaxvhPVUzMqaLENNTE4Hx4
v2B0wvpuRXfzDWIvC9AolhNo+F94VKcJXXM4vYWDcgn7APf3FSy74jAqEsXArC/5u+UrK/T9HJPF
7MZjt9LKePg6IXl1zve9nz+iaIA+D2W+ZAAdaXAGXiYOCiNAKtFeH8JahgCN1ctBgylwqusoY7lc
raGURLYDJavDJUbry8Uor+sMea5HH+TI731PXujCRSXVnBHfi0tHogG09IWzQwpqkWxr7oMJTG+j
ncRJ32YvzvgCmwTejf9gFff0eu7iyKCfaVsT00jBLTz9RaCanPozAd3SXEaCkhOkXBfzZHVeX/YN
iSmnJfC2bJUPmqb3ebCm2FU0YsyRgRGvKHnmn1CCiZ2zWJME1qjEsrdW6gRbBF6grviQ102OD6xJ
wWiUzlOMneSfOYU4Jt3Bcc+kaVmHg1NiBxdxaEglggNLaMqraHbCHwzKpNBcY3uR9imodJte116a
Pwh/OMVnRcsBB5wZbys8ureC1iyYJhYP63fC2z+SNd/KSjnW9h72bZgX+LigYTkDy3ZzCPnjbkUO
vwsn6fW65h0F3U5nVhr5MttM8fgvoGqtIHU+kLR7p3Jj/3/ptnayo8T/DtRDiCAB5xbjHuOgOdjd
PhY3jR4oFFzSwXdSnZlks2gM8+sspkEqFsiQRSGfAQhwVJHXh3HjC1BSUKWRVhELaF+sC5fB8s4H
mohZCsOIzWaZoEjqf7ayhAtd9ebMzM5q4+bynywzKh4SPxksIhlxyywHPUQ4nMusTy/7H73n4pic
SwcCC2ouUeIrP/kFps8YogdFvoeZVdYTY5/f5BRmx5b4tijNd32Zd25UekbtZUaD4UVK/07y9mJT
l8ufW/CDuhD1EVt89NVVO6T2Tv/PqviLDWu1kOP4sqOJQTXLNv/RD6REwX2HnqHVz5THD3bb5kmi
mIIdBjTCtSpMNnFpFliLIzAopwMkqA5BEtD+4CGJncpNn0JB9/T85nrgKBRrtGRmhGKPD4IMcy5e
nfN5a5EdI2scWhR8XZ79s0li7Cd984Qsid+blNrUMSPA72Jv1QnpZz/Su9zOY+JA3tSMfKwLRzuI
Nrse2IlP26KPGjdYPLR1pZVyb1/ogRixbxJHXFLXwWSJ9plZmn3oqJNIfUg9juM+If0QpF3iW8sw
5L+QpTGOZdYd8v9huK9JSFMQ92hbUoCfuGgtgniFKaCHFkkDJoO1b0G9KOZmOGEzbtlozAOUfGMO
D44xldvhEYnP/Y4DO3eCDTcxb5sUwV5pRmS0wzr1PUmA3jRgzedTVBUVM4UkhYrobzLUYstuQswo
Xs2ky8qw7wzMjybyJSpirbRfYyG39I053r+ClzKaP7G06BFEPC83+sxm9tMV1yiJWJhMsKzzOfuh
6WfMNYaEUFv1T/BZ8R3kLi75pbV1daSZqPtewpCdeCuZNx2ow1N97WK+QkdFAKzyR/1dVlI7pyxH
gZ8oc03s+etieTIO7P7BWfSjXo78JkJ9QC9+AX2w6cIyAUQrb6X4W6KHMSqvKhiMf3sCyHvYKPcN
dFzXpEk+mG4kjIqo9nHAjYipDxF37AHubm18rUwz39puon1T1nEVOdGpuO7Ml+Et+o38pmRHKZ8C
Ezr6oF+FdQROKy1Vg0gy0UaXkKE+44h+7LlwiaagPEn0MLN3L9m+6rdxZ5tsMnQkim0f0uzIvb4C
tP6T84wWeYpg+odtzFr4NpsqvQugEDeyKFaMpnH3ufQZX6+YNkdYCRGcbQN/s7jz4uFyCOJtkbkx
c2CjyfFPqMhPmU1sCurifZy9E5DxGTe5sAB/N/bUpjNCShF6nP3y7/B5t9FG1HAHgZYXpsrhLeVt
RAsx67kDfjLqD5fttPjhiSFMPZ9hX6RpL4MT9cPKHJiNs8Mx7zSlvOcmPyED1Xhn8QJ5G6KMY7oB
naObNX8r6UgaVsPaLoghnGZXOfx675wXj39UFgkM8t5EDkJ5igbHy1QsObsiDXx6GsCpL2ulRwAB
MOLu0DRLJeTc/gMTTe4/TJNqmxVWmGE1LVR4ENrD1oVBkEd5iveEk+jjSscKu9RWbWQScyAqTlLG
pC1u0vCCHtOFxi6qSL2gjP4ObqO6g8mfOhFdNxGzrMcN2GuM7b5wm1P2NXTaT0S/AVPV5y+dGHzb
UpgxZCfb0r2GMgAo+e2Ng4jVoK6QYkZTzfjfDI2T7pxgQ2yfcbByvBjrl9ZB6V7LUm5E3eWP581n
Y5hm5iraIS2+rXWKiT4Qh9aI6G1/g8yb3D4d6KbJ8PwzBxW4frGvwJr/MRZGmTVoUx6AjbTrzkKs
JqaIdb98wptZb5GWnkg/34xdmdJTWpXyjowCLrQ6/i3y5QUhTs+gYONnjum6djaI+zTDes/zULem
3jogE5OcamkN/DXD1/1V+0RU+KzWNL2rVHdtr0e6ntKe9rjNd1vLe9ucuyTeRuYc2cpMklFloNiX
j42k4g75L2okD5GjYM0rj4ta1DiwwKmI4PGqoGUMp1XcmUrNgloAPIE2x3oPWTmoQZIk4lRm/c+W
E2VS3OMjsRE3cTq0/wnbiywrt9t3wDSBuIrfDW+HvjkintEEPZ3oF55ULEkLpB60DPSCMPcCnK8w
Zpas4OVgSDS4qEVGLdll78Wvm/0W0bpdx/gk6aEPkTGWU94rOZMIHqOg1/EwMWaHbv5oQeA5HbOz
G067dKnD/f6++hE4Obnqp75C3vLm6Mbr4VVm3BJ3asMOp2/gye75UuXq8ExgetS8tLefaXgYsYLF
+LDo4uuP3lDA+iSR9ppEJBnuDrrJuO3U8B59U6r6iQL4D7NGj7n24AkU1PRQ1T8mkrFhirTVzou8
NNgjx5I3TvJZ3fwmrHV4ivbaW1pWtwddK89Kyfd5JQObY+qBEPDOJn1/wJNGerix7EJ0PCPrjGOX
Ds03rZoLDcq/449Zk/iaIwEf9CyjRGlIQ0JupgTTyUb9/QqMx+hk+Kf/GdmAVYhp/BY8ZUKqibzK
a455HQ34OtJ+UN9EpVwa6hsxke6KnNVK2UQBD8YpDFY3rTT3mUwkDbn63p0z3NuSY8SF4BiZ7vA1
G4067qv7K7KZStLCodfPbMHSQY/WlNjnNPyZE3rjrg3UQlJoV2DrpaYtbe+bcr2nEgUInNjUDWlH
a0e1NbSJCpWnPtrQYLK5LovwzaiALtSva6CA7nG2mZ+VgsaecvJFc+wRE4F/+t/IdkRntRcNi8WA
X1bnAGGb0gleT5DzBwS8J6wyMvGUj/WZne0pcEznmhzuMRq4VK5yRr8js7AvZgeNzihqoBxYQGk2
9nae/UYKfyZjX0g/HenWbgTaqMn9jdE172fP0eqXeeRaRIddetfgL4jMp8ymD/KNzN9kBdCtdMMz
6o+SjS6LJojrhHBRcnwFahi5ix5ROsaSmXMJFvdnNUuo3BHsJISZFwjUGYBm0XQF/o+asWVANDVb
b2bqHJq6iJxVV/hKNiRMIgvh7orBHu5BtCQCpwVROk/5/1WU00nY6DmCbcwfzNknt9Oi7lSjjND+
6+lfK0f4+S3ZyaiTtpUE7ApkJSafXVCxc1NdNIrd+Gypj2SxVH0OY4a5X79bjoQ10tt3R1hY5esi
tnRbVA7CEUIUoFm9j9PcyZCcOlfQ46js0dSTJoVqFH6ssSf+yh4vKpfq2tTLuszJoS3RE4LFqA8n
xf6QGg3Kz0WVNt1i2dn4phLTqc3DXl0teV8mFgfBI+XNgxG6eXFFweWV4dQhsRmXbpstFQ4nQQq0
z4E6TaLdmDTOW2MTlgczp/NczxpO0n16YMmME/AKZ7FMaTR9H6/J89A+Ht6D9YJ66/SIt1UG3sOL
FmkSIklCAfZ8RdK2rHbyAHD/pCNHlugb0GtZJgeSY2//knjjIrzLWnlQGowqRvumpAFl5TG2RWaN
ukgBSkPvUtUNOO/W3WLwpfwuoRGhNN/ukcUCjFrRdeWc7J/ij2FHuSvke5j6mnH5NRci0dbBQXB5
xqfaZxo/j/AAtQctEBADelgVBjFL2qQxzND8VfVXihc8J2NoLLw58Gy+QgKUNGlCq10rHP3ta6Qn
HFEc+qaKyiPv6U1LwPYTLDlwT5IeOy+b7HglNrzZfLwmow5yMopuCDN9s9kZk/QwJI1hb8R+trgK
PEoBrTL+rsSq++66IjaQy7HUU1EyvSAKwvmbLNOs0GpUATQI41h2EYA9M9ZCwMZSgrptJqLLz92F
Lo1DgB784S7qmKXs/INxseKBEBYXmu4Pd8oDiA1TQiZiD1NjNGNbzDEgnQ++pEktXTTwkN6AQ06+
ZXzLVrIxduhgPQBGSBX1loTlzY7DSbYimE6QAkKg1kNBfVChxi6UeDM8JgqCi09fiFlXrSsZIITd
xgrWAnyV1/Kvoud7Mm3c+CB6oofbolMt2yYcq6wNJnqjZWAcKZU9aQkRs4RGNidfirpZ+M/Q3Xo3
WH5swXdzT6XJIKKYcISg0fKoU/dEKVqgfz7e2uZw5oOOww/R4RaV6OIyroozNj8qwrIXzRSAMs1g
0V/5zKAaQWd07nik8utkS4VI5H2VRWeRc0oBkWuHIKKuDBTEMjSwaLQOy/U0WtZHAo4QOlwmGULD
wfK4nzkIOWVMkcJVx4+zMUrI6iN3zadNC2AkbzUSqBgsMRabA/pkc+t3FWbz9mYYqW8zcv+ImKFG
wZI/L5I1C2yDoX7q4z0AlzC7olBWKLDszlm69V1SAXcZQ98K061TPj89tooAjcEjfddMo3dz/Wtq
rhqTQGYb2QHK8OUjEYl71GKu7MQm+xvh5x5ZvNdWEprBXJIHAdUDQJv4MFvPkD/c3kLStUELWPBd
KFqHhfoXHyrs3UE7vWf+Iew0xVjnuDhBHF2dJin0TjP1bzZ4EuDEjEmagk1e+vWewSH2B7V8qb+5
qRvynq5SVjdnz76bhHC5Qq+0xjlBK2unVIBF1vvz1ooiAeqWUvsCRKTTHsO9fSJKVsoDmtkeGYb6
+6rsGyC19Y3S2OWBIJzh8CSssHoTNMi+QWCOxI3CquMV0JEG+pUGwnlEh9UyQU4a62Juzsa2R5q1
Rk3yX420C7oa8GkOtpFMnwRLpDUPkgHaep2JPpnVw8MDqIFob0B2QkTnysDH+juvfk+FVhHNdrtV
zL8AqRp2syPJ8F3QBIEbu3hl91U1VGEK8+Ducmp90LN0PjjFIcEsaueFBbYFPTg5UZXghywKE+Ho
b7ys5CxmNLh7AJzY3D4HHVmh2zUT69u0kLB7lgE7embsjgp2hqaz/mF+X3AGG2O0KD0rEGNbdBlw
BT0YqwCO17d9DpvInRYY/5FAPCe+IjWHIEpOAbWzOMcLdxVr6SEZvaBgW25QznEASIm6DeZqAKFH
/rGpGvm9Nt3k2g9HmmcaLkICSOKJf8O6ILdIjBFfHhhERWtYBDgGZOgm4h4DPZU8FjWkQBPNI5bt
NYG7G7+FBbPhKzarTKi/p1LfWYsGJoHAEV99D/EEWg8syigTdH7UCzfjgFgONcMSgaOpgdeaKZwj
Jx+ntbizD1JTOANG5xQqdeuXuOqIOAfh5uLcxdG/Hu6klBmbIVXZc8dxhV6O5Hp5nkgiHfulsCWO
NDL/GEVa3UM8rZ7k4xBFRzuuKY8nx/XVlKHaDQjuU7eg+aicAuBEH4AgOKPT2BjCLr6yuRKAQYq7
GjR+6KR6XD6YlBbAB8WvveE8wSCoMWwNgsAR1noWs96tsnzTd1Sv87IQ6vASExXlNSWAGJVRdOXp
qBOo34ghlKTvziaxRDn+EpK88Gw7EhUezMrfOjtHja4AR7VI0kVMTSzMRLdGFpsoLrvfxfcDOKfd
q8jVzRfg2LJgWFbe5hVDqZHPE39j8eD+R+eMrL8K+YvZsk1/zJBNeUcahPwl50JG83lWgURwHeEs
lR2Mi2ZtxlGgf67b4YEwu9QdNLjy7Q0o7jNqWfX+fEK5N1K2tMhAcuaP/1l5vIwc5hlmsF9yeZyw
Q6KBwgMRySsTHjvjMZp90gwH3Hna3TRlQqyiwC1g8Q5UEmfinPoKL9vRGLPQPapkJ5EyqBdM0aHL
EQjm+gj9pJFJYpIxTodyRDe6V6uCtkmdIhFYt7Wgtj2XwZWiSHiBmdnS/wwmH0LxcoInVkQsQFwD
ohu8mc6GYmsMHH1G1IHkcExzPUv6uEi77bdDi1jqyRjcoq2SeEQZX1LwQAXNnE6JXOlKivWxixcr
AHlb0xgkv6nAEeZvguQy7wE4nyFOIUh8DfIWgnOMNELSmEmKjmHJ5WsVTuwJiHyS0MWlDO75gv6X
euo/C8Ed/IDcsoFneIU+40qd1r4Mf8fmejuJQu/h11H8X1nLZys1zR3v3eRarrgHPmgfRKZl10s9
c+kbO/ro3lwUsviGNF+yjVjPJIHXteTHZWhISbqrbReSzSu7WSERa3wYMIaS5QAxbqTcH2UIP/Jj
xQeqHYwl8CfJ0abwCyMr9umTN2NJtIxzY6EBLjiSWdcjNthuWJE87SErZX08KsEEvGyabwc0TEPB
YZu9OGI2E8Fc40RlCjg3fNtAwZbkU16NJmWNhz3hJeJzgNzdGlaAGVCOD2dmekqMp51cyonnQ1Bz
S2bQRNYXL3IPXasZ4lV5qTFwEfEuhNyiby8GkS16wXH3dXtfGS+eEdgUtPs9+RcVhCCWYK35jfFn
xeEvb4AU8nXoK97ASqTGJuK3/8U/vtAy81Br/NOMqiMtB5yIKY9HeKiXvOEcW34fFpRNSMGJekZE
AIRd1NlEVlsyp7S/1Ue4zEagvAL7gIrwIxYMsVkUvvhWk/pBWbQtHRqmisLm+OtHJqbQ/1/ppcpV
NRCEbhvT+6ZDK8F1weYdReq6yQP9gE9JbnPqNOr66qrHj3rD4GoRHVX0c15Btgk8FPDsr9sDRlzO
3TH30gxb8Tkvtmr9jurHX9OLmp+FRAAgxj+EEg8ptSVM+axYivhynJ+oFc6Id1d5tw19Eji9Z6EO
K1cE9LOrXfIF7jJmVN/EFOMkUOmccW7sKCBmB+nu8Ce/JtRAknEbDc3IWBMV+g3TtXWnvUWElcAx
rv7ypkYLM3MYmL+DU1UvMMkHvRYRqjzLH+JgkJVo4ecftYFLh2Eku3J/DBK0cPakimIcwpG8Em8m
qd3tjQEBAVsvKF4z+dCsb7Ahw51ud2gK6HGpgGRuReCoxD+uvbiEjLAb1+p2/leUIHXlPiD8eY//
qtuK7g0whsN2pVFh4FB8p270DafLKGdw7mpYcX49o1F6hzHSdOX2QDtMHBlZE2HZpWLu/+7ofJ0A
VshiUfpBiW9jzYAZf5RNmMkqaxKF5iVtejfBxC4PMjcPEm1CL1Nfj1K+Dpa7K1TyXZ12NFyNGN+A
pX0sLBDNj0ylLcjwedGOTdjsYMmNdGtuT3xE8PeX3qH+JTvROtyEj9U581rThniXVAMuUL6rbnPg
nQOGArGN2sLpt3mqL47lb8yhtu2FrSd8dpciCCzp7hVXk5o8Km4UnqLpgnpXxjIcgRRcxFazUe4w
XPjONMJzmV3ZlF/TkPfW9cc1f3koiLba0xoeqVmWwlDyd+Yvv7SgCZ/OM0H1819j2EXr0SWNXiAn
CIkjF93Um4Aq/gpi/lESapjKt29qeQHHZ9lLdOqYoZA1EnMSdcN/lC+aIWpjb+O/umqLCXvd/nm1
nlgoy0B277d6BfOjEpt7GX8KOVNCosExxE600zdLoxXOKVMBwlpG7zpBSPBF1HPgVdYBchVZ/deN
BBL3G+G+BYqVW1S33hhq1ZLtzaaUG336dlHr2qoEx2fhygclisUg5GPfL4sORQSP8UdraOhN+ewr
LbE2XtxCm4tlHnufti2mAlp40ighl5qxkfataZLxKYptywNsBr23LlsXrqWBiwvkGREJApDNkvpW
FxNH8KLKtA7s/9xVU+jXOZZwyCewR/Ba7pTT1xdec5RpQbEc5888LqrtF+2e4x1E3HTnqeqw5jhO
RoKWQRWpGQ6vAbtppLhhUDyb+JXgYluBvXB4Dqzubuw2ThSdiIuSHmTrtUDbmtwZuEY+4jV4SmhY
SRyDobNFaioPLybPRULI6bZyeQVDVMZ3U6kPi3q7vZ4A53TyrftVcqTRWMNAnNoK/8wZ4jQhJXL/
5lrRF6yvBgPeGgJcDM5jW3tUwocE+pRcSTqOF5c1zPBYPGU2jOQm2oKlFRm/qdGVEEQCGPMPhQ2P
cN1iLhUsQ80KHkfGPkDn0Ipj7zCEAu3V8QijE2wsKR3NCvx1N3WpnLwcNJ5qvxt5qyNk8kgJF7qS
KUQP8ucCGO9JgsQ0OjgZ0AFJeNuV5d7JtqqYp7xS7jW2N+6ZYQzvb1rXrMmiksCiLpSZ8gtRyJYD
tAgRZPjb9hWMT4t9mqTFIMZvra/ix1yMjWzed3fPGPjrKpsWjKmvw/fgwiR1Hd/0TE5xOAyQiQF1
2uyp4bpnP79g85MiyEKbvZXRrXOriXZTBZmkOpFO+ptS8i0Vu/IsQu8MgGgYHcU+F3CmeLu1IZ6X
E3w+HXncDSJw8+5IRwiiihGiL2ZL/9Q24khpswz4BbS8kqjscNoKdTZMcsLu4PX11gms3dlOKtK/
bnk9250Y0T1p8nsU0vhZyIL9Z7gk/kHz97168+bx88Nj8G/iBKzhruDQd5N0ZvgCfH3iDu2n74xZ
3NqjajB0muzKm48Q8Vu73s1kWKWgTXsgIS/cbgzg2przZ3JLOkEQlSNk2dg1/l2udeaZ77vUBEwa
7J1QK5rIf46ZwPK5YhQqN9LTllIxZF6pycamb7LKFytGT7scqaa7rlmKS0lh+GZn2Giz5zttQCsn
Ep0AuZTS1HJnydEpyRvEX44HiEgfC0PVLuohYQN3lFf+Pjl2NYJ3zFiybcIun6yB4PbIKbXr/SHJ
bBk4Km4fVvN0SC4KXr3EHO2lAiXPpAViITIfdo7GERlVeXk5C0q4DA+NcprzGpOkYh14vtvHwVns
Hc7EhBNIgOOui4wY6yMU7mw+zP8WJ+JoVW348bpWwsvOxdFlxHJuYlQxZ+C5YQSeLMe+O9aslzx5
3R1EJ1Ek3DRvaqYJK931M2R3VAoik/QjCWaYHyoACmZH1MSWKppx/HlluIBckaeTKr2VXWxShRUt
4/9oWyNYQwFlLpUVnqG0DpDaaJXqk5roMQ+M4GeoDbl2ba/gJhiqFm9WZXr6T2zAmEA2r5GQjq/y
9ei8JFvBp/5fPKLDAKgujuGrU6ePHqzIQVnS8qvu5pdb/mnCIPVXXf00RYswRQSn8f6IOps74ZB3
0/11U2Vr76faqXqgdORLrYMC9KiV6jnhnVLdLGR5CEFC+hUiLqdTo7crkapqusobHW824aIYvQil
gqxzzav8QrYefwLr+mqQg5Pwi9lh0jYmosbIPn+siLh0U/Qz7K/39tKrNyaDuY6CKQKvXvLWec6e
iGyrNvYpJJef+Re3dKRTAZxp81kcSc8uIKDGsTEhHhWyRSFRnEfKbKnE7K1yFjPUTO1qeKn1Mtj4
PTyJhZmuOBHmNg60EY8wQ+xZY91UoFd6UYEEtQoE52dy0PCcueDE5OaXlV3eGabl257NJ/xUA2gp
EHwOoZSZDdKp0y/BfgL3I734XUYrIXm3NkMfhI+G4DWWhPEe1faCdNTHYVnYIqSLxlWITMMbP4eG
2Z3saYOv6fWHvmJe76s+h64c6e7fk0dnzHph+pOXjWg/TU34r4ve6cpnUwT3gDqqlw/qJqI4Bk2I
C+BYvQ2Y0ANvnQAr8K+uAoJu0MKDwJtv8+pq72H6W+ACOQxjnD+MC8+jF4oCve9/Es+MwzqxtTFx
tU0m61eIRhG1CvtL5vdwe+hGUqqfgObnBfsWcM/+TZa4/ziUJ+Jf2IM7YK4Q6yPMkITvTCHTGjDQ
5svA0ywJNaa1JOPzumZtfGaat/UXlLzUCVMbP087E9qCfdjpdeBhTi5G3uo8SYR7yCYdpL6xEVpg
mSY50fGzRTED4EkJqysnp6QvoHZ65pbIntCJdl+df2Fj9/oICtEM26eEP2++kbiLHMCeBpTcxMmc
YvuSFoZsd2T/2tPcAb/FbFd22UbX/M8RnAzqwIpkm7O19W1WKNcudNHy4T3dr/C6OSVnPiGWlJIN
HwJ2Y3P3y00WqFwYGzOijeAEIANZXkZy1b3OnW8iS4pGBFqdIhkEeCjhk5JVBrtfinopQrSHu1A8
SHCgb0sVqYURoRQpMWUCGyEpjHr5oxLr88TPRjvsJ3HljcMUV8M+T9nKtzUJSVngZ0AQGLt3PkLB
wQZOvO5jDgQ0iB8Hp8AT3FdfL/xdu5zVdK6g7m+XxFpBHLVT9etRQ6xIwz/yjROp3sivvrk5W3nL
WriHkBG4Wdr0dzvW8zb7rceZdzG9nILyI6I4LE94iohduPBQM1QIfAXzcmJ8xpBP6B6NaZ7zbSUL
3VCgoEQ4QokVCu8s3d8dEqNHQdMdfUN4OUahJ8eneHosxhUB6s4NssJ/fF/eiyKuBzKH2MhnI37A
KbkGwqq1cDDTahNIJFb5PgE30/RRrxFzSDN06AGRZiDNyZK3c5n4tjrwZu0q2C08iXMDuU8FJIQ7
90jB650P59jO5Bx+gjurN/yS8vh5QMCYEAcnthrrI9AdtZyGmo82fuZSR6OtHhyz08blxoBtHe6h
5UbT8PL4HwVVHXg4wLw2sQ1UUZReeOD+XrwVel9HdSIzIFrvSH4dK4nKomgHk7ThFw3d1nO04OKd
3jSr/qzmFjCBGKmOQ65rXU03y/sVMoh1JdeSGDC/nNoNasMpKkbqTnz1ZJpYYwOD+Df+p9xkGNpk
0rgSmY6OnS01lnYTIO0IlNPaFFonbB/9NwOeeaNK1zIytPHJ9pTPUpo+45AMeUe519UsLQV62BfE
abes0BYIT03GzJOcjipuanHGD/inroUvAV4EkcQksVwb/rcsmTSdbPe5UwkFDVtnETvf6ZPpqmiW
qpMjz+4fzlf02EleWaEtcJ+nKdOqu1ZbImKtqZrYhJYew2t1aapsgRmGyaXtB2Y0rgaaE7BUZXHK
Dhh3HaGEtyBXGypPEPdFQE8yttma2kHTk+CuWf072BTUmRrojWZWr2rLrQz27PG+obTRf3d8fCaf
Yz/Uiqf65R5Pu7qTXL2Pc8GBfK2qgsff+2or/ryUfoYwPx2g/qMa7QNj9z/QKeRVpTBJZl6texlT
DtmDqcFvcu7F9Nlx3Lq6IcszTQFTARbZ5LJnnnKdl5qDQxWptei5kMFrQN+fLrtbLPdBViJ1GEM/
svPvIaUebDJGqA/V2rgse4hWqlkuL/zSWch1c40tdepKh/Ss3lJI0acJLZEAMhosJ+dutm3XMjAi
wI+/e3eQ8Pvf2wDVG6EW3yS17Ex/pw1AK4EFnduQk20WHid0HK6QRlNI3BJG4z+QMQLTEVXfoMJ7
6v9MEsa1mQP+iOYNjvdozVyIIITQAqxwneIs1+RK0byl0JRKfVwR3huqbNoLjIi4JRNxLKmO22s7
7ydopS2XJP1owi4SXPyFKdTyDqbu1jfZ3TRtF1aanwWwcJOvHiRTcq3f2A1+4pp2Znf9rpR+tA3A
Z5c4olH6unGrSj3FBP20/ZAadDkTiBvFgCpiFIohzVKDSPCewxxoejU30RP+ledacCn2vXfPH3/e
kAFyQmdV1Z16lTkatOHfGr8UazEXo5GNBG17HWWDt/E2FIDO4vJipga9zIYduPrdjy7ehsC8xESy
5bXwa7MjjI6y+2wYGxEMOWCx6rPZnboT24LWNV+JtpXy66i/O+dU+DrRolkPczI4/3r9XJZzx0Jq
mfoNquSrCCT6CkGj9iFKQ2lxDj2A9Bxz/SfaS3eUYSNcNkislK/nINlv/DwCw3RpPEneu+hOjnPp
36guhXmanVCSc1m7Y+n2d3BXANJBk5Jdni2KBzsATICxaCrCPOAtVYQTThH0TxGQJ159W9QrGa81
IQNw6o9lTyuUxMCvCIUAu4UT9AEiyx446G4kxm+p7ZI9WNxLISZoupmhBE695OqbmFfaOb2PadCe
86ZP2T18TBMTkHL7UFPKpqDuKxBDvsCrPUQv4PK3JsIIH3FFaC3oMuucNCIFh8zLf3VC7naQ6ZCZ
SZR4Scghs9cxgendTpQZ/kV57ohaDiiPXIcIqeIpwMmwHCcyhI3SgKHUfROpi62hpSfdgdTLKurR
nFR9Css4YmF7jd7J/FF1vrIDcwiC+Y76pmmw7II5HHz5foWsRrtU4CM1Pq88kcYi3NeHi/nFt8Vc
SW2REqUouz9aR4VyaUvooH6zDQOR2zAEu30NWKyF2NGFcfEq69jIpeNXJXPsl+kj/ElyJrHHqU14
Lrat15sdnUVfMZD8UyU2HrMVZfEpeMFwiTwGZINb6XDV1ABQp7GmIKrlj2qpRujwAKyohfDW/Rwn
TBSzO9DyWIZ3zGkfTr06GDUWDLbO0T6iRkiyNHwWDciprvdIy95umnM59xTC1UQzl74BMVGcx59v
qAX0OPfapujYZ4nqmo6Pw+/atzMFHA/V5QxkSqYxc4RnV6ydPue8bV4iBPHT/kByMJ9NnJjEr7Io
KEWnyNdp5u0U9Yj+gsOXsIdW6Hp/yF0preoPBFeUPcYSmKKe2kclq2MkRjf8SHelSssgIeSBvnQH
anBmp1kK7rCw16tK/vgD++ftU+hWb/XTjpN6hfWWmIgWO672DbLjJcGq4BLIy0qxv/gFxpj4bNYA
rPlQ2k1nu/Dy9zeshbtqpBWf5dVviGMYlyS9Gqmv8I+/BROYap/6WPzKvbfUdgZSDA82SCeRLMRr
6zRn+e6eMfSGuLs3kS0u1Y+50SyuXVEfauUzV4S7Q5vDdt5mtMzis15QSsSTN+MQVIX0HMkUYFp0
/8Io1/OyvP6dvbpsf24lleVeJwCEo1HKLpPcYwR+SYS4AGN7U/qRpmoTMANXLssJIHFUy/VSgaq2
0Z8y9UcNFrJ2Tf2xqhghmR4Qw6f8tymmCEujPMZ5TbFDl8qBPzMr43lFLccLziWHt7Kvlb05bZ7z
jQhxASWAxwxVj8W0bFVI3l4DvigsraDtpka1BI2hsoijyItQojn9fgz6hXZa8WfhrePuyy5gX88L
jUxxmY5z5ueqFPru3Nn8UEzpJlKQBzUws9a2pKDVg5JHSDd2vAg8yVTzHdI0zmpVs3NhwSrrcbhb
v9dUFwA+BbAEs7mKC69oyNFuOfhoRdTbJJ/aXdVejyJqs7cT/TM8IOBD7Pobyxxcm/lnfP11gagK
HoKgZQ+fH3Ztl0kDhM5G9+xr1oFgB3rsy6ZUAJMznvgaNyY+gdp9EkaF8UtcmM5FDwnkUQdFhyuZ
m+W32Q3KxmN64Wi6g47/b4cOAMu7CrIGqsOJT5hatAl6qpyWW6GL/Kl4TBfdYEt4aZTFPN/O7mJi
U7RQuxzey5i4PJvKPe3N2rPqEKajwOMMsutW2TaIjz7FeEVhoX94gV5CEcJdKYabdAvXCCGUiKgR
irc4o147+DYTCjpBpjBIYUaUg1UCdk5yRmStSuFlzEUFCWNvI2z69o7hyxDO1DuWdTp4p17AWg63
/LCW2B7cHbihdzGmqd0yrRGnGQ0f0zEhdl9QNlh1qhe9rRf+guxLRrkZPDOEzEOn8fc3z2TFZ5ia
uqydsXQQNH1uBRBHVrwK/nKaWmXTE7+TnQZ9AuXGgd34QgGXd/c0M2lN8UvYY25mD2PWNJzvmg8I
hclpTCh9A50ayA/l+dehW5NwR5PCSHBktDioisWYnWUi8WT/657hON2SMYdLvW1OzeFWO1cb42vY
R5IyZaNxjSbR/0C+8DX4j5B1kQlz/w96NotoS0rSO6ybINx7sL7iqILjMbP6nV3sMkhG79NsZUtq
XxhuUz7ZapBMgLh7HBMamtRbEJH9j+xwynahc/x7HxRnZiMwEGn8nRLiGG+YB69Ydx3moY/a8wXy
auN2MeKBp344dIMlCWZOPIpMlk49C52yag5kmggpJA8vqBGOLwqjtONSkJez3FToIwoU7SihYF6n
e+NbFjTzqhkZ2iTUBIn5QOmkME1V0cjHWu0yxngFmCdk8mCB3bdoWMrBEtaLg9PFVrJWe+/SqXyp
9/SAbb3WzXfkHhN36yXQqqI3s2H4wGDeq5KUHaYr6p439hPeLTUWb4WkP5NfOGltPTzp0QRAnV0i
tD6e2nUQ32kjgWhb0v+pPRHPQwZbEIMaGbYFiJY73THjvCNcEgtsMYaxNavqzA3SPIR8VKLhmhnQ
DYi1weQFqd0GmlKO8Uoo9jzD7E2idrVAs9KJ75NoE2TiaFE98g6yYwFKswRRbcsO0Yy4jIqFe4zb
J5DwjQ/hAZ4LilQUKeA8XXfFgMr/gwLlm6wlw016e3CTL8kQzM1sQaQPfkBwgH6E7uyo5aiYHPa6
ASkPl9U+OUo0ewkrvF3cnxJOW0f7RJTNU09a3telXVtEpRPCmDPzJrpBRWIQAyIYxEzWEBGjcbbQ
vX/Ll48OGY0Nu9Oy+uFKWPM5xytayVeXy+JpFSdDODvtrDs54O8W5ph56DbU2mNgbA86gGekJUAg
mYMzjmxXltY7h7n5YxNF6NeRb03P5iXnoWU0JxxgeBELgWVaRyVbycbOYrRko3t2wOitdGqVABd8
uXSVNZvb0n4YF8pbel1581FoBtHe6PN4bMbvvYmwfoBYU6kiQ2VpJ0Zu58yVZ26leWjtg//Yoy2Q
NlKyvg7/z/Ik59qrQjSP+Pj3Np7XPbs4kgpl6PwBEm5KW9hvnd/GXcQwpz8qwKFZ1FWysgF375ry
8UVI8fS7qqab0WQ+pXSFDb3V6OWZp4eJ8uRzp4za3vh+XTwH96KnT2f9967Thu57V79T0q9vH6ST
k+8hUr1EKml13HLL6Df1hu9pPimwkq/K6ggpoWyGeOXBqLK4Tzpr53EjSlU7PL/Rlv5Xi1CsYp2E
5YvGw9Ndxp0N7BBYGEQSug3Kek/UdDOULOqAFoBC2B5PLzNAJzjyvHDG+MOhtY4wL7pzoAfmlv7E
xFVoKi5CTkm8Dk22O3HO8GWO0meZ9qsbzQoW81GXMMrRq7hr+caAuA7tG6OvVT4BcHQFoL5rc/Qt
JotgoNcNfCeccTAolmLwJVkgttrdYEM3e4l7ssbIauaQy4xAZrP3UQq9ammYYOsNhZRXbIsT4pAw
91O6N025kyuPLC7H/1HY9df7SMXisycQsz8cCxqziX85vzjmqXpPYHg2jOA+tmcGyDH/BOrCZ5hc
DLVDGo0LbpTG80vOBWr2SrpgwGlqdgF3wB093Vja4h6sYAXFPFxr9DpoxO0zYpD/ECZLALIjz8f1
dlyUJGcr9kvE3xPn2muiW84/qeHeBzpCsCghBr1h1ZwfFp642CvJSEGy2sx8saYFDylQurYkpq4U
mgfXKxX9CKwhb+o4hzqNEFmMamsxMBIaCgNJpiwYeDM5i+dnZIvHfabC0UGS7qsxln4esDALBZsy
9OXtZQsHfSNGksm8IHD4VBNHTZ5j+HCgGtZ2REKw5nKMwsCIKf+9HPVSSik9nNPvqJpX2357GcS/
3vXa0vTCOWKHwNaYwWW46SVviOei8Q4wSvMClcE8BSv7lFISNXM+sti6nnSEhn2Otzn8c7f+elT6
qDEUCllwcRpBr7RyBSJpIl8l6NZU4v5UzVRjQzaSBd9F+QDecCTNO4KX3dpIfVIBDXdJF8j5WcMT
OhI8ZbxgIfmLsCGtXrRd+4JUQrtEtVQ/HdlXMHhkIG9Nbr0LXKx0wI5v5MbKrglUPD7PQSP6zTcc
Oq8hzKPnY7FxoI/pHRVjoyRMyC3V9Y+t/r9VK3o0+9SFJOJ/CPdZ8PJiVdXq4lJElebHRzqgBKWQ
j2GtDVZh/hcHpb0GUsWejS5fuu4OkjIdhnm/fJF7WoUBXbLVOMU6HNNM+9jmYMtqOxrYqzXEXZP6
zeFWhFU2cMIhi6heeRuBGH4sWhAQLUWVYmyoPQ/ZGHIpbe8T+VPXsTNdFlUDsk+hApbL8kBqTJy0
5s36H1fB0ufpzgUHa9pZZO7ixQNadFaDekuchKM8Ix/tThi8O23DqbF83HUwi90BU/Ef81MwJqVm
OfkC/XbIfA/AuRyLgbo2VF7a7l/3KeEhKsrGyuvqWI2/avo7BRgAwe403/z60wc34ZC4A67DDwiX
2ocRhil41ctSMWoxf0SeaYKbOnjCml4FiZcrW1xuBFF+VGPhYaol3lVNo/esh+MfBsJ19mieZYrs
iBdMn7NLvKgmGCVugFQxO4FjQMosKwVMSgNftxsbY0ajGFVuHoLKZx9rmKPuQJz0XVBrqwyad7//
fpmJ0sVa0bhaFiCurz6Jlexh1MeLtrojbzsMZL29NkAtxnBfS6y65Ep5BlbMGDytZu8bZaSHzxYN
zaN0j7RTpMD3cnumzsBciOSwwc2cigUS7xQfrczisdrJ0/Hx4zkW3jsgGePM42dyuEhey2GuFuHH
Rp87g5Y/qZolecVyDaeT0FeSw/B33girAXPu9h0D/36LriCuKv8ZuzRGgMASt9g74DoT9Jr1Ix26
Dqp6+1n6YS9b4oF+St51RTLJs7Tx3b3C4QVLdmqYJ88WpyFa157hh02YeqXyJAmEOUWPTnfdIl1m
tt2MuRp6Gkwp3Md29DLdIy7VexlpUziCt3UFz6uIBMlfSlil5Rsd85/b4jzPPrincMpcYJ84ZAKl
yiaR7frJldtlFcrfyRTWllXusVCk8zxxan4LSmjKvV68ttp2uywb7ZIVbwruZl/MLniM2NjORxJv
iRRq6TmcPRl8VmYVgd04UmZQzBQI+MUlYBjlAPG20T0/yvfVsRHtZ3TIgiVD9tgab4Q1XhpSdlpP
4p6iEeIutHi/8nm+4h3cJXuPqxYUMGz2xwYmBdiaMyyZey4/ill9BfVCEz2NiTOpfzbDBcU6sr9h
rJwHBReGGMQPmBoZkDeH+006drxF1PqlFzs2VJNkwJIJXATdOUmh4S92f0S+MKEKOnhDtNkfFLQW
kTJmiJpAIyBBy2EIww6frF5qjw/GhV9LM4Sf8eL2+Y9nT9q6W5xW3SM/igXDVVEPAvD5Axl5Fbyf
niTdbJhnUZRj6E5Qy3jTRTMDUw9dLrCubCuvt4CamKpoYYzWIFbUm+Xyp3QwcxqXUkRPSCvezg97
qJflNhPEvfXZaGJ61Uq2LU/Ylo6oTUsyW0YiQkX2/K83fniTtY4Fyt4RSKaB0mJfJXed3RmU5cAg
gdUmQyY9T1KkEfCbNO4HpuSqys2nP5QL1svNlenQJjvLOQXKzBdpjTMX8VJawzH4f6Zvx6MoZY84
Zn49UktqjxJ0YTskZFsFgqOunTZqKvTg8i41TCV5ehDxdirBZETtHG7tFeSran4iL+yQAf6v+W8V
aw9knHGQ2eSUNb2AWz2laTOatDXH0oyr60uwa0GMhtYn3cr2zgkFd6zOACi4NFLsMV0PU8NobQ64
b82Wf5hjqcaqRhJYtBqBk/tERsYPnZLWC4qp3g8yjVVIq2Ax4g3Xo+7EE9mQLGXTCWSK1d4DYRr2
+wT750VrNLacRBqkmNgARPBwahBnQffDfW1LrH0JoqaYOML97aXtwmZK0THhmsbpVeHavpqETMkb
/CXbjKlLzsv3uiAjixTyIaKzWcReaho9FkQTdedamKvWlEMg2VX0dnjJCdaL+uD7TViAIwzntYXD
lX87UkTgdATS5+c/YYoTLDGB4u3qy0rYBXTK/I+qQU3w8lX/3PWKSRL75l60dYnoGr3M4Co8Ko6p
bRzyN1OViuQp38Qo71RC5d1MqzZOp6/G73/znPCZ2AbrnBXKTtOf9BI+Vwl0OSskNQ+Av3pEVPYA
criep0l1gr3wknYFhjCPrMyweP+M1VdEnyNPPRHXKl9UC86zm0OSRSMDm4HWv1PAxHYGHnFCtaYU
9VMEyBp4oxGDKeZ/duGRWeSdHyGlHyHmcOG7JuIJWV/dFuxGhWtYuXmyzdgYLXK4sIDyK1ZVKt1M
f9Nrh6DjeKPjGeBLFIPMajfrjcdn9IYh1zwefo2p5Au3dPXUcwid9YP+JEJZ+wYR+NgKFFHbo3hh
MU5U4Gu8EOuN21IiaafXh55BfGhrbiaEzdgNrLoa7vcuod55HjMnBm719FG1KE0Otrm7zvbyubnE
tMRd4ZvM+wTC1pJ/fIZQECumB4PuuK9Rg3clDzhtaLuqnCC/LQuvAcgHqwYBxmbEK23SgXSgZEe8
1d5l2oZ/K9OmfVBj68vH+Hdx9/f2ZLEg31XwTCx7izICYNSeB6CS/7k6NBUV19JYJq0236PQW2qH
yYj0HkrUFTl2G6Ipp+hFwUkF3KuoM1yfCvajSZZUc1q/GsQws02n9tBzQyaT5k3zym+X5Xo6sRTk
YhP/Z6LH/gQJNK2tRN4deeUum/FpfDY/hbZZP1nU906i4+9QQugaSynXKXED8vpB2qM7E/Qe6XJF
D/ZYHU91xD4rSlQvR5BsnwAljYC8wWlR3u6UZOC1hPOtLDtX6O2pIWMLVmCiIwxXTkQ3dG3bNqxv
gpf9lNpKL967PrZwPcP/7psZian7laozBHAG6Co2Bk4FOCbpuF+7IXoEcCa52WQQpDgWGCS726ua
HJtUtDNYKTYt3ZI2ebFrWgKjU9JcuwhCe9i44H4qIeOQ9F750Gd3OXPChWzKnysvl2Ye7CVu9syU
p8HJqxfARnI3MOraSAAMaCnC2Sy74SOgsmGUT7Z5U9lZ7ugGZzJ10ZYT76xqySR+cTDfGTGX1bFt
sXP1Q0mB/PmxLLjq8UK3pEvrSk8Xzg/e4a0IHG9+IwLX2pN6VHUZc30A6mwSpESRhG95Mq99e858
9ZW1iMdZSsnx6n/xhCpcIfOc1wXLAuBC6BqZQDNWliXuEPEZPET61/JUbZ+JVgJX7/wforch2Cha
XnyH/0Ymc/RhxcGhsrXSEA4nO7oIQS3p85jFufWm7Jt6XLNAWwjQVldZydxmtqYjzC/cuq/ZBUj3
DoInZt3GPBeCGxeFuRA7SEunGhnwoJWRl1n8JFkSODVM6Enfur6CFswpPq2LAs8j1dmeNUev8sl0
sTwsAM53t3yzTHB+A2TJg2mLmy3La3tkNmbkDa1ITmWjGLWlIXmkwifjT4asrBOOBUCPYlNk9jp8
StEYEf+Sv+gQdeO/K1pCDsI1B04HnjxspVLDWrThOaW0uSH4+ftmD/pJx0AyLr2vmPD8ySU0koO2
xl3ktRkJBT2BKYUMLYn/uM0gfsNUTUi1XRB1kvWTkQlXu3izdWS116CuoqdeEJT47v4cIxnKLiF2
GmqE+kRxDIEKorw+IfdNXkD3KK7/MII1bB2WwmTVR2K0sLTOIlRosVSFeZlQafYdZHS5SAJktaqu
No/nEH+fGY2rANpt1bR2Q8sQ42xScUuPEuJ4Zq4f84EUUajl9a73EAKAXCIZzcn+EXn/IrAny452
hbCPbSIQ/HdTyLry8d0UXp5OY+uLUvzcqtWg5EeATFYy+rxaQcxca5WT9mdVL0H1+IzFa9LiqeQA
PRLAbjpFh7RR+ukTwaAPllTWBYEJiVpLUIP0kQ+FT5EAGOvwITa2e8OkMntYZfVlHuI1SeWfJi5R
4gQRiBJB38FLR6vA8Vf9AArLPNzLH9M+8LBGuboEEtpbUl9vBOxL7HWN8lrpchiZw2NWvpL7FvSM
4VgwH7t+l5dDJ/CVzrgaB0990LSPL/72LOTXfT7BMhvaUf4PIt3jCbj6seMQ1eMkU1Ho11YEQ4ul
3Xa9I2HBJgpwtKxx39gWIYxjG9qUspM2pvQ9U8A5Jbx2Pd3TzVSQo/S0aWipFk/DWTHG/iXrKRxM
nZny8P5L3qHwLU02OkE0mvmDBhpCwofIUDU0AE9J6aNARkp0TLUxF7Z/ctWycgAEJn+Udm5ZK3Sd
LIW8Kxi5zRt4XVyq7UQhZ4KeW+7WZj+5g+uv1ofJAKeppVCjlU9YD2luFCcQrx9Tdwx9oT0E6KIQ
W3gtM0M2zSu3oIAQSj5H84Dz6INUdFxOTeb6VqZ2faoIRbpypq4KNPuGrqCrmSHuMz0fgAbXOcbb
99Y0U8nQ3QyUMUHK8tw5hm0x3rlg0PANhi5W/xRSP0INAh8n03tVfjWng00TYf36bEfwRDkThpUV
yAnM++8w4Mc/c5ntOUz91vQO0k7hevOQXBC4FzxJAvzf/fahFoGKYC9Nom7DCKpBmQlRRERHJ1S4
ufg6cd7fxfhsaIT7Wdup8oMCVoILTwLI9LhqTWXrwq9KvBYYFHvD7QQhaFtlUi9L2LsoOn4xjEOR
jQLKb4SYBDQZk75Bq4Bt4Ht9/uO0lltRMaesJl6Wer62rnHj7JE6d7lBFDoZWx7c8Cj1Gvbjk+ZQ
IfasQdm4t4O497p8WIw9rftCrSc58XOvpS7oMtC+vZ2jTj/McU69pz5o0gjnvQLKscIjiXVqhv6D
LjwgTJv4pqM31rnfxKC85JFraGqBjr51WcNANWjZiwX2i7Jw+Y17cXfPTGnoCY1/six74lu+Cucq
e3Mpi+JGTOf82q2RvGLrAWv3ehxGjz4trjz8bgHBkXkCcAzDpDdnLBKqkdoHpnUeVUcOIMJxpiPM
XW+nliu/7KTdDR74dgrbbrnTJlyU7NqLSuDPcQWdsdeohgBFysF+u61PCcQjTCFu33dWnPyPc4dS
AWWhXly9NFne84Cl3pVa8xo/aVwjSJ+Hqn8KVYU0GTs0HKDYkdv8tWupsHpAKJI4y/NukTp6wsYc
/+2LTulX936CxOSTJhOj3qlaB56g0SvqUtsc5jvcbEuck0Kndgp1J6NEXDiA+Rj2pT6OMyvUGNPv
TPmg1lTHV2FVNzaF6L1TtPif5XB2Pmi/ulpcQ8lz8tQ+Goo0Iy5R+jGOGnKCgxMXDDYy/xL1OyXR
vV6Bce4Lx7Grg9uL3hKjPs9VqXCubLkd2wsL3hB5knXIzQAzj0bLqPtPf03wYi9Q7l2+IrAlBGvK
FxW+oomgIIBtvLOwLUpxOpwXz887uS08RzcOvmIeFnaGyYc9ZQmaeZxewL4aD6VmbssrQJ++FmzL
YcxT/PknYGr/3G7daEIXnMUbx/LKZ8HBJA3bhfU97SI7oZcuGUa/wyo1XPgJaD453lJBF1nNjG+u
uCOrIAQnq7ygneWAnO2BzywQhj5FRMm6SZAX6SEwG31aJoaYfCCzxOFvayKLHZBSZZXWdPf06gap
2jaQbX0YODzvFDNzFHkWTByOlmEzgCsri9qpmH3kVWTyoGtDc63vmomFsqQ9qtc/+3mJeAy3F9do
bbx6Erex5MHlJ41Sl0Mr/b81tQSOymNZS9Zw2XR74meiGdr3+c6uX5c1SQ53E7DCw9S2el8pnkOT
WCRirQq9m/zWX81C2AxZyjWfnygEdQR//wAJNjTZSHdOmODiXMQlQUihUD6C1Vkm7TA6wodUKbbl
mJSMcrVmDVTX3Mv+Kg8mg8mFwLwgRkyhCKnRYiDwV0HHmcbteKlnLpWUgO0C3cuRupgflWMUL4Yu
vBv8RKBD4CQpwOWArqrCNevxjHKg9/1L20mlLuJKULIUmu6xHfZCXNZadhC7MCzlDPNeMXw1YFkd
F3KPv/xS/swQNQLSeqZ0sHZ+ARvRTJEHVJWtnu5PcTEn7Ge/TC0wRFsN8lZBAJMAgxQ5H3wugZHC
PTWF/RtBOrcUTo+TS48CCJhYPdc4zvLFmKV1c/9LRxQtPbe27K06nZ9zLpNrsTSh49SUphkGsR+0
M7rBz5XJmykAErSGytJKLN01vGpFbk9EKAM8K4nA5VteG6U6uoVq/5ODgeKdY2fJVcIz7d0eVZpl
3PAFVrgwz1ttXKml3zXoi7y/EqSPj4FQdgl6/OFe6qKfj7J6ikn6WMs8mxqeGg7P9hOuwp9Up0S5
NmrYy70HBzgW/I3cerCZdVO5rV3k3B6c55UobQDdcxWcQ8tKexth1k8X2Fme1SoQRuVoAkkP0n3m
/+qH5rau67RrVVlNvQ2Jm3ytdFtTNrzAF7HokZLzN4KmMr6nEhl9C/pT8CoU2o+q2Pjp4bDYcdpI
TQzW6OlffQAfjDWq5MqtqvqkFPPguZmAvpjyLZNqNoDsDiTHdm0rgOg7rCd5VEUKFklPIQ4vF5Z4
spMcWqxW6PbOcn1AoSQJrDWEV9nmSQmrCe/9tjs7itaNBkLPup3URuL8nqRsNooKYSewWXDikRDW
5YcBUf6hvwq0HLI7VXbR7PnTgwptnBiKnV9lplnO4nobXyT2/V3kHoJFpfJ/cuA327fMRfDhKWrW
SAkx9oMBztb5eDTdn5JBdCQ0kxPfKt+UhjvWc1UedOwZVcVcGn0zWrITRXPqrkfPWHaJZPImY4BO
rHnX2EZKp+HRCptUutnhIMqrlqD8jmaKmIjfHpkBHjEYX6nfYfVLtFkIvqVRmfneiQZ61Si57qwh
Z2q8RALRNhP1KPV9r8uPHMu+QrC4mTpvF/QnTA+9xnowzlZstx7JxBJ3FAz8PL8t4I5wM8MB1ZN9
WJsDi5GmLQ5brIkaTPiU3B2hrG7ZxWrxRNdfalpl0yE5Cktwu//Indi8/pMFvWYk5sDhg6U7gn/l
CvTt29PgaN6bhu77QEbr8kqW+kq2PSYL250+Xm24Iwtke46jZg9+WW6Kv/H7sRkyGG0y+h9H8RLU
WWRBc2med+xZYs5qNX4siL6hRD5uNsw7XOoDmGC1BQddskq/0Cw/5fAWSswceWDx5LcklX+opJcf
nZFowC0AArvyuLBvrjl0leQhtEBXnMSKx837q76tTCVOSbEBZyRpRiihW+N1PC8PdAJKW2g3F4v4
2Pw+kjdd/IVpU3x0sSnS+BrHvq2vwagqidz9Ni/jC21rTjN8gcE5Wj4sfAsSe07m64qF0RntOYQI
on+gyrTn1PlRBY/f+2Terk5VTQp2anCisfeXXR/vx6slxjZM9ocoxtfHPUP8VFnG2DWvt+tjRdEw
dUdeOUIee1jsA0NejiK5hxBP5L60eetkFOII7ipfeAef9RQoxQnPCZr60r04tqbWTMAjWycHbA+Q
+lg5G+xwXwJjF3/9Q0TTspMS7RBJlwIdzJ7xVkX5rKvIDL+8+jnZiIe6lQcBxS9artLF/LtqHTKn
CLVNk++xKtRRiyRIOzjEf5L5AdnKOSkLdZWQUKDU25KKbJ4YYCFRPJbh75aIv59zkpQDI3byTsc5
qXD8FpYD3yZK5+1ClLaOZICvykQufJgP/j8QhZkksN4JTIdv5q4/HbDP5s2AI154UEv0TonNLMN+
WL8a5bnZW/JYtMmh0rqgbv91CvsBGllvw168FAgr1Wy23cJwQiwWj1EflA2Bt4f+kpgYFqNEk0eO
kB7QWqBy2KjuEcT7MJyKO0Qr3Ik8k88VVWsik032st+oaTzj7C4QG/ayt/SE9diBHxFNv7xUBgJD
Uf6Q/kf6dVCem7RbgtZEPcgT7xRJLyiOYUdLPUQOP7X5tOc4kMkPbHhJ8UHnD+fuWVjSFfbPSy4l
G0ZBcr2f6ZT0bSwAAmEH5SyYMOEQSi9UrjLaP/6fxYrvIaq39885KruT1IR7InCEsmADvyYgMGNa
xpybRWtNSylfTTO7qnSwVFCiHb5rGNlr3qlSc6CQDrVYPDsy4+v37a4q6P6thjNjyd3xHuYxEJgv
74o5tZF7Hg36vrCFSAOONlZc3YGjBFSnQnxqOX6F+FS3Y7FaIdd3cFDl7MpC0U7Q3L0bmNWzCnn0
Vcno7oeW2AJ+Et7LXFoRKFcyXNV70kia6EPwpTd2YpXL6iYgltxB1/fWgQPTgaUWSoW/zlO77UxR
Gz3ZX6OMARJ4SLfW+LriD5EEqMlakBy3g6E4ZVc2tPc9eMf8hAk25bnKmL6xUI7Y7lgyi5D1Ziz4
PKI+LU5bgi9GMM+mne1rV2DkHSimpAMU3n/A7x9ERfN1uodXlXlyR4+vi7krPuDqZo8KS4nUU5pM
1JJJw8ZsbGw4wyi2ZL14hh+4oo/8ORaG0duqxZQr2fSus9+gavx1FexdUEUDTj+qErUDMtABV6MS
LgHa0hEcKLKSf9sgJYaCMNHbJBlKOJklUOgM6l4+p8VkGyJI7PC80UHk2W9D1VKUM0/HYMkxodNy
hpwMQV4EcRpYTAL8fYQVQkj/PTZ+RpRCk7ZnEJPW3HKEyYLw5UU5AUjkZopUvSq4iTol5lw5tAio
7pH77ozaL/KuRydfnjSrtXEht+iMaOCwqoBzMQsGCH0yeU7G5cMFKGz2mWywp7eR24OsNoA6nkm8
6x4lWikOOkdwRqYCTygYq4SqVBvHNAcLx6fUuyg8EnstRbN0ZuRr5YeNOpBoTepU8IsEEimNG7rB
iUW0wqJkUnHFGzqdbPBNZuCaRmAjuoNMES+PmuSkl6pHA/KOi3582XQnVic2HUzkoBRPhCBdAglI
+cHgsNjCrJrpAw75nHMDNYDzaaroNb8I89P7S4AT9mJMbjEbnI5XEypc/zGzlJJ0w5leDfdbdfij
6vWAMv3KmNqKMwP7T3bb/K9sArlHuFLAxRElEL5FeQ4Wain0SqEyEhlwP5Fq9YZZaYAsAwzbE3cp
okhhiIlwVN9mYj3Vt5WPC4HX5qEjz2/+02toCsbjf9rlGG9ikKZ4K6nJuIgSNu5n5/eR6SAIM4WX
TSsONy/m15NDStqkhFDJWlqClzICQH9UW38niU5IkzFTiZjTFfx3qsnunsqKwWx2Xnj1UWINyq6c
tMLAbBIGAFrH+4z94Nx3zywI+kUCXubTsIXZEgVqpXwtczVem15Q76mFncBO4zIWRcMs4WR0IYB6
TOo+yR5stcjjWpfB2kLHcb8zeTZGy7kUjAva1DfGUX6SJahjCNo8hOwL/jhdydwoodbgzVDMqZ0H
2aocvq9Mvo1RrEeJfjr0z+ZcGvkLekdTe+WYrpd6gQz6OWxhfom4VrWQgOVE0iOEsP0lZ6iFzewb
dxPhDwM4X29vd3S92wVVwk1i6mmkQYIISXH7FFKzg8AAPOsO6/bTTmx/JY6fc9+ZMX4gc4nAvCDf
B48M1VdB1x3rgcp6KlF+jwz5WHZus5a+vConfL9KwdJUFjVT6GBVjCPS3fRsb24L0yxq7xETh6RI
uPdpiBVvldp37Ez5mfiIAhUYfYBFJ9c8W51okgfbGaKOZ8W3isiqfDR1J0LFSyNOR95GK6wbb4+C
Pz2vvafRpLfNEhpYRirnbmUf5fsUyYOXO9vZOLLrgKxIhjEIfvYe9nKLWnhiteKGh3erdbz7LBtY
UaHHrpO06tbwfTaBnMv29WjA+lDPRqiK2PZ3SJvYlmC4PBkHCLzdyTTwTeGANrN9D19BnkgrobPE
TxIfXXrhoepI/Ru+aSp3KTPjee72/f66HzC1OiiTNrJzRRnIYzEiNtUslrgotlBurApbNgse0Wpk
8lXMdBnd1/6yg7uejUeyqTwLnNzG8vF1BIH2TPJgrY2AsdOk28XPdXrA8ObQO1jecjaZY83bgw+W
Jxzqxn52i8DDe7jRg7+hNDKpjGQGBCt2/fpcG9d8j9fRx2/qMns0q2wVGNp73yQuduXcf9Cx2/Gj
OsKJziBR1XTeanAC27tGmDYUwoW9D8GzN9A1bC7ZKqIk+1k71t0XixTcUDbvNlIZbW7EjqGEobxI
A1DOqwY/5MW3nQumpE7htSPn0sYw3S79IqCbop+a4TElIpuJSEFhdQvqN938eRt6smUXqsKswHXY
dQyg/PVZSVHGHiaZPcHtgIPJcQ/EKUIBBE5BINKWA7j2hO18B6KoCUSOEj6cVxJo+YAdhywdEYye
Jq1LBru85AgLgPSQ48kHFYdp4J5I0nyDmm3hH7/PaLeHDCj77l2/D11ExvYLU0IysvqB1NCt6A59
tEejyU2Gu0z3FWbQRF6pawL/nnDwWQBRqyyo5fiSJI2hYML1qxe4rbhopcSmXlGRx/PGeGFdhqg2
ORF0qmoCv7CMvcP185GjYZzNQAViR+zUmf9Ilx7masFbdyR/q3CXF6MM9WZkpZqy/LAhFmnpA/89
tZQsRn8FcphRkRDTUM7xPorbGiL5JJK7loAm7DjjY2xegLAXDJ1ozgAs1vaEE9Hd+N2pnkbDU+aT
Gf1muTTvNvWSt21oIUQMHjz2ENp5C8x4ZQpsFeXD1U8Q2XdgiB5ef2VOlpAnZkHo5lVoV8/NnYaK
gtGjne15P6998dnLHqpMJY3DWOpp25wkoRrkGi4yI6fpi3wdJ3GSciKkw7Ltj2F6Wp0vvRgHJWZh
hPtXYUHUYWP2+ZMY+C+hV+Ta5c2j/3Y01guhj4L7lpKt5C6JX4iXmi2WQI5JzezNEEILJxtWE49a
/+TJMeCuKWq/g2aj9UX7ve5gKJC9Dzu+F0pwwGBSiv7gmIWs5m3xdb5CRXEhqxRq2AakM3h7mPdY
fbh91mxy+NsjzQZyuS9ncm/6VJ+1NHMbYNKd4ZncZCC/MaDjQNoPMAEOG7v3KweOThwzmZ6eGQla
9q2CQwxfFNx+dI9AYLrCOe4rOCazqlaZ611D9mAhMwiV0v6AIEIIII/gpDx7G8dKxWZlN18vYGtb
rFm3etjATR8KF9JFLsy/S/NvuvaEn+fklyewJ31R1lA2UjmjnTBKJFMBUYPTX+94TDqgPr5g0oqM
qJiBs9pO9tiekbc8uR7A0Car2QUUCbnWhK2NbZwKMd6pnRRLSlPLKdgQPKpCMuT866TuOYvBqAkk
TVatABhQd8WoImJEgL6TcpngN64qQPO8+/4fUpovG2/G85VmwYubYwH4GOdbnwWt0WkgvoARqZDu
JczqEDgFlkLdb8qs02LkaGyJHXCS8dcKOl4TkTUpTZpgJdLD6pBPiKhXPcB2O+nD1eOc24nKruDZ
coUBSftb6pT56dgvGX9TeHebBHvQwRxgRRd1CFd2BGPOB9nb06wxQbwLHwT3OImTVHt7ahVEKN1D
f0y+qg/GRvr1m6v46vReQpaCMlgyWaQ01LiuGc+dAXElPWTpZCsoUJkWtqvAfhANwDiOzuawNA8b
f/7PrWLfTkIny4/k3o8jrk8jlY8KOBV1fb4hlu9JpHqZqIdZ2ldokj+uOrVgwDSGv+oWCpRsTxCB
ZwZepiMo0xrQwrvs+34uATwAgS3hbBErBJW1b0++BZ03+gz8LVbrz5mf8J2fegH5He6legHh5t8H
naZ27cCfQEvV6XdH15kdRYg4a+73zhlfO00QS2Jvme9nYDKZ/9P0SNtI/bmApugtrvZ858XN+DfJ
fg+WQtZpsebw7Ni+3ehPaBh4d74euHO6J+QTewC7X9ntYZwQEKowgiRwGQwsIwQFpTsExYPJVPxQ
27rKvLiwp/+W3rSu1JbmE4aipoySBIyepUIolUBzo4r+STovF4ZP+/L4UirM3vBxfkDWhnt37A5K
dLjHIAxT+0nuKhaXUkVADzSn8e3XbQVCtpR7I++BHLy5CCGFXIY8RuMa7yzYKFEhAchNo0BBBq7/
96GR53Pm67eXHPHpAro1L1nzIZDgs1mdOfw2mM06iibk2OYM5Nv8XUu/xxTqb+1DXuUHHc50eYUD
gYlcrIc530F/5MZAzgv88U+ozR+w6HwB0iX1oL3sAiPzxAPRRBhrI6N80VRbcFfoCCb7XgqtpRgo
lB+WgBUcV90yzykc3JPbXz0eNfYs6wPYxUHpwzKr3weg9JoPcEavMz1pQA3a4a4nv/QUDMJ9cX8X
4Dpi4OebExJSDvJuvEwvBE5F9HZbdKSAyEVLTyFEwWzXDWkx3JMeqW6Rd7iJb+0pxg+U8w2qlNVw
iJsFwhB1H+ZK6PJIg7aBYO7/W5hZuOmP1clRxaWSzfoqbE3V58wj9TN0apY5HmMM/pLogJ/Qwm4P
WjejihFg3RU7/Lu/jQS7lKsq7nmbPDsvpfqCcgpinBZYcoNDePoF1J0ep+5Nj1bIOjDuUgFlRtKo
1emSEs1XfP0ECAba5bQJqprlM63CCWZI6Uo9QfrU9zYJMx3CVNhG8695SvtdErHGiw6u29rtu9p2
b2i339pYo9jDpRTylA3dYmmBmEvCscsJqVfJaO/vt48LXhvDFzafW9wWh4e7UBC40dEFprIVzp9o
Mh41vk4arUVhmbGv4vcjDWqJmVUjOvHYHt+Ur/y6Utb7Ar22mgbgPGQtHVXccVFiF+tkm7uattzo
YZYfe2Zy22+/bko7TA0C2e6cwuHuE4u5w7O4A4aonADpeOnJphBEs28QrIstEGIHTVc1auJYtkfl
8YSy3bOlNdP971GHd3/cCqEa3/ePyeHytCohhCAmsfKc2DzG89VGr4yh1X0gMMinPBmHzAEH5rpc
widc5YQIVb9ksrCSDw2mx2fZ5rboSIoJz38p6yHFGAbjPXh5py/txUndDW8YpOVrXw40TAteuJbE
GPhS3ZdNO/GkF0KZhKp3IwKLKXI/giUmwa48Z3iLXGtxvLvogVE403/3IaCj0Cozf0gkkdhWoRWy
RlpoJCmnM/kf62ikdZgGlwC8w0lWx7ukd440jV9c4DAyIxOmPvPI+cOhl46DXHxwo7lRQoo/3O1B
WFA+Cg9gXTi8EVCqtrJ6H2CeJ7OFKOLX3CyjeTRUZet32LmdIH6gIt/wyDFryaLKncFuqMFZ0b5e
/F6x3Kv5AN5Av7ai8+HZBPjfAETGHK/6Z22YTjUK/LDipTZW7kCPicr8FBnc02qErzwut8XnviWs
SDeeiCy3UCItqDpetGMf1+c7Oe2S+ld41EEYogoHYkalAkX3lBA1psxXY9asjBmLaLidXDXeIdnA
yAnvM5o/Sdw1IT/F6JB0yhZUrevKxLNqWfsG1rCo6sMU4N21DypJd06WTSAnXbk401Mrqb9gF4NA
A+t07xpf1xfXXvoEcbpccoOA4KGQ0HdimRfPJqrTSFXiGCL3Jd+g9/NVKrB3fgcGw0YuqBmMf6GO
eSGHBZr3gXLJITSgZlaAx9UXmfuM4gfGqw060SjqzKd7uk1g/cQayyYViaalAjnDfzsyGW/AosFm
U4nqCw6XsIIfz58wDTd+uH2OzANPz1XLa2CLkvanFzkUHBa+w6E8m1M3GhSfewP923t4KUMK7JMr
J/9uk/zcu4hQiuLQs1juR5PROEGLwJV5sA2MAIISaFeVb9K3QBvV/Kvc778I5Fcx47WctAs92DDO
Y3sQdkGhiquI1RBmUDAIhaJAAGe3jQ1u1oKycUFFM+/YvaWZisO9CMoK9eEpJbsEPRTn3AnLahdA
svYWWmISk0ggak30PsXBm79a6obSeVS8UqFGWeLKKHNyowvAHVnw6cY7Xo/WZDbuicWztqjvq9p+
EpDe7fgjnAxQhipJcnkhKUb+xpngY/rCST2PD3APguVtvSzJXddYNrYocXiBVWX9h1ZyKgbESJAC
BXYQFuDD+5H96lLnMdf1w0czmsbfKNZf7tuKYCJQaqNwSO+Cw+QsXw2cDUOOPLnN0+okQAG3AVjz
liUUGsbQMU7L6fzjGtmgVU07xYYUgF/MKQevrR1eH6/hGNQyFI2QiBXJvKiS7b1y5nBUNJHcrg/M
D8qEMwB90kiSTwUSQNwQ+vzZ/HqVUw/pyoU/7hkp2u9xgs6QrHu4BUoVf6AtmRo5voG9DfInoXj2
7FlB236+SyHu1MYORQk9KlsOLU4vfHM827taksUmRlnfQ+MM1rXcO8mtBWieiIsKG/XpH/Hmuas8
aojvzx/UvUxPTdbhT0gdjFsdoHHTbpHQXDkT0cMAtoVslxdi1xPyqpF3gCuHfjrXHFcmBR3SwkzP
585ZLyb6x44Ek825mplCcNW27jQ9De+whJtlJ4ZX17Xfqe/SEsIiZOp8+mgS/1a8o0wEezksutns
AhTeMOfbuae0qpdrPqqyF9mMhXmcGH2BfWSmOZN8e7LEF8VhmANbhol5n3g9e9tyzVdeqgGyOFT5
zBUnYfGvZDdQ8IS7noyc0nzhgsTO5odV6sVYt1lm5SwvP2/ZmF2kEfgrm5TDfSk9ZtTzJ9tbYbCT
Gvze/n6l2qG38xsWxVDiMixXzuwvlOAtSwiprZLoyVvru2QUFtf3DQBB/FLRqaM6FQLHmeiRPeUV
uC5Jf6kDAZYLiqjqr1Xb6J0nkNBYSGDt4WInrVep7vHnhbAyRlov8/SAj3AChmVnd5fo0NpbtYC0
SxD3hL2xKh3pAOq4aMmT5Voc+kbY/oVGdLgD1YBaRRpU1Uj4ax7HeFc06fP6znELolmazHuvTj+l
btF15FewxhGMYXd7ARbxqO2pfAedTfQSCaQjS+A+LX9AXyVjhLCfz2mQW2ZpEmGzbUkEMrF+TjH5
hFvVz4JhT27kUUMj+vhKWsAv714/6e47gi1Jhqj9rdLVhLSrehl9DO3Dj1jMJS9VrIln9ewIVBXR
wRxKABl2zbUxAuN6L9cQBM5xjugXnIXdrM3BnttBAM3kGx1mKFwY4mKnaKTumCAQM7dtHGHUoc58
CRYw7bdifC08fpLXqBG18j4aUVFw/9JpCG/BkSDghN2hcVXyLSoln7JbP7IOf3JWRkNc185sYB9G
KOgL0DWxElXbqb0+FfcTrdusx6ZFv3wYltOS8CZ7U5mfkKnHmKVlc+6xa2ArVh5T7h78fYM8TFji
aYh6Wy6yRmufOMFTsrmZ0GCCwd0z13PCZ0+jZs5svTN49IPL3aEc2bGggt9zulAiEaI1YEFgFeRr
z1c0EIgQlufRlKtpKz9NTk9AkyuJrG/4okmlwwwVLM5RzN2za0Lo5DlDCvT1klBo2JJ51ennxLzF
p46NZUe3lHI/Vjc7niY1mogCIt5ndY+NWLfw1zMsfRq5ISa6+3/K3kD1sGnbW42J2xEVpEg3/6oU
nP4bfdHxLBpqYQuF+CRfGoanXu8WAWdeICH9agMLLhcxWEyCrB6m6ads6oNBYNfllMlo7KQYnnqe
8kkgGXG6cOBwaJ5ViK1wjuZm+h47j9dx0IdvO0qJ1WNpRa00UWFZFXAkfLSqhDD5AuYNSsPIT/Qq
0G8c12hl2NAK9ApV3kL5AZJGgfFZdCRJPmGT88c6wPyuiWSODlwmY8EsrSbhYAKfeTaBWpzH8QbN
vKPij5tUPI+87uoraUk4ik/XBVIJIVKCK4V/XAS/qYSV1fCZ4OVGDAQCJ9RznmWg819XNGm6AJag
DMpzHmOlt7ZeTpspf8XYAfcTppoOxf8M5JUXvnpRkOFcsN2qQ19G9RZFT9uzQA19WPLN6CvWHwWz
dRnyi4Ay03zFX9fuOXxsPFs+o+ydtkJyuZKhGHehjq6gD3pxrAYE3+IhEKST0736LT+rqBlbA3AE
JbgXADO2I9M1DffdsOhWtSGRiWqYWlAOm4yCcDIu5ScDD/PLAL+e41SyoXlrQUDYONzWwWIFOYNA
Nb60L0strapJSuinvnl4c12heDAo6N8shVXevI2pIALqqD/lFO2RNblDn/g7fMwbz2ts41sEDUEs
CWbWNeQeVoUyUrvf2EFxM5z/IOB43a2ALafITfaZXQdgdo8IXWffQ29J2X9H4kgWJXoU4P+yKG+l
2aA7Y4F6jTOSdbtuL1MH9g2gZ+nN7WkiRvfWUs2q082ypM1rn8ld1doG6XTq4mgWkHwY9KonsOvS
5Ba02s80WU8U1Fq6lqX6EGWgXryQ6Mp/TYRT8ZeRJxGxXL2OlOCmfMaa4nLWkpDcOesoLEETx2dV
XJ3rBAPADFBez2RS2Vs3gk6MGOH4O3/N077a81ZocIuqOWai+KZGoUxzXh/79rovu2azlXpRmP/S
yFJ7y4GyqN32E6PpX2bew8hDXJRU3w2/HCtRVcwewcSpGzw7eVYtF/Im3hjJrL2dvnX8P/tizthP
lvUGnNj8He2T6phgSbDMtF4huLhoR61kjRROPMA4W9CFUaQ7Vz3hq6dgjCwjBofBso5sr8Z4ql2g
c1R/uXF0NQPjLuV2ymUdPZu0hvJZtHst/0Ux8vaPsDnNqdB3jy5zyRXc/pD/Ix2wB8tvY6x7lMd5
0Z98hbOor4qkVah/xJ9QD5oSdD9cP674SVPTIt2SjraagLKVlCK2zb/r+3CgiMPHW65sQJH9Lojr
er++oxi0uVy1xg4z9g4VJvtgk7kbX8vIZMzJOLGJJO3U6IqsSDQZs4UorGBqOhZxQP5+aSUIie0o
ajDtVej8bG8tuAd/wXlaxkPvoERKljk8lS7EjSMCXLktQRmNdBP78lKjuT4Mvb9R7l7voJeIIbPy
90lQY4WhZqLPThdLd7iCAzpcB6NG74BAHvIj5luS+vly4xtU0zX+cY4nNFDpjwlhpKrzV7NcAVE4
F8CuYFgIn80xwQaATIHchnyUcvvoxLZXEMha3wAoUIDkvwiyimljRvvfivIx6tefGY48iSK8tzld
qCjowtJokDzwbAGkXkC7VcvXu8pnhB1PlfYgyPRf++Sg8/czeYhX/O0ICojLCzB+Cut38hOibWQh
tM0+dtasMfvxw7IoejS2Zzj1qbIA3snaqgdFRqQj8dIFRCqCQoW2bt/Iij1x7+0ciwbcZozkl+No
mx5GZOuFtMVQLATbWN5D/OU5whhJQl4p58tzOfMf6duWGsLR84i21iG/YntMLWB4cimHyjlKwAiy
2UUmQiPZTcVXkDGbFdGQyyaHzPsSPbaSWcdBBOggHuSG+pOWWmNjTplMyRa0YhwN9pT9poMmnloE
ABWwy6WluTXiuiUuVA4El9GX1zsheeAZLFYfMT2iew4meX2C3oX/doW94FGEgk7LUSo1NSsWVNby
3emuNqtsKqBxsGS6PSJSvWVLazVo5NvWBvcycAyBzLfzF5VvGVR+l9lU6jqauh7EOVzvJNiW95n6
RIQ5m/VbCRHo8qVMhTc0B8a4JIhES1ElI+1r7ZFCCK7P7kYg+lwPGI9qeQSoBXflssOzOVjMuwcn
sTmhupcaNsrpvRYWDbAqz3HD0Bw7wQS6fA1d7MPkSltdAm+ONJspWWS1YqAo9PI1XQfr329CPTPb
OXkc7YmeEShXOo3sOyhAWs5QCA+CYjYf4q5vJQ9oqsOHf/trFnr50wiu6XbN4398K6N3ookeVoSW
hNmPWdIPHOMQYFpoevkJCpEVoMHdwgEj3NRPkeFKLUV+stkAjFcmRkFOjXhB8v8z57aGV22skkvE
qIPG/IZBNIFdIOcYOxRtQA6fYcx4H0TzvQdHIrGYegCJZ1F8+IYkiBtWpzanmaAC9KWQAtKZBKUC
hM5zIBoOlDNGdIgKaBTlZY41+X0KjnQ4SZX5YyFiQHCNUj1WahRoVPOnqVSZMoHlVQR3yDLd5RHf
uirEWqpXp3k2evX0Nh2HwO56CGwO189zt5dnbeua4IEsCiqSbVFVBSW/oTZePaz8K3oUaF4UZDMC
rpZ6jDlUla5mn8WDfabhPk3RwvNG4l5vlNY9elhlkWr7FsR57WA3gsIwWc+qQiYNXwhBkic6drHd
nyko8KmPBKjhQoAiQ0vspmEqj1NeiADpWQr9eQMKtlLhCbfLhBNKTDP8uUimDqrAC881mIeD4T8U
BRs0fkJaWLcTBmcV/hGDDHqLfiLQkukadnieufOjrRUzCIZvMc0j852B9rY5pDbFtOne5uuXh5KZ
naUSyILAGFC9UwSaXCEgZtBJer4RUR3+oLoA9WdZU6+YUE2KdmcscOMw41ksomJUwZ7YbLWrbdRW
2NBRkBw6hqymWmytku64nAr39qunHy3ugvzZBpjyUWfK72brCtv7CAbRmCBHQHVOWHyhLCQYrJsT
QQ1Qum+pkXH9clyUCgjMwThXzmcqRANKK9B6VBQG7P5MWFuYCYmLUfTw5TrGSh1wtbmLUB9Sd/6t
prw7lO8qJ5HcVcv5eeTLkLLtiD9GaexoGzjWsRtJ4XSwcoCTY1HIjd4/xiwxWuurk2O+lWER3QPX
+dTinTa9X/x0M4TKcycahXs0QEXEowswZHbhuXrt4fgkP6qVw3GbG2xFZty1BS7NwgJvr1yPm09N
yBJ+9IYi9fqMTPV92AOq+iS+87bwnYUfTkJKdWua+FZ7U3Yaz1FB7ugmQToLwzBIHZh+fuVmxvvk
pDlBR/3kamTW45xotJt1djqbpVSTPJmVBvBVKnkS43ROHIFbzgxFRpkLDwlndsH/YSP+lUGB8bVY
k3yoDBxxzaZhb96/XQPOxT8bdOhkwpRmOgwoQqoRaWA3+R1Hltp4WmIb+Xrnu0S0w/UIVIrDp+tY
N7SFGdRmh+0/m7ohTRu85z0x3hFuk8QPhUbKNcoEKD4lsFtXp+TNnpU7pu3RVYwdnkwTLd5t6wvM
6PMpj6etEHuEYR813Xzog7A0FkYOWVOoHyWK8+BXMqq5COeYmysuBsfasMVTjQ8dybQLAtE59leG
e61HwylNtcT5Fj4ZShPvAUFBHbQGUgspD5d+2Z8FTr8R2MjMO036I5MNlQ/IIw+vDT8AdgwuYgJp
yWOSOhJvGQd11oMX4HlKr3Xc5hJqzP6KTbvOsjEeJwz97R5yKwGLdsl82IKZcymrf/dlfY6iY9LQ
tX6ebXoBKnF5Ig5+0gaZq1Rfs65CpgxsFBq4L0ELReBowzyQ4pQMwjXl2tFIQ8NFkQ7qLFl4A7Je
Uh3Pp0vQZGCOtxJuGDmEEu+8dFLyX6A85KMKMWRgtvO84GUM2fSRtuaGuN3EKR9j0boj67e2XHdE
O6AL3kqLjQtpHTSJpWCVceLiVx4f6Z2UZu0fouUzcJ4fdhCZqvV4xCEfjXdCUdpLRHbBncL+RUc7
lLCORlXhpJYD6pCiYNdUL2J0LzghEjSAXQJKfYLO/0v379ho/nzbhYrYj627pi1QeCtO9rMLfpmk
jpBa7ntSTzoQSsAgronVBl/9IKvNmIkNeNzn5ZElMsZ8gHFH2bVH0nhKds14pkN2ebnSsJFfnTFD
zuYRfM3xGKuoOS4MWV9ZqeT7UKzqCZVAw9N35bVJohElY39VohDq/jUDSlNl4IOIKy1Y7+IsrWrm
E8s1dswsBs/OQCWOgwsg5zT23GpsOCPm4fbMT8+6gSbm6mwn490/RHRDrZTmTOb5XKMWitQrliQU
ufBond7AZm6Xyf2NAXpW07g+qn/INzRAc01TJfBGDGTEIvo3ioYXUyLlV+XR2dkTMqH9RzcE7i8W
ADbuND1JlBwCWPhX8nbycVYp+Va1JEcLt8ELV/naJfMj9nH0fm+mz4M6+0yYgEP7Kln8BrG6c+ls
b/WlTywmZ5CFcnQ6WjyXZXRjmQOPtttD9Z/ffN1+E9uBcePgQ+7M2wfSValqxtx+7CbKHZTiwpuS
kabWCN+oX6WRa/Qps+WQCtHA70AlZV+KlE0sBbETu4kDNTC6FLo1v7UxpfqW/Tog0pZSx8JbOwn/
aIOoEZvt6lo4WxjicChc0ogcf3oD4yFdhAWXZGpRp4dMQaAQ8im4ilCZe5tcLTcx915+nuT9jjy7
WJ+6HEpVp51rnn2mSqkYa9U2l3JeV+szT/WRGh5p5J2Mz+AiIxCcPOKFnUldWFzjuYB5yeX8xedW
9FOQkOrDL05fRgTy4aKgZVmnpLSGMCByNhX42e1UK9OFFDdcAVnq65md8NX8P8Oa2OqarfIrOP+t
bScPLQVpWz19q5bnpHMVO3k5h6G3vX3uPP10m31Mbj0FwUqT5opzKEalapajfUClf6bWRIiHEmNu
TKKNLCl7IC2+AkwsVoeGscVzQ79uMBfIWLaKg8dGqyC4WGMmSA92/kjlX6Sw7al9kiEn0HEF1D/Z
bM+/5b1ED/VT1NsMWmFHFP4Uvng3cCBFStBMiHDj4O3+82WwOnqqgTGanvkeqPmJzqjqitSBSDzJ
p+eWzuVyh25moizlSs+kZv+vuYyOMX960O402PTbk++coH+pVPNR2mPERIgSs5AAr+N1YqmmsQmH
xXejUGJXUFyR/Ayvoi8UjYPVY9Ssky7v6smw5/rMMon5XeciIVsaI1Gaz3BHk/rLjuzF+rbV6c8m
myCHweQEcONsk8ffbNrd2xmEp1p8vWctDltRyQ6OnfIXun8RnpmaOp3WsDLLfAjpymZQKzX74I7o
ADciqu+bgj2zsA+izvtcwzb+RuuiZyQL5DaSTPzm/t9X/a/+sC0IZBPJaPEJGiAkHFekb/rm4jWq
RWOW0ez1QMP82SBFcReBgvyELASfDpSjWQnfK9/Lmr52t5DmyoaGQfT3CQBKH/pIaEdXfH9XvcDr
oYjZQeOslMZXZ+KqsDdw/0oJb2MOMqD2NmQe7KJE0QUn3AfJgTAYQ3NBb0YwVLFHGLyCNKMoL/Jh
6eTL2lDkx0iFbBOZ81YUhH+KMDl7pN/vV3LANZaDSn7tHOPngliM2c1gVh2Xbyo4hwhmCZFehrFs
HM9yZ/DLrhljk5fXLPLAIs0gXHHdqunevuNcn0heugli2u/UUXE7hvWzb4ZGq8URHDu8+pT+R1eE
k43u5Wz7oo/WPVBM45kor6MLERvngxTaJZRQi93Hh9l6mS7YoRv1fG5pqJof0RVjspS3+AHBYmWp
wX6P4fo7LmxBIPtUgwfeDf5IzZga2+2BGaudep/U8sqWU+b9kSQ5C6FU5lGhDdG9mNKMREPByqNw
rD+oY+oXeiHQ5Fwrtx/ono26WVS+c3JZf+tMFNunXc5YygbbevOk3SScuxMRJx7fLQDwsUOo3C13
bqIoqACqPfiVRDUKWj90cfK+LRDjORIqogXbk25a3t0FrkWocPQeosZxgcZ5Yknl6Ht1XTssLCKh
nEsopQrQwII8IPE0990Ib/fyQehIXf7dnvGPWmgtp6OPzdIVvLun04LsH/hEfmOJmkXY3deNInVv
SFif4vTn9K/yYcz3Bg30m6N01wtrQE8x+7QtY3/XsZJ4ZisZwLsLl7CaVoJFBZuDWDgpX66cC0ZF
P/lhSf2CdVjd08vttQMwULFWCYRZ9zZdDovsw4+AjehsEGt5rM2yoSaC2prI173XV3GeymUNsNeE
FrfwH9KhygjruyJqfBSpSy2DB8uhqjDZ8+Miol5XrOPwEW70zNDK6ak8Wk3d7Lqf0Vc3XK7hqNt7
u0S0xYUYxXBwJSilp9GreGXaElT8Fh4Ddx1wGOJJFyiu3CSc4I2n8Qd48sgPV+GArZ0DIP+BWbZ7
gbE+r8LKDwIc6DaixfAfcv2Sufr1r1TPR+Htimkv+Rr0/WEqd6cpwMkktKBCW26/INuRAOO1lQUT
GG+ew9xU08JY7FfvE8eVQT73xOH4RN8LDIrPhU14vDK0ENutqqLGNn18Uj+rlyGmrsuN5YF+e3Dt
PrownGU3yPLT8p+fIuAvM7sChxvY0VFR70YOAkLVvwCCzWckW1Ruu0susvohxHR7J0DbrhzvBCB6
thVrWeenBZUxMJvUtlRyMtwtUA6RM8H0D8mWoilnc8ncxLmfVEUH66cRPICiCgGtOs5SjZVhXCDT
Rz/Z9iw6Rifj54v4cJ/5QiHMQ7+wskNdIzUYBvKGIIUvJN0ugIxNG81gIpruTHIm4zVUlTyImqoD
/RnhCtEkd+Ot+6eEJm/lbX4zUDGOP4h3ah5vFT4KUVhYN6FT2BYJvQqNdArIDtuVYkBuMcfbfd6g
e52Fl7X7ZqkiszfHTmJm1ubQfnGeFVnlP+5duPDzWCqvvWXOlVD8jpCU6gHdVXGfbqbeB630nVZa
BhbN2KHSfdWLAZyamoRAO6Sys9L1ZdgVS43OevTJPhRT2gYWdVqbWVQzF+lZv0ApFaZMWpjZjVQv
3C/fraoYOW+2zU3eB11vnobJyJ8s7ZIE5/bns8cNjW62a+mXTxoZXiZtCxunhLnnxzcVNdjMordN
Eq/tu8inOAgDGctJnte0EA4dFG5hH55WB4BlzLdWaDv9lIp/5UWNX6cZmE+LVL1WSA2GKusT+M1d
Y1Igc3Ig2ZZNFKNRK6x9xsLxx+mzpzEBC6rh37MV06+fJpt++aFawEZJJX8ExiKfSCJ1cwL4HJNS
SOp94GSTZz1hNkXrI6/O5wOxUzDdDdQ2Xmztis4SACemgqbWv4UogprEb72RXaBXgAftEtsdEXpd
Jqt+GjX6X9EFl3WBBXK+wHcj7vYIgJ68WR7DVJRz6DCpJisviyvaAHmow75Ca/BJFnObCRpwZr2E
gnQffvNl+B0pua6EX4zzel6BSvrVB1dkv3/T/FpFfD7ajYoKf40i3fkPK3VYB7uvOztwjUS8vMlz
DdOZC15Jq95BrKKam+OGpEU+2oiKVFV48XVLpXCoq4NM7GSyzE/qJOooIklPswbAXr2xAWwu9TmC
fLl6uPWdDv8jCZepA8R2OOBDr/br3ZGybvZnZD6MTUtij+hv0eOZXhmx6winD3pb7NeqZRr9kpd2
fYAcqd4QYKQifltZ9xA4yB0C5VDxqBPo+2tnswhlfUPRytZBs8S7ZV7JLUjGRbLCVR6VVjk2rgep
mDxQBr5O+vsh5+8w0QLadBMfOUsFYz4AZi0nGDc0i8hjQMuJHbLzem3KIx/Q5J4/f8LD5mHy+Ikg
8aPKEw9wNTAUPKqQoX+kXO+xTF1bSxSidOFtxrOlTE5v3JdY17S0AkjWRu6/HssvseMPmqTLokqd
1JzTbK7ezZXVxyyN6b7emybdOu3OPk1Ar3C1bMXyx/4hRh9VPKMngTjz//ubi3eEIqv2b7pRAsnT
GJSMqyAWNixPBhT/B/y/CsNf/VRgHQmU21qGVXM4s+mI166vZCieTeOzBe9Iy+mNFI2Zc61M/Cop
8mdn8ZMTAu08FlkVv34MBu86H4La0psmYDzSHxMqvofIKfMkTwM3bqVmFsv0mQenlO6bD7j9krzS
tBruiERPcOAjPp1eq5NpySAVY89GcNFr9YL+0EaP1wEMc4sf3cnaXVivZWIdjb4eB+nCXGzSa3Z3
VoJQItPM+23RXWbLjqWF0a742zLoTGkVWdNwp/xTJD7739CaaHpwzylXDAHJHrb/lHtvcr66E5Kn
n7IA45GMII+XxcJtDzothQFkZznyl4A4qCUS9M4rEDTcvwZVO479uNEDJzujDiGmGx88hBUgs6TI
s/tmiq6vRncULgsG7r8dnM96m8VVZiV79oOb6wDtIMJAfpcyJBV8MtdS8bKMC++wP8UmY9vq6lGO
DCMo0Q5ksljqtmoPk14aYM2uuiMtCHdkGvDtOIEQjfQqVVU8bcn3wrJT2qNjLj3HIR00ODDIrMJh
X7xXkiCAGBoBHaPgZr9CAXb8X/RGMqlfCDN1sVS4ri+hm7nM4SGRhWX9JdDDt/FVMeu2LdTDzvON
/cl3XWtFV/aUvU0C+azKYyNMHKIaXjkd/sKAfWq3E10P5WWZ5aOP97/8hAE0qCHNvh4n3qK10wxE
ru6EZ2wSr/rUy28CHbdW4Vh37lDZ7d0aZCF/pLwFCl6zDlLm3TLfyduTYZnZg2WEyUd2/350cL1E
o8jpmPjf7iKg/RcO/Klec8GOzSS60MeffS/mTng5yaampo+VWqn3TqLzvy63Y02f3NB/jeh29kc6
JIws7Ipnaw3niq8MJQL5exKA0kyJiKT+BwWE5+cNhX+LHsV/qD7i21nje6cfpWmchqiA+1SNquzF
c/E1Ef/IzFJmA6QwGVaWyxlVtiSRMdxKL8/rEM/VZ5wHqfY9IYAf83g7DN8pwm839GKDspuUB1Rj
PRnbkh45w5gZzRfHxpJDZyqJjMNcRA1PyCSXaGYRg3pURxzGG7vl/zFs6DH3sc+qvB8f/yJNd+mk
wsSoxD1CCFo7WdeFFzWMrIGgMPkwz/C2hzGC/8BXEUVBaVfhHiCd1djpm5tQsAEiWC1yNQfyKSUi
ntDef3Rzu5W9ochsfCbBryB3wOxpPIWIW0sNbLdi8hcAV6ExtSyJmgYLrsh9gKd+DunExMzMI74m
u0DHSqREIcFZYIpWACfVQDd/IU1tC5PS12bWmDwVsZROngX+EvkXz8xsewIOZAdwH7l8QDsYkIxf
5uGOlHjXpG0uySqCa5JbEWK0fcVHPDh10reAUK+c3MMXuyGD9UJ75ibWFo0zOw8tm+1ZBzVIbcId
4frKK4rM3cF4vLFFSIhFhODUwh0IBwWjmopgz3J+Xo7bLmiir+RIrHty0aSY8BMKn4UdJTPSvgwZ
AWKcARkjL4/z7OlL+wwW75dyyVauCCSjF1W1jjXxC77JkRnTxP3UhwbCy2KCIkr4ETVHSpmUs3eD
Airrop4wEHlh22fTt8XS2xB5JdruVzczTWUYvfk4TXWencDTLsaGIo4+QVoDbNeZDE5sNwyzc8nV
PX28X/1bTN10Ypbpy+caqzwoY0NQPAuiSSKFxx81CdZagKKoRArzFGMj2VyAbK9pg3CjNbIJEsO3
0pdRyZKN/GDz8rz1B8oi/0ekGXAn20tGXG4zDAeYJXMFPKtKLRxb7eBy+yA0nbxId+PLpaJLtiaB
I4CbX20YT27MNcXtrmKsTRfXURcIlPQAb2WkauEEsO1YEOIaEp6FouVIfSIi5HJo9pRIYUwhoKl6
3iSf27X1iEGkbx2y/DH7ryEQWZsyLluvZjzSv9WST2jaQ1jZTDReBWLRGYs27HOGe/8OvGPVQEQW
WoTIWT/RG6izFqWlw+TF195uMvxuaZMeC4TnSJ3//545PZ7/7Op6l4ZTZu1yGpiLdsQNn+bh+Yz/
dRJmNSW21XhAEXEaREBsN4asPtWieBmOHEv/lJ4zuDnTQ43ZjNfARoYqlRs+q8WMl7brPfPxgCwU
pS/GUeSylGvuUI/6Zoz2fCQfRw758rps3EBkLH/NVQ4KFbUPU2vKeluI4IqdtkMxCy6FPTtetnXR
ohO6ZjSu7kUVpslb6okuacyvsOTzf0VS+RZVA42AidyapGycQcZA7pb80IN+J2RNhGsJhgYkES53
CwWhf/pqyzKF7483R1H5ovHI+Y+S2d6k51Xl7kWNNrDuXQdFU7UUTq9bTSTyaO248rQIDAUTiN0t
LL7HbuI37Xegh2wzOsWYfTDHjsf0yOPGVhammLJUhit1y9WXi0rHFSl4jmq8O030kKI9EdGBRLu4
MdIOt85R9sN0JX/NUXKgdPVDWwEhTZ/OSrj1fsZQHemFH/K+EfnaT8CUKqYLGOJBukLPzJwg+yW6
vL9q8sQ+fzrOxK0JubS42H/NmTVEnUhi38l1kuop9mlFbQnEds9a6/qk8lS+yeC9pWpq0fPaNz5Q
MH1cC/YL+uvhwY1b3bNMn8gKslnuNADMA7wFyIavg/NZqxfcf7HecF50sIYwusmbgM6SZ5mrr9+G
5n4TmycFxXnsBG0Yigc2CTx6IBD+EHl5/9wRTK5mVa9nM8aGZsy48xgee3YIVThKHh7i/JdAoIMJ
9A0frBR6O2Kk/wmWWRULmMP2MUvXGYkZELlYDLY+QuH8pFcgjkIhHCmTxhxbKHTLUTMQDWcjkJLs
hgFwjlgdX34EuByma+D78W7kbfzxsRO8S5X7gSDjnFmpJtp2YiP60MXJtjVdGUmrxuRWPfPe0lY7
Yqcctzb2zTtmOxZFQJ81c75VpPeuqglfAOgtigdaOlRpUgRfB3jnbGpvcqJv8Yu23IuQiVJo91+n
X2SCPyf//tzrHJhiyQZvqBSCORwce60IYWyf15Gbg8BdDtQGq7yAQZpGarJQS43e9skmqwyMi983
JEPot+ZrdvmhiQNmUKwhgyAVA98bqRcsp+CsCsMVAUrI85m0DcnZT7zs1wfihcIyx+pDNS8wxfKp
Va/f6nh4ic5g66pcZIZULqjV3aKUI2Qv/OAHKH7eixJkSe8JaBg9afcKB4Z97usC7ZNhNauZKamM
4pKEUyECiQJ3pMX7obKkDwSLMFMdrrZT9XuImezlIZ+xZM/muFnn49Q3Qq2QAcHGGiPPujhTvsW8
B6Bzs6/W9WnHO8Vs4gC2HtLFMFQ0ihbvDmK3QZpYuMGxHPccQi7btMhvlZ4ZDYtRLk4775KwrwvM
kCwKDfxvoiramXKzexRIfR4KGFzUz6y0w3Om6cyYDaKB1xFsktqLwntxNVLnaV46aKKyWry6fjV4
hXJIcnJ9ZkRckqcrbC27U1689GLy0gYVCk7guA50E1K2MlNaNSI9e2t2wlDrpSIcvwR9uVc1kxHX
rpk2YfCTCGC8EVDmXi1ZRPdazgOiaGVzQ+l5MlVeQmP8Hr5RLj6U4jtreS944qxfVNTZiELeHz+U
sZLTjxCNNBBDwRNtFJa5hmQs5mDIrkP/BmLKNz5p1L48byPx0QBecaaHZvXEEdxDqbi6ZiHXnlXg
pJOzWb2JpQ/8/2eDQIveTCPKxCv+HMnpXrlC/ayCl9r1RUMbzlA2pX86AP6D9nSbEb/+su9rG8nT
VWulyp1SQ/3OAvU0jKhr1opSs+/NoZ04EKGVLclzKS5KtBPqN4hu2Ru7hq0UyaHhXtexvvosDGpK
U2S/4rdReTv4m2xZueqS6kWNb5YRL17cryNFJK7Y0c6zvwBdEe/Iap6TOordeS4fqJx82eO1IdtD
X23UfFwaXbQ9FKIhrAxwcw4cpbXbhDzMzeRHgPyzdXfBAeP0I+TuuuQJBT7uKGcBWTQtCw2ZW46y
zXgEhf5Li8hf9fZx+v4raM9+xYVUJbNYJZO/aelp/XExGv4J3y1+yWgWerr2FD9sAP8FLSlgdrkS
4UXDbeGW7QmAAcKyE34pAgAw7j7C82IncLuYyTwI8bbJhwoydRa+WfuxIO0JlOja/ft89rrvWaNZ
AHhU2pp+bHf3PPz+MRs6tKBiS3kBYkx78em4fLu110TEHgZ7E8b/MndyKfgww0G2Olz+6rpQVXVP
bQzrW7Kbo/QYU58gkEyIW9Qxyk1FUAqA/TekKiccT4D7P2D1S5dqKe465y4o+gnqNI/wjCnCOktL
j7Lq4GotfYpxc7by/p0k4amuO6YqqyEfLaQOGMI2B7SjSpMDsYz82ZM7IBJd6DzBfsOEJFLuiZfL
3orQRkqb8QzXlZP4QVrIg4wY28pUQjM1KhgWRudZgR+7BbF8y/IHu8/dQOwinvxM1A5fbGg+Lzz+
SxDnZSoLzx779jbrA/xSrk9wm2m/3W+fk46rxOaAEWGGEMYBx3S9GA9N9OoXoQuUsczowOLNJLuh
MihvF9eC0c8U5Ukiq0CqEMBT1Pxs3KRGc1vgf0NQqZRp3gKGML2FHUVu4Vsv4qAhHuYijgwEzflQ
UpkJXkDGVHAWWan/utwlMAN6UhxdgPBDveG0M/9qfzlhU4W09Jkn69qT3bM834YbHR3KyG6Oda6l
BvsQwfKcFgvNJYjf/2jF4HR9Toyc0zqKXJd0Cl/2mKrB4OD7ZMtxPog7lLIHoF2zQ6X5cwo3EBDL
YJAZ7j0esgITrOVzwyQd3k8W62hyG5IEE3WpSMjliPTKJupgddlUzCN46pLUSbitf21rycY1gbfZ
5aYWUQAMHQybF3FoGDpq3ahTXtppNPcP1T2c2WV03jPDPcv02K+QjjOmTaEYjq8bQ8W07krfQlh/
HI0EjAAmDC1i1Zy+nVmZah87wSOkBhy0ehrQAX4PqiIZoCy5+OJrMm6p6YZl+JdrI8Pu287pWbbN
nQbroV71j9xYPAAHIurekIu3g+oWjGdbp8RKzFVUW79C9rsRdXj0m/j1DL6oKMVztji59EnGgzHg
F5Aiq0JvdLjVu8Nyr5BG6Xva9K7m1ZKPWaUMqnrZYu8dkEK5Amg6uz6OCY9Dy58pJcLKi8SbErBp
OVY0pSp4LXzCc5QmyTBfb00BYIxgx2M+w59MEscEVmqI8NYM5xp2o9bgadu6Ubj0PO0eSpx5ny/i
hYUUMqpA/jo3hjfKE0YXdHtDHPKdtSbHHBqJoy587MkKH683wNgg68rEfKjp8gRosG1oCvvZdw9/
uri1T+KCTBShY9ErqkcSZ9f0aQtfxpwNPnANXfNkNUkeOCuge8Xtc3sNBX193QsdClYYRjU0qz0x
i+CrpGaeWjJAyivQ0jF+p5ZDnZPjBQE4pwiT93Az8EKBa2Mj3RtSr895w3WIJbD7xk/AAEsU/mxG
jQJKwRDMvlw5vQOotQ1B0EOT3qw/26oqE5+G9/Cw4ZVTdb3yiNcgtQupy2ugYXj4AMgDQimlWRCX
7LVdxTawIMzN4c0NI09X/Od3cdeEnhic6VM5HrvVm0s99uDa1+T6VEXEhHVtWdQdNpFzi2xere/e
R3mOAV+puEYh7p1auXaiZz/Se3tqbpzi3M2hsDQ1SlLZVVbWISOvLp2wZ8Gk15Xww9/s+z5w//bL
J/8r2siE2jEHrxT35JeiyhuVLlpLHfchWrLy8kss8U5i8zHPc+QNvIWHaNz7tP+Roi0Kg0XvaT7H
j3cSPg7D17iM+EK/dw/DfCBw24HAaI1DMbXXTA2iGTt74pFfzLHo/wfHZxe8Tm4m1fKMa0cgIRGG
3EoH3dEV/FKehNi8LXg9gcqXbpgd4SIfPcKNJ0feOCHs3fyi7ReQqvbYopf8hSWLiHCxvl6wFNXu
06GIKAUSBsCkNc4OKnc/jkdjzlYyBynrgy6M8U0ZjNJ1qKyznTo/o/OCmMUwujPl475eSsu0clAv
GcCn7E5w9GcUtSOF0S1sqc2qhMvdUJKlzxB0KdjM6wpEwfudPh+UBWEPQwQePkJ8kKlbw8E3dvdj
toN24JntvHlqgh4JCwz7tpXhJ7Yl14VV/BBNlyACwoGxmBB2vV0E18i4zTpSq7JLUYJRTXRSC2D2
2d94hsI7oTI3r+K5ZAvklqLZF4xQS2y8itI/uzDwhnJuCRHfSAW/PwrhE1oTPuGovquCrTajhlu7
cOQckWrnxlGA9sKuEP+zyxobqe0/rFmP53NwEt9/HMQ0VaIQxiCXmdCcVdiba8lwBnBXOq4RkF7H
etgpXlB/f+o9n5To0UvASAuhGAlLOAOrVkzElyY//dYD4rWUlU35A1jdRHDMhQhkB/3YQsbSuZJj
9MbEM1IMxlDIUEtneiX7mUBNV1Ij6WP5JD0AJt6EMD/9htuM2J1m42gnWTn9ibPNr9NjIp7w7Gpj
6wPPjZ25lR37LC6CMDVSaouzEhTQDKpxkC/dk7agkQcEPvHQiwfiQPBtjURSbWOem35eRhcB0PhN
8xzJQXh33+3zomXCnxSG4FuEjT1xjLgpRMzcBHvQf2F3r29aqx+6ZAYA0COPy7aOUY9JnlWfkPZY
W57U4+pOYPFWvWzv71bc8GXZ/DP8LdUnKb9lcQr1RPNkikMOOkMqeweaUKArTrUqhT/HMUz7L5Hz
iyUTa+PNoZsYD0DafhHcomY9RfxtjRpOr51yE4wZj4XdafDXMz6we+fVz/EMaJ+JKQ+ed3LPSurQ
eVrM/GT3SAHM2hwvkyor8AISqZzWk0z9vkAEje37L1RdTD3TQ0vuKeFTacZ4QrumJmfgiJDp02s1
2UvGv4hv9YII0UdohpbYmRi8FAOCMPqS21x91P4/tuouUOLA9yYuHV3KG8Qr9DFwKKEM3Ynz9gMv
sTqKc1ixPqhbpXLGRelysFEUtd6zhyRn+e5EfSJoYMzHN+/Y5whEv4AtrzzmtwUO4+8OE8Hws3BK
ERJP4CSIEfysNSZWYQC5IR2xTQ6D07b5nvVa1K4wAy4d5Z7W8mvFvehIQ2CgA0fW7JJrlV6QdQjP
35kbyJoVxAu2ef+VcCEcPZte+e7K4uTdSGVP341qxJ1oeWqucA620Wuju1YFKLVGG8/ti+islUaR
NHndZ8BCja9WN8qJuFtI3+Vtyz94YYO5iIFaRqjZ9jlePBTAO4fsszFkdlysA96tJECcJSF9vSXy
Fjn6//uTuQnF4vf4BRr1bnCPZ2cbuCnOJXVKIbfhan4+VLXLaznp7dZeZ3Rmi0+SryadL/ozBVyV
w+dyHvzoY2Gni7DmJsCFNgDtDZE1XzBO2ijou5A6fegzqXiuzJDHJj/Tyox2nWzqpSImw45krIx0
MxQcJZF1PChUcx+cT0EpogdubogSpO1ms8AYFxblGsDnc39gHpuHrNMWzT2ojiej/ineYnhwReDf
4UFFlxWffkzLftKwN0F6nZRb4hz4XBpuS64Rl/mIaadLkjGex5eJmY6ZdNv90haGbEDKwlbmFQ2m
EO8s9WELWbzxfHMJUGfvz1En9+CE/EFd0tB03PQHVTsvf+tWx1U6kakP2Zm65uBd5aspSfj62MJh
qOzktjCK7Ul4CT4rodmRFZvhngeMPBZWkjSJKmvoKV2HB4e6OKrt5NWAFr650CilxryGBErqvQq7
eAQ5/3llza/+sgKpW1bHRH62VpP3yZI89kljM77Wsnbgd3T12lhy+vIJc0cTiPnR5TKV1YRlUaHB
uXUKYJ+Dy7KgK3BkDArq24P52tzRGp5aBZorn8WlwLYqy4k9l/IOSAsqO1A/a1AMlAe4opHmK7hg
rGPwFkJUQ8Pu6lQrltEhxvaMxY87e/0eeIff6Rpx2Lr7AAS/XylhO+0MQUjc+hFXb7kKaGx/iQ5W
dFcUNe+Lk2ukIw6CLMRORkgOAoBKpNdeibe2BBIHQA0dasb8D40OJ96YvNsUKptS49g0PBbUoUx1
3+7iuaFb3cEGHr2urdtQy446FPFQhtf2tWPURnONPLf7pSWVPjb3kT+krTm+soYc9SxN0dzGSQTV
jHfIY9mu1M2eXUMSPzRyMCWDEyL+f8d7jI7FrS70+bNkmslAzN9ItzoEhtFtXINnb1Y4uLSCljFb
VPJ6ni5VoY3P/VzrAiKu6VVTuZ/m0ejD4eVKdkjopomgj1SDZVz7AKYuGc53eMvhhoRR8BK2f5sa
yDK8r8dV2I0McVrXO872S9bVvbi3POr3VeK9FSGVDf9VHW6SBST3OeypYFcmA4Ofpv3ROxfGKOkn
LyiOpro6Fy2agekbO384pjsq8sDkoKxZJOOAWbpGOKeviowqLizBj6h3pIlR46Fd4qyXGtZAZCd1
RFgyuPWNqEWPmUwQwG887CGEL/8uXAswdYWYhhU2WPtSTT+5mnIXliAabaXwDBWbFe2RiD2hYYPL
eQeiwz47cIH6l8jmQXNiiThuyPTVBwGJXkq7vUN+rUZiP0S4/3BUqiwkrSXOqnJDoEgBUlLgoZDF
bNTzUuzqaFRULNqVBQD7iTf8ydGlL8eU43XzBGMt3EL3UQ+RbUevOs4PyGAlk2/3czOkd/d02oAw
6wKUUJGRQ99266QHcWUO3zQSgfmP0nJOFSkDl+BlbVkGarT55JNPF6RQKo8LdTT9hSnR4tORNm72
a0gReV6bOKAil4S430JmIOMeXj2tgw1MFzXawQGwhtyk7hIEEiiUNJ1ZMIdOsD0KcDStXBcWejxq
VSJjgCIFwtWba6qIxykkx8digUMdJiQDRafZNZYgV6PpBybnzeO+JZ7Ykrj8QlaMSTIIpTZOCvl0
N2h2SciYZV8xGZpaZVfTkEt96UQ74SZxa0MZ035QKPx04hWOE7VprHekDEpg8JS4LRnMAFsiSmN0
X26LzCtLJfn44h3wY2ixcqhhg9s+CtqqEuIbGutJap5SGBCvtqhOs9DCc/Rs+0f7mRNL9pcSXhuR
XGKArpMiL7XpJEiZWrehtnGom7Zf42yj1Qg4fooHwmRqB0vlHHfcMYorMZlz+plS4wWan2vCtd8g
4RaQYJGnFUgu7ITFZrtSqK8Fim+47QIhUgdUvXRYyRF6tv4Vkv9jipZQcdnPzAWN3cfbQgII72yn
8hM4Rp2GYg6KmrpRsOqOJrlRC+ZeEnG+1GPjHFAN+Q5VffIWi470xlEPuOb1ykpV024Icgkj3KMb
dLYbqMnnFyW/D7OFlRnJoqbKFxSiPq5+XQwB5vVjA9fkPHYRvQ43BE9GWqrhUGy93ekdtzm+vm9x
VuOU4XK2c4BFr21hYJKcoM6nKpiCPvEstUv0jfyonAgNF8y23i5ihGW3NIGsnMIguvwFtIvml287
wQB7dmqEwy5Z55tztVdbAcZtW28HLHSQwOeMiCaR8kM9Pyp/Hze3uWrdNLGR7kG1RXVGtTLV8suy
cBtRBS2r8hFFONA/J+JgQZsC6/Z1Xem/yAow/QQluAQS6vmNRIJOSjSMOzsSlGHnsxVLIYQmCzYu
XGnhMFL69cFtwYaax5a9XpH2LGsKNca7dkB0P61lvnZxWPEsiXRuozHwkwhpoSIhvfm3wdlsjUD/
qy/UNAVQPE88YlFYdq3YFR0n3idvu3UpcUBUQkArIo91svq40oWq/Z/Rgbdp/IQtYh3VtHDtQZZP
PumDfz+cp1pHmxgTypRa+Th15iRJ5orPc7OV/DL0uSHDHD3Faxqz3LIP9abgmiT+jDCNWefUF7+T
sNfwvGri//QzhzvtO4pyou5s3nGnqzZOjwI+YTMQD7Fm51GY3CzyoUlY8o8yRikQyL70ThaMv8/4
wcfGjwU8Q5G7h6Qegow32JL4AOFRB3S/suYxHpiTiIBKeW4Z79k07X3UODowQVxSRElbNcqmYXCV
QIygXpB8wESBbU2cPPukWJ7Gd23bZnztp7vk7gp2FJ8Ak3frFMDBsh7m6GQhGujEmjJEo8kL4e5/
t0oRvsNoOveLRQcAGbFDkexGVASp/NgcWrSNK26a5MYckOZBpInbBgQs0qW/j0woX17VQgD4eCts
nfZOGcdGHNwle84KJBNXQJNEQTkNW3J27uH3SNrYb+aOOV/qpXaSKbkSXAB+FXsargmOkl7zix/Y
mZeJ54YZXA/+hpXdh/3ZFqGrt3y49819ndANvbrQcUGW6PMI/Rkqkjh8dGeIbtVT7P/GLQgS2zwF
CNMEryw1PbQ14VQggF3mWFxkzxQQ9rKAMeC5by/lIn9z/tLe/DEZhg4NJPdN5xYgABGPe5CeFmWk
UZk7MvpZrxPeRoGQF2S76GVrHjKKE236s35hY4IrN/784EyqcGv/0VRM6cwNihFwrJ6toT6jjzR4
oAav7ED+5KphnYD6cTjm04qPQwbjIQOzPSRi/DiWtl3WYOPvqhjgtjMlGPtrLezWKUmOXd5L20Dw
XMALy7GcQtfINklxUuChGXBnOcfKGEk8hGy5RJVpHGyrK6J/zNKRhBZwgA+35RNz2t6c5nsIFH9d
+rQTglqCB7SGJl3OWFRno3NBTPQC1hbya3DVeo34TYY0mxyLzLQOXQXIEQxijmXnyEM57Tq2sXjC
P1D4KTnyjw7B8emZ3xC74BEMyTh7DcmBeD/NXtqit/synAvjHP9BfktKt8ZWUXqckIy3fzFWzIqG
Y/wjvY/53Uae+chicSH2bs+O1Yo3z2ilRYlW9i7RQM91h5gYZiCrFx6amwNpFdK/u5Uw+VRL05Tv
wb0WlPLu5yP1GOQcrqfeHQByEwvG61Ogzbzu+R+bILqUgdhvLmi482imrsdc7eINyhfJwcP8wVmj
y4bsKxFI094MAJykelUt23n6Oxcx/Kpi8+SqCPF5DjhFjGvhAOz94UUJW3vcaR9ziZF+DRiLw+Wj
sXo8l7Hf+BRV6qdPC256YnWnGs5qdHADR2NxQfdokXsF/1W46OO0e0Y53skHcljpOtYm7mAGPw5M
fmyrVIC803LlOZb7G0AZ95SQPtdmnk5F4xRtgmuw6Wv+6NlvKOpdLjrIwS8av61duxO03LruSR8J
37ghgooUPEJd/708s0UUs4Qeitjge8oDmmx7Dahoh2jI1IEq/QsSe/L8g6uHBYiCD/dT2+5Ed+kz
FIORf8mnWKOcx82QlaItcGxPtdX8e63yUWedunT35/L8nHoJK+8Gx0u80ULjKwjXq4sX14ByGOdM
cyFzkVfPhaaQ+pM5NYuYcKjlX0FNm9wB2QsuzSya6NFlURCCjbVAUVwZfdjPCTBGQ1PSyljKSUu9
zEIFePJQrAE5bu1MCuHdQVMCQTZVJUEGO8I21krZSurd34EW4SJbZPeYnwcXIDDXHk32QoWLMY9u
bO6Yzvzj57nnW70SDhYxIbPX4HwoSwebvhLzOqz9AqqJGn6Nkls5arFP1Lv/RGDpAhhB7bjcly/d
gg53hFhlHPRkOgcRx/+G0dubfdsffUeE6Hk/Z1qxY0+IHY+YNUa00410SgesPqMuBFB+b4uYRkoP
9ABoYJ1rKkP/eBLXkobcBdtcMnLQyr0vn9DeNbAp9W0vlavsSUCoW0X30uVdldLyNocmuVl5C+XW
/3u2PBaDMb0mZFXmzzrxZL2TuN1vw6V80zOQ+frwCT+y38sDanNoe2Xly2LyBkJiGB0d5YcWZ53Z
ZMG8kvPSJ+zFaC/hA+aJAXpnZswoufdqUrIJfuO+N4FdqnmJpSnbT7wRP1X45jsAPmoj1Sm9jTzx
fR/qPj4MtbURfb1B3EHErAr9ATnYB/ixUx2btHGMdeld4BdDy4/q7WnzkNXt5dNyc1AQwrwtM2UT
kWWnWP9FPAvDU5NLS7UeIFziMfbSyE8Ax0+rB3j8ILUmWB3+07xTo/f92tFfZJuqKeO9bFiHC0aW
L1rG4PuJbZ9Y2Pt39dGZQSLuVjqJgGAkPnz9ZqnXiFCj6TyAkXQuGnDMcyycsshJBy0NyfBFU4Ir
FdTDIzlrvgSyLRKR+LfSwCwShJRP5VxGPop/fLGsLCu84FAgsJBQM4iJlBv5WcK/vvuvJ1VXiV6a
8ZZ4oI6l7HOl7+LHH9HUK0hDnnUhX/jrNP7jo4cXd6Mer4ItqLPkfVryexPc1LrMjyD2I636vgaD
gNOWNnpvUteZWmzd3iS5pCxV2iwoIyTfwHTjNzEZlbngATlepl4P28lrjpCwoYvFeQwlc2Pa63LS
svtsbsxX4BoZSUf+aSt6Vk3mrU0JjZrJx5LBktRMRTMnmkswT0Iulwr3v5Mc63tgUxfRTaVnwVaJ
RPsKJqRdd6eFAjeuNnsMWZ0vlhIEylPrmOYOVFYHAy7qCORBSbjYLQnZCFNAvd450pLsqvVJPq5R
WWNpVFWouKFmKwgRiJACAsys3GMRHqFa4fiaZ5yiloYhYYI4IVBA0WW0WOAB2zTpT/PxEPmtrXMi
Q9bv3flTToeALTR3Yp799dt6bikmjGIYpWcImwxtfUQjarhEZCUy1baDnCyV+h3n/icFnGJzFATK
xI6twY5lofILPkyaPip+zyZ9RXNNuax7RCp2TuueKXzVuY3GQw87K8idpxHy07v0DzgajVm9uzLc
gHqhQzt+Nhz2e4kUfrs7gCA/GEjMVLa5PM0nFAFzJX12lj6j9OeaqmF9qYJL+bZYcbZjNxTh6BUn
nBypafsJCUJjziYN4kLs9SNGlxexU/fncZQ2w/ZAm2MbjhhpA+hToXtRNK/eCpyD9Y/GW8IAVUrP
6Ov6jehhR6VYdfTLV48qfiOMLF40Uygi1Yb4jW5bdNWLBiRWY43vsNebvbHW9dFqSMJzGOdzXeau
GRvbxoA/yvNkvlJZa9/btQozQ0A0vhtieSERYP2hKIJ3nog6ToYlIW3ch+ADIsChHO/pTUN1E8FR
GQzFtm+Qn9r/6tYZ4Wt/NL/oGCPFIBMQe20cl5gDmnUeod6O6q96vzNmwYEYvzABTxxYCyCCk7GB
gkd5kEuLo+VFNPoYum1ntLtHC9mqoM9NVuYtk/1miMPVYY6SpKhPHvKnRGeXDvHEDqrgWbWjVoja
/zOFYmfkunIpsi7rzKd2x5BVQTOqKX68PgK5Eq9el/t63RAxT7a36C6VPN1aU9ndqKi1Gh/aaEPM
WdhYduWxCCc8OG9c8qydbWZGnNjoD3ymFw7D0DnGKNzpadTTzNM3NNlfh1YQsr608e2cUg5fJL3u
iEImVoZ2fOi1hUWIMWFORztMz/cPSUYDsY6h5J1qLJm/2sdRPxl3TA6zZCpNLogBoRKE7Uy+lDqF
K47W6ioAOB8nvQqqcqYI4OpHqSTgfUXgmnt7dvW3vKU1y/MZTUNnVQSsJQ8jxqbs8wn1aB41ckrH
oJeYHprfWR0T5u/Yg4EocF/YOUkMgRe3f2/VnlMfi8tENP9JQvsSeOd6uFhPRBW/MP9ik8tbutLW
iw7QwIOD0qWvNmSiyBwdUojRdCN9tPHsiOlGzl+FYILa9Prw8sDulSgrl6zI1Z6Gw9tJ7A44hICc
5R+0caInj56rC9Wtk5+e0WDV+K8MxJx0/OgAP5WD2RhSqfQsc5SN4d8SCfUkn4l2VXdIPUPhTD6/
SZlZjmvLE8W5jBcL6Ajx7mRh5sSm5YLUl8xUKHD2zK5SQgStIf0jDwDZMI5YqkUBTnduxvZTsJiM
1F/EzIhfp3Hctmwi+NM7sOqukFq8q3qFsCuBaUMoS/Mg1n+o1WftFTS+7t6wARyHlfFetGjep86f
ckl2DCU0Oe51rbiJQthaN1TYAgYuXq9zmWUx6kwT6B5shErteVLIWrijI0J+TfBXZqCypxQy9Hpn
JDdP+eFI0ZpA9NTASbfjnOP8rtoj9J4cT6lkfXzgFlWS6UYH30lHavxsJsbYE+nx0sUFbL12l1EH
jgG07aaShWtlYXfwoASNnjtqR2YR3A6spR/BAZvUvBnIedNOwoKw7Rn5ad3GfW+/JfDWiYH5TgYj
An+9qndZnOwCqBau4Lg0bfG09G9BvMZIYWTbOwUGWj/deRui/gXZ6AljWSF0SkVWYM6mo0dRm92S
w8GdDFpocrZYcYPIjGTEqwDtqs8xUr1EGj5N6Ez3Tf4+Z1ezMeC4hpxjLyUgdCbkSw994/nP/wAW
3bU2BE8iGEz2w/6GsaXk1l4iy8r5lgcpo3Xi/vGacDtX6BDRq5D5pP21rHorHSKEw4/goJUej4jc
M2gYcZU63SsacViFouR4gLIo+BWby3pYRc1j2BoaOkRM0Ua8uEXhJ+8bA7KjyWA3KXzQGxhNtO6R
SOC/zFqC+mlXOYj1I03lhM8W+c7OQdVGSog7oHi0a3eRMvmtoFv1Kx6qr1oAmHM1iUhU4GA9/+SO
cbBLtwVwgxk4pykL5kAal1FeKj7dWqy21T5S2FRi9qK7s/Jf3klu0jrcDD8WePu+jWkGt9WtOgCH
zPfYdYyWsbYzu2s9AUzSsnkhNlLBPLMpSxWcSbLDlOubORL8Ndapm7MX/kL9SeQeX3F5nkOSL8Gr
On4/J0CRqbCiCoP8epdFR1UtMM+7x2wbis8x/dhvOE1zXtiCaiOrgrmlNwq6DLyf8/naWAQUyTyA
kfyQPZu/xxYacdo4qyPX8p9NKmKyILpXW4gJw/pP1hPqaApUXaillTgMcd+5o4ZxTymA4gOkmP99
BaU9X4s/hHGFZO57Y2AnL2YmL9AmFNy4fxjs7exZTnux+QQoi3yDFL3DU//VOz6wI8MONqC346yT
qIMOdYEpu31utx/TpCGjVcij7Ge8Vz6u6122mNSPbp/d4c76+XPP19+95dAm2LztyunZg5vRCTR+
2RrUglbzpBcGAl3Bjofk8WAXy8xcO/gzX2ANK4n5dxpufmR5AZufb5fbKe5zvX2sSSMblZIjV14s
34QVHJBNtIeNC4Jjx7hpWsxCUbAS8fNpY7uzxcxV0/tIToTTYUpTI7T1t2FhbZb6WK/rBBZOwB4G
jYTnC1fbfFyjHDZYPEEMv5TeoS0y72GzFP+xgQdoYDzdx7ysBCCZ0etRxv0x+nzvWMfCDNrtq5Fq
PcSZdaPIlaQADXfDuYr8IBL82rtZj070rWxm9+7WLz2/NyIPiopFwXGCANk722L9kl1N5Fj/goXE
uO+rC0F0RAviqu7t4cKjyql1P3wpntE2/gu9UDg1NIuxGt1UID634A+S0chXLKdlNPfqHvv+JqOl
SA+TrMefTpYbwvyakfodCTa0i0LwY7iPAaZ/O0vrNOEif6fdsGLlr8esFx0D3yOP7yloWqSSgkNm
/wGV3CEdZe7hS+CUXpTVhAEKjIHGVjJf8IQlx4wRDcuWU+0Gn6TlqdcrKgOwmAUBz7Ji4B9WzDOv
fSzlqdhvph25waKInN70WWQmPi7F2bVOyZb9Yu5zUR8zw4mtBepW43o1caZaF10Wibnj+uhhHS4k
Uy+OOItg73eQKoK73DpSKIadqCUt6hAQhNE86g/kwtpZX7yxGKBEvj28Szl6+X9zBijAsE79kx5T
0roD2mFD3Is0XPNynmYSEFDKO8JZsbbcpjZJ6vDRpvkDCye5iTU/Xxbp5DVd2iSbP9SO5dcCZl7B
oOaEGlDB+h78VXYJzO/jVmlEPAP3EI84NZSZIYVm7CdOrhSISA05pebtD48RBWMQdvU5GYvCVP/i
m7vwHit1MKxY9NY5TtlkLACyxP+6rbtNxBuoVOwWtl5Ub4Xoiwz/Yug6Cwy8ZGXPPaQmf8BBrSuH
vyhxvRMgXexsCof4Jf5W98huekWoSKTAqFwngODZlJPJfs25vorxBza/w27FciqYUF82V7VsmdxL
3VDoFR1jUNqYjlZN3I72i95ZefxUT0rAkJx+3stpUGueb6owZp8olkDoZyr9RnDGFN0JDyfWfR67
QSpkN2aDjHwHxdwTBvm8FORJLaNTwhABsZ3usqnxvmKyHG7cVoBV73sxQRGajjXAILYH4cHI6EGn
FT6McOYSD44n970FbZIg7czZGSqVDOGmy9qiXVXzKiWDhM+J44NDv94/aCUk30YmoF/BYP1vUTDj
P0hQV3LhdGp/CJyKQkm69ihzht+l/bJhCSASFPwZb7KUDxMF8cVBGohi+9WJCMy1LVhmEs7vhce2
hKCtLiNwXwrp/+NKeflICNHqLh9mO4kmDvS8ZN3pT0TnbAzNLio5NqmQ4AcZupOiC4tA/iLhsl/n
bHUf6LU0L2nvwn2jOdMBYt5LhpJRNVBuWfRFYAQG5shvbDbmsrMIaazwMRXRC+i7sKyWPoPOUtwQ
3Fpxfus8DVz0hAOoFfEIfghJBQcudxECV+RmM4R9G60oWSBQvX0WIDXBD4+l/7hQYyK7SiLjN7HP
jFuBnr3FIe8VW26DudMEAkJAV3UTgwr0sv/XpJz9YTYSIGfcr5A3yXlEx4USqYIO6l+/aA1chnW5
8lMy8igwaRceu1xSjBkEXEfT3P0DcOJd1NmVYeMtruFGDkJXmmlfCuCCPiZKAj+n0NXQiNPG5z4O
Kv/pMofysvFv81etcNloQPnYYJhs4hhSXXbymk+2b4q30rKnMqhYHBnAFKOCu1LBJMPsdDYf31Yf
D0Kyhn4P4zQgM6kiYCUT+Lh+8wGDCh0zj2XifQ1V+bh4FgElbJ9d4RbicsxLarqOkhlGA+ajTh5I
VpZdHW4DgpNicUzuF+vEGzeDUNbLGIPr0Cr+rQotI9LtByx+8H05qE/vIDz14RhyGn2ZhWXOwZgZ
6yi14kkaFf3NKc/GSnoxBOimEMxLJ7fe+4d0wuX+//BtgrqIjQeYWWgw/ShBoU98HNmXJlBzkbET
MC0KFmAqT7rqoD8iK1eDh69I/24MQqZUDjFLO1Srap9toyqsf+uWcZQWDNQn9k9FnoarEqvyIYEK
3LmcNTOisN2hF4a0ka9qEl62fd05enWTMFmdfm88lFE44la2q3YIeVNiHavnqeNiiowf4ULg8ck7
oIoZeXClO4aVJr/ti1dZ/rOo8BHKVJCAhrqMp9lgWGkyqV9c/4pIaZb3YvaJj5WeNgggBQa7GVGS
BsuKswRMNF+1XSDiZaWHOeTV+p5oC9AT74XHLZwntCNnsD41sNx2TxQhWWg5DdDpn0F3iu/YzHi3
bys/Q1BYSiKPEiT/pO+dcSdLLpfsMQcfbDcBA+D9+v4RREZDNgkiyQhlRaQK02kANDfC0YvBnqcP
BXRfp6C9TMYmppBa+ZgWvzdQA+ktySSh7EWM2Py3zdVf0FZY3vRMGVLKP5oL9hACuSx6+DHAFLBx
/18x2xEKD7OcgsOQ4zN7BSj8FBy+NlhLNKrGQ6IKUh0yPT4du++zs7XwUdka3ypdOn96Sv3QjKF6
G70KhwcB1T6Up5s6NCr83OcWOg3NVmi/XOf4oV9BL2Hm8mK0Fdc/S0vM1a4lLhHbhi5Ah0oACsr+
VdER1Sz6wqO18UovaVdjf3tRq4CW0arsi0UmkQiEOr77AOjSqITMrwPYC1GzILjvjkdWVO3Z+Jw0
ZbhnreegRRCdUVQtkq1DzlMEdpiv/Ui22vTJBSUN0CHxYAlYtklIs4ord1H+W3AGv4zMYS5Gnm19
M5geDlb7bgkaCFsYGnXsATRfknh1djH7rH36Vq9U2d45Zzaeo3ddUUaRqBWuNE6yxROgDofQVFkB
llDd0q6O6g2SQmSNfBHCvBaqLXfAq7BpzaWwHhy1eaPrAaZV4JjnbeOlpXVhNBVGQGa5Sc7P7bCZ
7y9Oq5/335yMPfMFVUkJrAzcVE3a4m6M7P8vmsWoSb8x/AKaY3JY4NNkTE/rWz1ps+6z5p1sLRbl
BJG8x/fwh/+kPur8GWdqVIgem7YOwX3FeVKZ5QhqKcZ5LQ0ilQc5+sYqcz72S7OaqiUKbgRjagyS
0VbfKSyrVQY+K2EdnidDkSCK7ouf8Jf7Nae7giUhhWi+/4fwAxn5EnvknNOAFVRiFOB4Jvr1dg1b
c18ppRzMspG5vQABzx8zam2gAm1Od+FBMYLmdDMLAzJfZqXpXq3BYKR90PEeuejVCxKsIZ9qVN3n
+J1ZgnnggVZv0viO1wk7ZHu63EN6uXIzF/E/D31WsBoAcbnhEvbh6VcQkrVk2iX1mjZYspBjvaC2
qhbo1frJPqMDYSvNIYZV3kWEwoNjukIODPtYZw61RmkGtdms87+1mW7dtFIKxbDDvnDFZExMza8Z
enYIlSJjclACcDzaL2Qq3Cez8bJXspfdAIlDkcQPnArc6E6qPcelcMSuevFtpyU7Irz/fGF/eVET
apvkZILv1oUaU0hTV0FARcK24hLUcZSi7RhPX9QtgWWB539uPgXtWp32yAAqrABakQjaNus7LE5k
ISSddUiJ9FhLaD9Ao429/olRHZj0h3qmSn+I1bwsxspZ/KEmGLd+JnRun1YepJyuC3FdANnB7AeP
kae6OzqIY1YGrLiWKHGc0vMZ1JfoPtzSNSNTqiRnTHtnhwXN7lRQ2ROZ6m/7tkFGPL+d+ro0Fspv
99ntJCeys5NSzYS86dy6Rv8ZdqVaFLWy5ibSQyhAM3JNk+YsPQZsjefBXWQnZ8kgjkTG8p7WMUgc
D2++d0Gb6mWQqs0GfMImRqE8eE6qTJHUZYTPuiEPrZq4dr4lm7ul/RaDiaTj21lrCIEF+0BSHP7Y
w+jEQPScICSuy1mDIurMy928J/+CnCKaD6Q1ZzvYNlZkgcZEZYOUB0UvwODvb6jxilfd//BuEmPh
qonJDlPeBbhnt+vq/IVPL7zesjhbM7lLpwOLKCz4fBdeUV5w9K8pXtPtTpC42ACpcBpmT3y/wlFJ
D0MjURoK6SRLmyZLYlHsS8TYNZvAsnhQgvUQ5XekQmrVDgs7zGUyyTXvPxWBN+/BSJgJgBUrFsvd
XITWMJPeI04O4+i3iXUI2/r58+ycwlr5M+KhBHcOIw4JZrVN4KL75KKYUDCu9TvdPMkS36xIo2ZD
XrFKFrKaLUCgFg+xjCbpdTEJvuYpd1xSSbJuItCKw3q6uxqYj1yWqbSFnOcQRHtPLxHvOT2K0zlS
Ln69U7sWm7IAS4ec8F5pEra+6RZSTm+oYXlVGCQBeMgmqLqviCTMxinHnW0Iz532S7qUmhtFmFdb
/Uy6JbGbtlJwhDJCYFHZmlqO1yhp8nAheO8JSOtI7ofKER4z4as1dJy1ZFh+WYrhNHvPyN7t/1+H
xJn9fyLjCrvP1lhAW1PlAVZad4c/XOYKTpRLCskC+C/za+RyQ167UhHA3gtgx2dMAl3ewuM5VtLo
Mr3ep5gYwwzqUcVYNzXx1F3lZZB0nlysv56Wwq/ULPpUULBW0ZFNvEOZmHabADe8/xcmpiCtzFpX
Ia4gFNSl0/5z1Hbai8bEPRQKw8m+034z60OZw3+tUFcCTrGpff7ZdgUJ/kEiSeA2k98swyjln0T8
Y1Q+Gu2KFxN7/lKe6ol/BUHnrY+U44pQ4QkCmXSnH7gYmZ7OvXx86xOvYJqNIOFURZ8rL64JDqzR
+YE+R0Vhkzx1CMPExW1XMOtl3wmAFxXDOpcOdHXKz1M692kOlcrplijz2AsYFhPzE3QvET6ZnYdo
hnfHlzculONRs8rwUsic0+rjvliv1tWSYAVfZu8v3rkGbcy7AybA1gyMxcvj7NDs7K26K0scuVkX
lMiuEruZDYqAs9bwfPFzNjpgpBMCFA9zNrxW3XacI8+OfKgxZWmhNu/SusBeLG897WfEWsa+M7gJ
YELcDn3wpGlkJcAHMDMYAQvpnvO4JgAgl3pjsLC1+XuTqVC/q0oakbBDOFzrme7Y0tPiRheAuo2O
fGcV7ZtJ7V5rT7oljd6jqLt/gJUMb9fVaaUaQUvXJuPUK78jSCK1ssSkpZrUHlf+wOQHz/iWtUc9
9Zko9XJelBM5cfM43K7o03Mg/laGxqrGZJSYYvkqGylE8tw0DzXPupQw6m8reozIXf8mCCyTSGUq
RlvWzAjyt6fSMFp+UohbOHHngBgVkOQerXAO33HK6qVc0aF1EAXJybHWZvnNB1Hh4+Uy8iUJI7tS
sTg5hj1ngjZSKQkKfzTJJO0OJpJJqB6tP+qaOnZaZwQ+TARUm+EpvHb1E+hbV9xbraALYhovybL2
pfSKkwaWdNsHSzSQUlhNv+OzEw1qsBSDsj0FPvVjz+p0qdGs0LJ0A3ompJxOXnu8byM9/kFQ/pig
nqgQ1em4uGbgnbysEMHdc5d7Xvsj1LCS04U5NZOFypGoS4Ao1lG/e86w0ZrXRbxMuY1uMb6LSfAz
/4bhUMJIlc44HP2Ulv6qqQTBz9q+DCeaulLUsInnnUdVcaec28KoaJ4EICdFFTvtSV3WACvSyas/
nx/EwMLEBw4+LKdEhGsdtyw0ByQhHsdwpG00wWJISKrIF2KD0XnvjbYGbVo2Wb9bCXf3UFayaFQe
y+ZQ1MsM6rVTZp0JHx2rxVD1XocC6f0RrsIB+jnOaetXEwOcPmU5lPKleMktSe/UeFA5J/Hvy5JX
hcS5O7f1yt0nmc7xiyZitHWLdJjnifkA/va/eypS1VWdYJRnMIFzNzXs4oBLEwLyLxWnbVC/7uZl
fPHsR0kyEttyIBCPNyN3TgDrHLMRe+k9fwZ4+qx9gvTJb+8UTsTIEE9nZTKeHNbNyxgsVP01L05b
WYiWSviC1e5i+xs35n2GBIGNDs+q11kIUFYasA2a/ucrPXNfvI4pvqm2ltjkMi601U3G2VrQaMYX
9iix8aH84XIznZXR74cQZXsrKJQPDmyBXiD7Nx0whXCVQhF4b5KBOWsL+JdOewbQJYWgvdP3RbnG
Rkp2+RpR6vIp0C7kUqO3GiNllHDDnn3dyJK767ohjKApsCBuyhlm0RHMVNRsPB+xVi2xEd5xxqHA
PWR4w/L8GZz19P3Df/fBuahw4H3ddkZBb0URMrvV7HybqZp5fe4TGV5VeLrgKIGIoddJiDrNFlQG
9LY2yF90+4xBD/auRYHDZL+VsvDA+u+m5QD8Xmi+BU4Tp9qTzdFwnXgl39Lx9NnwFmMoHRRteV/W
tmnoels8hijFJc2nitkU/vqO97pWZ0OeRMgfs226pjuRYTcz1o0SyE3PK4NCpsbJ1rNU3sSrP7j+
olNOG3ZpyUJPG2dAbmqMbt8+aoN635fxQNGTaLuv+o9QKP3MH0uS0TTiXlkPDeoDNhROcs/qNQwC
Mb1xaDuKiFfCII+V7UwrlnUvmB3LktxseNRP02uOAZ6Y98gLjjrbwFXR5ePFp4nrpaS9d2ZNRzfE
XOc3llXuNpobjDgqpyDrctNP0SURV7JDFJuuQA4lyU5tmYrUYBRaYZAhwX+ADGHZtn7rss/h4R9C
NDxUKsyImI2dJZa7u5N75qkZ0gb12ud8Z8U5ct7i/1NkeU/0a3PBZmypCcJtZwhb9j2YYH5/tdYQ
6AgqfGpD5Wt9kBZrkwgwWcKI0UV90oK/KGZzCSy4fCGzo0vgXUgsfv1tX9BlzPLQFjZXXugLb6qH
BRKzw751WPMN3wGgOj71i+uw8D/LkVS+SxQvBjZ6oL9F0xSzxEOgnk4K5RSzMfjr1yyCzTHOBju/
98FyMgdZ/66VysDl67HhteIC0nX3sM0vrG4/k9J33Rs/q0QLCm7DZFUB+kLDf/fOA1BzAW+LTd7L
UW9tmNSNqEnc59Nd+Fq7Kb0di19UmJ8h/Ecj129zJNrctMx/OklVzYVSOd+rz4Wx2ib2Q44Kw6Tv
BLijr1pnaaWL245FcBBzLk604Dgc/DOwxRYU6BRQG0gWoEEqiZmPqKmVmSidcq6rjWMbcq8KQdG2
iDaN1RVz+OpdPU4iuhE91DSaxwGYq0M5Wl6bKL29/BvXv8NTHJw79OvJHu2P/9Y99owBgehkCYyw
XjAiqLJyjzDoVYAMRwxkm0yXSbxHK0tmFldII2DbgWbuTxFLDzFm2kpPNNSfNi7e7C879JT1zVAZ
YUxit/UkKksAynEqOxi45KBjQjSYGsPkeTWbMOY30lVmrMOes5YdTBsjJz1kaXkufNFxQtqzhpZ1
8hfGFwvWqGFx39cpCo7ihblGY3n+Rzt7J/XIiydCSvRS3ZYYsME7weAIuF5ltdk0+V7Cnod2P9bW
KHAfpbZCq3sfCNH2W+FF6t3P+ExM+3lsYppcp1Brng4vnISIlkWp0T9dhrv3o+r/qfmVhUqNeT/G
LyNk55ntTm0I/KWET6QuLb+lu7cZKGuzrKZhtUO1UMLPEKlbgYn4iLkaMVMVYkzkVTwGJUcVV2q9
xcjqpyesSkhkOAi4vpi6eUR5LUc+6EvLWiMFtM1SpUNml6fXz/+SGJ1GE7twke9ZTymveC7+UXmY
BOGpF58hduPtM+JrCRQu0D2skb7g99rxLIzMzlWNN85eRxWVaSLyz9/sW5SfiA4eeuligaH8Nsgv
SiD/C9bqmS8Q45yqdrA70+KQQwJIpxrPCZqhDI4bbc5hsi2GKHM98EeHUTHiXSy1IGdhZlaoxux+
Zpmw7oCmPky8OsLaMCdoL/XhVoIidmGIcrVCLFR0hwRAIij/mlXvvnBvsvRHuc2HYxYHHOjyP4OS
TVvhHK/iVcvRIpEt0Nn+XGx1WXMO3nZA1GWh8UY4/I26m7jgbJItHHch+BxYJDZS2+BN/7BiM9EN
G5QrZ9XdWo+LBzYWN5N/umAVCV9Qp1KKLtVX7ec+tRtKw6T0ZzNclvwvQp1AKJvKj90Bt64Uhjtk
NFe+NgwmexbUGzFwAZxUEXkCC7pSvLz5wXH3Y33AEwNEm7FrOVmXrICVFcmiSXktFTthGD4i2WsU
MXGUroDzFYmis2O48TzuUtAjfqWeZqRtrTi6hfbIaUsSjj73XX5sV79wde3YAqSeZGIk9FYxTAEc
xzMAlXVItusXO7IZbpWYxszguorF04Z56GRv2uKofNToEOux9SxhTsA+t3yYDBkJl9uXb2w0O7Qg
CPxeDTHAHAAxcXxKY2K8FYQuQEVAbdAJJoYzWbn7ApKaEPxGVj32j8rE0yr4VbLbWI/0AAhqM9aE
AF0CNsns0LxGIdLxf31/n/5LgEK2hBDiauZFqLORNJkLWgFb1l0RiIMWaiimFHa6O+i9ZBY5nKOk
DYIEJeCkPFIfHtdkoer3aePT6XfbDu9vBm29UU/KjcgAIlrLo+Gsvt77nQPmNhZOvFv4dFDDuZtu
0Y1of65j9XVN6DZpbR0Kiouft47BynexNX1NaWvHFJHfcRhrIvRyhIbmxLermfCVzGvyFhPIGHpM
oDQe03Dj5SNIyKGMonHnT707p8YU6GiSZzM1kUNXNTZjA/mGZXWcQ89pmAE67tuRXR22ARsJqm4G
Y8016UGJITOR9NWQ6sM6TRNSLBF3QAb4W9D3vuBXPm4MAf1aZ2TO/WH4cicwzwHjQD5HKWxrs8Ji
UrB/cz9pyGnh4l6/s4M4ZNOepyOrAwlM+anYV+kriPVRlBeQ7I8aaGbyGEXlYix1LURP4rvKg8S9
lMt18s4vxyzkqx8Eu6VlI+6zZx7+7R07+8o+bJVS+QVo/aeWY2BaLFUzRz4pgy0sz6CyThIqNggD
BEjpfieU7qhcQcsdKb2Xdx/b/+IKt80dH8px1K3O22HZHMddcuCoWnh+r/CUP5cBJV8C3IK5pViC
BGQUT5XtQcwgSm7/9a3nIhUMLuzPz5b8J5kqwtHsomySZ3fY6pxrU9dBfOQqIdRGNskEPqyitXwR
fCfCKPbg5Pp4dysvlHSXVjm31ekdBD9W8kbOKrJ78uQ6nexWehTHqGwCo1HDBvGuyUC0tOUtiqDD
jxXsNunR+HJs6cUGMejq2iVtq846409sDpQFrL5a3jyRc2I41dTw7+jZhLsCJ2YR6TxDhXtvdgX1
lRvRQWk0mR4c4zjzwp24R291x7ZloEE910P3dtHRD5pUPu8t2Z2YPxIhAtHsM1lrli1eIDTKKPZH
Q7y2VrFopqgzCVvFI0jj7bzxqyklEUsFVxnXb9tSfo4Z6XQvOWDnsOOvuL2Fw9RXMPlp1cKVieh8
DyLLFQcWqmUrattlVmWNW8HZNPiUUS4+zahqrWSu35RT4Ng76FBLNnFhPAimy8aTN6X8z7qY1kwD
sux1GOiZW9YDCrXsjFTrFcFJ+zOS0yx2IZFa6tfOwjmzFVTq4spVVVPdi9TftHArTe8kK+5yQKCa
wKo/wDtqyBvaciQNvKVu+bKe1S3Tp6uMxP9shVKMvQGjggSvCr/MzVZ0HKrUsh+4ZpS44LRjb7fb
OizwbaO2YVHe5lAnwe/icmSoopLjNDPUFagUhSegHc9ss4O9Y7hfH+q+5jmCNDlzrPcM+VyJH+68
FsV4bDqzyrePMqloIifDXcDe5jLsdCOLh39A3CwQrWjZaDn1/rVZLx4gZ4xkUA48PisEbqE7R/O1
8Zuf3yNmzTegyFsz9W4GjxAc9JASuXwY5NmLFl1zWdYC5SjFfDIRTpXlaAHueIw5SO2BORO0lL7Y
7Ds18t3CgvnkppjYcf+OXHbh6vrbQh15CplVsPZKIfcEUZxfjQEi4o8OWSIqB+yOUBhazc2PZb1k
NPLbyFraqLCbZRj1sep5tZt63PwFSBDNc5oRLGm416YBRIMEkyJON13z9rMthFBaZDO0zXVrd6WF
L7UCToEmEiWpqHqaWS3ec1YOvO7p2G+mwCvR4dQXsl2fEBXRp7YnE6Q3bUBIAPDisA3GQBeu7Vxa
Vl4Sx1x9yihi/95EDInoAdYyDku38o3jgVw7JyszUe+0KljhE0h2VdPLeA0pcHR1GiGzmPT/weoO
MpECmr1gXjt7H0Fb998BdtiKaN1K690Ciggt5c3KsIWyERFMv8+1Y74uJh6je3UUU3GtewUIY6/7
ZEerKME18jeTbruaSOQPf8SJFy1Z5dvIwVRGdb4EEF2LQuq1vvtelkwt5gHcBp+jvP6LPsO9IVfr
CmBmNnguuLlLkmFovl31rHgMX5wdOJ8NKIsqZWWZpd5ovq4FbPXCCZd2UEahsmGGa3gdC5CjBljV
tb5sj7mq3PP7OhuxDW/bxAZbt43dqdLP4ndPttf8P412sHSrYISZwwXGJpfKKdbsou37F77V5VSw
PqSrS42ovtaHFPW/62gfgtXkKgJd4gR8IkzfQmbkbnnvFPy0bLcpNjV8k++6b3Fpfnm91AlNWrP9
+wInLZ7gKwrYtkl/sL3fi9n1QJARJVV7y7oMGmxKJPJjZ5OZq4thvGqKXP2A0WbPXKj4vpcevWI6
M4D7ePmAMAGIncAp6br2S47axgn5KJthlYRh8qGswnFdscOl5njP9RcWDz8yFeFupzauy4ybcUaJ
QiFMuTduKBrynIunB4p3KYR0BhHmbxjtjlV2SuuH7P+zgdi8nJXcukurO4CyhG9dYduISR/tAAPG
n9DNkoUcrpNlQR4jdBToofpmSFuA9caS7jqfne3Zc2dV4P3IMxgJ7C9KH2K0Gyw93fg7aDSPcrqw
2Y52H9/FV4e6rRtQoiSXv1c51Rra0NFxb00dh7YhsSQx/5fwUhCurvfGKCenghxW0/tCoVRec8i3
gykdI9dnFxz9JK+SGMQBW5bPsXpkEy+5kWNvgBz0vU57sfuNrnzkXUkgEBcfdg3er6d0HkxrViVI
gJbf18mxpq5xb6G3NxSODAh76kD8MY4UaRsFX5Zc6r67VW7SN4Oqju788BLpQ3NTHo08Xort5K0S
89Ry+Tn3ab2TSdOmq7TbrHfScxru7aYsuGe7BnW0BXn5BFfKLMH7bIyqJ+aXDUsShfdbkNnpah3W
pCLL9D+ZYr3h3Wu3lQC/D3eKuyQ8bMVvcj8Ay3Q694B5isl5PJdu62BfpqjI7oaHGJE5De4qhd7o
NwMusmy8pErVHLJDddX29teUu5KCUY6CGASrQBrvmMjavV3N54P+mwOjjNSXF6qYKsoO/OXu0Osq
j6N1WblRxxdae6oKb3v1cZ4p2zzkHnzTRFLXl3rV4p3g2nYqDsCSgCIgArnV5KFnbmvEGkJWD5VR
WFocnkmJdZN8tQKWdz0OP1wUqCZnEpJP4k2ddxsxqdnaKLFvjGzvHAf9oMhxFIxmXXTa5FC0YUcX
78pGcFaFUyXqp9ezuYDp9D8yvYv7vp70v9HqlIp4KSpN7b05H3TugykLYr6AplqTxirh2354gktd
FDlDSp1AiC2S8+AHYexlTiALC51fvu8m8BGNi5GXiadxttfvyI6ziTmfunDKe4dpV8ijt7Q5TnwU
HUx327hpiQ77/b1+ACdwZtK7vVRPXh/pjYMosXXEDiJ66ImjAYkpJh3yotaU0p7+CddBgGQgPC02
ScRhOSUMQRdXKMXEEZWVK3wiDwIU0uBU0qgUjScEG/clN7Ss2TGRBh/sWQEW8H3MQ82PCPRM1aK5
xlK6FZt851g0hWPTj9xGzKVtE2Z/jAa/DEbk/odKy1dgnsOKLMn3WH0lhIB9/YNl2yTzhI5xisdU
tONIRMkmSDjUtJ+o648nun0XJrE+2uGRzfv+4Q6tFh/wP0Ip9lez0vhBJ2ZWev2Fg1b4PMpgzYHX
HqRGUpLkfWEyuYqOyb96IAa5ZhrpVnMTdpFKA5fXP87GLJTmhKbcaP/nfiD6XeiyigLXS3OB17Hm
j/h8X5TmpHxz6aCP/s8KxT89kuSqMdeXUgPaUCWA8VH9ffxrfjCuPSGZbE7RLN+DQ4xoGxc5nJtO
xczSrIJ1LyMsJTMWkoRWDHwWXcbDT+vd8ls6tOP8xKu8YotMI/9C5xo2xyukjOnYwhJcEXlvlVG5
P/oEYRexD5AW2EE8L+KhPPNwXZC3vaXulxh2joWaMWM4I+nNmGNbC8dC9dO4BV0rUKRCk1anrnCg
6JH88fuyC5Bx15M6quSEgzOIawse8uoi/CYPCWyjakOT5GjVmUW+xV1hYIephPunRV3dr0eqz4jR
cjvCzWupUGqmmJLkVTtj6h1ry3UeTD631zixKVK89PL0l2280qGzYu47OJ64Q1vFWEQgw05uy2lq
xYlNn6rFrtuFh5ABqAUEkHDSxQSnuGOVoPT0/AWuhkBvqyc5wmfPR2myGsI3QPsNIsSPjutNGvBN
GrAYp+gay3JcoUVWirGA2yQDfhQ9i91+6IMprVdBT2iGeLcyW9RRfzazMzC5fOkArN+rCA3xi/Mb
xIwlI0BL1gVhKZ2OjtVjNjRo8Lve47Glv3rDQzblOhFGQq6PjNN2I+P7wNGI00Q7/E0PiV8K2X3S
lWlYiMxnCu/YW6tYNc8JH9J5FNfkx42POXu+wGCc1dzpo/lrj2k8Qw/PDHKc0yCSZuctEud7Wkha
Xiw6ls41+6k1U59JhOq7vJ7NA83M78sSd9nbeFJfL6q4ZK73V12Ca78LRSVznOG7CwMqmHAL58Lu
9bmJa8mxH2i4sbYiHqPQYecavWiJOXmipk3+Qu0MoIRNRCtrr8ASWMK1HJLyMkTqRZz+drzFzE4H
i4rNv2yFXwfcEdQo3rw09w5YD60cV4FyfWQe+cuqPITUsCaffUGzcEPoEd8DoUOv4oLGoEMJSz/E
rtL3UJo+Jm48Zdb+0igf8zhLCx8rqyUcHOw0/m3yziP/fN954G8tPATW/OUWvRSrZz2W6M3d+mVM
cRWmqFyYg/qn1f5e9HSGQeKgJpq53q/9lXO6qU9VXUCtiESLrnCY7DX764el/Ol+XTgYjVul1JoE
i037hSlxJmnhq73eNww8LRivEw2/ECyp67ovFl85QFPcxG+6VctK/MBZ/3le3Zs2O9X4qkNrKqWj
vUU+9gEgoybE6af9ZjmrM5xX/3YZrdahxcqIwu9CefPwqunkYpVstTEygrsvKS42vXNQmsjqEaeH
JGp+u/e3EYYwVomod/Rt8RaAV13Z34H4TFrtBcg04G+JTvCxUUO0WjJAakpTNTTZWrKu1PiQX/eG
l/yO/C/t1L1sYs79VUcNdSPnO1B1MBeqq9PADdRQqxLR3YBwzJJwevnnmKWCcs2nP6bQ8ZPlGEsA
pju3nMxlq5WxlHu4gW1PerydESpIDh3XnNvNgIvYcqQk52O17W6q5BMITWuMDCPlkI9TO8P94H5g
qz46L79a/eJX3Bs0wR8Ve/uVCJ7rsBkMpKZLpuxf1xhuNuURImG0MnhiClvw4wFC6ggeA5fnt0rU
Meq1vLt5401nQPAIh0ZP8/+a5BcVyix+/u3SV8yUlHoVYu4GBZaiybxuduQE7xXNTwbuUfdPBrLK
YnOn9OBN9gFOnsywbQNaW8rIW8kdidVYwfP9lheUjS+Yb6w0vGyWGqa4TwWDnhfpClz56XwgxnR9
WQSX6lr46jZMCqoTtdOcpH0E5DgOHfnwvSltA5O1ygHSIfNzWFIu/xqokLHPX5CXunZfLeBvEewK
UfeUvivDx1yhtjK7vVEPkswcBjkT/qSWR59LJ2wAtNGwqF+o+11OQW45ZE+I/fmmwXmJI81y3SqJ
lhRLbackIDJ4o+IaorXIQTxBXgLlotBEnUn6UqzixdIZcr/PLP7f1Syb/RXbb4GOte+iIRV869+d
2sGmNGl1T+mcHWFVc0ZfBm+TZW7mb+hvfVZuhHQirgZpGL79vglXME7SCx+d6bMvf446OG+G+Wbz
Ot4xMBMXB9D9AvWC29J40QBaIfYm80zqQeb4H+QAk+G/5y+tsppPzae9KyjKLUX1dwCndlfkg8JE
xH3eVYDfqw8u47X5me3kZaVzZrX+LWLrCm492jX08WRnwPsOqZKMywoZ4l3akyilvFosiCKRM2jw
TyslsoHadBNnzTqqaEfeccXZWjg+wS31NMJ8VNkevkvdoboRRwxt5Fu/mLykBvBrBE61J+YsuIea
s6hnWh0rxNSb0wKmvtd1Gbm+dZF0eI7iBuzWLDdKxCmqI3ogXN1SYFCI3UJZLg+in4k6Anxjq3N6
Rd5ky/C9XH0Q7KONg3qZw8qo8hsoYcjwxPZf1rSXxkvb6RoKYDHO8WNQqT1In3G6IFyVjxaJaYw7
SH1sHhZR25+sBxq8ooEK0jO45BoEVDEpJeGc+tBHp+EsUxJeWrXL2pHSrlbTSKsZKvFXl/mlPRhq
cM+Rvcl9WjMqA8WNdvtiYEOocQvGjLGv9Y+g9f2XhYPOdAzFUFjWFzgGro2SG6HYgNUWfJn+Z1rS
XHB1mbxvz7XMdHb3Agw5gmVpNFvr1mUAd3IoqGthWr2Rd4mJ35phgmtA4vbKGwoI41TYo8Cf9zBK
Dy70m8uCFkYt/WIzvUCE2TJlLFBUSpT+LzmhUKNAxbTkVuAQsseUrAg6KMIHgkBpQxk56X4hti7B
L/JiTeNNsLjmIoqV5xwRx6wi+xaJrhGqsZoeuzybWAw3qKHsbIovRKr7yXAeVuQmpfi5sAhR4g0M
W56HZkc1ZBAL4RX/lCdhOpRkmz2Wgpvc5WzEftpn9VTt25hwc2dWhFjAEhIO6co/rTgoXl/0NwIr
XZvaGodVTGvGkfdWCuw1LnwUuLgs2U+RHwcKP0AkZ4zqH7zIgDKqVAoTiZsupTvpqVVP5LtplWne
W4fEvJ7S8HCqy0OiFP698TC8s5rF0WPvwWc/huDH5o+QBLzCykDoGpFad67KfwlzRIm5XfpP0XxJ
GP42DJ+/BzgFhqbugKVFoWqM0x6JSVallRpq/6QIGgIXt9fLQiTnGDOAkpoo6iWHQTqNhj4KWfbr
P+FziHNn1/Yxb0aiUDx0wYjXD86vetXQlK/90wJjCHfp9qrnrQD/IGbnIAQfbQM02/ON9SlaqjBG
Fshb2sDCLty/VST0yo6ZG9Yxe8SNgPYM8537yRkWb/K4lBFkQTHH0J79PdL52BkZUIGn1BMvuGwJ
7iUDin5n4fTfPhRtiiiqohgxWDow71zPUMs4VCGnUvjOdt3+2OE5BN1iEiJqlVUKexmTY71Un895
iSdhOISW2ps9dJIJMZsPw3BJ//sMKwrEau+0ezRGY+yJhY74/BFnL0dcR9Jm4xPgYmIm/CTcZlSQ
NxZ/xw+dqxosOlELgcqN80Fl7FPTk+TkfJjw5chq3Lcwn2j3p2ID8DJ+7TwZ0ePtyz0fbmp6Iwdo
GwbuYdmBdifvFWFGYtnQsUwRkJFy5um0+GfyMmFkm3bA7q0voZzSP9+I7cFcWDQSPAfY6G/NwUL4
mtmHGpk1e4PrCbYq3jWG/fK/FlLuPMh7qaHkkisZf6cYS83pV53W1dBZphbCJk/xCDYRkkB/9Nzs
/Zx2Bm58JfeGrmZgwe8YZBuxaKgrlpdXBR6lP6asTscwm/OqWaBD5o8+QgaSRxLplPvmS7DOjfAX
uOow4+K9gWILw3lZMdPGomwGxEhOSayxjHxcKg03rQ7dsza5zdqtf7SJoilBZ6H1+Gr6Nc4kXDiJ
TdsZB6Ui42672GnI+n/mNgg7DI4mztwS6Q0eTz6opCCDcOweH/CxkuEydueFHs+po+id8fVgb87c
IoAhX6EbtNwZH9W0d7R6Kdk12dFNKF9O/YirqAvNa3og5Bxt7bn+wExk/FJVlUP7s8zkRtiU1gRD
2FiGu08+aOmzE2uGITVwPQ+mwaC8eDrVyCp183fk5o829KxmS5H8BGCEVu4JRhr2+MxlLWKbSXaC
bYlJ/DhBID5W5tptAwayEwqxIoqjeOmL37KDqNGKsnJd11gHX8RnHKVAenJ146r/pQNrWd2heacG
X/9H5GN5oka2gw5o6PGb6KWD/pybnE3c3WMwOuLToWDdlJDQao108R+qEMU6hymrJAgUUc+PAESX
eyAASQZ0Kz4rAJY3dYg0U3jh3nO1lTzTYKmROXIbVIqyYs44ouucCJXUEsHCs5TNv8ugkLDPuPvT
Ys5wDOc9KEhMuFEBNdrhP4G4Aq965G05MPT0j2FgdD+rOOBklJ/1cLq0DTE0kgnm8SpOXrUE0SD/
/Z/gA2N4jkgkgM19vjZbp9kpW8XmBLBPnXBCNecRGmXYmb8dPpJwLBD1dab3KC9Ti0mQaTJt/R6p
hE4s3PDSK3GgwR33d1+8L+gqLmJvw25BuFvn56uiP2tBVobkws12jnfooG0+hDQEfZsuKGVHTRBh
U4Zb5yk9zg6Rx6+C9sPA2YjTqHUsrl/upBm8oRGugQ661AhAe4+jip/f97xCFQEaE7aeeIwN+LlL
aXuDlYnvMA34BmnPtWBsT0koQ2m3uEETg1TKTXST8mZR9HRVN4lAFE7iiGb9/WXsT7yPYvk+wP+K
WeeobiNNyU5M9RD14Q+BXjPaStXw7vth9EPcziW3fFPC+fZaLohbL1Laot2SQHBYUpQF2S0dtyDY
0GCrCgSrXhWlznJRp4UgWxzyOA3vDFQt3lORVA3dGZZ2nkI80ivgqreaoC8DoBbq5DtlMx/5+zN/
01sNQiOYqnd548uvqt2FDWsd//nPXZmYfJjk6hLabQJm71ao8cQmM6YTDwn7yclWJKS3CEXlOGLn
zbzmrSCa0PQuNMG4zIReYk1Y7Yp7ZFHvHDWbybJyoI3x5sY3bSyVt40rp1oUNCyss+D5NBD8YTVo
zlzFBOGCLNNl1/UgQbz6IldJPyI7qzz1lyqjxwwKqSH85TZ8/ERhGtT52j9HkkqSgUv3OK5RFI7z
jO885F0OS4GBXSwZ4k3td1h2QfT3ZqNe6CliU3fTHaALckkIIjSSX5vN0zFbarQA57XkG9YVCj3f
M1uUe8e56GvvxD/Ye2ScSf3JVSk7enQyupGnIIGxvmTs0c69vBAsTavz7kMkWBKLfO7ekazqf/BX
sXc81+Gd+kFQYUROF2cd8dxFdH5j9NWwwtkRuYwMatZ8IOukImi4Mxzot6WPjmicce6SPIkci1nZ
1vFKFFNQM1pEGnfKao8y4X7GlppOT3mIXRzWvrsR8UEliLBvN+wRCRNRLW9G02GKckN8dCvAxDxh
cYNrhvO2hYkeq2pUTzTQNEgcPOk61LByVIsqOiwUNwWF0AUMX3MFN7w+11/qJTruDfmf6XrnDHn8
ChOt8h6/nbUl2uvLb7AdBsQG7Rkb2TBhEV9P1lnDOyOYBRjPwBA4c5ZqT7Vvz7wkewRi3BTcAgdA
fLqSeCel5Hfk4teltRvFWB3fhvyl/F7Q2pBeAuNDbbYe87leYTJb0ugFldKxL9vMuiPFwmY39Zh6
X0+76SOrU1SPaEca35R2IAQQqxIUY2mC60QxwHAvDPzzZSOXsFGOhxczJYrb3pcnp8nRAOi5Vcvg
HadPdDhOsvTwYAgnvwGHeOzVe8SjeACCZp7v7N9tfG2krKci/A5rf2grju8YuxMX3rwmXrWS0Q1Q
do2yFBuXIqE98HI5dLP1bzty+jlCTsUKNSAOxe9KuU1GPuHFEDdhqW+3ZJaT4Umehq0LydX37zH5
fzrrQ99rbOCBClYPqRJ3YY+ImOO4Hx/weuJoCCOyLEyeFd3GWmUdxU87K9PDofbVsy61Xso2DbCU
gex1R0bwjtc+lbdSNgBAKX38ddphr4OYK80VmhC3Zs29bvHp0jMflkDGDs0P+xt7FMKu6+Cu67U9
kbCHS46VP5sAoNDBQsR3m8UpmbCjV0V5o/aa1YIphCPuLqX4ZTpoIjkxOVZaRYUOGcYe65+GGrcC
qcoNzerEbYZNMXMuIMM+4eqPOzDVZSQpMrxkQhY/qSYx07NwDd0ku8UZ/YbqSMFwco2TNwQuTqol
P8fqXHCPTe8WElSX6mP3SwQfdL75jsBblXBSw4VVHNHD6Tg22D/PGTCWzzeG6D6aoHX05hAyIiU6
ERUuTGPndLDpIm5adKfiquWaO/XOXtFLodjDnhHIyaiR46NxEezSKcNgfHl1HVlpQYgQkdeNiTQE
nHZRUOTA0rt8/AXHsmYSRs8Lj803vDW/I5feVmy7wAo8SCj70ZonI37pEF0Fz2ves6vK+XOzSaAZ
OE63I1LZ9hD5XxetjKd1pPWzZ2jmMBfm0HRe/S79T5Gct48OLUFH9VvxGqITbn7WrqKWUHOdd4e+
+s2ctW+MGFAnwuzjLHol1Cfk+rfqpnocYZ8AbN6EyP3D7PmAeCJ7l8TxsUlij3ZgwJSkCtS9pBnk
2o8Fd7txmVMcM1vPITGcYW94K9LqTq2RlsAvq9KO2VPoQqyHS2oxPbhj7OWhpTpLmeUlZi+42lEk
4TVmKLWeOWyhUpPlo1f8ppNDNf8Emk2Vl/tMGtiR84SLOLqyiUumWjLbJa3uwn70XU8D2V3bglff
BRG2aamTpB08tu5Wl7mZ0JkMXfYhESafcllq9qHstxfLpj5ds6t5DnZ5QK1cS/p/678fxUn4wyS0
SO451Q2cllirYGOBbeBfzwu19uo0Mo0z7gxOtWK19w/BWFAppvc30fBb8cUL5a07V9ADNME8g3wU
+xmKLgQ4HdwwTM1Qqnp3E84Y83TNwMrgIihFUm2bFZ2CyBgEPTue219NNsEjQmLbnbncZshaC4ZG
XPUrgLRBirpUU1463lYInp6rWfV+o2tGb0t3O7bQiZk3BI9Xx+fC4dT+gFCwTZ6/2z04GNbtyjpR
wRRvtx3Jyk5CML84a11cQH7iO/Wfqcz4/htdQCmA3klJGPTy8h9gxN0rdqJNMADIPj3y5Lx3LLAU
TJler91FaK04Jl+gpGZvfGud7LkyEyerP+eWUplPrGRUSsMF1xPAHyyLpw9uvSCoT3iGuyQP4aRp
G6wpArhk9LpeWmarrr4z64tVf9SiiaF2oMpOfyUuVFom5lN2EGQKXYsTJcPfo9SSeUQuH1tk17oA
4RsE9NTlqWMerfBRbqZDgyqUN3o0RqQzrXX3xYJ4xDSzzsUXS9G+tuWFgU+a+R/YufZgr7FjteHe
dItFBrRePwQFtMJKbqESWz2+jnwZqDXwUYWQotLI1I6tXscStkseN4oHZ2QypDySh+Ptmz3xyhi3
fu5ANXdakLqyS6C+GTO0Ct7wh4xRbn+k3ubxZfSVD6AP2sqZoSDR4s+jOwWIHCVUqJcQ93co6Dh7
Bo7qdpU0Im0YqCBEdYw3qQjBVnXwqQ0cmEe+rbJnXBASFaLt7KepfJzobihvjWPbf6CgB+JmFwNS
maMnxnTevq6S5ax7KaFNbJ1+yG4D2lyuCQkHBYSc6yiDmMvDs/eFTogetT+vwVlZZ8Tl/cuhYN91
jA6Gsf/dGnHbjY2iVoRE1HjbohCRIl8e5WmIAnMRNonSbIw65BlS10p5DmAtUdA1W8UYztka6K7G
4V1W5GSIlLn3gZ/xF7t3+hmMS8e9OSIM65Fwer6nWKmPlf7GMSlTxmxtOUkljFXzqV/jQaGWrTyk
n0CVXolVmlN6yI/JDwbIgE0jrpUFMUkFoHZXaUL4G8vqArngla099kD0QupG/7b5KYG1xBy5aNW7
46vATcPEEul/YUofjCjjhZXrPJ65Kvs3IVoyH0PkjV7eLB0xCB2JpA+GBiiy7j4H69n4RRkvnMkn
9wbe2z2lwM+9PXy97foOm8mDZ6pEtUDSCBWXX4mha41Xvwfks9YXjkKHW+SbtD/MF+jexpOpds1J
2/FUhqrBt2iYYd6a19Vl086L9iZalhj9Wl5n7Bq7hNOFv+S8hN0FQkuQujloYRz9cQ0fPQWb/8yF
LJMH9VDpBNP3NBogglJTjbTW+yk0VzzKz8JfdgO4ppX0O8S5gsYcUzMoD2Pzv0/BdbeckLXzJ8u0
Tiy5e/r/FqH3apGwbg0y3TOZYwQ9v9KtUkP+//UilDvEdROwAImGKjOz/nHKo6C1H/RdWlLu/6xt
KwJKqv3JNDyJ0bcwPIUYgj9ZJMdzb79MI0+hnXnrW1Q4WbI3B8l3CtLFI7F7QZfa32IzjCtsQaMe
za4KxPo9gCa86db8W3coXfqXTO8pkKnU3s1SnWIKuh/LK2il6Z/Hc4gTNEmGZIJj9tqSvoaj+hPN
PkpKDOnf0K7PqyGGzRQLckXSPTH8LULdaMIQCmZKwbirr9p1CdZqaIKBooUGWrOn3YNkxahdq+ye
+MStfkJtJ5XYw7Dq73J9VmCNtjpycjTPOhbZ+vMlF8RiQHb5Lxfb2RTgbjjP7IKxjqlx3DfjkV1c
bTJO/Gjri6c6x02U1Vbk8queIuC0M4gXsu9hg8tpDilFR7CtOsBYhGjsyLzJg8ebycQ1SSxSZZeR
5NWTqedJarXJn6soJ3rMTUD0AhqGuuk8gxMYtMt3Tdh4+wGDSQ2QEfzfPFRv1cBGGolYWn2q9BnY
D7IB/T70V48PwRjvtbM2ue0b04gVJSJsmsY/RWU9zQhNjGNKsBL4HD46HK/pxTHXwyw+Fj4/gktd
21L9XDKV5e6W1CzV+VaZ+oLAh+UG5voTOobl2MWAUF3Sw5HVdN1+IpIBvxQo+dNqVpO+6g5oWOoa
LU8HcrD+241C7CTICFCV/+5jBrFb8DoVpSswfwIFS8z0H651yXpkltqSGDCGKgkeW+pDQzijkFQw
MGa36zuEKuC9lkZ20ecdhLmYsFvr3u2Fyw/Knbp4KsO8vlVkqPN9igYy/ZA9ysOPa1vJMvFFJzlo
zwxoVs1gEHso2Lo/rcSnfXHa0d9jsO1nRY7L8IxuJgtHQUAmxGA5LXj6YonzBvamTDRIlW/KhE/b
2aLgyN4VHPp+bwF6Fz0rGHboMyhDpb9Qs/xZAUidXzlp8Fq7UUtLtAjOEtqL+f2TaUPU7k9tWEN8
e1Zld8EMnxxL02cwj0yxZnwoG8HntLPpZLjm9nl8mgAS2r8OdMLnyliA909eN+PjNbezF3deNErc
pvq3PJ74YDBVxxyGRy+x+xWJwLRo7aaUY6jMXZa/kDc6XIg0l9uBsOPFj9KOnvuyFg3HTVZwkUH6
Npqm26SU7eU7GhZEyCPXpKa2UqUsXWDnCFr8+r7viEJ2+CyVlzXSucyDePWonotEhe3CgpxSWYL0
K5InFeHqmDNuLRBL1yl1GXluwmJjr9crTLYuciRu8XjVE7TCHKcoIQlxWiMDXzirhGoRDo+XCASL
neFcuS8iDFzGTEx4S/aW61MUnxc/fDkVG+KAZbsTZwG66mudiE6vsW7b/ebrTF62sLgq7FuQzmCV
rRxkw5qCgIiLVUBrMQoXIU5mAHcPioT3mjBaJ3kxH0vXg7BLbTg0rkL9wqK0Hz/4rUZqEHKMovEE
pTLbGwuniF0K1w3O8XgjFoJ5lehzrzuYEbrEByIOYXYmS7KFp4mJGVAgnxwQm4b4pU+gntQlOyZO
fzRrjE1tesXCnCPDJW6e7l2z85D9QVu+6x2vGBXfHz7iLD7c3ivQqnRwhkdg/fwVzTjvohJnP1jP
XzZ0lGvf84K7Rryw4ZwIwCLuC4J0Ucpqpou9zdgxRgdhWClULeaU6hQ5OrcpqjniT25iPGTvAEbM
gKnBBvG4aYMotezeuEXtcoFvVAmEbuJZGjgF10qutpWR3GipMPwRvBOjCOKMxwONNiJ3+omVMp9D
/EYRZhbC2uIKuKmqfSLDpjlOw/RbQQNEgcuHQAUB5ts5MyWxKSFLJv+L7NZsInX26vqpnsAzNfy/
UtXEus5K84uSfCj/jUXXrqYOt3jR8IW2MSyt7lgGmgnK4Fj327IIh7IkKMlbFf8kgP6daq7yc1LZ
uGvowFkkNu69lNFm3jmBpiv2tMDc/j9hww0FlVXLzoygLofWKujvIa3pM+dlhnLJCcVWYhRHfcHD
Wv++LEqGNVZWD0RB/4ivOSlEVjjMx1lM/fDbDb5zqThFmy5x1DSCJnFHevQe82+stprbBFwdpSu4
VAyLPS7Ys0BI78YTWgtcvEXBq4kRcl+5pmjwj0jmcokvSlEgBIxI5It2vLWgjipzGX6hYX4BvcjD
oE6VHkhFn2xSqb7Pg3Z+0r7t/WAuTSr6BCRDX1Wr6fvU1HEph7Wc8BuTkuh664HqNBIoPv3BItNt
bB32NAQN2EEk3UanXgAzDX9giGPlzvLUmO02+CbI7mKvktuiQSCeRngzofCrW8k5KVK/8Idj9ynf
tUb5q4PtAgoWunHbdVuttdJ7TCLFQoSYr4xS7uPLs+a1uAjSjYorILJdeemdK+MhDlB+IUXlSi7f
ptaDV20FjKDlPhed3oPb//t4st3+37M/JDHOkKuSzi0kk4SGJQ+HQSYFTI6AaJSkY9z70UFp5Nhb
9fsgt3XY7NxU/SC0X/A62ibHdTxnqJxBxPawTQjyrIZY9lSjlkk6CRye6P7N7DTLHSV1lh2sBaQo
3VFQuH1/1SO7QR3Ne9Sna6Fv38HY8SMbTLNVmU4nNdcg5Gtbir0LptRT4+MVK9CZ2NFmaWPjA/hs
bpWmXuaxGFwDevskdNrBra2mMRhxntTvXTHz79tfnH4L73E+cLNgbX6vhwpLJamkV40IV4f7I3nM
h34OqPwoutkVHugmlGEuI1RteFaI+cgf/66Nx5L84EKGqp0RvHSuSHhoR18kaQOdh4r4OFle3C9d
eiyamSSQHNd6Jl6RiUdY5ZElwZDH3Hs9TkpClMSkDOw3u7GK0D/trnDlN78l63qiskiUKhSPHFOn
TRepotNCpLPoNLTrCcZZulrC6/2KePBOlY7E+XDGZboMIZsZy1X52RLa3kTyQdCdglnGSz+uaKBr
86p6mn58NmzDmkm2nNI7vKj29ZDlmXjIHNowAuzX0hgPxS22jgdwZ3IUxvk+yjiJ/Bh6c0kngzXV
voL4ujpWI7jOM6a4Z+nmGlWGhJsInWTvKy9ykgx7R5jHILBya5sAGFIcJMsg5sbMlBrbY/94hylm
+xUUPkn6NJAuf3vzgI66OGfNyaOLUgI7jnITEEmExhb8QfcjxTxQ04ZS9PzZCIL+E4QiZ+eCXlbj
gt7w8XbRCaHRVis8GvEePqPpTLJbQS9YiaN1dPzyqcObL7+/Tt9GPPJLdx9bFu5SvWd/Saa57Idn
Aa1k6DrD+9sSShtQAmZcCrWAp5xREfcRlpIVKZuG6Nn40BpPaF+kDZurNZbRriu8ay142P9hIeuj
IxSfiLio2EFqAzjbJg4La+E2DMtlFs0XUxW2+bEva6C072QaW9MCP6wSwLvfJKa8oEV1Yot5b7vS
ZU5qllUPw/Hk0hFACxi1n298Xm2G3GMP0tLgkUkiS3dciE2jHiedyfxTN/MAxi+vOrWFmAspDk7A
7HXxsHiCEwzX8We/ON5u4EeOsdIxtzZ3/uB8ZkPgH6KMZdFtWG6DaRuHW856HMBxK9x9iU3ZvT7S
h8MvGTszJ4bfZ6+zY3W63qZstZA3ypHubu3kr5PKxPkHl6hGiHL1Cq6yKG1XRV/OQVabNUunvcze
PWGyEtHMlag9ZXc/4vNH25W/cduQcL2E4fUN27OVBbwmmLMKf5zLldjKUbEjPkjjCvHRrNjJAhF1
21z6OTuPrCYVK8JaLcitJSaZ4IH689pDNM/HGEbS7DDluOsPS6E6mBRNQ2obsJ9TmKckn9OLOw4n
rmJ5q/5FnfsVdrzEpZbKFSMXUGB1jOuwBgHP7lWEGmjOrM8wnW9GDiP8EI9q4+TCRTQBb10AXESW
D1wmnIP/wF5Ig5IfK8oDllPuX46d+1PkFcbPt21SEUefxveJQzCXB0yeL9/0bNZTutu6x4HSWlrB
yx1qShGz/5fbjsD2JVjDQ9ityzFex8Dx5qg1++Oke+ib3KtXX5J65arGRR7aOyUQR0J5zlo/80hw
EA/9a+y0LhSVy19wpP/4OgKm/BNSKies9xPg3fZTMjvMITM8I2RLQ77voHReRjPkpTZTtHZo01Wg
npP9etvdyHNUBfRJviJWbhIQ6bbWZ7hr7b3FpfC8R2oC54UZNGqX52nOFGn88hvTfkBFp5SJd7nW
Vhjm12mF2Dgp5Vi0JpZOZlKwou7LECgboccRoNL2ILy6XRlc17/uXJploZnFX+X6mKehSakGMYvR
WdWRawr2YIXjMcztRAWaUL7Nul4MiTkyYHPT+CMoilmTelOs/P1JT1oTkICjFpXIw9PQz1YR2OCA
z2dvxBvuJTPltJer/9NQQi2KZMf0bKHJTxwFT68sWZfi//Zexg95v5dTA/c3IqHwLThaXaeiZpdt
FNX7xPXzF/myRDi4BKjYMRGqyKYTTdqVed4Bqo5ckfImTmAPOVnHV9htu8qop13W4Ggs1mTdkkhi
kGx/q5+KYt8KT+z29I/rNRVibUFf44oG/qG8p6Q+B4WSOP40BOtwF+Mgjel5eMqdtAdkfH7x5yO2
bG2RZ7G6+oNkDnd483hKwi539iwOiUEvnH8G1gq646W5K6dgzmHRyoysni4F53zUF5xMs9heyeFA
QW//lnir+RQ2GMjaA+R7YtQKJ8lJMvqio1RVKIbY1RYMronMjTXE998/5qfSi8IJ1RARE75ngAeK
8AQ+utL9XT3ch4cH+l7m5Ofpurrz5NMJrorSqwRZet3kQ0IFwIVNMHo1g+KGQ3vvWwdTtrJ3aIrM
+q+EJXSD8Z4Bjnx3eCGs4d1so9f7t9FVDCPiHzv8skNSjDOwva3oHMvd6dQsDgXdf4vVC8ejXw/1
19dbv72UpvjWl/TNeRPTP+gtP34YG5bGnXaz0ZuM5RQnA0OHi2hlQT5nPRTBbaR60z3sQR4wiOyw
JPZ7naGaPnYZXKw0ii1QabCaJPevzd1sG+WPp1L801spXHVoiXgWdhRBZOG3MA8n8/Lwg7/9TDK5
yrBtqmrKnG5QrC+yM8Qikr6p318PetgKtol6PpucS5tNaSsWUOBdX/bX0tUIFjIWZXwN5jX+b7vm
KAGjds91WctZTUmq8AxKTbuIQkOhzViNkNGd6QP7b7aKPyKs/yuSLy6KX2pWa1u/7clwO/NDZzfw
yT6iWf2G49pO4MwuhTgyYIDDkx1e3LtByIsDvvaXNIf3VfwTCzu/OBXHgwLAlNGXddwxy2hjy6+L
1n0GES3ScrbzEClCFTCd+6lNjFYmrSE33QrKaWxoX9gLj8tZXgxgLYMNkBcEDZBueD4ChNSZH1za
9Aolixjvy0IxFDIQet49StWF3pd9Fj3APuS89OtZPV3H7LqCFd5dzqR10coPyu7eIclBUJBXVoje
H4wrzAO41nYV/kPlNEwIRRhy42XcCAhqPCo9FIU+8xWLzS8bLTcSGllIi02+LcPHZqD2M4I5SeTR
xOQy0FUCOJtYs6vRDFJuFlKA9rihBhxYmq7/roB8BOFtc1XQpkLokRsvGmoNuiQqY+m7tySbProO
XPPHhE02fY0zTW9SUlfDjN9A8Lu8gbts98/trX3ExIa9jmSJ/lEBprO0yK1p20aFm2WuBKaQW0dS
HecT6R1xVqMPiZQ0dpLVbRmbZ94Mk0/BLLNpRYtuBFaDC4VnP7VKVACu27TCYo5kfPbCXSsxnypI
Co4SSlqCSwg+qD14z51UWquRecNPaQM/Wj0bkygLwkjvOjpSSSkvj48CV9mRRHp/UPdwAbjjyeTG
Z9cYNRREctXj9UiOvE+F+97dV1TAvQZg+Lbfu/jLo0XGwaDZkGfE4qJSgRejQX0pMsUVxUIefoTs
V0/vnvkHy+sKiRYJJQXAIvRYoTOI4op2/RFG0i5V0msY0d4/glApfwJ8iva0Yr/YHxBf0SmQwbSy
otUXQcl+gVwEWILOIeMNLKCk2b5qdZIqRR0tl77NzYfHy4gRqe3GwQJWCepbZtXfF/UDUVz4VBFS
jVudOAccgGV2uaIRslXKQ1qF8gxQuHP6RE6ksfQBxphd6bnxSRr2oMJpoxVwq8+wzyOGOsj8VcUz
i3Wr4qnHLVebC5rcogwap1HpvpbQg5AGfIaTe+B5mfLjmbZN2g3xHF3oh/vUUkuuWM5JgzzKLwlw
lwR/CaHzRZPnjvRPvrKppiYHBjnc42cxvRxlxGfjIgqXOdwKHFWMOtgSwHaGezEoPme6X86TdXuo
EjuXfEqdR7gMjMz5Sqkj7gsJrPtP2Z1W4K/zdR6Y25hKGLG0bzeumJqLzboQRhP1GS5n4cBWogG3
GcLmfI+foL4U6xybedEuvjo/jvB1JxxBJgmgi46VTq0s7G4XX+tTyVssDVL9LwylsGpQVwwrHUip
RI9fVpkD4L6APUKXeY1Qy1sExQYSKQzMa8baVBHvkIGKc3++B7y74HdGsyFyy29RlfZOu4Z0AgI9
re6doDtq+OTaSymlvPa8rwMURZIljb4wXqeittc9n1mvLoXZjAb7Et/ZbC3V1Nlam/32EUyroXzY
vHTyD/jJZ2dtjQGQduLP+clT8JEbjs754vTiURjD+WdRLxzn3WVEkfREwp2CZvrkZt00Iqzr1kBf
rePNEprnxyLgJ6TSIcj5EIioZVZhkOs0K0DMsYLQhb31nQM0RoVbtolzcxBNwztkNIJeR1XB4dsC
6ZPG/YhDBX/KU/rjuv8KoNep0YvyyaCy9epiLSkjGQTfQP7GKZX3guMPQMMcqaVA3ef5395zos82
U1V0wlRp6MpefBT4wYTPtLJC/ravjS4xT1bNyJJ2keKb1T02rGSpljmMOhFeQEia1hjg0/wCHWG4
OVVBjOWYtuDTluwD+6stOz4s4vK6bxu2WkRfFRBUPBW+0f4+cKG/X2/jDAhdaKZ4veZ9uEThtU4T
sll7QPzycu30aHhq22BQuDiLTExHHo1Ni+rMosiXrOFzq4IHKHNUSRNpqg5dy/+eLTD9S4uDC/ll
LqAR1xRhW0pQd+z0zUOgyJSLVtX1GhHaQAzuuDHzSXO54wm8caNnG9+8tCjT901gV5J36an67v4b
/jQZIrBqvLEebl3MSxKN5s0iNCnTByUkeTrQL+8+bKoPEOSH6RPsQxBrnLPXIUGJ+81RmG3QdO6W
TE6QztMx5Dezref1Aa0s7klUPyBlgBhD82GaQazAo01Ychkqp4m38c3jbWcGDjtVeJzox7fHLUJO
rBXMZ5MVlqY9jpe5Xc5IuAyAoFbT61Je3Li2dYOowkzaqpKm98acoWjNU6HH1teAQX3qWnc+JTFY
o/EwAvtPmhoCAIkCyAaFipU4K3vhd4nwm5LOCZCCgUVHBbkUsvKgFUJBch2Ln5UxulZb8vesmi2X
uKOT6cunZqoj2VGC3MwLDRBg2fpEuIbBNW5BErPz5G/dISQ/yE5lf0dZ/op2QfsxcI9mgF/xbK1F
3p+TL1Ra4JAfPWOxWz1xkefzAbf7zpPrtVZDPNcoAAi6XmW829wrNZ4l1xLvcHmUY5wE3sm6Zfou
f+9T8Rc3Dy5FWl67qJuqm2h9PFB59EDZX4SRHGEt0PnFOv8oWFmSvoNBBeIG/i5DvvUT7TZl1DfC
FB2PA+TDj90RExtSBcd3/PYHVz0qPo1dADtFWTYi1DzDHutDvN/wgAHEXI41XlZJRe5KzDXW2++6
qSXEsh0bzKvtx8tNU34UB21+AGFTT9hBCPqOs+SyCM5dD5h2rjnaYyXIll3j7AWvmRl6yj4efrku
HLhkZsWRLKycXYBC1ZaZ8897bGwiAUGwZVT3H9/A5INCykQK7zbo7RWna30Ul00mv4KpTOC3GQE7
OQNm+RsSYVr5W2xGWYxGefxcW/0WBdTWYKhUWA1sqQfNyx3LQvchhnsnJg/DBtzVOJNPebhL6Ead
7n4IgO3Dl/17ldIH8s4QTgM6iwaywGuFjESKJt9q9Ln4zMGvkvzJtWznFCWh1Q0FREMOm5/4sAu8
UfY0JxGrJP9+CYMSGAtROW3EcvliCT9Sf3lzOc3VmQ3O2sHjLW0zvJTPj884YS6xvA0wDUWmTImg
2Mn+9RYQEBs+6qd933ev5b3Grh1coN/DQPf4Xbr+JGRHS0TP68M4tC9YY67Ksc/y7WMMeDdBC6DS
JHRHKFPtpfK7iU0hudpKNTH8TYkCBBPs+lwr3VsiDhovOSuGMWIo1cwYtO+sw6XNjRS6B9yJd6QK
cfBcVOs48Ol22uS5L0MBgPoQIGrKHPVoiG5/L9/BvR9fk+5FJqGq+/5epH0TivjGZfo0gqsRLhSx
CUU8RwS9FwhHavb8azHQCJ7bDzie0/tLYqugPl20mjqA+ZFFDaHKjYOOeAp5AUkmoYrD8IjEwRE8
3BaHCxTkA6kzThM+bwlFC5UcFB2H8+rWnlrE+i7NDTkbKrAlfXCbyHV0LQfDoL3xeR1P1WOSW6ah
pvSlYEp1stfK3Llm9T0zUr1/Ebx46HwcGtLT2vg3564LhQoSu0E6kv1lb0ClMpiHu7uFCECW8IuD
dhe7Ra4r58wzweRfWwBmVOUgQ4C4d06eF8qWlmhrFeOu+HRvKnxLsrBvoJkOE2ClXuzwcGQhE93+
VfVbHfvu650igqjo4+d/Oz0NOZCesdoUt7m7AdBBElbkXIXcvFS3kcRWH/nVuTDWTGbChx56I0Cw
ubuqp56gdRSbtQKFbaRJI7yr5kcVxWUh2/8w81fISpcIO0SGby4NHCX/pQIr3RBqccprs4q+cz8b
vbs2qUYG+Hv0tVYWgyCmNrpIbKRgcew5yUBiWQ/GD3aaKF0foGvHecof8P9BuAv8zaoWJFzvSd4q
p5RCvNMrk35wSWzm973wdCQmRUfuLkjV3Op5Ov1pW7QQt88H0qpgH/nW4wlMiSky/kQWq3iBH61W
FpmKm/WP9mL+7gSJn1SVc79HtHk9BZK11C2aaRMqlD6sdR3jqN6IsWpa9L8K619TVKJPcsvGuUvw
50RuSo4MMEUihvrsJHDzSRs+En9U9kRNYdyCKIySzZu+hle4+Qs5G+xBE3lxRoEXChdcBQdTX5Rk
1Alrzh2OajQtxy1cPjNM0VWu9+xXeC0lOErzpekelrMZPBikfUqedCcOgMluxNpwqlA/3H2hVWS7
NYyWDPpELRolTDBomPTz4XQ7uUil9ru8DgFnBRy/rR818KUiSflX8LRVeGSe6Lw+2t/f3GYbi4Gm
Tdoo+kI9rviXlrVMNfpJj0oNaThOz07BCUxrFeg259b29bs+kO2VzYCaESAy6Q1ijpZY8TH9C7Dl
Qo3fBtxzf9iIuOOzyD7+qNoBznhmqPpvBaYtucOeYYhjJZYEcR9NEcJJcbg+HpDsBUH/mmYqk6H6
Y/K8EZaQzPQVfsGcGTghAfdCanPE6Zh8RwL+U2pniua8SwsfUO3m/uTtPoYDk32T4g+21wFvuG5N
jWtZ6zMreeRDhDpqGn0JxPwCDDcRa+ivs3xvC76GLZ3JUXurdbjQktGGECcaQtSE6FEK3Wp++oEl
dkCD5AejYmer5TO0rFKypdXWzXjAOkwypWt3xhzA+VrsLa8QUVu7g+WHNGf3/bXStDWWa9fFZcoC
9FrdG0ur/S0YS1l3hPdAU1pIbsS5bJSBrgvpg4b6wusXOk5nCzmPPkEsQRCgPR/tBr0nNRIvt7GH
Kkdwh+3KwZfSG+VkE9SCBZMT1d5UunlQWWGizrgdWbEJC8piJ1T0nYoqio/ymcpKdWAh5waYzcUT
l2OTjY8GEcY/Bw+GM9K0hWL0uab5E74kFQpTKcx4GT+ErMJdfvDK6rLFPkp/Iw3aJVTq3/UvDZ15
YoqM5yV7Vm2nW6+U/BFNCrtzJv421YIUFpkhuTodDCEQGiUaCVhwMtwEaQ0X7ErW1B4WC8xSpI9u
wem340q92s9iUUGy7YFmmpaupGYaPYV/+GLVDduz7caL1XJjoFhV56HIv8bNAyVJhwpZC/CTXGbu
8qHZWZtt9tQN7oydQtWWfmH0omVwIU1pQQIqWciMYsMyhMJ9S2GpZ7gVG4TE9CZ36GdtSyofWkCM
PaR1duOOZYQoQouB/tHyoIO+N+0VprULXthTkk4MYnkc3jtrg+w7bRxaA2Obo+u558eoDVY32A22
TfAMh7b8wxwH66Q21Ni+Lva1WUW3lUwE8sSFOB0lJ/cF47nfMUOaKQuOamgUZqG18/6oLQ8x/es0
YpaDCJQfOhAyHlCTWyuIyJTvV7fwnXdXMzGSMNs9aFhi3hX8SGkKc5Feth6UJ8Ax7+X3+U1wqLps
/h+AyzVYrEpbcNxs9Kv99mHxnWhUuEv0nTuF07GJyIKgiPoSRufTWggwB/mE+H+XxKvNTASa73IZ
1rvpNflxmDlHKm+7rY8jUIIYkuBpbBxTWBCMxTi7h2FDRVsoJioc2YBZPVExJE1dSPFBr9l3LdDR
K4GkvBuv+VbrLEe5ZXvWuDy9xL2LU5ZMjea8eGOB61z04ZEBrS9VF5p1No7x2FvpDCaIWGHYUPoz
LoNyMalXJjRwk/HFReDzYVc6Wz8QFiKifyDijWuomnOgXS+u9zX2g8wxmOawoLHiQ+0sMG3xkp74
36hODpoGvc0UVGO0wTfp+FSpVd9sku+XF7K4aJE5pkO1PAJOI5uVff8zM8Gcm66ygrlRPposYAsY
OHt4QLZE5Se6npWNkdS88FLdCV6A18sYb8yX8Bh6dJOW/qHaCphDgFqhJ/3EcQ0TPrzlyiU2d37G
zOPCX9SZfHifDnWF/r9AcL642omon37u+x46N4Fjq0QGZ7TMOKCR+ryNVfOymXLQRf3Dpkt9xfe0
EIO+Zv+MVUb05d7JWG/oR+8BdhDIGxdTx5E/eCmryf1sU/Q5smH0EzqUfLIRXocsc3dYTz91pDmF
1l0M9tyV7N4gMe6i8cv1n8pAFIs/Hhtyd++es56karGOQXOkUI0rsgoSQqJzBIcRG9uCVrLOb/sG
I+Ghwa3lDDfYtEDHpvrPT/6DBP4lYtlg3krZXJQYhN52nHaXkgfzgdVEL9uNF6u0+KDYjF0DSppf
QzAP8uNGhOjaMDE3pnUDZODoZVslQWTG1kfJh++NKLoNfcFwgcWNS5jhBLAklCTRVcJNx41FS4uh
4UhrdIKUo1lexJIzZE7jSs/ef3ekXZJCTkEnv4gAbjEVorIOjJ1pLOQ/OvBWzVGL2K4uFtLVnD6M
2CMYFt5z2Z6ZyQfu1D/JacQePENCkU2LQvdYAMYInyDQusb5kHh23YN5zBnckm/g5PWbmpn6fgKE
zoxPT6DzehLY3Ixsfn2ShVy6twj/IuKLBlczSi4NpxYk57yDHvaO1wcMIeIW+B3KO/EMvOYoZXrh
nRZhFy++6k+HEq0fU9mK/C0ExoC5HKRLZphfSu+QyVfmjR11CvAAv4dRR7ROdPeP1fGJPjtIg5rh
KNxBpJcRo/VGn5TR8la/Dvku2tRTBKzw/vwWJKA/EC+RVlifZFlFcCobDZHTc57b2nrGI05zKFxD
N9z70KUesj5W9exERT3nZfRkHeOU4yLE7bw3kVdjIQFX6vLkSb5NdTtV4qXQXD6sG/7rUbfQnr5F
s1JZJmaWlR53ZS+I90eVvwdWdf/luOWq+8SqQIg3xQO5zETbvsMgPvHus69nuj1SMaQz/4aAj4Oc
gHE7A4fnrQGTHkykXBOSI2EfSKFdTZYRh7xPTshUaAjjzNndAnRJEQT9qf69nsD/TG+PX10bL+pv
GOsKEe0SBmau4ZGnMs7okgXY4uAhLLpNyEXjmSgFvjxApKprC6t62f/obWNMK4yNZsco5C3lUnO1
s9FSQFoZpSEgpSCPbv0i0PiU4+IdaH+VkENruyU5cSR1W7tdVJbBk7nbEp+MCRgbgEl8DPQTnwnj
v+tfye5/NrDNxqaUvke2PXNgTuD4AjHTVYaDyh764m0OJek1t4SUmBpViWkxWXwtUU8YfPBEmppA
Va2BAd233JkGSjiOkz3jA5L1tsJx3noBfw54cQyfsn3X0wG8U/ERviEiSwIq/aaA7idxKAoIPDes
hltwCMKsDd+f2675zyJTIwW4p5BfoEqMQemma0eeuSzvLUHxyU0xUfQowy1OJqtbPM03IrqptcsY
3mH7ZD2G5oT0CiMAkvdYFv6DVe//44VzbzCDKbDSr6DQkliJldZ5ZVskO27efTz72IqHlfijo3EA
RKB40ACyq4JOZusoumwJLE3SD50QQ5JGlxP3uCjeoVtgfOGZenun9+40qVXpITEMXZGc97w9EbDK
EYYywMlEZE/Nj3v9yTs1CYQ+3kuUiPkgiS2EMVi0Et7tgcN/MFBOk3fdu27oBEHwcHA07M5ygFd8
RmGnMZSEUPJaX6ndx1vPOYPwEH5aDlh04bi2w8cxwKIz/IyMaG4/WWuQRlM2NtHP2XxjYV2K/jFq
YfZ3cw7dJZHfsupmkGULfBteIHF5lm+GClXPp8j9AXttvylGiuvy6tNFPj4Jw48jn4oSf6jR4/Ly
FMqsQso/ac0zJnj1Vu293sswMcTKbqlOIIBqX9zv2HtkCVNB3MeZucqKPSmnuweSlsaBfV98mtAh
kEw/tO6Hkslj2cg2Vf8pud7RZDPL/4aCsIFMPHEeF+yKk9LbsE/GZMunKwdm8RN8B7uIUXoyBtK/
uiX5bMjqRrrgMc5lbg1G4sFKiyWH8sZeoAwBUDt+mk9mxbFL38X9SvPT0byjW/q1JUniVBpXXW8G
B8F8duk+JK+/PZEVbXOOMqwCAS/FYpczAfQuUBN9TQ4IMB5oAoIVhGMb6KblrHdnEJRZaLSXCcZE
VOyrRGgk5AVhNEtgMzkDKmUcOwtFfBa2+2iDoAgvepnI/leLCMwq6OpgNmTLPOPUku4rL20l6/RK
0Vw9hHelOo//aQybbtdcnSQavYfFNBz05BlelXiRpBBV5oBGBdBP0vTwgSlUqmPH2XMH8i9s+eL9
CF8Z+Nqa20yS+FGarvEeu+3u6vkYpyGDR+3ooV69mPLovlfdn1AE4B0pMQUFREZoue32qUJHsI5E
4d3Pc370G1ovbbQ6CxSzpHy05BSjPqMDVL7kO+Iuym7LvdfU9q3vysnuS4PTzMVmuRsVQKXIAxUe
b08YCOd1Urin4eZXjyhKtuq8CFVWbchMKCKEKLWRyb8jff52xrQrcGjuNHyb/rWiuQKFcD+H6VjR
9qUsoucJ+JmslJV8930eoCwU7CR0nbYA+yWMy5+6Jl55R3KwjpbVjJXw5SC0t55ydyKblX7NLqA7
LHt15/mIfNQeXB2KB+2Rq4KVTez2DJvYqYXuyXXMi0+xyG4qQZqdr1DJcH0Rfh8cm+cKxVW1J5pB
r9kR/ds8mIovdu10PpLHAPXStCDOwPTVAkT6PrwWMcORRCAoUh/cuy1ScA6LcygW8fwKMaou/lOp
FkbHMYWUz5qy+JB6Le9lBsREFkBzcmnzAyeWjQkXDnBNAL1MiCk568jA3XGK+3VvucJnT6+97uXG
c8/IfIXKioXKKL4kmXrEAuABFgonAhkz/JNn0bLzZjZPfz8kScWCwXtwPeRAN41RYKKtSp0gjIfZ
eZDcFuTHOjH7z4p+VqI6oK+PWC06tjzL/mL8UfvOJKYf++mntehRqgJWfmHvshG/fr1LLtUpXLZ7
YC1xqXecgeVAzTeMJ3pyQWSoFz4LoOXPa9iZ/JBQrj0dct1uswnCfiuQlAxdR6T4hRoNqairszlH
OULHI5CLa8pxRlShxtZzyo5OrOrv4Le4D4Qu6xErq28xVEXR6fe/0odsSD9Aa0fc2YyM8q4UJ2N8
MA/j734N1ZW6BfeR6zyDqM4JUVKByHd3+UYmLAk0tyebuzPuQt94yTavay8sAtUmsyNfXv11NNWx
YD4Vr0x9H4RyldfAaCMLp69AFLCbxCvJhA7r+lGgzjhaothhqiAHM4NI45+l/cHaF9L7+a+r/ewA
eIxTP6mxD5e1mu6hXPIqYUC7+5k83VAr6PbNli+ubqj1m8Mc3TJCCW87xEIVo2dvpAvHI3xhzmDz
i8ZSd5v2Ue8XelT7hGiG/U+1n/2mPUyvi9RmtRpWeu1y0YqLpbLvUQI0EBNnDtFbJZFMnCrF62FH
WMMtSCsg/H4F4rLmfRFd2vXjYfCE7pcBTCbH6KTXw5MsgTfymy2Tan9NNyuUI6beUcLGFid3jKJL
hp/q93pbsIO9qte7J3XtzvxtJM2x1LlZ3h6LvGceJYjXglqMCsUQNViG8V670h0a1WI6PXYJnRvN
oE9t9Y+cU1k6+Z/TP7k2pHYL425Uv3QusVKFy21lGSk3HFoUVmnehCn7T0nBvGJJzp+RZN4Xgsns
yEodlrFAiGrYwW2J3EM1f1m5eV1vqfPZypO/yfpfx3bmwN22ezn4VhcX4jUn+UjU7A8thyoa3NXv
MWbl6Ekkq3ksitWXSr/WEpG84GvW5lTgNMISKBYmUokAkOKu7BENPXXAHFloGAJBGEhRendROJoQ
+J3atB0QQY1o8ex83npf5W7lQEmQ3cvR3pggk094j5W+Pq6JqAYcUuM72fhEQYVHcDiAjv+QtlsR
p/PLbYddyHHMNaaD/iplptaJwqaDUv6gsuE9pmigIQQXkgQV4kEB1e88A9TPtexKPbEZunnD56L+
pqiF2ZNIEo+Nuh8Voxx6FgutotNic/qu6tnk3VxKgF4vTU8KwMcU0fKqbTJx2eaWTADcMjX7g1h3
ndQmo2wSMZ3VVwQofqwFY/hWzttCUxKEh10x02NE+ObRX03THUzRrNO0g9Sgq2ciT8KAAPm5g4hR
FJhiRUUzQB9UEBxXFJtP/TEUrMvako8kXcJLBciCuGnnlsfCdfnpWUrN3vLvNCKZ95cHG4r5k7T7
vjk0xHLUuYCRNZY1YRc1wH42sGNgKyYGxeAiWF08YHAxNNkYXSI3ODE2IR+IbZrz24qBGBDKNZuS
muv6r+9KoIagQqu/GBXS4DpMa1BAl7qaeBwrt7LaIVXuZU/drw3ZSifhw5gjF5pIqJQoa6UT/axW
I813vbEQlfr9BMvwgU4miU+DpewYaEHdVZN4JNEJhcZCaQEHg1Nv91QV1j5VVyQR3wKLkHYn2u1r
0+xnFBeNQ8FIxRy9iVqTjpHrOPliYLVtS++4NGwdYZISY7VzTdr/YPr5LKlk87QlU7mmP17flWgf
zT1INGhAIwk217So1zMyCSiqS8Ylte31txhyiSPRt0BPT8Boc2OWQJHmbUEqsP3d69wM9qjyo2KX
6BrPGKmqvDk4g9zst/Y7YMGbZHLhUsYTvhcrM8lgDxoNJXlNF1RHXnD+cklHbDGGqkmfYKvbg+qY
0k6PN3cLyzMWNUg0CRL1Ep5GKc0caQbO/sEQB2WcAogw8iP6BFEAdThXV5Z5TNt6ZWTJvEs1pTr7
d2FiiA31ri5Fj19q7jtruGvDu7YqSHesItEa722zg4k/nCAsT3/QZwsVt3+sH7juPMaepz7hrxa4
2u1mHen9Z5DW9LS3Z/2bsZn9TFezMuC0U+ZXvdo4YC7YFG7v8PTW9SvPVoHEvulfLKx8g31VUJyS
bMiw4GyXY9zzcztVd74H6Ox2lny3CRk+tyu3nQQonzl5q67tgcA+Vf87fQ39BN4o5oMDEnc0zZPs
0agKB0e69snQ76F0gXjWtR63gPDeqSU8Nvc3YbKCAI72rZecTI+PzL4KDp4RihHHWcznpJcohTI0
gDWB6YcvKJQJUmVQiz/+fYXH8YhPv1ZkgWyrAb5aeOP7CHuAdv0Zc7+W+ZpPbNKhCT8n4IGcnGYa
TGZPvZGpKG69HQ3rrDUHm37BhV4FnH/Q1Q9LAtm3wdyol/zrvvTZF+3HyR8z32nh/c8efXV2kqhv
TwpjOS3lfTJMYAwMZvciwHXVBqxxpO2wpPg7fMetro95VHmrFQU9oCenCFjkML9JPvZ7cnbCfoMa
rDYAhyjGFLN3Wr1L3oWIasTe49hTEKiL0QEd/9MGSv0/JRvVjbMgVQbr3jyFNHoHo7TYJSupALma
4FeufB5sQNBetqIAk/9OBXWgycOcx2mMSOz+CcriV8m/fq0HrhwcvMGYEB3L944+9J1+0+Bnw3Tj
tFrS97B+/L9GtE/g8NRS+WURLzCPmsJcIou5j4ZhMpRrJSGbQjhypOdQv39LEqW2lYK3sMykuTBd
9eQRLRSHKlh1LhrHVqVYOKM28V7iBl3bXmqGvfTlhMfFyybBIAjUmrPefKhUpQmeFiSDGtVDk3uv
+RhxnN2InUE02KwItyHxi8TjmLAU4KEAIY3d5PG4LZD5ntQgaDPPa+Duz4EFtPPXt1ek8hpBRpR7
lORmNsAVVa0oTPEAo40RO+rJsWi239lTT15DkZTw3tzypjQpRSLoffcyP4qxuXlWgDcaukXrLyK7
aoAUwNplbqtoDKq7YT1jtRONYcZK1zQsut5hCgna3Jz4rOMIdFO0Y0tyj49h4dhfZ9h080Wq1VkP
Fy0klrpa4AO00R5hwEVzxGmP9SwMqa8dCj9xZqPunI7ndhHQ/emRs69HL5szaznx/X/9xBrIoZRv
1CHlliA/aN3yIGb6oazE4DMwfut+Mk9lLhIrgs/kGxwqUc5p33RThOLi+meWJY6gA/GyOX9UTiyb
Ngeb+LraTkwRW2CUO4CqqO8X79ccV+kJBcqv6kAAHLfo+4WqHDcq/SwsUjBbH+1mnblpAGTtRsDy
Uz06ZeM7lwoxBaT4o36HNPJLpFHgNcYY6vI/p86DtDP4Ui1PwRWgjlpY5wJNDl0HS1wa+1MVyILj
T9xGtbvHd37Mnsbglzq+EudnUrnK4HnPXLGWr8ln3Src8HCB96ZTPG7paCcri1YLu1hB/ZpsG+M+
ei8XjI7VhFNhyU/VgGLP8TZrYrV+MyiJIvL2zHnkD/OGmfT2sKV+QE/xs2VdyqlEHP3xhoDGlzbo
VuZUKlxSNc77GDZmh9/3BUuXY33/nzChpVx9AiGD9QLWwnK7kR8PAmgjkZJLLeurpKPLTWYfUa9u
6+z515dwwjcQeVdoID5hCtL3bWC2aGGV/zCLj6mkuMf+9h2xmxfeKNJJzPy9b2vEjlsemYylux34
0zRWS5cbwa3g52XdXPeD7B29PORx3zyBVgN0ccoOCbiI2YfFEqonVeKxwu2NWhjW1TB3IfrDuOUj
wACOSSMlqGos0SNeTLJnBeBhCdbLmPFAR0zFWVyrmeJ/ptp1sr8LDMhoMG24VLEaMSbS1AerNRia
SFRy57fxXmhEOGg3dDkXQwN5Yx4mOywezqc5lTYUsDKLMwWyDGLktXtTc1EqJEzazC6hO4ijKPRU
AKIzVsuITHtEkWVOtJFjzkYKundccNbVYmT0/WJpiRQA7bGLLQBgwkxH8jiAe1CR44YYlmBD+Cba
i8VjJ6JHAV/onOY/PAOd8WhDvai9SOWC1sQBkqkrtUqHl12Ep8NotRKGt6ObHjtBOQ6aQbc7zKnr
UP62bYNsQHRxcoCq5a6fUfu8CyRtcOj6d8qJBVtRsES/+JdV7DHuikC6Jv/SJ8Ghnw7sShHrRNsR
6GrGFdlpgnpXCnxw4BrCWYcLMFlz/MPJD9jSkyvy4UTJvfGLOkfd8kT3/E7Vcaeuqopov7qBP79d
3+45DafW5PWwbTTe88Ke1PqR8vkW+JOB//bRozAnqpFz/sK4/YGPAl80ArYRowFyuKHt9JygJx0Y
zhb+gPXaD7sNlwng7DkkhKAiVy8W1ftLZLgSV/nNULmKONNh5d3bFUoZyAEjpzjDI3KKK4nXyrv+
QPmfk53x+amS8XEqrq8t0WvSGPJhtDIyoIpLjkLMFzptifvl4HJdu4KH6Zx8khzZeT3DGhcXG1+5
lWrQJxkwxrTN+brh6DskJVzBRwnMb19fHRS09NDS9kz/7tkvA7iZjZoes+WKqACO97zbLUCS2tO0
hYy1zlQENSIyypc1+6xeZNNCj1zB1teBHx6DTVLx4PuknfMmbbKcY6R0/urZnIAhM/B/dD2oTcXY
0zJ/z2yL8wb/UrNG5bjXOCPbwAmoy6WTGXsw2so81iaJZIulF+IfJD9I4Cwiebb56ip15SyltflR
KozhZNoiZpUKFlUuNoEkeMu/8ekxUz6rx5lErho+RjQanNrLNk/rblxROekCZ1x5WTw59fp1SOTo
O2rFrmH9E+nJJ8oqRU12Je/KhvOS7GQhDrGvR7gWK3ERdvHksKVUGNWtF8PZP81TzIeJle4hWl8j
lU/pS6Py7OL3Jl1RZgzzfall2DGw72sgaHV660/67BKLecSDD8qPD5sYfh78K0DtA1yAhCukS9RM
nQO9El4C8ejPrHA/mRFSLVgxRKB5GLqp49u1CQcdrrzwfwsdmJvpRtW2VpIxovVR7xSxq2EoeACt
0BWqBALtA8LTaMShVRRHEq2N7tmhSt7l2Ah3a4QrAnUrE4h2W+3IKE7O6FTDj3hzi78f7A593ccT
okL4pDaMt+ojx6yaVsVYj+HYq+9O1WlBRlbIYXvNRFsQ2j7e3LHs+jcz/OF9ntEAqUJo6qulR41E
xfOPaEklzhLnffc4I9Xvi+UnjkERbePHEp2BeIHoyBI7/jGSi84IDkwkSXCURfpbaL4kUx7hL2Nt
CdSN0KP1xU/gfBoP4A5S3PdKySUrRKk4IZFrbNmUFqo8Ji8RyWmxAr+nbCe44Kcz845Qci7dTr5N
ToX9ac4k1qRm4rLmj3cGk+j4HhR0d9q9+EyYNQ4A5QsCXAkc5f4UH+LaM1F8SEgMRvvxVZn+/Ca4
IOrV7hNFGgtph9DrOu0LgFCTW3Mst3OqAn0BZnmId42b9qgVUGImd1N82xPjMfAGthlAH1fHqSCl
p2gisRBDvusACMLp4JZ9GQsaU1SwTb/Ux9mVjTayi9Orl1kAv73/B2piQWWlN21SkjEXxXym6QI7
qbNWVlE6uc+MZ3+bbSrtrwBW8XMn2IpejQmBOwDdGZHQv/UIaz0jPv+myzNFq+/9r5Wjs1LYqQcG
IeT3cA0RNi0AnG7nJUbyUwx6ec4hY9takWMNzMiADA1lwqreXggxky59JlcEf5NK0ADn0ACgpcRS
SvkncL72nBRESKoYclDLoGAz3fj433fbNsOhU0//2XweXBlWe/QnGZU4yVMcvDlkU+pz0EgVdlAB
hObI1mxiyP25vwO3U+RugSt7LlSbbdBnjyyi2gG8uRZUAoJie92uiRf7Xv9rSVTNqMjaGIyIKvTR
HZEhY7lUE0Ib573LyqUqrKbt1yPGF5q5U8P668NXa5c4P8qEOObmp/chXUtFSi5B4l1vmGDshdwn
G6376MjOUnVXjpSaY96yMHTpRcHsOu7SM04vkcVDbFrABcdguKtT2Xg7np+nlHtMR1ms6d1wR12W
Mqd+qJ8a7VERFWMvVeK5bNVmE39J72cKunMVvT4ZN9fqz7K12JG//vOw5s6XAIGoOAY3Y1Rk8iDG
a1iTEt5wauyEoO6X9rr6SRGxxadmN/2AcgMaRT9BPOCDbWvhZ972bBKIy+Tqv/2NvCsaLrRl3gmu
sp73H9FrheLtYNQ5lqx+FroPgsa5BY2cxlJeYqSgcXkda1m1ntxNIOZluSHsrGISsq4EPpIAV8ZG
H5C5rnmiSTFR6MXvaj5wMwLUSGQTA9RX1djNsKAMLekNObBtHqS5nuot+O315Xc9/RBQ84ZQdXAA
CiTCPFyNvb3pmDJwDzfoS90zg2lRIdDgnDhTgSmCo9fenOzUtX1plAnMD9TZ/Ci+soj4PriUwXj8
Ijhl2vwlQl2zhXy/hI+1vGOhAfcXk5MDFlMLjB84OTmEwdhuj4b78JzEUlQatc39cjnqFCgZrW+P
mPaGen1HgkBpIZya5nNssAI/Vu39ZmVFk6iNKZxbLkl1wszt1OZypSgLFqVnGK0gQRXS+FoZgevB
cuPCsr22Ls/6ZuY41a1CSjQUE8FSRXyefZgxOQYcZyZ+0c3X17JwJ3oW5kaeN6D6ifeSUNX54ddL
w4h3He0znVKza9kNCwic48rldva9mf5qd1gEaUVbPcaGtNxUwtpefFtib3b8nK8fi9SiURCFCn+F
l2nm29C6ZyJxF4dC1dhoJNVPLgRQfPx6IbiWgQW4l8ssfwDX4SYOtqir0uQ22T0usWv8cyH8s8cc
tfhhv6Ekdxoy5QBMFJ80T3qUFM758pNOhR4HVFWj8QPls50aKuJY3huT/aYmgUnZ3zoFkNLC3fXb
OMglQRpU4RQkq0KQSfA4BRoMg4RBaa9Rx17xz4Xb7wgC5sxILES1A1ILyDeO7XoS8JoUJ2Xlprm9
e5fwogyEAJFwcGhQXcz65oMnBmQimvD4MyUjFIGZ0hOZ2nQO0aCVMhuAfBh7Ro/5pTLvQDpclaSD
QzcNSkjU/dT+8VGHilJYcnHcSfhVpq/uNGraorIJk3yZ5r2F4RinFy/Y0CB3m61Bb2S1eQQx/eUS
kpqTzgaq49K0wtpcchF67MqjGAuUhYKfu1bE6WXa33XtIzqSDMnxXZ5CGkz/x32SKsC3G9hn6GFn
gu6CuBUoQcSe5mUqiY4E4nyTjFhtIJzfJ8m3pqJ5Pif1+3dOaaRIbOyn9Zw++3R7qyVBzlt4p0m5
s4lgQW5kBnCtQi/4Gh6sv/7MnmrWTnTm664fp/bmyCjp39CPyjW45xpaz/z3B0kNl36v+74+2Jbw
e1LusQAXI87xq9/+24LO+beojilGHX+QhEjenRuW9YWywhOcG+KEDskG0V/6hmAahpTpCJkIGIh2
5BrnDPBrWrp6DH5MzGDE9E2rTGWz7mv6D9bysFB0/RC3HjIACnMkxvP7jNOK4RQb8cqV1b3gJzlS
drjyxDHlb9v679LSXEmUivm3WXsC9dhxSviUkFQy/IloUlrxIUVn+97u+T8lmm/Xx8ZPzjQtAcIF
uXyr2mRFxt0gHJ2gtDlq9e+/QJPJTNycVcbcleJPCZoL8wv4O/36PCBtPc5hic6KzFwrK6lzX7A2
YlbmqGPst36LcKzs5sF8G2Yr3tc0QjJBAcOS0VN+kUMHo7MDQzjlRd0Nn5mpUi+ycwW+ko14jgNi
okaoipbt0mBLJGKlrZVKY0Dgsa3LChEkNVAfBWEoYIsTyPvruyB2SfKtLEtF6IMARBx7iFxGFRfu
epCjOYmZ6EKFJNiQ3QH0xywmW1A2damp02RvZOx/lZdOk2m1oEqw8hET+VNBrZdbxsNws000q+Si
CakimWf6YY39jc3fuihxPwlfVr9nk/77ZyzWwHgCnoXd1a1IlLH3hZdGG+ptm0Yfrur467NcAqXW
AIZnpUL/pv98soDK39U0CkgK+JMil8DAUSxUepIyJctNDWcsx09Usu0Jp2BepHQs5QihAq7uHVfp
YWWtm9CDBc3kF3cgKy5clT0S9wE3o1F3szrK6m2k/7WQNXdVLjbXE56I9j7NQ8MwcOnhD9/TAkXS
0XyyxF5bZ6InSFd49HRo+34uSCHqnx+P0aGUdWgBZXhy09wXJkYCkqP4ZiOjPUEm9eksXy/cFXRa
fPJhj0InEyroRdQnlE4ITVQr5H3oEASIUwgZkZyiZK3yhhgXepuSJ8swA8NWeqA6DyWSaRQAkiNg
11HfNGO2j0AyhTcAqpclmA7GshVtpI0pCZ5c2rJRGEz0/PgkprKGj7ieDoeTVI0fma32pRjmmVaz
6rBphzGFbEnsrpeePPhxiaCQ1hp9zNzr3avSZP8gMPJY7TrQc80qOCRmn2raMZXa0gu/WDqGB84/
gjv8aay5DFqtG1I3WNYa4JZczMVih58THxuf+UpLiqjX6Cv/TODyuECVwuD96GAFg9s+vVQxaLFs
kvZnOLhGO0r9k0FxQ15jEuD1tx2ilZX1FnUT+TOBjsIKQI97Ue8eS+XtIr9ZccgTC5fVzCKlyoUx
zZi6MxW9Biu7gTBsp/3t4Jw/mYOCTarxoLCWo6tbOA7VCIJBm8T6s5+ejVLtjoDGL/5QICPPDKM9
v7JFEIe6DBigMTBPenkRCCwflv2aUtAd3UvfsFJkBVzkdN4rFKBgfV8OCjjOvhCruFPZZJvsaRZv
B/IAzvxUK/1tyuNFG0RGbK72oadKh88IwDyJ8ZuCV37YvzS9+Ym2rg6zvG4u5LauL0Ia8dOtLkX1
33T6msHx9k5p9IZrMxybIjj4N4OcFR+Z5N8b46wrHu8SezMSTBuDbE1WYVZGMfvavLTfaXzJqMvk
Qbr3kYWLqzRQ+e90jpMFjb6Le+ObExEhi/APSUKm6XsmpnLr7v+F6QaxBQ9yxg6cJtwx0dVmsNX5
awGQ6Vphe65zpByyeYbLAcNHofWXPen+/bl06C7F1g6YFZeWrTnwpFujIgZqUyKO0U9Pc52JHchI
jMPMaaYg49bbd6GaxPQoV6aZ33SuNSMxSb2f6k9tann4xBSv9TXlvZOILx31lNOEyGkIlN6fYrIw
O+IsPqmJAOhVypAD3m2LJl9GneXIgbXOdQzFxsbxJQXOVES/kfRTxMQy3lyE0uEvUnqB5JRbjZTF
+N8nv9NO+Ta3lYJUXi2kze9g9fH92pYisF3cOiJ0NoMxK3BfmDlDMIaYCEpu0iGY9mbtrFA7fwpm
+8809+fOcr9nksg/lLsStxjXx9U8YJjeHKhGMLvp9zeKm/glpGrVKBBdoQWdxqwz0YYgKsDWyaxD
xRRPH6ivnQT/ycER/rABbzh0lisS8DWKtRgHYrgrcyr2KJ4fqF0nJdeN3BZxvpo2k+5xdGBaf+WG
HV/jw0DPeMGZxevMLy5GevvKmN9XDHIVadZ9Qy/KYIq0masH9gGYQ98mWPrGpHMcEf+it8kFvHrE
K+EF1u6D8HhKv0ZZeejExjzsLybuLrSVuc0jF2MNYNWIuJrwwqCxwoFaqxrlF8dBriDoFbTjxdOA
KKa+mFhge34jyIizNjEUfsIlss1ohOFyrMiUy+FC2lEB4/gyF4iEgqZIC/868wMAH6pxSYSfgqli
/XfqDKUWzxsc6mhscmMrdN5fz524HKuzWjw1WfG0722fYrj2jBn2pHfCOxHkpOlXOGZsTVfU6eWI
WSvS/AdfHLMairN5LdmPVIERP1qaGgvjrvJvsBYLwHi9EqCgVmDLCLpZIV4Hqh4ivLbFJ8/Caru/
m9fAt5gtJSasLkQKZfKf92L65scVMw4+po07jtaE7lWfH3seccLuu/o3ECF9HIf+LPy1gJ0h8yYd
mXblYmRfo7fdFHxcEZ1x3cuKP89W3GHC8hZvJboTejJH6VYlqRNOlbo5xBYS+L/qhgiAzS8YH/Rs
m77HFuocb+SpkvrqAgJ9VbUgdSO4fPR+FVFQsZiQfTaO8i6919WgrxGfFz5Y5OpznrzwFnKiB3GN
pXGdn1YNaf68Gt9sp3cCSEWy1iENUaoKyALJrtOR/Xrqgf2qDrPsz7dGseSwbKKiTkon+wEMM/JY
FzS29xqm0Zpizm0wkSAfQ5UltHAMW7UpBz8SfgdwoWYSmepOPSPwoVw0UUunkPfF5xiXy3urJr0L
vEubQTueKDk3FLox21lI8EEskh4apnkr3LEasYlTXn7Zu/Sz2UwP2dIt87l2ynPlDaBBSfizZ8dc
MWEgG2EsQN9c5pBCPwsJJVIMaQWpHO1gekVyYcS+Rs0CoevPDCopGhbih9yo0rVeIqVi200wjdiV
094kLte0VuZ0Fq0xRdjWTsisobrnGvrIq2eyx+rkYv54i/KxzXqqaQHUAP/d65XXjbaKqWeBoxrR
rOa3loqe08nxJT4y2LnPl6phE3vGl5bEKUDvzAaruQqOuUu3341QwJZwBe9IC7R4ZVocU2d7A1mE
5dFx+RyM6arDMKYKlHT5UyIkmcX03AXpyM2/EXwF8b2GxBh/5RAZbpEHH/QdfxqPH0yyYtfpuIZ2
MaWbLq0OQWK2Yohd1E5UXBsWn7wfdQM4MO4bb/PziOcv2mfvInf/abc2m7QO+5rrTxWFkbq0W1Am
2/OIU1tmEsh8ZWs/jXm71RAJZWSY8zZMRGbjnXYL2eXQB/p/WZOWx6YTMmsBGUQumoWHIX/uFWNj
CgJHCgB8l0LIimi0qbYXv2GAk04lh1uxIuyNXkCo9nHkhtxIJZ3hWNeh1yr7BAjBLtuqGShWl2vy
VaVc4pvN/fK1Q5pgSU76zeOyVd/y5wKQ/8/6OZlaJtnjaPsP1SS5s9RuSAU9K83c6o7byFxaBCGE
x8vlk+LSnDHJL6ZO/+md92xQfN6GxmQCw2a1Q2H4JNixZlY/ZGy9YbLp2j1pfh13gaLV6/sF1/zy
UE+7ptfVY+Hhd9D6IkJ0BcuhHVWGXd3Gx2zsJyKdV1EDttfLlLe0RHkhgXn/BmIa06X55D5fnbpN
XztsIcn7ZAj7SwxgctAahwu0XlukhXClk0eNSi1AXwAmBjdX29uupcImIsAufb9KvIUUiRnm76OZ
R4QU/7+RrYZ3sKciEJh+OfM24fwXjmx+GVTu2uEozKVhJg0il49FNkv6Fn7OZC9RMRJquUHK6bC7
oAZ0yskCjIW7Pk2apeL75c9z7huoqaMG3Dnpn538Fz90LQGnkVI9BoePWdgUvp9lb0dQwV/1nbp9
Mf7GNuDYW1Mp8L02gh8bH3+8cxA4qUIoZ8/eizPE0NAv+iPm8yqL7FMGjJVoeTkgIqzo+bKuQ49P
VKxRicM1aIcKUhjoVZoBhmUNwDu6cy36HZ0pHPhoBgMvO8p6aO6QeVlR6hVV/378Ro4su4fnFxVd
PFtjRTTrlLHt9IrHjspIw6CQGqJpPQCWfiidhGNvaTkWz1Q1PBwZPxjrbV7JMIdVBWrwixdTAUtd
NbHib+r3KhimgCUljCFbe+5oVQ6lgA0gn5MdicS74E7EuDpKaW800bMinMK2vmh6YFg9fqRKcP9M
+XOBvBmR+PWsETZt13zUknwDzSqSCM7thRRhU2UC5kmxDe3FR9bonSy8fJwzaQlc5wlONJqA45Y1
qAZwBLFf4rg6k6bVdK+5Xs45ytrLrqzzMBpJar/9JFkPJq2wLaCYWKRnfVxCHrpKMzi0i9WjTiCO
YSvfp2vADBiUj3gma7hDAGrTp88W6CXMi4r6Tej25Mt8SsQtkUXiUhm60b7+22JbkezfcvHIb8d7
FJHWW50Y/8VrL1Bzp8qMWIAHxED2AA1ysWhdPVmZ4fsg6ibBthPePfl2/W6Ddqdm8/8pavDJkNZI
lLVuQ5ZkNmep+BpupvKL04OYh8qtEKN5kpa77jzNobgnLEvAjt1QMk2JLc7A/xt47IWltaTSPM+8
oqnjKFreou/QjgTcWeeV+9/371LlxFjjHGpgmqlDczK7O70HlOa0oh1ZJBNenpolUaf1bAbV5SZ4
aQQaA5BxcHFNoPNVBEQFHzPYcs3PpovLyNnUaxxDoPLxRnSDBplqhSj93XrK64doCpvx/YMeNtGr
JLXj5zvN6UNR3OwzgF8w83UoYaeSmYSBUpRnZsSbA7ViA83ZLSnDtLtL2gLJH/gITTUvT0UFGC2g
LrVqPhT5Tdgzec3xuCNoUlhLKQo3Xe+R4mihFgYolcO/sGvC2vILszUBUYgef1xe/e2T2w91kCKJ
3gtwyTuMZNexT8+l45kSbkrmgUAn6grVUu2qsAcv/wj672p3xId2hO913f2wHpPpPNw/vhqbwney
rfTe4GGpK+MI0vM6liF7kVoxivh6xsTjSaT2P54BcVBaPQLIEwF296RvK+lqXWHAEa8t2CbUZIlB
TvSoStg2+w0BZuuYIt3cubAu4eiLGxh4N79Pisv3cmupwVHFfzeGPCD5duZ9KRpS1+QJxmkd21yO
gcgFMoeCfV2+xC4+5Nq9OFmDw3/O/pUDwjPFVbi1Ki/VyZ2SoLPGRUl2SMeinvkYAKna2cKfZ0ai
q7CiWpRMQS4p9Z6hq1lMTzLrxBf2Wn3cRMvqMALTL3FVxtIjILJtOVebHL1+kn25F6IBDQ5rd8wT
2jdAKfKcAtDetJ5tNlTi/UMn3w2lQ2pYsB0oO1AUs55DZ6YJeNyxV4HqoWXDCdHiRfrd2AR3flMU
P0V+JMOPTm/zTutIQdSHsGWnN5/IfhIUimakzWaD9hhCzFGI9kZ5hMORw0LVDVVDT5wx4LWwrZaC
EBMHbYQVLvdHQJINsZDDQZ76WglqPbUZhVrSWXAr0wkRyu/66s266/pJzkQgV7mcSVKXcNI+wzZN
DvT142XinzXe1pbkHu5lnmdWtFgqp4u/YWggUijmEsoQZvLEMh7ncmD1p4JaBCL7olInEhu9DAfI
PdVmLAjTnn30C62mSI7DQOVVfq8EiitxQ1tWZiNomOicVOsYB/afcEwdvMM/J40GfyigtXqHcqyf
Sf/G5bCt5pYL6Hki6KpQQT0LW1acx5IA62BScKr+kktIbnfu1b4CLCF4GafAG5hIjQErTIPE20j6
Ar/PMU95z34x/wsoF7Li+xNjiDF3+txe+vvDaj1FdrI2BZkg8QUCuOdd/9Br9uU4N3qViUIHIciE
5P+tWcUwoVFAsDUpxT0Kg6/+jErrctu2JZ6+Mc8PHtMvOyJfCrthasuN94lFFPXuK1iE1gPQtX2e
Ce9PlHq29yaXUU/YqEi9i5SchYTLX/r1osmavRRbtMWYI0GYLHHGGPrUxXFv+NAvla5/G0zmw/Au
yhYE7pKTJ8TYWXmQuTcxxnV2llC9jW0hx9/WgJyvvW9vcFQWjQH9ma6BuCiW1iEoTctuNrFrx/2p
iMbajruJcuZ5sziLfMPhvYwoXbwTVBW2Vxektn054cluFUK7KHv9L+FFJY8cEAax76Er5W7n2Sy9
9nRgmVELlHjHfM9qtx2rd+kGjM0qZcUCl1mTq6oYTK96ZvzJzsjGoL6wpLdgYZkAoQyppMliBSg2
4VI6ay1Ugy9PhYjKEdysZl1glxdb3wJrBt18OMOX31w4DvfXMx7vlw/2C2v3SRwmzueVNIZviTwG
ORmOI/HpmKkc+//louRRdOYbruo5lfSQbFdE14uDWSmFeBAh3zklSzYjyhR9pFtxVX8H+/Fpq45S
f4CIu96rxo+pVznzZBSoI7O+NBL0+ZMt6KHVut/h2eK5WnZX0c7xz1sTUm/t8UO64t6Ql4EyBsS4
Wuko8udehjeuUYBUKVVv9b8JHejsmAykYtAd8+Htzu5RlkoJShq+6NY6X+WQuXAOdGooS5AAOUJc
gxI4dMhimuxOZ+CDu/offxdhkZl+bFyCXp63S3FyaxNqkP2pbE2l0rHaP0AYtTz6eHxHjRr5W/y6
xzsafbdY+CeMA+CLw2cdNX3shAn/TbWfapBKdOcpebV7dbWBWhXs4h76UfQGcFTY/K9U5+OCaUjP
Qgjdx920q3L/DxCk+6xf3LNre2pvphZvnSlcarj9mpra/EAQMsJuelCW4NeJNwv7RQrwnM1+zHei
0QIEXtydvHpPCaoV/x24todh7tgVfttKwJtZuCE/4EVZ8I3YPGRtKqhC+talAHSots9Lwax0v6Eh
h/Yl64FBfRZSuDSN5E4TGo1NrSDpOs3Zf61blpNa6mnZeLqS+0KGv+/VA+9VA/YlBY/ZD3MND/uB
GwEVPH+frR706ovLjSGDDQDSg0PMzsrzLsyWu0TmMrOrTZGjKOeXOB3m4O2Qp+E+WXgKi2uF9J1y
i6M4blPlkkWDVwxPwavzCW4yDa3z7lr21R2H6X+YU25Pwpa8SBibMIdiGs911/E55SjTZl3OERMl
p6jYEjplI28+nCVbfu38KSaLAk6GvsgaXSbZd3nirLeoDSc985mmFskQ+TIHBSMZx0XqLyslpu9k
/gCYDm2Mb+Uu9kbM7N+1FLAqc/BgdD8BrfbCr5rYzNRZYq7jGEVYfsQ7eNEDUVcIixn/k4krFJLx
tv4hvSWhLkmEhqv9i0y8/N/3R2HFOLodgzunCM93KNzKe96gsXDFMvYJObrbuyE08fFEXvzTC2m/
+JpaJSVlIbd3vX/Wa8eZrhRqN03JOFIWBoYfMCrf5gB9ZHpBDGq3zX3wJnm7lDJ6tAjOmD3WHN7a
aBqCaqWM79d893olCZyHMQphtQBfXrOxIq3lXzr7WqnexD07wTwg7j7RCoRyKfd03YXY0HDchJmS
PDQMbKySKpK/8pkJuFC0YvUxp5mWupqEifgqgEeUNKXiA1HRR8VK3qmXagHLbK7m+Ojs0I8QE54q
+0QUAVyhCf7/I8lA1dIb+iAKGT5C3amOjplmpNDtgFCn29LdO2AY3m45o5Pqb7tEfRHFjPTvPuW/
AiTOb4BrPZ/fNFR7/nfvnpIWaEnPE8VqH3zr8ZEvP8m5SuFrTpaTHVUIjfsLR/oRFDY64qHwvQAb
S0O4zd+cNQQM+eAj8F4+FUIoBXAI1C0wtklPiEz0Ml3xcZWGoYlbkdOwFC2/6GF8GdL7JPE0HmKP
332+Gaw8QcJiYxBx9EdpD7lLIKC7ZqKP1EEPMMiHEAAzYtSLzEGRwcNmgHrB0FJX7kwgqPVaNgiv
ba8nuYeT4jcXEWW5FW2Z3naFMy2Ajz0/dY9FNWax0WSccKKmBLcB8N+xuZK3WG5mxItN+vbZpNw7
bjRPBtrCJ02d0VHKG+3Y9Nafy1AOJfUoSdrbkty6qMPjNILPUSRbcEs6P7Vs7X9DOznHsN+z4cTL
8vQwnJ/oStw83OGoXHQp/jdaFM5PYyGMdeP6FoFojAZ0xl5DyD0DRhULF/cNcv+H/QnEEoLR6nRu
Ogezxrq3PBshSpu+f+JebXvCnNTXmz9EozD3T/9Bc8/4zR+7hlYQMooGynyupizxNVmPbpVD0v0U
8/DroPbFsTNiB2PmTBWOyM9NzXJmamxI/u4CelsJxLdDqMIXx9AwPmGJ2s4uVEKsvacPNlezyAL0
j43EJC13SLmpY1yCAsdJhcTubjSYoDZOoUpmrPMFF15sIIluAcjqiTMVDkpL2KlD63fvtvhZi7yc
/gB5M0vD3tF/cumZsYoE/eoPEaVQ3FeO/CYGQDgVzwX+MBFIDHVY8AcwP8w+TPE/FMQI8ebldY7L
npAdhZWb+910uuBi7S0a6Pj9zu4cIdW0fdLymBHHtDKGjLVUVE1DHH8Uq3ncYpBbw7jOkwvTH/nl
En7bz8Ja6npn4QtPh7m3hIX/gbmnUSLdejLKKu00eSHTKaxXqcLTWTLVIPZhSlzuBuDx2f9Yo1kz
sLR2Sd/PQb1V56tKi4pi26GrPBa7GUaTsQDQoPjtuWnktQC/Uge0NNSACJ5QI4sU8dEmD+gAqO5w
Evs9b2aR0HOkoeLcQo6QjKw0/B3tqW8VPpHZpkix5E7sqOj3ZYXy0GZrjThLoXc6Izns0EfU2fNb
vNXYWGXuhMZEVu2O1vxV7jGwmQ7OCl7TV8HPhP3QF4jvELCMVbmQz4efyw9CtKi7xxaUBjjEX9H5
7sRtjGcoE4C+c+AEwaP3xX2Uggjv4zNGe/C9q7F64+aXs7sh+VN0vfD3LY3pjyrJ0Z1nt53Bhsv9
3PwrzZXlQ4dw9fKE95CSc83yUp9ztBSQyjCg8Mstsj0CR2ZN4gCrzDrkbwE9yfjs0RRKDxVY/fkt
WZ0fGrXs2MHfcgZpqvsG8KvFWk53LyqQt4qzWNxvx+CWtVwWuY2dzdBsNL+0bxZBRGayX1aEWc7s
Q9Ge77tyKeBQSCPOZ4ms4NfZz4KMwmpgjPldd6dewun1P+NtR797QycXySPGnck9GxT2mv7WEQR2
vMk/+xV359RLaHunB7z/CdZWnehB7LEeYZVmITLUFHrsi49ZKgonErRe30aDaStNzJgywiNlMWYF
OuhR9xVs1hGkEmGQZk9gaLRP7Kr/N0A6Z0oYHS7BtwjrCYKX9j632KxUqRoh/YFNHVurOHgFy5jm
cfYmcgtXU0c6MYxwtHDl+pJjY0KSnT3YTymA7qquJQBRLgl3nCbnFBkyNVi7T12fdLAqNluOvNXs
49haBiiNU8nXrj4d6d7o4S0blY/fl/aDtfZ7JZLVlH5lm99jhSNItMdPcJ6T82RDEnojgfnjKW/z
R7JgaTHWGw/XgDwx0FVkJWW519b0w8qUzTQfchY1YkWODx0eK0HkQrPTX8g9ZePU5WtNYeOv2u3J
qT80c9E15kWm1VIwpY9CQ+uZXPk5ElILiRMxQwtf2ES3WjAo//b8cnn7YuWZ8UXBx9lnMGt/p/0x
x2zrllEuTXeJtF6RpHN0oUXLY8sUY26RXWIPigOBb+uW61B3p/FWhEth8vrs70sl+KOfPWoZaqyk
1tZmnefE+UyOgDAC5IBiog2heqfyk63G4qtlgT5k8sQZVtcQSTovkB7zQHnLKrKUQ03Jw+TxqzVT
0KH0wYy1011mYra69uletfgjW/4GYIvf+0dmfP9tCZUmQHjfr3J+vDuCNHSpu2+1D0ZCUBfDfTxe
nqODFr9ocCrMDAzONZ4kSbjc8o7cVobo20xEj0Oh5Y/gdMa58CmZT2/S0RukyAf2BTE/uo+UNK+h
/jKcUP2z81N3YjM1eOHv2dhWCGTdoXiHWcwj0hpQRVywuNASrhwtz0YePb3nXClK8IpvwQPcu/ve
Z81YqLuTS0YVTVfEy1CZV0wPTiSmQ8o7UpnKTQkszk2wZV7fEvD+aGuvZ3GBwoWBCXG+ugBddhBh
LIgE7cL/qKWY7FCkE3snHOTvm6SBNloC8/eenq0Vmv/DSKV3GI/XA65paKT7DTiPMZ2dYqNrWqA5
lLN2IYaqQRXMvY1SeHAQb18Ch880DhyqTaYU/W9lR+cc/u7SgbVVYpwL/FifAoes74f7G9Wge7/c
YlKTEXCQJ4v4M+D72+75vIUb1G/AlQztDsY+MDWughFzgeqLY3kjqNxufNvmMm0BkLBnrfSAypkV
GkcKDYNAgNbPIYEgASFHMgs/JGbjOaObVUECG+3+giyPW73u8Dv0ks0tDosoDZqRFPQ+5+USbqs0
qsQYDtVqWn8o1KofNnz1sKliLev43dBn+O44F1v/9W3aSmmJbjb1E6NYC+n7A6Dy+f1aSP0XFwF+
SNdg/MpqUP4Xdkda3MQbdyuauXCPgOcAO439oZBB4NbnlBoTOFQ86To1I+3MYUkCI+t3fYsXRX/2
hw72IfKg4HSEZ9pfTzHfve7scUDsQRE9Jnx1zeHyqLpHd5dcREYlAEOaZ6qM+kk22+vlB0T5d+b6
Cu5W3Gy3akK481XsP6AqZK1fa9avVJPsWq8mrikJ5hR5xexgd8iqrgxq9uDzV4svleTGMuuAjfMf
EaVbEAT290z0sYGIi+zRSTmVgwiL7elJshbAUZW7FSUyn+fqPkLgtmxqTXiagADOs4+PKRYMFqIt
iz3/urUIes3XbC75kT2OplKJGCwhSYn0VwizS9Cg0IzPhQqnDxn3h9R0bbrKY7j7VGkn0BexcraW
w4F99TYw0689JOkTr/E8RRMbwa3V6XhoLlkfvN97J3bi3G4cTNLLEt8OPDEREE/NALI0JrT3V2sn
Z1c5RQbRWPFUhR4+HkhNkhAwW3lHKgTtnAgpr/Ep+8UPu2dUe2ihU2Alw5bXPc4wANYD02DAN7Pd
IPJ5aWCRlnlhCncBNi0iPOrXIZPyMF6uempSvkqrOTF6SDgYCyLmGR+khLfg/IwYwjj7Jaa9Fen5
5nmlbxbuzWE0nfUEQTxfMMPPU62n5pPwKb0Cn3A/boHLLDsvmwLWzOxkfqr5PaTDj8E4RzYYmxwd
7YdUBQs5nBHl4T2yj1Kjrv2fnllmX24e0e0VJEyXzmz7TaO2EgKLEXWk+eHxSsec4Aay+A252pMO
V/8zRF9x5aY5LTKVWrzIP5vmgAObfatbH3SMq36eRQ5trRFU0lkNXbaXtSZ/ey2tXzrC+bNgUNad
UMNQEGOtQr1qbyhLxJiJ+fLaR0s9hT6ISZNV+ENtzAQqfEEtP5raJ0bvl7rjTSdw2XF9OafPpKa1
i+L3nKq1Trx7uQG23eJpuZdduhGldfClOlEGN/RW31qKUhkuFRzpNgOo6lusuQwKxpL2dQi4tD4h
McspiW07j3xQfLPLenon+rkWQydNNH4I8t/4ztci2Teyi8BmZdfLYitwMSajUfCUDVCVTXU7XVMQ
YxYpHOLvp7Lc5z3uxXdrp6A42dqkRYwPCN22wtcorA0YUH19xfi8r7QIfDUGT8XIkT+J8yo9ykx7
9cfuDN/YF01ztJ+o54bH/tNmsrEGuW2/mCmqErlkn8+XQlfB/VccXhSNdDao8cvlUQngkMcLIAja
6kkLSxoCBQDIYd97O8ccOOm6mgwJF2rQtDvYgik6sIgDCTlsL89j0EcK5Rk8mCOGvFwM/OcLNvF+
IoRRIEsrlirDtACdEhPngSP+zWpQ0FIG5OoSp8Y4aL/BvIqI+I5FIlpI8NGb8C41if8QIGoSaVcq
gpOWSFGNi09osLrB4IIyKRMQVp4V7JhYaZLvmTDYdFriRxDL67jD1tsDO8Qy2T1Pf2L9ImaB19vg
3yFY9u+brARl0q02neKS0HovyuXM1earSvd0sTvt3leK7hjErJRfDBbiINFPGisTvY8vs3JIhzup
6XoQVbsef58SE3hKyOB074oNhlHXLyERnsTbeuD61L439ZuJ4ORbB1htOVE1HJWxW3nNgB7sxFa7
hOkGQiJNgeBsZG9OiGT1+K+OsrAxezYChwNQtuK9fUDfKjUK7WxmypfZ5kofGciDcBwuK4pQNQQn
dauq/es10HiaNekGBCcI7aq0DFL3otlJrZ5pEaW8NscCKQGodXpEytAzcxpl8UnhIWagxBe3Ho+B
KWFE6KG6F31YQ1SRXSiACZ9DVV/LU/1Gz1OvwQygIuj3DJ8oIhZWlTlKStK4KQkeHQv2JHTdmgdv
IC0ZmLJ0duNrmTuOzCwUG6oSSOw05117DCoCln1BeHPB3rHMsez25sE+pS/d/kzWJ+pZd4b0XFt7
fAZoRDcqCQhtOQopNsZoQ/5ms3hB4+H6t2E882lTaAaZo5PdNsO2DQM5afWkekOOhee9s+7MB9UM
8B2Kh/dhs3ScfxfZfoPzZUCVyza/ovSO8T+5dJ/n67lNv3ZkGxUAq04lkXHUMz9ovG9ZbfvSOM6G
W3J10pVfBQ+81RLLdSLradHNJGped5kC6YlTC4/uIefsVK/tJKzO40i9pytrWtWwpGMUcx+cqYtr
RQ9iQU5VuaMm6+sGb8c7mp09bzUBUbOu+ZXQeATDt/F+K/aHa9HLAvWy1ujwDNpn+0FB4plXTlE2
pDP4uA7Eao6jaXOao7c7qNqCXppukJbXWR+mTXceciNHSQQLAvk8h9ZPlsBrSSf6hLyUETwEMG5t
ofuwfV6Ccm7Pnu2XhhgpJEFX0V7DRN5jyJ08jYiGEm79AGL60geI3Mu5JEdLQJj4DSI6I9XL9Yv7
hBnTejWVQ4djrMJJbCHy80Au2j/W2wCiFutk8WnOUbGuG3mUAX2UzzOa0aTyG0+UUocp5L37TuJz
qH7nSbT/96CWzgiSuxBY4c/iKUvfjae/XKvr4o9oklUtjwIs+VcQtl/cqDJmQfQSg4rP3qDMdNQM
+QWx7XhocYSS1fn4FMdY4pVocAUleF7onHS0kEeI3c5lNGFxFxKuSNnGUn6OlQgDR9ae0fDcYiNX
SAFjlF6nrfIfYQTXopLRHR1hl/2G70MovP/HGf3LPIhthPvYA6/QYTvaV/cUhPQ+BRJDWlFtyOTI
J3FnkPjfDJh6WgxB/v8Z5TNS2y3bxA87kq974rwYg4m9u/0ZbghobcWxR9kVxLcgg7YyemHB01az
WZUNCvezp7nkZ2UTEkjjza+/MFWV8v4IHtyDHgiCamOu9q96xsbTOCOjvhZK7Rqw72j9Lkd6Uld3
AWW0Dtc1aLnqcYcR3PTl7eg+I4W+O/nxPNG4ayHmRiaRQTjOjj6BjAvsp/IlNqxlFXkCWFXmTqnK
Ymt64JBuvl33hRVBsYcpMoU/kpBaV1Pe+AcGqVb31xVHh7vIZQmyS7PE/a2VeLDoX4/7JfHkzDQC
DQiomjPaj4ap18FbMnatnfm86jjz7JrplwsDo97k94lhmNwjRtPeFsA+EKq5+1v9K2Bbd7F+UHsK
6gqWFUSAy3yBjUd8/fKuE9x3wD0Glqdfqv3qxPAQPSrD/Gb5zQ/9OCfl/dXEjiOVR06FHXCL45eJ
7+sobhCy4jolBWDvU556Z/QMv7CySfF8o5U/xaAVRZH7v4dvS8V3DmcvymOkie7tDibjU3brUR1M
WqPUivd/dF4WxG/Ijr9pTchaAacZEi4lqDq3CzPAcxDwvtxKUwQ35oCZlYirWu5tEHstCTfGOw/Z
4VGc/YgdpHvOxpVWkZyL1TGl9znhsyowuvb0ncWoJzLXI9iutztIpTfiwLUYw8v/Drg+71V6dqD9
omrxDkwURwg74W/hZ/+ZP56zFAp9Ukpo3QB3DjkVn2ty8nHW6YPfyA+isIYV9fApEFSsEdP6mOzG
1odtp8hUmuPrr7DahRBsjlnmPNF0Ms8SU9KM3C0ETT4rMry3KxTPIdhPoYdiCvjpPYsSozscqsAy
fwXCXuAryv1E3BrtBoIjRZgoFVWCxV2HBdJrGTIM0ymaXf8zGgJaIq27gWAX4N/hsFYlYi+ONuM4
pQPJysKWyozMs9P+4YDsWKDZ5bwT9QktZSIGYnW1RUfF3OAhilwimDcVKUFgAbc9ADCxfBqQzKow
bLotolb8hx/7LFL1zms7BDUUxI5GSQ49Kwd9OwMoU4ji4N+xTlGPRUqK7zccIQ7D694hsVDAeb2t
jgSfvJwD/iopRYzluloborYhGAQK/ibvOyaqqLmeBtD3+/lDc4eX7prdFpRo4rnlALQdmUwMdmhI
4jeuetIbY3xsbqu8393SKXPsnn5kwT+zLT2NCt6qlTamHLNg6ivmbi37Sgcn14g1wzFN9iuD74Xb
+E/owt+DYKDOCaPg0HTbssZK6/9iweT+8dDwhY9abcU3F/qwI52MdZK9rCAMb6vgc0vitB21OAe/
r7NUpH55QDps8MEEfgc8MSurMxVMHgyo649tvSYSQlIu0Dcr6qH4/fFJ76Ev/j5RKfMK/V4pXeaK
kfV+Kku0L1gLcEnVH80njsoK6j94VH4S0SQ30oX6sP16i0BtUw5Sc2owjeVvPjfFYXnfKRaoAdz9
Xmy05kXMRbA0uKoqkQfsCH/1dWdpX/EUZ+w1P3b9HA3bAZILyB0LJ51ItRGFrvTFQs4+tDQfRB7s
po9nLKu4AuKdzHomDG0Oqyaib7oSBfot2wDozbHLr7dgkbdUJO+L19kHNZL/pKZDrLodHj/cZY3z
8keu7WYQ3VB318lwYj3/G9LfMCnqCY7BIYvUZI1oh1bb7xgyFKtHsL7TnA81SC5ha6kyCKdZIh9z
mI/6tH+XOTU4k8nAXGdh/433MatmmXS/1dIixCYcne8tfs/k93gZMDg6q0meKtXLvaejnB1Y0C6T
9GFplQjeUNQay2yq2H7Qp3gteXa3zUyjNt1b67PCjGCSaoxNqEYVHIdLZH6BJrkwuY+x/4Oek65E
nJ9zH2Sa1DIGSEbDY5X6bGtwdI94I0UXU0N1d/mlfr8vdBKNg1DylMKaSfrCle8rutNHNl6XGmsM
1XBiL5fDi/6Rr9h2TU6BZNLb5APo5FypkJFhJgXnFonqGz4qhWgkq7goSgXiPBM1Mfaywew5Rajs
LUCOHnIU9dZ2KaQrptrSJ3Ij2MyCtXiRg5AtWu3+eMdPTBgqg/t1NWq+bsixqUk8FSS1PPGGKQZU
hrgWQiXm0972hYEXmw5DO8DXRteOB0ORF+Q/6wyt4CpJ1E4pf+i/UdMzbwsrcbf52P4XExNxAXhD
EsDMcaik0vdd1u4mxc2bD9fmnyx1fXQFB4CGpo8oBBdMnbCX9+jUvHPxky+kThwOKbKts8UTS+fS
14zknGLG/AAzpqYqR7j03QyaVbMh7Bd5fy1KKXx44VeiGw5I5MHeu1mHW/z0gc0A/dNxslyH3REt
1myF2z1CGcC0zjVYHHWrrdC6A7Hcve52eWtqcAbF4sEJ4TgsSCc6PSz/Byt/enWENARHWwJ88n+l
qpjUfb6gpNaK8Y6STUbsfTl/oS+e3l0cex6E6RbIvAaNvk9h8x9ygXJtRPaFUGvAhMqQaGVyQqlp
/SJARftGIPiffCG3qA/LWE//ybyA0muzCeh+58sEMmlnAgbvdB8vNBURmKUvwvS+wqQJ/kJ9hWCF
jBc0jFCwdwevfscVs5HYNXdJazz2YKPcbkfECaWuae8/372u9FZ5TSDT4R3bYLppTAUWvJFMQw7J
91OtplwGO3YoKWpyecS30hQTcOsjCtdzrg+zdfp56DENB/7GznWLV41lMdRfajHC7g18n2Z0Luxh
gVzynuvb2RNuIjCX4GfzGoks8/EZyXz5ojmgd/i++hCIQXk/pQLu4b5QAWd86OxTtsvYiv6+LJ31
JYlvRR33mgZA8OJIWhI3Zlg2V38wGTrRu5lj1UeoqCz3xVnxI07Y8kvJnIoIsPijMtfvWOAA3usi
QflR2QdkSwlyAiW16XD0ppxqp3qvr3Wz+dQUgL0X8yGBjeVcY5p6Q4vSWFJWvS7Lwrvz+jwdi39D
eZ3ISDN7QLqJMHIDKMqbbxlylUifdwHaaThZrsad4ab0kcPDHA8xTIbBfWMJGcutA5bKYBlS8a11
DOSBl4/yNxkjwwym0GvKKeHlJuzBPT2oHSyvbQ22eV7YflkLZ41JN010xwYRVBcpw4M3kN4/qDnr
YGG4NIQCyU3bdp2PDDs/bHAzepLJnpbuniAPHyE6O1+xp1kB5Faw4fXtnTEgL5v6zhvbldSIUHzN
KVDw1Q4gLhpKOLBVSXafesSqDeBbqnoKNNOIDGhdMHFzC3vptSbY3s1JMfsJ19dU0dlaGWptvxiq
TTE9/do7ALofSTG8Qz+4+/8YN1JRkU/TOZMXa2uIdnawvynhp0t2mFDA9KdAlElnwDuWKemX7w/q
pSrolvAWXOmYRk+jmVt1m8gPOALPrcs0rrusO9yT/aqjpLkNR+zvokjUxw38akWlJza2FeZNuV2M
NWpksD1plPKrzKz/vlVvlaaMGmKcoE7iXCcpyaIX2YsDDYUmyFDSb1dE+bE62gE4QlsQwW/4kLca
aHZt4NjYPpRmNN8FSvhP+6uix+7jNoxbZAMHgDYzQv5OsGadXt5ear84oEJRGnRBAQyph7aO7TDq
C3NI5RYcHfiWmla8usAINHqsx2D1h23PnjSo47tVYIINYJ6WRg6ZWum3iYLV52F4weiY7SF0BfvG
STl3VMoiYahWcvGpTSUY7GHn+RGUU37O+ppYQT/w+B/UbiZjrabTKlraa8O3yERrr/U7B8HNYJYf
etFi5dcoWVr6iowWyNzHsADNt5tnoW2rtu+TIxrtHX1epyKTftr3/veP26/siAyR0emRoEq7UlKt
VH/Vd3cnUJWyfqNI45QsbP4EfvzzI9hNdmc4ROaYSjoXFhXyI+MopTAnjwLWAQoMOo7fSiM4fFvS
GoxWDK1n52LkeY0AJk6FLnLLxMt1oVeCAmvi26TujUr6OIFytPL8AVVC5JGF2df/779ZxCkum0R8
NgzJXPm4JH9K2PYXX4mnXAMN13UFKWhG63GhrXJS4Ey4HDkm+iEb7CP/z3YpdxuEchUlTHjTdwWK
DZSM51RGTRNWmfdk6qKh/GWTAHpD4s7X+xM/eWJ+II+DZlwXKAeTFwt8CPvd9XfqXeWzCiT0m4qc
LLGP36Sb5EWZ1WYcBBhrrI91hXBLT80S9eIJe8HCjmfuinr7LcgAEPT1kGBlZj/J5q+b2gXRS+zI
5REgM7N9F7GvWNnH25pYBLNH6+XBiStS6bJ/7cHgl4eHZ+P7PQVL79RLg4USXhx3tDkMAiX692GV
VynwoDYAO71rkA184/oP3/Rw58VMYbzhLKSxsfr3rrS/Pp/jWGrsBWB2BIpbG06Mq+x1qRt0PWio
zouR4HFItRPCplbEsX14z8UK8LLUikugMsrSPPp7U8G7+6T7R0DpRtF5FSpNuJYady/v1jRZC8rH
1lq2pq+3YcrIVtPMVxZ1kTl0Q6rZq9cemsn0ZOkYwqq32FrMP1HWO5yxrM8gs3cyMr5/3ie+FTLA
0RxHY9ktKkjnTeL/TeVA5d5bp8dzZeZQeKA2qIJbQJKr7U8Z+NFA9bFVMOKVTIX3zRqgkqw9MFqg
KNCI2st1XE6mvmM/vnsPruK9MYy+oDehrb5fG35tW74xz/N3Lr8EX8LhnWhjRBb/ocRLSTvRvuIn
F/A/7qFvBnFwGS+6a0erIoVRZ4w3RLVc0Vtn12GjEXjX1MBhZV0z3SqGr4vMl3fB04I6eaVxDUq8
TJnKVDhXmC7VsnsLz4EPti0i6/N1K08kSmoLYAh2um35Yz6Mv+YNZ3JcwPwIhjDusAJ1SuvP/2z/
UNQonCEC1XMCdUXvXAYwQ54ZEmPMXBBp/Cl5lgxjNFqhSCGi0zOUAROKbXTpbwemlplvAl+ZWAcD
jX+/KN9LKYbUOhCxdN/S1Tk/iBcihMmuDOlW34tFTrCFE5oknkrfj5M+k73P4lbTxvjJ45ieb5ke
2BKlNZqAnpyr+AqJ0WxfqUHLr8GUnSrPMx2hfPiKLdHeYEDZpNxaRt521et7qc/fZROxA0419nVV
AD8KzeXcaaKudl1UOsik16u7osH4PZaaTaCmxygcUvR38xpq98bhUxWeaSc2HRbEQsu88HXhAjhY
7bWcuqYskKpAMJzckav/ujw4TRYE2r1iD5kzrLxdAEkjnLi7QFK0DRX1W8fqApL8+SWd4p52Hq/A
5N+dlBtfaye2wscbl4GpX+HR9UNuAZ2kizIWj5aGL4h6EtWDeSDw4jeuqaE30qiXpDRRFwh4NTki
L2V/o+mNAOVVaPBTFQDU4x+AEUBGkVX5wwtGg9OtL8Q+jr03Gx0bwTTc+j0DglMEH8fFx2yOeXAA
CY5hHOq1RpL8JHswB9ffGWuoblo6/ZarALDxKa3zsuPBcYad9E5L+fRFl4s3nDuinb9XxicDkVeb
C3o3d4JjQO1/DlauARzNqEqhIvaHF12duI0SnMu8vhFDWu/5ICRSw3hXrecYxh9Jr8UeTXAGk/Ti
v4NORze8DYh83p3s3fEpKjGwb4lowgo/Hfbu8yyNyf+3ah3J3FPSt5fqx0DkNGm0kk+BgoUDQz1x
Qyoyonu98QPxejOs8NviCyAHmbm9gzzzE49ZqTID1ssUo/gVZR7o/2/zlUwy6VdORQNx9LTiHokc
w7C89uX6Wh65tLqKCvxVvhXkWgM61DZAnNFSo50IhrNwix2XhvgjTGdiN5XcdP+f3j4J65fuhgl+
cE2aMxY7O3k2Q7VH1NKdp5gRHmj9Jz6naSkQmTpB1suzuqmjAddbPUY9XaVYdf4jfrBPmbdE7ry3
l8LMjosa3H/i0WoC3NbzEihbo1cNP5Xb1tDSXKTiUZbFkOrIvx2BijcaHMt5NEhqJbkJ+U5yyPj0
JcnpIYPP01niXto2T9SdPR5fr4wRFSL8M6DUm4bqUqXI6w4kSFucellnvqF31J041IqNwLQEmCxL
umLAA/injE+nVbl4Oiv+2TpHh+vt5tHP/EXaU6KJinyAsysw4mth8eEjBFRbBvj4bf1mKlY7Zar4
QJwonff69+4srz5Ap9PT7qV2mSszxEbTyh483qqjUy3jl6s7lNl66Si0xaw0A6xWZidH0PTnZZpf
id8nlEBOrVp4m//rgfjzYaPzdTtuirZLHt0cBwe7qIfL5l0xh5MYfHsEo0H/LFX6RuDE4upk0ZdF
4InOJ1BQLyKUWgPRetxFxmNA5/ScBck/6cCP+y99Jq4pfJAuJfHImnFyzWHshlY+rPPOMY+eJfDq
87NQSc2gSwlXP94wt2RvTjpM6ROUqAngRrXCKzSSLo7xWWDk9FoyQRMg0eep4NRI8B3u9u0oxJ9C
ibTost0/XtocVPWj21uG7rAbO6mHFX216tNiT67I6Pfs/IwMtK8+CU/XYYvM9LLGzfmZRJczK8cq
kjG6P0DJ+lymyMj+m8gi3eriednVv+xtiW5WdZCrVi8gYCj+XVMQiqKOF8KTA0xqyerPAIgPYU8Y
osZRXm/jKrliNllCDSHA4rX7/oS36Dlig3KxaeNLGbhpjUcAOeDt9O7Ilv30SJaG7ch72nCZVwH6
nPLYxbjAmjrpKuyKfMGUg7RMKaqq2lLxSV9+Gd+w05DawbgggyZj9IC2d2up0LsfOz220mdrlhu8
d3hkHry/C1MgqkIWg79+hugaA6jXmsVagEBmhiw+nXtTBge7ceA5hV7d1LHUT+4WFi9OLPiqArRr
h5GoU3t24y06PMT+cxbh210HaSW/OH4oPl0BPJtkgLTUHE6uoKE3oL0pMSGZtIjvTQNdlkJdU57R
a3MjvGyALdK66jPB9/AjJRB28JMKllQ2k0E7nwP3+PCyHm8H+U01BSR//1WbtYP9FKi6jz5/03gj
BL1zIVqSJvd1ikLPQwOcSL7QM06Y9NrNSj+N5X5VktUh1s/aJwfYDKe3a0TZeHWJrKvEMVczrjml
AvwYCpXeyzyIUzK+e81V1pnA9secTBXABQd8K2WZlM8cb+IoySoX59H8qY6yzjJLkcfigR08Dupw
CZkuuQFk9VXEwtHoloc5e5as9Q708agLQdrH0ap1g9X/+fycmVzONBcn8dSS0Q8bmLNeNNEwadf7
ksDctu3pGATN56vLgV3CcUC6CefTrBfVzmrV2Uu54JUHNA55X50CEYo7OcU52gi7mfIVMurAHeTV
fkep3zSNPnimrO04DZIv3z/znMDolAYC+EFAi5UhBpnQX/WwLO6c6zomPMdXL4F/SmkwLSGafwjh
cvthUXn1u/mLljECxH8Pk8ASEOTQpu9ljewUBu58bM1/2BlPd0+AKQTTQVWc58CQSwtBsgabvyVu
w7uzNpWq+P4oFhVEVA/9i4dWFwoJmQJM0rJ8vf40uZNIIelPQKhgmQEQChbuag/3My3uk9uXgTDK
HfdmASBdQGoJ5hRx2oFZ9Xho+2oOj++1X/g/3stMpiMn8kMiK6petzFRxSUxxBR5apjguXU2+uIv
OBt5VQWLE8cSNbvQGDQfV+8eCtY42Afntk0tIvcE0pPAimYXzBumTMQn6FIPNojPwwabnEIs70Tr
5PvOSwlUrTObaMQvRmXHGYeQeT7LbQx5/ihqQ5jY5JL3UPTldgGZnGYGkoUPRZlHf+G6Fh91Q4YC
0dv/XfBTxI+T4xcXt9HqIuULG+iWNajyjyW4ht8M4fA816dMu1h1asm8DBvcITUNMEBnPo03Xh5t
5mbhZq9fGPESgoPK3xkSUqhKHfcRoX68JwKQ5nrbZO0rRvfVVY0/MGyx/Xhqgvc6SmnRI6L/pDF9
z1IkUCQ777grjFwQTMnMKRqx0Hq7xzFWDIzgCJLcvdLpsJYQQ3JMdqLexOiXu7NpvwD/2vC7pDRw
5Rdqg1CQGXRD7riR5sz/2IlEgCelBnNYgNV6HIN9rv7NRHWF7ttZU5PU5MjBH2gWQgNpiSyj0L6v
joS2kCwu1yTdLnYT4QfVZhLRMf4fYNVjlQ+ACxbEkVuDMqsIa1FUTOGBKNGcBuN6M9JJWQ3yybmm
PeCwEOcnak+d3K3Vq4YRZH9j9G0mOeTmyXn93PhRX4iiII0xDwKlaKoPywVWbRhzVmcDjRKBQKC4
yAcGgzHZZ2viYH1TadDE6g/xIJBOhWbb1vGiJuAd0bBxknX68HeUa4vvr7yGVhu0yLNnu4OJvQUV
ekSms+7IFCgHe3Vc0Y7uTb0byTGQBgOqtwjfSudbO1ud1TAv0JbMqB/1hyn9M1dboikHBp74/Ezw
TY4QEJ6p+4DLRqdvTl2PxmeI9CuPzeEM/Kb7bdtZlXqyUvQ5ZGfpW7CpnEGD9Ux9xdrWf4fYLR0V
VvS/enAUqLyPhV1luktOqGsjkkfcbRUgxln5GdYtK1R3FLXJHGd4evzvsOaVuJ31wtoa83RfKI/Z
8MkNVnRxkoz5NcUJ6i3kTq0jHxdtXEvpoxfZ5kzSJS9JlUax+rLZnN+PZtsq1t8MNqpBkx2Mrnaz
l1R0JBhtL1ywRc9jONo8SvIRlWqbGOJ5qtQi4h+Mi0bnrDasZ8OlNoXT2sTlTMPDKjK7swXMjRMi
06eU4ILdxEoM4M+h2oXmHqMGjfVFGp6xGqFbeT6P9WXlM9heZ/OnvxmVnboCPcuUZ2eZ/mZKo3oH
H1oCRr5vs8Ra3cLrZNChP7vF0U04qKxBmIszCGtKD+glPZq0vRch+wJ+LEGE5g1v2Wdm5XuaVDkY
HsmiPo6oMCTgmAFmfX7oARTrAhdWaF6oh0avDwe2AA2pEO4RH9gBKZcPbfgESPMQHcjqZSI+Iej3
7CfNI/wByKZQ0j5UF81Yeihw5lzOX2wQwqwuMaYNGMiCGyDDz2TBvcvmzfzlWcQyubay17yTRpSL
SiZyHLD+t+ERgLG5jBdCSO11SybUvAFtg6b0epE+CDJZL39hSgsq4xUqt1xcU2JY1rcNYLJhCuaL
/GOrYkBB7Xyhp1nItVCGSbdWenlewpTUfSlUB9jROjSCZ1hjAhShfYQEtXr3SFBIF3MMxpRKM9iE
S5xl6rdnY2J6EPxhf+1KR8LIJe9Ra2a4FmRDO1kL7cdp/61zauv5MZp9dlrfenGoNAub3eJMXCni
fCHphs0R+HwFGtpX59dsZ8M8C+CgC2Wj4vwZjT/OXTs82e9uy8k1wU8xiJQ4mX1N7sOZNEPIkN2K
2nhkxjpxMfdzsxlrlJ4lGNh3R8a8uGjy0ec8XXxyhkc3XC9v5h11xcwBNLq6u5M2P015sll6Dhwk
9Jbubh6OQeU0mil6Sr4zDf3DSbdZCTSOiqrIAP97kdExVb3CRTs5xrlIDU4SZVc7Pu6J16CLIL2U
uw1ZTvQi3BIJwsqt16BVPSdZ0M9nqN4YMHHkdve59TB6YIhEFA7HUZhNsibzRLVMhjkYMqfvHbxk
HzxFjudwn9VSTgsY1r02e6ZSNGD95FHuy5UXUGS6GCadVAVh2mXlUpJ/zNUFL5Padtz5GRed2s+s
jbjAeXwfPsY5sCpvJZUEdHFk0xN98S9iWVPrBt7NIUEcJDEz6d5J+x8finnkGtLimgttrfL/pskL
v1zvFZ3RfT+xHvSLcES3ixd+ghD80BZXhk9xWHsWO8U5w9hKyWLHxZoZo+5ZhPjRhjsl+CpbCT8i
vhg3VJVAfjJX0hatUMgXjggpFjNtDMu6fNjfyJygrrpXou4xnqb1ZlXr3OBYTMzKsVg3k4U4HCyV
n/92tALIpgnaXDAQYaPH1w1JPDcoqJu3it5J5NXVb1Wj+NXVYozEEH01RFlKSgfloal2Ua3DisTk
F97OKjn0QPpg1F7uax6+W9s2WlLD7NISw/HdHkwEH1RS9nIJryFJgTm/EQSZFldXjW0YfZpr0JTz
0NiQpiHiLaRD1VTFs6cD7Y7xeVp2Hz+GQoFMJ/uZVxSZz/19E70LxWDza68yjiatMH6iSJ9aD/AV
g8eYCN7y9nyvm3r+B7x4mJDRrzmmIqiM1fadkJkpE8XG5V1iNbmdxqlahHtUEklqkv9cDLsBZVqj
fvwxDhfuAfoo64hBnt9xaajjd0nsleH77hwlNci7TyvJwmY9Nx3g0bdEFX9ly6SiNO0svoKy1QBI
PyHq2lG/UGMG3aBILNMmtycvVBQzR1jDWH7nHOrktfYxGzNR25yL4ltkkDrGzQzPgAP8cBgRkaV8
6xdt0dtv/fN852MJDffSq2B4psqNdZAuo9sCctous8qOtART/y70URFxlMyo1VFTUE5vEW693XR8
9pFWh5B5hRj/k6uhDGiMjOSp1LCdHPirit4yHDfL1YBi0++P7pZI3SYhdiVZpSAqPIvXO3OtjY5o
1JvYDHpV2klfJKqrg6bm0XfwUapbXyBmvYNOJJVIDNWjO//Sa3xAFF9k+6BTaRCcJELUJt5brd4J
XnO9vNdtXQT2TsgLmOdEAlKJ6+JLGqsTjzyQsewyltjj3A/K5dzrfnmaQwl9lbut/gJR9/fRxHhg
PV6BKuWFL4zt7bkN5IWIUv5nNMWP8JpG+Hni9+/GvETGwhFPkQNHqHkmWM/oXSP6dwxjqni1y0u6
snsP/Z4b+KKV/uYupCpgy43V+gK/y+oSJ94JkRLapCcBx4VVw+dPJBfiDqJxSjuA8PCeU8S4hPqs
JwNS26uFhZSgnKeGxWTglws4TrLYhRsUmXWT0DpmF9Ph4fjYDKjAw1XVT6zJyDEejlI/780ZDza0
AStXEE744ZCFSugzrvz1LainXi5gNf/pjnjqT5ut93BpsGveBXrs48uV6bBCXYY65Fj3t7AXooNh
9k6jc530qYH49BJfLhTwt21NvQU6Vi/y55Gwh+NJ6VsLLZ74IJM/1r9o3iyuNRCdyhJmws1j5ZX+
QThau+N8IJ7GXHnOcGzHdgYRRBjJl4XJs+in3QncLhM4e6YAU8aXzAttv6mn5rUJ91m+LWmvnE7E
4aWOOj67YjJ+9MPWkRoKS47h7Ljj2dy4TVENHaka7kF9ZSEQZmh2PiGeKQZ4HRWfjJl0Ug0ZUQH1
DlLotjHERzcl7/piTUEwrBbkUGmxYc/H2XGWvgruQGkjvmu1Q39PnRxMcZQbqCw0/SL+J4SzQTSl
C5ApBWPWVdYQC6JO920+XUsO7UoWV/PBBjBMSDblbEq0GUlMaFKGUvqSWGWjFDXiUAFMM0MrLlYI
LwqDDVliWiUb0nxX2x6f13Osaz57C0PSOnT+y8WJ8S4RVZLXLr5dTXucBs64/9XlfghuQheW6Ceg
gci/fndPBdRrlC3WzQKRpvM6zJPQQMQ1yVIACxe++qgxcHAdaVsTsUsYGS7sgButF/iuylbS5bI9
hWdCvEj1s0sWiBGw8RdSKNSmx6V35wiCVtRKn0TxkejZwjKssMU15Z1B61pAEM9kA3OPriQV3mul
vmcnxANUFwPz10ZN/fZYGrMJeij0H8THHp0XbpO7wBRXzhW1OVFS56KMuboG68pY6yqggRhA+cx0
kPYoV/m5fCqRq2LyHBGpxF2lXhR1W5qXf2AQOtEduuQWna8r2j0u9xvWmyqiqLwhCU0MvzUq3XjM
h0dvoGN9rOFAmdjZ8+qgB+1OKAWUZdCtXip6i87rCUXus7MzicsMiBy1GFg55VPMObK60dvW7y8H
Z2SR7SRutFUqQQoFecd3OEO9MxDiE5Qi9mdKVUixyunKxJeY5n0i9cBpkCpnLUBV3T7tKrnkBUzW
CZqoIp1CqJtpZdZiUDqtITSkMQb7opGM444i9Xr/s4m5IKvrZLboibHZJQ89z/ddTGtYbYocWTeu
EsE1SBPiy10pmXanJ7a0XvUUHH4ePHTBYMabi2zabRRsWKhbUEoFHjnOLwOSvENZaMcwa7RXMJhu
s80dTKGvaSVkvDJ6qSIdCFFp1NH/pUg+WDC5j4IKs3lH49U4LrP9+JrLjFCTNg/DfREB9vr4sl06
GoJYDkpQTlFdQQBqj6zQ0/O0H/Fwnury0We0IWIAIRIWSAbUEbSuMdRBh8Jmq/MX/34YitSo8oVH
2EwywAshtRiYvLPuny0LLcJQ25sn4JCrAViK0J6l6ssGQfXGUzw0n4Kl3RYfH2QIHsmZS9c+3hov
F7Ueup4LnGIjycCV0kO/cTJea0g1UaHul0fp96yDKB/I3QDwybDHNThfDSExWCRtxoXJGQj6cUVu
vhEVlyrKle+tsk6Ox0AR+RgWPYN/vfo3yhPVO5DXttip6lzP0KmDDnlrFKH2pnY/+x2OqMgSBlDH
AC8kg79VV3c4gYi/xv9lQIOhOpEpQwDPC5YkFm1XgNos2zDBtHRcbYK/CyAZROJpEvLByohJO/CN
tsVLFVoMQqqnJ39xHBrEHBbI+sTQsFqQ1rQ2rii3+kT9chFSt6TqUWfPt1Ks8vfw3w6STrHhFcdq
7+BG/kzfPEnDmKVQk/7mTS2G6lIjXQMm9hyjbENP/rBd5rDqbJqgOAgccHELrK9uR12Sbkc7VO47
eaiyvUp9dvcnMSnZeRfy3yWt8i4p/e4aan5fUK80LCDQN2voSH8r5K1kx8Qhi+FAjdNKTjJQy19o
90Z+YHUp5jvSiDtQPW5Fs0QTp35x4gGlq8/GgC7AdR62lbzbmORJHt+ZyBCRt71xDxe817DPepij
ebWYy3A5JQKLtmFlbGDCmpynyvKEfjmc7CIGVu1hce8NUE2bIb6iXFwFH4vVk3bT7YAX0xlpoqnn
OLQdHnYXMYfSqe297HCqjfoz2QDzcIFwsoSyTgVPfkaHfMoPgDqDDkB8iJ+s+l7M11peKCkgupop
pFe2/dUxYq//H18aZvVfIBVA95nnF67QZKlBwgbPlRmUrwnGDsfIE7GsQHuJLoPG5EAmbRPtA3nI
26sx+5etDwshkB/kT2+EccQDULEyfDt4WjwnJG3rLirb/E8klVF7f96SkyfxDZazmpqQCM6kgibC
DO0cdoiakWV/jqR5F4Ac3CKl/AOss9PsOf7yKn+xOVOceKbnUkuTN/IpzfReiHQT+3ueWNy0nVMD
ZK5HIyN+XIh57eBsNn51szyZzHX0CClPGZN4xMBgIZhqPT5/SRIE9jFLcEyp5cSfAbyLnvw21g9N
krVQ8bqJ91usPsEgJuk1/ax+VBfKCTCxytwo/LEHJ0RtOueK6ZvguSIAKWVQgiV2QCX3fSmg98Ws
jxmNsPWQa4F22+iIbvvyxZkk7a3eV/B9WFUB8c1M43nVEmh3EGFeQ7QDSBJp3xxDEQZ9WUhlgmuO
p+sJo8VkiZIdaSq2cGFBJXHd3gYGI+PZgVisL+FvadvaQVrrEYMxmcIZXsprh6y2XwPUCn/4edvK
8lfzyNwOOmMGUWi16NfqA/OCYImcLMDLqK8Hmu3hOCsK9lLMtbdibAbfwE5xKt1t5w54E80PS1Uq
ov/1JeKlV7w5AllxSmVoMiOKU8+Cs+hXcCcW4K2PZ2bJaIQMmTBDTvtLneE4IgcLT/uy5GHy5mU7
/ZAvsDi4zkTTdwzW6aFMxuFSdT4uoFvR6MBe6rTFNPKllXVuoMpiSzyrue5/mguk1o3Jwzph3791
jLoVgkA9r31obtCErnMClkVuYMu/gnAn3YnkABBks/yMe7fOb+6KL9q5u/s/0bHjXMrdALDqZ0G1
PCy9ZQnGq94ciIE7BLy3XxN4dDlP34jaVNvVUSdlTXKWbMq76O2QQ02GUyLT+09y4IT9GSFdSkFI
QE9bJ1CkRv0f1Yppz6fkO857z5/E7509LWcN+Jy8WxB9vHaC5CTnKfGYAvvG41Lyle/+B4nP+At7
DnJWPL7vRqNFTAge3+tE14V6nppbKLGlbdkQCWiZeTriXEbBzDQ4IIWKe2zVuC+nhhSF24lad+3l
JRtk3y9gZE81ASv3ppMVhkrnjXnsMK0i3E63CY8Xebd6Oytbi8PZlMrQzXu3C/gU5Ro6C5nPyfb3
ngKX/Dj09k8m4gpzg0xIJ4KBhLBLjOACvJN2UOk1r1Vx8psUWzG7W8MCTixvF8KsHVGECB7sarM3
RFVmtCZKpZazmtjBssdH4Ln6l2s8+VQr/BukaaXOotAOQnt4vjlbPRcf+fTaeIy4bkPgQnzpUvsX
fSxw8e5f1l1Yt8giPV3MuAEsAdsqjCornHHzSvsqGkg5FMFO9iyUeuWlNfuTvug6HD64PRcxDY37
z4PJvQ80hD5gmMD/pOTwdgBmfL3FCi18jqrhD44WPS9iApr/bCERJkceoTaTM7Ef3rQ8AsSmNHq4
1AJqIFxlD+aZlozvKlBn5CdCQRq7PBzG937LwnkloYfXxL9iPjIM4vQmRSJCAjHi+sh7pTwDRp8V
pWJqJ4sUEI1Ehwr2dFchtozPVXq69i1NJA2AaxGciort73MkzDQhsy3Xd2xhdL8UKqHeRr1IX8sz
2U8twrHmLL/FDVUE59397aIYfRWQobQ9Jg6JfKPhRXFV6HYQvUftK8pV5ToXrkR8XXPR2j9I5JUo
tneIvinHQIPHNJgsXGPTWBpV62eXU00zPWZpBIy4gp5LmqgmhuNXFFWmvNZEGVQkdKcJIW5KX4At
Iqz+yzUE7B4YiU19CBSKdg+2hfA/90x3oyWu+FpiQCHC+IkuAxuk+wAohkKna0YaIRHmruvY2wmV
Jb9bPc6GfYHyYTL/waoL9BJKcMDh43TOJOqgYs8+VjmQdw846gt0uJR5kI9TTbBkk1DPBxctUaes
lyBwf6QhXEmcswPoyPMir6i8Y+ifUJDK5M7Shy6CpRU9343JVasnNZ4n0W3e8yLy/27Abi9G5iPl
Ij8PiPgqX37OCoRX+h/bJTULtkCb9vqRWoITTnmYK24dAjoeRoBRhCl23H+27KhCHZlyPz2IIHOI
/2Kut9ZOx/WvDaFN+smz8VyAl21PgIQSOC5KihQXDQLg4RpTjLyVVs1ZRm2pRTJKppRB2GDXmpg+
x2MTcAI9HG7K91TJULIgoFg32T09EmunfDxare7VdJu4FXO478isPBh69U3dAOx8xOM1Jt5nE9vq
kAY/0Opi/IgUEUFBkrNf+neeIkzHp7Zz0xeZNNVwnl32MwBbOhIlmy9aoCzAukNbzBhsS84OJW3u
Be5/EdrWUMQHfwdNp9Fwsmx443SBHmtQRmgHZdpLaLtdTfeEjEmaxQC/Fj9s5q2W1ZiWseLyxnZN
gvLIVQzhrxKqIWwfUN2veCmBvIt8R6AoQ506XzBdBF5yIKsDRkl1f9LevcDG9QLm+ESndVCB9dEN
I2RCCPn29o7XzFL0m3eWq4rVX3Xgupo7pZ4xD+hWjr831J1FNJMvkjA+gGxW5jgiVoDllrFr3eQM
B9mF1Ccvgc0DJtjUvjgUydYZdkwcpUXL94IGAX27hDzotklXftK3CFRwrEstvpfZb9Zrfab6bZ6Y
2H39uV+iSX0DrWiRJ338eyVWqFubKqQLt2TOR8yAWUjAEb2yjEA8qUwyQrQDS7hXGNn/ciV+vHzt
3VVwl8sWT0zR5OAVsggKPbBzxH4nawS0GUBjdxo1vH+EdVh7DI9y/9OZxT+FL8R7ZrA7VI3lelJp
AxPVuzNvrC96ACdSSgYLIYX2gRkUMBrmU4cw0hj8bCxZVjpostsGm9CtyI7STtPZGV8awYoEtkuh
4BUUQWEYFFdKq5RAGcW7prLIuA8bfUJiGATHxRtwERUqI9AExGWwnLkGh2VkHrWKJDHWX1WmsaQa
jX7TBtEJDSXG96OQzwSUEVUVhh0zSdfObFB9xrtxplxfFxNzRQ2HIJqiYf3HTouD90ppuVt80R+K
4A36OXOUfIEsJfimHLXsHsTZ9XYqw5hAMR4LO/38FrsRsDJh6iz9NeF+urTwxyk93F6I5dTPDElb
X0QwaCKANj8wzl1khXONjFkWfEdAImAknUUUsuUXsvrYrCo9jEE8Q0dAoUgg9mISGzIzOy+vuyfp
IZTTtusY2flI6oia5aOMba/gwxCXY3ruqNd25Gr4iGrvLxY1We3gt5TKW3W21ZRZpu/lX5Az4Ddm
K7qyZySHaTM+RWYL1Dk8nwXIp9jWjTrr8P0caLIbPlKRcvg+j0gSMuFuZRa+amfEfyjPvuToafZ4
b5/yMnDpf1w6280MFhmIz128ZWPIb49XaSE5bFQnDAoxgOxLBhbhW6WW12IhhhgQ5K2UpL5Hc3Ju
44thXsBQxBs+Z4eqEjo3QGScbAHPn/SZFkYcyFoS9JGsJ1x8MhSAlXah+QQgwZ4ajaWhwAJUI9l6
76TxbyHvGV8koaR5Tw5I8DaYk9Xfi7eehRfk87GT2z6K5MSoYPox4f/O3Vsaj4ilFkwoNq/kFoQc
wI6e8B8/6UY8QLNyjmsHDL9bltjpJWhq5VsSmcvsNAH7X/Av7n4zQNwya8mNC9PNzz6JthYcKDs5
ODY7eqjRztoyAWhoDBqx7whXvifr2ky/tvYBx2+0ZmkT5hVESXEs0FA4Zz8s4Hax6HbRdLGeekxh
O75NB7lzKl0JMU9ICsMhJWyYx9qfOWcghKJyftu1iDEUV+vjj30bt+sII8vJ23OedDHMuc0xi4dK
rXcRWrvCjUPbiCH+wq0bEYR/xzXrebyOWNegDjdWERM+gSTRZz+iHWyOQzIRGuy+JxLYVAvz36vM
2Bjs62ACqeLA2I28/wxlAwHyC8baePNuqAytB1FvyOoDeog7P/a8kGMdixgf+kN1PGbWlUnjq5+h
DSoBAZd81QAdAWzzM2lcH3uI82L+A7dP4+az8CSSl1QdWR2c9Es5Tc1A/yxjFviR4sLBy+89YuTn
XQJIGSl7TstK7KUzwT32D83apt7/fQHkL33Uq4Ngz82oduhqSBYu48muk9/imDwdwbLGaW+M+m/v
tPYTYMdcWUd2Oeo/tQBGmRvkWGOJwoPSA1Cb8v/zn1cj40/moCZ/y2PwWN7gZa0UlWysJAbEFJOt
s7z3cb4jCRkce2Pz4m46Yvn/ztApBrWoq/xxQ/SQpylQa8ZPOE5j7nXfm9lmuRQSn55pstEHQ8jF
yEkPxSF4hJ2sh5SsPi5TSE7KYkeuWqwWoZedXr4lcGdp65dlCc6SS/FDWxmQxmkMp2GQ6yPHTt5H
YjQZxwTo86/XpXcFaAqVMw6DnSqpqdNKEtFH0HfbeqMAw7nguCI/6KB9eCC7K/xp2vzX8IjlWOnR
BnT3IdmOUiY0vno/D7FQhwnYEfxj8+W77ZO6BNDqmLA1Rzf/YX/jw6jFkUWCprZts4xCk1reUx3q
LiYwzZoP2wre2kz+PYZWBmXesStu4WeUse7ZjFPLHBZNuXvjPUXQ2R/UY9p/hPjWfLfiwmginTi0
gKoWUYJ17WHnYV3CnkQzv9XAAFDKnGJByrm7V9i7Mq0KosNRJS+Chk9/Ilh+GfDePumOGpzTiNvr
VRv9NpWoSTOepVNL6FtkTKFk7ns+um9U2A+k+nq5MuxplDd4YmMy4frX9ClpL+MCxjzCQFMinGFB
//QKDrU1AgRZ+fUVTxjgMNg3V+8sNAHv1Eoi5Tn+ZGHuPM2AR53tE1SBbjzj8PPJW2KczDSbw1w9
onM60Ta/7YaUQYeijNbrFwcpNQGWp40YX62eAu2yz8U4zBu0XSrnxhDBqcGuqjo3CoMJeYb+uIKm
32dPpKPzLXchduO/XgbAMlABOwWiMv5IzFcEdQWrii3wJ//zJHQKNsKpEf+OG+4dVM7SRgVrCR8p
PKhyx94MinWMD37vJcUrhcqbi4WTg6SG+heH3zlGtdAj+r1WgTPG2B35MKsOSKfIO7823YwE5ncs
i8SRBocVz8TqAC9UXktz1QKPDe3tYh0rlxEPzS3CPmqAqXydOIM6p5uS/plFZnPy5WRctbfG0Ua1
QkxpqTnIoB/LRiIKIsh7vyEQAL9OFO5M0MP+RKOmM0A3Ha2Y+UhJP7nadf8hJqRMYlKogjCKCeh0
hqo30kelp98o9fus5G9C5As1EOk5/7wRrPhGP9CSDcdVfKQNqSbkqCjri9J2Qa11E2xgSSjRAEGs
UV/VV0wlUuMDrTGkVwXzaxoTIRcgqtmOvnc186SysTJHFi3IOa00TCd6TeyBCa4Aszvbl0nQ6x/u
12g9fFho6JIMiZNDlmy8B5UVEkpKOtnWgz1aLUnWQA9gTQ26GJOxX8mG2kRoP2/Vq+TMt+czl2U3
YWMLvA58iBG4Zp+O2xtW38smbEKL3Bh1y7IuMa1uHAvsMBARk9egZDdG1ppCjBm6gQ9w/KBSoo3s
9UN05Ke0NxOH9nNbw52zRFp37pVtB5khcCKroLHhG9EKugsON5LkiJU4U5sdyb6EpSoPWCqBErjl
wo2YbTBt5K3id9Gj0REPVg354DIp4czIDKLMp9oXnY4GH2VeWEl+hPengBrePn2pVD7gkDsaiR6N
Ko6giiJbaXMZfxm10GT31oYSIoCmvOTepklsaXhyGdipd5TBUWtNlgfuLIwU9GqZ4mQ/ZVTt4mbS
J6MRtFZSnju7Eqc+i4Vdq/evKNEeY6or5wIMA2WYEW8NZ7vCJWpH4VCYM3xC82CMz+RtWB2CxVIH
+QEGJnud5cNBxW25nzsDagb42CRMzvzbEF2T0UNmNH6PvgypTOyoW6FfZm8gqSjcreBquia2q4Rj
fKPzonXvStW/VzKL9uGmJyZuaOD6Me+moAtMhIU3SclAXh1HuNrhW7WuqOb0LsG/uMC6IOdh9ucs
/hfguly3jZZywaoa6ikQPOKzCFofJ1yJimSV/7buoiYgDNLgXfgZ9dmIzRyuVDM+Hf6xGMFfEGZo
Be4R0nzoPp6Bjl6ZZp5VdIbUekCIgINjbz5FpaRBnVcJX6Js+gCYxjqa1RtbWYVkd1rdwJp+hsnf
JNn+Txg/Y2rsNnB676uKtfTrHSy6B/Bd3wBiR8hD5s9VuGRiDtO2x+JZ4E8V45OoFLRq8GSGqFep
T+bctbSlebP/EID91Sp5ai1Pp4PlSFk64rtrf3fLKcJGVm4PnoNlqllw+b/QGIg7I0SuHiqSSIfq
zG+v87w9V40gp6QFM+OeSgfeclG/GB2+i/ugcQZDkjqGhut6ep0/DF4uUetjaepHbZ1+yj529eiU
wbNEN/FXTfL1TxDXA6jxYkZUTjDMda+uHcvGVZP9hW9IwT4TWHxMvLgBNt4ElF0kVYF4vwAR3Yuz
AUVXj2UoKvd2nWO13fRPY8kJKW9vSpnA6li9NTuOmkDxQdlx6IrMjfecxF59jTwFHXxzRcdpjO8K
5b+TnAqrVKoEQ6D/2zSCfEJRZmFChwLZtnzrw2EBfANwCUOdwMixJ/vYspMtxz2KY0nNkqz1Uq7w
ufeQHekVXwOHnalJfStKzYwfKw2EEFFXfgKAMMDniz41Hy+xAMLXw/xP2qrQO+gq/JvtsU2RpacA
GMz9bUoihV1+E9QaUXevXGZZJtqWXE0tmLyNG4xU0bx0qyIUOAXEuNno2XI1Z6l6z4bZnR4NisXz
Mdw9ZDXst+DfqOntqievmJ6oHXLy09jCpZhAusvfBIOE1aASEdBfPY/gXP0DTYGEmDWWyI6n3YpI
3x6pWRiQIy0CnuWgDXxqb938b5ds3DFimZAPYD1v+/Kw1dVRn8wdPu1OTN4qsVydY41XzLbKMppp
SbIfzbGJjS82x/vdm4MXSMgtkIlFSJ0M+SOQ1IAvbIdWDxEAaLUqvlV/u+R6TKSioGEZKnXQjLmz
FIv1XVvSNIru6Uitn3SdPMjLiRFDZyTjejS14/TBaCVkQQsXFKsCh2DlJUZlIMnQkadI9fq3U9he
RSennmLCsrUzMPTufU3qD12X09ZjXqM8lBu+eOz7ISjJOD4Cfg5Ve0OP+DiNNy014jaCD1jluRbO
t1upK22peiwr5UuH6I9EjRbxpHIKIUQMaC5cEwQgNshqydexAuWeox7jeTXMi7NOEu1jnLPTIZhM
aT9Ei6QZUqrj/RUX3fNwR4cKjfZfbXW6LC2Y78HjBY+9F2m+7fpeY5I3GrgQPcozQW8WlFdQf6LJ
CFODo3NDUmfjz/SXgEWLIQUeGTpx3xichYhq/EYQTI4PBW+ACSl0iNLm86q2sSfaRP0a5ZgYTMBv
+ECPb1erNR0q3x21VH5B8wjp2TcXfely1etOy3ric0M678eLESik771AzWsCraXBwfvYxIpY0m5o
MqYV3i5SjYOdftzdJ+C+OUVFoTlLRnKn8/b9ZIUSQRQKnVp8r4sd/dIWAdsgO19do7P68wWcoV96
UcH8leo/Ya3UnyqvhYAVcj2a7xRAiSrE+4XwJcm/VQ4f9iSqDuJVcEIlSXsrxpiGOrt2hW2ODuDj
rp2zhsM/YuAkTBw5OP88LRiujK0wcc2kXa08VzZ/oyRsEg4t8v3Ndac3zTKsgXB64/7WUrjexRZh
LzqcLqnwu1pzYSQ8NQZIL5UkA9vK7RfAjzctZRGeKiHpehmROuAKobscBR1MO1/lL30BVg2rnZx+
AYNfLzAMXfHZBnaSczOu/9bDUSGg2AyXOulj/wMhYDzylWAkux+7fJL0rlm3ub7dbc/X42YkJBAp
+IvgPq5exPyyshSAgWzDOK/3DuCEObusWW2eP4HzU5kkxP/KOXyQLDOaBIa0zlqXeuNpMq3LPWUx
OvhT8sW7DN8uiQYQOsfaP2pzdLkwbAQ1MmPMcImB8fPCABhNtjOQfolPX1sD8bPPmS1+dMaQiM8P
17kwAonvYlxAr1ukVLjaJO0Bqv1XTTSVxenbX2NEtqRWJyMqIo3zjLl3f1frU3l9k2nDkNUkOfq3
kDJVUSlv66InzFRJl+ZBMIzgNQ/GooIJYSbLIWwfbsUuuhR25eC+dsZXUbrsx6pqsyFnSlGyuTYz
eAY8aWzFYt/eht/Y1NFDcw3hrp8sVQPeWZZhZaV3sdRpJtUbIeNBUhHTQ8sTNQsnu/gjW9hRJ87f
dhUiK8jTvfsiOrD5hmlZy0lMY+mybHzWy45WjDPrZ5ph5k6sBUqpCuERA4KHd9xaojYkeho2lv/F
A1PnLFDyxbwR+PPRqcV9JkmInt/GN0/khEzLaD97Za9tsvaOfRHrfPgPnTrI/mzVkw47JoCaUXo9
DH0ciWpzk+pnBED7gNYuqzY0vz8utUw3yifLYXbbEWsY2wCULwR/ruBhCbc4vgYQsE/OeDUi7iSp
KiXziT1wnTYMaRtM3gRvubYmlCy66KEUsMOqXI4KnTF2Hg8zm0b5WUDJoVz7/KO3yEqzbQHoee1O
p5BcC2E7N/Zfps+/fAUSTzueMAJkFPzqBfS3IVBQLats+8oEX9eMoJGXTHfvmTvHo0iy4j7FRzHU
IrSMh0ucchWaoyE890iU8mtOFvQSxFFUPXQHDLT1m8eX9RdTnzsAVKo40pxv8IVCAkBzXeqxeiMd
IdZ/9438hx1pIqj1HPrwShRBHWMMNKRScS2orC/NKsvv0lqSUfIgqjkVXKkqj/tsxtTR1PQxPEKS
zf59kxXajvvzIyAAAG3etsInC4YrjS43e3g1Wsw8iTFBVVTNTas6NMNRFUNC//djOWfyx4TT5tWw
Z2K7PssJzOyetyiEXKwlhuKFM8eV1OhqKZH7trhrhIqwn1GlZcULt6MVERjjNbsuj7e5lv4xA1HZ
qezvagNUqoR+oqjwVvOXUPjyS1sbbjZ05Zo3C0p6yCfsif9wTLLyvsd3uB3Mvq661/yg1lYQW6T5
qqwPCwmz1CnRAgwyCo1/nz92qtWlPZz1BqHroUk8aLiOiYh/poAIIqTb4teAJuaGYYBcLiTzKo/j
SnJhvnUzxWkl8X+P+q1HbPpVPyESw3CKGjp0dWnIx1TtJQ4nKOqhtlx2dCgC2G50SPPznWPwLnTi
0iq1jSPNiuAJLRHgZXc+uGmPQAMK0vNC7GiZE6rUFrnXxi/MTsiJCYa80D8jY4ZR0dC3kzPs+6qC
x3YyFydzZyfCble//55o4jP8oWoZUad1/nigH4jqvMkxB1+90UkB3Yp2W3atpANVYdqv3dPuDCx6
uw9ejz2mSFUZMjBP7fmK//JmzIdQWIw8qrE+0ZLYscgOY7i3CeTraqv3YTyuZyg0uO1sPdAj1sFx
t+xvvR7ZPnIpYhcKpyt5d6BEXE6vwwar4mImDOWHGJTWbMyc2tj1VxlxZEPCXkuhgTJ6XfEF4Qn6
EfsEZURCSM/kxGsZ19tLgJP1stY+LfLWBa90EScfjckjOZIxz9VEg0ZiwvFHSPMeR1jcJZek5Mag
KhoPw33R3bsK3plDJf5uu1X1oaHYTcZmQMsM7rNHVleLRAkOvovFTGldCQSy+KKKCvgzgYY9JWB2
jKXQ8k0jJfct8s6+cPlv8IqdmV5mAmcVrb8nD9n1o2BCgj+9oTUHvpSMjMth0fhCIHISSPwwEjfZ
1loCjMJ0ugdgFauHG+NG2hj49qstsgBj8LOXBfA7U5aGIcXD/wDtdZRhZjAqr9cDMm8M1JIRL9g2
RV/nZXoRrCxCER5lw0jy3La+7nw0m9xeAtKs+gy2ygOzsOCwDIFQ340CCvirMhypQcLGW1g3DrnP
wc+x9lwHpgTlJGU0GXbJSPDvS514FhaeRduC/HVhZSLgTKYn872OQHZKlF/i9mOEVP7RJnljXicW
9+ByzjfHr6RNhWUs1IiZbaUu6wnGW+AGoSXj2Cd+Q20F4W+aTiUK/D/fWxZtQgpMqhJD2A1npzbo
ic5ttxrQIdfJ9ospDUqy8VAX2CeP4MsYHHfvsK24w9rby+ONsXK61vtogN2Ly3IEF6nJWQEZiY2Y
qOcw5sJwwGkDPLG4UP2hZ/PyOMwdrQghZLgD240161H1s/Sfdw5Qhya9d+5Ku3ewvXrmCVkL7PGa
krtVsySs8CBrzig4jNMY0HBkuDNiS7V0yA+DCnhc+vR3S1j+FM2K5ReRuEO3jBjS1zjXp729EdZp
EUtb2+etTIcPPpYH2E0J64qCCh1cvrTHGMqDlXln4q9A0FlvbrkUVhr3BZLYpvNhjhCseXSq75j2
FVmHXmKwyAcw7/uFM8PFSWceW2mBJ80c6crnqGMVJEY84Rwpp2FLMLNOfSVGRb1KydUfrQZsLkaH
K/ffz5Fh+ESdZYZVGJcbzoc3DCrpxGIuerDhTGIkLtsUVxwo0SenaaH0WxdKTmu8Blj8GEJqazeR
nN3Gq3eevhOwp8iaxMOCqGJTfAYVWqS7AiU1TKW08xMiA2rhYDJ8i9VfzXdWpoN6sMTrrDe1sAxi
n5+r0nMcWbzBvTEKkMPCrKCdDaLJYnh4Db9at0Uuzwc+bt1+iTZqxMSRaQEZrHT8QJXLTvVx1PuH
yZw44L2uVWpj69Bmmha4aivay1jwz+5CE1XFwq5QQHlmQqdXeEntCWhn3VASxdZZMzZHuV9ZkUhk
NFMSTPSYgWDb9qxU+9qgaCgC1ygqd+NNRg99dr9Gx0Duh0Duz4Myu0qOGT0VnDnKpLnPn39Yv5RS
OHlU2dUQIgxhNfjQJ7cAmAPUjYl8e2aSec64zkFIIEeZJTydddhN3f7uzUMbuXLHRNugbdK7DyXT
DfVgK+Maw6IqTPq+4GLiSNmiqCjBzKJbPuKMSi3Qd7ZxbFVLTa06TjlQDjWQLyU4kIov01PYm2H7
zCKXEib8tsovTYkJMlQHln4OZ/SXeUiyU2hHal7P1HweMVPYiZWHp5XgX8l69NKQV0/aVaka/Nbj
lMa31djalNi8DTbujSBBvY6eB24hc5nvFrJcSahA3RDHmBs21PF5xqddEe8HmdmZ7Amqs8TtgXnG
E3Q4+8CuLDBrQa7U80nlkntwVQ6uRacCaEPx0sXFLnCyBDYNt4KoB68oGVgN6RTaFdPgmF0P6FFG
HM+FIGl7kmm51ECJNOTRlcXk1Blqc19bBIn0EkoHML2WdlbsYUVg70i4E/7r1DVhyRPJ9NLuzmUB
GLWRO/LfCv/V3AO7POu9wQd1HDVe2zzEHeAQHlEgYokNwnUMsKw/2hYOldXCJ+HHvyiOkDuKvOZ7
nqARtBK7pOx5+fDyNDvrLo9xSpTxaxkO8iRR12p1TmTEZx4qikH2wJraSaveGbGX3WAd/XECYkfD
gopf69AtMT6yWuw688Z5XlIRwnyMSUeMCN7wHkpFOCVtXoisWNtvNWSspPs8HjnoHm+VdRSzVjwY
Y0keRhwZZ1CZGNR23Zow2xjZG9G23eHuRl3/Kx+VygpmaWD58Ym5a/ralmO9rqJNRUEU8f44NRHQ
DiHpz7T/l/G+//G+VGPhl18CUk5X5/s449SI2cZTFWA+BqXSd2KEdmKKh7Ceq6PpLRfwPoEJZi8l
tIUK6ylP7J/BYNtbaRpq5J5DgiOrL4Y8eyRKwHF/RpoO1mW5/087BlW0+C1n6lnvRNes0M1hgIml
zG0rtTkqQo4xNjQJ2GsejKIZRg2hMMRyQdvLz+CzJ/7P4gQi+gLCsKelh9V7atSsAcK08Bj+1RR8
1xSOlCY5OtD1EtNBz89/vYftngjmZY90KBU/HWYst18tt6f5W5KSlEFBCTJWXKDOwruC3PTh+LPk
L+K6yHZp99D5BVSxunpHVVehYiw8olftNrbMELiysFPJzQ2mkmeY2upVwJv2XZ14+GWTaXkCv7qC
nX9v1ZxrXPGMqVBLJ4po+z4Sn7orOmBfti4mcrPqU3Qn05hY6JT6xwRqL601Dh2mtAdX0qnuM7DY
t0KJLKyEJiSW0IEHzBrgoaFqH3OyDAbKLx7xitetIu1D13Ri5tqQbUF6neHWY6XvMx5gEbLYJavY
Zfgu+sULbI4wQmHOg1aowrD1Op95+XmMFcV4PVY8CLUNW5C5VvgsesSOfQCtCe0rvw+4sk7B8NNG
pdThvPk+eQ7kn/2dphQb3EFcEQKb6xUBFJ8pvfPDvQ5pbFHNhHZWBWeITE7txljDL1W9CYcKW6Vw
TME69lVuoBuyC881vUkgRnVXK4zzr/FLbQ2JaG1EGoCC0/TtoiBX2JRiMrtWcDlWaU9WMIWB2hv9
L/dlsFMBWE2vzghUKYKnuxkQXho6N81EmR+hvF9d6FjuIq5aScNcU6WgCQof5isKiTc1kudvGoqU
EwAgIXdDbk0sW1URnuBO2ELyI12/A6tIREm1Qa592tPw4GM3/wGXR/236k0ahVwSRROubAQIAt2y
ZBxVO/SskOJguMeRo9aWkR2COtNZDFVSH5Y9sO73K2ZzCwL4SL2GBODrU20ZUdaH/0TXE1rWpyDn
UT/Z/IGTz3YpMl5CmWiCndGQXKem0jKvKNgV6iMGqoBx0XxoTj0t9VmZgaV9FN5FsPbpIndGSmAr
sFuWFLAkwoNzHe49Ts/1+T8UD0TKCYMmR8Qv4V6dDpc2sKnxfZ4Zznllimyf3lkrfsw0eSzzYWV8
sd8NcWC1QdIGpZECZ7ciFk6BGT38rnKs7rjOxRjiEexRRJIQLXoOudDZYlfae2+Y8rjlEUcmD8gT
3FBdUNxNQSBj1RsgSfbGshRH5NKm0kUywHW+mgX81mAr218RrRMmWroFtdrkaT6seDBEssD5AEe8
NcaAHN1ieajpTg1hrk6OdFwXSFkE8QmvZZO5bW93K2PioJWPHYhNFqi28WFgjyImKZeiYeF5l0/J
cm8KYovw2v/oPzZhx4hePyxnDUcCynhe/59FVqzAgw3w0zNt1PllLBLilYKzCv2Iz15S7VgVWSzL
Zqak5KiD5vZjk0G2OhGQkUNCSQ23JH0SmDq47iBxzB5997IjtjqU1P0xHkBD74q0dyY93T2ff66u
mC/Gy/3G8YZfeuS1MTFMyM1QVkswgm1m+o7XLHZnmi5I2SSspJNjuorbwih77t8PVUuL9foT+EAo
eF6OJT3nLlRsebqXRjojVXKTM558qs/rlR7kympSJmDa+888hP+NDBPYq32FuJp2gsCD/LIKaimB
myy6K22Q5esmgPIsf3kjqdONhLfM9ypRgsInFx3fweeGQ7KyeMU9/ijGTgftURazmkcxiyIjtOUD
6JKGKd8H+hCUUPoGfEsp1xa0JznlUEG32KR+4XxponnvdnOmzZKJPnZ/2cV5vD9h1QyLID94fxhF
NmFR2+n2cNdZjcg31VGIgSIfhgAGm74bmAl7+sHfoANkF5CkstblE97U9xagx6vvU5j2rtNfDaWU
GCVvljKNFeHQgER+sPZ0O7eNAdWlWEpi05Uj7cxflo9rcT8dxaG8ANABcGsP2HZvccFvl+8Av5sD
k8+KMwnCtX0h9boIFlsbg6Lq0Ji8xAtV4bwj2CDNqhbRE1UY2hrh/lpvpQhA1WZUQ71QvsHrHdls
QXefG2HftqYRymi3hgTS+vNY+CqBR4aM6yL2Zngu9za2/kTUxKnaPiFUzCCtMwE3nOY5gvkpAUKm
u5UjJnyIJ+sw+yG8aHjMuZ+3IoaBq+N1EHSuS+4WgUKFuDp/5ggoxTcl5V5g8ZtFGkfva2K5cBoc
SPIZvvIfiYsUtm7ugWBpjsZPd6FZ97F30ElPR9UbG3+QKyq2D3yiz79oS+20j2Pfz8SYpdF1EQ+x
NKmO4cfI86j3i8SfNRqbFywI/sAQOrtMvnY7ghD7I4CnjH3tZTj9XKKsfhVPyCGfsBEd/T0tmn+N
7Fg53FRPtQokG62fs64EeFwhtQcPrqX4fX38sxWQP+lXe3be4TitCaLXQxHC7WtA5MP8n0Er8KAV
1R5miaN+zM8obHcPbv8+qtl4E9q/M84Jy7CL6q4VMXILA1QLt1yqc1jyYOOIE+ECAIJY+8pHDrRr
bSt0P4o1YvLhBNyFtek9rko230Ujs7K0XX1ffJr6vdHYeGrAYQXAvPYfHv3aCyQZj6GLAyObKicb
shv6LGfgFAeHaVO1xuJzbBzbOnIF1iK/66y6GF412/j/FZutdtTLafz2ts/DifdNE3wdL0el2mhf
DkgN/nH5b5EQ35/QUrHTM4bpLUdTSoeKivRTiT7Gj4q9Eyip+dV4mCSWJmLWcdoKUQ4WvvaPHtsL
PUxk7OGxJF2OAWzLtwRjazuSeWMu5xNRSxYsuNckOru+l8xn+XSa1ugp8wMV61epnx+u9Y3RtxZn
jbAO11lo1dU1J6A+TXL9cYYNR/t4GaxYMqHJFCioOWs0UHOOrhu6zFJ9dSaaLIcforBWiyNU+iss
sIPdl0J5dqEo4S9eD10l64cfaz0VE1boqU/YW8j6CMyQ+p1m4P5sbpF07kmC0yaXSe90dj1PNG+t
o9Cvs/J8a11mveLEC+vo9qOU5jIhKbJb+LRPkJYMm3CKuKKk3KDghDd6X8zkB9j4jbSzDHlXTXSO
CEkfSexsoLB/ZBPxJ9+nhuRItYa/zKRNOiCHi5lK83JkxDyJqtLh8yj5uy78uv871alVZgDHl8pO
4QspZur/ySq1euSYsS0VF8fgoTxisQywl70er+IkRZUMDLt+DREpdoTRpPkQ8p5dPxZAy/J6FSkI
fC5PREwr/zlMeV2J2H8Is+N2IaS0wUDM8g7ynnDNagQxTxhMCZja+dnpnaTaI7f/FzX0RQ4Tu21H
RW1U3/E/yY/SDbB4hwYwU1BJowFaekYsHqSKeGCUttls+kjKPv2rXI9v9hvYkm3Cin8m11DrM35R
QU0j+q1c4bsl+xIb7U5d29VydoDm7bUX68ITjv2mcylH/mDIeDwsOLQjRPVH1YS+0EMHr/92R61P
2XL4wklxlL4Zbzgug3bdQHaCnKgJf4oG3WE34qZxxJcCdVOMp6kpWYXUEZ3Sv9USGRAmP5qr9joP
CzPTAf3hL6gofybDRr39ECVpIt96jVJwZQ2ApYqNX5FqsLyat0diNV7Lj57bsPGO8VSP1/DOx+Bc
4+XRmwLNZO+Lx5MQhq3Pgt3W8w1Lv4oe9lDXhmhYyYjfNTWTmWzdDmC/hgnLfMKH8XP1gNmnj4pg
qF8NEupxqiuTRdBQ4CSdqiDHVKH0WMNV1ANg4PUDwqS4doznyQqFQeQaB3wyaOjqMJukRLD8gBc6
wd8+r47zRhvGyl3XKj/O0Q1zupEMhgjXfwu6VEAro0YpL+JM8q6iJbTjkiHrskZ0Fv6zT+3hLKqe
KjJN1tQ/i4pH35hb1OAMYPOb9IkpQsfT0Hof94HIelsJLWnKZMNu01Nui5ieGYCDrSHFBsGkDQN4
X9J94uIYLa0+ezike5MXIHEYf95lGMfUKJFzkitYWNgiKWRnDJUYshuHlAisLTVIUpNnJWCzPlZT
dCriRizGrb+SWefG3mqdWW9Rozl0pGDBnPTyobptwBXLBxEdYzlOkb0xBuGDb93rHJVdLdXdHO5Y
pwBP4rxJ04v1MmQMWjOCOZRE4UX4LATYHHuxcYupvqfeY44UPaPGqzYWrYjko3NL2Q4gr76M0rpA
2TJxVAIa19RNIEKsMNy7QYFZQznjO8DJxf8nGpg/aT9qmHVc+9CtRn+fx6ZGadXCrMd7gM6DVpI5
EEHz24e67xYXNy1GCNq66iC1QgsE9fWMRT7LjD6/22j7HXe9b/UPNT6DfuYDCiNrvPoFoxE84kpq
2UroGb3PUPU5AvKOYuxMC3Q+K503vellN3JPm8XbAGEvqkyl6m022Y7yCmLLeySsJCrbsepOAIAf
QRKL8a5UMo2gJvIMiFezjGa5BxubPzsrLDrJiFRyj57CuRVPhuOywQ7bJQ5uDNfm50pERa6NZHPW
l8ra6S3TtJ+bomZSWqmIWNvU+GDMtZQHnLN/exYULK0GKJkNJbDmuME3i6T1vzS6wPoRPUVmlAnT
dTkitF104cszN0a37h8oje0zM3B5aEL2Uan8HLrGfEkiQ/r9BUZpbnSdUqXlEDIGAfUOeGp8H+65
/o5hPTY5A413FVED4M07mFb9f5jnyswTo+GnQAiPV5uQWEvDuovRq+DuWjCplyDRENlU4gF/QSLI
/79TCZOl1pGWqeGQlbggGI0o0TsCYSU+Pvgn4OuqdQ0wkkDW+jl+4CCzobfN94vHaWp1HnAdx4yH
knPouU6kxW1iQHGBvdAeWWPZ+8Oy54SXDcj2sYcspRZ8eV81/ypXFMnoDKnClq8fKS2mOIhMR7Cu
JQR09MjTtEfpuAcsu/TeKlKkdTRH7nwvs5srekvxT7A8pvALmDtlJVcmErD5kg/5FWewB5nq80PZ
0YxjZojX5wLXlj3vUczCoxD8GE8cQa68+VLihy2qvEL2R0WDJWrtXFpXBHlyGclqOQCGKV6oPqbh
NwSEAZXruhHw+xxxG3QI1koEeoOY9lRx3kLk0a7ODP0pvMFz/UfPO+BZWCAuTrxWMXYPIHVLs+3x
zvAMESatPUDJ7SGF23gus1fDXpDiDyiiTCDLMa3bJm3IAg1WArHf9zWxw4zu1vAF/FgdzeesprnV
nO+PijuA1Kv40KZe+EtSeMMuze++hMooyERdqhCkcS+3yHvEn+B8/A8AwgutJ3ccGHubkBKquxU7
2tHPgml0pb9U4Us22Nw2596m7JRlmFBm8kimIocLDpnv6TGLBOeTkAwdtsRN3kziuko2nbNdyOKs
7j3woql+fWywuyg/8re1qsy8qfjbzswkQIrviIEVTAM7LiEjFCDcykryLUNhbC+zx/O1qiWvKkUP
wBYGEf0DzyohJhSFjpDUx6S/+NqYPo1ya5kQgLCO0sK4CL7BzRQ1C+0vAVk5vHgsPf0JDAYPj8lA
uNUErgDUdwYAu7qM8xEiF5nkoIAsJRkxsVghnMCZs+J5XB5xAfVJ89L6zzc5HLt8M4g3nOkEQjM+
8cPuNSECsjfeR3t9ABoWFmNv4iztVWh+xPGhTpzpNJELrMiqv8EO0mn/1nZ8dGlzb+wWYR1UxZa9
N2xU9aFZDziZsM7TzM2WU/5qumYr5d+jHwKjmFSGKyHPXY26Qya0kErpvs0b3aUcIrxZFq9V9cyD
6bU0GioF3h/N7/UHpzC7Xxkpok3bxAFCDCmNdc5mQd4g1nvfuKlvcQ3+TQa/dFwqlzdcPwrae1VQ
QWY3zlBOWdVxqNxypaONJsr6s8ONHNMKspAH3krNI0knHigXezZZStAcs7Xx4+tSAG2w9nCO+7rB
8+wpEmr9vwjrydIAQ4W54fCIuTRJuNNyuL7ODC74+sf+hnRSKeaYPU2Z3WQ9nJQli1T7yFoBRSpu
okFzLhfFTowyqbXIJ6U7LB+1PmLVrzSXpiZaT4IvxPnHbT6kkvxTSAO6tr5FKNdvUGR6+V3QSu8l
UPP8uCxRhEH/6kbsT1QOg/3DdRS/uXfH5z3yakFNVRn2HXX9wv8gVLc5eqdw/Kx32h78f4b7+hnC
T1a1C+VewH87CHhCypVUyyyBMLO37RzHy05s71XsDBCw2i/itkbavRLfETyrp4KVWMVydNbH9JQP
lnP0MJ3spCKFGIP3RyHoaunWCiEmjpbAhE1mbeBxIWqCySrEnTetQ2I//hJA2T0rPeOEp0dXaQrc
LDx1R6oIjCpmubCL5NeykFI7cnNH/j9WFnq53ySZqLPWItyfWbAcHc1ivTlreRMar5ssHQYbbx6V
b6MX4iTrQ5dvWuZJkaUx7X1oKjXwhK17uNd7l7sOwSW9tgsbtQaWt5nvLk3+O5tcJQ8ZS4UI5qhl
AHCpOPGszYYmWfHivtkb+RmKtY15/YyfaOfr+z7JSFh41EcGumVYCs3/CFJaVE3n2Wx006o7Hu2j
pbUx2eVHb4vx6192Ou+X7d7H78sQCl0eJFXudkOkgMI+Dl+tY/lgTS3OeDzHnmHVo0wKGx8okIHn
6IP73FMn4g2xB+WykqcmjHzQvCP7s10rKA5KOBdcKOXlSSVJFVtjj9BrI44zvXF4/+SmlWCY68Wf
vsAHhaTYURP1FzlPQkAe1PVG+VLGeKXbLgxc71YUFKL87aToQ5rGfNbXFQ4C8ByIiQCLafYLu9AW
xbZurDt/JVDOdRQ8eYSTcUCGv+VoqjsSKwLOKE++UirTzd80D2/cHPvz0uEGA+48As8XS48YTbdQ
q5RBWjX7q/TA2b0f23yC3LAvUQW3VsmMxf1pbB0y6zHvcniU1qcj/ncuhOLYGSFbR0l8XnBziBFA
T/4GSCMyV5feuZzeY8NYESYnzirFp9Lz1BFsevh3TYjjBpJG2mp3/GejH/78RpYJduOLwxr/6Hqt
JDB/3diowU+BvJoCQEYIyjzmUUOH1776wKweoKGVZYhRHvwo5fpeM233d37kViwQWxN2y6OL0TwG
ixjuqerqsLdsP3M7hWbNw7hr0MsnzaxmcQ+m09N49R+qH3SY5vtSsX9LFKw2Wdz/1XaCpJXKI/xW
m217vGICnNJiHCJ14qi2M+F78tHGLp/qra959rZJEbaOMfvRBTOEYrF5sJvrD85xBpkJBia1bscE
mHucjjq92phVzpVCC/9BwNVVKPrkaHQ64vDDx1IKFTvv7VROzjpVofDqThs6ex5+hSu/AC5yOcnA
2NW+UBVtPI+mEieBQKR6VjbHhHzWN7caVxuMg8VSf4T7Y+vjB+yAskuFy8kb00zf4SOSQpiQKxqF
1lgbuGvJU8aavhWslHlEdy/fn6YfK382pEslbcAix7CF+uvFXCJNUpYxG3rr4E7E3MP3r/ycVXeZ
RMChYu7zqhXtTTwS3/kO/IjSqrDqYXNF3BZSj9kdmNXMD3MDYtyxkrYHAJZ0sjRlm/2OCHNY8zcR
ZK6XcDTsIaYvhSgIaCJQQaDZ2wVuYBVNrpivmMq77IO4XjcaymoySgx0WwBNFXCy59ZgyydFG5oo
keSHVckyRPS2arB/wtleeiOOlMMT6A+4KyrY86qwOWQ1KJiwDj7mFJONMmq5G08IUlVErZt4fmzQ
jpkVpcNSTVhY3f4XKvKnVlwTJQm0NGYWiThkdfdfQbnf7h0ydZ/ntv3uxzZXPy5YChWZGlvmjoeR
s2E1OwlcfwSJp5el3g4jA2xXwO8yL239a5BdXKbxDAcmycY81h14/7bpSniFUQ/LKoz7VgGGxW5e
BHgLj9mGLAB3GP22NeFH7z6mdDKb9ZM0KFQnecVKPPcl0LgOGH//HUOVIAj7JGu4++kT6VxlqUdN
kq/Fzpf8wHAMXwMiyJYK9V87DVUqpW+DyBTZq98Us4Pw2GqhLgq3LUydU4216jl9GzB/dpSVL0V2
l909ni6RapvBmNKgSZDSccrRlADmHlbrqOez/O11cr3QISTn1PN6jWrBRPWjhEepqTFQmmio9tpp
rXndQrWSV6YalaRPzYfslgPZwTVp9muIj6mtCccv+ibrhTHF8Rs6eL1SS5kTTbzqFfDVWAm3/qJE
C1kxOv7Dt6MBwibO3uIoxihfk447/XdO60bioNCNCOANh/EgnSAApOIBvj51mGmTA5sbC8fcAMrf
0VWgdvV82YN9rhb3RexFta8sXg65Hta/ZnlarEdRAivI9gpKGEa40+DoailoDnaZhj8p1heJ840l
DrWYnqOkvQxqF2zl9vmAdEKNeDDfjoAb8Sr48epB4UAGJJIZH8+/AuPv9QvPHZLPEhekL9eSNDWD
hTD5JlZzQ/a7sPJ2Drs0H3JIegNAZFAMsEwlcJf/pCovbZIofF5w7BSLwGExKPGoBunts05XPALg
rgaiieErP8lUbZm/5ybjDZv/CMT+BuzMXStWLhO/6tGKIo5+GUWdKg/hOpGJLWk4JG1JaYyB2Al+
uEwcLJ34uQHYF/AOpWA3kssMiTP5NhJP/mAFLhsKty9d+fIlSfzphEURJeeZkJQq3lv2IbYEDqc/
NAf9XcKjJI9MRrPEdEZzoNW93O5dgznC2/chIAgGtWvKu2MN8u9fGlVKdR76M6qBi+SrKlrIu/dR
jc1HpPBIdJz6AHfOb5kAaUs3UMujhobjD1+Wyqv251001akdpimyB2xis8X4Tm7j0InDiV9St05+
MDG4y6aOXSlqvCTyK9O7rhUJRUGkUHoaCctm6Mqe+oKKXOKXluIxcm9dQDPNHXaymV1BfOmjMrkg
5s4YKqmYz6Tb+CDhShaSyTcEXDc4q0tV/+MJrE/P3m1DTgM30xxaH6QoAgm5yDZkNbqpvX2tSkxL
CuLxQUHFWTIMyqSyAK33dfGCzO6T/uJw6oDPX5LXs+6PBso85rJVKlCIsniT0un4S0zWIsINvqYh
MFjhTUBI8Qi9eSEYXBmHeGys6JLvnMQZosTQA6Ua01gBmcJXkAjUGEZfJ1E2mRVzwxHSkKvYddJz
YUQxODTNZNK6sd48rYY850uv9CmdlxM6lm3GIcRg5jpAo2pKmcokfTMTj2A8wi62+dZO1cyxdHC8
Y6yElE1oE1dbgRJv2jOAjFGU9FHHtTyquNzzJoLAbswh4gSzjIuTcgXMujHsfHBeBSxtxn4Hgq/5
M1bQlc6q9w+2fzIhIkwcbQ8Ij90s6/LmOxu3WFw75bwheT8FRgfOUDIKsJiPmdgb4yHzFchJ7ZUb
bTVKUpnesKCQQTGkwFcjychUiscD+rOVrEono7+HRS/tjcHX7pYdneJT9tI7xdR6xopVpSPn90zH
PkmiUnsQ/5+VpzLp9iIrFPvvZNCdB44R92Zw17e5uN4/luNgncTLxJ4YWzYlGl9QqE3OyAkhcYAs
qoJB+x4VKWWLdwKnkioG7r/1JTTT7JQuBBF4VY4Bt4AyoZ1Yqy9akhoUGg4TF9cazBwsfYCdxR8m
bnljrsesfVtdQZbPJkKFYwR5GBWGma2HfQP9TdSA7VTWsf/SGDaIQTiPK2z/xiL367ju9v75ViJh
Z9ZLXXVfvx+BexhDZ76/+hLA+RZy271vMI1Zf50IIWRBNOzBuC+n2EVdrV9D4Zn+JDPucbGSXt/L
Yn6O1MhBwGaz/WROo3y76Ue04lTAQ6CCgoqy5AjUyoyiiDBXKsUMk9KxzypPp2SEoGjGTE1P9vkZ
MAkakYBOTm+/688kNHlu+6jB2PmTHQbVKDOJ4cts6A6Tt3dqjREA7ITWZjkAlsGOaVmE4WuhtcTF
kWzlpG++jWpJ/3nL/UBbs4FqnjX3/K2tcydoNDCQnDceoDMRsVlzqy5WRl2XQhYEmckFpdWbiU0S
GD19fNU47xaYwl+VBdWCLFY2KTB8U7CmN81PO1uyE/uW455wq1HrxzYlKd/ZCwKc691ufxgK5TSE
k0n/xVeKx/bqCLPhLuO19JmIwI7hT5+eKrhT5/pfIqFmBiaxr8ZEqpcMHBKVkt2lqH2W0zQZm4A4
SJuYiNiQW/UaTBHUQKprHrgjYEvChiYIYav+Qq0luj0CR1N61eiwVhKKQ2BY2ZX+eCZTjYOROo/j
0slEQDCwF+oLErf8BuCjxitIwG06QidQKL4c82RlEcoMfc8v/G5/T9AWh3cfvpokuGBRljCl1Sqb
ZBeYEEo0z9A2JUQSiZtwLbnvKyhrLf45wNOOp1weSMusS4qtBbhlpqvAcEEODsr7kmuiNkjtiu94
HRILUguvF2kGAlpJvxn9+fH5q11Ig7nRT/FjkxcbSjTRvTJP3voV9LO/kkWckauKNPv0KnlJNo/2
3vmd8AuHcHQDrAwpGOubO7r3WFJod4CBdg3cxK9R569jmzb6YR5x3ADRYlNJ3+xN93g1aQ84bHKW
U0A9/OUVLD+O127rKyd0uzJs2+2nHd7s2F5+FXbucqkSJe9456+8zOVkPVFEPZgFSIC/Ul4CqiOQ
XG+2FVHENkbTN5TWtq86g4EWRN55E+XBu/wwY4ycspdVxUgnsGg4K4ykFEptnqmxWEmTrcdHg80u
HX6Vr3dYAjhNgyClA0FHvstBBvH8A35MjwKcQL61uDH9E/PCHEDlhzFJojYcV6VGs81qbiPgQpOs
vN2Cv1r5GNCg+HKCReJBNeyKrjb/32HpaUzFybRvjlTyFKo2CJ33lkEnJ9hgi9PYNNYLe/3xOsKh
+lGby7K1AzU8qqD0FVYJeivtSIwriT1ldkzQlLnLsja3dWmM+KNnO24M0NxDUb0+rr0O6Hlzff95
3uz91px3jgD2IBM1ccCyxmDcrH/u+yGEfBDD8jt46azW4K5AKSKemInz7SDYLItXCe8n/j1YObz9
dbTdpj0TMnACCgoGzgMn+wnp09GoJSMv6Tc0YgTgGh51AAqDnVnKQomfdOSxHGUbBtLa/VPtc6rj
M2rR3JMkVLJTu8uVUx1BbRey5RiV6p1Yjvb6EU473ydg3AXzKS6tUH+zxvdOjUnkhVdsFjHHCvIO
4U0eIlcY337FQwEeHBE1V5NhWPaUurpvqHkOojsv9sdORDZ/QJxPLq9BLb3AsM4PFpQFqu4arMZJ
m+VUfDqcm2qG6lI6rxj9rxzG+7cRToB3e7T/4taZ6/zasgqpIFWqMctf7hglVzcFvr6BspO3cN8G
nZVzu7AM1KuIZRF5G1i9UmNGaEMWIXYgTwNwgyyKvzCENoswoCaiWzgLx/03XxZu+Jufew8d9Oq4
nkBNNHq5I0iaYa158WJbIHhrcxSSkdgYHyRuGJLyk/bw0b+UeRrdS8SAWEl8lL3c1lx3/TI/QuxW
PtTb5qSzhAxnjvWGVBobqMsyGWyEZG1bfwC15XqgpjKOHwadrbTXSbxuvy2CD6BOY0yoBfMuUSeY
Kq40KtwBe8Dq4iGzIQRH7SmQ1WQUEWC9IzQZ5VqR4sYgxOSo031QJ8ZervNqLg1b1Vhu1XofU8Ol
Mh/ETO/DC44TnP+hO5Uph7BJiso3MoBnKhxiCXAjjljmFFPFl1q/4x/L/90nSODpRR9zGY3wZ84m
EzWupP+YniVeLfBz3j/64jO2Spba45B1bQZfD9/Yk6zJYSUMczRnE/ocvWGFuoMz442NZJH/c/55
3FirfoCowcnDYkQDpB38QU7zgv8RSsHG3FYuOu0qmjBS1FHtP+UB8pMkFn5YSgK0MwnnO9dYeHyj
IrpV6kahJL7ahKWDRx+vilUh+Lbv3gnI0OVXloPvkfv4A+3ENEQekcx1Jkl7Oh/9vVqoZmyZR3qG
+YOPvGqpegcEQklC2XMP2XugkKaChyzy21jdYXM8SWntpAkyNmCm26fU1I2Q06spckRgsbQoJmdd
QCe/dNhYkkDDht9JZYkpvE9IjQXaJIxvGU635KsESJjXYEoZ3QZ/jmITYd6JI7jOeEQeRAEWNVuZ
/A9/gQbDaMeWY8Q5R6+sIxL56q6iI7sVyuvVVDRIk9B0Z3XLeCO8SKNbFAP/O3ixWP8AqRVdkU8t
NidU9Ro992+Jq1723PfEDDs8uJC/YOC0Sp/hZIycjWQR3pmVtSwTu/+jwTJ1iQHy/yrOi+9gIHJ3
l7WxiQH+E6VDpf27SKEDbhv2tlwbjcKikboblwI7m9rDLbjxbad0m71UXSXWFUt/n+KiWI62sPKA
mxpYoYlUEx0VyJVgDcKSxEEdI6rURRQ5EnSxb+weFSyubadk8PwRChK239l5E7YBZcSfxNeWHy5o
azwKAcbvIMzmVdTXW+4rYGAIjte4JytzMw+MWKyecD9xEidjgatie8LPGa2CjnPt7WS8QRxdiEum
yxqk6U+4PWilHFYcXCYAbLOnC7tjOoUXsjeStnbnWsIGRwenhivga9X4GQCrHrX5/2j8a4D1ICuw
k7fdLUvi1CXddGOa6sD0dJSsmANRvwY69F67kJPASDVdx4rU1T1tU1V+GlH369BBR7GlvKo+1FJf
mzGEQ/j2vX9SvhKULPR+bczjHpv14aYV+BzBWoFhf2877zi/7HxV2vTaPms+EOth0RPCBMf+vlm+
2xc97Bk985mJhVCwpWugnO2LvUeZUtN1xmKF7QepmfRQdK7vh4BBRFBf+EX9BT/AG7U4Pf8CaYPl
O242ra1o//CNwoY/VI8E2QuqLV1jAvCyVGiKD3PSGedayxG4nIPJv+kgZcHbNZu8uxBM2Kt+JKPG
txTMQdAJlXGwv5X2iBV77Xv8PUiflKXBt/4Yq47tBXmYe2D5iFy+Yjb/IypCwUtn4JqWb2sWJn/o
zqLxfjHJrBaTF++ZYbzAXck/S2stElYMYdEiQwmCiyc7chM3LP49U/cJfRSzODIfQptzVH6+PJic
3lzNBT7aV6Ru87tscoKK30J1gFbzk8wcEiKtQUnk7WRx5I83v85tpiWXmQjrRUtVkm8subiQy5aj
7sE74yV4k7uDLi+c58yIfqJMzJ5dLyCMchoaIu4G774sTaa7buCyrBzLzDXcdiPaxOnsREJT65NW
NZZf0rEL08sChFVgLGN+wNtHQf6n4jn9BZBwR6qurL29WBv0Tie0qDw8y5ZEPbP+iZdCSqijZyr4
t1HgCBY5LpRRlHRgV+wjEqwXvnn+q3NpwVMfo6/fGqMHEdfJ7yFaP89w0HvrpTGV8eWtMxTp75zo
iI14BaU/YI8de6/z4wcMFf80Bj1Rj5FUi6cKzpI9J2Cp5CAqsNcwV9N+HNNWlt1iGOmfnAROVd7P
r9fnKdgKRc18JrGz77oJZ/0yRFSdJgTXVAsHQAnSr0H2UyjR9NkzWeAGVx0o8n2Sg+5HRhMEYfm9
Env1fQA03YvKURKifbssWVqtymaUu6J8P2VXBu3gpbIa5wI1WEcnVJu8+q85gAoBnsvDXc+rU6fE
KS0bh8ER8ZUOlIdO0XTkJP+/TH5ds7JufZGXjThXFWld+LjG4ovMIeqc7YmOkorb8S0Xhip96Sdx
QjUF1hvlepdO5PZh2VQID3QYaQFZPdd/thhLJremTWtgMfUfL9W8TeYIZs79OzWIkPsV2amTbNBi
NIagNmf2K3/WGEZDaxaqT1Dftt7PLD25KReWYPbrPhAWOGoDrZjQe1puySapi1aRVJO5V47fykXF
tuaBLi7SuyGNa2bUsV4rzKzF7jqLDLpY0bYaUEyID/AAC/+WTe6Fz68G2wo9wFflb5SWSAT0Snia
lXpW2ZJFGf+Vb2HYPuua53V34ZPHwlEJuppKaIx+XtaIVph3gP9+yRJ43S079aT/iTqotGOzkz2n
UAnsmlqMYObcw7SJsVnMOWDF/2aIPAKMuW5+WsET4QcFdJ16zueeGn4c53O0h5IoeLeL9aUYZI/T
XALvUn9fK/OlYZb1Kglv03lCGpOLmzXig0q4ur/mo3fZtpHnt12IvJFfEtS8uwfbMd0KVlIq+/5p
7I7dCNie8DGXpy1gaLkvuIDkP4xMVp6jku5MWu/LvZEuOwcZ0kbDigIvrkTQXLMzF8/m25ptLPWG
ewSbGJ3vIhWEqROvAsAJuTRRaxWYz8BoB+Lm/c/Pkze4AUT18y1cWphgEXngWpOXA7jIWtxlS9+B
kuj2j+MeTYtDyIwNzwjvFM9fvNeB4lzotG0Wazdup9EeLkJqn/IV2mOui0izNY5wqkMtJ6ZK1yIT
TzmlYxSw2pPqIZetKKUqJ0BprIL7VA3O69jZmPwsrQMuLChdVScvvxbsZ7SpDcAg/beSOy1D2fq3
uGrJ6R7liHrrPRRa4iw1GS+QOG16aEaApoWCb/iZDCHGxUfENb0Lm0hYvvZivlDtTaFUpBgUavDe
Fl8cWmeQEs7A1ZlEGeSOYfk78kp+H1Q0LqskvWqjvg8o86Y3Kzhx7ok7tzGMnUBfYtsZSVjklHgF
5v3EpwwhPUXfDFrAoK3XaI+zkstbH3Rs/TlclaG56ak6j/Uhzrh3nElqzYUaTjUpk+vjd2KIs3UO
NtrAy8hZO6FAfyE9phrwmBHaMltixAJgTtc5Fqxf1CvNvCZ8KjhlQ9uZmhiBnRLUdVTDk3zlCrEQ
YCR23AE40/Os7LslNIkMUHjZ8mRSmPUGfeTXWazkgIVoBbpTprfEmpC0k4VkjMcn/12TAactlwFb
qJEpQGIvzY2I5YAGHURv/v20S433NJIAd7nWRlxY+szRoTHYUSLjGZsQMyYA95V8xz6gkFNk4zpA
518N/0Q+bMDhYtjulS+3SncbvlHCer/VDlafiWBeMBryN0VTLPdkZfHxkV9DDYZwnocPWGIxvurD
xKauF8hlqkSoXDitxAqL/Rd7JMaVpVtthnTJQjcJ1qqKeYieOqoRS5q1/3mCLZSSdTSCnS9fV+Vt
4mcc/OMN2WwKPD31WuT6ZculgQsX7fbOD3NP7lFZXuJByWR7z6AZHIvJ4HWlALzYZ+0+ByXfKLl5
RLih7KOhJBW/aB2dHlTL+7WjBiTM80U3Ox4Aia9wuILC+eDETrnCfnE+m5oUIYfBmVs2pcm/fd8n
gS4CDuMOuoHgSYq0NkFaTOUP6aaRAlbozCLX6QYJr0PTP0KW/jjdtjsGNF0yOWpb6soGzAmvd/5o
cii/4zTTX4j/bC0ikJt1ho/e2EkSa/2doU3KqzdI7nMQBE8NQk677P0bN2RqT/BH7mCDngubnbbj
AC2cQxs1pdXiK2AoMlLT5Gz9w6+wsCGANTSlsu8lHcneXgDtLEiAWZ6zk8o5tDc0C7+IrSem0bjq
uFSviPuEtrsQYSuOgLlQ8QofawfsL4eS4MGlhLECmTnF+ts6IOUlb6vCsJG/eMaluaNjHCig0b/8
9NjAjYrX306nWP5WmFyvmC07rYMUEETKIS3YKdjTNqhOXAkvI7VLGTQuZ1Fy6CcTrFeCyzYetsm8
wI2k3iu6tAT/Z7rTa3ZdFjwqfiBFqZUYqNWzTKKjHE8FyRD169bsw1iNp3wilFpk/Lln2h/nXmxH
7ZLUrCE4X7BwaWKQpkdg/tTA1nrE1ffEk6zqi+W6iWiSRqctl97JpSwIkXEb98HbQfX3z+q9i2Hp
plc1WaYgQIT3UMT7TCL46t8hBtSSQ+FR1UfoB2cMEsCkT8gQ5gtp3zqffgiH+y15EHBslwDWh0Ex
YF/F1z793UBEpEp/6rP/H6Cdv2vQyKa73PMg9TaRJrmWOcZj9wNbkj45OJLiTZ/9DsSL8Ol0UtKw
0B7+15brl79TxZFwSlsD+YJuSUt4XYECpg85II7lHGjCi+xWwheySHd7l3GKmV/HQQykj+Ev4NaC
hxjKfKmotGUd6NATh3eQR4Swt5D6OiuWMzXO0P6gg1EyBRHVE7NgxodLzsPwedJtihdUhKPXi55A
kAUuD9qkqCr1a+p3wdg4M3BUXDAd34RKTAJn1z8bNHgn7mayIxAhqAI15k8D6GHPnH5sbhrv2Kk1
rUDpRDd6RYR/+iey54ryOmBXS3zKZtrwjFHtR35eJx1IeKhdFcWX2TzLUz596kqo5+mkEOktj4JZ
OQY1DzukzWbF+nLQKLhJfrjJXFGNzwHrpWHSOT1+6nSntCPKveboube2C6kw7OL+ALSZ0WUcSMy+
Jg0J6S/2bop1Mv+R5CmeVRUhirj5T96h1Vpzt/jm9NeDBLfhiwYOHo0KOTwxwBF1RW2XSR5rXmC9
GhYai9VVYEN7261NBxhneLnh3BdiN9WfOqtiw3nfBMwP/YL+LU3R3AMJHm7/k4c63212JcQiLmC7
eN27V/mg3+I82nUCYA9MQxmm3GkpFYyemgCqe0k7Os60QkLrN8YlcvMOjn0b+xNbePHfTb7v5JPp
hWMZZMRGwv7UmgJllJJ8BO0XPL1ROsD3N5yvEygZqHdvsfcjtjjr9yjJN8FOyH5ZZA5DrKCtHm3n
aeT/rweNnAOYN8+BwVrTJl2FRMhhmdNDROtXqpGiBuVWC+k7BLwcOxZa1CC81JtjZ1AALZ1/A1sv
HLWdlXDMful4sqhXBH9R4Z4kAr3mTv3z7R4E5LqeM10fwFZC48FeZyCpoIWuMZrMg8FaaE9VmYtU
SDeIKJKvz/MIAYc9PvcTmRlY54HGC7p3vlFHrnwPQGSCZctaImpcQZkHMIdr6hRoCtG6wu6ptWkc
26SdriKSfWJXF6zvJyMY8HXSWp/OzsaKSSYsmR+bjE+TeeJQP+yoS0FMvgioCnnh0YoHpRIwXmhD
AbiA32nMSNXKtfwOx9oG9S1dYa7SWkufrg2xETRhLwjmX/RVfqleclM9Xf7ultHzcl+fp8UcEIpj
Hdmf37UwfquiM1iWA2buq2WeA9fnSX3EF3BhdcmxA2bYlJafn7VHC+UaSnhhKCZJMrHtu6nGQMNy
ecwII3+IvFn8NM1lMf9fvlcj+PFp1mAh3YFN4VhPQUbTnObxyEfMbCZ0ZYgegISsFb60mOk0z4MY
pmLvORgyjaDd0lTMKtXOAp1K6ZLPA8YnOfk2XIh9puAre0FJv9Y9z0DcJyPoY5QwBTt9a/33qpNy
DKj3Nr2dAJ/BEIqn5X4GH3yMROG10/5eoONrM/PqKLT5of9ZYBKajhfWS6sKkRbhyLrm5qNhpiNF
oeU+gnur+EyEMC0tSW4dg3vo3FPfa2t98OunP9MxoegEp1Df3nXxG0h83NF6xgB0e5hfj8hZ2QnT
4NbVuDaaS/Bv8E1mIV4CEB0TTg3MkuTVuOmuySYDLwRR9wiKpUI8a8Bs2o06o7dAupTIU9q6Gy5M
ucOtO8wp+olpy56fsjktaT0Cic7Rf1baf03fmP9QkqUXCBZ6Inp5ou2k+NSE695MdmC5dLLOKuiL
CFqHpreKdpD5PQHhpKKJugs+fKp+FkO9QMdGNw+QyTZZJMmYP7+RT+a0cD+MjkWeiP8QQuLI5L1/
yhMPRWU4KCY5JPJB6kRacVUFjzbooHytiE7QMaHw0P5PTc1Jwh+GMLRhDluV7F9zs8r0oaylPP4n
dwldzoWeVkRqJRp5nZkcPuCy9FDjhDUvDBz114JJExqNzRNEuPj92a+KlTKg3ieSDGvKNqrwCQvW
eUBWUwCH3ayVyRp/2S/I+fe4WSr4L0Lq7QJtipnIb4NkavSu1TgxPI20uSu2Drf6rbkFMiZzVI5v
ybm5Ft5xvkFKqeQY49d4pscANMpKEeLSWlcKbc47OMy/twnehHImOOmZS7j/1LFDpaXtqlFLfzpx
dNFTnhg7u4RRSvZNuOwnvoAwVtnzdPRVo4Q9SX1h2D7HPC4l5FjFqGwneTH36wDTzmwTxxkLaeRw
OaZAPHn9RTEvLur7PqEn+pDFb54yFIyRUb/0Sgpin0uAiwfRd5FlOaFXG86bWHeGNEKiXPfU4h4R
b5b7LQtwQKg4c4F767XcZpzqW4gBkpBn+yzwwd4s2WiVUkT+6ZqNa6lw3yAGD+iUKcVOzglwAXS/
xwYgI+bMZ7aoTxxKOBDuxuo3QOJoYjtpvTgxqkVTe/nlq70WBTGnPpyKbG5ucm+zOaCWrYpTPFtK
iv0QNVu377qMq3/mrGlLim7qK3vthxP1wwllWKHzzS3pisLrwNKJp5AFelB9RYzwx0Q5+24/MQSF
jow7SupPebiw+1bKyj7jwW3VXz8FGmE+h3rR7IjZ+5FbsRqraGs0K955SN8DYIT6n36JU/jb2e3i
Iauf5sk7rQWtePuw9pdxiIFxWlW8dQF6qRIxdP5xsqOQiQ41SMVuWwQAQT+Sl5gvfIiczSrNvaw8
DzsA/WYZSmzbAJFapCbRajIIVfBpZ9mQ9zzvPafIDOEZLuoKXvAl+wBN7YUEY6GJyT4S9T+3F+Xl
owQp6pLG61cF/tghgBcp9DsTNdCV+IXfQHR6FDbaMIaL79kFHM6MZZqr4qv50G2L8fGeUMpYjQ3i
3yaW/SR1kM5YAC2PrjN3MQOUmde8jZKeuLCb0fK6QtZujsUPII/10KBOecJPUqXptct0KEAjTFf3
foGm4RDEmwFgF5VRZpQVyf1X8sMMXmUnOvvSMhKi9Yf2SVlpH6tGvBKCoTepZyYyJdzkALQrIxR5
hHt46UvGvSW4+aKX8uw2vhW0OxeeoMFZJfM9t9bs88y3SxZrXFx0/Wmw6jpGWgxs+nOk9wqOFrW8
PpHI87MDt+zsRaK+hpxubYzN5y7Sfap0QC6poeubqsD1gyOUEShT1HCQlkML9ZDGEaPccdTOjdTc
be/n1vgtNEo472FThJVkgUCbhBvVDZ0bXKCx1jmsLa3oVjNXJVEPjHNIkaxxL4XtbDtD7BXHudQC
5pJ0tEIb2g4laSns0MoVSvQwy4xTdR1npusDuyeUUiz2c6v5eHdaFwrydThHaVRu5pkjfbV4jBL7
7AZccZR3SAMmqB76jYCkxjR+2kr0nzblq1n02BSfE1uVa5V9CTobNZNWhNueZXlKyRd5mYn94/Ad
eTUoK1FsqszNWKMqDByeEkNe5wpLTf6ALBYcKdF5krNgARgFQx0Sx7th+51QXWfDt5+K0VVlyUta
41LGC9LzGjvGK+V5oOJJ/fjXi2evmgJlQTNwFR0zcS+RReUGii4nUgnso/sVeWmdnh3w9o7wUHDo
GaO4fqvx5mUCQckxcrNyCwRJgN+0m+cx0WPspKOKCExZl8h2ffNnHVxBUCaNr+SWCHfC8gqbb05L
3ORjKNpRV4XvwqxBSexapL/3t8yUvajkycCnP1DLtd2ECsoIDjThqCors0uWBSnV8ixurmJO1KDP
DwFokiVjbVOkgZmjIrOn2lL870PsPoEAeobPBaWwyMV52e/bgLmUF5+aNlBks5Wn96GoKlRleeSg
HKRKLQpHqcXAnM3wOqPHBcrSnDwieLf49a6Y/4RfquOA2AqgtlZBC6dNAG+bluncQhZ2Lvlaiyez
pTzqZApicB0WB9JnUNDJPBKdxxChYFyfKxjb98aqmzVruMSk4QlbErSYGTuU8AOr7AZX0g1UCQ/M
1CAzDj/4k3HviCB69ArQz0SVoI+zFaOZdWAFSeP1T1WnFXgyMVyq8esAy407qiHK2tRhg32a71uw
8+eByIMVZTGdLv7ssxeiRz71sn7CndZDKvs3y/fqrv1jNxUAMhsmg5D/Z7Xrg77fW3HNULLUgaUK
aqeKTfjKY1cbNG8zLUX3Rp8mbLy0dVdIgjoHts1j7YVWBlr7m4Rs8ZheuDV615tBE+cIHGBILDSc
vWGMR4WI5VnVTlVyIIJWuc6mOurtmcwlfGi3K8FpSWYeypgA/3enfuehQ1TdQ4hkVwfH2wxuAD7x
vZ/XH6DlICz8oto87dkF9/tpWJD8310maf7ctFIk1sJ9lFOnRfKfLFbwGyLmXkDcvWJ65ay5xn0v
gIKSyKUbB6lTG0/SKVobLiwAoAIVYy754rGe7TVexDmbWE0Yf6jL1tLsc8epIF9MBmmnt1zCgSzq
KHHALk6XV9SvDnkjrhZ5h05Bp71y4dCjGJQvmclf4XyrMWRsHf34CivT2f7aHnPTafnIhkci5uzW
8Q5jIYCaUjWFHt/XW7egXqVR7siZ5Wc9flNnfXZNUP3OkaVULw6/zuTZnXE4g/2msLGD/K9DWe8l
0Cb/r+LAw1ZCBBd+0H4tM28knzQnWkQdlLTIOxuRp7nYSz+gIL4VeCKQHwcn8IQO6/iJ8+Lc6DC3
xJfAfxiv+B6/1OMTe2kHsPtUBCyXhvtNAE6nS9UDCdDc4tfJebW1hnPL//5P4Ur4Gp0goLO7pst5
10jACR2W+L7+cNKnBx830SStJ4Ce1ggigw95Ecse/h9eE2mwG6wYoMa3o7pyWwKO4vug1G+y485w
V8j1wKOGTFrUbFS5WMpLT+CvO1cM72qSm8KoTo/VZNGmKW3hWY+eJzKLh6vqr6yUF5eNAdeOkYDk
Bzge/AAZMIN5Sq2EGCN473j67pg3toAGYwWuJCokFF1CMiOZCaprBdVS1q2JnekJzxN1pIndgYQT
7Mo2QBNohUllM0TGMNkMbLAsoQl9WDLV56Pebwv7xs1wbbnJxmWUBi1PMVlW6o9JWUtAkF6mEV/A
mb1SLQmt1XJssQFJ8/uTfmfqAWe7ZaJu3AV1nNFAeLltZq/7TdsP9cx1BupR+C9kq9uFS2vUhGIb
seIF2DlS5sQ1qOlJDQ/OS4FUruWjhW9VbJDZFUFzZDQl+rjDU7P7963og8qHniOG2S91LTIS/2P/
tEB3DBbhYK7BvbwY1xLCEANXupbmLTdbZcwU97G+1jTI8f7Lj1b2X/y/EOO9NCtjLfyLb8SUQKzO
kH6VbacniVKNaZVBP8Ict88L50nvQDO0i5fES/uaVbVSa5TfUkI/9d6v1TTGGxBZo0X/g93QwN8U
OpmEi+hULOWDaESGq8AbGYGK+qxEkiq3zGKB3VdvOiWe05FsdAw7jKSyu+YNsW43YJCntJrmFoDt
UvHdtUAN1EdNwWpZg+Lckc/gwmPeAUz6jgAsdj6sb227ddbkqC+BY1LaB2as5dzooaALLWhG9BQt
uqGVHHMsosTiVuj9HrhobEOMcHRoCk8DACSq6mBW+t8bOeRGLhHEWhyUBrAgTbRVIpmQSADgrOVd
FsUBfY2XdQ8KI5ax9/Enbxk02iXUMKQwHGZwxguuVIxb/K3cEJHeN8HoTTpAJyeU7iZl4lr7W3Ws
g3hGshhdkndGPnhbL3Ix7/CMxgEU+q8W6RjZ1BmMZoqfMn98V5Qi4fgNDQV+9RNYD6c45d8neCHi
1yDi02e50RqBOWyVamZmTp38t+ZlZKwL6e+qWgtS73nXUdFMH1GieL35k+NR52JMaUjMgY3/GaHq
bUHipAv6dPOMKRd06a4WnWYJLfpk+JxfZ5wHeKzEmwKYaHV9yxFBvNc61gU3H6tWNHBkoEW9g+Tq
0Zs1msIXwk1SqHBnOl07euzLjetlPbEo95KZ6PDCdMtnkErKKgmdm1sp43FO6eSorUeJGyZ1egVq
FUxzEYCP7k1JdIPSMMqsoJXwG9+sAJMAibwTZcdSAWqBBtKvkjLbrs7cNBDklCDWabyTZZWgSN73
b+jTBL3edU6KghaL0vs8WmZfQ3z2J4QdbdumUkImlXoZslURong2LeBl7kyqpM2Uqo2oiUwdz7Zm
HFQhCteFRjmVA8EGKPyeUEkwSTcomGp8g7RP+PvZ0iPUl231B2A8+biNCUb0fM4oImPUk/E5P+bY
v3/LJ4vcAcKEUfexrNYl+EmXccpBm5gUbhslDvy5qwsuWzyLGl8Y2wKXwIpJJ7RRfLCSYHTK1ZBR
9O/vxa6YoplqqDvyLwW4Kk54aheeEHYrfWj+IFTbxVBFRMbTM6aG/fjDbFKKT5OAOFg3unnRl6RW
3xISr/35gWietsSQkbyMpME15cN6yoDSoPTkleilZN97Le/UYiJNPzuCVikT7dwQ2siuJL0qVchB
OHRyjBOPPCT2T5cdrsydUOVS0WTIlI/HdiKzknvpEqM49unBmNf7I8xWs+uc2o1CRioRUtRWaXIC
4cG+YO5ruoteCFrQsq5BSMTP+Bfk9tzAhRv6yCLwFecGl1FUmVGgDo/WkDQnfwBeDBAsvd5rWWV8
wglmkCwkmpYyQQzkKXUtyVUMwgvY3A6AtBRTt9mKcOcLtfkGNEHwRR5acaeaHuh/NCL1Sl2r1AKJ
aCHinPph+H8WXqt5/JdvR+E9Rh++R/7Fxt9euU1rNofb/2viQhfWcC1sI9Thu4vBUtCEmPhnuO4W
RW3f13Dex0/lo76WYhXmmNzxfMg1tH1eDvJ9Iw4RDb9HH0Bz4yM1M+G0B7FNqPMpe/QCRsViP71w
/cZnsihkBFpfqZjh9DBDGrZCc/PFadIZF0WLGj/DqfyKN/utEM+y07iEf8Li/Lfbu5MLh4PWpVTC
kxHOb9NBvEQKKPXrd7q8AXSZVjO59rMT6kDchdVLY1rXqoxdHftbab2agY5y+kBQQJoV76xsqFlL
wv6jy0Lhm7L+vn/GS0KDWfylwfTMn3IcxGUMPxvOVRIJ3oNe6NHvtygJOOzLUpps6SrrGc16ecfT
kIku3unkreoTv8FyZ+TzxLo4tUxv9L/hoJaDCWlVgLkK3YPldgBo53zqGgI1OKuEXyJEiZke9CW1
TXN67bgzhIoHv1nbnF22vsfeOibSzZkcGx8UXqQZ6bRnUPAgzM1FWJ9G/TY6f7hnMD+ths0LKoS+
0t/JaRsNx+9G3SOcSbz6fvIEIsy8w7zdWfjRoU/Be3x+2Km/ALETM7PdqRhZKqh3cplph4GBrLZp
nZ+02bamTm1GAz5BHYTWNhk3B5ybBNdeRqLYuWr3aIZpUXANYW6Xr42bBMs8XgFWu3xAUTVF9czz
etdNTU8+f9N0HpSFo1EmkauSG7lojdWho8qLvP0HotyrweYAsmygB5kuk6EWEF5/zMDL6xstLC2n
JFyoaEo4qfsQPASF01o53L5Duj1PThnJ6fW+hADsv1aL2T8TfhJ+4djLpsQTcf3eoHIqmT1uj+H/
AoiCRpxw2I1LOEzTeLHcf1bq5cIre7iTO4EJmZIqohMvSkBImOqgNelINXp79jmjerxjcQa/nkbC
mEpSTk+GujzMnudxybwitOcMhezYR8/kgxM5iPvGQSEgr6NlRvwxdbjqRI5L1Wzcld8UbTCw+UyS
gYXQfPiVnYR4YTGi3dAJ8ijv7cI5TcRIGgK6bctBOV62U0s/1E0MyALZ5D83wOFFZPNWJp70yI+W
gimVPsimfPKu6A35vYKio3SVQxyMO4l9fKc095h4lVPOay69Cikvt2zFRZw8WI7p+d2j5w6BZV/z
YnlYcsDCfbYLpEfCdQ1V5h57o8Y8jje0276ax7ToqPi8W4nI75hxCG5tASAqxM/G5kpBMpRcda52
j/L+1upXH+XOm/35v0upPTAPwav+oFjqXtOXrfFLEsSRw7e7d36gHp7Dq2LCK2znbpC/D7aZPhyi
1FNsAbhSTyDRn6/XSgXBvL0QWmxbw6f7tCr+M2ABTYqvNfGqhlDoqP8J1qWebBSFUUUzZbv1QmWu
DaXfvpAO8d36txfFRcvTTCHVBRFxIkKZnzZ2qHGhXauHlTO2YlDpmykU435tp2gWdPIShgy/tuqe
KJFnKc6oJ3KaQjaANg3Wm2P5An1bwML0hBjKPCLC3f/JNJ+FvWhxEOvGwRfNraGc9ZKv9zCuCu9e
g5arYbKaeb0dtiS7+/FVv1GeyQYOP26If8CUuw+nWnCvoWrPzBJv+hLv9zbit4jUVU0LllptNkjY
LtZN6ra5kzaS1+wPG7hR5OH6vcWkgCTktjJ0yWGwZ4OuBZBTWHQffpLzIk6BU+1U82/RtjFPIVhp
Ni7FpWfHMG7QBQUEazW+SYMfxFkXQfJWOz6hbWS1NowQiVZ3EI+Ltd+U0aOzpiwCr8XwuhwZ5p07
Zpv8oW7Je04cAqqgmimteDSeLHOVLBFNtN+xlxw4A18YEFVQXvG6UctY3DDsAIYr+O9RKjXDtPq6
FUgFz6RJu5O97iSPj/9C9SEIQUPmwpkmkJejpZi8FnGDNfOEsMA8Z/oekneV/x7ofRXjgHg+v8st
pxgPQ+kV3ltItv3+ei0sZK2SX6ZWub+JoPFJn8DI6pkHBdqfnajtmbMXptJrZV9Gn2OUh7rqTost
EvmkZ1Q7y9uaozHjE2GiB74OlsVU7NVOBFKgMPJevpEqxCrosKB6zACgbMc4Z8l00QvNb9MzxhvT
VaiS7YG1i2FhCpbqCycGGYKvm1sMLvcnQWXKf/1sN9N3Rz396aoFFCx9k+mUKdYqlctK6hvZI6cE
wM9p5bYayPyFQt5Hs5Xqadx4SVTmEdgxMlj6Gpf+uzKIcFRR/16FDgYos6THeZxuBR1IaDx9Tb3A
ZKNoD8AHacZgs2hrWDIdmji6JOp9e91eeJ6D2EoLB7wM3IdMnCmi0pfSKKFAwXD7I0IgmMZ9JIqg
4x2lsSB9hgD1l7qEK7073e0kGXn6y7ljUPmzinLs8T9ENSc8vlFzO8s2Xho6mQJsydj776jYrKc9
5AApzBZXvpvKy0wc1gk8EHsU5Z1eFZaQhWaQ3xWR61I2a2Nl4Prl0gF61A3fdtkvQyh43T63J9c1
XzL6Hdlb7NOW8+uCq/HYrEStLKUWGsMK45GuNY00HCNUkd8HxqSXZkbkI2vS+0uTIkEwM+NfEMTd
+GIp6QjeGN9NvFkajCrO+mVuKrxfR3+wTRBOCZ6yQAf6mHGIF+M39gdFcCjSOSeo+QYMFpW6gWwX
8WUc6c73l9/ABhoe1UwF5okhHXGhrBU7zaVzAl4RAsg7yC4jWc8OpUNrqA29JNbYIYa1P1FObj4i
YQyck9vdgyZ/k8fNUn02kcXozogmJ7+o5cyha1CMH0h6zX4cknLWQdEWS1qfOCQAfPjqH1MUGtJs
SR+q6PBhB8h/RgxCAjj9l3MEh95YC+UCJZ+DV2NVI1WNM2bKvE6Dzb5iII+TP1lLSafHwyFHz0DK
6Hlr2MEF70Z3H5BXIIMRWcsik1jwlJt61ysnYeeAWgt1E2WYJcZthZGVzSOoXa+Lxf37a8JckoOB
WYK8UCyooufIERTXGBbnEZx5cuINVrJWTBgnhgFI/WNua4VnqU67t0bhXnqn3x116Yk/2EGIMjRl
ICUDWV9EgmZr3xDfcUn8AkPCh3if15h+0y/rHW9mSqwNEJAQXuWzDJHwZ/VDI8gGUCPTbnC4UYIm
er7XfnLcq3nz1lY9HHk77wjMB8dX2vnfnnaVkLU1gageB+DJe1ntEGtSuPdZL44mhg2HakO0M/II
VSloGQ3/yg7MnZBDtTblo0PSnq21t04BFoqEzprpjaKemgDPWD2LtNpRbFm6iZ2rjpHQ9N3zGV5N
WreLggOA+/rrfFVO5fT66V+33bQNbw9sx73OV/BlQn9AGFvoktXxTuYGVCO3RRZBt6gus7TZ2kvK
uoXkTeDKTPRBSnXcEgPayY4f9us35nptkuBdNq0z47rILucQIQ3EJ6gSAqfq4i+4XNullG18JoI7
QJ/o8t8LOzjHjr+prMPpuISEmukiLJV1LVTyzT6Gwm2cxxRn/DG81djd+6Razb+2rFd826uktLJ7
Wy9efgqBtFLKvOhfN2Ujy5ZaWWcdONXb2DMvoL3kX3qBQPjCf1Z3BYd2tJEDcVwYnsC4g56gdjk2
8x2JlHNMkWiy28Ke3sqp/RM1IZABkRulh1Z0UKn4zP5nY+oXz9gJYGrpBwMtjf1AKJLHuR/wUemg
vJUtlsPKHF11jZE8lP2g77snDfWwfl5K4K6MmtlqMkaOZ/UFVXBFzitGK+0XWT8bDIjAi8l9+GHU
E93Ih+LOXTTSv5vdPoGa5iT1THMAL5aiCPD014lIQKG1zuyrgEakcvGdGY0wmRiPijQEIpl/Q9rd
6v5KvmWdwLBivDdkvvhriaIhz5t2UeMSF2ZqZABqGoeUujsGPNkEm/Ue8H7sOSA4uj7rojyxmXYr
XMGR/x8rP+jnFAutrGchbB3+UKhUHrakSwvwJhzwYO77g1VwqhfmvTmoBY/WxLiW997PEXcy8GgO
rf/PF012wTa6dRMe6mxqfGyn7yW4dmwIoL5f5H3HPl8q+kga6UYgxGM0y902bFc0ctgQ8saoGTGQ
S2IetM9MU9IsWeu4u+fkbPBs46beJ4jjBilxxnaHXscOwkxnDKfB3CmL/A746EgiJL/GAiCas69O
EZ1SA9ZPds8KwQhE2nNSPfx3S/KB/Krbj1P3A6/JrXk+CkGWpcQCDpUikfntLWTMIilxdyKbh2U9
74vqDNQ7U6Nc7qk/oMT1Ss729Z/9QkpE3RYUoHcSKrCaDgXuJki2BLu8bzdv7BVd/zFO5dS1dptL
OomJpDLmHRUeukEVYAP3m5rEimfMhE7L/TvfPjy/Ueb6pgwnlEhKddXaQP9YRdb66WWclg/eSS2q
UBmlJYiFs4fwwx3jwX9CZGJy4T7XMrakgf4VIVh9J628RXyttl+AKNODHBzCzgNzF2br/IoVbHrt
VtWglDiNY0umdSkRjc0bo/KnMYvcrXcemakvsrcM1rgT2yY+Jil9YhGo7VBqI153m0Ac/pL9AARn
wAXy75uzKD4TZlsfNCtQmS/ZbwMvVMgk2errZDMoKnmGzIDrj8pqaDIfhNc3vTHEESl9XlsZbfNs
m86WeXjBgnVrV103fUc/ThdRWPvNHevDi+N3UTj2eehO9iQYdXMVj5pgd8Pd/lc0vnCc0GVdys8z
6EZS5/TLmlhMssxr3zTUQILKXIB7BtG8HbXtlxfexVWKYeA4t3eV5nlU8tKqP7r2pdMdc7/6iTzk
D1dTQosqrJsv3sBG/8DaUEwuTjS34V47qP3UY2hqbMQdBu28SsDrrEJok/T8WossO+666+RFx/hj
DfzYQT1H3/UnndSaN8gP6d8vQIveT8yq65BX16yAP6FQXT82GNFdF7X8Iol4Ckzp+xVEACUFDTcS
0HtOvzqgW1RvoEwOEOvfsmey5NfMIkYXp/XobEqB9hk1ZaafCnwJOQzWg4gAqQJBLfbEQ1z1nXYZ
Cr+v8Soh0Gg0WKTJ+qGwQqGb67v1pg/jnlT9sNvMwZYCsFTIxwjIdZc/wmZn6vv6yZbZSg42eJO3
FBzzBNsr7RpXXhdINyfR5ItHFN6zUcbI6a/MS2FObbWpCYcfealHqgyllfcuuEnptkgB9O96916g
6BWAtrtMG+UIAN9qGy6LS6Zn9pyyBZsNWtDHOmleVKE0tK7/2AfzVG45sMRS3TYwVkSCdu6WEaYx
pXhjvKdFlxoJnndtiW+kXHZUgglo2LwKpsiddXdxwQYPeolasTShzolRJMrE8JgUSRS44TmatSLB
nTk9bi16A95bqwAcH9uzS2GtxL+BJqmrLs01P+82vFh3emfXMEDfRQ3nGnzy6b1hVyXxbe8h1e1e
yDsR0B75BztKYLf8PCmkd3oWfpCxc25t4RZhet0qfWikOdxCAhxUi0LNcu0M4G4x/+0JY/JdUwRA
DdDyzaV2OFBeOWOUihC0BXcdeDr4b/ErQMxKl8snkSdBQ6WxQLF3R5IjPkDZ6IsxODrC68pN2eLN
qm8fK0A1ts2+zfM45PuTLqHXnwbpQJU7nYVEfR6AgcUr6w9jfoCapHoR7ek2+TH7r7iGAH2eTmQH
hO40kis3vUq2UDOHb+/b/0P3sFu54R3zBFMgTcqbi6B+ft4HHvQrfKYJgpDRKHqtGEBTPB3c+clt
uJSaqNX061daV5VFAJrQ6dP6Apl04353g2/Gr3t6o2yef2Oz0NO8rW3EXkOJqVRhbiSdw/sv3o2d
UX88BHiJHYT/bXgGCK+/Eccpdi9OVHkaxfIj+XR0YCF9zNfOo8lRt/2rDm1gm/pX36/e+hBUHiVh
lnQ0dwz8jCaKz1pl7eJxqccMrQOG0QKoVPLFAYkRu4hF6SMStOj4QAMc4XksrpHNuKMsbu0g0eJ+
bv4WTgSx3sx2ysfYAHYGC3dTMK1CJ2Y3g9qHyTR4TymXmjPW+NapumjmaHdRKhLL/Z6oSqucqD3T
fA8laUcbYnRttSBm2savl25GJWRZ86lKeXm4tABOFV/lefZr6ICLvbkpn/BkDGBG+vh6LfQylf7l
RSdFuPJOIwLw5S02JYGVqIe4yMw0WfKXgWFZ0ni3bVnVX5ZirNW4y9nMWCkgguM/WlKU1t73mZPB
cKzYu6/JbgRtndNgyHdP2jSJv1IvPFSSWrt7Ai3FQmkEsdTqUsjO8KaqqyiGjk37z+lJnXyvJFIb
Lu/CSVMiMCgt/I9tkG6SvBQXV89+91GCVpCPdfKlt63eBWZHzomQNKrNUV6UXGMq2/nn5Jce1ODq
Xg55ysE44cTA4qQasvJtlmiqOyj0AzhhcpCebtHVEUjVZDq6aBhpyhhlZkFkKZccZuaQQchTqh1r
SussYYa9Hj8pLx9+w3fAvWhMaTVllTEMDJU7ia/SHxto87pK92ppT8yhZgnrXsxC+AitWFwtL6gp
4+Jr3/b8r4xleJshfpwdt4UDbkEdWsf2AM6Bwpr8V/EneG3hPyZxpmdWsCYt6IC7ZOybw9hq3vHa
UeGx/yPp/212kKuAey5ndhJ2tFwFFAzzv/EeSygVqzqqvFVepxrVLzzL35WJL7eqDRfLtGHksYiN
V3WfFjGJKY87WVmmU0VgedtgCOF8S3iq2JrAO48YxGQQsqzqSPPjlmIgb/VZACH+ncouyPB9i8Bz
PJswFmNOPQ9wPJNECLiZOU++Dumv/JsWc0hnaf6JN2Wx77YV8Nyor5yw9FDff3nN/lxWiq4GOfZL
r7BN8DHKWhZ3cmNjHFqeeiEotv5CZcSnqKP10lPuXygHnC1pTLkGNuzRJ9Og74a4vi+rYDOwJFGW
ARsfzZG8da61BekAf4yKcXhvRn1fVlVCXpwnZx71Bit1lKXvPiSeU/JVo9iXajsCJFEtqTQmNSf0
wzi79ZreXMZ9ZiHa6vBfGiCi/xU3tVI4nMtjovSjaK33b1jH1384H5vg156xO9CwNeLJBj+o2oi7
VoEC0zqGG6u/RKeQNDjbM9jc4OZPXTYaVahrj6PjUWTio+O79jURSuZHJDasjjo7S0g7ewh9V4zJ
KCWIYt2KJOawM5igPv6xSivZpF/7PXlMrzdsvP8JP8ZYM2IidAVASpasjIvH4hrfR+pfXtkeEbGt
ZwtTW4nTI54Ym2z+L4ijtw7vwRvpX0Eu6EnqhqvVoDDbYeE5beU9FCECAmcl6lro6HQQDeK2NCmV
IeDL0KypcUKdB2pVrUnxoVD3gvEqkWwfJBifTbjaBi88rPC94wQoTeGYlKV9ZthoWYqZZBbKXGbT
nTsm51s7HYSGzumIJWG2HmqAPfmA7ixD7Vz7fGUL9NtZtSOZDOpO+BlRKE6jLCgA0ZvzXuh6OSNN
Kk8T0dte7/vbn1VK9XD0uMVkicCa1Gr3+7qmhwGTa4TSDnls3GEb4Z9Y01lHbMBPFFgTb5bUI3Vj
fiyBoWOoJypzuC4fDAO3zHJRrTVVlz0bymPvwvuajbOl5dgTzCcu9aOGrX7vhMAyyODMYNBNdH9U
4z75ldst1Xz1TkSxey/uDCb0UCU348lZ+GoTz058Ts/+SslsL6wju0+TQXKI9p+XuXLjzB/gz3NU
1N+EgxdURFiBIDcUZ0fipq8b2q5bGh0NGIVO+JHDaR4eI0bv9E8uMIRZH2JR3SAwGrRoD1Fogr4r
j6Dsr6/3ffPoAdeARMKAoZrSbUejnVcyBvChN3Tk7Rryg52h6D+vpSyJSgWXVkK7HqNbwriUewNY
PnVr8449aP77UGEHZ/zcmbHs+rhd3iA7lIj3gm7M0rvDPKMb/CUDJ9Ra9Ziz+u/jN33teEzJbR9y
e5v9r09oDQGL65EBOIDLpbWN6ZeIg0WfXXGjgBSsIyLTQZdaIzfAkAFvOPdiVEMP+fXhkTiVub3k
UlDEn5BXna2WKVkyH9PEZu+m+/IDKyXFDULeaJbHIVL8WysnIM/OxsQapRqKbv/5JqVlejw+Gqcs
4Ve4sR4JzSMMQLshmsNYTzQALxK2v4WgDibDuRn02m98Tabcoa3SEx7oSxC+pQaaSv5/93d+lMu3
egVanjvr2AlfHmrD00bHwxR3K11olgZ6mJEVx3QgXYTKHpLiPOa/Ex3bMetqZcfmmWOxyhWlS5Yp
/E3mhcfxUEL6nlEdnWotrP7G7eK1oEh1kzRR6MWePBFjtd0i7xydQ8B5zmvi/YB9tbWU96Qgmfy7
SJzPEIgSv7uMLdTxzLcutyMJOY1M73NxZTsJSZeQePXlpr8e2sPJHmXXLMAwCkUrNBqGPOhrgDW8
zfKQU2NBBHFzc+YtozrPJd7VWOIu94aL9HUXfT36wsmJfVtIUK+ipGwoR0U1ZA24l04E+5w4fjev
wotY+5MvH0TlUsLAmjWEbpX31wWnPOb8R0vt9laCtekEAq7Qaicet5nnbUR7n6V236Jjiq855Dqw
9I1BdYtacKQL+HQIEd1ZZBHFcF6kItGVld84Vtow/zIv1+yebU0BwI0Le3o3LuD/Pqkd/ebE+oa/
3OFkPhu9mvcjhRK8dOpRnYPn5hs0a7O3Igvp2z6T07wc3jw9uOb4Kdzz2sBeGnsgMWW11N/a8Iyg
MWjuEmB3vXF6jnCrbic4lgQm4sT4fomZbL2vwqQxxA46rO+D1cHQLCs1q9lAZuaA9J+20Awn41qp
5GiURbWqbc2HSL6dJQqjRiHK0G4cWQ5FCYm8hTaknPRq9wSfJYjMHO6alDw8qjTYdUelcjWC7ZnY
XR9SLs8p5RU/VcdjkvHEePTjZFblC+10pUJOMf0bw6ze3n3UrAB9pp1mPUF3zhUFD+iWWlXA6RRr
2tWj2groqZ/Md13nwjUlLuFVcwA8kGdA7BsJKDICIDQdd4u91L8WeW7LHqrf/b9fGTOtBz0KfH63
I1DifFbi20CYUSErumauqNkpVbSHBWEFw08jMBkGeiwmDtFZPYmkBvO1ldj4V9ra6vk+M0KysNRI
3h2tTs7157ZtEzlIzM3cfCourJTkNCkzBCokNE7QZF+K2pGd4ut/9LpI4c/R0NqSC0VsEVoz+Crf
63HJ/e6aeioAyRc0AzBzJbVBaQ/PwWskkgXma9H3XawaqDTpqoZxpRnziaybOTRx0U/7W9cibZln
f2Lcf8KCC1pFaTx4dav2QIjP3cTvWjGxTy7/pTaigp0pNwtRyc6RIrkWh0x98ygsXBAA5LkFGVcj
3mHjlRzktm9nBRPLxI25fVC2cyemEwTBZNbYeEwsBM2E1KCYMQrkpHD388nxImwn9opNB9Df2r2w
uM05Yqx55UhSN5SLVZkHsqiQhsRn/7HrT837YfGUyLu/ht5xql1FDSrreBg2nvCPsVPNgfSgzs7Q
JQmvcMcov8lx0k+TwDOGGEKXYfR97Y7Qy0AroBrzeCLIip0H+vikJ9SZAkUdv/iAkoY81Jaut6Up
3hJ3NEMJ8e827Tfigyfz22JTugVXTRnn6zUaqIKLa8z/UKkpscmuFdCqHNYNq0GYB6Zubee+K0yH
jPRLqiFwbunY4iq7S3y+vugtokwFgzsbnF7jdGs5lIdjnD2mcGk7tsEfbIKBEtdMOmnvUq1nQrlV
iPZFgK3/mgV6uik9c2bjBj9ojgH/CkkgCP/8CABQjDPFC338IjW9mt6V1gUos+A4gjsjTxUt3sr3
5yb9BaZ5Y9DfQVwcTZLzAL1NmiJWZIEj81sySxLPm7m2oBKYrHqIOnwWs7aNWjAhO/tnDJj9gedP
RgI16GvRtY1SPq07oN7cyPXW4fIFnk7MdbwOSNzhpfR3pji0MuMjShcdKxgkZurj+TOGwCXaFcvF
wyGDD1inSkVLhOBClc3rgHTA7E5Z8sr/04z/YOuXKXG7vlZvG+yCujp66mK+I60QaKcWHwRjCnON
R6L8lQRYsbpCJzbMDagiSLccm/ere96+UqlgBe5LOBMPRlyOiyXO7hWvhSuJdxfn9xM04kUChrVj
HvyMgiPHOukKWuZodATBzJsGWCiI07rpBFYvdtvrgQjdE0Bw5xZETL3LlUmAyBQZKxdkNmY7Esc0
lYHAVKKUkdVE60MnyZ/Vnjr/9vRGy/jFNoRH6A1xtVY4WNkf0C4qeYE0gjAdBefiu/cmBjtOvZq9
6KIMbHY6kJsPBDroSVcHIZeQDX42BKR6hjN+q/j2MzTs9UTbJQsBxl8CT9nDB+nfZRF8MJdGSRav
ddYKGvLcmJyzvIgv/2xIx03RlX6UNwkIKw1VlbllHDdnTi0iTX05jhqVJxl37Taf1bBMIPg+kNQO
ljTxvI6TOoO1ExB6l/Dvep+g0Qh8XI8UBScJ0TjkkhpPykwrQXAOeHRuTYmQuju+XZ/eeLFwRZ93
M0uW3ilYGkeG4wzVmwZ+tgUkUCkvTb7x+JnoHQ71VK7cjgMt7HOqNZJfJRFTtMnfOhGKsVYfH3oD
sZ7AP9Dbjm/xIvpbsyAkk/BX1pFhEjndr+Kfniu9wXogBIdvtlzkAwAkrw9kmyesT/HX76D0g5mY
RROuuRytfsbPHgTy2Nr0NpLPnZjPEpiUZWfxjAYfGl4EXiwkCsAaO5UO7WvIk5yDLoI/y2zUsTz1
3BrOUN/ijIEvTxapXXOFpJCZkKgtZAcxqzxP74ZHVtQJpORD9Xi4kYpylxvw1ekBS1+9tMLjwBmD
rHnV+/QwhWRwFdPXww2j4Ak+CJEit2aV2cuNyTBSV26JSCRZriSJ3666O/EHqDiOIL5kQpfoLvHP
QPrjIkTtINKAELggZOI5pONPwGcVuZxn/70uXRAz5sbBJeF1VkdeQP/5v526i1RiyB4mfvZLQXmQ
5PXKRLU2XDAY7vVrEOqhonPnSIbsBXgN3FXeYU6xEgBVaSMPqw3FPPkD2dxLb558VR/eYn9Sefhz
wIgiEhfjJ57ttBtB+RwJ3gOInJP56BUXC6DU0NgLvXwlJRRWGOVfwfcL48vXAhWtPSqPTt4gaTVC
VQBJHtPI6IbiODV60EHWxMBC5wQ6zV1SnqViCxirzEZB+jtdUG/93ImkbO55iy73fh+p72Dnkhh/
eGcbOh0QcAL1dKVb0H0BKjMfGvNWHDmFtEnCijM5gWKjZ32WuZ1G7oq7HE7RpISaYJWFauMMbPqe
Enuc0kPhYNPe8FE2aB4LQGgCxr4qLq6ESHiIkc3lhTjklr/BRe/KbXos6lSoMcI03o8m/31om3Vn
Q6FGPJmRsruufBJpI0wd7HQp6iFjhuCQOf1JVfHm9xJaOtwkrDTk/cXRweAeryHa3FZTadV5v1CQ
JfFtST2EJ+IvNGevN+FwSRZFcMbg56155Gdmt4XXhnFTGN/wPnN7fJRJsUw64PUfXRANvlUWJ9X2
m+5LHcvM6hVjfPoFavDA/Y3O5Fj418US5jgnDoih6MNc1gzFKkIdLED9ke7jjWK8sWj2WPON7pjX
JLJO5K0AcVJ46CSyd0TJFCZ5AmGLAtC9ROsCTD2yNeGTyQej4lsRpJa6qopIJbS+hP5ilcZtWcgP
H+JiRpcfa/Gz5Tc+gww6zQsz0toESAwyYHq0cmQnkRAAIC8+alTpTlNxC2kOa5A+L7FaEWmLCeq5
4JPl2CO3UAAac7ugvsYTY0V3zuh7St4vPFTcQQpvZ+nJ8vBpqHAHkI86dW7zz62lSzrO+CsD7U/M
zhJW1OcOzNWmIXTHvC319Nw/U2V1ExxWakDPzVBUVq/c5C2SDFhzEZbIodxGeHk/TS28xoYhI2NG
4lBakytT8a26CwGCy8Ka6Kji0AV90NKjAj5sNItoyE8R6BzQvmZnwbv5738YPW/gZBf9NzJMRmCN
v/PZwLkgMNybzmBZjnK11UNPE4Kkzkf5oQkQQccNHjfZtC2B55x8S7+I+dxYbCrJbflH8NjpBxa8
ZwQECpjwTjpyUTcS5JksOWc0c0Yf6XVsjURzdrM8wZwWyBEnBT2Hkl//xMn7EKou19d2hJia1oVL
/abhTujEODzWlpuy6Uu2ZkLPOopgtYWRMULvJjdB0o+A4kZ1QPqwh0/Y7o00D68KID3KZUNyytY0
zCtJRPvwI2OPKBKfVcPgSX4Lw5G55HybGnWoVYUcfy1O+0P2jPAObKkCt324GwwRyf3GwVXXyV6p
JinYi6T6D9La3IbsixlcAo1TV69gSYPcOy9dHSX6JOLY4NQIxCjcAVC4cR0hihhPTVZ3GmMwD1NB
EfTZjlusT3XSGShcOnKOU1DfE+FWomm6k1sk32UziOmz8ixMtgTihxMFTQrPHt4EWJx7t8LwhYqU
SJe5VDaNCl6izPZkAWCTeu39jshqUDQscHGW4/AQmUiy6WVzEzRkG49JlK7IzVp+qwaJf9KLSNG5
YplJk+NzcP885q0oa192F4sd4oj/mYOJ1SWz/Hy4BldsNLY2lqA+BjHmTfYmgd1ViYFD+qSwUNiY
UXi1j1KdX+Clsifh1DU18LBYTHIER4vPuRkNhcvfmUW81Op9RtcqYgBhKfRh4EHCY1g3LC65TITe
OE1FNGbJpp15EcWsIhv8y2Nz3nLdycWoJKx7M16iaTzuhvXkEKoyE/dmUG92RgaVyr/vNTQvNOkE
vjUZssmsKLl+8KujGEuFtgYQvQo08kZ3sYF1yici8YXZhuPJ+VCWQS0m0sJhgADz0vvk9yBSSDjP
RBOTjGE+Yc4niQolXKzzxHScZkacCwHYfVWtWJF1UdbOEGUeVdeZjeeAQqTgcCK7v2aYiWkahIKC
Q3hs9ezQmzEBNYHJhRGy/8EXwnHzyh5KW+ELV29LJgIlW/PrmnC21sIpdtd2jCJgD9LR9WZDDa2g
0wlioRw1Hc5Yz2UDmPsjYeOp0NrWIDalZQPzitP7a5GdKFB4E1ohobhX9lohfgoGmKq+0CVSS9gq
sKWVAImvoWZhDCEjzDfn3vlrgP8ZePOwGVG33YrseQjVScubjWOGM8qsv9/hJpqkoot9VUz2+co6
0hw7Dx64lsBc0Aj8PRbloUFVje8CqMPa1B4ZWbShhjf8wZtpoRn4LbJQebRfNqkDcntYUSYv58zI
C6ufvBP6E2oYzDf9GCuQOQT/osiNMQqXuAuiKH1KVLRMjIx8R6sN9kMncl61KSCA1qhtPn3Ur+rD
skP7ihSnIdwOHnKfmPfGk3lYS5UGEgLUTIfZVI7rqzLL9arkYPm7H0ZuLQT8fq+275NHLkmSAE6V
12YCQ07ieVGK7cNn/a7RDzMzcLv8+alYcldn4p5jclCraSymhVTMrxu46C5UP/AXIVvKiEXMIxOW
GLVrbofz3QNvUfAt0JbYgklHa4b7wIB4JCkHbnjC50o1UFU26WsS3+l5sbEVH9qhik7zj59fYgua
Xw1Mgqf4m2xEeai+a/mf9LL/GeKHS8VfUPuq/qz8Kh9FOwv7eXm+koQWuEXLdOyaVK5QMRFPouX+
ea5qQy9w+e7fu2v4ZpW4uj5yhDaVNOwv3LEV+CSPHxIYKh3eRgf1Llgfy+gjFpXnAbgpPXblbMTJ
i2AmSHIPqm+bZxIWe4CkQYgKmNUuYSEa7vHonKHnaeIqNOChEf1dEatbchS3GAvKOt0+3Q/Y5eQF
N82irui/TNCXhE7VhxMSGMUD2hFP+HMiVBamWklENcaETjbXpw1b2klKsRIgE3ifz+iXqe16A/+F
dflMv+RxUKMOMvA0BJnlMa8SfWfY9EViWg/o6PNpCa45brQYYi+FfDG2ZnsFbW8mBa5fKHoVOJus
/QC/sxGvnv8qWVtGa6rFkfo3ubPYXOOjyKaaHF5YKLEuaoQFwQNChX6pFU85mryIDzt25EYVvjkg
qezGwgOzYR7Q8iTo7ut4TRt/nYKHaLr1ps5sLbWagCPQyjFxTJUnsinCnLyUnLCaGhQ9GxkX3lzJ
pSlcTzu1YR0HnO3FsKYIh+VW/0dVnKEZSt18aoKEHKgGP2ElT9I2iyznpylWSjpnX4kd60+KlaAw
oiCJgRhefPMgFfiuUz2HJg4XByR6qmlrTgNE7oC63dWw1gZrPi9++0r2dsl7NuKCpbE78vocSnga
95p4UWMzJCG4XoAlR7vUMlIDKKiap9F8WItaHGIFG/MUlA1NKTH3gXbB5Li/cCqUTzsYyOXwkIwS
botXaE9ZVbMsRunjlsehTqhLl8dA0OkaFBfC+7UrswbFXDHXHL1DkPTC/NiMtaIJ9VTyWrl1JdmY
ccbgejIcewn+LolZIGiZ4/gBO7kMJj72iVyJZSdbD1EGsmrPWUyENd6Tz0GcQL3BFXrZO3D0aMTC
I4xAdUrWQq4SEYOornYmZ46aBd1muWauuG6m5uQeR0n+TpIL5imEPRekR2iwQYLiNPODvSraoPt3
H7rG/H8MPUin4fSdhF3ruBtT8z3yIdW9P+GjsxmSlA8aFII4JRwJo4W0vWhp5mcpmFrf/k7dDE8i
X/wgow538P7OBWVJMXnfMR7aoYTuhmOMRPiFWGmgLR1Ork4ck+ZPUrd7vHesvMuD0/rOZ/K5B0XS
xWBKJF3uniJrp2qgAznMnaPzlH5zBVgOrUb9LoJmRCEP+sezKtYLsc+twD0yqZXxwJprmf1ty3MM
GxkifXLp3ynNaoezSEZ9OE0IofhrcMR6H9VnRp0CUBw6d8H8XmjNaBVdSMkfy/ErSbButovTPh9c
tLNfgPIdS/THIT/Oqcr1invUlSyxFvtfvyLme1/bSSMw9fywi6IEHdiOUw+MKEgs0+OCN+Xg4eAy
zcrDWM3GSYd5HFJ6iZbaWKmp2jh1zAjYn+IWk9OILAQhJkDsOWYuWyJUvU2pbMUM+j6ZV1ocDU7Y
oELnp0O7sjWE0+Dm/q5Gxy2Fh9B2UVgHWL6FSfUxJhrPDnCyhSyn+G1QIiU8t06fu/d6gImuto57
mKuu6ElLauLX2WjEYFzkI6h60dnOIh5jmTru85vCB45XMUgAjP9TorrRlHVEUZhCARg392Raw3sv
CeszE7DXSp8CkZ0wqoaeeZwQJOZsUHZk1U7DE8ROf1KseNzTQMV5Rr9hRE/B3R1G1tdfyNz3iqEw
Htd35SSQO35Yi+FMDYnrqhASAR5Li697CwY3F86jndNAGY1O51C7mjHpHke8SoFRyhw36jNK9gVr
IolQWyWFpRG9J4wSKREdFqdofGHeNRbmScJzP2UTUNHK14No6/+NNd+aeBEbwUqw8YJ5dD37Svjo
oc3ibHCm+vt4i2JXL94tMYXmFnMZvMECcKJWuKGYxJm2l37tLcHEHd90i685p8ANpAl8gCg5xLav
OcDjfxQPVFsVZc5Ug55d+NSeHppVYbG8sZCall6799DnZpUwpId7dCGyURhiVoIUVOvgKXMy+wWu
erYvpSUdLE2QllgvuZ/9RH7zwsvehdhAiHvgSqG6m0AibTYZgoLRv7pjUWeBx7DOXSkmDPRi7OXS
9a0XYrELapIFq6jYjxsVafWeGUkBuK96mUaXKTcb3grI7fNc6HcWp8dNGe6u2Hb/C3vlx8fkseRt
ZXjOUcDD/mSQvpER0J1AHPOgwXLWL78/ulIwm6+mm9k1x3Yk8VyyV8dfb5MrGyBDbSfe5YgGG8gi
BvyLO8bCtJ/gM0rJ+LmJZ/B1A+ENu2Al05INWALbV3jfosz4CxJsENxVrynmHCFuHitPep0M9C6+
e9KjOLqX23IdnbT0sloFucdU5f14z014rVCBee2Nj9aqadK8ShzQ7kGUbirZQ6ML/xDOUgF5T4zN
hnvEnSjGqxWo27pylbDrop8HX7cmzy95WUF8KIRtSSADR/ciF3954oFztgszHzTa1arem2Htlkq1
eUnHmnOlUhD6JF9T15AiiHwJrwXlud91vCgEMJPdKapS0vIHUktqQps6Xsl5OdP4de1/vzlIM4x8
KaQZQmN9v3M3mO/Ov3QCXu6zpqNPmEmBf55OfZbS1xfQpkwDjUsfvYLzATGHJHRO1zT1lOMZQgaK
52aOJqxIff97OLv/fqchdqSyOR6zzaWX5WEobvmXD88+sXA1mIcUv7JOeZc7RW1/XrjrtyQM3bMJ
8yu/CiGps07JX9CdobaM8IcQ36+u8OzxRb7NaisVvjar0bqcQkDLgALxa4sUfIDSxPe4tpeGOkAB
YpC6YkPsYAu0c20lgh4TSIjI8rQiNwnUYeswiGYuN0VWeTmWs6TmZ891Hsyav1uUjiYcAr0Y6MHQ
3gLZ0r9ImTs1vT0RwJJnpEFefu+xoJDRypboyK5EytnoJX1gwAkwAJUSSkQnYIzWzkIeTy4sF4ii
mUnJ5LY0oexHw3W26AZwK9rvVT0HWYenKY7fBO19FlURTWoTguMAwXzIcseLayFEEkCVWxGdh+vK
yVidhYo41vvo+UxHh3XQEbkvkL68lOczhR6vVrjJtxn1tf3mfcGy3HGvx3KFiVex1Zq/cU64ai1S
OSU7e9FgfmISPo+LsJZYfuOPkLP1xh53PXB9wGEvTsXjSbIDeRHwilG6rwn/JE7VA2RGXtWLXZq2
isrHvGYfG+rHuCy6P1vmP4UQZF9s1dyup5q9sK0Tgbr4xqWcfusTXTl8jRBLVyP8J4nwtBKMF9X1
z98nV7dlpFPBb5znfpcvOI8qhmYrlxFvQpMY5R8ceslkZWqP5vfKo9rIFCztTXxO7pw6VHK+Getr
T6IjsyWqlkDswk/NRQdUmqWqv5osLVgJ/vfhBjdpUDgngQW77N3Wv3Sz7/JPvW8+FfCzjJeifVQP
RmsM0xRa8JtPzGbsJYCgoaZAz7iWvUK4Kgu1NIZjaGXjHmlpaw2TvTLWl1u4WzSs35T/irJXoDT/
ZraE3H+YWeI+nGzC0/+pZ0psfeGwukGiW+r2Dq3SzCnTFP58NTg5FNvgVZDL69fn8gCdCbyjbDAK
swBcaQ3K0B13rvPwdMRi/TpWyIQ6y3azoEoWAqTrved7NFVWeZMuVWCJsyLBoCABRSlxSObyH5wu
uvXTfcRPr9czVKjBNkYfvCdwJDH5hDtIttKk8BM6mD6f5sVCKiJnSdP72Y3ZBbC7KOKcbCVOZr74
v/njyLFoOsdCJ0fCNqMOCZwUPiw6hURVNRpgsdE8ZXCK274kM2xeFhjz+Ds/Li34JtMQ8DT5a6j5
28LK3BM/mfHcBSZU6S7E1VaURbc4VRHIAKtZtC0KccGRbVNlrVlzWfXAHzl150QEtYPLO4456HQr
Qh2oSQPAgjfTDKNQsVuKJAa6sv91iQ21GS9tK6KMwrPWB2Ub9V9P8WqbvOoLgrVKIMSfbwprQENJ
/GszwcWrzigPIB6lDk2+ZgD7+IMsLCWZyrmGhyWk8u5fSmz/zwXi+uQ6jj1McVfraQQO6WUKOk1Z
UDE8ptCXRSPIjKuf2ktZQpfp39GcA5sR4tIyTRFm9ubT5R40LxpGhgGVXWZ+S51VgQqZ+SaiN2YJ
KLmvkDmJRrXX0BN00wA0mfKPTEEyWPwv+56+lIQXSTcrDUl9LmSgVXkSAnrf4M7zsVm2IoWs3S0b
LaULbgzlN7oo1q1RsjEUMvJUj9RV/3gQJnM5adxF6wYdnO+1Nh70YeMB7oXFVGywyrYw7QrSCP8x
qP/ugrKpNjzP4vCMCAXqLSeE5kJoIKFlOvoIwVOlEuG6WzujsvvrSM0+TDbJ4MBnptNEmrYXISyF
8KjHpoqwiSIBD/+zp1IgrmqXgtLPyCq+5XXeZqoYQOLEiYm/Vep6Hjo/LfFmvxmuVn21aTCphMwV
B6SjtsW6C9Hbc/9jmML1Xyb5kyHR2DARUamC2ke0jd6OEgGERJ8pdXYmwdRMn7qioUCHSKGUMGNE
ahIHv2a+b4L2qq+oz3EcmTeXfqzOMWuSmgmqOn53PMP/onZrYbs3KsYCuQe2+pUWN3vJw62zGYoo
UPjylFZrRTP/wEIPz6M3gZtYLukoP8195sEVS0GKfKDDAyJLkrDewKLEGR640QdjQHRVIDD0wHaw
m0Xw7SKUNchquT16L74cf3JsRWLEALJAXsLv9bZyUTYHAZnKHebqCWiQpfU7/anXrs6dRQfS6EVX
z2NYQ6xval3IqL0q3Zn0SrdtQUGdDLIia/PvQbX1lm05t5einpPTBQXW67NkLBRn4a7SexcszXv0
kGI1nmTKqwhf6UvexiXZu7aSVWLDQp14Askt9u2cnDtwIICDETQp/IIcrwE7ie/e731VKXk2z+4s
3NxI/PTwzSaQDGMsfX3MYpzabdQdFBt/Nr0EAOM+y0QYVEqr8ew+eQzi5P6aB4oNOgx5Xo+Z870V
00fW32vLBk7QAG+VNqO8jcodIoUiCk2SOv91ZHcvBQYWN54kH+KC4hbr8B3OFy3bTFNZVNsRSVLw
Ik/NAis5h63cbAxwypZ0ct8Yx5GVYdhhv5wkYckctE376E6ugvakhhXZriLND1+WVcALX8FGQwG6
pF8sdNojDgOhe0H4iMk/uIVCCgg04aEQAvkam7a7oue5r8cTIjLUTJYJXSMCQ64BTyH4jc51KJ9L
v6DvZThyyrCDZofRoNVaKVvk2jyEUGOUoR/0ktM88xVFkjCU2FTrLBPCSBSZpfXKYa7YAqEtsKPZ
lULGsMuMxcQc5qqV2VMKKzJJ+jcVu7yzf9AqSOxGC2s9opFR/PcmnQ4btHoFMdHLEmesw8nI/Z8L
z0Uc34NzS99l5uRE4nlpZI8qYUifTHXejwEjcm1uscxW4CZUMySFZmntVXXpKdGWcrbmMdl/8wQ7
9D3eEQ2UU4PQ+360htQwvKll1poWbuZbt4U6mhQhQkXjAJoDLh79DXT8vQiYYL59n3vBqDwKqCxz
fJmz5WvTecd9ufja2TMYqbRjKz+Q0y8E5yuZMzbHouCNvOKERuSgSPiRSEWVMWzG3FhUrDKu/H5c
QxA0o4MJ0O1FbJVDWlShnII8Jgwtcwhmp/fSEi8qQ1+Ga4avtr0ZWkd2TmZ1DNHTFUt1dMNwIymp
Cj3lKaoYQMeT8bRN5p17LKqMbhP10rwWCydrKRIIIncwTleYsMmFMmV3xZLqfCAZcI7WmgI614mv
6BRjrcZyESuMiFAZ9X/F/ykPGRLlRhXblZACDR0q2/usvDaJ4lvn0uAbZnfi9mYhO9vAhh3Y+mvH
9AM/vqV9Gt42CQPyyvPBNjdAg7rY2M/ZU2FUOwz6R6J4ODQKZitFsieqez247YQzLvkbMat3lAAG
O9fg6zL99XEelVz3k8rnUha6bEsHurZA3ckQ2RpnesTp7CP0pqoTQBuqMe01IcMDaYn4eIYiWrYq
6ys+FQZnj0CowIp86Pdcq9AhWbIhduVkqiObIayFIwo7Ui5wsHAdhsbqi01Z3Sct0UplaosJIeeV
PZ6+bq1qN7vhN1YOqbUbXKXPrCwFQiclG5EiGE/apC6yOqIP66xa5c+R8spfyVwo8QzdV1kGc0iN
Xb9mDmvd2FrWmnWef4isuJWPN7UObomVE70e7ibB69Q76bP+/hEuRJq2E8hvRJQ3NvS5wsY9hhvt
J4cjGAYP2kFBADXvLDALZpHFxFRXnOqCrqP32UgKL8qiVI4lJaHgeT8R0nFeMTWvPgQxBv3pZHao
t+OeKbCn8g2p2hAjV/TKmrOhNnEjjQIGHZI6fq3BExoRYrgjqyE23lRHrSeq6MGoKysaTs5W9OH0
hA5Abdd3weWdbt93P+9UoJHIzdC2xLOG8C+tT9GuYobzqQkCPRagG/e8XsinXSqVfdEPwvqXBAIM
oIY/MmVkSMRmh2IFujS8VBll9cQ3bnhCRSTXBodwuabRRc9G7BcVUltpU+sUeHv0V/Rt0M6Ny6Vy
4i+lOSqGHhFWNUS3twsOkenirMpSC6jQTS30HgEsiHezBb86GLLobzj7aZ4FpVTt0NSQLUpQR8Gt
r0GC6ZQGQCQhL1CQv6jLMsIsCbNHKMXY/tcdGLSiqApMfvPtBvi1szkcdzkDacMIZoeskvmAdwFk
OCyXo4v7bWF13zC/KaZcvqJzkIOMziPRHYfFNSKsTOpAjd7TrOKCcWqfRCG69GFdNtyd9hrxcdTB
MsvIXkpq0awWZs9MqVgZ4efS2u5dR9uorUDRffPlg97jsdoR4uq8Em+oe3ajjW7O1XMpLDck8xcw
e7RNJJVjFWFeRnCOgnYmebdSaY5InyHq7oTxLECqTOfqcjlwyb9HMrRRyn9xKFoZDd0t7bpO1R6n
VfW6H3JeTRpBA4PhnHzPuq78UnOJ6jKRp2x5z6kevARvKsJHQTvQtnLQR4/2vh5IeZWCFf6b0U9W
ImJSUey5iv5eQxx7ivbCrCpaOYxsOsHjq8cgL9g/jRSOiAyiCTxmGacaLxB8/UyjiHIw/NZHomUR
RAvaecJFpnHBONhWgV28Ddr3iFb6JO9AVXAqoVMEpWawbjdccJpm3R0PSjOzztfkiFmixPI+ilvi
VPaOQW344XR2vR9atU0NB7FTCZ3jVpcq8NujEOGGm2dKhtNFxjtlLDh54JJoOuEdF1XrQjTNeuPg
vECCC4moCWqaNJreJK3MXW+3Be4W3Z3rmFtnGAX8upWyiDxWEOruK0IxzcikZlBJ51xMZV4z6EyN
Oaq1yCGNglrM5mEvP7P8hJGI9eL/Wi/sztg5fAqFKRXksK4VDYEblZNc2MOqykie/4rEJLAAgE05
TzFfS+Q6DoPH27WuQzwf23NJsbA0VFNrFNtcGYs/WQ5wXmhrx+vAm/tvMjljOieb8SYFzWwiFH08
FDI68cxBGp7xkVQFaZV+0lK+8WivFwmkcimsa/IC5T1+OJ/QaJB7M1WWfUO37rBOALWRcazCZIOZ
15NxdtFno8MWlcxLlvvfEdInx8ZwQX1FVOBSmxVWPxxA+vljth7TPzk15bwX1l6cu0SI4/DxOKPl
tUw+sqixhzx8NTRe/3juZ5112Xp6X9I1AXslhMR1q+x3A8nJrMoijRkDLZpO2gj2pcyQHnePRo89
ifQzb7JpHQoZUsZzudsaPZIL0Izld0QpA7WXzOman2kZPc17tjtJs7saqLR+Bx/+rSIz05J/Sekx
TOymE7pnw8+cWzoXkJjp+CjlhoPCcIvzLXvS3k84Tp3060f+kAUMcNAG9t+/mPvmkqT2tQj4DUYk
B7wVN1WQm6mMZbtbXAiSP35KVOeAU1eed0eWS9Q0gAmDCOeYtv7rzUFZalZuDK7WbdQM7IWNAgpH
sKr1Mgef/EBxj0XVCncMR1hdsAHXzgaNvFHPPuJ6nvcM082AJD/RvVO+9xLNi2X71PBKD86NEEyC
WdGYH1ftToAdPMxTvzXqZJcr2KJG7iZNiIEoH5fPMq6+m3rk8cbSXhoxW+uYlO6ygeHP+6A78tqG
H/a/fyd1LU9Xg0Mp/Do6Ze8dCDnaPq7Hxjbqq22UheXcsgkO8CJyJDUm5HvHb+TG56JIo7PXARy/
aowZkN9gduArkB/YfYjbauwlH+eJEaq4eBvdu8ZTCLFb/k8tsRLFDkVAxnY8bi3z6RVX4R1VPgxC
r/eJrdH6ZsYWU2bF8GlYSiH8d0+QhxP37LjFnm9SyqAEOCAtu4i1QBMD6p9TbFVa9OMACVlgH60B
lNUKN/cd726V2GcXGahOoSyI6zAxpgi2T/fr3I+/0yBU8D8N76n/ckTyfoyJjjhZVtTP/hc99x69
RGec+XN5EAuCD5f4gdvwikSQ5SOCx0os0FTAayL+g/1FDA963AsD/bn5khcy1ob2CXUa9UuKOQgP
/FHerY2dF5ZZiJ2BBV4mrXauQ+r78gqeeSJ25qO6Ac+GhTXH5rM/E+OssCGPpPQjsmMx8UDd4APa
GlEGPPrVahZMxbLwVXn8RJUTBjvALUNJkG4CoPgcAfqJh/wchFH24D8Fl2cMJDtki2M7ztzRaIm2
yx1288R4fkenR48xZm3yDb2dEaN3Oirq1cC4tAAQukNlojtxwih39O2Yy955nGIZEAg+uN5GXW2G
WS2y9asw6+wqQjXBglHYtI3SvCqQMrDpoYVNIFOrJzJumpM8xBFqLL22iRWgGoADrs4eUdFmbDUX
RO+j5f1D6SgvB6jQY7YPuTBqpXB7DluM5r1KfU2AVsCGh/Y51jjz1adJFl8ja0jvFxBImwaUwfIA
A9qzKnXDHz5vMYO+xnL/uUsGG+eW9jomFK0U9Fd/1lJ6+4H8O7doDPnd0RgOHktvPL+3txzyCwq6
/DuMGmnBPhLi157gJy8XGo46tJ2wPHfm8jK7/FH4ZSY6NaV76/sRUyzXJxbe+nDZon5P2KJdAFV+
YAXI6fq4KLdsO+mgaqQ85U6GEDr0uEcrTNJkBys53bO6zPBAbBQm86LfrZoOoJSNekTOWwUdchjL
IuD3XeNSUKevoKKDLcI0pFaY3m9uK8LMfFx9fPI0GI3RQfcq8jP8o2TUOP+UgsmXRgAkA/wcH2iP
4og+5aMfQhlkmb0GqHjR1n1K1t61LlPBYRdAAtzstXJMB/dp+1XZB4l9ZEdDfj/I2MHt422pZbC5
BRQSoO38HVl5nAr193TFxZG+IQMBZ4VHUHauuFQjOVZkFa19LP4PLcJWAcDgd5kZCVKz0x4AWCqR
q1hH1CJ+xT/Kj51EvPK1/BPSETUsYz6pLNFSKXgt1VHoDOnBIHKlPbUBbwd07Vz8EZVJmtW20Lt8
W84ETTjJ2iae0mczqBT9qo1xgEIy7lUf7qs0NKXQiUhLd65JCcAIl5/LeAf2PwpyGcJRSI0dyQWu
IqMrpYMYAbbFx6jhAD+OftVwUuO5I499Z/3GhH3CneMfrE/lZzE3DR/VK7kE4s0JFMdnUOCeFgKZ
v+wrd5hAZmBKyou8mPvbioDeKv/u1GGHp78ItSIi/Es/BJmI6mPMgzvf46zhaL6Ucx9sa1PciEDn
Fc1b+h0+GT+035s1Oi6Exx1Ku9UMzoGeCsYagKKRmWwzuE+boMwpRuzvnvK07H9JFPw7du/+Iz1l
h3bHUdw6F4O+tueMjQHtF0XBZuClOFV1NZ3W5FhlkcejRa4wg1HTulvqjH3EToXtmImWcV3FqQNg
UyUL0vzP3ovCu5m4fmxc4RaczMJZiDG7QpABHcALmHzyCPYRhB0r4+ORFOaG6EoRQjrhSyahEJvk
/C9CMDYYM3sXlAF2A7kfpPsZi4qsODp5GkCAbX6yv8dZV1n1P0nxtjLE43uZSsSpJ2wWRaqosqDV
0Fd4ncvaGKkluHewRjuvL9VrRXuPMCGwnV4sBUTXakk4oUHPhvm7+FwcG5S9hSpjjXPrb6L0UdcP
GGkPSQ4m+qICMXTLBKBIRGBQpDHwA7VpyOMuhr3kD+e5UJ183J3ArXL0Ol5OzDFWTvlIs1jzchOl
64Lmw1o8cwUfhGWxdoNjQarbfQQpmtu1cct0Lq6yzQ8bYnVoCXjA9JYX9fNUjhlSSVYvmipefwni
Ps0FT4LnBL1CrFLQzqebQOxUiUE22Ny6ZirlT2DoYEqpYkthf2roUUjubA6OHJieGcwWAefI2dOc
zqZoLDw9ONKCGbTok3Z/otvuekzqKR4aQ8gFHryOJ/bmP0C8SMmTQYEI1v4RMv1dV60Y36A9cmhI
GICWDWFF7C2ZZGse+PxWazNaex/OQA8g1uS6+ngb9HJe4YdKQfV0EYjBjyvE6uF7nh83ygKrxeuT
UMVqgpm6iQ6T5s0S6oi/GKlLX2weSBX/Gq1EJLJdqGCujCMWk93CcSzO+s24gIP2UwVRY7ibwDK0
c+d736qBYfB2+8tN2/Cb/lHJ6KnCmk7JKWWSWSHUTleJ8AX2ERrrHg0DvL59d6r7UE36PWeL9mdw
Bm5Cy1PmvWJ6sikkWupifw9LIVadttdTpzVsxL/5f4fpb/DNoPuNEbV8yURp10lCtBjEWncYeHbc
PLPUtshK1Qv+8Rn5fMxwsTQ9faKhx9rtAT2W/IY4nQCWr4DFUJtJZLZYUazRAgHk9hB7jfBwpdYR
Xq8oXyyDmGucnAP7EfukVeDyw9d028oq16hog7T24VusKPyoYQgs3WYm7EFwkHDJG+IAvbCrN0/M
zQOdrXCYxDGeeTmwu2s4JyqDyX4Deq4rMULJutjmaXdWz4H+8YcdMwpaVq25DlMulVltGliLSU79
08SsGeKYLdOQJbqo1+yLeQWwS/eAZJqVTExISwEqMJom5R84Qo/ezFDFuH8PxuSZyDrTvxXF0ju1
IGF1C5h4U/cdZ//+Cvo+oF+4NnFLyhacdkJTw005P1tp6HJG2xxz3lIBOZWz+v6OWT5wcOgBPE9B
/zJjAmDez0FL04ltPuW0qXcsXGyWaurdPs8ht0R0n4Zn9S3NUEeF2dGHgOKLUWUGkmp2MH/JPjoa
6pJTHvKJnAmrQ/zGnYYWGN8AUlVzR3sm96kV3saVOH/qmqCH1vEt0wczKLQBlBEidsYpu8q9KByI
9RCuNwHN6mchJy0dFT4puVwKJ5NFHo+tGcNf551/lzwLxVCrDO5cmWtN2rKwc4hJ9o7ViWDJPQdf
Kx5IjhUQ3ZrEz158P2DO4W5TESdV2f45hruxcecnubO2VrQPGI6dUvOS8NmrbtZYBwRGx3jFJG7w
sBNdSoyEOMwmEuSnxbCIbFzYLn/2WOLW9cPMOflYh3D7hLUHS4oKY5CJh1EIML42qh3BOx7629Cl
suCxBtHFJc1pX8+fMaGe36NvMhuoQEeeZf6wdG3niNDX/RUbR69ZDBqobDKrz6de1orUZtf2dK/J
kDNHa601wVwBR4H44atV+knQ4efViyyc9cXlAG2JWZT3reG+AlO9ZafUSmWdsQZ0x7JPwTm411bT
VzTu+EsSqgrYBqJQ9/WGcngbI65YnLxcm5DRCfSOMXzXCd5LGEDDjVID/qcnE44oNH7KNyd82waW
4CbtPR2K/CO25wlyywCRXiVrc3Axfzo8gCC2ycK7fyofI6GqffTP5is62hje5uBjNLUYhaD2W9eB
h1c6TOFTNB57jjjGG18ok0VcDRY0ZSHO299qjPDwLR83gLGlf8Agd7U+SSmnjzPiEJrlVpQcRlF+
ZfDQ1/GM0PcakDZbimSsyix7Me0lsgScWMqElBy97QLA+9uZ/V5S1bvy/lC73IT0noOoCJNj7VEn
an6a65uS72ypzoyn52fV5mH91mX5LdZYNoAo6x+89Lg/f9CHyvgs3cnY6Mb300EjU2IL1g/irD/4
hPvTIshHj6VhlAhC/jTlBZXP0t4x6lIKoHySpKafs35EdtiUT28dRYMNaRUgO9uysa6ejbrWkR1b
T3gzkmtw+MxhzQoqjoIXU/kdZ3H5F3i9+Oc4OXz3q32kCHHFTARQNqvGMlBAwm/BVvqzHBeLuPBP
IOklLIkRx5dTYWyltShn4uY0buS8EZcwKVHeE4w3RdM+kKGiq8rz96d6soaQ/pa6tIiUkvYXkv0P
N1OkI7eNqAvteTn6mLaT8KC+m6pv00XR10vI6A5kS7nVmuppwH5LLlljAz2DZN4jTq10ghWLjuL7
Fv8NJbiCUrY/fi4NC+dKW7T+w6VdHUdtdciaJZsye7RxZzZc5qfrQXicd/NXiAylgezFXGaO3l6o
ZALfyjdYMlxjGls//Rf9SAWvDxSbi1I24Y3en7B8l9fQ6buBc3Wl00GgpYmR2KdwdLAPJQfaGrRE
7tWOa55moKpT+jRRqgZkXQbXjrmQlKUo2M6l3H6bPIc/edb8LGg0ad23gjxfW8O46kC8+bixtCid
/+4PiiN12FkEW/TVt/3IfwZVv8Ci8BlZTEkrR7pAeB6IYquDzbrbvalP2+WcA9vFLKMFDMJV2MOW
fKe731bz26l6jaCrFAfDr4CKfwbHT8tPDuIAJIUZKd9tOQuL6ENi/Po5z/jgLiLMPjY0CcXDUtuJ
EcRqLBWDW0LpBzSbFRSJ2tYAlWWr7Wrl/ppeEQAqG/zrxlZFcUhNX5EgSgaeYgLIvuktY922xlVB
E/NrFNkfBryzNhIG5quAB7TZyr3NjS1vh6T3wmHKHojQ9Qu/vExA3pJtN7D06K21dqJ6uFC90fgz
4qyF9hMXt2+ragVJt54m3X7KZjE5MXSXtU6kw7EmeiujdviWpwb/+XMMnt2Xf5pP55mx9GDdiA6u
WOhv4XDTY4+JaxC7PIGum+5I92XrZLPgOrYZDNsiZR/mL1g+X10V+5VeoKe9/8DYA5kvssQDfK+w
KnhB9NJ7kzvLAo3CfGvTQj2KKrpZSTGKH3GD0QEIvta/mosIwIU3IQxhG+Ko8zSvowJfMQKPAsVW
Hu8mgHeF+y5ZBpr9BKaqv2CRiiFVrgZB8rZ0iKCThldYbp/PggR0vfyY2PMD2WV6ReA8QIYpWn7q
M8c3xAf/YAa6xEctguMQAToZ3kh4bcfg8OK2QGyhnSzzOIMeyiHFf1r+09nZfV6lpp9lRpjcBDWG
p+F3z45XIJvFNuX4SiAybIqxrIY1Gd/WEeSZFHzo7ly7QzCKclRLATLSJaCt4eOemrWOeXbeO4BJ
3CkUUc9G0HPfixVv4k7rg4yV0qXH05Qq7JnCYkry1b/5Bno9VUKAYC60H6oYNHbUwlp3Nx/FToWs
HLt3ZOeZo4Vp8LACiJ7fioDm4Q3WRuGLL567vWH2Yy1MYCueHPyQiZE99l4Abwjl6Nri8R4iybxT
Of3KKuROjsLE5YJZ+par/Ob+mRH6Ae9LInid9J17o3o1++6YauVF+2G6ufP4I++yz/IPyp70gBNT
YYrDKiJVWLQs+YoZ4SEBik85m/Yj731geWLyGng95ujJ/w/y+IumYc0zYSlR1uveteNunzI+Nwc9
DR5zBS9zcbAJfI/D5ErpIAsssGlu3FlCPEQ7/VZPgfiRkWDu7hxtDhIGqTiFMfFPD6y2HZzLOtoM
fK9w6s187Ef1clJL8p9aehj3uBuKH47nHSw4b3Re2Q7kzVdsAN5JmEkHhji+mmaUKDkDhxQeR21O
wqF1eKYE6Y0grbPSTYaVlWLzmo3OrAEVTWpKNuMprMnggDsjc0uvaIxWFD+1pRtD9Bh6tXkQsA9g
wZa1L8LY87Yww840bMldSiept1y544sYHJPpH0FepWcpsRMl+pIo5PbtwdYOZL2PmWQsEOjnJMqG
CVfdRNhs9cgiJSyE4Y7mlSNz8U7Y13lRbto6vyLhfhYC5sPqU70/B7hLL5EDGaFhgYBtBV/797Bo
TMXHPlEqB1m8UAB3q6mvD/3MVse0+E6bzu2Eyv5FA6Bu5aFu11DV/Rv3J1lVs7l8m2pGSMiCwLUc
5WOIpbMigBO86yXZjvaC6rBj/bmKGwOyZI0Gr/9P2lc3mAoMXC5iSNfT6NMQ0PoImT97CCWTPkyL
rxYGXV2FRD2fW70kTlsmE4ZBZXpmwmPEKVtFGzDMtpSBHhR5pj33ISS/6cOtdksKyTqwV0qZ/SsU
SAKU7oW73uEas/9c3LkCF7D0WjUOc+8aX1H4VgTEv9vUImGzpIBQf1KM0m5LFITldjtwwwKDDEFH
XLA0XzVm7Ib8J3vR1nteCa7FwntsJbbez1ZvfDpPRQb5wNm9RLkep85WIf3WxKpyC+hdcuXRcl6H
fSL7DADXyF6Nxh1JTCjb+gEnB+Bilr88detM+3MMkzPP5IR4Z2Ox/z64EAopeK3Fl8uT8YSCDpCL
sl27pKF5JKe3vnspsVpU/zm4fwHOlCYgXHvUmWMXvct/DLH8oSjkL8RyQEPPB+7kMt5ya3I2cshO
41VK8Cl6jOjHIni3lgKgPoCzAuQ+4c1p5q4j3MStnMIJsrAI4thlRZH4NVx6QJfNmWpZJsEhdv+c
IZcfpzpuABuSs4QQSsLgycZYG4U9RkedS1Ey/47FiiuvQkdKPnt9B7vqVECC5aVcS8pWsehKVYIK
xqRFOvNgDZXPbWfuUXgb3TiXjwl9f6dSWgOKMsbMTIl05EcQrqdn5I9ZCYSTDwUexPR0dmQn/jAj
XZahJ+Uvug25EFASO7n0C1AkiB9u70l6Qw6CEnrrMtdnH8J2mtVuA7AAnspRly2U2p+1h0napcS/
TMq9Cr8+TI1lhznSgGhzUcWHE+ZdmK7qcUwJDiYoR7sgPjiD5OzjzRcwHNRNp3LDZ7xC7tJT+0qG
tgt7GeL4GT491Ez3BRlJ49bsOMqUE6PEy6YDsfGmCoNaYy6vqb2gcX1rgh0qn4P3KX5tJ4nAsqW7
tFVIzNFNp8USDXJIPrExAjiJ1WvBo69Gc7LV1dcM+wv057Oswm0lsbWMYcAoN4+WI5wmFU7kiPiS
62aCQznQ5XC5zxYOcoeuT7Pr0/pP37nbrC6UZQJggso7zHzK796krRfpo2V0gfzMjkCsxpx3oBDN
boz2i817gxVyygHrF+JzwEyumJASLvVf8AluLB+cF4L1EmUFsSY95qLFYAbHbHH1h4oy02wfJ31I
b4gnyODhNbUrKfmVRASkjutus4K2FScJiPpOlNwqJkHCArYDsmNXOIA2qZRECHKQcUozTjruOTx8
LVo8IuWF4vkQV59F3ghg/GAIglBxNo8h9UFmzIPK4oLkYsmhcEE33Jc2qN2FhQlTjoEFjLcdiWSn
m+T7zumFfCifd2jkfl+IL4+1EYWIvD0OQnnnQashEgNhQLHdcpRiRF4Iw/RB22oWV/2gjr16rMtL
mjTqdtl/03MQfvwlWY+74Zq3uRUPQn/SU7bBl1T/nr5ffTJJYNJ4J0Nsz72zSVf0oKrZ3LMCylGY
bBYRO89A/klZ0IzNECg38fv4ssFfltsdX9Pj77IAo9HO+dDlWwuU9gzJZ0rqO80RCy2pZhk8Gtpy
tqXc9QikqEUc1FFmDvl+RQ5mcfliZsz1dNJO42TbZbNydyiUIndWI8C9VIwFeI7wJchxKI0aOdYU
MlZiHgvvJxgZE+03rCeuAXwpVXchR4d5VXkELYwlA6zmb/Gs4c2A6ifFWgcpKWJoITre5JXtwU21
GP+KkEKmKdCiJbur1kVi4rjQ7TyCrbawvS2AeRwLkHFYmedhAL/waQihEnTWd3vD/x0jwM5Lk4wR
kmRsXF0LW5y6CjgSazhMNk5Zz0izXUDkUwAoC62kbfuJqmm/wExXpWI0qaaPkXECoClKr1rHtV+A
f37SOSme5vEZHMwBGghPrKSQ2EK8YL3w8B1mVxA4fBbwlfdpzOszgBUGKJFc/4WEmHL3Dwo/ADHf
3BTVIClsAxTqfjaJlQeAItE90Oqud+icgP/JFHcKd0Mfmgy58rpr67Ijn2JXp/UUUhHHPdD+2tlL
dM+GUNB2aHsOMio98SMdCfwzaoA96HN+WXZnkbHGLRdSwxhbCZfnH3B2zYLmJHMu8nucs8luMTLE
RR+qTeeNCQWWTS3SVnrgTA5tU2HAypPFmZll/TgjrKHosLjIXjTSOlngQic2xRIOjv8Z7XPa3fsy
fLBRJg2rx70kGraxwe20vODY0pGmw068th9AxifWyd9ddI3/GVD0Dir85PtyhZCHIBW36DhJYoqx
V4CdGE+3Zgt8OEZNOET7YAeNVwDw1RxbbaTdEH4mo2R/Is12R+CPf6s+lC8lRxSq0Q4O7Ntx0hQS
U9LfMu07c+504m0eu3l5nR+YBP5riFWLfFZpymWAZlqdkGUmgTkp5S10R/pIRjfO2UtSzusctiag
ToKqo9QvzNw3Uce7A7Cx38CC5UsIbvwicokRUf6Z8GK1HflfGaYgijWGcYxQkk0eVsDdrSV6Jvs3
XO9CRwG192IJIff10ArV44vgWs5nK5TJ95Hr97Ne6yNYU9aOEhYYDQguW3oXxvSzAApW90cdUfHG
OVrRV1hze9bjFCyXWTeBB57Gy9JZlsOst7wLezICBCYHVw/h9u82EhYTYEJ9je5oT8ZUJ6idlI26
7Fnlhz9o4/oyo2cKkuho52tdciqBCuFXxk5wOnZqaJ0FN72aBqt7iGnEiYxgcgDT6FMpeDxlZUFo
DEOEDEvVaXWGmi8a7LGavjru8sMoVW3hGkOzIcibIeDyPTPvGpk+sUT0+NWi5KT94A0yEw63FYc9
0ij7wbYd0bLtDgFtrFAvtISzxDQPGyzOj1QU/lj+LmLorNWsvBh+sNUaKXaoa/sKKP0bnpJ1DAuQ
AWK2UYo2Jx9LWlZ40+QNPdcBLv11tQQuKqPWKK9DxPJ8fEp044K6BMKxvPzdfcq/zFvJS6tCUj+O
nurHc3OAa3TvAyTXMgUKpFWBWk3b7zyI7aasT5WbNDPJt62Yx++CozS/7mbCnAcv3sYyuw9m6+EF
xY2B8IM5ns2lYTP+ElvXoEuG4JcTmP9mOBIb3llcOGXYg9CqQ+1fow9OyiHB2hFq7HCIRnGwkgrd
YL+ni6YQ0WxYpum6FKLWvIuM0Yi3rhEI/NaAwj4oZCwtqVpjJTWs+AcSK6ar2rqDQZIQ1nZ8k0bF
d+odwFL9p8KtQ0PD/0D0TRIuYTuPYlpATXZG3KDU2jrfapz8waOh8HR5OG/TH4J7JdFrnWlEvkUw
029zHc3GvWedkbXTi+cNQSIzQSgYz6uIgKSwnVCOG8nxoxImMa7S5QisGqLwMsEwK1FNNHv2oOVK
ZT3RS5qlTIwRy4pYXpGrIAtysK0mHd7xQVbuVB9RWHjJYPDfP2Lt1rgoHYnG7UOZ4PKog5T8Hf91
YRgtVZu1t0hunHpOsUb7NolrmAfZGqjLpKnJpUGuY/mcHs0iT9DruBdqR3SJh/NxonhjgfTs550+
rASedrb8GElEhI9JW3Ff7FXJdjF8zJMzVAuWY8mx4CRfeXADGCjhywBef5N++jM9TIAOPHDfacel
BE2eDGOEV9+1BE/VnTV7lfWWtHZ8lCjc/cniLcXOOc4hnaYHqTkiErzwa4uUe3akSoc4CpyB0i47
wpyOGRlRGqfNV0QRSgrQk9YOAoQ6WHY/2vGqTjlXXEgBqwtALi4adpCmdzY0WuUvL5/2fAdWkCXo
IdkFGExQ+5U91I2JxiUa8gB0gRhHxO9G7c4huWasjXjxqgMS+JQFD6/KJ/vC+MEXyQeuTfd1uLbV
8dbBVsu+3XLU6dA/HsUEL5TtXweBtyiqihU+o5Q8r0qpQy7q/gHo3AsccACEIcx6fV+I81fRVHR7
Va6fDdokMgGSENP9jmRVWMd6Jcij2prfMZpQxZmagFhfXqm41qoDkHWuBzVzbKITKKWtD5nw3OOc
y5DtaY3cMCHYwSJDeuujQGoZ5tSCj8X7RRQUWtrKHl4MejcFtaqiDMu8GY8Zfic/BrMlW/kVhPmf
4PGGJSdOJaZbAvLShDaCeagg1lPZ/ilIXXao8VdIxoTTec6lrIzBzRB/yoXMdXE0XCQ0Uz9UKVmY
6oIn3yOOGmBU5YPMq5RVU6A2xJdf76zThdPXm6rbPrGTDugpHpOqOyZh+cjAT/L7jkA2bMVv10wO
u0R8oRRc1kuB1/N9k4dqlWZGVgJGExdIrNYDDKSK1otsAWaX90acT6mFOshES2+e3ncLao6US/D4
x9uUvQItrMAwFcHGY7Pvfw3z8MIXBpjo2dKzFNYLVVrBxPvQ2amYxYaRetv7OTHwD0BBgqPXQCq/
GzOIQQc8pkFLS1FR87ECq7jw0h2XLS9ArrXqnUNTtcwT2Jyrrog4P29G/KtAJp2P15dDje7z5kdF
o0zSpMtx5zhyjA694ewTYrYXCop5q5Zlcju03SmmPRVHhbI0z0iX6cQM60/Bo3sGG1zfvgNehf2W
4Ba6qtrJmXVbzPf5yYDQzGpygL5Uiw1XrWMU2abU6tqWmNlFzejwnQe6uERvHRJ/OaesTmSGCtQe
kHR1IjLd2cO7/Xtc8dXG50OyyL7ug8WzddhUjMVqMjDYBvID62Yc7+cfo+NKPyCjyZXy2tOECTll
ve0ATbne4otiAVKg+VBu4bxKEHBDcAB4BsHmKUKzM1YD4le7ZA/T1sRV6TWDLzjKaLCfRStyA1S3
xlckAj3CnqspTl65Rp8N7m1dMSMvTextsrFsX5AP/sYpC1l/rxfZpaYlWOD2o7iKNydkOkEyBwIC
JUAx1anICmTAgLvE+PwMG7WDrjmLhVgCLoaPDtCGQo/miGnJZA40D/0rws2qZqMpw6p2mqOD8BkK
JO0lgfwDuRyJ/TMgl8eTjAuRcqdm0vTjggWUsZuID4zBwSmbr2Tan+I96YwYMruRSg2sTTZ734cX
L1ZJn0PPCQUvm6WfySZkNttlzj/ucwIxsRVpZ+bTyHx//0v+Z2gZ5Tq1S6ww5yPxnXMKN4KsvbAC
/bejT9ECFOw8nja6TWtojxmPRJlSUNb/XcXjniI3akiClGP3VgZ8ib0iCl176DvlR3B192qqQ5zY
SlDhBvRfCdKv8Sbu1guRL3YRl7hj85M9zljNZLvVzFoEs8MUE5BDmm7iUnQf5/XLOcB3AquiOmyf
DrPDSVMzd+FkZ6eevV9pLFafZG2w69h+b4umONHVSTanwNzuyGcTKTX1gTfvCdgVlhquGlY7FMdT
CiNO0pMCN5gyWy4hZ0rPJcQjwxQIlEKrEUcuFAjxYcD0G1u8seLI8dN9RkfzK69oT0BHkNL8FiRb
DE24cRcOE7Q90tdynyoh0LUAljKTN0/pRH8lcuNpAgjrh2vSjgm8cxSkeXSX0rVeUFKdMCKANlao
9LJtOPqtQKXJabayl1uDfz6W1c1iRkUoJ3LsxE/8+6YhodlNCehuFP4sR+zv29TGgrtBAotCaL9i
NWhA4SBGumW28MMVV1yEbSXg4muSyL6mZ5iABAydLO5SbJPI0SKyxNcoaPUadOQ9GhVHxotAlr+t
CAXNuD/+OsbY13cD2TdTwcfCVeCV7LtzmBx50LtYW2UMlSe97dFypBOd6xfSQwDr0oT5bdHP2Wnk
/nUiO8ia8z+ihyw9BJqCJmFgWm+ME2nLy9LZ7w9cJs0j1JZ4+vq5kmdnuiOU/orAIsbqwBD29u3P
Rm8iAm3UVcQUZhBhn4FK+x1vpElCMdCjyCrfNMOK3Dq7HWgJydxWxTQvXhS7Tj4VTgGkxxDeG04E
7cv3SooM2T0b37NooS4heodMl6ssLtB/ei2xmNjT9ZdaA+R0adAas1QiSQNh0pz6JRAgQzLIVT68
NsHA8KI/uHp8w07WHPmLYVipMQI3aovKmGPVmwe5hLdBRNTi3SJigo7TAyaSOUty1TiP+plbkNbr
QO9wXpXZNpR6T4AK8mZpwoEM2DJgRisGsEM+ts0T+HarXRMmh0sewtaAaC5gNCj1dncL5c6C63I3
uf9HP3SBrb8oBxFPIJ4fcqBljbxKRO4od8yjPfnIMCrWlYx/gzI9JW8a8so6NdX1Ap4afIBs3vwk
/uUo3Q/bUfYFcWdNBj792/4+WAqJ5LVUG/ACcHMCJjWfUZSH+GrYYPyaqZtOyzPdY6Re5nHOjRbq
z0XdMwBcTznNP9XXHu9Ku7ZWYcEpKl1YGeb2nukR8qj1UsHXxBIwRjUuichnfX/bD0QTpHC6nXZN
Q+UTq+crSV/8y/lVB+H8PDKT0GT7SDhxawvoH+jpH+/grOrZAxwzjkQ+HRPkisjWw2d8r5+ZBPOb
Hma4F0nICyV4FDM49hCgUnZ7ASj6wvGrLjqgBEdAmfKcSFhrlKwHA4apUragZLY14AHYszV5Yk6Y
0L89KT4cOpYpF+WNCUrzI8hD11nrf7LoznSrdRMfKw+uOZjzNfJqKBZ/J6jXvkPREKxJd5J0Ax+e
l3xIhLP5yNI03FlZa0UUx+cIcHtV29HNj5d8+bvofiDDsHL8Y5Y/Ix1M5caHd/IWcKkfiPO2B/gv
ZfDKYi5CDZqQ/wxZeZGLirUsxV00i/wKBAnVQdoxWlgTTp3HinEOfg8FrKTyXXWu6cWxKZHVCETI
+wkDa21G98MSAugNAkFqqyxk6kP2OYvskOMEhHkcbHebpGIGGGzk+Uefvcbbc0WTcdkkK/RkNfuP
kD09w0jTcA08VOt2kSrFaDX1pBOk9/nOS1hBSaUHUf9M/BJL4KluLfbd0qASY9wJjUAWO1yTc7WT
Qk1DjnupWGxn4bc45qFiB+P9wcv9m4pdZeSmxJ64FdLw9InlQfMWOD8/AraWuaQUP/dTvJZIJBD8
VuhFqnUJyl47r7poS1DxDTwks7rdVWn64sVm967K7Nlwvl0ksFPj0LihFzX83fkxRdem91uCAAJK
OjTXtv07a8AV2FJs9ct1lHWGcSdn/do9X14jRXTIsGOWHPZjD/tVywTEC6RxzyfgtbDUoM4Nu8Ke
GaZt2Pp/SHeWdf0vqQq3ZyjCHrA864drh4VfueDVTBStOQ8cT5i7WbUyxn2iuUKX7zUlq+xBCont
EAIWoSXrV3NaaKVik04qvGMD5ZZbF3SkZeFgXRlR14eRORhEjpXFeXMhlnaNi4R2/5FbVJvsW/x2
TFDWJUDIaHWzOmHtxilUOZHBY/avi/1kf3YF+Jd2dSWPIYoVhWpWTSWSvJOXXwxovyovfx4qvw56
npCX51wiRCsTEFDi0Aa1orPxNbLzsFAgIA1WWbSp59sPciMT9I6l+2+yUBOx5JUSt+P6NtotkBZI
JBTQ8hjFizaWeLXy02MkWk6eeB5gKy/DM8KyGYOXnESXAPuu4nV7IkY/vTzRFsLVKq1PdgNacCVa
M/+YKtY8y6eMfVeVzpCYDTlNtG+VvIPmDMutLwhec46j/cpuRH8EFY+4XJrFGN4lr5Aml1R9UcTU
8dMvjlKRNkChlJVCMhjc6YPeeHqNmp1CXJH1SP5/oouiiQ1mhpaBq7YSvxj00cnfmWYFf/E+5oI1
z+pw+hQdl8CbETJe1lUw975/a2t3xx7rfrJG9Z5UX/r4V/wvt/DVNe68bnVEkOJVmJIvoO5gBGX7
w1qHJbzt7L38HDzxkRaAXBpLVnq/HHG1wbmNZt+lviG8BzrBjiP50ajJ294l1QLMJwdi4u8zaapM
7HtRyYt8UJIvJvorOMvSoubAN7i+l+ax5ox3zLEU4kVWk6ov07LM44/HndsQi/XDiFsa+jHJwWY5
cVievDmwb/WgR9Xkp0/G/C/1FZS5tBL2mn2pf7RN6VV8zaCf8HgV2/MRg70wTsAo9WMepvK3URD1
hCYJldezfdvgqkK4ebdO+AeMinBVd1SWcNWW98JYdq+HkEtBMTQRUBUhiYLxq5cflSG7xaES61rS
3mqNavsdqGi9hhVhnMaGWfxFDISjlL5d6KNgozag1WUsKxt4cHchXb37SzcvcdVukM8beaKH5hf4
m9rx7v6li5pfYZlbwkCXW+VOixl+aYyuxwKMfEZ3btKSDiytW2nlUTzjYsCfrudTbDxhFFKErzHS
bdfFVeEtwRufpMs1vUEXh48WG0nD3pdIu68DxGz1FZpwUDKWlcGj6AkzE5ACyfbk1ARC582KiO2F
wGvwMpwoQ6AfAgf2BWdJfDAE4p5fHKKjlME9xLzO09X03+CjQ3X9hkV5FR2cmPhmx/17WQSmhj2l
oQztSYnQ3ffJTp5lemeX2hM61HFQgZRcxKotV+MJHBGnkh2/yjYNo4o43rWXQqF80rhZxY6maxtc
71J3jHHHJjNSfuJAO3XN8j8x9kwFU3d6P+JnYPxmxD33u5k2YzZXTJq8cOpFz3Rdiu5Q1KHMvAxO
Kir8UbClrrvZDEQRMoR9okjM7AwBM3flqJpM07rJpts2s2MXwLhVIuQHe6HD/pex7HORTp14BmY7
kYSODbZ4VZY44cU5isKjlVRUPbVSjeBfB+JgddinHcKrSTvG7+L2+mobzFZxsfmesYg2xNxq0cxI
EmXjHKrMp04BpYdO2XxIOfmekB4lsN9BLjKH3o5ctxFpKJg9A2KDqbe4HLPWQXTdgCkZxhK93PRn
VRIQiYM+2Yhsd84sLO3aII8HPotfh1/hTIEyBb2mBCsaaacZgGKI0R8s5yXLdpIy128wTiaea/hd
/kxIfC4kk69vXXGy5jbDErVL/NePDjwPWLYt79uahTmlWBQ82bOLDoQFGQn7kZo/qKf+/R+QJv88
heSfLKYhLq8J9ZksbH70GCHEl88bl4NoEX94OGAW5izJvfS8g5IkGeBcfMSJdefeyskz1BxUkpc/
/Z5WlhWjD3gq7ayGRrxLgSg9EQmdVGGjt75iiUts5Fd8YttDybETOtiAnhrZQ1BKv5Qm8YsIu8cv
+9M0nxkHMWWfcehLfjNarANXlmIi6KMRcXzfoqz/zCqvzkJWHHr09OBOLZK/Jbnel+UVHKENNmK9
NNMAvBdxVoamatUZIa1h8tof7o5cr4+xdp+IA6KvtQZ92ODvSSsYjj3B5aq5f7Vxkw0dM+c5oS/w
m2kleUqz4R6UuxkL7+k0dsESR3V8OYkIZjl8ZODwNDnetqayKGnhkSGiqkY33MRFHqRLEX43SeK3
n/TyRiRqUqdDyYEIpAZ29GiZUGQ6u9xRuacVpa28MAHCU1SsHz8KAwFIFN3wvXwjm/nuzFr6ObGl
uO0AKjC3JU3pMQVPZpFUlfm/ERm+nw44xzLbjZCNMRJRWcAFxD45fc1oATuWgwLc3lbukUWiJIvK
EIbVLvcMrWDZxr1BREfwRemXhogsy3dCAY2wv9ApfbLWTQZKZRHFcSR6HJZP7Br//3RpOZQU0r5U
rGdQodsVokt+hK+jIKAVBXTh+c83RtNIgJ+1UuNlG6WTavFxZr0UUNkVTW7ycGtUbQfNHFjrLZ7Y
EzqCJ9FW4HUCmK69nDjo7Kaby/9HomgYbjh8HzFKuUGiiUOukdSHg9b0dcyzb1uOAFfk2N2QJm2D
o8CgOOTeB3Y7jo8nhwONDhgIRJJqaO1m6kmEpiH0H1DJ6nFoQ5gb7jS+EatlPRQrLw9Y4tXLd2lZ
kny1tx6YYeWLjOC3LF2q3sgQsplleXICKVWillUSGl4CAN/w8S55E7w0lrzg1UAQm6vvRXltA3KH
AeD7T26NzMPbQlMObbNCk9XFMZqsZ72P3CwSzl0PsLOzEjao/DjXARIPjvcA0GimRgndMw5DNW/4
Myar3T0/vyZOMhxTD1EevbPuhJDyGi+LzSUWxGWDiXjXNykVEB16GrXo2h1fpJivkpVh38VmFlcv
n0fAImeXraAraHTsMvKKGuJhTuUmmBc4KTgMar+4cHy0Tx4kl0afxdAQud9cTDJ9DAHwdlXrDBHC
WoUMx06AvtmZFt2djqT/vHLCj3hs3L/41KPyMMKwMzzzUXscx22cEle8vEkhhEA/4MfUAjEHqhoP
i/RlfJtQJZg8dQarqY5yfWqa0SnjvwYt749zi9KhDWJTlds4vw9WcGm3jzpLFX5FIawfymvzN8ga
ZmNHP3oIvbB0zhE9tYGYPTJmOFh56d4+AZQvZj7SwmB+nMtJvdx2zc/oBAy5wOmhS5ji+i9vsETJ
HeweD9gt/lSCnq9VFumZ5q+YrljFnzO5gKJwMkJm1rzDwER21N2sGQ/Yh0B8GVWel2RwH52G784r
ehmDptFfG5JyRnNX0A/dEfTP8uI8OKFLwQSe3WjnBvjPaJpUmkkYTteOGvILTra29uIEXEXA2R3a
LHwkra+BM0rk7nnc9KxdI5WECu+RWbbBj9veZlUOv4wjqqZiTWCsWScv/LjEFVjfCvnLoH+R8Iaq
LRRbXFu5tIcxS7IXlV2Ps2Bh/q9uvBSL264xw4b276wJsmJ/OhMKwS1kRcrRtmdkuLemGtcLPd8a
qbF5Ntddm+crD5YSZRjVCZp2enEHKislSshchNAVrBMiHyQ+aeWhBddK+NpX1TsTv/Ov3WATgTC3
a5w1+3TU1H+qxPprmcTpN5vmXe4OIVCszws+V+99dI9eYRMP3yxpTe7fa2RNKQ9+jmucB+jcL2nF
0r4roLdd0Bu/lkREbyGYtO6ilMSLIXGEYs1aQZE8ZV+e/hFlJBUnM1VZxOl+qif0YiXvE1eeAxUC
vxeBn4PjT/fgQZsSLu+bDtHmYSIalc3lasfZuhxBtISWJ/OneC9Kz+eLHtiyxbooVGXqVfSX+EJA
HBkL1FArP/lySXII+e4Y/2l9rApSdARI0asAidt11Es579Gqh6uV0rbx9uzH8/21/126B8m1tWde
WjcbzSl3Qs61/bizyAdBaq/tcYpZGbkdye6ih6kv7d9VWnTv0yQZfkn6QqIPPSC3IBYaj1BdCFmJ
Jq5iRP79lsEEn/vgXRnjQgsW/iTzC7sD+57mK6nkmAim2bUABTb4okNHNahR1h6OwCqgWiTOfgWc
Y69yvf5yBnWysmXCQ74X6wSxoJVefzCdi6R5NnRfoK65aNe6cPCDq/Q1+3Rao3WMG1jgqk/Hh05k
Gs6w2DXLbhxjvJ7KSc4/5jDizR+4E5BCJ37U8wwkZSPZZDuBz1591GSqvuG9ubhjdBFU7VSQEE5n
MEkpbnF0BsJKi8mJAK1KWlxsmoW5JgXU3ofzpehgIf3DAxLmvR/VKvf9yOuRz+AHAmeI26/47hdL
g9fz0WHmzht+cySnLmZYuHOuM9WlO+ZXdSL9eNub5qPKD86i5DbISEnwhbnQyaPAVdbeTvgO1bP4
m21uhl53fOSM8moqayxrYgeMXRoslJ9fP3dhfmywCRniCqYNnslcj+ZDFmj7y4m8XoaBbhoiWSez
/0pKAPl1WX/J6FKWfO5cJapa/ZK5a+uMF5vSSj78izEftFR7pOx/Xmkwr6+oFb7S2gx1w0avKlLJ
LswEJY75uREd8LwfcQczp2/N6a4OU9pTicTbzlElHYe72ccCdtZQvKinbCk4KEEIqzHfp3BqmzeF
TsuftjdsGffjDHOBi4aoCN/F9Gsx2qTMAr0WKPkMq7fMkD5HvdCf4LUbztLxQ6b15ep71b1tIWrA
EehxsjO69OhzlUo27Lhwcbc9HZ4C+S1gu/Fy1H2XaiX+kfVWoCkA9iz/1O8GsYhBJ0IeMeFm8h6r
pqXFIQJzQmiDXY/PI1146Qz35sOzQ+T+qAwzg5yk0B8LEmAH8ga2Je9OYwJX5F2VenMz39IiwM+8
Db9kuo4oGVXXcTJeYvXEbRYMGypopshQp8tldMh3T3RJtz4Bie3i/0XDp+YHELYONNaZiQZ7p9pq
5wrW7P7u1phfaprGjvlGPHQzMgVHUqJny7FgqrCtnhV8UtqNjLttuMmKhjZIf8cf1K56SiZo2+qj
exJT21x3M+spygZagBw5y/mPmFVdmA9K8VsZpClOG7CSCjzF39JWx/IqOArN/sIIXZip2M0KZEci
GXqxnqaQzI0Mco9STMDaadUMM/BTprDalFqseyZwYyj01upbyYnkc7yrV0Glnx4YBh9DNoUXFGTC
7Jg3hcpRceInBZhLVr4K2kkVeEM8EynFtQY5+5kJ1L+wa+DKuXJlcKPD1bSd24pgoUoT+tu19YxE
ndb635g2TqoZZ/fOpfG3wvz/RX6XYXytFS9/qq4FX2luKwnTUDr7UHUREypkq/sfyHWwt7FSICN6
SyOakblo2tqSkBgZI9rve9EHOeY4/lr0Nar+ZW4GXi5OYemurU0OnSckOscjTL0qG+3ojz5Pv+en
3OcJCotTTcx+ONHNS7M3wUAPUjpd49HihALMLZMXSK5qnZxGnzN7K5kfftigfiTJzwzDucycDa3A
1E3OrVH8XqeTZmFq69X3z+i0R/ALw4p9NYLStriTl8oQA6Ny+CqPPnN7OTInJjTg/q+VTSLhae/N
WD/Iu2tn8LAQfdvXAuxGPomXsEtXxj/6JddCJSqHvnOTM3NnKWiKjzhY56/9tOT24TgWRLhm/Nq1
zdXGNp6e8/WL/kbf2oSFeZgb1VxX4Xe4GPZfpHGhnM2aeD+qKiqMpk2MVsiyopdyocHsIui/U3Ph
JVOhEt7ollV+jL0YoN6L0uVwedULhiSo8/Rc5J8yHG+zPtc8PayxduDAPS9iLTOlx7hvIoQ27emY
EaGySb0w/6nHW3/ijvpA7zDk/21xRsxwIl5/KRUHevTbKGghHrWqbnVg3asHOUp9FXfPKPsQ//9o
sQxleidAv4A9BR5xF9d50wl0/84RodBunDh3JdBuYZhntpv9cPm8UglwkPRRgrtEE9o3pBzORgUY
YPbeqUS6oboHoJdGcnXDWHyWfe8DyMOugKkC0yHP5dJqXI44zkqom6o5b7DZzkCyHnRZeqCqF6C1
2u+YErit/wnriS8NzLNMC68n7QfFUN3C+so7pwr1g5cCaq9jJMyeBrEpzhcu5WipY2Vya3m8nlGC
SkSyaMuaZS7EGHpA7CHyjVR9gvFZKAnuNXnEvTGHuu0/tvoBi/7TFmpPeSKOdj9kxlwHmSPGNZ7h
rYzhElaghw2vFjV5TxtUKcgmgF/lt1IKTI5cPkXXMADjOYjhY7sYf7NgsH8sOHYGLUhHRdqsV2F3
BS8+QKLC+QRhwqok2fGy4y7fo419d9Cul33O7urIYIj82yy7M0TwRY7XbtDhLiw+BOLNq2ciqeKt
OYY3ysQSSIQJ37HvXJ5425e075q/Mo0t8GTAIQ5wGwp1E7PtPkSQtcYCfLF63OOZQWrjAEei23rN
qmjnyCV3DXq4ee3ySG5qudxgdNTd9TTAGhiHFFUMW9u7Y/d2Ei5Nsnhft2N8qsIm/XkSpoZ4QPSJ
rooLNF5qX9CDzRc4owx1ifd8sJAdu3dWFBmPavNRg+ap+ETOvLCLoUTMrdoY9MKiePfAyy+FniL4
g2rktyXum7UWzXxIJ0SihzgnAxZ9/S1DbXdt9FaL+lg2m7v4vXuZRQqbXXYu88rkXdnz6bi+OTZM
ISxL9jJnkqZ/HRDiorJM3E+/cdmLqixJri3M4srfzblUbQjkNTznSrT37+safvsi30CyohaGckCv
TK6ypEvMPHqfHxW6CBxoEhBjN4tbHsoBY9pq8SHNb1Tjqe1TXgaSrGlqCOvQnHvmmdzNoHvEdBdS
qkvGHk/AM2yxO5fPsr17SFzG1cMSRY2myGMp+J+B73wH1W1KH2xboyOLT3FcGAQoLKC2YLr3F90W
rLm3LmIYzrUh5Z3pHHU7UuqkXShXr+L/R/PtM7W+1adn5d8td6kvjulcZ9Nr1CLY/9GhJGzdDXQa
PgKqI4glG4ljp4IfLZwl1cT1nyYbyfogH+BDKqbfxDhWTGWjyHppLqksElNLhAIXDG6W8bJ65a4R
vCdYa+yJXpI+XKLD7uak2KTeHVmFKtChka7jhVSHHhT7XYrlvp0dM7aBpT2HdHX1ZTNLtYF7R+sN
xbLg93HvUB4BKSHmo1SksSbtJJFZ3aXgVI13Xog1IG9L1KNfkidfz1cQO9CPg3lhMuxkLThxYIKD
dcT6BMBdNdI8ZFacXINOxDvZPfls8P7Ug4wvNDGWap9ewzM9Q5TODI30RLhT6RytgyzgXLw/FWbb
nwI3IHmQlq4RUxJAyAiCfZl7qw92uap0pPsMSKL+k2xNBOiO9bRuXua3zTe1ZtlcSoDhnhv0hT+L
K+GT5Bf2WzWSi7A2l7nug8VmFyhv0r3OkFa6V5NL7Sd42ta3CPVk3nWWoZ2tTI5W7YnpNeONeLGf
ocBo7MgdW6ug0YKUk9daPRTONJNjLSQFUjVz6b+Ufp/wedI6GmBn95hPVKcQTZeTkkjHHs54NSbM
RgNF1nyVfiaZFmBFc+aPQrZY4HwzKgzK81YlAhKq08524+Zj5pbeEkIm8neciZffgZ9jvgxsh7TM
jy5KdzKugCVjiqFWOl9Jv5tzIZIf7hQNbEiowhtqb9Q6/7eL0Ttj/tVCJ+dG6ybKBC5c7m6/6zzX
yChB0ISsp9veiYilEVNgDLe2ZaF7TCnsXCUcpb36IXyObe+26qDUCQrdWOexaEUiqUFiS7pYloIr
chBTmDfTstqw5Bykrmch0wlAXWN+HGMn36udqciBf0UfR7x4FM7S9U6SvRRBpOkheSmErdSWBGnQ
o0/STNNPb1TFu9sZK50D8+e/m/B9pcfxcWFF4PWYGbcRNeOXQUwskB2/9l8V3BPG0EGBFjAD+8FT
p2QkTJEttesp6putkrCv5jKnud9W+Ca5LxaIYVgo7asNB6MZHkez0b56QOAuRFl8OISoYw8pfKkX
aIfjsGboQYbtgMRMwu8+CSwRhA/aeZVU5y8GaXm3yaTPqa4UFNijKqjr828Q4tLOjVs+lwZwhOeL
o94YCEIuG406uX3shv92CPOkuqT17ASppJctAR9B66h93TSL5izdRSiAXbECT6EnoFawcpP/Xn4m
Jk9+wv1jZg7aECiXYbTQTolZ1Ak+1Gn7yNxby8nOOUxaLutRwjuuoskGgv/Z8tfkfbnRrQ+3fSnr
WhTGaRjwNW9H7bcEL8kZ8yRJvEud4Ma5y1CpMcq4TFvnRB1OT2FrrSipv92L/sSng003GX87bmEY
H+FgfhcqQJDgS7Eo+FGXM5hO3mYBreIcMHVsdVS6N8RSXTXZsvkP+GPWutWDvHT6ggSijJyB5w7o
3Ef6eNYRwVb1KFEfRXpvYPhYkw0J4MaNcl5RTF7g439CIdoxMS7IPiOftqX2SdOSwISjIFcZQlVj
ya0UaTRFq2Fl4Nmj6KoP/YHGt4+sEl/eO789NBJPTu/9uE6gV9I40+RI30cseCJAjL5CB1+KkoJY
OWYYTMICS+xQuCw97h5U2TsKvHHM9zpvM42zRXoVcqAfjEdb+1ejoNs0OOV5TK8BajV2ZDhNENkG
41lfv1WQxg8GBZ7yp2dj9tF/fLthCKgh3w1pC6vyysAgynJXc1oI1oWABfcBTf6aiyz2r7RJB42Y
G6ufjhkVcJk7dklUsw8tzEWqMZ3JKcN2yADd6nJqKfLWbcqEUMiEtaM1JjIQe+KkPx14QU9Yot6R
nUZGHY0E1McVWvVlk4QLwgTr74Mcar1LCqxOQH5pjKxofLRnBMfsDCLNQvimozLGujo6OvKdaGz+
qWEr6tyDHq/a01mSUzAbRUCEu0m7nJ/0G7XvXQulmLEkSwE0eCM5OV3SzgOgAqpu+iutx+Gx3Fmo
70twLHZU8yXmSo9fLxJZlFdVn0fjwZG/rtDkZm6xrzH62D0maq1+1QCtVwxhkFO5no3bRedP/1NF
1XOZFaaEyoB+wnIkpqx6VDPpx5jyFzzTVESMP9leYD42fCZUga+LNsiayuEAgG1PYvaIBhjt71uc
csK/7/nwpEVzIhtM9sbdjrvBKaMJ9Lkt4+ra1GYFmzysBXf0Ciwma7Z2MtBPmst6eBH/1BfWEJ9+
67NN6f8VjaAQX5gJCYFkJyrlpf1SqsVwgIG19KiUc2GCt64EbL5ZQwEIfaSS9o8eEkgQZvbZrY4N
BmP43eDal5jA/Rmcrvkhsev+Lyw/9YC2qZ38iG2gNVo64YN3plbUG0O/shxqBcNlrY01w00KFTG4
BBlHM/xDHNFsldoig5YckGcqNrmzNvbuW2CmHbzS4ILl83yVEnN1SSWGXeT/SsLZc9iDGEoXK6IY
AKwg3lWQkWTf5uYCI1SmcaRD+kDL0aQea0PJ8bkWZSyzkUFMxWlP8QV1NsPEZbfDa65kwjp2nQxP
wIAP25LHbdbDBDXII1NyKR9ffU/KCcmNrIuoTzas6WFKfSf6fkneAnBGsZE3gkD7aAudq77Ih4ih
CN2gRKdPjm0bsCiV7pSlqJiuzEhq98nZ0YmEhbrz7sqLwbHxDKXCroGgs2Iq1ZQhdcKNZnL7OaYC
6FPvgKw/wfibQAhv8w58lkPDymZonxMosGzRpLB/4BHCdpK1OLWKYmiPffowgPlbZoH15S64FSPa
mkAPVFDB+yHD3LlGrayNTcHsu0BiOjSXNqsAUEI3lKpcyXApRrB/3BMIOo0KKpejbypF4vpUakJR
6HRPdbyFg1EbDcAvOpAnB/c9zjSp8tiajiqQ6r9K6Vb4u6dYj6oT65X64EQOek3ghgjwdYfDoTfY
rirRdhNdrrrBczamvhKEQ4i254lKLDxvCABuFBlPME8WsxboPwI9uOCn69aLUbJutO8iCMSXscH1
oj26qActuzFAVQJ3ioOgEGCVbyEEyNdCGjtz91zSvKk1ZJ7Vxseb4UC9TNIumIlcXMYcfSsnIong
xBhqJzmseYLEh/ufR64MIQoRvn6D7PLqmCiJA8uGrINbTX/kDSQpXFOKVcRL9Lea8a//6KsbC8ee
yKjNo5TPfNdOpKtZEOwkTx8DIi/eFacrsRkLgJU6EpqvhECAiQgoYo4iO1RWO3Xw2Lq88dQvAE0S
pWFmM7Wf0IzNLzIS9OWs0KgsdYsDE04P7C/dMA+K4ZsZtS3Nees8cMV7dditn7Dpg1p5TmpaiObn
w14hup1/jk/pwvYqlRF0SGhCg5HaUzS3Mzoro7rvvDUIYlyGWhC6h/9pNWXH52ZjpL4zsuVhBC4o
uKydelGTRFkDtyjweaOqTXiHFcYvEb41JVTak3yGnHXIWSypZDz9gVNFaDIPN/jN0aRiVt55Im7X
PXuNhOYvEY8ON7KRT2qpiS1E/7YPzDhys2vcQwueN4GUeLk6OYUqxbEMW6eXMMrG3hW0qA3eIh9L
0F4TLGO5k/wrcDX/g6Gb7JGexzYkFCwEm28fr1J3jDHiHYdDqaa5IwCxycUTgdH5DFcQ7yDbql0P
F//OGYv3ndhXlv6oehBaeidNA3kPwhpDUcRDw2tUALrY4Tch2tDibkCfX6NY5af9YtccKdRLggGc
6q3YK6JtHnjMQz9Mff1+R4+jdSYZr8eGefj3t8BJ03ij+B0dNqKOlTviGwAy7RsN1Sn5zPzPFYRY
kgA8+01sA0Atn/rSguihQeKR2VTXbeBZnpwWScI9z9/GuEuLZDmNznve8O5FW3uKBPzVwWLHapq3
n9kkdEXSAo/VlSRjE5xVA/neX4uNYVYOrMt1RgUIrwrRTYGLGD2qPnhi4kb08ui5fyyGAus6bMct
0pEqC+DFZuhRjx5ODSRqDF7G/bxyu5s6SncOkLyRUsU/PZRgTchQr8UEzzzcEO7yd7vtyH1YaFHY
zb2vj/qlL3BoqGYM1KVemiJnBdSPFVtvDduMOI3UE/jYwnIjv+UV4rHWgEmcjghfAbhHPYyUZWRx
gkubS7KNMP3b3zIM7J0Hr/m5PV/WZ3rDAOfdjkeV5cqZeJFeS3G0TUfdUI7M1x4gd4gFda8trhc5
XNa1MssC0Ygt06NNVQi4butAQmLVeKdB/T4Dwys2Sm66TKILJd169bIuhtIkUXWb0iSL/A4E5Tya
xTOM7Kh5Ac8Fbt2BzKkYe72IbhelrsWyS9qhk53SLh41E24mRP/iFLqbXZA0X/Rei/gvVUt5WnXQ
jD8rilH6ymB2T8t89g55hpnuGaQTcaDsIhBlBB8kUlTf7iRhA94fQakx0GbdJTzKxLH9wwJfw5iX
cqdpt9oXVkXd/BDBgfrkTvwptKyi8yNtrusmG52mkDwJSnPcajEylqrBg95Wejq7a0RN7FHE+VuR
R0qJEXrK9x2EoZoeoFxuM5OUzyOBmv80ua4zF3z/C1ADh7tdU6mRj2MEO+JQpKKn4onvVbGC09X1
v4s8TKZ9b61zwfy2/E/Lq3ctIVx7gmWb/detMbfUE+Ylx4CTI6irfu/TlhWUIR69z3fJPSeJuZcR
AGIVwqpejr40wYTOjzrCiUSbwx8Wd2hMuKxbGT9m3ygxf24/rKFM0WEF3j7DzFxR4/9MRuOGvo1A
HMnxQ2XUkwoneG1oFvkm0nj9zI5IjUVEyuBM8UL5TyoRNKvte61dQ+4iPUc5r48KoRzpPtg+6rot
ZHBzsBtZ6LQbe3KeQWsyqW5/Q1GoR2HnZ3SI5FpZaMUPENnmG+qxod9GtXc+DaJcBmsg7OsOgeGa
S1v6BuN8oDR57NSb35z9no+z2c+vViCLwPZT5UAwXAcqYppIDD34w1ekI46Cp/m+W7OslBMfTINC
5TPO6NMBSp1B/+klh332jN4jaDgV0pJ7eOfw4eqeANOAPC7EGzGSbdHrcJ7JD1NaUuNt9B5abz3g
NqIhn8PABgFTHwLa5fIfu0PydyoNBNF7O9FQvyJprJrvmUkoM5/uzwU8oY9TzEkjogrPjmJZshXZ
TWkFyt4JcWA4OwC+DFAzCrxIBKBBW/l9G/JkbHBUa2G6VbQmAuVIx4E4hmZMZXaFr6gOE2nkYJo4
uVI2ZlgNCGQQTRNQ54yAURg/j2hXPRny4QdeBUoCLrLBLFgLs4CfD7wfiQRe7XXg/UkimdWl88XE
iJWcGm8StlDRMHuXO3c0hzR9YpVOxWfqhJRf8sVi3sIiRiMBywWEKi9LNsAbwT0tG9TcrKdQHnbE
m7/giBbBjpPyuv05IACaHjQ5kiFwM4kIXbmZmRyWj3sc6+QCE+Lq9AWtio/mHFJGMU5at6aMNmnE
Rl383zC99VxkIVV6JORYdN/FBovFB28rWGc/3C+Gp8fJJNlDwyQSRECBWgwUWla+GniLX2ehDvtb
AJSdWB6KMwS1kk8HDR7d2zgqysy9NDwAgoy6qUgUAG2m3qnRDISnb6AWarpM0t46UgyUmJMfyizt
X6RFqBf8++TdLH5G/hqQI1DVT9lOxsi8wi0rNdJksF1mRJOmSkmhIBKmLozJOIszR5Fen2l9BEuF
QLb0rVjjhTfXdKUY9Pk+ARyfyDzDVJRXTbemCE6SF97VRxHsOVJpD0nnDx+tDVGF8fBuc7bN66Ta
AGbYjGaRtTECCTSwlZWMgrmyeU65rvw9kjZsGFfYREKM4cGjB5l7Zrc/3oZ3az1rWE2OJT+SQo+F
2zRmdin1aJFfvaglPMG126fHyhwkcjoUJzP2WZsivW+9XBXHhSsZxuSSWCedNl5/dzHCHF61d31F
DeauN/1PaI7cRGd7eELtZHrseOtc8nBDrkhVLMlh3QMi5qHOMqGbvAWRsohOvVuTKF3GCtpx1t6u
zCIMJObO5wvqZdQZHOzKMeRMxpauMqVBDHImKxF7mtZRFB1YZBQmok6an8Mnnex5mIAb2/txLHcv
wEfw4JmvNFqeACF+8urT3RRHq5eXqghageTE53J7HfBCfX5wzFT06+TxBn/3/A2lp7yvAO/q24Yi
QEiEgeemsYcKQsn8Z2cJU0FWs8VUCKuUadais4VvBqHqsVj4vO0r/ZdvW4PfV7KDFCx50sMatq9F
Pf+TVHc+YMe7qT4MT0yAFJUkNCuJaQuHc/BlqjC9k/XmT+UhMin/b3St0rg5yJ4pjeoMaffVKi05
4ABQ5VqqDZyF7hgeSe0UJOMJrwFiCjnOo5X8Bjq/84d0O/bV8Nt57y6rzcwcTkMW4zu7JOd4Q1pW
fxpVI0VV8dQ/cBq6Y+d0KAAWvM0LP1CVolzC5hfjZBLVxy/C2r0fY5hLZO4q0qsWgzluKXwMxhKn
g0fzTcacuk0EpoI4dNO4iWFMmMPUsnUZYg2z0saaCkfaoOHjLk0cfT0hGQQUBEc0vedlD5JyiHU7
scNKTkWBbBTO+La5Nt9kH+tWVghRHzhriyGTMVt6uamYyNrrLjdDhBQjv0N0CLeBusEjRn3Ru+Yk
huDV8PrsvVQ1oL6pHjMegdH7FoBybISgkLcOSjxbDFjZiiwMhoBZt7kxEDJquTvH3glTWFaJysYZ
Gdm+HSZZP267xd6QqZB6Q6TiujOI2On9Z6X69X5z1JRN+bR9TUgjp3b9RB0nGa7XGWKyOYa79HVd
yieX6YizjjlVpOCwQOebywAs3nqOqSJRYhot2NeP1dOBHLv5ZrrC9vmS277AUDOZEGc70kricXYs
85pEmHdOs50zysUBgXIGk0/GpFeXzwqiddJfSUVK4qNctwCeXyIo/WtZ3z/e0V/hMrY2JCT0fna4
hjDDyva7pblgCgQd+oLVpuc/eqD9jPFF2F/635OEsuGY5JmhodlbAd+sNMFX+agN0DgFkMFKSHeB
LowArS3rUFRmYEpBIJJhecQxsoSqYgBZcwh4roBUV2q24gja4mE8jDEzeqpO/3rnAqV+m/xFh/ip
bDOQLJgjuwG1JY+GXsAxw0dOqK39Vdzl6qh0cnWnH7LqMvQzX5bWC6qoKd72On4I3spYHjGmmr6k
rItjrqJpRmR0LhfgY+oiiHwMcUC+JMtz6VMhQnqBl84vpDZXPJrJLh3vla49LxxzR5vfgq51PTEi
0OtNUaIj1PbXgrylD/31KC98qOCKgazDALFQknNc5QNDCytTbRffzBxA2dvZWWK8C0uRdR8VK4Tv
xZ/kVe1I06N8DVwhez79AwyBB6kcfIhWnE4iibUVHLWcrdfXFcDojujQNqQB8f059KV5Og3eAgS7
Mxd6LqKzbeWMOn0L9BOBzRt7pJsmxUQTFqVSFuYIhFYNMMnUo9Ea19rkbdcqi/AUC3I2CwLxWynp
kltaDLDiQtaNZhI7ppo6Sq/h0t+tE7OrZdGwm3PLUx1f8pz98pWVkEbc2OuI0lg4vV1FEbmPT+US
40hsIsF4WX2/+4bje1DrLT5LPuGqduSf0G2TBwXm6q/AeHOZ6bHUkEHz7A2pX7TgqvCN/tj3Msml
eUE79Pq4CzV2Jzmq4lEPn/L0CqQEVNPzT/i+/sDc0SNcCxVVIfAXhmU6RUag7y5LMVzhmgYhHFww
BW9zWrDVeAJ9U8sQ55yMITQfqncOq4LwM/0OAQfzBD87j8dsKXF+FhkkLF5f6dyAT2c/Bl4Zye/c
ZvS8O4l/bHW4GKF+4mNKSyTCUJ2UoEWbcNpt5By8dgKJ9NVBAHLR6uQ3n8wjCwpyBpV9h8c4wvfq
MGFZnlYAFzlorfwb2yUyrxB9bE/7HzDoiUBjQ34RdY+x+BXoDAr2hDL/qLr0k+ttMrgCflKyRIIr
BXkZof/aZXARvAI52UYnihmuNAbKBEfH87fAiu4yJhGpBZNKTzQb2S55usQQdu8tGBK6bq3EUSb1
c8W4T370twMSDuU4dq6eIcnyObzWJvIr/nuTYYJVtf/gcarC0b2/h6z4GG/F0KBveoGAzQ4a0x3t
sI/TACjK3649whT8jcTsu3qOutycD/t3wt2hQFAnMMuK6N/hDripqfq3ZToDf3Xs5WSx//cqqSZR
UkgGYaswJLFVPtyFlfFRK27Nbe5/7J1thV9Jq1/Yh7YDjHVyJog5H0tw3stcNzaPoqtlEiD3mjG2
DGypk5can2Ikz1WelDCyp4JPzC9/ql80ycJNXWuOij4r69n6mN2X/4cMK4S2bpL9OsZ+Vf5LUMIa
59iLBItkQVHtsAOY93QsZIEazsbr3SEhU6Pa6ffT24zdW2F2ajQweQlCfjdgZzY91mF7lB0S0nNK
I5tjS7syfI6AtzGScYpCBFDTOs6DGeUgs7IVjr277FEdile1jvDcPSsIGEaX75UaJAFJA2FduGCQ
qAxs7qJz/cSU/tIJ2rzoXdhV7Ua8zY3CgkFQeh7Y85f3+P2qERoA9Ysln/enms4aShi27Z97WsaW
Scm3CLuEBRk/Fy33LNS7c8oCkMImyRjoBziaZmaO2sf9mrfRERSezhToeaIvLkucEKX2ZEhYfk3M
tPU+s8c76rcJu4jg0X/85k68fUAb8hUhYGxfX/2UfqEED6xOoCKt6qnccqNAnxB0ETiBTgVpZraa
VXVt6GFEKnQjOmxBuOvhedstDCUaae7y6gDBIiCNmfmQYs9drO3S31VR8l/EZ44YIcSFkwckiyKV
/e+JWCJBlxOST2dOVvDK+AjSJdecrnwhsMWn0c7n3h8dMgXU4LW0amghHsb7kMQNsLZOFwX60S98
g0Gt4uUdolH7M0OnYgXLNp9PxCX4cjc/WwKwVMiHb9cV9qCpF0q7cmsjWOR36AsWa1yhqgGIuJd+
2rTFnlHAzADZLotCIIv+Iesb6o7Pmmf6AXb3Fvc/LjruzxwPB8XEGSo6pyNofWgtJiJdIhPMJ3tI
gnTegrwovAoy62utoU+yre4snXZ4posKaqGihxoULe8A72wqmAvG1fBje/5UesY3FkKpSSlUAcR1
cMVuIhN5/xotCHjEjoqHxEAcpJyoRDe0x1fPLhiL4mvbGbbIZ2VSFNuItivZWBiyVoW8aBgSNIOD
sDvn/ZNFDI9BTqmuRQknJn3F9wwYZZvrqYb1ZypCGZm0jJYL0XeUcsuQXWfXIsOO0D0p6LfHRfba
yTZJnsBILgQKSKkxK99o3xNuO031ds4PZpgL/juf6Gs1QFUkGgqsxVoM+5/lulkTSxAIGY2nv3yj
LwiZ9VAZsViw55gbLDfqT8PAF8sgg68FgMJY4mOz7ANzeDc/DDAvpzj5HotvtyYVWQ4V5rx+HMjW
5LPPZKVWgr9L5Mmu45JHWaytrvhJePk03fFN5OnOyOzjolKJT2Vm6DfwCPOl1PPo5ETRG8zOegEo
PzTOwriS3hY2rB+z9f3l7MJ6A0nCEy5W1fAUiOLAFDmyt5byGJ9uFFN12CL9BIdD243wJ54kSTMx
OvOOjnNDEU+GaIaJmOtQofwQCeWxryBTIizFqe6saiOmb2ux+tX8sVGx5qL7mwVlIb3yv+IEeuxC
hf0hKrAcbe+SOkLLwtWbxlOkculUS8Kb8jfpax3al8jQHwWckmdVxjx5Qj+XmPEtFTA2599oHiKa
mzupiBnw03wqoF3wsDjFAHGAcRU3Cp92dThaMsx+7DfUKvxKXh7ilc7E7q+1ISs5wmCm7u6KLWlj
JT89bur4q/TGdPoyr7DPbNmgSRGqQ6G6Pi2DgYhmsTWOLEXpZ5kwLCL36pBWQfCUKPU1xJswk86q
wYfETh3qR1dI0jCquHEyZbA2VkXaBBsZIIrr47zoFkYEXv7UdmcwCugkqdDw/iwCfn+QBy4W6ztK
tiSkZsLQmZbEJm6WrRPxoLVe2W//qh+tSkd2TjjrgG3pClDfHJIWqVQHIUBnvVVUr0LCDloVOZNR
t9V7krXAYL5054phS4SUtI94TmofnJw21WSodel4LZvZLSvLBQ6ltC2DgLnjxZ2oGaVwq0MIuzJE
MZSEKJ27WRFox6OPq12LTNsxgglf+tzNmkRzurFhGWMoWAeofuNcUUY9cbJ+soAoAa3J56lVTBUX
rm2oiA+0pcKF9RxyaOy287bsRYSICPlgk7UO+PII4keZ8fDyExfU0D7IsfG4cdGD7ggTtSkjiMI+
NixLNqThVVvuEqXOdKYQUK78sKfjGpJX/GuqLTyivBc84pLDaG6wCeWU4i6RcHxQFoA5VKLsL6SI
nwIxS4bn2BU45MuLiJSP5hRO/BXRrR/zFbP9V0+KA9fucfIZqETqvu8nQbpmyzHuzS9+obU6UP9Q
hhFmz3msoYV1ODldRg41ipHdFnCV+XwxL6mh7B8Nqg18mmdFJwXr+BoxpBi20tOzAfelYH9kAv8A
gQQz3Lap9o36zKr0MT3tp5DGFJOMzQ6zKydoc5zfNaO5JYZZK0z5wIdVWZTVKCk9xInLpYNRqj+E
oAP2OKVe92C8VHNGQtP2HqGIiGNS9euKW8xwKzwmaj6lpPTb7RryDFXdUDgweCN7KnQChSVNJpuT
Nj5M+9OD3z+MBvPb3CCPUjZVgdvJWQF/WJ7sAX++k6T6Y79SKcUgJtVzswk3y//WzsYCJvPbmVLe
XAMmOvQMk4TkveT0E3sIc6DtrAYTnnCFzf28EPLmHwQMHpqhvvotE5wWoi6H272FJl3NPT2DIC5c
9YpKunq57Wcczt38STlsvpQpunUbGisjEjjGtbc3Kvap2OkrbWOP0SDD5VC1/aa83aVwM3nlXwqO
Kln6SAqv1JX47ytOzDul9vNRDHDq40jrDy1u1Cci5FeSSrZezi9KsGEpUFbqLjIYAgZK0KqXC1f+
06m+f4Bs+tGnGuoPzzy7qZyxIPL65Zvs8eashTove5pr2+6jI2ejfWnwpVHz0uur3mOxxB0XIufX
ZNVu01adAWtFxX55BSy/gCaWXWLlVPtz+E1C9yfyX6iYR67vlOEpZgfR973WvlUxM8p7AYAMbJ4l
pJgnt/cAXsZSJIxw4vv4zHykUOlxThbFQibb6802E87oMiQcHDijlngiI3pmfFiGr/RmFgMH7wSR
6mK0Xve9ja7K5Lf8Wf9igjCZ/6Xf25jjBpfUCWHRa5FLvzil3mBTkqIlzxgG1fWa247fC3gVXlMf
CmyjBdUcOfslFXC0CvtsfutcYkn/nMksy6sbN9cMux8+Kt5qv14JVsVWCU4CtfzAqQRZVmhCfBCi
zha8+iWE5QMOX93nwkTSSGENb7UywFT5hgMIwsFQuGDV1rgaJQ87F/QGDP16geahazo/rQcA++r2
X4m338UCoxiK6q8LYwSMq/j/afxopVMVxyxiVAFUSRf6k+WbA675ZGNxuQkyBvpJv6swFEyTrAkt
kIiEnCvuua4ARyOl/nnP6va/YmMmNC4xBYOkXt+OnTA0rSq+kNk4aDVBeJe1Z/JMoKjWTvSS1L9L
5QG4g/8kjdmgd58HD1DZScBDvggYDpiPL6xINgWMJdHRfmOcci2rtMHZSuL0pUiW6MviuXEqMis6
CatlouTuVIYgipuhz0TPGQSsGVXycOnXgPck57L1kfC7TsZrEj+QVLSz0OtdkCgTrhghKaD07b0D
k+QumLsPoiv+fbevhSDvXr12Tg+q1zTVYiVbrJNLXbB2vBIGH06KPv/nL2nO4FAnY7wbkj17Nzli
mdK8t50OZKHHhYCpMfGFMOkE0Z99KB95htBexUPjUd8hZeppTIWhWA1Ppu02kYEg3scgK1R1fbC8
b6R6aDSjcch8DCQLQRR1Lrx+476y8+oElERbXthDXLzajV0lNdFo9r37X8XxYYMKbgrfRVOOO37A
gIraOvnJPo/SIT7I7q3/kBT1Ai69XikbL+tN69ktQO8SPRvHrWnbO3cQf3ctbOvbqC+jDbD4dTRL
nJN3CpqepO3wp8Xjm5OpzIpRPUUiu+35BSqhupRmOAGqYXm5UBwVXAlJY/OD5fMx+z/8SlkNS8ax
FqPRCYQpN/c2SlCSwdwEN6Ktbv7Iq/Ygx7zUpYzbS/ban7AzyaPsX2JuF7SQsnzUqoG8Qya2eyG8
2z2RCDYeWVkfSPJYZYWEBCb2A/MToosACTzOwSYeRbFfEixQevdUJDkHSJcg6HJOleYkQ2h/3YD0
O/RXgOO+qdLO/80gbwRmcJnlLNb/AEz/4j4jdO8TqlrfhgshQDb1oa/hwcs1FScy68+g+Tyx+ABL
liW10HJHMzsOeQue72G4BUgy0ksokiobxer1X/yxO4uHv4l5phAnZG0+Ncc3GxTal0oUviFZ4BA9
lESESTy2m+TvvrX9ADQzMhz7BUUtyferR8PFv+WQILxSDkFAU6hhEEPW5UWFhYuiwzUiMhi81u2W
S+ExTSiBREmFeaT84xdpWQohSJdwzV2GjBQxjUyXJBZrcL+bPEiO2Zd3FJIJ2q5tdw9tXK26O7oR
DKxHG6WKsJC1wiu3b/Qc/CK3oHkQcVpCmHJx5Smg7jVOGTa+vfC2TaQ+aRgBtlJs8+CJXckuMTnV
SBlRHFl0iLOlyYACjcuB5RyJRAe1/p//b4/UavPnCeO6Z/bO0z+VqZJD5iwm/Wu9N4A39VVCoCoW
cpBx4Ds8SmpHzdM6wQwHfHkChPAK2A4McvPY76CAvZ74DcEemCA86I2TfoU3dWK5u8vBizvvnq4U
F+hh72gelcegXKiN61eF9zbU43gzDHssNAvimiMQ36bS9TYskS8S4iHlW3YrQiyQ+zVoIrYVl2My
a4Klnt0J855xAgLoog28b8ZMoyyjSbKOjziGBa7wf7jpY7b4OCm4dFGGJD/fTV/MbkvG8B6VSgly
0O0bCghsy6dRuQb9+nqFComQDZ0iHs/qAIZOsDzkldheO7mAqnypyrG5AOzG9Ph3L9xHPmvzFsqd
mOg2S5Y6YMuU7gvxWfJThyRCxGbF8XtU3ASWFsCfz51VFVSyfZvTqSUDnEUM/HePW3c4RBep87Kw
w4/1oaq9CjGlPSFED2ML5N4ShWH8a0wI2ByZ5TKZ9toLEQT4dcOljxNntm3pXlbziMHO2SZbQgCW
a3sYPQqg69X6lExP6stnklHM4jOi21QuzZVGnZtY+9vnRuBbPk3cEQlgNEqFrOf+sX432XqHqwbI
iYsPPYKNrmeIj9naU/vPeyaxhbGVSD9wgIjbJPVDEAfJeheE93UtJ8uXHdXWlyO/8E+jdW7rCPS1
XzNF+iMbhf3B2Eeg6wC6eCi2yHwK2qiUrOmsn7fs8SQT3TM5RQ8O8QA03+6SWZ3C0uakQpQ7Deqo
glx06IItI0oOJs8LP5AX43cy/mhqvm++9tkiNsjturpXRmjiluOLNCWxiKNN9ad5QqyhjNOeba1L
WOAuqFsh82hVpxy/8na/sqeQHVwe5QO25yevNQQCzX6S9ADvVlR0sPAnpjPAv4URGHWggRWakMJp
ycodJbWU65FAkKz2SWtMaHscTcUnsy0TB/Ch33Q9dPYqRwZQjlgPwGWvxKjjRkGJTBKHh9ANgkKF
pbOepkZ6tFDp5xSCJRie/Lt8cd2WcR6bjdEXhjhcc/xg8/jE+RCm+Y5TQVElocpdzIO4QhjvwqQG
rb51DM57VezifCluu/SJHmiiUVu4FECkTOhzr+ZtAMuRSBdmKFX/a7Uc85JiSrxHE2jBcROyUS8G
7xkIKxIGqqcNaJZO+lRPf/J2BH10Q+Xs4G6431knxYdqqNW6rWFv38jDONCG/8vPM4bUEBcNuqw2
vLKnr+2ISGA01YJvRBJSKT2tVQTtUkbxVjZg2cc71j/Hvvxgu4E1cFlGgTC+arcUDF3t572VhXxo
lKKtWhIhgB1zXbPEwJkKh3YaZBirGFdH9woBVK1AR6ytiI/UXAgu7MvamNT4xmil2c9Nvsk/ujDd
wOY45VDRzS7WgTjw7LM77WvTxzrEaELjBMXUm698LjqfawccZB7Acwm8SK4zxRNH/Ll9QId6gD+l
qUT2VjfQGt+ZFDo9LS6O2YeDl5QIkHLTTNBf6DEeJvyKM+PI7P9N3rQGWJ87iPAi7q5ytRzdwCmO
zPjYzbhQfbJKiBzad+anX+xRbqoY9EuVXJvSvnPh5SPO5pzT3llmM93zd3xFAMpJkPXQ6Lpn+7rB
ul20GNKv4hATW/qkI6mayeUOi483wGgE0N29D27iqm4+mln8UXgcaupnLbt1Ig9NolgIZI8K0b3R
on7oddTvwFQ02ESE3VcXaFBLuh7W+rpTvjjlM07rujkm38HPOxON4pJsL7F7qL4ysUzFTwjOFNEK
VIc6mbDUq1PF1w9b3In9vBJSRdomi9wZJa5pJBp+kvm7JxGP9rgQYEDrp0doJ336YNWBF1sYo7S+
7xdBNxjsQpG9d3YOrRqV9iIUH7wZmeOjdzhIelUDAeFSVPoRakceHTehkMGdIEa+a1l8rV8arZRe
MaM/uD2puttO/3r8EcukmPd6AEzUdBXrGLFIz4blOHQTLE5rdIrHuJT3jSK9ceGoX11tFDTYA71L
6KhlMvibwUkq8H3oqpdbiKkDqLDtlcneGmjhH1X7T1BZmv+xsAJD907DSMzGZMMMgMXpS6Mini7h
HXtXHUT/FtfIYk4MUNZPpwJjsq9NBNVYoNAZPh8QdKBPXxUAwzAkJepfjVdPueymgHQKotJpGOiW
rhxpUcftXsAfcnm3Ordelj4EmJCd8lVRr01s79BamQZtVcjF+pcYUi9niG7cUqPzNE/KhHRkVCIu
MzTWvsbtNACotKOA7YwdO2/bmum+g2tBlwdSJrrOyl8xUZZnHi2WAYLTZ5IK3L6NBsFNZBv1As/d
4OCsrjSiJpbZHPKi4yrzRCreTqksNjJ5GagIL4mzugm+oswtIREyh9wwABsdnYEkwokiOvY/H0x6
osrQresWH7X4TkJKmJyrABZxHJO7hRHzEnJAbtb16TOGEmPSSgUCC6gQOUcmjH9ZVBDrBmyoIcQr
bYBdVfsYN4N51BztrzIgf7bxcF7u3TmUoG+zak7HgyKQRa+dEcsiOuw7Hl1PWCnkYz8jxntuS5Ma
m3EBmZQwLNeiwm6acX1r/SpiqDzs+J0wv/IYJmpJ83XXH5UHlxQzzQu41wQuo5lfz1QhQAfA/o4v
hCVC9HHVzP3rbF7qpzOSzih/Utv2w9CDdIoyRZDzqYhIajxeveORXj/gWYTUKhnmh7q+mrolurCc
h2lP1ef0rsni32Vx5nJfRbMQoIpmVzFQsqrvaYPqgpYnpJfNP4uMSHudY7M37SJoh5Z0tKSxB+Hh
1Yk4zCyOwRpNxH/fYZQZej1ULz9dwNK7fMGJXxgQepcX0+0xHyQX3GKL1AGrEFsY0nC1bD7tI9xB
yoYC6nTJWi4NkROvrSm6cbcclZuZLp1huhiUzl26mSWUsS6eiqKeihDQ++EJrnErLN9knGiJiugy
DQfOLGA1iJ//a3djSCwvR6u1ALYyf4UBofKD1PM5FINZjQdKp1SK1LIUD73DH9YyjfaGdI5HxTWX
M+8KBapErGBi/K2dHed4Ipz8V27e2XkgR2kBpokrp9aQZkZCzSoS8vY4NM0CArAOJbcfGbfkJCES
UlYLemCNZaB/iUbv3V2EGvww41WcRuvywuQr/8OJPhqZA9TZb9fMtXJamaS3T2/04pKHxr7DsOLr
70muGgTDwxX+b7cq/fWpeUqY5CxhT4o+GTqvRpqkaUj0qjfSDy+kjrkibeIWA6jivPI+la+tQXfM
8Dowo3lSH6MfKEjdJQc+rQI5xA1T1kRJTp0qdYBx735nCdGmOrUJ/4ZawkJLC8KHCyVA/qAHgUZl
7l2dbTKabHMh2R+GFnikiCS5GfFUPTIaHyUGCELtFzBW6zsDuQshX0EqlCdCariIxVHFJh2IFREw
jKq+Ca2xnHrYI4bKpcZd/YmjwuJp3J0gu63+xMOoylxYsOYdH8UQCe0Bs/jCoksQJ2czLWgnNyOe
3Tb5TXtTyfm+DurvYNa47c7GUuCgC9OlPcdyyP/TKBPUOFeZfanw4Ru5IaY/d/Xh14byldAjNrvG
4VuFpGtw20lakQYULmGZ59KsbYi3lS5gjgbJmBGGlT6NYdsGAjxqpEkDl1hBr5Khe31Am2BtfoOu
YLZbmibouk8SKL97sZYFAwn4B6A3zyJMT6gAVLzALa2gZzoCVbD1R/iGlB5z4QvFekiL71eMy049
my1U03+NJ1lv7RTePL8H8srCBlvrO8vV0piH2r+bw547uQ2XImQdjoTt3d7JOBUefIulx5Q/bOVU
RYmHlzJxrhzH57Ghk+YCQB/lsFJVK6YxBE4daPvRQqcfreMQZNAxEpLPqUS3CMJuzJ12rfuJ+DlD
ZjVJAzgSW5exG9r3lmOUA50UKhI0XOZkReY8iR28YjH0Lv++hV76KNjn33N+YZ0YdZjZCfj5fbrJ
haC3YQ//teLQdq+ZZQxRY0HBLidyAP++3p342c5SDu9Tv99vkLmi6Hdkee0ABc7FVW0fy34uaZPv
5KFlJoQi0QmpMavOCwMqwjD7lb/hzZjrSg/2tRnthPJo9r71tdjftc6ho3FLBqYl+FP4SgE0ivkk
uKIw0HNy/lzm2zt/RIOjen4Go8oPUJLPn0y1sDQxQgfTf54janx1tD+r54tkqRnF04jXOuo4q1nC
Tq5MmA5AEhhP8hxLXI1yHMcyCRkdaH6OgP3fTOdSOAohaj779V0jWYBahAal/8ofA3nDlVqbC0mA
9NypG1m4ARUqz1+mGQP6+0RdiSrutKVaFyFjNB8mjlm9t44jg2I7phxgd4GIHogP30IeVOeGY2FW
YK9AdA1RzemR7qJ/ggQ3t3xD1hSx272HPPVLPttrRUSS85s/WekbbmBSNCew334PXJ5xOpMELGLP
s5dMfbFp+dYssKBC5GWqI/pYxB/Ps/ML8Y9aSRk2QgKfNcoOSwNR19peJYY7rNeEZL4u+uLYGK2C
6JJ+KYLLEWLWsDL3t4raDv8IvjnIvfD1v+c9B3/mYGSNlxSTKP+mnbI+2lwHiseLV9JThdmnCk4x
o+qDWMkV1wSMkyclkCmrn58bBnZZcYMIv0Ks2Qs5FjB2I105dAEw7nOG1cC31ZNU1IsOdAzqIK73
RPp3i6rLjkS7OXDXt6ZUE6PFQTwE+U86hcfVY6rADLSyQQXqn6rZqAFZeN6hU3bfrcVnRzKo61LD
XVaKq3bBWrxS7JaTJbvuN+TP9TvZ/5lpcmnZMgqau5ze8uXVW55JKsjbdjRYg9rVEoMtQ7Qt1vgR
ekn4f9MFfua97tzA+xOL/o72gWqZirxirxWH6MZm9Gii1IO+D487hI2B7Jjueu4UlZ5oYpdj4aYq
Ku4vNNkI5+mQtota0CoSqmxGl25eihEc0f2+xZKHuI3Mxb5mrg15s4KWLAVdQ+/vJgKCkrrS95jw
6yB9iriCf4YFGmd72sWypjO1/RvK4VvSEDCtM4AGyQpA9rvzuXAH61vzXIxAneTAAJ2/OtFhVblZ
WiP68MpiCkang2JTwPN6lc0xvYtgXm4aNz7iNCKSytCNzKYRtYhtojf7/8gOPOJWBuWounuiXqE9
HCL0u9E0oHgvvqElxAJ/RNjIsTMrG/uRbgdmE50erOWCD/eghVe08Q+xfwyU1WbibgRoi+xCicSr
PFw1G1w/wSOT04MsdNWRAwaY0ZcIlkT2/LokR5Zg/dJNHWsJg/d+qWYGDTSLC5jYZxK02ZAsKGVw
m9m0UkCKMrR/uMCk+q8ueSJbjEz6iS8dlJ69Q1fABjTi3QeJ89Nfx5fjApim/Z5IylrHcEUsmMZh
rfLaDemU62/z43i74ECNV+Uf+GEMHJmWCA84Z87P3UCZduBSFiXcu3i2wlykZUrBMh0pAK9m40Pm
lUZBszK07oNP9AnUttnhhDq7wb0EKrrUB1dnYb2dj35Z83S54n3b7LbV6mOg6azth5pC3QxnYWOK
n7afFYwgElWy7zupZjjj+q29kqVChX63DHbHaoVHMeffzkVpB7+3/ExZ/Gmp4HTFpZPk98o7Eagx
uCgwteiZfjk4UPqs8qLMEA+r4bSKmKNQl4RxvPs32t/dIdjhIu/sjrUOvsM/bORBfmE76GPBR/0B
wcFXt8psBe0mT71HoXkVghXbs5GQzgNedXnkNvA7FBD/unwk0WCxIEfyKN7yU2j64gQOTI6Civui
hV62pqxP96xsgI+BuN7cXhfpfH45xcP1FnbkNiUKt/31gDzPFCa6HgNhOAmRgzGP96RX81eZOBTN
HWeQw2Xy6iL22Dv2XrOGgsCJzasGwvNC/sHp4gJCccKV1CQFnCgPJTfDd408VK1qHiAPkWbKAzKb
BF0C9TVfAI2E/Tiqj5C2zmTkfyKq/aeG+1nzuOGiEM9ra9t2Sli9/+256CF12regz72mjraOeMMd
Mm/hLXKi1CDdZtNAUbk/EpOBfm9PlvUvu29tvSoeJ/8iloffhp76pCxK54MM0x8NZS5vE6RzTRG+
+aeVOvsvb5SjQPLoZRiiudnXwfW62Mr3bFUGdyOMI8xIpKCGkC7SGjNi4avLyyKHGayFgiZ4PSkR
pjQAYokvpqsrZCSHyzkOZR01Ko+teQZUZfZVnt3V+rbI1lnWksZqigehRbSU9bakaq0dAJ7z6CRN
hfXkmqRJWsNeh/icRP0C28+flhF4NqPLc1wLGS407rCihZo8JMqi/it1SsaV+K0O3UhduU6/lmEK
ALW4UgiglpFPorVJErHJS1ngAFVqFqvKGAgtmOvafAzZR7q50IHvhvOzHS9iSUs9CDs7JgxLOcIg
bo3WZTZg3s/88iuZKyd227bWqiBukR0ZM7DJj7jSmbEMOcLTl8JfKBKvndEsFOhqf1gIKXliRSqK
YDlCeb7c55ibL4WU9uvYr7pHfr6o+z9zqIs2J6UVeB+l8woTI9tGvvUNE8VOAO2dWaFWloVJYu/1
mXO+7ojsAWgTDabbfvaur65iSdbOS9R80QdR2b/+TBdt9hJaxFzoZGGB5ls1YT5Chli7cSA102SU
8/xbxCsXMkwZgkPOfvgw81roKd0JNPG9Tx+3BN7fbThLZmg3Ge3ZPspcnodDpvKf8cu7rPuLKuQs
9wDD0o9aCQsiOm0QGmsaE8bN+3PD+Mpg6luYF3ZA62FAuJ2mmQ36rAFRa3WetukdlH7YdIO//kwT
WUiL2nIiAoy1DvcdyWZm8NWAipJB3dbY9I/FHbnr3utPIjeVghILJhPBSkjhFR3zT0SbzGRbp7N9
G4KErLZCeysDOxYjR1OmVvQ6ieUH2Ak+FQU5zJJezKBAC755XHaJOWzZRtGcZRsSLlqMmxs3uj++
Fry2BNEBbPYJKhho0rt8STRlpzjZltJHq0kYgMCjUd6ya49ejwIBRcFjoZgo6aLRsHm4w7PcfYYM
bkPyMVa39LEY8PwDl7NzPloGmdwJeLRYADWMRWCeemi6cRgBUSeMmKiQqznCNJ+0MxT78EUl0USd
RF34do2EBLxc7RZ38EE+iKNEVDv/XxahGptIWDoBw26Qd28xG6wXy+9RnMYGiDzhwukABNYkv73e
eDunWzaBIofLkqPec/kuvi6imNjcSmNi/mm0tQ9U8/WS61JAgnkQBFSTXxVk1KN6TQPYBYZbHouZ
YRophqcrDiyGwcc6X8SEmVIcRy4kA0b5L5gCjICYUJMGXDzabXa1eR6LfRcxFaycXiTsVIRgJ3PE
WVrpL1LiNmAgFcuN8bHdJH7NiO62vAmGpOkpoC220TRvlbWl0JE+J0rO5fPUlYPKG/xdIkKKUh5X
INGjUpdlfjBGeodwq9Lrf/3xnlfSuJbMpF4kkgK6TPg/PMYeX3JAR7vmvnWGvS1Wr5FNdOrQDGdV
mfF+5Z/p28gzK6aG4XInZrtTNuTzdYYZptlsbAttOjDPTjcPbieWfZXqkdedzMmfnB658mYPsxUn
jrzRWhTyJZ0NOd4YqdBWZ8I0yuwI620NPV1kZKJIsEaxO+Ngi3pRlQTw1N22hOx13hiO1SQ4TuzH
grHI2dmOCi3ZOfd1t/o/Fo/v8Q7QMnuMsWU3whZdn8D1aiLWelfqBJ/r24WaUEHImgAbXymRjfll
57DfWi5mGBvS1e6OwwhsTsCu9/+wZhrS1+1dtMLj9uj6JDTE5clqff6sK5mKYnHvXLLaJqbJlfs2
kdYU0PWRGLZjHXf1xbZYn7H8cXvS8AYur9MBApSTxjTWnG1bX3Pe146+8tuPqqSlezBJqcyhziqH
RYFCX2C0v/qu5sLE/x48vDfnsB/Q3X/eicdEptVAGw+cFY6Hg7/+OFMAVORt8hQ8eBZAo+zUz1UK
IdjeCWA/amT6LFwxgdx1fS9fvdSXBZebYd/ZwoZLkIpDLZwBkH1wYIsOSTAlOYdAubgvkAE1oy0I
u9Ap+eSOwIfDY6xB08kG2CITnvwXP4IkZ4HI6PGb0/0q3q0kV056sHo2gr6GtVFzKXui1lmdhNm1
cQlNHr32VaujTs5VZ804AYEcWl8xwv5mdUs/pjUZObzwmT/IthY8QQeDQxMkySt9k7M1EjKCw1Y+
g0o0f4ZdDw+ykODRUJSThZHWcUWqf6fms5VaYIK8fLYLr45BM3Ui6fAcdNhoA5hQczEkKbdiJBq9
MMqLRheJNJntumq4fKqyDkeKvqPHjDaPRxwdiuiiVsWW47wTjQdeQAfoI23HI52wti+gki4XmefP
dIzSUbMWob3HMqM1styMj8xeDFkD6aIoDCMOAVvQ1KNAe7bcY47RwXF7bIbYJVr5I7zauPuDIDLs
Jjp27NpsjcmPXHpFwa1vmLh2G/IP5QsLOETqVMZm1n3tbhRmvpY+lz3dePy0/XIGjIXqTV8hjSrk
yKsaPH2C6Wd3eQcVW/1no5CLLp7nyrhBAf8m7/Y0xDFwpJ82LBogHtv9xoW7xrBGnPgAlnge9cea
2jYLVV8jDYL3gPVSAwhdcuoe90ShUbSu2S/dNf4JAYHTT7aiQ9nJEC/u3/xxyIy2oLBMYxJcIMd1
0ntt4D/z7AetCTMdYH7IvFPdWvZbQfQoUO1d4Y81hwniiE9I9G00PlfWRRCSFlzfSzPHTLlIXc81
Qg057+NxjOlvdjEP3aos8ik8izS7Mo+MqAMB/EZjAdDCFnIIe2M4oDM7jf6E2YuZBBOAO47QpMZ8
sgFX00J7b1puADyk62bfy/pBaOhptMm6p+x7kpRnlk0YZzbadLEecmVCN6+Dwv1wAROfqglt0Pj+
F6HqgVYoPSo4xUquQTPL2hhDpXnqLPTrkBu9+k6GxyPT5k5ax+85tuQ/IveUx+ZxdFoAefmRCVF2
SNTvB9pULaKjp9xCLI30sC/8nyNWpzZOZ5mRLGqCR5yX8J5qT73ZM2Utx8+zj3+gBV4i3mzEcTDk
cWbp3qft5Fq/7+av1353ZW0mP6nU2SeAs2m5XToJpIZOz7sRm/SsmFuprEb9ZPVNe1fd8whzDvS3
iJBtxXuwT3XF3S2wFC/Dih9BW62/2HArpdeBMAodsom4vNOe8Db206cJa4K871SDyblrzWY2Nxbl
cWZ8uyCSYccKsZlAwswrxHB5E2fIHYLxp488z1dNMSmNm/sBN0SyNf9SqP4Z6NB7pd4xC6m1UkAZ
1wGhx3KxVOPEAElPOydHIH3Rjh/bCcp6vCU7Z7oD0RsQLJXmX0s3TBhzHxGTpKMJ8dTk1ltidBp9
ec8nJAEh2Grsm6W1S8GTZZFKSxXUk7gTiyMu7mVfsU5FCHmAgL+bnV/FC3jlIzOYjSOYXHSzc6UI
sp/tho8N64D+k5NTEVa8LpPtgEkZdwwGyBg4sZvelrQGSbkwqSIoR3f6v68pNDM/v5P387RA/HuI
nlFRJkFJICkJIWSRGKuwMtvyPRzBt3e1HXJ/pYtJlwTqbDan1vx/T19vFQpJ5XmVF+g5iiFr3BZj
ghUY1YaoARD5OnkCN33Xs1vrEya28umlirXAsWtWBGMsl/AVirVWZ8A+zEW7h71GyoUZKQwoxalL
KkSVlFyIkSMe/CoL7xveqqbxGlLlx24vyFNxd+y7L9OQLWeYbAPYLhg1E9DjDHdjfCcSOvRiYm8S
B6oAeyit5/4qbaDjfROdVyPd8G4QG7hR99P8dzsNRQeE3El0bWza5H4SlCrU5mmxWo9n/q4T6ekW
Hs4TRxWluPG8qJ39xXdunBBp6nIesHLVOYPmqPN1kQA2wBy2IIMPCiSJJz8rcUbTXdtvdZmvR6Wq
biaPTJN8CxPgtRbwLA/0oC555H9zm76N5ApkK5g2q8XzlJeC7mHNRxEU6CudZgMStc0fIZm0721G
iaUPGORcOnzvSXgskUCzcVvoeT+X4VijqPZHZCf9H0AfPj6Opu9/EsB4WvzRsCsPattr2TJDQcMr
sFLmLrZElW81bkJ/hh44FZa54qpI0CnJ58A6qwqlSTkTx9InMn2wWjDSfFR4H1dyo7J33CNAtAFz
3iBAcI4hrEh+cKNCR5CqkXYTkTY8nKOjeQC4ZK449nYjeRKvd5hFu1UkheUJlwF2XStAoHLRaCqs
bH7Uq9eBkONxLyQoDbwUwZSTgHF4YVowcE1EMGHey+SLgAGzGbatoQ3VxC5Cm/5LWszUmvwBq57N
+jKWokYlnBbx9SM1nMorWC9qRvBur2rixV71O7xpqQDFnAsdK33TbMSruMyfyY3JUVQ+ZHZb5U1F
B6E4IJAaRhk4zOQTxLD072XW2Te7cfbCMdiukvgjSObzuAkZxyDxCqhLaA9QZzNaGI/lygGiuXHt
wwZRBYgKME7gGYJmW1ACuPdmo7SAFaMcmWIUCSvd6Xp0EMkwoG65ycUHFo82AxO3avklb0xOGrin
N1f2pHnDgqd/e6XwYkigy/D9fBxKEh1uSYABimVTqMcH+Fa/KZHEdeJjlIbwibdls6eb0QsYKO1f
K+CgqHe/MDlMLpg+o/66lWhp68aGKzsTyA5Cajjl7bJPSj8HqN1l0wScG8dUYBD38bItD/2U6nIg
MstJoRiMQepQ5WZntiGGXHpCB3Hup+lnpZDCvFy1urYC6i9q6bk5nMPQsJc6eTZllj3qb6XkJe3T
f7zNXqESLWwBbSpqRYTvn1aEwS6ZhbnWdZn1WZNtesCvIURLbx7aNPKSlepMlF5+/3vW6FigVk5C
x+75MyHTTkNGiLef84bM95TXqeSms3pSdue0WC1+WtjuBUimZbzsk97S3yZk/RB+uN9dSpHe0dj6
P3d8ISEcOKboU+FfASmmOOI46KNLLI8E6Yyydxps9/C6sbNDRgzZCJGGFjGr/R/4gth2FdUHDyUE
18ASfVukKEXlbm+XbG2xWtVCjN0Fit4+FnQf59yInCwR2ExvkG0y25HfOSzJ+ZrfkjzqFoES/6VR
mf/c5b9+yrdcSmK7IahxdKu/U1ovhWa9tRvviyH1KrkCtl6ggNSphWf8Jddo/wUtPNXVYi15gFZr
D4YJEnXApc2udV43rUPis0KlsAPtQzFuWC2KthDxPGNBeSw+no69cv9UnnzHJjrZ1OI9yzfMmQHh
VisgleBjfQc/jFWgKKl7Nc0+ouLumjY2963CXPzd5EjsMRhA3TldPRP5NssTOirOWg7T/oglG28f
eGuLxrMA4lQfceF5V1ytyoNS4v5GiHyVr3+el8cOLCGig3NVRCgyunmhVWpRgrKRX7ZC+M65P5jQ
7F7wDKbgTw/mA5yHzmeMgnsk08GNrB7s1lbB8p8ftY1akbToomFmHYdkd5I9pxt+LuJmLol3+DR7
DtoTa0z47gjNvYXOnJOlTUI3lEWTSRvppTQp5mv7+h4F2scayxpNr4/K/hmcJVr5Eke5fkNNahoX
RunLaEzvDNsq3i2cD+44OnBn2K+DAGqoAlcAAfhzZB0/8GfUfzw8fq/i6FiM9XEghpfPGkUjfKez
ATqGS/nMwvpaPXqB5G19LDNjRtMH4noIFVoTsBIO0KNlHwKM+ZabVnixeA+ZoG4I8i/ZTHTTBe9x
SXW7YoA/LSr1qhRO8dPQRPggJg90cEOOLfA7jLcRToRiA+iVNDDAlTYnLGxox8+SBK3EZ+QTaMtc
jxDIz462YTukbY5QTMyBKzsC+zshmsjMZsOXO+AX8mKlP6x0yjIkfo7EMPUaB43o8wLL9lG2IxYN
l86+yvpvxOgOMTm/hRZI4kMioeLLyFqbtEtF7FogF8grmwEPncdOcvH/XNNvxWbThAsIJtbXX/d8
WQ1IyePWc45KAnj/6J5fwwaZE1hO/a0F49yuKvSb3GjuD3iZyBdkUQRjkx8KfAySHHlZujqXGJrL
jGVtBIT/fHjIhQDEwf3qYiJgzRx6pV+71qAdY0m/xe1zvwoNnMifVnSUoR3K2KMXvKFpQiCyIE8A
2A3Md/5w6c2kXgykZAuwIsObPofmD2sBmnmtpicsDs0UAC/mAJ4Fx5VE3rjQZUsuvJ2dua+2ScDV
juoY0ojjvD1AFkZsImxj9TGZ4fRMYSVzjKQVA91UTLmXSsFE+R0Owva0kmsX9JM4C26SV8YDiMla
2j5oFga8ftU7bkZeqXaiRLhiUm2El2+L0hioZAXtbn2n0Rbp3hzTJQuyN3M7zlJns2U0H3C2Ba9s
QXXfFVao0qvSDdTEl5rR7GxFYyHKyOCPcLMYBZgmV8Rmoi4u3Z47gWPPMFriq6OSbhn0Djf/WUI7
7zitRDwS0t4kBBtqA+o3WCe7qpZ9c7SxFWmJZYOPoF8Upb3rWqAE8hBwXWzbuJPH3L++GkYgOip5
8jTBA5TvVRBArj441+NqbeH9nksurknQRp6wBG6wTsJAjxt/T08ZmlND2FL2vgwthn5kpLSktccv
SIcgKkaILpXT2dhcpZY9eZTV/10euzbnvwjNt+s4gAm70eE1kHxOnOqqltyiQNQ8kXZdEIs5kzuo
uh4AGMlM+NQXjzKXJVy2wzGzklXAfraa984ylbhJzMAms+f1KWeIbMecSQ7775coSCcpp2qmDrB3
OVllcNVGJnOTA9/22v6uS8wW81epV5pxKUsCBf2C9YybQUQUT7IfXZ+mc8lGBbapXLWTb1bGW1bR
0xdYnVi/EqRbCADvl1r7d4FLtlW+ohyD5T8uRZiJQaCkbwzCnnQU0PDzoOyVUYXlWF8hHW7hKC0z
fVdgGK2Fx7syOs9Owd4lT9RsqINMSF1oeGvnnUf39YircLL7AuN524t19m8vW+Tfcpn6uX6IsVUh
q+5zkudpL6ulqJY6mIVNLQNP3vXKwh6odK81ynmRcM9aDIpFr6r9rxysdbsfMARg8Djz23NPUOLg
uaU7NrXIj11ofw1BFTARYU5ZTLjXBaqUNfqFh9PJKAfCnxaMB/BBISiVDM6km0x5iUzx9WxVsCxQ
C7mKBmcYUIHzGM31lxLFrDdzQE1wcnHWpB7shJAKglK7DiOJGp/uHGz7OmYhJFZwyWP/g9qqWfx5
Soh4PhNaCTl+Jmj884qx2/uULLGvQpRAOJ7C9zN3ReahV/Y6W1E7Nb5ruPeEaZ8yXw0o3HmamWNh
Ew4DdWIb2B/1znd6F7yY1KK4Yd+yEx3xsRsEcxbZfmQFBEqJAc4gixDbBpMqrM1DGD4OEW2chwlY
z7/3n5VnzIwy88j1WajRwDmg9yqs83x0In29QGGZPbwNr6d91AP4t8AdXCjr0iYshGSWA0ZwS51M
S1TW0ZViYISGgEfkhHNwxKDZLXJIfmpyBnflEIHwiE59OWjOiFlmaYadAujjXkYgRzPmckDmOO9c
WXBTAwlSSrn7/KKYsHZS8IdyhAhgRLYgARGc0ZuDs/oEarNZ6iNXOZGnqz42cXtf/4xHzNN+xjps
92U99g1rMriBSXEXSdPcs5M0kD5LEX+87d6Sx5BMxli4taq6p7DEBH5mCmqqBg/Anqd2M6klsANn
1aJ5JnLX8M2j7WvSVDVVCFtadSq29DctiKI1Kw8MQYWnwp1gEpEmQKf/cWo18hcpeLgLWhaEWONU
ZW7zZq1XqP1sru9Ncdo4uJvlEkglkg6r/RjHib6+JDYPnG2aqAH/AF/ou7Bpd6hkIRWYK2fNFOea
v47Bo+LFDBKgoYrxYkFC5ZnoQSD6TBScmOVqZleJbjFUQA8So951Klb0+GKfHiEUU5aQL04hdwZd
Gj91Gxm58uZlWanyih/ForoRUpvm/gjCCcNFp30NguomQq218P3zUtBdk1+7pJlGFCa3uKGosT+K
G3XfDQBavEuW0Js8A9WJwAc91bwPt5qtRDbFy4V47qQlNGYdD1fO2xRdEfjj0uk9g0q4R6DA1IXR
7h920qIblnJ+PelxBBw9WxqTq5iJpYbQN0pFNu6VIOBUto7Lb5fOg3Ou1MsNSMjH/DIVigdHSW3x
+WHejE1ZT91M0wennwyK9spoVssvLjbTiNq5tlBnD5APWIUXgRx/4hqPXiRpvaT3t1d6aQZIfByM
KsRMWTs3l8cQoicTnp2ZlVoDxXlym2+OU5rRVKtm/e7DxRtC6DgS1U3q8JZvhZW4QsJ96u6hVZeI
omX5ecVC+mNyJkoD3NIwEkTr2xU5y7OfjeB7P0517CG5gy1r2lLlkKRGNejPmawjUCbehEF20W57
+GhRAXJ546bs6dC06QNd3z7KgYr6lGsLQGi4XnguUjJO8uhKa0nB90wB/MD/zb9UNaV+4/opxRGD
1p+uXBBvPsnV7aGximIq9ASDCvXgQxERbQT/ev322xrkNSiV9MP8HAwEbNsZo5se3LIHz5eokmSX
3QBYlSqId21e3nnPu0l6wtQIx2mpBPaxwnmLSW35S+Q3RH7jzz2eeDrieVNbcE2/5hD3I4wVqyyG
yESFT7bxN3YrM1wuuT9yRzVO3oRyCVsyWGz4weckTrzZTkC7diaM+PQUK7VjyWYWETs5ZLSYryaZ
ZojEhFCCdAcEuHnVMqHjU7l/lSmGFNI6Euz8W7D296yjTv+tRQxmU912VCdsIQ/LO+UKcWO8HTno
5x8DIczGcvA5asULMUf7DtQrz09rkK/30Jf/qIWST69xUVWsctsi/G604WS4g+9o8jk3Sq2Ozans
bg3YTi94uOUfhsLij1NNY+7t2JmeF6Z0ng8ZxFuLB4BBBVX95ZMAHd5zaRf+4aWHwXHQooSGbbA9
QKKOXuFul79MnZUbFEkb5CTdGWoJEUuoWpQK7m58oCuiVFkuhdNHc5K8zUB6DloUyAh8KhZVfV4V
/s0LE/5pQCqO8mh9jOsoWSy6/Lhuk+v93WEsVhdShJa8G47If6kKJNotIDH5iv7kycJmxmVPhOAx
QelhgNj2blIhp+wAWb3LjtNUhaOvWLfwr4a6yXeSxL+W4WVkGBKuwn50fUD56YU5xMAnfVXoBfgX
nE0XA/kx+sHd3DoWALUntRu2Bi3drZv5phoApfunoQpnnFqUDn07hWksVF+c+CQVE+3BcsdjYyMT
BY9EZ/sEgJaZOtV3tVEgV+KhARFqek8fq1t9x43sIqYISYv9s09AdDUSY6GNLuhchq0wPA784SUZ
8HL2jXwCZ8sJwQAs+ux3JoILzfokJWOcZZARoSkM70V9YbMl6+UAh7RPSPD51Zndfy6q1kHzH1FF
z1lpPzrhWdKrfhYT8MokUh5SgjftiDLzWqUthSzCsD9QDGB3DGki1/KfgY2RWvsakhQs4Oe3PtFF
Oh9b/I3MizcnU3Nmjr4/WtUwa2yUhBH5E5S9J3s1g9/GfnqP7JpYwY2Ixfbb9r7uR3uoNZ4++QPt
wreLUEb5p/cQVBop1rzN0cVBbT9VGJQSaH4mMGsu/6UsMf44mspqylnyb/BnJBymweNMr4MmDAAP
Ebuh2O8QGu/m7HhG0EaMaZQ1EGsgupfZfcgYdoB+adCLkFEczafFpW/wG9m60u5PusTFfA8dvxxi
Sju3QV5YSBZ3Juy4x6BVhKJyxCeGscfQQ/HLTtlTtwov98W/nkZzSUSGEl4aY7Y7zKXHy9TdENh3
2OPdYepyKa1qOzG56+4om5EiW2ut0eagms/vMDlWUpdcBLEbU+QANM0tyR8MeXxaQpk6jofGNo5o
QrtP3KK6j3TSu/br0UY+Yiq35CSnNOqi3nx9QrhAqt7Yw92qb4CxlLOjQRJHWeY+8tNoDUV5wK5k
FQ1bzGx1oqx+i3JW+fAsNTkSMjwKmEk+VAurOoWR06vaegnFfTbiDr5btnE/DnAz5vX+iDglN5Aj
rkwLqZuX8g3c7DWvL8DxN02zdIobaEWAuwOh6akpJslAzMi6ELFZHinD9kBP4FxGN2YRJuoZPN7H
odtjc/yMtfysNBUt8KYrf15NrjpB5BIsGauZ7MDTNGymgiiLBv/I7PH6IoT3jU5S8+cdKcIK2wiB
ij0jR4qrAbrlxz3i87h45FhMKLIF+DIQsyS5VjavggtzlQ8G6XUZa9wEPCFfJeh901bgZHtn7x9p
U6LcG9e4346uPv/VAdulgkX/QzrF9B2jj3GhFcZQOK0Hvrq8R6j1cqS489TpfieInnh7wzJsHNkf
AWMpyE6JQqNf1lALZguW/SWfEoCfw2fBc9WkFv6W+IhR/fjbCy7BRoPKMrwgjV8lAAxuZirlDYTU
0UC7DHE2jJebEnpyfOjVXEWrHkH97HLkS5kTrosw26X+lbhgILvl57sA247VwyJ4CFdfPUBJaUA/
jKe35PVZAm8RqZB2iaKP/gO2ELKKkddkJ801cItyxDneq+b0oViDWiwFiEolR9zFEUll2ZW3ituF
vJ0f0GmMHdVmwShgTlhCglMjxuU/zuadxDxII1Bt7g7KyUXkrPVdoOYdAyTkHwu8+15y2r+Tnoej
BgnW0mxNHPqNt6dGjPDTPVj42EREBLA12xKHwkvjcsV2lpLMmFB0LG3GD+MkMoGnJNlSoqLMO8iL
ik7s/tisgiHyN0bbC9lw60t9KEN28k5OY4banw163RXA7vZOYygGwMjDt7nQFB4t+OfMNtgn0NNl
4sE59Of98tVFLHay3WdBrm4u500PH8riEobw1iBBgASUVSji0n/UGOCFcG+Q39Tn80Goyt2itaN3
Y3vLDnItbGmxvFE1eAhHHO5xUSIxcGPQzsNV8zpK31Z/k+rm2/kSxLj43mK9RT2NpnvhrQ9s86jk
/bxkzuFtJy0s5i2iky3n21KLq+Q8PQS7dh8sc6tGRjuEXYEbwJ3Rw2o9z1cQULm+eDnlMHoV9eVn
qMqGommCP6YfbUl5bwl+BR93I6yDk3BdPK+AZkO0/aULiptE2MLrfdLVbSnqtWy+ZieT/MmNaLmM
VKzcd6fM6l2xE+7dz6TQKex+iua009KdGsqrVSFGPVVPo75Np9s0BrW9faHriIVtBsRfQa+deSws
kwEXCcljuhc/hkcwnbR1v8StnBWplmfKAIFElICjJZJMn78jXcA5Dtfg1G38iSi1KxRCw2hvdOSQ
OqOYU3OtyqXf7bknNFMlHBrogvTGkz/UFJzrQ5NagYLMzeXlFCzRBhwOj2FVQ+cuSlunEAAFaadw
F/7xIPdB3/wWO/gmCzv6hd+ZjCAZBoGnB+dw9V1cGkzd9pDa/X3jKYH4ZSBqss3bP4iQHDBdtLFC
qpR+LbPoVuzQe8MTZEbb0ReoCyftqeQuQIz3uFYkdmezYikgf4rGoVP1KSsZjdjfxaeVrqRlK3xW
3Ys7K9bj7LuiVz/42izBAhhaSSAmDXwMJndtcVhu1k70blqhhyDfBll/PfPE1+zNIuXA2cf7ciu7
yTf3xk3HNmIZqf5wNa//wwBAb8R0xhq0yj3RxxjnPAcqgcWn+jLvJAGczy5lMScomSsfjhEF5OfB
gSWiPSRVWJiDQmwWPv3z2yNVT1lQGbaVP4eZVOlswAIDWy8uptpiuvZB+dZhfsi5o+IqT88k2QHf
ayD8AtdACKUv3aGx9USH3ylWj+cDq1Fegh88fwue0kXyfCdBbdoe3BKNkdB7z1vZdqCKc5TVETui
MoqDdxRS/QLwAp3YBJNLIdzWtw/Zh+4jSh5V0fIJVpckhE+ZVy7Sc8BicEo2EBbnUx4/67PRZKem
HDy+dQi0Ua+HjcwUDwlf+JQKn0wyjqj2at0dVpwOO4PMjENNEFERHLlakX7hhfCJ7ctN/3bLgAse
0fk/HT8T2Km82WhFyOaZV1UBDFc72AoDW32dObLPMCqao61BiyUul5++SxrrSo51NRH8oMKSalYS
n4QX01p43/VTtsWC6fIgOrIb9Eugux/fF+18fsFW9qakLOLsF7P4XpvwihKBEOAbpYC0mB/vbN5E
dkyBl7v/d8DhVQrYaLpzj/sCM8pswWy9iwjhCSEXuKCtQTpRC+hAQfjXb2sjFkUPcF1NmcpcjrJn
/PvvJO2Xh8EUfOrRGX1UbmjX8MiWUQlsJ0amJKv6u8vpW2zDjQbfQL0MwN4u/1eBROKwBffwWf6H
yn+/wCILzaOj2bKJLg6m/K4NBXA9LjShI1patH4k/lG3XHOXX5YA6vpWfSS1QYicDiALnuYCXaGC
E1xBZx2wL5IwJSbRYVdVUFF0CLn33cpOfCjc1dqx5Wq270AKu+V6zaLCi7vFe+KYkP5XOFvrUy94
6eghBzQLvBI0+BKim8Q0l5eXcKXw6Q0dVUw8HWxzSgET3yS4AejfQK/GKD92ETZxD2OArYTH8uf5
QlmOQCAecGwebyJZc/zu3bHsFu43Ym7lfk1Z+KPnDI5DwZY5FqTTM9fO2TTqqe/HLYX5AEWArL+j
YlCa9v8GIbu1KSqzJ6qHd9puiY1hjNWsjHcjVBQNl0wH5jmMsISqIYQYSuKP2MjE0+1fyvo/lpxx
uKO80MADiYqzenXBHH9KrlokZG98ouf9xH/mpS8LzypASkYHsnb3dmT22cYhklfBIXzA/Fpq91+H
kRwx0nrJw6816adMcBl3GOD6RsOYyVhRSCmLyL4Dk2+HApeyoKv3CPvhhpn0OzpdWM98Z2Ki7XHe
TVehRGzebwH1QnJj0xuBzkEYcOFoJ5RQOVitgC3VS8thI+u/OqK33XOTcmvJXDaec2+o+3qB/m2o
1eu0NCVD+edZB1/Sj/w4SNFMCJi+d9JnPaLMPDhC/Wey+J0CJN97A0MhvIJkwr6RW+s5mQPXPfPS
pD+7IdpE/DvTYlezStApNbqHCmRxrNaT90WSelsAnzKxyc0iOCLE0DouOdpWCDg73pdyJyio4WTc
FcWMInbVGMG89zVlqmRnycHN9ttYfCwxsbwsnE6bIj7h6aNaOvKZtiMTVrrv/ZTeUg/eubQpv4dx
0dNtKnKBVQvlOKq4k3+BUpvC6LGPoqX9hO+56bXcNNqkL6eLhWfF2S+RqHExSnIpBnDPXiA9XbLe
IbWDJoi55/trQAXcDCaFRhjQE5UP1kTws39lEixtmMoUhaMTmQvkrfplW+iLRrO7lA8S2uJMRfye
omPN7DHGc+sUxgw/JeyrYog+ZPv5EFvQoQmcpTRVm+kttgm1s3l2U561iCikKIm54Gfb0f+O7JjM
g5iln8FO9jmQ5PsOGYkfq3fTg1BE6gWrKwex842adbyHJZGEOkNbzcCsyj6U9nyeX091DHx92kkP
gv6+3l2wNFeWzrY/b6FTQrRdeERF7G6VwC7zqxdBSHjtmS4qO8rXBQQg03JBqnlFbWkqvcpd0+HN
qwI/d6JcVQoORvlQm2y+LETsA2nLQd41LPAuJh2fy/ADVlQQ9q32GG9CK04RV9YD4vAd5A+YyhbB
UshzghGw/VRkcKr27TdcG4XYeqfglaKOmjBohhrLP4+KYhX6k8M6a29EXNlniGry0USW9aYZwJK4
n8hBuRNKfEW2jXxyJwai4Am6SrpvTOnCNZ5sVwStLFYW6I5cu/E+q04ChzLFU6dlUFIoS6n1psGs
P/f6LlwnKEgAJ4Gdp0nPumfQv1l/TdckTVljmwfnJRYlCexA9snhYLAUa/eZLVTRvUY15yj+hi3n
VxeJuDCeBP/NhLb3MHTKaZnZCkP5OkjPfJYLDODwpga8X/aFrP8WXHflQskCffKtN/xbSI0stvA5
lrWlCueWke2jScVSLd9amIvGs3/tDVpoFYXthh86bTRy/+eWgVbBsiR/p8FehKxDigRcz6LhkxpE
xFpFbPn/k7wj+0k1IaHpTR/RC4evSjiu4FCW6Kc1S3w7/Wz4ntiq/IQzZhmq+Ib0hF9/5dmy6wo5
ef0f0TpEN51qGnFkTmOxjGgbHQDeFlgibFhwDT8jTI6MFSLJ+q05+PUGWIxGpnmLT1uF7Fmw3KRH
NVp++ayHPj/7CrxBEEVmXBG/Fiu4wxvJwq+0eZttfM/TqH2bbUSEVS0y/bQYbmL5AOH/3LCDZ8lb
y2AY9/H3syzc0GeSGbjZDIILWfL/a32LaiOH3I66D0+nCpIAHJJGo36poDnLUyNu8+p/jxl7cAPk
laacC/dV1htEeR8Y3aOHFbylbLpZsoZF2+QbCmrSsxmyWPP9Zedu5eg+w5nXh9Ole3/Gnkf44hPF
zrt57n7t+T9vS38Wbfh16nZieRqy4RtxyUTKEJ4DOJCsgidAzz/aXOetqfxD0g58zddQAIduTKYX
l0m14mPntdCe2RACKSGZp0ZTaOaRyt9hY50VDMSB7UhyYx7zaJjFqlcjB1qxQFCMdshG+2D+Ejds
RFpWMshlTPeuwS3daDx5jkXPwWe6VkCnXpMMJzarY8cGJVGj6kusctu7+kuZRdb5PFpHANc0oBz4
llYxQW7HsoCBbIfngY33jJ8BpXEorOHMucPT32Yoik8vJM8kVkAzWwBz5F+1pNG7dGZvmszJcXWG
sOk5GoM1rVBBYkuy5HcoHiui8E1rBLCbFI3Z4dTejYRpmglASi3jxBDE3oDe1tbnSsnBLxUCHejn
xcNT1j/l1vZ8bBYr8xsOLiWn/4lQ1ozx7RerERanSfgXR+Dhk2tfWqya469JC9a+JhwsETnFJj7i
M4Ul1rmNKGXqGoyNLKjyOxYQL5NEf44/ILvxMZqG5oe3QfVuODMDrg+rxSyTuZVVLbM3Vd5nLEk3
Wt7Zv4ktOAQ8QU16IE7Gm7qVyWH8lIJpBqXh6U+bNC1g6a+Z/78kP/RF+6y36AWWF4OXDzqaHSYi
pBFqj4dq8FGnIqQjpCD1o/thULsqvHUxey9cECfzXGEEvzdQf23peVy6mnuM+CF2RaoMtpQ8PoWy
JKSAFdKQ/oBidVfSSlan8tCJ9KcY/WktpY0QrgVzGAGh1K5bWHnLsjEiIMbyV7e68bMXxNGpnhqU
88qZ2XimyeZ5p4rYN6PcMC5y/NZrGXBww2RCeuobg+nRZSAY6P7PCRysAkWHPdqexoWfWCL9jQrU
/Aaqco0yNS3VayohhksatTW3klk67FAnSJy3RcIH64xVv3vmT0fIDGOgSTAQTHZycgPBsp8pcQGy
koZZRUX50iX/jp1MGI7YBi3jxrjZEBaQxS/y+EcHa3YxY/R/UfnxBUdBJz+PI+dDnoT8pbrQbu0c
ysIHohCVqoRJrKJzLg/ZQMpVAu0lkNIhiE4/nNaaq+FVUbXYXBi5DLwrvC5VO7wH2RPrNeVBtml4
UfvBrcgKzRtnGcn/XiULggyFGuz8rIoPpMqWRA6w5m8OxrI+NBYSXg5wg9bjy4l5pdTFADz2ohwZ
I0OEUBmvlCtc5zuIEDtIVcafrzcQ+yN5E8eleMK6HD5frOrbtJdhmP3QycXP/yEPhM6hDc7krs83
JvFe6uw9nFFN4I0tjA5qL8lDlZxYnb3WYshQj2un/bdBul3KuZtJ6bo7yNPTFu67ZH4IbynaMVT/
xk1RzbJDzcOJv5fQ3hGh1lqd/gM2U2PQHj6RHOfqrpFhXJq0tmO8X19Ew5j+3Wz5V39fRphmrsWX
JUHCXf1710ORpwUvYbYZ6iR3ze7OOXFulYOeU874/eTtzOpbuAfD7eETjF7NhEcuJpfeeM3yjYP/
ML3i+MUzoh5MzlvTTLEBqCQTf8VNL9FsHqSKPa89JjyYyc4SLAppEIP1Dwb9QPAynQIXxml53tgV
KCJnja/JzfOXpklUkD5ll176Uf0ySNb0SstaWxdsiPvVshkq8yFGeIorYfb8zaEQ0++0PNcyIqAH
TW2n/hPDCQ7mYv67lCL7GS3l8mYyVWVR1PKkB7i/xPE0QcG+OBlfPGCcql6PZ1RC+Yubngmiuqwh
YHvp/2UUbg5bAyvOWpqriaPhPHPUP6AdwiBN5XkejazyQJzEjmcoFfqgta2X+yg5ifh9QO5gzXZr
sdLudgvrRVChFn7IIu1p+oySMihlr3QixBz0Jn6WaTb7s//rEIxcI+xdoJc3/NDtpcA42IWfz8lY
02P2ByxXDwc4Z84ItSt4AG/QizgCDNfNXPUgbHwTxTtut/y88+ZDUu30dr6gLYRWX/huB0I38miH
Rc88YTodlqk60f5CMC6J6T2bN/ia6/QcXIsxLDSTWIh1wtFVKMwbCvQj9lM+GkzWpIdMEiIb9JTH
6UAX5vrVPA7m8pu+cy3NPJ7XKxougPjrtTEV4a2NPb/9ZTmSiftIMjSNTytPEVOMBiORZG3nTwU2
Ar2uq6Sb4G/I8jt0woflswiLmrk60KZRyaOkZsLqhbasRHIlm6CN6Z/oZbMJBDpe5xj8BUGaBGXM
MfxUqwS8SSAJen9If0zPiv3xy/x+jaFoyJK/kDGonl5Lp88XMB3ywES0a6tjn8Q3qLUQlxbtezkR
CT+BHfRjSLl0ZB2b2uvU1CBUHFAmzFl6BvTg7e6nxfy+p8OOP0Bv3TBdW7Bayhevq06tnCVI6c2J
AGQRYamJEPovGZLggE99QEbSwu/0+vsQxCT4L6SsOdZvknPO5syD+ozRoUGOUhfSs0SsnwO2acmp
40gTvuZCYhRaxZCDcAh5sEBUxk1Jz1Ettwrd3ojlfctxc+3I7PCV0BwgDBlSOH0VKcVC4gYCBUWq
u7J3KMPITimZGBhM4JMuX/ZUnKOZla9SASZUsL4AWi5Kt0mJ36155WHw0kank1AHJ7dvXVKEkqUN
RfiwInOYnEgol20nWndnRd7IdXrdwbMuNgrCpgHgTu31kwgrQOmuEpnljlxQrdJSB0uto1Da4Y3s
5DpV2MC9oevGfO5fa7IdfwUWhDx3lDS0G+mZreSLtNoGbb9h/rzy8k1Z8Q/cwiv04MbwdZAKyKzA
hqIBvpAZzr12ikNk34BqKBBwGQfDwebmiNCCRhrDhyqou8LHaFSnJHSs3Ox9+9PJw3FPMgIkBA2f
fC3LSZLzvbTk+ImIo2lqq43tlfNCug6/PTts64Y3BovJ8Bww6BZSEtgzVfX7MM+ws5k/LFPVhmQ2
MP23LZUk7cGjU7Z81LUYHHttReevvuWtQUZnNgpShRBdZTro9OzzIcYrs8cju9vb9tGI/Kwak/hK
1/B9gU1lPqcjjpB5ancD0aHx4FF4WwQ9p7mBYFV2ZG7aOKPQwmjSDDyNh2iGuGH1FgoSEqcPxwnO
BHSBPyJYcNnG3VUJWsJ+jx+9R8bAIkJwtALSmrZvXFaDSPaDcYmJiGjya+vHmllbTSnmapfhWrR1
me+pUDOtk7+qQIJZ2fz6I1PXPYsgY8Khy4e/pL4LjuJNgPYDgEP+aLF3PwYKf4vShV3l2wWD9RSh
/nonGDwF831el6tD+kmib52qY9MFnfKlCkfhcfDYDsHKJh77buaHCz6cURWV7lvjsKctUksTlhBP
ElSvE8EMavsyMoJs7BuTq7eOaQjQuAVyLbS37UTAKncDqYxpv8DmyAKtE3OY7FL6H3Q2OfA2pTo4
61wnI1UqMlaIvyWz/paPZ929JKOdSu6ZOvDo8bJvDi7TgwMoiM3jHB0RrV+CQ11ghvLcwIY6MkRe
/ZYyFspp86rJzokcbGWu8Qxuob2pa3pyWfnDXb1JQDaQKt1L2HD7mIpNLfVvPXU8InIiSj7U99Qk
rEnenP6o9oelf+nGUB4O9jggNpwY9ECgiagEdACf6ibarxbfbqsmUzJ0UaDk2io2UDT6o3bn07bf
kCoUhMjV5wlb9iQaXrMngwSw5NB+IZhmIufnM1dAeQk3O+GU+yXcg0rsVrwjIrfn+QGsmeChaQIz
BdG7AvcTxWFKIDviMIn2qVDYJ07D41iy+MiQNqPMR29EQHbGq7VeqNNAJk6nlxq2j14m38dT4ESk
VcQV2T6jyzCCix6i+FWgqJ9Mqr3J2PruJwg1fpC5Np5uU1U1AtpLhLwKPBFqZtmR016iIHDmzCHC
JvflY0yhg/BMEgRiwGhta3ffrn2/ZxviGcIiLbenBLGPD6HoCZPpb+LkjOmiM3sPtJA98nofaUqV
pq/1+E9JMZ0NHMRHeBYH/DwI7QyN/G68ZYV//c+V2EkL/AmBRG4zvCfEVD+NVTVv9oi+xLorNjcr
wFeBv6QVVR55PCECh66AwEJJNgxI2iHv5/aGc/yELrTPaYO2oHGDOacT7diqxihEROyhRxQUhO/v
hmQliZWph2LZwfWT2VfNnwt4w0NeTgvsN1CXCDVGbeMaVZw45zwv4r0sLIppcb4S8l2YFLdCrFkC
rHnwXr0PHqaSCplAYG/Z8Zq9O1DrRhhumE5S9Z/55lGVaKNDXfQhKGPgOtdoTA2Ww/KGmWx5FIVk
PWBlITId2xjDR5IZvxb31ASuxtEjt4jJJXVqkAcuB1QfpJru8SrZrNfe6cJ99Mnq/K+LT0IIqrXe
2QwCXp6MJDHZBwZBffnuAxXAqiHR2+Tzq0+Uv58Vt42rB+BaxdJNFyg5KFk9Cg42GlHQv1NHmX1V
GaAunJMfBHtKzBAerq4wizfYfvlHixt5ujiIJWRDOPIKu6INMOoAb4z8+FIPLPprf+FfYZhUy3BC
UCoemtNT0ClsRv3okJ6T9oLbkA6AQXuy3SE/UyUYkKpdvwlMw94o0ygP7gcMTpwvJMnI501ZBVKN
CVCXmxWtIcL00gHokm3ko6aHAXTz3FNlxPmvxK20oojRQzYkHLz/wXNeB1wbzF+qxSTSxQT1/NQD
iCx2cVV/P2z+57EklON42pv3ksCZ0xn0oRAj+IH2S5khas/55OO51Wx1BFUna+VcQ8HeDt5/n0PI
u6ag082RkICQYbIoiLwbsBqD6JHmGxDZpuTFwLaua6KmKI+MLCyuT6o1EED6tr3uM+LGfXRIn37Y
HtCzQvF92fX6S/NwahKf4YlLiVTnXiIfHfoH9PcLfRON35D9tcKt9n147q6r4LOyozdZd091iV3X
AKPWkP8mPS2IVbQOBJ7+nqSjitjhf0/6CzxLmP9HmRglGVKK02UcM91xGez13934Z69mv2JOsKpX
AIL0/HFcruiqSBzswGikFrG0OSq3EwaX3WMZBuIsaUSB+uJ+8DQu2DKQjm+j24TpTYtU5IHKVu/+
8dOee3LkgNhCFvcMfLDuUOO5ot+S4W7ybLfeVaDX4RLpqHXbSwHC04h6XE2Vf2au9akilMzNmdUR
0k1pOXWdkrPUVILBSNdKLPRyUPZrQ3IOqexmVxiMGYwvXslzNrwzf8Ygk/lEEgy5k9M4UvhvBu/9
wl01q9wxn0zYndk8IbBLxHr6YA6xAoqImdS4nLJfHNZwTXVjXXPAiWqe6t8NUUTyhh2I2JD5T3lF
72aifSQPmLVOaOfbwe0MMB9FfQTdicJBA7A++qhMHau1YlPamo/EHzeSNdMr5STdilipqFr8fcEz
8+bBqsqblnQyEylS8f5n2/35Z/A+rM9XGo2vDALUV3b5L8Rj66RMeILLWMybaCwNBWNUep9ElJYr
WhaWT2ZZFvNMhxYwZapj/ZE2sfTo+CUw8YfC71lA+MkKyaUFp73uilUdimBfIejDTVu39IlIRF5Y
GsDsppnWgl7UQHvbEb9pr713/t7cYRbsYcFzfsbdFaMKHc148d5DFz7faYLmgaJoyvojgFaK0Q/h
39lJ+/kM5lb0wUJ/C+YCi17ElaUyoAQdUpvFp1wnAmtL5bqNfHaqQE2hWWt8M0a1rhUpi4vbKYzy
iojI8xkU+AmUfol27kUy3wN20hACaXzLhPaLdX2XOp8p+YK85Hq9t35Z/G0QcYf+Ke9r11bbwGdl
5jZ6Z+7ap2TJrA8YIgOcUjKPnoG7vnslMCw92qA1osn1XWXgImwWLeX84Fcer0BJjn5mbmtInAXG
mizAZsKQw9ge4seTOhwQRj0K+YJj5sXaeC+r82bm3pnhi+VPhD/SYt7LJ9kiO+pxVkMCd1MiTyTV
WnmRoRBCGt4Jx/lSGQz08SUFnlH2tOw5EuwHdjCcwAcLNSsWSnTidNJ8f5PZBi4Z2RLJFGbpRZnJ
e83OTGUGT7bIlnZly0GdFHM2F2PzDu30VvdYgLkQR1iVnw56fAirBHW6ex27NIMvOy1XRtrItRHb
t7dVQsQX6DLqSXk+Qi2qC5xLBcFGgxQEqm5VhVNtj9s3fkX3AfIqmMqVk6CE2hp7KoIkHv9WCkUN
+SG3CkMGi/vndp8n2vPCAO0v453dtUWItALQP2JfYw2dsxy99Wpi6ifonwdTSo06Pu6utLU0SKvX
7bYGDCTRBiaz8wAl0Kb47KVAOUmFC/4TV1YaqhjFYT1isTgF9fjEEvPPef0nrgrZwwabqgG5Vqca
PVI97LPBUjD4t7180DIAyae+gZjBhP69KO7bYle/3zzQYGMQMvliELkb/zo175j9gMKvIfz12fVc
CyufvV3Vd/oo4p3wD87M7Q1hJY/9ApugXk+9mi5q/wT6f9BKyDhvv5HofHH9wl/zC9qtUhG8pmyP
urJPzkabnh/MlTNUnIp6//P9MFog5zKtFc9Zw/CserxXMPupp87AW+wYuQ+khUnUayN/NTTKTk+d
lQ7K/oHkXF8ZAkIQbYfUtXfSRX8mdWpWwAr8py/O4L/IrsVYbLuAkiS/bvr4UqxzxjsyrpQ52iIZ
XAQz6+OYMDaKtOxua3U32OM1MgaCAp06tglqGxKOaeShIaUTR+M8MX91JhwGVKsuE0ZWagrPo0kk
h+/et5ueaK5gLsajMtyf3bbkMQY4BuI3Bcq7bbrtPBd0zOvRAyR/YXXfv8NiZ1wbhj1futueyq44
8qLxXjva9cMyAxQEmWfRHdl5P/l9U3ctKwdlO/Rn0JrcPBb64a66ZBAJdJ0dozq8FyTSESGyd4rI
DWKEP+LaOS/l23LrIZc+PQLuj/kdBzpSPPBBFjO6dzzX6T+YwyUmVT1hX7rDaiXGM14AmiSFgcT0
qMEQNBzCztQVSWjYRuW3KUWfux8AkSc0c0m8H9AnBtvHt5jL25Msm6ecmGePZNaxNGdF0uzZLr3w
JK2sj/oVD9fwzV0GvnFXBiMyHSLYh4qwW5mQxpoZzJEeh3u+EYUBiUqRb/FvS3OgFQsPtoYrFLD6
vxDT6L7ZUKG1hqJZLxK/TrDcsQN4zVBL3TpnGNJqnFAmS7S56efRQCG2tQyCvqkU8n4E6M7Tu/xM
alQ5CUlAT+cEcMGcEdjFhRjRRPgeebBBP8LN2j0DtCryPCC3t12aC5grtR47daA5weSj9FleeWgx
xiwXhgX97gYOxDeIJw2Fckiljnfsssn+7AzumFSBq6wDjVFicX0jZqc63obOnDhTM0j4G73QjJSF
uwW2zIH2N9zIz2AOh41eagC2nlPociWmvJq5f1wHn6/ccVqo0+wMUU93HfoMasf5m1y9xUZzLYjh
3DIO0ztaQcaYtOXOh2tLmlzyrjteytzAzGvcKah+zlr3yh7YqjE1t95HCkCI2qF1WLfo7p2R85DC
k5NaoR2Zfp82AIxmfe9E5QZBdPKPvO1SuRdLZCxYdzZyhFIubigSBE9jfP5LhQlHjAGUkYLm6WnM
Lravj63x1vgrMCKqs6rdoqQWuPnpmu4DKSD7QegHHP83jAn0tbeXzd/Em292Y4QyB9jxJuUs4npx
eubTKX+aSuaEwIqG3FVPyrgqxglVyHY6KhkqmOqjxkuJquPg4KYGehBqKrAUQQg0PBNNg5XcuBjg
4oxo3uYQupAok1JIE58nxVrVZlEVfcLihRqbSXWChgYQL+UgGB4wScHGrMe23r1g3vhCHmFJafit
OnZcup7Ik1GhWi7J0STtM6rrC/tTmOQfvIRSRTJtQZmm94RZFYKbiooPBROwy+kpqKI6vKo6yViV
DFW0w79eWTlpe2x8qEO460yudXdE54JEIMfIsh6+mP6DeoW9yvmBhB2vFtuv5S33Lr4WBi3mzpyk
G6MxFiahKkZeFpSmJaoULQLVlMYLxt0ZreEf05Rfsk4SezeX81Ih+DHyhlma3my450fwclGX3d4i
zrXCIle/hysjbXyMemQNxiKoMQN0ZzGcna1LxP1TPsRUWoxr+HwZa83CvRN67Fz4h5LoLM9GxAIN
fMiJYhsHgRRV3HzUfO7MDxz2ey0Dtjk8NIOT91xC1XYtsublMml3suvQkJKAjHK/fqTyIatfWzh4
AuEGg0dfawP8oRu9amh993s2+vOTEl2YdfSN53fRFKBjKTRfontjZsP8p3REu26VqCQwlUccdR8y
wtLLEZUAeXFkmY5I02JK1reHlmIOfTlZ5y461idJ//fi9jivJmeG8ibhGA/nyam7DjP8aBXPMWIp
MLxZsd2kyRYrIEvZYA4wUOQd0E2a4RgCV0fHAn7xCBXw8PB5QECHEGm/m3Oytz9tOKX/XKWkAbLW
HvZSIgLB8NTbNvnXVXMDlg5U7YH/h268iGPRxZnwRtk4FovtsQdBAly6XvQKENSh4th1iIyfTgWP
Y8mnzyjV1Fmay2ckhZuC2QL/mSHUDsn4hQeo17BgUNNzLrjixsWk95B0QdcKVkoiSq6jl3u9hVWu
UKZlDs94qMFA8PH+JCwqy+kEAq2YECBghUNuNKqRaRTFp7FedatpAA2xKNR/6sUJbQm6CxAb3DEF
WBXHDtAwCyQ28IMKonVNOjShefHU9Fap/ATGEKx2wkZz5vJbgzMPBbQg2ox+zCXk7U7K52QJbCGP
jk0yK7IPcxq4uGmNitRImGlA/RbF/ZAQwdVvFj5dQ7lm4TTp0vsRusgJI62lhsLMv0FeXptQK/hc
5kQopvLFiKBusoSIIlDuPb04CFW6Q5MTdI9eiDY1BRzbmjxvs0yUPiuj2178XhtSsw2bQ67CABJC
3VImbhcUtBHpzggBzV1m2OG6j+zef5i23nNwmzNwiKmym7TA2MnQIpPt+leN88z3FUvchLC1C3Bh
92ot/MqwAkOsWRsxT4b+TwVwXyVy27khw9i0iMYUDqugdlL+2mzjAcPaGKdWuLwSHpu4pJihJAQK
77ptRgRb0pb0+W1zdcR6L6nrfP4EygvBg8ryhVLXlf6ZWq2/8/I0CZ/pPUd5xa7yvIAE0RuDLY3g
JVtKo9M3wGTge1t8TrAF5YFAqaYEU8+Q7EW9cBZXaaRY9RfRe5gvPQy8MDp3zDzkRJbEWX2JGLi9
5w6Tbxd0OZtwH2XU9exZgAyL5ueEik9C8Vv1cX4FAJdz872x6uCotXH/mjlaWAoFLf4pAuA2pfuY
CAz2RQmMXVlLImGCBiCID0CkSawOrxyKppFzD8AEynEjVsMM1ISOuWroIMBRcB1c4VxiDJk3G/z7
W+CoI98qBv0wIfBKEz+l9XAg5ed6ePbIkHWvDm7aqVYr2unUONVt3N6SY/ecsFBrW+cwgXeD6cxM
/t69VJrqAOWl6noZhcgJ/RwD5KgCWkSce+LxBBpvYveZDfLMgLbss2X0yGAe9iV33mBPTefIoO7N
ot041m60AxJtTloBDKzc5FjDpNs4h4ISzMGdJSfB3Nn3lPhKcepx7uSG7L+9PxlufkIYygaOGXhe
XpSFFkePFRkfBrX/wL+UCYHOqYqsk3ozzmqGIQnrBKc2hTFbJz+ayGgypG2+Nti1+sY1V4JiN5F8
txFrQrKYAP50pvhYb9zwZEAuigzJT2rPsZN0VoEq+L5e4q5/jpjEjCCe9BGyvQUz5h734yuuNgxL
iDJ6amjGKvbO6gyqfz6M4iDEjkkjQgmJIrsKU2tDFK9h6iZ8dunl94Gro5IOTUWQ5oEUbMccszXu
ACg/H6wO9Pc1Y8FtiRe8JcgfBJR1tLgcaDL9/VczNwI1+jUUfs4KKF9BzDxEots1dsJ6ZSTui9Qz
WlrNAKIfjbh9XCeAPdSiIPYY7FHJskbb9SgkrR33eIhU3wdP4V+1ckMx3x3yg6ulbOd7SLubBC0A
VgT6lLbgWVZhU2V4VVl5idkgmsfIWk97C31ZqGWD9HF1v2RlnWwK07boQCCLYvaXr4OIijJMQcNW
HjST3t/1zPPixjQ9HKRMn+CiFN3Nmjp3L2MDqVbtdbnM/R1v6zauhC6xtbhJxW9N6v85YetatMW8
LnVEBlqq7YlFgGISZxM/FdWZeFjzvURUpwtKg5ociv2u9Ql34qrfv52IenTbqLPKrkdPeklp5B7s
sytNu32/P2wXFGLKaHdMHyhcPR0z+KctZ8EncEhEUOozgy7XG20Cv736mZHVCKSK7pO1Fjnb88WG
e/x955UIEwq6GXBFowVwheBB6X0lvaG6FdCHP2tQoWsNZ9WDb6SL4YrR101xg7Ig/rE/L7s+llqF
6be+ElKLascPPGahfk+yf7IK/av1wTlkE6c5pxsN7griE8H6/JT38kiOU6ZKZN8ILuvtMGQab+W6
NZb4Qdr0b2h/OsnKymLXHzrwGDrTen9mZB3QbjhmTy9stwdNh8fjz2FDx+fQYqisq6zYTzLOuNch
B4G5ee04RgFC9xcdwxRjg8CZNzf54Alu2YzFLvX2BA0P009V6CcnKLbqXdxmIieg1/le2bcERRXn
Yi3/FQmkWkE0sHHGftfinDvFugaoQM1FJuFNSQ/YQb5ZaSYDHthPNd5mD9LNtk6EDDQGz2AgSPGa
6CwZd9jXLOMlTitWC2ZNV2tApgdWkJRHmXazsu/ycUBmdospKEDUSFPtrdI7pn+Rah8iZhEthau7
1h93L+7Tzrna5nOFdJs38rrYe2JJVTqWYWwsffVYjr2bBlJN2FD6m6mgNRiIfj+/PRiBTldwx+eD
tOSK/n69SiIACov8jYD5/+EiXJhhJ49nlKQsE9voWVWiHur+9M/llHHCSD8L16Yek1uRW5AQMNlB
cPKBiuowycEN/Ls6CbwyWpY0f3ti/MOz4PGjzkrmMLF1dZ9MoR+AzyJhQvn6k6IBSwPW1BQjojUQ
ZVcFWQgfwCtzdiE1Y1Asrql16Zmoa7b5Q0lPbj57b8H02WpkrIZcO0VLNxHF72CFJfhPqnPL5mzw
QChzk1ag5jWt6a3tUAAELJY75qXKbH0XXk9L2TCFYn/XKl/dNf0eGeGiWfHUF6JDf1cyiqsBjJrX
LGmjwqXPcuDPChQIpQX+Er0/Xk4Xs8QKmM5RhZOiWAbYrwkWyYf0honRw07iwbpZoChNglwgWpPa
YVYERKSrMoyE3RfNoD6Bimm1+fgk+q+fO09RvZ1C0s/Fy6cnm77M6DaOXHWCkdKSZLuICfezS94v
S77/Sib+rBgQle39sh+pOe/oJoRT5YjxiXOzzXh8vDVOok3wm7yfx405DJ+oV5FbckW1iBD9WeWN
LSLhkDnUGy20JmHq+1gujMY9nruCU7f67mc41HGGHX6gZW6BdjjmfiHXDUooHvv9zWBy5lSVrjzn
HGfJ2dd/6PmO4L2Tvpn8DYvsjX3PzTghAJ2N+UXot7x9v8GX7mt+Qwwk0O3wgjLrRWm+Kd6K/JcZ
7MibXBGI7e5tUSBqU4jcd7l45RB88Jr0jOiCvxr+vdiQA3aiBP5gtAQzDRSdRsLUkmkpiWlI3Yll
FFgd9S+zWJix4SQ4WcStvXqsYalili5/kKOf7QjpaQpbnMPS4DUJ7bciS7QByU8xXWKpnVD2WkZC
eivjDGoPdfZF26xycCnDSV3sxa4/r9J/OF5CtxhYUy2b8gIs2u7W9VWeCedrQFWU/rXLHhhINrzz
DjA5lrR5/wk4J6r2NeBLsVITgftzYY6bo9iBUMm9Wg4iFvi66U5EUUpK2qFWwhpIYRdNcnFJNZ/2
g3ypfun67MXvdTA17Pf+cy98X9Eqzrgx3Y9DbXwT5AyDYy3bT4PrtEbJcCcInZkiwMdd8KUf68OI
xR8Fl1TbBB9lHSyXg3fTD2b2IVZskkIeJ4snitEJRP7LLrO9MF3027QFN+YfQkCack+WqAT9x5bh
q64KkUCTw+fsVDBcmtr5IJV6auht9UzfV3sY/CN7ao//oQ27P47OTz1a5uX94449MWkr/OzozkbB
NKeY/HuQTJbs53GfSeBZxd2etNQiyXC1tqmqz4HOFuWEP4U92UY4etqgigSw1RhxNROaNd2+u7fA
YH+Byxaw0d3WXBTqEHbmYOOgbyQKc3QhZ/NfF/31fjDdM22GP7vZeHg3RFNYvJsA7j6NfhitEB/P
NpkHgmPLNqmJ5QEw3xPrgECoJ5jxPajOBKZFhYxlgTd6zge+aiiDsxm0ZuVtZB5SJG5dIdHTj5MU
JaYyjn9sZ+XWGNhUJLgpSivdlcpL5GLiEHWeiWM+eDEiHAZ+76eElVXrAmujAD6NT7iAU53+dVjO
3xVErmGtIdeAMsKDxK8v5acDYBL5kfjMoY16chAxyV17RnXNyFSjk4kHhi6FgrkYtZ2BrsCPpI8W
6tJC5HgzfO+HJtmrpg86ZkVxKgb1QRy8R3IX9a3vjEHLul9uaQ/I5idF3eGfWO2aNrfo5gUzcAHQ
kI2qol6STPeYEAxmGTHNno7q2VsP/qUKeBNIoWJ4kQpkSR+W0H6TnGOsIJwIwQDK/z6EamIB0tem
lxb3jmYXECoxPJtlwLtR1ZxuvO0Ve9lZnto9GVXEqVGmTlf8kppG6cRpWnWuaFmdAkfZFyDuAZnG
55DwGY/mjE48wSG0oyftkfF63iybsuinFB9WnfK6XvKLclgS9Dy1ZtfHMWTDwGdZtSG0whspfNPz
aK0NDqN4Ig6UuT0Jk/H9N6X32vcrTqFJ3l4clwZwOBUwPKMoX14AAvG16miVJmHr3QRBJNyWbh5n
f8SniPevtUY8U3J7RAib34fCv8gz+7XiJtkr1vCSrjeuW5z/TCGeUVvP6SMUmKYcM3bW39zGklAQ
Uv4SIPjHTeQTYtHM6UVnIVHsABcyPn92+nQ+dKT3UmZo5hPp9eH0oEX3DTv9HqWpbb951myX2NKN
naMTpE8EK5svJdp8wTb9+jpeYk2lmUKHue/HL9J/bW2J4QmoEDpvhrY2/vsCk94EFw+Je6MgjNJ6
0AA/cATKqw7KLGwzOV88H6yYVqJ57V9ygsmgUAkc0SZ1B6A/5NZhNsvPLeWW1EStMlGvRoRFZpNs
RK1unUdkzwWxPQaXqQsC2Xj+g3aQLuCNlwOj3VUCRwFnO2hteWS0b7Tm5Hj/SHnee1hyYay/0lHJ
hJkttDdQt5XdPhfMlybjoM0OGtmvGkmFPQNNuvrXeCKALOLoP0eULQmYAvkmo75Z0j//GhgkRM5T
+A3KGNzQbX+xQtkeziZPCQfp8cIV/7jURMIgN0aAXhd27GZoMV6/pTBEtlgYVh6fN78WZMkVABgs
3K1O7IF+OmRFQLDtpHB7wgouBZpklyFQGF4te4yeWgDw+WxJbPgDPatNsSCJKM7E65923vAKbvaQ
YkCu8WMtdqgu6B4N6Rs3TycY3vD2U/hF5o5icGNF3/RErU11mpxMJcj97Etx/GjvbcSrnIsTjpKP
Wbowpko9F4vX+QpAsh3rNw3OMe0X8z8wtzkzfBqZxILSVC5iT39bdE0/IOTs0f/yMKKD13tVC5t/
Can3EAQ8FzCDfn0tZ3iT1xFzrB97JSIvtHBwq7lyuxGja5DQIKgmtAN+8RGD6zXSm6w7FAns4VxI
cs8vsSOYfJIqwUMo68wtHtK6wL/gfyjPyt+YR/BDfaxeOwnRjR7EzA3RbVDo7dIhj5mEqaoCZjzB
Lru/ISr1AgWsdhj6OoJdlINp+cRyj3pqVyZJV6hRZ5KirYZgS3LoFKjJ653NlCMDYGFvhA0rHABv
E+ckIZhrYuvV3mMuAlJjLobxbGLtXRxmix+LcPeM5XTtt/ozIqusaRPhxOhyeNdYRpXkS1RJoeSn
H1nHfZybXCANtZy0SGaiioJ0132r6c2ME1XJbFpJ1v0GQvRPSHQzvTfg2PvnbXKpocBQhL1DLXGW
hOsPj/IlPAhNb94FE/hbXJ404eNwFHNT7AmiQx7+u6FFU3hzhIxsL/q/R8nvz3KYaJVyq13t1za7
ysLihy6TPHMDDA+l2exzCWl7IvY8tFFTEDqfqIKormCG1Aw0TWrf6QIofJc6ymEkvOKatXxycZ1X
NVH9jc1POv1rVQPgIm/MZsz1Pkh+zMfuZaQh/8aR8xfRAGFJlh2H/nX9Vfd6SPILeshlsFUISOJX
r18YT8dnX6JjIByJ/x8CEywmQzYdx9cvReAb2fKzj20AiKJihYiAl+efX6MxI9V/qq5z1CkDsqhq
zk9ANOyeJp22XoULSDBXAvI3Sr58VCm/PdXtvx6zYtT+vf2+shjRbWILMUFTHrZOFxeTDEJT6L1H
7sF13VhA4Z2x+FPKUa2yt07bG5ec4cUF4gPOcbOVNUFaSFWGI0HZRR4lZvGRqOx3lqWR8o2V4Tom
BLP5iKBNPLTU9TOeIvqnIMT/xGKva/MkU56TDykE/ePNtwVfff4srG5ZC2XKQyozIUr3Rqk4IcY4
l5qd87NTyeHQYD80BsGx4VLm4uBX8aF+4s7Ny0d9YlEA2eRaZVCkcdL9cnvOSMtEqtwkrz2LDUoO
TWrVW+FU5Wuf03NxMPbLyexuDoBO50xC0Z5IlFRUBdlnTAj9Wmazz/Zkb0PHyibmgeKONixqiPMP
GUia35FAGsPe1uI4IrYQKKlEI9zLB9CC18ZBGCMCA8uv3c5jwhjlTmDDoIFOzsFqYaj2DBXQ/Gkc
cUKX7gGjL/NMFU4nPKKKoLVrA+ZlMYcJn7tkIZuVeTFHoDOEzsQS5jzqCtH6DTlcRaQ9qjZJT7xG
FRaO+lsh1EJAnzDtiJDqvR0AsmzRrYufISRfe+RCgG8GA5yO4KixJcBo5Ka4ewu8oyiPdOx08RPW
Mx0HElG5DdqRoMmrV5HjeQxRPRwVS4ZahVzFdoI54M668z+adwldZT7Xma2ppEHEoi2zmW+zyK2M
U+Z4fMQrVX6HpoCWvMTo9JtsUHRg9LQHytXpRqTKuhyltodmFM1T2Xh9bMWNB8Tv3+kXq2bjFehp
2CfBchqH1D8xQc5LLRuGjyjND0t4DXAurPWQestiMUwJVsqgOBvyEVjSEuejeUI+qIEM2hOldNKD
DXkfvbjtZ/o7I3vz9ZSVz8yT1KZSVeAbdR7IXzf6TzpZjYWvbTwkvqRyHhbMIZ1jFCRRzYK7cBb+
2blWj3z1VDDN0o/iaIZq8YuZzzIoz5Hz0oj0lv0thspnrSddML8ayVyE3qT6CloLNMJDevkCnxCD
+Xs4g1GMD1wGXy/f/l4Or0QkY+p4k+23hEw8nMeMTvcOw4q0rxM1DiEr9XyM+MVh9rgfKRd7mKfM
xbiN82ZvSzPTaBC+eR+bmYNDtMbyBiGMrCyYKy1sT6F50LqVEC5wYsyjPxZL7OwYx5CYsBA8lDnm
3M5TOQSQjGWwfJU+HJ+/aN4SGUG042cZMtE2gs2dcH13Y70pVow1u4QqBG6TOpppn9/Zl9Y+/af0
dYJgoGyCxsE4czBdMgJVljU7wLEWcC4oKeUnrLzOo4mTVc/RRzEGhvA0XNCfMt3t8A9otlEAilvJ
kOyO6IrHdGbsSzGVyvwH9xbfhOFVYWwqIyO1CGTNSQf8zgx8jIbITS8eZYm4xMLDhmb8sdUdqhAR
TitnsDYPBq5kMz+I6hyuVv+iQRpk7eppXVJAqhv6bA2n/Q2GDqM93td/sy5Q9mEqonoSy/9zSqja
gvmZZHbygq7IUG36wILK6AkiLTzRCUSxOkn1ilB+kavSSCqR71jtJWnEADLRlI2vXTQxjb1CGFmI
Rh8R27ik1xk9pQEw8on3d35ZogloeE6elbuOb2ldlwUApD4D2aPTKZh/LqZrTfNB7qAjJAgw/zFv
9ValKp1yr2RJKqA1Jeij3BKFMyM770kDP5Prmt4wa8rqVW7OvL8iirg6hkrcBRjCwToCL93ztdJk
U/G4g0Ty/oGEwbMQwJdY5kyxNz76zthrlnT0Y8lvHjuI+oA6eCZogFGEQnimcPXiQ+9ShMA1IoUQ
BajJoDD0GZlnaNXbl1j9xqlCunno1CscaVKQ/s1YKmKQX45Mrp9KyxfVfVTaerDw6LFdpB1lT/Zq
jLFbZGV33TdYI+Jih82qnFUxbisk7nLb6sCqu58tvxLN3/gGxa75A60ZIrgbvdq9TAvEcpcKdg06
GekbsNbeh7GGr7swNm0P3Bq5GXR0Nh/RgytfygpRbwlLnz6xglU1oPj2HL6scwqkN2xFOXdBwW1Q
I0CS7AmhNa6ID34n85AFq63pIr2Qi0Vvw6vtlJ2/28aXtRthg741k1wwucd9nb1rOlsOW0eUg/Oz
wgg77RjZs/aQMpUhNboZZSW9zP5GXDtpxQjQvka+BIIvwCVv/Y7NbNYZQgz9u7C3hISEt0qLQ1e9
Zqs0uR4uAT30VbdtdOJau7/827NSnrhWoPZLvtSOb/OyRMcUNDEo0ObEGUSLoMcjNFJqUVNFR8e2
Up//acdMD0hTfAFxN26Grguyfg6fSyeN7HFI6Gup+rFDS75Z48HMCT/gLy4+a0zjqhBexBJva6Ep
dWqjk7XLa/ibGZl1U2cEiSC1tir94UXI2q7f0h9vbQEPCKqgJtKKIQxSmQ1jmwFhQ5jhKbUaN7K2
VDtLc2con6NpyHy9Q4wn1PRztKrjo9NZIJ8HlQk8CfVanlJHGlBZ+BGTRaVCYMqWAfNFMiQxthje
/D7gmDaRBUviR3erysc0rhR7mkO0cj9XMZw4jbiyfMqUpsQmIhp1G0fw+Du4yqnTp1kdnWDfY+mB
owvJjQgEOrIxUOlNgxupPVkyTCis/baglNWYmuwkupn862wREv0226jPdSP7S0nEbvtMJn+rJJWf
u11n/EZJ50OQbCQY7Bnt9s2s6j1mlAKKyB15n9kZeH2TZTlFmpWiTnyqotLvJ2dobIC02m6adCFb
7mQiujJL/w6h+ICTeHXgG8CG1tuoyc6AY0tLrN9nfEz6muDRBCRseJn6ZQGs32LNRe+a5qW0Ufts
Z7tMpT4z10XNxMMCnby0omYW21H+rGV095Aj3JUUmCVvdhfpxdlFjyZlBpYicLxSaWLQFLeuaAN2
fyAG1r8iB4aAnfv56gmy8l+bKf6M1gpy7iAHQKAR5w1OfMunDmI49ALABn4mfigw7cwx6AZ3aapD
PzGgMti6PzASD2iiBnijWtkOLzhwpjRrWO1E6bt9j5BCKVD18bkiysfnTctyt9jafueruujcgJif
ebT3Ix/AhWljMQ7yLvK/6z9073LcH86vMPrtWJd32jFC8pLaiQ8u9UXdt67Xqr1MJXdIR+NvbHKj
NUoVYpfEhU45+ZjVJa0JohgzDiB+zdbnO5Whdv7pEio4v4qfZZLcJL6DL0DSg8mOVeqkuhMFn/L9
oli64yZvKF1Y7LkueTDy11/63Aj5LRLs74HXrDv5Pf7B7fpyb1kIRgEyYY+u0C/ghYX15Cu7ZOsr
rb44cCoZYhFI4VoeiikkUrQKJnLjEQ2hPFPAYjW4fdTibfzXPDKLtG7UarmoOee1H3wwHrxZp3cZ
4q+RhB34v3tedq8puwJXGuN4XH9TD3l78gwDGJ3NM2CJuRKaFnc+4+FxJXzOhQYobK3A1HJOZvD/
TFPKWvsgBja+nfnDi28ao0xshJrw/wcMOj1gjw/Rn2fuVF96+RfKfmL5JppS3OTTo3CWS9XLzoCJ
X6tduZz9bUDABnn2ZHzHqvOW9BXg2J+RI757TQlqNAMtDykaGYeE4QvaAFQxLaHYC0m7KJeKkOvE
cBRKhxY/Tnp4orQyZqahUQDQIoBFnxowaVAMFGGHI3jmnBoOgJFqGV5nNqUwGuZzulB4TvD9v/09
1FfVGbCkulo81WNpfF6GHpMlMbeoy7eaUaKu7xWq8DQKAHc9B8JHf1EwzXmNJhgRywTZcHw1ZpAn
YeiBzf6Rw/4BTphopxXxRtOF03KRcHphyk6QKCwFR2YirtUF9zg8cOaxXiTs4muZr22N2tkvnLlO
FVYiWHG3K2VwfrBK9zRU+/3DGbmAXeXJcAOOJox6jKoKATxDB545Uqvzg0bLnvGIFVG/5J1tM0rL
kqDzUCNjBPavmEAmK+J58xbPvaw8I0XBjDXC3Tl1CM/49/CPr2CRcZ8nS9q5ma0iF4bxqZ9Y5j+w
vElk/Q9u1MpofvyZKWk/DRh8ffGDK6ifeNWwCZtcX4WEM0y8Q2yQLHcq42LwRTU70ASl+zV+1Ryv
QtgYUgo1vtf0VneQGYA/b1zFfVftHkK6xDjoLmx2NISg6YSjI1oeva/8OBtST6s92FiJEN7GuMho
HfMd3g3xnLVhCLaKur9Jisv+cUeCnRgGYM8TpxiPMqG381ISjm9Nfw8hOS7iiXEt6KUKULX4ihsR
Cr27tMqB1Oh/Cx3LKX1Kd3TBHIqoF90aBeHJA7cNI5Tro7Z1rikgcxSWZXuR8mVBvFFJQWhveCpE
BAXCxtEmQmbrSJLib/EM41H4CzEBj98v4HjIr8YFwe3QbmK66de+XMLrr341+WfBEknVTfxh60+C
goP5jzCRlhq4r53vqcmoo7qTODIpxtx7ur/4PL/lhsNHNtDM0Rnl0JXJyqRfuEJJH2WhimRs3frj
JVdUAMzH0780Xob2UmViKDF1Rx1qdFlZZidsu7MeBv3vddytcifoMXj9h/vxKeQy+mxSg/1b8/Xh
fYVmPgWjvzrMlXNyVCo4X1XAMfjkV2yeRMO+Ypq4SEcJnYX+PGtTrmkEZHER/eN4/rXGiEYn5kHA
TLmCGBWM3Av41Wh73gdMPRs62WTYqYHrTVH9gHbX2NFUfnFdfNSe+e9hVd6ofYZzVgMlf5PNrXcs
ZFZaQq2J8bJdI/vkIl8IzcCiUSmmildHJ/X75bldi750F8Fy5Qv9IrqKMU52Oag2BbRtH2bCIk6T
mDF2lh5NWVfqugIEWZPSusvXdWYxPreIH51NfR8GoFaNk9LAxEGKJmGuttCifDoOqAh6cNuz5/OE
cQ9+aSnQRfozVAOimiOcrTJNu7g5ddaqmWQctWXRGfdnccJ0vLGclmAm7DYa7Y+AFW8X89hAo9WA
2J4JQNRhJCSMd4K3O7/JUTivp054Y+uqEU0JkAOWw8Z2jJwKpir4KuqglgtKkxwjEOjz5D/vQsaC
uWd4kgjD0x6SpZbDSEHM0fvSg1r7TUTDtRy66VMG3MQYFIGQXbz2OIHy7nQnZyOd0zUMyZg8DOX5
zS1TKVSRF0EerRRKjyEzudZUXvs2xs2Eia0DDI9ul1TNwBLttKD7PfhFmP3eM77ggLQFYHL7YR7H
FKmlLyKJ4Vg/AS7j0eZCcmGqLtuXxsnxiIbsXyx6rwHlnm51EgFWjwBh0gxZ3Si/bTbKCfAN2Y12
xwUBxVm9xQ2oYcWoLDVPUqzJol2Tk1w586oTkQxIOBn5HzuiNtjSedrpl0CZJn0w9CovSWe+RENl
IG7ovgSmjKDQNCG+yG0d2DTw+gBgWrl2hCVqJkZmw8KyHwS+yHMn0GqXZh14qRz1g+zcUuRcq2Rj
BvzVFEtgzJrptSz+5ziRF4a9WWT98XieT28Tq9ke+zuIKhUnJ1VuUaoqvvcCJtx058h9EcfzZ/VE
QZ+v5KIsaWVc1myEoZWNKB+3bDUbtai51OEQClZOdjULvIc/Brz3PqqFnaUqH592yZg5Tcdsd8fP
s+gdy5bZsUOpFllNS3dYumWdd71W9whZ9yJy4E74IDIFlLAZ8TUFs56KXdqfgZFIfcnk024n0oEc
/xG4qht0FGCgHXV5476+3ySePTXppfMs1OXHLBl934wrmnodN+qcoRPJXZYvcw+Mam4wQU1OxQxt
Qgk6+FI58tA1rbawx+Z1ESkZFxqaH0ayFA5S5mOfszhUgz4sazBjOKjRmnF+klPFnM0vX00h6Ds1
h4XoBaWLe0y0H8Z37W8AvmDO1XxkP81BxJ5AamNdcpz5c12su/Pep+SN03GVUVAccQESGai90lkM
nQNef9PWFWhNnJzv4L2t8+8HuIp2jg+Ie58yXKuzbFqtNbs6LjyPiDPz1R+ayucvmOaORDkIoqnL
78zHRGwYbZvztNLUSCVY+O7XfcRq6gkF+BsszKBlqaBD/MxdMHIGqahYcDS1IqLwwHmx2dkavjn3
D+u89nsD9f6cf8vmwpb8xCaGuzkPIhItNnyYnatTPPjUmFvritjVk4526tcFmb90Jq3GLOwpfXDb
BruG07X2QsFXyNbjXLQj+A47wfizf8+jfV57cAQZ/FTobE4ee5DX684832M9b1GDD0/uCvaovBnt
g4Nbsc2rDlXCUoA85o+5w1I64eL9Uz8X7pVKjp3jAtgemvUu0rRGZKwORc8dDi6FkpuZDPkbx2OO
2UNcZp2ddq4d0PxK8CfvZZNuHstilvP9PBWgor0RlUhr8IGsX3gRKFrKIfVW1y1SPTnAYb1i3D/C
UWSEumxQBxhN0q3W5W2zytOpDydUmHpVw+lUdHgErNaNcq148DPr3eAvJ/lc8N/zQ8qkBizxlHd4
whvp7aUn+TO9mFGT1K6ZkWYx7FEA1fCn749R7cu3uKvrpzs7SBeBSGXOYv6bHQmX7c+E4s78x8tD
/fZRPZ9yOurFM0EC7j0Z3JKAXso5bDp0VV2Smh5SDAjzMCVGCYDCrpXL42dCC152F3mf2aRruCkg
q2qeHJngwYJg96H3sKcQiTrrJMBdIRqO2+h2yk+we23j6Z9KObk3Cfh7WJuoM52L4DyadrVbxQdk
BhTGSIaFsDPQl/Z7Nf2FbGlmiC5b6VeNqSDNM8Xm9zK2kXzCnD8PmzvR3nDGQmSX5gpk0vPFJoda
8c9Z52K+b0EPy2EzYc0TIKHcyJXkMfT0oduZz6t8A9zCByjYx07J19T+sb0sQPxGohKK9lDJnLj0
nd4oMabvQIJkQe5lAIzR65JrR+HSPLyYvaibNZPxt/zHAj6lF93D2L/TkMHia3laRpXjSKyJeeVp
NStA3LLt17Jba6JybUp9jlgnR0Ze8FsKOwVTF4qKiQobHWmMRU+ab0F+dX/p6y8g6E32fpl4SHKf
hyIbdAGFf9i+xwK0KeoM+1IWOlusna2InSqy92/Iw1fPT3wsKuteTnsOBtfMZT48FPNOYbonvd9W
fbrTS6NJoH9tbFb0LD9Hszo2z7j3z9iRn+jDKXmSISbq4VFggKbZESSMV3fR6idnIGjvjQI24e7k
yMZ7dMa4pN3LUsQIXbi3METNqqLYxMJDHMOAOv3RNjhWFrcyuguxJPBHYolZgZ/5mJ7/o7pxkaDS
usItIn45FLANhEVrmdbZNjBKjf5+niWi4EQbLDQtDrzfgbCyqZUzAJNnlPVxgusKapdlXzL+GPOK
Mi1XdYEDAw1gIloC2HU13KR+B59x91rXm7p/dEcPZsk6KJx4wljz2q6Gb3xOrH3kFYwDaH4XX+DI
E1cIcMgAGcg+s76ABZHTMWK75hYnNyyYLRwiUBrAQPIzXOECIRmOO5oU3CWB/mX+JivuTmLnK16s
BWmflS6jhP3c3M+puZwYVnf5x9vX96nPRyAfbYyZ+SBZWBhTWBXs4hWcSMoyfBOjOgT0In7Z3PW0
pDOy7GrxOhLhJniIJV+YC4hmJpAtWsZF8G2K6HfJm0xFtAwL3RNSrhNWCvx7+x0OK1Urcqto7IrJ
7x0HhgedgMyUYXVryKoxmVfrUiSCinNPX+OvRXLtwCRKzl+jCGQr3dd+4WF5+vGGXWU3sC48wZAz
Rn7wdCY5rUob8/qN2e04OBRNBhgZGLMELTinBLnpXnjm6XvOjSbMTIYT6mZC+KViNbcXRty8Sors
hRGcp2jeP+OzJmD/XZJD6BeFaDKYHlCLUm0cj3sPyr1Avn0JqI3clV4HjizYTTh8qEMtqPDdzF2F
PjBbS98/nri+oCuUUaar9oTGWuT+OgF6N2/N1/+3RyGCrlbvpi33KWay+P6fIBObZrHT5AqkuGT4
oIGcHcvhzlqJHdocLCCMiT9NY8OG/PGhboi4clvw8szXweqtpdvIfNTSA5RqjI322Qup3IezGyQg
KphlHcIOsUdGIYt9N2eGQS4Hdvp9tKA7gCj4Ui2c13NAKVoGplvjDbzO52dyMlwemvUINI4mBWET
GhoPjst/ussEukbjk0D4uJvnquPtYC70i+Xv0pP4SQVqs/nl/JjjcTtj4/SkXzHZCA4OIhsw5YFi
vGBgLwguSSvOfmCSkOR+nF50qwq2XKqVpifAw05fGKhl3JU1VoZ+IPjm0YD5bxIGqav4LCYDX3Av
QoXUGqrIY+YdYFL7knuVSAHOGKu6dEWe0PN1wdHfq22koRjX/4959biyOMbCLTILzQuX1O/PbKQq
TWPg/RqUyHQI2N8WOVdjYxC3Kengk6RSGNk8JYc9Ds39GEzmUDTidhSXAVqxsVa7BwojVwf5Ai3F
VpcXrTFX6ecFm+d6rA7ODwtPkqzHWsMAvqpf7JXV1BKzterDC68X7Uev+ux1xpVNOq+aGDxcoN5l
KgeT9FcVztIf4jOxgvdDpyCDyAcQce2TCIsnzEY4dJjsLr+6KMU6z+gji9/b6UDMHleigXkd0gJ2
zy08qLvntCQtcxd9dekRBVPZq1kJqlm2qLj8HicOnbnbfb3NyZip1WZA+KHk0JBiMO86zTDRKOMX
apOOhRGLBqVc3YmDLIY4Cy0tmqhOz+iXyMR6s8Da/ucAwUw7if/yU7TR6G/TWNTbYYvQ2yEXUpoM
deZoeILKOMlBygFhPSqSc3P1AEsZVgId9izQT6QH9YrvQjzwRhDMrx3v7bj+kWQPED9JDhsPDFAy
w3FZ9XtqCGSmjF5/SfaZo0gU32QXWIW1upWdEDgFwac8uTzHl0EliwY0rLMYEs8PpTba5+AAZxGY
Go961pXb63PPxvSFOlXiAUvEeBhsb36592Nul78H+QmXyitfsx8fCWw6//mAYHUEWKlhAGZv3xU1
GqXTwKSjTUaTAJJy4HQ3WBguY6v+FeIbJaCrVDywA8soHaXgAlYm+TyuWJchx932LmuLIyZxNnHD
RWz9lBlnH3mYbUnVaGi1u3E9iIUC61bdWlpfCoUddMWpaJrdeOemRt1+H5QSJKo/uxK3nkD2ISuA
4ru3Vq48kITe8c/SZNTXWSoCzN+EUYwNIbDrIn6IKWKa+S0dS3NTBN8Nxo4ekUAaP6xQktgO4HNC
3v35rdbCJJ5DAQeLdVEIDmTVEJMGmDhYlNJEfvhYLeKP8jyTrF7bBNviEiXwGapSoQJ9IZk9Aq+O
+zl9yuaIWHv2ErsDSHunQos8aufJcd/kqivGMfGywC9Cx3v9A86Bmr+Txa3I+3AgB6O8bn3xsuOY
/pCM3Dn5vSn6nkmUoU4CFXe/dS+O/g0mXGC7TAPVUhXpH2tfBX9F6f/4iv8zPwaB+XhXR2eh30hs
pm3BCJ30AP1PP2+ygForCGe3H1jNRSvshzfEpqLyAHbag3BR7RAKkGmb/DDA7qQf9Dy6J9CNCZJT
I4cCwr9w0vKc8IAH+s3hy+F2eN6V2UO04aF2q1Rv6LSKfCOEAgNOJk+mP5j58rIcUaHJChX7Gs7j
yqeaQ2rIqiW/6MlGJiEIFGUyv/yUO69SJ7JyBWiPhNrnTU1YR4FOvs9mKFfrjlmZrnqBQp9ONvWI
HKQxndk1ErxmeihQjrTxmbpTrSspuQ7XVRwQ1zl1F2zD3W1g0xSoHtOb/7Ahoju2b6HFopsBfLkm
rY7VsEimbz//cfVk+j+GGoU/6gFi8gB/rI6yLcRJegWXGhnL683ad0osH1Ncr9uZX2QTfIdP1Pd7
evZs1SzqDT7TKFSyInfD1tv8Nr3OkGBOeILh8xJpUfn+NsSTzIR5vVYAuiGICqgTkbwn0FAxX2dY
+M4Se6KlkksL7aAwK+5czbI3/ypJi+2f2ee48YXjjObvUI0gT7220iZgAIQZQpvUy/YG/5Dm55sE
5OzlXtyfmYN7mEiFYMwBA6u62hWZ/3uQy+UEkhYnp8LU1gGccBsLl7e6z1gfQj4pKRXJRotgx99N
OnUre6DZWU/wDi1HUaE8yW4SJyZjeGd2LPb60gMyrCc0Amth4E5QChxHudDKNMfg5UvMDaq5ZOxe
Kwf9icsAHaU4dCcQB9eAPi4XZzJ+h2ais26/n8Yj+EVbbXbz0Z5f3ay+qdp5zP57KBAOGJqTs6Ua
WVDhM5xOQNT2eychFtn+QFPFOF+MHkFysrlmInQNKb5jfIPKh98MYkJ+XH7VusYNKMRI5XjmHJRl
mBk62bNRpc1+1XGJGa7u7+YTaOeGkINeb4AC6Nqj27zQrcYkJnwYd/TveuQ4yPC91p6agFjKtASj
UFJ58dh8ecrtLRpyk55+WgW8KW6qpZf17s/XDffO7PDlpp96p3+wz54RucNq0008xXSw354SUR5E
gSyqtAFYmu3+9ipnWW0nwwH5THqtEW3V4PgiMsZ0JUDlviIE4Gxtg2XEpDyZpFGiKPLSWpxBrgSe
Lw/Hh1YZWjJTwweNrby1KckkGUmIsC3UGGRYvtvqErXRrD+x+eYr0czoKq9czIJb4wyRYlbj4n0K
ueFauWoGIn1sgR4tKUhxxUIES2vYkZj4DG5rKenO53fu5Wt5q47avPkr1atDwrj1EkYov7U1QsY5
ISvf131XKlzyVCu7QwJThkMgh88wDxI6o9YAc82RYG4XEPKiT4GlwxdcfnO+5w0C5q4sBhtfhJi2
7r8dtV1jFXkh6JzKFiYki4Wxq3D8wMiFKQDOIil8wh9FQsPdCp/YvHNNZ29IJu5VPBnJ5seO8ETA
VTVoAMLfqvTf3//zG8PZDvGDfhBPJjNAn9N3aRLFmKG97m4+NvAb9VuyPZZa3q4P2Y4DltHVaqLm
TuDjDfbTD2TTbwbXJx5sdQAj1KryzCsd/QYpfP2bNDk+J8AwwZWyA21EEqffOmNTFR1iRTseAMxG
Tkh/MM3FJQnxH2NbRUPL4HBvnYy/uHvGKtuR7jmK4wqFIWoGCgelgNvfK8FGB4wlm/uBoYMpd09x
wCcfZchUmSSVrR35WKb51oD8ZScTUwm5eLL7uX/CW8wU8yLr3e59BHVI7DDgOguWpNdL26tja0SR
C6esEUoNb+fWudUKKi7dsZseTqR16ns47VUOupb7xyLtswrejv32JkjKL2Zx3bjR5ig1kp7iJkX0
ot0fNC/OBHxqpOCtZ6lsovoiUHp2pTpY02g29Upixzx+Wnq8Yi3n6NQnmsy+kogNQIR+/ZPekbWG
o5Zmd2+3wRF+zdyZ89H3jyjkgPISdX+0Bt5GCn1VbXMhwlt3TR4qeUy5pTGIdXctJ3XcHdK7KEFz
MSAi96YvG8xi92UDbAp2gbfAPBCICRHFEqur/tyWkKJHXwEGVW9+KYe4Muy2UEp0taIWZx0c8gk/
FELqB8EF2k273MDZO4nrNOaLHkFA1z6FVNmXBEKgDkub1KPlQTPIchle7ZhwITon0FJgyBDQ0ER7
rehuVVFbKfmmUj8ynFFkO9VMcadt/4L8/zumMOocVgNrqLWBrkp9++iVavc23NxKYvEPKDBX4GiK
gXanUDZEbVKbS+byAnvt/qvFeJdwkPl1lGIIQrsEAXWwClsw/Eoc8VTxtfgOVzUIunPXWRieFTSz
dr1E09K9uZtganFjj4SfdJdA+TaWT30873GY7ViPZ5JEfyMR6Wx85HSZUXfFUg8gqPeH5jdyjlyF
Ga+oLrY/uwFHvFQMJLB+w5t7ewEC2JHT3IMWsLG5lpR6NpsSvtCPiEU5c2ryhJ+7bitF26zsEBjJ
mV1gRcwie1veLr+yMk/tj4G1zRUgWKB2GCYZsE9fmh/L9xMySe9FaDRpHTgv5VooKywgsDzv5jGM
zkZTQili4QeTKz66pIdCCdhiy3eK8owOuc9oT8EC5el1ByiR1QGNN7DWKuIIJ3czGcDbvMNUrSDv
40ug4qZT9bN+bytvLhEf8Igk5OCWDSZDlNySEE99RiaWfcORGWwHkzOb2JaXT/W06jQMR55dP2hL
gV3MSXIXeWNCNRun9tXjjjdpwLICaQFlE6LYHPzXBZH5U69EMj2zUWABX85CCBC+L/3SrA6v85Fg
fZpHpFV10sBoX53Dzy4FQa0u79uqFe5pwDkaOcpqbsV9gjGmJnmWyH6bX2ibjPw0BElFfXe6/DKt
yvjyW1x3+cY3cXOJ2xK3MEcv1XLIbEPZp4sNDmDmS5jCSxNH30cAbDwyx4/v85hc++7GfWG58P+i
VQM5V76n5SZcEJz5V+/XakovuhwEaCdLodjrxP7ewtERcOHamnTZ8vMzZq0djHj4MfUeTKXLFnuS
URzZC8WCfVcRqkrR7uUsb+4zvJap5L4T2Ee7RutdvzxJH8IneelnVh5dRoTb7E3bOHx5vr4586Lq
fgsBhCqoPTPv0otMDy7x0M93tuWy3UC7ugw9mA3AerE+RCRT/NtYaI+D3opGWy4H0z/fBUQYiusQ
O5A/+CGtT3WnTT2b0WY3TTOaYQv4is1puj5DXAVqZZIWjiTXJzzD80OE6i+hl/FauPol7QIF73f6
s9Lcr0czpb0idUhPoI9ZoufV2cqbgyBs/nF2mENGywYUKGyy6uHm/ZgDY45qV2gQIsZrRgJV2NL6
gwk0SkgCHcNCjbGsRjRCWR+HUZxzqniYfbIl0GUu6uL8gvwTRJ8aJrYkp1zfa/FhSDWdwXKyM2vs
n2J10QPpxOwvb8UtqmiYj9s1Y0neBZz5SeEw9SXgiG51PXVqEHDNTydinA5E5vVs5WULcxfZFri1
Oc0G4d97Qej+qis0rZ1FvDWYzfDa6RbHXtvtn3Pbu5kuhgX6NqgkTqWXgMSMQxQdgYXFWS2SyoEf
YmFM1rphHVl55HruHwdOn3VVjJkql1h2pO3/JClyxWOcpx+eqPv5/Obe3iBuzlPnIO9hEWkfADDe
OoJEKDymG6tfOC/tArEf7y9y6EYIqhvaeqrsGsapJ2atARfKu3cujKjqRZxe3yHKficWNHAticoB
elvnykHOBgIDxcoUoR3aQxS9/pxVeG1FrVH4qX0AYCsNuTvPlC4o1lhy0ssc5UUFKLUoCJXChWJl
Xg7Haoas0sRaTqmjzQAsahR1TgB3pkuCcFV7X212lBXtiQr7Z74AhB1k3tXqvjJf33WcZueu6Zil
FKABPwqRaogN5UHzT4dPhrpm4M9p6J9mYqg82Eg+izyQvcRMwk5X2E/EaSbJ+hWRoNUA65ybSzS7
2tcf1jBaYo/D5DE5F7M2CIip8DVzZcH4kJUBnQB18eCZI1cfEaTRdlEc7JTLcu2hkfmUp4N18vKt
q6stQnswMuAnWXxqg5bw/XfFmUnAHKIvz/kotSLz9deswl+NuvzV6sxAAWSJp/v6UdnSavVwP4gT
qW3V2/R8QWVQYNtpAyuFgZyW3WKXDxVcbGBfBdtgaQOtoPfC1gC87CmtHF3L2cEbdyGXBHZop93l
zkS78UERtFXFy7eZ3aW7+LsjgRGwmW+7LEcrvZk80KfO84HaimK7YzvdZJkgBiyqmcAc01UkRWVL
7Q82WBecBKKWA5EV2Tm0Uh2ygcfxO7wFWBG80MMXF+FXOsjuI5PMYjExIrskUBcrtBfC3NMisEY5
X+7R4StL9UC2MYEKgguKYiq0FyMjnxajVA329uY2UEzdGvIWog2WY1sJt2ji8i25LYBYRBPzUAo4
+FKMs9W1MBOmKPLCzFPAwC1GJZ56M7qVfgC/gzdiXzt278hXuEyvmBFwBaM4FovHyOcoVy3EcpfW
L2G36LBhgWQp0OCKhkuTDmBd0JziSq4VVuSDjgEPGCADu2zMCLSmmKThLbyRX8iNhz5/D8HUgVUA
SM85XT3a8AICSjL5wzWbneSprXYzgjSu/ilzWNMXEQw5U7BZTS84tSv/mgnvQrswpPL8RwJfSOoC
OJZCtD5q2Frs4mBwNMUZvoaOdfusafovSS77mrbiFpn9gTcjio+CGkudYheBsQSwbaERzV00B9iu
7ls7DBSYXTNuHZn3A9FWArnO7OtMz1qRiWdKREl0qOgt3FCXuJJ5RVERYiFSuU3iOS4HS/J2wdqD
R6cK12cW2+woHDxZUMGw9Z4tlaFCCEMDmjNIfzKtJYAyEAS0XCL6ns9QSnaZF0xCxazCu0/iAUz4
oqbSyVvB0parWTrnuP1v2hArEqowjV6G96NieMUpYE6rCbpsq7xuFR0uMc+KMCkIl/1I7Z0zf8ea
mzA1ioFSee3J4icLYmdZ3i3hBi5afcF7iX2qa2hKfWduVKtsmntj4/4C1JVcCkHO49+taPLm8y/e
d8Gud9ghDBRCa1yJ8PjqLtu2b7/5Btnq7LXH+cAdBCKyg5HgkzjYYyahycjAm2QSA+QQvctfO1fs
EDuG/ZzqslI6poQ0e2SQ4Ulnzk7FniOwxEG2CZzANFKh+uqMzIlJWzt+MqZ9eI+4sI0IjvWWoehw
a4KIODr432f3y4ypviEkDOIb0+pv3rXA0CUFFGPx0NuljxOYzH3IVCSfhbKz31cV+T8jdcaqF4bC
nzTFsDWsIpX2fJSo/AYTFRJIH7yqDuCL5xGHFm4GWx6g1K/rTIriGAQ42ftrUCdaKMr10j7aNo0f
1q70+3fF3aKdvPbnzMyCW/AorU+j5yN2sl9ZdW2rbPUp3XFm2SRHtDITkfjZiNPHoA29b1kb2BlJ
3tmLCdSUiXbjS4doaNRHgyf2fGsx6AioCWkBYobd4ayLVQiq5p1v6pc9gu0jOFLS3CpdCDc6kv/Z
dRWFkHGrNHWJlWebA/Lrx7zrruW0c9KG/YeTY7p/Riw1noX7Y1pYrOUpO2S7+ZP08NC8+wmFhZcy
ZMhlqh8tE82QDjDAsc/nl8ySrzZjh8VhA5mCDZv1LyHs/Nwy4CN9C+pX5sLtVMT40rLjozZn3YZK
BMYbC0EjYR+qYuRJ3GUL6Z/LBZTyXJhOm16+wNpFjoCBeMjvZpETYEHC3vruL3ECji2xljeRGMlr
OQKK6t5ZAZ8O89Tv+63doPg87s1/gZSlUnr8fONEUMSM9bCbmLiyuRCZ/2yRBg5bhMA88RtUPFm4
S7gDwxyY/zojwgfEUCCRVb3Lo81nIfdrRrOCDlcE7lt9/2GT2fsHl0hJC3CBT6tEIqVwn31gebsX
YFYIwzG5q2UArGu6vGJWfWpIx+aq9XrxVyj4oHU+Kz8Xz3dcnJkzEc9mI/zbmmafw9kUQyAUqnk7
UWLFkjNd5lISZ4tVGWwdGwPlKUW9Vf/J+4lnDYmGM0QyRrmgyeFdHtw7HqaD4i/snXfQb5cV0+2j
rpPJ107wnUZeOeguPOcwMMSRov/n5lZVblbuRP73kZEIEePFPy4dxkYbYHjTU8iWBEcvLNRppJpT
zgNl+lshntpsazLYumzcZRuaFMjyfFPNl5jz6p7jmF4v885IGoe1iC9gORO8YQu3Mz6ozQ4udqlZ
kDz8kusklb6Jn4h9EpHxpnoGrOG/+5VkBiVJ0etpkZKIIT/TslDqQa/ZjsDbZjiFf3OTbXRhRA/+
KkSn5eZfZY/LgcdJTvqcFMQEBFoum9n8ap+1ajD7mTZbeHtpVTCV4OKOLGE3UnqWuuiuujxQZHKL
qibEUMONUdxHDFwo3y5TB71tNJROFg48G31twP8qTwbQIjJReSfkqB5FazYONy23kre6YtYC5Xe4
rhVuTmuQWi6NZ2cts8ZZWo1k6qRi9B4eh6vK4AmZvQpbo/Km8/sYYWnFAlo1yOSIiKDMjNF5Noox
X3YLBWC7bz2GDDBI0KNZz2n8B0fQtvPwcDSkjHeZ84YZt72arItFB+G2yEaRC8Li90TlDrKcA5p0
QBaZyvR7o101JMdXmsnftFx0pVs1T6H8Vb6nkmB7lr+saugRP/HimdF5ZI6zTzJiLeKhuvCC9977
+l+Rd1uf5vzJMrS8HI+gO30sApp5JjHfMkAi4f8OHIshcOVBWPeTnFym/3x04pEcEXTCId9HgHts
3zYoJdlm2L6uK5ouA1GmPZMNum6cLw2A5lMl+CmbYww5cSOMnvNcafJn6armU/VDsoDvZ5J3IsLX
sQRW/3snwsRLyZD2dOoxmREMgOUk3nSkkk5xy/gj0NJ5CV9dyiJ4b+0ATNmDRZzr+WlRfn3087eP
vvq+MW1WIdVOEaBxJbwmSX+aWrSq7E2GUF/47gNA9v7/rNY8wo05JLBPlFt9u1jj75gRJmb5fp1B
YYzHizbqE6vZ6qyMjm5abxfhVUAsuOvG3MuutILLgw0OtcKt506lfl5gdbYl6InpB5Ibd3f5YcGK
N9n1vRvayPjErDzjuEcUc3aMEXAABrGMQsNxBfC/BkHxmOOq1wEAT+I7PTe7hAdlCBzYj7PoGyOL
3gEZYaQZORGKrMDBsLloAzwhmrJeS4S1djkMVn4BXr01vaaSNPvrVGU4ZuhgwSamPD2IUu6RH6F/
FrLQY2oRPwHtWVH2XElYN77wWevfWrY5Jta97nHtOiEmm25eGdILojWxgZEFMZSyXQ0KzYYg0Ee+
gErf9CU9ZXUg+AIeHaKuQeC/PccRN0ZhJgYRJiw6Vy6wa6sE9zOKq4JO/ZcJ6eDo7V+V3scU1wLP
VsRtA4K1vFJ6hAxb8jQg+Ad0+SCCd3kTOwasiiXL+KaHqLCSZw0EIGwSO6ayVTtQTA3VRQ1XlxZ3
LscuOk81QqRdgKfVetXNWUYPDI9PCVjwCkw+VqgxLYQ9ODrh5wd3NXNpJwkrYs2lpk4uTipZK7MM
K9cVZpd+nMLB/c1WvLKFNpzhSUbDHTo6wxks5qkOpGsrQTySb2yp1U6xeTVuMT9gqDdN0u9ToY/s
e/G7dC4rBdTQJzxBsT/sL8eGOCTiAkyMQZZA7EqkpfTc1FeGEj0aFcpkTIn+HRwndyszOVgtIkd/
8hdwwKvYvI1wA56xhP2B9kjlt5oeZZWcXLWzzvtkjkYUT7Jep7IoLAWlLmDr4JbrV3B8cn5qoeX/
6NvmMP3BhraDVfXEj72Z7EmZ4FyFECbnCV4m4VCE9FW8oMfkzZHGE5VnCg9l9MoASU9CHwjYp8vm
eBt2lMm2BBp00/GFmdoQONvmEFQ2ZJ25lYyoLM305rQEWORilwxsjgbiFg6sxWwwhzFNqaq57jol
TKlWV3hAqPApgd+I+x1lIHn25vcjIZZQMV5qw1kqmwdKasraZOyuWvyc75Mv4pDzvdcdubEu3noI
NIrD2qajmj/hjgE4cEpFl4Dib8qBqrcNxmYT3yryPSlrAHdCnD0NFfOzUNAS5whH7BUtTXdioE0p
hU8BMtijWPBGMxWxIef4/Y4VISaVr3a2hjzw+Lz8yMWuSnN2oVMwvOpGOyR4AADvV1Iv5EVWiCic
IYPZ+W63O6J85fp+Zfgi/JuaVyl1FJ5qqrgx2l/lOp9cN4LkArFmrbxJzcRYoozXg0jzCBIOtmum
bR4uDwx6AKp3c0FDTcMoZVl3BawHz+IXkEiW5iedgI54zt/IRzqckvuT0hY7NVQ9unKZRWoTmfIF
D/hocxaZmfo17KdSYCverVae9tOAU0JDhSPKWk15duotdG6pEbnt+WcJb66iYpOwm7pazQ8BLalN
5li5B/6y3zxOynqmDfTJ2an0rcMBsczLcQK5GahRjEM9+YmxRHIOh8wNLFBBPfQ8psfKLaiS0E1j
rHOvoOZUr8M3mhLav/PO/mbGAN37ioFGxKBV0m5B2F3Awk4tAZRZlSmzZFw+HOzTuFBxf8Y4F2aG
kPAH10+pxuvpF7GhZf5kfMVafM/Tc1uRI7eWboAHKsH4WWmA9KKmCRVKE9gbd90f1vcv0ASsEzFq
TIdRdY5wD7we19oQSoB9KgcIXwjB6JdGMCCkoY8FuRV5cAa+nUwIDw25lfkQGkdgmeYM2uJISVKX
Bs6E0Wf8cOX06+rjMme9OnXqVj4BYWcGIhsIIVjvW1dUiAkBpWkuN8dzUvNCQig5FreqwqQWMcqR
vs5P7JjHq7WejNpe8U0HUm8T3m+tWGJy0Rext9IKBiAwkFoWG9jIO1kRNqhPbfHXA3lJvP4i/JLV
ykDnD0pUrzOgDwPFR+/MK9pvI9traF+e+F0t279HL9qhe8ak18C4v7fLjevfG9RliFDJnlg/i8rU
167FEkxh6a/Remne04bqs/lkSJ0dshPvrwqxS4jnghNp2S0RCKBtA+BohEaLLt/olr1j7RRr+xIf
SylZoETlr7oPiFAbzaeUYJ2zxn+/i3MKoWA0PuHPrhgepQF0XHvkugmW7gImQoBLCOcONdYiCEy4
0TOIoEzBU/HpP7iAvU4LIHNjP337mbxg6UF5cHP6iaLehCqlHLpsDGa80piRT5jhFU6ZLQsV9+CB
EWUEF8HkSY5AuHB+4k3PBZF0avN6rwuu6YwlYG2oCWUxbXhSqwi1rzJwG/ML/8Yylf/+5d1oEpyh
PtSiuUJ9OUXu8d0R7bxjhAO8LUjrwgmgSaFbspP3D2AysXR9spwbLnjHBiNJHhWaRtGoPucPFy23
C8gf/Ksxtz/+z4vnk36ATWc3+lodjJIxmz00TsniSsAhjThOaCe8ETvSbmuRzmLM/t417tLobcsd
DAd6dwZ+F+DuopCImRG60YWOYVAhaSAlKDBaIcsBWc19jpmsqjdHF4ucEbz+QvBRVVAAKV0FRsIT
vk08dvjW5a6YoTlED7v5Ihtu0aW4M+0d5z+yRdifcUnAV1rQBBDEFswy4j2LwynwT2+n4z5c0vhe
a062WzvGqQpIAaKVzOAPSjVx3bpyXRo8NGTdskHCqnGNo6WxLPvYLQR/CnCOA6uNrzK3dcFCuUsN
mcMkaawXT4LzUOf3wiFcTdKLP+C7NhNnuCtuVReK20SOTtIwjRZPkr/Nfw/kJVLemW9Ixo1KVtmc
jy2XVFJZ7z4nFIF3oH8uqW6LdzOhGvu/+RgNyoiHc+LCmuu4IRfe78n3B4hcYx49DjfU0w7AtISN
Y7NICaSxf9P9CXy38GpGrJKIGGSZI3tTPUtiBGtAO5UcEIVZpKRUmMpIRVblGreBc4jJQkX6dPJV
xEbZISbamdNwb4PpvI5lZQifGDaHN1hkuNEVp2yuKnbbc7jIWosFFBvXb5VDcnVDU1HmlWZ6Xzi1
B3kj5Hj9dCZytxSzEvSq1yILWf5M8Lg4jQt9KnrG5L80UiFmjAwSsJr/z/riCyRLtdQaqkfznEVm
KU3TCoAfb6CRcYm5EKviayem4F58n9eIA3LeKL0BRSGwJ4AT+empERQSd3VqhTdR50qxjYf3m6ve
nRJ3VMiYFiziAuMf4FCsXGQp/JnFoqf0QJUbmb9E+WdMQDnVSUp3v3t9CQLDs0c13FTC0zdPzxG7
i21mwMftUnvAq+P1nRHwMDNjOEO0nybn0Ebzu2ok6jXlgrslNVU0scVsMNvOEu9iDwYPd5oDU5sr
X3BkAN2E+dnxcDp2GMdtFNhS3lBL12i9QNhrXdKR5pVfZOUBYgmtWylsXxTfrr54bY4LWrod5a/Q
TX+TM+xROuF6RPJaXLIKYSyUFAlefY4JuS9XGwEPaN141OcTctwqmhTll7yUM1JIK0yAW++Ac0u1
fSgTn3IZrXJZY2SVO/RmSGLEZ2QA4nBSBVipPTMKb65tjPNs4o3NCf9N4F8c62/B1HKRinANZKHf
/IRs/khmxkxAMNXpQGA+QLomw+I69fzbaoj3mxG76M/Wi5SUk+dcC6BnwvwFvKj0SDznBZS4yJh6
u6RekRgIQ4LIDSmXDB4iFREHteJT8HQwD1VYiqOeFQd0xsVKo9pDIj4zbBNUUQyd6qkXc0dfmBzq
COyEYUsqHkKO+OmhFbN+iK8oRFawc+OPdL1LqXa0A/jn17Grjv818OPpZ4hHoAYjkhBwotA+JWev
a7DKHBEB8UKzfISbH3JNkEtRLT+Iw5U4KoYxEN8oJAPZFv1LeDZ5j0lguylyoHN3Fs45/QT9bocT
A+1CWWbdCIO8JscksrN+W3+MiJlrWH5Ue9JvNIvrxXaJ3WmxQ0yzG07YqjNLh1zJItXxqXFFcp5Q
RE5mWjT8iBzYePJKbtI9aAJfRioojv6Ne0dA+3iXPEBvHPD0/SGWtAJpwQyiuTxyHJJWkZVRwOlD
Zd1GO1dazLVjIdaYKc+ZOiHT7Q/8RsR9KWp1DcDYAuHiyl78G5EuaVe9+qHyxu67YTtfKx0jEQ4A
EXDtFx10x8FtbADV4E8eAO/+f4/pimnvYgLVxNvfHvP2ZtdcdTUGtIBL9JExWQVqvAEr2hZqaIid
WoN/3Cgr2QJ3iJWv/goNhJ0EjBU9O4nfNG9Yl+VX+Or2a13WyFJ6yOoeK4J/j3T+kuhj2WP98mXl
ROrHRiyI10WbNanSIhcZTQPO4BlJzXySr+2EMslvg79LbQ1OKdLx7sWRzOtLUWzq1x4fZ/r6J1/a
hfmmieYzLMQU7pi0X9SqU7vsl0HaaUCF0i7jh/R2N7a++3if93WMPYgoFy02DhSqU+3DpxOF1sDQ
1GXbp/3/AbDE3wdyBiaoNqb+krLUeUU4S4prof2WLo5+rUS+iVlu8aHwBAl/3bWZGb2YE5bQ9JO/
W2807KF1GlQ3y7R61RY3TBSUBLewg8mIwWZVRg6a2ulpOhHY/liFxV2URvoE0KRsq7eWvN0xr4eW
dOoxmnqBS+sbgk8u3dzW2Xv5iTOXaSecVhRlMZRiNTrzawSUj3oABKuCy2Y3M9jbwjIk8W4+m6KZ
ht1GAAfnF0wDdPSq/sa9pMAmZIF4mIZjASwHqR+jUoXTpi4xE3cT1ORU1cK3P+rhuQKrSLZudRJl
23C9r+nLlxYcN2QEfz9m/ghsIsFoiAlSXSsVPW8eGAca5dGSSWHoLVTPRt9kQI5uo7MeMhSNmODh
f8hqp6RCTVI1TqrGULRLdFOED5yem+AtSFOtMSXyGbLVNQpglEW/Bk8/r+aybamnjZphUTEn7HfG
arAHRfWxfdl7zRu50JEu7zosqKtJk85Rgd6wxFOlS7FoQfU/LicUkaSl6EB97DnpeRsbgsdc9rpy
Vz/EyLwuvIGdS+QtLRgv6c+kBv6vKRuG9tbaoZJ88pudepR+P90WV/R99ChL0vtJZanaKpJvewFh
s62zq1bi1ZETptVfxA23VzecIRK0s3XzGJ7Jt8aQzNsQ4DZ2dif0h4WapFzSbUJ8NkW5vlIqF9z2
k9UyvaiWpCHMnZEx3Ub1SaGR6OEQ4C1mLm1gQkTVyP+xWdIF9OfV+N6PNQko200nDG48nLBsc/Cq
4qxuo3J7GVEpwb3sQ/+EAEnk6dInIInbT/Hj6FH9hsB+u+nZaBr//Zqpyz1ijJieSous8NYyy1tQ
L2Qret13cuSe7SmFbVAlYV+4e12bzh7SE7RxlbrGX0mnFFq5rJ6rX8490yqmWnLV7ejmra+/EkQq
iaUB5HvxQ222tIWSt/WLtFf9e+1KwUUdlj8XohnDbwRe53rARuLE2C8XVc6uTdZ/GlRUF3BY6vmN
K2iRVKBzCauRapBY05komlNPpWWtIyTfXLEAfVWuFxRMx863fK4XRNmBFTsDrF8wWlzsznU15sc7
xKfGJU1jkDEjw8zWUYR5e7+cNW8GDzix1PCGoPVaBNLbkNwsBnWMgQ5SiAnZ7czOVuMdFj1nXHc1
0Ky6gve3+C3yC5yEjOQa8JsydQ4YlwTplzyyyOgke3tMJBYkEe30itGVVYulI8yk4NJ0gqRNAP+3
N7GWGUDaNXZOxTaI/5f9ZfEX2FCKE/t14UUZgYPmRPXJcABKT8dL4JKRf0FmuYGrJOWnnS4BldwG
f17OXYMQgQtrPGthUlnx3qCkfC9XrE1qiinIz/tuG0Wot2yiNSkU8WW9wj8j1PQ1EZmowNR+gzCU
Vl5WFpbqQzcm8ML+TqnBAu1gb4bAI6XbHSTZ0XaSnOOdUx/Hj/nzyYR/fdlMX3J6AZg5wuToY3/J
4umzodBO/+2dypRXOC4ajT0gBapOwVApG/nHrlE5RKY4DelLvGPJPd1D/MihFQ8NA9DZSfJ+zGfU
5g7LbCGF0dJvLObXnXllRMVw81Z2pXpNr+5byjaMvgHScNah1Um+yKmNKyBdKr0IaJD27bqZAOxT
bNTySJVy+LKaF3t0pql720/zV1G5zxzz4nPgwfFEUhlONf7vxE3s1zZpr826Zatb2YVzbfY7mbgU
AhWxszN+TPKK9xKDdIRtqTjLrufzVaOdbOfWaBJKWTQz7uKBhe+30PEwaVVn+QvzqB+NRc7xPurr
Lzw+77YhoJnXhrgVvkhjc6R14OaC4PicRQzXk6wor9lMLvMMFRnkKqsIPOY5AotT9xuCRJoYWqXb
J/UX9Wuf5X46Qc9pXc7Inp1PH6VVZ7kHwL+LTS0IB/+YNs1cIhSECwl9NbgMyF+0anyVxYPFhcIZ
B+PqwZWsuRRK7eGAFMuwCpSIIb8bvdYYG5qGW/BoB5Is0vya+UJy2UIGbfmSPhzgrf80oCY+O2AK
3PZCzbghmkffc5WDnGX4SdgFgoDBIXHOtHDSvA8/3BKvjJnK+DJQI2qEcqvt7Cr292kAE6Fwq7x1
59yq8q335es5PRrYVEcZ/X1a+Xd8bGHnErXRPPp5uQ2GsnDpB8QOKT+nF5uvkhjrX5FkcnFGdV44
p48GcCRb24NWe2vVipjT8FCCDNyHnAfEy8JbzYWf+qHqnT960qAxj36QKrkETZO5Kz92OYDrcBFV
Y1aEG0gTYGBCSIEH9iQk3Of1J1n8UC6R++GysMXmy6pIIk09/a4dZ+hcFGqcX6fWffJRp6zyFL3k
Kut23YkPAZk06gy4BfP2hVnoqBKL002DjsH3XlE+B2YLouIgM8UJiyvgxTUU1U30cQO2SXcg58vC
gPUgXzPqwz6fnaXMWajzWTtzVnZiGXo8qUmhf5UvYQvWUggrp69i83Vd6F1xNkCLd06HsmJj1yqf
OmT7oQh6ljpwH1zYw+bTNOuYu9Y/CM/JcuePcYryzejtGPsWe0W6ZU+YqmW2cMC/yvgIdUMw6Pjr
5zPDHgWqUzQHMZSQWk09J4zxEaGXoj4w1/gVwni1PNkZBLUq829JVnvNczJuU+SoNEqBeI4imB/J
Jbp8iODAxihi8FaK2PWJ5e68KY+PRTRIUcN8hHJqbXQ7bmKJNSKbWNnCHsQ8lm9IYb8hQGHOA0Ik
R5bHtUFpsvTqOFfQ6EmwZ0ZoU5QBNFz2h0HEZw56Voq5z1TZ0YDfmbZ6/xskpH/wmpdIXmNbpqnw
epQfo8elTAIEMEiIFh7VSWojPWdpVj36yVNqzgbruI4/GnrUuDdGaQ0IWGEhN1Z4828PBxU9fT8b
Q684wvTTUGVEFBOEpPDgaa+neWnhY/mPCdcz6Vn4XLnaOSDSIX3PeY+YgnV65GUL86i59INgyfkM
UiD3lhXuaXBRGHH/ccw03r/JlyHZZqHOYqJaGJYkY0/svCzl/ZTm2vvHJ0tzEHbW7Gb9wjI0RICT
4Bh/puOn05TwIxywy5RKKG87Jg3/tq1BofPcD9RGuAymGZDrZB+yw5wyKpmVwtY1XX3BXXGt5fjG
eyHyWX6XRxfdvyFZ2oUYlvAXRuOEkGoTsjBUJ5wBcUSsO6CkLgqn2k/2rNxae/3E+MzVootaEXjW
TNoi7XMDOwgJaRRZqJy5uUXlxshVHdyI47hQNLGt57PQqmpWbxU7veZPoKhGQY5nI6TAdSmvwqAI
Ssd3uq2F3Oe6zcRNsELNVa4127TNr63E/H57WIZ4QE8jpAoTrFwtLjRP7wlW/RGsdW2JgOdHXgkD
jBx9ra8mowr2uXL7cGu1Of+2apgCdBj+O/Qxa2qwMaZXErhkICza2C1PCTQubyGIK4l25MaHmwmo
bU2t6nDyWLd9DhxSOkWrmVGuH+GtcDkOMpGII51sD360G15/J+SkTAEiqZaEGnmociJBoWEQklWf
3DSULLMP5855kw3azFqNzR8CVYzX9kVi/FFTuNTUJgx1Elodw6GfFX5dldhoPm9TbmQLJcJEelUW
VbkQWtuGWAZxrRaTlR39oS+af3Y/XBAlfPH8v3KN5NH53D03KI9YPReGEUEaOXvieW4VGQbjqlAp
rYjOx0BcPOAGeBvV/GRA/crFe60QwP8xVWIeF5KoizLEPeeoI7l83qPZO2sy5u4SRA4X+kd9WGfQ
RqcF9MtB5qmSQhD/LWKwoR3+GgqFBwnOqQ+Td9sijy7UubtifPKjj8IGplgiyVi5XcH4eAl2HfBy
OViW3rE4rG+myKT5brte6404gIJ1vpPtFVSwCacJLRPfuE4MuCDNNYTBeqQa1Me6kMIkhJsg2dWB
PTHSwUY8G1de00KR56U5/rhy2FXLqqw4rWRh1C3igFANXJCrqduKLo5CbpVgY4E0Tx9WFytkMS4q
wbfs47SwMupXN3LycSzgPBAYHzQ9Afbn03w1YP5PtMcytIHOss8ZBVr6RqjJlxcyg1xGiZuE3F5W
tuenK44ghftp6xAVUxEnUYrQaaH/wFtPMm9kk8CGMoidO3P3hKp7QH7LfHfg+ZPZauSxjAXktczT
Hyp9vNpdvVv9SqSnCtM5xpx5Qx/F2jmvIm1AB94sznNWeTv+o8VTQQ1j27PTiuLT+5llOoGt8RR9
j5dwz99tRdQ/GiXSvgdtbyrHPQ5pf+/9KyTxk2vIwkuTtemcxfiifBHnfNg2TDC/E61UlthaFesB
QVhzRv1y9jrpMZpI8rgaAln1IVauwT5SCaSld4+OIsRVG03mXd8SqgQaxPQsiGomGuHS6cMm7WN+
ky1KdvdpzJxsAuefjIQBkFpwgHPwWj3Usy+OuJhgT4CNTu7Kp7EcsdAHbti6JOKiNGEnksOTqetS
15+xcgysav8SOpAJINEwzgwrMu6MdvKxSYwnfvpwXMPFRfyvQrR+daWP02PeJIM6k0Q9Vlhgu5xM
VPgtogHBRXN0pJPV2DNu+xJLSkenZH54symQMgGM6sUEdbtX3B86+wl+UVhSf49lu4xEs0QhM5eQ
0Dc3V/oRsJRJLw1gB2GS3Tkz7K4OI0xobnJJi/Nk3nojE5rc0YddGmWHEIfk9/gJk+mcll3zphac
/GPPg3e5xxnh4C6A3p2qz+ymucE2BaOLfkU2OQYTRQNDBPQU09ktHR7NNrEQH78aHeF0YY+mLHOO
/sC3DbcUAvSQv307/WzGuHSYWrNSbjpJxtje/HaQnVPnnjNQBIFzp1vdX6PfyqyolgZDalmQ9UsD
C0iAPtoefWV1BhAnfkFYz9K0/Rb0sLkBdkMd7oUhoRbqrBEQ5W3lt2YVH8cUJDr5asO5ciQOWGe+
2rqwoFTIdbQLjwGdVzuw0bYAHpAALZPM9gXYXVvJJX0nsLy7PrrW+p4KKPwV4Kl5DbYSCl4hrpQa
dNkx8bKpbDEwn6dN6g/QWy0dhzohfUDZ+qvesBgH7aM+0MO4P5+l5zYtU3lc3u0PG19dDYYj58iL
Mjp2zI3QH0e1GcxXh4WAyOEjOt4OmsbAUr9a4utbWclNflkdqOb7JCq1CBaYX0vPhndwMs+v4aA1
HYArEBskN6y/DWifjfAkoPEh1Rv6vyoUt3u1MkGGRipC7Laprc5vmhZWxvVEDnzguvgUslXNIX2m
JH6yHkr1moX8BVz2zTiBf+0WDNTUfEuIjlFpMTpglUkQD1kf1NjnDnqh9BtouPk0X5mg7gLxz3mz
Y5B/l8lDa8qg8cQB1O6YJjhTKCDWvNTzpKXVP1TPtJSnCDTCk8rYzUH3Ewz/nCFGywPKgxcPT19I
bl3cYUvA8Ad5RHjffKBJh9WiEmxFTQxASrFFf8DrQeMeAb7sTY6pbDpAFQWRNQ8pJKXiAe89jSLw
nuxxCSYcpBXBsZ0n82bShSXY6xAAg05ksrJf7sbUUJnjAz5662QU9xdTC4jlX3ckxQ0baSTbpl+c
XumK8JCqI/dI79vmIVi8Lt8ncH7Wwh9yOYa66DY6SpM4Mm1y6NuIqk/4lnPYizR8G231qVQ3dlOx
9ZQNM+tjxPPJdd3I4FekMuUPr+vVvrH7Sd3gJ5dXU7JB4LMol0sFvx/jDU9maSlFQbM1yW3f5/ge
uekaQ4pqpHH9jl+IKJ1FCgBKpHy2C81tRVV42ySQoompoof8vspQw4f4+vk2uxMycfFiBGK8xDZk
elVvel+b0A+smqAJKJwF/eaSQu2TMgzzutRDTYKGg4VyqcsMgNYTddhrtLtJIJlErIJ10IXK8f2f
FEqbJQTXXtXhqQtjlEnzbs4QWM+RJLXOQiEVJ1jLat/8peQysXv53Mdny1cxbYONwHGmES3tDPgN
zHX+OdYLRCST1/BuNb1MKgx25iC7JreFONRDJLAutlNkYHzwg7i6ToCvB1JMvOWVkzq7GHsXrLZ8
dNXy9d9EQddwm7iEXzRJjQcgUpQlhjMoJKXvVIpy0VyYHgCvzKhWhs4B5IjAmGVYXsTi92rYsEnw
eLDlNmkvJNRwQKadnnviTDAgv5PjQ6BaFT5NmUXboYAOZPJ2rwbwcEIHvZMbuez5dnmnKWOmZRVu
w7nc/4s35hiWLD2DxH3mjJMJaNGDWV6BNHVcgJNkbEdBCsPir1TsHFuF6ZSgCHmbq8NQkV4JugMU
CPYT9xsRdXQwYEwuGI0Ka5EOkw2GNfPWC54zJ15bGp5aDaRAHPcPA7WMvdRC08uFaTgY0zM4w+E3
wkFwQIX731ass4HOWi2iR/GSBitu5EykEBo1mPmUECbjqekPaXi4tjUa/QmjPs6A1azNTMlOAu17
VDo9Ee7LFj1QOKxj8cNDDQjeMR42f7FNNnWr9YUbO2I95jJU7xpSWWM7BsGcFZvtmj7qJ44p3zuK
qH057lBU957tbEs3eJMUWVmsOMol50+EnYv83CvUDAOHpMw5YnA7cywphP1M/3W7i4MnSJx5bhGF
RTs0grjSgyb2uyX9XtV0T4a+bEwITJWDtU/VkQtJv5F9wOtYiOzw/Crl7rAtx/4iUlEAlRQvnoSy
FsuwaZ980Oc47/qAkrQS+k70j7U9+Vre7b4GAD/sFy+E0bGyeRDApsC75KiMzAmPvBQRsc3mUHT3
FhZ+TIH8nGs6ZwbmKzi7/egXw7WXavQsTnkBL0iMG8wucm2LTNx3wwr9jjXri5u1oTFte2EEC2vk
EnHO/Pg2BkT/EpKmMhVR/WwBB7HjipUChWFUBDQyBr3gG/ni6EGrcHtTfUH94D1WwaprZmxBsTsW
mqxClEKNNTiHoKKQmU9MPJQOSZq5LzOjbnZYYUWfxQi2XgYL46Ny3ja/IvKnbhl1Wa/IjpAG8d6l
Ni/gHAwR0LTgsNsf1TfymE6aLHvmkuXtTjy1GA7fTVcjdRSXaBEr1A0XdysDfwZ/4ww8Q5Kp8K11
pOurvMo3k69ALVj567itlF/nao501Ire+2lyiBw+4iZk970Qe9L/okkivL2VD1npFCkgmaZti6QK
KgEb6LhwU3+ru1xZc7Aq1KhUupGA8ilYmNNCfbVj9yOG+CD3bkie6nR10k/lCYTahQjSx3JZSYbe
8Z/uy312Qe7xUz75Ujf3WIB1+/qvEuY8HsJAagDfaPnfVyiLfM4wIVWZseW2TJ80JY+GFBcekE0c
I3VVuvoSVE033/R1JDB8NO/j7Yh0Bcf4zzlc8NdzeUQntmh2i4UF7MtXxm3nYt/aLU6GEPHnXq+n
OH3zwM4rSCYw6uVllIL3pIiB+YJrz8+8vJoZ0+9j5Dscj9nW1TmSvpm9ClNVsVqlBWIByWy+WNIH
f5Hws5NUEcpNc8PL1MZa+TF4PXLWVjFC0yGUNxzuprC9WtTKxU8Ia8dc2QyDJajLjoazo7Vpk0t0
jhYTKT+F3uexaNwqLg32mNt4SXbSIJlrQwLandygMIEtqWW+aDQ0cwNrYRa/hLCdATuSN8RrmpEy
9sYR0KSpINfNqb1v/jLolRs9IuURESRhXBYp/qWJJNznRjE4+ruV0fug+IBnWGDSD72pPqhIIl+C
GkDXYNL0jF+jqPI8NLYql5LU63cx2h5vC2alOXtBsftO6ofyEhaWKHSQnVeH76CyXsmi2tGoiy74
ALNQcRU0yZuSEyo1v6ehgmd3+aNiqLhtSV3SCllxt3GePjrotq5y7qlnreMhA0qdCqSp86sPnQeO
3zFr74yVf70l4fz6GfFMqjaGksLDKIxKGu7g0IxPvW6Qoo1gFdCiKO8hFOOocUPXwhr18CcGiNDu
Mzg6TnrSrrKTwlTF3R8um0OyHSz4zEQAlSUABKw5osNta+b+dqE8118eKBcWG4LyQaccsaOn7RUQ
FQmwSDr2nvxH+LznlqmgPv8T22NMDoIzyR+mqmy0WZqOdD6Kcu68gh4eTCMaLgZ6bymIyXN+4LvB
0xFG0Lg9OEzfbPGETmJ3goYdLr0b6Dxca+/cFRwMTBk16vzG5jB4xl7ReyUNuF3P1Bz/nosHDrnj
KQRt/fp3r644TqCGILh7k1HDydFcoW/7FEY9nkAfPEx7Ou6z7ljPH6Ouz0xtK+A4IZ75jEP33ewU
fmCR2+UJUnA8geWWcgLj3NaFb/SSLjcRIsC7R4mGcmIv///cLT3jUqCIhOjFUTirSIx8b0zrT/jh
ZMKgirPLQ1oLYXPO7PXt+OaEoe5KuJtlxR8sddTbboeRqQw3PmPf+XwpyO3PBy0Nz7KV7HB1ukP2
AI/hyoGz4BzN6A90qSlCBO4XJy2YgvG4ms/bFzP3U6ydHTkg7Le6YFuuKArJzF+eemdBm7Vrb5nj
Gwc8BOMmUUMKNfj0TG3fkdmo6R16HHEDsAtZeJBIWnVYmDX519rufrIyx3VcqkQUTQdYydx8qKbz
t4JY3AJr1vQGCt87a/WYO2dKd5x5AAHmx2fPlnR1ylSMbcpDLqkW1dnn1aYtW0uyBZPnme1UQnVz
msyD6RZbkp4yxj83vHOlBzRBTO6xRDUhKydpTOPlrDNp9tMuz9r79unNODmz3ddfBDeM16lQ6UaN
up2E1eazc1BfpmXBmGGW8Yj17tTRi4coWt7MNXIqTlah3M5NW7jdPP3TvIjUl8lf43KP5GDYYLa7
hhUjQsKSfbminTTKOvtUFmJ3NSUXGnwg9jc/slS29Fn3Kge9jnZdfvFZqB3Nnnprhdi9OOV2gSvP
PrqmaO69JWEEpGr57KXpI7CGlpdhJvstkH0SeYwab48X/MBBrydNU7QBMGFS2cSnHu9MHjTFW3/m
Nfhmk/nB3cnvx2MwfIV8mZriV0Ed49DFVeWFNJzDrkiJW9HiEv41DUY/goqr+0pBmiU5PR6Smk+s
pnK5eaScIoXUGZcVrvUckPNWDy6dTflbeZeSsWBEKOvkAVKtxIOsG4ez4WmI9e9++b9m9QVhdp1e
I/kYPfvPxpM5ATWqalgENvRQeZGGL2czLjWuJmCIRFBUJnM/mBbA6vihd2P9vy+n1GgqBk794ku3
LdXlBn47rRVoVPdNxLFIPwcuB/O6uravDD/9/G/yXLoBSACD3z22QXKoWzjhae4rfjzahWQfxIQ/
oWeFWuRC203wdNQ1MGNtkHx+eCSNPL3WEV/mseOc7kb3Eys344V90UAN6CbqlY5FtBeYajHI//3M
iSP/T0QJQ9oY7VCirAY7bumyEw3E/6FVAin+jd7f6OpBIFf+deNc99sgQyqQ7X3SSJrVGUgFxJCe
xLukaN00bPKZVmvRmCtqtZvO0Amp/17YoJ7zvdoJHF+b95cb1C0CIRF0wT/+j1k39Hblyy7YB1o0
chTnC+1u4Kb96AxgeIDMdP9VOe2yGbijdS78HMbD0d89XF6TyVWg7tJ7DdVhTWCIfgRInEMFUhge
i6HnJ09llMCqPsRJW10D80OZ2tKH9fsgQh/+PtN7TMiNGoI2fLeSTU5poPyWTudkoufPk1WzKjjq
xxHErA0as0b7/CGuepiKPDI5TvimiyF9MMWbw3/JjxWWsdrnARTj3iUyEEm2yhUpQAFjtxtGRJ5J
UJGbNsxs2+twFkbtb+Z20vMmRV5Vxz7UA1nUTxPrKEgp3ydcp/b7QsmTLUslzY9UVL18TcTPgalZ
291BBeEescismhxSEpue2b/3UbIv9zTg8SecrFWHawS8gCrEzsANXF5uMZizyPPKLT9PsoNGO13N
IQtuUb5Fet90pOGZ8zmfvrlZL9j/dFWHjaCii/YCEzVxZmuYOIi+ZiddcNECvAZI/w9lMW2fSjQm
Lv8BQjqJs7CHLuqm+xTaCRoFLJ8+EE728EcBE54bNUdvF8YM4Y/HaRgfG9Ki4iUp04GZPwYAT+db
Eozr2EbpiyA0GSiDxL1abzKdFXVlnZoNXtxPZzMhlQgZrNdd7N4W9we2D3fJ05EPLF/jORud2ER6
qaNXjb4+VZJRsKD8bmhQ4c1o/NBJ+TMM9mQNcaVH0QiXc1YJfsw4XUWRWAiWDjzUwpYmkclQ9m9i
+mcIHtGVDskNh0+2UvywDOPUjoZEVy4qqIzFVu3f0GuEnffDqhiV4gQNyc60jW8f+i3nslFqs6vm
6RYS2kPO9mZW0u8QqV8UfsGddpkmIv6VFPZKeQIFkbDD1f4AVZItre+aCa/lKmLi1arpGVgwoiTV
GqI6/sL81+RhXETg/qUcPzzc1MvkMj8DQkipQTQ00vEyxpgXidh1PbPcymlfMGWnugCvCVZnlPPc
QNE2kp0ohZVl0T8hJVqhM0n9AV+0pdD9nqeH2L1q/aJwRSCgNZExhpK7YWTPmFLqFLrcahjTzzeA
8DRNu2a4aWqXPEBFniJcAZiXyn7NmDfT6oJNp70aDAM2tckVXPxSS5q7mww7/cBmNFkpTmMf0RO6
k2TX08EALlxlNh2kD5cb+boabXUniHen0i9KRQKgofOWsKlWdYJtyrKcCrRW2nssvywwkQ97RSsz
7vx3eOfXz1THBUH32V2q9KVv2yoPB2o3FAcEvNP1WkC1oTmYiD++Lhftx5BZmT/JoookDZIkMWRz
xfNyvPGzn+9uA0mcPcQMwikyH16jtglPnSgL0RvQBJ2j/fiCsfUoge8g36Axe4Ztq64xjzeH4uqI
bhIqzYoriT6Y6KPpHUQ4DEyyGWIY/NGrXPIdMf5T/5ZBdO1rQAprO0Nx923nOkhSAYjKW+4e1K7n
SByuSfPWUQZjbp3fjUrIgKoMrPfHRVoEIMKXiNaHG4wy7p4UctmI+DhSHI2A7gFPXPv2ivBsNHt/
+AVzPwHVd1y1OddjL5fDzQrhSM5bKJ22eC2di0UoK+yNK1CpeNF0uLNCyLaH9NACNEKCWRczNg25
KXSASbiklDJuzmlbPvl+wJ2/g52634Fb8G6ykl4wM73W9gax0qEr+ehexjpK0PVibayWod2vvBUv
s72wIennn3KK1sWWxUgEqUlfuBKKdtTsLdRCAntviD5pTYM31Vr8fIYE5VVg168mXiHEf+0fTEH4
J372wb2t3vyJDfOIVzkhXPwJBgNYawAuiy5bmDoH1vz+8gGCnz/SCQO7K31+eVWaD+O6s8CYxrXf
Pzitm1ARqYE/W1s9/NHRnLPRWzguvH8VvMid0VjMr6rdet3hsGaEOroxv+7TnkGjaj/PVVk4LgXi
PmKlltGPutRR++V4Sw8dTMHhtJz53SIiaQy72TZ6L41MfsIuk/61hzTEstacpbzFG1JhZ1b+jHZg
Tfp+poS+aFDWMhCPtUYwtVshol1oXh+VWR5kcwT8h4bAaZ1tuOunVrl8hUToO0fDkrk2+v42q31M
0kYjL2KP4hPyMgjmUmIYTonvJIxdWfqRwA/ELfXl+7FDI9LYPoTY51LeeGsMUltCMMdS6sgfKZ1K
Agk5mmuL0e2Swj3Y91yIwQFJw2O6mKGGgQ1/IgOnSYjOm6lahFbu9/m8yXeXvcfiHE5cFZ4maTVG
zEgUB32ALLSJtewgVlWt8Ms7pRo3HFrI9j6kWxVceM32QUm81CBJVBw4OSVmIBD44pb9MQ32Q+yG
u0ucU7KEKGCKKsQhjhcj1UhHBoclE3WbEXNH+4UXQyRpiDelburvivYl9kEmb0zL7/5EwwEjUeDN
Uez/gZqFhSi4Ju82nvT+hEhnnG/fcqLNQJ9uca0b3/Sk5DeTHioIpwPg1ncwDCxRuIfZZ/SN0xoI
+G/vt8w23+qiz7Y8vPSsCKZ0rvI7InYC3xX8lvxY44ig13Q408QbgVnzsYqh1xGMms0l670baWr9
tEFNoUYDXSgfZEwSpsaNHJi0yvUpRaofHJqhL4YjAf96puAL24gFXNgNs9Tndoag2L6pbhomwRCF
+zumNd0l4yhMtgN4AP5nPTRSBD5f6V4xJ6mKH6S2pfDlF39HMiuFEc07J0JTvDukROCcin/cTNUE
fWDFwliYSLt5fhefu6LemApdnjqz9u0WbbWB56M/vNp4zsA19IongkBqWjM4QHr7sIRSm5pH4jkO
8F9+Wmol5NTS4MznYrS9LRAUGslKYLDsrrxpe/xdP/6MgiWnYDzcIGKEtUmLGgY68ISHoI/1gZxL
0vbPStket14nqMT9b8rzN236Ch88gEhnKChR0lyTOvJqvsDh6Z0YGhIG1KCK4UafKWq1emjMpTgU
H8sW1aMVD/B8c8Ar+LRDAlEDWc9ntdFco4BfebKGzVJQiw2bFM6ePseQ/cpbZaw16pdci38FdOTR
rXEiCNPDuctQBTS3kUyF+f1jLu4bJsXjp2MevbH6KgcuJHWZyDUChbceOwvkvP+dJ+vBg3/kTXLU
5FshK2nBp+ym//4GP/Ufj28z2Ot0jcaw+PZ/kOUF52Xblfp93l9VTv8OCm+N011+9jEPDOozT4UL
PC/KptELgJP9jktfJ7aWx/E0bRqF1yI+Xn7FCk2/f08kMqpFdNySfnDhg7V24i5rEOhlY+eqFaV0
wUM/GJ/LWeInXzlfw8yDgKC5FbJCps3481goyiPumkiP7UackfoOnk0PzruaD20p3+lkyiEkLvp5
7dzalfjXUGAr4QSN68wGFEexma0iEog5SJOc8NNSrcpspSzKL2OT+rvdH9RhqyyDqPP4Y9PRPTqg
qRy3ylxAh6S5mgl8kq3SuM1ghsLRSs8WZ5ruJVdAJz/UyzYV82xcNXjcp9I2kCaDUnozq8JcKqII
3NLeGBIHeSyR7lJq9hQ3lTdr0M5G7Ow0I4lZ2mtczQkBIc4IR71Xv0BgW2gtdSDmdiq0uq71wT+Q
xVu8yM9gTOHwcfl+cyeLlnzR3W2NUcS1/vXp//NirfQnjXAVlOoX5+clj2UIA33A6qAMpdwZkaL8
oQD/Xi3zTYFHqBGHgloVykBdXX/FgBjVcZCbHUTzILqVQSXeVnwVIRycPOhIGq9atiIv+HaRDexc
SBwya5tqsJ3JavMEnTwbnMmKMxFQdZxnGl9Hd+Jdz0t8H/BthCjh0dDEO9z+5W8P1MpKabfJlaVC
FZtGuJsbxVoCKLM/Dt+9lmqoU0d0xUKmfPcPKg/+uKfj4QXh43C/VCMNDxzACEUW225wMwqPAcxB
iwHqqNrgEFpsC7946a5NyQJjNqjxdnhv7bAGwEwea9kQPQ8wVpQpy8rYK1GWemsyfHK2oXIWGdB5
xobnYVM3rd9nkF0QQsQ7YsoQngEn8s2/vz+3GUxXw+MGVHJ2mnob45EXIi6pNQZUL4cjIIhovYKb
mMAKNPZhnX6cDcrcaQMn+tc51vwSdZXNeYACtDFWtSK5p5a3NcIIJ0DCvV75W2VAFUpEOd7hkBth
JCVg3UM5N6EFrBe15YXJWxodZgkdkUrVmMuMGX6wy5gBSOXqYorqMTp6ULzZBgwGRWqK+nMl0v8B
CmEN/ECOfv1q985DjOjNB8BeT1D0qcHndu1t4c9MQ2eGwlqhNs5Ql3Z7a1XeY2EAX563sEWAP52W
eUMS3qy2POdxPOVvHuxdlH4LNfNWyQL4MmoQOf9pWU751bi/3Vsw0usT6ASzgYqLSgVRMLdNsTrw
S0gjgeNuoUwmEqRoW2lerHaAIFPzxXTbRTjFP9FcQwOT3oXBLkCXaV+Akxinh4xGi9pTvpB6vqEy
6mKV/vtlYcvrwuT9Mn5pon3tz55SXRDMJT4hDROJ/38uQN9AH+VxV6iospKM67H/QiXTQq1QFltY
4b+Is3lZx6XU+wEn8nABsuU/COwv8BBa/1OjGppIhWpCmB6mhRj0Ef0mXM8ndkFtgZgdASr/EO4Y
oqz7BuLsTR6tS1xxygYulL2TpIDd9DfNcyZ1olH19/E0bwnpaEbxJmGNzXygtoBp3KKA6c+N2ro+
PVfqdxLirOUSkONdUum0P5SldvtG907EPIHqynC+1zbtBDrRxugxoDg/hg1si2MpTJyfeoF1i26+
L+qaVBNwTAnhz/wypRwbUKwN0z4bpGY51jM5aJEFy0lvx3E/bpPoiJkeaQxmDAgs3Ll+u8hyM5rB
CowWqms9BSfo+AFuYM6MLob1KYsyR7SZAMLOzVHL02RPKUuP805NaIjSjSXL+v0puA2m17nHiFVH
Ss+7LN9s8NQ2iSjlWnjASF3pUNoQttEMXoZH+qdKnqpTiXoV3E4LrwSXv1acsTgzvReuknh/yyWs
sNiGFhqnZO9uuCgWrsMv4jVbTJmRO5s0ru0/JLc1IpoHZR1+diOyKhaL6lNDYabp/GeniySWDAyP
qTeJeord4C0ea/ljLojbXoFJDAGMdW+98iucr0AcvwZbzzi/ZFZIm5tJ6DHT/nLrYtdhd1+5QzhW
FgfNZMNF+eCDRGDhSOn8jnqd12ZGX/p/jx5Emj493mpIZ0tV7/uc3DEKe1E02gTMms6FJoTi93re
Y51bFL542ihDhm9C2MVNb2PmVHbjrnSbVqLSFTuUY9OLQHBnKM8myj8FSV2VdPOJgQ0XELUmrK6p
h2bXjUxFl01wa77kLCeRaLxCCotWB7Z7bwH0r2H6bZOQ0ZAZNXYKuEpXKvg7ePQoBqJzU1w0+vTE
VL+gCDV9Y273kDlA3ZaaqzqN8wrF20bQbaDtYsMdUX5ojeTDx839zW/TL+EgViPvctnRfJWFfmRo
B5PVeLg7GDz8jwGTu6wuaIPRhqtI9AY6/KQSxjluYYq8Ghz+jAMRrYc0oqCgwhCCruT46isqdtfW
XNu08ckxaSMaeVecZ2PH5qlFh5blp59+L54Kso+GcXuMcmfj6inj6vuRZcDCrSH5k5XuDuee6ubt
u+H4ANUi7E9oa3r3A48vHNRLaGqK5c97wiqEH1+A4fXtmLs+8+L6X67liqujhkM/APDdQRu8SD0w
V3BrxC09n8nseWmD7H4jX1be5AlmWK1o22xyFrYH9UmvBJPwBIaRoFLLuVCAApDWm5oAHkC+yf/0
5bMmF1fLBma4no08ZCFZpV5wWYVg1s1b7nOCJaAH5hN76FJw8nBGZHZMhsKpEAObw1z4U8yc4DKx
tfJxSAyqcGFfn/+IX1t9QBnGpTZ86c7jHz57HYIZvRq7k0n8GypVxHSjG6n73vA+YRSQNMEB+D67
CtLTlvWIr5lQvnLOm2f4wFo6ddovwKy9AD6mwfHZl1uYHfazYAEFJsE+ESIPt8RRZjPq0H/T4Axe
U9SkCGoqWJamAXOjlO6DYMXFQgMA80LOeQ/WwRbYr/fOhYUsNaIRitu/nG5hlYrk4zmKS6U7iyvg
y0UhrvrHxDaGlk6eh7OH2psZeZyhwqqHDmkXFFR6E5V6nJMOyMNySGKhB81WUKqDDV9z19/pW+sn
0sCCfVBanikVOCPQ5DOBQlmVte4ngbpD87y2PSLT/OtLgFe3Fgvd+3+9LMgyyIgYCyqSRjKsMm1P
FrcyAFFRzi8avtYCyLbxxawQeOyoQpQQhiKrvg+3UDz3V/KAaVUUSIgkwy9ODNM5Ym4SxTCIb9OW
8fGnozgJT719E6ZTiEtUEVtpZ8evxylyLrt+FYcSzxl7gjOWqCgh9KA4yM9OadlOmkRJA7OG+B/V
G7XTw4hdn9Bqxpqe3nBAnmj6bV9dprhUvrv6OTxOpMeePXme7EUkR6Ws1Zv4ZXWv6exAYLtW6aDL
uhZ5IdK7FbOVUz+a9/HWifdXurgOVb/oSb7A282m8QacGDvAfkmIxnBOqkdUU34tTzULVEUIo81A
qv8YjKnbyEfFHKFd4LfHxV9OZriTbu3foFR6G25f3nnYKEh6XtGRvsPmPWgKYq+L+SZeURk/ilXW
uqlqJWjjjwj3SpM/eezCB2okd9BFV1Cm3/MbiVoCZHNriZ41q1FXOagE5JqqvrsNG8VLFc/PZsS9
SUGEmnUFyuZrLJAtV96pBsm+7h/PmYnIjYWzs1m0qoJ55gT1gNMtBUa172Z/OluiAQ0eZTCqinVE
wB4zMzWJ/n1AF/6vaKZxL6HY6NyfQJyS4xQD0UFnvboEhl6pVdNmRGoKqT0zk650rIHn0OgE8v0u
z/c7doXOHg750yYMLkcAqCRQOyPUNnnJjtBTmobhEgFOOVSouInBxZr2ZeCWqlAglZQP2BLRUu4c
8E9haiPH7WyjOv6oCGuZ+Qzg8jf4ap9u7ZZQ5H0z+6jvZP/iFxe8WQCHjBX28RV6vOcagLCJNK1w
lLej4yAFJudYi4PF4/dA+zePZ57AsKVLuCwuzJ1dln7M1ZmjUC7OLLzG/XBbDeZRs4XQxvR0Q/n/
9BX4yJRRsghRpLDDM9sUItCpzdrXXDGdrKqTmKeKBXO9rhrZmAg7qN8LFa3cyN3fY8MlR2uX0dqu
oNYwudaa4QGOs03cmMfqG6co+dN/upeFdFXN/qDNrmWj6tjh4LtQvjKTgZWnl4IdIHv2IfXFN/Bi
0iYYTe1hvDfCYzMSW+dhUPEmPzsR/RUGlmDYkeEf6nANSqxnJO2VLnjzyA+NkMpwtQXz23WUupSu
BHCrRpROT4nACG1TjCIrLyoRkGze9YM2XzQYzchjdjZJ24hBxoDMbiBOqYBDaZ/7jAVsxXJlauy4
gAYTf5GGxa/dlgt7QPknZL155mYLO8ez1UY/B1+R1JfJg5tmxGr9JjOu39U9rUkmuYHhBPkrT3uW
JxKroKI8sQknfKs8YI5KtG0zBmiibBCEbk3O9DiSjJJnlGZ8lk0+5dv7yTiM6/qLvr3kv5fD963+
jKhsebGL/nXTBsVOrNnxxecAZ2tdd1SVtCxbWP0aIWZDKCZOVILEAJI2EEDpXPhLJqUjlUqw4x/U
BguXuoKxWQqi3LXI9UooAnr/St3tazGLasybaLAMqh20E+RWddOE7IdYPNC0ePevI/HVRU/efl+e
fVWEJaBZxdIikBSb1mllOv+4n2k75Z6RiFnNqn+bFbz7OnRsOSX3aDSnf39obYizzpwsB+EKCHxb
63Vq9jcjwRyuiEf40PC0O3QSclt2OlMDIGbZ9egA15w9NMOzlPyqYKkI2KhlTfmrani3qJ3IrVmn
/Fc8wpWj2Pfc/dUSBdp5dnaJzvceJOhRgya78jq107ueOkgRoohpUWxvlozBeQcZzca4Dx41vcdk
wbnGre7EjqlR5OOtxDmDVkYjOq+ZwgCJkeKwo4p9u1TC++jpDwqbZSvkW/dE540+ldCTTxz0OHAg
wGGBjrdcl2UH5MEVanMNKtTJWr71TNstC06zdZO4k/8DvIRCvU+wOWcVVtX12+qe0nsmUZmllcNg
BOExATGsDUnAv4rJRocMxSRK0YMAyk7INc1p+EW9UjdA9fJhq1PP/Box1F9/lmdzZOffyTw8KN8e
6POJsxWOzQoWhNqB5JTQetpoGdR3IU2qI8MA1z23uWtJnSnkWdildMppzmeUt4K5SdoWTCWc3h4c
LVcWbhDzIVt94UZgy+AtuuDZlHUq1FrFRd3lYJsozkUOAgXdbAGURQlMBh0Rs7PG6GrgicG7szYJ
qt86tMsr9UW6pLv+GiJev/+Ozt6CLoSvUFS2Lbt3V2EqBhyX58kDUi1UnRLqeIG+FKXzHE0A/U7Y
P73glkivrZBgphZvUcuFVue6vnp/LA/ADiGelHR2CBKHPtTvx+SA7C7MLEUQng+Ui/I8MdgB9u3T
9+XHrFELTZ3TCd1i5PC+/pl6dvRKmv6p3mz8ecehdeVzzES+qKXsF5jJ/dZm5tI/rswmhEFE89rQ
E1bxM5IL73PlyDzDLu8nq2Vca9u8ECHsqiF3QFWYKojzXuY3q7ir8F/U9Ui0Yf0TUY1JtV/6ssFM
jJah0LBg/zHp7l4ssQV5Oc0u+Tyu5EUffvWMvGwD8/hPL0TIwvXlg4SkTMZGtVCDqw26kUZGFFdc
z5WzE7szCDUnB86/386WqsVrUslb3TcIxvQL3QyoBGwTj9o90L1AKcrRj1A5PhY+9CQR+ODrNo5T
YFTVJ2DdTjPay5KiYNHGwt+W/ojYuOx9/4p0HYwe9B8Tm65ORXf6lEuF6rB9e90CBT1hD0MSK0bW
fnsYuELX3f2tLZTUrW3jRp/zI/ptHwPmWpSdvCanIRLzapbYwpAlZe0dKp+pfQNiK0UrEMfygQBQ
7jl9n0fR6EQ3xeH2XmVEp2UNzyGGyLjB4w2MJlBvUuD7NWDQlFLFttWH0aSKvBSet285iJUKz8KI
IRCuR6WxjZS+4t3BrWYh50UMDIq9bzQ3YShxqFCU26EwNBLHqRFbGpkO1uCSgsziBts2MzDqg+w6
aTNjfBltfqWO8Vj+bcvh0IJewavYxl2/qHTdqJU/WYCPjS/fnjaGDMo7vC9QJBcntTe7u2242Spk
cIrH/3dB9tgZnOLFo2At37FMGw3I3vRStQ225fn1LbsI6CkHM3R/mhg4ra1doYXZ4RHEuVdztunP
xnUFeE6NUl2mdLZQHeOb/Hr1kB79hiOjnj6Bd7msoeCf6+u48Em7D6T9pxoPTzNstvsodHDMUb8k
Ijfe/cF834/JEHVled3eyDm5P0QHDhay4yxIjFw6soF+cl/UMTG/oMCm40RkZQCg1viWQyZIBFgb
o5s2n7j42w9T0D26hHD7zhlP8UxZkjjQaMR2Z5IdBt2HXthBvMYZHWJP/vd7Rbnib1oeQqq143ej
t6rG86wMCSbxrYOSZawUqNYgy8ZeCjFJJ4LKfFXwnEE/zvQlACxVWv4x4p7iqSkKdi6smsJ/Yv1e
WJvXKlf09Vp/qd0Wu7kzHCgOhTAXbou348tzuBWZsn8UkJj2ZDUfH0EHAQo2uN1z6HVll5JiFJxN
8PWDPJ17sdkxKQ/h+M2oJMBXnWyFSZxqVd3SvwK1dSq/RJf7bwH3PzV6n3fx0BYsER5BJVm3w5Tz
TiB3qS1O2KktWxOEhJ/ZPR7DS8HMuXakn7uw/ccJHtnhJK0HVq51E4OQ3CoNcxQLei8cMbGdW368
KhvRroLNNUC9NBNb8BwKtl06h1KVf9xlLZk8R9GeEt+sMGQkDzdP5BL5AICr3GAFIibTe7paHBS3
aN/Uezfrs1bNhOv9Rn+A0D21sQvxWUnz50euvFr4C56niadAs1ofEMMw2G0OC/GUUVeW67fP1NeD
tvG0T1REfQGuF8amLB4n+dBP/mUxmVURpFj9o13JUAM0jv6EfK6BAbNj489ozdPHPz5QTg7xiSfY
DAPGhsJ2bLDQWovGc/5x+ejeRQltJ2bfz4JhQBjC047lujoaaR4zHbCmGynkFn+6b2T34B01cckW
Tzp67QuHRgT7LOzOcZilnhwFIKds2HEZXHIG9mlHVKCm2Ca2BpKqCWtMw37aDZqniOvPb6xDy0Ag
o6q6E3srfVjhMiK3/anUPjMrYMB+QONo5OQJ10MYrymYX3F+0bUlj9B5RcTcjs4SNs2N8aWWrMXU
NSXliXJAYYsbNwUJpzfvB5iTqdTPWRSeZuHeIgl8OGPnnSDRw3ZLPUuPVmi3GM3Px2CM6zbf17/f
TQCmmH3GWF0Nkos4NcdSPipk01VJPbplP3BmiF/G+GR7M8s2Xv+1PXf4yZzKsZJ3IiHAMGGThe5v
WybgG4UZpQedI+rx1L9rZH9t+6B7TL90VyTKxDHCgeCsSrkLI2Mfbk49Nx/dePSJJavb+jxst1/u
1z/Q5/xMXj/ViDrEt3/eUEsu7EnFkSyXiOAMXC5ARf4SbRGYIZ+8vj66BonDOq608MjmzyOgU7FL
DDyEo8AiyQhK6W2oahiTTVfPb3Pa6IitJfdVfNrgSfpLIssmF4wZwhaoZ9VLiHvhKYt6lVWP+0HA
i5zpW7kFP4dODqfVG88zofJ1v7p8imQltI5/uVpcLRrdwgBOl40nEr0DWezqutN0pB/u9bYQJjRN
6IQJt2qnMcPR5RjiBAewpMMzC4T89vMv8je0paOnMnCbk3BA6qVlTwdPdScpfa6K8TtWOn+ND4w3
v2fMOgL0LXEb5P5h5/hUSue5LQMmzUmvxWlyaCne6zLb8mPI9g4Qn21nsxO0g37n3qsiXA8ypKw4
hpxx7d2wVcH87iQlidNuDZRrp1FF/HyDsrPhqzXNm13aEOegJkl7mSFBOyI9flpN/SVXB4x3IpYi
3tkZNL0WKjAuLPfoDPGA8z97hcCksZEg8LDBnSypg3+D3EDjG14XZmoObukSPh4sKE4aWKkeArVk
bEHwJm8DFhR098reT+FEiVPh0iFjTRI26rwrOWmM00xA7jbo40FWoJikAC1HxY/4a2wB6PtJ58+I
JfVBJT40gUSmDPVuMZwam+aTrBiol9iU5VgEG5/GlGzXJ7Vlq74KlNn4em/O1maatI3//1wF3idW
TUHX9E/9tKolndDZt2Y/QyGQ8zJJgjmV0iSSk/xliM+nfSxq7pNpYQfg681JQIiWIPNPVDzbKzca
JFxWMZSw/QYz35mFUGjW/vtg6ApGalX09X8DcU0NUbdzFwBcytXFx5cRbU/iZGx7B6Je4zkS9EAf
ZqfNjnM2zzJfOCCnluygWVrFGOZorblCfttkYIhwwuDH/GH7LWI5jlwNsAVVkvSG7t4DzVxuV6u+
ivHRYowGcClLaB6P6ctEpFgLrPw+KKO3jik1X9TqBUqmWGXTDIh/OIWKIPHjzpmO8ULsV3pabGyE
kt8ug2QcxeBJawWSBWBtwjNlQF8MiGuCqJWj5aSF2hnpq0HnzAYKg43M1kVwuIxNQW1z+TeTJyKS
pppZJ2LYguTPd9R86puvu/ZXlsEU7v5PvPUc0cFTjLzDD7Z4gkNLDulUFpzshT13VPHU4aouka+O
uy5jHvdbEr4LSP5YzmKOCaRTCNaBeaJn+C/s5jzBlFHnvZx8Rfa6+Xh5BkOpwbdNrZG5i83SfSEC
YivuG8AANWl30o1E4UmuJmTfH+/CKOauxXbrg3cBW7LaYkDFInuXL3EB+v9fEddTrhjAfFKiOl/L
GLUt1ZvxPfNT7NnfFMxn2y0OskREglF/7C9+1IeQJPG/989WhXnoEBVaGb+40FjZjSFWnH2kIauC
sfUXlkAdu8WRI+0vnlOhHl17yYGBGBAZ2u/WMVhrSAwGsYw0bFzW5MUdDESK0ZAkHJVOLCwCHDEm
K0TCGkAxYi2EYYhxwgpDrWxKvqyAJy6ke81Quc74FaGSygIYBTQP7dl+yQOeTq+NgHfcT1fXL3MW
RfsghzNtv8tJNbsN+tkHa5ldQ5P+cVZJXH35Db+6W5D+RsYUTLoICcfJMqUfMhdNrNIs4c0UfzSC
CL2c5Oz5MHXVxqeJlNLy63IcHcZSviIfBrEopKeDiPwwyY2KcDWMlT7osEs4q4TqXoZms6DGIL4M
9sXIruRLoG1fd8BTYI/CBZLXCfZ0G6SQxNL7p7jwLabduMju7rPj3DxsWgEVuymQixXGC84v3FhD
YwY18dsfoFeqHzuTk+hbRB89+agr/Iaz8ocdjoyBzYkJ/+aBxaZ8vzjgyvtnCClIqGPPIGoRB6cN
2dr+vZ/GkAJtQC2FWrp+l/1c7DiRwLaI3dHU36Lwp6+IO6QcpbW6JPIm+nmqA8TG4rlyGRNvTHcm
czOK+hnMYA/vHufxwnpMRbtXgkbQeTnXe+k29yXGyhMI2F20G4jYZMqhxa4ZWsCN1oeJjgQ3H/GO
8JLfPfJyEp+bUz6bnvtxhqxtHBxywy37jT/qO0cExQgvbREeY9ibO/aHDEj8TlMhsFq8XP5GTCh+
EyjnigdVnnoenpaQo7eboTDiTHfPRsdP3RBI+V4OMUK+Z+UaNNUs0IJcfV/sZhegGybxIoqZQQnr
m/MNRGq57Hqrelt+Wuv2yQSflGlK9l1pFgBow6QKjSfCygzHLf8YoGj5jGcSbYf3TEvsryQel9LH
Ry9k6R85BcxFtYEWAvgLdFnoS2pmQuTQ+zmk3TMZRPY/8dDJNjcMC//Pe9a3R/YO7C6tL90WinQg
ynoMSkUZqqeTeRY94WtegF5xRodOqE+F1pX9hAV4O8ikvDFEbsZtheNoc/J5s+oCPO7YiYv+WxGj
cVpoMZGRPcW4KHDBeMWj0MaLDzu8zUsCb6FuDLa5FUzAz3Ae+o63gfl/21YuXSQgYJ8CfrfjDZ+1
izBvvCACv+3F+9YXWaTIQUcnWhEAclcsdZbrOnmqPrL3l7dGzCyJAMZEdpGmc0OZ8z9uomNOKaCW
xWEr+zYkqF7ue7vPoG85hvLs76o5oHmSLFRNy8y5xsZA40L39n5TG1ztfP+XRc4CVq1JlQaOJxZe
bQNtd7BY1zvPUHt4NC1rX7oSJpPDx5EXg+CidyAK0vWJmqKOtwg4jlri5+09l9BYiK/V2oWIVuJV
+7/VB/kjKi+B67QlwBauwGg0XkEA0bPXmlbzOJGTvnickhEy4XeMQ1UvGndgsvSk9Goe1WmrdEUv
W7iEaRLCveJsT3TKNoBRtLHuqEs2BRt12O8N05LNAiJvRL1MXloEEPJ0X5Q9hSqw+SRMYZnGuKmT
WoUL9aQjTfQERqNYUC2pJGmuPCVU60nbVXIxzPVQzMzhKcSHJ6DSm3aqZ0PfMBkwuGJ6u66HZ/Be
1NeRyWCAnF/5oLmwK+GncTZGikXxhMbPVIbmcpSS4NRuDnWKOaHlUB11xXzNzXFiLs2npp8zcXDb
46I+LV5LlWuBzM/CTnyW5c64lo3rkb7a0EZcJzRa+Z1uhv1gUk1uqjTL6ECjHz8Lg79SMZaAu7+1
UywMMrLOZTk0l8yjXwSLejo5dGyWmN+nHoWeYB3u3xILq+T4SHFTW5J26GyLraM3WKCgA9YzJcCZ
pN7QBAtGD/ths1IUC3VXwrSX+e8E70pM6r3A2sHzf6bia5g6yHoLXm7MmJo0790yGx+9P9s1jY6H
LsLMkQpxuba/dyYZM4WWLMGpOez40/9c/i1Q3caR4/L8P7day5NM7l3tRYh0jYSNfVUCvx1uBcTO
jzHYULmQ0UIf4K73H2S/PmJsstuRrr/SBoVHS2EyLVMUmZKdGnVbJonIHhoOG4ZXiXUXV5G6ss+7
qd4Jp1vZrYNwVMCMLYkD7d/rPSG4jhBv2W8i+H1jIYC9UeI9/tJGfc3cvMQl6GAcmUdBhdlZoXZG
4QCURm0RX+SctPYfnXcB21KAfAYbfqOpmh2twjGHww5in5M2Nypp7ecxp0iTMjEgAy8sLnEk3mt9
ZFq+aYlzceJ+8stqoNZWvv8t3T2TpIJ/bjZMKqE0OIXRHJQ7hhzScIByw1MMTfC7B/hybfXaKGN4
aMOdejryZYjKrhr3Y97rIObn+d36vLuY9TYnC6edvGgZaoUgNckDJDCIbvfkvgHjnKtiaKwiZQhh
nNsJ0iukjTFrSgtRPup/U+yp0jW4c6dCCUP9lv+5Ppgjn4hlLRHqUG3+PhGhKwKCyFPbzTHdUdis
DQk/F/+yp9ENc3kzX+UqLZ3UB4jPmlBoo9OZTuQz/P4k0Mmw/ARdDJewQ06mXXcEt8a4gmNLXFxq
4+kiLh1KJMo+R2GbWl/gmPsiw9pja2zVxhzyzeTg8Y2S0qgqU3Lwv+7akVqCncM1CorghDUMXZaf
AzOrlkYzd1KDCPvchaRlhNXuM2qmQJ4HNXqe9g1pKYLYgbMFGZJP+LO/MujddoXDz9Lf77rASdS/
qn5Ma5HJDvNI+71tKF3O/1QBQNX6znsopJVOrBKCSS6/sjO6CThKIp4ims2H74mM0bIamI2IxHZx
TsoAYNn+u0czSjicTEK+9nCJVuTEbbYpEwnD3mE6jwyG+4YV2WPzRq3K5ruedgYpERVAR+fL7Gzd
X/2+FXd1C38Lx8qN9CW2u0P3+Ztgkfv5o0DmA/oTfmt9ZLQo7hSyVZyPZYt3xvZsdhLYNEkR0Bf0
kT8oWVFG5zZhgqf+GJS23iuaADCJp2rkIFLkE721i8GNDyY/6HWJbRjxz5BPvOp7rvhTjZ/4I2FY
e8s4PthW0PV5LuGRc3gVtx6w0jFDHsYQ1N3NWmKMIWgObXDq+iJVUHvBtNOXuSucJT5u95wF7aMk
YjXRq2XAXlw6dAtWdtn9E1hpHG8TkbFIRXkPJEUwtd97vPGQV2PqONNZ6YBUgvZAnsCsHyydw7sp
v+9RC/XVvUu78DBxUygri3/iaPdScgVNIyF8PXx+oqfbM/7CdTCjn8w5w7hGblKLnZxs4pPP7qe+
/lttoXaabTKnk4y9h4yvuX108EGM48OWy72P+mVhGAdvQHcTaGhLm3BelfLBSZXsmloCD6yieA5M
fDvS1Vc2ozA75MB/del07sgjb48RsuSgX3YV1J61YuTshg2IfJ5uncWTx0oIYVb528cMsB9aVgWL
EwdSr9kDhjJyFJ/k+KJocYulWJRxvAs8dIBMYkqvy9lEqRFkokVKzS7MPoNucuNSaIGruLZfIIXE
8cduqBa8ZkYIvXpDX9vDZaTVACVucQ6KiHc+QAnu4vuSeGG5cvsnPlIJv7CPdI+sDrKwtBdL+G+o
ehUwqaw0bAMlpodAFxvglTkqmUJFSpmK1uHe8JmPKIiQ9t7BkdFXx2CZRdgk6JTgtunOljZErc/H
zZNsaQ/tFrpJQ8oW+1a5I7M2rjKpfM+j6MmM5sZtqC5Cf7mvfuHPtpp6KZnxEQDuCMS3ZlMBgbYM
f4x0dU+7Sgl18UDNU+7E+Bkm5nZdl1gzdCtwFl7tPyNSpqC6Y+DPUlv+ejMyLm0zwkfbGxG8rC7Y
SeBR8IY1uxfdWTO3K10gV3ejomUyaj5MJwuXB+bXgE5zNkIyHM4o85cnlvlrIyA40DdZkyD6TmAA
px4MSFtBvW6cygL7NLHs4ma0+7UaNdkeDDvnp7rdVCqWNRDReVP1QpsvbPTm3+FPzTUtX46TrHd5
oQbaIPtDGViVzVqRlDTJI49sHGZ75DIxvEJ0/vdzbh/iTuvNNku49GoMrgVlYVzBY0dKqem9kz0x
+wX3V/UQHWUonnk0/P/SCddcn6IZd24emj0xjeRvAoCga4r02LauGeyZLkWwMn63Ca++knylYrmK
iDqdDKRVCw3x69Doy//ELQEEUnaQ1L0686FzJ5yZ1f2xactkvgoZbfePnYYXC+vabSoCleEphL00
mUnXwtXEnNpi+zHkZeeE8KAeApC4g4BY6dRVPM0aYy31L9tsBeOzjHSVE9J6+HNI1yQ/PafiiMGu
3SIzQhFeqDgI0CjMfyJjP6LABE5nlrvs1K1up1DjXrLZ37a7sU7O7Fbjm1jQZzyOvBpKZOePI/1N
oeFWTfyRz6OWBaMxoYFINPbo1PvZDVjeXCGTFzbGkoaqn0LHgrxq3A2c6i9r5yp/3makHPjXNlLE
yVzA0TO6qm5NvLzi3fPu5j06wccptE1Eb+WY4hdK2ME7dmn+EYcBDj2d0VXp/QiZ/viQ8U2yyF8J
RouDJNriIfKL4jvOhTtc7NPd9s8etv4KpGbEBOsPynj734vnKpeGHmoa0FZYKo6ElQGakMulFTQB
HY5vbDPCGIYGkEb2992qU1A/AfmxgPTm1ogmfDPoJ+aNhnxej09YcnqfozuDcAhu47B68svbEKJ8
2VRbEAmj41oyHzExLO8Vg2TISPeonBQ99uevwSR1vRO7RNrVMG+r1eN3Am1A/mZPOGlZeS5sdYNa
bdGP4WKDj7RLpAJJFv6VBMQxvz0ViAmBx0Z3wyDK96JrqCCB3QCiS/3f2eO4s8+GuNM6BVYhDovI
dd8/zlyQKa1jrOGjDtwPGc3l7TTqHcuA+YBO7CgomdF6O4WP1MXDJ6t6rrTzNEBp+L49R973aeyC
tyAVYsdWD/4i1b8lk3kIOIAuSSaUzG8Sd4O2w+Xaj8RU4sZgulewxOsuFn3ITkFG6bAFCrdfmfRA
StcajPpnhkQPfTLh/ZGr1uxZFjcT8/dxHA5DReAS3U6jSb6vgbbcW/XE1WsSAS6JpfyBMq2toaSA
90A1yLDDEAo0RUsF4cxziHMjiOqBbYu+JTg1OJY2gr2MlnKTwqAwrCTOpWvS5ovu9JTPEV918dSe
DQ/f6IVlar2oCQ+ED8DQZrPGAh1HT/F7eWyOag92e0+phFteMZpKqozzji1SOz2IfqzlowcjIj6t
A2ykzAeJCp+IzSCL+zdbIwpUE+WIeAquImMFcysxYPOSvzowtsd8ZbsUR7W/TvkXSoZ+8X5ZzRzi
J0garUIl+Pz95hgL95RLB3A3k5KOOOKOyIxOj0xXLGuwDHNKaMWcWUCKtrIUqR3moO8REz6yCLOm
OQo3Kqr8gTAm9lKKsTbSdviWKj+dn7Iif8Ub1pTyS7kgJ/LDjAAPuQGjE9hon0+om0QGxkskVqHu
QFrBzG3f6KRz5wloYgU85VwdK0U/9XUO/OFvHQkOoIu/hDDIsuRe9FEb1ftLxKrHBAzEI41S6Z/d
XBHEwqLyLwjJkNFVzwNpK3w/w3NCSCPHzPOZRDfo1Ihy33cuJu3+W/Np1VfcHDQNCKMkfPKTSi0g
Z7V6RMNt6HPWg2TvAIzdkx4oW1VbovqN9/qnrmzdfkgsCM+Xx0UNNWngwoOAVkLzG9eZi3NBUC5i
ny6QIFN65I30uOYerkhtVPMS6fQZ9NQ3/PrETvNO71TNRZqDuMpUujK19cVg+BzxHG6rpvH17H6q
11ffFjzYN5z0jNJJouhsxmW+D+W41TCB9qs1pak9AFdQMjKrX7xLovTg3HTrwiM9X3KDoZaspsdR
VrqKgj7BJbG/Xh1GNBdIzinPXIb/do838yaqTrL4eWXQk2bPqAoM2vboq/iR29N7QgcGBNw8tRwV
Vhd6czc1O/Qo3p6wjiqRZhl2i85KYu7YathyEqnnlq2LQ6mWVRmBBYHWi6GrhMibPYAhq4wboBre
6xvgEKd0hYmzk5qcsvxiIAne4iKcsgpeCQ/EnI5XA3KWo1btulyykEZxF8umcbvNNof7SADyDSiL
u5VQ9dkvlxL4eSyAKUA4h4zL5J/lT715aIlSxL2c8EzKZwb4V4JslR6E2bWu9CGk3SYru2Cun5je
NnEibRARrH5SyXkuc+H+Xe2fXrBB+Vgy1hN13BufsGxTMk8nJwK7Ibio0CULXc0UNvla6GYlvytp
rC6NXI7n+5xFM8NVLgA3P+jIqKFQg4xIRjSIsHRgqEuM4JbocLKTweLQHHwnllf0BzxxaOdQ8iHt
s+pCxyjzcjtZ5FynEsYS623/1iqSwaoZ36mQHlAK4NeiAjV3Zd9LXyE4baytORAPlhaBif+Otsui
aXIDQNokf8bKcN3c8jFaXV5Byllaf1t9A6BM9HBCJJQlWhdMNgTSRYEZPM5UNto8WTECIOyYeL65
5rew2Yzs4oC7Ubr5cI8XpMCy7kUXE0VEJn6MV949omYD1TiygT7XG8i3QeIxKTmilSSAq0IRJMpa
NYnppKHvQQXJtgeSaj/g+WCM5MIYunVBh8ygKDNXU1rkpzqvm0sMETVMpWUkgx1gL5wTgs70Socv
xppE1zo7221mQ82jtv5IF/L8kvJz1zxLZ2/0m0h6wXGu8I8Q/6G+zTsSFpsLtEBtMVcg1SHF70s7
X+JZsUVaG5csqs/udaGs6Kb7DqGLokGNt02by3nj6uiC0r4+z1V50S8Q9/hKzjWSpaKBScT/D4WF
GwLt5Zf0gzl1018ogWM6DNF5//wLkQRsK1XfRVrc2DyvRLZO8aS6U8tr6QDv9RfcCJ1gEK/fRFld
owJ54yda30zHpDlR68x2XIMdaF8yubXUBJmMj171ZNKyLGRKXxxsE1I7mXArX3ZCHzGAgQ9pO48u
yogdIvQTGT0U7wF+S9gWNF+adCua6UimaiD538DoTRGLlxt2NkqfG+6OnSbdB77pQJYZImFFnuBq
JtrEIyW+0oGq2U4mHQPW7CPK0O3iBpuLvyt4GQbublhUuJ5sK5n+/4u0rVJAHmWOg4vgLDCb2yvn
i4fo0VgyU2M5eBVf5mA03PWb/+EtB40NxaPXDbxt2D/kV1NrSVrOKHObPC8ibXCYn+rOTXJeUHHP
/G2Wr/kISp0i5BQK2eMJiEETSvtXius4pa8xr8ejRuCLMwlfeGaf+Wfm5R3ci/YiDk6qvAAZzkCY
GZpbkYyGEYHaJR79HHtWZKdhBzm1R4sEqMjZDIKKsWZnyRGJsFMULSB4NaE2iTGE/Fy3X+WuueZx
vu+IfofZyYZId5mQhV313MWjtDPzrwDz4A5Eb8DZbahBhg+Jdvjzia2v7bWWKDkmv3iKzj2eFVFH
JT0QVVjuOxWjM5KzJo35NyC4dqn5KB5meySmBSVeQ50i5uXazFMe7MOUAcxfiw4TQ72EpinPFsYi
mBXBLs52+XSv/YdQYE67tOyZAFOXQWzdFdtIICw88MuXf4zsfin9Su0Ci2eibXx7Ym8ik1eJKdw3
DbuCWWAkxVGWDcJAuf9bZEdrQBgnHKTQv3PSP6c+h29ZR18YojaEo/4D/cTf8jPbtzIZVq+ApCnN
AFi8IoC4zKIJh9Q4ApeFSHtvicJkligXwbYr1rN2V05qrRgSV52WxErLh3bUds+R5CXu37t2bbMs
n3dODt2FUGcHbB+Q81hNL9dKsw48GPLwxX7D//Yz6OzPcy/r6JWkZAeF3VKaYpoKxQE9qbDYvbAp
DpQSCn58VAnxArUrjnthm6uHhtjtVe9GvFmOxBt1mqcIxSIDtCMp7lDwVHnMzfYPL2XkP4H0RxEj
atRaP38V6v0kmMs/slrKtyjjqdRCQYVja4xinb/8P4kehYhq6TelaW9zhOKun6uFecFlalNwJW2m
EkgssKlrqgT2AgQDZXbr8OH9ojqklWaEe++tnqtubllrLk0vGHrGe40rNcLrSZyb3+EhlqmYE4JP
xK7jEO/JwuQ711ddEszen+ieEPM7TQcGRACJe/BY39EKFuz2pCq3LFtomzjyp7R4W7BSAOFGsAqM
cBhSxEvmLQtPRA8U99yQjnKc7xUSqJgNi1PzffSiuTWPlb3pDnLzk1IU43TG728Bu+H0U70Vc2q5
tcZ6Zh8CC9OnQcGw7o3urB9zCdlTyRNrVWEpL3e3oCPKsroila5bSe/wsEl2CE8xaj3NHn9plEbQ
EiyU0Xpj6prXjw6AOv0kYQMRNRNU4Adv3mAAe/Kjr2fSvFuU9Jzf9jd/CaZU5ZQHzwjikKwpsacb
86r1/+uovKiK4qy5fFZxB5M4d04OF7tD3KW/dBTK8aLiRBtiznLglJXpzE8DkcQ4UcGZPdr7JU6w
eODllf/quOSjM6j9rLcnqQ2NHVKaLGZatL/fuVNmwpcj6OCHMbHLbTvuCyzuRouifcC0OuoBwMQ/
NM7hwOiGm69TDpUPXvWghXpf24zTKIIjeOzfBB032h3OnTCibZ+sJtxu4DBDA0Wj5vhRyOJz5JiE
82AcbTuU5pTc9I+TaoxwgwF7R3OD9boopJ3ijepTrvawQfrBonswcUc8w+0g9kjNtVdoYpzWFHEs
o8Cu/N3b/UXiCXCEcc6UyhAljERHK+BUvT9H62jpsloR8tljD2ailpG7evm2BuEWZEJ8WXyV/Zpd
zBgUHFQDaEL42kdN8YlRdyaCUNb36FlMdqZWRkkACXR73mB1i4R+uYeXyp+BtqiY9VsVUPT2ZubK
mHMAUjrewc0P2J39BBlnT7gDD8D4yBob1XA8vYdXWIO6UA7SW+v1Xf7VNURX53StwvtLaT5OGgq0
GxOD7v3YVrAFSEcGbrozznjQ/Ix4kTfWbjZmi/vj6ZKrv/4KvNA97IXECyv83xLy7hVv4MT1uc0w
x8NU3nv2bW9KvbFV8d8BEcDYk1Dq/39Q0ACD1PEfCzA3xasrnKZE915WmcVslwPSlCfAMqonCxXH
leQmMgfzne6SesAH5I1owTH8a54uR0inGE6ac7gag7SldtVNa8H2py/ZF0+dSN8p35/TS1DbZeZN
TovORIxa1OT1ZTF3CTGY1moAGag0RalsWw6jS1JYCs9gJpCDIKlY5yBo4c01G3koJ1UF7QXpE5zV
mrwGqcvl9cyvw+olW8/yodENXFnnRa0k8eD05f4ZQSazR+XhdKSc/gM8rWg0NFeq9kpg93GG7rPc
0wXjrHsP86bxufTl09/g2JJzPcz8fY/hzf5ETizNxZprfj1d81X6jttvmc9lt92h3D7d+QqrAXjs
A9RCzhvg0Rs57caQ0tH822/RHOWfa0Ds4pPkJ7DrMvBaAMwI+8pptDl2rZ8i51FkRQIp1u+QkRtZ
uswYUnQm9E+Rj6rPDnz4hG+bYHMRdCe5x0wJDnxDd2t89kkT66YpNOlyPIP7zy6fCDHEOLkPQA1Y
knORdaTYERFbxjq9F8PPH4e4B1H1RXghtfA/dRMSskG0njh+BS526B6Sk9/zaHI0OUkvdVG6Yu04
4oCnUirNv5XUWVqHxO08H3QKJ9jI9gbJty3ErtsCE34ngZ+HHN9oJtCH9ASYm2ETmhhcWgVDEDdF
ZbfXnO7pN4EO2PmoEe5COJXK8SwHA0WiW3svvAKjPPLX/pGne9X9OLdd2YZquDEyFoRfeYu4wIrH
PtUkn9eVx39TqKFORwmrLStism/VaJN1EV7zSRBsIQbO8MuGlybIv1hs8drSk2YyHaArMsysrRh2
77qYtaCD9g/Y6Tl4vbDGaTwR2axrlFUKIzZ1473uFxaQhSYeFdH1GtNL0orrB+UX2qFJWqu76vqL
9J0/WKpXJxJ3yKoueu/pEo4Jyq5ent6BSXNgrNXvYba+sLNkSxmeO3UOuN4fJ+1T5d9GCWH3ZmFf
qnjCfjW4jOczArTD6PhgcCs+aaUUD99FOqlXTdl1M5SoSHbdN5w1zj1Vzecsr2wkHQjECWHZvypn
jmgYDiAi2nHyRi/35MhxvTpvTdONGK/MqnMCzhqv67CpL/8UWXHCSxDXVKHNbB8XiKPtQEASCisu
89detTvuQOeh8SRAohezBeLUz16S/SsoDNpIKAsxkx93ev5owaj01Pwry4xS56iewmxKeCt4OuMe
qk2nsEzUghHkWjhiP0PlZsXEDjvnUkj9gfbznzmnXSvfpbmIYbgRuSaCF3et+Hzeg1SjQVj6AHt7
etKncVpTwJkULv0d9LZ2RnkTrtbBhsxbRuqKfj7PrD6nAC3t5yvQv+2FjEH5nczMfaI4xJ/z9IHR
HJBY2fLky9LmkJ8wKic2OCR/IPISw75QO5je5bhUQu3tcNfjFQXM2gu0FqMH4NA7dL6rs7MEaAoU
p+kajzgDEYAdR/xGtjvnXRAc26C/to3H5bOLRWqmq/A4HAwfGLsPK9zD4uu/+kJ/7uY4oEIK5FgN
98of1W8ReIEMAZ/DxFY3ENu8qlK8C8AcPT2woj/SB3ZVv/dkz3I2UT/AZtrkxRdvKJLfPxlG5qA7
XuWUyVW9LX7ZpC2sHN4hBQSrAv/FVy+7aaNZNmjlWImFR6GQkoRyuBvTXEw1+hiCB3VnruEnrsBp
13ZS+IHPVD2uPabNB2LFsdh90SuBp5UJK4l9QGmCyZWPGE1JXhPWkC+7DXPpryszlCye250YEwot
ArdfoMfLS3LFoR/93xl6W5rMEoAD/fwAnyxtwwetakyceaQJxh58O6zFw5X7AhRu2Er1YlG3QCDr
mWkZ/JARLOTmcWeWu7RdiXXw05gabDQ6rkK6/S97HqRswr4NK0DVqgAdpA1gL6pepx4mRKQr3VLg
ADtbw9DO6NhymFcrqUzwK526gOidU9iQN3fSt+gmNO2Jp0b7dIU2Wp0apOL6E/hlo77CyHkFv/mQ
SVATvL0MrAo3sybaNuIufcOHiFEFntlSZ8lEY1q6I2yvPA71n7t3/IEN11NKEIcDRlBYj2yILswP
q2kxIy15eZNHinKpS8oAu6E/IrsbjWG31QYgaXIz/fM6s1BuQeQQ/byPhM8YemVI5n8E5YVes6eq
Z8K+nbiwmRq3EPb8/CoDSALjPZTZiRxwwAY2Ifmb9FOzTPTyhpBU1IyW+5aLHH0zQ7e71KEIkuiB
gZAORMa/6fzZ/zj1/L/Jc0HouEKLUl+BXaMsqb0ENBpl6oMigc4Nkbto1VXN6bYhZS1M6wqODbpk
Ak7YmH7oe8SI7Zn91WMieFYPcuQRFQrE9L20poyz6duFpMR64iPJBsgaCblpvY8MePTq9o8LiMQY
O+HLBYXFKt109vgn/XttbYZudbQX0BaSe3mBAT2lE9LJJ+Q81fne2+BzcE7iZVaZrj73+SM1FRiH
zPA1Owm5L8EuQJcF9nUdjaZAUcYSVpdh7b5DK3zGuR6QZryO9s6FbW3Gr2YAZKuz89oEtLsBNMYX
Stp9Xhgyx7YwMmWTG54iIUpcrA5qg+rczY8xA8H5c/hcPcNr/OGFUpmHfpxv2qMFMdzGz1U5xPrm
YRnmplG7Ucus28zS0XJnUQJnMdfEkpFF5akZfkVxcR1Q6R7G+GEiU2/2YDBrKM+VPEOMWdNK0iUs
j6bZxRUOCIOsf4Vcwd79HEh4Bjb0FOMBEjlwVPv/Bp9VopGnt+85G6ouubiSe7/R+ME17UQ1jLij
Jd1KSTzCfy4eL8U53QRPYAKjwJdDB/V/KmTNWdKLReyAPQpJm+tpSvXH6onJutqu7AvAwXtZ7DNZ
AsWr0qvaRsBd3X/RC+JJzuvggLQ24mYMhEjp1qNUgFK9qlZ6B2CQT4fC6eweYtH9n+9at6gNn4ED
zxD6NSccWFXpMMW8ui/qjdfyG0dHCYZiLjzFU8197Eym99HzsrmiwAy2dOUc1COllmBRoYdWamh3
P8fQ2zfBT01VnVCyB0GqSXpU8vceiUCcX8NseXOJq/t3N36AI44xatMUh7SEkzRH4JMKK69zO+Rq
TUHcuk6ovcrJuYXpc12EPLHtuVPuNz0SNZUAPlGszRel+jlXOpZAe9ZkUwraHQEClUJCGtIL1ynY
RjGZS/Cr/xKGR3VQ/KcROQpWMySsU0r4Ihg4JihhKutiyuN7MtGtVO05wMokyboGXeoQMTRWKIcU
F5Y53KLLDf77gY8lOy5gzHRIMIZupKYHqxY2dikhEjPVPVP6Mxdk3xgct2TPcz0Th10UEHpZWNBi
cafDdimQqOvPe/xhxNnul2jVzo/MSVDpJJbsoFla2oNP9qx/ONvlSXg6MjkbDSYqvDT17VFaHSs6
Qv0e4NkkiULQZkfLWFoVy42jt8f2fa6QYmmhrSkmLcyi0uEaNyThyyEmgVJO9osFYSz7MY8dM8QJ
mU3Pt8yIaUGUJApIbrn8ATV4Auk2CsSmTpngxPqBskBoDUnnDI3e2MHM1j86ixrstZzyXsCq2KGb
UImYEzuyzqhEmPjklYWHXqP4/p7DKyt9bHEI14ALSZO5fTCSn96bmEBIlEBZIbnA+pDCM9J9b8Fl
sU9F1NibVb4yNsiEVIW1S5FLHCFVBddZbrw2DxQqbHBoLcTlbEpMuQxASrro3avdkvWt4XHl/YqD
NIlT3T3cny4y3HPb0NqBGvEm+FfqSuAnaklb6k57soCD6zu0Rs5hG0q973OeBe+Ov7gSBS06k57Z
whUsYXMdpNDcBtSfu0FIsM9PI9fe3OI1oSaJrd0jXLrkYwqtEw9KirwXe1NUHIVtz9EJsIVgTbcs
efnjDqreJknlRAqngP+Qe9lBv2bk62b+TpnCG9hB3EylfGFL+psr5xOyzmf/JCVUhww3TxAB460G
KWe07GXlEPbX6XNMyHKY7vW/DKDNCzE5VY2rBzF5OaENJxLQostOsnBvTX5MJ8N7jRfN367VHKHk
fdUYa1tZqdoz+JjW6HvVO3Q7LVOOwRB4GR1dWUNZuKtGOH46VNrGSHtIJfnDQuvXlBmxy00M/K7x
Qwd3IHKiJp93D6POYqT4GVjI+HzBr06QKcgyih4Z5Vsz5zeAdrqwZirJ7lSCcxThlauew51YVUcN
VwbHypiM3gO479TEbrSrCja1MoFX7vlRZCpW3e5SOOFuW13QLNaE5xwG4yS7yYRa72VZ83Q2xlMd
xRC0Nymb1SZMRpycOPLSx9pyF+LVcjMVibWu690ejM3TGBpTKQTcXl6cwW+RyHZnJPr1x/MQ/SE7
Wasj+fw960OUyzYoMzc66/YOfGt7C2LCF4v8POVz6qz/rN2f3HYfUjT5zTFmOnDiPrG8xoXfiJny
SXcZR6j85dJHiNog/1ZjpQPfXGEjXoZxcCwS5AbI0UwfxbYqyiQRdWywd2TLFrH2KSwcCzjyhDTD
mMRilhrjRa9wFB2WqUc+w0ntCUc2lmwTdUZ+v8Q4byuJ/PS4VGv36Q7v0fbraVr7f+fIZwoMO/jv
GgabhVDdRsuD6a+1lHxTlMHX+u/QZrE5TVHodYQnEtPxm8yxbqvdb473d+nAvYuc1wv9lNtAqjcc
ysxSiS7XPR1PnwXmMcI8UpCCeQOoXXUKnwoH7a0HkoquTxcoE8SGUd8V8jKNrCL/v3izhX9FYgON
DOlJx41zdElOLgHqKNz+1In83eaxiPOiv73378/cURpDAkivJ9CaQBOP8h3a78ZkTUAOQZMgwTno
zaEXDFMg+WkeU4QpDHcbX14ZlisExpAiK5oFgtQyIGqv5K+hpY8JTwPEiwQ4fDszAjK7hlj5v7i3
+QX7049SnZUcokwwcRDw5Fa6lSssLA1tmrKO64I3DYVEtVhaUWkdJ7yqRA5xmZ+9LaErxqNXEY3g
nI3QISEhpUha3mERvjWK6FBE6BN/ZKFXNuQWTIXleBd3vzN9JS+QkUfE3tplNzlJjODWmafRegvL
4Faum+KVGalg9ohh9FRgNcgdIR7bulExyt9qTiSW7oZdKBxQPgPJ3hoejkLPkIMP0OHMACiZVHFj
HRs2bTWA2JMlEkiXfzZkxUUF0AS3zY1o60uT8IozYXSrRyXjjRpboWWCZrVjr2shL9BoEohG5w/w
tr6yZvJObQrCC5ywJmONPOVF4jJk49IoJxeg/AGnldNkdyuzN+HgNO6jo7DN7Vqrs64/J+aoMZIY
79DzUVayaYmlnhS6eaJRpDJrCTf3hDGsSxiKaBwJhCRNE+tjftj12jHzyM1lhe/6zzGslcFjPyKp
11KR2/bZv5BmVoACQLVfkFr1VNB2RKuVBqon3VlZTOjRu0DjjZ4zXylO9lGfTC1QUXmAi0alReJb
Gv6NxmTiyPmBB1fPEb2QTU+kSqRUnK2Y+jWrBAhBd1GFbGBPiZOlDkrs4hLN3IXw7nipd7LJUWJE
YeCkQAZktg0jGXVVBYexEaLicaBhnbNCamh9YVA4HlPlE1xfs04ME4dn3Uuhaw5MxY3ogtasKjul
FPXwFViF0K2zvhlndPoT0qSfCEHAy6rExFPNoQcl3Qxrfx9OFvskSthhkwYEXR/DQ8l9mI5nCdF1
M0/CEmjSeB6DlOVLTUJJtkz/p/X4VRk4sNgmCZT8NKrS9yvexwunwr2HuXD2PRFgAuy6k1k20ubt
58R6RmFv5m9LvUe7rbCgjQAfF9M5f5Ugm5g1U1xMJF3POnRNawrdJSv603jYqddK8Q61af7dzGCm
ucCrYCOqCs0M/uhKs5TLq9KaNWL3CEvutRtWev4EbGKj1CUzmPHlX9aYdopQ7QGvAY/bs8CCQCvY
Axjp+QsjVyZuELSPFzN/kVrSHJGDz3jEpQEiJppOw0k/td6NKo5O2rSn1hwErLMuPGyvXLc5hbSF
DgvsgHdyykTnEOYAD1KLUe57cZUhSZIFYYH/5QzCIYxCDiypF4YA5BgW5zBEsj2mbhHiz8r1ZqbA
DnXnEwBkVoyFVemlS2zockY/BOxne8O/wMWVfMwk9QQzKqjATCUmCN2mW6h6ZNoTj+AO2tI3mxBg
gP4h26igZlRh0XwCrmCC9+Wb2QnxUGTQegiUU99TX5QEIEMgaVL9J7+2LmIxdI04YVzoMd21aPdH
yDjE4SbzpJ+65cbJ+C9CqQun3LH4POkU/ukU33NQUpaAmiisjhcPix3bCHn2TGkn2MTToDeomLdK
C2ZYNNyNikhhRBTy/RPUgt11jJdBq1UYcftQu1SpgjSE5sRzhRQe8xDlB79vgEPzhSjdpat+js3S
pGZbVrSY2MLaidEBMn3jCn84C/CdYTbPLAHCp9nFZnehOsCJo2kRBMblcFMIh7vIq+2CAWR+hcLG
Zyp5esXZeKP3/835zNWFZ+G0G6c4/zwHwUMuZG5UOIwkp07W5kzozae6Lwtvkn4yrMYUskLzXOrw
qVAzMChALIIZN/q1KySP1vd/LfU7wBFp+fp+7QKP9rdt53w+Ud184XkV53cl1dCCUGI+C3JbyNjE
9w2wSk0OvwUfUgsHSTF/OYltoiZT2Zpaax8Hwe8UVgssiDkDW2o5OART4IrVrND2Ql9Ntq8HWUt8
Uc2v1OMOWgmvAIpAzl5RssaP0dTlXBTCwg/Qn0mUaul4GHz0JnxM+/T4i9J3M4kdH3+jn37/Dr7V
+XEZBcjzB6VxuS6E4xNgNqc6CQUqOy6Zsirq/v297ennJmIyEApQJzrcgmNDLITWCuctbvkg524S
4jYHaaY+VPMNS7akLlRDQjQA4IRZWznPonG4ASTwVMh/gsXYqRc269/qQNbQ1yZN3VK7yf7GL0gp
6SCytxctTHhWecTq1Q7T0CbLeNsk2tP3ciDctBj/CJvWjxLJgnPjtv7l1GG4zN/t8ZoSo7Y5UiiP
iy1ZiyCkijyScKtsELl6gMktjeVQhslMCrpaAXwegj2Wjx9Rkln5RRePFXXPbiTss1AgLgofUayK
KgNfnPP4DVv3sgix/vvRHJZWRZdH9iT1N8XcBLuLfFuGoMDCfl2gBgiQ4w+pp2lj3yBdZ5Nx8Mz9
DAzBXQLe/S6DDcfuggQXESBEzLRoRVbgUmvFDqhPst6R4Re4KzYdxuQyXiSZuT47BnTikuUA/1/V
M9kVcrKZjOqM8j6gfFZ4dWQcj86jEHMqx8i1lrLFcb57agp7zBIZltJCEYFmILeEo7EyUS3TVqv4
xyNGfN5xW7/2crPHjxIe+wxaPbG903HCNXdSuVIWHvclPJnKfPB01TikjvfsZliljVzO/+YcTuUc
dd5eqjThdtWgCFDMYJNJUXn+ZpIoL1f3EuasAXsFbI2B2tjA8taN9zHjThJB1u3/VYxOvrfT48R/
kGTi7KGsq6doKDF9aGLeRV9/2spwaheHXZQhizIqhcglsRoeatemk+flN7r0kotVQP5UkthARBeK
jDgfXZb2wx7YLE/UPhUI7c12uIDsA/NCNqPXi8Rd5XHwb02JO7WN53PltezdAHLEoy3qZdrFYEXN
HEc4/EJBxITqX+BhQ4CZtYZCrP3mYIOD6syj7kuZEGPOV61MLKZePcHNuErqV/vALUowUQ9vKd1c
THT4l+wQCKAeBQELKYi3BKfX1fffo8wSg9BbwrrJe8nWpzpTTHS6hY7ljDnHqv0QQd65I7+lhAaj
/kW1cJtmhqyebpT97qINshgVN5HUBcNz3rakSKCu52PRuBQoadrEImBUJUtikAGrFcMS6a5ulwKT
xhVuEXet2EvPIftwuFe1q9jLZ+pZ6TMcrLMoCi51b2gJPYL3A9hQWJk+y7/t38CDOU9Ir37Yf7m1
Q194SmBC6qRAScPsr4mg/U+QHqff4KQgFVIjSI4xl/FhINOX6zIQemov+dDgLE5dmvNAkSMf+smd
VV66xfsTKnpJypzErn+s/n6zakH703S/ufEYwXQIhf3P/NNxOSA0nP6ZapXA47EvY4MMMegUYHt0
TtLNdMrmA1NYlFoGz/TF2utsVYSPaYEIdhf6i2W+IKkHz/KDDIofVg77/DxUUoE7wZ7c/peTVA4f
jVpKaJ0bUZ/gHiYT6lXaSBC/EqzyjUFRz8UWyutmD25H0o9PUog+Trho7iD3crJvq2cZf9W8lG06
5063pqwQiRR7RG3L+iQpFqJpUUxc7TLbJ/rZJY8cfepO8g9KEfyNRnPzSpo0sDptqz85qcKO80+5
rchjsFrP+kVJ3sJluYLEaXUe+/f1XvBfEvTnimGP2Nz2+00NRVklDrHGyQDivbOdFEtivTFTXb2T
k/b1sKd0RZAMfpNboGbAGP/wIAw7hU0bJ0ARGn3EZ+7d+OoPQAa+PiqK64HECLAGFqKuZy/nMl6W
5Ka6slnCC8/SubAXToMCoZI2UlOUnrNO9dvCn0vUpushk/VhkKGeCn4rTxhag2X4NBp9ishJPZUV
hgtFnG6P4XSuVSoQLhdi+BpowqFAWAio2uP5QM+PKFHTcYTgWdXTkY7RyqhaaJgYTW1qUWIBspze
5PxPbg7VAc74hy7KbDP5LtQPe5qE8ehgCD1R6XgGwdvQbbkZ5tjmTarWY+9evghE0RwvHBKlX5GS
8Fq0rzy3+WkLcXBedu6SRsPKQdwscJPlVCU/QXkrvsLU0xhx1h/d6PfGwSEPtQOmEXZ/uCzgqiil
rOmURnnffBKOeWIk96GuKWIt6166A81SJF4B2PQ6HUlLyVKgVKEWxkOi02orIaUWaZfc9OlxtVuE
XOVrhtPZTIF4jRvnQ7vk1hqEbaIcnp3sqw6lz10I8CIxjOY7HuUStstVOx5+csGQzK+E5S/BPnq8
Ej2YJ9ZooXwdDlv0RI1c5CoODhu0HPRzkwUh7Glmm/C3msiebVnxZv4pZrsFI82o9CJ6NL2WTUVh
9XOpQXClrjZsGRDQmG+pnAu6w9ECrqbitDasqZu62fcFmceha9HQZi5ZZCDyk819Up99o7jq/GVf
OpANyVuDceblCIh1Rjyh0hp5DPJTocpmZjMJzWZFQGyuVU+q1EC9KV35X8HdStMpgHboD6qrVtqR
k/CljlVC3D/JhFAbObOfn7o5MJKFS1m4MgVmkCdkpPXPXY4ZDNFHq3V3YPyW47ZSOaNluZiXfZD/
KQIwbHTb/A28Lq+HLumvafCbSHxqzPYgSLvnpepa1fBcrJWK0CllKrIFCTpsqLJIwxkT/nJp3k++
BcV/iqpKbzT4DVaDCgXuAVjEMKtL45RvAgAON26ZgBAwmMKcjMqieuDtWH83wFi1akmYI4UDvJ6v
oIhLHWQ9BX9khhr02wzcau5U3AdDxcIuS4gofQwSyur//5sS5ab/g15cymeUD6tJSG/YJZAnHGOR
DgXdq4xDM/PF2x5RUPmeWFUEkm6A2ke7oNHKqt31LIcVUcW00veNnm6uCPk6AxRfYdKq2Tws4Atj
f2FgQ3PHsUlXuOFZGWv/5qBC4FOmyjKk+lHURdaVbyPXEVzONAwGssO0ObGaxtbcnftYtwOhFcJt
/bpXZQazqt8JyO3SBtsUSY62Zxv8HNYltH7h8K5C/plojfgcHrAohuoBobuwqbU+e7HWVmOKscTA
O1M/mduKKpVRAGsqw7GsxFw1huyAaQ/V8IdnEnHX1CST4WsRWiQea6NL1YjYl/dMmAilwsLVC5NA
tGOZ766Fs0xevrkD2Ke4WdIkan4P/ycjxQyuLDl5MwLXudU/f45ak+wAZ7Mqni2C0CDoW2nVZqnQ
Lx67a4lYErBJ1YCDwdhgXGq8j/UPkcI7en/lWDlcZxgx63g1JkWyEXSamc5SrMVtjyTUa3vTpMHn
u8/1lkS34hWMIWqr54ox6LCnow9feqfLrYQ8dDZ0my/8mcoKjBV38I9SWGnKVtvWleZqrh8sjr7I
1yElVxpyvsVUKTO9sVd3860oD/gM8tFin6JnTzDe98C4lUbnme2O4AZ1dZ3megHL7+5S3UFixssI
LaxTIaeuQ6BeYanjbIpdtW1poOF8wtmOo4bZgTvKCUkACZjRRtepLSFpROa4bESBaAiUdWWrUsPF
51KOdueJRB1LzjOKTUhpDzSxHy3AEgjvj4stskC52YoU5uhpxBN2J0q4FWOUpxBnN4uzvSSneCEu
iz+wUVcqi4qTng1I6hrfGoUYg/ic0ZUiv2iu8BDadxFhliFoPfRlfaq27ZfAqP2qhNB45xltW4Ix
u83elwuRNfOT694nEySU7+awxI6Bw6fEZSAKDhLgxGFIEhm5JxsIM0oN4ksqPzzq3ZOxQqH0CFNX
l+96ZWo1Yv5UJqPmbY/9gLJZPxmoOWtE8HhEp5ydQ/WEgbZ8CvCmEXqpHhE+uwOLbhCNVETuY03A
1VBfGZgY90Q5SS9i+CIVHQNC6DVQ+7utqjk0UQ44aiwn7sVZ6Ea594AZUtDc8Z1vhgYIswz+T/Gy
nMtXs10u7sRqQHWsJViR64UI8nDunSmS4E9v7EXw/ZD6bsFacfo/yPQNcsOK7x8t5l5NGWgRqWXc
Myrx3f6leUQ8xMwB2meWPv6RwSH5l58JHoQk5AwvyD2vO1PwOA2QsltOXC00wUxi9hFIecJypgQr
1jpmQE7WKkv29i38MDpxNl9OhjotgQZpcygiFyE8pOUCIF+LGYz6IP9S2jV2PCcNuilxI8XtTw5l
omyRmy96o/RParxdFKIKV21mpYGcmbuVibhzVpfT7Nazpo5dS/C9b6li+fEGknX6Or1jMn1nV00r
6r4Q1Xvq5kTlDaWWdsjw7uKMdauatkNBnmDsC2V2PO2P5zM1b3smhsBs0OJKfep3c9GPGfqiZKbF
IyPzmY9lNNPKbftUP3h6QoSw9T/CfkGu9650RD+uEvpqxoX+PFMBfUl87xTmFpIG0T8kc6sMcmYQ
D8xF+nSuaCD+pMWYhh6xsnhi2/+eQBWduZhXEYLnN7JbWL+0KA7HSx5ZmFMhLfd+/hfPp972oXLW
P7cxg/fIe2IG8ciPRWoUADWjo47ha2l9wtVJzMf3Cu3AWGA0wBFW8uwPsW6VmQ4vP4+go/lkRUuK
59AbihHNr3ei3kGfMUL+OD/v5tXlSiMLrLSshUVutlEtZyie7pL7nNrZI+9guZdghijg5YgpunZf
XEdeuEDjAi5TyubPBdDNLX6JBAOo8TmRijui9hWQYCxevl6yGKIU16ZfAx1TVHDxGdpHUomG0OJx
KZaDUOAp8uv/jCoHFUIiyd1amq3xJDCRZHpejk24okRaqbrKxMfvU2as/UV6gXkoNABUnzqt4w45
dHSVEccopQq864T0YdlCHhBJQOEhQanN5MPGJ1QixBOdbIM7G912Am0MAVM3ycuuuoUk6XPRWXwz
s1KNo+Np0ltmC6fRqLPSD1EEIGlI7LdkeIA8h4PB6IcRLz6+tNF6pnN1B5UhE1+eoIGcmZIKUutE
GrHNZUDHVJU9Uid4ms0HehcVC/hf7MGYzI4oJ4YSn4QnFkx8BrkOUINYfS3Zea7tz3/0TegDIV2H
PSDIBxHSbPXtFfb+Z9VBjfmvszPT+SSYXhX0khDjsNyKxWWIiyOaOwt6oEWwyUSyaRkUPaE8R/kp
r+Xd+H/6HzbeomsxCuCRVNcVr1S+T/AM4RYblwUVEZwweBie3eUV847e0EujKMq/HQqCVYdOcrUO
XkVZZvHrCDX8oGKpizt8j8xkZowRIRm3xx1IrKudKFBFq4nNZsGjuCqCGP0YPueUPebtwCwzYNgT
fhTWLYBR3XroymZmJCBVCDMf4NkuODcUiMCUEo+jHZraPwsmLL5vDIPFgPv4PHApxpEjAcpvFSSc
VqhXvSgJDecUNPznIPakzi04ODPTbCTrreu2VA+QccHPPxSKydOpFQWISKEwYz9wbkXcPxt7l2O5
vNE/2+J3yVKC7TCsuCXU/cts+ZKHkQDkOJ6lqlyIlol22OnNFlZM8susqNNukaUDlR1DFLUQebDR
g5hOwT9G2phQpNAvOl2o0lj2Q0LB13OimeX/RzniDMntUrG05wUnDkvYhA+KttoDZeTuCCknXIar
HJro8LT4Zbg6/cv1R9aECzVMP5VQ2QhccR/Zz+wiB72+21fVwLFUe9CcgQS/16gsK8C16FMP2h4L
m4hiRsLKA7Z12a+FnOTBOkmPVoNBNb0D0dfgUeGzeyct/wvsUcAXSGp73pXlXrAjx0iN3e5/6GBX
STsBg9dL7cwOQUap2mvdQm7TpLRz8CkdsSSoZcMwQK1gC+TZQr8JQHnx3HI42S+oGrNNoRXE6k5l
7TW3Lc1lVkhupjnUoNPXho8M4+gzs5DGaDrPKJQ6ITYdtv3oCJEbRW8rBnylqTieV7K8NMaqyEJo
08rXZ2cskBcyjqqEab1/FXE5+FhlxTaB9RNH95kVhbX6rgwjlJngk7S45ORpX2cfzLqfMIwKeVfs
fvjoN9Vjc/0Q05IIWz+vV4GP83Z0xsMSzMVOUsO0R6uIL0pWiVZkmeWJH0rko4xwfKWWhTpitOtB
69Z7AxHohIAMgqFfPIzqN9JaIuNkzCCo5Xd1NN5DDse4KgSVi+0HEakzFOMfN5W4B4TvVwKHcRpP
fsHjIEx0E3NG++IJNIlEtsOJZ9ER9XkZpN4Q24kRF/uko8+mDO1M/FEknYhRmMJtPybcIWkT6b3h
Eq6wKPOEyOqVYOHUt5e2U+WuxFfCJmFsFHZXSmgpn4l2PtQ94YAhYTOoR8CGCRpstnlgZJ3SnGWc
jgo9ocesHxnTPB6oHXTKotyexMUxXKMq8yrWXil6BUjKHLb8Euh+d9xvO9ekYLIfxaq6SVJPWWqg
DIMtPcZmpfUG3ybe7SMdP4m+C88i7YFpPxQxYoBm0Rk9OPgwzAfK99q5raWJOeg1csxcP6lvg72J
1Vxli9NX7gGLvaPuDpOE62rMC1arr2TTuNDcfurvAHCcX4jchZRFTaRSU+dbDSOGHNEzlyJneXcS
qfS+sf0hRAOcIg+1tk25mYXLSymu+Bj3k1abVi/+uioPscbc8/nAhwqY90zLbwYZj1JXmgRLS8oK
De5Pfg9tm1nupk4gkBXgjfIPmNHA8doW4BnfVqEiA8AS7x6MRs4GHYMKfv5peOnVHxeNor7jtbuz
qK2ucg+KpX58og8WCNuMlrN5HnDo7CrbLpVEE0ek5Gm3Ad4vV9lHyz8mNLx0DrmHSQ5TJaSbDyjT
kDHYuQ+Yj8GoD2vqEozUPZJyKgzKkl+dVgUdDu5jSWMdHJvT0WVIWObnBzQKdTKTaxMIe7Nc+Ojr
U9IEepjTZ1P0ADHyDPP9CC6wXfWVsgYucUIc3BRY0xFa+5JoXMmjm1645XhaepLYsmVaFbFNYVTz
AsGH+YFjQSFzZ+0Slg7Cp5zIZ6Rqw/WL2iSbI4ZHqkQRVaZZsAh1pW4Wze2qbjnFOqWTu77A/Syp
iZK1qMpzhXs57y6NdDpl5NsAYbtIVK04rdK6DgDCfhpZh+3oSfilYJv865LSjBSWaE8b5OzMX8gm
1cNV4H8+GBlwRzdq310HuivtjruDr8yY0vSexsvS9+GiQYUqkv29BulUEV1vORF2AeuNzjLPXgNt
rcaTFZPRmwmRhjM6DtAtUQ4bo8lsB1iTI4RJ6eZ48h6RzjdG7WmK+les5EFyjc1gK1+AqKvOvbh1
CoW5oJW16fbUphMtDSWcRDdnV/QjfIHEx32LoygPaieI6YV52Jgyo9E7HVneotflNQBao/N5Tdab
547irgT63Mjaqb/0UEnFcr78MdBROozSd+y3ZjyldTT9dY2YS6Q5tK6ISVNZTD317Z0BIoVlossf
EiSPtEUrx6wDrABpfNCkRCWFYQit1t92Er1vwfHsSXg0sGAL+snBZPwjsgDqs95DNDgG9GsFry7v
NPgXV41BEWzRubCFW6XEmKMULjgvzO5ZsN10p68JvI0rb6Dcy31EPWo2FLqS3I8onceFrTyByj32
6P3jTEhO/pjPIhwybqmVobbkpm1VRnKcFegaUSEdowBqjwkLPTeCHBhhLZJ+9Ec8ofjptECTX3D0
aqFkOM/OR/doCcs972qUq1c78hXQUVChn9rBu958LjCG0/DXK7p8kd27yLRfAqH8eUZFhJk2qGEH
8h9ya6G89AL0AuVdUfFlJDxxUb4wT5MPeZPOVUCL4nQuH7Jz6ZR5gvapFWb76/um6eE8N0nXZsR5
p1ifWLIu5s6JGAvuNuDe0XdtZUyrMof+A3QUWI97duGDQs5qgK/aVgvuuRzx9iooa6WLPqAH8omS
iXssgarOrzpz5c8oAyBcBvaPXUBy8UJKF2GOUcV5J0cDuOdaQJC1a1yBIVvHRmqz0cVhadSXOofc
O7VSEzBXICBMPHTSl9ElA2o1WmAfKljuke5+J0lGYc0jqdVd5oIV3K93rSHcv6s5Q0Mis5FkJaYZ
4O9RyLb/N8d7xMtjAA+C+QZ2StkH44M0Q8wVNatypJ0561akOakUrirMMfbfZOb/uL02w6FCYsoy
KIlAtZlhlUJG5WSp5UItw2aJowpsdXbDdblaAmhuYUIcEAKgg1YjhCgAO6tPVYlV9YsYI5FDJT6o
+m3eJKj6fzkmuIXRe9gZXVGslV7Lo9YPi2wRrvcc46XIaQqDVI/kaOcYzYbnPrIkXcPvwECHjh24
3blQl3o+4Qy6fiQJfOGM8hLxvGvEqCGOw7RKqS/tpGkr3FZ3NN6p54iaq+bZVBW1jZG9MzgQY6hM
kJrAkN4VxBCZCzM3V5uRpRAgb5dJFqwWWfsruiSOWiVeZwtZMRnnSCkJBFmHqvAsG124n9iZ8RsT
1bwIvhoMhvLNsUjqmVYLASMgkGLPGJ6M6Dxm8bGx+TvEZtnGgJVHrMAAhXIVSxyoBy4SfycVv5PG
8Ds5SBdO7Qc9ytld8tVtTKlX2jh0A0S178iBvf15zCCVrfTcaVORM4z1PsyxiSPHFdeNUEG8tc/L
9uO9vFGcl99dwKpbeLE3rrcLdYE0WybdIIFUJvUi04uut7c3y0BQ4XCnHDRUJlwyqGLrcSFNh0ti
Rd1+bRSpz+gjzd3MJh4s1quiXas0I172cZU6Ib3W7AajTjRhph7CRfwNBeXPVwPwhyEUCTexbiz9
Rjm8UrIstmq8maxxDAfFa1nMnWaj4Gbw4btOyidbtdCGbGaajt5sFyKp8Vkdo+ZKtcgW4BOBLHbp
VcFG8brQgwYiM+yzhIt53nRJCktjxZVFgMY+gGJOdfHcip80jX9/zPHMGyv2ja/h52/N7MBKVtB9
yHm4sCN2DrRH71MhPjYNFl0OArOrBQTAl+jjhFRq3uJ5kaOtEs0CnjdkXfBLwXrJXqDe29WrsEbP
3UHYO1CDoQmo9E1tpNyb10M/0trrc6Qw1TNzlnu5zJHppu5mtXf0vKZKYDa+pStEjhcTeqOUMrIe
WQJqXqcEpTiI/yapwtQCwHf4WSmZ23nl9sSd5umuQY9/x2XUNOcuXqCzdeanq8x3YnjZqY+nkovF
kdXnjfrE6Q4XnbiSl101LWx/9KSnNxV75OjRosbYIUzKOb+a0ud+3kANwGxR4NfMb1/xFrUufKEb
pzx2GojKpR+fb6I8+eR8U7LLc1BaxKS5Mb3MpUdPBGE609v/Xedb16QxXkw46Sne1h0gmZdSc0Ag
N2LgXReskQIiJ5ZeK5IkKwhjpnuLEgeCa/dCgoCZyp7rMuwOFWwpE3MO3UZaplNwXSCLbQlSZ8pV
XQjJ/Nbkrxy84FYqgENq9w6Fy/Xb9YIKbMX+t/JJxDb8DQ4M8GG3LQqaIJufMKW0hLz0NvKw72qh
RRUkZ8O0+Sfox2bS4lfHzJV+z5GfrIojC63tjq/m8ZaOk9a8iP1pxWvIL1DLgB/b7Gc4J6Hbq+8F
3s7IdZ1Ym+XqLHmKhyXnsgwvqBrjDuVxNKFJ+EwdJiL5fuwW04eba/ZCtAdjuIuhu7kOhvxGKSja
eUknpAAr1Zs6LnJcE917OgDqPKLTO3JqNFNKEjo06nkaKchhpF1SC7PdPXZRTCSXuLDpZRQfFxb2
zieUQHXwJ42qFnGRlgkmTaJVDV9DIgQcrcIKzXruOsHU6kxU/rGX3QWYYjXyViGTaYoAIgCUiP8i
nCAPvt09nrDcVf4ypC/qsQ0ubATElccNN4WKfKS7ZZ6vHv77Ew3BwdSuiu5eF93Owsz7Me4E4vXK
8xkxsVpujjda8Ra8s1oMsMM/AENVyKK8gZixp4qhmmPmVPnewyG64afEWdBLZvg8mMpwQScUZ5Yr
knVx2BPBgSiFeLmA0FKIQWvDWAGgCi6sOUqc46Hrvz4FeEH2i3DJzSqOmRDXOl0c3LtxPM7gNOPr
8rbIhWmINhgONifejA1RudYAdcta+8toe0f0ziP41XyQXOHOdHKQSXXGy1d3r7SQ1rIsieAIYDLs
iSTaYFc6mtg1Z+mBkU0EetVIeUwz17uPYbp9hdur57tv+6UTTZ9n7q06mA9kfPoIB+63vNJr/5dJ
/8T+NQ6KpG+MGOrglGzDnMgIjmTJgk78PpD18NFP4YaNQxdXPKEwIh4/Kq6NIG8S5zTAOrWPy+F4
oz8iTw26ECyrwpnANbJBUY3BhOn6KfgylHuliUBoEH7irVsMegyjx7WWNcl0LvENSePehR+yscN7
/OYPebr/87Dq9GmSNW/YbEuMG5JbePQXzCynGq+klGCsbSn0GWwv9cVxABRE8BcsFwIv+1yIGkU6
zsReV6KZDz31eHLLiHtc0dITXytMIMmSLF4MrazOGD9jkBxRUDx7fr0tVEu1DBNRhpEX14zFXXtB
wgDrwhJQg/xmTVBGBWSyzKM66ldQ3DAk9MYDPYzP/YqCYpPFExVIYY8yZpFzQ0CEXQrHfPJi2i0z
JufaRU+tS1sUFinM/PqsFEvAMnTfbkaf3VJwd8BUlKdg7zJ0JDvWWE4Ff6KaLmdeG+5e7HsOpjBD
9a00QUvv+AyHyLdi25/GHLa7R8+GLkpf9vU5W2kRAwPprcFTA/uoh07rCvSWttjxliy+gWOKS0gc
g0AEadkdW7DKZPHZFPepLraDYbjU+OOEGvGR/cCdOx1pkmgR5+B1SPa+yGtnIG0xFes9/7xzOCtM
AohCnuoWDGOY429S6/xtqKaLVDLh5YIXieLyhE3y/hP8CQODpTSpxH8ZAkhsna3r8xSVa7m0Ojqg
d4RA/R1H8xAZ43qVuYTcIfygkXhZ4wCIw5hmNmG5hZHkQircel5DMvtMrfDbL0twxs1ednKQtgOY
rJOcGCXNn40frOPLDb6RhrEyDjGGnnN8pyspE/m3htwrF/pVyXTZ1Fe1+ySNPRs6GKfmYXRFppig
BdIVr2pl8lSxO78Og9Xy7/6KEjYrsDqst4LD33NpqTUsLYCbmCm6ZhSfKc+lwOOdtcnv4O2RETrC
A36VfRMz4pYwsTe4deHUiByC9W8F/1v6FGCciG7TaAFl7jcX4FD4AXM154C0TGSmg8JliGakf4an
5c8kKdZ+wPpyrMzOtIyknY1H8Nt2mtXcsoP3FQCn58A86uvt4YwKFKLVPmW1aLML9PPTj63sTs1y
+864gNv/hHMmAHt9WoGuMGznwMSPW+GpE5CeAJxTZHwkOQK9bCqbUv94bnQPZIzqQq2sa+KkEcu+
T5vF2IuNOgsd89RskvqMbbUf8iBDkBRqfb9zyJzF9w2FQz4RJQ5+23N+46Ce9VvJt2XaINNdU5aP
o4fQsj2EXNvhkpF+naWqIJzOCcjEQmmuckofFe9Q2dDv+Yt5JS8cdggN2U0OABffaKvvgHz5FN39
wAKcyfne/SFGEEiFMqtW1elDrV6F1w16Z9KfNkKCkJb6H9JHeQLKUvf7bFw+CuPSvHX0kcbcaVH3
WC1nw8ojFg0y6vCZ/eVoMHkf1nq0m1z/TVufq5DYy3GGCPcCc+QQ3S3Qi7fBE/bZI/Uy6K+izVwQ
n3VtpI9rBWvpmjaFw/MPkDDh/qS7Xz5veDqquxEq2qEtFP9tq79MK228awDCqXwOmq5tUDNKY80e
XcWgYnvn8w5cGtq2AZBpLWH/Ym1QdYegs3pN/D81mlY27Ka2wdEtqZ6jDQ+XO9BEFTCFJ0JoEcVD
5IuVKTE8G01BAk4ail8HUDfytESS0kijoEGxpg4lWlnqi8TrBUDcUusoJJTZ8pCxFyGnEA+Fxj0+
kjj7Z50dLQcxlvdH3quyjVAyQD5FYdmDGqYVTHqKjmTSZOPuxQ8017lS3BwGgLK+NbseUlIl+03P
kwGj19qsIv2Xindl52U2kgq1h65JfcCc8jCS8aBbtNlO/mOzVt32KWnTXWRASUWgfWKURed2Pj9Z
9nEeVh2VIE8vvy65JStK5GvDIiaA/3Gvyk8WjLgHnpNU5XqteAiE2NUXGooWMdXzvzPmgR1tCJL9
+GcA6mKK7kp49+asvM5Fw4m2ggJf7Gl4qzyt9HKucNb8OL92l74zAOq+KTDIp0vOxT4Lc3rGpgtV
hBdMvHXw7gGrcb5my3kaK/mLFwUzgctSLzVwa8eLYBYiFMJnjHX3rSn0LAYFBZQTWwa9Hy1HF3YW
Y474Fs6fPBDVYzvoaGvLvlbODvtnzmfYUa+Bt5y7LyfxwLEKst765QdP81NFffvyhm6xFZXJa73W
qZNCvXm6cfpiCfoyQ3Xb/A++OiT89DUtyR4IYRht04yyJKdowAazqBUIX9mL/Rw3+gBrSfMSH9SK
SufhDUHUy5kmg3/gk30EAlEcNCA0rLIu0ySt62h0s17tVz10PgqQpFLkxslSY5cAS6DR61d/4Vlm
TO8NIFUB8a2rcrk+ahmnUP6iIih2jUe0oVejgbV0LNokl3QSZ1DYSuOO1rFOc80ROg9j8sOydAl9
S3QnrfZ21wiQmNfQqmScjAEjB7e89JHrAn/ryH0jt3+47/Mx7R+ekhd4snqU/gWhLpsEP8OUGxny
0+m3rOWkUSK2M7l5JzXY0wnndgqW1a2cPipTJ+sweP4kpEOxWe9PwwN+Camzpb+44jOeKNA+KtLk
mVtDyC9PtVi+ttVWt5i4XOMxf720NuVNbLEegSwQXNLpVB3PI3CiOguQHXXAW+ayjXMkE1f2aY49
8uL6SLzuuhshQngOTLuUIRyiN18EsskIIe0hcnNWYJ1U2IGWfL7tNNlAYbOJMN+2u9HveoSMZLGh
FNs4iDeP8dytF+N2VSVPp+beHnSC4LAZYJREhYPyNBHmV5uGSmR8yyhaC8mqj3ySJ4Fnf1JMMWJM
WRIgz8yprdhUkWABHm1FWlKRjFaKXmiZjwSjqKjUslDO5dlJK5ar2hDHI32dESU3P1u9eEAQoBuX
0yidnzLy2XHaT2AKbB287NKbrqnWvXVWp4609zRaIYB4vWLKoNkAirKPcENG1kRnr6nGmGMGBuif
o3iwfq7HREFjvePBLBfvSULhkM6WnJlIC9EOmOxdEVFfFK0HJEMQ+DBSJ+/2+aVVBRMM7uCOqvf4
607a5p3miG4at/KjmLh9WQICWlFFbMv5qItOV6aBn43kvL9D0x/XGa7npH84Jjw2y33ZR+G+vS4K
I2Hy97ORymG+5wRi8gVaQWMmx6vZJ2gy7oEFERmFTsb3EAsc+HsgHprDnd8PrqpPNS80970Rwx0X
M3hv1oAEKUb/v8JS18YZ+rWOUPTbYKRtojdFr1nimnzjELO2cQy14XVMWKi7wV6J3+wkwFbtjsLd
FMHv2lkmDuwozNg2CiZ4QPS2Z+uuT9j2VmRhkHjUw3tyRQpRB1FLcEhQlN862YlRqi+HW4Ej4QD7
p2FXqtEHVo1byDnI3jDGeFcSjwDSnZ1CfhGa3PmWEqQMPB8lvP2c5sBK+t67imNQ0RRAY25416sh
yauNv+XoMJblBu+aa2ym448rR529vCahgz6o8JMGKSgX1B+MG0PfGjJ3nnFlvdGRHNOcdY8DI2Qb
18gogtNcCS2zwGtnkfTWsQCSxlXHUpmqy/jP5JGIEbbH43CwT58Iwjr8hw2GDGsveJ90IC48pNT3
W6fv4UEIydr9RkSFWDEad7qvyuqudk+dzOWZiyWu9FsqTRl0ymlywg0MN7je4iYqxgazZ/zc8HJ+
vBXm/dyq+e+vtf95sZKaifBKtJoVMz4WYt9uZRisNg0TJuMHhJoKlHbT8why6MCHk0fAQR5EkteY
+Vd91QTrSiBo+X+XtKk1yvtTBqZXSJM4WMUJMHXztu8ZGXz6Tk8LwZaMjpq+YGz+KMs46bBKKKRP
PUz4tIuX6K/Y5QT2c2JcHaV0PGpyuJ8P0vdYj1WSe6csmFZL2jAIoRoJK3NwwWr2m9VWtWy8HNJB
LvkmGz0LY01dw6WVAE/+aGuL6ZWThjw2cnXmWw44R8NpeJr+I6WYzp8ndPKTp/Lu+ppJUGTfDDAC
E9KEHGJGzIB7UM1gIo5jLhTsSEclnCrlN/90e987cHPQJ+7ZXeeO/jdmPdPrRGApsY1H4l+teDWU
Ffe3blqvOE751ti9XUZzGjIpghHQAFM2+LvSc5fxEJaCMohm0v/i36bDUCFppMi/SbKPma0eH1JS
+ucz/Oq3ToE5+dMjq6ud0LGpEiI87bA1lOLmTX00JCH0gSxk1ngmpbQtRkvvr7YnwYc5fIioPp5W
D4YZX8AUG+lQVu3MyABg82+H4xCzPqzNTG6gwmOVBK4gYT6mkLjKCyOewitTfIidgZy7CEvCx0zh
cq4odGPwhGFuy4NAkUMkaxToVhxYxPS/el0gOdR+o9euJYPFe2cawgZ77p3fhbt2JAEnS4pLsS1o
faRa2kD7pAjwQ6uuB7GdP1wAe2BdvYa+1nz5aowdPdto2VB6S/KuV/YcMvf/5FyZrY25YTiQkA90
g6eJu6kkd252mWEmpc6d0zoiVfi/QjraIdOQNDSOtJWmH3i/iY9xazn51UCdwywpZcJhgZyeJIlM
XbqxwkZlRiJm8lgQOwFqI6vdhLSnn37LnoyxucozB4TCYcNQvP4uw1n4vwjzh8//qjXKNKaC2XTm
NYxK+XHEHMICDYCv/6caj/Nthh0gNZoaFpZjthq3zNKs73zUtL+6TyDOaSuRNKgg8Pb8sP/KF7c+
9BAklrIxH/ij1M7AFl4784WL5d/Cw/pEAnhDq9jcbC4YJy905eQ9+Q+m5hEPgUxi1Z/R6S3BX/Mh
yoneeSf67Bg/PzJZvFYzlAP9jOtHPvvZv6YFVD7ljx2DTDc/bEz4XXhNj0MBCmw+xO7v1ScrZbdG
fBE3YYXOwWV3wPTGIaSK10HMcFBcSpTK/RrELC0mcnHs5ZyemGozepzDBBRzl9TSjRH3z90WvRLS
g1KxsGpSv5RN/DPLeJt5U5QH06WS/ySi+Y2mttEJiQgx8QyQN55YnwwSudT4vIyoEPkvS7xTLWE4
EojdQddgoURz4FZ45+bvUJYQ7QRboYdbHmFCGlBjlfrmuniuxUCTJ7jcuNXkh/9ijTYmx9YHGRwF
AEVtCzeFa5uaNGRtaaPFlK0n6AQhRcS2FcchgET6HSl0mloyWhYlXETQROkyg4VNfasYrWB4DFD1
25B9qQ/yhg026/aqwmrz9w2IZBVSkuKH8awFYk7efTL0DJhk1R37RavJapL/pcHZbs2Dn9hqP/e0
xYV1JdeN9aHaPaKbJcj6LqTHuFG1ix4LIYGu8QorugVNopDD9USyd4Ll50l1lf4owAV8/1lSRQgK
r9YvcM3ZWcqX5I053V8mRGp+jHJt/q0HAWLrl0R/2qj6dC8hWX3xuJVLrPDLzkRmt5G1K6TC2uD1
NU+lRgdW07QuBTw/dQ/pT7eAlWJMEfvFuqeMYkaXplAFSw4tga1FTYQp4xWmeEFfDoMkBEv26URa
saKeE9VlH5DYNg9vRbymP3ScEVYCBFRy3Z5JN/Mdv0MATAVimuv6uEHfXbZVD29ZsQ1aBQKR2ZoU
EY2F9oJCSSpsfcl73cnizpJj4pupTiAUooLH07KMONCZWvOYUGOuF8MX3teiFcNK0ItchIP2eKVD
SkFgIwQfrV8OlDyzVKucTFDYoiq7glahoRHEosTTg1/XLHONTmYILYVcMKvWArMPZK+kuyA6Cq3i
jGIrBikFY5vvrlU42zxYTc3GQF5il5g3KeoiqCQAXnXFI4MYpzme9ghGyLIZP5FWzhByLxr4g0IX
WipOoJFcVMdmec+18LUldNZIQ/BtHwM953BkOsTUd8t9QjtmgmKgviem4kjDaA7gOTIxtjnrPjI3
GK2EmRq0t7ifDsgQSDltitm/EtyzjNpksGoMS6TPwOrs2JMWkUj478Gudn6iCwM8nogJYqzLG7Di
+Fpl6Yp8HJ8yJyLog/yaMTgU9jd5g4PLrOnW5R6thpCnNa5VdW8zKU8XGPOMXgFA3QQ49eTxTNMI
bXA+dDQma8qsrQnfp/Gw2p0skbAZJe0eizCKY8KnlXf05EzmW7x1kPtxMnzs7rYp9Z8bz5G1eq1h
lsTmg4jPfh47PD6UxfNkwMYYFWiRvkYW74K6+MlOPujHYu4gZFsZrjj3sBOLAa+fIKLQh74fwEnW
M/hFZHeQdO/gv97rF7f9C4obm3k57ISZ9FLX0I3KWuKrXyEyWfX0158INbl2Mmou5qKgEvNDpCKt
/RIxXCIcdTsBIwn81GhiyFV+DsvReH/WSjlEJnZWauFq1jme4rJchZGBlUfT2TqiB2y4KSqOpwe8
F7twLpTc6eil2Ad554bP4qSF8esOV3cdy0KqCYir53k2/jk9KtH3MXgghf0tNiuqF3Ud566oZNXn
pt/mCZR/+JvUYiG0JED6ziS9BQ7c1qOLgafkfd4IFGnIfAIPulUYVhGKEvGiNRnpoai7mHixYTFS
IJLvIvuqTmrtvV1mN6REN2owdWNc7ixZk0yRkuA91h5pCkDG0zEXWSxQjbdZcIWkK/ajdSrPDo3l
HsQjLGK35JFEzeicxDGoyrb0YUNQrgEMXoP9JHJVKld5p+LqQvQRwcm75zDdsgYEXFfgVhnu+aG+
UDiY/59rp5HluPhguH57Kl/RKNf7i0YCip0jOEMeH4rjN2I6rsiCZc813ttd/OZ3n9Qg4g7zd7zj
eEL0hpYDJQ9Z0/laLOdadT3B83vN0LVZcsMO2+6q0+45JL4DGzKxvrCUJr/sWJw3AcUnJ3QR9j21
ECojJXHGU1RKtBmQ1qFwt+JYKNowhgUOsQu+XKuELumppEPWx/Zgl8I7y7v4elCmgpB7qr4B9KoF
NEbFWW7n5BvVQFqhKBXCEAJNtyKckAP368yuMrSymJiAJZEsIsczy/jNole3m9ozJT/x/EVuSTb9
WM8QgBVfjOBlhyaxb0rvVnxCWTQt+unhq+HvnPOdipGpuHil17aZH08dkquTJsf5hTQn36pMK+h5
OkBJeVKNxOjGhX1Uck8tzqo8rAGI/obqOOKUoribhlBo8jFw/YYd6/vSSTsFVWiafFkzOJgXYgCb
A17Y5Q13FRce32QTPSp6V28kSxcq+JccnVhUqP7sYZ0e1sENQ12UErRF7PZ6GzhGz9Kzp6oh38Sg
JcmE8mHMeyT8D1Vk0Fzqe31VumBtU/8zUxizZfDbZ0H2fB8q+T0j+mlOYQljcQkCFKCmJcIgrKjv
fuv+32w+/ldIKzxCclH5BQHYPM/C37RGGJXo6DVHHU8ecUiIAs6BptOD9AHsLdJvMoUmZiVWyqns
VI3bIVZO9nByfQZSFKrbempvTaCQs05q1fAFubKVaOjXMC7h+BXGG2bMsqDQsjXH0g1H20LQ4z0n
Et3exdmfVVz9h5D2O7YqnE/J+870nXljyIvDcCAXkf3e0V5hT2XCb3s1jN8BDKE/XRU2UyqvccaB
w5q4GfUvYYYh3A7S13yDJvUAJiWo1QvOqLGOwrnV70eWiokpwxebT/PUR1G2+9Wl+eW9UenqdPFo
REAe5PUjXUZU/7fFlNBPpc6/n9hz9IOK8bRyPIMjoXBa/ZYfnYe4LQDR6WT8E/zYEUIrZvwUsQpv
m88JtXhZzis/NTYVkBR68oXz0EfsGeSRgxN6ORpBZWRLJPcf1ka3pMbFKCefhaLfr1F4xyXjW5RK
MB86DlnmlMW65QFFC72ousPgfSeF7cl71pAy37n19q9rU49bRsx9bMDrH0pug+koRHgM7Jg1+MNy
bUwjgZBbThYkZMrniFOr5lchUAQHqE0Zup/k+YCJumf+9+QnQgjs2EB1iQzPbmQcnDLowQkYmbEp
t+9HfAI21ztqiCXo6NqkP4EFWRcETG9xVA4wdBa6BefukYx2pufwy5TTv9VX05QoAWg7kVbAONFQ
ZrV04zGcwS/M+EumCEgcUFgnJUNIygbDoXIvlnj68Y+Klw3IyGnldA+TWansT3v+HQJDQVWe/Egj
6uUnxWNqorcvVh/SThyMrQBkUWMzsXAyCPj8JqeMLvSdivPmYbvk1Hsfh6ZVF9SRL7TI73OprQrt
IEY9CnUZU0WBgYkoXqcjEwJgkNMrHLYqw8W2LsIL5nrcuZ1RnTc4eq1AkdddIIizxj2dyONQfnYj
/ABfOuH7Gk/FAOL1vhOWgG8ieK3GfPhjpLTczugwFXGct6ZfqMHPN9g7Myap/zNqAUqDr8KCZxOg
DRGeiQhx1Sk+aBtWD/ZBPnerjWFv58mPrwciWLV6wjl7n3EjvY9dbygw+C5f3lMw+ogjhZqqaivX
T1KNEh7gpGAMGBTddNjzv7DkOyeIVaWTApLqD/XJl0vigxa2fiWE5yGSV+B2IbtRo/sX9P6Gbog2
65HjzNka+CMejY2i7qq8Ki4butfCEGrPjTzN5LaZnb9kbkWRUEL2RRvy5dVJLsr798K0V+pB0C7U
j29CR9/ejP0o0+zquHbAtBG46G84S0mKFgDwuXkDIFa94Vr3ngO3Qrb15YTn89MAUSLCA8EczJWP
cMgoMkCrgP369YH8GZJSCE+CUlfuX3uNIjHMhV6njuGzt8wtw8wmRZ55vqdp/fB/893EPJ7hEuNq
hw8KvHnycbon3YxPgc79agEmdGP2+ogE1BUiKgVToOIMWjNmeZYhegpQSe87MkUVJB6fyQPWqF74
l0RbRTqk1Zwbf3CXbuXiGiVa3a0b++uWjlJakcsa21rqgmsSXgopLiSwYMC6Zx/XU9BWhNuNu0VJ
oSDjpHvmFGDofKCAwua/5UVlARD1HlSdij/FM/MMaurAzLPRZpbIuZmBlFFAnUosoWTbDF3hneiP
J2vyS9zm0UYI32FEVdJkobedTeH0Wq040BXN9ufYG/d+q99nRoE0ysMozddswM5Tm/vcX/iuTxso
T1ALrDPST4zHUX5w4s+KFDzEkrHqGrzbjmFQf7B3e0Ql2fgzHBv/QfZl3I9RsVZ5FXMR7DncLyB5
VmH/NhaDjVxZqKRQaUt8ga9w1/ZblS5KcvoZLqvqd+Lxw+HUL5FB4KbqjKxHKpmOdSpGyNvHkvOa
ipP74uy30QXMfhz8w+Rf2nMiLPSrIiHIITnWW5N9T806kE9wjcQhfjoIn2un2v9mwVvPGV9vT6qP
zvLrjpJ+JOnxFk5YypCwEvY1AZEHIg1eTdSo6XuSWvBzpxOwj8rw3qO8u1qyb+qcMHPPQ1JC84C3
SjtgPiuZT+h4TxUdM09k7CyJwAaK+Zo0eGqdTsz5ApajjapYfGNZ0IUB+7SOacTcQw7jwJNoYFxM
RWMSR2AVCKeGEqYW2iNBtw+p6po75ugpAcToaclSpSb/gT5OyJVTTbHEhrIQHIozCByEV2xGJM0X
1p5tObQagnOE/ibzt8vBP/yOcMSHBa4s3WUsFGbD6aRyX0ypcrcmwgOrft25z9zcj9623hUaGoM7
OCMv/XYzvDOsS5SozlBKNN2HoLObhYSHGjpu5dINUaqwidMCaY5QydKITvu4It1+9IlH93eaH9qW
hiflsB9Q8pRiAmcKdJm5+hs1NW05FB0P7ECcv1aJRbHJTIuaCS8vqcYQ6HxOVJwXGq26e+tzo6TZ
oCtDiMQciVvhgcN7u+QK7m+q0Q9HwI57XvdBKuo5owJH5htMVj9WeDNfgsLGYK8lRbCTlY+25CFn
4oaQT9DyDocK1k7xeucH1yzqLe65Dq0bNBsd2E0RuEg8+9oVOhYc8XbQM0GM7ZSeme3dJJYUcx6f
aP+dM8o+r5nTcJ/n/SPhxF3K02DoF6uD6Uuv7iutxUpo0tAqcjTryflnxWzEFoKqQDqrPW669wEb
YCALIzVuQCItE+5XsQgO3GYalbm+2hYF0iMk+8BKPKbmaKqFrZgXCfUhGlkBOIOX6Apke5Kbuewl
TW1vsylnVUIJ/wXvB04ujl+I7XuX+6RZEcDPoWgEc825LNSY2jHgdFweimit0QIwIeb5rUeoY4qn
5Fa3nVvj+uXH+HDi1l4HszmXhc69VlYkyFx3s8iOjHMseIwA//XSCtWfmI9ogQSIhwKr6/VVl9hq
oFR4OlpMbD28xjQbkiYfY5OcYZP5AQ/79MTKRrDIsLVVI+sUV92G5mdqJSd5669xMzfzNgtEjcaQ
C82ulPYLgqTqHErglISyN4kBNffu6XwqqP2ZDP8hcupCvR9h526y4N5cufnRiLnFykS+G5CeIra2
OoF+NJeVmuqCNaqKOxbdwT5KwhoX32QW/mMuYiPYJ2QD09Zx2Ymo1AJ4JWRfzsd86JjdygARkDX2
byhEWPjI4hM/hBAP+NZXAoMiL6TGQ7aGHB6SvvoVttTsoMUwCDabKYzRvTk8thZnv3CSUUh9iaZO
xTdryK1c4fd+Lk0VbOefEwicmKC7w5YBAXDQtK+/yMpc4ohvFA8mJkikXqpmXyw2x7lWVpF0KHIr
QlhR9Py2iv3HDdSChQnPUN1fFAcauWQ21iwL1M6ZlWlT7H3E1tSJbBDDEK8tyVOOU4UcxJoOstSs
tBS/816ZUf75G4gYIjigeHEcOd2M1MF7vK3jwyQKCrzHfA8fIgybv5xBjfbWHK9+v3Uu8HNAbTjq
pYWSdQeJ9Rnanygo/qO0onV6MhfHbx4doTrqc1Naj0hfx1FuDbiuqOMv07P4eUJUlSt9DA7Mmkt1
BY+ion8zTTFmCzls2nXfIVjAp7++iViIsb6oXFR2Yiub4262hbT+EvSj9CaKhNHeYGIbtu4Uef8k
QxKnyGU8jMerqkbgUkcFFmSesSMfFKMGLxvz5IGYWk7VRK2CTE++bA/B91fX72OQt9/FaVVFeONV
PRT5YoL5w0w5ZldwlWc5Ky7kKzqVaj642/LOcmXnQgEzIVGpHP6oVZsI4d3ZfT/4jcocoFnyyxYH
Q8R/1J8uIGTMJoW6L0Hs8iDFr/0lbrevePZ/+Se28keZl3Q9uKJUl2JsO5OHkFO4a/P2J0PmGmdK
9iTJAFYp8i+h0aniisaMoL2qKxcj6y7bWFguwKDwT4oxgq3qbXvHIve/KYnQpqcSpYu7iZWUgP+p
vr6ZV2BTk6ELXfmAay5kvbQMJDGxQ0dTV2I/PZnDnd5/sU4d61XsYSmOfpFbnqdQW9nlHBE8ypMG
Wqj/7dbuT9kl2hKONTVq37bKWcwh7BHrAvVa6u0PEWTs9EsO/CNl8/alY55yN7sE0//02m/A9JgF
TxeM0/1SvNCXKSB4jR2mf24ke5L+akg5oasf2ZXAvVP/OwtVgZ/HmYuR6wTO1X5aBeti8GA0sr9u
72iEM4Xr6H/Yr5T9V+5WTvMJDgwLkV11jJT9F9CJhwsxQxux51h8GBX0xZdRC05oMx/irzmKYwW1
AOC6w8ZfdkgvI9puPadKXDn9+b0O3LarWZO3g+LyPX/npbnVmTr43eVBsfwciolIZdwqu9ShL6QP
2kTy/3E8uupbZUqvurzMRO8WWdAkQ9WGImcebRMa9blS5h6N+VfIZ09kLNu5W006DuPou3p5cuhC
NQtNrzBIIVZQgiX1jCbO0re8TpU1sxiU1j4/Ni+a3eA91d1IzQzeOlLD/hvuXVE03+UT1ibKk0og
G5xCUvE7PektJP7RdfQgYsi1uqlg6+QCPDrsSS6yxhVZMIwki0RfEABLeoKzsmdbPqEhjViHE6DI
Pgfz4tufbn7NQ6ZMXQcVU0ZsQ3kKMvkRskRwEepk7ojCHEv4yWJ4mLh+oJrw9Qm1T5cOq7WPBUyI
oT7uDMDed64qP2O0SyPo95h5R7k5fCi1aedDJ1TP9NnuBKjvuLDAg71MtU0E4pz47ZAX0JMWPsn+
icaHdLl2JFsyGEMacVOEZcIaM4jeYbojSHPuu4gpPU9fbXQ3asFROMRToZb7W7wjMCBEqoEh+0r5
Lke3jNfGOk5KNjwAOXtzouCT5TX25LrNHPhabKSlFfVxV5Ek6CUs5oFEQyUQ/2EelKkNW8vM9rp0
Uur5nWdO/dCofzdEG6fas8aktKy4gfFA3mROeJqVpmMpFXcWeBIUARlOQMK5vUxjhp3k+SedKuqS
d2d8sA9zuFh9PDEKuAp4jJIa6G0QecchP8zEvRxle/wLbQV33NTuR15CIe2TkKpBkks9pWEgQhiY
kUb1OAbOM1gaKGDEUpmQaUjYpO+JZfrIvD3ZAGIP55izGvILz9WUH5T90KTMxGL6/QrjtRm1+WE8
UTa6iPxNiBHPW1THqAlkIEHsY1KngsZyy+QytguubP24nvkjf9tEUAeiyfG6L7RvfYgDqEWtd42a
HWAhnSPG1TTMO/5t6oLqhuoBg+1klqgCnANrRGW6rpAYfAt7yqj4FzSuXMM9qfRxklFmfHA4gKyC
zXqqBJquuBycFpkPh+OW9XNLST60wyidgaNpeM27uSCEw0ZAqG8qeZcMtiTYDTaZQ6LO4+t58x1w
rlSBx8/WmWGBLgqxlkwVsRqG8JUj91RYube2EsOQW3unrIX5bKM+LcFMz4dS9Jem0ULXj4a7h57a
S3RRMtyurCzlE0Dc03e4Wmay78eFDFIw5tS9rZWGKViEev7IK99hi1ED2ssXcnVf5MjaTn4qB4KX
6ufNFMeJ0CC40Lph0Q4LDT6frWUGKE2sw1Gkgo7SUasyLzSFgg4iBtktmIsrTrr9mQxAioA2brVW
56WIvAwanR8JVK8oYSo6dkvCopd1aHL6/6afBHZBxsR6QP0TNF5OyRG6BNGkzoOq3HWOMJ1+JmJ0
f9GBZp7yoBHsGGNRYgwVpT2TNMhNfNb2xqJrjJSwV4EhIQgsSJGhMSevtC2I4SLSVL66GAcyU5cb
Wz3UVwV1JPvkaiCm2fltfZdVZKlgqPMuX0J9e4Euazb+cWCLXjr8HOPZCTN0/dUqyqBe/ETTjz9Q
AvIhK050YwOme1i7pAcOuk1uzoZVYaDE5tWCj3+c6gnsKB9TkzIEpfcCoOLSeCIVRiW9GPZzwSkL
UES3PStOUHXGQjzja28hYsmxs56RiaAJyKwQSsRD4naKrtuoSpa19D/wERAoUddxpUDfluCF724a
22wl9a15SpQmCJXCGHZiYhyYNZsothvi08o1uCMqtAghRgxruGJy7TuLSm9TLbpi691mJLkYIE2/
Qiwfllmh51UzfhZNdaFQc/d6uIrMaN3CidMMJb7QeCuEFCH4In7nBNcGYXsr8MFMqm3Pi1c7RkaR
MMLv7E5ywPIaq3VBOj69uoaOzVLQ24KIQeHc1yi2RuJHRdoREJJsFAywUZOY9QjxjI4CJnpO6YOz
TYRD1XdSSslFkno/dhPy7zrNaQ6WeFdfvKO2BZp47wqWxH8t73NbaosxL7+PTFCOpXq2CDSR75XR
S6f4r4LYnvLHA8aLVHfo8mPy9gV2W4pAaQx4xXFO/kODch5kB/ZGufAPWuLhX3ajyywFIcCQWIwJ
WtnHOEQZldSqciWvUvl73yvwy9veMMLyIRfrdmUkSn1ZMj59gbH7OgLhDGcRwxTetDu9Xvj5NZY/
fRJawNL+TnYGlnyX4glqXBUClSRNzJTz7bjB0d4xWC0olIEbyvg2vkjPrkpfWMI3P3dA5oo+vyEI
Rs7SZLAU+nw0P108t6ePwtVdApFRjAmUADxrQTTDfscoAbtW9cY16uDwIW6m+JGZf6+ybkaYkRk4
Y52FEoybcEZE9BCokvL4YlhfmM7usGMqsFtsA3VxoU+48DwtGmJup3cfWA8c2I0eHMgOkkXChNpd
thBTVbrIYzQe6TTp04ewOrUKwYq/BbjaqSoFRe/G3AVvr9EBaJW2A4vSdkhvcwXBJuUg5ZXhauJ8
BzD3RzxMnCX1+cY8Aag8bi78QBpIPfKPYmTU2O9sEU9UA+vCIh9rNewkP6lkjpNzGY/ThqfoHhKG
qzGmF4KODkxbv5xJDNJcPVWgUstRbE5bPQ1RUrE24QpAphxM7aAcj1XW1N7R8rIPPmR0NiPePhaw
0xV2q25XUA30JQzYSxpwqD4EXi947aHKdQ36KbNvYL+sTAv+7ZuZY41NgXmCNTqXVgs7z/U2Ab5/
cGipOU2Igz8mhiY9sjjHyMaxbmsgdArnAr6TkrtPpA1NCyxa0p3arY+gMlxATmzIbGFz2CDeeSyb
zkLFj0NiuoirkcuSTrPfElvKDxge70ho0Wb/8UUYaRVNPavWOAEQFqnRqatT2T1YJYOnoL8Z2ND2
oSuHOXxG3XefrEML53ACFg7JMgXmRTPA+45Z9gDECqrWf5JuY+cZGScWXxnte3OlHShIbrKUh9GR
1QotXkKPjTRkV0HNF9OgXqWE4Ym5omezel2ZKL2rpa0gxTf46MyVf2LwED9p3AQdNFC27c+Q/th6
iByukrkgmWVKYtGn+wsRsnOP4a6WzW+k5T2tDcPv4qDuDARvVmyzu542otP25eyVEu9Fkq9p6731
jeivnqJDODB+YYB8whvlyOz2gPbcR3gqEVRT3wt0F0bV4kz6jeAswMkXBjwhpO1ahQPr/93SNPu1
Xxs5V0XjSrpVI0eLBls4qU7muEROcNqsIvyPrKHWmhZ1sNitamuVBxaxcFqfFkzz9HroDAiFrZdX
GB32SCGdsb82n4wGhIpKExcYou1tuSDMqN62zuZgn483wTmz1qtHcyWx3OzspvG+KQYihJtxYmlS
yLMYmjBAEeU4cPaErCj2JIYuNhB5BsHjjvxx7xhvd8THd4izmKW6IqeRSoPjRQ8RmpIrpgTaZzMj
ymmYqhXTGhTDWHqt/EaUHk9pQwU+RmL2hTYsoIC1W9UyilJvrgXcg2NoQMrLFlYI94Qff0Kg3mAH
YMRDANeUwTULWlD+Qu1xV+DaRn6Wde4/AabCQNHBLnUiZXgOdpJ5OG4K00VZa9ojZMuTJ+1uv7bS
MarfDiq7SqCfJDlEwPXm2WxYcn9JYher2y6CgA8h/5zjEtXDyQPJzzPubc6JrHCOufOYKtmW+q6R
5g+7yVaPiHbVfEv0EmToyKW3ZQb6XAK4vTEqqFqNDofe3VKE2IBPXSKlRdbRE4DNDChkbCsjaMlz
aHqJ7RBcZdbBRwiHlD4DQjLbP4ZceWpYU1EqreFaK4PBR03WwnGExFyxkySuaNa9OkDqklvtmAHi
igOOu7IBuKIZbBk8i6/KkYz5YoF0In0/0nF2XGGO7yA9If1VaJUADcgMRq29DDGvuH3sNyrgQ+uN
eNTfSR3buCtlfMLG6yCelFrDa1NCXb0Od4w9SBLunx+85MaVfFhQoAx2pxraoe4bpZoaH07XXNoV
rscJULSxVZBaWsMMuOiYUfo0L648LG3O9O0VeD+8e1YbPgyPGh2CnTZhjjW8bgXxLoezjs3dvgFp
mS7O9LjX/wUrrQ9dsLHz11qEKPYL1BG9FmyvDwP9PdncTqXrss9TAq/wmkf7F0WGr3QfF7Om8nvG
asokygWKflUnYipKZZatHEw0EnF20PPOaEFpiJ42SS/suJ+ax/HCw7Ga1z9efFRiVXvkGNdEAQhH
zVfHghs0ZRp5iNi85wWVKo7KzWxWw65eBIO3nWUa8gxuclUBcCJfWTa6ZGwcJeBgyjh4dEEIO1cD
v8Tf1jNEy5JQ+xuRo18453R3jzMZLTq7RmIupV7A+06AY5uKt6XdBXu/2zR1D4SQ1Kp399fckov1
Z2en/99dfnc17KcvcVr00psQFa5ieKUw5LgQdfSeGNwadKdLWw0jZngwbjDd3MZYPN/ymW1fLiyM
2MjSFJthobAF90rYIc54RfCC/NRQrhFpiJVsjhCW5gPfZ9eoSh0yDNYrVmLIwQnjkbQKmhdfrze0
W1Rt05HW+WT7PN8EL1Hb8WlW4JnE0Kdr6Z/ApBJ/Gg7S2Ro4eEpXTU+oWVdcFVQSdrX42VdPoUaD
2Hs2w6BMuIJE8UIKKtH5jvvIxTRMZ1z+ZZwICxBizcB9KWTIifUFku9rCJlhR18bxSEw80VA+jJB
GROETM9SXVyX3ucz/JEdBIL8SLD+9SDBQNcAdGXaotz3PgaKaoVxpaMUQJ349i1pM5yGr1jytawK
JP4RW2kkE2sdu2S8wzkTapAwWyOvceF7MJ+AGx+b5ptRT9aw7lxmyS4l3amTBfeNP41guAiFFw+j
3xW56volL2vYfkXu+EfsoNaFnXU1JHC4/WytgqsL9ghFKajZuZLEaqh28vTgA4Gnu5uwx99K9nkr
Pc90SAERH8CQlABUUuys5ZVwniWuwsMB97JkQ2lHU0FRvEjYt3BiRLt+dAlaRdtBOCC4wtF27ZSK
LSB2y0+6PAdk5mxY70NW3BrsjZjDe9jjHLDo2ikyCTHci4BY8bw8CFr0WFDs4scoQHsOckLIkXOF
m9Os2Uv+MCBniKEMiUAPyh0tfBYYYLiypZAp5Q/4D9yjkeMTz27VOgCfzEFCDHlle2jK4JKltA31
Fv/Zs28nbY2qgQAB0999XIwTesbI56gsaFQGieWHxM1ThWYtI6Nt/XkRgDpyIzm/8Ps0BcRekK3V
4eK9sO7DNpEsQC90KYN56Z74LhuuWLHRH+L84/5gsAZQvPum4gR23Z/SbHI17yQ6ifoHjcWU/ct3
2VpGwcB9tOloHyKRgdnU3w/9cU7YXwzJ9dW3MH2N1NJyqE51g/0cwIbWmHHJKVtECjuXza/kdPq2
r9UaQWU0pp5lmC35uWp5HisklkTFt3nzOC9sLaPx0CRkzL88TwodXVt1kptxGXT3ChvySssUZE7s
lTwEN0Om5Et6XneBkB3LJvk/m3POFle9Ramhef8/s0tOBT/kzFClPHyTjiz8BKjqytB72vEKgcIi
5CFZHepVssKnGAiEM9tk/HLlDpNkf6l0Ul3JJBs3eHShxOsh+2sWDkNBbdIJlJk6nml+yplpfmU4
hRFtDaY9L5o8vTXTFeniQtmsTv6hepkc4VEPvOJ0xbwN1DMWkCbd/aPCbFmj1WV9vMGQGbLNIHfj
3lRbONuL4u/If+xxflmaT0f+nbP6lQjuGnXZxWlFO7Q+H8WNBDkWUpXLEUWKLXSPh202djK67jY0
DT8EA868rYBT5hwAMiRsh4cDqslN9bzR4kc76c9n4/ZzIZnJuphqM/IrALqel8lJLCLRfw1nMWwm
c90+I4Ie6CTxasv4/1ZgFb/C87SdBlVTpIRMbKlwSy66vCXpG2RD1VF7e/jo0Fk5gcp+Dpe7Z42u
UYiPekbKZfchDcJaoROOCaKywEIYYpNWI7Gf544mh0sTdx4VGtzQzjeOoRZzBNtX5RnhGTfxgbmi
P/zeFG5ZDRaz1yc5mTUule28vZ3E5IGrcN5yU5l0s3Svqraol3rUDomx3fjpUKc/P+r72IaGen+r
SB8Ww6HE+qpbqMFdekojTXPp7IJg5Ud8Kdi9Oq7MptS8Dl7futfM0D+6aZi/Mt2n8tIz0EAKfQvD
eb7SQWkpThVcjQ0O+auwcM/YJUspJDAQL5Mj8+v2NcnXVn6Io7HfqmmMJ9D3RDopwSUJaXMr9kcP
VsbEZuInEjxgtv8glNg7f7JJmHlSOkC254q0O/BR8JBxD/xZj3Ahju2ihaWYud3XXpysPHRqZoKK
dpjuYdwLQqnqb0mCL9A3IEHDyDsdSAJ1NcEITShJ3u0YHTzmPmulnpvptcZmgArw+uSJcXXiWx/d
9pGhqJozsHLeyllScFY+gBFUgjMsJvlJzk4MP4c9jWmsAfc+j8iCCG7WH2lqm/XTpLrzsfW9JDU1
NRGImzJZ6tiCawTQgGNOQ1IEC7q7rS1Uo3I0SQhxB+d5xtueScZW49R/fs0eQ57jrfcvI1TkEk0d
OiKjabd2RAQ4sm/u3EsiA40POGr5ADsic8xPiDknDYQI0wK7TPo3ll+8qvkpAUJb6zhaL6CrzqxM
xPAEPH1Tn0SgalX+4AlRK5F4Wl1Ag+a4hvL0/3ZWk2u/QmHqP5USkfz+vzQNOkp0iFGgu4rS5ts+
bGEpTsAzEEsgrlljam+GN74cbPhCJuAWaR/9mi5oC/+3XIeNOIFLvNSLxJHbK0SzZUiUsrU6CSS4
rS/1Nz3aR6/gB4n4v1jio3hM6kZLjVlWxB0RqEIlxy+qo3LI1bv4RoRb92SRkMaI+Akg9mbSWjSf
vwxU/ywtZnScv7TG+N6hYndfgI2B/xzgbH+Z8VcOJ2WL/FE5/ORFltlGNQkEPf7Zbv4FJIV1wKy8
279vqD3mFXySQxebLl3jBmJGp7fND/2zeARkltQwn+luerWyoCQmC4kTlF2yBSVu+SNsd0eljMP/
TUHjvHZvIiJmk8xENJ4jOf2I9/33oT4wzy8nrC+aIVwHU/QJJs7yoI8VQaYGfbuw/Vf3vvYfJJvU
5E4pAI8dsTPbyQc/d5NBcA8hFMpTsGXdAqF4qDZaQr3YCg53idfhAXq/ho8QoqsHbX6RYFCDB6QJ
7iw9E+/Lcm1eywiu78eIjMQU/ACHGA+8YLAdnYIP77AhyWL79p2ltVIKQvMy/2SKovAAbRUH93yj
VxCAiAC2UuYx+8HqS0jvcFHEj8xzlvuP7KIGjvAxFLebQPN0kVKI2WH9/mJ12ZEuszgul0q8Dgk9
h74+SEzZgUpTf+I+qZG8I79xKxARLkbY38Lt/h55G52tA1LMJkcUupegHWL1Agr2NZ1p949OnG50
0tW6nyJodXpMnxr8c/NCbY+vU/JgEKjLn/Buw42QiRlUdafMGuayFWKeecx9WBandXyg+e++HuQT
F62oFJzXytNBOtNOb2LqRY2tf6XTpkBDKLV/WueNQ6jfSOv9cRipet8zaFt9dXouZ3C1thgB1Xhj
U/RkW/3c5NDSNQzzCk5R5HQDM4bdtgYqxkZtH+eVQp+urkxxa5+blegygeAoGBU7naqjC+eM8Uo4
/hu0sKfvAidN2+KImSk0eQQbnffJlP19OWthukhsrbSJqFkyyxRws6G+RBfbLLka7c9IIa2xV+AW
IMhsqgRwgUi5X9v6c8/0nSiS3vzm3ahjRe0PXo1Ex2ODS7bD6HeJm7rNO7DEBcYeW7Sbay2v5Gue
ki55E+Rj44cF6SxZbztX/0xoSmM8ap7IpexkHOo0hsRmZ1gfD/UQvawGpY2C/y+MMZgbvcd+iHYE
hfCY1xKuvQ4A4bi7yvL8IFRTIVE0hlwNFsjQBN6DoT1MQH78NC6UFP6o8JBZXIVXBrPShK21/elq
vf9SYd5URlRK+6pQfZ2xfvq2B44393dB9oeBLqVeIN3L3p4ZJ6aXyaB+zrTQTucrGNQZYKAeLc0j
P0FmYoSS/qAyLF9BwzoQFhOPt0QL7Ty/03FC+DHVRU7z/rUrxbtqotcMv+gpPU22mZFEYFpXjKM4
VgNjoWnFgHUjY8BKbaWQterF0+DSL503qOIuIhFJP6C43kh3iNIReVudBUCK7pSUJXFe9uoHx61v
UYcGBHUI9FlF52+GdEW+mygVTaLGquXqBDirK9FUneJKLJ8fm7LqqEmjnDlQH/n95T9yzP74ODqx
zaApE7HwMoTTKqETgP8lOV7RH2IJ7cEgMpHz3F5hLxjKMbwR2jaB/3TWTHheJaSl5V7NfkedX5Mh
ZtdRkYPvLo8dAPDVaeUvbm1l5C3mLrg6eKqZFLXXzuseXkC2ytLzf7CHbZUOISBPKm3MVgHr96Cw
T57jS39lUI7MzBoihwc4RqzzLNYA6OrnKAjO49ABZK3ISnsHJA0IIU74t/ondm+BztsAiMc92/N1
cljHIV6GKo/Uqo9gq0izK9PfpbjOzxoL6kqrnzHhHUmLhPonOUL7t2ksN4g5Dn9G4SNidBN5Iym6
+PGz84nGI04DdXPQXHSXAnQlanvCQaD+a12slgXbcb4FxpAiH8IBWIpc33wEDhrqDD5UqimlYDwX
AuUK0+z1vcY76WeFnxFqywLXX3X9/aDMk1arEwNKfE6ZFLy/lWwGglZhK0KQ4gcAgfH4+o7jTMuY
PfIGgd5UaN+qGMtAfzbn+mXcutRrBDTDpah/OXJku0JlsSbuKSgLkoULJLA5AqzAr65TdQZODoyB
Fiee87HwqGaOyXls4SHEuXxq1XKNvpo5/EUK67sIRIMoFpBae3YuAqk8LDIxd4Q5ryDXeDPS7iKu
rADHLBWNfk/4glVxEm0820gH3dBaOeZKQa22JT3XKwNAUoYpuxajiHAC0Q7SyrbuKEeBSNjGNGjY
tjuJE20VrOBsGe8YsQdoFwfGEReOChFlWbNtc2bPR/GS1mvRACwRkA5B9gaIzIxIB+M7u8meht5M
TxbvW7zeQrbp93umQaG87wWouOyALbYZOFBcbGgx6cN3EKTGIh+PqcpmPxbIDylQm3+kA2ADXQHu
aPMx8mTN8WtT7vrWnk+dABrjy60Gm1QOk6tL2gsU57zipf9kwxHhMinVrRVmgFIZ3S0ETFB11aPp
YmU0F1s/LrxSGgTze8OKISKG8Hnsbeh6jN/ifXcQvUztUw4ZMVcvZJ3bIFKvGt+pL3epFK/AX/lE
1tFES7Ou1X3Kc6NEWfvs9bztIagjcIEkgsQCydzXTIgFF8pN/snqw0ztwFCLZYgsCkhZD4QOWxi8
Ek0eZLDgYJ6wWUquoh7sAiF44XnYGJjlhqpaqnt3RwAhYtszDPwhm9NDvyuQZ2DMcB47O4QNrLTh
0mALkrJjO5Zjd8Z14JorRGnqEflHDKN37OQcmF+4d3PfdNxUJhBCmovfOS8ezMLijk0GpR77nqYt
g+YFoBUFm6h9BAPhizlpKBgmqKu3gl+AOTF4dnq7QqB0xEandOrjM+k9O8p4/SEq7wZwdFMBMLdw
HaBdo7E9wuTDGfcPZy6MRD7na18X/tCIlEa8SY0aSOImqqTqywBfLroTCaVUk4+iqGpoBo5tAaZc
ho4OaZd62YamELpYMMLmEH8SkQ0t0shKKE/xefvG37N+MJy0AdW3K4nhWZK2Yge1qPiWNfxy18aI
vUhRRm6MPVrEOorPhHiWRrJgDWomaYgGQ3/OA6TvbSnxBq9NtLlzGDeWAqnejNirb16Gq9M+iT7x
IBveQu9coEFu0CGsScHxCrwYVn0+hP/WFsBxYpolsKuYyAEK9e/h5g5QfJRy5oAtWHBOTIhRblUs
rPAOSIau900c77P2/qzJRfvB6L8YvtDYAIU/1/3v93t4Bg2rRbBPNOyzHmrPhfxr648AmTMOW/9V
qRZHpIsp4Cn44IMwKkuYR/k4ohoT4J/XbDSjI/vD6U8Fn2w6qkSehgYvcZNDERt7RX6nVclh/iOr
FSPopnSFrkFGaapjSpgPOadRNTFXjVv6uKcDhyWaCQOt0HvJZsuX5bjMPoqXoCuUBYxc63A8V5Bs
toX98Z9ys0qk/vuuPgYj9LssJorOfODt7h2fAEyCGBkMOiFuCipukw5kL2i8LF5LZcQDoeqYPJrI
00bweH0x14LocD4RtNpVfvjbG9zU/SKZ/PCajRtriWkAhGThdblTtEB6+UPy9k+g3nev4uV2Aabo
HA5LbPSlhaYHvly2RH2+lKLh3WtFSWEY+0gwiXNJT2l4qoinPUoLN0lYOm5thaMHFsOLHS7ITdtf
56wVo6KCvalI+fs/tDbawmL4UC740bGHSfcggDb6Eung1i5AVnuC5hHtjN7Yaaq4ptLLvFz+lf/6
TQ/VLCFs9uqf2CKpa8gVNjCkLRc6Z2ZKse9Kkht3dOZuMgLth4GoBgIPhwwubJnElC7/lAg1nkN1
CG3EeTGJmX2EjMOFxx7BJYjs87PT6xarhFolhDEJwZAReKcLwQKqm2q2md6qgopQYyVuBmDaZQ+N
AOdFlkQbdbZgOJYDQzhgV5cfplgnAY08et1OT4EYiUdY5CKkGlpfiGrQ4PubCHpeWy3rd6+E6zbI
R1kjj0pkXihG350gAMhWPvFthPw473OKPLVK1NkedihuV6mXn8ifwGoMrTUEEB5clhpLHeyhF0Au
ORbflwHnw1HNcAk+K/zVqM7BgoqtXypwIn426GMUaMhI/Y2PtRhN0nFH6fftJIqwngEpPBC1bBj3
V6LRorfV0lhI3FzcvxNzWb0M8bmXduHD9vkzHrCiIiUhri+Rb1UAsPdMc3kfUT6/LQ6oGgnuTpxy
czpQ/pN+bM8X5wmL18B+775/lEL3mcRJlederTLukeCWpAiwzxtUeYTzP87jnJwHpMeOAQXjiYze
YDNTJKIxB/yGdV6Qa6QflqOaLCEmMsCTYvn/GNf3vQD1MdRzVgq60iusWh2PNYO+7Y9WNgWOX5kW
Kb5cWF3saSK+Ob2YBDIz+bdd/2AnqmFgVbD9CM60LgtwxV4D5wLS1B/K7IGprREpeEo73A1MBcMS
T5TlN5Pv7azlQfJb/+6zuCRF5R256dPJS2gW1Q9bjyeodAAgFsTh35PnLofiFI68xNsTHWvGytEP
7ZyzSp3AMAlSCJqD+vwSzFNB+JglIIbgHAbs+wmDBaiJglcOGh38tlsm4edX5MeOVSb046AUbORQ
N2eM2yfGsEzwahYh9n1W7+DNZUFnw9it3+ShJiHRKbymvBFinDf/xvB2oSRZprXHf1YOGIm+tn9V
0aoIKkf0LjYXnabxw2fRNsV/4k1EodwFxGzdvCz/pTCnzMb0qW2RyoZEO7TM71AFLWecGUT6zSTU
2OSfQPZcI/X/pTpTJhtlh80KAJihQWpzVs+LFGbMZstNPx76z3zCAujveFlJPOH60PxQZmlSSFyT
5DnKUm1otivRsDd/h45fRiAXcaykk7TQBzBHmjb1FZ1/djHTJindLxtTjLId2fFxh7x9BgFS+RUN
KHCKp3uq5LUEvAdufgPmLaFDOa+i03IsYl7hk3ti33El0Kl2m9gamDJ5rTV3vmUN6c0QubcV4qFU
T8vzhzqm0MjVFfSVUHZwy3Tr8zHC+EIEJN25uhqhc8ALrKJQ6ILxvHVC0SGehU8/bMopS3CoLi3p
WmhtzP0JpkePopTvAeRZIn9BTcdqUTDn2ZimfYbhXL7wXK4RKp5NAG6Pgi9ww0qSOslgkG2Tv+HI
jZaMKcqH+6jieuPSzVGZrlyapVS4SitDo0qAA7lxetjaxbGgghz0NYtGKsM+Da/hFq7H9wWdALIX
CpjsbLGqtrHGfjV4JkADOnD9eLimkB+qDrgo9sXNs2t+VhToUTebXKzorJHO+Paw5v6lfJzMWjuq
0gQE8X0LpH4jtstzEvHVhT/yPNlerPaBsfStI7xKyv2O4S5ienNrVgORt+6ATeN4Agx5AFuYJxAV
FjS+NgH+Dy4EysHkfGZHuC5IXNCiBp9WmymKq7Eq4/3Hz7syD2JEhpR0xhO04IIYOyj68WYTvqan
KBgpDZkBhFXBIpN6Y2HAN9ziWxvU/XYDq4DU0bNAXcO3KMbX4kmZJnd0AEBlmPHPxDh+rhVWld91
/wVGM5qJCG0VoLpikl2YEVpmFi2bjWUfcxp2csZ3QMMzCpAjC21MptGSeZ1tBZDzmZHomD5eGN5b
1dxSEk1S/ktf25/ro7dtTbb99dWGJivqjEb1JZVBCPBSz+sBromaHNigGjxwhOBp/qnLeG5uNQzs
6Ls2PzwwmxO3hCA3p7InivvIEIGUy+GEvpUCUiadNUucLYW/A8ltwF+gw3QIfPo45Ahf34EwSkRI
xIUO1Nj16K7mjBmZ03xdPe/RTVwlbxwyyVQlZuaDe+JCeBQKAc59zDFwnao6h9K3BG5CCscZ0xy1
Rtr2CmYjot1lFuRsWxDVS158t+Yva8kOhITokQUngKntU/xfQT0aJaZXmXh6fihHI85FWTfsPf88
VGkZX/WIWKMpo2xFXQMpIZe+P84uoJgeErdY7XXOtQJjUhXzjxr3QWb7lBdKw12qPNrc+6S/rMEc
RgfAiEagKvExrRHj/7JG4TgZ9y0GY0WmfVqepuvF73Za9N68whMQfFzeretr3w1y3kFEjlqDVXwL
viU82U/6Jjf+ImQ9jXgyL47fJW/jGfgOrV3mD4hmrCJfZITovXMvReqj2od5dNj6GZ99BfOShoC3
KlUZ/uxUVplf7ogx2i90x4RcHIdbU9cES7spAMOGSuBL+Jd2oG4m37GmnzW+y9g80o+Wjm4t4c2f
GnaNeiuw6LSztshCCG8UVB4opDN2HU691QLYTj3bI/7MzJU60FEdotw7HghOz21vZV2VJvH6qpVJ
Hu6i1hHixv87vHJYz+YGBjDRANoMeaamoSPq1neou0+rrBwww0JNf1JfrjMy7+uVRtMJw1fZ3FL1
uQszgit0zH/VmT6qLo829BGqJDuWFcZyT0z8dIEKAAsIsj2vCtjT5AMfIpGcNXVMLA/hq3ZWt1a0
jlFQ4lhe5hulFiWOSYqUNM2NIszMZesw8Bs3024alxXXBbG7vyXwKeI2Ibr7as63q6oKBjU4ozcN
Y6ZGJqKXSlQYbXlEkf8rwjddzpwsIaZ2b769COpvzF+/qxiQy4JlAcHMb7QKX/D4GNPMOpGC+Dmq
1tTyhe/pIAkYu1fbi6wMaDlYohY8wmLxnnecKXz3IKfKQvbB0vMgFmJhTwh0p9nDrKY67agsaKPw
7BUeRUZ7LakBw37mTiQTk621xiY6olym8MMxW8un1wrJUJSNdLPb/taWb8As8t95Vqd/s4EYle7G
bjf06Dace8WF7s9ZMKCpiTl/CaVDlAA82/v1lEBF6VF5m+EMbAP106PIB4AZiV0b58gQ7Wc68yWE
VyzuZ3fs5Ky6L6H+6jstMuOZ7DE7wIeufcnfLL1LGSMoBbtUv5mCSjjHe1Z1ZRV1s7QUJXavKxXL
iewzP5rpM7/mWCC+SrgYowBDqhutWPvJnLp4OIw0Z4jMj9gSUtFhyPSpv8T3nyUXoE0PBstV0F/B
FeXicwajaVlBQpu+5Tk/eqxJw8Zq0byH6K3BS2M/vZRSdrWQpPZn6P2+E2GW2Tj87JFgMBUkxqfv
4QoyK/ROr81DqHFqATOmiejSIqU/Y/wD15SVK1XuSHlKZgd9QX1prCFxfDyOmrgyPa6q0NFV2+nj
Y1NxDbNOrUS27v30fhfPdQIeVxLibjnnpttpSyATqQKEvIhTAJc0L9qpZvTa/4/bR4vz5J/8ZVj4
zQU9ovY+rcQvmaxDMLFa9gneKU7xtk0e9bDhfXDCjVeLB1F2zz3d0SF9r8L6EiUSDx5lZPAbEnWd
enCJ8fBESQJRxpCq0ccUTQ/eUo461cy8AsXoPBqsjx6B8TCeQFZsMUobUbl5OpsbeWZ3DnEpRGds
yIc6JXEECsJ37Ld19osyVUYdxcK3u57wjGdUA829IAliif7r2y1gpPMQMYYh/5NgLchQZicNR//w
gDnHI0JQJKGMgkFryfmb/TOYTk7WbFHpO8n1KvELKYQFEldqyP6V+Io+4V03adClfIcKaV5KBlq3
FwKnCqUNN0+Z71/dlIdJPOnWcQJEqgleDN1tGe3az21oq5Qs9whmtsscb4rNghop+wzb7Dah7ttZ
+AoTZNOz7Wo9/23qAdRrydnGFz9qCt3vgS2wstssn6O1NiNDBlHi7/a5wczv1bx4O+5sJz6fFFun
azMzWU5dLVAB6iDnbh7M44JXdds1MggoNQtvISGPNvkpXmnsVnieN5i0HQBZeSM95DrygVk+cSgQ
woTr/A7X3OBzSa8owKJQZHKPUOkc0nTh7nWVaXs7ssA1zessFSlhkBWtftG1o17w/r0cpnbue848
PVELkAUsxNBnwBFUFUMGYhjujnDk9DuCRvrkXMit3ZOaREpChVMM7wNrC50q6tk28/dNUd5vnRTA
QATAPOGaTYI67ePcsJ4c9NOdJWqQoRlVEVjwc51xdyseRxc0gNx7qXxc6gTe01dz1PII3UxRZ2Gt
m0R0GVeOp8nt9Pekp68xHWBAPCGcN+oKxt7un/mZtR7v1Y3YXthOGr+2DNd6JF9c0/cFgKfBN9AO
QIDgd162j7qKoyFYfyUPKqmKndv76iT5nTL5wIFsBvMMvYCNmc+GmWgaO4t3D6aBRnYOhwooslQv
J5g6qlzTMxxRzPDMBAt1MPBm9Hm7CHOyANn3jeFVo3m0XE04ektDjdCio0Laft1YyPCIQOaLUvXc
emCjEYra9GbfztnNevrONiC+DUp0uYI0nCXyXIAgUifj/Y5ZAW31OMYWNF0je1nRVMQ54sKWUD62
oatyFBNojTPm8ndVKSFyH7hSez8s5GhA2SS/sFloHxL94rn+MFd035RQrl+e0bztDP0O5YfVxVG0
LMq9n86D8YuFmdYfrp7QyYKd75GhqvvuQvQUISlNvZI0TPfOhDw1/EM/PZA1tUkbnzxUHM6SwwZU
A3Rp/4o+R0n2RH4pOlzlscISr5CgY9D6UFWXC82ilWtJlfqD3pwDwGgI1nNA90dfhGX2aW0JJvt4
tDhZsbDEi8SlqewgtahseuVWyxTH0SP5Byhe6FI+TERW85Bt75Nk7jp6ZRokrnmg2fb9Dhzcz+Ek
rNjs2BMxN6nmUHbU5uFMgJsBYnTqXCvLwirMkQhgmn3jLwjtSFeQFiKjDzbWLWMPVd/WXRyO0z9r
ivkao7qDWQUaYFxP+Pl5AomEQYJzwmV8CmMiwt1+adeZYIimp4viZ/x7ZA8gRfF/iGKB/oPB0+NO
uc9aIoMXM3/KSlWjWTeUBMsmOCKaHaM2c5ARd8e/ENE8PYTmlz+kZ9981PjzyJVX2mnzKLHSn3jw
/DAzJGELmHmz+TunaNg6AYOEUkFUSCGysWXavjh4W/xvL/2yCTdRjaLCyPHLYc+uVcQs1XWtpPYF
+f/QhKaD7ri/gXa4Atsbw8p9Be6sLPitGZnYrmxkgtCWtoM2/bAXU4qbGGa5BrGAJlgjc/rKCWza
bLxhO8ZpATdFh4cBc3MESNfJAOfZacuxsI03/GKUOtPSgZgdVHDRwCebX3ak2q66+lUoS84LW3Eg
z+YjnyBnXZFotmPSWsoB/Y+LL9/lsnIaEEPH6EwtAtS0pijQDqxPm4kl30aMJXsjEhxeGwLwT62v
KRJSeqtB4ZtlY6hntncUJFu0foiklB4A/jHGLAKiSn7aRfuNWZN7FrWunErL4oUF4HRUNqtEHW/G
Vy2qQb5+lFgwtW/4GDjUNnedDNO6P+Vh3hJQfWn737/SOo2b/43xmvVhZdtsHquaAYFDIRRNEcEO
8jZnb3pKnazuySxvkGTCwoKvgrs6zCN4rt5+onhANfWg7jZYvHa7CpIJyHq0uAkcP1fWWNUWHB00
6Bl//+JcdrFPAP2iFn++2z5S51UiQN2ulvHIZvGKhna+j93ANmHG16kFhhr0969dFtVHMGYsWslW
cIljh70wrmxAFigeA3tKQZm5TGqTACDz7Sc44gZ81QqPpTz7lQjr9nEVpy28MOm+rCbvrLMas9tL
kklUFWbCTdy5YC+pPrMQVVFs8jo9/vW7L7OJefMMZIuBolxb7IEmyGGHZlTeO4qfaJiL1fGIyO4M
Ww6dRz8KpOAhAQ3ypFlCHN7scPcI5rtsXJWnE1JV+J1B/g7mGI+QpbJK7WfHaeSxYm0iis3so/8x
0If8ZG3TNsa0UQ3hjtQXczhiPlGToLeNHa5vVpHZSyRwHgt501QOe5OgRzCFuHQo0P3Oy8vhGJm2
VFaTgT9dlPWsClm4twJJG/1FZAM1MGXYEQJAW1AW/mdXV5txp6ShqVjJ1l/R+goCjJ+EAy9RQl+n
H1rSr5DtX+rAXDz91n+0rj9wjNAoq4J/oZgq8MzxnRqoqPHPF/NUJYFuk5u/yLbI1oaEhhPGJ5oi
OqQ0Wy4uSSSIaq45B1GaH1VjeyRbUJO+7hZgXfpWElchtw8eCJD1+n9sETU+uR6ZZUbEhxcTwtGR
BA/xo8AWen4qUfE9C6grLumBVWBQUeGYg3uqlug3nyejL+bI3ksLu4k9Dr1hmp7UUS0GaP/x183K
5+mvUBzhAU6AWX3z2eFgvlBePqDr7dny+ZNt4TP5wVCvDcd+8dH412dxg51MQ8VRnQ/JvQND7jTq
F3lWrFlh9z3UR8XUCmkIjaGIobjOAs8fLz8ZzF955oTDqfvl/dm5hsCeMn4D1ghb7ZyJiOX582th
IUIBoGR3WK1b+bBOaiqfHCmK+xwjbfwMvuLT24K1VPqM/ioK+5EfuTY1eoOBiVSFzircmu42DeKL
P2O0CVhxVgjYJOZT2KvrI9sx4c1vFSeK8jZjnv2g2fh7ntCyO2mhMbBjmFTM8ztLzhE6Emh2f6NI
8END9lkJYyQCRjzA2Asdt7om4IZ7KcpABu7Si29CYr4/v1Rf1fdByRGQzNYLd1bW4706NeTuEf4R
bf318yN6+VH6lJZv+fnAHPz2B+cAG3YKoGA7uTQz1vBVzHMTAtyhBQmoqgHq5T+idKRJGxmREWwg
DdsA2xXkDRQGdeqzip/S7sIL3alAWryCV02hGNtK6qjcoCLVdqP7dQmX0YVf7hu6FDSUh/ZHLqAt
QGHZJXHlh441uLZ6dLyyNt/Q4HiV56I96ELbAqY/Qh9S/fFOafqxFgyvBfaKaO0HfNWkchrUaOJs
idMo+LAJcxwO7jchMKfKfsJfRy/1wpRTLig7Wv7ZsUhx9cLlRFNj5MfgRc9vgy2SWGukGr2/EjOq
d2DrMEH8lKUqn8bMqmAsGaBY+eBrMoepEqXUt5vqygtKadY8mPTaHaj1O3TgwjVpxADMBxc+UE1c
S03CcdNrIIS18LcTNwCctAQ3RsbA1cu94UoK4/2e9Xw5NlbcrJgg7r7af1n2OSR9MAEyHRRj5RvD
0go16xD/V4ZWskZTcJ4BC78B8IeRTEVd6jrJxh4azh7S5lrAgt1SjQ+iSaGwMRnAjr2nVuk3c5M2
3iDdfXk6Mlz5GiEhrx+ge9B7/RR4erwwVmCmnhqll6YmkAq2a2p3vFntLr27fu71IzHfnknpoSw9
jaIiu+/Mq/LaBZMkrC08tpBlvHzl6nEZBw0dY9/X1iKxU/un3RiDcQF2FTPWMsLxe8XiGtZRypCm
D+e3grSyaCJEIP8tnCClX44910+AHiXbfNd+gYIeYabH82ZcIQFZsM2n1sLQ1vb07bdwyyXA9RVc
KcqbJFNipbtPDDwu2bRHeZUS+QYTEbeN2B3i+H4XMqi7lrYkMVsOlFJIO6cj4spq9LnpqA55D2GK
UxXl4J1aivqrEb8wOQILwJVxtGTCVm8ljf0cjQ3krhO9DcmrwHJBrIHPgL7lpw4u+D/ZAbut0il+
dp/9YC6/PD3pypNm8fmk5CapWLf4N7sJeA4ztchEbSaxoS6phQagusX6aWGIxEbj+sD9eBYaSUFp
9Hgpb2SeB+nELRRp5+7ZBXur3EAo6SpaZOs38/PTJU0g6I+gQDWFZHT2fUVpZwlpcGbK9/tBtDuy
M8NiiXjtPD6UxLWmCWuR1kovTBai6Pq3yOybsYybG/H59rAYORGUP6cKu2NvRHMNBzvKSE1bxFHV
84p81VjWurRdzhEthwl3vzeUgBl3AnbYTJRAANzfcI1ef2fXZ3JWzYuwli7McwCxFfQJ5K+xgUSB
MIBD4l10UAFZ613hZqmqKf8rLGmeZT1BNwAG3NcsW17GnEWrnbOSL9Peo5tRuqoKfSvH6znxku7R
WfPgf3OhxBKkYfhttRcWJqyurvXqnjRd43vY1n91GVAkjmvDKR1Ek994QgBoVQxTs83C9IRJo+9G
Et2AWRD6uoCG/lS31ZBIpV7zTs+hqX8y5/AkV2CyQ/XFUeouJ5ba9BK+vsAMr2Q9ZFukOMXOfvFy
WbdHXdF3YbOFMIt5yrPiGytZX1Ui63FBY/SGEz/jkCxC2Q4gdzZd2h7ALTbtx7UAdx1n0IoxAnK7
W1GJM5B7mVDwAmBehflTXb7gJ+DR7Nyc18nPc9VtzHn4oIChpWAPxtjY0k3L/oPujryNMjL2Vxe9
d05ixYWhKyzg0jL44GnsdULcRudbJmlnq90G8Z5eInDbnmn4hDkaiI8M/duwhh/qaY+7ieuyuwyv
1fKunrzLM95JUL2CU4C7MOkK5uU36EyS7VE3GZKhVfGvyFq0T5bQNpMjrqBKCp8rAoFy9jAovdyN
Dr5Mwvf+ykfuBLvSY5hXw7BxjIpwTlYFs9ByNyrs2xtH9UiPE4c8liuVykhO6x47BJoCTxm9s6aU
n8/BXX115t0lxmKzsL2V9oABBdaN6VapI7qqArX1uSgLmgUMp8T8S9VPQyx9jacHE5i6gsMDknc4
gljQxlmqZnmILjUvUKSCzGQaOVkauUzosmtWiuhFD3AMZHJF+38mnAR/oJztMRvFvqhv9nB/9Thv
uhokvcJFRBFTicaiGuzTlnBYrVQzidYn4u94zVGCUqefzkUVpEfy0oRTCm5m2lAdfg0F3izmyUoB
UYBJzZiyY/v6TFOF2BtAp86ijntb8uViCpJ7ivuArb6vJJ+mT6Tlo1NB7dOVsgpJlp2AsgQPX/73
mniCDvrDZjRdzv6nUE+fol2zamLBFHhLBvNxwOhqqpockC7Q1q3h4gVOVICzA2yaKUtfWpDUJpGK
1+6kWcWCJ2fgo4Ro60WTjNff3uFjW1Kl3V4qR7+6Lr+wBmA5FPFNOJKyhhdhzCn2qXYHQ0dzH+g/
sNanKol65K7yHdq38/cDKU+phY5xqEKEhiM9pbsMDyMvuet+Vw1jalKIwl7pmnlQ8JzDU4/KgKh+
tUKgF8uTbqKVwOXB0uZyjj6oL9vr7n/DE12Klal5GF63KDiBXLG4xbM0j37PV0vB64BgsVPWuINL
WPNkQCaw76ax+78FAAZ6mvosIxpc8vHAEAoDjKIPC/y7Gq5sNWjfb3HMtvElgdmQScl83ecIYSZK
1Srk4/GgWqcRdB/pZ12o3EVag2TC4FLqrg0lpKVfJo12p/QMk/E99At85OdY2m7XFH8M2Xl0zFgQ
g2yh8BJK6f11OY6VkYhjtLoe9MC8rkzKxhtiN3obPIoWGjwN0OzMtLalCO0Lj36vLI+41ivxLiys
PhdkZgb9PJvbCHCImi6jgYkVe+n0KskgHtUzk/EYkIZgFLnGumyvxmwZGTVYOrvPIshVhm2dsUNv
tXYrEEXACJkAR0RGP4B5Hix98lU6k+kZwIclyI54r4FhCnVlWrE7EhtHVMOFV13T7MrZ2NHYoRSE
CQdKw6uE0ZjoB+FK/uIJ2Qcu0y5hxbUuD1FWc++hevxGv33CVRPpdyMwXG1aX+wS334P1Ga6trV/
eM9B/eNDlyjVL5Iaz9HA1hq/2VDfgGADjhr+XMUjCwDUcumr3bLse5HlP9hpFN005N6akIdgnfqP
V/I+1RzIU0IvOCnquSvB69bCJCPyWsUE/Kk2js3+WmCzQ1jAXZBSm9htkqPYMx4eoen4zWwXoLF6
Zsgvlc1w+7oa7mQHT8cU9Ahy2Esh4Fm6SEOZZ6EMWo+d1wPQb0lzF5jKL53wQaxcHi4FZhK4osXR
GeUBx3UldLRVHYNk/kjzdjEu9JcltRI28476+Hv0+puCSnXggVwUaBNnxoT7/mmJlUl3eBDrJHMV
tZOlQiA/qAOyJA0ws/ubqyqpe+QR7lJcxrbVv+0yjqoBTu12bicPis9R1JKCVn1kMxohvfjE7rtc
7uzZy49fasVc4Zt0NC4KgJOAAIH3OWEg/UtcF04o/5ryQJKqZvqvW5q+6/7aOXA791WBs54KZpUd
LTCVFH7/omffDI3vmXMFxxmulAfLHViSItahgHEHAj0hwyRZHLI0WtKZurF5gNbzxomdotrW98oR
SqV+nuuDYsYW2EeRGm3VRSINDZiv5YjXQlyKKWxyNYKzpQxXKyeP1GBGZEkOuiW221TQ4HMW5vQp
nZPCbyuW5nYOcA8NBIKA0pagOKPmiNwpkwl8fAeZkN8lBrUk8d+4LTph6zjGzOYJNlEZulQt183n
St9dPBJR5zhT6hKLyxEk2CVJuC/bDDbstQTzXFCH9a8tnKXRp1VBzsL0B4uIpNIviFslQU/jvtrc
cqOHUhD5/oRh+g9kOuEvkXReP1MgFVEHGL2huhPlXdkoD3tNIdFRR52INYjQYxu96vvBlNEkhddJ
GQwYZFN0+wnRk6tbxaPFJ83xQFBIB3H0FBmlE77KR/oJTPyOw7ELOfdtvA1QaZGCs7U+pcUWZGtA
yadlJ7dmL1mFb2Nt9LgWVzYOWe4nV0ttsYVYGhfzP0Midjpkd+mbMzr8gEmLU6R0472n2E51b3BO
IP52BK/+qu5a7Od38nJ8CtZlI04uEcaYqqhiN+qTcm/m+fn6AgewUmWd26a527fDxPo7PkOIbelO
TA3P3vG8fSRf1+gc/pCxRs5/tQo6nwrkr8tpSXJqvPmAzZ6zosorzpvECqTFeR5lPPJ4goDT6W+9
csp3zA5ka87vJWWCQJzW6RUHHwOZbvujiXd7y3Ct9HROhNoNoFbU7p1lafF7qNbchjXbr6/qsD6v
87wIVyaLtBPYBcM8slggPbxSmilzrvbJg95UgnjznQ2R733P2OYEuheBtDN28THcZSzwB3LrymNd
InyHUHdMycrpsX3CEUlGksyY7BDlRBsPb39xexpU9BmUnMwi/eYUZWMR925GkXF6z9hMON0LCMSs
71dSVNzbicH+cPNwI/XLjyVo/Y31eFeRjNNR+zrpo3yRrwP3IK6/vDLuaHMhVVg4KE833A/a6g14
cxtMXD8lkNLuynzj3DU+n3JRV8KObgqlgxgdsuo8xFRgu6QMg3bfyudKSBUqtrjLrI8EHSd1lv7Y
458t+bbIDzLqW5+Uo4DhSKqdnuvh65D9dsG1GpenzSWMOAlQIPZNWL8dTYwlu7Xh+5hkp1H5+HOM
6Wl2cF5kx7HDsA4u3HS1yq5zPa7zFcSabbsFDmP2exa6qx7x/3O831HuX/Vk/a+uusmJ55R9OxZy
9AVo0Jwb2FfovqqjOUeNE9KCVi7H5uirCwItK+aLBRQ8qQ9kK/kEtZ8Rklmzz7JBhWOnydtctc+D
T83RxLlE3fceD5EWlLWqPVFsUmECUVxqhRiabkaz9QlB5s+/MtSsVyujKCc1WSNE2yClnmKZUMjn
DKM+5l1Yvybl4182Pu5lL5MKWDrwgT/AZUFoiYwqoEVBihFJkoPufLfssADGfT5M+RC0V9r6Iry/
ZwyORqOCkATyqozo7K8lqauIYY4em2Uq+lUmBminfCzPdXdgmM7LvhlhsjVMlTyUdT/T66q/0RBf
7K+u3caNrmgoUgj5n5X5uZw+FztbfA+VCew57IEp4BbkhxJEElk4UI6o6SE5FasYksRqpatxclWM
UTVCBHtMFFFm8AZ2EMRYyqUC1RS66yQ+ejzAP5bHP1eekFEoSn6aA6awt8ltSWYc2NEHEtm4VonN
EyRUVoxHVo+uQnaVdCh/tHDoYtRxhZJ6It+UBhz2pFKeYzY2fXzu7Ki5fhZBTWQlOr6fEM6uJZTm
3JwVTbKHGrLNaJMxtYIJyah2gyiWyh1AETe4pbOlPwIgBejI+UmnwxOyJHD6McQU1SPnqPGIVlYs
uY6lZDT5j53depRqRzNPsxHkdClCcQ7YVAu5RZzeSPgka678/RS8EtLBrosG2Vvmvl22skvDscye
oQSfTAENBK+QTaPZ3ov/z9JFkVxDs8RTL/QBxYoIA9t0Xl1+T9PrjVV6Kaqrb4g70w5vGPLMYu/o
3RP0eHMZus9AiZZRrJmnvpeu3+Min6xShtTxc8VtkJda/6M8/SeETkFiYciY0/Upim4upYdC+SVY
XG5BhNN+tjUYHuhmSU05Z58BcV4jOhZPbkoaKgrqI0jjHysX030yrWzJQwAOzMjbslwSu8UJRZ2s
6dmBX5ZWwptB9+RpPp2v6r7qniKhFtgI7QrU551vkDymvt7n3Y0yIevw6sbP0yiatTYY8JW1hTQK
NW6UENhN2ZxHPwzNysYSIFwtz7+WtU3g5NewoRthB9hvJAKEccMFwfCPdRvFHfpDYHUOYOu7A/Ln
R8RG20wo0OJrxHfkLOH655BjRpMNxAqrZVueOLIsHVExOcs7SiCymK4ebpzN86fJC7oPWYNrFmIV
07oE5uYB+I53sDRfEQHcEIdOggYNFHYC/lcoHnuC+v2fpftXXVSG93mhfLQo9Hi8li73IKEDitO/
eXxUj8hqvnn46+emDmUnYk1rNDpradV6mzgp3fIGOOmes9vTQ2b8IRAtgqOkK+Q9oKLIrxRFMi0h
YyDZi+eo8xzm17BklYWIdfx1BaPYRoslOtAL8QlhCEbVowDIy74uKkAFyD2jgcvHwMcU8LgTa+4P
lDyE3lh9jSizdKdzfqNtk8OPTnhBrU1MOrHMBU2f2kTduE02FxGgo4GtiZSJhAPDuLpSKWI8aUHI
MvV/8OQ38H9+CYwXzXD0ycGH/YIGxpvYsCYGSMwaCmkr2AE0znQR+nz8NvtEKGFL2VOeC7EVzgxk
lYNET+Fd9o9lcr6dhm+UywU1k+1saTzlKTWv5l7TlDm4EDg1jbZ61jO50a1l5pcJoMoeXoiSwHuL
ykanWmLrfsWojx2hiiESRYpTyBElC/kUA/OCsP5XReWrbxKPtgF/aZZVxF0IIbZ7y7ce800APkeJ
NKIBN0Ard7soCc/QCe1af6SSGMl/qUSNQFs2XPkTkPWuAzN6MCnaRD9NlAiE4C5rvSf8Atj/2mRu
7xbkUagagIfNfyzSafi5Bvp1crB9rPznbVzSM3pncIaxcmt9I9lyY91Jmh2GuibADEW0TNXj4fP6
scuzTiO7++t9AvXA/qyOPADywy5QFehmffIKgcUEMATC8t4W9GZH7UYzRq7OfDtYlgg9adcMTj4I
DLP/DXiAhzL9gIHr8OSd0lbBo3YGfD41OzThy0cykKkUFldTxtwcPxImgP1nR38PY4uTQnQiorQD
0JBCyd+att9AqXUMHRSzOR3n1Afzz+ICrPa5p8N51UTLB//NAS3o7099/QPMjdeLiaTdNY+gx9KY
8RfifSldlPL+4IH6EmnzeMu1if7JrWe53qy4H8GXxT6XbbtbLVdCyYnZXLvJ1gKDAwx8s4RFHfy8
bKdlBhmaic46I348XyRZHAfHS8PPVV6C41MPo0kwEKAGdbFP6tlcZsoLCdTl9lv7auvlL8cVbC7R
SD5QtXSLb2kWPwA4gRoBEh/aYtpuDP02or8Kcm+0zt/62W9+UmacDPD2T/DrEICmjO2MUv2c3yv9
gafM0WnWTNg/5NzqjfBbi4VPrqm6BzyAT+Ag74JFxbGYyBpH04m4WeSI1Z1bnWmXoUyWHXB2BfKi
BQBQbr7V21LTVp9q9HrhnlTn7sIWg0e+81dUZRFbYJhC1AZYulN9tcDfD9LO1MfXcpLbfi3OOKp0
45AZ8UEyemKk5Ux3yNeCVEIV0cZ1AmKOJqO/SkibfjbhvzrwEWZO7sPml33vz9CROq6YMobGuZUv
nX89ye8VrsUop+vL2MS/kUwgfdK+fKc2lWc82I/taPPUlzcGdsZ6lPA5eTwT+OIm1MCpMzD4ZL+t
PntmwcGnMTxuVVNEuz8vjsn9BJv5co52S1aiIpt1b/NiyTCmHYvDVRIR8z4BNi8lPlUdqVn4liKA
tiTYN2EVOkItJqVyAj28hKkmLEhPSijBX0Vt/Qwul0kUnlSxglw0SUQHQh3efUt8IjjY7Z+FmhhJ
r0f3VQGf+yZREDDsDILg2n0O3znAUt7/IIt5rHocXkm2L38dmv7QBOlVsLtSlRa9ZQ/zXxhXL9fo
kZm8D6NkBAnDBI8rfQQc4xsb+ed2bkJjtvTea/Ygk+fytX6hG3B8sXlSN3ESozzVLtMWO7dqmoTA
YfjTMvBKbpD3HKwuMJNO38wYZOTbSS2chwSASrATdZAFjNxAORLwcoYRJk1A/ZVu57SKeLvFPxfr
+zJQxVz82InJqQAEFxL4/wh6m92Dn/psfCBzRt47rtVE9huCjvyiCksUcWNCaQxkWjP55GZKq4nE
BHxYUV6hjwfqnlVApKVR07zmCE+N34Xt+ViumPj5B7DDHYXakXaDIAiorFGJNA6jHWVzaeIC8fh4
hrANfyg0v2f+5agMXXLsOwbtMYxb3fqB6buejXci+lveEx0XG3XHu6nsY7UwbvbKwLAR3aczogXH
7QjjgCJgV7yC6klAlRe+EVROT1Bzwy4kcpWAq00txUpR8pemceTMSkbF4hheZG9F6rp3bSFIiOlZ
dWbuaQbouD4a8KqV9suKVxE8pHt3Wc0Lx5EqqIA+pi55lkRWa+K/nvGzXBlHc4CUJMQIXcCX9dGO
kbNNJazFKzZ3OJ6XvzirJEwArUMzFzbIyGnui1bFfOj99u69+Epg0GH5+1VxmkvMUKk+ngqJJm9x
T9yQx6/gikeUlebWcwBgKSXljAGyCzPrJKugJ9NqZCd5nWcv9SYTiVFAmgbckMtlhJyXBJTEIs0T
ReFT4cpwF+LfC6BH03qHMA0dUJ/8+vNlkO3GLc76zgzk0Kc9R34GJQrefNWajhVioqQpsFQOgZwA
/QOrTT+EZr9YJuQjM5iFkXqy7YdfFt8YXX74EIBgfX64kPE+dddoZ9UylhhvpJ4HwFhebdANjFat
z+eTPGp20Uv0gqZGdQ2saohBnahW2Ds6GAydgAyYyXU6B5VDSvupAmdco9nUgAZSNXALw6fvHI7+
Gb6TL7Uqh6suXsdplpYnJcPFMHmQpIxNVY9kQGDb4SonNFJT9fac+sK53Lw0W5ke11n7PzZf324K
anWf7h2b3uIZoD+LmBzJkwX1uObuGif3wofjMaJuHypl7Zax15z1PbGnCAzCGf0pJB/OMcy5MUCI
utmEnrWwZn6e/M5lGcfen4CC3dTBoU0XYtCdZu7wa1+9E1izSTgHxOf5jijR/sx8OEDi+slzntdB
dHdctR/CGBdPcQfikwKiaoLj7GMkSKIXVihTxDE+iaFm+Z2Ojq9Rh11qGw9YgOlYLqzTIKbZ21NE
Vr0j3DfL+e8JgmW4zbPgeDFlQScCJWLl6uiq0R6fmQGecQP13Dw7yYEkykR/eml0sNiMBfCKrmzt
AoWrt+mfmPKfArejWUjRtzzt99NkBCJtGAWgsC6qzVwjA5gnnSdndoGctllZPiZ5NYd7QqonXRhU
bOQ9hP2yL5YIzE3Y6Rezo6ComNuPgUOwDE1pCOo1avWPkH1aOTNgIpNs/FWSwZQUtjJ+B95pJi+r
pGSGB+ma+Qdiu/BU4+SfAgG28/FdLEMefffbm2zzPwPcEAP7ymJXUq2fIBkcpbWKpZeNf94s9r6K
CS5hGzcEBA0VHyDTzu/en0HYFodyvvDLTOajujSOkr/LR7CvJNy8duwpMgWNF7yq1TEoI29y/SPP
+0/C/B8fl/WmOC/etDZ9lNRq536WnqW53e4K4jlp7wlrJS5hBMZrnSFEdaOT+7bBeD38ETRvEWzg
PyirshVdk5dOqS/BUhdNswwRmdbP7HjaFr2k+ZEKE0JwS9e1v9oUXeuxP3mCeG4xrLSuPjHfqMSf
RDj1TTip7UYlmKhQcn9Mx6pyxfSO1j7raGRxWcC3zUljO4ogv2B9D+XcboRK1z5f+Ukf4sAyeEo+
u/sTh/+KG0uorNG9hMP5vKO+tSy7ml0g7ox+GzxV1QuOzhJ49vIXt8XfvvTV2f3+R9kWVPVDYPfZ
vJeyhohwHe1hlEsuk9R4NOf8e5h9E1AHJb2FhxE/VW4gGuGDkUmaTL1P57Cpti1ZqSJnS8n2RQIE
yDMWGCI837zeYsRd0GkV9SPoaV/CFdLuL5VxXqVHTrVZHnMZ7E57knrc/AD0lY6+us/KJfbWy3j0
8tkhthMFVhEmWjEUU/Nvf4rUq2jsL1jfcoKTleQSsZwq6VjycIAC5w2n1wBN6+4LcDpVj/J32UCv
blS8NjXRAFTIl7iZtJOLeX0GZvJMTmHlCgSjN1l9mupLN4iEWDpLgjrXc4dCi5tjckHBZeOOOzNo
gItWmxlwkjudPNIxBBPH7Gd/riTAWDHt9iuWSXvRBqyk7SKyyE0ufJVn4xhOWOb59cOdjbB1b1iz
a3+pbfifS2HEmV7urxq8ql7UaeFsjTWkpIB6GtIBKKxLBRn2acLsDPHnhYSNvc54Jj2hXFMJ5xkr
7wtY/vSO3apMZxgrAASLZ2l7l0Yq8lDdmJryo2Bwkh0QaGBRpL9ZoIBObsG2wkQlFRA8nNylgb61
Cv+nBnhV1c9MNVonjx4G1LUp4EtPq9lfmpY0nN99S5h40wvHLk+F0C+hBakDQV9bXkHbfBFXf4pu
BVELZNyS+mnOvIuq5IVTcfR0kjXnaNwWmMMjXN1ktnetnac+jAcUdNa6alG5eOe7ubgoSZkcIlG1
DVqExZS9CEK979PYsO8tAlMLdVdxIiPDAZyEjEjMHW8XyiAEbxq/9vBHTO8EA7HvoPD4wgIuDF0V
3rypcd0yCSsfm29XZ1Sp7cvmRpnDrUWk1pXE7uUq3k2TyOnTP2RBB60TYNqvQZsSxkkOI1YiIwc1
wpce6peNKpL4v8rQdll2zSS+8/ZXoe0NAcfhvEi9eL7CrKbe7GrvEDR2FoBj3UcCMCHJG9v26Oum
Cz+DdJ09iedMYGxJUahnrptw5JTd+QCwWU7TEURqImOf+Cjk+es1EgYiCrRCCMYaGBhqnNT3DQ4J
tT2juxLy/MNeiXe0/OyELsHBJ+xyNGC4V7zMsI+TN2zfceqFGUKUxXpwU0FVhdCIecgk6pVcrJ+2
SlbRwLTWz2W42gWr1ZoXSAoNWRb1rI9CH1zMQHX6C5BC2oOX0JrV4xV3+lecUeYawS3eHRIt3alc
2MY6f8Ni6Vc0FqU/83zInV2PFKkMh1cuHgC1ZAnfwZe5Qed7Zh+ETTDUYFVhZnt++g1kHVyV4RTi
6dabE9TWQW+A6gszMK1/gUQDo9+dGipabKdOk9PwjjAgFTeodIxXPm/2geNKli006LXOpsUvMrZK
mOhwhXQh+IEDx9hUtMiQFXdRXvUp8Uih+XUqW2DzB0NwwEodv1zf3f1Jw587uShNnWWjD0lkHNqM
InSTuFrxooPC5sgFfW6Yc1xAvgzjPD4mr3gBUnMQWSvuOKr2N4FnQwj/JuAPlmFov2zdeeIQ70bE
1H+zYKqEZB6lAOGcgepgxgd5NGbOx0oS9D/stltsI8ubAC4nvX5kwvbjdfHIkJLqKHB6RbQVtwfs
CqBN6j2s/9lQI1NcYQ9nDyUY7en9lUdRRVJCnOrOEJiooX8kQ+vWC4gRusMkR9XqL+k9m+1Vhsu0
35ol4ESrw0LhmX0Kg5fqhpD8tn9Jvo8mWEJqlNbqzZoPDuU2n4M+yKoLWpixonSc7XGBoPWL5qN6
4dAzW5ed7TCLBcSWKYKGxkAlxmFgQq4Z/Sa5xf/GdPgLdcQ+tM9HbkkGxhQTrk1Y1Cm8XwQD5nqL
KyyaRdPWiBAf0Ns17lg2+lfoHpEF+77b7ZQ2xxUQdxWAPRZqG0JE/bWv3HpGmwfOQ3adm73k7wjd
/nt2Xs4T6Xl+2rUbMB0ZcQYc+xea10fCk6Zj4IacKJSg5p7AcS1aymUU179x/2zaNkRgQdnB1gnp
Q2T0Gbz4Fr00aJghtRl9d3BXYPV1THm7wx6v48NmCywbvzacHETvp5RqGmD1gtOWuydZzlUX67ni
4vA8PV/+6s83I8ud0QLDhRrTyiMI1Ln5M7Rt0w/QJVbKH7wUampe7JIcgz206j5kfDonUtOZ1fBQ
mds4syQ8Cpkw7VZxJzLZ2UWtDBEdfq1vZMrgKcvpp5Fvmu/7D/yvE60OEhdcQV6GSw6k8XUGp4fJ
JC4PW+9PTmyeYjLoTgz6ExKib26ucA2oqjJxYuC2pX4jekp5MxUvvzRJ5wz/+stkfZHRo4oSxG9t
C7HFObwMSnXf/Wkp7M6iz6dla79E73v9L1gPtYnTVqkEDcbEcMMVmpj2Zo9i1zG5kW9fwzByF68L
nVEcDgYJUUcJMUxxGSE1IAEUbFbkk96ox9lSss9o+Yh4PJip9s/8Rb6jfaOOc/0SbY4sjw00bt0A
JwueWwMQbCm6IiiR95jCnVCssm6dJWQD+Pv0ZejHjJNyAxxhEnvuCVqMJDg3iZMrJr/qa0E+/cbW
pUR5/8vNz7F1Nvh4MwwAVxkFigkrBro65Kl0H3NzQJ0watDLPOa2FiSQtU8KtYeq8l+XZMzWG0wF
OWm2yf+eAorgIfoLKO5ZUf7hlxeAXrKm50Oflr8AdZvPi7zUxXmtnBk6y/GutmBqgbI3b9829ym/
rHYhmtBSfRjHAxZ5o2pLSL6GikDK4Im35khPD2oTRX5Q1urO75tf4SAo3SkqqrYu3n7+pCJ6iNRR
9u3MLBfkQnf/BKALaamQzDWkDviGLDDiUMXIC8rwTyMZfQ7m1kYNInnk08307e/207SPTCURPDnD
BgF2qAYU0NvEl5aitZzLQIpJRpikWlc1xE4kRyfAIm6Ykz7T6ydnEdN6ig8GeV2mJRtckXEWgoxq
QzSJgZtoedShCoVWs29h5tgi2eazK9sri1IZ28fdsb6NH82vRKrQrPNd9tqc2NAuzW2cyS7GnJew
0vlMwaS+shfKncknE+FLNVC2TeWuLi4sECEDwt35FHMMfTZig+O+O1WhBQtg+q5to+1+obn3s1QD
3J5EglRXY+jF93lG+zkruCmyfTgzZ6hwe8xIAcUKEbt46Ck+KPv7G9D8Yi4TvoulkjUNZEPvSJrh
gpFdchAGaaVMln6PKhxRSLp7lf8u9T8Bhg88W4YO7e0OZ+DjrrNREG5vbPWUvKM/6TjyCMZFQitV
ptOqdKt1qUADBaipcGwQloel6txuLcPQucaDscREI9Kq1npouoaM4gBwvzkqUL3bZv+HQGtaW9fA
X3DQXOH4T0047EJUIxXWmRx+MnEWIBEn0PswjQ0y8f48M7pvLQBdxqjctsT2zOalDvXqMwB/tpmT
45CUd/vwDut5oynFeaW3q9BKDtOt6J9FwBn0pYSyLbTOZWubJzeQ/0pJMFsbZ3um7Erdrp0d5d+i
VrnEw5FiKy600BpwCHEcifQAzMR0LyfoY4sTfTf4KPCVk3wwg1sEJaE2xdYa90R52+OitbwjabMC
ZLo57YRP5HJuUM7Gqq02djAMxbjNiEJJa9L8ESCcxS1hskOKD+epEEvN/6c24CNjyP2dnFhrDNIb
5r8bplqJnu/DB1Z0dEqExN1iFn9n3M5Z1r30hAHz3KJgoG+Dhi546fKDGS3CUqEdazqlzVkCpWPI
b781HfDh9pe0bUPrqnP0pvlEHuhsNLvHOtXlisMpjICzvSBZwoJ8cJnk6bl2EQ9qTxK1TMbx/23T
K+yW1UXoaCxqZopmOItUwCQXwuNiodmgsvUlqov7DQYSZkPV3Mo+Qr1LDeaYmJtdVnq6D7yFlXLm
pvu80DTcLlm01VIFAGM8EJ1vAcMoGNuJFFfu+qty8bzcPQDTJF4RLKF5Ut5DEBdxaRP26l8IjqcA
aiZnZjB6uJvGf3Z9lpl87F2jOLGjRNI3xsh0XnT1JlQqnyD/9pHSkRzfISoBptK7Zuqsle1lBVhq
nOpa8qtAYihw4RW28dmFXd+J/I9+mQrq5wbxoIvnPkyubcoBfRJgFs7kDEhD460YR2p6nreJfNIr
asYwgHB0AwV1/CQ2gXQRO8qzsCrqmi2exgMWov70auQK45qzjQwu1n+GYHkc9LbM/b39J3jzgiKv
JWWdQrE4bpfoia2IgL6UVhF5z8yz8udsUu+BQL9RR0JdID9lFF7xtx+F2GMsCu5i2OyYupM0LBWC
O6/0b4ZxRIyJNXptQr34RJbWER36unPv6ETNyot90lPOV8e7n3XWfNcf4on6/lkhEH06Y1l1/IXg
PpFcUOLkDOHx0p0oWAym3FP8TMe22z0kCAWKQ5+VRLsOspeCricH7vGrf/7ymQMgMhvqlQD38SVW
GvTXSzVWVCaxt6SxHTE/cIkYLV/qV650CxV6h1ySkPWeaRjMBVj6F00ZTK1GZNI5jwUVIVpjd4U+
dLN9vDgDbG5/pcc8vigtSsxghi9IoIKSkf7hGla/7nm2fbY1Qkp1/NvC6E+WAgg+s9mlKKXoKSU6
1g17cL3/KkA3su+L9QAYUi81NFyuBARaxzZMRaX97kQvkGXNefGwJWPfgMxfgVEQiUYNSbldlS8e
htyhYaRPvHedWvgjLoIDcVFIWKfWfRl0SzgI3LGeFcuOW4P1tojCd5na+WS2ZSk8qEzwiA+NT1NI
5sPqlbATu4jOBiPtjkIgcj1WKDmmOvOCLLvkIZXC96kpz36ab+EXyhM/6hVHLbrFLAYUnjbIqDNP
VrEj3ForkPOg22nzskxnuHM9VDjMVquMrFeFjXXOJUr/YdmUs7WTRHIL/npuwUAzdXZZVw6/wRYP
WuDRcT+/y0l6U0VI0luHzUgUI2tYotrzTpQ+xL6lXhgvtqe3XBJyoS/jtSRceiKgha4F3n0SRJpN
Mwd012qLZ2vid8oMl8OnQBsTdEEkGST1YGhPtw8b8wY3xH7bsqxj2xjXU6uL29MyH0mSfZXC7Bk+
+LyJQfuRnceLn71yp520C4/EIjXWz/c9nQY5YUH/4sU9VtzymaFmjZewf0cf9n0fUbaEPK+floAq
7JQURcaPKOw8MsqzHnDpZwG6ImGZU17q6cyVzJ/kLerK0xwGc5pnbkuBunY+d+eWqNzTXR/eXwvP
4PY89iBuL0P0uc88Xv27ecyCNCzfouq2IQjsIyK28ojmrcEPqMnhhy9g+Z+DPRLIm/qSoUrYOdj0
wikh8vq+oZZ/q42XXd7ydzpNG+LKph2VZCbA4B4dGm+kgyBKFLvNZ4Jyjeuhy5ZJ3jmPnLql/w04
dZeQGjFXGIzNA+8OHT0H4i/V3Fk5jCXRgqmWCRqhqiCJtW4MB7kpKGRwfuvpl9VFKU43y3onVW+1
RsaSMIIw6RpD9RUoDecL726BkBl2bHnKqSIQniEirlyFmr/IjsXNs2OZa+vJOgC6V37rAUuKt1S8
jmeFYi0DUUBjrM1klfccdhjq6YvXDLoy/5tKq7cW9A27qHWiJ2alaH6qnoJcXAnTRarjz60+TBf1
A69rdQQQiLnoyTA2xCx8hBbbvrZQO3ZbyCS456EgQhbBSKAUVS6ZFHYCPU6QUq6M7luaFVg/N5g/
EUuLAyqzfRa8tVJR0WzL3QZQngjwzHUA7JqzpLtMYXfVcnuxikdfEJV+Jeh6ZS9tpLtTXCFqKO4f
Oy6W9c5kFEh72JrkIksNXxPKp4ZwrJNAeGDtU6bvptFb6l3kIK5qUVRD6WkjlglDyjxypVxplUIr
SMtUK7rXRUG2HfeYev3NXsQ6RRaWVfe7NebDowCQbLZ9l8mOj8Z8N+E86wjEcjqLn4X2+7Zk/aln
WvGGK+KgdOuf643UKbMEmHX4VT5lHbmvYDEDAKOA5/raNLJ/sjGCAluUCA956AN/nB1rVbFGhbNm
26YlbfJSPan+SLjM/yPWd/y/AExmDnw6YTHhJ9tsChUiCHeQPjj8foXd0AIWiXY+Bv6e39zvEKu4
PAFgjIh5tQW/Rl5c0PZnCpoG36EbrduRVXSS4cdAZ2ZO+TDO7rvD91F2ZhP+ammAZ7wt3qSEwA0J
O24aRLpc3cwIfCtp+rfiXcNjhPmslJS11EsAVfrcGtgFk+AoyT+x8ObsKXI/nnZ3ORh4bL53S96L
c0lKcYIsXHi8VvUh8QZyw/QlGjSMYM4cAsi7CFTGmZ06VQjBI2zgQBHDRdyd9+v4/d/b0zU2HHZm
/4rpbPX56m1f7U/vgcTBgMpnMRuFm0KqYhpYAW2tP4EajnQ9WfM/ke3viptZs8rSGF2iVVqDoU5d
5vyS8pcGGVuHnYeDHxdSol1ctPptpt3lAR4Ws+Kc5Ksb306/EkKF7+wtk1igw32M6iUF8/bIRyWX
A0iJzROBgQ2xtzjOdjqe8Csm2g7HPMLo9VVKQA4jZfHzGnwjFXspE38+dWSca/6Hwmy8yMUQET7i
J+qSEeZmQIMVjWluHBbxTpIsbSaILzxk9P86lIwflVVTk9ah2CjBo8aqFDrCxPdXCVqXP3bLbEw/
AbbvvlABDnN40/JyETb0GiI5hoz1VjBGSg/2zvGeYPUuojY1llWCKmxXwnWEPM0bBwhByEDibh0h
b9lYXgP3RcFmrLSQv5Grsd/Lm6DKpnqB+WgE8Q7uvPEXcaZ2iqoE8hVrkP+VrnS/rQC1Scwp6eHi
NcHdbSB8rpk/1KKSyVNift570kfzox/JVlIj7tsJdmr5KST0i6ihn8zT9IimxlxrfSy9IRi9TRJz
LBTAVn8svo021f+HPK8+edbDy6no4YCptdV6rz2QDxng7a021FE3RwiTEOoCEKFu1n5Y1iYQwE44
RiR3JRmgOBI0uMnGhVvkeno/nAaPtHbxuDYXvpbms6wsSkmKX/WOM0AfHy3K/TbV51VWxw+Rupg7
oykCOyGwQA5HRHoIVzMp5Q4DF4HpXDKiz68sqMKUXJs+5rO2K0YJDyanekjKU6HpoNwwLLUhlvN+
tNw9EDR2wmBkIWksU6FP9aqTboZ/VCjMgBS64U5sAqkot+N5CxhHgbe1Lf+wAV7PpPuOfBMEt6Z6
MA8Qbe6myZXwnYwMObwkIzjO+GAyXvhi0mQxKo/Q7reHtrocJi7k0vc5qIql06CGlmTv/l0oNY7B
uFd2NRsCCfpVgrvTI0+gYF+grKkpK3QkKvO6B5kHqSPcCzvHhTjZUunFpM18Wmu2WDUALBHCb1NR
+UjC/ENjOpxolKjRCs8rDP972m8VfnSv4uUQIQ6YzpzvYC6ggTg7PCWMgswWi15LnICxOuEJ5bcB
b4cxfWEYTAVLCbqW1Hd2mA/qDSFsLbv+xH+drew5bQQW/XxtK9cARLB0Cy/RULOv0T3iQFnPN//I
EwFfDbeZejTBB3Kb6LmRKOlAdOAUY4Fvxl8pkSnUuKKS7OZxsQp3XWZVeHCmH3CicZEQmBSfxQ8D
1UrQgQcJsrqZrWD+HpKuU/rSg5YuaC+MhQMSBMUwWt8uaKaY+IJ7QBfmjyfiNHYmPZ6doGqpm+Mw
nFZMxfyBJgsHJT4RF15EBf3x7r/ZBcB/9FSeZAxB5NIma+pFuubT0TQ3jvpv4Q9/LY81JfbpK4iP
bBzQ5rQxXhB7azSmrEPwYSuylFn9PXwJf+oEFyofOQdRG0qhFaio2lIYxlXf7Mf7/8ZTdAcv4pCA
veAzcTpugY1vKxWdfWvT1H0Uh4cHe1y2vGbPK648jyfqyJLNNd8UZOHsQ0wBq5Rg9P4eVx/S1V0M
o3g1CfK+q0qSVJVgDcsAbBjEO/vhl83+GESXuK1otMFVcQFzuEQ4oyr+lEoDSfkGnLEyA5AHqV3G
uUfiYC21gX+02Kg9wHkFdc49t9jOs1HQ4o1N04Z1dlTnrfox8ho1IDagkLwuKC63jzPRus3BFM1s
J/X6k2aJyA5znxHeVht7mc4RNEXXDXwZ+LMEsBh8jqkTMfhKT/UEo/BfDtIztbwvRWvdyEP2VYhS
ON0QKA8ooPhqnoeXyFy7QfQJg9rXZaw2lUq8EQQBIoQsfdTeuLVLzWEYX4SsxmJ49fUCcZQ+qMEc
nNbZ+jZ2s12a0czevGW/74rAiw1Wz85+hddokml7kOW57vls69xB9h+KRJx9p4IRbhK97ZyFbtf4
RzwxtGYA3JPlmq70Tw7yaAAI0qd0F3K8doQ431jWBZjT+XGgimafPfyBB9Ya54FTMK5xGR+V0iGO
JMbXYFm/WGuE1Ig02jCuKv7wVno7y/6qPkD/t+f8+fNMmSGyhtKbzypcgbsYB4mY/jge5GmfGN34
4w4airU9yikjquawICGl8m11e0I4lu32gk+SIHqjKPRjbabMR6a4DtD2Skzlli1xc2itVg/wr5FH
I4l90WPPKFbi5ayYctEm9vaBz3VJ/L/79ExuvSlw8OKSs1PxoUgGFUtwpofLr9AhNzROjxY+DO9k
O1scJOOWDTpGR6Kr6wLhoOooFQ4fSjXqHXKE7HfT9BAhhtmKzJTrr87FbofrIGzj/HsjGK3B+0s7
hAwbC1k++kFqRbnV+lnFew5mVBkp7a3UfgRZCb0QXYKlCgdmXIofIO6Vx2wArYv6tvlWgt5GsFzA
g7FJVjD5LhM0Qm1VKOahgG0g1BNbO2RpfySO+LSNqaMIDkec0hx8ncY/NCg64NfOggRHx5u2Ru4S
CxF4Ct1pOp4DvlihnQ0gi7cLouD5E8WuPO6yac7h4rDj0eMvtazDsKN/MHAhNJw2qtlL4vMjts1F
qLwPMpG9j8sz/OkGa/oybeXams+aaluVOlh+OKwCX1tqs0SbCud4OUahJMScOpZ5FAvhkU/X3UoP
jWfept0YbbRFDnSxXHWJouC5GcFfRaDWRnVklzU0x46a7oqzrh6+QEC/FnrYq08GfFOQKHWyi3X/
N4zbebeneK6loGwV1AOqXEtJAgWRAVBBC1YDBWvIqlPWHP+3Zy4L5fb1j7wpxvhCyOwKtfG73fJb
xKAAOGeQTni1u09cVLHX3zgt8MzwPAjJ6Mpv4xbnM7mww+u3tGCJKKUct3GLX3dA10bWYZWLpG+S
nX/rfa6Q/0ck51q3g9v01XdWLy5FryqOxqZPWQvLwly8tfkHNkGMoAISOnIsg5DWZRed094WrUeM
aPDsEmuPCOiMUgoj0Qlopa9FSOBY3ec5301oGvsQZYTc9o8qk2FkAX26ZyN0RyaSvsxx/vWeljkU
wmwUg7ac619rns1OxqI2ipmXgOaZATkSjiXJ1xU/IEXBcVNrh1D66gnvJYgx4Yvbi8Y/Bw5Y+T16
2iBhVO7jz2PGezWNJJQscfo39BsBCmGghXhweqPWNCB1jo19GSuRBYFQu5v+Qaxm2K8HLVopcUau
PAuxfbxa0+ST2aiec+lH9F163LmN3YgbsU23kBbpmtrCriG45WnL+LDkaojKLJwAPhQTU34zU9V/
sN/ICy1GCQqq1T61Jrl4WQtt1Etxz8GR1iZMaZeaq2NlM4lSKEoHx0Mf6Sj3ewzOoerLGNgD+1FB
RK20VXiGRlpfJB3sDZBAqbtaTsetM2/omaneC2SazoyqJ4Aq4KJ9pDczyseHy6N41VfEAGVU2X9v
RUChBsP4Do9GWS81UiLmfWzJPISDD85V+s53RlKXUJMe4fi6+GtRDDKsrH7EJAwHLU5A2oReoxrS
XW31CG+57UIiqFhFuwr7839JvLq+ex+76/b3KR447zkcgOlSV/F+ci1T85gSSCKi9CKESI13MmBr
b7lhYO/uN15xd8UqtTLLMenHp4zF8FQ29WH46qBPEOnWZXi58l/z+63DbDeqiWy8PXI9JJ5MJ2zy
OXnCuoXhM9MWg21zAIArDXFZeWgH/MzD+GBDrLEXusSs3kYgtUDLe/rGCcrXfoLLwL+hCsgMJuKb
4YKW/93kFyjFIPFVs4ZSqmnXGr3i+m64hX5cvVVOqoz/SH8XsKEJvCjXmPddi05NF8PR/bEJnIj6
MVHgG5qqLhBa/HtoIFyYPxJIYuzUCpKbmVlOwzcNpYxrmnaBJGKBWL4+lrPYYUVeRs9EdN0rQ3P+
ST6rob1cz7RNwlp3diy9LaCRtxo+99NM3Yg6rjepXcTrFyZubTRsnkAleSJ34qAJ6m6rsQrnz3xz
PfGV2K+CGN7ExrGuI8gJ0xfeIkMF3IP9YevxPR50htn4z2SAtFAXeCJojCy6D1zQF9zMCorT6lPy
au1IBvHhup2wXLsOlyoP5nR+bxNX12mr2dAV4FGWxfrpJ/iOhFuL7R3qJ6qcVudgd6+JXSztytuS
sC2GmVIQUuZ6skppIaN2WLszRBpydAyzNChEqlYoxmj0E4fzp6KRLH2SZPOXktO5vcHodmV66Hvt
IW+qOztc8/9zRPWhLBfTMZvyHdDbCB1myzJPzIZt+YMGS3W/6j5u9UXKL/6Avz04S059z2jh8TPu
cXEj1AkgsGD01Twp7IHvXKdzc3lqqXI/sHxdr/WkpBLIkv9ftDeCy6vFPLYp4mUkbEBTB2gO1ri1
vWt/YsZ2v0sgEurJPagZzUexSjTmq9wfRM9YbNcVhO5lNUfd4Ra7nsSb+TkxcAYo9juBuP3+6uEr
NMTQ7Pf2Sd5l0sNVx7YzOjn2xkpkW7EESgCJM+Tt+iST4PjMmv41Alx9nrokSxV2yVL3sdhZFPX5
fAK8TMLj4NvKhcKH3tgjks75LEJ+oheez7W0OZ0hdoMMQFpNH+hayZRhJSr2S7bGgWgO6ZuV3Fgr
T8xWSzfx/aaAUVGNOyYxB5lj1pbVyyILqTHwZ1Fq0afN13Z05AwgVyv5ZpRpWm9tJ6lGWzFwaatQ
lzhzjAXE9nZbFnHN1szuCCXWrjLhcAO2vk7GS22YHitjF3F5pDnHV1LKMpBp4RqyDA6aMKm1XgCC
jkeCtNaysUNauqovUW+TE/ryG8an9nOtf9upWUbhAHtTpaAMr2mcIKtqJlMlzfBmstpSSg7erxma
93XvnknCJag0w65rb8Oeb5gwCYSg1RTtMlfDKoKtXFCd6lMN2PxvF4hI7ftHtu91v7v8n2S53ns/
bF3keC91zMp0nB14XJ+jmA5GBMFMybC8EqB7hGyuESPLidMt1oOwdAkobhFNhvOkGSIr8aXPpJSr
mbJSm4aJq3oyvQT35helFErqalAJhFuOTmDQqU27TFOAGcv+euGbqbc/TbrEEryzRQ2tAFfuVErb
1QH31rCLt7BccITiVB9AWqReIoTz5jeVLoJhUz+Kkgf2lKzB/H+At+t2lH1qWmJikOTVv08vxJZy
RfRHMUEBmKcKtDGEpZhOc2bMvQ9gNp7B1tvWU2SgtjcxKQUilP84QgXtFSMi+ebiMJwWt59n7AY7
w7QU+pSUq25zB5F3gTnskjYtRJRMfCrJo7+yRfuql/xqQPlEnMAhjZRoSNVT800XOvg/KYZboGxF
mbUmXOJ3/+n3IG6CDoAX+iUqnMnYHNYcdsQbdPfWC0A8YseV/Xq/W79KkyKKFW2h9YPq+S+f5Aa2
Fpe/mQ5MjWhwjKFcQqal/tt9HvmZqG9IGvZVcOxgOzsRr3FCCZeFY8HXf5/tDjk2yHX00aQqAsEh
cAoUrAsYmoDESIhyHSM15mbjMgGoS7kxl/C1BiMe53axdcuTUKQISuZuJHW89cHIICXjS7AhfpIw
RxxneNfpOGL3nW/1Sn8Guodm8lmu6ItofrYwffCQbQf8JUCeTqZ64MVInqJecyqyObkiMmo7/qkV
5E744GtfmqlxxfYFElHRHIRmtNA3LkKvwyA6z9XHy5HLBdZ7a2DgxsfU9LadFKVdkaLvFedTV65+
HDhB0+nX9npWvf0GczX4oPEnO/jR8CbhcwvRFGNpFxcFFhN511YYx9EvPulrPnQlZSHpaXhKYyVR
U2ZUGmapL7RVnl+BRzleeuCeFyo8CPMQeYCZMtPOwRkuFjW2qG3UYg6HkQ+2Gt0IT5uijtmyvQoI
+mvqXgKH9M3H5KksaQldax9jnEnTsc2V5iv6sB9wMby9lQp+WY58P4SDGE5PPb3PT2Cw4zGC426H
W3v5t6D+Gd/LeoYmsB36hT16ERJzVISeitP4fnS/gae8vlo2HvlMMAu1z+ZYaS/Jxwoc34wWCEPD
5U7vbE7cHDYIr6JBjqMSxomrSw7KO/v0aMWGrqhuzU6NQbHUN2V1TCt8tV1Fyf5sYH/QpfEQFaVp
9JtQdhpfY1YxwBY/4mAXuz4I4S+0x1i/EGN1tKjtITnqfSA7sfv5CHHMVQD0TJYTtwu7VHpTSd9M
tQQM5sPTRpEm/9NDobKNbkMJlvoIHgShO7EUtZ5gObL8rgpcoFUTdmniMfdV03Ckev2MGbAmvMIt
tn6aWMW94TT4NY/3Xf0l77yQHXV00t9dCCPAPuk7cu59l9PgcxxoCbYKO7IZKwTIsAkHCEyudZb8
E6IcL0KY41Zb2EaTg3esZ7En7VxkQXOIcYpgAdNrm8f6F2Ex4wLAN+t6Tt9WZ0Nmyp+Lor0bF31+
vj6yVnns9e+svntYXBWFwQZp6fxSGzaey+DXb4CJFcQdKD3yAEZcFKGeYzTA5f+MYefCK6nbWl4C
DSxRuQ2Uj7Fjwyq5HUOsHCJDevolJuQTvQg8KSKM8poAUefDf0sfzUQSqcFlNclEML/bUZDz7Fv2
hXUk5H4JhDaz39ayK41FW4yvtiB7gUtjqEHmFPnHXLQnwbax5ZLRtrBCxTxkHqa5ueKIIHiTY4H2
xiyB8nUkM+GfuRg/KKQ5BaRsxnWeXOdKqs2Sk5vQ4lkfOKnxdXilBIPwmGbtTzuYTB8D1+tppJK0
LpPFCqqx1I0qhSDfFNuc9l9JLs6LExX4WZ0wYYEA4jJ2dT0QoGd3x742Q73lhxC1y0vldlIKhfhX
sg8p5vVdRqu9iuQdnnEpbJLTMGsWYPKQ7OmsZ/3TqtNKvE1gCPpKsss6knAedU1fRnoL9B0yJ9bL
7wejxuLRQXLG2omjg0/bovqlTxlb5x0QKB1CmYyxhrGqUjOpPjoeomzpf4tknsb3Wq7WHY5CN59X
Sceh6VlNYfysBvIya7uZgJvT3my0KbvBYRiO4/KSgS76euXF1E4iDRleONbY4q1t3GR2SB06fCtr
JzOSJ6Rx4vMcKOvokaoWJSr9VL4hMFytP7QFTTUi4HMs2l5IKg0q0gZcZve9ufj10KX+eWJGSCBf
jPWutW4cIQFInK0bkILPh8ADWHlhbAsNRU9SLPFHKfuiV4LzC0E5D04VkbtAg9TmJz70WY3KDzcb
YqZUyUgBs6s+9lkyPVYafO91EQTue/hI3QTohEhczX4G2RUbfRYLB4yeybbaQPvrAxtzXLSs7+LJ
LBIyFC4q4D0Gs+7Srh6aITtKpRW+yBn34HR1MLAzVWArBOOGB03c7U67tQiRIOOHCD8xg+7xD2fE
MkRU8p5H1Vm9EYrScO0LBofLkd+6yQF5DrX0nhZ2PZqiJDkJel8gB972PgUvqYkF8OGRrbBtu+UR
BLVLnLQzUtU0P+z64p/p19o6ZSWPrzQN3DkHDVfH71AUaaBunqv+zXa+11k7rH20Qez3J9UeVmPL
wW/leJwUF2Uw4c6X0EBhKHQTK6SB60kmZp8GZkJBNxP8qemAKbOlNBUY40iFlYp+uKKBTgVGPE1x
vG/zJGXvGKSRPzjqBoqO/Gjkoid4vYKL4DTCFH1lqFQ+NnzHj5tEOFhQO1oqE95d938kihc4QOnz
VJ/9PAf5OhpHFw4PjrXr11azIjD1bi3+dl2acsEZ14jGzMdMrtUcNwCVfKT/neRbtktnKEl8nJe5
vVxl5aBX8weiWxJubYzDpoNkTrGWKzmpasDgpPvMY7VHIVhoAZWYvnbIhJ8/eKE61vmeDLDCzHXc
4+mJcoPxN+yxjHlHFmBoXtT0WJdpm+qOkA/E/ZJZBnW1ZoK/DuOcaPfILMWy03B8d74PMpVjeYye
PuRp3SruIx0vygVrBo3xr8a1vlXWISj9aCAFgMGyePp6zQOEIRsYeznG8Q4FVdP/b5YiX1i0kCBB
+cwB6c7dIZXwrjyvpTfydETb23bDOpfATeC2AInxSZubz2oGEOjmsay6WjA/aH9X3KVNvi2Qppa3
jSeLjJDlZ83TorluB73LgBAHAAyc0pSI5WY5H47JMUgnsLgt2nwWcgqi3DYVUhbaE61LOMbpGsdK
YAvAASIckKmwrIOZ8hyCiyXd+8mrFg5x+j1hmmyM37oh2HbGge3DtjUMyEP7Z5Hd7UOJpg1a3cB0
TFVvLtquCZl1XBRXSOKnJ7JbjoEfPaStrfioL05s8GnQjG3IILTIjJIrg48oF2c54TUqMDLGj5tE
npc7xWYSTMCK1pI8zk0fv1bnivTivsrtKaVyoJ5rCSCqxslfP0Zz1rdqF5a8Bj89+e//L+pyBifX
ThgKvxTZowEzdLNiuBCuv/p1lHfMIwaeKdxCruuVqjNHGNQIf+yFnqlgjirfzi2obDGpGQ1gt4h7
j9jp0FOPeTv87DlX/VsJwpcMdn0ulm9WhpxhelvaVpJifNhL5T7rQgMJv0zr+EvbqdyfTBmf9rBT
ovx4Z8wd7caaBVI0mpU9DIQMZa5I4ny7eWc3qlGwGIHe5fPGX5FFz/pbtiskLwTqRNadLaMGhxjy
ejpaY6aZMpmtYNg/rCPTLVJPt4x8XG5f94KtFB1Bidv/T4ywbEWYbEgPq9aA+ZezpEzmhZy2Um1h
5kniNkQNVhuR+mvnWY3s03854OQYFTGEmerfnTmdvZFCCzA9YXgtMXKzfZC/Dkag5h9/cpZbGTwu
ue83vl3fEa8ZlMa/pxCz6+K8pEKQyN2jTr1kJwbXzWdvSwIlnQTasg8yYPLVRR9RGuLFJ2SiALQB
cIzL5Y5STM1KbJwbTEun7yLm+Pz8CezHjQSu8JSGfdVhgOpSv6ZPs5jeQcDYT6RFsSBw8LoRVVA1
a+WAh63UbSBNbvXv80BsbLLm/PGxK6rtzU7qSmRVU3bl7ePa2zJt6scHEDMgCeKHrf1ciLaF+oko
1SIyZcg5Cqmj1/LXbYbGSda0ZGL1EjCfZPYBJuLK5PbW39oi9o0TeZcrENJAvZ/aw2Zkn8YK8bLX
/AnNIXkK3FB3MQQNwURnXU2Osh1u1z3JMG5aRdjYEKJaxUoGQAmMHIVc8r4odEAgm0AVXDI4rWwq
jV5e0NUGPPTRHLOs286hOD0vWRIBrfriSInnoR5j+UnJr/vSRQN0M8lyejKTdaPge+l/T4s0E0PS
WolSY7PnIL19bwzogP7pwZ1Zb5O05zkzoLzVhOqgz9g0Ysss0dzofd4IquPSPOKT23oh44Q1a/5k
9bAuBLj196jYgCyGhiA7Wuk1i6kb19Fk/Wm9dmnH22wxizBFIh4lsvFiM4Ok2LT0NeYb4wkNG1Jm
XtCHTetM7HPOjN2jT4fYl9NhGUcJioAWeY1RhxcDcIDhSOBb/PEUTKBsq9+Vd4kBzewcBXSZiCt7
p0wCjXFKtir+fHNou1ltMO9STWLtj1rhSe94cb2dQM9dlZ6Mfw0xnttsYek5iCHY1R6SK2XLCgmQ
uuMBIiIPxQdxgdtjooXlG+aTkmHLAuuG6Z7As5+u24ocPLDexaJHDT3kUn2R1nWtY+9ROI1y8bsP
4BNGt/+8shUgSBYSXaiIIcDfqFF00JdVUoOsQuMnQ6xTx46B9pxSQ6iMRTgtvppZrZkEwhtLCxUq
9yuB2t/t/bAysEZvZfH5MQT5bi/1qVLV8TFuqEnHsBWEclgPJaI31v+Mbq83Jk9ewNY/ElmOEM1m
ENuGqOrLR91bkiPw1Fgn5cgdKDRRLVoPcZ3T+HNDG3Z68uM35dzdDUP1jensYPZXkhog9necU07f
jjIg3D0WKxNBK3yEr7OujXyd5N5onUi1bjIanpzlJp4Dw4XdHK2DOQDPH11mqC36ILiLG6oJABjz
XgIik9HFcujE0Vk4B1O84+Wmp1oUokfyABt5bBxJdGXlK/UiYmW+HN0nbvq2mrLpGOoDMrgx9/IB
+6li3mWUI7yi16M0pk0bVnTI4DhkNhiVa/Y33PVNr5EqIbsONl5XW37pXWyplnekz7eg069PJw3n
4qC8/O+LIucTJXe6/7iYNGddGalQv+tEdFWkCSWctXPFIMm9hsbH5AgK8h2XYT8nYokpKweVIwhl
TUqVfaD3+GxGcw/EuxkDkQsvIoC2SvrteZUJtJhgf+WlWRe/7W8Y822fBXOzy3VLEhaQlQFPKX4i
iONJVuz5Y6J04FPLkBPj3n1/rjPMQUZJGtGaaIEjCAc13TxKUxzD/0Q5e9Ptc+WnwOiT4hlXA0MH
RPfQ2AfmvXuvfS32avyo2EJnN1hZAU2I+RYgcLjfX9vC+IaHkE8gWzGJyZspjYcLslkn6d0I+Wxg
MreGj4zNoU3uHzfULQlbek9u+1LTzIuEfxIy+TOLWCOXOwSk9eGWbMurLxq20FDRyLpY/PwFDXWs
SDx1cTgA64j2/nxwJcvlCHrLg9Uvf9QGbrkcRF4p9dUM26iN88EDuLPk6FznrzXZr+d5HP0qeECe
+xsH7FkopDE+P7Su6xvb5tMOgplV5rm0ZXFPlY527yj2Fzn/FsU98MzqNE+DfruhKRg8btUlnzvb
29r+AXqyS0Zk8N+k+LlH+/TUcovpD9d8KhNErY3rzyQBss+XJuTcr8fRZMfA3f2h2GiDYqeLqT+z
vZrPQY9RA1FAv7+vR05oSVhPHUIOvgEQlDyXzZuJBGSs7h6hXQquNruFWHUij96vJujQvz2Zc5F2
oGK5oEL53fYUAj58SMLZeVyWNuE9SWYNQZvaBn1VW0LSsz9glSI/x2GdvvFVCBbws2ZT0eXoCRv6
TgWpt9lmIyTahii105TSkvFzbnqVrGhAYsFKXGPT8b5ou50n40nAwuLxpRp/s0+BfW+AnwsPPJjQ
Ux/QGAaRXu38frM5ZIOy/GMsjDfkTBiJZKiBruA+Oi7zNgPRgaw7W/WPi5Bz23oRezjSIQmEku9k
eG081in6jJ22K2w+Cgj7UNmC/PERXoXUq+r2vNMU6GYDaLf1Uj14/N/b5NvatwABNWLFpQDmBaZU
CqGY8TWL4xLiUUD3C2RBXvYXOLjG0+GPF0EoJo92OF8DtB9OHJiRxcx7XJ5ZcQ98BjbkNe6ix0Ph
Z+Bz5KyjchmZGGlJlsWvg6GqH+bB9vI9TI72IE56Sh8rJlSd8AYYHJYiqWd3ZgluP1p7YmrZln+z
y620UaHgv3+0BILto7ZZmvbF5LGsp6kX2Mp+L74JhNlzFwxcBpBT5Z251lzcX5rZsZg+wMgu599I
Hj9brwVW1vmf3qpoXknmwzqj6L0Tpa+xq5L5EFhwJSo9yvYpHWK3eIuF9WZ709LGo87lGr/0g/or
CbPT2bxghq7ZW3ONEHUEPEZdeTUkgChpNeayradltx8PBe58SFq3L4K5AjI+AN4z1tPVtn/6w3TO
l+VPARBtn06jMS/cokqEwkl5H8f6H9OP5/qJLfGV4/7B6sCoj90eEa87V1yosym1JumrdrgDsxVM
JAjU5RF5J0Mq3zS/xn4DVV5qFkkoZMStGpiSMi1lS6Fo18XbLvunKeSuIOcJMOBo+ACT/JNvqRG1
ocjatf1BtLiSWRg4H4guJfiP1938HiX/9dMPU9aT3Havo1quLXIb2hu8buQdxzARVUhmB9h2R7kx
/czXh0Vi5GYaOQmpBm6xYkNmykU2vSrfFPQNwpuNIrybOz9aK9I91JyPwXFAsUAL1J8YvJdIZPWz
LhChM2jqHUYVigkBrifbKYTZDQBGhZTqPfqQzExZKNlTlkbV1ypsSJ3a2htbSeMqlSOLzJw/krvS
vFHRBG5Q2UROj8VHrtutrD7EEx7YCAZAil82loFDs0+11Lxm6a5W2b6Xp3TCEOOHVGEPg+sMEX56
w1dUuh8ilG8fFHsZihUq7KZE709cltlT1RG4Cl6EO435gG80Kju/cLJOrpVFOGEmWuFyJsojh7uz
3wJtqvi3YuoeltXtesPMnVZ4hljMUFINV0+xEnNlsmI7JNU3WizJfaLwK7aUXi7pCBKO5zG58Aki
ztD3w39ckToOO34gCsz3CkEi60H5PqzCXuKm3nW2dC2fwinI06kQh3ROKHrDfEd78sB0QwxX6Ihr
J5W3tSLTtO1ReGcE/JbYgDL2B+Rae+tD0Ivk/u62NhHxi03RM1Tm7ZSrxPDSM2zVV83+QzUlPNZA
jEvDoZX27gi4HOFlFSiiwzUI3x9cRxzJ4z3ckUkqkN8qS53iM6AP/fM1kUW72cmfahOgxmxU2pvV
QM9oyDpck9I/bkFScHzKSc3YxAWqqB/pteq4Uileym2QB0tQvkTs3S1wo8efmW70h1hwcT0MhSmt
BCfH2F6dEeFx2Evu4jz/PPv93AJcns0Dxun600rO9x/yZHO4zEhuDfKJoBGtY9vX6vx/VRVV3RqK
aalYXjvxSttV5pUM5HSH/8bbVFOa9Db7qMBqcq0ALjlrrljc5iuDdwbK86NSklqc1useRgdaTa/e
G70cSbAq8zZOhkaOoY8nXe52N9Xg4oI6LC9GRH05hbkNEgJMwWnGTzpj/UFfDET9WCzUAiNLonGQ
v689tipI11N5RYedg6Zo7FZOjO944BIkeSMTY3MsmWyLaO2pygwPvRXdMforWWPc6MRzVvtNSGi7
hImX3LPSmaArJybH+pyIXXTClTYCnrJJFguG6nFw8DpmUcBgA/T6gHfam9obDd/020lVM+G9oZ1L
id9kFv9ButFp2EQk8pYTPvn6Qlq14sSY3VksLmbEgXQg5YByg++Fntt3MPpZ2L8VKhCUMnOVa2mR
plCWKCXB2uhYqrGAkJB0vtGPE1p1ZaB8Wtm26F0qAvIqtzULXyLPvSZky9Qm+A291HDXcgUJ/7Ss
yQl5pMD2EZFuTztCvEzHIDJPHnSQOu2tVt+BoaWmBbtGcvDkBgPugnYJavpIsSN2mI1VYgYLn1/9
wBUm6Uo3pcaxo/cpapqc+IBup/AYXPciOesYxOGvWSm6sbnobzqWKV/4CPVvoVAJBxp51B0eW+sy
q7i/i+7yh6VMSJ+swM9xXYjFA1SylhCz/TW5raHUVkOGA+M+/dzuwy7AREAtU7bzP/gqurHv6Bqd
oSgTdb8Ad679c22wOwMPvKEGX3rinNBVH5RTzzLyyHfsUBMmVd1YCdW3/yVnX42gigId1bonGHjd
0huzU6fXfIK6wMUHHiN6kfch92dnCB27GKBdm9eWkb1d+y6IOqv++RY9C2V51WJzEwLdJLy7WViN
snIYRiiGVPpruum9wY2pg3vAX7D7hYrw+3StXTepUBbmIK7yKoeTGbNEC+6yuhc77Qg0Eg416SvH
icMY9U9czblWV2gG9VzGn8Y0AAom17zJaso4dbh0zvTLDZEa6Dn+1jZF6xptwCbGHRGN5Id3fq/4
6sUyRFqk3wUEYGvs+AVFZ8EnVODfn3cQCFF+1RitWfK9CSG2a7ySvnRgWKlPLR0oKE06rLR2bj8B
T91a8Q1Vg5AZOmGzI3Tf3K+pZZCEB62jUm5gwKrru0oOmb7SreFuG2wDulxGwZ9qc2+NSkuExlZf
MJiuTveChw2O5Z8p10BTLKUlyroaGrhKxJQmBiXBF4Syjf0yp/uzfCbmXHfsa3w//QtPrm76OuVO
raYSRrhh7vII375yXQsLCINgppsoBK712Lg7IhL/85Tor5pig9OgsTEhkTq5hfOc23nUyX3CbNqs
p0FVEU5HSQ6T7fBGgBI9/sMDUQd0T/sZoF40+er5DOp6879hnRS4g0ijsaiTTnO4KkUU9DmtzfNI
FQodQ//8x0fkpUYKlNclwetEDw6LXhLD5k4RLkhKyF/5rLyjDfL7KGH/9ljyfP6PB/qJI+37hwLN
W/t7ouXd7VUbCdFxlORN3tsooH5jViEQIOcwu/kkSRQjVWGsAElbnOltUaeBgMwgKn3PEN3AYjVi
oCmTXk6MTFpNwGZ7lFwQiemf3GdzwYzFfxowg8M2TpVhjT+y9k3IjMBpOGojoCXaBaZAphPTHjxj
yzxff7VOCEprU5BLVAo5IRkDAxbeXa3SoeUU+zmG7M+QtrxS8WQV2e+GlUf+zApvIhJKW0c1AbnE
wlir5o0v4f9cXab0zo7nX9uDdbf2rl2zBmz+6RxDm5SXdv4PK4KpaE45TJZne1d3uMbnBgPVYOI4
L2VmYpd2LuzO7AAvVlmxcu+rth0mPxd5l/2275j4F6xF7a1vLL8d/C11qdx99Yd7E3oFCxtx6wGL
3j3kFqzDC7cs6IPN+q1rkr5wwCcQBdGNTCaWGNNI1UuexB1CpCYBuzNrDqxRP3pAZPSJDFldnnwP
9KNBWafkOW/jSrRrSK2NN6gxbauiMeQcPiVimR4FB7KbVOzof4rLBN1lmPuzO8JB4LbCY8Sq1C/3
rqfffJEtvMQgWQi1CC+to6AO3zy1BESnTvoO1NKA6x2O8o6bJTq0ZZ7Kv1odi0BlYFqUgDvXMeOQ
UGZC+EPEvfbVkoP/FN0IWVlCC+kDacff0D0BKmZ2otTqD86y+BpoFG8xyUtx22OQvq/WMpId1cbf
JJGt+j1CASgni4Sg+KbePAZKgNal5F4rlw+H0W/37PEGqxy9z4JiZMYFIDBdJWbWSquqtfVRs4MK
Qw0SsjLpwdddKE1vgT7O8pIE6Z0/1IQ0tUR5rr8nm7NbtcpTqHtuv+i1y810DOWcezCLq3f59ihp
S78UyR8ySD8wdVVU/xxwk77qT4buew9v0EJNYMDZh7TcOf0QiqQBHx7S68qIKScknqL6RIOJYoft
QHI/ooLNRfOBfe/Ye4ivz3fH7EhvZPOBU9ViPTaIo7/oY1o4jnodCQJs09T3lngPsHrO8RxK8Nwq
eP4H8nCBw0LfIkQRD5x3xHbmjT7cVWSoPrYwP3Y8JtnpXJDl7K37LZRUrc/CMhOZsjIKCU8Wmwk5
sNVUNBtsj1Yyd3AZf/R/V/92J9FH3xQcqm4EYfyZ8a6Ttri735GpuD+Yvjosv4BsusVclT9Zjwpd
snHtEhKoQDAiGukXjYJef/n8/A2k4PN+fz0RsgKJaYpVM2wRHNOOwkGp3x8DiMK/mA91UgCaqpoJ
JGtsznlpj7vjxFcDl1ZGAnXk4sMa7JdmQJOCQ2ABmaeMOD7zuVBNwlQpHf3bkA+LjREip1gvlrJm
lyv4Ruh2sVXjKfKaFwRtnf2tuselsERRitw96FQEnml7dPQbw3Yth88cg7d9GgycBIPezQFm8va3
S+s5JqN3prRsWt+wVJshu6AjyAnKgV5wqV7+OMGcuM198gEF/3UGpfXi8WM+7110Dh1G7FPQ2qlK
KeRt/D2XYpb4dxWvG7+V83K3F+7inPGqsvExxBPv3hXP4E/YEWmtcJ8CRHQKmn4dN6JqfFDp6BU7
fUe851yBXZXVr+Z6oW8iQjswz3WjDroQn5wSxlFLm9+0wNofExjB+yyeqwZE9q8jGPWPhzrJ1MR5
DRkAsNZSlu/ydZFwQ/tuWZ2jfJnp86dn7+chX8NuUv7GRdZYUQfVAs/BJibyTqrpbTKRr7HLbSsf
a0+TUcUojPdiycuebyF2I96F7ZYRpYs3FuA0KZFb45lpWiTlK71EKrgigtqT6be6B2yXhY0lgU6b
k1q6v4Tl28Lfa029xhSy2XAdwYlklj5rwYarqn7RZh1D34RXtiFugo9DMxlKx0Xp5WQT+HvoRGFO
tZURe+bOOtLLr/bM/4aKMe7yzfyLqvj9n5iwpbYgcp9b/PWZ2f6DZZlZRGm4fDl4unrnb7nVlIeJ
J3o6VjAaK42ekcTYBc1n9GqEIFrfu8frFhjkRYjlyY44oGoJeEeXS1kN0DcapYcIDMyAXz8ZowKg
SRJw/Tkk2rCAIeNJNS2QzyTyfa4iF67BpVD3sct37miZjIcGfisa3kjdX3vRgOWjzkBDYOZjgAdN
AEsagIgXTPxVx+CM4itcAdNIJHOyi4Fvf14b7QSxWLXHf6e0cBcmFKX5gVhZAXcVlNdmlH12Mds/
CyGEzSvisbPgZ4XtQfWqn4F6O97pOWst6joJSUFDEywmY985/8+fINpymi0xiZo3ZYEB5wI72t1e
6RdoI10alIoFqwNHS6wNvb0cfuvhsJwqy70iCYFgIThtBjtl0I7BgGc22kfybPgBr393E7agfgHt
puLKdAm2AAZO7sBrvAn++YuzuK9WLkxE+hFLFj6dznnsWg4k3AVp7jqXhbOUwNmoSzMnqBBT1rZp
Z0GbMTTf2v1KbU6vMG1+FcrXkztr3JpFzSUx5uBKvYimar/RNxUPrltMwuBJyozqYW9Ps+z1X6/3
NOTZXRDa6eB2RAs+v49hCXavUO7wbHnNdDZzdP90ZutXmPxK+FSYTnlLR5D7Shl1ORtqQrYZ9wNO
2nNY8KPU/urc6UDwPUaYPN1kRfNUYohg4jNh052b3EeQN+ol4ZZfNZznP8McieawuTbmgUa5kObR
q0oRf7cqqhp61OdsSfqzsiDTEnEjeDr/+y/Ykf5dMvLHBQhWpnpJwGg5qSTwFjzwS5JoGdH7nhGy
VU+W50jL+R3XvZWJFjBvOfpm+M4k+EMDwoUYHn0mRSex8T4xISuok5GrOMZQ7InOAdj8xIAiqTsa
uBapYWDJOhkzarIREX7Wnrc3a9Szyh32Lbduwr2RBhfBDgAVxN2qO/nK83xl/gaqLjEvqMiAEPYm
mBcxIQ8oIj7Ng6a+Zq3uscuvoIO2/4pdFeajB92Dav/wSVzkiFdxxPWtx3ORDGGlcxALVRADo4Xc
2wOK87x49+08iuJog2trz/id8+Oos844GkNJpjrEBHa2DlC64DmsDLsjzqacnp8plTD4c2JKkS2d
lkcWFFKD3q2Yk9aUVOKNqxkSXRaKFVz3uyGsh9d6E5N3GJ62qbWAhbsrHEzr9z28XEYEJmhbuA4v
dwN5tUrb/UmRYomLOqInnFnfGk+K2mlEmLR5K/QBO1vc8iFizbCkFIuiitWvZac1HR35inUYlrhl
wHPK4W3asEWT93keEgzhdit05Se3b5rL0iRgc5yOpuguwD3f0mS4GERmQOBzurVlK/PJUYtT8aaL
Rm2BT3AFGlkZ2Fzk1OuWOc1eO5tzf2+O+i9ubwVKvuPCupKomgKzBB8LKJV4fzN0zVtiGqFfiOb6
Qh7ZKfM9m1R7cLhq+B3hameBk5iaG2ejNkflrZMaf8Be4CcZnas152HfLsEoYdYXT2jtZqQkVYqq
KMAp+wGeSsxmtTS/Z3MhzXOvlBn0nUwxM80sTH5qjM3SrhRdSxBIXEoTuYomjM/8LRZERGcLZMPi
/zHnKRHrZ7IX2e+ukVvKzw7JQOwSFYRAUPuaF7vhir98BzEEv4UQW1dZmm1O5FjUbGW733dS0XDs
JNok8aBesGz4rBYCCUNBnAtBc25v0bcql9IpjZgW8MZnJSMRelJKSIhG92c6rALE5nPZqnibFpvY
5mXnC5/bBnaf2ZHtiJOWpBTdH3ST47tZxRuDARWpvKIHsPeg+vtEWAHdJnNlKHCYmKt3qx9h2Ne/
//JKpcrCWBQk2LvA/IbyeFgcylRPvlHLBTRMXqhworxsHTt8b1MIhzzjpA9zTQ2XsmFQs0fX9jXt
ti3wTBGMB4E+rh8HhDPSHx+8MlO6BpbM1xw/4eHitGXq3LIzPvsy1cpCH9QgdWIOp8shmjjL5xK+
J2yKxOYEHNw1+BGDEfj82u+HH78qpxD/vtaYhsb174tZiBhbsnf91sfTm5yqizMj1F3lKt4tl7lc
s1hxv6l4mQt/K8ZiZ5mSlPXuVtPIU6kntfPFVyyOEqiCLHfOJJdRRDLziXDa0YPZ9Iyz4PcPfQun
vzsSQ+Gkp1Y/JTrrJv8EwYiFu6/HkWDT3FTO3aCOmEwgjJQjDYIEH+uu224hY+Zs2ZH1SWx5pIuD
dDExnbRbQOGi3XEAcpADR9Ke4zCx1O/+eILmwDF5sZQD4l5/ZbojbQRd+b0I8ulWjAPxKrElSs1y
sfJIasUrC24UKDVfWkcSvOfhfq2TIo9h7kF0NodMJo7PE1byGahAMaEOccTcgAG/cm5giHwxIEvW
uwgadE2i2n/iII2Cjc+1OU87ctrSXUY2w+cSVWHA+KzCkcuUavOJ/BOUY6Z17zaC2SlGsUbgJ4fk
lU3IfOL9gTS/S4N7aan7w8TV1tH8snvzis7/f4BRi2vtlfvQqR7Rt5nfCWRRNamzVRI2uj3LtGjZ
gdoipjtdQYdKgW5F4ob44JBftVQYJ2MjqUFhg/l/VmzQOxiCotoXtU0kLfhyUZiNAyLAOCCeo6s6
Hgzrd/gNaPER6pjA79ZFeOvnrdyZVrCpF4fVIcV0QGOOLuJ2K/vo90F5uA/RGOiNf/+rJ1tyqs2Z
OSRKvqh2er4B+MOpvfDFjHt4Ttr932zGAuia3rS5KBPd+V+BwgCMxgOuE1xjWXKmI2hLFYv/0CS4
W9r+MIg7roa8A65+sM6AqOykBrbeorIQ9T/3lkqjUH9HmOzyesLEJ9KjInhI6cJELzwIK8VbPH/1
EN5d1N3CKfJX+l9FqgZ545Ik24wy6LYJIrQbAiQgUTAupEdzuAm2BWpK/cnZIkNt+VnteCSz+sf/
2H0xPKCkVqQ8LU+h19iABXV18KPhUXvPHXzZSutjBJRuBlbN2RE2cNVeUelolniFYdtW03/tQ5Vt
/vTuRbwspp+v50kmDxFmzTbI51080PsJT0O77NbU9YjGGcsmGAELdWlrhKiEgAbXcxJUoAASl2HH
qJ7cvyg3C9+YXE1z4lKeiGDh1PwshFZkciA4qJd6U2yVmvpBpZWiAyNAlU/BEzozwRr7iQT8kIzh
+l6dMZJv5zc5B3xpJuHkT1PaTnpXv0LVjdN6jkvR1Yy/NVryK7kWW47tlvFVZLEIf7DJHn9rEi/t
euKX7trix14PyWwmbNpvqMZmqo2ZjnbPEaAzjmoJp2eL0oEkqPp3KqidkT3ojNLKLgQs7/h/hGbz
kAeksRUMsvsNffKf8E93YAt7Rmvpr5R7E7IFMwLyKOa3lWjeKpvaSHDH1lVJGdj4kNmYay7DVm3h
OYftH9xagZZL+Sndl95nj8KR82vrJFw4YDsc9id90QbPD3pgtBe4f7F1cOHJxEgVtL0h0l1PQhwW
JYtnMfOvgEWMXrjOiYEq22qSYq66jRrgsMBtYEznR5QX1bkk37xW+FATHHIB/Wgr1k9fFleIH9N7
JjpcNFRZGFCb4J9TjBW7D0P2aeLtLfxhmf9O4/PB37OA8Dn38tIYMkM4ijXEjyM3Tsbg2EUAJZr3
yIi0vpOtNWr9nxBIDw3Rdg/22KhJBG48hDuMV6aqX2zJgUVS4hHyjzN+pxqzzCql4jksGNF6dKtw
E7R/fGLkYDO0pWZ45PsPlDAWGlOsdAA8SGeiebMhivO4KBZrwiDn53Y0hC/sKaXAOhC7W5yEj2YQ
BQLBsvY7mxdSx7Gxr14EUW2IemRmQz9RzrqvVYx+2p9cgkj3GsI5q8kXlfL2Sx28HO3mdNwE+6U5
lygzVDZe2rZ9zsFnTiXG+sLTxURIPbxpurv8v12yzreqfllOUbyMr/sTPn5dBS8g/Rg3hOsFaBHu
X9Dlm/Qt1hvkvbfBEfepX4IaN+oyWTPWHsny804pBIVQlKUDXiowaF4CHWMlsXdmmjQ8gEjyFd26
wIM24NtypT4QqO6EO+dZp6hPDAz0o94eb+e4S/GnUfQF8lTzTy03WtzgyHJIiFsTYql32/zhz0Ew
SIEQhh5GyFjoEWdOBE7mVGVdT5gO+a8EmyHbzOe1Hcmgh7wpa8G3isHCWConFsJ4M7W9p7N4mr9d
bdL0erMaT6sjPV9Trn3PMp837CzN3EIFEUc05yL1dOomYNI20TlgxTL8ZwRRRli9MUnVJ5aG2x6T
Fr8L6mVQ+cvqFEYXNtFm4zXdvWIXHFy0G8JV/3XsfRubeSqwL1VvS1YUEnpCtBqne9M2O2DTK9Ag
wXNqlyKUeUFqVffa7kkw6RGU6gNVLTypKHPh4I7vP96RGpmYf8/UMngulMOV1DB4R8VKXzIgc+1g
/UjWJprtg5CvXIUKOV+Nq4ZXZfS56SPWcRQMLMmDvtEFm4eyhp0Mj1ogwOAemSwTukQKbc2m7DGy
PcwjWRlYM4w/kvj9tkOfHldqtN0wIj25q1rYbrrmYzzUZcuvxh8TtAWfM+8umlvBvB/3haaw1rbX
srypow/Mh4pjirpuZG6ILusT3RkW/VpVoYTR5UqRHxGNKsyHY76VuqNcau7EfBXEY7V2Pm155F9w
ATaOsfWe7+juwDNaMbwTmpjZzsHJ+PIoKXM28K1/pmT2tyHrSZ2kZVuLxwyMpnu3TQVduIynjs3R
oSmsBxca/nYcuRLl3sJoMLNUs/imZ5oyS/RFJjiJeR++7E1bhTtEhhrtOnty7V+jO+p2gih2+0rU
CYLOe3sUfO3hUJKBiU5gIi4jXwVDuT+K7l2FSRkticGo4dwPjd4pxA3z1ZRNqhCDQVKuAYzeceJK
m7kZ+olu+KodvNyVmYk7v7svPIiOXsN9a5jOnIPovKsI1w89bOVi+lX/ZzHagszXXfT1O0Xf2MuN
lYMQGW2zoO7eeN31Rxi7JupNjxL+d83JWn8/Hfeta2+cpndve5SXMvh9GBtsF3nL5pFSv3yuRDwP
I/Cxldb1IaKS5oq2KREmJEVmoF1pEFEQGgHUdo86An6lCftyRB6yEmNNnOLBEIkSIaPBwuSS4t9D
Q6k55y67S68mcgbQId+K7u1xYG8YEXQV0Cfyx7ChufYysngYKEKFUAm50fUzO/jrFrHRnfNp8Z3c
L//e0vfxMKkVemNk87wQ77r1cwLOC26OnanRarHVl/kOLSwpKtDCUG/RuWMGVRje17vUx04A/b7/
a9++CXyRJH6zaUUyJK51tEsiy7tvdKEE29KFie1BmK8rjvGpfUYJFotmZkN4kPJQje7vW2TbwxsK
Wfs5YjTg3v3abubXsmeVhmL0NN6j40D1NkktvjBkKc/3fuiJVGdGJiYZ2zMs7CTbSrn2l2JzLKlT
CPBSWIePHDdlv4UmbAc9VvudPhqw8a8Lc4m3YfMHV0VqaiWUA6AbcHMTsGPeD6jMKuT/1tWkvDzZ
2bl7Hh+clPpkrUAxxll0OO1y8zEq2fikuBj5vgJZU1kVDl8l5VyiqfAIJf8bJpTtJLtBofEpkFTw
fUOqz1U5BE2D1y5+cfKwGx8zOvAWW9rkvxpuCfA5ms3Z1OWWGzCvHJ5Xrl3EYcYJHkY4gc1tS2Al
gMqqwhfBDvKZGm8CfiehJKPEeD+/uWJzZ36JIYbjPtw18s2f6N+Q0l6F8kaG6EFpTAKqZlGHsNnI
O4wXzq20/qqvBpy25uxt2BOUEq8To5Y69sAkwRmqbO7p5eCdnTcCajrruouaGb6mgNumFF0SUTO1
mIjYue8GRluaYN6X2scgnRAkjNgPIWnb2LrmoAZ2GUPFTa42avOKiYaItAnFk6e7I3ge6TAWNNlD
9dosIU13xr1Hn3miKsd4IaTvQpaEcGzAkrzYzs+kSV7sVY8rFq5q/b06KPn5sqmM0tj8aVeTwMzD
px2bgRWAcEuAw70UraUn3+GnvlouE9jBURiMbX+qFC6wzr2QsSxkQMKbD6vF+5+A8iHb1/5z+Ga5
HSSLBWrEM4wg3nM+FFCY1nWruuof+1cbAjXarRr2OFTZJSua9XnPzpHVvgf6u5j/SLjzukJUtgB3
3P2hlr3ZH2APmhpZV4Xgjci6lM919POOJMA1/PAmfeddKrggKSb3Mw6tK2LrUq8bDCMirpXur+gL
gsd56/2avduov5yN1n2FOzuXlltu97TukoED5dqrS/Sgg3k+n1Ku6CmJgcY7iYvdnQssgyedm7XE
UsInQS9Fkm3WUjgrFcrSi+/yxsmvnhqWF9ahMWdZwemKYXmW7dLEe8MHpWFceJbmxSErIfVH/W/T
HqzcJfFhw5JvyQrClD6jFMkuRcsU3HpTLPS4tV8hH/tKqSgNA4tQcPcc1Wzp5kO1S0sJ3Q3Ngv2G
CM1yzhySw2G4P5zIdcDSyFYZM4IPki3LTLlVs5Cx0J8F9m1bcvBTRiSL4Xtl24pPkvWDcvBRQBNx
jdGTnRAMVjUk/XT/hkhof7ZQAnanQuFv8pjStuEmG6djmgwogOPZeW85zfXAasJ+Q/Zui2nfeKeb
lH0TDOY7PV8WhMhqn7JkdUgE5bZ4UPM/KhpO/CpN/LuKwtukjbBrv6Cj+lIL9ywGLO8EmBDJMs1e
Fk92gVuvvGVsWB2xDCR5RPuNWpOpwtfT3Le2LZPoyyhSoldu1G4MMRoErbhoZXa06rmeZIAtAj6O
z9VWzkyq4FUnFJmIoIKp+vCHwza7wl4ztDrDMCgVPMBeUV0f7E2MbvWB3egXTki5mMi/g2Rh4YLD
1UVvSt1G9UKi41ThyxA5+adsIM3+8Rw2IcDDKpQwY6N9BvteGP/agj9tXtPcapnU+0vlPT29Na6v
8HplvpOKXzR3TlZSY/Fvi4UmIbVZX1yADWNaq+2WUkbC9US0ZuzShq2WEiSER2MilNE2BYwAWRAc
nBkshtIZn8DRTVefCB5/UY/3WXrwKgCzlLSQi72l//GlOoVPt2gbXE4NS+QwVNPIOKGw3/3fSHQf
riOw+VcJEVyvqwgUDV4b0QLYzcKn6qXyaTyUIdtu2W7UoZ5nvgjA5Dgp80lrF5f7pxlv3PPRdlxV
hv5tQsL8ysAqrlzgvtPMu/OjyqHBNKJdERLXCY9R2ksbElook3zkrmnPxAl+Adh+2MLS2F8CzixA
HTWdy6B+ixESRJT/ufSthdEj3/Kx+CcoXIdmwcbir/iUqcQZ7wVNj3jTlf1z5Pf5dzOF0tD6bftL
h8lbq5DfJlFi2XBuSXE2GcwvIgRijDlSY3C9tJ9BWM8Pc+EskmZQ/4GKfqxIYQlw8tyAPPKmoC1A
ROUfPmtmsk/vUFfUL4YNYHe2Eanbk9dRVeoFf5dlpf9xWNTetnqnvvVKLwP4zKWsm9uGVtIOObnj
cWwl6ZmC28shcP54x2FuUwhw1iaZnCO80iz4Xap/0L/+MFFM+8UFpzZu9vIzuxUYwV8LhViZvh+6
XMYYym8F5ymEhBVAEcAxDW37oKJjOOmc1AYgOVt/44YU1CK72YD1iP4CGAzcXPkler94Uxg7CFQb
wZqQxmbzfpR65ELflBn9KBV3r1Mj3mArnCWxck5D3Z9z0GmojXils4LmMu71bB6db7ZSF2cI9i88
YBR4xXca/kxLhLPvBgfZaEmFapI1kuUyVqyToKno44xYhVHTEVxQt7Kcwq0OhU+U5PzxGa1LchKH
ryXsfDE8wO3vwwK7RfGahwM5nSsoWlzkPDxDRz3nFqoOkyZUj8dC9LGKyUf22uRFfATbvlE4690x
lGnqYZeNE/KgyXS9ITCYc4T7YcIkRpBD0BbIYHSxlRRTDUWRUZJ5RqGiP5tBqO1Q7OGMn4R1GOql
4xERc2oIKmTQNA8OWVtsGBJbMsiu+XUu2MfnjFYpF2unEc2K5muIin+HNHU4q0V3m00ELCebTblO
F2aS4vnLRaftmDjAJ822AiqO0ebLVtEloaMUZCDZTpw7oFioISennyR+vRopGw9HSFXtTofl4pVT
5YGzzQwDlVLMQIaGIsi36WunIT4O/dgcmttYcGT9Lar7XpVKx5dnid3JNSbvg3KRiVq3rwFEG9pl
Rv7vrYsCnzAVYezGhCW6ck7nkj+ARYQb0Ph1P7HBbpcITWo+dPeOGEjT56gg4EIVa1wDMU+Oc/Tb
KbMRYFax64qE+TYt2V5hx/7+ft8Vvkyr93jRLL0n6R52Fsb2RJ7AadsLBsRw7UROqbbBSV2kttC+
RUjp/pEe8lt3p6wavt5zvkj9aZ+aUAGGo72F6oRW123CZB7quVbSWQ6pjjBZkfJE5DZ0cN2URCeC
iXh/Ce4EdWpfHX8HdhzQXTlPikvhLX49oEwKEm/FQgKpAgnFCXuqvJcovUw3lY/kq6JVB/Oaycyp
8N6N+N8qUo/DL/8IFCLHoypgbyFWHPp+xOcgHCHswHSBQhTnXI3II19VT9pFIpcYh9NmU+jHPK2m
wIn5QSCq29oYrml6MAj2wTrt6yHWfj6G29qe0QLR0TtnN2vgu5uVOEC37yLmmAINKuyVe4CyaBqB
uxBOIUkX2uNwFlVmK5n6oSUQdpA3ukvbSlAZTTaoIzB68ApA9vtcNrPNa0/yRrjBt2KerZKMVCFz
4ynb7l4WsZp+envfL5fbeLl/lFR4KU/Hw12XRHQZVIe63BZ+GLoMfa6kMYtQK2Q7ZHj3UY6R9zRr
JELPny4Xp6QF/H/tNNiyPtjxb0Q1KqhzzZQnVP5r2+Ajg/nG+3odOFm90pqEk/wOUllX8uMkEg+g
vNS9xZohhYAz3l5IXCvQUumtR4ufnPs7gdUcFqYevRldQ3+GiVRyWdIG/yNd8uesXxo4Oe5k4jHT
5NePMBMj2nc966UHG9K8hhIeSUARsF0nW9acQMoF8Cc5gAtf1EhLkRKcUylePnRzw482ZbtkzYaR
P+O+mJ+r/5wYTuJPSRfhUfoqNaxtbsB47Tl+0HfVIBFGf4UCZ5s8sgUjK+JIOjEa1zM5QvK0U3MX
fMFUcjyPG5ia6wDTZUophABmufoyesz/8+nk0SCoXIwjYaQr00+oaJqANtcEBVXyOo7fr8ra0tsC
3Xh5Ja5Dn2hRIHfrOOIqYXQ2X53JM0cOWozf4WFHh3fCbnu2O3JGXrM7YuJaSa4G14mWcPLU5SoJ
mf4W1p+HNTsLd2Ie782WGDvAVxRyZvBncNF9pW5t2CYenZGBOm2GlNtENAdNV3IbyIN+R6WXjC6n
qmr81aX3/P5dG8a3UbKsMOMNU8l6RwRd0jDR7lVfrG54O1L8vJgqP75+pLp6YaBDv9/YCL+xIFgf
LE0SOiCvl9ftKeypDol4Mti8GippNghC8cTLUqUraoe09DT3thWC6ZputrLLlHtPwquf6urbJ88J
QrB/FffEQPEpzj/JyJ4zOoPJJ8AQHwEz7JTCmaWhviG7EK9oqhPrEcssVP50hixeAXOWbjUs9HjV
Qy9RZVZlbu8VXL2mxsyR/dWd7yEzIsutD64LDRfjI1pva1512cee1iKHQ76xX+GVdxqN2pRKPVEH
2MT0UwbdiIXo2M68uRoqJyxgYNZB1b3HBX7OZaJFGDaa6QWfOv7VlTN7wyl1Cqz3c8flOgwChh7e
I+Jf3vMK19IEgpCvGtMwCAr7e5qOymJDEnnKJWon0b7LPyb4TG4hPOdn6uqv5+f2SfPqqj5x3paJ
+mJMT6YRl9cY8tFvYQb3ahAKTcxIjjW01L5bsWzx4PIbxroPe1rSPN8xqBidk2wYuPwXbfbkr/l8
MLqr6fVj5j7RO7idCMNVZvSfC7sA8SRYSJzmXi8PKg3Kjwp5gjw7DKaG+ec1enA7s/TxBm+t4eSD
cyE1bw+kCoESiDtk6Q+W7/suEyXTCzz3UAXrmpEZ7056Vvg17rkm5sBd3JpgyDnVd26YnaDs06b/
VEbC21cKd0nMqCrpNWIpjDCGDLlWxPrSqbFqEaz54bBdSpiiIpDWojdh/rfRPX0qkZBZkiZlXbbv
2hBzmL+I1vJ+EU1p/pY/ePMHsRQGOBHAnJhzyfPU8IQQjAX+OoLenr+7mQNx4U4KLcREvtGQidhS
wsVd0wHYmXxJMKLKqUKzhIe8PmF4cqFHDWzqAQdzPU/0uYCQs6l7ZJ/S6eH9gIU1O0ST+uqwaCMa
1XOHj87OntN17sKhx1XAhJsbqC0Keh/WFFux6K74UH851pyFHP7EUWZ8x7RsLT8eubWao4O3ba2z
ZmFdkav91iI4uYsd19mXzlP007khNvqKiLB0tKZBcyJOCRCx7nDoBvqPMUMgRT4dRXoZSBI5kCWb
Ft0mzoRkjIRrZ0KfoCCap5DqZkdPXNMGAB5ciZ6/pKWCLZXUxWAzdTnRsc7ysG9TpPNWMlyzXUzr
GxDisjOkzTSw+bxZO5mltjgoxscLp4IO8MeXul6XMVhmsJ4N2+0oAfGdknNM2Ntk6nWvpkv4VYuo
uiEflcktbFQYdwZNOrMS8JGQ50nIm0n1Y4INQvMrI4C2tBPjwuEOuJ6aNZyP9igJ+YeknLtvxt+x
Q76NmJMEmy6ditojlqBPN7KTxoLV4ucbz7UYHK8ojEfvAJ6mJd30fv3xpHzLh28FtTF31ITL7uCB
T+GfUyKX63du9k+/m4+WHZgF4aQSBKXR1TW39hFCWNWP4J71GFI8vBeScKhosudtfBydQ4gB6Zyh
dwYBnYy/RFxQ2pS/sW9/exTbAhRVqSYucHLmnLunLImNxc45INFdQf9pwNWhbi1+hasLElQUG5rN
HFK30/hVcd+IjBEGsHdVTdtRBm05cjmD9XQoOBHEYQnXQTwlbkaQOTlXleYrqpehWd/snrG3fo1u
wBmbVROVem5YsonDE0owk56dpy+zBtPSP28jfk7KPWtnJorb59cRpbX/rTJKZe/2vr37IS8EkswK
gc79XMAaFUotBPwDr8LBleJ+eNOGpLS1xSDY2amtVBtDUUyWizMLw4sjzOqGi2HjS/k4ISRg2zyr
JuD9n/LGLV5OzPpdFvUZ31uqL30d1zwC7eI7AoiwUwm4cMxCsPx/dJ8SmDBJ+O8IYjJx/RvobGb1
YY3iZxASEqdPfUpa9MkXHbe2fJwRPsG5OYLcP8W93na5+sOf0zLu94qSeg+MUrIi9iXrFlpBHQJT
WMiIlFyQ8CupVtnmQbyIlG8Jztlm6Frz8TElAe7zWOqL4z/Z6cczIux1qxCcMtuQrbCqF1K9JSaP
96C2b1XhOmbCkoQ2Exz1Jn1pQKyoNJtbCTNIvQdGmh9g4AIM6MDbPpLd3HIrCDE8Yiot76snzM1o
XBEVAON9+1+OsJFEi6wjY70NepMJ26ciH861yesKIHMLcaJ1clyzp8TGKuwMTrJt/BKExiScXzaJ
R/QBlUdj42rcynrocQzWV9EqK5eqjjTCYAjibvpyWYC3ZY1Htdo1aOMMZ+jWdQ9D0YB+FR0srXfR
VmNBrLXQZ+mdSIGXHFRUSrcLEB7AT9bdPDhBCs7+80x68Khx++upuZG466pfuZtOVe8c7FFpo5Ab
S3hd1lDBDc7Dx6C4v96UM/T3F0lJNFMiYbsIc2wNya+ExPG73Ul04YLmR9C8dh7w8J7m1QxgFA0B
JizyFX9bg7FS6qTJ02qw7sZdmcODhfSFy/En9v/TdSXm4Q91PJF/h+RUKL0xtyaC+VtsYl543YWy
/Tx50QYZXmyR5woZQDlelifArCQKt2dlXjAvJzEQAgEsKHywJF3hbJnqKFe5tmyL7pwjYe8EKaxE
4Ml+jEv6Qi8vFXG2DPdpiF6Wvngehn81rwM2iYnJDmoSRwUFJvFSZ8kVC6gCrU/XdLXbd3XroaCW
UZIU7jCqFcqgvqlmVw0zYElWt6NFPtxv5RLpfoKkC3yVQ6QzBJCj1yS704KqqC0yzOapNyRUMjE+
QDYieAH5euKlqWq0vq1XbEEmodXP3wqCs0aagS9ik3OfmnKBp5kgLVpfPQ1tYn4xULvxsn9Rieca
ZmkG+sGh9jWHRn68LV4r8r+/79zO8yCTOOIY3R191GrSL43b+p/TVmZj0N/8bDAIBRTRBsMYiklc
qAkbjmrma0fA3qSX32FVSDIhuKXzBTvn3iPZgeRdiDXyvwpqALmv5c+KdV59g9TminCNX7Av2AM5
Dlqp5YjwycrZrz5rpJMZqjq8Ba6ph+vXlKeCVxhBxk4zeWw98z+v0A/bTtvuf9uuX4/JbGFMoLFK
8WoedtU3qxlL5q2TJTLO6oXk2k4RU/00SETxrUty9whwzJVo5TpGoivWJUv1z28sGLUhAVpf5Ccf
Fw5JW7zICI9MJvnB6RIhknlcLmGc5Nd3hFqz0Mqx4pkFH0it+9ERQpNOXla+JJpJnU5S8z8GCiuM
z0IsvRJ9l94dwxJRKW+UpsJncaiRG4m+Pv0vGk/NHlem9PQWpY7u2id+eEzYxYOKOx77tgAqFvkJ
zVq5CRKuzD47MKNIfgcgv+3I7q3u5ZawuzN0l0qjX8aTCtkf+EikkHmW++XnH7DmStc4xrA1eNSQ
GldLhvhDxkwCz4wcnFvyYiofwlCReNK2pm5QJWIg7vXC6ruT8hm9OiYm+nLm10tm9fAsq3ZjP+Cl
cMqNnYnSXhahlgAIud8r0BxEl9RgqB9yPatSGvztVWvqaU2fzBh+z+dp/A4QmvgYFBSi031UBNc3
W94QuUf3Dwvj+0YR+OGkgjlPi5Igcf08YzlId0BXhcEUjw1h4WdI+Jl9z+mS84pHqfr1CeopBEGi
/GVwrzH14Ke86j4NAHWewCRYwCTyJGtZJE3ovNtu2ah5gwEb2mzfu9ZZsHmH6Aj5+/IIqwD7etUn
yt0jUvgE67Bqa3nQS+OMr/VzQY3PBFgc/oMS7ZDmLhdi8zwMAsf08LdMlTTfSdXx0Hkjvl00QjdB
wIqpRJ73pwbzb4cR0AHioyI3fTDucE/4lZ16LRxlytLXDdcPdsNqRSFj/vG0bC1aMyny7px/3qBu
T718PRmPXd8tLJHnt03J1wqhi2PXy9tkzfRJoVToNq3rY1EVyL3GnsjGRtQlUgAlfYc1dY6PydBB
rong97yrSnXC2x5hHyGYjinZVyLw9wXpQhFmRaD23EeYX0F2zU6G3Qkjs7BY27J60oC6h6ZAoIdL
DrfxH2te4rISo60fktfyVJrJ814a4DYVHulNbKEcbX97RgA6CqemeIgQ1el0E2IoslY6k/g+Kd4Q
A6PLdSTeygs29vXFrZIB/yWnpCgOgFbyU/xdl5gOvPhJO1irtdCn9PTSW4mnweaQTjuaL17nn+Bh
NFYrWPZfAju+LrGWIHlXfRFr6hAwD9BymL0jEsXW6J+6wrN3cVqr0dbtjV+7hs/1fYEKoowtFMA+
6XlObV3jeJAJyiYdTj9l2v5EdtzlvrTzMd2JqXAn/ebQBv+RncbM210aqnBIMzxD7r+ZQjM7+HQo
1b6aJdYxy6nlMT5cgtACN3cGZMIJ68Oqe52Ujwq0yb+QYp0sIDkEOWXrBx5zoDHGkxRZ3cOswZ5w
27tjkBBXt/4nMiHPKfOeeuApAJHEzew9HfxEFiU9AbEBTVu3nc6vyy4un/THO0/uWiVvAdVGLuUR
nszOoeC9JLcx5Kx+S0zRe6zBlhwHjTdxra4ZCRd2TkKLWD9TeoaDu8dEqh1xBdLu0+8+u2kNcJ1B
PHixj++Byi676YY6ciVHT1XzMttpToT/B38YVWbkjnxuBTCz87aEInsusb4A2YDun4hXBCP+ysu2
qRWdgRD4Mv/H7lJ+yFUg3j+IysUFP42rk/pzw5SHkTxTTCBAI6PFMntF1S33IxCwlCz1yCE8Aefo
Da2+JSZPi50zb7V0ijJCjM+YhpQ+9kYmk9mIml6rg1PBlYWQYqnSMyUbJwGLrlwLKL3Gs8hYT8RO
DM7VjcPBJO0twJ6e0clKFAJJpsDSU2x9x069mIhYVCKIdxCuPzzil0jR/iyl52C7QKke6fA/rOyi
xZJKatV0G8b/zy/U/tjWFPOkw3LLJpvyuZ9lgu7jWVXaP2dqeEExz7Po4+sTL7+r0wLMFNnBZMWP
QXdiKSWFMyfR4THys03tvkxiJyqCZi7EeWVXnumcM4PZuOJpe1HlXEbRuCNHA5Vb2OGNiSNDLSH0
syDPcngK71uhOYMyxDghnSQsD0A/LX3ulmEzDK78B2z+vrHrdq04zPod6AraUIhzrP/MD4dXeDQK
kYJNgSVoaaNd+JJVKCz5mULxhEi7eusplBwWhbjuW47opikULnTj6g6sBqtk7Ho56XfLRX03rxVv
VzP/2AySgLYhl+7x9jMEjIQXb4v7pn7ke9pHJXwAEg5WoQoDj6ZYK2fLIAK8rH8NVaGpv4RgcAu3
4v+Mn3ec98wSHy/cXL39T2cONnn8573I4ZofoqVQz82YORN9Uy14HGoiSA5HS+cM37HkTT9ImUrZ
1B0BFksThR6EgFhRWtSHwQyUhmlPpl4h7vMJqENQyqtT4kuAzjp5MrVFnRscMYTI4UImFjW/fl4U
WKlV7DvdT17W2l0MdNErQHtXibKkXRJWvSvvXQc/yhFjCcbmmWb70CEgJXfo/W3jc63NsuQVkc4n
2He7xKUOtuQeiHHFs1M1Ktasbz1H1He9zo8TAKzl/ECriZfplrUAb0KkJQ7NkawTrkvqPUMaqtB/
urAv/qXnDbDwaSNRvycf2K92SPo7h1cF66sXEPqkDxqVhFACNAhGDXSUgey0EuGFsqsYOShYMCLp
pmJ+60XnRkzJXWOHTcnGkn7+8P6KqbCYq5r9wE3MVYiur3uZuGXJFg1fmkUSE+gRq5rWROvTRtNc
/vz1GISCdjxz6lPEwYr+TiC/B8NqmBCtffIlTYZChSd284EgE2jokiYmw3u0o+4Rn8r99NnxAGJP
GtWVlpOBrSIKhxiYCHpijoWcMh6UaxNWHw0d75I6MF2eLTxCvGb8vF4EWpcKyrjuB8uvGpdWxsSK
xUB+maLsWTRhTYJ801eEVhooq7GzNt4SLFvTQ1U6ACqBmJ9YF/VBjbmZtaDSysEaWTmDGTDlBto3
r+b1XvN8iEY/PkK7N9kRus0GWsKR6Bf+V5zPHhhUrE2NEdJhR4yziWHAz02ZVTjUPdn7tzmfSUsw
OOZFE7JikwrSbu8FUVHQTONV1KNLiQBsbyUxGYbbLHjAqXLZvDPXuqvwQn1/iVQ1dbXkdFkdW+S4
30lGYabs6/r4OtE0D8HKSbmR62G9DqyitckuRwU2jwF2JwAeSoIgyqJ4VySymx2Qn6AKc+v6W5GY
FNMraR9vKDurpfE3TZp4qgNTP6EbOLfuuUs9ZUOtrD3pAZhs4TXD/cHGRikg5mbgkW9L2vMTpgjL
mamlCi6PxKq+Q/ZEUgPk9OPW61O07+EE6TQZM+4GtSlI/SqmxoR/kDvFk6xeoJKvq39J4tv9vy09
Jy4p6zC90jkrOZWL5A9wzZy+66n1PPJjpkAGaBoKNM1P8YRP9EvgZgecT1HcKyj2QIcGfbdSPVRp
30r3okRT8yzzvuSApc7RJTdcYhcb65RxOguiLGfy4Zx4V0FJgUfS3fJNjJ7vp3SRTbQCkyBnbbE2
od5Q1PPpbvyE3gom/mgbd8KQSmYbsUhI3sUPSTg1OkI95C29ZuVoXSMVOMWAoSy8YVs+7ZXU1bFh
L4kqV9qg57JQpSxC7W/+p6sHLIBnsYaWbsiFb0pHJqszwUxcJCpramDlnynaGogD0bRZnsxPrDDB
tCOx7EfFpUImBhOh9LUpJY07OSo3L3kJcY0J7ELnbF2Azjs1UUXyR9z2TVdAQMx3yv2pr02m5srA
WQFFu+JI3Zgzcp0opPys3AAi3yU9k9F7owThsxPih2i59sz7UasQtKkKVwZ6Arbi0pm3491xUPIP
w/7Gj1vflQmiMQypAMBIoyFjhmAmHb+h8EjjJTTEVXVJ5cfbOQps5q3UMbWhxTV5Jzz3V6dGw7cU
ffM4+ZpTOxms1KhHB5mR4EgN2t8FxrEm7pCoerrETLM0NmH+kbOpin6bODzA3hQRQ3YcTX4a/Gm5
qj5F2gLAni9tLCLtuf/jS4FW4GtmeN3QN0L+tQssZoWxfCDBcpwDGARBoJd36oBCJipE7RQMr9g/
tmAihQRrJCXtSzXXah5Gq2ZFm5ZOYw9iP8FRxIHN6WVm4C9eqEt+MpfWNPWUOoIV0I76bS6qJ1DO
BYrYkiUkbsI/mGa0++ASJARU95gNZuiELxkkyazsaG0VlTgPZPtacyvW1yFJNfkvB21/NTfJ561R
56d8wIFbtrM7AVPyE31tSJScKsbmwBslWqpcZ59sJsSTDTU7UsE+ZGgObfQpzgZPUuYY6XUr8wK+
Z2fh0ksqgBk04ho32VDWNuX4nUYR5iqwlnZrhVxOjVgZLYO4aDgfuAbZ/8UzFRcDdr21GU68hGKM
SDWgT8C//OQrnDTD3LvrcTLKp2ylGo1+vgcTSx2wZgfMxLqYnld7NOC+r5zuFU+liqcUGgX4GL25
QtuiT4mjYNLwCG7PYbJRKG3IJ5V/8Fq8Q7pBBtoFvtyOOgufhOyBLApVFFnRZ8FrbCV0xaamquXL
BrG9if5chIlXhCWRMVV9/8ZFEoQMkkNhbd7GcWTkVNGzmSbPKXjqZmopTa5mDlDpL9LkDVV3WNUv
2kX7kLfpDOUEeMBN/L5gycRurlv57v/eQ0s6EgQwEI2vuEl/NprI/tIqiEbEK+iYtHuxHv7M9TVR
z+ConRdP++0D3JRggS4vXXz69zqexj+JuC1B01R8s4JgQ7XfwAgDdXtfN9QciUxy8NJ9DI5uN7S4
TPtPdD+AKnZ0ubAoW15DTyOE/sGKY/BK/2wbfvb7s1DZKlXJUNBTP23nlv4lEWEwc60LPL9y8qGe
/R9RHGdGPoTmNxwUrRTtS50d6vVjEKHR+/37kTZTsNvTnt6/1NpTHCkvMRngdfFA0s0vNahwURi6
c3hVZyJbF+qlQINuL70s8e61iYewEcOm0WkmVgOT1KHP4vjObnvs52uOi7G9TldP+5DmZ709M7fQ
9PK0aFClrnC+0mWdLJsdjaYeC6ywyxw4Umc20HO7JagQzZp9AMgGqPPgyQ5s3FZyL3lEc93ZWCsR
oNFj7DracZuiikGak2AcxUUBm+Kw4FRxUv/bXbLneaQSgVD4+9C2r51kenoqji/QKsQT8Nf1sSE5
aumxKsey5E5rmOSOG4RJWK3Fvy9ENzE1kE1DqTgcNGLW8qMJX3fxYThM2P/Mpy1j3C4X2zSTcwk3
8G0e5a/ZohI8gXGTqXVAuoN1oRKFpA1tIlXXgtWQaU9QPIFe+JTOjNmP++u0Gk+Kj2oZhuBX5Lmi
jmfh5qHwW4gFIYt0xPvL4sgHJXRoiW4cUvbxYkYJX3ErIYTyR/IMfOFogCb39aWl0C0LtY1KhXMC
me+qIvDOyeWhr+b5Om4j0sR7vfl8tEClqaeJfua/tbC2Bry0hVPNIAztYWndpiLxhEYsiP6AO792
KN11JuXBn7qWfEw1wWfXs2M5pk0zL2YJ+nQf1Sg7p+VMOOPPoy/XRoCO16+2C6iCwQ1cgbIlOpk5
77Mbca8ny76z0vOiSs5w3MLpa776PfO4lOWZSK1rN6+QdBTwvON44jkx0D87FdosVl36fZOZzFDW
rlNj29tjN2GmehyJvJbd021U/SuCW8x4UDRpH56nrxOOmBMOAsrFVcwq7dTIdznJskzwlYbCKkrS
mdWNt6P5NFzYdXT7IplCdodX5QWEyqgOmXC2qFv6stLuvxXeLa3xEp6S009jYgzyne2CocD6yq/e
iLdc3VPcoWTyDtagYFP42kV9Y8cH+gYAYy4hA8efrTpCoFi4gIVy8JFQAJiHxw0fpeKmwJmzPIaB
IhI08q0Al7Ltkf14LpyEyN3V7ijHyAL9qyteM0Qo0fP3on4kFtfchgIZDgpO7HMXPRIoNGUNEXAm
x/nCUPqopgFeb9z0uHOpPDOdBGZsF+3Hi5lKy5L1nrLKJcydiNh3In9cLK8T/JkSuWbUA1PQ0Wna
iqazg4DIZYq9LEDN00wGUWsRBgzcGnb+LUpptAIcvian+nDEEjGMAdZvEFnbIG0Dh+Xn5wwS0UA6
yxTcc7RXPbKMFsOOuof5/ux8hv8/d6Sz9yLomTqCNbZVN91gE26w4ZzI0tHyHAQ2qqBQV1U4BW7L
QqAMH3Repdc9pczib87mAGVs9MyXvyIv1REHDLT8ezOfEEow6sY6MXrzkei0lM42yq7nLUdbIKKS
aILxXDRGPl7ZLIIJYoAWjeTJ/4rLFgSLzw26OLQfgG43jF6Vhrp8W4pEHMhytleqrj9WvbCnwtef
xpgk3L0WnGPuod1E4YX2Td/mvzjI2P1ezELq1ehJSIcg2buL64coetKIPTXJGr76daSgOGKkpwhW
G64szUOWbhHW0ElswmQWqxSO32N1SW7mbmlsv/evvykR27qTNXdRlEkkQ3z15P7FRjwuRWpcPmUK
UZwGquWx/2TvPQWkXElqRDNmU/kp/D7DTJrZnb9lvl8z+OuTODirF8HTgM5cD+K4HgWV9CRq6IG4
XQn9hXikI6oeKkpkDcSaK7mCQShX/jLKrZFYMiLOf7oZW3Rcjl9hQkQmDyXLI1anFPHS/3bBNMrP
qvJvAI0lIm1DQeM/QUQn7GpoeaaHvx/DFISV+8QYMTXbKrT9YIIpbFn1c5b6YjF4eEUmZy6V7qGz
m1jsMXYbOlPymQDRExl540MCykMdZ4QZgwSmhgz4gDAzX0IvAmvLzd2kmEpjWALwxTK11Q2s1pyp
xa012h3SyHILWzum9BfcKovjjCKJXhAxIWPmrwm0nAwwT34igzt3Sp8crlacsCFDRIX4F+39v1+l
KomJbIFV8/3QOoaeSP9cALIMp2Tjv+HtFD9t5ZcYh996KZCzAeXgICzsZOGKCxmmvTn+ktfME5hk
YkPmplqKNQ7745QGtstkwkIVtSyykRM7GY9tSfNlL4VWJ2GdZkOpHty3tQB2uZF08FwjNk9qh65u
4yJdL3emvxLAPwEkPla42R5O1M7H88jb004u7Fzo1wLOdDCXOfKquJmStfc6uphD1IkGPsdvTU7G
27C6fcJ0OuNPyKMlXjGUwczywfeVQGJeMSS7o8FiwjqPOrWuBQgRrGAdlyaZ7kE9VZC3C6cJmVVa
AAr0YZt7c3n9ZyHD/UKeYCYTx+veI/9IRjaKDbjVYWcMMNBR9jLHRVst4I9xWph03DeiRp1pXYFg
B84lys2jnWWSprB/mpTRluedrq8hsn/01vCTdrls09VOD2yehKiSPIWEBJNfofOyNNJX2Kv7+Hd9
nDHUujQBw+/vBMEO7hyW0x9ASMWcXCP1mZWmnNM9oC156TxJze2ZglBgaX2qu3Yy59vz85bm4c0C
AjNMlUwVvU44z0Ap+gaF7aM9B+gC6xLI6flyl+ZXxgW1mn1tJnjIjWGiLCgcf3xbmlMviaUJ7I/d
KTsA6kbjvhrw82opgKjP6Rsua499mtLuaQXE/crs6UpPwM8Y/iyCYXjFriG2HV362WCemAfNMvRC
l3oxqvjJevPrO8gIi4Zjfnf3Fur++BEs+59Y3+yXb5nHroisnHx1L1ojvHtWRl8v2mm5sfB4KxWR
Ysx7DluIHQjcBzlkZQpCAtfRzyx/Kwu8lLyEwqhb6HSYzTaevA3BF5Hqu+7DWB5QrN/L7vJxHldi
HwYfH+KtpknDdMJJGaf9i5BNd72OrcieV0m3RcNJ9uClK6FMjyeYpBIuPmpAn2y95U46X/dvyOwM
LUyapqwY6cF23t8WxFRKFpbBWgiEqJ8I4P74iFHx/QFN2k6XRgHm62qBU2w0ZwUSdSC9NVNDQCCQ
15qHOEik4RLk8eFWM86e+KE5ntjSSg00vpVqS7ekTHFRhz0ylvD1u+wYrlxgKZQTWGBjE6sXMrs4
5DSKKH27nkBsP6TyDBKe9NFidndvcGq+xB+L01fPHduqS+w4bGqhfMcE/KEqU/mg6GSsmJrOq53J
LUPqpkd3Ac2gVqVbIQtyBnR/8ODS8F38FQatm24BaxJsWzGo0cjhCCbAjHAtZC0EkusjJ+3xq3GM
E/kXUHHH9kI/gpLpQMWsWXRhuh3Z78gkSBm3HcqgWCe2oLxKC7FM3G4zYvm85RrAfmacTBv7gW3H
aF8jOnsAJGehIfQHdWyHaPD7RDFhDXMWdQGTiouMMrvoX4Xn1RdxToLActJ46heeoXWzBLyrohH+
us4U5T1Hx6nIskM1mK/ZX3bUUPYPkhiMcR4XyW/7JFd4DAzdChS2XrEeB7WLzJjPMqMjtWUuu6JG
KM5Ic7sxGw2wgqTgyQI5b+0XLMmeroSnB9YfZaUY1ozmpg7XNDDJpwPyqDGDBfMxjYM79ZxTuO7L
UN/vYKyic7yLd2TSvkpLrpOTN/Xy575p53Qqe/+8LN0iIXinZslGJSUsMnhsxOMLRBFArRcLqy7d
nv4IpjwbDhLEvV+65GjoLOZPJ0lLBweYwwAcADRelQjnleRfCKQIAkNOSiyjTRjY2LKkaOWW64x4
3c0JC5W0KR22OPSZajjGKkJcbQTlEt62OdFQR6P/duk/+AlGO+O4s3S54m/1Ww5F9OqyL64n8kI4
c7csW0DTyfOkvHaMma+Y9lxZDIShvP2GBNqTnIPxud32kedVEnc12R6nE0Tj7l5zqnbRknKIJcWR
iJmwktPk1lsQbTkGbgDp9vvRYMan55SpbIki+uBKyLV8TCbhJByfzdIyu6tNpGc814p61slUaDjI
tl2QRbx5AOm/67QUOtN0B8/4KnWJwwd5zQcYWIshZbFVQcQ2oRnmu+Ok1Rn839YZ4xOIu3jck8QU
vxxLiAm8H8TLogdOezmYdo+j9G93RFzL68Qiu/4E589vDIEyvTzXReUuMbohYaxZrNEMRWpcJNHk
LPhPg6DSCCvUBaIzsb8G1FrlExv/SKnJWRXStLZvfqHx2YCveMpdzRN/sZ7cfI966TQMAQAXrw5k
Rl6cwbn2Svuh1x3SWyuUHCDtpHgrNpndFCruaejJLB1W4HpOOYn+SeUeX/lpMkmfqNYIongm7FE9
Ry4cgXOkDZ7DFkkLau6DHzKLsybN0HkjD3jbXzkf9NmTXW0hSSioQtaLKdNaH5WZozNCQny7+Fl2
Q6QQDLPzTfN+xt2VzrxDDt+VT107U1jjnlcN7Ul5LNVF23iq071vriJkQZTXx6JxhcQ4zYK1fNfV
dPzz1BLRP0VZJSzLot6tE7aFo3btjfeidOLm+mVNHeTCcIRyhZKG/oIqZ2lDxQ/8MCC+k4YQjeri
bKg1r1U3h658m2+rW3+cJ4Phd7wQyNM2KLCdzjkbIrkXdzKVvMJVo5wxPWtbElx7+xWOWZ3VUApo
IXnBy/38pHIfb4fRIqvT6GJa0h4MHm6/VUlLsEe6ejH04gyHdEmky1szDj/BAcK6W1w3bpXgPHNA
2C7/n3NqO0k/Io8b47xUdoma8p45maM8Zmxiu98jgEzR7Bip5k18hGOV05c1ROn/trT59V632Cxw
s2CWl9LOHe4POEShdWDNP0IGLXGKewDU1qIDPUhdwNvl9T9Rn0454YZnTP8Rd2sZxWGDZcBAfmIj
urVfkO2XNGyR630ayTTAufDHQIXv5Ao7jJaTTV3x+enWFZCotfB/u3O9913qZgx7Y05gDtABWFbn
cLNJa+UlHjDY9E3sSU6eMPs+OEuIY2yG9VdNxlOJqN6mk4jhb2fLwheuZJibgwLGrcAB1EM1gnZ6
apru80mCmht8CnZfF2bfx/UsKdzy9KfpHm2jor3N2rYqo8Uww7G8qDv88tbpORS1NRl6N9ilWgwk
H4ej3ISY4svFbNKyB7uU8Soz1BoW44raPG7k5hXZBBu5MBQN5XLbC0OvpwWQqPL6gE+wzc3xyORJ
qjDtb/VwYFI0m8Q6C1qj+D9H5AbBd1CxeP8aK3z0BPv1Wdv8Bjw4NnCmwIIhScHFCLBOMZhaS7nf
e1B49gWOhVGGeAhOLYKZEvTVvk5pXd1TRXaeZ3lPEl7+48m9eriTBeM1i/zFdWS9La5enYL8niA4
SIHe9JzBI68U1Db93Lp2Ot4VI4iPEvzczNY38SGTyHiSQHWXXVGNOMKs1wwk7+bMNK5whynsgXqc
WFS/9wMLZqjVmGN3yPRmsV9tkpTIpGSJ7LBbzZhU0mP7klJbcGH8j003FDa9JtAMrSND+bgamGI9
DX9fQiFNZ50QQDSSzeXmay45mCpapg8FyofssQVh8GOLMHYEg/oaNwQJd4X3J+fjw5FtT3Dwe1xW
cM8RfGTMRM0Nr1CGy0m2mV4pD64z2IvGoi/d9tYxHzZSuarrlSwzbsDEMoNJkzVPJWRIIIgTxM+E
EotkEHXBTGhRxaLOn8cSvwdTFRbt6/YwgmhVjMI7uqMsqa6vieQZHZGZ7dUrsWrwIOjpv8rjIBLU
Dl3aQH+S4wsCXoIqOuuufAHVybQ+C/TxsZQrrI3sne4NBA61lzrCWwh82CyoQYEGqss3TvdPlBJs
LGijAedhlIhe67ZlKLN7s0NkJSGN5P4k4Nlxw/6Ft0+RJUeOb4G96Rr/kOuFL6OAZYYhUi0vt7eg
Jn3XfLM+g5sNMUnuDG2sZlMLnnv59zVdHK7Ktk+G4XZExnhmK0Cm5COsM7cqtO0rQb5ce12JsN6C
nXmHIHAuWytkfpMuNRtYW+PyAdH87bB87q/LQCld0XkzL95+C4w4e50vvXnMxTrmj4GUpn6waups
GMfo7M0hF7ftI/GV0vDC8L+0XZe5TkVUllG3hsZml2TW52prpvdjYAkc36dVxclxzE8Xlx9fUTYi
hgIM6Aj2iXx8HGpm1VyqFclQVMbFQq8wq0p+1gOqY9kPJqhsBy7ngpFxPR9zp75vvP7Sdlw3/a6i
+9LHg6XvX8DXsCdbo3IrEga19UWgfm8EmuEKhQg3M3iJ4X8/KQPly/fCQ/wQKKcncs5/zg5ZeaYR
9SQ3wTXgSdcrjtrdW6B2nXheQBs4bt1ZRw+oTj44LH65vpDALiqU361Wi1CuaU62v+dMzbwwKnfj
EtdflTg92h8cneauQL41sNTzqlnQhV9NnOFFEi/xTMMniVsiGm157XXmwI3bxDfIhUIkvVj0kXIh
0NEe6UoGruNWXDLXlb2eHjoVrKUVOvL6OLYMi6t6NzmdsnESGs758d9k/r5KRc0NnMooXUojHG8/
On4xzx6XnJttLsedTA7oOsQmz4Tqibe8Jau9e+6th3jU/ryspnt5V4/E9ikukAu/Tm3+T/q1Qk53
Z5OW0VBoYECuQlwDwq1sadfz7NGbcm9LVcsByK92VcF+0gtz3NQpKY7EkfoKZeGM/egNe22vPKi+
IsaUxBFBmVOqQdL2iQ4RLYdxh4fFq3e/sN9Chrdf1F+ZdOpjOnrTRUAAT1/VrHoTWJeVQEFvtEaU
FrZg+nb/wUGuTwyTgx1nAJ7Sx5EG2aoCLhHmtFgV+A/ieerLitwaoe6gjoZwvMlMlEDJPGtOxred
Ie+CsB5RndJoPZ7Fwss2Cx4Cq530KNgalkpH1HYsQulb1CEPO71uconr4Li16YJ/yHnwlq9ZEjbE
ktnZJztLpr5SU8+JUdYFuEGeOPLyJ70yJQ8MegPDhwzaLhR0ESP2si4uuLMln2RV32d56OezUG8a
ql3CRKkUXxEtRoPP9z8/RE3KGrwfkMbCV6R4IBdPDL8wjA0xTfsGmK/XcbNvvn1K1m7D7KrklS+E
VP8MAK5uiWsWoBu8dxnxyL4kgmBWrWwi/nNBp88wUujnWQ+9A4BK4RuZMTw2Adw5RpYy0OLyfcf+
6Kf+GGgU3pebGV589f0lIzhSB8B/+3rodot1QCZZckKP/hOA2OKhc6yAP9DF9qFYLhisjxctr59O
gYqAeyv2m8mWkTd78uPQbkCWMPCzeVnBhbZQbF5Z6vvwj6AgMSkP3vddASEvfDtuw9Hf70YcDIob
WLnebh1Vwhab3Qjws1UuKkxEZli9tAA1HOnmzvnYARPO++bHm2tfJJSvQyCigL39ybnm3xRznlM7
xaqW7/jS0VjiCQ6KmL3Zhz/gj8Lrl28DO6Eam679lACDcn7f9f9yeLMpQdawJOds63c5z0Ah7Nqu
X7ze0YyDH0xHFH9OcWPrBL4btkZShVSfShc4G1x6Eq+NUJphs/c5B6egr4S+MhiZmrEdOUwVDzXJ
xiV7uFWjMwvwqYhYdiqupvPw4ZB/wgV+Lu6oJ2HF3xeNq/Ui3R0eud2mmVNRYi/5h6Mj6C/djz1O
tuCUdIAeBG9zzHTovXVfPBHVIZ45YFYoANoaz7pRapUjWod4PUG4Mys7IMUg3WL132/MPsrQWMT2
UW3X+gIJz8XSMnVyMvnwhIqqp0bmkOM02oYvVqmRgW60itPKWk2zv2VUrdAjf42cE/1xxKTyeGWD
VvFXVmWZd+ZhjePiIof2+Wcig6YA+KFgtdwPgryX+rlQQs2ztUdlGgSTmwe+y7yn3G4VIGIwS68m
VFsGSxehmAQBfBMg/pb1me6PF+/jmHyPHCGMPDWuBtLF/GUnLB0JsRRUEhuCUd46tLsMZZvRnVSe
DUPBhXfzlIAWfqy/eF2PdUskGNW87gTtZaVXxvAsLxVhiHB9kwmjlJyGWGHL5d6HsH5Fs+XObj73
TkHqIWZsNWtmCUdgdak6UMXtpDCGeb1w9FEuD+Q/kmj6wJXwKoxl4l35DPrydEd/+GkGhYcmgvHt
v3p5gTrMRtzUylIKvULTEFLBtT95xjIkvQvTM4UoK8iYfXzEOQFAclKfKZig95ljOOH8BMGW1xE1
5dBXWvbbb9uoMJcfyxx6VRqTEgRvEMbEctBo3izWDB9+yRbzrS00+Ah5WGCL/wyL6YoiORGceW+g
L3WOWNNF6e9uoYl7yBbJ1RO2aeW/GlQCt/CKy/Uc05HXCxu1QzJrKOwyneXaH4xjT4Orh2FLJvyu
Ukh4R78xEz1MdPylzx41u4vJRMci2PcHjbML/EvrDEtsm0YGpd2NPtUCogtrc4+YU0W0BJlfZpWz
oW2SInJKp7Jr+PdV2arBCR3MFwJMSfnt4klge5k6hjTgM1NMhmpQwpjcTmikPGvsZvCSLxgrUCB7
utWYdeHeSX37fivs8B8h+WcV1ylYL67IMpUY/7cYzJ0j3xnYYOhReXn2G6gfe+jyPbIW2Tpi3OK1
Z9XUzrLyXUxQlKRwsExEqJta34jvbtn+DpU8L0Q5jv8kwwIhBYWs9q3nV5bNzZ0RfOVZxYsFHWg3
6GUsw96+/vfzy3/bhp+BcS8knZ8LF2gJsQryHuDDcNAKmviAtr93+ggtengvGGlRfCDIrtzGv6LP
MNiHRupRASt/5xjWuReE6FA0+KaREaUqMRV+HJHqT1EGpOhgsOP7Arf4n5CN2rvnM3PjuwugdCJH
r5JLFrVcgUPYeWDbpMOJZ3YdLIDFhtgAQoKSZ9DRJkgh822C0+rBk3QpjWN/GkaaR3Ep3P+33/9K
Bd4BaQSqwgyLz2bZDEJzSDiNQzEmyQYRyD87ZPWoX/ByOPob10pd305hI+i4eRwwT6bZdtCbcGZT
/JlvNjy4fARWXcqu3twpp2sddEzXetsGLCAaZW5gmzxZuUblfys7jMaA1K+VbLtlwW/G9sZoCpNl
K5iPDsoNs2slZSZVez8aqHHvBCPoT2rydJuF2wMLKdgZgg7W+8rubAIrYS/aOYXn1Fnn7caio4tc
Hdi0kV00/IsvpxNbfzTrDoeNj3BHmgg2OuO3UtALk20BtbY/p0xvFFPp1hISDfNa39LL66hn5aCy
FB1p9i5v3ChYBiUjj3E/z7LcMoTzfZ/pJJhzPm09ZR+snJoQAP9JqVrBiK9gOP2aJ43B4//P1YYU
rtgzt4nuGRJJnWaj3EezZA47gakfyi0oiaeb5gk6s7KFKaW/QWBImLrd73WQUmJ63cDS5tuGz4vU
T1He1XocGHqwwcgSMjY2EE9PPExRdmmhNltxlLYvYF+vI9ke28JRrCbRoePqvWCXB7FcMDjEM+SM
/DIholXfqWbMY1JTfozrnSrP8e/nnvqAOSeQECQHZePSY16nX6sbpXUwCOn2UFc/UMezc09QQuhR
wkfOnyX5sh6jpfHJ5G4rpRRk4RHOzbKGJemec5OnIdkpQ9CC9sIf9w8qccSnAD8YElMirjmYEQuo
EXG6dMlQ8LnHxrinuh0zVmbhkgDQHm8H+eHi0FmHo9ZkYlBo+t0HzM8Efv31GPLMAy4SwiYK+hx4
JC+K1U3nQv1gMVJ7MyeXkBt4K7WMetfNI3IendAx+Q0XvWBKHLjDJTn8YTNY29jhFnCnEKIXp8VL
djMFF7vWBfQgZ9FjxCCfMiIxJeu3x6pb774z6wYbaAW1yEkGoH059YGs+LnK5kGwozr2Hb3JZ8TG
R4hqAR6mzxFVsTrasvsle7D2bfxL8M4RZ7fwpqGRVQZifUWoMp5vTSfrbAgetvTj5UIXNAJ4gAZf
RJkBRMce+ctPHYdWIADKQ6qb3BV75geCr/94/E/PlxpbLCS+UQkCyDDilMOnBcO0Ga5chT+8pLdQ
pzW3ZwE4E4y9J8Lazqc/g3w1nr/MJWi3/gdGcg4TfQR7L7a5s9UDT2V9IIpff4dM+VtgMzDFvz4G
C5k572w+ccxLFiA6zTzRuVCpXHWOX67lnski9KnfyzHKwjB8hDUjeylwHDpfvr/zum9ygW08nuJh
wfrS5jDQHoTRPhwgBmZftDKQaBN31PuwCG1KVXMMfOL9FozrOVRWjNrjm6/wwrpk9SBJOxGA2sTu
G8j2d1R+mMUAz7q67jcbByDP1SRHXm2FphtplAl3D60D8GH/wqMLSFt4L0WfxLRWodjxUL0OAGlo
nxR0PaFipd2Q58ahxkMOk3ukHZfkSJovGlBdMQPsA2mglEPQ11z9lwVRbJJGB4yS8Vs0IgS16mwe
X5OyK67PFMk96C+aPCGWQf8qHsQpEdhodoV3r/eoIpBY1NXdE3oUcibixph93e0rGLQwisb4kds8
/7jH/jrLi4vFfKDcwJHpOivkaKVeRsYNzhJ2z9NrVSvof7Atkb7OvPASZ3CF086peT/b1hlgCH9j
T9O60CSDR3NGEV0t8GVlrai/7PFtv2us2/xMNGk/dg/9kdsIVhZHY9+hxG5cjhS6pMq8lErkxCMD
5ZScIhP7ec3PbLR+/aAw4D5UXBk4c2ZuEABKQyXRw0jHMXpTSwiLMP47gTly3y05LBZN26LdNFoe
IKiBij/5dG9J74Einn26MOd5bebBCGhXxIQZKntG+3Tgey87aGJCDWDTSBeojYa/YCZ1agdbcPYQ
xYm8f7Yr8a3cXFOrgbzBWV3Efpftk1xzjHTpLlZBKqBuNQaQ7fhYcJEwsJhkk+ZB0cL+5xg0HbQ8
N2RJkTw6+pXFNyw2n8KrmdowWfp1HdQHH66qzsA/x/NAqg0sxU6K1eZrxyC87pfUv5S4U39mpuVj
pG/Z4b/lZRECuiJE0O5fo89914k9FbycIMXokekE7cZCJN8YCQrSbpzS/SwrkgRWvMdGQGN3Qn6l
B+FiVUt0oIBd9oQkcjYR7F+5385ZkYEbsrrfn6m/SARbKGj8349hr1iG+Fx/5lmWf3hZ6GHnXnCW
fxJ7AcI+LHjN3UTEtOsC/dLyj7hiY6pVqanIhp7bE73A8/Kj5c7v/FWRgWOeZoHJPV3cl6dlExLJ
OqodLFOmEqWEaQHL5wdnLiHxG0N/u+7QFTUpqG15k+oyxvQfGWEhXwRljUGG4LmezfwFt3vlMX7n
Rqwn5+pI2gNuJkFFpCFGGvRtkGjbASmI4vZrog1cVGlSCk10Pj/TxHWnhnT4bxoihBEA3B/Vn8iA
0AxmooW4DbJpZt1aDhHldZ3dOTtRQV1mQKtDol1WojhRbMCtMZrlAQhA3HnAI6DmLnFSKyh4bfgN
JuZqv1A0B3t2V2Yjw1b8SfduPBYvPzkD3Qn2J9L6ms0lOZeENZBa6E+4/p5ASQss9rjmqqXBsHV6
rO7VP8PFeRSgUFrEgYqwBMGvpxWx4ojwWzyxTS2IbkFGjKn7uMAob6ClBjsxBwc2MwFwxlQMs6T7
0H57IbL/9vZfCR8ES+622LbL+PFua6x1UosorXqnbP+TBrTSO7hR52+gyCs20eeCOeQcc+al3k23
QrNcUnVb5GBBC+wnki2CyE+ZlGwAhRGfqxHVb4p2341NkitVbEPnJ/g/mKEjlew+UABZvU3ES/w8
JG+5rxS56KPaIXESOLoUJzinyT3Rxc9Oq4jDDo0F7El0RnhNpFPLpfuoM5baT9ehrwz+xkjTvZey
DFySM0MaoLVfngsAx6HZUblcwmosop2veJE5BGt/I+23MuYNVEtcYGznelSFNIUSZF0o00CWa4+D
JsCMXsLcjAnKyBv28SC0H/gorCGN5E6SFVnGn4Ymbnt2rxkp6irXT1j0nng4Wvh+mI/h7PiyBax2
YyqrS6J9TWTcFD7LskF2K/pHDM281P+sfCrvih4fmODHQldMr0aW8lHraQKLhaRM98l0v8a4nfIu
+aOqo5dVao1pvuA6XK2+kNUeTBnd0Hjba+Kk6fzZzDZoP9FgMvHj0+x/RQJU5AW8QTChuWm43uaJ
WT6I15hVtlzabF8XK9Y9DpHZANmnVqW1C4Jl3EQTku/J+YHHi0pCfU9WnUOM4xrmZm31JGtkd9cM
q5f7N/oNYeVT4W0M9CuS/cLOWQXe6xvxcyw/ngsAsjqqFdANieNpB9kqIMc7PVHi0A93efHZrlLN
CctBDR9EWf6TxRWQRWR4Bou4hn9th1wYnoGc3e3g+zRstmjnJtlpspffEk8GcYgsCEUwR0EDWvN4
aFqDRy8RMHHpr927qcYLCN3zSNV0U/20TVP22IFdCPefL7bsJ2qzwJuXHAtZ3rrMnNCz3fBCkqVI
pBWBjUyAz5FYslCeSJdCkiIzpR4tT/yvdRx1VbEawWtzbjW/39i633GkasXhaoTLLE4SnxI03qu0
5W6W8iSkywSsX8hbrnG9n/r5kGeTHP0c4PvorZRo3Q4S4eNsaYEj1kxrDTbFGPZHxPFQ/fZAidFy
tGuFtZHU94EbvygEUW7E7w+4jF2GiobVrgKCKaX2GqAZoyIxYdfSPaXMP3VCwQeiMpf5I1b02Yh3
HfYGetRLAdJ9pynLv2Lup7zG8eY798t5Kie96FD3mTUsEBqoFBxAKwduaqP1SKbcfrQu+PbzHMqp
L95Lb8v4QcBprtb4DHF285f5gwxbwkub1DCQEAx3uaxOI+qrWPatWazEj+EOFodCrGWtVKnpSTGm
6KRKl3K2yEhOV1W8J1FRmbY4ZT1HfZKx4CkW3VkS+a4A4jsMXF7n0OgC8o5D2cVrUltKbrdPiMLg
cHa/UScIDrf8Q9+hS4zBW4QgmXY4RYu4pfATrrlg4XLQeYLi9CzpRbCz5txrVCqFyH7tiwRQf6Wo
x58KUFDmM36zlkwtELTwyrFd6ZA1S6tt9xHjdjeZgyMpOQF+NS/CFqGqCESNyE2IJ+F6YiWdD8NX
dGrxBsFUeT5+jDHN2J2zElF6+Idl7Z15qABcCSRKNDktxDJdEWCmJ1tv6/MEe3VkQpB9/wL7SNdZ
70ZdtWNkNEMRTYKGpFgN4Sm8Aj2P++6GYq5/+URVlORNRIW8Al7XtjRoi/96zqQvJDse23lqEW/R
l02XlVs4crj+DEngEGVIvVyvv+mTD6jUS5LDHtLZ6uIKMasrJRLc26zVWwWv6HOgfJwS2gAUwMfE
eamS3egBQjR14XxA+G4paW2VQ0a1L/hMl7k2D/fcTRSJH8L6uw+Q5PqiSejklp1aZ45ComQ09/xA
2VHOlH3+QLlZW9F104uI7QkLCBEz50ooFcJSuRRLW1P59v9YNDxm4U3mNhzCR9PzcNJMb5UjVoTe
A7K3WgPTCzCkjUw+kRoh4HuYlev7zSLIODGE1s/yqP5wN0udy8Lchv7oiLQfZPAkuiyuw2Bj9Y61
axIycPOLxQeeDL3DywIn6twTnsFU3Y2EzB7P0OW8WuLe1m7q/J9bP1ac8f4IeG58j6gDGk9NyTAF
H2Do0qR8lnYdt6pPwPzoEQl+cG2mOpQGy+nQlYMq45KGFU0PiwDiNFq3ATtqAfWOt8JZcKbfLmpV
8hRCr4OGOu832ohkrEzUSWQlCv8LSeglA/OFEE6NuleDiHvSxl1AmUJIAXMX9KYyLBQHxqJe/Xd2
SEhmrjBGJwskiP3DQ5ipFObzU/EgZXCp87z5uy30pvcJ/Ja78XZqnmIyqndwhVTQiHxW6ZJ8Qvyd
FRDNIW15nNgyomOHJmgvTvAs1ctMZ4cVwhCBFuJtwg9aPTJG7IwI6rVRf9nT8Yn4rgg9bPyGSfsx
Ssb4NVcZNiiQAi3IrkHln6nokco6iF93x//xGc+JkUw8bJVYayd0KFmFNyKS88GlnfbgzurVRwrM
9Xuq30/R7nMPRTLeElHpU67bhwUcAdx/YNgg2nmDWHT67NEKI5u/b44YqrQ7hzmahDwiRHNOb6gc
VjWH008JQagBbwzXEJsqyDARGG9qK647aH7s1VhKRLJh9jlM0nsHJCIOA3BTLdWHjqUY5N7NdR60
ZRbZ4ZkjvTnHBVZYA1pC7lI1MotXR/HLSpYaqSnFHdHx1fOlF2JWWhYW2ol1Dx1Gd10/G4wOObk/
9eNKzd+dV9UaE6lrrEs5HXHlqJXRz6d68W9+idExXOlEf8fzddld8rD9ggD/HHW2AnA1LCKeGnKY
IjXL9/YIuplBLiFRZS/n1zAyunlpJlAgsLkDWbZtbmbUl99tRZdh+8VPVt+1eL8C0F39QYpff3TE
ZgCPA/+sutRc+PkBKXWf8VOicEGUGrrVvFm7r3P58eF5CQR4kCWkeoT5qcTocrgr4QeVcKx6GnUu
129WWka+09tQk5b0eKd2n/3kzEioWM4H5zhpqO7AXvVPLSz0oDPcQ9b7FnMe7bAR909LWY2wUN8s
RMe6I+DolIlttlEDKKSIIshQXknmsZOGIdS9H6IQhjF4+Ip9cXcyhSWPLowBzW/ZLrqmNbXivvcA
pJQUbP3EAQ1lhlEeudlLlpQiOD1LwkdzoIU7Z2uLpKSq6FYperbY4mJS6GV2BWbc3y0cMlxAzQB6
e2yjDFUIvpHalBkrDFL/DuCkaJtaDP8MISUAlNT6FHnPOqPHV8PRhT0UYk0XZccGn3mVw9eIPB9p
YyPUS9QIVuLyDoC4m6EYR8ASCz003Ulv3oS487PScRLMBvtI+b7J8AXBCySNwKrQE1cHhq0hzheK
WwmhCco8rnot1lRDiCp0u2QmC0DmvyYEdW6aaJHBVJEDo9EcH6AcYOoqSGen7E+hIyMFLvNw9zFc
ULONCGw3raPfpAuHNw3Ty44Y7O4l3Au8Dix3OwdelC4QZZtd5IAQXkqKmmCUN/jr8fgiELpEmyOS
zWYajXi8vOrIcovg4E88sYpVHfEZ6FMwkc2/hXnb9WhdiYhuJGmfb7V+eEti/N5kgSpGpDk3u/5d
fGF36orLAFdzSS674drnuhbvHlNhmluihpc65EiII2IUuAGk4dj7Eyb9OYlm8vjpQHhegNAk/S/F
T1TC2lvrU8L6NWNDJNHzaoOn2srqpcojSE52aX0AAj7qZuS88OYpmIIEbrpXotbOhSTtHzuxSGfY
Z9JM4hr0dQVyu2SiVFqoZXg5j3NbqBHCkCUfFKkYK3EtkOX9zf7gBaNOb4Gb/8t+AWysEtyKPwtQ
+d8sKJSFIyBBQrId6nZYS7q7ICSV3YKIJqquUGcW9XQunsWHzDN1zQa14IU08We6wdx+GWCUz+qk
8wADBCoYJtUIpa0ia9nbmuYmEN0gHdkr9DVhd5IVknu0E36J5HgXl5AAk63Av99/BetdcE7EEyd7
+tk48OQaXLUOpSCF4hbMWsfTn52qWsyJPDwahwALVF1WkkSiyIheUqkt4U1yZIZMrAKZY3/554wQ
NNp0ghiMbZ/8SpWsu3QEXj9rU/1MZnOVHSbmgGYksvFY9wmQiyCVhzYahrTb4F1AU7M6DXE9qChi
eVIKn2CPrjDa7DrOWI92RgXNLMPQyd830ewpl3vzyoqagxfpzFgshuJBHPiobEI1LR+iU/iwaTx6
mvenwgPikmjlNpwSrRsIFEU+OOOLuCl6GMGsyCBBzD6f4YINGMDOKWEXz7Xq4ZOtjJAOFj3roGJd
p2DCxXigormVs5uhDZRRlGrpr5hNvTKOQfh5iLcwDcQHCsYtKIjsKUSS1szfFHkt1r77jijMqVaR
+jvZ1/8G5e7zhA+iasrv82oJ0q4XZ3hOJ+L81kPJRxjwB9owO7CJomHUba+WXXBZa/IYUm4rao2p
hLlaMPvdE9iS1DvCfNxKnL0eY5M6d/iy/sEdoTesN/EfWsljLLF5s//lbgg4tg2fwFg0l5MowJue
iUh05tx7f3BQJaZnbUEO2QDTOw40J0hq7VXeJP7CHb0sFRephztXLq39YZa5XkXIpB4xVzYSJivn
pDrTBpF5OXrrhdXgeFGqSrk41C3pfWvemdiLSkxZ/tL7lKyb+3FkD13r71+XpAglJSiGU39mSz2I
d5QEfRUhgo1ccp7Qj243PHK/JJT7IGiLKhILh4+7KlDTXOT4o2ImS+SJczi0tWOYZyxFbFlKJIK3
6FLLJv0U3ijsWaOdRE6TlYU1dJ5NAXEczVKl8L6yJ2bw8eyET712qUPt4NAk4z364XyKL4h57458
MQpzqewPDwaBsu305y9LRRcfILmwPggQsBsRJ4aNqMXyeIdQn2sDoSWjYkvfnajNCLAVYIXBlydy
A9I7FAyX0dkbH1gbx6mLhQiVLZIX1rPJUXQ/vhUJ09Sef8GBM0guIs9mMrqi7Xa+3qPuAqh5Yyp9
Sa2WJ5tvpJ8V4v58AXTMrPyAn5GY9u/wOjy/r9L1uJeotWr1rYDd0N/Rk3QdVntDa8H1dGNcn/XB
a9I9Tf1/rqnHlxHiJXqPybu82tNFFmX1FzFcG1v/fE9NLZKRQBNnFjKjrWWfTffQNaerp/EN8036
er7hQlaX3i6jR5xX/OV1IBWneeubfTS0WFv2LV2fxdQC8p8BjZ15HtRCG2dYAld5d43gqCxUESfl
YVb4uf1Sfku1eNk4rTgT2YgapDSafSnSFJxf9FfbnyqRfMzDUoScfqZJsma+NWNWiXAbpThNSStL
6yo5NhZrL6tYpjgSGzsNLO1SM55xjeVgVDc9s4/+ayJ0lV7qoRs9LmCsdlSGh6F5AXn9knQm1/I5
zBB8ZAoQeTg5iog8RhWLIxNeBqB0znI0YhKp48fIuf8AbxfmdEDq6WeaKb3KiPcd0wGHvvOm8lcx
ptNV1rZhZ+Kq8w2dlmBCnHbQiiLdDMF4g5SvZ0jQLxw+FwyLjk/5usAy6m5IQqe0MiYgu6MDbrJP
zeF1Yyz0bifUbPLiEB9sU1e4/STs0Ze28fJPfVA1SC6I/Da7rj27x+lbTPoK5gjn+Eb5HdyR5NM3
laBIMjd4zGhOsK4c9m1Jj13KVs1G73kg832fdfMTbyYxEngANGvFqFgHm7jPvR0tXWca0denqqfF
teknBgApC517Tsi+X+fEapyjspg7TU3x61/8pfVxjhUrrWpfPBn6BB9+nIcY+jAaDHnplGwgMTEm
9Nmz+Es9yTWHVYl+3moYyBqs7DZHGPjmNL5JYIXeoY23MMhLdVQQmWT7WXXRtpS7EJ8N6LeESMg/
+DPV65ZsE6R/EDvaTsnD3fy2q4NvfRbXAA3SXQfiVMQ2SYEoZ2YA82pYQ0O5oaG835r+qX5qoG1d
+yax5d7sjlY+uPNCuf+jtrLwSi6YTehK5Q2u600FuiFtx5OoniMeUQd1PMLc77nOOmXOD8mKxCc+
WgMw2/i9SD8bMVY0FylEcaicKq0SMq3iscbP7ZMGkz/eCxTgrl/7zMkCDdzO5pdSAp58cw1uswu4
jEGJW5YtLTKYcLSXhRuWyiXjE2RIj0nSfCcbMZS8XYD+jemt9mdgDCaX0qATquNn+9RqxjHoqHUx
3IoseGzen/e6fYamiSMCGb25DWkjmjbp12vKLQAPhDMAOTnvUbmN+3iLWqw+1/TGTAQstbE1sBa4
Cwpwu4PlSzL6YHhBOEIW4kX0LgMUO+zH7mq7k+noKXjInx5mABPkPHano6Tjg3Ws0n3yLgW3rnSu
Pzg2DyVXcc6Vge25MkTMpfMZGPEun5Lz5eTUgiwJw1SWWN8HxCavkx37InDKz7+4niz15ag06NOv
NeRG4VMLc8sPIMvk6yixpICyoo7CzdHikj6tJKNTReWMoBmxidT1gGjGfRHR7/H8mjBrYiOwloq8
d8xp7L8A86Zn9J9lNXsk8/oT0AAzCPlIl8CcTR5WfWpnuW83EpGQCiFDgn5Ua86rg/XmTZarPvG3
Erx3qa1HKuO9ZBfCxdV715Mm0WAL8BVzK9TklLA6GkxumaFbPobMm9iwODfjsx5Uip9Vh8Z1RLc7
AW/KFxfrSOJsOog8KoOw4XcYsPXKRZpdtBSeFVPvXByoZo+mT+QdYsu5J8KI3XIDd2LccJHizxmO
2Y6IAXiTsGiaiOvfzJ40f3MHBUvPm376sOO5KQUq87Y9XYYWzl2bdSDj6QEu5jm7JKvf00WX1OA6
w0CkZ7myuwETCiFTywe4aeO9/FMQrNo4wc6vigFPm9TzcAeyyi/zmGogoFfe+ZH2gazE8YQYx2xL
A5Ogjxx+bs9dY0sxTzyVNE7pWTofSMUdt+ldoPtZCGQgEtpkc4QOhKs8b6G0aLqu79kC6V5U9Q99
vZCF2Le+2YR4e83jruKomFric1IVS9DyNuJQ4nnrRwaYY3JHJQaY/G4A6/GMVcmlqrcHo1N+VtCJ
ckQEZ/TG4UT9JuAoGTNxwrA+rmwyBfKb65XvUmz70LK2YoGaY9Iaye1YGTb+zrLHDb/V8zgwf1Os
7bS1aFg00NAuWopuw9MpC4nZ5oCYC5ev+Hhzv+OIf9ol1sgi8NQtWrJWCMx5XMWZK1YwzBXBLiCs
A7+a4Ds3VG9RMNG4v26DEFvLpsiHfFuT8YXHgHHSG/KntI5sP9v+lYyrfKr6kzxYG+tLyVpv/L/G
0e54UtAjmX4MKFFVzKB/4A71RvnAuTGLiThYMg8FsDRKNaIy8cDo+yMgrH9qXeA7Nrfgdi/6DEJV
nfMb6g7YcLOhG+rQiPwu7t8l9aGT9mraDRyPIWk2Fi2mfUAF1l35sRwJ0tE2JY1G6FJNrfm72vp0
rN1jzX8qePBx7zi4fl5zkUAAqHxL6X2j3O/7xRBgRArJOS6GlErAD/PEas1pXPqolu6eKfsO1078
BFP0g74Cs7qsKMS1YyY+5qOWljDbqYWdfOHWsJs5mLX1pyAKP7WVAw6M+s7I6wgvvlHgRGd4GZu3
6kro1E81vVhod57Gucgo/gQzdakbQ5i6s5cWbY0mUk0fU5VQc7jfepGAVKp5KH2oQ6JLzdqPQtvd
Ugbd5lo9IhqbYB4t6x2VkEmkj07qLji2dVb9KhfHiixRuiQSUo/pzyIE650YKwVD59uWdHfwlOwo
bqgAfbZ0/pwf8KMlyY5aZQd4CoFdoabR8G/boxWMjruya6i0vCNeOt4n2Sao3oN5Lh4A5ANXK9d9
LVgGyP1iMvH0oT24gYJKbgBn/hUF6jGuOvtybzRJ3c2lVIivlrdpmG/sRQYsYPOrZEgiCHXYztq7
cgMrPFKDb84kem9xy7emOu4tKWNyAgrTvtBiU/7p1CIPOuad6H8L/+HKywf0+GzxKjA4Edj7XGkR
BGvbUSQDDLfM1LRBQtcJPqLWz23G/l7y/MqFsd0acp0MLqZoKeDF1hENn9K5diYcS6rxfhpgbZmb
elosIHZBAYWFZKbt+tPtWXQAgnf+EUt66zyUIoDy/xTKtXOJ366l0oRRsADvNs+GTDW5QG9joWU3
ExBjYh570dPXNzTPODe/yfiIA9MKElGzyxCKnN6AdEDmpOnTfaftcsRCHoWOrL3lzQ/jkX2Wd0PJ
IS5/4Fj8Qv8rfPh8FxdjhjOBfrq6B/oAGjBtvnXQAx5tnALlC7hx52yoiwL4iTrWUi4pKIcFuQdT
U+iziH3pUFl28xiW8lP7baQVd8sy4wSxIMJzc2zmGxusNAazqkirL/69gLpoR/Iwz2DzNOB4MCuw
p618Clwb6cFYcOOZVx+SIS1KOXP8RLR0gaqa/6maKJnxrPNOG0EdNGwtmiDvfnqFxWqp8ZDVBikr
4IjkhhxnQMKZNbGM9cTzeGxlm/0B90BY7swgSftF9ssBmpURfx1GkD6f1pPDAKAurjL7BPZbUUzZ
FN/RnSxKojg3lcZaXswhNMFSYJnN/1RF9+tM9r54kdSMRrisMzmPpsURECgMbC8ptlPzYmjf3/mc
4j30SOPX5cRKtqRIBUrBg6J2Nwij5IRKtQqNyaD5VpV2SfV3nYY/D4JlAq8lRBAbEJKYJr3rweeR
F0wBIUB7BYkjDR4ACetsDtucE0BCOTz2Jey4IznaVzVsd/Akmfgds5f1FxmZLqz1C+2Qz0tlGAOo
D0CwHElJXnIBiaj2VDiJih+b6NU9KjCC//I1riA1sqMRV6BO6V6fi5T/AKm3Hc/9s5bTAGp0M39V
A3v0+xJs+l4EJa6TrdEiUigyMIJS7PLn/XPnKsQn5YkGVzzEEYcz3IqTS+bE1MzfWqAzmfFE1QIf
LVv1+bV42vnCHtYeSRh5JFnuPYNAW2JWBDeNtBOZvbC5yGtMd0B7Ru3+xVtdGXCdm4S0lvHN/u0O
2DINF+E5q5dfyAjPR4yb3fWt+8awT+l+C3VVa/cc5mbZVk2CQiQQm1w4AW4k6H4b1DZAxEsOzkn2
cFUtBz2XLPwzMgBmpebn8QWLB9OPjp5CWNYMMveLmXBPwxtkxmAeJQaO91hoU2md69AljdGV+Noc
PrpnlkkoLaadIWaxbZEY85aBZ8Ox1VPpLi3GPSGqs+E3EeEvrM3lYBVx9r5wTmhJOlUnzYwEBt7c
ka6uenPeF+BcMx7QXGJs4zhTaXzxIZ5cbrV+5usrjgdoDdVUdLRVfRLeA5ONt3NxCiMhhyNLsR8+
X6hDd8zl7O/wGRfRorLofAKR2PY0mdqpR2cHnGcTaGQkxeQJJ9Zut32sBpyQ7bZNkGRrVGhTxbek
g4TKx03YURW4EHaTdv8GlMwijOx1WLLN7IpqPC1k7z2icsKzVMQdaCfz4tg7q/Udz+s1pdo+k2B6
V8XkU6FKnWMzMiNiFmD0352SCXApR52B330gTDAou3Y7DE/EusDAOdfWhEVDz8cGLx9msyjEJ+NH
kCrLQSOEwmPrNkBcj3k7UTzDOw1tNy9fiQK19YtEfQck4ACC+N1dqTI/NgC6ikKpYOszK7Tx+dfb
FBq1skZOejtubyfAyjK8OEtTA7zIN4MLvIhuGxuRo6a9fgtDfjBHWZFMMATAVF9Pu8kz4YWOZdWL
iDX2esMnITQR+rtxf7DnVqrQtbYteLZKbbqP/hEhK0fxqRq8llKolSYkor0W8au80eRyE9AE5rHv
0W2BItewBDCdjIgyAWTUqaQZE+//gaQkLGSxgYEa7NoSHPB+9eDuKqO9lgbqIoOA4R5dG7BulnKN
XkmSqurnnFJ3E8KK3NMEhcOQhY7t3kld8Mtfa0m2OABsLiHytAgWzkzAG/LX2+SkZMBhfVhCufJe
jT0XaC0B/MiU/R8MLs+vuybA4TvQXO8rJNOi/iXgobOLrWVF7P9QYcqRFv8s4ssQHgxgydJqp3ah
WHk3RX+wDhMMU81/m2bNILyMWZTjMtm3byYXy6jMjoWmHFVl9tQxdURGc3V1LbzrWaUR/L4zEkhb
RsICVhTojIgL3w3/3MnMclvYL8rfZRNCoi5fGnlCSAHqzrxtucDF9hNosqbWR/ICuUE9tPxXhDyN
qVka1Pab1JcHwgFk71/ZmhajVk/RuJdj8XtMo/Sgt6k8R4i32p/xuTQUYvQImN071+QYsIOLxwwW
Rl1qsoKpfKLKYvGToO6fJ6dF4g9TrTqUgx1iETPHF6k+GoZdRp3GOErTX9JGLUaYUbz81YnUSnNL
Gp2Pl2qGEi43PdSTWeDJR4GVo15ITBxaDdpX5Eh9zAWF0NAaQC2GtH27eAgXiY3Q2CAbP5PNV/rg
3Y8DjIPKAqOZlWI0x3ZfqGWlkn6Bd/qR+R+wYoSwuCWSVcD93hG9KKlbNmfWfU8zsOh3yXoewLX2
6FnfeGMFbC++b8V6BKOkwuUpnz2zHR8vcJmgFYp3nr2z/OOMJj/gfRkY8UQEUkSUXQzLPuvHJR0M
pdlPXQCo7LObPj30OOYD98lRgSk4YMgWtPmKnoC2DkpLdkA3+Xuq5P4x2VsJmr4F0HqHQFjIwI8m
1paMawD7TH8EyOAY7x97IzqNr9PiWa5LC5RuMcwIox7Feo2DjMfTcQeA/y80lxdpeckIjIYJ+K+Y
ZwJs21ZXaXQSAz8Rwd83/kZkTJ8gspk3VzdZvFuNkLUDoTIdyTIgs4q5vpkrbFLtRARw9L18WEKA
+XTQIxUmgesRqpg8rvtRhCM++LRqHODRIBCVLBqxF3SXK3451W9sp3X9fT3iRcUB/GrSzafFg9SH
mXcwE6GeyYcEIywglu+gk0BYvgziVXZjsxIRbpsaI/DWNErZTn/ESKLrrxOj9mXjwR6rxPPDmUjS
9+tdrNAe/2VAumlollxRDq2tpF2l13l4aDzW8H09J3m+E3rPOd0WtIQgVqrJlej4lXQf56qTT4aS
vOrQjr22o+r4z2eiV+3cLomb7V6kXqXRD5Lz14VY+XHEJq94kUfElyzIPceTUBPYrJfdttBRu0EI
40hfO17oPx+ojAWz2Ehdi15CyrGw3RG4D/LYPD/ErkIvbwmG9fNguzz1YptdYEDvNGmmc+jluUvM
w9Ch1NpCEtaXJbv86hb5Wz/xT8wUnILPYnIEwI2LezbdsXq/Se9ivJ6zPR5gJydy2txW+2jS9Ys/
S+ALwTjJl9TFtkuyLgBYg9VZeaf+LoxYo43DIXV+YpG3jWwCfMrO64PVsmzNbXLL0q3VzVVTD9Sf
7g0n/fFVbUGxapwLN48SWL5zMsKqdHE7rZggc+aNeDQAGq4vI9p/Mw7QU9ZKBTMzPmQE/3JVFbEQ
IQ+N38DtHL7uhDKiuaExzQ1ZQrCTUGS0BkwL7RlHpxWPugdEvN5ibSMjdBsqTRvEGyRYMVvG6vVF
n/D09LLarNRf6fYNvIcPdAxmeeBKu0hMdw+o1cqEy0MeJRJXYPdUzHKP8SR+n0IgDzzry8BtYvOr
QCjQfs3sGYhd1OOU2+FsimzgN+WWeq4cmkXH5xXz13qF+oFltiWrimNR6759oi12ySGSgIVe+Dtf
DfhRw8yTJy1lsxJrYLhw/072VpFHd3KSx5mtyhSHEopGJxo5M8yFZOijryDPn/zrdYi/z9+ZQ9h9
+tOl9XF2sUL7gI2yxY/LEZJj8IXI8tzQXLs7KGrm/YwZJXVU5vmQruOPZ6Z3G6QDkw4ejOFSco6N
Hz4YmDSLG58bbNFcGbVOr93xldagCEx5cGIhMMvAW1JtE2hWmepBBFVX6CuMgID6sZTSjYw73Arb
Mjw5YTRWJ5GVnywF2kOUHvOB/bXIvUJ3oh0gvG2bEdHbzvmHvLdaa+tzydVU166X2v3drnHXZEA5
lwIDe5Bdk7kQa9H3YUNAnAEINWMuZpvzE0oDF9aa+UnVvy5s4tuCm1M29roF7Cl3SvWjtxWUfEr1
Uu/say0xYgimxlT73pLNfH68C8BWYQFRRDiI24PFWVvJmEVhafhtPSf6N5bj6vYG07+6Gwe1S1cv
evKGfrNRc9XCcUZeuZ77Umc8cRYH9q8kx6JEYL/iLroNORSoPAy6X/5OEqOavqcYzURD1ZnPJf0J
ndT/zFrvAPbKhFGLabnZH7U//ATsklY3LTfwV78spiGIQVCKLqDmFdXgFYey/ASkz3tOIqIByIsW
y9Fc898NFMyzLIVTh5bVyJyjEvktH7TRKyy7nNk35ZmhS6mkKT/LrCMB2xhlF67KzRzf3QjYLO3u
gvTVy1uS7A3DeNxsHwc5tOFZAmVFhMo0zoryUu7oqmBwdq7dOMx4C2F2i121OwxAZD/fP6jUmprj
jGNUB2CIaiysFCDt+4Y6CTn9elChs6mQtap50OHdawGYrol8MWdoC7+7OncvkewYqsv24wSeLuxS
dxyn86nxt4RvXAEJQi9moTEVaTA+oww4AYj3w52ty0QnjHyta8vit6zzPR85Qh24scJMDAHI0DvY
pys9KKSRkAKs+7+/F4pSAl2m3br9RsAHpnxaNNyTTf8a+AroyHP5VEToNv9XyXnM+KGQeZlEeymk
LhdefVWCfupincTmfEAWwavzaT+Gts1MRC8t+VVBoz39HSF49YnWu5uvjf8p3SHbqJt+TwZ8jbHg
xv2lWXL/z1BsSUxvh1VP+xlq8EeJjRY/KBZmegtwzGtSPGV7wHbREWXG56xaMcHAjirKCQSdkGIY
Yw4Ku54fWhpcggnzqz9nib2qJRHq4WIKRerUOyfrnCX7X0Npl8t3Xq1lFBVGZA84CCYj5iTK3Oyo
J5nEnx8HNtvGhft7g17czvTzBWjWksEoykEdumbp7X7kpWxUu+m+e5Ky7mr5YGhljSgc4KJgvraF
/3HE/xassZROWpNEpXxUUIcKmejccLkIaSGqnp7kp3i5sRz0lNteM2f5aQ8QS4rO7u/1vsWwvXWI
BML/3zzlE19zkDuUTVnwydGTRvzk6+TKddpb02wl6RhVBVl9TXcFbVWvQrrYyK9hJCyEteOmERxY
B6dK9S3hyWAFRT1bHDYMa0rj72x4PP34ksldKjUjYRbuFjVwqrRUMx6xBGZYPt6U9Jj1ItdBAoma
WJxM+q0YI5Ewuo3BHGqaTHTkZe19aoTpt0/593NaR34sz7CFZEqCDVSS4jBoGoJxbCjZDYQZgV4y
EoAuOTiWiuEYZpeBWMw1a/Wc8jprZEmPEQl4XkKxWsPFZFWywz8eJD8+/Cv1neEzmqu2G+tIIC6g
Vs7dviiJXnN1eCcb4HkVM5SqnvUj1TxjfYo2CjZ8ZjPrssGAX1I8OtDhZOwNgFWq4FuD7wfUk27Y
uJ/6LCW6uiR99VoLa0hSqn06hUiNCjzBb3rGk4Fpd1pIzJRtny6+e8emJaE7o0tYYiGFy5mIHJZR
WOW2Igb0Apoegex/36C6hoy3yDtOZd9F9TVzoXBi3KQy7U7vRT4caX6WDXttuwx3+Y6rxnrk4PT9
JS2QG0JYDclVRxGByaRom6TnJIWUnzP6BtYfKpyQzwKT7spGqE57hj11WrcFOs7uBuD/D0dWyR+g
chR9PBT6FOM8spC8I1P4LYndpmXwCuF5J5lprwJpFVufB5pq+1SUyib6VfC6tWOZ7WPEmGxCGOH/
i/PV/bbsSLBOaOyFqwR8ScFSe+Lvkl7fnEHSDrpL92erIQ5m5S5ukm52p6AA5rbJEhBu5m9Yb0DP
eGgOifHLV74z0+dBktyXJQftadkgUrF1k/l7sLyLP+ssuCUtZkDZ9EiCYCjcGseEVrFV5b0N1VZX
z5qvChMT76XnDb/ZXrt3bw9dBgx+PJlo2HzjfJKuaJcmeQSCfuoofTcULg+KVKCpCfecnLwdJdzB
IIeF21POQzaIf0//rbgyN0xTkdDx0PRSQmqKeh9xEnOF1yjGTWyNFPlc7v6E0xqV9u67FFlDYood
EKoA5jWfocohQq6CYXuw3jnHKTQjguWTTUPDCI7FgcCPP5uvog9rCZEDNuvxZNs+HIIwFyKrUhYL
NXq7371GORUzruybaI6Y2gLXeavN1tW/EELE6/LrGsiNrErwimyTHzpPlCzWTXQc5TpeNAyhZAXw
U7Ad77omvXOnc7Y7agmv7MtqKO5KK1ttYHegA8ZV8xl69oR8/UZdr9Um3QNpWEeZQf7JzK+ew3bb
W0uux8ULP5x1RqqzXpdm8zUsMXRdCQ8W7+2BViNCBUBZNyzMyaEm+ax37hvUKS9kkCY8uQ8nhZAn
GTkO9y35cEXMp3pq18uudk7i/zab+TxwRTZjoWB5V4TCod+sr+Z6aPojV/+UbWApzypbOk3GXxDO
uA2KvJkL5LPzaY0y5/zJJ/Xh2snkaIrQgltUIPOEv5KuVVvOaSW7syEl7dDeGEbDz2Rkb49k6vzV
Rokg1IHucFI885jUxceKht+kGkHftU5oI+X7C6hYpcwIiM5vipA8uDBWfPbgOAFD7eXP+jH9jwWx
Bl3MJ15SRWYI8aKEDvuh2pwJqtfzQ+9uiZxUmvlJ6GGTiei6mJR6zNjss4HbtoPsXrSGDl6+lU+2
iOX1k7kpASc5TuJUio2Viuoh3KL41gyH+KVOtW1xuaORpy5m+/CJb/je8H1/uBgqVe3LgHSuhUUa
yBJ8nOb5k4f8kfUahpJ7S4104W6pB4eFSpL/bZvCl3r6uQK5jJo9w4o9ejQvy4hSLtf431DrcFZS
4meSN1cmnR4KdyDvHk5y+K0zGGub6egzL0uBXS+Um9vHomi3xaCeIf+G9bxqivt0h6i6cmXd4aop
ZDBxXguckfBMldru794x+mzqgsLyBOEQGJybizKPV89neOjOCjgQNtb48keXANBNPXZ9QoOFqdu9
WksSiSvtw/R13Ml6uaQkf892bY5TNbBF+phE/ZJE9jmaNCVZzK6rjyFaaIjxGMhE0zt2Oc9CqvUo
MGnrjdk0buZFUFZhIBTZQICemidWAr26EXnMBoufO7tbTtMZU6FZRrQX+cyv4kODxo/LQyVIgH0p
RDhkLgaHSPznG2ZwDDDZxqik6onKL7M41x4qqfO3zq7GY1Gx1DaHQBS2CUvX93aw9VqkXgoTazs+
ler7Ph4aa2WP2WO+M47chk6Jf56bcdUPYhWFHMMyt5YypXNaFhL5UzTi5WsBL21IN3NI2/JY6wvp
nxF9vP99kGK44AHWAiQEjDxIyCMD7r1KB+uL62aMtGQOit6uMrEXx4ZXR82GOFTw1OFfv0hTFC2W
FsPFFoImbF+YFuqpBrEd2Rj1zaNFXu409e5FC/7fOmfl9IKU1Qe/E9He8ornShmIXUgYgfmMcIVU
t/qBxyUtVuuHMlyAtK0xBwqYcjG1Ewij2p+tCiVjAC1qwggiDLF8drXI2/u9JoMwstmLVlrktE46
A+YRYUAH5uArH5D+x9hWQgV5AAux8dYytAFJpJo8MWdj62TWQ5QkZ5uOksAJRu9z2t9MFhlhXkto
5hH0Z+iOcvXs1sjmXXsG4GVS0pcmTs6mBNaKSeCfstH63HfqrkZyBSQ3fdWVvFifyyxLgJb5hCBg
TOCgP4a/dcfmrrqYDbqhLlV1sr+3iC9UeZPYuApjedwk1Y2xw5DKDAB9c9QGilb+pSBZ9qsJ+2OV
l5YwE6CgOQC/8NEVQvDbIdI9wlrq1aboRfI1iBiuEwRxqcvpWSo6E97LIzQu79dedZcmhzXij1mF
r57dbNYYE61Fa80tSFMwtjB6kcTQKSLySN7sCIO4zHFFJr2tpxTGDBw3UC5IlpdvcGYI0tWwdA+Y
1n/08SEn6Lhx5TG0VE28KdV4SvEe5a9F41ZGK7fbDBBIckTtIwU7LUUJsvT3QDYOgeGg+EZ5CLZi
VqkUBmPOFhSh+rvmVzVKC+TGiRRTptY/ccsaXUCgFp4m+wX7fTDk+OM7imFsyIo/rG3Ru25uFsLp
VklIosBkm0QlLku61qtAXZGL/ouNBU2hK/P/Yynst/6O6fWRMCDLwZFHtrkz42ESWCh4RWHr3Oto
EFGJAZYh+1MKQ1+7tinRg56Qo/gKuUDgKM4+ltkifEuNYIi4Sw61D+ckJE0qKwy2mCdZ7JVrWrhY
ByuNWofCTPcUobZ9/b1P7K5x4taVdepj9sWSq3C1MlXPWnT7HSScxfgra3ssT1ANJuTjJSvfi6wX
4TKrWHbE3XYQNGkdTilN24KAO2jr72gPFBoyQHorypZypK91hXBYxPljWvjuU4tIvZ7I3SxZWUTY
sY9NlWt9SZIOK06jWSwrJx1lEkIkE7fxKS0p1bur5LaN4rAumtgIpJYpMURx9LoduQpNbRAENW/e
gjvhLfGwoNVVrc/bUOtjpRcs6zVYMRfPxcfWlJ51LO+yZP/63jIhLdDdct3sNuFEqn1B0/EwSTw4
rqZU3DAQeKBJPzkjYaIBRw8cujrYjapb1jdKdYDs4se43ErF9AKTxEaGKEdpQ3H4v8pSzT84CSvo
dnnxnep7D7fGdboOPV5m6gZsOVlNn1u9+qEGWGQzUxLmBgFEK8KUsUGE8FeX93z2dypQF5RrKWsH
NtL4+FgKgyxjIwH3ka4P16IyT8irU3Oregx9cdZEWVrRcyP0BPZOy2KrU+Z9NifzYmaD3oqEGmjg
rePaRlkrPkkd3bdStU5iITDS+KAnr1OJZ8vb2njq5udtpxooxLkh18QEGqQmjuqHsDTORXOCSrUP
gXgFDCEtVzRJIlXCiAb6lGbW+iWGdiJ0YBWoC/Wt8GhpQDTh1hL0taawf0E/1ABGh7r3PcFZZUI4
ww2ErsowWqASwzzUVeXq8JyEhm6flGUIj/TirJXPctJ6j+TdEnDklWHoGtnsCieedWgRCJAW45a4
TlxGuS3UcCxJjUiQyXMuinlDlI5U9S/8TugBYxnXnQlfYRGzs8+xCkjKyP5RjyMv6mYp8i36yin8
B55HtAtarjNRumNEB96mONQ7UJsWX4Hpppk5IBQbRhYCnZuebFMwGx0NyT4D/PqZEg4CnoKk9ul5
zdeVmmIDAOUAmTullE0VdtHRJ0XiDXhcFS0YHsAx9KAteR4SxbQu+c/X/EXSAOIn3rsohEZpL2Ln
OL81ZQNUAhxlqseVSkCsREh7ztcq2HUdBRmt94wsm92BCbAns4bO61clbSNjPml16XRiQ9Whada6
C6FTac1sN5v3Y2q0cCWVu4KMFhBeH++wZ6mySJkD9eDtCHGR4GLNnW/3JNsTzjBFafTFHulIXsgH
nVqmvb3PpxelnqS41lbMSPeTM42/iEySGOVzZZNyZRCYGPKLy34NxwP7xzvH5+sqPO6STWNeuv4g
OIOYgSNeTuPAIi8S6OYz1Z2RplSaJtutM4pEnpGUnfKr0BUlKJfxuS0zJm5Q8JffPDfnI2KpsCmb
mQ5d7B4qfXhESEB0f/48lzxQHL4gaCaVDY06orelZbz2wiaLFkdfrKLSlId9HdiR/RVbzIFziHhz
kY3ZVBLZbR6OHFdRHNZAdfy3rVrqiWLdABTE3Hg0G2rxyFf3QthZyZUIlBRNOvQvYBU69D1HYIsl
s4ko9tkwXawnyKBG4PwXzK6YHldBoV/oveokxh32nRYQd+UQONM5r8cM4RbI4QHGWIBHvzxpfz5n
EHWs0tjo4JBE/6evv21fppJGdczX09wDoX6BmfPPI5h6lbgHFzZySCDfdluiYwEzaPp/PNbfBRrg
1BU+HcPzfymrov0GN4bT71fk8cIYsQxUk22vWjjBdnaEfxGpyVQ8EZPoEbyYqLillWDPueLPBMcH
gZvz1wAB4piF07zwMz21cztqw+rtiLJgcEH++PqaVV37WHWhitmIknJtjSJJrIxV/QpNE3pQUWys
NvzqgnQz+Kvay+PQ/UhCZyMvXXeFQdxDXa2awiZo20ywzayKR6LepMzsYwrrjlKwF+MF7gx7KPNj
wbZr3kFSdoeA8/Iyyr6JF2bDF+So2r7y5CMZMwBu+OATVCUIwwHtzN6qmM8Z/8ks8TVuPI+lK9S2
8sbUah5pliPubjic3/HGFhcPCj/cv1sMDoE4kvDSw43dvvEEG/pLRlb4kO5ODj6dsjTKAvYXzvBb
O8aftlLwVG0tq69wwF8NqA70j7QAnX7XYt35xtk8VHM12D5mZmgZP0KFopQyJRmDDoqhzteGFBC2
rBL64jEfi0s05FYtoz+vjdl30vnF0HzN2jZK7+B2GYzlCRJddM5CCLanUPYzY5MkbsMDyc2PRA2s
5sSLyiIx/KLDMSRZNaGRrvFTiXo1fogiaLw/L3PzrWrxvRXYWNiyfiEEfP52JIWvAEC9lMeEk022
ytIlaXlwFP1MMsEdtIy1WxxuxiyU3I0WQ2mGxrpu+s7e6JKp8vuR9W/X9WtXGjgx2GNvFn6K7OJ7
0MKasCBMvemqkSQ08xNEm3mDGuHd3SV+je0jgA2r5Eq14iswxbypxq/dPz7wYaIIkO2l5XpYW0Dw
TZj06hpFPH9mJlQTtxPHhEkmli0Q+Bi7f2ZzCjQDIHnEOOKMuZ01sBqnEsaRgkVZdGfA+ijuiJSb
14AnVfh9XXkPLO1NstADDPyzGs3qMbL+Bl6sJfuHTDWF3LgARPRkefqi00iDE9joFyyLazM8ScoR
BSZ3T+rZatY9Nbezdh88V6a3ZyaFwK6sH6yX7WD/ooFIKYh/rQFp6GZc+4B4nMo2NdAkhHBL1MV+
s3rDR3I/gd9nXOwNWdZMkYyeYaLLg/xLZtcWStg8tsNR5hVnfow2QLKCgC/Tf9UJw2xdSTjrw6fn
HqZ8HO6oWA1mtgV+5IucyjBUNalrai5vcBeU0DW+sFC1f9Qrd/aPyxMnhz5WTIONkFYOytajq7mo
Akny9oKhyA9VmOVDKzVAQWWPkN1BMm4PSXjutzwZ5OD0T7m0e64RGr+1Htag6mtSQY3pr8KubH51
xQqqUlEA+ozpehf8REM9em4BCdLhUIF2E8GiUqIb7PX8Blsu8o04iEDyaIDtDq7v/dj+iPe6ssMS
CCG/7iq5RSdtNfIPrEw5J0m1v5j9ORA131BpI0lYdU8AXxVL6C4qT0SYSrHnVOc1bXj/A1KIPlI0
3I8yIulHGhdjfo38mTrNTsxzwdP89Jkc80RSlGIdiU66tUjbAtTvKrn+C9kXyR9WHYl1+rjvDvLN
wB0obrrtiKOfKRtlihGE1lyDI9+SNYhF1URaMoAQUJUwt6R7Hvp2Pp4Ic7FLotoMkx0TRfVj4yWU
spr1H4LOmJOuSzz6GQf0Nt8fBU4J50SHLlvhvuIergGaPu61l7mA20xEHc4nWa7woEgG6QiRWEP4
vWJBjl0HzlgiIQg6RYkG9XCIKn36YlU2zTmKJy0Y3HomYfom03c/ebO5TWHidI5dndxdmukoHNNr
T91BF+SyY7Rzx0YqkQeIa2isygMMiHmd6YC4a/tzKSplgZr1CGGa4vzVH9yIJpDWf1gMmyjWbraY
XlG/VMG1QHpkrZ0kGpaCsbKDNQnjLJPi80Mz67whnsa+n3P4wW0VicZZhHlcsX0lpcs0bGB/BRzg
XX9SU3A8nSHkmCsxW/TChWs2UgXn4xF1ABZd89o4ycGrTj+9eK2OI8K2PTVko/rjubiQIPsO0LfM
WXB+fDf6jj+rmxOSN98mGlihoaURsZd95C+gUZR4d7YaJp56YeauoUjpLFsueSnaY5TU3ZZupt0A
jFWlCmuc2bFTmIgoOGGa2SK9UaYcM7hthKOZoXULkzLU1GIzBy66di6+dYSE7KeDxnT1Jzlc10BU
8XnWTK7PbN+WjrhdmNq3MBBvag7TjIPA3Ngy55aAfj7pRc35EEaB9W672lp24oT5I/gj/PetihBb
QGEcShRZLtq/a9wYrak4w13ZIu93g4OjOslwpd/h3fpi4B6V3t6b7NNmFy/xCoqmKU/HpEI+MJ1F
c7XmX/zE20oQYwUop7wviZPN5GNxCG+pJfNTiphPn+Pf0KHKcV/FGru5TfYSyik2WM3ZIdvXZQdw
7i7+ghtDaHpqH5/FcbFBC56wJO6mt2reewKSWwrHwvxXrqeiUtPiBglUTDRJisVuCsnOU3M9a+O2
4X1t4Rniwkd0JmqPMYPX4h0QHGuyEdEzOSTIrIMBwydmDiYSs6ssKBrMYybG7k1YdGSyhS8O2Pii
iJ93oVUpwVI1PFAPj8zEvDW6kaDnidFOBLY8QIcIIN3CeIA0+Y32lFQUUD51visMAgi97oDeGVNi
9oQRxWPSq1+D3zSey+pQqw3skfu+HmH0YEvliB9ttL4jj809qpygBjh56eYfKJ356Qze3IzjoHL2
eQox6KxFXZxGf3J+00VNQea+SGTRfitnYoX5uewCSj1E7hkdatLGhxJ6URgg3mnGQaYTphHJLdLT
jx1J8AmqTdVcJwMwZNBdwNlfvPuZWQEIU2DC7YFHZFpXDZHRyjw8SUgM9KzVh4OwcOBN8BGlWAWq
Gpe59Acd7YQCbDelpqfPZdcur98WkOCM1bNxTBbkMBkImPjBx+FXbUiz3+p2dl7kyv6CD+25NExS
dxoiZbf3FbFeosCF7esgjT0mzNn8S6usyXJZHm3bHuvx4mwSV3reBqFJ9N8Yb3yRHmBzblTHPNKu
OJg/+xUpT9G2KDBukrFCunB+Czfn6UKPk2jK8dhQljA1iK//jpGzMwJrPetEELhZbGYi6kSwzr6X
mhZ30I4h4eJOO7tFoUEh24Bhnn1pujVlZsaBokiLdOrLRXyj/ZUBSPFjYu5FNUdnBK7mQ9nbIIsE
6kSZgsi4Wre+auMb5ZuauefSZflti4qWWcKpSYUDC9wHZGKRGEEea2/9m6T3QFgD7/J4jPlmt2aS
QNFdHH+Npg5NRBHkgsdxNgHYDFARsKVa2B8kAoyo9vSsCQE6XYq6marUH4F8Vecw3iJ+nzzJUh28
coh1JILvmfQ9ClR33X3qmAa2LBi/NV5ZNNAQNpprvayck8+601CYdsXxC61lCxUqI8LnKoSfBXjP
9dF6Gdjr3PkynYvvwBtAsgMihUvj4mIwlWewK3jxxg8JmCp6FcKA5O4MAFmwkYa/mQVgCjZCvjZr
00Y5//5jGutnyC3/ee6TcB6iTb20PVyYGC/PQGPTZfxAViucQMPMTlJTwyqNWbx/eB6afgn8weCi
crv/OzX2+PfsqWtPMFCrldrjlojMlUHlGFS54WNEKP41imiRbQy+cSeHH0nfuRPuWo6aCrWMmVvR
w7MRfpKU/xcohiqu4kOGT/VTZMkD+7aR/OM2NcqrbJvypM1FYUwfvdCex1Q5b54GBJ3DHZgOeWbM
UaCbDrB8R7sKskdJpudKiTlQyOt2EBXyBQHxpkpGQr7+hf3SDG+icy3nC/x4bHgjdFvPa0O68QSE
sY4JM9fPixLB1CTq7eYYxXER6T7iWPL7pgiQMI46HaI6hO1pyBBr6g8Ic7nDH1J/V+TA+Kvq6We6
580KaBDufV7tO4LcLLZnZ/bavb5Hv4OpLX1x+YZYM3MsR+QVlWFk8/n/ujSN5j2BPXst4aTR5PNm
KaBP10wm89dmXvJHtetaAscVu7Y/5KHB2ZTNvB8M7q3j51DYXtGbpC4S4d5XDJz8cqDFAeAvE1V8
pXxXG22bgNjLr+xxVGbaYg92EcGxRai5E4qc+nj7q8v9kFIWEoMEjapabKYiBV9/jWs/wpKl/Ixn
TnBmLC4AOn3+88AXz5foj+/3ru6nQ5zzm89TLHkuDOzg7wyXAE1mcBmOEypzkbPKyk4Bpl0apjvK
aOZd5p2TE3H53is3cwWfcRKkC3Dt9ViSSkbBJCVqTTfYLslMtDhzrU3gtyoxqf478QnqLF8gnnbB
Ec68+J41fD5uD4I2c7pW8kPdy486cQeIMluwgsLNFs38sJh0+dDufIFDod1EaUgr+TJ7/wlwTiUu
gLsXw+x3YZRpiva4cDOG/8kr23LNw1fO+9iaPub8SHirMKgvDbIY6igdkcTTp4kiJhbvFco2+U5Q
htCMgyz/pkGVvPmIz0brACjTbZ58cMTupTcN/aUhZPw9d1lcuID0cgMPy9oQwAlT5yupzTkiPV9U
kItWKclNUWh7IENWyunL9AWtayD7WvWKI9iHcHWAxSxlOiGOCMmdo3ZhgE95S3V2O+udaewX2WU+
bgoV4/cfl7sfoVOSp7UA55+eT5rDcKx00IDvchWZITQfhBvVAArF1tCW6+hpEs8lZG09wuR5l5PE
nvNubZidlO+/XrEdB9Ya3Y9pXhCKc11BZ7G9ZNnidlaAxhSboK0dG8NAp/1uqYBcxBP/E2dECgGG
9w+pBPzzjumCFJH4tBpOIaRZzxH9wzbx/bP8F0qtjz6sJpZnOO8lbHP6RF3RdhF6IggvydTCHDPI
dnk10JSzj9v5pL5wwKHMwt5pmBEFPzg5PI76oJ71Ijq9aUtexuJWt33YcKbr+xB1HnF5gg14EEwI
syuQ2yRSP5SBgYSn0LS5Fl9LIZLF361lR6tGLjNP7V2SxVyUCNW2V0GZF3jAuUw9vsFaL69a/KW9
MD2RYsE3JMOcEb5R5VfuOHGfY4faG6hcVhFNoaDOJn9PfUpgS+xJYp588WE1Nx85yhBL3ofmbA6F
UGEWQlTdePRBpqrjhG2R1tV8fknLhrAOhBOEPOBhA+T4P71+4g4QJMXT9MzNU7q1yhu7n5hAi53H
czQ9iiwdX5zOyWoJbdt5vCE0Tl6zDk74OR0u7zExgNSSsj5Ix9vUA5XhUe9fO6ozRGPHiH7gkzKA
gqTWfqOulF+290RFa814H4b8xR4lcOJ3fElqchpHkSeMBOJg+45bULsFxnHhmK+mPKHH/oAohNAb
IJe2LRNyhYgn2zaffmtktezrcC8TrzgLmECgg0/pQN+//9bDvmhdhlcrEkXliF2l+5EjiQm5cp3f
VzOqTju9TsB4T6UCGz+Y37h/4e0YCNYywNodRPM58XdL08w1XYA50X0TbLDqhXZWZOfn+vNSxUZu
suRtSBFCTOPlUW4YXUIsY4HDd6iwxNTHBr7/BMJGExmdrhTAW2C2drSa1yblqHERu1724xUY1Qq1
ZpppBAgUCgYeMnwk+PHrdQfOupaZrEcHXgx7hjdLt3H7itk+uWJ2EWFvpwYzR9jnRllgv07PkVEt
iLj/eicDuINS0w8LUfEscoOWdlZnQvsPmvNwkPP4645qnKXexQw5D+JCT3OWu/a+nQp4aqkHhm//
GHa+b6AoS/zUnOG5SasgNF8BNQ4qhMw8UNEwvuBJo6XW/OV/oNvMwmn0xtSt3TpmrAqA8HPRuhye
kLihMIUc0bD9pdghnOyoRg47bxpRsCmgf7/QzEjM70RLHuQuloH7WoPtqyX3kdpwbpaH6ENlZBzd
i5v8j/XUA1F6M4RIDedm/0bwMuZpePMyTAx9GI3Q/ubXHqRWlJ5JWeMkHLm22MBdzuE40MwG5nmz
5trYgUxUP3SbwTpFBVW/Ene7gLY1jt89a+L+FcHm4/vtyvHx9JVs1oNx7qwykQf+0h6j684oLMaN
auE5I9Ak91YdFEkCXJrDA4aD6zT0MkL9qgd9TN4TJ6u6zXt1XA/qXlJfsEct+dbZ/J/3LPVPbBRE
ehfFYp2i1TiR0TPZiPKRmul4RWGIL1Bnk212Jg4e/WKzl6VUF8+chUiNUV3F04SX+p2aF38Hz+Az
l3q3QZcMugfedrpIj1eZ43ADI9hTpktFKTSnayJ7vlzWkjayvZzrdPWEgz8Zd5QJXWdy6A1sOknV
cB547ow7313KV2ECt0PdPW+fTkbnEyAIzjXHa0ocTgE5shFSFVPzLbtOx9TWDetG3z/8pHaMkRnM
H78A0/M1LKuk6vmvDS3XlIDzEB7hofVfb/j+E9P+6qoWzLOXnq2qTlca4Q51Xm0cjFjrFtzsE/vM
PTVxLBzb6HyKVTaJzg3vw4voY/d8r5IY0Sv8JAsPsuOKjDb9WWmcLHlemG6IS3nT789PexSYb+VI
Nzh2c6So8As9SpgrkoduVzYKnX8in99RanZojLh5kOa3rcVEPOFYrJhdWN/3xYC7Zm8ul35obe4d
WxfqZthnvO9VmoXrb2lHOfstknk//LYNaCU90/Fc6UzYYuCA4PzAQCNxwX6TV8++R5sCJf88ay1D
B3aEpH1gQ5yjpUwWv49z2LbTv8sw8piDCLaHKOte5UD/FT7GkLbeWtsOJBJMEZ4YZIISKAkZO/29
FC2Qjjt/HHBPnz4UOTvR1bxxz+7/E1RWo//7nf2Z+vMIG6WcUy5zH+SJ9aT5+OqKmxPQ5KBMmFvR
QBd425sCI7L7GtDskzknRQ1Fkds1H6vXeua63IxI3bJriFT4UeAd1JvDinjvJm/BGJP4022MYs3O
1bX+KMEljxYJKd2lq1s72KZf7EBEM2DClfMDfUrTxwTleONOeg17lahtYnTvXYkRveA3K4o825Op
5bWW1/DvpoWdPMFTmm8AnBJtl4/E1gSOBxBlz/xpmBEQrTVHKvD3G8+viXJdejixPTDqCPsR3O73
5CrgG3BJ0xSx368irnFQLOcRfJiOyI0JL/Zxmn9ylmvOvkdZ6qJwaGYrsdb+fHm1XUjJ3biadTLr
TMIjtspXw3qAdju4dGFooMR3FSUfjPMD8ysPGZxRao9D2xcZpbAK0TzT3CBwQS8NEArmAJzPiYgj
85H3cBemoo9lVqTA+zREyksgd1c6X5qb9K+kafbZhZ5XEu1Vh6PMP8UxujHOhQRaCmYeARSpGc/U
J76AVFCP7K/sDBexG4CQxumHjyKnFl+QI0mYAUhst4QX1415/+XDczwegOBLQd62dSBs8k+BfeQj
7g6diQm8tmjWkeKwEFPProEkeOsb78+MWbi5CZiz4teMnaC+dquAb8Iyb23ZWfAfo7FYvHI4uaVD
BUuaTEBlqfjs8TmLtNejjCT8NR81PxK5JFgGfJIbt/n/Dkk9SXTad996tqnDDCDfHe06b/fmElEh
+Le9XKyHFhS3Y3ppL97CX4jFdwirZ/r8u8whVwgyJQcHx2YuvlNKuO41vP2nJwU0iKl7zen0/v0N
zPDDXkRBuT3wvCSuY6dtmu+3qHSlK+EGr+E1N9jfJVbl4njmq78pYZtOhVroqwxoicMxeumetxJs
qb3q3nPQroU3iTu3k2JBqmV95SZ0xe9g0BCfFa4l8IEnXCDqcw4QFtEDOrA9WVxkK0TgMHBzRPyB
QzXhbZ4YqoV6KH9+mgKDoNkIwWwUhWwCd1R2HuZ4aqLinASMYiifCIyAZ2aNhn+ytnM9XvXXTcXI
Fw8+RioqTONYv8jpQf87pHlP345dQBwcnYOihdMAUeMtLAiEP9XKCfVwcGTeYDJHYKfBBVlcMX0l
8vez0iFcZ+bNJ4p1LCCrqHE2OE+GSPwYJwPb6e0956e3dDZ21rNXfI+7xjO1cVyevTmhd5vsQG0v
hFHn9vE8A+pLa53qiRjRszvildnrZptkCMNDzCK1ebYqNlIOFC6EEV65Ep4GhuYJK/hJraE77HOJ
/MTLwEsomMlloSCA7ubGE3zB+cV8N+XWquMdgemLAVf7L7tcUKxQfSeL9gEEU/QH3wiN27nj6602
QusvCOcEAKMaLjNjqsRCzjfFzmORNSZM6k2Jlb4HzIIHzVsP4hSUJVHZ/PLtAKlXYgCeVj4JpFoU
0gvsvahT0+aR/LNCKP0FLnWtzlhBEULUXUpMqmBsNB4PFt2c6MCjn4ANxzw4rsHta9cRKU95C9/6
st/KwH+eujBlZ/54wwIYiPG6nynEhVf+m0tTbealE7MWMdMpJwGk+1DuM096n8Jj6XVxY10Imqei
YrWQGZCRVzpbOZ3h89SFCfiAfn/TKw0cJXaVO8zTP123J2uX3IZI+drtn2OUlrAoxEyaJitopVY4
700g8oIPxrt53bSY61QGDvdmFYUjUoyuKyZQAA9xx6ITVzxERxOC5MgaRzqs5fhWNOrFZ3wtVG3E
AFjRep1AQOw5/rC8kS2jFApW1gI0JZKoO/CX97VFud/qk7PQU4qpULgFl8KpLRdfkNxGKgBzgMrc
lQTSWcQs2APUy/PYiKPHk8Pz/M/UhqT7sn1bmx/S2BY7qSrEyqbIrki0wzNypOjuw2E3X/40yrCD
feUepqzDaXHxreWkxhLCMlkJqrKgnHnWWkUZdz0JDAcZCNKoBeCgfjWHhLvNW49K+0IvycDvad8C
4Esy3Bj+xOunOQjARNVHrswyt1FBDj7Rbx/mZrwWuEeOcXb75JnxMmaaUvQdy5+8aHW8gNPz/xLQ
K3BirQkaiGjF1Vl0Kp9ijKA5pgTAifwvMV1XpoxqXqfSjCgZOx4i6dCH4cQL23aI2E3Hq4lQhtCs
397iVu2cQP1qQsWEHyNbdVuvBsXisGBtQNC81ucZ2z+BKWT3zF2W0p+PpnSF2anY6UJiA4GCp429
cDXCB+ryTEejbxbEoivTB+tIov5OeZUu7ozK0UPyCI20oQ6MFrVX8EQ/8AmWvDVr+Y5sU8Bkdrjz
h2vPekvLWGjeDuhfqgH2pt1OpGZA/OpPhOE8P6SVhIO2500H7PGZm15G06Vo9N1oebr8id/sop8N
QzOd6Cg7lV/uWiDIl+aq9MUpyzHoNTgieV/ABY/AOkjQWOAW/kwQabEMBuezuxbrl96W+bMQ4Gtg
hjhAUAN4M3qRFl1j6Xhs60L1kFh5Ilgc1LP9OS7qMDyQ6A5xBms98EwZN1Nv6yYIYH17ECjoWGuB
UgL7aOsQ6NjiR9muBFl0HcUUfsIi8ja6h/0qpklqLCraxtn6wxqkq6CmUnIz6VXPy4oYHpoTjq6P
MpKqLXGL2L1N3SecI6H9y2nvtJl25SG4Rc8jHsSz3Wa+lK9jqDIBWYZNF6/qA9l9gcT+2pOwvcz2
EPcQRVeaUq/zhj70bmscv9UdI5kCSsGjTNPFfyk2xJy5pI7ZXcDoBiskS6emQ4HXkImTmZcYrWVo
EdJKNd/oVK/4qFVnKQsPfEeVphav4XGRB172E6rGKIfakrr/eYyTe5TVexkR20pXxizmZFSkYAUJ
cAY9mzCAX/2v1kAJC4wiWyIXRkQV9DetNBIVGEMupr8DwSGRt7YSdxnQ+G2SNDBhVDd7PvzprNkT
Zdq9eSjppXW1sH999DsNEL1htOYNmqrCmWKa+OAVSjDIvMEL0M0Liyf4kt0RgEZDeIKDakxqtqep
bYPPOjlin19qF3ul8snk2JU0ApQE3BP49SQ8p7Y4kjihe81IOlBHAgcKX+nehnJqhALZfQ955FsN
CyIqz4lh80blf66Ea64dEqvCbRL7Bb4wC5/5t+k15Wn8YVW1+Dj1UMklU8YJek3lbuSlB0S+OpzQ
xDCW7WgqUoks15cP9K/KBSxq3E2OLXDE56rUSFzdGwArtj/MyPVEOvlY+MEpOqcJaExc6bn5wDhR
zfAzg9kkDDQEJnjpMK+TApRKpC0PLogIIOBR7KZcRhudW+Za85ZQ00WmKl5fBqYqvWEP/WamdKaC
k7eMnjTFFFTQQcn40nN5nk61XFzqLPZmjxOvUeEURTzoCrEMbNTU37kDbRhRRcpVmqW0LigPMCw5
bNsOk7CuWHSZrx3r55x46tPQzyBWG+scPFWn2TSKWJyLiC8qFK8Pv8lq/Ni3dhOUOKXQJhkn71ZO
aE0J1GumgqV96kCL+FDAXUx3Iotkeyr5Bxj2nFKIpW70ir2YejDcrzYCMjbFWcDiWZL+X3cF+a52
uCAHr5u+h7pq3me2Zhfb9Q4fFLHnR8G8ccjhZPn1Nj0U+2337sjyGPkQYFeKRraBGOxgs9Lpr4tW
HBJBJs7+YOlf+CqDtu70dnzxp3iACmmqCRcpvUVxPqgdDAnpOAqL5hcGx+5LHOxSecAr0k5+VM3J
6w3STlaqwltOn8gMRhwDeYlnzZluimY8k2RMuiCNDt3QPD5+NvrJ1KWIW0jocCmlpiHoKwlmZBpU
pSdGfxBn9eZNlIp2H9sXMLpCW/DO1YfeHFxqbqyoI8oM/6qmxOYrAgoOlXucLscDiOP2IVIwfT6S
bt0GRv3DGKumPGYp6dAfWJo89vBAzCeNZb+ccC7vOM1OpIQxSakfkOk6crIQsH4jCUT2sD/o2Wq9
ssGdH1i8s12A2nSoZ0fQK4spHhY4daNwJw83cZBSX010uUM/risa6vht4gmm4BRTYZpvXV3AbUMo
pRoRsdyCoAp8ah1SIIYCs6l5EFXR8BNbBl/M9Smo/zzcQS+2kaxqdNPZ0ubLRzTVW196Vk3n3jhl
Q+AqaHy5U7Wg/t4CdGeZZkY4tvu0mGCxJgY/ZO4olzGAv3tNZnbuSk9lJHv5NcCxqoqyOx9Ua0dA
1MrdaJEG6Q1qC4lHu7WohbGkq3qw09/XJ3hF8TddPW4AP95A78k1RMlcEYZorwKbmrRikirnd47U
SjdL0uRq1DCR6igRBOfnU27dVzXddhNBODsMA6icQ3g6JJT+/OwN1hNOLGPKWkkK3RHiT6NJEOQU
rsPmSH9KphzciiruNBkXCsBkK7ifQtY0iR9uCZer8HLv6pUFnQlZWcn5vckciaKJu28g3fLBh5uL
fUOTHBzormZ+w+IqBdk4y0B4wbUQcysNl122P/FzIODJwuItRpqKDrWkfqtYomPbrkrNAzKOk4jv
DByrXA4LShDg2R9FPV6HhVcFEQqCANmLwL3cxjs5mZFr6tX0j82Zo2+q6zKEfekx2W/ejmdPeRDv
Xibkj2nBk/lGdSgVwVa1wYdREpGCP5roiKBDRvT+Iw9Q2HDjuhp5UVaJiO8tbextkA4G9porR5OT
m7vCV/l6fizDwBciXA/h1U02PFOYBWSa1olfC9Aivk6GJuvuH3B46MBVyLG6RK5jYK4uU6oCuf+j
BXGj8OnASY9kHXsYQ7nPcMaqUP3B9UmJ1dh0kBGrZv7KPwxYAhLpgEJDkVkj1WB0Nyq19pH589Dx
HH2gCUc3Wg1fewgWUo/NVAU9PpoTdlHAZR92mt+bsKkV3UCAyk0c9SmZCyubl7U8WscwCbLNyHpN
TebLcVxPWBQ/kXV1U9fdYXVTW6Ia5UFDUqIoY/rwh2XJNrnsw4q/oEZJSXOGfq5xFYvqmTTVnVBI
2+WI0U5Z23ZS7nZJthucFeBpUIU6+V/PI0iDN1Rd0rVVzscaQz7OS4Ic1t+EMa0L8hCZRl7a4oRb
eaS0klwFVe/mMtVq/sPtCtHj9F4uhNqs/d7sdTZISVCLXzMyGeL1l2g0OWsMcm0+BVWbYfSMsToo
HJtUhWuThv00Xae95s5nttkJYFJR83vYUGyYYTE5aSGzMXFOIOoNq2Hzscm4VReo8574V9lFSNY1
nhaeOMPo12SklLsFyLeKRNUxP2nukTQZZSLZLQGuvzJBU3dJ1dcqGGN2TpqPQwPjOZtU3ikoZMT9
9FGf1VB77d/tKmkuuAv+hkTEJp+cQbcVE5cQin1cridBKim+D1TM4VpGlwdwXuiSvU0JxQgJ/vHq
PGc07R6XUSJP5fxp05Y+eIovDjgooKyNpw10gAKpX7WUFeX+ovLzawizPwQ5/YwssxCA/7xT5s2h
02AGKrn9gdHTHvDsTPIM3iIm09+5BjkviJLSdPoOO22k8GdUnN2j0Cd4cn7DXc1gRa+C9gnIaQ3s
ZMwD1pO0n4/ZOQr2MFxK6kJIIdyYuYIGmIUEE5ncYnM+ZDbpyONRjZyVmBensl3jXcIgDaMERG0k
VxJvMXhgSHWfoZsUNsHC5nfZqxxr2N/84t9+ewmh9yc3gc/tMESttMkprjQPKN9KPy0HkLLWeyUM
YZAIkY9FjamhaG3EJPU1C13YRNApRXfN3ihPVVw1ZBJb/ER2cZ22+piQ3CpZ1jZ7wAC9qjifZFYf
MwrrHMBYE5rL1M5dE5Ea1wptCCVBgrakRIrKeASWPzc6airmy/W83MJf+beiWyKssYk83NoGai0V
y5E43is+p59nZlLvx/cTKTjqpq33COwbzD2Sg4dkdUQTJq9u6IBhUHV54q2mZ6jb5hDBbYCEVZ28
NJKKZgfIYQyg/KyYveu1X3CA+u/SGu9POhkogc6M6R9bayzKB4wp34/kIO/qD+nRdKcvLJfOyCwa
ohj14M/MMFuH3y24FBgaRar68JnjEILKguLDObRdSZEtomO/My2K5pIbSimPaFr9WmHGVRRmQxzr
8a9fiT8MX2R+RSD9gETxEGn9caWR8+knVU84nS8MTa5BLvBshF//258fejDwe+nSFUyzgPZ6K6fi
dJ75zFqJO3+PXopj5TSMS4QJ214Ha4TGg6iVF91olGHmlpPy903EppIhwRLRrXUrEXfFRDq8Bpkr
SkWPpkzQips4U/gHm9IlwV3/G4dIh34SaV7ozQUSlDvLkruGezdnGGzcQcuQCFcG6eUz6lqmaqwb
pXspJZ4s0F5MkxYT2on2C53EDR+LoixHa9TIJzlkTojQb/nYzesqCou//VAZ5munkQFHMOiSUKHV
FS96+UlaOgPh/oWaS/NPLZCrVg9PkRKTeaduE2ajVFUqZP9sysdQJWVnvhKKue0crmuOFg2/TkfE
kT4lgFln297t3xeJVn+aObBWy8RfBUZuqTNGtDjjoc+EM0WdgG877AuBeHkwb47ibttvUpn1ago4
PfHoVJXfMCQV44xK+Lll/L5g1ngx0crvkC3bGiQNpRoo/YC8Ng01B75R9jQEkQIosEFhDrmX098Q
Q/ARWMrghdnuwMszCHaOGj6zyD3mu5gwTQunBCS+oEpkt+eJ45meaobujZZXosUQSuFXCor2cm+0
NRe6WiwlIDXK64Oa8onlYxktiGMpqPP8HccQLiH8O7cCDEt1C/AoYdGpiVacjIqptkCZ8D4jhHBq
VFNqhu9PJwtSUW6oK0wJ8AlCgLPUkvPdrHntVma5j5VyXc5FnQ3EKXlltP4AVOjGqLhJpanfC8qK
6gzvgjOxgIDQgQvJIkaBBzHT92Z4GTYbv46FTFZ6NUBpNloyKrx/wooImRTz/QTCjDBrA7OSQUP3
4mx3+4l8a1giqdxq1CXYOmOLHq7Yx7PMIzxsJR9THDsftOZ++AifAZQNi+U9/QLsSh+nIMzujoVp
boLS0/R+2E0Xu0Uk6oKNzLZEdDNzfb2/QGjpFrxO7j8QWR93iYdFuZFNxzz7nW/17th6ILbV/bgh
MsIigqZ+iJ2bYbdSRrPaAZ7//tKs35R+GNRZEbQfW4O6KDOWxENHrBoRV21Z8ZnY2xqCXkO9gSAU
8ZBSuWOsd4ubUqT5INPANr9uumvQvdnIgojYFctp9azOU6LwKjgwZyylL+IvLQaK030iiqgDQ0z/
PqCAYMNzkFZfcsX0DT2yAPCqNentvMFFImird7OhVHssvy4Roj4JfssUMMBF5L8gxuGdXvyivwFf
a+XckiJnQ/wh9JHkRMz6g18im7sOC9qshIZboNGwH+1JIZ9LlOa1IaG/GeF+z/hNHyK6E32xgNIV
vTAgpzDvolU3Gko30pMLW2wj5RYcQPGSf88tc4xc3KYcc0xIc65dmaG6Hg7JpJxH92JYBjQAhAiv
IrzsNWGgxSCd0mNpjPBeCRYpp5N/RsGx8CuKl+Ewx1MVX16d/yzw3JzslO+5Ae2Y/TlNPDEhsWDM
sOvYHsqpy/KB7hsP69msq4dgsEKcTpUFSYMbX60nfBRuqhw91qnKG1yp5OxvG72qSL4LPybo+rWf
KSyrcSWnfXCtT0nwCigBBRKj7ubbx8IBfnaBFwvyfcCnvHBu6+AnCX3TtvKttbs95dFLbf6RgOi1
7dEiYnQYwtchqH8ZqLhIXGEiD5WAVbenlYa9EyJ3+ClCIQ0uX15W2OnGOgQCapk0IkWl01ifa8EA
IuxcCHCGDkG5RI0XgcM8NjtM/C91+kC3lK5FV2J/fbKqDKzgT2FVFhdURp2/3ewjMVavjLRhNr/v
ecUZRwtgVMspkKxkCyyu/X32AhiOenL80haHD6ItvA3uG+6IpMhy68mUtDAWxxFFsAI9kZAbmHkO
KoqRazSGg7N10e4y2ergnmqQe5JFkwxpZtL8vNo+mOFu0CEuBPo9fgrx8/6nDV2exxGspGDFiA9u
XApwsJQEv1mAX+J8gtFB3NRAF2dpc2ngGHsJW0S1b8NLFvXkd1aYzs6hQGr8ezTC+NCPSvR+LPTM
os5R5o2BUAfVKyWHV584ttvKhIv1a7CT7m9Rf37VAEFuvPCX333nGBYWKbqPwzi9sOJCnnJ18+yt
otLZ3ZHN1Suy5OrBK0VT8Hfq3AJPsFMEwxUjXM6URYL3XSJVz1knAkGS92D162pf6SPT4AsbPfQZ
PM7rfquBEzUISZRql7S46Ixjkf2aMeYo6d2dLzCFsUSBdbc3otM1DlKSZC54zyBW8HlxIScRtY0t
o+qSdBNAZp4sqxdhJ+kerP+sFKA0PNXOmVWQ9Y0mNpRZHvKR3Fz3928l55c5y51LSqppvL4pNtUa
DVMIyplIzUcy3WrFkvowJHKNwTNWh9Zgtj2datn8NPHJZFC7jVfrMVC2genCZ7Kv7glReCbm4Vbb
VQmyTomJJKDVt5+YY8nrweOLa50OBdEl2uGo/udBBsn2gPAVfeXnxfVQgaEqaX842yTX6jtSegSU
5vd+smhA/MepTtPz/AHr6wH1kl2WSxfVSsz/OVbYwxk1ufXUjC5Xx187bvtevNdz0FQFimN4F67o
VBuaHpgiGaa3gnm6G+6f/cESVQMcPPyDOxHbi2En3V7dAK8OU2+cx6wxRoczziPivorgB4NOzDAf
pimEhJ1ZivIG2J+cz9YQILG4JyUzGD33VxdBl4rqN/TdHM/YbK0+/aseRKmt6H4+oBZdVGa1NalD
fno7/SreiUrddwQnmCIb+9FBPXpeu6HvIeIhi6Toh9Iv3Zp3JzJ3vdau99Il2AsDQzVKzPcx/Sig
KGrA87ILIozPopofX27G2h1xz/8R1w0ZlsQIejtguxulZTqOxBgs73/tqAdaQ5vCe5Ex5n89sEOf
DeWtTlH/kzkfPm54XXM7kh+N4e9OSb0VVX9c4+FR/pg/YdkFS/SL33JpFTILUceHs0CDV8/P8KdG
1jDNRy7pF2z4hEJy2pnIRD9EbAxPS6kdLagzOx+j5sqPHCt/rL8Zqi5/x0orUlTc4S+SbeQBERu/
3Nt3beegXJd5wtT/15pgbt2ogc9Lz5U3NLpkUIlw1C6zGkO48b4qg/mGON73iODNm+oXW6/klHrD
o4WNtflQjPiiRFR00Q/sFXRnI89d7PYLb6LvCHQSbFyv0zAsKNUr8bYX4BgiWao5Zac6Aby0bTRM
BpzRJNeGZ8KZNY8EDjA1GKtzwi+mB96jR5O/r7dmr1/QAFdite84i162FeNNPapD8ylYi7lpKNNc
FHW7ExQbYy4xNVg2ip+1H5lwcLWfemYk5lLpcudVuK9q8StetxAdlfs3ivSCmnaMaFE+xeEeVS69
SMKrA5SC58gCbPbxza/hOLrzwfO9z6ShoJpDYW/uUNCtGpacAn9ZBwBPPer9qznVlq4g39Fol7fm
hqn26ERolD1iRAm9Mod/aYQWweSU6tGFLHIhue09NR7LApMtUJc/eP6MkI92imkUnQ4PNODBdK1y
GwJ7DEb4NNGRSqowVNO7g66gpJk8SvExgj42xRSbeCH9AwGNjc4PIWgwKN1a8a2MDbiE4fliEyxA
tRu0UZkwpOcsRLblShCuG7QlldtDGz5mQ94/P8JEcnr1ep0R5H+t5Kdd92gi+2NHh7j4KBPYSqz+
1258pXHeMFlY1FqaQWSEEfWDmavEcmM6yu8URDv2rFr0CUzR7unA4UOI/NV7PUmmJvpNgVK2Kz4T
LVHB/utfMH/Acj6Z4tMT6W6kuGamIF7Pqj1VzititrexuAtBnlw9LeHT9z+qYqVdSYQcY6Yb1PcC
XOMc6dshAKYJZK4vNoo5NAvV6OE/dZOg3WsRAvZCuh7bAVEEF5Af5S1dmJiEJ9pOkta5OWVQy1wm
dW8QzUwk1Oc1kMl70uKVVIy9r2/aeOtF5HSxc7+xNd0FAWhOFMopHypy3ad1AtmmR2STkFfe7ZGz
zB7Uf51DjHvd8EHtYavfWITWxPD1oT2KDG+PkNvnoke0HuSwh1yTzeSyjVG8Jyai8LCQbZi9s85f
NwZT+DYEBojPbDSu0tMta/EAYj6l8tg8xeHUbEpUkLf+jddTBrBiJHXOQiSEq9s0U8TZtoqHJbpx
1CypmY63YNJ2iqOWX94J6FYa+Jo0mTI4Xd0GAwW2VoPl+a0Ss2LU9pM1cE+dI1T/B1ULJvByce8n
U19h9EhYUJ2hFM5WsmL9pKA6CmOAKCs2A0JPanV+TcnVuOZGgQ9dgHOA0MP8UtSPqaz/AuWg6SDA
z3mJT06m43w03huQ9N4p7D1FuZyZYk/U1VHMI5d+0yXtqFv96234iKB8+13NV9zGwxs9baUf00me
V5B3BdxHaspkviq82kJMCtsgql/e17X/pgj2a+CH1kRWuuMaQ09aXN8dMT0axRfZS+Q4qH+3f7LD
fVh13PhqAmkJCJXEfjfAI5Ot3I6ZOnwxomVHShetH3DbPmpZg1FXzt7Egj88MSwlIbJUgqNFTKDy
4cPoD77WjYRXqXFvkbdQGMikaEXNd7gg7/x4cZmGsRRB0ub24WOnr6ifZ/Xvhx34kfiQDiv6GihO
JcU8R6Ctw5V7Vb0hdJPYNhGcg1hnWsUZGy6eJfpr14OAWb09yK1j1+9FEMVWuaeovYy6sbIliSyl
/wjvlsswUAQiv0OXcxYzISYKOHCwRbwClhGFVMA2X5byoLUV5Jou3YnF9VPUdg610NdN2TcAG3fH
PMpGHFIEW9mmABz3ro/c3R78tz/JYX3xU1Ehf5WfoG+kkaGd2vfrX7P1PwXpDgGQoCWtjsKduwhe
lsIG7niS40f+YEg6/epVj09epYhVTUDAcKl2VlVo5Ye/g7qrWMqo6TXiy1i69Swwy4kDd3Q04CsH
e2NMxWh1KJ1HK0SFmDl8CSFjWyYOsJBmXBAK3G2DopBBBLG5BQu6HFSIudT4AzpEc8cLLMP5vM5A
0kGBuMx/u2qlSookJwcKVj8FjZZAQ+iE51gDc7+xyZohTvyPGvWVbnVqxBq1t5CpNFugdqzGOLSy
dZTgJ7So580rXKVYgN+0WD5LC+dMjfd2WlnRWcoGy9VOsV37/38S8VCMGhroylp/B+EWyVpSPaUA
/8/fu3iKIbozP9FzesoH5LWDQuHWU5x6cY9APymMLlpqpWMsgb4zgWzc5kxzGcvRQf50Nlqrr6Ol
1bANAFBFBBn/xAPopb/tJcFEbHmKZ1ylBHziWfEnjDBLIhA1lWYN/C9wI8oYDZ6yo4XppJCyP96H
r39V6JPGgwMUnx7AIF+qaN2QQ59qd9HhBvewT2lKkqLblJcCDUA7VuKTzEVb6gFNBXEhCaqBBYED
kgjpqbVZc5ld/OXWfMfut0twOMCBe4f2J3oqwGtgRd7je9oT7dSSQW7LJwSdkussj2KZNSWk+UGJ
poFkaM7vPvpITPseh+2CCXBbX7brO7aifHDD3TMAJ3ZlGN8vJ/+8tIW4FVBHfNJ6g2BS8NXW/kH/
aXPP1tG8onMDnN79HG65a4PoV7Cr4B1EwS1YH3r8nbVXYp8wo3kr2uueaEnbdavz4kZix//9SWi8
5D1stJXKlK7ZElesxjpuies9pgBSfcHCYYxATNQv7NtiFwPnlpeWNY1Bl3gfaQu9BT0jf0BkzEDP
iA74ginMEqaxtZ36OlKXBDxHveZgZpl4Vp4CScIabAghbeglHMwzAP/CMC8UziOx6OiK4HoICoJM
WEl8F0T52KidjTr8qudEQxihGiohXP2DNYFUBzVR8zYMgoP8D+LFNZoHQR18k3Q4bD5xsMcDh1sY
0NkDFiFiqiSPycToFKRz/mPbhRrYle6l/oYbGf4etP+kaiYMRkXflQNIu6hBMhZtBV9ijG/qWcE9
i5FXnDCsLxDFaicWX0jVG9rU9dTWE3PQb26WpgGhGZgo5d71VcUL5ne0MELkXC0ZoI/5mXAo9I5d
XTpBnS4wIwI9KjLDA6kYIXbcAlIp/BJW4QcP/arZWrnpaRjwpaELesPz/env1TnH1S4Ip7Bm946I
Vk4pTjc0DmV+n0txgDkpH2IGBaRnsRfaoocpSKTZGzS88fWvMC/o6Tzsw32AtPjPZclPFIirRSaB
WzI0x9rzbTEh/mYUvj+1cuJT6K75Db8gLFxjcnI2knzgQWAlu49+XztTBacOPec3fAq78DPjPLi6
dhFoU/F6MGKMNMYD8wzbZmiKoqXEu0fMkvgWB2Men0Tfd2UINuEhRlNtWDJWzLlTgTdokd30yFN1
bnGXdgF72XkIejgK4cX2Q9d+YMzBA2r4VZSrMl1olMZDyO40O4LYIatFtJs9ckv7V0j4+BzalTza
PK951jrAANQFb3mPSTYPCq08wbyPFAVHem9BH8CY1JOEEN6FOwC/vKLjTIOIiGNSxMV5IGXQNkGk
NddxHx3yPPP1LGzYww/QjMWi/p+j/mRFuxJe+FgrRn9gJqrBUSHtOL/8WXYNiVbFRw3CGsT/m4cY
jvxg7iVM3N7ZfFGx2Kc1mNuh5MVIjTKzsK+xxjsmVRFjoJ+5Gxopb6abIwiYMDTB1j+Z5TE0X1Pw
Cd39+1dHVNWu1eB+5pcJSIkLe4MEv2U2CBlF/5cjLPv3YZSX+7fClODbyndCq9Obego4iF0Ualum
e/XH6dXwexxdhtq6FE91ys42XeI29xe4wcbVU+IYl44NZRl6gV9wIHJrMSH4xOPsO8wb5Q0eARL8
ethhwW25R2c/qCgYefA+vtpthcuwnayCtld7pJiLXaOvlpampw06B18qvApTNM0FS4goojy1d71r
MREmuMln8DRmzpkx7u1U7sm+khf2AfjzyeRwVztD6dwwwI7w96CfGQ9LX2YEZFkfivxyy0cmoxvH
xs1F+BVDoNHo+4EjUjNCw/GnUN9CsclhO7qnFH//rBq3uUC0XmE1LkcLfJk7e+j59kLMaGcyU0kF
wn4oeGnW1hsXm02g1trokWlGgXDZgEXp2kFTXbaz/v3EULfUY8zY+NyuvIpd2WIpCmh+kcGOgVnj
1HXZMGhJpHruLQVij0cS6BZ6W11mKC4GlvXshOhCUiwaU/Tavk2LoSfPfXzeoMwp0XpePx7u10iv
mwb9/lbDfzpeWu3pypClpLpuYB/Dd1xLuq2mcsf1KKgaiiCv4llD8VJASDY2oJpPOnRzxCXjtf/w
/0jXfkNFXI9M50XuXSLAlz+ofPMq+UsqeQSsikh0hX3LAFb3sqG9LD+IMLnM0/VNFd12B+D4La6g
zjqNfYkYFTndjMl4nwlGDYbcbrhjOFASupBFe9dZ6Z6zBXxnw6TkFzxbjzY3QjFKlGlYEzKXPd0t
rJ8wUCrKobS7QhmRV6+870TlVnbwfFQSjCjHxnfo5Qi8qyeoSUcw8wh9eNpf5FjS7l3LDciXII8y
/7ULlchmRphoBLdcaouSDmpch02nz28ordXvrHiXrNs00LGjOb38G5Wbw6wl+/MqPG2zjfzomw9M
/tldOVLYIXtC2+iKIV/Nc2rdxP2f3R3AVjtM+ylc2hDu34FGc6YALKHbCsmnzF2flY0sxi+hJnZp
DfBi0i3s4g1yLOOoUCc7x14IkiTug8nEgnUKpNbB7seFlZKsBpRyGwADQLe6m+LdGp7FaqSApQ3x
GmX932bsiL37HolIYMWc1HYu4GuBtwVTsMyLnX/3GeGZdFSTA332J1LjWSe+6NFZCnX3JI/cVBkl
0UDpAiurE0tkJ4vfTJ6VhWYF/8RE1Pz8BjejrRmZg5foej5XRCBMDQjVnBtNEk+WHTMOeP5CRGnr
MtHJpKyJlJK55bbhe850t9wEdR3Wbi5bt32I8vqsAPbZ7+6QTbTT7s4yM419nCh3YfmwrkEChULp
Ce3AVuQg51Rb+Zj1lYd4konrT1qMYLLwSBjwxqWDj60Lhh28wBJ7iQaznmRQjLT3IGCfK3sWfJz9
9xdypYCnxy3ZCds0xX8C/+vNm780G6KRCTiVr8vw+L8PDHWf7IJ9u96Q9+PrDa4gfRYBaoGhufS2
8upQ7fCl4uHw3tTjiyum42Zxxig8cvoeRnLGA814yvo3XWBAe7CVLmVVkGi7rBthQt9Cup9oI0mu
xt0CR9ettusr6vlUDxoCmTKXRcrPDYWa5EHDCoyWNjWRHLzGO6vqAk/U3k1vEQWoBqFqEBigPTsW
LoAbo4PIck5E3dv3Cy0ywodkO+gRsd3nfxjjr6pLzSZ9JwPFbykNn42S2U9UOHuYr/UTTraGAUfH
uTwgl5De6VKoKsSiOvBmlDF1HOrZPdgYfu6KrL2XTcr2VHTLwA3sF5fejFMWcpQsIokmpmDpyoH1
W7C2mL4nFG/TWEllW/MIv8NofNhA4sQgty/mqMOPYtNwZm4LRB7S5bFT3aN41IjSVdKyZ2dCd9w5
XrzlRzJ9wwXl5IEC+VgWgRaEzDvJfWYr8E35o7uqZlWmKXKbxkQnFSILUqsUXa4oc34duEAUPx4B
V5becB7nQw7kO/UfDMc1qi84OHxHSKL77U11ZLFa3JoS6cCBlfca83jwoCrptCS+tUAepwWqJdCj
K0gPwPhMNaQlBBfLH77JzIluusCJb4Rkd28gw4z3anUQKzCC/USVRlRTHMMC8nJ1zdMkUpJmNFUS
vbaAYNIB73voOBucXNPJ+064mSzkvNet4xHm8+Q1X3FUWvqNGv0AqsWutcPqnI/0dyBUV6iu4KnR
l8nmGpO+L+EGfuLwVmlNqRdOYBR7gndpSKpu7vPHp1BbpV1fj5eVyg5qm4pXMWQMdLfv6BcNbuGa
dNGWLeIesDQCFkTBrg36VNu1pRSg2g/efaJuEedZOEEK0sjtQRR8Ed1hd4Xxdiide2vCgutZyuy2
RteoPOixlL9dspG9eBQWZhere2OrUYoQPuU1gRZUban/zi3NUHmfO2tNI0efsM+3brc8vhrfqgXm
yMIrkziMPtIlrqEel5JA6o8L9cEaHtO8blXC7lusbZmUwAurotVuh2Lwr9cQbH5SZo7RwburGFXr
6YLQqiVIClkYNxke6zjojOBaBU1AeSCM9UgN8F2XpZajQAlhKecfSPXTrFBhege1NbkqzzDaJ/WY
DoQYBWz8imdVoyKVskswf35sLo4l5NhBPbnHhY+v7lDHaKuewBjyZlpdNwdg65xgTnZKbxlRwT/i
4cnWQnhj5RdBDUXCWevNKH/uUucj+K1SsWhQKmmligqwlGGqXU4PybusTe5JpteAHXEKhq297aRy
n0YGjOsbWOt9zRp37Jt5gDm/sX4bfvAFwfxeZrJSCUoibUBcM9Z+CGO/08QBCNOFY9MnvhE+Ab46
PmILbCwtiXUW/sgCFYk1rZDvBnIgXzHtTz/EWdIqTBttwPmfM+NFfKFARE5hZH062HLORua+XrrM
6DCix1w5sG7iCT6NPGwDWeo/+Ve87rkOfs5FxyQmQ7VqBb82O0IDEdS+lPOFu+wrmLttRwTB9iPP
DEyH61aAfWjBCKtDvG2o0Tqk7S1eG7bhMy8NA1njcasag26rhzkNmh+sFyAbQfW99DSj6TD+Cd06
x4tDEz64LUSXuHjWInVQzgpgMxMtqUhYAZjVp0AVTOWOaCcSFNkPtTlbxKQIVmzrKaBbV5ObeNXn
AGZbTq0MPBoQOzpGwp7GqQ4gQTCIGjdgdLjLAB+5GVcN6TAHKrM3eHMdfqYdGNBKAZjueBeUhkUR
PLGAT1370wEF8a1mzf+HfshRI7BDUM6NqmbbniZuuMHjFVruNnI+sFtCEvZ502GiJYwHhsWo0XfC
H/xfnZuRtRIdf3EwF+C4/npBZX+ygPnHvE69YpT6A24PZyRJ305zilKj4xnYq1qVIpgZ/8yPM39r
LmFL3aBoPDHQI5Imbo8DzOik6C75DJsr8iIqLYc01RLz+EKsQekbgfK17WVFmKL5B74hQBP9FafZ
cB4yxOvBZirSqEYZKckM2675weKzFMQ+29OpMoCudj/zpzzxD/NGJI7IIU77/9NGsbKB6vdFWmkb
OUEE3jUayLGEaCyAOwF/+zIX94a8mqtRK0GxFDiatFUYV+VcR5BEmesYGKkmvxBVf31mgdCbMRwy
4Vz/CJCQP7igM8VuEwPDOg1VsLxaUHBNh7jR3OI/k9s9+HAkSdW7aseNgWo9LJBht/PENvDX1qrg
+vMaEh+OITdpPqbveDH7OQvTb1u9IAFlqi98E9Wdn9OXe0VbznyEK0OKsYkYGAV+ahG8XqLwWZO7
dFqCV2pH3GfOgQb8v25h37lW1h8bwoIQL3uIKaBLBoVuFqIgQh1apPo6GPR1PNSEKVTAJzulssEu
VnvdeolNVBaddUnLMytMzzpmCjdl+Z8xGkOLchuOux2bJbM+huHCBtqmOya9P1j/l7cABpJBEjE3
jWN1xHdjjXeTI8LZi875gEiscGPu7bwLuwUh8uk0CmPpIP8Po6vTIZmmY8Q6qfxZ2DyBMQz9d83s
RF5r75b2nXKS3BseWwPS5zOkBn+cw6FktEiAK+r8JsE1MsSxi6FCN3NXhtCHc2sJgF5/O1Vr6Ofw
BFgajg3flsexEaRTl66Ar5NFroLZCUH7GP/EfNs7y+BjZgfynGMmugWd51xm2TnrqKNTVhZhbnV/
bmqQAqmb4cBdFZxtb9Cxe7eo09ixxgks8wkereAMlQRwBawRmGgbsQh5Et+e7zO2o4h+GN0UuTto
HE7NPrUvTLxaF895PPXJzJ9QSxTSf60wIW7mypdLHTriBOkjE3TQ8DDd15tQyY03AjAujIe4v5Rv
dMVzc7OOWxCngwJgrUBigVFfstrvnnjtISBFWjVEl/ct7R70qUyRasaXvB+JuD15X3KxfPAIERs+
yIPn/NcXojv0+tGmZjV1spnTqGZ9Y2Zg+mUX6kj2OmqYHz9x4NtPFyZD9fFIo5Y6vUZOo5i/IFSA
e78RhUvLKTZrSglTVhVoorLJlJlCTB+jaA9+09AC922zPL3nJ7g5SeAiidff7RkcPA5yFUSPEuDC
3zDWqkUH0W+n6+6GcBpr36toS+cNQH+s92SfkBgsIU9W0HtN16VgKV5+aFCprrFmc0U2LFtkjqfJ
DyTFt9rV3emBpm/K9CDU5EsEUSd6v4H8TLcRT/ktytE5cmpjVBE9NMupNY8h+zh+MTt4prfM69Ji
7Y3gCX1v/jyjo1flLaxWmGhJSHcMLSgP3JHSY+lhPIlsFyzJPO44x2VOhPi2PInmxLJTme2vKIIH
6F/lJ9LZ8gNM5Kc/08D3XUw9gk/SHQgjNRQZ3dKZEVWMXaQi2uz3BzCd61WAEVuSV6KV9UXu1gRk
yQP8+6KpKhGwPwF2tIITDjDRIsKa0b/BtvJbfSwqurZ5wji+t+Yh9W9IsLtxtc2QJ3/dYvjDO3j8
5LTcQFQnyZQWKnTiVv2lfgzJ4Hg1j2DEEBAQOXlC7zlqmCbsQaetvErIkV6TdSGwJU2XGpB7i5GG
Rw8ci2B4FEAas8Yn/0dAiAcn7J3wYhGEuTO3LJ7AbiMnQxZbc5068NoaQV05NnYuKZaOZSndsZa8
rg8fsC4LX5VHglvBfJAoro9QavfC6wyilBV1ygCOXXy+cgbp+INRV/BwBilyk9HcIXUMdgJTfYyj
J4+evpaAN73oCX92gYKxOI2IG90ncvl0FZVyIUsMnh6w4X3Qu0FsVr1IlhoYzRYEXmkXNA80kH7f
RPS3M7eVrJe3h2t64qclWvb3vpuBtn5S53PVTWgwQEVhRmG6Ht8GPQOSVxy/3nex1IQA8Fzj9hEO
8WY6inWWulbeVnCFw+i4J7Zuh3nlAZ7UZdlaFg1NXrUj7sPmboqygW/D5HpkWd8IJDmC8bQAefGz
7fRFejrqDr4q3CX8x2zcp7et5st3bpMeuhazcy1jlOFg9d0S65c5NBDNFbkhNZ1Kwb8PVymrj4+5
01qQRGwxvxnZlqcB7DrnPPAyQ3Yb1IE/TpiLAWr5IPnzlHIkV9wAIpg2nHae7af9slbqO7RZG+uu
Ln6X3EQxj01lAqbhj8IZ/opd3BPj4Ef8Kd+gYX9voe+n5q0DWJzzkgaqyWbR2dkTm6DGN+BHV+dJ
11kikl6oGYUhVKdZfotP4s1Ooi4m81+W5y5MyWIfiUwgecFzCk+Rb+/s3uWeOG69oXLEPWh4j2G0
98SUCg2dvbnQ8uuKUcs1wGOpIpB/bkylDIYIPbCP/+NQa6v7haCo2woAoSMfqHJdcNfb8JLsXxyc
a07XB+ffMInTex04HKspsTYYOF+s/lIW613R8vHdPTz+esKemmTfKFNBHwZpomtDFM6AYFVtqgPb
tAoEqcupxzgfiLt/GX1qmWfjF4/4j+ypNm3y+UjHLDkOdy9EDJP53amygzvy9m7bP2269QCbhf+/
lAPvQFq9NZ8aNtgSqXIA1vFfTGcLkjpWsMhZkMu4VDpFgY9UbBn8H8q5v98/hqc2Se4ynwVnXdCa
III/MjebHnNWrbnTTH+R/Og8xOi8PQS0yaqnDwHncgGZqzUKKqDLeMcZG3wKsX+R+HziC8/c/7EO
A2iO/4wuFQOECBI75nJWP5YB0WSuwNhbjLKSa0OGWL8dttr+H4UHphYBMQttIeAGWwlV89Ll0oQF
YhXlo8OwOq6XsWeakEdrv2YZQ2RZe7rvw2KDMzWi2Lx/kSyPQ2U0MpY40doxQ6qtp5ZODQRtKdqB
J7yt1qU0PND1xEOdWzC/oMCuJHZBpNHfJWyZnIz3FzPEKfkQNSxp///elST+jp0tSSWqraAST6ll
J0/wWKdivVlHJf84QP18e3zFBa3bPBT1zO5JLOLrLmh8gxsi7HLx0UNWzRjkDcylRh5r2cd+BP3W
tXvlgnCntQ8YqI4+doJ1e+dz9V19iCgb3iTGnratPYAxm+kV+drLoP+ZsIKBc2HpLcqKPl1TcUE+
udlTRtqLBbW96xx7gNJg9rffqrmAGTL0amzlErQdQIfeenU/EnPyjMemUhCkjnbxqOZTRM67Yvkn
54z0U2blM1NLgzHvl4VGMV84LjgYQqSVhvh1aolQhRt7nChuXAtbba/JgDDKEFE9l6kfi4IQVev9
EIG6Z/1zYX6SnRj+yKRKjP5gfYL/LSYf3EnY+gt6uL5TEEwVP29lMhtLfdso809Dk+MZKd2ixFWe
crXg17WiWSZIjXU/o7j6YsOO+C4CNwcPaFsJV7djNDqt4zYbJFUJWTn5GVIqri6jdaFmaNZGjsFH
RQczHEgz+5eLK2FBKDQq4hgljzlhIW5ZI9HQz/lsu3I6xzJAigpzoPUMA/dujqGH0n0e8CqI9npR
Hny8HWwplo6u+E0urP/RbHIBYHA8BZOEHFrE79Jvpljn6kUO4X6hBNE51MKRioc1w3jqe/vWA5EL
EUrpWUnHg2voq0esuDlt37/RwgJhHzjyx1r/i6gsqJQa1girTBSym5iQGspd8ujTYULclwg+HDIU
GqITyldxEwAVs1PwmKw3qEVBSvMLT0y9AnDmLmU18heF3B6jXMhmfLnN/aAx99KLGhcXxvTuQcZO
dApdT9UBjikriM6EdV7ojlzUEU2IW/ESdRsuQXt7ZQYWFcrGISWKCeo2eSWck8CihRK797bWhsLU
pOlR2Gu0mNgylui9Y/9oOy9I7zmF2mEJ6wf7ynDDyTNRi0XJjSLsEo+VADhFhz2q4F2Wkv10kq5J
QQb90JmBdhp5dicZIQA2RYqv5QG8xft5Jb4eWMs7z1VZGgJHcsBH/vHV3dYOCGFOyufUJhSoyQjH
6Ltoq3mdJk0MIe4s+bytKWlN3j+vok+4e1/PiSsCEaCkGVoHGchBSV9Gpd2HcbSzJssO072Whl5z
OlEPHu43RUz7vwxz/nSm7X06lFb8edJJb1WqwQKTrlrmM29pMDf7g36la0dk1aDbUPl2gAbw/Qx9
FZ0iyw6NR3YLhT4pw7iS41YVXr42LI7benrr80gM8jKRezOAt2vfBzmie6S4TVPWDybmpJM4QJA6
2Y9ZjaX3x8DyoIEsTJqhhCXDb3Fp4OgOLi9LpfHZRCRR0e4Gaik+f04568dy6+yCSqiwx+9Fq/Jt
uha9Ugh2XRtppitrDxiDh2WHeCAG5Zo56lZY3ayZihUkUC/fe+ED3Fn3ogRn1m7z23i5mbzWF+id
YBHB4am7cDNh5qlu7oULGX5IKzrJ5xUEALx6djAin/BGD9DZTdN9vmC6eAB/Zn00xPUoq++oKpm8
MhEuYwT6JmuTSi8usg5JqgUDkvvmu/mrzEX2iYUn59zUz3sjik3YRyVJrzCMa7qE7g+ApCIsnsL8
ZhRenzQMqQ0FfIteamjTZBqLzq7npxHyFN7buc+g1oswrmBAQ+2e3Hujop5RbcjFUQx2e1S1WLD5
AiWlEAkAFVMeswiAZCjERwv5XU5WWukiZhunhTvV2TX65rf8sAs3QFV4EqYWc0K1GoHbfRDIcPaV
TLjeoSmwtK9PBkkm0y9Fl89saLGZT4U78Wx/cOB2vcP67Uakqon4wMySyvsZwxxwDYij0LFo31yu
qU64hfLxUbWCsHvI+WAwzpaCwkiXNObO4evOqvXAYU9AV1kA+97dXXzKx2goGs9Xc/mxT+gIZMfw
4Ic3IKg5e/t/XnriEM/xR8h+0nBxzG24xzRnqW8jllBjIVtsuVFZ5LKf94IRq96QgSwhx6JNjsxF
SdZ3fDO1pf5rh40BvKSaFqxQZAu997CZP6el1uHINQU+eix12dkZ+qFKh0gYPPH42Q3Z7uakLHfk
tsmN+wxjEciCadXn19C1y2ZS7dpsIRAv9M8fu560mAB+OERnoJLtR3mJ4CkTgEPHP4G87kiLWFk7
fBfKIcb6a2QJiFP4+u4NBTUB/0DnNzF5u0DS2PaRLfEI1WPI3eD/s+TYjL/FjUbI+chl9JRwXp8N
M65K0X50PM6nWekpOYw2CM8unl71zV23d5Gy8sUvWf9mjpaqw2Lr+KSS8wWsqsMid96kbWvN3qvQ
fVXSTXE4Z+heaiZ83LtBm5Ziyu4kZ3KNDiM6VLRmB3wque4uYCRgpj8rhFq2t1bgBsD6f5rjCoc0
8LtZ8wYEuFEH9t0pBNHCGWxaG4Hmg67GvLl3OkDcuMVVqiI5+LwUZ+5+nwmhW5Aaw5PDIQZ7KIHy
fPMu7HAAx+poaPAk5H1MSGLh4MyUvM59qQ44P9AedKAjOesBJpum8OVbRXV3FJQWXA8+GXy+g6zH
lzWPbuERjAsQodMkhUceApUjkU/CmffVLfKfiRQ3HlbiV+NFuF5EeDqC3jlTQUH4GVK+uE5J2lRK
pPb+cOlCNXGS9lwVhQnSD2aHBVk8l7+aU7nTnf6Iagcp8Xk3pWyNuKLTP15MixAP/80QAWpxK//t
6n/BDBzL6g2irrb9FTrLN4tdj54juJDRlZ7uXcXXbaY8bKBKkxKo4Ajdur+JzPvO0/hOjnwtiIdw
qK0XIDy10iv1BjfNNq5Eot7BUrb/yimm9biyuXnk0SgVMtmzyW3GRYZyevGapWBmtf4fIPGl4uiP
pZ4LcJ0Kkz3b3HukQAnMZ3PS6zAFiEqpV/3o48M3vzwYPMa+vlzTNeXsLYqVBYZAvqXtQzDOUbqM
z1cNKWEKKj0W+oNhJrl1sP7b1FNUjy2CRukp+s7qR3EzdsmlVbsS016CpVaDove3lJN6shaRTZHi
e6DrRipWeXe1Cja+syp0pqzQf4dGroZCXqsYTf17IRFBOlIG9f6rZjrl8ItBwzMsBXysyHGIxs3Q
yG5BM8YPQtKLh/KhULwnmppjlXb7J4CjwuYvucRIh/eN3hlzzgZmKucAxhTTHGv5HoctTWgn/j05
hsS+sbSG2UbjAbG4lI9pMrvXALFHDGhqFWlXLwQedJhhweB/HQvi4gEu6jv+S0pcTJ1/1qEOg1ti
1s1+psFuGfQYQeeJ894U17JgVM1y9+2R3srdbauUvnF5/b/Pv5jeL3k583Qq8fQpaNeF+dRhiCMt
3pu7Sjx0r270VeuKMfY8n3ev/WB4XGgAbutUrrEBmTl4ZVUGNNjRJ7wvBybe6AbSA5sRg/YS/BYU
9uBvIzdzWcq1GJ1J6Ym8lpryxgYBb1ywYkmEX0q2wm41cDhMSRqJkh1dvBbBe0r1uSwFuuL2kQjY
hHUoBe1ZyXM98WNRXnDQ2NfLrkzx3ddE+6/ShHjh4nKq7VG7luAku6DGu1ozLQ8Uk3HKv8Ts5s+z
ITCPf4gk3LVCbXjxQ/nJRDyO+4YamKfTE/TnlY0OSNKgiSqZ9mUfTGJmIWFWcp2A5ZjCaaYR0qkq
YEADeF+2uVwPX8OeO/uRU4nf9aaLk2sHSdmqW/7GjytG1aNKZ1RhZIaVFS76pOq4e8kHMA0IlsMS
GULleYsiRA7MDrIdBXW9R9gLZOYF9fFOr498UfNhSyRMCWr4i10RemyGgqtxCUbObmzR8Vg26kRe
u2WeXdOd3NHLv4Hrxubqz8Q6T+Q9fG43+daCnFkLIaxiSBS0GFm5PbTEFCN+NoAKwidlj4tII6Dl
NiJ5N6WDIx7U/0bHpb6rZGgEAWi6g3sctSo6OaoBE0oX+1XWSJ4kxPdDamCAEarlxPEKGeQvkJ/f
N3wSR5GTeZcq8bEEaqKLF19Or0CYHh0hiwM85/bqEz/vtwTrq8X6ymgAkDEvHGfzx7ZIvB16Vz/U
TPiPnwXTrH7P5nAcri401R8NHYLmUTUtfokdnvBMmS9vKlYmS7Vpisn5xmRgL48m9m1Q1sTYolve
zcegU1CtVCGQqFsjPiCaQTkjx8jbKjvLBO38TMYxhX6W4HHolDN26Jiy17/GlNN6eRVE/tFfkGfr
aB+ms4W7vrK940jmVFSIg25BhUUSRz9O3snE/p70tDD8C2WwhTrxjarudbfBALUCVOfv0ddvcUf7
0tuSqgQ612ssemA/ez7cIWgwvHYRzo/em/jcvymPqocxFngbtWvF/wIyqWqBRVvTDTWA15Y/kl7j
zY62FeoMmo1kTX5ukvbHfXxS6XYQEBXLqRc/qbSn+I7y5XzJhLWCR7Mw+PtbWQJZ0sp0XmlfQI9U
DzeEc6wX58pHCl8Vp3pANn0guAG2qNkTiSBi4yFoEkqM+16dkQa6hGlbnS12LUh/THS9REP08BM+
7uSiON4z6iyq4huX0DqLycT1GrcqRwfgQ5iiknShKj1Dq/419KfThPWxK2ntfmgIlLlRU9eYvs22
QPKi0gPEfxwe2XbRmoosph1QEps3eR39TcjARUqy214S5zWtkglk0JEWYSA4U+wHjie/7SvTNn80
eYt3LrE6Xn98L4Hn3jUGCUpn0mXv3XfMokQ7ujiqEAh0UwaSS7wT7G8rGqqmvEyOkDykU2b52RBv
WqHZy1iQIr5DdRSZncaTFHoq8o+bEp2afTsKaXnuNVxItVmefDEGmWaTBr9BktUhDH04JsA/txQ7
RrYvbYgFv0j+wswLvnefy6Aa7+2oqoD1yTVjMCHRBRVPRLC/TCOlF2Kdi5TRzAsO6jXd+2qRdkAE
LtSXdgpam4njHHZst8vMdZ4bQA5SFynR5bffj76tSV+c7J2LSJx9UqnlKtd4wyPzclbAIdmQhcMD
g9iWTZvVylEfV1O6csxE6Rn+bfm37lgbBbaf+8npXGe6oRG+pdQZr5mTHtju4AO3hVz/Fz9NC8XC
Mp4AVTlj+Z/B6KQoiVG0Df4FtA4j25Bmg0lYNky1n6mbR3H5RFFfNynUpIPwY7SPfKFLl4izx2YK
w/frX55UjtDYywIpMkvu/QHQOhKIvb1FOlO2cqN1B77dW+0X1ibroRcnGMk4muwLWXrADwTToK4p
VY6oN4HjmqjBYCEhDuHtanKh3BlOlviHAvLbKHQczPdn9/ZhAE3BjjlgCcM8l5uedm/vDMw/j7we
m5KYD/Tui1/1TdXnf1UsIu8Eshzd/giK3rYVEy4hn5EtsB6LdvIBeEF1QbQnGU9Kcran/aZk47pM
0JkBT2ne6esNLwDYFg2lms4VQYVPnVUNBntJg9zy9AjxwzGkj9cL1LztDqVJVDIOoEjdXA0a4XEl
VMFpjbIZsgUnph9r/Sqh6o7LW7UIuuk15Nv3jIVHaqausXNmHYDJknSvpKBvVfk/z7VYt1Mbg9aD
S3JdLrrY9ButlVDSudwzA6HTMEFEMssm3o+VwiCmAAIrsKjitbgRufJX5HgoNFFr0U2h3GVeDtkl
aePk5A6eI5w0yYOVHiXA/Y9wefvqVQ5b/RDLJCCegWNJ3mC16c23Fg8RaL0iwEvsv3C0uaQOKoff
GyGME4qrtAkzmtyJyYf3A6j0hTgGpPa4G8J5CIE557ouDLOpcgzgRSGKaTltdkoB+jNM2zjSfadn
QyDARMOn60cGXflbUqEHXoEh8JhLhSf9pwo8PZsWKjcSJidRoIp2eTVF3fEtal9T3IOvFaymbyjp
yRMeaolqopJYpih1y4I2ZPS7/mdoFGFN4HMKcqmF1gzijMYPfFbNJlt9/+pUnIbocGt/T9f0X08G
oL7PW+orz0anLQhRXzTG/obqNHs6eHvHdamkgtZJYUELOHbOp+/I3neUn5MaVks5nzocIvypc5DK
A0jBGas4FPKBEqbPj9e24Vj48p8TK7LK77WUMzuRvNbNuqQnOOKBMHJ/pOrx5/WDJWZ+eLzQ643B
A+U9+FnkjlwdRooDJn0+u9L+1xd/kPW7Ji5FnsXaX1PuXa0QPvqRBSaoknto42FmFGo+rsT6+y+C
njC6MCORY9yhbPjVHZXuysKvQC4F/IN2FvkCeK2d6bGDjI60BY6SRetkG008ogxr0W77va6QTMai
iuexqVorqtBizHvixJx236nraB247uiQH7pjpXZQlHpFM+hX4j72Ix2DLLtzqmamkRumeiFNS8qH
sRqq9GkVzrStMPbrmW5dlScQyoSRe/esNB0JrsyduJ6wMYyjW/+G6FvhE1e0s4dZMJ2ScwkWuEoS
G5B79VTQkRf0cVm5T1SHoWJZDXfK0dUxJSH66A5AJ9XecqWmBFyjkLo1NxL5EtuERsUjM54BE1B2
6TQTB5aIdJg5H4JlD0b5sjp1WqblsFQFOJsViId46DKdtscouHFqNWqiocBKZLtVg+deQHYezHdu
sqLv0ni2eJrozW2phNJQne8JvQyXMj85B/iqa2tbYVEx4IkP13BgLvm7YzLWhWFVZjXDrk/lMJbQ
KB8upgBZVcpu8vFEj1MulMgUZuArdkiMyc30Rtx+2c5gR4C17T4gsuZeAicNo2ynNow0Ac/FXOsE
PVC6GFtiMCdOsyhUR+C7VyTkZk2B7vwdM4zCDXDtahcXo+E6O9XN/TGOhrEya6DZcgoPKL1XGULz
WkRZmtMtbd8X0ldIVcF8EC50CchTs2ZiXKJi+izb5eeVOieQIe3ML5R7W4iQ/6Z+75VT/nl+ufjf
mTnjh1rapb69NT+hbUnP/tVYXK02EjwjNYHucj7LoG0jvH/pzcwCploS6dUsdkwmukG3Elw37Mrv
JK1ApxNzML1cfcb4S4IqF7TBzMI42Bz9Ek4s4gyqRJWhEx8sl3Bc+gHy8n6C52oiP9shec3wkuxR
h7HB3HcCX1LwTxBu1PEbcMkNMJnk8bCHxBqmQTl8ykC6RP/LC6YakZfU5Nn/OAz+Ta0fq4wqDZBG
XGDKssJOPruzTb7naffu2EzwQKyM+TxaJIX4ZQJ65BjgBtZf7NZLIbXl6xdqNHopt+1BBrivzBDh
NsgxQHv8NjXt/tUPn6EhBwa1pZvPzAVKA+4+oKegN1OUUhZq/ZXvaG2OEP8o364yxIQJrMfiOrGG
Jp0KHmtrz2dLazhszXhiD6nr9KRPtRKpQjjTP75fLefSyG+G5sArKbOYofyKRuLAHNnV4x9eJ/F0
uxlR9wOp6yzpZY1RXLQGeQ63iFAKtwIK2IrF35iMLcn0MjSlH7uutFimpkTdvi/Hb6mPwWDtnn6u
qTnrZDZ0jYNbb+i6A5yP6tuyqLMJdGxzcn6j2tCjq0J6Oy0wWrgD6+A6Ce0ZnMuenLvb+LTRg/Mx
LkyxpJtgSGtW/YR7Qvdz3uMotdv3FPeav+1iACJZ8/D+U2q9+/c3twmr5KJ8VWAyrUTTs0F0SbMt
KXGlx6IjQDJNnJ1XK2pMHuAv7V3R2P03T3P7mapBiPfF9axcXwPQfoV7A4rPh1ITi2nJROHCSbe5
2JIFHgL+tstUkYmf6/GDCiytskW8Oj0tmFwdSC12yrd5WGdF4rGZVAEooXWgPaqSfJ5U+DV0fJQ9
naOwkV9N6oTJF8vhQrb2WWSugx47McdQsAfskF1qhknfGPTdbwFdNrZ+UQ3rpfR9c/wTtxsNzSN9
CUK5a/XnCTwtzjU2i0TNxpvfhrDftNlBQrnTGFr4yCT7pthQdFZZJA+vY5SxeoIhDrf7AGomKlsr
2U7xw6ikJGRAuaekFX80eVOVYE4hOsAQP6kDQw/HVsguKSRvtfoD4up+LBZVvYB4jVu2FR1HdcA9
xVyQqlYZ+KsWTfq/cexqwLXoaOYa5YRBalp8qenR4zSnr/B+mtoXTz11Aod7JddipOMpGm2nOiNe
jNdxA+cRAYLmCf4H/FIstRPmEuPbwxqVx8sGeZGB3ZZblNdbjRjW1Xl+MwarYX11FoKftFsczhQL
x1uwmuIkZ3nyug9Znbs+Ez2wvxCngsxMLOE09JTB0Au4l/Pn2XMdXP87Lj+1zlU4tjNTHnaujmnV
cddqSF16gev7Tua8+c6bWc09sEZ151uQYnJ0VGsA6zg70sc5L+A/iG5hD4yeY/UjQOAgS8ERhwmV
xIGrtFhI2+FcTxgQYi0MLOtIJlda/s2DWWoxtkzPCM3TVeZq/cpAqcS20tETOD7ETQxkBfr4WCnu
w6AleHWicOQTYOwxldK/cAJwkPWgmNt5r8/m2T0W+BjJdLb1wFqz1xHr3FGDmWGOxe48uVVysWn2
ltc4CwyhQlPFub2XdqdHbKTfmuIwIUWMAbrsETnhiOXeHSwKIIHNwtCV53yBmXvbV+GD5xVm7uO7
wdQg7CQv66Em/nIWpRK0gJgg1IKNcV88VqS23+/6OvwuQefuhvXiWU97+VTdrYVjA68GLiLrdGoP
pThYGMfHX2sndG8C+AXrT9HKyK886fyKZpcLNLHDe/k2IkgC6jwNZ1MpQhGASOhd34WGX5nCki9M
nnZB+DW9WUUSSAGemRREG/Cv4ynowTALW7KcniTNFghKRZ+bhwZga/mT7PsL9D7DQDxwdmjWeK1D
Fi+3FEVUs4rC+Uj4d387qvC3P2nRgNpZBZnqI4RHjLDfeJBaGn7cRaHSF0IqCrFeqbRi+XIg99lb
tGloGnWC2j69PjQPk0AlpXMF3NLqBvJwLOaCsTYVc+HUcO6sdsXRrsd076Cdd5XHRSoYorQN5eey
h/8xfXFoK1fuaWHhG3Dn2oNpk8FtzDLp9A2jCefyclNj1XUKomw6qI5t25ltaWN7rlyoCnjQmaFp
0E9ttzlmQd3HUfmVN2fTMuQBOC3E6BVpW1LNfn9mV++k2YEdVp9T+LvG4hJdWhr8hWcTqdwAU5Db
vAqHfKmoM2c3L4+6DJDEsjb0yKzZRo54ITESMcBIVw6usS9o5jNlFffoO67ETrCCXxR6d6RbzWui
kgqtteJy5/jOs+Ze3UWigPLgIE8PfczyQg93p7TRPJ0pZHShjdumxYn8eT4mjeoU0RNiw3wM3ptL
pkbVFtZVu3MEkT/Sd9IYsOm0FgfGDVG1CVCAxnsRlAK78yQCEbYbyF0ZLmgo5t/JMCjivqNZYiFh
ijdC8UuKLMKqc1mUrhiPSgN+MuLsEP3UnZ1GJmQM9hEOw+4vmh+pBfp4K++RVmknYBmhrxzwNlFU
zXO3z1V5GwRAu34bwtNh5e4DG7w6R/a+Ht+VoG+7vzg3XBUb/Ux0kd9wg7ygI3axmbPAPY0LVtez
QzlApf6lb4HVX23qhtfMhkj2kJHNB/HftsAuhx6e4Ldqc7/n+8oW70xj0NuYoZ9qVoaBDk7iv0bR
0gM4FgknqJ72nrNVjlEb3Dm+NXPin4WuJbXGJb60zyor5EAoaYDGkMF3svk5TnkK3Mmp2brt+D5O
etCala/U++6zsNSJ/ftBg2SiohY4VAI1uPp6oaOPMUPj9Ce+KUtmqentmveDuTmh8btr2/B7pyJr
8ORdt5E2pj5xSDlfaX07z/v5yj91iHfk9rp2XOwDVE5lg+LjAwhWQ8uAmyPzl0rAhvSuO5XCjGx+
v5TpDghJLpjdqpv5TOQ351U3K0u4dYFDV6yaY1hZMwLV0IPU2DyaEByf2/MGKWtPX0gaDc8oi61o
QgPubXk3F4EpoNUGKunpqGrTtflUO7Kp1R8p/Y3Qz/hKjLj3Wmm/AjvWx2w0QeioYEiLB3+34H2P
jqP5HSP8PZkjZuEEjcZ7AHa7cdmOOg0cPRHu5p3nbFgNjzEsymqAoTIIQs1YuC2WpH7r728QW2AU
EfS1KJUVgGDHh0O531qSmre8Dv2Ywn8F7ZY5CzWOrWskBMKCT0ugX5iCGvaphMK5ujHiv1AlOznn
5VxR0Xgkl+v9ukVDmu/ZM56n9YTHGFmISgMuFUKHXTyYJC75mfuJKRL+kIg5RscjZb3lxTNP6BWt
WyAA07DeogZpfp/zUqKdsuW/w5ynQXbibuSPvGwUIOUGgLdpYifm8sH7bzjay69ajb28hlq+65TM
W4aT47v28o0RkMK+W7we1Yi2W3qmpWr1UEzGSBRg7vP62mg6Tu2hP/qEV0g/pGz9Ga7+nmL7FHZo
bjz9RKEdK21YbEVkUBTWdkcVenQjB9iIJpDSCcP5i8lpJ7ZylwJlj4AyJd82y+dfaUlAMG7ejGCr
B0sFVzAdjyQCHYCk6Gfff6Fmk9qBsaGqiDN1Pfd2sgFE9X+lMaerkUe7yvw8fEcwbI+ToeFKXf9G
J/91msaH54wLevH0vfsGsId8yp4rabrZG/GiKZGFY/iT1BEApKbhnSPrRHMWR+JHvUNQNnbaVi9R
YtU261nZsUnjE6mFqqJP4BFuVcqwVp0TKZZXuoHl1bPXhE6nv8jvSm276//vvwSNmEJEDmTRsmmb
kYFlNOc/Od07Ts+fqJoZzrqufI/zHYFsjNDdRmzuKzEGYHeTw2eCpRDi+y7a68MbJ6uhU7DCX37v
7mMC+KD8qOnd9ky9euEQTm2f1uAYqlx6zr5RtXnNcohPmIOMPMAXa7HfL/lrajcHwuQlF5t+hEUX
0Ye/BloHK8d6g94hh++BMyUxLSMGKWkNT4Tj0vDXA2cmIUKhCNSpy/YAAaaA+iprbsjyvYf2Q/QG
rgFLBVqayza03eQa1eeyYyPdNZUZ7LZ8ZHo19JjUghqrIPA6BLf/iK3biFwrMx/uewBqthyoCf+K
XwULvEXNceca9+mAmNVp7vTdCgC6ySUhiRQdxclhpkon77v4JMF3z3skOX/21gYphvgd5W/U9RwW
9ryCASBkE/cCFxi5Sc2Qa0MyMxIw57QyccehrUTeL78ECoj+fUjdaeYMp8bo9HDkmvwYxSUlLnjg
4fClYVgA9hktth5uxqeBhGXmOmmLQIrJibDcF41UEZ2jLYc2wgLObTjt6ty0SJ+ptxm3GW8trxqF
x9SDkWcyJ3b8zv8AF8FAKR1x0zoAFEaTzJfAlWa0bzaq1MRHPJEUMKRzZa8elG6lj/8yeS0zD4jK
7HQHOFQ+Jj17b+jNU6wMLgWyL6aopvhPu0Qa4100j7fF3ORVqyz4786Kg4np8HtuianaaHZkq0P5
7yU/3NK0gQA7LPwJWY1vGafkc6zg2qyTw0KiHwJuti9uw5dYaiXC/XHXigFqRYNhYhX7BsxkB69c
YQNtUDsQxii7M2/d1zoQWKg/RHMpbnrBwrx2g/JgkBabYqGs3QwGAqjfUsZGDMCcldfBe6Xye0Nq
DUj3UJnaLrl9zospUqA9pnbaFHCiIDT3SeEOEsyR39/PWoZA+8qWVJnv4yXwieTFM3jHt8796EFh
pcpkZo9nF7K5x8KR+QcOVN76VbsPDuLu+DDAt67qGOEFsAYR5osO/40/UFYeaLECenoPNnf5YxGi
KJKadEG4kX7jjvT485V1iDs2h/E4metDW3X9zCbfuHIvu1SpvIjzQBPnwuOSXN0KFnvclI9UQ22S
5QLrtoxG7O9HPgNndZ7huV/rDeB2RieiBoiLtl/Dq3PdjYPDBXBNXuQvsCTeV/GDHRs4i9uMFeZ+
J6KekIQK+RRCoM9Shx8rFLwAqTXRG9i3eMt3lAI6tAEDxSt2mRofhXIhSCD4WcUDNZ00j1+P9UPe
4SbGvKx5PTgfdNo50ircAr8QdgaS3Z0WHK4z9tOnCSPH8JsrN499VkLBWYQXijEqHxCqof7zlO2S
DPbVFNl2pdrAw00odJEJI22QMqerQ7483WIuiUoqd+XjKBmGzVgUAkCtqijJo3B4w9bE+sYVTSN/
cqbXoRXu/kVo6UYUAup/3ceAiLAnfUWUXaivs8QTfKkEZeoO1Wmax/4QH2i/c6ZHLwavBs0Zm9dm
A/Y293Sbkl3Q3TpJGzk2e9EUkUTQlPuR6Tw3CQ85GgLtAiTAK2hL2aTACdhZwsWV9/fuPJkC7PLh
SUUrkTpfjbdV83fGUcOZtQZATspYLqwV8hOMPm6JjIc1Fu5tgDM1z3VKWCGVjDLB7fdXoJ4ogM6I
1yNeIx4ZbBeKwv7qtoqRj/guqwgPY8UUSXtup4Cs9tUnmuMdj+cy5SxNLH/s7BK1MrFpAHMDBM4w
aG+R8EPW3F/F2ICVOwXgIw2kbYrn6UgkBwEE8f7JMLflaNoatS6YMXHOIBHGyjLnQC3CgFJMclxc
YQOrLfhy5wyCYbBPqBg0jhxzDLPz/VmwWz50jQQB/sBg+qYHm4ChtPoffjkHKg0YkPjwaj7QRkCm
fnUjWicWXPM2BWgVoMg3oro3O7Ducg4teeQ5Jw+LoITG1ZBO0dfmc2SgOT4EPSknNQ09a4+89pa/
Cp5YT4tFd3OmU5YReN9Y6LvbUOgl1Im3XPHXENmg522ztSBoEvDz44QjWPTiJe39+BPHQCYEu8b1
glajl7GhA5PcaS7SfAhHce2I1GFRXd38aPcauYuQfk7rybGq0ZfbyAPSOsKZybggFZ70OEvNoMAr
qdBy+RTy8jy9TYeX9LrfGER5O0fdFGn7/95aonJttLJRI6mtDD6cTlQgr9OYcNSpSUorHPCYejqU
UKk6dqdxWXLDxh45DB7eI5nhhmkCecfKMlg6ID4MgBxy6a2frf1QitEjNDBNwQBy5umFfrAUEx4f
OZHxXA6MBSV9B7HNdXMkyos5RYzh3if4pgz/YbDRYreT1WMMRRHVY7okjv7eDRTBFRbQN1pc5wtd
asHZDPKqIdVgoVp3md5y7AepWoBC4QaaFeFzIAnZFp73wGfZspZXPJh2tVfgsCGQIWrlojIQ+Zdg
znv2rDS+93xJKUm7WKYSd7NJ6dyTylEOAURuWOMT6tyhtsROL8pasmDQEqi4zgcDWGA35XS0iD5A
IjMZyiw9EXInJSZVknbCa0z0zaa+ENiM/OCBaB7dw9iAsNg+ENDR/SWeaGHWka4VO6hwRADxLeuH
Xr0kAkXT6vlLx5YYklDBTH6InIwblU4mU+wZqf2wi3AKTiASa/rfwQXGAoAWEjbnjIPtSDZ5aT+t
LP7m6hGNWWIbzNXQ59QuTOr1mid+QocjcuQKyudtntFHUNU3gjcO8a8ohY6wrqKaqvtlgG9lNeax
AWAZAvQkjM57FS/2KiDxWmezq0oMHWqHFWoioRth5CdYeslFnWZdqmdhnmVJYJVftdy1H7es7BNm
KgYPrJmZAy3T7EorzvSFUJ4LtXHjgO9vrQtqia6krbByBgiwJjjfpQxindNQFk8yyKhJArNHdFse
c0jH1eePIwbwSdlU6Z4riChL4yNWasWJiIMEMqaWv7Bpdgyd9XzNbG4Iuyv3r8dpdPW2dAVXAON0
K8oMJAVrjU6kUSKTa6cWVrL/yuw63MXscjyyVxDXCYmck/asyrLfD/oAZ6jjXtmx36uhvAAlOBu2
sGiJkby6RuLElFsyD5Q9ry2yvQOgANCT2lN9+vTl/aSUN8pzBhcz0hq8jaP1F0imWPHQghA9ccqI
2wnMLjqhKTLt/PkZfTei4bIZF+sXcnrNoKotgSzNjrXu5mKyzzrTH8cMTjc7bPFsNvcbnzw8peOA
DZGIiBWuCGwQVX0hPCuBdE5v0n3lQYe9JFGDXuh2oRZ8R924+lULc8lANY9rlRYS0qC6ykPDXjIK
UgDe6kSDM7ugX84pFPP3GWRInueZq75216IO92K7ySuZpOXFQxr72bXpVw7A9fH2PuK0FQpwpBdU
vGSSZUWXsXWtN9/hGlqlOyPKlohaUvbLCM9kog0+w62z9bDE77TGhhr+aXwlKmi/3H+Jk42MRxtb
ZkmEj3B9Ozs0kZKIOHeU9dnXn8j9PT6TfxiXQ8VFkQeSiGCXGc8Q8EU8Vtvc6cwAcG7/0ZrLZKiQ
1NjiIKrxPhPHB85c8+yHd0fBJz1kPgql37MaoK4bTJPEUHYoXsFdBjJcGnir+SatiIaDTXb3YPmM
kEQnQL7dEi3iWqMLFkqVF5V34huc5PKYj+9rLVld8JlozobSpkwrHZgGpsj83s5qQQ8BHejc49t2
xPo4esj89cIULldlHlFKYwFH9Rj09oopM2rB92Tmwh2rsPT5Utfx1w6W8Y4vPfODnJC1+r1/yTFe
n4KdQwbCkUezv1nHjRFUGlzM/w19m9Mqa7R3fHwnGcRrHAUCrYbrdKTgoCtRR5X9OOu4l1ssBLYh
7MjsOMegUpffRIBfUIsiRGYWubGx1K9DdcM60ZSai5UNW4i2rtHlOmCuzAIVaZ3Yx3YzXXaQLjjk
pFl0T6X6GmFNlRMUggT/wi3V2fmaG/zHSgn2DQnWghrRho0LFh3taGuWTbUWJMqymDjvohuAdIe3
nenqzgge2/s6RPHm/AWCDg5MXeXbHeRyKGNmWGih7mITDgZHsc1MWPiEadTbfrI/Cb8G669HYlPw
1vevVj0pQP3Zby0wD8QP/Lb9HZyn2rnsIR6vRrIIwfB4AvqU7TrVSRSIWrEgP+rawokYHr9Y52NY
eRabwfvVmxbRNJ1fJlZfKbZ/1jkFKiGZXpRkZhYVbAsZo9j6eFzo4aSfiJXjL4ewWKynPi+j/mGW
OIDOMH1fM9QP2ODdE8zX08DGxSe0CLiodzzQHRf95M7DkOdw5P5f0iwoZN7EvOwYR7cbrNq8PT0C
iqpBnLr49frWtx74ZWNaeaozIbYBLjevBvss6xncjRKeWPT/uVs+3tvyZyE9DHDE2y8YWOEPbZ6O
DTophqTafmConXgU56ZWH0OT5dvXNxACDn5itEuWGGxG0BXfLRFD0bXZp90dHKi6W7qq7iQUXMnV
G76HkpM6BcMXNyYbHClN0W6IZ8E+PMvPvQtao5ibQPE4Fqgqu1mL8/CJTFiwiHdE5cd943VeCJym
OxU4B2qIy7bBINdYZV7JXf4A2b+UHmCNBCPP8J4nxF4JuIlJZfVKPH1Sa6lwFgK8LjlNP+iEdGG2
DFKMEs7yl1DsaPZz++mh3FEghGGmASPVis24dqVHASk4xwjLNxTpn3A6fZOJJOI6ybM5aKJIJgFT
ucLh/dWBw3a9NZRk4870VVzJTGG32tfUs0K8qyOzjD637y0/2rCcOK9wCB5In3G8UX/7kgIqQKwN
DsVwdWsF1zG6gle9HrLwa3V2+zy3sZR0minIAT4HjQRkgBtwHmK4cW5CHPkdJRSXGjwav7ogJ97K
CqLhv12uyux1QZPIIPxyNddnDzviPTbHcO7frOz0uzCEWfiELBKiVt2JtXNtRfP7FUJrBasBsyhn
6two4Tp/a1laAt4AyzJa74iuxjhC8bXHyRc+ge8yso8mU9H9PoRE+5ROQKt414pzk0bSjsAwvAkH
eXpc8K/M/ud8shmqB06g4R8tDFGdZImFMTauUGzp5GPHFvkHbfrCcpFTZEchLapF2/wi7pHUxOfm
v14TSpPRaq5Yf+Ygoi1TchXvKLzO9ap/ixh6B29Vi8WCv80VzSDHo0rU2TXoK3MfvSAo1G1r3ax9
BKvqUXGVoxvHpMnh+ktmbCdIPRSjVDlqMwO4KkFVftiwcVb842vv2AiW6Q4gMPjouH3OsN8QAPxi
2z6hSIjffBasLKo2FUuY7+m9dTi0QUYdoe/2wOEEwEpjCtLC48Caz1aQnprFTPmREhLsbtFF8r8/
jnbxsq0dlPiut60ai3NGTsj0bzw588Y9sHl+wCB1whlt7s8pUigEEEY0MdCgBf3ZwLQYPq+UhAXS
MuO+Gd4dH5t3/XdyanApJIzYMn3AnHJ5h8xfS8wasafPCluj6NVlzIXmn98bCz64YSpjP6XaOYtQ
9h7RCCefFy8Fsgow1PqkK+bgYpt3NF+Qghgb8GeBVKhhOYiBh/J1JD6fuKmxleu7RMHiQQgahuoF
xra3fjWVRoHQblivWj7abwi8QGsvlpJDFgsom03b5Rg/WFf01HU7hhpjih7FYb9d6vHjgdLUfYv/
8IXeykOwqSyZDAyEL9H1bbpD6VNdKye85cVMmoUJSSifMLZmKr2ksy2dyRYUya7/5vqmIm1CHbao
wAG8VTO1/WVU693IIrQHddtEs9nK+EygU8+aM69tasR/GOhRq6iGLxypVF70D3Ni9IaYjTB8EF1p
7RS0RY6gF6LjB08S6nWYeXEQMgd9sgNWoVhU45MIw9Jd+wzf3MoTFc45ughfcDT9O7prJ7Jxef8+
BCeJz2i9uQ+pczM4uvJen/KgaRerhCwit+/03LJi9HruoCh1Fj8F2rVOhugw0+VxpgKbQlruUTTD
T0aw2ZD5E1jrtf20FqrLEWaEkJhtygXenpdjA7G+QNKaRPnAkkPmsZeGzkYEuMq6lxXmP+ZtfMPq
wogbpNa1dMCa3DNz3EZb85+woLsmfSiPn/Ll/YHpuifDRFFKUK/GcsvxRzE2RsSPTybm9xffLIBy
XQwYS1rX5J8OUGs4Q6WtEPjK3hP7fO94jtYdmkc2cJGagRpNV5OqohhaV8uSNf5GrOUMQwigjqKC
huXyKsJ71ni39tsYpajlWwgOBwLxeMdRbG/awqdulb20mOay5l5f4sVMJ66vSMnt8PM5dMiC7mFr
/OftQql8/zi7piODRe2rRRljHW4do1BBkmdEaF5YY4SfDiIjPnE3pb2yvRSxu+OvFb2VvfJxMLL9
pBwgxbbPWxB+j9ZKOt3/kISePSrh7MEs8XwYyuCpEA75I3LUKsg2VGJAsjTNSnwWjo8it8HqVuED
Wrt/5HYOsmpk8d8xqPBzyZbecmkDr3Shsnj5UQ7o97X3sPHznKkzyRUVv9k9mrp0J8mwx0V0Ltlu
mnBQkS7L0Z/Ev9xUXcttPIUptiTfUt6zvTud7o6dA0qwcumIEa5ApV0WO+vDe3OZOMg/8M35/hxh
sdmR6Va3BXn4vZGxYYT+7Mwhzr5g39bzTIion/45ddLbZmuRxMsAd79mujvWRy3HctMvRxmQAb9r
4vGjCQnZcMBk1vkyNgZxFk0NEwbcmyLZXXdL0IbERkRvcVW50Hr81wczLkJHkPCW/zXHR+0vd1oM
e7r81k8H1RZGlexgorkz8xj/DlfDqeGp1xdhmv0sMiDvN39pXTndJUBuvfnEi+zkM62F2Au/xCAO
DdyqTTX9dUMCa42wJJEyqXq2ysMVMnDJC09/2qRd+5yiM6itymcE0x7CsXEdGlD2BD8pppPpxsuB
peqbHzKJLFhRl3Scgv/D8UYE6pv8ZZhMKn7Fg9QjM7yHBfJDRdncVQQx6zo1vcvgFWSdcZ+7rhrB
m26mOZZa/o5zBrBAAUlQoXd1RFPh4JY6TTbyT7AsFZ/rfDXtE4GNFdWtSQmPgKxAXG2gkd7Hog1Z
EVuaGAvd5lcGf9Tage8Cs5amCHLwmfUwBKA0swwwjtJjWkuvKH6i7AeiH/jGsV0JHdFEQKsOKmUk
XZAt41nSMmpVtGGBMpercy7ticbGpV5OIhRB2CpEN1UI2AFFm2BL6o4+9Ai5ho9TtuIvJmUokTJb
DffX6DKGu5Bl5EHw5dqo6g/fp5SyZq53mDrJsB2Fm2SCSnU5XEoE1Om7pNksuo5AFslr+Z7mACUr
o7dnQTATA4Wo8V9c0Xd1WpchAJTBq1XkSvWth5c2zorFz4/SCmNp2444UNdnuHUZJbjb/fDFOmhr
ytHBYj86CZbUkFoziC/TpKKmk3ofklZ5uUFKou7fJ5X1PQpogvcwSt4Voir/Z62VYRLueAnQj8og
QeObQv36gaTP+9FeZzZ9hgJ1FZDLsjoFgWJnOz+Tdpd5s1omxtNhmJCCWrcx1t+Ni6BVvHVNa8js
xgVsPB5xdhHu4lBAY87tCiIw/ruzqZORDhoJ3nJ+MSJ/VLZFKyDkvZLzBoOY7JaQn3sg7rpxFig/
B9u8YzaD8NfnfB3OGxTExfXkgaZDCIIjcanYVws3wy2+gft4GYi2KYh/QZVW2aRdgOKwMNSsgYj6
RoYyMsN+7Jbnit2Sg4xIrXr+6TKVly+WlZaUxa86p7A1hWgxMPv53YB9anHdj8BvFfc3JPvw9lX4
uvf10OR9PjUgfIXLSQlCgQ0f6CnpXSaNjwUZVAhqKvhfHv4q4mEvMbsqjQRdUbV3RNcI1BMMavP7
w/ZWEQkGtDknDF8NBnyfi9Kwjtxd5vCgiaduux66taLnBNOZt0HrK16/DQmfOTG1ktS0dyc6kCN0
6semmTn9elKp+uWT7Y3McQS56OFr6RF/S2noKd7EJm09mBt6TvbMsc5eybH45gtscxtR79VkWKfm
tihdR+CtVEGP5XZ+0I+L019kOMj000rM05e+mCB5AGix8ky5QMfBq0itvYzWTVXd2ex4vY06q92T
yONnm5pjzFA9HOOHhkB39dCykbylEubXsqGQhoQYqm60cThYmkCA+bYCzbfb2Q3bSd6TiHcfCQcb
7se72Qs0iFjnm71PwggAxjMHCSzDSHUrtcW/zsQlXBkcpmMBlrkUvHHxEY9Vd56LOZPKp0mp8Owr
N+lMMLzOgl/7SXmghSmPSr8wKzAKUtv63Gwwskph6IOeZTxw5Ju2GXBFWhpJINLSUG0Ieqowm8u0
oaPkC6azy5DZMY7YHX1Gx/hD57XZtdo7uUYnuuVYXMiOsBAZFeUGUoi8Dx8d2VbOFqdk29J739Yx
lhPSLnRFo7K6QZF/dG8Tn4dg9js+ri8pkyREmG8LPNynW5/Ke+oOQkE77OjCJkgkFOUvET3MO5ov
9npuDOE3y+GuqYdWTlNVAhNPhd3W9Ecojxmso9XUN5o4Zs1aK+hTnOU/KaDzB49nC0LPS/za8W1R
3g70Erz/I+4m8HtaZvKEThr8mAOjnvRe++rgKN1U0zRqwoRiZ99kd5Kv/LYG5y03EPyUm+j+DZ/1
dekmUTQzxYiEb4H7PhVY7/5qS7bCEu/roq4/1dixPoSpTzafqJ26XKzQXWy8H8cNxpzNn29UtrZl
jucthWkSJwYBvSCtLZWjIupz1unWVfGaGZFC+UTfiYOoFmksV0/pp1V8dpujEmEj+hhnCQAHDx/m
YxLY0ZPKkx6FBeGq6YInN5qbPmRMTOOvNwytElY1hTTqrYWejUCp4Xt3wDaII8VcEvcioCiAWtr9
aN12GjbP2VCc8aC+H80Kh8Ctx9pHETlMQVZzWQ6ej/nAbyvEcF4LblHxhTydUo9L91MWuIfC97Yg
4jLvHGCGvmlsSV5jGD+vQ17a6mstUVMK7fO7ny/ofxqoQvzA0GBrqRDy1hRwp6ThG7g/1k5g1HOu
ynXmBNeGB0AQzgmXpiLP+3MqebwmB70X38agpaEHzSOKos9L0nSezoYh2uxgH7q9ZRiNEuN6w5MA
2hjgEMkEfw4TmbCTZbjszjPnbcxwzc0E7rmobmmy2LttS7pKgF5MbbncS62bdXrOS5bBSk9nkYrT
ZAWtXep4Gx0dTb+qvSoiG62vG7E7Ie9tJ+up8TyovyxRHnwK2NPJTEHW+txT7FoUU6k+X7em+mX/
UmXfroD0m5JM2dBN/tLkgJkwTzzyZcS/RiNRacFiwmR+4xtHgXXgFIdfy4KsBh/k5mR0fpn5u+mz
riSmjQnRpQ0q3Ke0DqOV2ZErvvoGcctLyv72wlt0MaplxJR2QKHh79j/88mYcvcKyYblZuGSJbKy
+/A8KOc89lVK5QddtBTHqVSxrn6koBFBpY55Ix04DUfi5Y9TducqSKMh8I5Od1yVLsk2yNSyFyZ3
9nzsTDiiEF1nuN1yKohN9Mxkf12Oxe+JfoE4+kNugPCu/wU+jRyxd6j/rZ8/dSLTptLvQAWsyjWQ
HPF2T12xhqMjr4DN14qyC2VsEAsSVDIS2Tus+/XA/It466fRpUvln0DPkegdrpDFiPuA16n2UIwD
brUMCjdONxeFqgZN413rOtvK/OXcS2PI8lbAVqV439rURT378hlQZHOgl/N+PsYgVKrMYSGNbDWp
TbAqwCkpn6CaRNlxjNNIbdmnFoIjJilT3I2AOuCDC3RdBuZI+nqMIgYj6R/gbIEX5wZXACNLsVTH
PfR05eGJk8mLOhTDWEyDwsq3uN/FCEgorCuJkhgR4OGDt82m/frQKF2JHujx/Zo9eoZOdjOFhW0W
oeJakjxQA8hmoA6g+8pvHHgq/8H0m1+UaaEr/jGirlG78eqh+RL6JTqEvXvOPxvI/hRQ+lacauMQ
y11PckX1ZqVm+DN1jPMwDRFe+tkxcqTBIwzUAJuxP/r17z6vFNH3rRQg6IAMmqqNJbsd7eeypGgd
IrfUmHJDCc0PI4YoZgxtT8gRBnj2FAG//ieBPRMus9kBkKjBk3K4pjDu7gBa5iB4qAGZzjTdr5G4
jbC6bNGsh3tTNs2EpF4VEORSkMuJEnO3QYhkDS+O8VABlEH2kXgAJ5N9+GqUPtrS/gk45c3GTSzh
T/VcDGHRja41/r9Dzy9rJpEkeAb0oI9LqSIWj1kXIyWO1CDQCF42AHJgGFGFgjBL0Kkmr/4piZop
egNrhC5A/Cl0S9soTda+yVTG0yvMkzNpr5iFU7aESvzcjceK80LL4rOhdWUADmpf8Unq4iad2MCS
FYnHFT9MmfDIVCEgYTdB9H0XnOBs3sKKSK1NGlDEViqjo8SYze9V0Hsv4aygqRu6+Qn18maPeQDs
yRksV4ZprYd7SkAOkwMZQ6jUX6lDlenFzYMZnd8DobS8Rqs/MOsUludxbgKj7NUHJWHbgb8MqqdR
Pk+79svHuKYGIXmVV2SFqV8xTqyIurWxKv1dzsyJQmmBN4kVXpvRg+BRvcf358PMWG1yMdIqd9pa
KujJryM0GZ2UKKT1dbJA34giyAxeujMzwxwiYpogTMDl4YN05jNKGGko/uBeWVS7luUINoftCa3n
12ekdbbIkEQW8ZWw+hEOOUaYFDQLV5FZ3oaX7r0O6//cfcIv1XojV7msA+O5PsqDW2jiidvMEaR9
GPa/9LhN74auUzWeWbv423QMAyCHrE7fElybm85dHI1uHq35euXU25E01lZd+HLliB2zB7PlEcEE
AkYWANxeprNkqsbQMFjtaP2vE/h2yCfCbkSkRh3YLyi4KYr3W0slKtbMJyekc9bRF6OBR2A1n99s
tpD9yVd0SogyeKXq6eP/IrLLvNz+pFBpf84JK7bqlkIjOITonEVhZR6MCpjbzlule5mYYXkITFEY
vT4ChMA8wfHnjhW+ukGhBhutb9m4JmeLZ9udBMkNiTBrUE1OtVMLS6WIaXJNB00Z6UVV+kZmfM88
MuS402G/Jl2j8OcjZZjSnEmGFnX6WdgbLlucGH/RJqhCWxbEk4oegrG6E/nq6/VpKcnKNt95G0ON
/ETNCgOIiBN/u3ZiG268HECjHTOTUdf0C3O2XZ4xgPiYSHPjfpQiHkWab4tRHZz4bBUqfZCmoyvE
GcH/8yx1xlPHYY0j8G3Rslu6afZlRMNrbqzmgg09vyWLZaJU/nfG0h88bucThxB7k7SkiEPPoZxf
njcpaPrcpz7ZHsSxhE4NqRBEAjgysclKWVNP7MDjL0kJmKO5CSfjp3YanJgIwOfNvskGlH7KIqox
PSSlGRKp+HNKRKvke0aHGwXPfrqhn1UC+dKQ9/G1kMU+raFpe9JxYHM52k/TUIBlsMMxtC3xolhu
ywPNdPVy6mzDeWQBxjhL3bIdIaXuz/AdXVqcvhd/md10X6yAZrVX5cvRZdvTyjcrzPktvYHnihw1
YEp8tIvc0DiKDC/xmQ/h4+KMbafbVRRI0UoKVWgoNi6nWgZJkGKzZSz8SIPJ3ST9g8yc8RyId5JA
pmvhQNsglLBk2U1dFeWb2BgI7oS9UEN0iR+wx6B6gqNa0Bk16GOhIYwPgboHNoJdJkUzC0jaR67D
AQEdMVaFc94UVwjw9GO33SJJIN6x0Wn0qSNvMi9VqN/NEC5kXLZF1fCrAA162UPjRH/vddEjNuIQ
f+mMnozi+eER4+TSR/YtlxZ6xyQIllXR//54dqQvP0wr9rDqiRkO6mlss93+ZhrI/dULmstVKSX/
IjeCMZaRKlEMHff9RryGYBndnUOMy4c7nN6AOkrMMIuIxrgM3d3URnOtTptWCVerlCWWmSNzHtQw
jk0IhJrMK/76ORhq1Wv3/3rNfb5eNh1lAhXHvP2IPbde3sfpNAgXG1e9wU38OOHINOLDGrtcEEnj
OHlASsHQevtvbwLDTia04B+Ndv9AjcFImcbzVbuBUWWduDRr+yjrwHQN2VcXVFJTlthMnaJEg0JR
0ow/rdBrH8p/eWdm5EUOZB4sHepn04tjuroOeBy0dchwpg45NpVJ9Xu4Do90x1o1e7/8uUzvuAaq
G6NfBTkbVWBxUnMQ1aZWNPojlHPESpxpV27qgOFCZOvBMoAmTUteJCQxXSNyrr8lPD5cJmxteBq9
2s5WG1YSXkwQtFUiJlo3iHkeYT/W2VVdnURoogwO7litx2U+qaLpnw3lBdLHU7X6UUDHwrU8ECdz
DwXrKJ65rZNSiU7nIuAnrsTG4LCsQvlcMRXQHABbeFNk2vmQEmFxhzWH6u7ZLYSP1nKKW9OcjBjv
/mXbnH4OF0y9voEW0d7xVmFNNaBQUW9O5/iqfOnwqbDQVHrmKNjQZvgEu3AMLCo81WgwDQLlnaJc
QkIRfuQHJaCsHwM9ig1h7DK02MK7xynosbsaqoyohoIEGK+c87QmD9I6U8zsMVr2+YXx/F/tUb05
NzY9KKQj+//3cC6cAkll0gFeIxQ0CUzqbGRrBXJ76QXRi0tL75wqyl++Ny/CyxNVtIXIXn319l1Q
FVBE5wzSJS0inII8CMpBtpXne98RunjUgOi6xSElztSgHvgFlNreqDv0RdSdLrsHZN/9rdei01Jb
HgHKXA1F+UF7jmG0SX8xrXo4/Dvr+xXjuaxB+VnymgoZL4OQJb6wuZHhhUsgeCYFqgoqvVUO9rgT
Mt51Ia9/g0FjaybqK8xoWolAOm7mJ/bB/YiaoYr24DQ7fGLn590AZZEEnf48PP5jGZ+cInKKATo9
6Cz/f6rlTzbRFgqxECvYIqgFFllWcEsyaJxYD6skLf93qZ/GQWGlCROjWpuHqVHB5gn6PqQXJ/cf
WBGOx3V8sdK9iwXDQfQHMr/e42N6e3NJuuHRaYm3U/Z6f+mSqKUx/5Vdj6ZdHuXOHGYzHn32stNe
inOxLYC2d0haS9MHCCsuUcyWAMIfd07Vftj190CE/o/afplQU7k6uey6TULBL840Sup4+iRfiBy0
y6HBZ+GYp38L/9eubh5xCyoPsrmaO1latCYtiZKzrSCuH3Mu5PBOFWf77rLnKccBYm8Ulj0wU8bK
UiYvdsJQ9Rk/1+GWndJaiDddXcmt4RD1Lv9gParI4l+0B2IxkEqwxuD2OY1Xaa9c4fDZ0Ar9oSOm
T5GKC/3nKakKy5pxgBuMdLtQ/sJs9dQMwOmqShEFj+6MB7PFKQFrPzQNidO4dGYMHMYwQrp9z2ae
1Vz/fdNlFf9IVfq8DaMi2mDhjEeZHNNf3NZ2DMNQ2JXKG/tMDWDJq5mgSPin35L68tXvFzu6ZQEL
0vCbgEu5lEtNmj8WZG0XCfDv76zgTdL/sU5G7y3FO5hNRh+/rL4ZCFcDv8dMqN7vcyHPUtVDju35
3OVxgoRiwAVgcJo5XWqJNXTXxom8zzhNntjEZ3qg33rEKzgpWOERDKQTGMO21W6BDAO+GG32OkxE
RXQ7zgGSU6uGmb5hqvZZ7OiXkMH+xG8KCwY1xueKAkbNYDkuWuI9+dXfSajw51e9VKysyJ52ct+W
A9ZEvIjnscLb5wMnmLIFMq64UsNioXr4xWBo8dmY3Q28k7od383land83vA4D5xU4uEpCRvUFY5e
TLaFo4wmD5Rw05uoGZRfV1lFB46z6tEjrBg+wLlIXgK++L4aLMiPeinu2vTApaErIfz7xkLaY9JC
nEBJXhyP1ODZmEAWKG56r7wVZ1Z41zAzUb+SPBZfhD5SUp6s2uqf++ApLYDWSgWd94znAJWg2eLo
OpmtCErAcvy8m27ehdbod9INbOaZhgHsXxf1J7Nt2aK0jCeVYod9aAqjWTqthgxhgvZBnrcxpp8t
mxKgs3DdHjbZiey7K8d3ePuh5nvBiWy8tIWoNEI9yAnL0ds+ojyucUcU7zDKBbxCCemIRuE8OrF2
FU4REt9c4ZIeUQkOxlpN5q4iVxVDPxqMx46ytwyibcdxTtVJVB1Jey1Ru8OGDOD6vbM/Dddp1/K8
iCFLhnIhQYoM7XUlIMriOEV49+NqSOXw8a+XqrCJwCVDdmcrgL2Yrwo2ZgrvrTQqaGtsyJLKQDP1
bdiNoU3dqqgvNrAJR70Hf0FU2wCSASy+nKrVgLuR0FW5fzCVHb1jGkxlpB4qEsr3DoJB6mN3UYmB
7BdhHJpsEAVk5el7yUEyZ1HHfmb0UnktVs7lAgBO3KKUiVStSr0n92hLHl0wxBzWby/2I5jlp94B
1NYvn6m/GCHbUNYz/3W8pC3w/fluVWHygUtHKr+eIWKmYGNkkOfFq56zA7BxUXhzaturjQZf5AVX
WIdGzo+b5W2vltqGf4EE0eQ9eEszD6jpOCMSfudM+zQyoekYpU0LxG1IePJebDbbVGWOxTwC4guK
EnvcKFvn9plLnlYyckFM0S5fFAkoFR6ifg6ZZpfo6iiU5Eq62WXRfHKhoRWpAO8SMHLshKAU9UVl
fQ6/V3M9zIuUB3Q8XdRH5+ZcRmsvuZTgVqmRMFJH4bXaewHs5usEWud3x5CsG13B/snnPHlp5vgU
k+2uCHUDhc8oj5+Zcawe6eaY53icUBBku6mGyuPhxZKomBCJo9f38ATsCdgsOnoE1yV2JUjSuhsg
yELYvXd1UH8bKlzQgkU2ukJ6D/xoLXDL49WNklFsJO7mRf+QVMubQNRNoP5L2g5EO9D8IZOIRVaO
SanoMLPJR80uf59BFei+pQvxqody8l8tj/uUK8ebXbRJ4gJmDT/DPHiCkoNdQr1JShgUAByz+2dY
B5+UgyGXFIvW2SVuMqcdR5Tw1DxsTcDyDXsep8TwM+bJaPuQjqQhGCEuJ7IkZ5uNtO9x0HsNrNKh
HEcfDgEK6AwZvNjNXDmqfc8g9xJ63Jp3yqd8uyXpMzK0zerAsiAaO3fVvNyl21+WqFtrUOtr0ssZ
OfHabZOFmvfGxGdIc0jrhXn38AIj0mt9Ihhh9MfOoZ8oEKp3jA0rbFX0j93fy4SapsuRvbay0f+L
rEGQP5cXJwxp9OOC6GfnWRkwx6Vm5PQ+SOAZyncW/rs6enNJIxG5YLl/m8u2bLUAsRd0aIfoOc+3
OfcJ5ow+9Pdj8rzKTzTbEKIXVuxdD6bBinZ4pu6qlUqIkV/aqdLz/39TLUr2661i/wMKATi9jkzi
scLXUP9UP97RXiH0ihbiwTTkukgEWoWJjSLwa0TbeWOw8r2muWDuBNJG0PEbuEIRn1Y1k55pl8iN
sjsmoaQywLGEHEcyDusa4j6lG8y0+J7jGsQZY6Wv4hQ31C9PNp9mVZd+v58JNb9CiMtw/MzE9qnm
G5kkO+DTiHCicZN4JndHis0EP6atTq9GVpnhivOD9BcPyaHbFw8ebLkTXwV+8ou/uh1TtQ0JSmLa
ocLc7aFs1B0AM3sMxAavgPrK8FGZ6460UCrBJKCE+K6VhmUJWfqSSwrhM4QndUjXR6IBdhjyk2xE
/rvpok2Vsru8pkCcTAngp78Fxg8xOCFaRmQjQjWK4pvIZOFEhM0GiwoqUFk1nk1P9gRWtZ+8R93+
+9LBU5t3Zv0PBN1G+W1Xl6nm7sAj2tQmxACSAIddQFwDbsaeg9XPX86F36RIabLxC3AZ7txBf9cu
3hSNEbJAy+epDATacNGevEXLRBm5eTy0xg2mEotoJ96pX0VXJeRoKDeqts2sEf7VgDZLETqAxRVD
rkjbC1aeoIDpsh1LCAa54JxwXcE0xWqDB2Nv5NngLfWkOvXscthwn8vDmnTkK37C6PpLhXv4nN14
MvoX2uHn6qnnUNdA7ym/8YSyn8CQWB1Vu0eQX7C0P2EHEUj0DpzFD8Tp1FVY2OKExmLJV1cF+kyR
uyxcsNhWGOB3dPxXglySE3Sz5ZU8oCLifWvbYCVJt52eo/cIFM+N86QVsSeruN+rAGne3RYGFpZO
yt1Bmo05oF7uOQJGQY5/ca0jOu/zZwHYdoey/1D/1yaPJP+YNDdrBgp0grLRcZpgbLkWxRG2vT+N
r/G6BeTL/u+ZJFjXPlbliRo7XMEIaVSNUEsOoGBtZriEDTkYmLVMmraWlNBDSnbW9+s7BIqxvgLa
ByxqjXfNoUJgaWlWunm6eg0asnkaDO4hGYusqnCoBHhKYUPkU/LleeNnxI2b1BrxxMJCZQb1S4VM
MLCA1iD+N6en107PolSZv2Tj/muMsO/2g3bOtj1lkZWoHvUJqUxaqOAobZTSTaX+ET1BoAruRwi6
Q1OEn7pa1vQmx8FV47nBCCZX486cymkidCtUWhTRUQJD9qZ6p3X0BkKsYbgPBjWe4LsoBGUUNm9v
SRxnR4j0B/MlIjDXMYPqcj/WyQ9ACSHHF3yVifwBbJ9xZndhrwWSd487QeWqGLJZPMsqug85coRY
w3If+fDVicfhWM/zYcP+SRIzdWD8Sg5JzqvJQ7gBsdRHmzFWflLDGqCYQYXIUMp2RhOJmpMf1mrC
I/wIKSY8N94JXjw3D5iXWF27biqbymVe2zdL2lyJg+nYaMaE6n8+RxPL/PxaVkCi0XUALkfSe5pi
JehenDGHySm55xOJQ78TRQxZYp1SkcQJmxrLSwdh2vuRkfDQyvQP+T6uU6lt3uafAi1GjiqAcKlw
lsgs7bAx4sBvSPkMxqqyLxT3XFzFpvsOeNjgL5IXxWGwUEOv6CnoJfz01QUF1Y4XOLmpU1YB0txw
iJnmgiwTefQxJd5WC4JbCRTKtwViT6UItXQ9vwOsC+UxYHO5PhID3ePvDKB6/v3CocdgD62xl3bP
4zkVgi8edL1aERQU9+7QXHCDxrMBw6d7QKgvTd5z5oH4s20UFQveeoSmv+TiF58NP8HHVFKdGKd1
hzwIdp2yJy9d4Tvz8sFHLNCvQ2ZTbqYvniCqhyLZrDqpgLlIJ5kOX5/jaIxK3HUVhoz6e/ftoJKl
f8ApCIwbG4SPUJxq/P7mG9Pmh/6kommj33ssGsCjFMz5KfTT2rUqau7LJ7Xpj/RYSq6wnJHRvJ21
K+UI/sXFKdTHogZalP22NrgMDaRDfH0NqDILbD06khmBGRjQw0TUO4rHk186+fQD+08yj2RoeTid
M6mrRVs/m3WFHX0nhF3R0xLR1R/wf6Z1R53wcelf1YIozXe3mblXGOq43/MIbTRgOfynSObU099q
bC0h31C9m51bdzgrkxjH349/CaDhrAyMfzuxMJSEEKukKPM77FaPaV4ic1X6EcBCIacm0xk2Nz3G
i45GjvxuEDuMMWZOCSzvMer5ADEj1UtFAw9JMHvZzLQhtE+DbqHVcL7ngI8ao7PKemj4zrmkPJLq
Jtou/b3QB448k7xxIO3g0p2J5u7gnXyaEiVcNdP9E234rS/oyVCr6o40YHJQ+Od+tdJMbjMuKUrW
QFbpg7y4s6c/NCTOSx+HESV4eBf0vdf+N05WFr4TdkfeUThCNPoq96i6jRhf0sRwk+27ULJKRq/1
VhCIxsVXqrIm+PvbhUiCpUjkrz3tt4FVvnrfhb9j16eh0NolUkBlZhbSuXd/3WKKPzO4eDtOnrWG
Cp3wETbzVHIfPXSCRwkjOIejt/XoMlbljVHD06zBYpHhTKQOnN88HQpfFzPvzWZUeNXgq5KvAWiS
gbHzeKwB6FY4BC8IT6ixfN4XfvkSkOUnQXVLTst69MS7mLHaSsrBaLWbkcNyz2TnHSMjEfZA/4KH
brIiqm71ueTASskOktpwEj5MGESKvGB/UqLH2M+bBUj37BibaD7iUl63qY5NSleJjHBULtyAcAN4
C1nmCSp20/XxdCGjU71RmBZdDOoqzoRbecsQt97zq2NkR28LY21C+i0eEPYXGM2mKA1uHK8EI1jc
I3yH5qOZygaIAe1AEARh1XtZtdNZrW202U78rp+vTb/104FL3O8fP7Oho+O5aAsu1yza4fEhBV6Z
BeY4ccmAcHz0WOMyjSl5bBWaV/QAy07wqvLgRVCT9hRe0bZoxxuEAf9RR3v4IgG0nJfKjpg5icS8
VI+dYW2ZTznKVxX2yzzy3ppliOJI2lIhNfgkNaG6Omj48+LZIafYBNSDVVgleal35zhGuAKeIMtQ
0boIQ/M+DNS/q7H147erusCV0MnAxvfraITb1cSb3jBu+So5Z1E68EhK+1ts9bo4JDcoRcqfdSzz
m2316SSLiB5lJlbG10HXf/3+pjcTa1E0taL+KtLEbUX9jLEsDULURFkxBuVDa9eueNTtKW1WfcUe
PjhcgFSOZ8uDJ2G0UUjr2NYkIxb3DgKyeYxg1BryXYd58DBYnCzRaqOotIYjAs4Gl6HT6DHZKZZm
2lgoWJVTATuE5khZow0Arwda7lqXB4HhNhGA+zKyMHN4QMhTXwD6YHo/7KzWcNx9/aKL7TZXb4lm
KFIHBu+iRgtB5B57v8IOCP2f4eHTGKrmxuiiP9S+bM4IIykV3Prj2bBac2xDcyKv/ioQYSNMmBNm
Mr3JXJ2QojR0ijhty5lBWRy1FUjBrhOOxUSqb90gokmK3qAeOMDbm4Al3rgV+GzswzG2dOHiHRXC
Bajt9gNdjjNBZf+ezi99t4pRbbfA/VPq3xIQNdO134snkZnlww32eZtx2vcj2dUueLx3OQhw0xqr
oGaKbXEqBGca8nfE4qKU7vSR3c798g0pRdG/YquKOGIT05LEg8HGRypORzGNPcArWBr3oUoJW+SA
AeUkPssXfx5+PsasaPYhO0Omr/0cKh4TzPueBsXJM0wjA3MjFZ7w8jlYAvnPg10XtOMG2Df1v5JD
wpzEn/3aHZmf3zGtPfFjCd0SVsC1xiP/ynjoa+DjoPL8/cyNyBMb0mEAbCo01lhBkYbJLwelnHn/
7gIqD47MpxSIwEsxyypQ7W7uHSmtJ7n19mhqwsxfaXTHxAebvYBJYVf3AhhxP/uQxO7PQn74Lx3u
bkajPoBmyt2l+C8vsGwSWS8kfu9N1RM0szUXHbCVoWdkEBjsCfqIbJRXM4w3ytJrSgSiFPTJ55q/
9I58AeoF//K3ywVFCVaIeY0nAiOJflgeGX+jePod5oLJgu1fAamer3T6TDW4Zq4W2lVRqM0LAUro
mp9OVAbl5YNmLaUYgfFRNP+iiyEdMDUt3t8wKS3G439Mj3wnz9/oDb7JeOpW38H2FqFwVZwSYpQF
gvsKNdDLmdGgcotx94jK/iBplh61dOOnOwmtqdfd4y4gFQAd47CTVAyqHTGExLF0m9YlVVJ+xCFX
2IIQEitKTzdR/c/1mBnmAHhinRLE3WVglhUSURqQbScGVT/Fwakc8kiEhMkcAWYyjxJiM3eNnCjX
vkBs7ymbkmzbvvmdXsulre8+/4xF0J69+3Pk9JF6JPHzXB6cZFFstUxp1T+4ccpd2es3EFd+br8q
y51NLO8YoqkgOLZGZlj5QezG3DTLbbBvLeohc3Fc7MxEzA40phUtRa44nGHLQCiC7MQGxIZDzhv/
2EvIct/qhKcsgkXqnK3Afd6knoHZBvmuTfdLkUoI0Z6apENouM9zI7EFRa1iRfUc+Liw46zHOIS6
8GCPOfZKym96g9txvw0ZwRJG/c9A53VwKwcA7lJA2eK6qMaIpEtzejFGAGKKPZntedl1pHRZv+Az
ossT3Hp3sa3tPhUf090sjmlW+3ER3M34Vb3oTFn0LIk6hxaW12Z+t+BjoDHo1C1bypcn2/som+Bu
HSuXq6PgS5VCvs/ojjCTyogIhJ3QNHvciKyXY94FvOkG66DECNJaGCKS1gceuCYMwUc+C7YsBK5F
eTU+I6TCjN2Ao2DFlVjC008m3P++iNlLj3KOR4BFKkO/ngZSH7YwYgz9ajGB+/BoA6EfdPDrly3C
IeRUHHs9Vm896j27f40gLalsbKzM/ECAAbv51ql6v54eK9Gf4DTqM+vofItogCC3EGxy9iZiY5p6
4IWpTmj/Hurl5aPtrH3YceE+Qauywp1Hr0IfY0ufGXHhXGER87I/+qT9U5N8IHdKGUqpt6QqlKBC
PwhHlKcSlSEF5et7b510BnZDR39iLDr3rFjAK/qv4Akqnim4JJDpVnEODOGI29ZI9fiVoYj55TaT
9RKkwk0DduiCBAVmT4JtP0/8ZUv9VGwi69tQor46ZlQzbtxQGEXMrNZ4aq/ULLM9LhMjCNcHC14A
5Gznp3Dx9c6dv6QzTcekK7fNLBqFdr313LneFIdfId9tjJwbMeJJG7o3xOxnOBZ8vHkoOfTXnIXd
v51RYP7nJNaqSBHe8Ka7htmM5+D6L/72zOAAs/LdkFNSHopWCVEijFz2eAdPGgIYyO2v83cjWfzR
NvS+Jc/jQYyNnKNF0gytNE7dfy7Ys3mxZYq6fpCQFLKVYJkN0QonLhzJEVnwjPKSTBdeBi7OWAjU
tG6iJah6ZOUEqxJztUv/lzoWUuXKlKENi9hFuBS7zadURbAk4JU4ID7UX8LZEs6Zco97SKjrWBT/
Tm1v1W4R+M/0gHPT9mfFUEHqx4JcXd6k6pP0Q8feZwbgBBjFacdWTz2BE/0mz6QrexwkZ9ZFjJL/
bkRPrZSqOv7TuHKSdJaJ2CoPsVkq2iOAcDj+Lch8zZQwrxBmhFjC3jX228q6A6kSYG9+B+WTS2gd
9JmvG50xHGZ08REgnxhiUo03mlbeIwNaRQ1YrMZEmKwkW6uCTtezQYpST5lFQiatOX6uVPJDT4Hf
6Pc5KuhndGOasH76rKl3o5LLD+et7hhuIaJh1XjRBSCfHo9JlD4kQu51MH8EBFsRCvxB/9l4JSHL
WRxtNVkQEyNIEylWYjH8ZhWdOmI8VzoT2YZRJgi5N1H1dpfWmNCsF+Js6KTlWH1NkhhkNixW5ZgV
VRSEA/x+a8rggWL1VmQmdZRK768+B1bDTbwaIQPE6X2WYK/iQR9D5eefGxYxIUmlUag8tl7LoUlj
JgzaD3VHigccufPec3EMr+VZM4UeS8WyUUf8RynEUOHX8nemEWmAhyGQDJOOfGdN0+PQORFrfGHe
jBsDm9qHg7B/Z7ITPXNTlvz5TCaEWg/mCtWCWjuRadVq3Jzwg5Iv+RebMs1WHJNxByA4apInF4YS
RDIdIyJEub0uZHy6yimUq2MUQKBXyDSleHupSlkH9Jo4l9V8Yyd6ATEFrEG88Z6BQGwk1kHvF2Z3
VO8WGsbf9VGuqPmibeeNK3QHD60l74P0IiodyRel0dY734zbfqvjdKFmOoxn6WQs2k9sDfW1fNSP
1H1e9nHZ5du6RFyt85dQtIeEDOMznwVawtzeYxhOPTi9mQ1ZTvoSSoyu2cQ5Jz6aebbPKFwZWAmk
7CqKNZFtVOELsITPM7M6+cq0rcV9GNKb4hcS2DW8iAm6vlv+kG4fSljya9qk55Oy37TCNCIpVwP4
u4Fg+7s4DIoe62GkWf+TZGUy0pIDDdFwZh+sEHqCPCVE4a1y/No9VcLNhruU+QLg+KSMeKD8ayx4
trQoBpJOmFc95YTty6AJn72b6mGKp674uCY/lBtP3JeyDAWBuhKWLb6X6OkO9OinemftlQil53Zh
3JNIShKqzGvGkptIRoElwwle6y6GAWjrlxxCpoMDVSvLwjjlunUuZYY2+PecGsa4ch/5/J1NH6hy
AF9xq++ZfwTr5GuZUMup9D6K4PLcNPHDPjx4CZk4hpgUlJyyneh8swCcj+uv9pMXyOpz+mkZsUhL
c21EAa5mFNgVJv47UHw6RvvFpYhRdW0PyWQFUG8TKlouoedsM+ckMzua2+L+2SF65/3yOFjmBYbt
m5MPGIKT1pxvh8GSeB3bL3+CJg56+9M3wyXKfS3EDaRMQraD4vrmGDHe6Pu4SpuXViuAVsSQoILI
Ljbt8mXwqhnxUandkVPmCvJ/cFmLktsxjIvv3jK9A8qaoIpc6kIJpFUDB7szcGL/5fx+FDkNpmkh
ZgWvodD/WJ+DoRepzgea6PCKX/jfhEpQ/bsxGKOVNsFc2OdAiHmRAV8HGQm5uFXXC1vOriCAk6XK
fh86baXqtARPOSGb3ohk8oB6Qor38snyGBve81OobfEMFH0zcTI3MoHL5TstkA6rOky2TCZJJqng
JrZFk8666PCWaSz/aLGV6PBNJZISQ52McWTgALa68tobjLF8wc6KKRaCkZAFHMTfuErACVoojS9p
Pt+fg+igYwt7pTXyjQOkKZ+lnY8nX0k/FvW8TGDIYZFH/kJzF1FZcgixRbtVuID9BRSks4UyW2HL
j1DYMeDQeX0T0Jkm1TTPHw/1tCXY8NCdA0vW58kHxzRvk7ecSSc+AuxF+XY644wC7vq73AabKSLB
PgNqxgNDTT0gGyWJdDwzia7SmC/EOED64UbmczFT/DolFSjjiiEnIJSti1+6zAzvGgvd7DZvOPS6
TWmflM+0+lDUo7LfWzCggjeb6I6peQCdqvVGXltnxycq6BBZM+3+Z9eyMHk7d0x+DiO4m+woYxMN
zCqBHOdd0K5L0PPPkiB0tT3QB3T2LC5hQbI3Yx/uVmhyYDtfmK84h0QKFz6YcT0P9ATyj9TA0I0B
/Q7O84Nv2RkWELqqfGxKwMVKSTjBECxF7k+uhjAH92NvLO0aPut+91gQZbfQm5woL6VSqhmH5V6g
O2HIRqKP2RmXLLa3VJbkiq+NorliFW8+Ce+ytTI2gXkPm6TfvuNiaGWvadudKUp/RAm7s+Wv/x55
n1qju71XvzG+IomrU0xQj9FqrdI12Hi/OMmkgdYMCEnb2uKuGbQGDOnOBO3aGYZeUgjXRpSLDqhx
eDBn22f9BPO/KF+oKZUTqcGtc9sq6qV+PF4ln0cpB8IulxxNA6iq56/9/WhhDkrQp7cFV8xxQmll
Z3vL7W8rEO+0U7nKN9l64hlM9mV0utUhuo/1xd1jomM3iE7NzVkGmrJUSW5GRua+yaYippe1TlNI
mbnTJQx1F7pQZwmRosGbA3zt7CNJhZ4NXgcA644BVJ5VwS3uBh3lzqijiXfFk5IbmJAVd33UTz1K
zOFpQvx8DkaJVYeTBedPfAbeLaabkBtOoWT8dGPHSpQ3NQyd4BfZtDAQHNZQ6UezNR8Tr0Z+J2WZ
ActWb2sJZFYdl/nKkCWkx0X9DOsN6RrNJ7/Q/my/ySz9EugzDb0rXDKtrpdsyFIwIW0EM9l/4tLd
t86zabI9Dbpf+n++wM7+Lr67zWpnnEvIE2kGr5O+2gm9SnqZw/FgNr9btuNduYiGQD/3lQli9BmT
GDmz3fUkRz63QU7ytAJ9YjWmDoCN6Aq1m0yeTaAhTT+b6kkVc7lkfwQyyMHcpKDzgV+VYbu1qwnW
4G2Y2uUBdmIgvPWEiExMN8Vy9zdKiZ0T0LVyVcoWKJdk4hoODNXETwemJrQv0NGtiBJO35i2SEJX
zThC9PUsa37EZzRyiio4NjlNu/S0MxMqneHyTW8rxsraJzXPYRC1xWKAFUW/nziwI6q8WfAvjNQl
wEU1jpK75ioXQ/hAkXO6qp5iKvcNBgvTpYFuUthc8V9m07tNm4jmsug9O8WClHpe3HSkR6ufchth
Kju7uvZun1WM/Sxu6tVuvY9EIEkHmkY7A4x1eqGX6s4ZoNm+4Kt6d87Wjc7x/YvhlRdKZY3bxdGr
Cws2gSe/X1gw+ERxW4EBX30oeXFoAuZr+Hc59D5AZUjIg9i6uCvqX1Z108FfFQ3zjsD+DKRmt6J7
3UOBjmPysBrlL8RFdqWB3c5TZvCTtxyjbMdN9eF1ROoZHy0ihlFzGNXxEN5lLoc771AVwZBIpxXK
ToFp52xcAuDtONODX06dkR5vog/8XnjcY3v3zSV+BYpijP+DyijXxFW06LZ1RkdNUDwv7RtYpd4G
SES7mIpgxbEl5ICZwqJEDslKIy6FNZnePF/QQUkosX7z9hUK7c9/pAdPLMC/tpWf1P9AYQCGKUIQ
0e9GMoCyWhN/pJ0mDwXRMpHUcJ2L+tL4ruvqEl7u+X2JosDVCrBmAD6sPYiAeBzRNx88P4BswND+
0fvmZ0wJ0YPpCn/BFmJKuXfGPgUlp7niGq6pPiM+iN2EDt7OIUeviO7oAmR082b2zPjBfYZb3XwU
AkdHGZHbCPvam3XpReh+umsu3/5j/q1iTVmBPTsKP8fTg5TEBFku3b51cyT86LpXykAerXGndyW5
t2J93YvzgDYTM2Bfkwl6Yb5umlOpB7jwh2SkMzwmW2/2JcPZCwj19F0SEgbWhlI1vp9O/3BfD+Hb
h0iy4nm0c2xhgDp9z4ETTTtyn6QuNtn6GHxeTFuY3VKRK7jYiWqM1uCHbia+af/hWWx1LW/bn0Up
4QCz5OFxLH32PJOd7Yys26LJI07vw2YkyM/y4HV6UFsXyd2qzhGk+SF/XnXDG5ifIBskVgAQ/9T5
+FJTYn0jDoijs27AY0U/W928sDWgsLnww8em32cfYN22D5R8irjpV9/yq5qmhNI5dCMG6c+JpGXf
DdxMPEPsBWQl+7J2Ed/Tnyo+Xqmh6+snxSPxUTKRhkdyDcTpgbLC6zDi0qUFT8ARehy+gXA6gFpY
fYW9aEGQPaWviiEeRJwlwWYiC7xLkXt3NJ0HQ46OpP1ELhS9tryCKcEdUUftzhb/EXFqOSdJT1vm
XFHwTGiZEYSSeOOKysF/XBXAHTFi61pz7Gi2NXhduqpaYiroHsbmWDnNTsZ6QOkpw+u07uhQmgiJ
RNsWv9mfG8x5km5XGkjE4p4tFpUV5jVPBDyL8AKquQsK2cAL/Q5cI7SS1+g3bn/sT3DIJdbwBHeO
VQU7TLFEgtDPX+vS1IBsNJoZxiNQM4z8EpO24jVWH44NEN1mN861P2AECiGXuv7AlkYFZuii0J6w
F/XIqoNqTN3inNyy50L4x7NW9E6YwKUhYvTgJfDANuUd5alnBth8pa8lMImsgjLcuurYt2uvtyDd
NYwqKUoUlGvoI4JLqgQIujcEKhPqOl1tux4Grb6LxRVf3XIkn1OVa+x9Aaih34CIYnhy3MccPg29
xNqyYi/3xmc1SkrNQ9cERG9+mo2o5TGyr9i8/jwJbygN29YZDghmsjTlxd/XSG+Zaedz1xS+oPx8
usgkVuAzJjLNBBGeMhsVHpIWOe9GZfQIB0LARhxerakEViZ/yyp67q/8rUzgtN+esDyvSMCe58zD
OtFnj/XPfZBQx5pZodp8soqVdYjyVvx9qev9tF9YqJVSPIR/oo8GUeLaU+bOHRzhpRtb8cSwltwx
Nb8uoXVS0sbQKbAAlwlscNwnOeSd5A+p8VpOOkUO5JQQJCzM4vF/uF8Gj1Zrafd2H6QmU0FfJgXl
oQeUgH7kG5XEvRquHHs+CK4WE+0yCwtnW/CSuyGWABfnTBSuSln1tu/GfWy9vr1Z8ZyG5+OqPKbK
62gH0DrO2vO0Iya/JzJ50oZb5/x46oykb1e5swO5f58UKaro9AJcM0XsQ4vflnmExn+q/DO844WS
A9qyvZo7aRhq7AGYu4azaRUhdvEp0exRvKFbzVkzolBeIRtCqY+NiYDY4EMLhXakmlAhjmKGxoAB
vHZ+MF/hHpasafaGh7KY5WGSDhe5q79GMYSfr7HNxGZEaR6wk7QYfqYYJD2AhpuiK74HWyWQgFk7
AWNVfcCmTmAH8rxanZizVP2MqyIoqUKVSDA5lDv2lF1miC5bEE/XKAWS9NxO6zPidE3onHXRi54w
NoUH7y43kf+ypuePHQ9KfSYgifxXIvg1QVdMjOpwuO+Y3x6h3nn3jaQJrgJkOhOTedRvlTqTapSg
/WRSiFgEX3T4mshOkRYj7itY1PHN07un1srwvwPcqmRrTuwdIFv7ghYW0HC+X8y2Cc8Mb5N18hAj
ClY+d6LoVu2t3IftMoH/z9EJiT1T2MqFryLmaMyqXgiDsQL6UDsdajoSaGq2s+mlXS4mPbhBu/RT
urrmEEEi5PoU6OQXy0zFaElqST5yylpzk9dNk4rYmXq6hiT0Q2efVpE/qd1xfkZHBO4cIBWZd7Yb
y0wcbI4z8JMBGx/VO1+2d+Irfv3l7iBeyFKzlM8WZtwG+UrQ8TJSTS9nGeuS0KQ7W24hI+I/gsjT
KIaJpY2wpkS0ZXKyiFbg7wDCykFAZRXR3V8sn6LN6LliBS5/jeQhB29V+kEwZBJqFcTAKj88dqo6
DexO2R3cbWz1qObO8ejTAItRYDr5tZl24vhmj7Men7kaPQDgHZO6oABE9L9Bmipke/Uf+APv3oQ3
0qAIbCfs+Q+Amg5HXo6gDgLBJNXLk6yPmQ1Zfbc+Q1iCaNtxeIRtk9VzcnICLHzTl/40E6Eu62sb
7PvX8EP83jAQ1Lrxecv6K9YETIACdLSaSoMgv0jtwKuvM+8fMWaohZ9EBjZaf22H7/tIyVRDLAV9
/p72xzbYobAM28+tG5a5W7veHJzi6gJMpJRlmLLcaXu6weZHWV3ZeAjqgiiRkdKdl1GUeke+uOwo
VBj34Romc5MiTJtPh3sft+bSR4Hto1O4/JUXnbE8QPsKbAu4yIF7q+CCRXc/oBAW/hNGpVFazCKG
u/Z9LyMBbNfcTG/P0E8C0K9hIzlJsW69QFWJx28Ivl8Ecd2mDmV1bctXVJcY7hNc0KXhinrIs59x
NqwEyn7wBxitz0OifAZz89aJBT/JOnq2AOwVYTQXclqf/n2cgAxFAbZHQ6mO7AjdpuGtv5whf8Ah
xKBxl0EwZlE+TCx53VvJvheSdAcE7JytwvA5YfPnK1MTbexLDwcJUN1GvpFQE4rQlETPoQYMADgG
SYvOdhI7y1FjRMsiLwAlyt5BS+5qTDpaVn8TPQDvVEeNuXLsP7wxvr3L3NwBQxH1J48YoBZ1WgYI
RdtqpgmDTBZNXrILx+2Xom/1ctlovXmBarw8XKNaiJSKsXGR+O8EXUrcN+O/8J6Cv3S8szZWMDOU
pFpq7d8DI7OdnnNrLncCw0qbyCTJVj5Jh/8SLfYn7y52G/Ed686uO4AiA9VgISTnuOmDeJ0FbJ+E
WVhlvC1R5sI1/CT2IqDCxX/+XEhsHpHfv24UUBymG6EvRQKS2HTyGNx0gr1GUbKPLUYHJa1ARkbE
HOty8xuutvSTNS9CMgeo5f55A8z2ZroRGCnGj8oA6yJNVSDErHE1C3yHEMrTGLy/SVp57xqsrHDL
S2lre7SqcmIllheC4gI+VcbculDxnziT//DeGTPLkTFJ6smbq9x1WPUk8nt0viBJUjpq/ccpi6G5
d0GfU6N6KtxjepqMV+iwbk26umpcX1tZSwHLDkBkdU8aPLP2BDP9Ry8hqZ9mukXvifyVCFEmbhhT
rTQIxxjLWnisE9ptWJkzX3j/6kooJkR5/qStxxAW0UPV8+R3P9/vJmb5do67sq5WqDiXQfQ1ctqj
ATc+cFVqMnzoWYMgIA6Ejiweve94isgKvCV8cG8+JBHPWidg742wwnxIScC4fSHY7IHPjW17+i0B
TGRHnZzBI7/Ma+Wgv6rJ9XZyQ32Y353rPxJUnpseeciHBSsP2Ucm4HCA13FPjuo506cK/da5oa2f
YapuaBbt7ZgUIY/7l0DRh545sUcte8GP8dRsyMilN57wspEatM5JxJu9CMr/IE1E3lWYOqeDDNpm
m/IbYTW38cdXNg0PdD3EzUitIeRQpuQYp1w+S3bPkaKWE4Lzgfssmd+v95O/GXIKzNUVvpO39u8O
a0BHzEwFTdrfPc+yY7ipESMN1g8Z9OHrm3PshFonYrKV9K2gS/MyaOIWr7/oEbm2YytgMts5z6dq
bOcyqNHWzI+iTPveLSWUphzG2VfabQRMmRI9El7BjZqXAkJ+YckteQPUevgnNy8Jcz2p95jip9Jj
WmX2ww+XD7oWyR/GgXUTAHMKkQXXnAEdt2ZCZCa1hZZPWFqKS5QmJDXNHy5Qa+z1tppOXRTc+zYr
XwgVGHWwPo3EYYcNpdEt/5ZlnT6Y6HYfSMs2nIJcqKLmOE+noeINSmaYhqUNynAmgnJR17ZdyJYw
kXq1AoT7gueyWh8XtbGCFSMLoWqPowjeLhoZ9oCaCi0jt6dJgRFwCK+MalN9S56mk0OECY1cx6Fd
iacIzk0DEDvykf/gkuDybjWy7RfhHvxOOXJ7oNKRJt2FL5p5gZvF8xFENnAymTgQvwWivxPTn96U
KkqnImzynrVwGb6xparfofXC0Two7bAR4ujlYhXWBsDmmqIh7WoqHJJBtY7achRu9RNKG3Fx+0ex
mXx2IsKTcJYoY+6nokAWdEPffyiupdaC5vvxyPVRz654OFVh/x7ndpm4JCS+0SXE4QKDjP62U7XW
7kYLl91oFk/pNxINKFja22DMkyZtt1TGEUQG2Xas4NeoXeKUPdHKsmp4zjWthsXtkLdrPo4KUeg0
YwruZxQpBTqt1kMrX8bpYAAp+ewEGxyWc4o2EduqJ2IdDIGXJxsnOwvZgFeeY+wvLWrq7ZLJW6JF
RVZFHg9GZp1DCQKAuG4Iw0yfmPWLLMH4bqT24Yz85+fvf7OYV7fmSet6C2kBERhnv6q2tz/kiRBP
m+l1OCKjNZwfPBQq2MQKYMS3n1tUv+ZndW+VRXjdJzL5MmU9EPMBa4g6JsB+az81N28JX73ZhHzI
oOTl6WVQ0WW5ip/N97Fj1bUvevcjxGrkTqZ9QaCxav66Yy+O8l6wiWDE0XqP4M+vkOdZKGKsfet6
MeKKtPqt6sxHZolCOVd/7j+u+MREBzqUieT1T6C+2PXIyvvOfbIXyA3CN22y8b5HpUcuaQbVk6p1
IFddCdNiLGgClWPfF0ChbwA4bHqJQJnRd7MZP4+gnnak2+X3sVF4AWjQr+MYAS8PqY6+A+DRHX4q
nGxu0TvpLhoUuvvWlz/yUbIgXN89dk2dZPEbHkE5QtA/rS5RgNkLthEDLjU1h62qO4y4muGJuntV
iiWjik8p4pelz4jXnTRTig4rJ64nxCrMsTDVVEuN+tkOwvbtPK06Id21/zc5t1FzxKyOHOJ8BpgB
Q4Ov7sK/mQRrZk+gdnr14g5M5TiUQdlGpyVRt0TS/e3HEi6V1LTVqCmKg4/8IYA8peiyDLziKEGF
MJ8sji9c9nbJBvMpMQxAxUq+PpUmE6SZ7Zg2Neru3i3eeg5+dGgwyz1kCFAGwkJwqqOrdI4vL8dn
TqdbDoPqPZdJzdDD+FekiUtB4+zjbiGX1CmYuyJMP84bTX9Y2bdytoKCo82DaGB4lRaoOChfobv0
Mezt7euHwSC7a4T+of59mukJQ4GSfmkAY/9CqA1UtcJpzXdZj17E7jUBStagH29b8ouPkrNzSWDY
hYF50r1baSvhZCaj0B4ik9rAU5V4BMzQqelLmsyuS+gK1f1gz0m6T7y0wMyNWteFpZC1417gGD4L
rbTodDdwTLI21sz8A05YNPyp2kTpvAIa4GGyMNASVc7wi+v8wpRtvrJ5FNGKtbtTdcRf0KwNHeLA
anUNAV9RKoMe0TD8y5/o0WFglsiZzJOceZKmvPKX7pcb7nmEqeqVNGHSvJCO1nHydHYko6eiOdPS
x4WCyjiJfFkKIS6Ay279HUosKPSwbXm/XRGwcjD0541MOfhyJBIzGvn9z+Ro/zudZ0BmNjNmUH/5
6mjm1uXl2qOeShTYkugg1Mm4PywSuQkqYY9csoZwwVyj6XaDvRSllL8zQnvWE5IvwBf3lxs8T8Af
Zqepbw+5K8Tj502cV5xItAEvf9w+4sWp/VAhDCUSc7NlDV2Coq9G87bLVVEDbwItWUqNIIxJ/Gg3
6yXqobwscMm8v7D5yjOL21fZfT753kNj7hCwQCvh6rSlupsVlIRIlixa7UFesIzBbvYGUufzUqKT
/Fns3Tj23ofzHNuoAFW8Iv4TY6SyP7FeAqy5KeLdBZWBsQSevR0xyfWqAoxGYaYjr445M/AMOrQ1
KsrOza3FkxNSuVwQ9sgsGgm521RDxBkgscF2T3f7CUQ9E0mD9rtT5RYB2Z0EnOAUpqIGfLDMfNu+
FewIspspvM98Gt9orKnOdriBk8+l9/EPHB6kash6NktBx+XyC7WthOqrQtflTuuLmwrmNLwszT+D
wzmogvc7mMkbqQSEumGSge3vU5btSJJ/KGO6vpA78zxZVvbGmukAu2Ijb76FWa9k7K5/nsG9u/SS
SIhGEYyU7AFntPeY50wND4Glgn/cDVBpVs4hsP5ALLc6ebmAVtS4zaAOE7DjdLZUqsa84SD9bWVB
Yg17tTz/xJtBkz46+pqGg9gRsO/OXbGjFZuvzvUYkdHVKYjac92zz0aDbQ7bFdaqxFP4C1HeZkm+
XJzx/7Tz96XRPNLAViaofzhYryUNE2yzr77XR9gESMUMuAWYQSdAltuKopOtmdPSmH3Irm6QEAZ3
XvSvmSlqlJW20bC/A+zS/VN6FQQPSsBEYIyS703k6WZkmc8o64zsd305kVXat28mgIhB8zuB2eUG
YyaIuY6l4dtMESi7H55vrWzxpfpwn804AKKg4ED72JZMIwkcohNR8TyE0F5XnTO64c3G7cTVq53R
e5mPXDns/xjvBCToxf1oqzpsiSN1JpNwt2YZdebCEgWx8m8SKJ3yxHlREJ/D0KYo0Xz9oGUXke+i
e/wrrpJ3xCNCRjoCtNQ3oPvsO3R+JB/IpDR5G07WISq/TfNGqP/TfU+YhlqrGAXKZQ+PLUFBxmr1
iZSj69f1VntI099i4mI8/9Y4zeJy8jDFR4SBoGQmKdRzCwEpQZB7dSBYRr75Yye0wDCh82CmFufj
qzAdMAZZxC1mfXPta2i34sq9V5hpYHgestT8pIkR+zUvITLFfiHvevzvBxwVNICEvkPl1dofYCUH
hF6oS6KzM6Uqfa35/x3XM9Ttlb90aYsAtE3+xekuXGDQvfg9VIHDHNkMM28Aw6uiDNPG29NNx0dq
cI0/6cSKJjgSV1fSxJ/cFA4g91fA0mcN8GLOyVq0GYhAenHqE43FSaEh83gC0OzWf8Ugw7P2Ay+G
Le/dy0T2E/k4iKlWUZPolHxJUc4jDPeImcjWe1Mf7N3+v6HLu88Mxfs7BkDpZ/YnOJ3wXWhoXlqG
oPMK2s36rAeLOTDPtrf3Vt/CQ0PajBUYFjEOdNFEXo3b74p329NOtZBZ8Yg/reS9zGjougp0ilFt
ULw7UgA4UtKOZhbTrQCCQHZa5BDd6JOkRnVPKnEkR2GyjCmnMNDtguDdjUhQkAMHY8UMzBaLvdFw
Ot3rdMAijCusxmDPouLFRmvYk+QBIAmgPemeRpj0BqBR4K8McwdCgE1jE2x6nHgk/o9/LzJ6CNpU
WQcUJro7vjYovO9G9cstbZ20yfZC8x/LpVc2F+6B+6O5FhiK0SZcsnSPHTcavOZro4ZNlrW/0umX
pIT03j4iSA8GeNElvieOwdrrwGW5PaKNzZ3FHh1Jy4VzF/yPHJGrlcoR+JMjRNHtKEWyYmpK1mBe
I0rJ8LylzGem10ajtwVfz+oBkaDka637H+qlniGYux+SeDfVS1wspeXJF0fK5PVWrgE8xY03vPxG
TTZBNSgNjAVXNR/9cu592ogKmX5HSRofccz8IMwdBDlpHv8QMCk69PVZ8QRsniVkQ0SV//ovnQZu
d7MeuHeASA8jL6HHxUtoPN/iKykqomeDFgTi9e6xQK+OtXN1/DUfaearLGVfrrSpS8HzyMoBWsvt
3NUE6Qw9XYDH6u/ARuoCd/cQnsjpGKCkk4y4TtNZIbT26F/TCuoy8HgDl8RuDV4jYdxR1DHzPn+6
+QIji/a8o8q3wpirkuWqhw+i+t0UeocvoBucqaPXdYsgXzy2JbhIosYlVnqFgOgWBBB7Dv9rpZfx
sotP2nGD4zWiNEgeEIE14B6NuWfMlUfCrZVnLTc6aEOv5XpoNPmhQMg1JYSNr+URjMwwXvHcxvBP
BSrKc+giUJSP7jS48Hjv6nof6VSQCwsNAUnJFI55KIW6DHhNv3AgOqJ1fleXh6AMKTEgtfWVsa4N
QE9lnTTl1mmspV49wS4n4EKx5bhKDnlSnc/grYCiopwMMaobp1xhyyYXPaJYBA7sFkN8Eshyfti3
ZOUtLMoQrN8maa5xM4Iq64hel8vCCf1ZQCYVp01VvxGu17Xdbdwa2j5GxabwWyV8J/yD4ja5XZhV
duLuY8PkRz4l3G+9bXLnmVGnNNARoy1VgrHVfioI2tgS+Zxzi/tUGbpg15d0yApETrciG3nNajOB
vpA9ik6DLUtPPYGXTTOyvZC68QY2JsPzp/w4+/3kBQ0YY9msPDFJk0e8DwlrZspyjxkH25Q4VzBX
w1SIVB8tx8bavZxXRjsRMOyZpWOA6x0sl6wvqSVGLn2SSwF57F8W2FPZdrIURiTfUAVQ+a3prJ3B
gmveYhK6MDsokVQfHqXXgQJIzgZF9cB32AFsHO4D19A35CxFPFH5jY21sT8A6AH2O+cnGjobfMxt
xxW8w25QaHkZvn6iO52QzP33pNkiRySv+GbS2NJ1Hsadx2V4oExvyHGpMX0zz5/dpbzm8XYQTEpq
FPYMt5QhWHD3MWlqiraSPs82v2IftbZBHHocYWhupnqOqsmx19LiLQDX7dAlHOPxPMBQVwAlaEoz
Ozsd1gTehQPXGyBQ5r+JUQZVaXL8uboKklsi0VSUVskEuB/jxxayhLSpmwa7v4KmQQ/aKFxQyPym
he5FqbCFOUvnsw89es2P2POLnlhjT/n6w5rNUlNWiAdy2gpRHjcXDg1DteAugVgYWEHYlCLkbrGW
cJzFxuYgcsnI0mjR7CVB3bJQUiywWnwB9LB6Lj3ULLCfDKEmgkbNOI7j6ag0ub5JtKoE2Zn2abnM
NZw9u+2UHFWXGF+qZWapRQHXUYiPz4ocY5hhWbbDMLV/dnH4AOSVt6Vds/RRVIlMeqLTxF4r9s1L
yoC/x9qR5eN9ric99y2YEo+mPZOD6e/0PqtswHYxgT/TURgYu6Fs57zjsY8flQgioXGtx19rxU40
enWFS/h1o9JkUriBR36x2WFvOdBP/6NOajoymqDrQTYhY7GlJ2Ru85le8whxxlCPMxCncvU1DGEK
9lUu7kXHaMKlLozPWn+nw9PCqI5Wko5bC155lNuvhcKOfvqbc/rx2LXA4U7p5PQz+5W5cpryl5AE
gifyLLm7a74rGtxH7wWAa9KuUAA6tgf28oGMY2Efhzdio8GrSOHfkuzoRqujRKK66nMZGFxPMVi/
Z+8TmB2o1+6N4CLtMQoFKkc8vPIyyYuLjSQa1U+uNbX+wM3JM7pETbcNMGJ4+S9hpMByi4BW7ol8
6tGi55Lw6RVWnFJG/rXSqLoapmOOVrqYT6l7QKu/qzHZh3TG9nfTiFXN3sZysJZEtHbHLNI7zDPB
X3VZa1GltwzvatotCvIa//eiDVN+q4Ink009R0PKmWwbiXhGTCkq4yVUnrxR55ohSQCWef5HtAZl
9kXwathcHhJMVJFE4KzRoTlgv15LsnjeJz9WRfcKlRTpNAOxzLQ8GvBvzyqsNLKcBbf0t88ORPK+
VOiznzcO2TfJy9T7E8wH0aEOho3vn2V36BxuobjLqTxitUmNjNFhNkwKySm/hDwGbPXVpiyycZN3
yeuKmZGBQImad+wrbUmjjh9nLfWiA+aGWG9xLwqYOnQDFx7dRG3vsX3UMSVi7q0uZFjISY0RPm7G
XbZrWBJgUQb6I6DHDxq7MPJUfCHu+i2ifXCgiUaj8HVBnoqNMOrOPuq/u8Fa1I2NEVaa7x5N/+9Y
xX54sJaO/UBvpBgoB+fO4GUSbMCN6Efh2XRgVrXrKQztjAKJDbCj1pY4GEH9weQG5XJ14n7d+5fB
IpRZgMkHo2NO/WP7WVibahRO6GToCFqren6MAwdytGZJ/sehbDrcRcSoipRWQPmcOEIjhle0oVN2
wsqf49R8FUbYjCt5m4zBUPMp92BYgYpaPzUcZh40HLtfRH53N6Ooodp+Wn4f3fKm3HqQqXPh4jph
jsJuNrUa1XJ4GuIq3j1blWd937YgzIe+eAZgHJZmQ0uHLH6ZaZm77UTtHw9FmWdSaCMAe1xg3PLK
TeFiPByaQApeIqlEqy+9o6GKAFRTNRspX3g5urWDKS8LsrT6X0xfZBcByfUPYzXEFnl1X1DjFzgz
AHdyhxCbRht4tvhV6tjztR1sJI+uSWhKWEMzaLbmzVG70A8GJdPxmftqOFtfpaCizJ7iBybhGFLV
pt+lwl+dnfEvI0u71qIGiCh9lj4oX2hBaRvKuyu7SEDpMkNbhfCOyGByB9dp2z8gt39j7R5UjLBg
ak0QzU9ZwFKHqabA9yD1r3Aorgqqx0qoXy6sPsZocmUuVQkStjjcZ5JSGEhlTEJqjOrzSAPHtJ9U
pu9UxISLgyrzlYE/GU4henUfOhyHAH4oB6/J1BPCbLXO5ukMUQ5n17mGQG970cBw2zCY7cuPbm8e
otDqJ8GmliLDDAczgK5um80Iub9P8gmfhjZr19DhOXADNX2otx7kle5YPgzLv63Jg0lrdLj1mwKx
5XcAO0sznEP4/dnM1MrZPZW+Jm6mo/Ysfz8ATZZfbIFNE+wNO/m+m9YqnfK6STUk+fOZacERt9kT
TJtiRqFPg1LLMVxE/+vuRqs11gGvMEBjx0mG67VXL5rmfTIY5ZzggzDlkM69By3zexPHoOpLntcD
fAh/Pv1iOyy2zsd7G5w2jE7A3S00I+pjZ5jg2yz0X8XjnK3+mkhfOQKz67ZB0BEzzmj3VGOxxEOG
Uq9W8A7E+Jh9M0yciaZkFhGetpOALTY+E/sVicfEG5DetXtdMtp0rdmNNEx27RiSDgqP0mIEWAh0
kOXspr7lH9+fkPYh6knCLQzDRJSs0mYGo7fD9TZEsqjRr4zgwpTUrnOB51sDhO/LcKOgJX6EtzrN
wlRb2NhfMN0Ni/swzkqAjZILO4YIE6HwUP3sTzkjPk2rYB0GyXFCXFGUi+yXch3PHSwZRo0gyxH3
q0LoqqV82ZxH736zYBxQJ0W1TgjvVM8Q8KgvoEWyXLlZ/mE0ULZ2TW+wbafs4tBJg/kGL7Vs0YTy
dLFHwWXeytJJd8A+kxuplc4ea/wEwGjVmO7htfkKNa0uqX3Cs1WyR+PBXWdJUGIaUnkr6dKR60VX
xWzTeC6liW60tdNkcBWc64AOUrqXeEA6QeeyukNsEeBGpRe75Kj/qbyvKSLHsKj4FKzDWkow2QU+
C+eun+r7p0shijp5n2s/TqaXkFUfGqnGgNQpOgFBuWjhtVIaA7HTkgpMSClpD7lOKk+lngalOGY6
dISJT+GJ/PoV6SbEA9YGPgyUYWlqiLXjyEu4Pujh4f7PC2ySmo/xxHBcZPWRDUpnqfEPX6bl89WR
AjB7WYlK/ksZD/CpQfYToRAUPCBFvZdhWYS0frF0PN3oO7KvKk+QR0jNQD3c0cXToATrDtR0cYrV
5ImHAND+1wBsbBs+NGmbtZ69u8QkpSVQdq/AkBnNcjTzbafHALKwZiRyWrDWFKeHA071jCJ9MmjE
tjmreZHFmgoFjz7X1iJW6tcLKz/KqlfzbfLnR8M5YCfE4OdrtIDp+bvpSTrglGv9vygWPMFg43Uf
AUhtTMoHdMatkITUN01h9+vwZbZLf69zehaCfYlVG3apELbgv2Um1UCmNietehbns2pVYObEYxom
aN/oog7T0h0xPvx6wIN76nlSMsEgMh5vCfdY0ih0YmYTO7Qdi9OzmR/0LW7I0wUIq7AZBPKdZbLZ
w428z2OXGknlIknMufw9lO5G75m18yTgiAtM6QBDOe2z2IPEN1hyG1lIpbYBvGnABW2LyFtStxbo
PY8YX9dpxxxgOrQIP3EVdd+4Sasljg2K4oQPMb1vsBvTuhE7F7JaO03tA82f6croHbWZEGND/s2k
k7q0vjcUMN2n7YQ83ivdtENWYROWx0FBmA8sj3jQLvnAVflZPVxMHCE++vT31Q+Way1Q0COPMrwJ
hjc+YkIyfsZ5Vs4kkYdU708a1eUM+06OQ1Bn1dPU4uvaIvIgZcGO7VcwxE2oXTyeqpU7o2ln/cgu
X0MDIwntVELuv3zrsynWp70FS7FDAg7TVd7okPkWgQD1/sLGUmL1KMehuYrExdWaAicnyhcAaRMM
NduXsdp1pAZxD9GHG61V2YiMDoN3CufySzLkI8ar37N8ht/MCCfInd2Tea/UeX7Kmwpja49giJAK
g5i/yRXL6TWm/ZA5hem8o2GFgzhn34MQvy0quMOceN91BRtGr5nxiiAsI8W4UwixE5KaLJSM/gHn
bhnrdiZDv8ZPIpH9hcZydHyhUHxgZ3DTymlFg3Mt0h5yAGD3hO+saUbhCjni/W3d9/rPq4tHkE7p
RvCE4OTe2yJKtcqqEJjwoiOi3hh7GvRpcRuc1b1SJ6bK3Rr2yIx+qC5ZEwZ3vq8uqzrOe34ERWxX
7Sv8mIC4z4nG9YyQ3cYzmfDmXmzOfcPND5QMle7DxDpQht0EqJISA/h04+WBcjoaQtY5HLcunymW
jPzmCVlAn3lZF7liw3SYWOXTrg90OpVAEtZBUPIWfRPcG0JTXc1ikxcETEUFa+3guqacCN3IT+Kd
+W5DGWJh3uLy03aCrcuD+VKrdGTrve13qEriSR3APTv2nQm2b0X7XeeZ7lvlJ+mf7YcrqS234hE7
gPkDua/gvX8Ymf/q53i0Vj11LOXMXFAk5T9Vlxibkm14t7TgDrxh0S3fGG5gFUn1zjHxC1c6Rxt4
1dWAb47+mcCg0v8LbhLV9ak58/+2MYgDLuV3+dK//70yGLjBlsV/xc7NxJPvnCiJhZJCGbGOpQpV
64SXvUDUfGvK7eH4fJpRcEfSnolXgka8ByS2ZYtf8ZzjrhPtiHItLD8ecQB2ctT71cy8QkFC+mPc
o8m7FduCeuo1W+Kk+qN0QtFLZ0fiIO2khP46q8d1MtBGgmwYCfyvEPx6cLAj0+69Y+yWadLJKP5s
vM/x76yU9uWLqTmAVHKaUjTveAAzPDWZP+utxci3CxlmJsZ7uTTvuUyp60njo1jnmOgZBhPoW93l
Ih8tUUoLgTuyYGbeeAQNtr1JPTRaqSBfIFBdGOF7A0VMZEmxXaa4oSrt3CI/nTIMnVScgoyBoy3i
CyBq9a+YQK2IZGnho0Cug6+cRJMXC2jQVC6gw0R6ZXYB4FnYf77UHtz4ZM0S9k5YQGDtrUDMTzRz
LsCmPdG+1xvPMn7f0AIetRQypP9FQ1XiHT7nZzZeo6VSSTYOIebmaU/JuvfPIsklibyCtdtc4bJz
Ajcaq9hHNlDGNJLJJHH48LDLky1dBVYF2gQgLm2GIfYc3iHIkrZivZTjxii7z924VZt1hOafpnjv
QbpEiGFOopNKlUf8bI3NQwiL5HFnkJKwsRIMhFqodwLcBFXcItn+iWp7ftJxxKn8r9FB0VlIuZ8e
tDH7cdGxDcet5cnDT6LkRFYRYZppnOqSsOwXJoJQJ8ognq8S79y3qzIFLjpUvTMuRejKjn6pCrhO
T2fKHC74quhi44TiFuEjrh+rwV0kZ2fQ9/AvkL++n5Dq1gZVXrgs9U/fKd9zoAWBF4zMU2BX0EIe
Naqcxc9J/Wm/Y338Fln/x44b1dZQPAvUQQ3ibVrjmu299z9UCVGxYwpXjAz7C6Vc9XDTQnheo+kP
uOct44+NmA6f9H0ZrGkb5QkqIxJ2URGgbvmx+qSxsWWI63088ZkImTZbECQDc/lpbq3QJxFK6jtI
VTnw+RVQtsISn5/xBSNtZgdUv9QGrJBhEmgcIpVr6O0O+e13GIPyky/U6T5KoXV+iUGzC3bAsxsZ
JlzGmCtzTo1e7krc2wnhVFjVL4sVGd2W4nKRNY8jEKOX1NxxBpHn+Rgg5H3VAuYG2yJ9C/Xh7RrK
wtXRDbmG2N72QBUpdEZg344/M0k6Pr7orf8L91tWLDyD8RZjXG2zntQQtozFWQ5itP8gxe8z/+TY
Tt2d62OC2PAydtauR5WNiqqVhJo8CaC36WFyPaE3Q7Ff508i1M9u/fXFyC05T7akm8MeyyRPZSgH
sR1Gxlv6GfcBiWjQNIuPYJrG2z458+CicTzvfvTIzLVldPn3piWHx93svjSEdq4q8OfXu4BrnmjY
CXUC4escKtp7+1ZtommtikkZIonq8xkNQRNKmXN2adftNhuL8pibNRDFCEdWOh1SDpF3nU8U08k7
o7R7oeEnedXXLG5DVzwwK32qpjALnARXZJyYdcWCpo2VQXyCngDTfcdgN6IjOXdPRXZrIBrw/0jN
VBU9gaOx6P9VPcsxvGtz7bgUr3TuyyqVP03TPdvI4gURbT3wv/dV3E9DguM8/zcjEJxClDFXtwPG
HSSIPlZagwQtqPwGgnytn8TIwxUIlcyIcZJ7kv8PdOcSxVir/eGmcZWYo3OVksBHTMbzNqQOI/Kr
wIFSThka0R+SFedtLwDYvzbCcrb0ZNfJ698J0E7KOOrzSq0g7ft9+YEsuGMXWEzH6ezhZFKozGgk
9jxkhVK4rSc78ZLsd8wPit5EaqdeDBEFqB/2TUsYInKnPI5u2zorM2qIfSCVVU6TZbAiTaWquxnF
G19FqlrukA8V4BdoW1kt5hvdzb8Ni0DvbYebdtz5l10wqqyWXE1ir3SkNCyelOwq0avwaF8qUqZB
UFcfVlZJnFxs7nwmLVkKjoYm1PZn5NfJSObsp9XVZcoQ/MrZE9rq06spxmMDha8oQ9iWRJwKKTPC
Y7hNa8ly2qg9gikBG6uH+x8fd0L+Ycybues+pvaj226cwnP3AVYqTdcy6WluBAFwgpd6oYXFGGyc
1qFc9Fq3xrKYNXCSNZVq6b9D9rNTdMqagX4XTE9uybJ30AJvQAyPWRylDD4bggBQc7uqmWjdyQ9Y
cAip34f1Ga89Y9byG1x07rCRWduvJoVYBIRUJ8oa6453s/EB0Ub1NgkUBHT7yakdcMT17JhmoYKE
+3WvpSZM/M6VpnTgd/ioMCBY6VFfTOYetG+zKspMqjGihQDFVCSwl2eHreF7T6MKFkX1nCazsz4q
LYkyQRRzS8GVu6oZh+MBrU2wTms7oAidLQ/4ZmMtZTmq1wfWbovjikDlf7AGdZ6UymrHYOc0WFFU
L3TM63Lx6m6iA6jZsLuqQfzi1n2Fs7Q9ry4LxttTUZmki/NgmeQ/jy/5iAA0wXyDib1ErCv6eTHO
id3pUxGGtTIDVB6QLFBOCnQq+4gxX8kktJma1IuNzdS0xxtR5W55wAIUwGlvhYcg7SrsDJ2WbrR1
rVPUkLOeljyv86ewWJbKQIgIADhDjy++Krg8WGWUQkyeCbcolb5Kp5wR51l8V1HZgbJB7jCDCGdF
R6j6x006igvAigpzzSKoc/VUzrLPUeZ6gh3fPIApkR+Ua+fsNfrOXNV9CBmQ6BQVe/sR6dhXwivz
8BUJfnAR3Iw+uYhcRRUBgg2CRvWnSCXB76V61OdP7ikKFe4jtCBfEVnqnW59R5o9Lj0KphgFl3Jd
fyazu0uqPCD90eSHTNUz1sMvg+rRYu/iW4OrprpRQCRBIH6MuHOHhzPwQGASl4QTXKA+ips47L7X
ytW+4nuSolXTl8NncHgV7eMa15kIyagoClF3qhoMX/RZwHrs/Lmtvr5kuiU0jehTagbz/Ev+5vU8
QoCa7b5DAREzQkEGNF13QVfH2O3Smx2ayCJsn2kuzz9hay8+PdqUnY30PvTfZ1agm83+/JJ7X9kC
ahBjScm3M7c5CSt3GViP7Rbx7XhRWqx/4EFez3S1itKteaZO592odddux5oUp6w+LIcbBsSKxJt0
wzp+uJnmMh4Vb2EsYf/mWSWhMt/KqN05ATY25ZUMNXaKg3LEekFJgLM/hPk+XGyQqh0/1LnlJVFr
gWf2STR0YZNo+kzXoBz35lEiqtZAX7xBRdXQfCGmx3e/7wWKVRBpQNlSoJZsYfQaKm8yYCnKO3wL
rFpD496UMj5T7Zwfiatop1bjZZk+v1h3rKCC/btFron8efMGVjQskbV5768wavyehFQrlQ4R63/q
akoQErRbktju43MJqi5C98AgeBxux4GylKxXgkubiqtx6pQOBX6Fvi1Jgn4F7rXGlhs+eJJLh7iG
jW8mnJuAT/qVgbBC77Zvg8SARw4XlY5gUV2Hr39R15X8fNe2LpGFoLearUQPfodH1gaBvjrJ6MDQ
hCItKspx1/Pu+/ipgw7Qn6ToLkvGtvfS7ikGQ7n8exjoMEl+OtWfDht2si5dWwRQT3SkLaZdVA7o
lsnjX+1fzfYEGL2f33ZUXw+YCOIr9NY/bxI02Mw7OfNp3uLG1IrN5WLGjSXUYRU0+DVbDCTJNXrP
YJwwE5/DAQUvc572sa9qzJkZ6mOVMIFb0zICr8NtfXccENnBn61UTmgrji0xcRxk5lNPUI7xBL4X
y0PSxpxuwHK7ea8RzHv2SjqVDpMQP8H/ZHPoJ65G8EhC4uRsRPnzl+kZf6WLj7Z8VeJgAqd66hjA
LP/o4ecnPni24CVo2P9tvDp6HtpS8yCcG2BhthXoB8i1I7l25ozZNkOj7jfPWTDeCEOfE7j+fxq/
hTZmWDfJegCazEzS08SG2rhsrbDjrrSyyoUctUNMl7mSiq8Dz6PZcv1WIHB04Ew8/WTl1hNs88gs
GVhAYyJD/LcvXVHyZTtNkdwkUlA1pZa0PxPZRhAtDzLUMb2RlK7ZiYkH8vdvh+KNoYHHToqWtRBJ
vu3qfmv1SPIAuJdLobuDU1N3KIUUUZxCiuv3Ncy9XdVHhGzC3NnZO/kZkIll29XV4e1ZX7/wOqFP
8HDfqpT+/578f942biRIO8rrGDiyc2B8MXIDFiCUv5sR/3/u5fkzbZWM0FzQvigCL/Cl3jziVrBI
rHUFjhcK5I6sKDPDj7n10aI8fuuf2erXBk93t8gHRafvBE8IZSpP8fuhKch0GUi6T4yx95gL18iC
21NpYSYrZRAib2gd9Tc77DmiG1Fz6HzN+I5ch1o2kVQ1vNOwBxFBRb/0497rdqfPKF+faXgOfmQ+
qaMy0+1XN1qhmZRUS41BTfaWD+4bLOlrXAQ0u5CyQrDtxXAfck1oz3V3BzPcXP37l4s8zC6jDHCW
4ZEviQ3Omq+C+tw96cplS0zr88VYv8Qf6HGLySO+1OInnxz/qX5409SSeIplMWWIMhN3KPZbQicz
E5PZNf+Hffwzm76USCIQOnw221ZxPK55Eoc57nZO4FyXM0ZMgzk5caRcYYfd+UfeLy6kWSVj8i7W
GSy0HtOzTXNM87HzuSViyu0wAu7DF5+Akb28PJ5P0Ee5cKB0HSTyxXk33KNbMWjq2Bu1vz0q/Vqg
ltetbUgg7BY2hmZfafAosFrEpK6ARoXnMjLW8k7iHjlu6mDlnltcAQbiNnfUB0t1imcHG0Asm3ID
o1wWPe425G0yVWe0oaEabm8zjkijU3S1qpbT4cTBhewmQ3Y5JkbKYcAsT2DrjV11WE8IUEzMre2C
G+k9e7VhJ7K2MCWHdI0r7U0OdNA6OVhmQvZ4vdBulErvBBGlH3NmzxPVmAo4Psgt5g2fNFevEEvs
fuMRtGRnG9eDgvpNSw6XmA09fOnBzOc/Er5zD7G/uqVYfpP8y+Ncx3nRsZH6gHFeQOti/PSfiwQx
W+WW2FJAdoCMrDTkx5IDFgSYzMMRZdqzK3Il8WMt5zQOc7aMAYO6WnTbxw2G6bdzNuWeYFL7mY+2
PTt6DGB6vN2w/zWpEAXJjz11qMrIOrLnYu+kMpIKc4USzIk21+F//eCBumLXzZd+n9tQSRwT4n1I
s0pYOkrv5IULmSVyU5qVHmIfdKnlrCeUl/lYobgbly1TyhAaPBpKLwj5pbh2jcaD//GZeG3lbHTh
VZIvQhT7NNUujA2xsCw3OqlPhyRPpIlwuN6oIkUE9avbLbH4l/g/8yQVjQzu8Ih/myJ/UMQoACan
AtkaLmRkalSuuJhZTaduPb1gc1nUcI+oS8xp3sqntcri5Dyf6PX88QkYVZZetNCt8+sLF5Jc7Ip6
yavsNfj2bVdQbEfhnqhNVbes/oy2cbwRtoxf/SHmr9BXmRZcpBnsgF5yyfH+LnhJfR8XEW/5sGpB
vZoYvsqXIK9oBb4ZL0bVgxuW15PpxIK4hn7APaG1nrYLYenxeW+QsopzoU87v3uJj0N8YS5GspTF
vEOk8FEyKwu+61A9eChZmmEpmfQLeyFvsS5gFrWHXR/G0We3EdZJ3w12zoBYnsvqrjFIK6LINen5
wlaV9GIJZNQXG2HDwahMwauputkrcN7SGNIJAnlz1WZon7PW93KvNE+a8vpFEeZX6Gsk9sLsvzVB
rkDj5PKdy/5byDbGD8KPykn1K2b/U591Bn+x981PBF9Z3X55jr32fmRM9d4fmNG0TFu2I5EOWvdI
oyqNw8PdgwXwNALwF/f3naqYmeEigzyWGBgNi1SSx8ksb9jpNPPwzGKzJc2L0Lu8aZW0yOfHDHFR
A99ANI12NJuDML4Qzoy8jSCw6RfpDf4q8Q/1ShM+HJOSjRWqMhfDvrfPP208SO7BMkz649ny4LaY
4NLgxwY5go2MliV8i8Z8lqliorQt78TDtG2nVt3p+JOp9pBgCz+yi3HFhpwryv11klk06QuLruFE
2OVRKG16a0bnAyQA32yiZws3GKLkRh6tFlx2dsrpPQDca1YXgi5Uo7/tQJOxpiEFA/9C9EubDHbJ
PWOE0WqVJn/CNoYzxqSnIK6ek7ARQKz+LmEhSRgzco3TLRHJUZoPg07DEm/KvNalNjKXaQQ56hyn
abJhOMmcLioRK2kf7aSskALX1XpwA/6X0VfgeIGgY6atf6ey0YeJid73uUDyhzgqswcK3yRbjz/k
T3NT4L5GirF7cjXASzuhuGkoXcqILsnDhsmYYJ+pbkV3dxilKz4jwKlioTtu19aZy+Ybhn4RRJfO
rUkZjxAcVy/aaYOwUn9b+jmWTFlR37nxvjsah3eI6iNVD6sfp6JvibsCk3jKCZe2B5FYK1WRwNQN
1o8W8FJDbBdrmwI4pm/HDBoHoCza6Z7Gc1YLvGWScDsmEPJF6Vf00g0N4/uwpWugLCZ5QQclhD77
gxwZ4jr42VU+VsMlMRoKcZ8D3w/j/2+LufAFmOR+pmCeK2ftWjElkzxJqexz8qb53ROFAU2BwqDb
RQtjxlTegOWn/io09Roxt9MJx/ZreXF4OG+Co3yXnlBARg+FwCRuVFnt9OOnhVoQ7RE0oGDXw0mw
hcAmZSSI6plTdNnDuCM7PRabo53zLLajo8JgkLnt79m+GPQ57B+lTkrH/XVpr5I+NbEY2h2EUuoI
HzBloeegbGqNG/vMGVaZBGoZ8q2/q3yvJUDjXWMC2xnMw1BRCYEu0jXz7JIUEwhVGaS2sZQHH8RJ
4u408b6n7owQ7Z2r9xJejNCLlvt/buwRpZvLNoUJFE+jKFGkB57s4gvNS2qJ0wVXFrtbYe0G2B8Q
mf4u7432wvpyPlXWZh0VdXOtoxt5YcoaNjaYMZ2At+JAhm2OoztrlPbbYAaJL1ri+wQo2FzirP/q
YH5pTzeVNf0+8PTBwImPZyT5jqlHnAJhv4g9k4fJEm+EY9WcxooX4H9qj9pzfJ5+xtifg0r2BJpw
ltV/bliiZ0urbr3zZ8KOXZl87onBYCfcfFsQtLWJkwa/apVSbJkKcuyto7N3sURu7ANqMkhiXNZb
XaWYlQ4mYzNnUFp+CJU1BS4FxGZOo2jlb7TK0Nbdk3lsZyWMVGjCBTqimNKc/kD00PGwUfIgThXI
wStIQt17OMYEdpq+zhyjyH+RwkVMLE9Ap1eSdFXrwrVlTBHZGGBON3Oaa0iCjRw59qDJ53eMHcUy
4LOWxbClI02bXeY5bwp9hjV7Ufezzcoze9ygS1gtxEy8Wu3MeJiDoN8MrzynkkXj7uYZkg33r/mf
ydeLuj1Q1DPxsCKlFUn0CX2oBgm2/SZXOKcRY5bTr4t7N/dMaUot3KKUDWlsscA64vMlr4Hg6sCM
GKGk5iArjFeZszR1q6Z2m6NFZ2gBflT4kR/CJXtZVlLkgccvtC+ViXMtVvTJ5V4zyEYXOFVLYoHB
jXV3NQ/7iaH0UEHXoEiyBgjtTZXBD/lh+50E8E6f7JgIBgI36ZJjNRxXXgCbqJWm5Ex+0Foglvj/
ySB+pMbW0uihbzoTkZbXt4zDio1uYAdraYMbas6MUZlzylLniIG6JZLg5TIr21wYLg/sZL3p+qFA
OX7UIpYOR8edKEAqxqG1/isRjPyrGLc5LL2S5kCJB7TrExCdRuFtrcXCKuHg7Fp63xn7ORumV8ha
of0Lu57eodJCEBitfhwWX/HhAnzqx+nmjPIiF9HNwFrP6CaLDwIOUnuGJXXPbUqHZ2xjTs+TV+X8
SB8eFOYLF0Y0d1AwWXynsmrHNHrZcve9uBsKtBJCf2TDKpQI42pVjt9nLe6sR+bvuhK34m/S7QEF
PGsSxGZ4n/2/OXFNS+eeBTohtX0j2ngm4yfZCf/J5z847dEtoaxflk86ibxlNc47JNFQs5qXKEwf
i+yUd4atJ68+5DYXdT7jHInw+KTyn0pA0ygTkRBDqK8YDDG/nO90Wfe+Ad0EocOGWMIpOgOKZHoj
ptAjuVYO5fJB7XWV+wbHMYjOfh+907DUCnqDHUYLvh9Sm7DnqXksFMJSAjrCEvcvLFTFv27wrJfg
SytDSt9QMIDTTDLup15NRSPAxNcOG5tBQdMw/xIbd58J/SEWHtaDExc0/ZKTz+hGS6xpPLbnO6ob
bbRWj5AmBi94PvOVouYYQ7zn4ckBmpMWFnDzBKtB4fYFcIQ/li+6iGAsIZVOhcY8eYwKjy/KvwDC
bcVzZlgwSx5dS2DbeIUH+pGH7H2tzXIdZeoNjJB2pnMnkdGrWO0TSUgiIDJclFAG2OaBd8J0Q/Hb
FW7Gqyny/awO88ANZrOGa+C0XwaRVc/vD5vOI1hGuf/16Vj0XIjeFsgvS2bV9JCZKmTWMtl9wFe9
ytcGHej7pXjCVJkl/EyUgTs/wAZ6RarLNVlXd08U+PVuo5yRZchy0Sj17zS7tmp5NzEH3gZYj0ZY
tsdTc3RLle0JuoDjjRlhY9LczRMyXvMSdKuKkAMH1otPgiHbK29nhcOrKbUw9hNRX+ds2Gvypvkv
MPQWYgrQfUhgfEFbQGzwdtRL4pkvF1Juz/7/uY56HbqdZH67jcHqy8qvaN9mu0simZDVxCmxD04U
cD0B/jxpvw3Z3jwc9Jp685NyrQBEobM63LjVnwkPzUMnqq7wtIDTEz0/RWb9k4EzlWg0W4aR4FDR
a4t6n6IyIjgBv9nycYRvBE6XGnpZ+1nPQPEA2lI5K0OlXVPhRPJ5n3hjhq6qA9CtRhwPqDv497l4
sp2y1ksw4B/C826G4T3WlXJMc1zUM1n+3V52F/igd+zo1ZDtHfR8eKkUy4WNclPlUMe+7SMYC7HN
huPGzK1BMpuRegGdB0fBzwSnaWADx33f/0kMLmPq319M1nhohwDxONEoo/tWdl7WATp4eLRtSQWj
AojTer9ISh4Tw1kbl8Ury9sw25v26DR65/D5keR+7mFtHVVt8OChzRFs0Cj5or58H0veim91SGBV
0nb0ItuZ2xiTFZ9+5grXiXe9DNzdXC0VD1CGXx7a3zWgWLtYtAT0cVe8k4q4VL1xl6Kr8f4jlRF4
TFk7sO33N+Vo04uojc2UWPzwwZ8tPnIogRcvxw5ryZpl34bW3bLjHK7tkDBwibkdl7xkAvFWfDIh
kUm/rcsoi/lv5fDLQsrOQpM8+bQTvUbiSgnma2xujMFCYUY9/YKnDKKDlmABFH1fpbwRIOWXUUBX
AQYO35fBRhW5K+Dwwu6ZPgCZpX5/gxjYR6+qLMaJddgsZsYSj0C14Gby0f56I9lQQ3pBJy77VCjb
azTtkCKo3I5ey7+LuoynjcygWN3lsW/Hd9wf6cp3lKt1svF8Ie0ECrbfzLwIZtbwuGBPpAlQiEFr
CA0SpiJg+oWgRG120J+bNRDi4a7GIWlChD462h0WQRlqQro4f+ExDRUOfXhfR7AH/8qApqw2KoQo
NqFKcqvTlhD/l9GUTytj9kbNvuAlw0HNdZgEoOZX3YOuc6E2BkZ9sfy1zJJiqiqlZHlvFjLdIdXC
9wzp32kJ1vX8CGCP1k+iwU3amgAj2P8ACxMT9WHAlree6AdiLfM6p6jP733lJvmpbUBSW0D2npnB
9in0nJGFHLt9v/ojUJTLLIcDs5OxJFYLI2TUcl2XI7bzPNxRBKIq7KcCa1dpagkvwjQnXyzojMgk
tkDljSrZHpajLUX+/9X5mrwgi1YViMaalRUHs3W82zMSw68GhlLbkbCFcznavGagvjs+uqbuTbKa
qu19SYaY5S3AdEo42hVGWJfcN1BObRGzS0lANALEsSgfoZeY327UDMvLmceWEKbinwDNd/gVsyKF
oG+aw+JkG3LWH+NXnX4+4Z2i0IekSmvlMuGAvRqR9zS+zkRc59A19h9w21deKf4czMV4ZktNx/f8
5fVW36SWgx+up2SKxowaGkPBSEZ9HYqtdOxFY2PMXwTtSbv/RkHk57Hij7/pwEUBefGEkPXfTnER
1EydeH7p1Df8aeYLxIjC7g7Nwe92yXPKURO3qPE4G9tgESRXSjPMpPZ5QnRe/+cG7W/orZJisa+d
xn2iu3CwgSsqJXUSiNTK3Mfk+ba6/ZBb4ZWi4JXs+GWn5Ow3PuYZrc4AvNGJiPeCNiioUEfzIh9S
L/1Dy5DOMeU/PS5c6q72c5DM5KG7cHgInqpstai7uOuFZojSrLsX3HLNnSIvmrT5KKvRI9n5SX/e
k3pS8IOnvEAHtgDvBTpOy4TvaV91dVBAbDzDnBjMCuKs8Bpw4Hf75HDRVuAJPu1hI9jJbpDnJNuu
QXJPCDG0FZAHvRiRW57cxHzetAtdjpplXSAAQfC9fwsBx1oBzQqWGaugycd4ZWhsNSJYiZRWuDh9
B11LzhjXfg1V7DsRVuqHuX3dPkPu7ltFixTAhany+n+JfaMNMVdJGfOh7wOYSsmZUIasju+MxmOv
IMpwr66hAw1YEVJEmLtbWjnyn7IaxyweHbAr94BXT2Mock2o182iKjY16lTu3jTgkvYPQ/6Kz0Bt
dBgoBMA6/QGsBMKSJwLPaCCkFW35XXwzvBvodfZCKQtpCLpvggfMpDNlRK5AJZ9lQRzqdj9SYvis
qUYZ1xulbdhxZrabLnE2VaDESlaMTpfzKgO+0dAI9gk3a2nlnd1/EGQEDDjMD1Qi8a5V4CI3Bg5Q
6hqQe79d1CqguP3Xhhnq11PX/j5UxHCTQLoZFq3iMBSZE4pFQIOcO26comuje6hniOTloBKbvWD3
mBWbbRWyfmjHN/hwclobyBHSnAuvOaBcFA37W4KWoeJn3PVN5wd8alhEnKYofAYkgiG9vRUTYzSa
kz3bw6RWoeURpp894oonpJily0c7YxUCtgsD5IqET+A1TxCWM4nL3o0WJ+0i3h2GE1LcrD+YxTy4
8ETgHZfPt9NjNxmYjf32R/5UNAEswiZtsvGDe2mxkD/lXOdPng4hz0NreTgBFPzngVjxMyVgJD5S
k3vobywa0sgxEc7xuuNLmj5Zzow42V26eH+soOq+heuH6VSdolWi/MPYfytRwgzJFNK+TwDqgPlP
41j6Qd5X7YPsJJbQ1hTqelPe9qjONq8nvZqYfjtAOa+IcSgTZ+g2cnUPSDQ5hfFRZZ2NXaYfW3md
RJCQmI1ZsWRTnrTLfdQR24iCgjcKzzBfy5Cz0sqCoJflYidHMUFYcChSzQcJcNVEpiZfM5IwuVZ7
g1MoLU18G+8v3v1joGZBYFC2FyQx8YdE3az8Q9ey0prLrzwyg+1c2M+lWP/zFOpJJexq+tAUrGTe
aMz6SK7JG9NXxiFDSEivFCiEWZKr1aPNuv+sIbjPvSf3cyc41ME3iy6ndfVcZGxFd3AzN16f87Zu
rdvLrhrd3usJinc1ZmfygoTK1KD0Go7ruY+mOhoWetEQWgjNOqxRuk7HPCp3JhywKxsFlKfuLj30
hbj01kcH3D7S5TRI9YrSVlzlhp7/Xs8q8hHXcYhSfY4FO2X2ARnqJVh/KdkJaUcOECs3B+R79YZv
REZKRmWkKsMMRy9fPjJiAFP1FkZpu2jj19MCVgBRmlVqQ8jpJqLej+FinGwrtW51GjRoovMKoLFy
8MrwQdJ59nx6PliU0yJt+6tvSnybeVRD0y5BywnoSJYKKtQxJRAyYdEipGy9K6bCAbMpQjKoBACi
1hd7JM7yIh/pZb1my4G3o8GRKe/DVh0SDc5u9D7Uf5GwXBYXKPRRE0EINPaeMv3fEBj/8Mm6+EKG
q58FiJ0fQg0zyJ49wZxJqq6bGV2zD8faUqwbg154H8eTzqkQX8L1C8aCTGYuXyRAViqL6HYXb/6s
hw1F3plqb3BGTnCB5irarnQtqvqrzCXKN3OJfBhSiVpmMLGO9T6vRNDRdysNDWR/Vo1gZeJ1jlSK
snO/zIVCDXOzShyqjO4tAzFJs3WhWGeVDPGmBUEPoDw4evYjHL70KSIKPWRGRCV1O7332VUpuHQ2
ouUGFdTZFO9QKu6544WsIQtaYkCoXQY2INlYqGu4Eyo3LgqejIiz+w/isFGeiiRkbyd0vG88/DxJ
G6gPZ6KKfT8dMqNB9q2JoFXLsnYhHmSpw9AO4CtAnBS7xBVb+t+m8UJrLtTco/kRBzjVJwaxw2Fp
Ea7AFFXuo6JMrjZEt3pMNvLKDwu40goHKpA7iOQZH1JkmdRdizqUpLANdX8ryTcsITR5U9PyL7nI
9N8o4QnWQZaJMtZxereFG+DDUnZXEmekjCq3gWSiqNcDAWtxNotstKNQeZ1tRjP1l/FMWoXP7Kit
fA/kslkLg3kcTaFvOCEdiU0E6xEha/XaRiJZ/OrzjjKhKWB0nHYHaua6KqM8/T60kfmhOezIDbwO
q3aiNyMllGBToqnkXGt/fK2tq9wXMzl7LnNFt6ULJI7uLhhuGolSc2qc9VHZ4+d5FX4h1u5Dp1Y0
FhRxbpFphgWaoHkVSgICnPusbYbQzJtwyewR12JtSFIGdDcblxvFOyloACFEuDvmdcX3cDv+r5QR
g/nN81jrIgct37+P/i5V17qwPxUHWSPnXCMS6cKxO+wISt5JKCzi8hb+k4Ui3uKVFtdCFcq/a5cm
fQDVb9NYO1D/fronYJCqKm/rgtyNh6xRk43FEetH+qMKe7442zYIiM2J3GySCQfH6Q2a+NvI0ZwD
VsFe94naR/XB3NP2HQi9niJRT6qUDBamfRVtYJJFdQvoUUaBNz+UD5lP7pkFybL0S0D1nhDUGUSJ
VT+zM8oQksUdnkCbpkzg4dWhnJrUZ+2jkkxHc9fJth2bE1zi5IeHWU1yWRJs8Z4+tfnD8yVpao4a
JFpjXYbufQDLayvarik638tjqeb2ku8gyzdST4hwdBfXI4fDPE75Ec++B3Kt37WAbeChsTeS9kQn
DGmaTfGIRyQXClQMsNvDDXx+b6DXgzc6taG3VNG35U+98zLMgmeeZ7LJverZ/h/gT6pWOMv5Yt43
Ew5hXgteb62dEZbC+NX0DyxqO67qdAaAnD+OnAYvig55dJXgNAh92KUKEmGrO0UKK3GDKQJCEOSA
A3eczCcnsB/JWmZY1kXbH+pNuTtTwrJBCCfkXat2j5sx7euQhqXblZdZDwXRSvd+aW426XZ4c+uH
hlENUGl5D5753JIw03pvT+PhmirB8IY2StR+jiB2yvfOYZO8NdEY3/nz71vUVASMcB7MagzE+oRN
OAB+bQJi77utp276rMgcrXXE0IDr7PqUFJhBcCUuljK6r52KovdF45O24TsfeS6EzZMFAUxs3afF
4zRKmBOUu15b+f+atfc1Xq4UjJQ2UhMj7FColhHuHUk0urai1QLzx0nxnSkp/qjvBDUHEV4szDr1
8oe+mhHrOVnMXiRYPcGC56UScGsW315qL2DkKudD8z+OMTKDP6TnxGk1if3YKRqRUgbNZFdcI3Mx
xA4EGY/k0nEHVtfA99mhXlfUincGi8AbkDpSkHYngEJiE7BGSUa5jIyXl3kV6sULgdXgIxAf+Qyc
BQlzWabvQBvFdS9x1aVj4HxBfBxDiF20fTUuZdMHnVS+ff13LJBMgYtQactQpl1VE2KaG/6m3PAb
oyEX4d3ihSePQEGHLIsLm/nQ6zsyjn2IMYRtvbY+nDUB5Cfpw7BDMbNjsdEuUE32qGcO7mKV+VwK
QzrxyGAhr5+LgGRU+acXKJkAWhcMS/92XINiVK6R0kW8Mtu9ZRkxEs/F7tIFRwa7ResDrr+eTbx+
tlsmD1K1T3feXz5Ene3EnWiVE87WIFJe567ZTse95Kx3gngCAjqwskWcx6+6iEhP+zUzK1YbQyDW
KVebyKVSl0LF9A942+JeoUxlu+TPXSZ5Dh5nZ7R4nKcUQeyFMW0zOoQELfSQecByoZlwKs9LagFh
kog2IEgQamPTMP4liZsoAxSsfs5lLNdkW2KzjFCJIUUtcx2hVh105VkiPuBJ0NT+zzR67P8gExnZ
FT2+T87xFVaoyA8iAswRTzPNY4mvRGUJPxOWDUpS60lPl+AWeftFuWvWlJNfrKaQN1jcOQduU412
RSHrq2n8XHf3QppBZO5HdAjwKBj1JfAbyix3RECRUVXD53/B1bYlmdvZjKbmjE77h2aJQKreQqum
/XkoLjfTIJEqeQi4OLFIaEyHcabEXWWa1BWfY+3NdYZllL7uHusXdAm+5gkpJEmgImCvO/O0VMIO
vW7OMMO+xl5GNIjPe9QW+gn5c/pFAUINkG6xXK5RNjzTWRTpRJW0EJXmopFcvyicF4RPa5nlFE3Q
EXvZ5fy4wlww7I76T0Oafnycs7FxlpCY2uBPdLO5mg+gc1Co8+Ch/Atwq9bDzLKhFYkfl+EE5r01
M/KvvJERjCq9EFrHhPJLpqDyTSH3NuAdFvi96fIlN4cKczqyTng/2Gs6RNf3QSN/orkF9ra9dM2o
bc39x40Tvrm6an27RNPf6L6CjNQ2zzAjEpoRMyYru55xeTx1kkhSC5clg9Gy5n+t2f6F7aWT5LL/
1TzUUEwq7O2J0MaOKyRPpuIjmqYE72/OywkUa+/dhWQbKj4wnjo8c2l1GqQ7udzqYvvvdjbksthy
ErLqEuYuWhMFPNQppMxDDibAej1NA9W4T5dz52jWWQQJHdnTOUtmSLuF0zGGl0ImqsGTOrYoIZvI
4A/ZZlyYbL9Odx/TtaH/UFJHhbRXkM2ydEOCY98gOTpLB2hssFILTmkxiNogUl2i1zin2l601xp4
DZBsEA48mjcJ0M87KENTyP4Va647Z/Q+1JWX16h0zw7Ju3ZZSveNpLbMmmJ3WKIYgFobfttyARtw
x1wwpDQeSXfx+Rk8v65CvVs5DqReU7aWR3BpM3Q+bFc0s6gW6yhBZJnpKIRRcxntZSjx6g218FTF
A4F7xZ+lwQfLDUogBGNZR3kFS2Ar398n0jN4+jfDelo/KClzx+VUTmMf/Zn1uPkkn84XJ5slYqKg
vv3Qntc8Oa9X1JzNh7VWZlM8ZncodqOqQHB+g/NJ8IgKqT29kyIanmJVzsx+uSUtpbn2NNGg3v2H
sWFg4M3ak5ldh1cn4PM+NPxLl88K1qcITFCT2B9kUVU+wjTijd8KSZedZ77Q3ZUZAMgq/YXdv4Ea
0xe5FB0EGZOC/0Ug4Z9+Vw2tOCV4v1sBPvWFpMplnwN5xtOd+VQFPz5zxAW98zzGmW771BjLOQgx
7z98gpkbayoZevb8BY0u7BW+zsCAIKaGeaFqb88tm9oIk35xeScNjXLotlNUg3EDkDtgeU0+iENd
3EoQab4qmocN6g/MA6UlZEL8sXdKSNbGZr9WrWUitzJChZvF3m1fRC+HTUBH0Dgmfh/ubGFoIsnc
D+oMTvYIHz4RjfeZxDyG7tFyaVDvGsgQ7laDrZtqRHIcIkwalZY9fFpap703kWpkFIrjmCJCdKcV
+pN4W3IpuyYxFieDjkYpw+vwUsOZbzkPLcIXx9hkGBZWrKjNz8bIOuJ+BHZXd/JJVGNR7WW6mlSb
KjVYYDegHdPw+6sfCKsnrfNZ9jD4QNtX4vB4XydXOpwSp0MczfzPUCXzrscEeFhOsrXtIX9QuXqd
CGgH+ONxCEfBiXtHH5zzpPEZqbk3vncviRZH12MK23xLKJS/eVktFxHEXVAvZlePHqj1ACBM3jWx
9d41Jq4hGGKvaocp7So1YwMzfEgao3QWrXDAgy93bR6T9sPsnbHVfOYkC7D7S7eEotbOVdSOmqYX
TQMKFMm22JVGPtj4dg9lcW/2GnwX0lkf+rPxK0IlxgCWvcYoVJwB3wOMfsCQLj46Ispd6R+99pAv
x6jZtn3CN8tLFJHbRQgDTY4Xc7TlmpJR3nbIPQwWOjPRU1yGr/MKQXlfYoHik6dS0Vh9J3RDak7h
p0CvTCwd+/4Xsc4YUqqYAB70gpsOTdc9qDPL65LdyhONqOAGBptSbObkAfBQkQ2e3zJR3PVaNtv2
n3voIFpO1mwS1K450uRqq3FBRt63J2ulX/jJ9vntvliAOGtQ+Rro02mcR6iKC2f4zwEJF+4vuEC1
AkDewiPdHxP7pbXw5dpebo/oZcEPtouANpOrRLwh22lcflZHPC7mNrlC7BniA1wTcOnsvj5Pl4Bz
MqtzKBqn6bM7vSOkiV3zAKyMcYW1r/oKZ5TOj4CjJGNsFOhqJbGaDsYwxTp2CWYxLohTn3jf2v67
rMj6UwLVX7sbMnmRiF+LOL9PvVJ513A8f5dxBteXvNqFA/860cS2qLrJVHFRUAZnNPmF1ZkTblRg
+AtYCXWm/srHQNT7JjjnQx0+avMxwNTb98DMYGJy+w+5mA6k7UvFROs5V5dBhea5Ukljz9E0q4OH
8KV/9B10IcQCk/+AzfVtQzTLT5WlMTFJhDm7J+U1UWOG8k3Wnm5oAh8Qux5zV16FzBh6uEOGozQe
ZiJIngq/KD5KZS6mSqRFdNN2dP7NZdqlfEW/w72LeQscjzynRCgBTDeVIQHotTzrd9l3DnE6XOfa
EBYXswpMQJZ8N4jHXxgg2gL1PH3WpUXg/zBdMyRvGomh8Yy+jkXtS8UIvVJ7XA8ccZm7re8ACle5
ivd8gSeNhEHEr4SayX7ahrNPV6TbZWhetwOnttFnlSBAjwS3GUUpi/9OsHFGLPfhwUFsNuTO3Lu4
vqeWNDp0wUiGcg7IlWYEHMA0E1VCKwuDQsRVf7smbPF49wIVfOcQAw4F4/rqOkZzt1hotaSIeNlm
aUNIk/sa6VLnVBDR1NJZZ8uQDFE8IgaTDIXuhRPj8xO9CkNYWxUho5zBLv914tobrjOBx4SvqBAD
IldOFHXKG/4sKjTFXtVZLvVY64sLxhT8iBDROeX31SKGCrvl2d2Qaqibf1OBDGWnyBefr/5zInJY
0UEvEnzhj4Kg0IFp35axSWuK/MHLaL+pN+LxPIim8xQE9Gj1bPzpRr6dTjJk53jBxlPRwC7bnjEv
Q6ehKtVQkoNi6lfInU38uZ9osMk7He9kwa/mVs0oKB9Xv9KdTQvGRG5WF8HbUSlv3SIJ7Vl8am5Z
mcTSju8wH5xIdO/iAaj9GOwRXUNu3YI06lmpLC9m1KEo9RICimUfDMs1ukJtTkiMqYJxObDiCeEE
/oshBDtDqoW05ggN8fk6K6K2r5QDaeFuPVjL4z/dACeprAPJURAAM5WOlezTr7rLib+c+9ZBcugu
CpoTx77PunjM8NxQmRZG6hpyaj5NvtOqI7IdNFc3OX2TBZVkRtYsTlXmwgmHMFLvARFNLYHkziFU
Q9YyoD7xztX6btKO6Mx9WD+j7fbfyEL2Ocn64wxm3WiRbWaC4064bD74ct0eVdYKoSPp/akjE68A
KV05BduD9AS0dsWUqmD382ejGKNU1hmEPWnvYjT8ewINkxdPZnswySWzjlviHiGfHhRf5UUdUTPE
YZMd5S1YpSDPFDrkyLQbxS5DXvSqqVZ7RCACO0aSmpj2jXu5t2V2z0wwehP0sNKEKx6AB3xX5cJG
Umn/yHdxo9vWkq8ookvrS1NS0VUaj36JzRQi6Q//bohKenN8XWZL3Exi4luyIzhyPXTtufERN5mH
W1tw6oGtb7zAJt8xYcqMgB1JGlRxfol/GFaBSrqBI80k5NhDCpHLnyaoGGq2PS8fj6gNCK4n56Nc
G4kMk8Eu9psDOfNuCPMMj1zqswzmzTbzMd9wIXlQ+9z4nY2qA3OaerXMC43lOksCWn0jMtJrbKFf
zNEsbgEFCUMx9BJ5Lwzoam3JLqFw09gKdONxPRCctwKrjRZony6PJPabB/ErxtEPI7iHhKM4JRQR
pJ9H7Oadps/8Mwwqg6fhyuV0ILi/ymxGZWLhky2OIpTptSkenU4ZYAs0M3WWtvIoaeCrXEmzsX/X
A2e1YatiJbDCGDwRZom2QCGtaTRNLDSj2PDZ4AJoWT5/OKPjxDroWW3ptFOiv6OANUtBX0uJOjTa
WEisSrEIagFsBaFIU/zVmTJTG2YavBuaUP8FNMuHTwB5UTj/ftAV62Bi2vlItb9PgJHK0lF5L4tC
fnwxK6FUQcTYaKv3kSsAoVY2uIIrnO0wB7gm1ftwQokG0E+tILdoVw11ZhbJ4j79/Q55AEFeTjEQ
y3S0y3o54P1mHASY/PJb/Ei5T1IEsnAnh6QufiH4qnNYUZprWLA5JcXhGX4W4VYiZlmXNYoLUk5e
jMHrLCbF/6Nch8+CwapSByB2QP/fEbt+nL5cJnPV7+RwFsfPkskOw2tar0/iyq3avtwp/7FNo+Up
3PbxiOyH7O98qTXy4PQz3bBwxClkSWke4BP8WIZUf2gnh31NZAvie5EuLVzC3b0w6TbC7ZOeg2Dq
8kgT/56oPJDOvXhRyVjYaRP7o0Czb0F7jPE3cuAdrxKaodDQL1qewmM1Z7G7kYHWL6MrS9wWolge
CLFTp+MM5rbs7egK9tEnFgXwQPNf66bhs0hbljzSrF9XDIfSEIumSQadFYFYQosrfNd1IMpXIFXn
YnG6yjT2YYKWKmGbtquj6t19o38pE8dtz2spPAk4qqdwW3evEjgDVI5dMk586CYMGIBR90sFhdnR
CdXHGU89Iacf3z/ftLz5cZdVKKx3Lu/o5smpqtWn/+EMv5o2H9cUzah3JYA4SqAc/yV/ouqJy+O8
FuTeCYsiXQ8d9Dw5XLcC4LAh8KSUvb9PkZKvOEd3czUQvBDallNXij9vDXZ54Ste7IO7CXhXya+1
jKP9JeAWViJ+Z18utyXs97a0Jad2elxfLPLOJ0oFWTjvOo3GLx6BExe5T6XeJnQDrFwpsbBdewMw
bIEzfc963ZNciCcRpB8owSLZr95SkZq8eWKIWNHqI0DT4xHuErqCpA/fw9gcbh4XyNtINkEKvxx/
I63lmo5SwWpta09XZ06f1stBEU4h/Y8+9Pzri+RayJbZQqDdEj6NCz2Tlbhzou2LCyq1MtHKN8g3
i4INR1K2J/kX/Atee5+ftRUAy4WYB8eCaXs/RycKgeUbtZIINZ0uGE4QdMSfl/n4C4x29Kfax1Cr
impNd5iyA8Dja3uqqb8Z2mmKRu9mpELC2N8WhF2JdbdlxU6IQDp96prKPTvYkRF/E8J+w79/OGsg
i3NwqBEzYeIBcbhWi4UrvrTib2GJCvaXjvk6btdM/aVOY3GYSQa7KWFVFseJAF7t/YOfpI5zbYWN
NAV+03/n00J2HtLOaNMFpyE8S0nY/hxgN8h7+oGkYetuFehi1GEhJoSAd/NX5Isv1f6rEhayEDZ8
U3ppJsf/es74NWKvZMztUztqPpKifC91RRUL4A57W9M2b+8QlPf1N9dwNQQbS/4s2QJzF+TknFbr
uOy90NIUqRdJwmKEeA3H8l7QqGnT2VIngUdZ0LzyQyJq0kX/w1j24gDpZD8hBV5jjPuzH3IURSmi
xnJQkNoN2mAvabWECf4ek2ps9LbuRMpyQnZCc1U0VCRWTrEjbabrEf+oqJvdO7YbhrokHNrmCigD
lM2dl9gsRaIbcLvKe93TP/PMd9af+lNBSlx+9RpEJvBIHtAsLk0O2p27/a8GOJVLaZoMR4ZphBRq
Iq2XQudpb+C+J7+KtcyVGKBzZhZo+koA6+NSX6t3XihrHuNj9FnvVL+I/P/FS2REhAawLHhRuhss
MWKrsSOzxmpZf/C2W+jpiDmlfQ1ZrmXOr7LV8ZRNxCetrXxRUksIVOxROneBaasYuwtI4uCMT+HT
uOiwfD7Y/R0ikmlL1twP7wtmy3YazjRoCJzHDm26MBsqpekaKXJC0aN8+CKRvaqADL4vsIq4Hle2
/W47k1d3IZIjr+yrjX4m3/JXMsrIJW7Z4GRiLpBk5u3/IiqQKYy7MAIYkvaMbsh3XX+8CnokkKbX
RotRMay7fijoWKBOcAmbtD9dJ+OwI32XdvTGHd1JYluhR1w+5mI1FCG1JK4xXfbXh9o6HFCT6Aq6
VToiqRhWxF1dJQ34Udn9UKr4nUpfbn4gQUOKV6033u0ZAiM8UaQc375g1v9hjFe+yWoGOqbDwLLj
u4/jONDTKOPU5PvOc+0rEG0ZXdSLDYWgOHA8XSnixGjxmNUCPdR/gVBdPbm561ngpfgocT92flDj
QwMkpFglzQQQkSt7pBxbYGuUD+h0P7XLLq1lM7PE2L0nxaZhfjpc8ijdWapZ5a/Z3MaiS1ETIgpa
VfnXFCDijL7nr33vXmNBMTnVsmMAhVY0yb5Bw+F59yjJbA9dcxmBvsbBsvcGNMRfSVYFPEKBrE6/
HDaVukyv5nORUh6UiAwefQnZPFqRseI5m0w/ItY1lucSu8ZXVQxUSYNHUwEWYb0lr+xAYFppaUKS
7zrd06jwP5wCd94XFqsilj7KeKY/d1UEw8bFxBmRIXExP95nxVidKRx1BxMUgmktFlL7ASL/6aAW
LCshmaMhSktYK+wmHEkcC1fTNdEq7F4qd0mLxjv+fqAxVTiB6hCuVaGUb9eQ0qs4XenY3t55TfIm
pWeyUA0/mG7pE+50XtYTYaknc5n+bFtNCPxVsT5s9Qf2VRLnxBdlw2PxvW+4Dmdat7ZJbnXhVH8Y
2RhOARDYDBfojZNY2joMeAxVxlUsCMR7GX4Fbr1Sbk0fhlXX4Lp9wMBCwB0QQ4flQGPjoewnMmb1
BIoShyXJEqqoVvebCnlbLngJpMGxYwhxaiq3/BjZzMBzUIJfLptfOg1qDiaV7V+VDw34wpzERvhp
zodU4xMya0j5PO85tO9TpfxK/cNxmRqogrnw1XWqH1JrjkIfkonAjovrTKZ6Ttzve50DFn9RjmbQ
MoM3Gdix3YxJisL9QW3OgzcyYzuXMtJE3Hg1mDkVcuAMA11/EXu3zCufz3jRYNS8UaGwY66T4wPE
mykDLRRGYgfDhBPLGaAU1tBHWQzsmPndxBk1A50NgPn+bpTUIj70NnkcQHctHuxaDi/t33PGxnQ0
ipmOf44yahfftE3cHnL9AEISjsPeXE4phKzCQFgDnIRHDVTiRSHLVKqxbUQARd8gGGiT//IAh/ip
jC++HTVRWIurSP1WXKiAmhNvdACi56+ENdLvEMEk52BsWOE5qiuXeg72AKuLhugboLq24x4bCQGe
R67a9bIqPF1ha9yNu7aqxIlkbLAikXZ6qbr0u+gv6oY/A5jECAyxMEvEryQ2hGi5T41Zz0hpCDGF
QZpjDMH0cH7/h7zhqB0dOckDft6RZm8HsJ58rmS7S3Nv0A9rlfjSF0NKR7LpAD+YlmdWyFF4mTyz
Dbg/3r80lf5dZmIzCGBsrDt9p46Cr61YhVHhaI12RjBXjEjVjZP7505fwcsOHNClHwDsRiHHrgJX
j8kMfVI60gt+5gMi+bjCn2tyHzFEy7DP5tlrof23+WV92VGoTM3sW1h7q7GDufBT6vuEu9UNdclH
Gl4HgjpmhecvYzj3h6jVtwIzNGwtP45Rn4nF/OxLB4IhfBgf3k1TdTHaFIp9Js7wA0TyRV4bXns/
PXl7+gF3MJp63YV9bv3MxaAG1gekX556nXm0Akiz1g95qRutK68jXEGNnERXpORD5meGMylCjNx1
IlgO1CGGpDIHg1hAwzZHopaCu+eg3f++z2wP7hi6i9RKpGFKX4fQj+j4qQVPV+ukl2kCnJhzQG3T
0DH4D13Wbm6x+Qj/0StZAbVZMIEN0h/ul6NO2Ux6m1catu987gjhPaOg8qF/3O75fi1kzcLyGKfB
/RIc4Sf7ukzUfrcH5NPqHcx8omoo/MFmL8uT+UK7y5ERm6+0mxWfoWvVMYFDuytM+ahpGTn/1heA
6J3hmv7gjSBnlzEUjnDbL2ElqQ8+PzYmxRTREYDZihLUkT/WTXnDLvJ7IAM5+vjNKjpP8oRSyCaN
5JHt1bHLcu9JyMQ8s2Ij8Sl9A5GBqnqLgS37JqMC0UT9KR2tdbKDH1W/BZFjvSrDAOu2hTcYePfo
+eex4eqzXrM+3Yody+gDbTTl4LaDx1TeBFCDvJw4jIUf4noby7YnLlcskoE2Rf8eMSWDW3LGDwsy
VmBlts5nCbq3As0Alth2IhPzidBxEetAn9nJgxGHLfLr6LW4lHSLOGclG6LNo/lDwWNDdckzh4Kd
MuRUNpd9qlmxTKd/Pn+Q1/XT5fjJRVCVQTnqvq+RybnOnRd2dPl5nPF6De6oxGuNFb6RNIFWrrw6
SHltx9FrOo73r39pmI8nFMRwcEKouwLTo/Bi3zUPjnZq9uSXbJUAghmsEMKsKbkf3pp1OdfVGyye
eOklI8LsPn3vVxpAEg5yz8ZCARNc+vZXamvywQXLrxxPqKrXXhvHdeVhSPZDMOjoTZ8/52iY67GU
1R6eBHYAdLPF8YoN25WQkeLolYElWSc3gY1wXmTggqFZ6PQK1+A1JnVsSN7eIpXC3mep+dcKFR3w
onhriQG2u/dTMKXzY2S2b6Kb3eSRlNs2RqwqjhUQqS+a8h9Ll1+QzBI2Ilwf/ChF73kiWmDlr/vu
4rbPGOUNuyqJMY8YUHxvppZgwUaxeKw99vKSlZii/rTxXnoGPUmY3lFr4XHEz0HCPXdLBUsX962M
dZwo7mAON36Mz93Zca5PioAHEO0AlytRoSAVmLgyxJFooF1LkYpt/zuCSHzPd0MLw6WLsKqTiBNf
8qdyuuaKGNUbztisjZ7sgYFZhhk9vZnWYksqRY1JSXLheKk6zCykiD2wMXQNSLlQYTCrAeTOEUuH
QFFwZiAY/UrowmrQf3SJPcmfCF5QHxTMzTzyEnoa3ehapyKO5C5W/8Iun7UtT9gyt2YsiVixe32d
mmNDcqVEvSjhQx3/doxqqR6gu8ocLNX4G1NLPfhw7fzW4rZm32xXvAq3ndyPny5LHYQxZdS3cvAq
PlkkWI8PwwmMUJoTesVxLRJ0Lxg3cmDKlkCJBNfwPZBKshWnRNqHsuV66eqOHzaRA94YEKRAsM+H
Y9lQUVDkdB4VHBf+ig2O84dN87A4kFQ/Cmw9Rs5iin/oiX6UHrfVTWu/f0dLJvBa+mTlflV7xTpj
2cvSeT/Qzw6bpgz5v/+56gFz4nzj66f6t/FKze44L3J6MfpNBrhH1DAGqsswljjjHciR7nUI/oEx
WLyrR9mQoThA+JmH+9kkwLNWcrCfjnEltAqOz0VlPDEGp9oQlSw3hRv760Qfwb4NGqXNkY0NcMnL
j2n9jhCD76m0F3R9T/4+eS2D55O0adXynnhYhvH3fCEM037QVm9opmXJfFY5TzKaZ8LAlh8fHbkt
O2sMLevsb+os+OMAAWYpaQ4OAS9NNcuR18laU+97ggBHCoNcRxBaFugPXiWcJJEmi2LiJ9hgIaDN
BK5aV+M+c8ozYrbg2H9klssSgrOnlqZFGM6NrTc4zV7Bwv3fRBTL81LLDxCe1T9zA2RT8/yfOs5r
IxTJhhAPSvWTGCJXLSRCY/o+sreozTHaX6ce6CJ9ufSGfcatD7ru7rT6VavWQ0CZRqwT/WmAH2pi
7wefOmRvNk9KoOlfJwoWuvEOn5hd9lxpTmmLayVfd19FmWf9Qc/hHAhvajxYIsXYPizFqVKveAvy
0r866lIHl+O6f4U4shqm6yzMMV5ICcbqiTQgyU42D8FR/zW05PGG4hLXQ5qMgpGrxINJDTGI6lyK
igb+dOP7jMo18fpHZPlaCX/abHiRf2H0+FBhONRUbp7AskRL1AetoMU7uJIEwgjlBbLs9ZGjJKjz
MLy37EuXRL5fhT0c6LYcVBQc/VvUFGQupMkaoe9C30fxcK/B50wRa2Nwb7nIJz1X9yAbhDQfymqq
v/YH3KL/Xv7Qv7+EL2PonMY75J1ASE9TrMCNRb50MXyNQIoEDojfPKg0X4yUcBzQ9EKE89dw1kl7
PiAaWXNMBGhC6Ab2N22kVEvfr2nAPykKYPBDm3GqBkG9PnJ+X0lnZ4pqDbtb4aT/1VFB7hIqhyWP
pWuJKcqemNh6G55bJPn5LPtFYVC4dio/aanaxiH1SZOuYu4G8auhohUNdvwNxmvXsqnoklkUg7zG
4u6IIJvIZ2KuEG7/iSB/U+5CZqadEy6js9RHdPazDhyZ19PB1xiz6LJkF+QRAEeHokcBgBWk9/eO
G86wVhyvpLX0WwS0JZyhnL2Lwc26IIVfuzGlSjxeGmkKj4vJBjimcaMOeqNnSNWPmp2c9NFAJAsP
eZA7tpKEms31J3642IkCubSVZznZGOyWgCeCZWPH5acNwhkcnlowkaRUZoVkEZTOFsyOYpFw+7mB
aRmdMJZ9MtDge+k9Gs8ciRkAocyS3TFAZye5sd/MSjAXeMDIySHVBpgViYIPDeD9F9p988KIeoyV
TYVX7p4jWc5hOA0XXvLbVUUWSV3d5XhLJWXGynTN2Aia+ZT1tpaGprlke7W4044E3UpYlkEhFZWn
gjx4WGbe+lytGdoerfSvNHIg0gvX02VJni7ffBe2r6fhedafI2Uvqms9NM5fga+HBXu3OHu71yZJ
g3Q+JnE01RVI4EqbQQk2rIyD7FUa8h7Bk4mvbiXYqlC6jRjPcEYWsBBB4n8KrCgZIF0HVbiSViVy
1Cpk/gtzqqemtVCIYpZbJkAJicl1RFPyqzq7lpWl6WVZGV8EdmnmmEv0vAl5gLfVOkvfQ2KfpTiA
r+q4Gx+gZ3mhH/ZrJJHKk/cyZ1AYLn0vq4rjQomHQjKeC0S3CWtEKKSk+n1luBIsfhw537kZM7i/
9loCr29dg569lnvhypsfRxZtMsEG9lCGYZ5NNtfpl12FD8nvLiOYV9NduMKI1ErbgpEY4lPRGenX
jHZ5/dJu6zmuzBLbH0/o7m/PAibJWT6siV4KKCwqgiIBa0MX9rm3geHoeN0coWq1zytLMPMsmMCe
tG5AGLbzw1NCTkv7DhppLv61CHFkQSE4okO4gapXZevYusovea7NnSSv8uuHfY2tvj19lbE4iZJd
Qu+DPF6iauiQwWJmwt2AIeKFSN2DdRwvwGFbNNjP41LIKoOTWejkOgQXbalk1/JW4m1wx4bnptrL
8DzAvA2OfO72uDTVNjQaZ2gJ27vziBGO5NQrUBFeYY55KsbTjIt8Za8tIzxc+Ss18X6ZXdE9382G
hD93pBtm7h4ttBiveA4IUctM4+KdBXvaoNNiFRNbtotFsHDW6GvU/nfxMsCEUZO4iHaVUKx8hIy+
6c2PILp5wtk1b4Whk9N2/Lmrh/SMjUA8ZEfVn/L7d6B7BJHBzY0SBLcGJLsoYHpbTISd+LvOHC/n
CAUiKEaZKJJfn/JzUxheT/uWkEb4zWdmGyUFpy7Q6NNYH2ROTzXSkuFUkayLbnK63aS5Yv8AZTVb
fwVWHdGDX7QcAeukmFKK52KvTlfuys/iGIMw11K8wym+of5J/Ac99q8Iy/n2XcYGBEhAr3GsvoW+
Eu1mr6FmshaTw9kH+McKc98RoponEH/OeZzSW7bgPu1D3wX2FCAbKPRHdK3TkkCNEG/uSyBTikIY
WnUgNfJii0AJPN8ib/V0u6YlopHPxfHeYnt4T5UcfQi7dPpUSJOH4yZuqehiBgJEBRjWiTeA7og2
JODyrlsQ0tpPQtMdp6+3oW5S3feUzhAp+m25PseI9TiVbffMHBFeELPTzL/Y0Ozq9NqOYXwHR5Ks
55DCHvdbqoD25I7oolXhBIy+z4uVEf9XFIRncXhTMO7VlqM4K9F8RLIgzotJe6gbADPtv1DslZ+D
eUDRA2wXXmSLeWNZX63OoFoUC6g9WXOlJiOZO+iIhnz8d/lMSl5a8tclXnwGrmw2t4jVYtoAOdPl
kMG8+t43xui7WfGTXbKLmID81YbqUMQQNUnTPkTE6Srlw9QCbzkamsaOHl2w+HKLw/bUJ67Nyu6o
yaRzENDag4L7m54ngvEmtLdNmIBg4Y6m+Czk+mn4+s0xnvayu+N8K1KWR5F47YKZMqyrRYbuaJYm
hm/iYpQzn4QLOkqtVNDGa42gieJ/FUHLdu7EjMrKzySXiLT4nIIIaZJj+o6qdpbdCgDDohu7TiHz
LwkuXjwN2F8Vd3Ioe/0jKp3FYVhliHZPast6wIDKf96/M1iXWTo5lgyBUUlgy/p9dYSus4eCjORM
EC4WdubXZwOUluNZiwHdE7ih+Zg6Y28TXlBbUstSPOSG9HcQVtZuxSJtceIwG9640cikxOqyRfHK
7kX9VBI4uk0U1XiC02CPAgApx19sHbxt8GyIW92Qs7s0DuNwxnaolJJWphLPhPblS86y5apLqLpW
X77UfnwFluNmrJHBpUpNXA09NWFta3xNtbayw9keiAhDOcRC18Nj+K1Flg8/9RTOJfQ+H7Lz+C4M
uDgSa246f/ChgYBvI8hyDSBVCU7nT9XTndEFgo4uUzIvnotGfMy/FKrESUPezNpikhgKNPZBfC/u
cALpE7mS7MqtLSZmjWEUFBUBo+qL0ScLsdR7MwWRlPhF3kv9yUpe1tiXqvIyH8GdxlVv/eqaMtRX
QbzQI8yK0I9ajlBWDC9yWBT+i88MTvPUybDyXF28XLae7QfTvugSUAJkU2JWoYT29+nVYvkZCXmn
Tvc9tYpWgDl1XCPEWJthE8adv2Q59vu3qhprECHMYDSqoXx/0ohKUYOcxHe7lblw5iaodX1HdtOo
BwsECSlSZAGGivB2o2/Y6tvAVEaYj+M7OqkRTWLMEeymZZ1jxEt5Gwo8A/gQTrJK+BNj1d/wY2KJ
UO/AuU9p0l5X5AcT4ShuodXchkfcvNwFPw6E4r0q1ylxxzc1iKlFmVHsM8VcQ8mcLCNLLHYpzkps
5qjIN6OXm7NXUwYRgbTeX49/NODALbUjkCyU2IbXhF0LUaN1TugS1CD3xLsy9K4gsaZ0dwMUx8Ge
FKmX1XOkVt+yrs/Li6HlhOA+9S9lqB+I/t0JW5aUyUGck7krNpJ5NBZlmY6qv0uczM6ED+tst7VZ
Ozo4L0WSYm3dkPy1tlcjbyRQZZakflb1U3nHInh5oF4qF9rWX/uxArMCYBYOJjbJrZhDyA4GkQvu
pBWhiCldt+HddzSudQDX55vzcnxH0gq6idyZrzhLNjZlCOeY2FHi2D4BP0cVEEbs76omzoX1TKjZ
jLPcV5/3rcnp+NGSVhaKp9me4y01ylcDEn2mnx0buBwUWrKaDroDj7cg9z9QDgnwmUd5jSYg8Y7Y
9avNxFd4cm+sL6w91PURrQzMyiRuQ8oTbmSLTvW4Kelj59NiodrSYCbpdYgZSNPdVqBKqVRF1rRR
D8uNbZlxGiAoFIkMibwnHFZlmmVfrTVOk1EwuAxCP5GTZjYYaNcdlNTf8jQZnOOThx/Z3iQBVP+x
MYabj5IKyvxYNL1yZcqir14xbqWY62TW0TB3aUfE5GMrUTtywmxcXnxMpameBPyxARFdCum3N/eh
f7LqeC0H+/nAigoEmMjqf9nPP6/G98/3Md+Z5Ji7ExIoDwqkyhvhXJe9uidgVCrml1Zp0WpfSvfD
jTnE7CRB4u+luhckwXAHrlUPKhAV7ztVs+7T/8PibnLionC0HAGQfJunXSZ2OVRTQMLFIIccdKjP
7zbsFZ75JfrkVWtX9EnehkFnlhgK0HsDiDEQfW+shAFSXtI4gGVlBNV+TwX3IeMZcmLtyThf/XMy
kDTwtHl3k48/k7sTOilQMwgsUV57+Q1B+Gf2QHAlx1skVw3Gx3TNwKaU60SylAAIlWQ08Lvd0bb5
0fhEJ1GF9dzcO9iJ4OIAImmuOvK28LSBTFOYqmujrOTRjTA/HzK34/xMvHl55F6Hnm3vqYxCDvrN
XHUb3o9oCT+wZ965s1gAC2JxIu2rEpAUVVzcJo+5EQbuqDQ6vnQHKuXPEKPymgDXRaslNZIBv1+G
ISU2vAwlECmoK7M9FqDwAXBJX6B0Pg6MbFJ2Jlv+kXQyyOUQA+/HMj6HaA5BqUF8w5ZCaIWcayYK
4JoO+UNvID9gnu4gisEGFAiJB9w7xtC/HvOTzwLe3JKfkn4WQTBhV4389ZY2qahPd2w26pDMcsC3
jiIiUzMwQByQXj46HHD4Oa3IXBhg4GTm1Hah4ocNH0h9tMDXM3RGIxGlAdqRE1OMa1nPteDYvTHC
N7n0Bc/AHbfUlBP3xPds+ai+uekakXB4+hyNRQObBM57pHEitE/NHrr0Ct5ysKCc+hF7UIgz8kfm
aFZFRZvdw2Fw3yzAXjBsnkPP7NRjL60Mdd1AoGIb23XW479e2F6vKeN5GncGXLpPyb4L2mxiprRZ
g10xDXFFB0TWkCCk1HV3TsHyNu944BELL3daHwiQpsIPd+q0aS85xphTa/dDyJubYHU4myAmaD0x
csDo9yUp19Xj/hA+T/1pxNH1hAHNvVgP7/OMSrv2PWrcF2sOqFvkokXSlHQ0dBfjxBTJDlLYzP6+
pdHZ6uFEtZk6lCgZ+lxuj2ezuLbFRnOYnrdxWi9ZS7RWZXylidsP9d+1ABKAXoBci7QFJRwL3J4/
EyYwbTB5+PsFcjN29uHe6Sy0kb9o5mnfJRCtZnWgWXDw7mqNWNvm9+cxRfFtuQVCXdyxoz9DcmPK
VwgYLdf4vXlarA1jDsEtCJaLkLrg4w06b7JZuZYY764JP0Jdt8ALpa6GQeaERpVX06dyEst11h4H
MpR5QuwfwWPF1LqvXo7+0aza1+QcQzuYCMYmJGbEs3Z/UF5MubyD8ziEJiLyFQ/1Cr5f8ktMjb7d
mJQBZrN0UMumKQaMUB4EllM4ycjYnnpBOkISY5F/u8wnaHMIKjpw8FllujRF7CvCqDAEwBfYFPMx
3rPP9CLP7h9ZjFMJeKhzB389oedyJPvB9246adJ4LmQVfikcmSbqlbVKMPI4bl4sA4YENWvGtmmc
rczlMrmmnPe8+4PMNzdejxiw2V2/oCIBQ0Uz6NdrdJkIfXM0oLfr+HlSOz298tBLKkBIr7kFqYYc
B+TBPHJ2XrnUv/NArE1cUdpZQDPMHRxxssjyHQjBON7oeneuwDvXmTt+ML8LUhei0xlk1H2DZv6N
VVzklH6M/G4Szng38NxWdrC4xQ5QQqlssP6usigN0yEJcEfX/jQwR7Wgi3STD3cQwlCtDJi1mln/
r83RUQagngMixPw54vVfXb6KijnvxAN9v36eLag8HvX1GeXy9IBeDjRI7Gp/HvybvQzUaplqe0+c
LfoFYWR/b0WSbSch0z2N9/qHQVzdSt7bK8W1yL5c/qlafrxqwSt75nLEf7NM6Ir7d6Vte1vZCTVD
S0jFaWSWjEgshWIm3Dd8pgLsGkve1ND+5XeVWxGxWMWYwqHqEBE40lQ+WaSC2nTzi7/878YDjRBL
XeXcqDGZCR72ydsRy/bEUn7T46ayisMyQUWBz1//xsvjYmEttR6NnR9g7QI7dPQTOn6f/L4OUcqJ
+DZakZSQQS4ncI8vYuWUdbIx/2E+GJdGHJJ+jfSchBsW5cA7KmgpyZTNi5lxqjbYatT5JG2q2+Ra
KQEoZkBMWbSahyCx2ve+ejr6Cn/e8/HunDIjwRHTLoFqbVPTbRg8KS/wATwYQsxRVDQGI+yWkmEw
T5OoShw8ofdFgJyIvzGT41v60cFiiy9eLXNomcXUPU+AVvsv6ANaKR7ttLIdET1ObpLIlPZrZWFW
Uc6tHoNDwl9SAzEN9mVBvJOT7m96D5q7fY92zr0VZtE9bjSto6vGkmf6cvDXt9Cdr/cFotxDDc4L
LC5pe6hEHRkGr8w/HZHAVL+rk85jmDbnvuYhafDk6Y+du7vgSXX59eO1dXM1wPocsEdfS2Ifiau3
eOyurQrX3zoJ9UG+10dabYR8Xs7dE7jQ2bIAQ0ZBlFgIvh+tqxVWzIeffqAFt3hydbHHUbYCaa32
savu1o7rDk2zz7BwGzZqQ4K4XnWNmXqDuxVWceoZ/G0lyZVwGXtLNANt+63I17N2anF/3/mUvf0c
3EY+WokG/zK1CzH96FpYP6OgrpHki7ksp9xgCiKa5RpXmaHA9t7JGUkP3g90Rz2Oz7W3tPuwkpB4
BAuJYVrAsUZ0S2+UdtosWp9fADaG4eLeGuU0vj+BTRYGIxwh+Eczjlwk/6jaiP+9aU+fzm0tc5tZ
ErpHNdum+5s2hBOPYhzi5Lbv0SJIZBgHPFuWZ+CJPE9y30470RxpU/OIhmXtUkCRTOtI6T1pb90i
N2JZDMzDEmfEWXeRrWvMiWF7Er/bGQPqpoROA8b3hc5NkuICHHyv+S08gIeljQh9wkku0ylOENXG
3p6889kYnOKfXxElgXRHeg5Hw/2Qp4v5LkyN3lOy+uobrqDko/9GnNA7o76D2QBtTiZ9gtZ4Yfdx
10K3EKV+2qtx5G+0CKHCIo5heIMHEcpocTdazyr2BxHXcz0TArIh8/7W6mZWY9k3LObGcGd+jTEm
ZJL+Okaclq+cz6t+KTKABqf2rVV2O8wSDk6qyWjgZqmDWWDpzhoG0tK8CshQfBsMKcW9EdJgma5d
+V9BEksa7nHxkxtztMJIVqDUvgvyeAiosjWzkGJrZLOuWbspRfj9BjpPJZlTx8V65sablfjv6Xbu
HeeTewkq6+9gwmqQBMbATBHjx0ROHmO4EhHcK1q2YvWFMAtUCbMfrQlvN1R6wQCZwtYnPoykM5AH
rTUw0UBKtz52FFs/tG1Bx6VZ8Q6gmmBC6Ix90VL0YtJYFiLlOhqMNsXD/Fo2E7F5rfzIWGhM+XGY
Z3dyLpje8j65tzHAkkqaMoXgMvn5IvXmcFrxbChvZ4gG04SMYBLoxoTY5mYXQ7sMtDjSff+W1nx3
0XAcnwr8dM3aI90qEarA4Im26yzJN5840iHZz9kyP8A0CkY/VVmdyrldXQrpFtpuUzWwQGD9kQjr
4gVWwuyRO8cP6+05dPEnKUn3ieRk8IFTdz0axGCrGb5wB+q7fvc77N2gT8r9BygFC3iBPj+Ae1Sp
eo0aP6CdaS6G6LKvQmp9tyhPsD1FWJYwDzMJ1LCIMlvNwNQwJ+oQ6MJ/JltN+QcddY7c5QHBYUBz
F5Ek/TitdUYaLPrYdSTVYBfpTya/VBAwMuw419QUPYgAztEFPt3lsM+NWJ06E5xXnJgbBN/qh3gs
kqu4D4pMINoDr/0TBmXuyx7MiQj1h3ZGyCO0D5Qyg4uNJuZE5cTHNBMOVGwVzElgK0nEJ2FmCBB9
OuM+j27M5KTHvAPoFmXjHtHbaPhFUe/q7b9rRo9yVlTAWZ7DJpnM0MFXP5WtzCbyqsFqZWFhtVoE
vDrbTlr5QxZ2N2OARXBOaNpzToj3YJiOTDDYNsEVs74jB7v+wrF86PQeKUbwFqz38pmlDBHj+kN2
Ij8qQEogzc0nbGnnFIUhKqIMKZQFXjaUXMZ9sI7snJa3Cnsn7KURi5waocHbWcZvziBR9dsGGJo0
PpIbXI8njILJhvHF6vdCrnjg1OqqmE/SEZuSRnWqaVc5o9JK0cOVZtvjNadP0t2kvuH2t0GxHZFT
H2jvn0SkFBOFgXu2Q18KgGg7i+inZmHBWPE5uD9Nv3tZ2hHIcmryf3NCIPBBo9Q96xtvWTTeSM8p
9QsJHiM1VXQrFCXJNeX4bUgXsS8k7hFcPOqDzwP6Y2c1stKWe3I07qPJEaTlZ2bw9pl0m57zD6sc
H8IpA2bgJTTy/t3YuCK7KcQdcSHwdck+e3tXTQymRxupWtiqDoQlU0h37c0T0wFPJvZyDSMR5JET
vzedbdLPg0tw+/YHvMaR7RT5LALJNedygZ/bcULZ7HNxio9JP0D8s6iVMzemB87ZMHhlg6XLzyIt
Zbs0PEdNj/u5UdSBeQF6nquNbMOhmK4hKRoJ7gkDIt2XfdQFjMqDfdDQYqwxKhEkkph3ggmjL43t
FfdRsginDdbD+MoD/ItIZXRNCiHdzsj9xGbjXhBmoFIaA7qP2ti5UgPlfZxlvsZqEoYmf+uuFa/v
HfG57aGNaLzlnijY9VfEd69aPJCT8fL4nP44mH/WxiGUtbHsA+t0q+3IWU6Sy5IzDzkKr0WoHOAG
gOWcBr/NU8PabcVZ6Zd3cQVtGl538+GyN7b0zOxSdgNvHw+nebXBNn2I9Xc3+kndqPTCO/oImCvB
3BR8ZzQuQSwhqCwaMpTuffbsObdzcA1BUAJyM76KFv2tlaEFFUe/KVz+N37zixavECRZjvfy2Tva
xBlL8H3YRtcjdEYZ1zwTejOQTCNhljMGzwMwexroIyTjVr5ZnAb8nRpNAKyhWmRGYrFAf3Nj548j
ZbjInT0rcV74x7z0Fe4dmDwKsvE0sdavj/pFltgQJBbDt2+Kmwe+DfkJZTvkrX1jAsOONv80iGYm
mSRDyA2EPOm3LqZvUQL+hY9nVk0fy7RyEXEGkqKSnksAVgaUbx0EIhEwS5UdmPt/yGHbbw3gyv1l
FqTqQtGJvccYdOi4EU4M+/7cWhoTffD1NUR/pfafFU/uB/WLSrQQV1wsNSgqursLV605zzL64raQ
6tQTa79jt4ptV3qR3rt+w28nbSXSbokNU3vCvsVIaYzEQ7lRXaeFFFAcJTrOiz7rI56iE2oOU1c6
VXDoGudqpb3GYtRCNd+TrpnWIeDve73O7C8y/nOJon9wBQpCKScc/oyEpx8vnGyCIN23wk+f0WMt
CbrARVbneLLN/EriLx+fsRyjLBw8eC+E9lpgk7gq5DU8pXv2BAOE4yYMF1FnOesoJ1nUsNsPtyAn
BBjCNJSeAzvpwbXYtvbRtM6YEKMV5AXnLz1tf1kBF19Hg+jS9oTloI+h/myQsPQhh9FI172F9D3w
kxPdkeZhZS4/cIpdT7yvr39idgmhVoHTPI0YzkyVWYQ7KOcrGcOR8TJem/mGkkcs2AbUQTnC4yVi
U/WwzEn7FVpTOen90cioUJb/LqSMG1X2QXgf+UNZnsRzkVbEE4wfi0YbThEUNQeWGgf6yZxTYr5M
iWVnYC/myhOsFTots7BuIwsI+6dUc5u8q7TDQTWn5aZEH77LegOpi3/ELeLWzK5ss2b6/cFz7tn+
MCCUlzP+d/exoMQCrDmdI1pnCqWyM/dBpp28zRhi5VjUWbFfRbkfGXWivy7OFH4wESaggHtrWm+t
vTdK4kl6rF+lKUssp6DHRvHn7BMWa+V3X/OjlJ2V+ctrilJIW9P6JQRM28Y4vbzIVy2RQlhjfp4P
RpK8MMbO8hLL2CiSWAaGIjb5vAOmIVS5jF7gG+Td9U5K9qdbkiexyts5m94LDZFesbUKlZWu7h+z
CjHHhaHG/duqI6mRF0N0vweHfeSIwQ6/orK4QCmH/m4nTSbSL7OX1hmAhmWHkmCuFLpc/EeqMF02
CbZg8m5n/U9YK7bjBg/WfQfC5KJgPy0G8E5ednWDY8SPgNUOdAajOQKCdDUdhivUh7uZjdEDglsG
5DphQWhu/U717nkAP51NKEovisLH2HR+zHph1PhnUFpWmSlopG9vWOHgeDRX5MpF4rtsxt/WuNF1
s/E51YEZFk8t/6zWhmr8+xzlTRLy5HCeVjBvstcEHF1WHzEeKt5C1v/laZjyNb7GwvSkvGp8vwD6
etA2NtVFZcX5IVoSI7ltnV30mg9upgqNn24ykyLckgh7YscMkJTCYVqsEWU7jVCrtjgQb6hyPd7F
lHjHG1NoXxOHpgJRmGP+nhv8EbzW/S5TSbCHN0AYUDi9gaLnP54obHlD1vTdZxRFc0IjepO+6SCI
upLqYCgL7eYLP7ENyRjyXK6nVudNZqPYCkGKPBtPI6czKUtSKtLuMlgfPdmyA+1VShMjW+teEcWm
spcPYFyxuwzxVnFUuIQ/4t+5PHTjYXJjbwR4OMhPP/QdvFFE1KaDgqgNzpx/dQ7JaJUMjQaTlezR
AIzMZARAtHii/RdLTYBsQiURK9tKragpwcBs22W18a6fRNBTlqHZLG4WXabauzuy6iuAKU8OBi7p
AIH6VdnKJ2P7sCwrQilGOt3NJbyP8K3lUAiANUFQmV6VHENKSjpfw6viMfhsW7MRbqa0DGS/HO0F
d92ISBTrXwYtIjmNvTzHjQ8wBpM9gAF+z/ehg3WIhvFil+ucwCx1mv+9BRYTlTHEdXUhCqDpzX9M
AJuj72vz7JaknMd/PDxL/BDiufVaeL9B7cpjkJAYdn2uEqppK39zr2VG8f/4/Nb4p36xolRi6FO7
k3hjeLSkxY1f1AHcXriO4rRrQjNmOKeW0tUbPpT6vTTq8HoFK9VCijSKTgBiJFrCxvWlLEDpvR/5
/warE2Wy9Oxaop++5m3UDimz0HUGYriADScMTxJ0f+AE9p9UuwoiDy/oLnzberua69QTfRRnJQaP
3CnMt9VXV1ySJ+7y1P9Hk/7s/RmLGM8Hn36AxsAtdjwnn/AfbMQSb3LLqJwjtE99Hdevfx91BXtS
64bvyep9gb+4DM/TJJ7b5GV34MrKnTTnGpgBr365VaMeIk6zyuL2GFfreijgqsx7QaX7gj/nOgeK
ovG12lLvQjtfprm3WhBsdsFlrCz0N9TDAZ1Ty4MgKlLOSCuMQVFfal9tywa3NcP+14AK7DMKNCel
yh9IZGfXpgueIyw7vCnA/fM5trWt5ZlV1Qsih9Deh0V0T8tPoWXEoWPFFa7hk8FpCx+4oP+YJt/3
qAeMCfRa/LuUndil0cwsPYy9BH88zz8GcoVJdKqH7OFKqkO6ewRnbZ3fskqZl+GF9jLQUgOROKgy
MmsiWQ5Y86gvqn09pCY+BXp0/vh3ugWn5YegRSKb6B3B+o6BLZR7TNSQgOx9yW6GWEbUHwLvFT2t
v4x8xLmFVlivcYF7uP+TtU4Oc9Y0kFpsidkn+Z2Op2oAmJYx5Lgbq8fn4LHTmpy2guPw0iyO6Fey
XyzGp5l7UivTirBzo/664OycjDP/wL6V7hMf2SDGSoQwQnCWZj73Xaqy2ltGZ3HnaOvDD52XoV6y
Ok4p8PLuYxtnvNxEEhJsLtBPlgsE6oN0fKjsdlRZHkqQjE0iQklTgVZfBNLddvFmgMj3XunxloxU
Zta3lrK4gqtywvgCbQPfBi1lvn7Vh2wu/+kufN6D0JwrDR7r+djCCVz/j0E2NlO6//q/9DixM37A
f2jL8sJZGqS2FrAbQqnHjCuFBOVwjliGtwUHv9XSU4xXzGMYgkiK9OwpXEA7FJQayjaymOUOZyur
qOMDEFw5fYY95QujZ0PJz9Ac4ShXL8WO61GynKwaQQlPQc5Jniw4/gfAIbXByLdVQspWq+nb31Y0
xkTRPbMvBOjA9KvJuoyCxVlvEHzoEj6FAwKfOHNT7PjEW4ssrSMSPJkNIQ3IxlxWMhXcY6TtvFob
5ChferozJMUnJwruejb+JCIxlitzgBLX8hRo24mA2ErrtYNDrMJ5Jx/obGlgaEoa/wR6RPM81Ixf
d6nzdojEz+KiDc0HnyU0dMPg58UfoZA8fPdeWmKRXuIfudcceGVaeQgkNzhQVogeQrmGzy44WVhn
QNKeJWdlai4ojIHCoarhkZqmYBUCPZl24MI3Tzruoo9GlgQZh5vAUtroyaEeIbVo/gze9TIaXf1j
osxCo6DhgPEBMQgFy2HzIhwD7kIfe1qZV5/uZVKAqiikIImizigX10qOagCn0lDOW2NwxIi+rQcI
TQFoWtPP7UXcRKvMN6YjrxH+AwAVZrifgOLNA2GZImUS/HSObST6b/6vJksxB8h/OaaDPBQ2rgdA
HTvJiSts/IedYzrlWRkqJeGfCdDEx8URsHvRiSW9/9QfK5sLsaH3dcQ+t4XckDvon70C4IWzmzN5
4riYbfRNVlv8NRN4jCzXNtHokLhiRoa8V8WLxBhRbc8TeLu4M9XI0Vy2iKdcVSLFCIldWAWJt5bN
70kFP/8rROXs/79lca/r36HlXSOvqCA5yY4PmbFenWesMiRM+g02V27aeHyeuI1fB63ZMA3oURXD
krJjdZiMsPtugauPVwkZ2JPnNRWeEvp/IkVScoXVJKDOQCRBhDMHev2xPImDfQClZ3QrQMlIwYgM
6jAdFJTY40wqwpmr1JcWeCvIizJ1Pdjfc1GKkPJVKduA/WWh+kQq3uCj51oxMMkJqclbqPSp46gG
qDvk1oYwFhBWMdkk/fpI65J/qeYKX9C/UJ02vraHC2r+Pv5ls4+u8lSQBL0R/aufVuFSzvFlIvko
/k4sa41GkSeW5HsOVlUu1iCPv9gObe28jEEh+7fiO31BgjqUh4CXAXAo8rQPZl+XzcTSwGO9K/Kq
+6+gH8vaw0l6DwXpzo71DlwAAsf06j+qE3S/NJHSBNOMWEsfNrvWGHyqdmp9YVAf8TrFILCR+xW5
9XWXENS4KfwfeIbvQJgfdfaIO+XrUwGZY+7yrDSNtfeeJKc05ZoD6fLHEevi/1kIszjhPxBmbQqV
1L5BnQo2MvibZWkj10Leci6ukvPAGlzFq0sHeWh1Gl5yjunpejnbNK4IWVLVU48Ou/u0w5/H9k/2
JMfgH5qVjsH7n5idbFC9f2WSKEhFnyYMNh2vKuNRTrZn96Xs03aRF7JLxz7VRkIWfgzPq8+sGAAb
5iCMm6ek9AcbyUwUZgRO82CQ8viCwxQtGaTFxDYkGxxnJZEDN3Ue7PGHwYb//ZNnQSN0TlSZlHlZ
PyQINwByN/sZlkxywPwSsoZ8VFSfsfe6h7pMM8HH7TEjs7LIyR7kSFOu+o8jcIijQafKIu8pR4Rg
z3g7mVthTnUL6JpUHQzZOoZmJ4Au2xU12bQwf51q8/yABYUpwiYuL4smPR6NSCSCDx91ij4egEg1
GkcEZULA5RzXN90+WqNNnKowciCMQsKGUn0prd7UTZE4r8wR+M3PjhM/wiymvyAC8f6eVkA3nJg7
Tpv+hZ8uC5P6RbZREmvDoS+uF2vdUA3bAemnCdmjErTRAntmGH5AlfikDwMXWuFWgtJMEKnzjN/a
DC/gXjCGZa3o0lmxRgBsoG/JzxYLsmHPBSpcm9KviBDDacogRkG0DxbPVFBJmfJaAnx2Sx23sK/9
Rw+/DkTOla4Mj/g+gAlTLMABO4/7lhy+ftqbpS161DUx7DHdT7SoX+nvI1teAf5zVDRu0ojCmqi/
qD04HGIlfDsJixUrEuws4RIzts3ZO34jS1lsIRRcqp3/dQBHuDtavAbbRpmTQZhbHg+wTaaYaxky
UL7uXcwe/Jms2RV3flMIVBxZLIv3FhTJ1kn49iBo4fklE0BkONmcO6TzQUa5OmKi6P4VlmKWYufv
1TixwL1MGxUnFc/lcM1c48PYZjviqLeUp4TYu62Gd49P3fpScM8ffWGHBVyUKKJpYXMgbN++hCwT
HeD7AO5CUP85JGcaznj3Huo6OyMCQII6giavfQaLT6lwll1/lbAPZ1zHhtZ7vlKQTQGAR+Rn+2Iz
30UuIs9PWIvQn8kj1nW5yWm1AgmKIIXZ544bRF9NIfMm0v5nOokiu2EptA2u+g/9K49qs9s3uasV
lZ0gHo5nfe6x2hDOI5J4Fj4VVaMXFGTvtGnNV8Mj1N07F54waEDeNQ+Wa/iuz39QEQIhngbkKQTM
unFpzSnsHlr3nS8A3dlSKVck9txo9N5RBuDd2nSmu5BB7Y/w2xJX4CBKW9jBk8EzpM5ZbgXxZYD1
uxEJ+Q027hQkip1FqJQX8w7nE5n2wwS0XyellQCPoX/SO4uFwslM8dY/1GHvrrSzDNfBXCCtwO/P
uGZi68pKu96TILrNZdKuQDStF169fpoMxZ1F+RQ/N6573efaUq+DL+AY+7yL7I3+KdFuHyEWt5ol
pQtzYV4E1y+oy3+1pyDalHuIRfxNxkqrTV3EbQmM/TpCFGopIyxeucX6da5yuow8w1rHVozFFobL
9dYwMsS1Fu4COeQc5tTwDJagorrKD/Us5V4gvd5Y+R54AUjRM14mWQUv3soevOLo/Ohknz5P+7yz
qTTQWlwOOlD69YHCuz4iocgD1H3KLZ70nvbPNRo5R6k6++sEk8JFvo3AfYhBupUuGCwSibm4BhrL
tovGDU3Y4BzbCSAYIN6uWlduuEVFIHUXGbKWqUuO6f5q/J8x3SkAxZ4WeN9ubxrnnI/FLCJi370i
Wmt0cpaIIO+uy4xLjsJnLj0upQBWBubaZaKNK3v8/L3Wmcs3ZaK5b/PatBh3CdKQpRyAJo5HtWy6
yc4wGnx0r2CvStX0nYmVhiH80Bejpo6xm8A5D62uqL3iBGmePiKnPAQaXaQbBg4pEVAxpAzJ2mct
9Cv/ZdqZP5TtEHY4ch08+nkLbHaWQ1H5rWj2SZtlbm/N7DjEAj4oIzGCNnC/lMVbqgFTJdg0CK8y
EAiVU3nJQg2TPqy3xOPU62HPOo5Tk3hBkSNVYdfrYqmSJJN3BLt+DAudJN6obBt6kLcMIDfBIZHh
QXnmX7fgcPsGKeAg8lxS+OU9Ep7u+2ojuaUWm3OwGkrbgKMvdLsd8W7EXL7XIXAvuwUDeWkU/JLc
Tval79vmPKhtQpGAKmfHEigNcIpvHSvXXbN3ibqwPzklS1QyCDqfM1ZSk8hrMxlo6cnDGPNBI2SB
61mBYYxCx3TJtK2+Rny7pGNbbUoAe4fPgxsp5CjWtgV0ncYh4os4Aj0ZrCh6rb598FhA60mwkLp/
vCyI0+6xvFI8Zx4EzfY2yz/0zpKKkyDKkbeuadkoPkNSXFGq5iZxsLT8HJAv+lOuxqqRfJB6MxNV
vY9p5AmsZcE/qZCO+icjegaQzuXwbmJc8x1pQ0j6GAtzhHBDwqPm5mzHN/n88h7oGAWMy/OF20bE
gMj1M1HydyRUyfrjRHj+o+C4EhttviQqRBkvONq/+JffAnFFUHYwKd8c9Ix3B3pBjJF4ATigQ75l
ZHrk6FH/5xy7krah2OhucUvlYSrbgkCYFeXAy/W8RJQh6w+u9P5+8litJr6GCBxdau76aJJDPJ5o
X7f/H46SIIVniEuorOtprMbskze/fXAnjk/jqna8eUMs/AQ0YdiEZdQUyY3wy542rOKbz0U7vf2u
AEQySGHvOopRjrFNu0e2j60dcMTMJW6mOBMl4KlXgAJw7mmT04NQf7hjkAeV3c1X13gxwa6tzwUw
lS2G/FBKmuAAthHn/pgaOAUrfsm+FCYizqXbzH/cSASqBeyZ4a1R2Y/GtgFqyQzPDJIAJEenMjVV
d/f5YcERXG8pxFdZYH9cGrO2nsszuwt4RTBSepUvS86UEgEOAxNr4nCJDbdIYROyc2ycn2YrgoxK
dDE66LLnVBbk8/Pbz5YrO+DFlho2SyVtgWKCxbgj08cfdISHBjkwBOMzHsHh7OWJjDBy73t0LzXx
NzzcZZnnUQyv+6++RXtS1IM49bpxX7XolFbzlyFdO5EogNrQwjKV3TL0fhW3+df89BXSdMyN92mv
nn2DYUVGEX8eEV5j0h0wAeI9QxuEbBw9DiZFJb9r9CN+EdGsFfKMfxoh6ioeWXZFgwU7sjlLq2hP
Oow95qk9ArR2EJ0VJ10WOpmPXrr5xePFqi8gmGWE+q1WEvMDoocb+j0y7dDIqWAKXpHb5ei1UZci
QU5iWLPA3aP8yQFLnd7wMzrrZumCmqA5OwcPSyc4eyOV6X6GO9A4qPz92gp3SrgYYccWxwk7J/PU
HUMF6t/5XKOc5hNKPrn/sXXQGhdtP6js7drA39d+D+IoxiPPYrQcxWbnRXWe/niEt0A2RqbppbLL
6uFo22HeUD67zqwk+Ub4asxnc6wbDyPgZB0G2/2BUA3BQQVT7cw/1h2p9Yv6es+ifR0yDWbgkbcF
pQyyKnyzs0+NZGOj+vge/o7eKx1xxJ+ZXr5x203CJWhiUGtH3sJ6UgCNv+K8A2qjMuMJLKCbiJRt
2zhxCfGw/A5L1RdGy2EZeNokBcL/9Hd9Yklm4VeTuS0i/xtTCXk0ISXIMrt98ycVpySWksFQAWA6
tdMKzwPczAJmB4IOZJzG/sKmVdKJ6qINoZwgh83InL97oNLPDuEXpzw6LKwDlax8OVP+Co/LkpQQ
0QEsQhh/z3QcbOg5JdonWFGARWWVRT0UrjCcPlnSeqI0O3mXOkjp4cmWeegxuenlmKP20Z7jBujd
1LplwkRMmF1NOzRU6WMF4l/GSVMmVQzP7u7xvKFOutgihlDEmYQ3as5bORewny+ypupmlaq/rSKe
MmHnMzU5Z2hMFD/ImZrPIdAAuYd+gCBTFxROhnEqwnkDcL4qiLDVdU8MCWoQDlcuNFSj0oTpwF5R
CVpOEs2UhMsjK6invUf6JTt2gdOxOYvolQxQA70aG+Yw0LE4XdWuFagmmzNUVdacHXSdfvg5Ioh2
wJTkb+p6uI/lwYvENeCa3kZdT7cskvu/slwqWPzrMZOqhPeY8BO+b1GGt4ClvixYlflSoU7KinYm
rsdVDvucH4aF5v+ubk8dkRepEAu18PYWMYbZ78g543Btk1N5FSWCF92UnaOpxA8b8uzrrJmDPlov
CkJOtfWbEmib01jHk0GxcXZ2qT362FN6ZkdS9IboX5R6cPDlr0BQOd60T5IhZMdeE1Kl6M/YR7k8
WU/167RPpFz4qQ3ENxYDQam4KPaWq5YgRSmdsnHHcA4DuAd70mv7QSJ2QKClQ5fdeFQMc4F3qXc3
yCSq39KP1D7faEzJW/+eEwKcEuv4pK8X7SujdGXx3n2apZNCyE6trIdidpWx3GGJ7dEekDGHJ8CF
ZEp8wak/XMcBaVi21bFLZVtdfAL6Rwkx9KcNnor81uC89mezPoTBXpFs9HinDGkzobcagh97hIRo
Gh1UNL6Vnv9vkaEUjT0pb4TXGMfVUTyUrfou8iLS+kDmphEvmyHHqyuhvqNCmWzrehSkwNpT0O5H
KqBXwb8IIU48wEFPFZspT+mv766KUkFaVdcy1rav81yohZZ+h1ykEut5wVngPwRYxM2iUudZztCz
INkkfOYNyBm4o+ZJjlOo8W0fxwVATTsxjF3HiFvvHeswvycdkU1uvBf5qxnilZyeJVkd+DA9nQ1C
MZZiaUFr9g14W5+JRSTkA4wUFsAaTJfYVItiQj6CjRDIIPI+LmglY5+luoWuFFTOqQM0XB2xyfHv
8ZCmkgN77wVYrX074SHSlB7rIx33ZYWsg0Y/yIS0/GXBAYNVAZ3VHB17W6z3nySx4zXhTxh3vm6m
pgFL5ytqZBH2L95lZcKPp+OomkmGn57a1yNp1jIggsRZxq2e6G4r5ya/mhCBHCPSw1obWZzEjYdO
gKetqtXJc7ICjwwJVnhhpeAmB5bCGlPZyDGZVVrygNa8j9QMchBGrhgyl19Eg62IUc0ngGBGP2OD
jHFPOaoLH2ig8Wkut9bQQUvDvRaio4N0AkPcznoRKUvExIX/IfxjOevkGcnYYHJWgTD1ssyp4Tm4
T+FzmVtgoIHOg3Ul4MFDdr5jjz/ymxQghgfnwQiOp89WCxmxDNFORqCI5zn9Pt34f5kkkx2JwCHl
vYXUEB7UK3lmvEzPKDtTcJe3MDiKfzbkjcnMOmENxc7vziXJB6gVG+NC3lI1cEAGLaz0Nmd9sK2D
uC+pHGcub1+PdmsNuor53K0hkOz5U31pbo2fPD2m21ApFIXfbfQ9eIAKzP2BoIxfoI9gYx2+y/Yu
w/0cMfFriYM8jlyJeroPsn5XSrbaA2fP4bvlonTiYgBGGoxZm99+cqvXada2udPFcwuzWCCpbaVe
g14S7sI7gMNplNUtjsjhd7SCVkqJ1UjpswDqqQ7a9LLkmH8BAqEeZKb6fIzdAY44HH8xoHlCWp0Y
Tq+w2mrZoAghpdXHrLINdGg0BPC70Wer4UP8Zk1xugGSOKHn7cKZipnJRZ+l1Do8sFSZePxrl4GE
BAXd8FbQWQZpn16q4yAwDFAdgahfXz6K4dDgzjLaHkf+koalfmcRRaKqeeT0yTp9Jb8t+a84puFx
JWvysR8yi1CCgWJF3RoJUVg/efYlOIECn+tziJeewBzsVBJ2oAp2stgd8nIdvan1dr8QInB7/WqL
vFG+DHSTmy5QZEGoznk1H57M1lhDT83XP1hbvPzw8xZH3heD9R9u1Eo2IGijpRjkoManv+esLyr0
SUwcnQlJAbZpnnH3mwRxM0yxDlCmBdj13ToBVhZ4VSEZaSXzp9gMomWW72eN/YN+LrSP3XQngReZ
cdCOiBxv+4d9d/KZLUoLuM56fbxPJcL6Ya2UIN8PPYru1b/HWvefb0hpcgCahEfkwqmot59vElIZ
wM+7L7BEmiC9c6mqLTpIdcTaL35ie4jCODvIsJv1G3bNRFD5adeqTZXsfW34/yClckZWtCbU/eJ5
ixC5V3DAbP/25SmZhibtIAEdvDrO9xCMeGJo4xRY0tFlhvtszHq2wbDt6VHl5yxtFBY6i2bgR6E7
oxL8txzn15mtzVP0vygD89FtDMFfsRYJ3DjTdwQJEKUkCDuOJvvc1Zh1ohF6/QjgTwlRNURjjVgf
ERHCxbzWstvjqa+oasANCNNRFe8jgWFBn6Q8NKMjtx2O1bEXcTcincsIy74lzs0gOAfDUmeTBrW+
JxO5meY7McYSuBbetj4UPKo1BtkqOesOPmHy7k1tQUd/dd4SV+io3sDo1R5SA4W75vXlOlTXNtxm
5WyRyat+MSPPd1SW2lsvewTlgw4Uue+Lvhp8ZTvXKbCGVbxyHxK5EBHeBp9vx5cHrI3aZPq6eRLJ
fOvl2PP12HoG1dRFx+5WBEabeIDvKoeg2n+bOO05WilHAecoCGXHjyd5fBFscFHyNe22Yxk64BlB
f2xxUqqt0BhMETwvQZiBpiIkA8h++2cJUfac56MOy5WXaoXj1umJlHM+ZJLxI99MK/rXo0OwZe2q
A6hKrNFYiwwhZ+VSYX1b/YkOEBLAIqKZ61DNdIBwd+Pfa9a+OBgHYWAvPiIa3/VERK1UurXqvNQz
MSzmVHF/O7u79m/udhbC4tiEa4T9Fj7zaKEhMRYWuXYn8kcfPY3nuuMYy7G10pfituzihcTENum5
riG7as2D/qaJx1mvSzDOUD1oq2Gaj9a3kBmo4PupZjKn3vIj7szLOpSIxLkOtiVdkICe2NNQHOMD
JBGeendD/9x4rr5uhudu7gL8QnwKp1Ip5luh22njFwNs4gvPuiCNWH5dvyZlvMLaGiswpP7iJBH0
IhPeDabzP9LPhO6N913XhfQhFu06y6oRkAEmQtik7ZI4KmnSMxsz9PLbBWFoKC5GT9DRi3cElIzL
X0NXFV0Wbz5AjLWumPqEZAGQQWp7WNovrisDk0hF3eaWjq7HFOZZEptQRBwnn7eu7oqKtKS4brnS
uDts9/lr+lai4YhO8rwlJ+lvp9O2JpOW+IMC7PAMXiB5wrs6Te+8nrjKA9BVwPZfVfiVYCdbb4Lo
18/XyM5XiwegbMsV35GOfAJYhVM72piU1YDitcrxr4sGOz8C+QcIulb1Y8dzPOryakZkQ6emDPCV
+mV04oPVAkD48cvrvtGRDNZ5SCHjCRNHKzL0yX+vzV5uP5WANVBn+UEW+Q3QDPdyAv0jcTwDs7H7
Wdv7uPaPwxp3eldp8bXoIMcBtN9qs+fOIy+7sc6NXM8Ac/zCeVdvNSlgN1q/Vo8Nye8Ikt5YkWfY
Pv/fI5GbZ2Zpo5ye2wy8kmjn27VkEKm65715xLhPQpPUwSZQ1WfsFzrP0rfaIBArGrmbqy1xyJaT
qTmHZYBOHo0oI9apJepL+A5rDTgV+cPkmVmo8DbxFhozgCxjZaijJkQPpKUx32yPIP/iSnlJ1r6I
f5x3gbZdDaEJvfeeb/AaK6ZfORK01Wa2QQY83oU1eyyVCuer0w14DKQBXReogrirDqX3ggXdd3oT
k6XA+iry7ZJIXdhdos8XZ5NGPXBrlFTGgTe0cBGrfBwFs/EAe0F0jVXyUy2ukqBAVcZ080zzDS5T
abRukgMvGz0D2GnPjXajKkcQRiUmjQuE+OxQP7CUIZ1PLdWw5B8qSVI0Ej19R9NdVbnV93FWg5py
nMafaQwQa8Jxs4Nq3u81FJQ1rTfKv5nuN8RPBrfiEbpXfHzD67I3ip27F9XO9MJRY72tYsEp7jdA
p14KHzaFnSTvEN1QMtMXj+u7dW3g3YHLE5L79/ouyAY5obHXo8ZAjWU2RMl67yqFyNRM2qPX+w66
mUmtIkzbcsrVmk3BoZVpxraJN7J6o/GgTcgrMTHLbl7mlkk0niR0i+pR1N7mMAHR+AbCxS4USKOl
TgWlxvpyvkMNml4URwampQLNre71xKpLLoS4d4Nq751uBINo8P2xBeMtTug6Jb6swcYFz17UcKTc
r9JO+9Nqlgs8ZwNWfk2B+7wnuJ4Hu+32GX34cWjd5LEu27BnEvGA5FgSwjIvmS3/S7+GGJ0XKqMg
wBPD0nwhSQ71b0MpIywzwZ6TFRVRdcLGTMxuXtpY9yLND6twX8SxtmXG+1VEwo7V/o2LlB9IE6rg
LxbZ9QSB4cQr4G41dPZZL7HakIfQdCvJ8HW3PFyP6DMW+Zo9S4I6wV54avtoji79kz7nE9msS5OT
qfvCutIjTCHHsWJ8MS9Ql8Y+D0iCiSGzBc9JeUAEYBVhEfu0VkPbGUE3fdTQa/JTzdGCaAqVVnSP
j102UezvbnQkuHo88zNf5iZ7sI5lxZeBf450HWo4kGcUF4670J0Eo7+obqtO4X0zZHr4N2AUXXM5
uBGg0rfkusy4Os8jz3uSL3DIwPDYogM5o5PrudL5xHLNN2Mm837pQ6uJQay40EoJdCjvGjLfi14N
l2c1VQuL00y3ppBR4T7WqppgKJv9S3RgIHQy2gA3MrvRB5w4g0fbfqCMciyy7cL2HPAJebgqnjzZ
6qrUDHcoIjZ/vFeM9LnyuwWF8bSQG02O/UAcqFHkRP/pT0EY6o56Hf0GN9+4ExDFpW6RkRjXjZ0B
a0RNkH7hpM3uICdwt9gXuLYQXGJN4DLAFz2OV4iUFt1owhS6iSRW14Dk7Sfc9WqBtkPU0WKLTEN8
2sBcSm/Cw1xuB107IhtHBEdWO9CscmPVpBlqRT+DOFh4N5rFOomhXl2eHyQbecZ5KMEvwk0uEpqy
dVVJtvkmI/N3hy0v1yWBYsR3gh9WCvF+bPaKyxhQ8tcLZyyskqm2ppFdyVFZnB5cDcIYb3zUeBzk
dhW1Zb20XLW/onp667+12ALHdShxVX1aWxqFiZT3wMWCBWSMx3J691Y2UEQ2tajgLkEKHE9oC6gy
SD0RPrYCkNvIFp5KCIT1m1z4fhkarAPbW1FlIicWwmqiTqJ3DxTZjlaLEXA5opDt0aZ5XDKn7g5d
JckviZJQhEQAOtEkDZcscrBslpJEG1inTFZTeZnAt7FZfD/h7twQNdLNyHDs95mRv9vBJKz4zwG3
/u0G1SPqvPB0v/Pl2Pj94mXBqouomN+tZ0fnOhZT6nij/cVE3thRI+wANIXFtQKl7GPRuN+6cxLj
ET67pBpJF127V3YkemozzLkN8V3gQsVRhfNTfKqjux1ezUew198fDdgBZCjjmCj4dr2MdNM+TpKZ
lHuBJl575QqR4HR24Q/ZcTpdwKSGNRHHhaoK+H7wB5fkl1RNj0EyQpXSEK8/eNtCL2N7FY1LCSlR
jzpmIxTnPdey0bQUmh8EaC99sVbOQg6sG0GGUvrowmSPfRGBzfnyJQ8tdXQ2QgQ4Sgo7smEcSWFc
crFnrlv7IsRLnMzcX0uvgDD+OHXA5XdNrOObGkCpdvWiVv8X0xa6W9OudzHUgtkRXX20eKWh1RQz
VOxBHjBUMLC/e0vQhGIPMoOJH2FYw5j/Ieu5Lq4shnnZj5s0pMQI56DNQahF1n7F3FRABKWhSMSb
7tvcSWWwbZHlf/dAwWvbdtQLo1uVbXssvbEwrmVYjQTH/UU9D4Pv/wu97bvnBzGKQIPZKj7bHVVU
ctrCc99MUfy+73zfyYgZiDKwi/o4wVoPzRKc8id/0iMttFCzhDJ7WI+M6ihwNRMVWPOAT0eoxoHS
HFvVTr2rGpNGGDWDyOclXyjN/54/YbKWg0JszgyVYFIDoKBTeKXwykBa5M9Mrs58iIwFrDzPdTFi
DOoqOAzbSfiULItFsN4ZAxpJpueufSxwdnoU69LKsNaZRTqOnw3WetHWkE48c3lTvzB133YWWGET
tjWA6E5AEw6DQPhX/IJuLX6bPt2iLhal6oIv5JfK9bMU1B/k3n17bPmq0ksdXH7niB2q80Zx9b/T
naQVehsERV2zeZW+4+/bfr5ns6Flh4TG722IhF8Eh49QaZWDK8F8+MTmel5fssgyIcM8v+HsiNlq
5pK8eqzQ52iGO0nKTln0WmsV9Y/BG22VBQ1jQSZnOJMKLXDosHkda50HBNWibWP7NRp9C3XcKXgv
uyOOV/xN0K8lrQ1rRDLkJLQ4SBImdlKFISI6izFsW+GgHT0aSzltN93lD/CC3w7usBsZYF+dQNSF
CFQc2iG4LQEVti37+brz7y73kcdO2GSpUiTZ8ga1W5S+xosnaqwuirBAXUXGOWmCIWsydqgu4IP0
7jEh+HoNrs4wdBtq6iMViP1iK5ri+cfNxK4cRRrki/hcIUBgG0bbmTF3YGnxvZ5hubNBay+7w5ss
sw+mJndNj1fBmds7efE5c5X3nnFWjZ1o8DcExwvQ9D6GHDRY91h8vgcyXwHctU79u958syeW2ima
aickN3nSctWDb4IgcTZuiD5X5HJZfXVEU9WlFgMuMvAyNVcldeDoNXE1I1bLgLs6TXhAZcBH+BrH
96o3e/Xc+vP/hTEtJwENaAO8tlDgoomXtqmmUb6LmhPnXZME7J7dscF9jTzHAEgkP7avHa3q327D
Ng+44z7nJbJ4HxcDm97EktteV2rha5UsBt80uVZoJDMRi1vHFe9kh6qM0DtD7kYn4Pwo8E1bMCH0
jOc6lWLT4+6GkyCqTa7wqjp5cM34bRay6zP6ZyDtBmr+Q+gDUM77mhWZFNP3MgiPVdmXkrqU4E0Q
dGiU5QidqoNhR7O1SFhNqUtdDeNhbkghYUt2mvtKNaKhFseCH+rhSoo73Pgheg11xt56N99fSxPP
gq4cFanyVSTBBTnx7A3+FNKrVPAHTb6PFwnS6rp+CA1cn4bObz8/Yb4PVectfBo9W+fatioblmd6
hch/ikws8vQrHeojP63IhvxHa34OzP0YbxquDs11iA+oi20fJU3LnLIbjl1RkJ15FE1llc7Xkz8L
aeUYTb43JCV0k3aKrxwplbMLTWNu3l0WRldxb/g1XaT0e80ABMseSP1D+41MSJCtEU+F9cDYjSej
hNHs4TXW649w6a3v22QYQ8R4Kgwq4MkUf8LVO96D4id+ELNdrxA//jYlfG9H2z/bZ+LMA6jI/2h0
ht/owY8sTvyYYNCLW9hfrtygHhzAHu6kOMLPqZ/gttDx3fOGosbBhm7kn12iPNCjpU/reF3v0Cuy
DQ4jXjvKtxI7RZqQkl848cvlfZDN//yGLWxPf7RwGj6mTTvMo6bl+SAQImMbcv9igSK/lnAfH7CP
fx/KX4R0WLXKRXflYzdtuAdxKHlyN5IKP3V+XbzzSO5B3Bm9Dpp0pxbGhBTx6GAOfgwB3gLXkgFa
Y2hJP1n75Leh2IP4ORGAJMEokAMkn9HXsl18pN8uCNGdsvqxnbUlQ+cpuvEnBr6TwwzVJthF6dyI
veuAYMXPzwVVAAx6CrYGirw7Wy626lsZcEfe0lXv279yWjjSdcfYRgZF1fZVolTyn+PhHZXeGpt8
VKE7F1gqoaTICU8qi++BBNWB5XZBfKt3v6UYg7pjs0wPLldGdLJGh76PNrMv9NOq65nGv6+ExMUZ
cKenh7YSB8VIQyM0mrE1/aMKvGnu012IvgqQEmhLqiOnIUoB6xyqpkmIJ6hrulzyUMyke/V5vcn1
GX2alaEbTiu8Sxq2RRwoovjB2TTWrGBNg2I3HDXaSHzZLC+0YDVp7uIkK61xOelr2ep9osAHqjnG
vOuSKUBBn+MNXcf5InoUakT69ZlAzYjCHdDjo+slGa3nw38WbMY5kMw/PUW1WxhIbpRibnT5ODEN
9EKhcjE+g0oLWVpG+5rxK2sTLtQjR2Wkg6wqII1wVFI2KrpUiUX5oGyP9aP8vbUtgZ1s2wlrJ/xF
H5+qxkqlw1/UaVIh/tqtecnN+7WUrG0am29CzGXZIqGKGYXSxAG5h4c5nbv1HV/e1HOzw7IpIJVO
BYJ1CV2Vg0v3ltSJmg205AibuHKzFTHfVKUkUZX2wt+xSw9t0FLxapYzzZUdzTRZ8KfoiAmDAzY5
8TfOPCSPYWPuoeRIKbckMbXfE52Rze2sA6qGLuecxKABo5v3yINVl+M6LNyH7ziDYaQvNgGjOGor
4AQYTFCDQaVyR5TesZBAetvH/4vb2BN/Qogn1WN3bGsjSrGOojxhqX/n3pRiEDkLcrGyDGo4RxJu
ahOh3SJZd8z/sEoHiRRQQRqw8kSRGBCD/qe7WzzPFDg5ycsHZKMGH1iWptG7WM/ZZM/GskfToOsW
fQOp3gNhkViP4UnWBrJG9X6of/1Y2TMLv/b2Qvk2xYpF/DiH3BehrVc8EdQInNQ3ONioxFzQBja3
+qiLO90m2mppXemnoKUQQX72LKItkpZmkxBYeYRHn3r0Fs3Ch5vZa4kU5gfxeQunn51cJSmAbdTE
2JiQUqlAFI1xy/3bhKu5na4PnZEj22sNmEumMf/+oQ+NLem9qSMCkKs1mkxRdfMvIluE9ubZYXb5
u7w8cVg7XktUM9LMZoU3NLGzePkf/+CKoO4s6zt/iSGYQRogDfs5sDfjM0cDGuiWygCzMiqPci3y
jfwfpC6LgLxJ7NGH/4B8qaf16QF7moJi6ugqoM7/QV8GN7LsR/24WBe2FqTK+B9noTJ1GoeGnKT4
dlJ48HFIr4dnA6qlUcNwxtuYPAyCtswnsJbngi/2yzisxhU+Ozzt3IHsCyr9DWEmZ5T5icRQYUB/
fuOaJ8aSxulShpur7cep6wqQpIbY523DTtc5e82ouGn3Wu4O6ozKPWY/xftI5URN2jYW7vcdjCNo
3OTnBrnjx622GZg7wzDO3CA4V3IvPcxaovIPcwkT27vn6Pzgn/W1959MQJI9l2opZJZEYdWbIkT2
kZwSuTq4X5LMML/Q8rU/Cjb8npu7ZkYg9TpxQu3ynGeSHIN3akHM9iHPSLkSXfF38w+S5PeefHBK
Wjx/3Lud7/aHeNGeamxIimwY+ectZmILMI6rSLM10APcnfbbM5nuGj+DDVdCLYAo9O/w92CMfzVA
3GBIXpWij0TzFoglFoQ/gP52SXFJY7THYItrTvDTRpfnpAP5VNoo9le5qHy9AVNcLXZM1bti3PfY
9UsMQay1Mk2/59r1uYgJKRUd8JrwRPlUiN04IeaNrxD8IBe1NbSvCIgLA0NZZ3MRp702Px+boVEt
CuIW+zvXNFK7h0pV5Sez0qQBqvq290dhPL6eup+S09M6OIFuKWyR1ejNsuidCnEijDqMYSrjPvaL
Ezc44SKHqM/rTXfSEp4ZV8njyiKc6udvLx/NeSGJCee+cSzvJt+eM7mvtLDkzI5zIdAdRUlxap9F
Rt965VsdyXHTqSzYkqhhh+PDr3yDY4D5ULVYQMbgLA6qQPHNO4gzmlW+fSXSln4PnyLUQPacoNHM
JQUqCPil/qR3kU/Qrh8397SYAA/Rj27x4yT3g+2/v7zGMKsZdE8BILW8/Z3iqj1osniOfmKJU6E8
OZ1Fv+AeQUuNME7Ivaf2fpd03KeqMUBwoc2cG58SQYWpOLPc7ZwepO/lbuoT++60J57HuD2q5VS0
dcF7eLH9Dl2k2zSZBpsCnYbYwx+TDWqfSmJ1KKiXa5y/KTgfixQbyVyfsHQJ5oa52tY36i5Hzw9G
9SXW1Ra6X0mLCLR1nY4/UgH3PBxs3qnLdNMs6Cxf7AAYnPGz0muf6G/YFe+uYUf+ZLzQckA4EFbR
opMJ9Beg0nbLeD2mKdYRQ+RcWQDK2sEvww+qRGMG22Snhsr7n9Ke7qpxHcOZhay6aFXxEOnbAh7J
mTnuC3IOfjIgZ9pso7jW2wcssgtVbwSkeCXojCePEIX32+kKkIjAiUWiHKPWWDNnVcOooU1TeDfH
dlgG/6YPJHDjXVL37zPZjiZCHu3NEDKNjy2rvySUIICcghPKPyt30H8Cd92mWU29IS22AD33PYtz
2EpO57kDOSYaZjxaCvvxsrhq2CdX2wVH9NQP6pJWtOw6oSpfeuQNzHbeNPdmCc8iyFpigT1/Uo9F
qO3hrZ3ZhAZl5+34ZOlp9pQVfkN2FSuwj3cswhL/jK2bUeesyIFMnn7cwomJjl+I1+KzDEzM9IBT
MfuQD56CSmj8owyqyQzwmCC/qWJ+aYgQFUn8e7RK1S5Ef4GdZHUEgcHTuqaEzyiM2PaFv32AsR8I
R/z7Jug/qPxGCrfs03xE+amEgMRfrPbkc06Jc9dSrWF68+R6TjCJFPU/j8UkRy6SYV162+tEmcEx
3sO8sx92mCVG7usWa1gLM8WcG4C4gpvkAXG/0NF7Wudax4ayynoZrl7YOfe2vwnsJjy6uvcrV0OA
N72FjefkHV26W2u9pr62ZmsxSMiDRzf2PvzHL7Aw4YKxLJQRxazjyJG2FQpj9CmCTHkN0lbTW0wL
/lo76WuziES2fgw8QSkzCXzAUp2sjSLBkV5UqV2JbT7duKf++8p4msqhKzVlQD0xKsoZyAnYN/50
/RRjhTXxZfRpQlXlSkoAokEd+4mNyC5J9rgrqD0DsDnicT8q8/v0juWO5UmNdhf+1IjlGE475Js5
AoLHN02OmB5FAe6T8/OYaIrALJc6/hsM9/OY6YPTogXIpScbABFYnsTtJzuLup0qvXupCS/rvVIZ
g9dUEW34oEUwkIYEeHbuY8UxgoHHIZBHMW8It82FlZhFBBZ18d4ESeT6uU1Wbq0WtDlkGmX/lMZN
GQby9G33/PQM7IsT2xKskbwiamkQO9xGgkgQglIIWRSyCHdr2yvU0W3VkYKV7y+wzze5Pdv7qCsM
GA5m3EuuoFYrCpaEx8aYuImHtU2Y3KTc3RdZLHqCjrpGrnAenVBcWQdzUbqd2BbeNI58nhOmemFo
cTUSUlH9xrQMP+piBY92fiOCM7Zk5nMKv58Fw90QXYhIju2ug3dgqCbFxwXgbBA+gdP7SX0nHtLu
T1Ic2LjJqhedspqLh+G/zbykYpyD7/w0crqdieXp2Et4VAXwhb1kH8RBEI9sR7DSUCIB32Mqu/zK
/9dnnJlZmOPZuitIodg7A3tbZGOeNTPnqCuO0W9zxfHxi0RAXbgbOXijesX8+3joopyPYCLll7FS
nUqxX4wQr2yaXDPammAWCzDMF9661m2hxxtMDjX2s3s5luI2BCF+1tRNp+hB+M/s5q4mM32Uh6d0
r8MS45FtQqS956gI88onLyXQq2WYe8LUDcc2qzqEQkUKELktZHyfv8U1nM7FQ6mA4HdOKoY2dEFC
SgbAkr/c+O33v8A456xefwkE71TUwfajbpp+/KfYn4Wk7N5+iU/KqiXM0dgApMr6b01Ts3XM1d4L
Xc4fEPjsv5zJq050glStzf5DhUfE/LqXsq+qEErWiv064Hbs/cGwCZaCkAKVhFK4zCAiZfRpUHPI
QnCt6Mg0+0MZqcpsrz/UD8kS0IgmYkAEa6JlL2GxinlgPr47OjL50OlTQR5prSj6cdBTRkFi1BBw
BwlQwguqkgsMvHUZqfgSQ86Nuva+1qds7y88tXfBbnpwM3ETt8A1OgXvVZjf8Yz8ZfRYWOYpoBbJ
nyYQInxYKjfc4jrcTbRsZDWdNv2SCE7njXhWovSmR+rfZq/o1BC6G0iHxkELdcb196Mr/KKvzr3R
gcpzp0OSIWj444o9A3oV2H5SN3FX5OqF5LcXaNjFn0QeuFMn1M0oLHtvJOBBoG2t72j0VFgJX6LM
MNCTA15poBgvPb2wZc/aS8brHqrp87N4kcU02tDaeIxk65WDCxTFCNN4rVEMlymyAb4pvykTpMdc
7wIQwiLWxhuWKd+1zGU4WMAKrY+1N3EkeXeRpE93Y4Fn9+F1izHMjFfTboDe9YHoyPS7Cnk3Y/pm
7w/JZKv6TdeZTovtlNfP5LrLjR6ULqfLU6WXd27LlEHZflX/t/DPmN7kQh7xID6AsvRg+crOqQyo
npo8MF1yI1Q278UwruCGyGrbtvMdH/8oftPFcobtoo0KsPZ4F31/dl8ZkP4xo98eRi6dOeE1OYii
fjYKf9G/2dpzfOAUqpQhT6iAujnsApuqeDdazCyAKg+G/8PJLE/xc3u8Ec1Lw7RbIKKOrLdkHbaO
9BF3Q2Y60YWkNXoiysG4ah7j6AnNWn51VA0lVCvNhEoZRdzkbrGp5oTgJYe3ma9dvM0YKfIgLNLg
epY/EffbzDGUmzD30ATN7OL4265sPLDGQOe7pujZmuflDQd/jQ2CwhEvkG/ysIuMenK0PsPUAtNN
3wPIoIGpg4Iq8skApWM3OrqUm5ptUVPKzYFw8ZDnrlAKKoUiKNqwwWprUvkybzIHtlXV3kZ7015Y
DENmOGvD7q8/HMZqZIxgY1GoooFgDWl1v1UlphacwU80hBlYHaKbQa7vAZFGp3oNUXj9/p4k36e6
5ljWvfzHcF2cRXRB6svXuUoeQxSTh3ZRgG4RHs7WqcnvY4TSSk+Wc+sgznzYQZ+3wkbBGWvbVFD8
XLoMZRnUDx5bqq8lmro9xX61faP3vyDbSi48XnC+dgKwfToD/YUgbrCs6NebskNB+h5vfoFOdP2a
2qUvy/Io99jYsU2aMOttW0O50UVsbWF1Z7gsWv9kFsT9cmXwss/svLgRo1eQF9AXvsXbSeHzPgzI
Fr0lENHv4+qEiyJYATCh819CnfRYj3zubS9lxkfkd/A3r5B3evBmVrJxS1UAkF5fgZz16mURc9uk
BhTh5ltMW33AgoeGR7KzrB2a0+yR1Jayu3blUeet3KqW2VlOSNXc+D/qsX8L0kME21cLhlYa8Wn9
pQ64R6p7hrigawysHVRHXZZsS6rcppGlwIqtEyOAKhxz4oan23scI+Jc8GAFq2yExbv+hXRSw6Bh
vxas6Z8x9rAsvpUYRnVR/zMw1S4ExqXRbt3RVqyw11cIyHtNv3lfGRkuB7KM4ji0XPBO4PiIHGxU
4R8KIyqL/GmjZ5W6tEiZOSyA3UD6O/C13/0YriBz9cMGIoXvS64756IynNtjkPNlDYA648UO8V21
a3pe8AOSh+22R+W05w3HV7mCdiHHOE2JqOCc7dNCvn9Kg8S/dSao5pQmc+2FZthGNW/gvMTBMSCe
LiFwzcS2pvIWB3K5nxObSngeix9vpMr5N8MrN9Uan/jjJmlYyNc+OnuZsmajfP5MnCkmNs+OHOV8
Gec52WzBAkeCXTQcgflaMFJFAkdxY5YVc64vn8djc13uVHrsSTRCCxvsZrOS+m5Zf2uym1ZFpIw5
bpizgMRth/JzieHu/EMOmsTo64UTT5aDaqjW1wfVHO5BuXz181YXQWHHv85ZAKhA4FPVxULHx6ES
nzSr4NGNlyXBpY5vyaI4gCkyr8E1vg0S7Io25QCFUCpEOAwFmyzQUGtJ0XDH7jDzJzgpY4+24yC3
6JfxJypWqsRk5e95R2vKko7pDJJ6Q5ICYXDwywRFRdeOY9qxZm9qxSw7qFsJ46Kc9iFvh4EUGXDi
AXs4vbJSigx6fn97P9O0+HffAjJ7OdIOLERGia+zLrSgFPL35iD9zyj9NBfqTlhAZWj10w/k2Rcx
Ny1SfOuZOOj8C8S9E8SpX6c9XTZ2r05v+I91yWQIvoa++BZ+8ea+aLlj1hy9xLS1letAOdYfAKBO
kN9yQMKszVDVJ3U++8c80gU6XRTEMQh2qNW1lAxHDWKQgymnGrxheSve+LBGuyTHOyQb1UZeIBmL
pj7m/gj+cBgRzjzGRFLAMWEte3yZNu+0IChXcE5uTeRJGjpmLBqNfK8jxSo4pJdz7IR0VYf7mkjK
RmU/oYWpQx9gPFrEkndSWai+oE0VMAHOvTK5DidUVsOTocMOhd8OEDAxPmjBMVJLKyXAWT5Ptawv
WlJnsDspE7TnTMb2R81CUVUJ7QoU1dVhI69iwkhpB1SphscEg3+Iwb8qf3TKDEmztPNR4F6+oihW
rUBZTO+vh1DlOMqkqX8/uv4MmvoOvdP9l11J5zrmF5oZGdcxfFXB2DR7zgpTiokexc9y7zYReHOd
uoJnQk9kbBWd+pJKI9gpfl+HAGrOP6Tl4SIweGBWYLmj1WSo+BzKOA2x5v5/hxPkW5fO04NNjtT7
9Eqzc3OF4Q4rnJWxUlzWoU+FByEKTalxS3ZE0WBWYly1/2nz9o2JBm9CRXXNbjR/gRYPuTFhk6/V
Y4zRsTE04QifIHOlU7VWGgAvkhwQsag0MTsZ9Ny9iFxq429khEgNQqiglRt/mn8DDALQEgHY4H+1
o3tgpu8KpMW0vqAVAnxgbRkhRwtdxQJZoEzFDoBV7/66d9dA2QrwEC1oDUONLlyMRg5bcdETr+uj
fJI8m9OozI7dvlZTNcsu3UM7lT/Lijq4ezGuvFpPUGsaWXugjpk0y6hm7k/GR0ZlR/pLj3lZ8A0k
BKdOwABEMmp0beUQi6PZtt25AUfZ/6KgsWpUA3k9OqhHKi85jgKo1Qx5ZN7WMHdwu2cSSx4yKkoa
0oZkOOymOLdk8nkP7AIAwQ6QcR+OH8j/lfTvuFmN5HS+jKO1Zr/BYwsmJov7cDG/w52J0qSsIR6B
YO+sSMifTMpsnLOleYS1Ds1EroCuQeE+toyoB1VUozZqMjCdRdu9+GwJphsom2neBw9NPvaGxGew
fNjYIrsIT8/fSQOl7pawbfR/8EKRcHGgDI1+ZfwgyyvT1a3fgeOL8xziDsEZBIsE9eVktC9fboNt
vvoJUm46yR25sXWA1rvrUGkqf5UlgsuoU3cqzRMyklFXRBKBmbGV8lRjWX0WQw93KrJMBu27sh1c
sKHdQs3FpcjdoACJGB+1NM1S5SpDoEEr3uphhrfzbc55TSQWZysZ+4saQI7wsIiByw4Pijo1UOwB
3bZs6xgaBn7oeZPw8olR47+f3pJ07y3VFbeNGzWTggP4tBpZLjBX7e0mG0XZErwHXot4sDCAd4/k
Hg8trGWKAHqmYxvqym3qMug4xGGrK+0Rz9VHzm2PqcLqxJSSY77gNJakPaSrCH1Pj4GiWAoZUEFY
EvkPscLyx/uccjycYBbF39bgAww8ijPogJTcU7f1r/tj33pgO+Y/7RDQhIaqScLJ+idf40tOMNfI
a+2bgNy+6IAjtrBW8Yfo0Q0lIYWBjtUaRtgOf/bZM1KFihHXYwcX9wkRLN+AVvFElj46hImfx6Y+
IibwbsuiRopQL+if+LO+F4eVsnifqK8h16fEfc6nc2Td0i0r+i1ZXbTYdidoI3hxYanhw7ulysa5
vLYq6So2TPfUB6+OgxfJf46nDqn1BEl1tpICFX7WJIyzCxfkIwYpASKD3+uI7/fa/QsCDg6roFtC
j0myb6mwMmf3VO5+Rk3y37cQOI7vMmNXlGdM8bVgRnKSMKIjjberm8ihtBpU3vqQg+WpPqkpOIfA
Yx09Bsej2DmPKAMi6TV6IwmGlMh2MLDMR9R83LyD71vxUc3glovPKzAdOf5fDF67mtapgUNtqkxv
D8QFEWjuo0Bt+eWyflsyz33I4xYOT4gc2OQqaMQekcZtOte4nNCv/rZYLVREcpQE/ErIQxF3qtwG
DgDFnKG80O6zrYlqhnTBxJtn37uIFgr1Mde9PreLXQTbE66kQa61noofyk3T5yO1EHfYknsdARyz
7cZwF+6sA6IyX5mXl+EthZAHjhioAz2hieLcBqztH61Dci6WcsE1MmYCHyO4Ok4rx0MKtxJBHEUS
8nzed8PcYCLex8MKiLOIDpG14O9yjluXdgqn341oPsDbrOTOYFCypkNxBss12/yE5kb7hnOst8Cs
rZpCK5SADffIAx066rmw5p4t7bmshgajP9iEb5rMjcKDfEDV/I5yOao8YMUPawtFkvwdYL04RPzd
KMZQdBVhZFjMVbXI5U1EefGQhKY1STTxQqcBY9XMiH6KC8z8ISiIPfPqjTSA0GvHY8fEow/ReQuh
7Hfa6uhYY0VgbKeK3kVceohdZyXN/vlH565JZ4/eWAYXDF7b8exmcJs+N/sxQAv/P1gJRxXtR/SU
GH50k6lS1ehKdej2N1+r/Y61xLRczUS1aLoQ0CAmqnffgxOXAfwjzlSv6kRPT0rWXX4DgKEBFxW1
7owVokFrgIgHvsDrg3AqawSYjBT9ArftDGh1WLeVTOafhJDNF95ez6ekw/MKD4DYinFxx4CPblbX
x9HLk3c7JqmPzJvA8pA5PdWzrs/Kf0iG+w3MidK9keWvQwtj8UFZCM3Ss/8ZMcYf8st1oZC6WCIL
aFRx6nxnfj+tahB0K86eSAPTGQCvF0GMfni3B1Buq5acjzxhxi7bPcWP0rUNoMA3pY4G/PqtI1RD
wFkQI48es2O0mYhthBgyVSGEbe7wwC+SOVHNJvaaEvVFwHMUl30PkcFOaJmZ9Nw7jCJVy+BnYtwO
E43uMqGV4+ZtdooKGW3tC3Y03HGmDGtzns3tAI72KMCXBj0BgFmyCiZ5janfWhK9j53509Ow1JJL
NmzZIRYFCkjZCFmSFZRujj4jXH5NXxBcWaccZJElAVHbGNNEElf0R9LO65TMR8mgL9ElSOc8Iqlh
kgAKxxtXgfqBHpkTTEcvgkWmmylgj8v7AcyVll17K4uVNON5qM4U8GJ1oBx4dYoCQINrRq1A7k5z
9yik09MA1KWOxsV798NkH6cHz8sGkPUjSdQIN+vUQShQE4sESwUl3jUU71xiV52JTt4cY30tXqgV
EahS9QapaLJ7EPm/YcAsc6itAj9ZrpaMRUvf6ZkXO0sKZpUUMWx2DXyt7Jz/HZIywB56DQjRfJ48
l4uFVckrA0NgAlQvK3VrdDuo5KnHV+V0fsiKYlNe8iSyJzdKtkumyS3iTrtfAO4A1L+Fa2pktD13
Zli3pSjZYZwqfx0a88vuRcu+pa6A7TLZ9wGAHUVtuKO84jaE0JmYqmaD9s/bv3P8s1SIwe35eMdI
mKGuLCGY0vAzxRjDrX7+wVM0O9r8jtwUWjLTHXy5ODtSYU4EdruwgIagnzpVqFXuu0zPMpTIN8IT
MlASZkrN5iX7s18O+G6lVojzrZSZRFTglIVHBw0VfC5CVU1kyOYHx9ZFJdZ51BLy36y9qLmNp8GP
kQUBuQ/CgPLV8ZKnZHFBEgJZx8vlTXMYQE3mEAXGnatVkRwkT81RcWe2rDUgJ+EmO4xagIsipIzG
Uel4eCp3NcPGmslKNzBIw++LsuHtH3edpi+szGVCgjv6aVO0RqYJXz7cCBklxFRAp2LHprzVzNQp
HHpHk9Hq9yFp4nwdK7BnlUQpWJGvPpnwptizO5keMAAP+uImc/xr3t5kfCo6g84cAA+fP6gSl/Wc
GyfMiFXTHqiGsw6jgt8tgi3/bvsx5INvTcYxygqeOaHOQCKSiE14cLEkJjs6rMJjsMFxiSXinzj8
i1MD3vvF6RhPiCI/LNdWBnmDw0iiDrNh4qnEErMSykGMkxuzVb+qRdVtiqksP8C082mYS/A2M6Jf
jYe2bl1WKIdtCUMcNqbmWc815Mu/6q++w65yDrpTvI/HTMhibFQ8PgmVdmdENPwjp6gRQS2v/SYc
mW7t+xLqPbDGYwBzta/vWnKY5Kj+4zXiSnI0ZSA8l2I8FdVoyujVBwXbk6Zim9HUksJsCdljOXYA
8j4Am19kPE7LPQArRHif888jjuxy49Zo3pu1OVwRx+DypRPl/EBFmjQlnB6aG8DvXLUbSBEvrXhP
F+wSpjG9MgXGavqcyyBVX5Ts59rAu+k9o1ji66pv7N+dFk1GPT+rVLv8SR4cUXcIdJaYOdn2XtzR
bABBucjP8qVEOXT9FbZjcuHTfhFgpZDWwo0F4Lyn3/VWrpJRocxdQFWCh9dLXZDxO2uxorzz52od
QR0uIWslQob49LJqo0geN0YwQ1/Qd7exO1lDXc/Ks+k3W0C3viirin+DIZe2horvlsjopvGbQaP0
Kz+c9YVTuZioYErjXjcyeFb6nXt2Eoe5EtdGU50RAdVsRq4W8SHg//FuvpQptkm89IAHhwxvrJb5
NKP040pRJ+c3kVAuDvmlWL6jRTqp0X8GhRTjemJ+KXYVqsjrOoKvxK91K3HdEXtPc7A2Fb+2lEMz
qjuv2WA1Dg6VEQnW2CaMx9mhEX6zHFXw0FOi1eL1inOOFRrL7UB1lrsKKjw9cG4gMYCTh7AYj9q3
vreoWLP+MQHQVfKLH/wj+YX0GwC7Dr/Oe2Teh+eA5OBVXOGazr6hZGKT7zj9wcv54QcnzmwDZDOS
0VBROR3d5Ar7CS7MnLLEwGR2dUVENa+ziNIZNxjrRm9Vu9Cd768X8oo7KPqkTe/6EIeHfTKSh2wa
A9+XUUOPOwobN0jOpib2bM0q/ZUp2Qzv1DI3ac0Shw8bTFs0OsTf0Hyt33A5fo9Lbc4dk7J77gKP
X81teg4VCJktLcqt8aeie0iKTeQkWwWFgIhOadBuV10fccw4SGOJdlzA5mXYoiw7LLAn1vZt1GP+
BoDAxsYI9bZWCv8k/NB6Dskl1RgXuqQNyhCgVtvXwYzO15ZtEBFTqtk8zmU7WHQvIk9qJ+38wPQx
ImdE73gd7ZXmHeqzT9OAufY3iRirUMaVp1eizEAVzW+7NAjVbHHrNX4GgqlBH1YphvYenPrY0Dyb
Wuk4EAOoaHnBgjuKXSMFSdoZm6PBrNDJlMsz+t+O6h0TsL14LmvJCijcYIsdYXsIIxm8sh7++CZi
0lfOTHIJ+rwdCIymhx3syDgfQ3l0XD5nUGRAWjxiAkBsuCvwqWLsZrIXH9i7lUMWQT5AjtzXmA2x
h0b82qFZ9lyzSCfOtB7lUgr9o2sI5JxjZ/nkfTBEfeIjsV1sT9E2yyNVOwL45DdLss4iUP7SC5Kl
5TZhkSDLE6YC91uHzl/Bx6Mt0PJ6AuXCqMIw/G1db3K8het8O3D4JQFR6DWpx3yfKkM5Q338PTil
AZ6AKwxzo3wGZmGE18/rVYdhGAgFUV+EHZVKiOb6jg7zW7/Ymv3rzWJgf9GEylJs+TT77gaFF5KW
kbh0PzV5Kg/zzIWJ5RZbnQZpT4CBzONExPJGObWzgU878Utb3c+8rYvsavMCehFrz0x4m7v/8Kcg
81jfKKVNQFVMarvSSJxxBlvOWY9gPYpTfL1p9O9NPXy7qpYCJUvbLbqY3wQ+Yp44bO0eqeIM+9xY
F+0aYfmXIcju+Trnt0f4a3++FDvLYm9sfWv+fLOTyahmOoNQzQELGkEs8vmKt+oTRFAlRF51yYM5
DeyMAiVnJV5lU9lcZrQPL6cGuvA3ULdJ+d46rgqfM23BVYxEiCDQSBh98d5zZgaG7xsfsO3Y8B35
igMrV1va/apdH6TgmfQRb/RhIQtUc0nizr40jkboqCMzLmNp/MetXqaxQGvB7B0YL8MJ+71Fv9Zl
xiAfKN9bRRV5y7qGDmWRnvxp1gseIXDPHfQxxR9VIb7gYptcVWwWluic668sRvYgIXFRdRFvxFkB
vKdDskYSPpO+N4p4LjPO5QLTx5q+mlXoqozByROL0VCaBtcsgKAlsG+TFvCAan9K+QTTuVUneM8y
L+a++IPXyxdPx9GSsZRhRW5l9CrsXMWUK91257WUF6jmfl8xUCe/F13sxYsCrJjWr2Xj06OOgyqT
YIxhIazFHXNN8bpa0d26SzODwUamsVMwr5TPWyr3mGWqW0Vj5UlGaAQxaALaH2qedBPETJjZHM4H
/2QXl4+diBhX5F+Rg8aNrQeWMPRWwCwmpN7Zw1+B8Xie01KNXx2YOVTZZdhNNEVIr1ehSxUFkGge
BuQsQPgwISA/FdT3Ja/balIBzVrKw7o9dUWDH8118dEJgPkunwovt1/DmLyRQmAngjtOGaPuV7LE
Upoy+quwUWfuXt4NZJKoZvgLtWJVPidXiizgEM2I0nhoAe/y2ev1s97ihNUucti7QqfocppNML5H
miO5gv+kKmor3CzIj8yLPYzaJeZPyjXEizB0rfqz7rOS9GyO9W2l+N7mW7tV17ROQPragOORWUE3
oee8wmY4Ne64SgQaZs0//nldCmlwLmsBw1WylS5trn/JnWY73mLePiKoU4ccRZA2lGmtQ0grc2dT
rxPU6BMlech2pvDSGbcrN++LPelmr/AbTlF608X58fCTAQtjCZ/IxHCyhvDO9n2fS3tZnCuxcfzK
xXt04PgoSieyHvNU2QAS4E6YqymE3KcU0UmJFAtaTDtan6MWVB3eRjwb7jwTeFxbmoYhOmMAJF0F
kboLZ5CrG8vSr1ZHxn1DGzQtWvLNR8qiC0eSDUoewHHdqmTr5YgZr8C/ECJUv6YQJiEbL87MGJ7E
9onxTH/OHQVn+kNaPwR28Dy5W0Tb1Jki/AmbEGWrBJG/mviEqxAmiOVvSqgzWNO3xeNPd97faTmV
5gFqebFWyZudZlC2SuuPlBbQ+d0x26/APUAXqC5P6o/2NVf6TxKUm3xMqq9UwOIgnLcy7kIDXLwW
vG1IgPmMiyZKLt/kyIbBL8csyrf1ja5c8C0uNbMgcitYnWHRBo3s1EjGU1A5mFeeBGkzoZkqIgT+
PablW9bHe+6T3vWqVZVyoxbmL1k+j/Pzxf8butfwlsUiJfJB0Ju3sEjr5FkXfxyL36nLR4NU884I
4xJSp4GTMMF7I2rbef/sNL2OiNtfp66vILxPAgBExzpNwPNJlpuW2KY4uUWY8BJvl2mdIt9XSRFF
lEmJ2s0G8FyHv/nMvvCe0Lp73LHgoAtt+OQ2+oJKWVyqZ0R6HpodlYMYKpbX4qBERTnlaEiWq124
OKf/aUd3O2NpBympDYhmfBWr68hbKC11ZW7CRjetP3vzJeASDn+sp+4X+OGuoQfJtCRkDvlogmiM
NcgfeVPti2fDdvyGJhWN6pdvFE5ycAe8UNA6RnCCUfYF1GZtyVSA0Puv+dJZ3x6QirEAaQQ70vMb
eFYaPrHx7UME7P2hlzrnaueZ5Y0A0xD5QJ0JIH43WSymu1MBqOoatA5xnQo2WMnrSXA796euMwyT
xz45HCFCLteoXHZkkRNOiE3fzIzHfcnDRM/bmRoctSqQjfI6r94sDyKKE166KApkp2nkA+gZzA4n
2QtNWltH01M2v2viYKgyQ3+LRcL0OAiHX+pvpIi+5tK7ACNnUB5BcLBqlsAqCwMbLBXZi17fMswY
w7tHNwonK6teuR8ur+yO5HQydvlsWBaPK4TMU58vOcpTiJjp3rn3Uoo0cu8JFs9orstGc/CuUi2W
pO5nyLrpXwcmQzZjcUsyfczUSHagbP2EpIiL8S2VO8Aci0t1Cc1WyQRUvkECV+n1TVxDjhbKZdKo
MDA1K99WQx0mR7kv8VOk5MzvpH6sscbfo7SgmwiWcGNOodxdPDHsJZBagRC1yLZ5jOgAUZyviGFC
fSH+zBFUGV/W0ecfE1HLdpFmK0u97PuUt0W5m2TdME5HQh1VBCWkAGZcBMh0m+rPfcS8Xw674qX5
hpNnOUy3+kDMWXB+vJh78grRAc3hFftR+k5ii0MIGk4odznvMbNL6Fo42r3a6UXIkCdbX0mXUQrU
jjkjfMLw8L9gUey1gupTA+UDWrMLsfrOsLf7r6DWl4ZgUxqU43FlTJS13aWiT5SJYMefvZ18DFJv
RvSzFiYxwpMpFDghZDyjMgmSrcUPvA7TSb10m/ZS74u5IhuhqzgB/87cds5SW86q0o3vfON6Zxkc
VS36goDCCe4glim4sqfUTrdcGGSPOGmdZXhxROa/EiQulAlNNdekM4HgvWDOCJn3IkHppe2MlhhR
vWqVUDz12NdWwnxpG2Csln1Fqd+mWi0noJtNFzkMD85WPDd00CSpv+ivrJLhS1JCoPPDb3zhMEni
QjIwLlukzz+ngFTIH7slZMpF1w3cc2h6V789Z8ZesuKb3ticU7Jhu6rBDD0RzLiRN6OYyfYdZ4s0
qab3Y0kroXQQNPLa0ocYl9DB0WdTQqt4tOE082X1CwFMSYKQZ5GM4lFrSNppIvM611Yrf92BtZb1
7A931xbTczHl9cVZ3O2K2UojOlCxASmUndTxFbZ+qAEP9FRosoYhggEDUsXwzQNZSJXWaNic5NaP
bo4nSt33qb6BF5UmkT6sN8IjYpmNcAsXnb6ZgMB7SvLEqcnMhBUwHO3yzEdLb1opKTZL7dLsfwTl
0Ze83/67PD/lrjJZevW1oo1Q9UJlDBBM0W1zsH+HRgTaC28G8jZp3YK1ScazBxxxr0PEDmfIEu7X
oJYmm/eQHBhXfvwqQ45HLQWMig5r/rnWBIMi2oD/LZ5oZ//7i2KuIKSIajo4dRvMAntSNp8hlpIY
yPAFaJZYnSIZIqoywvTJQetV+wPdE4VI+ShzQEt9oUNWvAZYP/ARXb4IoK47KFmaBcFIXcGRDWIH
uOBRYK8TKL+GKMnzMPl7hyFmxOKvSQiNOv9GfK8JTq2/AxBRNRKzODVAFl1qWo73nvfE8pMqdw7u
YtNRoqQ8XbiMtnL/UxuEh+0SLoyFyHYaTTdZRRBCF6C1CXdUpxldTWEJPBEY+o9Wnl1QEr6B7hjj
w1dz7ajIAeVYO+rx0G0Dhymc82MR6DEv88qZFeluTweg2Q/EvxHpc67GZ5bCaNNzfcPedoVJhJhF
RYj6FWBba0LDGtTjmWSb6dTJ7MmKr2YHOzH2IxXkk7SncsfAerqMLaWjzj7DQiVE6f/iEz6vWu++
WQdluBTy1k21s9EJ9SMw3eB+2B+n9SOazs1TR+DyK33GfQblDscXuLziUpInGHVcqr8nIusWbVds
EmSfADwEk2ZY5zOB0TX0KLdXXfq4Kp1vU6seEkjTpbM/KF/TDa/yOnDCEKjhT5A3hd1XDPFVtzp3
S6T0kfS3GAX1MY8fXOru3eZxZEZKG4Pxz21ZW1EJ4d+UyAJxFzM3tszLgONMJ0TrIm+hmupz5/1h
NSlSGgJKIK3V+sC9rD4RryWczyBG2zhxflRv+ARsKHz4wLiCz/8KFPqByzJHf7RsMu4iRDs3kiY+
9QYRP3MZ5hLTh+tXzLSuNJ3GsicsLkXqxsrHnipaY0R9ulxzshDL8EMaqDrz65pqM9BviLdKttjw
oZbc29ZzcC3kos7U4n2F4VrFqpdru+FgMVaNj7URYN05mzfpk2/nOQRAppK/FPYnOficsRwcOnMb
04yg5BIp5HlGcv22JVb5IPHa0coIipHyqo+qiTKeYxMAJ53iNaYz81q0VFS3otJyiLXwYe5xzXAT
Pvh5Pf762LGLdQ4RLeFFlviaemB3NR/tBGXt2ReFXp0Pvr2TOV2Puv0aBDQ+ySqjyxsJMNu2f4qd
aLt/GQogpTp7D1u5OkXMWjvRKvAoWgKVzwbXosxznGXcP4WntVqcY1pJCKnGP38rz/TjKYpSrVX9
C/YjCxr9nZH44MkfaZkY5HHKLR47nn1O83XPRl4X/cLWYCjjMZu/X5cpUN1bW7dpqYNDCShvY3Ci
oWBp9Opkv1UWvRPo5LZuSaXGjR5oXmtIzSfRSwTkt1FtrVeku6dE1VxjeDnuBAddTvq6WnCXT28d
SFS1KgMDofwU1p91Axq24Eg7aTrJ4+jSyRxCuAwuvLkeR8PlgVrIOkM4Nfh37aFp1iFCoO+fyxLl
qI76wM934s90IBccTjR0q4UiL3MFX9B2zxkTZ+XHLnaYzMd6kPPD1KinOoo9HJk2bLq+nU16QdgA
yj8/zJWgNxU4SrWuuDqKnwAk1LpwCw+gXiMKovOYxxukQy3avSEaNi5dQ061fRekqvC2ULNb1GZf
RYSTF3RVcWrAZd+8EdXvEUaItDfrLox6tSFOZ5h8JVKtCyXTbZm2iO8tGVXp+mfLE5yEGL4rEK0x
t9dTNHQb6hqvHOEmaVObSkWpD3P9ku0x8XVY4KM8MR2dxQ/ZsOseYCF8uOn6y5KUZqpngHtRjdvh
X98BCw5gJ9wdUIdpwNOCoFIs4HqTuFLIbnD7MRiGaQPJiHiAGA3DWfziYYWJ/3GbJ+wx8KjtvzC4
Dhpt8Q5jASyWLjaxbnjyuDXr6WjjQfsgaIcoTNhhb+1DLTz5nsfw38kblGEkdlpn+zzhXhAFIGN6
HN/nuKkaUe8tUtAH791+oJ206X6JwddjTbYuiu0lZy/6drSJfR/wGS8KwrYuSK0Xk9UDBOY5ZF5n
xrwlaICqtGwnbO1b1Rde2ZPVU58T7RPnZ5eJ98u/nADOyYNg9/FMMW1H5ELJxdE5Sa6aWRlvI+7y
DzmIYsC+kDHV8TSUb9ChgjyCtXrpHonOi3TWATyDgVQNQgfKYuqFTXwFIn9A5WS5f74DlfbxnktV
D6Um/sJ+5LHkO8DcOrz941e+xPeZzQdXVrnR0WN0GvnYqrYIP/ZUND18W7ha8tAQZoi7+PTqGiuv
fq1WM5xZlNFHRoK57L/+rpDhTDsZrnziNkXwJRyDKvo3en7Kesmm5FQXvQTyGe9tEi0jr1wFMcFK
/Iy3+RXzWBixy7rWLwDe6Z/drWkp2XpJqOlhmsG37l2l++w+I1QsnQGr62qy3zNv+tBssVb3gNjk
XRyUwrQ8A3IYqimCH1+6IMHuQRk7l82MeumV/BAcSbu6auwOsBlf4GyHj8jMh0eJrDWMmhQ5vDAT
TPJIlCYhEbXaicCCCzelXlGPUjuGlGOdfkiQpGO2EHdN3A5WsCvW/w9BE7rzg5DoDo2pebpBNj2c
hF+Ur2S5hQeqnvKAe2b00+5RS/TOX+pydL0ZMI9lWvDDBkhJZIetYfCqhwQAHyHg2GBweJ/R95FE
OOJifvpHU4ldGw32yBN/rxQjcrnhu/2GcYdGQNN7x//18ZvuN5BPSDlQAje+qc7ateKRfPNk6sln
j8daFOEvjCSGPb5qjUUqwF5ZrjMNnjpGWurrpvYwASnQ/HZ6D6+DGDEJK838ut92xV/0I3u16VsO
q9bhPu0ikEisI6L+x7QVtEvNkf9aBkvJ7q+1F6Xi8Bk6U228AMxw7F1iEklsQ6iweIdeWpbKYfsC
Hc2tWUmd/Bw/QiBGLJuYnoxLEse/rI9p2X7KiDbTMY6xpEBtx+GFMAJrqfFlNhUTBVgp/oDitHIx
02Cajihw1IqcPMvWvGG3BPs0E5z/RvQQIye0O+fIBJ7Q/JHGkN65IzSC4gmwZ9l4VLUOTteb+qrM
eFICJDOnus+0wOGoh/tIFC0W15t0Gc1Rv9P/xNWjk2QESVUdNqn/1r6RJVt0EJX0lUzdAB7we/MX
JiN3ZDi3GCXwHdtyNHnMM0eyHsZhmeQKTaChjFVrIT6lY3FyNxrrVFNIOvnom/oYMrZnrCVPMFeu
g8bKm0vmQAqRUxV8xvEPCnVf+SDitXkQkl33V7bsqgc+J44fOJWNfH+GtMZdWkxtoFSWCANckcNm
Skn8en7cyCc6TnyuNuekkVthFsyW0/94mJ6qnlMlgS/IW2Y22aSfGAJr2r+IA/xzAhGL6cEFsVPw
Tiypun72mN0bWECTYHkSQT7xO+ObAte0kiLGR7tECXa7FRP+7iSyX/niZ48FnDYGC8NLm3Rj7QoM
5NE6MXq8CvF1cQzZG3PPz60iraLtkDITGt7AbiOZmTQQfGupFxrDBa3dQhUjrulIXqQt1dNU4ckS
XpPYHSNaDYB8Ezx8zhanAsMw47UHQhN29RJdkeD8nCifuyE83Av65hR66dh29uGmnW11TJsTFShc
+U1rRSRz0NJDd5y46Q7HWy9HHS33renfotVadbTARRGac3WwHAYXsprWpnH65UMhTt+r5u+LlfGb
QW7lwRYOYJGyjdbhE8glU1OpQxnQ3R5Kxz5BzpQOyjtW0ppnUgps+bs5zdG2XX5LRfL5W8ZHLPUo
FHcvboBVayjAKuZAXTPpAEVub7SSNfXO1X5uhSA82Lwf0PDtZcd67WRAOTp2wTFknjJEh+NdjIrW
3riPbLzSlswijV1lpfXlE4KoV3qyHk/qBE81Rf0zjQBq0/AWyIOdQQ5T/AiF2UkdTs6KIFzZeUzr
2TBaYr+r6eZ+Jh4BjLLrWpC5v59r4TATLSFtPASBsImyBQBKm784ScMcx2M5JpxI4hQaHHF5jwE6
y3+BmxblGLxmPp+sccZ/X2KjPQ10w5/DGaJ++7lHs6YyCMwdyrUhngyvIyvuTcMAemQQYentEysh
Q8jB1fUOedLvK3VmzsJUfvh+ymWr0WYxBa0KhIPoqBtvN5HPLCEHm5D6aIy4TaeZH423px702yKl
s1l2vkdLbc960GuBw6Q9BV6euvJGqEK1N+u3JJHSraPRiVcB4MHeQ/s2fqLryQqgC/40IlJHWZS/
crt5hpbnQcgg3Kcd4X+NpL95dbWhhr+Ci9XIi1ang4Q0Z4EPG/7S+Wufi82mKtARLFx6CZ2VBSh7
27pt2C4M4+ltvHNl3WFOve4/YNtY5oivdRghq/A49eZLz30ahrJzbzSQmKZAivYIHxksyIr2/M6u
Zil9hbkAb9BYfMQWsYx7aF/4x3oRCccKeOuiy8nfYRq+BGTdkKTkTt0MmiUzoe0PJ55hCpdwQy94
nL7ZcJ6mLuHiB7wesg2wzVRMOdtBSx70etKoGyBENwORpUbP+J65zHLs74rfYc+Ru5Ux6pHbmffe
esd2Jdy1dPk2VYL0iKt+pB/b4QNByaM9ChA48zbkksPT5JNqKvsF2BJzMS7lRLCrxBWlgQB5PHJD
D/qPCJISgoqdODaJPj3bAtvLrSpAwLjrM7hS8K7oFy1f38fxkAxW587yHghgtHVZ+aqNwpLba1wt
v+eI1Jpk9tzje9XST6QxaPX1wHTk0xypnpG8KZU5dkliTS6UtRzGeopB4oDZ9Vr7zx6xq6jp+swn
d/Ysb/SxlKXIPiQ6dWQeQXwP35SjL3oxycebAu6ebXGgQNspmCWv2jMVLxAsLG1E4fM0IVY6dKsX
XnRmf49Rpr2ZOFXXfh5iDik+ekX/nbc8AfeywQKyHdv0dxA8N7bu6h/ghTKRUvriAPbdUfooDzUQ
9TuYOI6OuMbndg3vqAn1SKtcCiAyXN/DtRmEegJJUmz2euq4aBpA9eZOdZDHx2/aSzS1jlda9zz4
ITsOQTv0RyZmAgHNYdjWyEQ2AlFzDYFtktmyt5mRsCp1ZE8GyR7sUmF8VSFzoXEJRyoT9NBshYHd
30vuPrnEASb5RwE79gtTglNel+S5Y61gLGt0r1p1HPN0wOLHuFKFbQK9Kcn+rz2gwNVEqsJc+uBK
DCo0BWJKd+GJTfdQ/QjuLhkmcoddJdbhvPUyQS0BzDaB7f0pI/TvGG1jMD486ks/YCd7pVU/r/UJ
thNYcW+MOdW0cjjNJ/euPFZruLVUWUXm0SaQYIT6/899YncTyh5Jc/R56/3jbDaX6d55Fpobd7dD
yUYgOyJAYZEJMar2P/BD3ZkJqut+KD+wpOj5dC9BboSiCQiKhA21pAbbSCPamj/FQiKHKua1SYTr
NmLMmvUTBEKw49zpDNcyc5twlbPaOqvSKEOwIGIt6dJ8RtY0eDhhpt8kiA/oeij9W8PbFOEOEN1k
kV1fJuOZibfjo3wwaWUYAuycVGxnqavVjsQsTktMQlz0P1y4xxNXjlCiDHViUde8fpG1DnzqTUFa
1BbT9PyQj2cf+88gdw7Pwq5KkUf5VGs3mb3aKvJmyTRmlpaA64Abs5b+1knySTKVMqGxTQOtc3Y6
gEUhMZudyEQOkDqJaD11IJErW8VSpCBS9TCBCJ18ox0ovtDIOtldJXnsKWtgOk0PZYttV2K4Umi/
+LxYZfYq9WHA7D5S2R2aFjpN2UFWjHEg6Q+t9yEsylZn7z+17OElASusX2DkjK31LnhEIbK+bjzA
KRew9jSdrCEh2cWNByD9z/XR/HjQYCv5tQd1tXm23hwVOEeLuSAYLADjD0Du012jA1sr5A9BNt7l
jRi0zN1/J/TXs8IMMCpy1qNYvTn86/2osE0v5zIJ6sOPfOSGFFk0ajrlyTqwzAIKjUD6Yu9Ml0qF
IT5KVoyB6huXcgO+E1ZK7inyyBICdpTHtGrgcs9UNRWAcAWz3E47t/jExGFVgAA5mi99MiJ2j9Fp
LAZkU8lfAl4uKHJwnUy6xbP10ol8ega2LMCNo1548jIz7i8+0yvVvTQlATJJX5A0wDD5p0URDyJG
KsF/CJuEfS768dkEqN1XPWj5B749stPXB3rBs9P3ARw46y8XlA5dORtNhLCW6aEGRWCj/rOQZRZO
uSezlhadETd00pClxYa/YrJcnF6kOzgG2i0881cFqjF88KRrXUH9TrXTcHHbchY96rPzjNgeLkYn
sqS7vBO20yzm9JwZ+VBf5FGfKhRpATz4yhTjjVWghFEdS9n5uop0ytw+SmBv665tgsUHcXPRYEyV
bUmMitM206eAMfiUkhu6thbcxhyLbBT+wFAxhNRpwgSrax06CN6KQ+o6Cn6sLZ6GVJahcc+oksAZ
34jMjCteLlSqa77BP0B3jrU5qIxfyM5pweKG/I6SYOMNGsIIx/CWIcrCq6a/gqfDfKYi4+W2CeCv
l4ZOo5ueknnrw8SW4vrZa30oF0xWS5TxdPdhl2+PcT1tyQHfF44d3hzrLab3jawi7slBpBDnV4UO
frkOVdbbfxK7kTbRhRERy4wbojIqhlxFk+bypJ9FiHf1HpUFfPqCzyDoqgoAE4xmi4koUhQfKz9R
xrGzUXNKiYDawn6e0OxcXKQuFGIbiBQZ5mU0RpSHDg9gEUo+aWJdsbSPP8eCYZmBdSOrHdHO6p0b
scL3ti6igikTO0CjenQ3zUjRFRwtlZiKl7YOts+oJMdq9Yw2P4Jw3EQmMsW91YyN95A28TJMy23U
e9N3sN1RtZ3HrsnSO6D9ommTojzonACM73kK9LX004Fysru1y8BaALsIxXCz84PKVvJp9bsJ9EPY
MVv7vRhyEBdvWsP9m4KoO6Zmi6rEWK7qKYa3vf0o2cDzeUO+LRdWGZoG6QI5hAtW+oMDOF/vQeKj
3Gfhirw/SZOZBmd0Xk2Zs29ToFxTfEIKUs5+9IOvzsPbD6nw76uxloNAVKKqSDf38NxkCsIVynFt
9C3jt+V8m+i5Ci56VSTy2XsYMPrQEcv/+NisUlaPmAYC3jpOcwqCHQq09OgLQm6ztOMH2YH21uoj
3vJpwxt7IzGeHp43avgYyQZIFsLIKgvhkUE4zj2HLqW42sXICs8968KfT4L57x4NXLBRzdSdpLAF
ZBggCjYZYsuz4IDV1uhZ86sVctAbWbj60HrgtNl0VXKIbsb+FDAb0X2CJlilZCOZVvKDrGoz3Nhs
LXG4n9KmWiH+CEu64ghKWQSJhoqcXO73cLytLc81O5WoywBESrzKpWn3OCMdiAvGtAWEAR8HnV6L
PRsECRaq0iRihRV2XptxFHIfbqyLK+hS9NPqNhEtF6aHiGaGTnwHY32H0Rz88/BD99RF0TJh/Fli
FEVz+YtPDdgndTMkyt6Gs43hNYMp+xok5iJCcaVNyeTlu5HX6EJJGIItdup3wkHJ6dLuAkYIrQJ/
yF4PNis1Xxm2kQBN41vOOnNDr0jyA4CLNzzva4lQKTZDRhwYL2ZLt4iqJAmE5GmEmeP9Qhs1x1wo
v+MlVZkN/VojdQeZgV2JXGwhDKxdDynpZu8lXeM4gy2FFh2cK+r3sjVp3p38PFZkXXf00xCfKSwy
SBPeuY6lxJdfjistH1EtwCH9B6DINjuVmAGXJIFnTUBOhZ5XHUor9i0TcQjI3jvzMfxx4xIaCbFU
KYZgNv0QmBpYMHl7t/gZ5p2Q2LW+putdZnndVeZKt9zCCiC9Y3Yv33Ct0c4Xukh5auBBdW4aX7ij
imLuPIIqvs/S9ArSi6TLSJGfujCgtXY5pNjYnJ5VgoKzy4FRGBY/eBLXDpW74bHdPVXxayyUtFnt
tr8CicuYH9XsR8PGyuW9S/NDcXsCiwQ9ZNt5jnVWjIhHVXWjCyvW3PKlMlUxrScWNXpCi0A5XATM
5UqIMv5bxAsEhYNP9VLxdBqhxbAdwql0Ut/gn/WUfQbw+viru382yMfzwFPtgkmpmV6tH/npHLs1
UUZMA5z2erRl788WGeQuJ4qXR8oqGDL+N1e8DRcoPjuL0Iz6MgA+jqyXPHhrY4Kyt4bobmafkDHm
JP3rHFQIKAzUMVUDR8jF9JVGnACITBPz/gUCjq6M5VWHxf6dgIe6UJ3/ulJb9kA29ws2fmt5Z0D5
ETG8+nLWA6ilf3pA3+30RlsP9X5yIjhssPBBWU3MHB4eSjWfeXmlrB7gC6xUJtjLZAdMBiZYIQ21
xioLsWxgP/fgcHurPUO4ppV56kPm1hZJR6b/9SA20EjMJKkssATT/39gP7x/LKfmM55F0jZ2BI6d
z3pEgDuyzI6vcd+sovj9o60JeZM1C3Lg4H90iVQIvJu94gxFyjyXxsAahObulxCUnPXLBmq2wjcx
NbqGnUcgzlpDP0jqDLr4fFBPHQZzXFA9NrkcWbI4zkwhnx7YKhuOtu6WBKwO0DWb84pMaU1Tmlzp
D3cdGIGW/cq5iUpEibqdmbYnkIt1/3wcG72o+aeGjdkwrt7UOM3bhKAx/S0VPbecgcAGAMuxY2nI
c/0y4vuIKsbrbaeZKo57zi29S33aa0ajJWKMCQys3y1uNpHyVY0ZO0ZeXmnx6PCzSwGfkJYdpbyH
lVbMY6emwqPRv62Vb8+pVtgv2pppY8Qmeqr3lJxgQuK/+PlXGEM56BcNEt1k759aEx6j3euCqxRv
rEvOv//o+K78PC8VJ2beLR4IJ3Kgr+onOG3Zp495Wsw/b6HJHu4jqbkbgF1SeKbnolOHVRuRoJi2
hFqFBj9AAV2d+Z71kHYciWroA9q50mb8KqwHk7r0/MD5uV0lfA5J267jpMzA1wx/DUGYZAadTASE
n0gcZULGzBO0Ld8MzM4hgsq+WY0W0/EiQf8ZOgF8gxPBK5UtgStDtAjX2+Cdi1I0OaDkDJe9cgFJ
Qy15qGvKdSdYCSEafNx5iBWhq6jZgY+4sRyfOrqqFvU8pCLHBvpL6uAOBwvBaNeQT8sSDPMAM4cP
F/5tPZ7cdFDYMM8y/yDgNA4sCfItFSS/UzUFMuz2TlPwfY0I3b7r0xaSNVXrOKUuQS7WZnpcbcxc
W+BdCx1OKSzMdjXF92bsbkgIQ+GC4PvTv65RNNtzXQxAWjs9BmjLeb1RWC34rNQXMHitui7ZvH3j
Q5xLPrkGCvc4AqOqMfdZsqwtD3U+W6odh7Zw9WQ0mBWjq/ibIyP2NCRh0LEHS/r0ZhR08Tb0X0pt
IK6XN5FC0K5wwyHg5hMAMiqXlJapvQ83jZhDOlE6g0iCFi8LjRkNQPDo85CnWJdN35AgkAhfY2cC
JROZR3Sa5sOeyAyVR3+QKlW8bDyHrLuQTJYOV17kfJzj7dgTeQ+ZksOFuyFtv9j3Pk551maapUTW
C9WmNUeOPUWf3E+Mfu1SoBTrfvz24yYHCKoLLaaHBl6a+PuhV9dVaYRQdEQMRWh0iuuF2jHkIIeO
kFJYMFoL6JJO12EJlE+PTeYSw3D8N+0rmf2r7ozN+cEA6WRLhlOCkciBD8GeYKTYnG/xmP0rujqa
eawxs8DL0xpdNwgIUacOsI9qU2kvIiN2Vt+oJpS38SUhMEiU6M58kHPI52thL32AnpA8uIOtDFeR
f0nh4gx17z+aqEP9bX6LaXpzJDhngMNbauHR4bFbbvzKx8V6OPVsL+QUdbgNzA+nPvw2gLjIv8LX
y5WojlzEWyCL4+orh3er1PBoqVKHihgowaIKhKDmeYGuX++pHgsfdsz2F3qs+T0sSUdIiWQAv6L1
UqfUNBoGoG3ghwIxfvjJyaJ2cH/6Q4ub9DqH91C9uqPZa+TAvXoRbK5Chx6agloUf27RjPqLSjCW
NkQiK83yCx8mNEaok/XUUGOD4PPXNOYVk1rJl5MD2nqiG5ASziRf/jPpUgfBeQFuLldgu//aI3zD
W5V1itM2KX41eQwGgtrZ88iahQOBbs6gmfFLOTGeSxuxt34LidEaGkK33ZAlugGEHV0Cz76dtN9M
5IvpvgVHqe46w8k32BWuN0mvQpTVwMCQJBQfepEcV2+k4Uhlo9wYm7//1Rbfanm4iJP3EZnE8YqV
DgQBAE+yX+EMPpNTtWVpdtiTD3Z6ckCH1ZuACtIm9fWtArHyUm5uvkjpn3mPwgJEOHho06FeMbi/
nhzIGS9YAt4uWSMJPYGC1ueD+AsntaBD2J+4KUG/UKZ+PcEYgPPegMExon9UrVuvJ/CQ6RP1bPib
GVOpQyOizMuTbyVgsd19d6xGtOzMGoWPueAq4hF/YYx+DHCj7iED+w8pCE6LetPurMOS6O9Q8vnI
Ns4XXBSebgBfIT8V50kExusufrcbXi7gGf6BnPlx8k39rYRoxnXPSKpO5IcQ/nQ0f6Z+5gZgFD4g
t/okS3aLecW/vJvexaNKZf51wRfLQKEYkwnmU0HivAv4O6TNu8GIx5fQxivQCqb91E1JBZSi+J/I
4fAaqiX4edJIkNQAVmt/yoSh16ahDWIuN3QUriVpazxz+7fEQic1nRFr8v5VUJ7wv8lNEK9Tbcnx
zIQaP508GFJ1bIOvncnildPZLz4TpWZgS4Bq4FdvxButEL61QGmt2gnAcRCO8cGf8ppvhLGBBMwK
rmMVuUADIwIudOlOWdX0nvt2+XOLm1+EkzSoFpYNPCvRF7PglSaugqLbzJfyNcEQK7idIScU+7dN
zSZS1DHTKU1mRxYvhi8PU+AVgE3pW4zEg4BBb2N9pbaBlzaUnn4erJgiGDUHybGvD4trNOUsGuJB
n68+7Uo2mr09JIqfWoThpxUYvatfic9hYeNglMW7EBh44nI35FGkqi9jew9HuostPEtngk8HcyLU
8t45AwgtJPFAl4N7RoL1kRU8QoJ9h0UMIytwNfuqEZMBB7k9OEV6IaoR6RLQPa1bsUE0FCQF/YWF
Gt3LPly5XpXywy5sAqLaKdPDXwgAcJ7CeFw3a0anzYIV+E0QHGsjwFwDeQRoQxGDuF1ATgNIGBMt
4YRwspuBAxJi0oqylOvjkXh3m0RpVUOZ/7PMznJ94CR9+KXm+/AuY+AEKmrIHkOeK+InbCdcXcu6
uEsCNRNc5SKtIOKfTPtW01Zd2XPHBSMArRKtbZ6AwXifK9/Zd2+JS15zHf9cuU4LEv5h2jpUype5
CrNuIpRC+mMEgQBFJtmzLhx3BKQV73zDiTsU5QIHheuzXSad0eKm4wXRchUN/+vJ3Vvfk9dzQ1RJ
HckEKsDg82YY2N2idDmW7YWqoMSaNled6IwKQZGgkf+cj2M5hQ3KARAghND3WSAHyPykShitV4/w
DgoUsXt1TxPLUCnD7N4bdB/l57icIbr+VhLlahvwERVC78Mriqdgxc31LdEgFb0+vVRmqr6/8m6x
lqYx/4dTDQo0ydFvWBgDmAr+koOYMIejgNM3Qrxg5w9urkWiUkgLahGgY4Twqj7+5KNwk5/e4umR
ecyt+elZv4jTgpjOTRGmQ/+v9cSSfECPAXphRXZ7NhtuvXt7WqWTABd02Jfa/fh7d9k+eeM0O04L
qfII5rwEX01pVcwHRIZpizl7uw7805vFK6nWH54vj85LTbmwIHW2v6V3zQWIbb8KmntSszILszm0
xvASKd8SKFW9rEEV4IQHrKrt6nbWZt4hEJW9wZ6g0d8XEaVFpj6KnaLVDhNjTiAJh4kW/DOuUIsL
HTxweB0hilLKBtOfe4SRAXG1qQfsVc/8sQ+FTecuv4Dp+Hr+vDPA5CEpXItInDRecIxWkiffr8vH
NWmCxdxTRImRaeTouVg+aDWV4KIst8s7ED20RqMclGy2XL17HR0smrmbgk7OEAZzhwRVz5fgtnf3
5kvXIrYzlervpEQ75KRacAR3zPJa85wM11yjIKK51EMs4inCzvX8/V7QFN06jjQ2t0+60AbNmG4v
OIlGtlrrWSLVczw+8LZ+m05CvMnQIxoxwmzcAHOxU6L8t7WTxJsH2KaQ4me5BY7Qzqe3SFBRc2i3
zqxwM7o261mrMEhNxl58RKid5a+FQV38Ndmso2SIPwEF9DRYNmjJcaV4zu9M43pg5D674DU7poWy
2xkP5w3fi+FUQobtiofRs7LaLCxZ8GWkavOkM/CUby2EXdWXscR2QI8Xh1POi+SIq49D3x2MMQ8V
qOFDNgvpd2piBFYkJEhfRRM5WCBhJGeFryz29cWp/bQGTxPcPPWCIomvLXZlESyK2SXgcu1XNZNK
ecjvcLWuIkMEpM17T6f6tJ5x9sQITjuvge/MkGEU0BgdK/I5o0bbu8MWbof7g38C86aUE/T+cmRl
xbEDa4Z4r1iCJki8hVL07GI60F7tx3Eac982sniIjsQ24aBGKR1VnEy99Kqp6wiw5cUr92l0Bim1
fSnWZMHZeiqGZFkQYcf0iDUIuGfhaMd2/pRra3XE+IEOEBzbHCAZ1+8abeLoeKUi2T5a2J6rZ7Qj
yBOLd5O7W6nofreEHEEvWgRcHjKx9K9YoUQSr0rOROvOQ7GYimFp0T/YN1MDyO/Bst5bhFP9UwFf
xErynBoFm+3f1xgBnvf7GbGkjHuBKQMi7beiuY/CI83GxEMDTnk7qM11eoM0vD6SHIE3/34gaxkV
VL+IdKDqQ57UlI9B/zIsPVZD0PYt2wejNcJlgdW+E/vAK+atghJQw42W6jyumizGeALmv8t51/Ye
pj6KglTl12TQHAHzphTjgSxrbuelv5R0uOXOzqVoy3K7SvgYKqa0YAjK2wXdWWmG5a0A8U/1A84k
kQUWV7zXp/suoEKKR4JTy0ngGOg2/7rYM+w1HuEsW22GxNg/hOZjeuPJuj6PK1KYLP7yU+jLe9+b
zwouA5zUyHd5XFAUO8IXhOKOkLcIL8+M9kBUNKPOO1ReT1eVTiUnhuz3Mj3iSibNhuZcVP9pI0FD
q66PrKxKuGn2/cvfazqFWs1ShUkL/Ps2U4UsyrJVoJ4Hl3OjXAyrR1cZ0qaNwDMew647H9eldvjH
3fsWOoIncTf6AuGKxrhJGc96jUMe5xUKCRFQGUNR+sABLi9gFxetZpisMxTfx+F8t0qmHjhHQcn1
kFg34IEr9Ny4tcyjoL3bTV7R+neUv4FYFZ9kRG6iLn9jClwHYB0IANbJGslt7lKzAcWhgh+g1h6+
XoWYjkprkHhtTR7VxfKWZE3KOgj1wijsLJDCgbh9Y6tSzxN2pD1DAug27jxrVWw0krPsnJ+c0iel
OMKuMHnuN2wkOCaOQOKMNnPpgMo5ibCZn/3xoeV0BENYjPsEot9pXCW0p0ZKNEJbGV6BbVoDL0n3
d3NfkmFFvFZV2usU3OAon1ylpDzSIQ+Aer7s8GIGYV8oRtF6SZ5YIdjpKsETqk8uWhSmAMCBCt45
jzZB9s+mEROWsscyMJW87EnVvyDZzpnGxz7+29riAyiejN4yguqUUSEtGqTqS3+WS8ICf2Yw4//F
M/b3A5PGfvX3gbulcjvWIfsXBeIm8e/pUMyMOipkyvgmHgS4GPIcJLDEsHsUj7C8rTyQhiIvq1WF
h4nbd4hyuXFQPYL3B6jnrSHhSCSetsmmGyTj69phhuXDw29y3SomNi/ajTwq6Y5Tg9W3XS17/rB0
Dd3rfe9exGfGjp3jDrOSWFESzgSfqr2VpXPzNX906eqN2CQy5j7u/fz75w04nvAaa5JOTJFuBeLw
9xERZZYcPr3MRYquxdECrab8JgrNcT18f0O4k+o+bygXfd4zywn51Z2FOrzeXCxl1kPP6kpdVHiS
hs6qIXmEpRYwhwdawFbqkaiVPYncrAExHqq6jnNiKl9NSXmtnORFRyA1/vuoAfXUIIc7InqmBFbk
R0Wh61eApCwcBtP/SQ6lkzPG+xl1ZPZMMKqkiT/Rs7w6EIgr5pj0+ebkzDHgBkHmMOi6ECitl9yl
95WOKJ7yxP+dz145auk+1LeH3XACgtFZiMNmjH3vc73+buqy7PsP4nqU9v0KL5ucW1BCY+k19skj
sSoUe5YALLAoVNKdx8/QdZ++FAbPOmcqk5DL9CScVX2nMHENcfmkn04HzvBwO8cYHeYFd+iZsrnl
8RhWHzS3O93aNqczWoSMpJimFj43mSkoKGu+OfPZPuFQKL+mbFC9IZ0xZcHFhEU766PK/X/XzM9x
9yiyM+OEOIGnIRXbT+8jxXo6KT3Jul5DegNV9T4WtNUFbfXCJMyPdr7zoRGThn8AMnN/QX5mH2UH
eAe/+TI5OM0ZsZkbFMe5jKWSwEgZbtVDoJgShmySkGglhszyB5iZJdPwhvNAwGjV1qcN1Pk5X9LX
LkrTQ18Fddp03NpTGKxQqFMjV2EWzdFG38wlPDj0No7FjTVTn1cOVXqVaz+P4fSINjw1YkpF4rIZ
UNjbejfZ4zG/S8BZabd6R+ZXpX5TG+ILEpr1+VeUk/d+V3YLkXZA6KSzeRtEloJoAbdcDql/dU+I
8PxgWNvInfK9hmfybiUX1gWKGgdFUryerpU0fVMLsvGEshGPUlUjRgZuZy9A3cGyZecU67I+5VWI
3FDD2WweyXlV8f/u8IfKbfgtdGWHKTevzXwg504rYlyVH5UuD7HuZQBUpveU+516NBAwXN0fSOBN
G3TUGHmD4V79h+08OS1p9ueyDr+zRnFBxWxdHhefdBGdpy5E2QI94NaXGnTjD7RRwsPSAryLrH2f
cVISeQ2rP7sI9UCtf5dzgS7TTr9r4BLjgEAA2Y7xFp8iznDLVZOalTe1/bq0e8H3nVC6+UUmNVTv
3FAWd1wzBq85LSbgl0RIoFvxt2SOmK7WiP5KDOdY/niowRdzm8okUbAgL0ldiKedVs1kohKU/K32
zkgNVpP3ohiO/Zx30RJF2ar3iowqmNy/ocpAHmqa99Bp7LFOZfhj6I1oHcQZc4R7gc86O9/Di8Z+
pTM7MH0+Yt0HWC1b6fHunxndFiKH6vqSvNSijAZ+V6Q8HrO72vqZ6iOiecmzcI59mGu1TWq230Rj
BoQiJyah5S1tc0t0WmJLZyQ2PXMdwAKSekCLypxyRvvCIiZNHiucbpBL9cJilIlDVPhPYllcPg5W
i1TatXJCnPlj8IIqpA1cnV0HQzmWi1jNrDLya+Spzy4EqbMfKngAjuJx3Svimbq6IHwNBmSYwjQb
+NiXvUMHmgzJBArsANthhCCJGbuPM7UKyrB/bwsM1Wtk2q4Nx6f5i/UMZsVcaUugP5LpzAujc7Vy
llW7aWx9j8QACneBw+AVqYS8InmLG5s4rWMxm2KcmQgi8I2MULLgDCT82QwONVQqY3dyEbv90RxL
V/IM+pdD+v9UHZ3Z+2JlLjad+u6T6KHtCCCR1ztKJ7uRKtxnr/OaZLmu5hezLVllyHQ3w8Uh+eZq
IBQpkHBQmMQCXjYHlAzMMlcOKJRYPW42zGBu0WGodWy53gHDDeqHEi+Xh7Y8XC7t/FzSfxVVk/Vp
+jIUejljkl8qNPVnVJEU0c7FGIYdbHJzXy30VkwLcpoW8Lw+Rqa6ceKGKXDfe6n6xIytHsoTl+AA
CnCzQrAyGRdC79lnBmEvBe8GxW6EgUXXCt3mhGpBsVJoCqj3GR7nDAouV7zJvhWjcGFS7n0QB3TG
UrHW7+g4asjn1Kl9uURPbrA/Eii02BB9WDNyM6Ut+G71pCHT9UstkABXvhFSX8LHdicdhua5VUZM
LicD4HpDvdSUEe07J8DNrYXiQvhJwbYGaMf68R8HXwpZoGLCa7Esf8noqNNBDXULyUVf6i7BPK4z
PmKKniWzKMOsN6v7P45v1O3xNMT3LG5/+I7hM10p5o+jfMLF5EGdh2PPcTEWM239Mv9bK1XVJ6w+
qv5JQKWaLgSvFUlUAqllaDXdF2V/VHjxivdnvhBkONzZJ5uJKO0nBZ9aUhjgYekjtjjEXVogtDdF
y4q3i8m/jXgut4r0/qi46q8MLLkJU5rn7a975OjmYaYtx7E5ckotlEQ66Jxi88xtcoblRWbV3qwT
o86dorx/8yaGYkNYgqqLrwBKgTKsWK1YbzGYlbMjBB9cfSKygC2cMUTyEP9BQhj6tTr5HZrIfKZl
yY/UPsr+cduAjDCuFo8GPbNGKco4y9GH+1WFi1uovIqfs/JpXHurBh8fldiT3o+yI1+XGAieuSFK
qC7p+rcVHx0T3dIlSSnv8ZxsAy35tuusZEcC/byi7muSlksG008KGuGGtXqNavuzGz4JVIZWGUaT
i2rm6O7L5vsYowVTXoHmFK9hJfB9fg1BaV8ireb1VMomx60hF+DHKKsYepqZrTUKpH61iBXJPPUc
/8Hq1mdwMcGwaB8zofbI7dKOzTYDJoDemhRaFdPwl0LEpwN0ZMqx1Elwnwvfnu391S0HN0XMFUWJ
VYyadAiSdnSLWHce/SFZ6RJkQm0azq2TeJCfTpwr5jzOZCMaDWajwxBHgNdPgTYPoMIvDMtuqOyz
tfhvx6cFI6SOLS2jdqaRsJRmcQcoTC5eTf9xZsCeoN1APU4rqUXfc2H8uIIC3cpFXtTG5qnQsgQ/
le+0IqQo3rG8XCVrYKOpX577WbaIAcEdPrn3yIcidTKYJpTVEYCs9VeVNoZktDE4tUMnX0pa0IZZ
ZOSaDHMbOeKn9zwSU15NiEf8RpkE8zW1+qU0Nh770q34kT9ufStGToOfGdBUQftA9/rrx2v5I/Wt
fvZW5/BuG3fqNyY3mSNYOn07ube7ptOgs6I/JkDKJoR/n31Q2ipEG+79XuI4GfZqLEy9CFFkN9N8
uQoB4y9DW8lTr20Z9NFNr+1FaH/RhhbDRpxyJbVBc0RjMrS08ljEYok/iHUY/SVbhbGB/TTuTMkz
ikBpeK4vx9QghJsGnfL12A5mMOzrt17tjJJGLR9ObySpaxjd7evxf8kwKcKnsN+EwqAJC3Z+rNZZ
GDSuEHm9AiMBphjCAZMQbFl9vU3immrIDvTl2PftBkMWNBeDnmZ2vt1r93IsPOj35iBivJglheWM
ym/NaI5dHOmorPEMw9+e723MfS3GeIfJMoSml6pYL1lrLa0FBAoj/QM7QUMyEv2h5kUzNts0mGWS
5qPFWy2rNRFBjbY4FhepGfdwYlp9vSKzjA8x7l3Tze+b6+CdpwrrUoLHtqrrLu3/DL2xRmzhyKFP
d8gI5kR9yBt5XsExON6kys8ytrJuiuIhiaUPB0/C6BPJxOsqXtJ8GuB51XwTWjdNiMUIhZPpYiQr
aGLkyT3l1Ts9AfJAqeEVz7oCrWiQ23Ej9MPQFlU+gJDV8818HD8uanxp58d6oRdq0wXC/zA/QtqO
Ra4HbZdIiBnlWU8FqPIIFJ5gRD0OTT3co7xegm4Zu7JAl/L5eD+SlrGOQXunY+H3QLlDCOvFU3k0
Aaqh/T5gQty2vkoz0ftSzuOIwCNvFF3PR9UAHljpYikPOPbZxWkQqiO3xMBVv6D5XO3XEppX639h
vEyh2j2tGooyiT1oiT3SuvF5nOmEo6csbozfcMrQCSOOqr+jJq1uTBLzsu6pec4I0ED+Nb+XZKAX
8UVGUxQLSxzxNoqeS3o4gXKysimXLOFo4+o5q5/WIYXu0Xyb7hvdBTkp6B5alBLqrsP5AQavsBJz
Tw1gxyWtdigmPTOUzwq9NP8cHurbBVv4yxtdW5xus6m1nQq/uCG4Zcb9aHXyWGxO0vf8LaWj9y3M
XqpJ+c/PH5+QK/x0VVHXNj24aXQln09ATXfQ/wm9sRQXpXHOSqwmeL0TZ+3+Q9EO+f8ImOBj8LyL
9YW6xOGm7rr0P6exDl+oE7swEubIXgB5F6V6NbbwZ0HQNoVs8Twt/gkJumhhh3Fnmjt8f23eGZt+
LtktqY486wQKANDKzTXefSGz7RDS5eXd6WFligGNB1yHDvdAaeg1G8wSsM3OKzP9Xir+NCuRl+jT
ByLj3fKqx3YtjSmtuIBehkLUi9dz+R3I0gIziudNnJFPvatI2h2606v6W3jwcgyiQeQzPVxAm+J2
cT4fAmaDgZQjWVSU+YPI4Kn5XrLu9I7CdfxjuD2HcAMFkdv7Ej4pExSr96bItJDCryMeno31L3M5
c/Re8Hy8gQGi7i0A8VXqc/ReZvkcebj2FfQTiYKGqHEwXSm6GW1N6vCFImdVD8MEv57Ym0fAMoIZ
DU4POsjhE9B4QpA9n+Xrn/AEXHf672PdXOQb7/JAuwXRiVLL0VYqLUWRTdYkaFA0KlxP0jpry0ZA
46Ef4HC2izf61859gCumlavXm0vXKPUFgmF5hAb5zYQRz2UvbMKR9gHnlhnpHgS9n3mdM/Z/6dsR
6UZcYxpFLzk6zk6MEDtNCx4vWEo6e7FEkwM15kniS4ZAbHKqWI4s5uqra5IqVg1RE7ClRdyym7Zc
0lDSWjyH+9bjI5CDWE8UnXFk/LTz5Rd9taEAiXppoKUg10l4gFlp0Lo47UJ67Nhln/ApkSob69CI
k20HRczDDDkudwX7H5edwbw/dgoKdj0VrMhE1af3Z8oOlUP0ZcnbqDita3FNX3pkL2zcb5mRhiel
2P3+3tHLampnuvb8Lth9jMC7IuI2H6AZydb/jAxHhs5tmbQze/SncnDKuC1RtJFuf1oE6F+ldjdD
NnCSpDkGrUv8rwi8gQQ3t1wbxkfAyli5Pp4i52z4nWMZdIcQ+W+GJN5vb9ucjrS2o9xxIGAGdP3Y
YEpvoYaYsTFN1ZCbHSdyp2QVbFjBBjwrgPxW/t0NaQAMYrjjNpmOS85K6N2lNWS1Yc91X/cHm+O9
ZYFAmfttxO3moQCjsrXgM6BLYUp00HWaNLkwktqCkN2H3F45lJUU/uIdR6qjfi4VE0YYz8UJUyAV
wHVVH2Pf2SIo8zyZ+aqZiJDRQldlGI1AsybHe4DyvekCjJWTvpLelGtSDDXVBNAZAxaWRB0wqRyS
1ERPOGYzkjgjCZVyKq7/d/N0Nivi7Q/hkdnW5gfzmYfwA1gB+iOWRY7/2TUk17DuIljgxF0hbH4z
34O/PAYUuU1uZ3itYF9qRCy8XBqHrU2C0vA9PeQwDkU3oKkRWgNc7v50fNKCTnH2dMIKwGIkhxd+
Aqcg9o8w075AfM4Ke0qw/V1/AzBTV2JyjUyq7QvXxbr8fDtl3Rt64nxetafvZUziAcdXJHJ4knRs
Gq4o7s8yVM2iXoHl24zx1lvU3vVwKKyLLgZ0sJdS2okWok3qrnhs7KI4CAgEmvj65ONbagBYieHH
sLIFHmFv3BscgHFONaUKoM1padHZbBBW4DRKKxGLvhS3OVu8XGBVu2Z+Yesdhp/ESy44KploI+Ff
tpdpJp5mmHIvSBBjyhcmnskWAMYCWqjiaaNA200BawjLiz2blbrMsHO4y165VlPgrE9nXYlPbeu2
TKa9UWaTAYR0ODVFtcpgHCYUeLZmlbUBRPgHAZWoGeovSmjqS4XEjf44Ok3JpeKZ7dPoJkcshEcC
LB0hhAZGf8IXbWBMp5vTsu5+7+bBjw5mIVxQY5KzQR9OnoI0jUDaPLAYxHdNJXJ5V2PygFvCV3eD
lQt4SbErxA8Ex/2B6olfFBfwTSk9sEQFuFcP0oNmoildA9A9neJscL0Aqn/O0wluYZ1Zcu3fuxDa
KjtLPemuwp57mKrNmj+bwFGQGb5ISR34BiyuSQECX7KMRRa1bXTdhNw38uCrefHmbpQ9OBoOeor8
uRn+lRbtSyPYq77wezFZQiSCET1j5zYpbm1Al5rNDmolPaxwqfertNwDKbPUi9Kh+a76IrxEVRYa
smVZ+qbGTm6VBS8xT/+BLAMb0hpCfr87t//DKgIijkre7y3M43L3nhk/yczLlDoe3rttnzxjaA2a
IWnEFnfHLHtKtRgCl7j20QKzCpT4JujNqVvxT97/idWmuBC2CbFyTsY5Z1fpzpnls7ZKCnrxRCCr
PJsPvIMTxkX7ghGekarvZwiaz3mVrsDLHRQcDV5cbVkNcaOejaWf1E9ghY4FlGrpxXQCSRUHzCfL
84GRkfeUHmZJFaCpyIEqRzrTP/F98fUxjAObmPBhQ6l4Npz12AtQ6PiuOXJowrkab8zdHcINUmLQ
5nParXY91n7t7rl8wKtkgxDukEMXJ6uvzXfQSLY2EeV+dQk89pykbKfuHLaSpbQqmg2v8FaOSf6w
VsFgFFf3P6tLuhlbj2sCW0PqFIz2+7fy8ej0nfjvRBVymqQqS37QDm1zNR9Ugvj4rWyMi4KYVLXk
+FJwE/q1rX4NPyYnoli4A/sprbaLhf3apd9KsThwm8JzwzLeCK+eAHFS6+V7S1X2Psnug43T/Sgk
JfKe+W7Fawjs925fXtpaAGbxvJ3S7IQQLyNO9KDuaEdwwOb4gQV70sJ7XxAH8QTSU47x6/JoJNm7
ccO+g9IX/RZ2J7NpRTEQ3uC5SQJHME6NAg9Lr5crgS6dfRIRUauAXa4iNHPURxegYTk7NmlyRL+f
ZO72MsT5+GvCdvNk2AH2EROp12aImpOQ1HJasgeHUirFx1NBno66ZA3cq+8OeKt7UxgdJx0Bxu7e
8aTzQgjp8VYjEYuPHhZG9qqFfQSam6PdLVFAOAhJeL2lVYukFQVaIsD35Q33eObG7QH+Z9EqSLS/
wQvOi0ufPe9ycChwo3xxE255Ug7bHSCKhwr3zHaNtr6TmJgpb7MtSOwoFpo5KsOsalpi2D/mE5d5
RnMgu3kXaHoSX4dR8OZMBwrd3A1fyqGdUfr/o89OopYD5bZfLZSZfbg2n1/Aq+YBsw8EcrpfwLgX
qfBeZMUEt2fpd68dxX8m6KFoaSHaGlZBnfo9TtH/+JtJYLMo6lFYqk2/nk8QItYeeBZOvJX4Qnac
zhoWr2kpQUMIPlbVgwIFTHYvwlettEkI5OhFSZ2ZRx4n/F/JwAGlOhwVmLG3ttjlysfjyX4JByHl
E4h/1iNMXlZl0dmrxjNypi4j1ErAC4E0TMceo5LoG7AyIX5qg/W/te1gdWTOGkMSbfIWCMFX+VNk
8jy1dhz8GR6oNkDMwGxk7jhK8WusWffnsC/wgA2ypyOe9BPNznsXmkQeLXp5co0/jDW5Vp8yUGls
vV40L1TRw2K80OWBUMk6J3wf8qmNGNftYusoeQ6SdgiRwDs1TuxSsK52FiNP4+LkabL2hZuTHPfi
/dORUD+hyic+UFEJBThCxpKxP5AKBT/2Zyh64Kw2Yjg6CB45UzIZvfFPANpgQj3toJOTqgZQejt4
QGh3sgnW2aLHm5a6FNS12Eg5/EdqwUpxTk3XxlDCPWo7bizACScI9Uc9Y9BMLqAeXbYz3lDXAgXQ
4y31MT0Bh7xAR33KQclTvdQPloLGNaH07WvMo7x24BUyEQc440PPYvjzHv5yoqS8Fi7iBYnbhotw
/517BWEnaPhUQutwT1Kdy9ebGqEx0Ce37NzKdDPfnHpMo68l6616mTfCESp3e+LoB+yvuAADeJpL
vU3ms69DMRXSEOpB6CqCQt6HKqPbwOahqLm+ogcKTq6tPphVqfw+FKamt6Zkew+dJ0jPNgTxUoX9
GKQJGSfBK/neYVx/9HcI130Lzt6mgdg/rGB9mrXfy20f1FvbP/mVY5iUh2tGXvC6zTILRMiiZ6IZ
KWIpYqEaF6m2twrQmijhBxPTkIZ6BTp2RmtI/Ktv1WjeZJA63f+nmTficQLv+vGY5j6ZA7pepB0v
ZKOBa1JdOzb5l+lsbdn3TOlMyGNxKvyGb5bE2HSExmw0m2urug1LgEG2a7vigtiYagGrKxDN1OUN
pWtOa+sJcI0lzu4yhtNoeR2mgAGfgnp6hcxcN55tP7eBmcTOPnmecOqqnDwD5UqwYdRXf/wdwbH1
y4Wa+yflcqa8ZdH8DiH2inseBq3tUZ1QfJYnxu9ymh7ZOiAeJv+ysGsAr3IyZfLXQaukdCFN2a1X
uXH09le+mEgTnR9XXlA3P1ZO6LthwhjfJjinD596nByWqeisTn9+fk1v4bso/ghSoCDBExZDQYFe
2Kseh1/Cb9DE3lveXS05rcUhB7t5q8Ciog8hvhF8bXjaFlIi4Ivb1KziXNX0ehKCM1HZvHtweKbT
QKcLK5Y4zwQYxuNMVB9e1s+HcOyCAMeEIWkcmHjp/C5AHVGeb4fzQbXS2/3gzUqXiyXmDAD0nzpQ
Ghl1GnvKcxPUc9OYPHS/pBpbdgcrJ2W5K+7QYHlUZoT6YpYh/1uHtFSxOq6nteR6euPI0u39DYNy
W9eRb4jgbSs1HGJkTvPg86i3sXjG5U2y1Pc/TUjTunn1wFBXiXq2flqB6OiJ32nu3LT1C6lspStI
0fPW1Cnra8mIzltaOy32dXG6dkt294/b5VNx6B3MGlenaf+8sWWOBqoVSKtdtmjaOxwQfSPTkNAq
2RwnCbSjhSMV5x3MWx5xuOMFtr0DdBlqJO9P+AqKP2RFQXw/hSQNbcvnaOE4M00LcnhnT0RW+BiR
yrI87+luzgB20lYSzKnMYmhBfySathcRrP0CCOfUvql0TJxEa3eAxsWYVQM+1VFxMUO90l1AzfI9
JyI5TGQWX7b+wJefi/8uyb6HzzI4fjuvZ7I5nsYzZdKSIFtVDRTwv1ulmgmYijNIewc0Ucvvdbab
EwOCvlbIdH33OFAWBduxDuVDrUlbYXea4ZH5YZ9akqqJ7CAj0WZH1C+SjRz9dDQgiIjwJNg8wDlv
ApSunACVWWYich/+CFuCoMszL4+wpBBy5ndAuBp6pasuNzeqj/KheHX461M1MXAfjHjP2H8M+Jzz
NTgrBM1/188YyZm1lEvDSKkWSb2PhqyiFggoVpAc1GzpSYqzTkbGbjOsePwFlLfiLN24lj90VmWv
KDVDc0AgnPlIyRhDWV56KLXfzubJgDuoDJ5vJQGV4aB51kLba3Hw/jM2fFjW/dY1+Fif5Sfsn0Jk
Hdm2QLuQhNBZm2mdADhxXNXlw5XlLAC8AalUiOHW0eyJElLMthf3xPwY28wsx8rmVbMku19ETr7u
8spNZv0w481lnzs/8QzoqS1CS1OjX0k4pGOkF5qPzS02NhfNmwxCC+FXQOzRJ3VErbVhKNHZgJ3a
2sb3OkBNQSgtLrHAmAmACxCFrGNjllTK1sQOSx+e+YftqQy+xXux8QZth2j54VdiNtniJGVrkANG
LulPiWWKZ8YcndomIQrwf/Sk6mJM1z1pKzA4yiRB0RQYB+6D81wYf4r7jPL+oaqDpATPvz9i9CQg
XmCO3Ug2HvIWrWaehnQ7gJdWo3K1K5bgRYVAUdLbA5RrFUR+hwuA5e3hq1aLsTAz7pF+LVU46S5q
ZAxhLQUAIbEfTLs6oM9qZwsZUn22jjJa8lWrEbyLwnXnBauG66sKjso0X6kADxe2ujsIepL8aFuj
n9+jrQyJs4cPSN21AUcDq48Etzse4O6dmMHBki+z2u+ZWYdElrLKdErbLVfFSKAwOs+zCiPRhL/c
NRrGktEXw2F/XvSHeMMjrwOdXvvnFK5/XGGSDMi2vwXBtc/GqC4D3FlMYiahi0OA7joHnYianpVr
IJ3wST7jvvGlpWsYOC09rZaTxFJakeux4PsvinzTBXUHvnkn0nt3gh5Z6N3wr4S4UAxL8YkCtYEJ
MyyMYcqOMp1kUK5rp9pm5zkTv/azlTY7maEZ/0K6v/G7kmCltWin/iQ6zBJ+Bboh4PTafuffG9Oz
tC0ggUuvblRRby1tnXwbLmFSNGYbt5rBOvmvS4eBfSB2JP/o21fkhdph7By/4jXKBKSt/gwZBvN4
lHiw99SGC5LPFdo78R3i60rRgaaImwCt87Nc+n4XDEvrlfilRztoaZ9gjZqRUs1k4AIytMnSgUXK
cWwutmZ70anugUpn/qzdJcW8PO2FFOiKFRDpw5CDFnz4HQ3bSjzSqGZ1ypnqQpcRNZLMJ3CT8lgv
xX3yyH2quDdKnwFMkhF3L3nWsQjK6ChBep35oJnzVFo4+KuAKG/euKYIR0SDGZz4UJ+D4HirFpsU
OLNmbwkrm6DtBOHuSOfUq2AHy1vDbye7N70hXFydlvfrkfH9til+K+MMaMWz5cH6o6U8epYSkLt0
sQ4GK5MjGUToy6Ri5Jl/bpwL0D03iAM6V30aeWy/U0j/HZNSSUnslorlMFpOPMe6LtQUDDfVF7Uu
Ud1E0w+APkgi/tsgyXIEpMYTb123rg/WWAaT0x82tgdWHyOFYjzldwGda52VrnZ49BMhQywZEGy2
6TTecGI76i4tALw0ftfxB+G8gHRIKSHSIhiItzk3+cfJvpUD5qEMiyOcQdOfaPhlQuKKzGbKNvVc
5UG4avrWWp/Tobc2QM6mGkTcP8FetMoZCU8JCFii0D7LIeMTv/uKCO/6tI7JnkCxJhTBwwCn5gkl
7knbOUKtMGQnojcuxEt64qs/54ScsoPBdn10CVJtq7wIHhkhStW/C+2TzSkda6CuNAQx8DL3lFja
jjcUUFVMXaj4sC2vtkDhqt3e1mwJr1HsIc1J8KBT/IVCt29mrZtf0n0kMc5bQZZg+oRAv/+8GFOe
/rS263AEu9XQFZmTjD7uyt2025B/5GDF+xI8kMd36/7FpkA9nAUt0sVjiglboP2TXfT6ioPNnrA8
FVoI8WUHdACzi7Zo9LMtev4LAlZOoeubuim2yQ2q74GQ69cNkNiQjS0Woklp6JkjTgwVXz8/ARKK
ELPZtkMJBR1SvCPWo8S24m299iA2XQpUhCoFStRIJtoSK747cp2EVPSNib+wSUFdOoOIhc4GYQhU
IhT73myWLLMPVdGjI4EEMf6WVt+xPVPrMVSkECRE7fssXATa94YEDPTjznwYQv86qfa2pzThR4SB
8/16/NCz4zPPRXXeC063Np0NWtMLiPDo6VCmIv6o0lXHoyVYogQlRq6dNK/nyFtFgAN5fY3aMFh9
tJaNT6E1B8wjpoSIUt4UshBHoZFFkT11w5oyR1RDogu5wdnWKcN/8ge31DdysmS8C+VmvRBMAQY3
KuEmYVyuiakPYa8KufMUUVuOJOYaY7EJWM1d/piFnD0bs1Nhza7M3BONm4YrseOc4Rva4qiqoMVy
QduKdhaug07QFBB8wRRMLO7FN4XyZ1zovxiI6h36I92CrqLr9UNsTZUpLRo7vAx4L07GEjmi4wZb
PA5o1jnijldyIAxP+unSi91YUm7EBsbi2kKNifA2FASofRVCJDFloFJrXuZLxwVjQIMONyxjjnd0
d3NKiJkpbJdz1b2uHvPiiOcZtbzh/zPlbyLahnnVcCTSgzsO8z6w2z1I7xwu/+cnEwh3MIBEdCoj
7HCOuk8V2HhJ6kimPBW+fDQBjs+1nNVEQN/dIuDaCy5cFt/p9qEBycA+E9flRbFEuK/1SG7BiNzO
dRg1Fvu2jNZ5oNsTathk57WovmXFXP6HBKQO6KXsJ9KQrP1XZJ1detNlnwpaFcxPkQH0GPw+XM72
QF4nEQm3P4/74i6amYDRlxEQHDIVNIOfJBz4WnRkIvryglzgK9AC1JBHLUQQceKLJWSx2TzkxLZl
ctvZYxjki1VJjUMAcLx2FSAziU53tabsyHN8Bcz+RiGtGevMxRFAl59ax/bpIlgrHQBiV/CurMH+
ccfH5IAe0Gq/zqJSSyX99eI2DWdNCrztwVMqI0qY6NQj3dkp+lmu4McY03KuPyU2Z25IgByn8/Ir
eKLXS7BW+JPqjHgB5fEGhNIUmdXqOItrgMLKSTF/XSnSw9cGjrsyyXoTt0uoejHutumry+G6tPUe
lVQIyiNS7U0CgcGXd/fD8KF6cfYqyw7AHn+/IbiASnz9HNCycreCoMiRSKaM6mNiSLJTrafBW2kL
PkbcRmmWktyhXJvuT4SnyvpVnq/9KGxC8I02B+y0dVKzWCunogyLt0yYHjjoNF/Qvh9h49ALoQ4t
Q7fCWbLcn39xm0ounnDQU4HDPVjRvtwFWQChFhoVuPhvWVRF8GD73CiUB23p+F0oDFwnn3xxQLJe
38HO9QZCVDu5p/7I0s/IZX5wM74mbgjP9mi9WygNVLH3X8ej0WqfLFgxpLXs595Q0xpoPu4aZwXj
ExWfy/DBvlGoQEyLx/MbKEhvK81fdVQ3fGxPTIBHiOYN2Nf4ysKBL+akkAMFIqFYmLC50gGhCBIW
2NA0PnEKhjpvkFfiMXH8qjVr2YGOV9PgKZbm8ntMQuBBnkFY2NMF9/CXDlu5BmMA1EXIsam5oPSb
QkQo5UmO3t/B/lcM2ooyI0uX18ThT9AUL5tvdvAvK0rJ4h1KSoKBT9LhMvMjcM3k8O6R9oak0/rC
zKlGPAbX/ogEKsWirw4HQMj2SA9AEKD/RBdujIWacdALI/+aSuZ0imhbLhNW4N1oKqmCIhSEW59g
MUXIIFvQ/iFWDe5xVFJIfBAq1wUNNF4G/0CRB22rK48r69LBGQvmyHS19Uq72aqPdUL1GBcNPWAc
H67Rfuq+2TOOhsRAZ9eOZizvs2yjTomZO86OeW8XwS4DG8ge4QVbEBy5IKOgZMae4EBjs1itSzcW
xL6+bMaHPlPy4kJlaA5lSOOH5mlbmCAvV6WC0A2zSALhg6VpVakRHP6bZnm4LDPzt11jOViN3x7N
QQTIXsUi9U7zoU958qBfpFoHPMSy0u2y/Ia/q7We+h2F7Ez1lJnPHyVoQxJXHLsn0RNYZOkKfhu3
esHtcoaGH9s4FyD99Wo58oHQ3aT7Ke1ZQYFYLkB3+omvc4L2ATjz5r5asZi0bz62NmlWeal7r2bN
xpmrfb5JpuphFCH1lWM1n2GKMx9fFgFkhcUtD/PFKDdgkycvCSwDDk55w7fF21EMZf6BkBSsy2Ri
2dd4+0hvtsC2TBtmyPKnv3TgqhDowfOxcGvjae/eZ4eyy1Sj+sG66cmmV95IZhoMxsi0a9WTBYtV
KbicIWeHqYTFCwdTt2rNrP80mQ6pq1XRN/oTZ26FziQ7fULlr84RzuXH9YPCFtrLRss+hNc4QCgk
u9jYFdki2rK8jCHewx6DUxmGcxCe+R1YZsAZ9lZ9olTCgg3M9ZdvvfBml/FD3a/sHJOrf5V8nu9j
UpQqFR5yyTL2wT5K3Uu4U86EDD9RKRX77Ba/UBd/Y/1/ULCo9ne7KImzDVRAWCIRAIfPhLnI4dTr
9vmnBKUke2LfkiSeUp6e1YZOqw1iuPtCuCivGgXqkHWX8iKITBpbnnJx+L7MN1g7Ts3+Fd5yLeqq
N2BXHh/uYYkzIa1pwVDTzLRBMNq6dMYA3Jf7qOL0NgK2JwyXGKb54MLpSF7LFBLKl5NvRJE6cKXZ
EDCTIrrCGDeHWaIBJuorNPomqLTyPn4jO7n/3xhoVUnq6FocCudaUcNwur7jQ64TYYWdlHjvdvHK
52RBd1pO2KYwnGX1ywV3ESkJGzCx0MNg/0vm6I8vIdRC+u26juB5hagB+IgQcZMeu7ndzv1XS0Sm
MkuWlU9TTgjdkdne7v/mtYHXWp14z/8Eck6hlxJi6B/ra+L6Y4UzIfy2mO1YGMnEgaf5YQf2Doc5
/X6uD2yaQns7Wvk6CCtyIlT7HfHtY2+KrW6bLSYF+hzrOUHw1H5t796znBFF93ufIRy+yh4R7uoz
zafIbult+SzCUuL1Km19jfQQva5C19tXOpk0rvVbQPAmNIuM6loc10vJUYqfA5aDWdx9vxqWC2Gj
vLjaivxB//67uHj4M5SAV34+zxZedxuRnSYDPLAHEwWG5zzRVcDWAmBxuF+zhHBTWDYXvZa0YEjQ
QO09w0uH+S9WKVyvjU6kTXtgkMdTADIGKNol41YQPQsmTENfgo4a38vkPdoL0Cm1v5MI/LfJepC2
/v7CxRDaskmKtf/xDFiEsLkJmUJjo8ksi2TsJ2uDgn0P8fGnZM8/4yS4Fmo/gNfoJC2sCULzumta
7COTv9843vjseNs/gh8GHrtIn1bdiFg2+IAlrsOtuY3sPy4Acp6RHkYl8pUhlJsEOkTRsbZqQx+Y
Y/YWbnfxzgIDUh5fP1DHxTACoVynrlwPjGcOenSGhA3iE96E+h3g/cXaEsN78elgj8FU/sEJm+3y
YPpgpNqj8NQBDYgrNgngd0+qDWr/Xc4Q0H7L6BNGJUKLgSkY57t2reLAzJfT7C9tvU/5H8iulzrx
4ni6LYG7ilf9hFd6aikndil+pU05YBPzlb6mufYsqASFI+1ElJXaMt3da+tp8L6GcipzGLg8t8BS
5970LEO8XC1TY90YzXbAwrMjabX1Wox3GRxRC2mt18qW/4y7EX6dlArKUAHQulKAWbQp7/hmM1yk
rlxeA14Sm8ViIR5AW5Kfplv7embJ3sFNauLFfcm0HASrFm4bgc2j0a6k93tQmYE65uP+OV1qSf2b
zDAQDNm4ha7qvd2IQJYlBOUXi+EX+051hi5/ZESlu2w5chM6EK0zlWBnlxj2BzYr8AjUb86px8Uf
pBvDcxty/Jhi/4JLLJc35TDIobiQCuqIClAF8NmvFy11zDNamER0fw1PhXKjPW5kLm8ASBgzQbXg
vx39bAz0M8SnFLCEKRcQgwt1+knAPfhhEZMqxXmTO9WN/ueqFyyDM8DL59wIXNxh3lpB3vMJME7Y
rX2VNiWGAk7cBGnhJ8u/RzMo8LLhogZNqukhQVACi403LblgSHyN0PQN0hKY9XoCDixXTO08KJCh
zJr3mAH6JruTAurXg5TiHFMPzw0flPRn+MNmr458Me4CVaoeQU4CZyydDGRPB1Bmd4KqGpM+kJUJ
dEJFlB2r52KSIPtayktCM+k3Wt1k4KZn7nlvsyVhr2PuZoob5jrcyQYX+AtqMt71mYM0peNjC6LJ
TaQRF97DoHBD8T/6sjAgux6NCPEAaUI8I4bGjk1dG7N77WhmliplHqUdLivIo5D3jJ+miRrI1GB9
aM3P9GrUvwfyiLt8TdyXpfmavK/vYQye58K4mqMK0mLyQWO4C3Rjhdm05qGkjAnOoCnYgxY3j2TS
7OwjQXhDdnVMcd2x20AdJgp4OA3PHNWJx3ep+a/fEpMtI5XQAbaBgq+Odi8HUCvzJevRce89Rwxa
nnoMXmJBL8CR3+ZqhfGb1SXbo3+F4986pjiHThz8NOer1Goe8DwZjqIRIfaiCe1OIyytigG83LCj
KqXqL3mYaE+uU8F4clzmXo5Tz3clV+lt0Q+DYVhrAnlckI0YtCO/+YcXK9pO/qeLbgyIUhC7SEdt
Yfm7zYTtTLPlkcu13JSOyN9L345csdyZk6xCul2ZWIBL3XbOQBTh0KDmQmWH2R0soAGbsJXrbxun
2siuylfJS+bXVcBTv/xwNolS9BbDu6SRLRA/BsxMHR/zk0C0KMjkXQxWYuGQxOMvhpx6OIC6ejDd
EdWKQ71pP7d/G7olMpuL+gCRHqBC3brrAihpF73NtTuEiLz/cDwFrqIxVvb4fRXVZw/vo9NPAYMO
QsWH6jC1MKEBVVjjYY+SmK+gg4U68tqGd8m7UgRdWnEiVbUd45/2THSD1JRe81fO40Nf5Hji9db4
Vay6yLn+St4J7cyJrPm5wtnB6OrkbLQdpH/0qhJpDIJDfdwKKZejgimuCREezDDzc6OSZ5symd0a
CLhArcZKufDc/SjKMemd37wgbKB9m76dgAuOg9VyN8A12dZQdmlbbo6ZDyfSq41HJ79ze/ftoi88
cka8oReUtngltzhQNWV9nrmX9sUixWj/6eIk3M/QZIodtUHp2A1Nk+CUf2ike36XhWYXw2YvWbAN
LLmL5MOKPWAYT5XvF1UcQm3MO3gQChz/TNJmd5VFQHTmP9fOilTft4z2W9pT1a5hkcR9w2jJTJA2
8edo7nkaD9rkbwJ1LwLoTzBJLlp6juDaaBHuPhh/5PiAuxrQ/mDWDXw7OerSyUqRwLgzqg1Vn9gb
f9naY6cBIKJD1QZjbBzuL+0RMgJi94nWGTFaqpK6SFVsIYbUGjSVPIdL297PjkR4v/dBEmHkYq8z
TbdnMiAlbWz+6EFTecz6EzUaAGY+jpUnyq8rFeVFBJJ0YuNIBdbQ6FkdBLiAMU5xbK2JSmYYK53Y
4eM/Q4f7AwO6urZg3m9dxM1IJkrBLF8r4GgvIe4g+B6Z22TjK07nea5I/keHN6SUKQDiQRtfh/rr
0w0P080nqMu55Q8r828zn7qpyXsaeyokDxKxCMqqmGU/1FJFnIJmZ9OPph+UrWFGChALfes6wLbK
47X2aCkVXczM81lx+Qm5PBatHmy/RBb+m5ttDRnt+Lh9rbWUqfo8mPDQx5phBSYGApiPa7CzYp6m
idZh36+6+fwMsLz9rjCMNwmRGBAmGHGgSe3dlHFCVUzZGO/U6AkbjVATw6bVSKyRz4SrlhBCC+tq
w5aRZFKeUdp6GqoGvusFgSYPmb6ccAS7fj54YhzH9LBdRqHJ88QOj+X6X/wb1ujT5YYstuiMA2JU
ynP3FSIeZ0I/kNXRQZhRQAMoKDGgPxNSzizipJueJLYBcg7e4o+63DP/oa8OC+gEAxzQGnJVgxWG
3z1JrZaSJ3ocxJyCVXZ8Bf6VBg7axBkO1jzIHAzEtmy9wmMMErIqve5gRAs0hHbtf9E5hdtYgwsO
t63erIKEOqnrDqMwPJoZoSOTKxC5HP4XYWt+ue/xI6MIAgXSbdNNrr3lfBzg5DLtgB5kx8fSEPwr
Sq62rloC3tyS/UA1MquT/n3g+lmvdK8eK+lxMRMdPEZWrLyy+694JLXAR9P0HATunASIJdsozbic
UQVEHuNP+hliHcK/GwjBX4/CI+LjthzqubkWb8NmxR9R6vzq3ib7d0a1RmnYX8uzDHr7dNCRYzu8
9xA0MqKr64ltT2EWWmV+LS1sB+4eIojEOdaSeCyANcR8r+f/y9DkRTjZgcC0clHNcDe17NCxvoGi
rPXXE0k5SCFzo3SqtlNvX//LWq28XOQ75XuKhDZT+LQBfbr07xn/k8Ks0W6unu5EzfEntdRzqc1u
kOGrpL488EVzE1ZBH2fAUR74KSfqjQDcnRYIlgcD1I8QS0Lm7/eHIRLN393KACWnTgoOuE8OUY88
otu4LVUBPwxz74mvQtb9gbNkul1I7s3wwBdYWUvWHRbsyHTVC77MVNc+ZLlWAq7YiDFmr0aAXrU8
iBXeT2blDSxmu3MRxjeR+quXHdnTlgca4d+bgzbqJL0Rgq35oV3ps4AxmnGxI0CelZxKzaeLFhFK
t8e0brRVQqyEXUO0hbBZFRTDeoxF5ziyf53+WoW+Yu38R51X+46KyBqLjbdPqtGAEqO0d47dzOYw
1zlrNgr1BKcu6R0aEDAbRanMOglouX7Ew85XamN1iF8+WH79ZhOfQ+rkDvWyho8lKclaXdAUv6pC
dA7LIrEDSG5Ia7ZtbokGDTBLl2GDhZKjSyDQojzxv9EiYhVHakpibo4yqQvPUFMU3opJRdF682Jj
CQfBppCC24cKQvnA1HRlNZZ97D3uTZRv2MgV/aYB4mD2oq5AKIsViPdP/Qt8hzvzJtXE+tPJIap+
zRybwdjbAf4Grtd+DgFCtc0SBn9JOhlFLbX8Nq2rFWjFrOL7DVx8pCEVLcwU4wWKQiP4tDm2hr+J
H44TPchSy0iw3Da9xIpuih6e8JF/yxBWGS4AIzKi1KovnTi6HYo4NJ5mc2mhTWCKwcDQktl7aqU3
JYKR2+TZ2Lk/aDR7q4lscgqM1/YaQ7ugUbWn/jiz/DkvVoe4XJQ5GbSw7UQsIS5sqvq1grN7OAis
wKREeTIZ00lniIkc+gpccECVT8sLjhfG5+2Cwae4uiU1NP2SnJiE3SZmEQc9Z6rmOHvQAN+RVKki
toNHRQY9viQFSHHL50G7gs2zMsNFdwRPkRr/FZHOTsZlusxs4+gYvD7Ko8Dxqh6uamjaUObL6VjJ
lz0Nvi/LQYhJHco200ZwuxXyf3gnHx+SV0MMN5waZgCowURqgAJnqjQj7SuUhvxE+SxpIe51gdb0
eK0k/ASDxL5Zn+Uu8rTxfX1RxBSIoRmEp7EDyv/UnmkAzJ387YHFyiTTh6QmgCHLPGn8y72Wld7b
rYwMwuwelxPjwIQk2Xapgr2hwW9ecgPvhaCJOhdNtBypMSZnXZr1jxjAZcBf6nRS3YWvcOH2F+ji
l8yRR0Li3t2CCX8fWYTYmYqbjIhBsJiOFIG7jUTBEfc+mV4JjE2bqe5rM9w/Smm2FXpeUQ9Bjkz4
bE+XP8m2aaNwf9OsNIK+5x8NQ79bznIAV5+wg2EdOIP3trC7Bv5Z/9Z7MyFeD2UlovHCZfH5wS5L
QQprYVLZHIL/U9e2q7ICjH6LztczGBQWagEtuirk7gF5aQXsgshwshUBeAqVKRDgz4lJbOfqG3QB
6KLUAI1gT+qjltcy7VjluaXnBAv8L70xK0dTBWajZvmW7qRpefhLVyPtXynCH6VDwtnYX1ZOoy8C
sk2j57LnGtcPlp0oF4k8tiggNZgn/91mFLVW3lvcmiVeIvHPyM59TQ2n1LJguSCP2PejuLSTE6KK
gRanQ1tmH/gSJl8lRVUSfNeN/yYftoSCoaOcteGefql44g/YmUJk7cCYhghzXekkY/TbGAGI6RnK
fFphWFyQ2xWhFS1s0f5gcc5+hmeTbijNkq3EpmjCJnAM6SJk9XyE5EKPKjJBmhJwYWT592Ccf95u
Pf5GuBPDFe5qEg6lNT/MH86G28pVmxaR9Hii9GVDvMnHXFq+PTsoQBF8kmMkjTz/1yvbp+oNtk8v
EFgu0kThhYKesVDnhnKH7WlEr1LY8S0jBmS0ChGWEOtfr0ZZlLP4g0fIYeiu8umXv25snGf0U2sC
z9XSYe1+e13o7aDM8Gjy3PVMoEef2azeaj7yhf9vUIWappQgmQOqgWxedAE8He03hZZDtgOA4KQc
LNRX4JyVfFSmG4b4+hl5qbNb+6TtDFReRyl/qJ87dEQtT5Sb+sdMbX43SALUHdXA/GQVT2u4MWHe
3nw4/MENGvPCxtZN9vLoPMvgscqZyZDb7pfjrOYJMmmXybqebIZvvBnGzKWu4gRNSQ4SmPFrP3mb
uqY/zPzFy89eehBCS0Uwea5aLtHYH8NtW6TnYLDZfKs79rAPK0VQ7snFFMxJbM7OT5YLOIT0Bvzb
g9O39GkbXzwfvT7QL4dVqoU+eQI+4pqZA2OCzyuE3zEjeJqJFf5ATl/UE6CWRUhfN8U1+a6Hng2n
JR17bnyM7LT2u2mHmtVc5EGpbHdg+Xeep08Ds+hwk9yihrxL5GzMF/95aJKBEogHlkawR3BvfcHl
R80vWpoe2ENHPcLc68QH8duC10M8mKqv//X5jVbRyvJiqG9kLS1YcQaFprtRAB392Hv2JMiiuD/A
E6tS1um9lev3Q7Nd9ChzKGVl/oBtwJynqwWW2EQKqItlzeV/G46DUx40PUv4m93BqzJVcjNUW7Eu
N/sd9mt1vo9Wo9bULajs1DspgjzKCELqluGmGvCiLMZhzmsAoxnIF0BCLa/IDZWBH2nLqosB5Tz+
E9lfo6oS3lZ9oo9UAJLBlGtgLSaag7T0n0rx0VmCUqu5LiRAxtgnhc/EKwfrQ+MWbHOdfgubaMfX
Br3nekZUb6OqPIa7Lfok1+x6Io7Sv21MZHVfadCZ36xM/aSsR3l0GgM1ptN6q7tT3GYTAtecGM8E
030Jt3ZGec8irahx+pWzpthBAykpJT0/aMkkBbaHsq5Ox8gegbxfvO7giXHOOWeG2T2Yr3MQ6N2U
hW+t35z/av9AWtdNmxh/HMhOvOE4pp860eSiDY+VtP7BOFlesP6+vgneViii2Max5xsMJhFVNGtV
sQpXCsB/XzjpV/ABONTcrpoRMZSLlXIWW7NQq9MNbbLI1kxMfn1c1IDLBu00r7upB4EHk2ZLCxkv
KC4ii/1ZEjHAiQ5VzBfcjmIUNTqQGsVzoujdvudtTWNi0r6CBwvS37/TZLQoMpPcgPIcdPWxoB5h
l+FRGXC0tBacLYIwsZ7CaiaxY1yPPJaav2wfpihXCg4yU0bHJzp9PWTtYAuPOoUIEJxNYdo3+Coe
3oDX1HmjKyQL6I8WQNEbN/Q0n9B/dhYO7BZ7R5Kbllgiv9mzFKaStYWjJ+FyH9f78ILrgti3YHNf
9b5hTHk00oFa0/83xad6ieyemf2l6ceoFGVQiZqLTii9KPq7xGPtPAH40pztz9/B01n0yRvz/88Y
p4SuPkgj6kNBVjwT5FPtD9SlrnE+ZXFD3S5uMrIyCOi6VKlnikEWCjRGbjLcPrEBQGaYEp5rPvbS
vQgjndBgyLq3dsm+ZTv5AXv/wHq3gspdHrsyAtn68iBW3N948240Sl59ojTvCPDSp7rwAGWJS966
IwXJM5udCyIO0u92zEjMKZGsp/y8e765mt7a4nU1R33kUAlS5b8c4ReJbf3pbFBXDuh8XvkTV2fo
FIj9YhcU4KDsBmbU0DQnG1sgRgsM0JxzF6KIrmMNB+9roQpidICyyg8y2eqxnuEe8QnqYyaG+ZAx
lytw9DdOXqvzCIs/fdlFhsKkVEqKgsTJzcT9ssVwJfwOcG+eWmMvd+A2n+VSqNctRK5izqQdkK7t
AYVp6r1dK9nClZcvI/0IJJw/Npdf7uKR1nxQsrE/lMo5zSq5PQZq5lLjOt1AwnOlT5tLMd068wRF
JEKcLHkiMQSVULYwWSRnaqR2jvr+lG8QAU1hD8uu0JQcrbYTwOGdhRN9sdPRlm/AsGiWxjkkt3Fe
ocBxCcCTI8jM9002vQwJzD8nQv8U60xW2Fzq3AGhREY14XM0PvJfK1+Qy2ltLsmgKuJtuZ69qPcf
2wjoYDu4oL68on7yZ7rDkp0ZeGxxc4keVMXH5nsx+FLk3j0G5CXaljhPWrH2zLUDfxjtauGHVbW/
i2v9/NB+6oZvzvWb4jp0tHdKYBlXC47s0wy8+YDPGXQLKhJMDQYOQNnLF8Ld4mz/RwQUF1BrtQlQ
8SfSQolKYszILoza5jfz8g5VyuEvW5I1uU7r8A5ifCBeoej9XMjL5A2E+oH4TcNahUnWczVb6DPI
m3abb+32vbBbAeYWsCxe+VDGwacZ6ciP5NiGNKEeI3wvP6DVTvT74oN1yT4P/zpQ8G8KQnJvmvMz
doqc8RN+e/Ue7W2a6fcax+URSM2wl9yAIXkjYE9QTL5f4864Ai5UIuHXaFCjQgHSIENUM81455ZC
AHh9JrD4JjyYaEqbaAoBfAKqyDNb5aO7uSYs3XXn7byEdYPeECOenK461F6cDHzV6n+RCGUL3Scv
9CQVFGlH2gMBNMFlmEoaRgqnLRIWwkWvb/liPH4j2xJTNE3708hbp0rlYs8r31eoeQOqiO7N9q8j
Mi4fT+IDMncACwU7prp6x4smSxtSzwTM9uwTqU30wtBeK4WeOMC5qmh5v2KNJBGX3+R4b9K7WbsR
WNHvZSljkymYC4Akj1mtazqDhDVwABJYuzkdPWE4qdGe3X6sXkgVfI52Rq8SN1VDtlWcTZPbZg7F
SX4K3x4jt0hvfzYbD1wTMWohdoI9GPTOeurTlTRZjY+x9funF8/uuELVb4WQjIM4tG5TU/Oc+y4r
QosYGaaRCFH3/slZqHmkd8nUACwICHDIJA4a2BWi9hywdimyLMpFuqzLmqpnWGlGajqjVLQcdEum
HaayLMc+d0Lv2tLk34DGRnO6aoNnC+zz5r2xZY9AjI72MXZ8PidX00m2RfD5l/pDiw1dlM7bFwq7
hiD7S2YWLsqzEYqe5H+VOtxqhUW0oJyMoYbUJDE15ZRAMLYYSCTF/d8+9Z2/jUoHYQOsu4I1T8YR
hHg4mjwPurxOyuEOGrgCNOPlrIyqmAz5tiqbrhjEfrWDHvbdXOC7v5n3tNqpaiFdNQh/UpuhGWaR
pMj7Qkz5QFOt7Waoq9H0CeS2astkoKcuO3RXNU3kZ+1blUsUcsicXVTb3fRjhLeqX46XVjdDviHB
2xE3XhS5mv/nnSWEo49EmeON60mQaL+J9TxUzFbamIXotzdxiqEzMm5C15nox6J4+Jc5ZsH+6P10
HCOxvVueAaF9/o93HkiYTc7FmynGxZJNuFU9uBmwspBWc4O9otYgIJ84bcRxRXn37RlKsDE45RkC
8v1xQYS83+aC90SQqzzPP+we5/a8xW/JrsLbQM4rnMsJdzyiYBs+H0eFjRCP13UXxLRbFVmwINlX
XaW7KLIp4ff0IaLngQ00/or5nto/cZAt2lAn30rAqlbgm+Ce+9RdsarxjbFDcZZW1a07s06996OB
OJtCGTJgdEB8FaYoqRZY915K53GsRhymaAlegX8lCVCWlg/xZGnCGtCHdnyHlSromxYMZvJWdfiY
8aHw9yYet3aR0Ia2Jhfk2EqlQ4U6Hj6zsvSf5k9irgXhYBNg8wlTn0kR4YGJrZ6m1+IvQ9Er8hrS
KgDkF2owLjxRWyPWLWckN+URcd6fkCUjgBVyf2xa2vBkr4Gum9q9zz74YmCFGF2r97EPDiJCLEiB
C/mrzuge44HDvRdbIGnAjUdq6VfBZ8s0B7NaSHWZDLMKomcH0yGPqU2DwsKFp3QFJzwV16Zd+bW8
lA4NxiAKmxzNRmcWIipjLCblf902/zWiSM3wRPE3X09vFOReqA83QUuXkOjsXd/Dt/+LGnKF5TVY
T0zZdgD7WHjWivYMHnlZArS9XWEu3WtTTKqJZ1zzriG/fxUCOCRU/+iDTtOEpHZEdFEFkCMlIp5v
Y+tTxu0KabFD05znz0E2j0g0395HVi1ND8PtunDNcEE+BIbIVDrvaOWGdXYQVw/e9bl5qqrb4lm0
YDEwOfjexVQsEn4I1q2qf7KW+nawlBrOSVurYsewXomgL4ezmdi7jDL9dQHxQV7WftKc+c/U703J
nozmOPCIUZVqiba5XVh8AHUxC3AVzAj1kgzX7T2bP6znPOxRYf1+ioE8IN02PPnhDRADAWccCe0z
cY4wF9V2EEJ8cnzl/CxiF5Ay+w+res2ql8tYpVG91vvmtThu/e+5Uas719ekMt6BGT6SCDh/l/M7
pK9WUU5JDGrIy4kwXttXqQKrrAGTnbjofIip+k+oyvLI7DhuzBBhqFd9AZBq15p2y+NAotgeUWEM
dfQn8zsFkEPxL/U7Q7dzS+CF/lhZQeeegUNF/C9TvzEg9bHGPCxQPURkQFeMsZI5zXeIL48BRduX
vWF6Y6kLvwYY2B1BE4tyZPnjp6uxrMfsq6MkCFK7xByqt0t0sBxYwTJ/Xgx+8mGEd4bOVtmMCwpg
DcsSWBiEPNGxfzvrvVKqaJnm99WL5jIOeurqo668McKYrl1iYR4eBAVDZgeYfORqrpa6pFANBRdF
CLxnVD7oL3l0KJomnsNprf8mYp9duOpFU6ODluqPrxaO3zR3Gs7atbu+7aDpo9szopGciiD4fAcp
1Reeth5xmna1mAncHxQ7uTxMTiGVWtdTp9wss+bZ0yKcJkHJWEvuV1JdQE53mdX0zxJ0VmG//Bkz
dogLwdRhBCp7Gs6GEEP7/hqlpBHs10ms8ZASLQjiZP2OGYxVW7axa59ICayzcWWmiUqC5vD463ij
yao2sc3519z7EIyxfWj4xfR4CAmUTTp6RBUeY656dsPLAyby4VFqPC3Fhew1UE3V3aAJRB979eas
/rIE3pgp1OwJtI4qJl06YHs5gfZrMhRcO98byHNGUrY0FKf2/g6nAvxulxMR6haIk3rf5xUIQH8L
c8RxIZdFjjKUZS2AA1juOxbNA5pFQ5WwUAk0LYVvPVUsFzh/pM710Y2+WfZeZuWrXwc1UZWg0PEj
OI0mrSwEEPIYdp2OALYZBoVGzFpS2cmU6dYjW+6+Gq5GT9lKKFDGn6NHn+xLNcQkA5lByRHEQx2U
MiqeQVp+cleJL4c4VaJiD+8NnWsLLsYZxXD2mlE1qwZ91yrmJXlMps4dQdwt/hHHKQQwj+lV+QlA
nnfSH8O5C03ygk8s1OwxlMtiUlA49wYst3Eof81feKlloBYyJUq7dqXJdqeab5nq3/owahh140nY
jELEgWPQgfHfgRFMsm18CFo6bAq289YAX/cn2rIgC2MJxdf1AuDW86w25T7FhCJRC3tJ3Pe2MGzc
xNCV4pAqKG2TcS7poA2xvsq30f4/2Xi8R3i3M5DWZgOmbXo0jH4vdyfWR6qR3ZVxw8a8y9yZCkbp
mRa2h8tCoSYlKtusX2iCtncf9TUiDIzBejXepnPnAyha9fU9/0JqRcBbQ7mCdCy64F5rc7m6Ofm3
q/VH6Ool4CfsvEZtVztfdAlc0RHsPsMz2XSWHhwKef6O1hl0rJe9IK5QlTLXV0EwJlMZSYCJNVs2
eY6REwAJbzj648xzWe+vFBMtBBYhpsBjdWQ7UebtUmQ8X7/lJEZxYMPMYXl4scO/2gXrw585w7Gk
nlnYVGL7rOQAsiAESPI8I/+j9+ecgnl5aXkw4q/iAlw6nO8PznMpWg5pPCBFUc07fbzEf/UfO+0/
byCZxXim2nub6dfF7VtVEMbIPHgLxi2nM+O8jZjgHoVTguUDq5sdRrc8dxrSN/ldle33pXikhijB
EZkMgCgfOVoVt1sz+HYMBvUi4id6qucMilpdIVbdDpE+CEYIMZOiWWheVN8O56UMXpIjB9nm5Gb5
gwJtBIZzDzJhXHm1l06K6bicVjFfxBlU/leoZFyIogAiRPsVoIjN1Wc4yJzvcgcgoDCWls2x003g
/D/MyFQMelQ0gSA2ONeBIeiosFcBmJ0hB7i2IAhazfAbUChtle9pwv+k7KhE9wycIE2Sig3ogl2O
HaHSk0yCMSoTod7ovh7haTyzCN9rn59kNWXqxZxw6K7yA3/fwuhdZMhxXgHyLMr1x3cFMpGo/Tea
19eIDkeQM2GvtK/z+WDMXqYar8cMw/pxlVD1vB/+gtyKb3H8sxcD0+aQx2PdE2QijxO5QQQoiD3z
jH/uMDrpoQbx87PlwPdwvR9RgSE7gUwejL1caP4GwKYSeyhMKnmjRr/6cRMkis8tUiTGR1yez5Fx
cFtfxhWwWgVx6V6Iv/6Wx+J3tqJn0Ctjm7jLGTnn3gmkHPwSjHcd5yWW2Zmt0LUUYAS7+fqL7xnl
Eg87QfnfSP05LMWcIYLJQ3dCtkbW6IbEhVItUfUGlN83jQb/5fcrstK3m+joj8UqkkJkIFx+788p
mRqYRIJrNSNeRVKyHoT41/vCzj2QkW2Vj+Mv+NtLphqLQ5pR7OtoqYZaqI2FEmBcw5E5W5tSlEIE
qgP/YFacYCiSCU19aRDM8fzn12Ynvgh8AJoyZbN4ptPMKE+9+QmjhYlOyaR348ePVu20CEtysR8q
3ls7cyULbKtPM8Mo5rH7dpyq8ZWB1ApskgPJUxUBxbWt4etfAYUou8wETZI8Py1S4VpZ0+AEwU3a
qUQyLXdSQeADFDIsqUjI47VXXYKIIZpJF2xYQ28ujKOVHc387KXk87w8xmeYgpyAfpV0wniU7ZeU
ShyZKzz+mQFXsEsjbVFrcXuP0Ov01wBsU8mx5a5Jdzk/3lGsR6TdGo8GkeKngi83T07kTlxFlrrG
CJU+03BD9wk1KFXSssRS9wnZ3gw12AGWJG6oeODNwDzzI4RVJpWgcgwnSgqQiWBcUnVSkLspapsU
XrqaMZb6neDlJ3UIUxGE9TDuAwd/Is8axvH/a+uFxPbBd0UjRgcdlwaPWJ9Z3l+RUx9gpsRp+uQi
KTNwUEWni5ZoDTv+nn9LOS3IO9cXxHXHbnnKz6LBLqU14FGq2zGfs75ydxcU+vQGRMqCmoHbobFT
5wXjlFu6182yWQ4GobBBMa6t1wcRHshRNeMxXebJMG38OvI68ZhM6BeFk+iBgbIJnaa64uWIew8z
KX9rKkn2j3EuF5CQxBDeiVMfF9gmce87+rArdZtFHzfDsd3J7cyZWSGl4tNR+FlVA3onqtCq3Q4a
fAYbQvElyGmiV1ai/U+bpF45qRb4GdiWsj1AudhLHj+WdA6YYOc0FjEQ4G+ca+lVyqayE33U+3E7
Xi8dvFk1j65xtVdV8XI9Np9FHmOiywbnXXGTwDYgDPrD16hK+Sq8/zRpk1XgH8WtKF16UE4wNzW5
syuVJSJzbLAHZPC5Sf1LMFOnElpTWTzd37nkZKyciELxccXRH0Lp+pvO61XQfgPLrRrHnnWs/iRn
4eTJeSV71Ed4Xn3v7mWLwM27Q2/gVJgsFvYjvpsOg/CJlgh5hCMnaoxPFn1Jv57M+hZKlbt003mg
xBauiwRYzwTlRcTwydXPXx8UQ7sF2v34u7FhjahEh8xHXmiNZ8O9qptZ4WqW2yis059HUTXW2D4/
45xRA/v8POoZc/urGfo9s85dqS3W8vM8SE0PJhBf4POXN3baK3z+E/aA8ADRtfmNiwcXLi9DJtig
RfdTdzAfGu9z0JQcS+io2oeS8XhA466GXm2cinG30ae1e9IyhUvRp69NOawh7PcbT66jvFZ8CQND
jxh8f67M9k0JCHmzxwcS1eMyrI0m03tFrg7EO+zsVyjwUMOpp8HbujWltCILd/fMh88MzleC3uh8
2kBgI3S/tS7bVHIacGLTXPFUs3OUY+c4SBvuYvPoMNrsoOwD50CANRjfUk4eEXI/wnkE8DWkbeqW
JmZTzmdsmJ96Q37Zodrk9k9sAokw242RW18BU/d1YTi4PjaIAn3R+dE57+fFFbXibdrbOGCLaxGn
9elS4bL1fVTh4kNj0o2STAc/4S26eaqz9TAC21WTCbN3K861R8F2/RD+oVpkeOmQ4JSGCxFtrdBG
yXYI5Dt+C7Wr+ldhVuN06YmK9p9CO8CCCN8E/ioAKTeXdTyjvtbSz1yrhPa8thDM8AFeLCoAB5f6
kDZuV+Q8hbE+rX/LEf/AhrIHLZ12Kkqf75sBu4zmPqEKEjtfARgfDQkJv1Z8znpDotwXDN/M/7ik
8J8CmDG1AtUkU8BLno56itDtLDf6QYezyaV8gttBzjZsikVNg3MbVpsH4Gdl+Z8BIgFB9K+KLpmh
HuRbDfpgcfCMXLCfZRzLyfiDO5qtMLRo8eo/bUcXw8INUq/vsGweoxeubVdxoEsC7d3mTgkdmDod
20wmOu05kZxnpGyJ22ArIAJAzA8sjpBWySl0ppaT+6dWWchZtaOMzX79wq+rHGAE/c2T9Pxu9vst
Z1k3dDSja6g7xpFQpzb29sDhRE617iLa2+7NBaAWgOqki4TT4s2xCkdxYPH8zUTp9Vsfh2AhQRlu
1HAIffl5+76K8HCnOHvz8BWYkm+/cv/Jp6ueedM2Hf0oa3/5RkEyigjIN6qDP8pC8ikU/Snb+AcV
LdJiH9XSoK+oFIPHrFoptxEiNcAvPPnXouauwcFk93jZ8aGC8L9SKJZI+uET5ntbroME99EGBpnk
ZaklURMGEMVsEXPiqq9VDGx6alp6lyBAojfOWfm96HkL2h12aM42APJkmpPB5DpY9/l4Uz7Fq5Le
44KsO8dBkbZcodSLEIYlkUm0o2vz5sI0ElfRCjNMjxvl4M9TsdVgL7jJaGRjM+mFWHmvGh+2rlKr
uFlh7SeOC2rGxOLJI8zzgbZkXXByPk53Mmr3v7dykleL78rJpLsCOKm4iu7EsHuOYh11WjCQXwoD
9m8kNG3/Hzmz8qOCD1snrPD4L9VAxLAGlcl9jqAe3ZJdV60Yb1bKThJ84tdoPlYU6CRsqNATnwc2
UKH7Vjy/As4ZgEXsy1hoHa5LYA69+dv/RIpr2cl9eHtjBKztII6mmfegnUJkmglbvbEt4wlc5eyJ
tmTaAB9BUGx32krAOw/uyqZ+I5cNAZLXgrWHthD1hNd5Jc9ba2Rh+of0OY2Dvtf85xT3YUTN1fib
OgeP5SFm7Kg6hYF0ZtWOMnhQ0ihMRd3vBas5X4/dIKqBOufEOSDLPFPbixs1wRfHfaWcGsDohA38
sUbTlXEdrFDGoI5FbsEBGwUftyPq1UYgi/bMSd1xREhu5UbjCY/6Rcvr494AAFlkS2vt1eelw74J
xi3WHhkYuD0drcmGjwwnbnKO8fKfT0cKsBHFuUoSgd8ijf4e9pPQx76QBOZAnYGxpbH25qPxZ/ej
eYRZRZc2zhyyizYzorSOOraa1cQiJmufukafLauuMrVX5ixErbwt3mSNolaoAsC3QnSJiTSxF3Ym
ySnxtV+7Dvqj1Z+HJIwuEeIeVfjaDuAbp/a84CY1ue/4IAK0R6W6v0KQoAOaFkAzste7T7yyAbZ+
pelHxdVzyohPk+XxrQymclM6gV5u1K0cGZ968fIZYuX0I7ijmKsE5rOtQIdvYPrcy+gRVkFNIcd3
4lqoppk26OmgEdGpA5xRZ/42Qd14/5rJJgmDBAy2CYTf26HKTEv2Z+cDdkTARyosLTtSvSARN6Oc
gni80YmMkYutj61vRQ9X+F2PA0QCR0sl2QywLzFoAdUzp7iVy4wBGMBr4DLVlgJOItnT2tAgq9Dq
4E6JjBgOcInbEO4xYLPuVoqxPQbYzwVoTaA078hO00RdXsA+K8i4IOdSH+ewcjsQyz3gIB2OJdke
CGGBMWKVpotx7d3nZKYlu2Whsc0pj2YDTlKlc68FXfKkPjbeKEAz01c19+SvInqzys6WIVqMtN+L
MClvTst6Bxp/cEzwYcKZ95xAql2PKoz1OoE/kBkJ7aWNLSXkqpYkodAcX21Cq+ODLU7W9K7rqibZ
ZyCgDQpuAuhbQW+OMMflFkJRu3kM/VWNhibMLP5Q02UBpOkYxiwrY8K/k8WkqWjNERcV8hHINJSY
Do0Qa+E2x9T2zcBGbgP6dEAOc6RJLtjPl/yLuqbO3sj1SyjKKJKlygZpNQ7mi0BeDZF7PZAlaEs8
6V8H66EB+nZ1CkvUZ6C5AGw27LAnLqPE0vFok/FdgXrVZuwsZA0ZnIYhKHMt7o5Bag33r/fynE2D
QpIefv4N+CTURponzFHDsecCIWs+rChKed46BaI6+5eq3iRHDk3gGtXyamx18CF6RYFTHLdwXJfZ
tILrD7TDObJ9rHhIIdx8qYRYy+pFe9gxTs0B6blJdhbULI7T9LV7mJLoZFMh5mXzn14nT5l2J02n
4Ih7xWix2vVx7hu82H/C3ua/fO9Jfu0uuas0VLuXEUQL2q4DmrhmUPHyHpLhVNC5UvtVKax7low4
COGpuRSxN79NJEvSRkpHUmZv/BR3cUzEyIFHgujlkdA46r3I8u6WLvCX0c2J+lfCzajD1iIoHkSd
he5CTwWjSoBHK0O+/QJrThGznijpYjwO689SfB7Lt0BVVPKXQrS2s0Xx9ky5vSjHhGX5UrUmTrVo
pPcHnTKfgegc2vt1pUrFZp5d5Jpd+K0Tvvtzyo8YYUkYKvq/+T8iJWxN2s68t2W1toFmPy3XNaE2
pELqZbq5ox467vX1aYTT6IGc5iepe/vLy7ILSL6MUIF0ohnICIRocks0CuMuI9J7vTSUPo1ZxiO2
bvqOLkKJwDrrydmG/QJCJqHMt0Oos5FZQtg59Yu8Leozu8UVJlV40JwbXNaxeOByMwBxrWAAR3GC
r2MbrHBotwShNylM7pgUpPIx4dsatHNwcSQbe/syz98mDrGoSqBqejwQPoLuV6djeSKPdy06sPwc
dACTaTF28qYgRROfFPmlUPHgt+GHTz77yif/ixAYqkPqWq2aV5kfboxU5Nfy8inKuguOOtTg+Wlf
pjuIcQGWjo0HhjNon2E7pbROpJb5zd9wiJSHDjAWvUSMp6lhUx5HwsTQO734eDjtH4WRbJsSA4xy
vYzDYQxjc81t9rlSqNstQFdlKNK0FWecMJWj/LNEwme7YTIEtFMzrqIPjj1dOF9EzZm1XN7dyESG
tpo1IzSJMcnnJhhQ3vdAy43aQi5zJl2ysHHJygOfPV4i/PlnEKevFuXMeEjQBB4Td5+/l7XLdTAS
75kyXgm7wcRJHkzf/1t0PAJZ0biR+CfdZtYK4xTmEW4JQy//kWUTz8m91k8uLfaiyR2nCUDtum3P
pZCVBn2v2KnvviN3P+W2LMErnqVkXBjsJyMgSvUu5klGJtvCUuf51KocebFXhiENf93QJiim0vEF
eWo61L7S17bBFY5urUIVuRrBUEyCqp4wNd7IbzIsFasGMeA/rxUGP5+1wNKq3/RPH1ginNcFzjWO
ramNORyyMvgUX+jHpDTzqdypJXjZ1N4Li2Sg2xCZPcK5gxf7tufgKNza7Cn+2Gk2APNeP3OLiGEj
WuL3qPVgO6qVU1i5FtNvGukr1WBuDVoU5N5YrpUNLzAy2Kv8Fb+kojBQ8F6JhVlihiOLNZdVN5ye
TFBH8ftXxzkdOn6F/oy7w3VlxgTM7o5yc8S/mgWJ3yATNdA2E+zonCIklh13MTfBDg2KEWuEAdBh
aWJWRc/GGTcaDXmasdg0XESbFDtVaezlYqfqdfbIyUjGzIHLWkYkFVub39u7VGbCBPAtVS8RYaxQ
DHas7pIxDCKGXhu99y6SuFlI4fupwEZqVOwsLTqs6FH/wboQc7N7gZBEFXuT6ZeLDhsTQQszOFaL
G8KVMuTZ+cWPYtU0fcNWe40PrOoCTIPO/5nT8hi8xDlAC7msXq+w5CJRsyDkyL0DRLMoMtSvA7jX
ExvO49bw9pbsuAzge+3McK9203qVQhOdtWnON3j4Ar8j3IRdl+HIswsQaT5trQ5EfbG4V0+tS6tZ
wfbnt1KnP+B3CUaOUeUJCvECkrL+bhL3OF8zjDEHC7pcvnSjdoHlW7hPKtuKZc04NkTOi5js7I+g
5aWKk7CLutKivjku44xDpfNUpNtkN3CELuK5/jlwO29WhokJ7q3Kbo58jRYlWylUSdEokMjpxX4O
YGMYS4cKNbspSq+WJyoyqymLXX2fF+RCHLAhsIFHghr5qbBHghoCp45Vqw+pmd36YXTnRAoyEHo4
5/aZMGpP3IL+OrsBNIh3al1OTe+ws3LMJnWl8L/45y/e40X3A9Z9isCKHLvCer4ohC5pyx/d7X2J
NdQBzLNHDgvXO3WMURNDlyFwfNxpiHYzKWM+cpCBrs3RZnOKJrKB2Qde+t8NpcRX5DSWCXdqVamS
cc0GS1BeFiQB8N9Xq/CgJiRqEsVMel+7cMfSzlIOFRGsIN83Xp8DgjrUsMMgerZWpruz7i0tE09m
hlxTDf37Pz0aJUKkISWFhptilv1VjlRBqGWSbf+i/nc7z6e3JP2AVfBrP5BHzTPEKNl/HAM8Wu6G
u77iRKc7UW9AgJdSn/XdFzE+9Tz0wpM13pgmzuiS9cjFpwPE5Ip4unto6YIerNkNi/NQqTaPvs/m
WNnUPoVtXlEbTNVAjm9edi5gL3No2eLxO0ulexFCbK97WmNTqACLETWwdlmuEJcT2Hzys4yCBhTd
MnqFBOPr0mBO48JY6jyAty9IUPjhWj5AqQjmKJQ0jzVvWjBFNG60DmtIzhu9u8NCeyYwdtzmxcik
1SUHFdvBN+V9rynlKQJDSr1XxB9zUoN65FEL1kJxsWwWuBj2aC3bZYkWFIyUVUXRhq8q8fbkWvgR
UdpX3wfy1Yv/blZMFBXHAPQ42k/F8QcpjWQihjLNUtJjHw8mddPe4O2u7pBm68f+VTdo1LGT6Eeh
Npo1DLgmOPtjJt1gdecuckWL1cF1kWzrJNbWeUwIR6g5EHhksdBa2Phv13SBkNbBjlzdbF6mCiS5
f7sPZLplPNINvw2CQO7HxFptetDemwmG4sG5ohXNi1AdyVYe0QGlAhbH628V467BmImzlwfQRGCh
4o9WAH+DfxhMt/Lmknl2uP7SvySuiSxbXHiLLJunpdRxGYckV4BF6b8r9uBh5k7ibLa3sWdGxfku
KcTcA+HbFmhBEd8hlCr3Vycb6pPWFQR2ueWp3itKOmKD3XLjZ+0EuCYG2gKauPZASuh31A91soTB
pMNAqP55CSkkS3B9bsnyiAXjuuR8gsPdH+M4jSirJjZPhIrhAcns2oqRdWvp1/+5ligNJHm9nMSg
/rnbBXQLVaRBgUN0/QY8diTFAJmILvQE6f34UHBELoo9TT9ArJTH2xpgZSS28SDBERUp98nNfIzE
p3Nq6cXTfyj1xTLSzxuqM8zKiWwNH4QpdwPgGPfXPtm8lrPl1Y95N5BxzO3Jhc2WedRc+a/UjICQ
ztME37k6lmC1mTJ4OikTV0xNLDbI98CoCPlC/lbpnOT1ncqqqh53Qnu69aSBUvSqpiFFBGu2CJN7
XxsaPg92iHJp74ak50RYw85ZJXrSzmWCdTM798ZMeaFIb/sOlRCE12/iP+ZfIqmyIcy2H2reExKN
1CIQuvmUJwOYGpyV4ezQamxcmUp+abFyzSHDZvDHGEANsBWkOwKY8ENIS9MqfIqCuH4pM0ysysS6
ynb8gGyDkSWDNvwPJC0oYKgzK4Smz48r9zQehWqrtUCgxkREeCTRMktdNxmej1iWdkZbhdHdhkmc
PI6tN/FK8nEWnKk61Tv1DOrSvOiNJRjihATeBSsf0YRGWVUi2lkUGsJ/bMil2yDi3EmQzGQjJa5+
CCikU81a51N32rc3q1z3iKA3OrhYZrz3D4M387AOVDG01nAHlKiZF5a3qqMfew1KDjJSkHmAVkVY
b0M7koHa0r+9VhGvvIh/84Zn6t3uzi2UhsvmROgk4bXawUK7+qQONgsq/UNNMF+5mTdkwywwWszg
0BTECi26OSdwevMZcp5B5zVbDe7cSfDYZmDVW0z1B8uNnkuCU9RICOKZnZlOMYph9+jh5MmYt7tI
BLFTHOvvmdEfJxwbGIsVxHq5kgyv0mFjU6A4y+so8nMlA5atP1Y6ApzYwdva9Ee40sZbGZtCO2+o
7FTyfYVnqYUyMBwisF3iP/ChCbCTzgvlpzhtRJc2VgDIgjcyq3RMf/kwyGfRwfRe+ydiM4csybm5
SO3N53auURS66/Fp9bYASsNvL9WkXtmxpstug7F+jKWptyj/Y5FMleUHMC2pEUpsML3GEZldGbXo
wvSzyqZUs/rh/4JBG/ZpogwWvMnIyKgVbUHgqfDnRjYy9rmUE0mQd3nGiDFbqXAxA4rlR7SlzwFQ
06CrcUCXdXSltMTWKpNCtPJmlprwulkHmO38S5jTYE6pcq/Gv7LVvezDiIs+B5XtmzLte32GIAXq
qrIBUZxj8QyliMun6qV4rOwDuQDl/yBnJLNXQ7OZHXYgTb3hGO+TK5Vo6rNpS1UaofNgT35mrhDR
tOsXm9aQG+i+/hc7mqgYcKpjuWxZNiUs+wUlpTpUBPE76dx9GQzqAYREqaSDd1HwNYC4ut+vRiN8
SjiLkBrexLEGnPv+iqmnLYAomN4Xe6dlzkWugRN3jUkJjzJlNKTD6O3no43hkLuMBBKLn+s2vK16
rWsKvHuwUDftJJbTSP8wLVrp+2ZUjKIJKRwQQU4doPIly8fTl5SeT4z+fsxGQqmRKKP4oahwfFN7
sMyA7eM24xcu1ggz0y/UeYlWSgWZL+g1tMDARNCFXHVzJO599nYqs/0k3kkIeLuwQrj8oVtgEccQ
ZcaTNTfktmnnmGprGOPzI+g5JB1sXBR1LJbjEZaBY78/Wok6trd0MqWyjZISWYkBLOUPtgs+r6On
flIaIvqNFTlYAkkvf/6OuPqqhxkYOGPyvKpxcRouS1L3Xbzu1tGIHKP15rrTltlU9XD5gyPu+abg
zM5fb6ijsMliBR/wDIoJrLPSM0P4zuI8Co4t9X61Nm5uZuGB5oBXzHXs8Q3QuDY5TImr8YdTS4e7
5NGYUgn3DSovjckaZqkptV89Kkx65kMvv7GZcO3gpTbJZzNsiyzQC6esYNjHg2wYwzAK+df6nY4P
UsEM8vbjXb5xAM88pp7xQZQ2EC/5pRR9jIQObZ1RMSmH3+aLbb2z3SZ+gGalzFnhuQgslXpsVXeB
x4dTjZNp2NBVTV2wbHzEccO6xxy4zRQw6+fbtFExw9a9IFv+f2np+rYY6J+HSrnDAZVsCUwxNK6/
h1SkuhuJsqG7RTqSVv72D0oAPGaQNSgsPvKTLSlxURQasYcey9l60/97lzOKvjMZwF6C3vr+FObE
Imap7WdayubvDneI/gcq71vmUyVFHEPiWo4W2iSYybFCBUyGWVeq1eBHh3qWZ7f51JPjAb+ZIia4
Va0aWaU60Olp13GUZ+FUDVUiwXsLYwL6nwdF4VYx7aTBeahlOHZjyszSSEo8N4l+SWMfQvV7w8ID
28MoGzVOEdmKTqS30HZPdlQNuzo48ypFhpSrFnH8zyrcK6D9Z2pKy3kOCtnsV3B6j5CH+lkcGuoC
Y65giuVso5AL/qauGttkB0+Xj9hJyPhGyFZhy1FheBjwGjyNF62Ub+iFGBMhH7JSrfqkJK1GIuU8
nx7y6X1MlI2ZkA/HwtxoPpLfT9DWFZtzVbuTQYvadMBhft+wrZnVTeR3aHE+vw/K6cYOzatoej4K
CBAlCd9ZXddskWRu3zoJk6x7JODI6yhOlXVH4w7+c9O8j8gCsHy5cNMsH/M0XXjqWK0bmsW/Q5bQ
vte14074ln//zo04EgiAWO9D9V0md5Q2wT27yPRJ+o2IbjKl5XlHe9u8V+djU13zeZ4p0rUfOUa5
HZy//vdlyoXM9aIGMn2oiXqFxpHKpC5Y+PLkkmbnKKVOhhnhAFMlCKJtBqtNwIWtLVRcl3J/P+04
Nm8hTGJYFaLH4KIMzDQg1CkjG3VDthqaQl3HuJDJc+eKkqfQ0TOL+lMTDvfbxvT8O5l9vUBp6bBp
llUvKPK9kxcux9d51SFFfmXtLUzwNVSO39C5+evCAmAy7pZqxQwvqh13Tq2q+nUGzNSPXh5rJuF5
s8li+yAk99l8yVc0WQ61Q+LwSe1Hgyt2ZeWAbYYmDnb5YUCcnmwLBIdGwG6BCwc4Tv12ntrPkjuS
KVuVeri3i2CpmPSTcut9+5ogr9MULBlgUcr/JcXAxA87CW2FmZJyX3/ykIV7x9k8jIT2U263Uw/+
qUQHKmZKspVdYUz+FeOeOzn7gNquxCnycphByIqG4FrS8OGH6OCpZKRJtb/KVbL8nDsmMahWU/ts
LrIYcsQicqCspqnVpjo/zWDlwh2KQl0PVu8sJ057lOM03wMGiK4SBZ1YnnBDJ+mQOMjqI2uRASmi
iqhzcyEesNao1W/ZfoiFFzLEX6HugZ82cQL5HJn4xRF8ZSpYUqT+3I/FWIlRyEbhmyVe7wW3tnua
enNT47fmDjSG5BOJLzvZE4cxZfQ3VWmQl9BZ50s/S8dIGWEbMds9XlwS878vR55KdbY1kQW1T1VB
DKQs5O9bDoug1B+L1uFw9S/6WHbc6crVdhS/y8mF517xOa6aLk9MIgbVc3fwwwu/UCVq2k6apc8h
5E026JMy7osGxQjbywKHWluAOIzLCe0KHiLIuN9oPGdxZlstmV6ghMBRTTfioS88oJ1re1xU+NZJ
3CMXHmcnuhUyINpyr0jlUDLHG7oxKoBIvmd+Z8nWZhsJty43Avm4G6267OTyFoMYF5Yoke/J/Aaz
htC4uFA0S082s0VL3YEPUKCUB2ypjpdoWBed6p1AN5+KVtBF689hkmsKadrgSlqvhpI63OcF0EIY
9/R2H2rI8hua1mbMBn20B9uGN5lLKxQq74dzRwn/ATyduT1Dvo9CerC0I49Cc0lHwu6ZwK7WndC3
/3yqlONtg3Pmm7R6po8Nknpret3h4N1L3DfKDDknr5UROUfW2l+WlYNrPh/svPeRr9W0o8o+3aYh
eQ9jY7OR52oJ2dU8XWqjA0C2qkbES0zqLfe85A0RHGWJGA7DjWYqGf9DuYKhOSGr85TdD2rgiOxZ
nQD/SuUv8F9nYxGIgF8KKta4zEMrPhB6pnYk853z4d4CeyjeP6SwulNiYi/fM3I+oE1OJLS5WIv+
HvhdTSwimEL6rFiHh5atzzz1g0pQQxJnaU08biMguoND4Ld9q602F+Pok7dHwJAZ9Ictef9jv76M
PIryuF054JYO+9DMoG0DohYv7dLCrrtmTW8ngMv1cDAsVQYRUKnR0Gu89Hl9g5xRHz/VNRma3NWi
939g4Vw5DsQiylCokr3kgDVt8MkZgFrOMcTxixKlyNs1sZqsczCKlMwNFeH+Oi95j4M9nsa9VGrs
ECN0A6PnNufUpYWENdGc4h/JLX+No4qqmtLNSlpQx24RQqcP12+FKlKVkFcc1eldtBYBEeTv0787
d9c9ZKH+DkUvf4QguqZJe+TFcvKylZ4I1gbXc0B1h7u9M6KPUzjPeFMVLnF/PAq0h5bgIfLGXfLJ
sC9IypQljF4yFzAnbCWR6GktFelIosGi5ItN4wEhj0N+b1nXWZ1hLy5UeM6zQGLVLAYBukoT0A7+
VBN5mqlpqQQi7QC2NF44H0eMG10JB1Gr0ERHffNJZ5QedAGR5+3h9MsGNDs87Tw4A+BX3beVdWKO
VAz/i665cd1KPZi/wvZQwvy7ohHMYqIgO70zPvQgzXEMJFouVNBvHm67Z41r4tyt7rmZyHMPhN0o
/Vm2YxOJQdd2HxVvtpErxO067VOOxQZABCWSngJXkPOTEp7+pponq9yBkz0ugX8s2+MeKoV0PwxR
P8UYvJBtogCj1/S0CD1sO0uxPxyTZA4/Q4IUb60hbeZcGGMdONaHMeZN04MQz/Vsm8Vy7n0hB+YK
hdo6KHC8I8PMUYdA3/jX64x+GMehZa2NjWBWTqHWbcByZ17UHdEsisqrqe1AQvPGxHawbfARyMRG
qrZt8hGs8V7sAvm7QcZ4P4ltk4Gdkvxx/6dAMYtk3Ol9MwRp5vzh7RDRbDI/LUg2xBGzqOntRjmM
khijsJOBnWJUwkQZdqsM6G3pwVk5HoX8TxnuNM/v4gX9mjK7wYSiCwMDrzkSWcTKwPIck5s0x5Rs
vpWAs4p4k+X0mHussX64GtcFIgirAognkE7glVEnU/ViPbUi2nuydG3vpK3hoJTjxtcTllZ5WF9D
zeBh9DHzeseRcNwQAF7IxkKO6OTE93P6wOi0j5ReRLkk3J7/NFH2hVVtSSy/OLnDt0WGUbY8buti
ylBlXkOSzcaDcMW7uNJVpDDnu0OaFBlUsEr/rCsvpEnkcjreSM4jeLp55uzNrHZM2cb/lRHkxgLA
NqUBfX2ss10AGZLlO/yYtAudzjPi8C4BQEX9Ww22C97Ts3Hgp1GRDW+Q7Gjw/b/WSZzy3B9GFvqR
6ylRhVqq0ADQL1sHO9JOCId9kix4rgAS8OXsQ6AVqRZnflqaqG1nFzc1AYVwsl3jpSTm1Wm3HpiD
3sahfivduOwM4JVn9Wi2hBhVwipNUxW6Kgli1oHBMqHLmF3a5u3FCj7yIqcqonyZ78ttA4/q0s1b
2rNHljFQFAepz/pXry6mXFiCYTcz+/MQlXYzJpqZaX9jw+ndxh6DyGGt9w7LUJRaIEQJ2QTP6ycu
RrD7S3Ul0BludpmpUWIDPWw5PcZaSb+bnuM2KhzKMxSMFxRg9vfwKkBp5527kTS8pqdh7jU24iV1
OKiYQxACBkiiF/rGMGQPYULZACY+n9/Kkgn5H6mIrUkthEpsePvKWBqEywusvBU8UZyLUm8R+4t/
tb1r/hgDtJm/v6aT/rHJl+q38tKKbve8/e0Y6Y32o7aRBZUQQ27uLXDHg5P1LHwK+v5oi/hd7oui
idBwuhYCuxwluR5sQjVi4AhcwQfSW1kuKWwp/AgHoJsbCcEr0SnQgyQdrcgPKQfR7lsdLteObuzr
fIckFIt+DEBRcJxo93DQPXTudkyEV64B7DcJ1q1r3eKw2i27h43KOhL0hgltoEpiTjhe65qwPEUn
isSQPow+CupNEutMHrBpSIrXepySWIif4ik4BC9i6svC6pVvBjlWyE1DyHSBJxecu5K2kTSCfrry
Eg8HfgU6yu53OmyyfNWmMBFmXNbhjLpgEqns1oiCNNd8Tq5dOMt7++vRUNm5Y8mF4BUiv1pdNGvc
QZB2r1/baPZ+K6Tb8aQ6bGsPEXep6drJ/nF4MuyhxpplhS0nk26KfScWl0JA4q/hk0dLamW8ClIC
7LFCLU2SDLaKIV59/yCIOyZmqyG5GQKvrgqrVxoj08B1oY5N/NpYMNomJMHo78cmqpxGy831EElY
aZgo8NO6oYsanl7RGV2BWwM/rM9X1e+xcqiubUPtthRXahzhH2eiSdmSNyJuYsc4NfVn5EqUDa/7
APYe5IZtzvvta1+gDKbdcfBiBGAhAPtHLQQhsGaguGH43y/1bPTo0uQFkNJogePWX52O8T6Qwaar
tXrwf+67+x8Fh2vC+BpJ1gjlyOJIuB8b2ZRu1JegrjOV6hFQTcBEUN+//IOMZncI0TgdEC1esV7E
5n5Uz5SvyRNmJXKMuGML3pn2PQ4EHqq+GDgqNSq8sDlWPsnShL9RD/GCFqXgWaet3q7AJoVGY0eS
jnaspiYkRZORyIJ3HhHuAg2vHjJzOd3mPT8vJoydwJJpaP6lx7q2bipyd3RpNMLmmJZxPCttRoNS
ZWkTxEQynqdFHZp85Ac8HDC5W/0XYP5dPygAVsuv/s8FEOrtRuY69z5Vlmpr9nqX28VRpyI5uu+5
bikvuxSkAVG1DhFoeLBc5jWcwnXY/wU0P5uid7ghBdELYhYcB7D8KAPt854Jbm4zLZW+ZQOBeLUS
Ox8HBMOIjIlR4sw2h3jgfIrzyNHYJlYv6xdkQWaLrADDvZ2jnH7ovpD8TVSbXVWpPkPRrpjeZtSE
YZNQ0N2ESsFQ27axJ2X0Nmz0MNU1gN9uumw4fzlabl5W0Kuu75kn9qDMo/5wd3Bm2D7MP/sipXRZ
1CJqSr2Qf0DLIDvzGF6btvCTTzKM/OlVp9rpWbT1QtrUNTtMhxMSnyFBnseZG+Wpr0RRdnXxuU4P
2knS18GTcxArI3Zpchd9IvwHgumUDWLTaUJoSL7YtfqjtvBw1wL/9+ultJDEvpyhiLXwSW7BIb//
UmtfNaBYdirh4BGFq8uz6s20G0ktyLW72Q651iOAnKmj58jzpk17I+s9mDOvZ4v1PUQZ8/bU7653
AVNEJIDF8ovnhcnVS6HcgKNLzN4c9jjiKiBaxM0vr7cZ5TAAg/sVdreNtCocXEJrpra1kEdI46hO
KScqRc2mrLRXDnAi6gsCP7lT16KqYGTZVfsFHPvBf8NKzf5zqxYyQ9JJjoGNcwMkc9RzHt/qP44l
xSrkCaMP1odxUAtn0DN0Wg60LakI4Cv3cNRphp6nMw5i4fnBkz7H2GDIYWCu40HSkh2HceRG2m+v
yN9ViSyoS3gB8r4u7Bp6Rs4Vx0EluOQc9AkiHCVe/ogd1FlyRhGavw9BXs3WVVLT+v+nYxkTLZJi
UgiLzTTFzLQtduEQ9WDtZtIrZMrNx0KKMGoPdNHzHOrUzzAJT9EB/9MWxFuWFdC6ZBlcugpsyoIR
w1v+Hh+S9S+/Ruf0XCqnHoowqpkqZPq2jvFjgIZpD5C/beG/fbIkgaEUMCHLSg/S89GVpo15sadI
8qOQ4nOlt0iNpQc0Fe3SyU0PxEGybJZLROBDOj13ajb0aEmhOnr3bIbLNXj5okq8xELrmehNY1Dv
52+p3cvI3sIS4g/9kMXoNzEhyIyrAz7ZhwsiZQxV59e/PiVHVZnjrzAkRGlVnE67nzVhtHO9ggrB
GnQ/MDtAcGs4qDN2OTt3i5XdFRcYWv8EqgOHULD2rCOa6sfYCdHFn1fsNUIz/UJDUJ0LwdM0TnRg
SLxLJ1gej9QutmjXa/Gu3LNbDSXqmRqRHjnrZbgMitWiqasyWDKvuJi9iHhk9KLy/48K1oQ1ri+V
Eqlvi05apJdq7LDVy+0JRuMADzeDcptdp+hYVAg39rdXYFbsghKb/czpEYldrage+8dTvbclNkql
fqMRVugaN9XRpgZ2dgQo7DhnE2wOnXz4blb0ZqiUd1Hb82O+EQJkqvmG2GXo3vySFrLx2/1RzdOQ
ROPML9k+K+BUsNt5o77tOEqWrO+UiSY3MLMQJAcprd5lHSBH6n/EROlKsPdbmeJ4xuV9fvB0iZcs
PL7EwkUGiTLEWm/GPEwMht1Rg9RT8oh462o4fgCuyCP2rXxmgLS8GMq3MluuoxSWl+mXKj21NcaS
024OXB0Ci01Kw/Y2QRXn6K82/De4Hn1Dv0YvjShGlWAa7cVRRKIpD/6F4qItGsfzCTEZCZoo45JN
P26C+gOmJsIGrcsF21uHoy0ZVvsEeQ/mdXRaE5zah0JdHE4mxrpgItHt+YtICwsyE3Il6HxHmZr7
f2c+RBDpYsg9xb8KWa0yul6USPNVmsJ+SQA6XCeYakFgV6cKr9R0BRCGdAD5movLKbhOhyMoAurV
U1zLXkZW1trXOnIqO1JspRcrw6JQ8hWd9VvtP/rethJHFvget2Snflti09mvNVWUrAX3iP4crsNQ
SeGySsh5kxg/ayvJtbGvoFKjomoAVRc+jMG0BEptFzsQKVsHvdpq/4wb1gEzHS/r3T3dyBFSwXMc
fYHqgWPTo4BL6Cjo0oALgQFrTkme6jLreP0cRACC5JEl+1GWniqoQsbZBHU+uYfTzo0UEj1KqxnE
mb8KZlBaiHkzTtyGpCihvucGAJEE9Q/4swWcO3FshyfkvBC/3y8Fc8o6hTm57szcrpN7pQYLRrU9
L32BO2W7I+lXKmXymasXiX+MKctJc5ViWGg23fetgmRrlMYZNanQWrDD51/m5ZInj/CqQtMsVXzi
Dzv16D+73PRZzsTNadnaBSN5QfHNxBcgfFQrF8WcBjJQyLzUhfnJIoRHthAgWqbEI+71mYmxZkIW
JFtt6SdzAUS69oEUYmptLBdQZX+/1s6EYErRXfT+qNaCwzjWYFYVwFf5exjyoqqMBkCVUFrJqe4X
eoHDLTcNYIKZzNq1jd1ZYy5JGRNQJ4Td+aAsDP24cpybsPQoQRueaZafLocbsehmu464hLWfp6Vf
3Oso/jRlmfy5JEF/27aXdmL+KVmvR0LyZ8izSbvlGqquguIQlHVQjFglbXQqAg57BEQBCG44Jhs4
Ty4eZXFmjurvMF6nA6H31IHynnZ2po0XJrcmHMjJnpuHR85jVxNzMhjhANlESEfnSW6zibygG1yx
508AQFIufMne9zWgFQTcIasXBW8q6O/h/ll1pmn4BXrOn2njO59sy556UCx2k4TJDPwNaVgJytu0
mLJcC37LyVpLIT7IBKX5QrPsfVgBFno4lDoOB2PF0N0m2WrXDwEw5SYBWfXlrlJFvy+OR8QVVKQI
CW/VQ6Rf4085rAdYAUzDAdmjSTxMAPqA6JB8QKCt4vHAO12LNO+d0GVr0tLjk0+8XFpPFg9jfRK5
Pxx/EdA1SizCNnbR/Sl4llNDy/ENpuNWJkie4uib/R2gdT/A/ZF9QdU2JG4q0P1Viis0Ha6hVum3
J8zAbYAOR6G/OHYeIzmoMtsWEsXarcXbaREtKtIYYMP//wwTd6+fmft+qZMX6G9Q8fvM4eBvReon
qNTSOhbFcrAy8ePl03kZmQAE23E60YgfGLOr+3NtEztIdfm3HuT2Rl9edbUhB57R+K3Vd/lSG+NN
gql+Sz/OMo1X2Eao6oHuQM3SPT/qc/NFj0XlxMBfgv+rgKyAovygspthk0e3XV0meOlCvv8+Ql7f
a61c85iRzImHuOHEBYvRcPx8fIBYHy1OR0mDOIP8V5uLFeIjLfeeJdw7r4B/E6rm8jlwyFrxM4y4
42sqQQi5chzOMZ+SZDBp11/nLOrGywryU2FhcJcD5ZyBsAqzaIOaQyw39cRVrMvQaF8aNvY92Fzv
EJqY+N5rI8a3Ryp592ew1CzrndkrWPSVf6E5K4aXED8UjCsKYDiJEo3nMbXpEb2olWsB3Vhy3aBU
SNUKPQXz1+66xKxMh2VBfeWDDla5CLXnsDKl7svrxc2Xzmlpse5XQHiNpyzdlW96mRDzqSR+nBPB
TD0/0/C63OU2DiTulpCvlwEB55TQIMNCenuAMM2GvHzjQ32hPUIvYO+bWYE/sZ+pn5efSFONe5X1
N/IG/nRw2zPdtsffW8xq8c/tKifobrpaILCcSMR+S8oMMR3rmvTNs4KDx4OOnpiMRjnXrQx4Lv0K
wWTEH20KY8slWXJsDndkkqyTPgIY2GfRaCIGHzaUSUuDx6OkCAIgjD5aGgPMWfpXxWbOq3w1EkEE
8PkjBQWPxHUq+eJmYOsAIlyykOwUEkfHyZ/2HOYCdmKBviDUkbtmCczBuq3ft+XygnY1zoSWZ4/j
uD970m36Zu5lFyyUQV7EbmV+TeacgdNh7v5tHniEsBeGTLsuHQG2v7PxCE7HgyxR2t04LoRP64XY
y6HnF1bFER52vqZ8PjVO+V4FnN76REyBOHf6h06gv6nkGX1ueXEybJlhjUaFLpDhbQr+23Ku+0WH
YdhpvK7x5a4uaLb7S4evETAsrzrSQiOcwn1kOtHHAPPDwRSX/aqam5lLQPSzpMiiFR9LhE7qTjXb
x7eAtxPfF+Bj7xwSmlgNQ3S90NuYD2k4+s33wl2CKcqQ1zDOOhu0l9IG3U8/xU/1AVJqWLTkeSjl
5cXSmIiDvk4S215vuCwor/VhSc+irdQj0zBDi36lmMBGcl9WqBMDCuzLB2cmW6NIOfttxl1rCg4t
WTOz4H/EWs+peLkWgbp+pxPhicR3BufMyxTdft1/coizjX11FUtZzA5McRa1A+TDb9/DRhr0o9zn
deV4W3NJI+noqf8lkfJoJWGQx3bGM5pGKQVdO9lFeJQlOKLgnRvlBZX0Fhx+uaUSEBmy1l96TeWQ
mOqIlFjP7vK0/NSQ2Yycy97BytXEjBTgn2Lo+lir6zM9rQj8YdmjQHo+wrucBBUqMYZTMbnSTd6T
GZ05N2XAaHZAzBAzcerhkdiM7aavbNyIr2SkyTifkVBGqjqfKT0XZNM/n+TEcajaKKziDiZ4ca0J
fFcq2vx3aFWY3KGX4UhVxbsTMFpO5xnj+KmRLGHb9nR/Cn5V6b6e9ErEMl2yTXxFrbzX2Je4HjGq
ydml5NHEDZOoTt2k9TeqIh8pn55tXhtp2sD3sYGCnWFr0raVYz3gA+a1Eld3zZJgTwIDDBQE+es/
hJRZFcKFhdVv7Fb8AHHJWZBTXBLDIbEJeBBFjzvzw937b1r66WLsYNL7R9u2N8hZwEgXMQS8aO1t
f0jp5mm21ozOfn0bnTH2vzLmjylLz6tW1Im2dsmW7eUnjaISHp5sbZe7ABU0q9FOraxiD+/wiPd6
nvCcMeLM0cLZ2pCxbVPTsXbvoF+cY0SAF3uMuZj7yX7DnZMqOeM280FE2vt8cqK9qGBvhLbyPgTZ
RHqlzbce6CU5WeSzMpWw5AswcLFB9x5YhIW0SLmEUO0vzh9z+ZC5n0nAA6frr71sJbYjf4TByqfQ
lMK6ImUgB4A9/xkf+CKa4R7DiX9uYrVUHNR5Ta45KKGHOrWmiRRFOjb4u6QOuuUypAcVRIyOR+kC
KAsc5aB2LSNtQEXFXw1gjl0PP6KWhPjlyEORiWxHJgNoBX7r5wsfBR0Dpx+S4zYEJhB5V558uCEP
bBcyGAo4fFAd66y0/8G6Sa8EsaMaZ9If72dFbztb/75fcbG3Ka8jwJB7GD0LeVQTr8vFxZpzGBfk
lZfIxN7tHxEJcCH2fwXEi0Xbh6iTVKLPxcvvSgzid4xnGKrvuChut/Vp3QKpZuvE2gjbpYZ9y03k
mYZ+3gZk7KPend6N26+/+CylMo17uyAvcN1AFZP9iva0Ki7EKZodlQ6/fjfjtFufdaWDC60GjZxH
TlZqoNDtmbZulcOlYwY0go8AYxGx2Nw5sFpY/hpogCzsciZiFMYomY2MQb9v2T0lOkPNWbAwp6kG
W97i6HI9qZmL9KmJsG8LJbTxiUhnS2atHes42N6db6XVfc6UxQDBq25eULER9+apsrle7LZIAtsn
ZQIYGbdbey5chQTA2STKcq9UcyIALSiUi91HeEvpJv6kVniFxlCPjbAN01wJiNxFT9D1hhjH3Qm6
VL1jPzCz7KUKcHJ7Ud1Z4C1YJgHajjvWbaUSEWMj+SqoZCS/iho7jaMktn/1QJbX60BJDgDpLmtp
9UI0EKypF1dEebEonE2rvPu0u2h4RDW39b0GcW8GuxS6VIpME1REhtbhAA5VE3EYth+oUBqT4hdS
cbL1I1LTt/ZB7SmDaiNHCH17IUEpmSwQBLmNBDn466BgpxyN6V7dGW5rEL1XJOtkNwYpy0e4fUce
EwbFUaLzfxYOtW3b79A++x4SpIVkwvLlS4/t8xdu+5+Je6Mwk0OsR6ooACzfZm+c24j9KbMeNnUI
8ovPL+ptIRcNK7wHpwg2/4RFBTy00kcBU+i7/oyS6ZS0xDjvA4fhfFcPYU+NZRFqTbJhgU6ASuaO
bqVN2jYvBB182w8UgLok9TzhswNoAr9ANqIpmOogOVPd57w6ACm+sDQ/pLLwzEcHs0LY/PBkciGa
pwsvi+kq+XVU8S3agjYeIlp7Op4doCKu9bybDaTcaEUHk860wqkiAjIKBhQlLye5M5xAngg7odgJ
HatEmiVNpdNoFKX+rAeFOJfiBppjfj2DykJWMvWMDMQTytZUNYrrzXtcZouxLbF3ZJctX40oaeSs
UoVhthwHqkWjY9OwDFUjJv8bUVtfPnSXqy+I1dwovSEeKBXGxZZdwm208NVo18OC7d9rlRTdsF8Q
yUe6IRYRL8E15aF1vdo++kqY5OJPPHtCJWiQb93Hrxdtko60bq5VTakmSkm4GnDBQ36iBzC+CoSv
+8w5pB/sKw0DbpPkbL+T7d3EphYqMvVQnFUFVYbi0omogFarta/fLZp/jWuFzLZv7ASutEEmHSm1
JO95VfuOuCkG1g/wClQWJ/B8cACEoB6er2TiUI7bE45wjygEggP2JiH74lz0hcyAuLWlvBkXb05G
QXv4dc6XtxvWRYSktCbq54dk7pdrBrR2FPzduuilp8dBS9690xaJ3qgkhVxx4po2CjVUjxEfzkDr
Jc5zgoHZzXembrDFGnQPbV/BUXybCsduty9c25pMuBQb06TDe689shey8yVUcmHB0Q+8yw51MCKr
cavAfruoQuJIdlmxA/OvlW3O2jB9io9tZFh5W8LtIgJjMCIWc52hO8v4Xskc6BH1mIffN1du9jIy
yqBQyyvbpvVbcOqi6VdrgUSBb5rUxM7wsU7OZ1mh+j7dFD4kTWibzPEVVVz3pnj9Ac1od4yPupJU
jAaIFlm3mOpHnuwV99bdLweikeF5DNI1w9iwXZWeSEERfvfUqvvI5YIwMhkaElQ79eYHcWjpQglO
mPmtq0U/z5r5Udm5lJ9uRrtz9HyTyOozVt9Isrz55fx1FkcZBMQRbwW4KvjUtaJjlTfT/dquKX5I
1pjx4AfdLPumCCXKb/8F+T2J6m5r8uVI4jRERg01vPadoM1A0RXuv8GH6g2j52MbQv7V8Kw59JuM
uft2EfQr4qk6ZO7em5a73vtgjwXtxSof83scJdXLckUeKNLyicnskl8gogfVXBTCaYhGpVjLZSN3
hPph92+92kAuUX6BNnmQW1k3buzh3z7jMX0S+qzdy0firsAfoRutuR3B5gNX78WtG9to+EA4EqKE
C6PGnK6ONFDfsl8Nbo7JVR3F1pQodTxToiG4pVXnCPo7RIup5J0MrT0RLtIJ/j/UrccrU4l8h2a4
N9rGvjVu6jKDPinn4rUKk7b+uTlz1luNYoaS2I0T6xZBmYLSy5XES2QD8xnKUAHzmSH9uMyh02mt
/T59I1wHFRpxZ6yRHoZsdLSTfIrsb3jKNpddI3mCYRgMxThHwFAwwGwhsZAEgNvxbTvC/PlQhEVS
YbpF/cS5gfbRtdqBuNUZmix0qA2EZOKhba/ylzLb9EeDl9PY72wbx58BdmIpQw3j9wbVpPG2U6gq
iIwlNoTvhe+ixPqVEzMBJlnDi5KMu8OPNQFhhzVKIcrK4KKolL+6q9J4SxZCtQiLtY1ZWf7RktMf
8PtyiPmZrgCOcIEGPIygC39szEnRbnD1VJeT7v9o6graUT3B/n7Ee3nJSNTDBeFYCYhx2GyGO6Vh
jBTgFcKDWBciXI3rfqMA6nKC8Zhwh2Bezpt8rNMQKRBQ0udp6/UpXFrqpkPi9/xN3ZLTbIlS9/74
OLo20MPnxNaZCzCh4AVKwheNSCqJBDRGBRZDI7DCNBnnsEjZubPk2KM83zOCnvc3MnarnJLQDM54
ks4vSgGgrzD5iLQ0icI4r8O9hkT+lj4iIpwM8aBIDH1OItM1tcu2ns40gCVq38PkfZsP2+f6JAAu
eT0zRtMQ9JnpkN2ysjRwkULNN5H1dWfFXhfHOqajaVw4EtneVrfGJpTSKzrWAJg4fSlnefHdGZMM
3t2+DNoIgQt/Qw7seHniY6SS41EF/lv9jL08R02WU6vTgZo0OmAWW3Pbcf3V3SsHoPXkR7CSTmiz
U2XKjx35/KOfQjfYPrOfEqsO0/UY/8QLBAs5fxg60YbcqKcD2NLAMIaIsLz7quylrzzackvz2cTq
7W1qJKhn0Zbsv1Kxgl3sl3SXExL4oPadb3gNfWsTAyTzD1HFBgjrje1fr4wTVM3mvwk0xNBtUEYn
sbFd1zfG9tKM2Sgch1wWtrcIYTPh/jkMRDtCU/djxWHsd7QsguXQssIAeCklbj6+F0VsUZBGZook
eGuK0iGdvVejTaXcIdr/eV/gOLP5MQ1bGwFxIrcWrI6ePebAWuA2ToT8clvqitHhcsWnlLFd2PLX
vFze4Pxkohpw/mDn/0DkoXjl55J2K61z8DV6dJ9JAzN6T8ORgG67HeUkPpF3sSnpzQQVJbrixb1g
An9pUd7I/r+Wosfti6D/22y1cLGfjQceZHNRYCcGzyF8Vuzd6d5B/5fUd0d7dxMVmW/8M8JvEGIo
WgG6EN1VzLB0+pY70zF9hxHeKAgnu8Nm1XvqaRoWGlkfVdDk1fWaQaSzr8gRafJiaNN9xELpy0/s
fU2nRYoepqwhSF/hitahX36rtd1roNM8y+6/b6Cg2SSlhHaG0MklL7HRhU79xavSYUCX99OLW6Uc
xhA5CJ1kUvEsfrXDYrH+8UHkKz4h3yOdaf10FDM0vyewXyfcQXyg9kob9w6Dr6UnSkYSJ37/HDhb
bP+HHne0K5ZvxnbqA5qujJ/lhYZZc+dJjnRgUizX979tFChrKu+lI/xUewaSqPmfct4FM7S9sIgA
iAmlKIZFax5GkKMhRlHkPW3Eek3cxhwzeB7nBINxr/Sqs+2naKldQUTOAGASVItVUywCHw6C4ZYA
24oWZBHBzhLlblK0zrTTUA+t7G1sfhTuKBooZZNvPdSwsVkIg3TdYB3mONNcllmk8RWsVVW6lDYH
Gpv17KYeMk3E3xpNJH1dSRCNdKo5psqrRv+R2Ji753iSxdexk0qmcR1r/fXaKi0qij2kVZB3Jw9K
nyqpdv3+9z443DPheEcJAoWgvAX+2ySvP7qt7K4wOzPOY1WTPBCvabh7qP6s25U+lm8SWEenYk5J
6ytHdOJwWtMbMZM87rMIQO4uxNTGCQEVY71Q+gutEsXy1Z7lPDafPJfhYDCZoaXWLj48E1I4X0Z9
xHEjOu1RDFEYXq6c5bAw813TyTF1lPLkLJDS3eVqReup1+eqBdUSSNbti84Yca/1Xj04Xws2qQ1l
f2v8Xugyjo/4WeTBONzFgfvB/oox+58eph70zIOTT4whCF/A3nKqwNwx7Zaqhy0JRvM8t9OZ41on
/AE5dR7ZDFnke88Aoyp/8I2bGdlaOpiGaWr2Hto5m3zoUOXq1t3QENuE344bR5enATOzGXoKIhP+
oat8qu98Ky8d4kid0123ha8n6lJOwicDSXWgwucZFhzyUBqUMyUhyHwC/MtOgnB85PHnBHPPxzsf
f6yr7E0gDKVnKCvBUoavrxoCDtJoOKLEZJmWRBg4LcLDYLhaVHplXCBPIkjCRNDFQVWhoOqVbtYQ
In3RJ3zQt5zHpievAgpfYU+8N4J4h1+rYjiX7AkBZazAAe/sMZ7uZbJShiJEz8NUNdn+ofRBwOM8
8fQDQGodvuVrFmEBLSPElOxXEdee5bct9/6a1YPEN81xtYN9f37QbneWP8VAOId3oXD7D+22Fia1
ub6kb2nUbVYBMcMI1hgUZCKyLEInF/nWzVgaGHYvt3rDSi3QSM1/CvJZrKb/P+RC3DiqXJ6qQvSr
VzrgubgNFCgk+O/97wF0O/YfFAXyygN2FWIw+nFbQHD3pbxnntFQDGvR/PqoCPy3MW0vvgcnj8FK
nXbXZe7AwfiLGx/fHlTRZbp32sAktcJlm8pcNi1sI2hJtZST2vVo2ulM8GYL/OhcMtJR5mezMeb9
aHt6gF804NMeXqrIY7/wynTvtcNCSlQh2YKrKvUJ41sRsREgown/N/kNvEm3fLdXorBMXQ2JQoQu
HxpopX6lUPPf9Vgar5UwM42bk9YiU7ASV4CCG/aAVEAEAeEh4nrXu85aQkL42Wp6zRVdsHo/DYym
c1yGYWfd4CoXgV//E6CHcOd1N1wqp4B5W/slJwiNZnPoq8bpDJjMnXPq+yHX3sEvmE/7BhITci38
gEPnCUd3dBQ4dalUx9S75BJmE5WrSgn5PxQ7Sn6R3FIF2yWLN58tcU2aeKnr5NYYf62VDYsaqPwP
gzzdrkC0rF0iQtNfKgIuu9xy7o1wZT06xCeQiywLiShxCJaCZMS+idY4FYG4b1tCu2ES7WuOY1Pl
c2t2jGP1q9gT8Q7E8FUSH9ef0UpCjdVdaLbZVByoaZSwyn2QsGjJu/6+GdFvTvEG25W8UREwsiit
8zq1UFuHSvM0kuG/VENX7Yt+XzYwTPF/88fImNd45d8P1rGr0SNe9StI3QobXwitchMx7Nv7fEms
ipoYR+7Hj/yqhT66dq1Guk+vjI0uTkDDR6GGY+dySUI3+YSj+VSqriJROY9P/9rDua5DaCKsDUkf
NB0f6/XY/EoXJlMgW4tOVT+z/uad/96Gl+I23SHfSWqbo15lqxhR5kpeBv3ROmcrBb1RW9iyswle
vFuyLa/JF2vvzG8nP3v11fm+Gf0RVRh6i2/WoLg8gbvgPlKyzLKebSmmgsImdsJ5c1Iqrdtw201f
k1/cjlKg5GihIHfMsWIa9mSs5f0acrxMnqoaL+whZAYKKponAQ5N/s/xgl623vBeJOzOe4ldMyQW
rlIe7kJLPSbpNDNDGj0w96I9+hJTthZ0g0caBRjcEUPM4mF8vTDTj5GcaWwyy9BwXBDx5fcU1fGB
Fqk+c0FNPfmNUZx6Jf4qdOcE0dxtnB9Hb1MSgyZZuFNOy830JvBurUDRwIEcyH16+/Di8ZBroYi6
kq2swJ+12mOClZ6URpHwPkUXZ1u72LjxPfaIORS5WzAXJduqsDoH4UdCPK09uOxhP4H7OBtlG3RK
aPEAy0xP5mIpJA3WCAZxrptVpfngA6FHYcBfqIS47OpP6mQym5sdJ7jMGFI9mF4tT6+KtAkSuQeX
nfh97qq5x8dLNI7eQ58PiuWUJF70Gr8rBMHJKTs2EyjMp/F9mQ3nJ5hTRNzV1FGrRb7rCsyLozIN
QyhaAa802QBi6Mfocfl4ftu3dWsheQVV8MSOlNw9wbT1k5nN/wcSKPsIM6qxP/OFdgdJVC+6BPsx
hJTwg2AaS676hX8n4z51wdhzPm9su1QYb4i50GaYlTB4EHZa52JoLmOxSYqLXy+1fTo4TjXjiNP2
9TwfrtR3BzATXfofX491GZCzf9Ou2APJTk6CjFrOZl15LCnpAqfDkTmiJWljTqL7zBOGtJlz7omk
U3/p0YYd8K86hI4P0ui7STY4RnUt7uOIRACZ2ZWIdJTtfVohjP4SRuHNJXWUTLKNRHLK+cJ8+NI3
XY13s6yfEpldEe8Gmbaa4eQ85ns6b2ipRsJwll/BJJK98hVtVK6SdNZ5i0iy7Lf/EVgPJHYtooQ3
sjwhme3UJF9+tKe1jzRMjzpvkMupvNuJyztfFQIDoiiZCREmorzv7hFmAnLbLcuDzG/G14HKhadx
+27l5C5rSZ/jjft2nzcYQ8vB0UBaZGc157Uth6NZBuWhtaVKzll1Tn4t1pjzYjmGT1WRyJMvJ0yW
Py2ehCMIlMHkdH/pT/qF7wgUNQ4oAf1tl0P3jPPh47ODjle+uEHc6X0+1sgQpP9ulJGMQj+NzPKr
MYRYJN8W+4wzRjB4ZPtaiZvKwO2sPsRMu2XwK5hHRT752UhsKnfq2Q4hvYuRE//gkj/kQpX0AwLX
PAWfiNNx6YWd7V00ddSD4gUNZDHCcPHrmI6NANhGiImlREiuFB6/CQFzRcasFoA14nGhzil8zu3F
DvCj/qrt9w2+Ce5Dy9uTA2DxXTTO+4gjGQ6fuMmh2XNInqOpXlzmg/Ljett4f1OZ9aEFuzcKPjck
LnfxRApKuKHWDIzT1mnn1UDGq0m+8mVPOZpvea5+0/Ba59M+J7E6qSAy+mqmh0TvA7JVlxfVhkT3
dEDHoFEBao1WOdo8freldqHWLwxkXe4WMUShFbBjndbxc4KGgOeKbpy4IHlaq5gwDZIN8Xnz+CCG
oWcWwXfzurRaF9yQbUmwsTnIgcRULv/Dka9XBMJQwLY2mRbVRyna/U07NTkfoge8nnUOT3tAKeql
OlWb3H5+s9r9QLT4fSIjx9McygI4jbaeduNzyU3ZZexmrVkSf5+emWCb/u8rvaZ33bwn841QC/zY
rIKE2+fCDNO1YmPRqV2HbIWVqRDBfjjWPsp5UpKxVDb+v/UAxsyOfXo3xvjzdaHh6n6FzWDLLPRm
mVBPPFCEmIsoBMM2Cj9A9/wLUTHJ+QAnQcShNgoAns4ck+46eHyfY99qGa3QaEvANtJWNFJFUn7R
bnOY89nGR4n3F8DJ3xcQEWHW1a4+gf9lWI4iXtf+arKZw9ASdsNXc4WqBZVFIskx4YVxLyxvZXzR
CoaKQc4GJBXtaXkza1H770QeWBDc/Na7aq8UjjJgPeNWm8Z6w8HxCShMU1SAh7PmU9QJfJJWcYQQ
ZD/TyWLTOGewUfrv0EsoSUqmht9l8MKa26NZkiwmmVbKOMLO88idZgGUPZZjaQbAyjLkpXEJU7Di
i+TNV3luzbdi7bpDwOX5w7LT1VjYPwKp9XbUlRzWFFCrrx7OLEH750n+KVKAjB2ZkLqRpYNKii43
XK5cZ2h6i4ntqbvcA84oUchRedpFet1aT9rv7iKXsqU/UC4XnnkLPTUuzQwUIdR3QUT4YzZQ/+m7
ExelCztz3gM6luMP8gq3H/V9uDLVMn9gYomzlR1hJgf3WpVz/SljMQMbdZlxkibG+ZPe/cME+isX
FvLXAue7JM2k6gept6FGuY3iu3kAuFFaPVPsqrO0nvgVjX1/98Iag5xg3LJdtWf2son+lOz3SIBo
0rpCidzZIcwvttxgi76MF1J/3SKqhX5oSK5Z8H0FW2S4cGjMoqdS6uAPo5o2nbCyQAtmcvBQhgJr
crqCVf+HQKNCWLw5tcNzKcYbdYiJm73kTxUKBA4+oqXRzxcemYwBbTdKxnb0WlmGPyjDfX3MCWsI
wKcgI+ev/GcIM5/IMY85FLwO6t2r+LgiK1+uPMuOoAnHchcZ9YTowWKzgXnzw9MKgpe04VX1HFBS
ozOWzu62xycMEp+Tf3dZAnCPPir1Tz9OGf5BVuHBKeHQdaaYShNAkjOfxPaTsIfBC5GeVwT+su2J
zi7SkTPMJxdM/FMMAci2oH6HO66p7BDWW8ihGKoiCItEw6caxKhDwIrbUj7N4n1bYPPxllpQZMyd
A6ZKY9aeJayVy1CHW/hDfCUIimLd9ioHTwk/cPDx/THjMNBjpX7c5fT5Np01Se7nArSCaHn0JpT6
PxeDes0O8M7fCCExLclKBaJw37Es3ijMxUR0OMjIJFYJI8pg89lfVK2dUSZ7MI6MZEZI6vPVl0fw
yLwFfW6Q24XWtNFrDl4gUV3W0GYYA1fyQW7cQtBIpmvHMf0U7syTBW6hIwgxRy/jyy/8oTiQhFqo
XAIv5BEZ/X7q/+G0aEHNRyqVi/QzAWWz5mGTBwgu7x37Z6xRysuUqRl44XBk5gROHaVfUtoEqm6Y
Y7Wnx9KF8viHjnPrr70YCuCkzGRoZncyu8MbOXlIy19qVvLqEAJ4twtNVaGhbh3IuHC0WRdKqRTx
dorbn2iurDyBwvNq47QzVEteW+BnvizCYq0ubQkm1ykJfUEChrljKDBWdAcWBh4RVQrCF/aJdbLx
VpbV19LkOd3T3G97SPTMh035ZKAFyCY89X7Y4OSlMc9Mg/p2h6t9anOrfFFZR2Izo7IW90/CzBHE
kSCsBy7hLol6tDtgjCJlphqX7ak01zE1HFA71cFuxq9zsFtGKqEh+YbktrXwa6vmO9eOlE+H+zPy
c/7bcmzwtY+w/I0M8/YQtyxAB9455KyqpsHB1jcdV6MOXH+vDQVyDTdoXbW7SvJoxuRsqYrKuYmW
VhohzhBLfdPbW3pMZ8e16oNQyPrPf5mPdGdJYip9qoefb1e07iu4T7Si9aKJHiOPicJbxaz8mXsQ
mI5GHdQI/0igTeWuylH1ZW6O+0Kw0daUejE16Cyje6szAtK8D3RGMD2jF0WAAeR6onCkOPODsfcp
DWolBsUOnIeSsAQTF5IW3VcUn9r5Fdx3Ll0r9W7Z+UpoMmKkl+m8Fpz9JAVyQ3upk6LrHiYHIN1F
kdr7fpSux8V99nW+c1iVaiG9ZSFDqVtIjQgBK0IL/tcLTg3AYu65ZDGjyq6nTLjJluJHJYxoNAwQ
HXaJLa4iiEURzJCASaOgrOY7EReAJQNEFAosmLk0Q1FTVZ6nRzC1ftuqncDat/p8Fk3amHaia7PN
9ZgJb6mQtDOh/OXBGvsMB0dqBzd2MLjzjm33ppA49xnoT4i+TfPpScQv7dTzXFQim1E/y3dZJVZD
AAc+2kMbUhusTeO5T/hQOJB9Rcqzzak97705phn/weT9I01vuOBwtclvGzgSkoFPvEzuiJoocqp0
b9HyqqHFaqyDt2ZIEqEE+R3pI8fnwtJp+DPzN/zJqRasFWTvyxPzzGf1JKr/yvMWPDeOKgm1mBxc
ChjT2QD9klxmR6ubjxxfqo8JlmfQTYcH+iATp5FPuPOeQn0wzVZMx40NI0zJu8ECOpA1pHzty2oH
MW3qkOq44yFAvWX7TYTsOc5upDj9wPp+xJq9A/2yh3C7/72n5ckOO9tWRe5qIX4nBC67Rl2bK25A
P37ehf4+ky3ORezYm/ozFkGT/2DCq65keNhlJtE5p2MAv5uf9ETahWy44KHJ9saMxTVyD50ERifH
1g4LN+Vi+pbXhPr2j9zQRjDZWNpBkO7J02NTjUZXu+YDxkJROcVeAa85quhHix5S+uukEkORz9Ld
kxp+TGy0YBdFDlmw1L0k5gPnJ8Z+NLm8OtH1klJOvm6lnUijq1Lb+CusCgZ01x5pmglfDYPS9ekY
5/szLslVHTrrDb7VvPYG7EcqsavaQ+W52opf6QT3fZvzjOp5nmuF/pcva2JYnjeCrm8JV40cH7ky
sD96R2qXHQKqyomyDteAagJTQ7GOrxLRIm9dJY35rV2edGQ4qTtZ8xjkJeHbclmrxs1YLH5pQKZa
gDzw6mdi2BtgXp/qOH1YJO8XjPTjgAscwabhtxsi5+acKpfFXkzRZNQFCFsv7CedK29QpbISenG5
OkMVo/v1WIYUD8ScYVv2H2h5RCYeqfuX4G3XBm0RJMdWL1a78yWfmWq3BZ/OSQEdLELfwsvj6tjr
hIYO3LxVKadAYQIwEdi54JjNpl3eAy7TS06z8RVgzgDfUS4oTW6s27gO98EkJ45SbC2/aokqMyLb
qAsd/LQZLPZMwFMsdKX4EWEPnrwkpqZ+GJn5bPMPO4ZL9Yl+FIqi2Xy35wNs4X4OqgW4mWdPKmau
QuCQGr3a5q3lq9+vlRLlkChM6M7asl6XoTxwmIYg03BlhQLRbWBzc9QKXEn3i2wQik/n93ePUnQ0
4Hzp/E0f8BwDdhRk2sqvhAtXn+HtFjWeIWOGBA8LhBl4qhGxcUoLk/hiU2PukwNBgTd1YYTMh2Z9
J02iWxekg16hpAqa2IrRoWiWkjMb0rby5BQapV9wa8cCPiERAzIym40wBZ2gHxzy0XvXm20Zm/s+
PVzncRWtBc5jJDE3gY91tkaXyfCQrQiCquesuDnZW7wzqbO6x/45Y29wPakMe208b26hR9uewVeg
RS4rldhltprsAWK5LK6BkOy9hTdCViLpjL8Qf2ho43rUEI3ElzsQddSW7qePSWtniih5/B0eR/E7
dWg+Nr2XAu+ZPbireu7Cc450DylB2nAjcU+AcGy1L6eUUNGOJNb0nXNZ4bB32DRj3ch++HbdDxVR
m5fxEFsnP0oSdzsPB5YqWLRezqIFRjaSIkFHd7ZTJOW7f/zNqrf6jiFk/aA6sKt6uGIZisGQxBZx
H1bsO+/DfGXCSIIfH2JRM0HYX/X5g+MCGikP1QNAWv27XBvXskQtay0sxdDBXweMoszNChiBhHs8
tDij06wjY9XBzDf7Uadp7ZACXJEQuViW6F+zuOGULLtrf0ObQGb+4ynq3b+cEswFU1WGhsizyHp6
eFYTan9xJHNj7pwLAIsL41tUKhYgbKWl1j6O06BLaqcuKwGqSOjXmebnCCx+zJN5UizcKhhhDhoc
xlN4DfrO+FowTfmdnTA6xIrP5qTc8gzEDCy7Ovl7suQrgyFvpb+VeQYfwrFe/UynL2tCcWOdcdih
7F2F3UYttlFC95sUIMf7ggkVQyRia5dK1rzmSAV2CElOwG12LZ/uoLAs0xkj1cT70/dha6R/XqWn
hb99AW88k617W3WJrsonu5wzgDEBHHSFy3P36StHBcncJ6QmMlx/svKL2PQ+xLV432W8RddyA5fz
kFNvccWSFuBRcfby/OORGwToWKtLhbVV9OhYVpKdini3BKlMb477+5qCcJdsW5untYW6NADdWO2J
KMsJL8EoWTouo0V3dIOzDwxWRBH3FtNnzSppSoy76357+5K5KrFs3s638nz0ef832xZVo9AeUwgG
bHMw6+muLcDuyPY61lM7Tk2raNWKrf5Fas+MBwcGLKpNe5aplf82i+ZBGR117rUkGCs8bddswNAt
+ecC5rBsE5oiYCqzyZb0Jlk0JekswZKocT6OcaXtiUa2GBDlKWHDrR6zG/jsBueIVLY5oTK82do1
OXTVlBF49jRpzY3EcCQFLCvmMUkaxB1VjaE4trvbWucNcpxKSxyGABVThOeP5eFOvBfoGIR4eXpV
kpFRXoLF5neINmC049sMufGBL+GAQ1pp6FTjabrDNoHyKtYA7wBQ5s8hYUreWiy06dsYENpIjIcw
LZxMv3PcXSRwWetn2o7PDe2QPaGLJl9cK+wAJLNuu+QILplJMDcYuT1Tm+dmFtAF9wQTF56jIFaz
ccwEF9kl+loKMBcGU0W24vHWxTdoVOCSPklKdESWPWb7D2Nimtx76aij49xLBWfogNIHp9a+3b+8
ZSa0/GOYv9ITze8+eRrKBDbb2L9CAjizvCG1sMzQV027u6a0gxEL82aod897RBpb0rGrR6eOPlqO
6fuLV4ZankSHmZ9N2TAs/hMvynBcoWQfVc/irkVG/u88b6Ckpi+fHffMMzEFRpPYoMx198rqGUCA
/3ryuEF5Zq4RDFlGi51qjoVSVq8kThS43G+q+chppxm28FwS523XiDfbeO4L1ht/CcaduM+lMX0a
PRGNxDI1hw0PPrJpX3NgUPuKoNIzyQV+gxErcZ44Pu9YZJ9Tk3JhAUPBadEtF2j//95JDPkQHQes
tIreBgdsvJuWkRa1lUSzhf7coqXnNWsT/6/if4TFR6Wu+fjEF5L2h3k39Ap4S10QUFpE469skLf/
Ml5pmmppcQCZAMy6VY5tTW/4Xm2lJEBys/j06IC+uCZpiCbuCuWNzium5PeS1GjHDYN5zkE2T5Ac
drePFHatLXiThVTrOzeRGad4VtOYdAuW9Qrtf9ykZPmExUOZP7NoJwmOvRfa3so3zI01pKkrRLfl
/LiBlH8jQBcOnQ026m6kIfre73yrRyZiRLXvGt/wE+JaG63NTLc0h9Axj54/kB5elIxlxBv1P8l/
dkd5L5mlVvK7rL2RMsx3bb79hiUtvC1XkWkJGtVfCHdf6984BMtsFP0YpY981xvU3fnXVVLqHS4l
ZjF1gDJ88FjMg0Hh82ebB4B6j9H84T3nwoj1l633iP4epZYrr/FlsqRVTDs7VUiSOobqeF8+HXoo
mLVg1v2I6EcwHpjNtsJpPESbQi4tcm3w792BgQQiNTEqnSzAxA0hW5Mx7ixWWuhLDA1IO50CLTj+
4ZMuf+8e+/ZkmDkQZ5ZBtQWEWApNgsRpxdsR77wBLwfeN3NqQsTMZEGD3DuaoBYiLzja/b9TWrGt
ST+4vQIZ1PbD8cGk9/NFe8Tns7o/dVFgmzEaCPP7Iragw78L9fc2JuBwSmlnaIgMsNLwOBqwNm1h
EInf+gPBFnuDynmsQmNQRGj5lS5ELVJpsWkYegx0Xm8tAzVij2EfIPgdtBs75/vK4JvUVQRB4GkS
asUymIKQXNtlumPZnZy79gRNQGd5RrYhxEV/SI+/DDBj6e+3U7bUYXGA9EgxBkIhyDW/iBwHRPq3
IZqS53wFa5W5JYHYGHfZSNU65RjYnf5ehOiOsMCNGCC+BihVDK4gCwDelgei8rN0Q1zWgWPVHxzH
c9caq1jtghPqfl/Haip25SrySjmbKh2QHuqEJuwb3bdELcS3yrTMbIoliEuT+oDKIAJH9mdFVKl6
b4c2iEu2MQD1US5QFtRBqWwelGgg7o+maRZigUGnCb5adzH+aDsXhBMhWpETD/UwmFVylhH9TIqy
RRwKoz70fr6xUMSTp6+orwPrYXE4ZLhlLBjw9/7z6V2u/Q6kJy/cFnA99qQIDyhcTEk9LM/ptSnn
eDdFKjY6Hcxb4B5qvvaHB2SZJE0JRRcxS5pWQ8qNPmW5Niq8jYjoWE+US6SuMLReXygpY3l03b97
5iUrZLBEM0cra/2ChObE0yPpSYoC+wd+91pKepVZ1As/iVxEw0CjjwUO+OpqG7RyHIQQKCIzK52q
4vDvWqaYDDyppwgBpG/A8S43bdh3vqJT2WU18m5lj5y8I+K1nkGuOAECgYIv48+cXeTg4vzSSgk+
1yX5BmtWixLGRU1X4db/x5+at5lfVNMH/EvYPQHihGP8b31Ys5EDwNYq0BQ1DpmWySSXO1Qhj/Zf
CQT3nept+3Ad1bjdrpac/VqpxqHJNye8+znlJPXKkXbdOQ4rUC9zIfTmmMWYKPuVzPm0vtXQvX5k
+PoYuvv+mgrOJT4OOWEvmNjvLJE1f33wrVb/i4dMRJ9sCSBuVOS5CZTT7rG2ARq4NV3aIafFVCU6
G32nX1sSvl7QxmNxI28peZB6ovq4y3HyV11JdhnoFqiE7o16MbsjI4gDVC8/NqquXY37QRGGyLrx
54wAvxJok8BQXT94okHfBeoKV0OB7j4jLh3CITKElYNgb4aKxS7XQIkgK5WC+izLghCOSZ8rwUwV
n91uX8u7UAX17NXeYbj10bmwVjEX5DBEDpzNthDs5YO7veeeU+sPGWb4WM0nFlA9VmsrrFTuWmjr
lks+8E4LxKdju2Go2vcJl2yzFKHsfvXQje2xoTr5RhxTlhxQoTO28C6cYhfqZp9/GbyeoTZwq/sF
ZsxStX3x8KkGn9AJc8a8tEfS0QAhI8J0FLgnoEnsLLU1EOw+Cop44nqdq56NaPBEVeB1kCqyoCUM
54O147Xs90GRcjfPH/yTYgUk0KlR7b6cy/AWaw3Ru3MNgC4KcgtNdP3ETjM1b7aSvqj8x1xdqJJT
A+hV9TVTI3J4niaks7tYbGFQgcEVUrN+tjO/fpIW9vxLoYSpHEJE9mr3gnrKGZlgHvlGrN5Jk4j+
L6vhSEoKcGYWcJagee8uGOE7SrzTUeUOZBlMgCMRfoiZkR2yXn76Lz/CGJLZcBGHbiZtAUCulBOc
F6kviI/PaySumIyimkI/9F+Vhx8dEgnEAfldKdsLmJ68PjgeM9ZPKiQAttGiIwnsWrQzuGjwauDp
9jc1gZCSiMu7QkMwh9ffUYzNWn/GMsVscpzC5PqQ7rkcIwk+xFXrhO3v/lWHo2aLhQjcj1BRmD6v
tVGSe9Ez/Lij3tY33xpXVGAFP538CPdaRcuFjhpnA8DdMtYBeZhLCHDCMwidZ6tK58Bu48e5q3n5
LvL7QwiPqn1PNBP8yiT3gGzPJTyE7RrFJ4Z2eDHcTL6yLCM+WqrimcsmcIeptRZBhzOHLJiMBQjk
h1QDQQjyzWaCjHqH1/5yczsaj3C0V39CGImFO9tZr5qqhSdFaRP1qPgDlsJi96x8fJjM/swxnNXK
gGUUqSuu1bLdhrr85qhfDH7f29WcjSTHSlAsXi271de8u/W45WrV1jzeY+122kcSDX2PEi4Lk9TW
xVq+eZ/YBF3QpSrTSFkJkyxx49fgw18ND3YTAXBUqOBXXen2Xs2ITceSWEblAkB3rNNqexO+8CTd
iwASgak/8f1BRoPHZE+iDZbv/kj5k3MbJUZvgVKbrlSakfpQDFdHehFLp8FUeRHkVmGjttJiRBeu
NAGINJEoiONLgc+bnI0nw01GBX+ihyuBl/468tcp2Rl0ozPCEpklqYtyrcILHTSE8vZkgBfV5KYB
wbXZHy/ViLUqNluron/vvnDGgLkRELNIxs3fRDvAXa3AqSq34raKwg0wuC65UIMKLJ36UIWU/EGM
aJ9dypV/jKvkVyuViPPebKL2AKpzLwxd45HWP6xRcajSPWjHcYrPy2EWfUPcTbnEWoIym9zDtdTQ
XpEDLVgufN7NoceYKCKVJ6VoqLlOLaa+bGKeb2xlPd7t03Zx8/KNpY3Wmy8IU0MEdovCUBd+/zVJ
hZ2F0CETjr/7uaurXnNxRVp4Wp9DZkr6Xawvi3di+8FSu90cmyonH64IUkHSj+v91Z02y+xggU4P
pAmY3OtBXUL2REm8Y73Bt5qXidCGH/ls4UNWRgxalUImJHotJLoSS9Z8IeeyANTn8peIjZNcpj5d
JL8TaA2HVRjIM2lCqduhR+Oo8RgXid6kRoQcApUXZwOOsaFhNsg3ZP/gMQVCCLJZfmeL45c9YMGg
sFglLPR/dWn3Y/HDH1ad717qCXh0hMAOwuE5MOvptu8oT4xb1wMCfWxH6XFw2fGF+4QJPt+kQVDC
5PrEyVZWLQec2hQU0ovkG8lB8DE+30uK6kf99hYM1v71gBiBMYRJ+QOKLqAKXUXVoAS2W+sBz27L
SnZ0yRrgbH17QRdZXDarnAOE9fOIWnbHJg8yeu3gU6qaiqUw2lPKJscJ88U0mZ0XDzf3Vbt9zbw5
JT64zynLAAZPUrCkT9lieJkwAClbfJhATdYmpB6YSm1Z+yKkw206sgQuQq2IynuuE+BGSQJdIbeb
mbQOdJ3LHDLuiZHr9mAjMO/KeRgKbEiFeIIiM0Pk+thjnXKfZmcc/DynRB2wPYG5pZ00YxUCsleq
QVLRTm5GLkjEP6SO1pnbIqUw8caGiMWwSk7DEh88SFjmjnYcr8XdBUHQRdrw8lp+nz4bz0H+bTLt
Cg11tzblqNgjIEidVtgfGdDpoKriQrV1BZJYRFTo+rJBdmxShlgbIWttzyUZeNcpbyz/LiF1zMU4
MOCU8aJXJsBvDQxUt9XqhfwZKSvJlZQzHr9Ohz6QpnKstmHu9wzCnPxd+XweYMZLNRw5BaHQ9rMM
8CIYq9UaVdC35vA0vQZUOfcrDpjpqokwTlU/w9rmLOqIAr+jfwWBDjHlHsKUJEgxma86lC9Hlc3h
Ntd1XGvES8aIvV899aG/gkEUGt+C1Un+ZQelUOLDDw6wG8UT6I0m8O5EfaBn8Kf8/JnaC8shJUKA
WuHcaRzZUxvSTGJh85CM4ANMluV2EmU7+s4JO1ulCmEoyOQxMfYtpPUn+QVdBAg7pHL3aPCmmGHZ
EhSqCWVqvSVWk0uIyk9H55e5WWZpvK48O69ikhcO2xlP3dlN5FdCmyxdOMLXqYsyxuSXlqkMGYie
HoD/Gb8MLOI927oKJ4R1/Zsrgi11d/GlO9ySv9QZ7BQE/zNMmU/vBPf+xPNml70sGJQEH4Hov/Cr
qblvO63SlH67CJz5P9A2Lcz80yyD+ILC9AaYIz3MenxVG1B6SE/+qxWDK9nCZ0+NjS5r33Jkapyg
xl9vaTit3AsGxuIARf8QgXSaIv539RZn4nOQ/BBTy6Bab6mWUcuIcZtDpSlMbAeqCIwsgOsF2fMc
o2qf93zNj652vq5Y2DF8fRT1rIcyLEWewV8q7lhfxI970zmgUFw+TiF+fd47v9aE6/8h0UjtfDiz
bXOBebt5DBibms/Qm34tUaT7TAFtd34Nu42GjnYfa0yAsQyHkYu4eRkt5jFeIaJaF+sBV8SbmkGs
2bpx52gSSUU5YKceRurb5LyxjLuWqzjcC/QMS2pEKFJy+HOisc7073IYBQf3E5Txpzc+Y67CobQW
9sVATsuj2X6/GTlPAb9kYBvQUU1+wczTziAP+92KmVpYUHyg/TrrYJ2j+DGTpRuv7H7a20D0R3Ka
HBcSvAvD3bs3Lmcb+NBw9Js5CwQUewiaT/yLz4rwhjYkmgVcY32eHoZKMwnGf36ryi/OX7B9Dh/C
OmbpvyJ9buuu03HZ1lHZ+iM2xzZFV1njNX6hqRuazZn6MqFwNs8GYW9UNThxmT0EiPboKGyATN0D
ScQMTFPa+BzrA8yaMz7drEKjeA9ZqQ4H1qTkoOyIr5f2o8BXUGllaYafU1ZZyifA+13ciSwmoHJr
tgAJHmzsrt2/z2B5DfnQDP60vHdHSrbjIkhcI2cD0hgDJ/bvlEalH2hbEviHkPHn2SgmNgc3mgcq
xP4cq3JKgQ159trJdI1JmQs/Kh7DIFKlXz2HoZqibu0TNWne60qANGGdgKSxwa35SVNBSDU1HRIX
u5jOuJPFAxSo2qKcOVUFuk2tZDLj0f/UIY0XnrXnfzcmcQXKasJol9gT/jLyBp7jgn8gNfzA0NQz
M8grm/9ah2HZP1R1rQ1z4m+sI0BkTrnGN5yyL6SLwze7SAgDRhyT8dCWLIdYd+HnjBuRsHEZvir/
A1Du8wiLFo5S1EfMbhfTAg2IBJYr27DNyPma1BIGFCrv/mPUAbePD77zMo0E5kzj7SlE0Q0YrYj0
2Xck9tj9qRn9o5WdKOQXdB88oIveB3dpbFsH/N9MXIu4iWWsjjGDm34NCcCvcdSc7PX+w5SZP9rg
zYYo0bua4f74gkbOm/R++u6i6GKj3SXSqaPIIJlPS1YVXcgB8PwNutOr/d6PGnPgIjqgaDuBpYuV
lcBTFPQNOqGn6+0zupQCd0CHtW/eOtfvvgeBZYWj3R9gcGOdp7kNIXSB3wCpo42UD1bJPuMroap/
opSFX1oD2zFYkvfIZTt/xQBRATufvjEwCRG48nwTKGSOhSi0TLtxjC0NEI4RatBjmxwy/+aXBU0R
efM3DYEaTCDzGcdAeBCIlyYRJLznQmpMn7jPzDl85a/lC54SOWxbhaeVPFJ7XcpuvnkqjvOjiSaG
K0uMQteXU38wPB0RswdxJANy85a6L8XTu+EHFtqBZFMIpfaRR4zjyRvqcsHP8bUBDvrKQiQz9zI7
B58zMq+UFZ4ZRzHGDgE0bzgFtZKmYfOL0AxQu90/llG35itKwLQaA1AAB1WUONT7MY9JRfQWmyUZ
7dh7i006hlpYi4oPvH/lbWyNA2Fq7EIYefdyTVvXYtvl0x1V6dSQ8GzGN/Rgb2owrkRIVWtRCMJF
JIlXj/hLzHSJR+wIRAiN1N2t1YgNIXQGbgGvLiUXKRLezmmz4S+4ZQEj4+nY6UxhLpoOQ5OZs76d
BAXBzi8zaNtUilzJq3q7KeL7F7cZknnauOSG/vQIaVgLpM5CMi5LrCt7TW6kp9PLX0bTUcbQ0o8Y
ou4aOuLHyM3BrpF7DaCv9/vYz8S/uE7ehoaR/IsQWoJIz7qtN4Rv2/UqGsfqQonXEQUKrBLTQmkQ
4z/Lcx4BDPca0AP5uWlzqmVoOWEns7qrdOwbmWGrAR/BXITLo3mURHb0xJRqxE1PPjyGjdSA8FFN
Fcbk3PFYJivwj0Wv8+91J3krhTha8o11qOCYFnyXPN+XRY7tGTvkoVILsPmGSpJrDKJ5Q4R+V3ZK
VsoUoUMxw1EWYu8GbgS/9BJrvrWqPqBfWRBBCL+Qeo+iwhmoO5KZi6LYMtqEe3CB0IlG9hlM0AOQ
9hXxxZBINywhufEZxwVtv+ItzL5Zy7xbDrXkNFBmVo8VBtu5giOfigiyCBc8XVbF6aOFZmImuibs
Ien9JahaW5M+eqRxtkDjneNzyScHXSjxUfA/en7XKICaPPO4ajMrIx7hA5EoiN1Gs/gveJtxNfGM
LweTJiwECCTTaSEyIP7H3FBSSw7a4BdibTPS20AopT74ILYXIxcoJcyf4T7gVO9ENW32Nf1Arlsx
Rg5Wq6j1v1GnlAqpSy7mIYYoHHeQf8EaEqu9oAhwCS01LGWMaIv1w8k5REPxxyANA+yEvdzGySV+
PsrHvjl3GYGkQ5ae+8g0a4Wp3+PolnMcVKMDS02z8veTMPB3brhVxwwkUyhWxM8o/X+h5vCcKZbJ
FmwXfWS+3vQCq0Fga42crUNfYQ633PzcXG3/hSpNq0yAuLh8XtJ3Pe6NIQEoWfeYza4ouzxi5iXF
0CTRAWn+Br+BmAHDSI2PaxYQOD7VH26rJ1bIGYekl+vGly3nxnGmuVoYIt0avgM3FsKtoPB1LQIf
VGdw/sz5odBk8y2JkAgz7HikmAa9GwIadbA4Wuj7YfYdnHcTCvBwWE5EfQOTpmu7cw8Ycbm7dlBR
kb2QHkjfeiESSpUZtRsbsB3TTPn85A8YshKuZgs8N8q93XM7vajcy6mU0smE9rd0r5VlsltaHLjY
xNACxIlVuAney8WdV3VqvROQjf0zClhX0leaCpfOd9H6shpbu9cg6ZwG5i/3bHoErsQyGNVL0lIZ
W/xahqScHDsYGKvJyBkwvgzeXdAEYzHvztbtrErmI19/7cHIuLYWxcOnBggw0jkIfi+PpAPQDvb/
OYP2GE1e9T3JjN02T+CKerdIKjAQPEj7DU96W7TDKcWHO6s0TQKcQjeKQYrW7sCFBUtG+Y4D8WMa
7xSjq57JcE/269tndghaX5G2rMFhK9ixkmXaO68DNuTOpZzDf+iIxUNL2gnzBmtbcrnSCEu4MCKZ
YYWA1CK8Kxoy7/TZvzfoFv2LapMDq6q9ylVYzHKRVFg8Ngxvo94csXAujaMkw0H9oIjOH1BzCOBT
fIv/3Q7P72i4cuuP0/mTOqYo9LcbPZ0njo18+rgJ6eSh7nNT1wTX1Evjh9+Ij5dS1HlshVUlgZRE
MncTHvmbFIq83NsJRmCLL4tHWKmk96STGxk3uQ8yvZB0nTQxaCrTFcNgIzF4kl2ARXpEC5wjXcK5
Cx1BzUpCpawrri7wKZoeLZhg72bHd9DG8aFwxU1fjBZ7/rqOcV2mcouGTWx/7NcPjcLaRT+zG6e4
FXGfRByu7Gs/T5cECEHodeGNcZOIMeQS5T1DKLjL3gCBh91/5ozqbvTqTIJgtIhneg0YjfUSqi02
eFUeaubL6RNmp7VKtwH1TGPUmTkxa8XBcr+lcoypIeSqcUkdm++HnjnllIeHOxiUKVaruvq1tqfL
s9cwmtFFhLjRRrH7HFhJCkrcya9M2gtvwwzuvnep/Sks8mtDyr6ICWlOSYZTcD8YSxLz0mUuuCpp
9AvcNkhJWsNb1q/rQQSZ0c3vg9/SkjnffYhrv0CdxHmT0Pi5heYw0xD661VPpDhDg5qI6iGbOMBr
Xbmy3VCxjQu3UV6CB3HlSTX/+JGN7C/bqKYMpboMmVabM24MOSVXu+b+uUjJ7N0iUTfgghG9d9mv
nAhqmz3m3wYve9XSHY7tA9AM20+OD/e+1PXLYS1ivCnfcJNbxwqQGyQRB5ruyo1ABr5wU5sd90gv
YRr6mB/yzgYt5RSu8Sfdos9LA3Cfh9yUntBcDKR8JvaFtmcOYVeTj1IwW6JfpeIWQkQQNFgFgwDF
psYN12gbgnrhUTQvsu8+ZYOrpxSXrOxC8kdMjWyEVzvKJ2UV5YTjvzKNd6gZIcFJ1XwwtDNMgjit
56kdtW3Ii2ZhQJleXRrjrlkJKtd7ymnFNQtHwu221oxU3BHBp8A4JJD6LRTsYN36Nm9prFcb8A/I
nunTk0hL3RvymvYKZGmINv8gaixx0iziFkh0/yBh7nemrT0DgHb3ICbFx1YlK9wCxtusplkcd1rt
v+rGo7/+j/1WZAOHV+/O/sbBL48PsFSkM135CPWpfML4we5Q5wlrOfiHBLbR+iSQ//L1xD73oMgE
fgUpLfgXipzYQeNoNGn49EX3uSf1JPR0mVb81zGNfR1VCF3FjDqnmR7cl9VgygdoFE/Mq2dHx1Xx
Nd396rzXZbAW8HAcvB2mPQm9pOw8XOpGpnboju1XDEkj3p/LxQVcwoQPlVhW0qtz/EfjI31AKt+i
+ru5fwPSPio4XZk3nFc/wfJ4FT4R6Za8oIeGcj9M/9isZa8ulPqb47lnEpaJGiPyQ1iC1MRY8w5R
WHZgGQtQLbfmbrHP2fog0Kg4BIghizqx+XM2YnmyWdYDn7f1JEuJ5ORvn3KCbVDyl2P9ydN0tqkQ
67Lp0t6CiHnUwN5SqjhPw9PE6Xiw/4C40RZnc2TSL+LTkbIxwO0yE6X4TuNKZ36Nf8jOMDC89qI9
HP10oXCO8IgFdbiE7CQqUKL8cVyCxtNRVxOKKB/Ygenz04qOAMWd/cYTuHXWTl4VY8xZx0i6skhx
dnfzkumBgYVQMZ+o5F9sbEpPoBqrOa94aHduj6fiByC+inmugc0+et6ntD61oNk+89gpN9hTECAS
wg7vfp85PEWGJSU9djA5SzQwcUe5FVDI9EztWYZTJIDrOKR91BSPx4bLnIOdX/UpyqCXNTF5YUYN
LoL+ZpefqsPpaY0krnNln+thGP8+VxtN1p17qv+Z2QPRO+4s7pZyQqIsBdxKr0btDdJLOy+iIqie
h2PjmNcl3DeEEKv1SCqTz3jYK0jx9D2z+BgE6nRIg2i1c82Gii1hvaBDLi7vM/R8QYOmUimtZkaq
Vw2xDMkZpNy+BW5lZAPim66y+EDwzegZ4mHzAZP0kYmeMyBnkT3ObK1iUPwHedo0Q4rwXqp5h2Df
bGyr2TIYQq2lPYE0+o/oAHTYcS9c7fh3+6AdosRBBWSL/TRvbtduplj1gMdf9APMVMXrY6qUVOJG
YkiwHfx4DuTKONTY9mSE6DcK9OhvbwQprM1/525wOKLQY40g4Ekz73TCrcETgoA/LvF+QbdysgLi
On263yMP2VDe6c/jnxAis2UDHnlJQAzEQZwBD3MnRpnXVbM3q8N8Ar4xmKxQfG3XMVNV6j1w48f6
z7kMPY6a1602rKydo3iOqxGgIGjELqEO5pzXxOstEHhLsp0kn+mloe2O9+W0k2hm7MzUSjW6dH7o
cpQEm/DZ6aimBvjp/MbcldNyb/YRsaVTSUF7SoibMywqgbemGGEw7Y9cewrN7wBn+zRFe9EvFcWQ
VW1j1n4R/QWkujoE4lLYUHEnC3JkvcaFf/b0DeGSFsW6W+3wDaRnKxw8sez6HhulyJdDOzhDt7F/
JcL5sKyRZIhYjq9RUpsKBrmg86oF2jj/0leQjUTgeIgqxQY3yuoJElF8RFzYl3YIQi9hviJPaJkx
xVq1shdld+UgOWNfvkVaf74gScNXccvrMgJYL2q4psVbBi+3+WulVYAyg1QlBPaRXaIFfrn3zxfB
jugMUhpUXQ+RaKoVAaEYMAb6xQr2iob07wlx8fP0+mTESeC2e3Q1A8F/4dktIo0X8ji1eCbNRCze
VcDiIT0Jn+rmZ3yFjUdQuTx6uLj5UZ+pa8Vg2Zb6wx6gL6xnPSsqoU3jlsUN9BuqcB7ulW0ap01e
hMqcorDfoamzLIsVo0b2tnSOfXl9N2741hvr4kDzS6AHWVkRNdCfz9mrfAhfInJ1kpx3TX8ipzn9
7OZ3RMjM4j6b953geBGCgNE85uH1JdQt4v4C1Un0eiRTs4rmyx+CN00+6Rdgx9FcppA1AljdIkEU
EDTj1bI790cz6WAQsquyqJuubRr1kJoBeLnhwGTxgizVKc/9NA6xRQySH7aPQqiTLAU1UhzD1Jkm
yazXDUCRBxe/CHyIoHqFzgigv8I+QCOHZo2vsIhvtosE70LCQfhXeO+ft8gvY4Vc510AJKfxuIRB
IXkaUatE73tO31siWYSQ4oepuCm4U/bPae9g210QeyXfVgn0n2MrN8AafL7bWoHrIqcGo0QjLfdp
+6v3nuiqtrLaJukUmN6WF7117TtYWO1mxcuQerlk8GonAqatEHzhAsBaVv5xjOzrBUMboovpaGYB
ChnB6iy8942ijyz3ouAVKmMxwk1mUYBK7mNKfW8HFPKOAJfHDCXTwUO9gkYjrZ8gxGIUtV6Xg4j5
IY55xtpNB/czJOLegAu7bGkAXcoekdJYEoQ4HOYpBHl6tqtOtV5arsDttgGVCY/MP5BMgE3N8xVV
Vpn5qhwFQ+AqOBvYUBMMnw2r/flA5vHK5G8JkNW4vCbaLLaF/92OUTVaOpsxF6zPO4aHGjCGVchO
rFwc56o8Yl+c6A+ID2EXi62BIkKTu8fBgKuoH7YA5Ziga8k/uJ5liYZ8ENgi/DvcCDzvxT566yEV
ME9vpbALJyj5zV3MW+H+3I6BHaHS0HaBf97Ujr0oyPMzug2XVCFeA9r1FuJ8mzqWsJjEcVcg9LqQ
Sj9fTVxUCtCqwkrZX6M5Uv6mEnwK6HLbgaENHXfT6NS1kZZUFvCIcDZ3+Vx9YTkcqh7R46VzN3DW
LXDyqrAlMqW4lEPAY9fk/1rYpagxlSwd5lbxVSiGRHQNLN1x1LJlbjY6bsvAdAJEDN2VdWUOvFN+
GzeeT2oZdis7BwpDqnSqJhEyVdXptsq3bBLRSPoG7FCmt9OYGPBS3tNoLO5N1ZSDqqlF9SkqzzuE
YsV9OF04MK/Mc90IAQTEOkVNlhOOzyBC7xXuA/pbmgfxEeTcXiuiOcLs/9Q9HGCbLzZyuVMy+QkO
xeVWxlmE6m4PMWdPGMNsj/0N1OuWU5yzXhwvcJ91307iZAApQ0spY1FQiNsIe5R/6ccXPJ/S/HLG
Qj7eSErtkyZkNyGOer0B7mtimPD3vcCJkESv42sm/u7xnoZiawqKoCB8WmYFWceehpwtZuQU8Om9
BFAD31hnMKysVm8n1hzxSir0hmOxRJVAIAmuZmudkNOPxRcZNLyUO0nNRGNipS7v/2EQlOj1CJqc
9+rHlJog5/99vtNiB8dUfJMtGKXu2N4IHiB7NJmOZlA340VdqsudmkwtA3Yiy7dxvpVxXcYNlFx+
Rdv2htFS2wJHi0TIWx3GiQqtN16a5uC8TD+XapqANCXbebfRXm9MKhPafihrfUNAYfxNJo6MD+vh
CXpQyK2vaVVsKcEmVnaOrnOtCMUv+UAFZ/b/4+FUOfCchIHWYCitOh59z13cc2N9Qc560/ThPd97
lLgqO7BblgsfXCO6mK+Tvz+cZy1OWLeYoKN4THLQGSKEF1AHPrPudTbAu5YZ3maMMc32Xb2DJnsz
ABqtpP1FXbTDoE+Q3tP5wOozCPdu3w5O7NL3/PDJlcZsQnMiin3aRvsCTW6HbuHhRM2FrVbMnEyT
E+fOYQILHJkRiPPamGfZ9jJsv44t5s1VDhjztfIFCUBxZewy6+JeYQ4wTWB7nktphMrduZqptvEm
ICU6aZBIFTEnpZf9p4S6G1vq+fLIpu7V1Bm9fgfDs2b280mhar5scLOMj1bTRxdDT2Gz8z+oAP/1
NzA6juW9t10CPVQSLf6Nh913Y9nkOFmVLrmRwDQlkWE49hsigY6EFpC7HdV0FYALzWQtG93ixgcv
KOt6WU1dO6bD4jb/d1pjKA2LKqKNpl1Cmll4pWliiJFi0t8JSbYitVbvnV0UDYCczKTBnj+jK/Xl
PMupFjqtlpmJaKDUlwwm5a3/ZOfhvqDD3PHOzmBAtJulflc3wq/S0Soa9+Luud/3L5sVwYlR3UDl
hKIqrT3SazjWBHycteb8GOgFyQY+tj9OW3FFhYe8/7utbTnxV0XNS+NPYg+47SUbhIaRKB+sEc0p
076/Ov94NOxnWndnLzZOHqDiVGjKvGABt8HFYuwpNd9ZnNIOFna2yNuwf/9U20DTc9wlS0B+7wFh
OXCA08UCGLN7dCO+JCBhobEZ67orWMVH4nQ7/nVJgtVN0IvXL+XVZQgcQM6Qr2F/vK3dRxD1SJRp
GIua4gbPa2uJ4BpXcAjriBKPRERfeDzMB82tvpZvZ6Tp5TFlsaBIIzol7zVsR6LRDagjDJr5GiLq
hLEADVS8Z6PFooLfCo2pzIrXSEOjwumus3GXRNn8WFSiPSiSFT/bPYii5PUpK4j3kOUTIfseGihK
6Xobt95lLq2+LzI5tG9FaW1uiw1MudAb01KvmX9QDcArRbF7xdnCJk5hBcj7cVVxevpfz0ro5rUd
9hY354zAb5lRie/t92NzDOkX7orAWf7LfGeq5W76acvnv8AfW9lQNBBITHZ74ZU3XjXC4mp0VbLD
IaaDHWW9L9+iFH6i9vyhRRDUh2KvHqqW91iQVxtNJLYrjdSAmBwjK6Td7kvAISYhcbDesFrEs6zQ
qyu58KpFWbfU7abk14T811Z7d6wi2h1DrKZoxxXmNXjTaQjC6cLdneWAjPFz6OYImnhHCaJ2kSWP
9a30YP1zYkEqs2o+vQV5nG6VqXygdn51HmdSXunJ4hehhCW/ZUsSy8/n4TPG2ThYa051N7u0DP0D
2Gg++9CruEpXUlHWJ1/WiUiG43NUEXCyU0j594ugjrlDj12ukmF8QKE8pKQsLLpf1gPqIdWqCsq8
4FIWlrRnH8aJm2VGFKUSchvQ1RMnZJ8B/IkWID+7KBqNNOVAOtUnTwEtXL87TjwAMDcoiEYoj9r1
Ssu1kZnEFg3Z/i9Rmr4u1J3hyDz9t8dUWbYavkDEBYmVmf7d47sPBYrMMxGz4Jyso8KC7mw/QH/Y
7YFT3AG0GpGLfihCVAmMJQIXG17R0IQWOfCEfjoI5P/YxxhUK+pg5aphQtLCAPRI64e3CB7UOB5P
swSBGlSOIZ/3uXnc+vQ/qdmZzdp/sIYp5QCvEYSku1i8cHbgUGNd3qQF4SbFu8ynQIeOdaiHXMLh
7+6BNXRQ4Fei6rfzb+MCpPcZuwgnI60iUb5HRfuJ3TIti0GxonLVsklfV+BI2lydxwUaOdd+Y7w0
1y+t8Tzvn/VSnu61fX2n3DGyqFIkygNR+wwvdZYYANkcr6zAF1/9GuF6rp7GoG7JwpncjmmJojad
wLrhgtDFR6ChH4rBplhURjTB2Z5sZenx1X0oK1K4bt89W7e5Jv1FTegUhzUsg1oSFfGGzs8Rv59Z
JCFZGGg87zoLl8dajxFzGKTgB1yovg8RYTVwlO3VTMoLIVpPls4EEkaJC3H6D1fgmtlqvGsZgGA5
kqieWvV9vUc1kHGfXKKlo6Iv7irUQ3e6dkeuRwbqFTCI7EH6nu1t1a45L5eT4asfmxf8sKn0sdgN
j6wWN2KKy+B9Ntgn4ALqWrFm3Z/GIlm77vxgj8W7FcQpMSpZ9EZVP4LzhwxD2plZeWyFV4srqXSX
uHj6+3oA0iZTTh8v6g1MXbwzJhb1dUtcW8WAczpbzfRH+MvkqRvipCaHzMvgmThSCqlKVrDgtgaZ
HtJWpA3pChiYIJqEhGhIbbYGXNj5gq6nuf9kRkirUFB2p7ryL4GTvnDaKic6weP2jVJGOQHY54iK
Ap8/VmOeB/W5f2uv8uFSITA4m32wgEETzQptJKXrD1fsaLnTuaBv9C/ZtXmXe3WQ/kKBILmv0Lqe
nbUm6RZgvE9SCKm7Y5Googodf+q2NeItVcuJ5daLw7k6Sc2B5DXal8B42pdbCrKZinR6TUocH3OP
9e5ZMNVuI7qC0QheEZnGLBHe+9NtxP4JBY9Z/hLBzYVQC8KVxQuy27G1IyzIp8tbmWQ6XoKTyDRB
phbGXSMsK03sTK7r3QzzM3oNAmvF2WXlYidkEAuSGKGvMS0wXvicEZ/cek7u4W4Y5GwaleBM20+X
t+kQVTJFXe+JmyzMoasHq6UMmvDQCJmBbJn0mVbDMFYihCI9/rrfkkQ3KT4NwODoxMpMIj5+W+Ia
ZeqLX/0IYqu8lbtViul4NMuDlWbKXX0UFme+pFB87WuzsLDcu661L9Hx8Vwe52Go66qOmjxUt/VO
N7vwlKPVg79nBHUuGr0iK5xZjlu6GsG8zU8/R31Uh7er3hJ+UUqRqtirdEi9fAXo2imSQcDpcOya
YKb7aeKDulJYXd2S/xh9kGyPBc8Xg38ACHaViqWJ7GmE4vQgIwrj0Lmkkg2H0JyW3fKasB6Bl1zU
6x/52qzcCkfK92RCLERmc/zM0wN9djEKztwFaa8KXExJB5UifJ/hzLyAXWgncwUStfsmqvju3UMc
zFf9PgBtZjx/YEbDp5/IUPQbm638roLMiCinjtn3b7OZ8LMvYWREE2v9T3rbJ8OkfccsXkiVZi+v
NhzgOE2aqOqxg441w3jkQqhcBWxXrmdyFMT3AQL9EuE3P1TOADf9E51Tr0J13gjiDzboE+e1DZza
VnypfwrcE3aqFZiq7haYk9Av/MgdqOaUZSNkwbEnUaA+Tqc7yFfypWOx7AGu/lhOdKXqxekWGvsO
I3C5Odg7FcQ2ItMDHPOCt47rN6jpgXbfd0F89O/HS+zTHDaQgPbHZAdKloHT/uKawR4w1C5u9Eeo
SLX23AU4VRhciGqhwve/IonQOpRQV4UVVihxNijZjsoH/+jqamFWXSFMwwWNCtL+3IYinZPNNbs+
nanXkfsSup6QWvk0nx/PGCpH7x4lBl+uqJehdO7naAp0k03k8VP4VTRK0AW3NvIsYu9Bl9/D9zIs
MvCLgc8UlVSLokIjp7R8/aUE/34avqGAYzMGMzn/ZXOy+jVVGaG1D5XzeJ9XGBsF+KjKmgNl6jMA
4Y666lxH8rhwTcdSR0yJKhUR0t7pjYpARMeya7/4bYuKEsqi8ANuL7yZ5Jd79ktwhK7Oyizs6xI1
/keRkOVY+5kz2F7AWnZygEmFIuG17Bg9cBeCsazuIghgXDirqSWqUteznreJ/Il/i3Mu5zOOYMHh
Wlfz9+qF5FFCx6Q/kDvUM3otJaljP+JfxNjS753eFURJAEovvdI+bStuXfrwpg3lSj1jKtB5JmWN
VtLL3jBcLz0+TzNwk0ycYwM/g9pNoyWnv5tvESQL9CbcSZgOdXhpmA6XaA6i2dywnK8ramr+eRqF
x2ioMe1zhzzILxJTQpuzWygpnlugEUvuEFTYnZuhtt50VvtxhoQxEJAVy6aXOVYJFYgv/j5Hy80A
SnJYiWycLQWpcbb6FTrGjp4j32qW/SXNs0S9bLiNjXuoRw/nTPk23pl0z1Uwg9cFYKHEWlvEsvVj
va/CZRYD/cRdg1RP2d+YZ/m6ksi02OAL/MmGicOfwQG9zGB1gEcLu8ucpigPzgoRPIE0/IDEL5wj
rVDfvCXmAM+MIld/KClbhNnSwsJdOdyNkoG3SqtERynV0W8khxhvFnaxi5HJM6Abr2zTYUAPFPNj
XCOuqmFy/UT7WBxcc3J+YjXilBgwwPirg7pPZnALVnE9i5eu6A1a3+2pbZ9+dbtFU6zfMVB4/Czr
CYC4Fk1/Qm6W3RLlgY2tn3dtQfeKZIdKg4mTFr+BW2LzVY4C/InWuh4N3ZgRiUJRdQhLIJGlILzh
1eJsuQEf2BYlHY/qgN2x+c9bN02BLBeW1FM/WGcnGd+6vP1pT55BAAho+Eik2laYbW9o+VvQdRyU
T+LudUH08tmB3FwKZfIOAXUMpNUwKeHaiYIgv5QoJRykTwvKWl3Qkq84iFX6Qe2xWWGAXLgDxNyg
LChE4PF9Le7jIuEO/hqH56PMmOpN1nI+Mtb93hwrVipUn5kSsTPiWt0OwamDMmbkRDSWUPgoRb3l
K0uG3+XX2lxNY267BogOqobMGugIjtsYUX0z2h6dXFn4+xtlDMNVX/dm8j1XN6d8OqJpy8i+bLIC
2Auy9LE2oO0Ou1jGlTlwPdX02/f9ydhxUmIM/cE2CYgdNxAi3+VJDP7HwNZjRfoV8U1VEX9BOzbb
zAG3VCYngP8p0z73Y/i45BbtNFxN3t4Ds4auFCvHdyz41J9Vldt3SzpFAX2wR2dJtFNSXAqKK830
Zgwm3FO8HBanYJ7anmn3KT/pc47ZBynQdZVl87dCf03bBWuqeiQ/uYon3YKJ15l9hrHVKwBqiCaA
L5zZzs1R0BWtZ/3t8iW/b8/FwN/h4WuU4boN8KKQ2gO3bnkCWnUVGbYSs4sA/GU5X5Gzq545yCdV
bZ+vu8K5BLoQSn1n9WWGS01GHugk5RwNVVgVlxRaCh6lV/+/S0jn7Nt5Hq7NMq1JfnpHOXHLKgT9
L2tZwzbuqI+QqtSdhBp6q2gilYsWWP3vtR3p2oMQb3tzMO2hZPLDu+t7FdDlzzPVdBjWepQTDwGB
vYyEYGAYhnFvStwDb5XjkLj8vgU1mibv+NWcuYBj3Q1QQggH8VV9yvLl4QJ53l+JIjC/DWVMh52z
7IGT7kinIoDTFV/Rz/5acMvsscso+Plsc8q2I/Xg26GfYeZRuNdEwP6zQYq+RVpP4rq4wKYBal8x
4ZhAZ4o3ZKkBKSGmyNfoNKsWBHRPNES0Z+CgAtDu8nvVAcpx+U+4Xpe38hsOfWecceRM6iUa/7O2
/NJlnFjrFfrgOQ7Q0DzEDRKFxGzUOgyRyG1XuWGq+gKeBwH7xAsZ5i+GJ1Ks3sz2D6FWvBlQ+jjf
ALkJqYaI8yV2MuV+iOk7EFTHra0sbd9J+SqJ34ZUg8sAUxiCj7jzawEvNXAEPNqqlX0PQCNqaj4o
AVqvjGG2xl/CU/ZgiPnhLQSP1cpx0FD5tx5/L8mdEHN4d0YzpbLDIrLrO3zcMoYeWiqFrkKuZ3Zx
5FOjg/1kwvxwi7JPfho31BshY/7l5L2EaPHAOrj5Z3Sz9ZVRz2rX0jQHTCS/KqNVZ+mYOiqc5Ayd
mY8upxlCOUJxEB4845//ZnzPEXkc8psEL59lyaAYpfWFkHu5gqlwQTP2sRHmfhnpfeli4BY5gx9r
cpbbWS7b1qc9A/obUyvbURQECLi+JRB4rdc+JRRLGXqNSU3/TeCyPlxX++vob657vDVymdcze5dR
imPiebJ0GgFPjWpY3nn0pE6TAx1q5dOdQDI+WHTPyaJpp5dV5x0KwJTxU+sswNOEKAo6SYBEv2jE
Pqqrm7SbUYJJ1/ppH0Oi093iLQLWKdUY605Y/ruxRr+khyYWNa3vYtubfmZbeRBneRmWMKOHZVIP
oc1O8QMUXDrZI8hm0O0bhHgRMdffvn5pxBxsjEPL2itrzRSdza2gLIuC+YFKsJ2EZJR1gsaEUsu4
fh34BYtkZO+9/DD8nF2kmbix4RLRt83vHJHkdF2t4r49DHjm8g6lSrmPYWF09xJcmHRWO1zSCJfr
e82GUJxI0/k/f+qRDej+uz8WRU2/mdrj3hiWjELoopUn7dwjyUaptG8GtemAXOgnQ2m6kAL77RrA
BMEAAqE3r5ShoWwK+64DNMTXqrddFxUX7Mn7jUbMnQU8gfWLq/u5xc9AgKZA/pxrio64xj/fyVoe
SBdUAOp9N0K56p9zmiS6NLgvKtWyBA4Kyj54KUSbfSXi4c9KAjYp0yb4EQTOHcX7nr7YXDQFqed9
L3T1qm1SA7jWcd944uRgNj7bCanKhdvaDZRpj6wk9XtTVGBvI5RwgJuD0udAHYRqY9Jb0atdJnXf
hERh6UNGDfUTOBc1IvYHUjiD3nn6QbWYRG3p9bNeoSLAQgzux8kO3tsDyCj9DhV2moQ/sfL9vu77
1sNbTYS/zDQ5anCe97ICiWzyVr8h3owQgmUkWDhZ3Du8WD/Sb85AsraJH+IIwhwHLPSu9FBO/FIt
Tp9DgxWPQ6h0TLX43S+UbWcHIn2tHu3ht44jQJVacmcJPa+bkfnXMz1Zir5a24QjAJG4S2ABB2hl
M1jvtP6bci8r19CYTaNDYjEympUvQD201aCM2rc+zW7CT75hWzWIczDu61ghtEkTKXxFqZzFWKOx
xqwR37pXjX8icSJiukcLSTmlK2Q1v5BQJQYgVyNnX2fbG+5d+veVhwY0zs7xmC0Q26VIiT4Hr/zj
g/nbNndlvmGJ2KnfEVdm8QQMS+kLiF02BPSTwDPCmg5WRk8Vmk0VWhVP4UGJ/fuequs5vZwEalkg
N+gB3MJWvfflWGIG5ypVI4aWMWFrvsTMM+gqwZoPcBRLn49lf6+TMA0c7g6/ioaBunoIR9P8ISfH
rNfVZdMcB4tDq5vam6lscSpeag9cdH8efgvYKOSMZQj2MSQPIlv9APFw/vRuhvmyCHLbox821FQ8
PlZqsZUKtbHvG7O3h54+CjmgnK5UTHiTRboRLRwvb4rgcAyTcVzcWfICViOsT687MzXbuZNPvo1s
57cJzpALqTuUv1mE95vfsqiQVRpotH56Nq6FCQQzJBKCjBghHWdQmdlInA/f0Di+ApikmtkfZbAt
yxrMBRMkbNiDA8Pb497wfgO/Gb5quy5uHeb4Pdb0GhGjHsEXpNrTk1k87AF7aGFuwwoo3L9Ea9n5
qA38WHqXYt1lPgoTHl2pSKs1ls6VMx6ia2BVJsO016ktCy+X//xwzED1JmMj5AEVcSHNKlFiel4v
3uWAvKYKPpXydpgXdqh34+yz6V7qkC4rgnH641iaLc1D9N63m+VMiq4dKc9565RZEwMgi/HRBDSK
MvwXm2bTUkebfYlUbpYejhOxFq3AiwZgICvrw/1WKps3GzUESrSA8fC1+0cef/1M151U0ngwshbu
e2hBaziauDP0xmW+7jnskJ5KqfwTc0OxdvKgvUB4wC1TPfbYFngw0XglywIOt0ED/cGPe9JNXCDB
Yc52y3qU8LBR0/+kAowXmcZ5qZrZX8VMzlcIqf/uiYJqDvtkNPX3ssNZqhhmY2Pe+sI1sIGGGhiZ
ZnCp+V1XYgHVpyfZt85aLVF34tLGPbejxb0/hl5RekL5BDaYW1Y/TioUJc9179yn+qgs1PWeT9rA
uTvFDV2+9kkpAp8cMnXMAJm6QKNc5rfI9pzUKMiuYRE55E1Cq+23sGHje1ZD09SBNM+Q7BfRdnF8
8K4zLLSbXHzV9KU4tNJK6NhBQo2Uj9lbZsM1F3YXL24oGeytIuGvF6a4dh33mqALFsFeH/FRzAXW
adRyv+f31hZufQiCHP5vWnLZZgNYvXDqNRleN8Tno+hC7i6O+ouA9/MpY4pn8JDaRIKQy6q6FOPD
OSYEbu6lgi9iE8xsaeGcPvQH90xARcfWsYvSr3+fef9arXQv79u0zys97O1uj0XUroke6T6F1LjQ
Xk55Uo0i5DlfzsgJaKxgmCGuAHfnr31shJLo/P8dCF+ICYB6Noltk6lyP3VmGRi8RL1vJ0uaDhWr
OJweHsTYHZR0MsuDqrA1iw6hWuZ1R614og5pM/es6z4jBxwJZrC2WwzYnQNZ92kZwG6lGCtq6ibA
AKK2E/bzRmgcVOjoXfJVz9yyDV36+gJoNL4g9lzIGwhhYFz8yllplQfBJs/nODmrR3NNMx9//Mwv
lCTaSZTkLyGXf4HQOoEyKWLu2r5pGyNtWWoVYQa9n9ivO4V7dozHm4J9TzizGEf3qtjpiIfkMKhb
yBUQyiwrwMQQ2RY05Z4bEXgCWnwNoVXMZJRVw5Vkka7/kwHocZOhI5pix9Wq/G2cqo1tnFrWAvJK
W2912eAbOy1yfMMgygYzTl3a/c+l66AdlbRNXs5eXHwMHFhWRZ9drAtJZwUIyOT4tcIN6C++Xr42
zocFV7/RcgbAbO2OC+DllLORjWsmweaXYzMpytEculw2x26scHOnlGncNtwHphYPG2+fnvhQ/JCB
I7xtbBss64j+qLP0dqE69B+cVrTcLX8F6X9aquSigCUh2L2fKksS2CU/RVDNaYjYVruIo/KOZLg0
4npeE8Jg3dqo28bPWWMDm7WfpgOvSISVhSMlYWWe96/fbTtkIz/PQs6+RJcPyoeN6VZzoJAbHk8v
GZBIF82O+UB5D+RLY/USabaVt5Q6WB06lqqCBhrsSQe05PUDzvOZX+RN27g2bZixyjkOhVspN8eH
MeOnOUxVSZBZb/0F9VOAZkuElkc4buHVr1zfRfqAF7gfIET/g/tULthxcJaVREfSgXJQwonG4WbU
1VyXUhiCgeLuM+wziQxK8bA0r6PA65ARrRt0P8fcsQzQ/ZdLTyRC1VSv4LN7P3ZINZHuKbJTFkJ+
U64Zv/QsAHrKR+osjvy7b0qPBBHJkBw5xdNMk6OVzHlepBhMtdlii29UCs5pLhQL3zu6D3JIDGpV
jA6NPaD0mR20HyiIWNtKhNnunNLPLg1MMYDh51MviTQtDG2U1HNoPQTdivcqSsKe2q4t/XKDQQZX
WZu5RW3Q68jZlEjRX0CvDyaXQCTYu7SU81Pgm3vt1KZLWXeMmv7cArn1dcQoqloTt72Cwhc3q57P
XbhPytRhpCyv7fpmtLTQfdYOe/iga/of2RIT/P6pCY0JYr1lgdqpuNo6udwZzH6MSuSGfv4jK1P7
gQvMyCL9eN2e2XSOX7CY9t4LeSi+103eIHesAmTMWp2cdMHnRWLoS0s6wGfeGbp/EeHahoSe6KzY
ROKo3Ngf0MPFWTex7vfn6UjaOlVcE6pHAbJHfGSRAys3VOB+14EDrvHdlU+Iqrv00u5ITR7S7aBJ
7Qsd05xg8EGEYlEGvYb3XYG4erDZxMAdUiTURvFsOlQzn7Aon6Wthwm+uLKQ+uCizlQxRgAPcNkv
ThjEl3ooAfWJTsA4Ri/P3oS0iNzZUNpqMe0WIgv6ndnVxCxSZZbnA0nESEDfSbvI8O+FTKJWKj63
tsQFpm7E4cvnSqbE5/8N8KPMc3enXDkYiZfajScwy9Ly9QvLgcLYBj0moxxTdlHMXW6r4RNoJcUu
ei6D8U8nTekmsfJVSwikodeKo5etJxLkTaQhmx6UTouAE5e/r8EVAoln/87sgsF8a1lo0vH3aFrD
2MC4zCRbGf7LOIsmmaBW0UZ0UCSHMT3GGKiJJeNmp51q649uGvJnzaW5vgz/VhglbTRIjVc6k4P5
HA4Ph6UCx2xDVhyheXen7NS+aopUUZXu65Q0jD8OZgOrDL4DGlQNt0gUT0pEX4flsSfNEDyklghd
uP2xTH3h6oxrj3lLUJ7N1YV+cfEMiCIM0k/1MjwAgcR7HtM+3mpAMNQgdsnfk88Drh2TjJuSVsxm
FRJ3B4GqbiaqIWANX7EpVp1k+jg2o3zaVD2MGpMUdFDy1ZwCbG3iVnX1J0OjHGG9ZBgFA7bMy909
2ykZ5/fP5Uu7scf4lawgGYZiDYiXCyN4O8uc/L9JMEKJyKTy4JTCVnDYhuuIv5MV0jnehV8M5NZZ
rCx8Kni2lndab37YqAo0TAbU8GHeyR37KvBTUa5sviPYaGaG8kylqr+mNYI4/vGAd75/yLFQVjmG
lcan0laFPY4+UmffyPySODVPtNhzs97u75rVoTrKO2EHySg5mv3Pc3/VaMKDOWwKyIJA8Otu1tPD
q6PvQfGY5ASf7M1SUg3ZvgxneMspsZCdHbh2C7jNr/wc/Af5kHz2CVYLhsJRldbHwz+IROmV9ZRU
rKx0NRrst73B8MOZhcJfCTI/51G7OYpA970129l0cPRuLMCnmVpaVxmm/sQv3i+Ssnjxj5hdnTtt
x+lCJBioUcw4Y3HWnzOpbkd8DqwT5/KN0ykHg5r4qzJxIuC4Viu6ewxg+l4vpbAXpGCyZ0oLi3Qd
4Og0dv+Qif336GIx9+MT7kd2Gs9FRfQuKYgtzNuz9E9iz+4Cyyge//y4sbM6lHA0TLQ0rrn29nCZ
WBX1j1MakdTz0s8TSGJ/9TNos/y7aXoMlR2lSrVZmCBlCSc4st/dmNb6opJMP7hrqcSvcPe5lQ28
J4UQ6M1CAQJvLmalxn1K1zZiiw2lq4NgBy6GZlhiQshN4btLk0NbmGEt4qruVib00E4JHF7uOZ3c
x/AvgWKclbuYTo7ldRdhhjKowwBbEB33KT2hMJu1EdjpZHLaYWMeNMZkaUCdkDjJA6XZ9bu4dhuM
cAOUE2uAZvehqG9rhfHXwOFKY4H2hw6pL6OaCKl5juaSSWE0+GNG8sb4qZbB1jddoRaxVSfby4tT
Th1BiEAAcNBfodtkwIDb9/yg+hk1yEvmHAsZLfCuoHwVhrQoRPks1ChktR88LiwF92hB2cvoV1Yd
uIFShH3pO9ksWfuYZcQunfQKq0UVMFIZAs/A3ePlZt1nYyr2Qb/Ng2KRCK7sydOJd1aP/aQcwcfg
oVLnO+4MraC5l9XMYaZy3rk0PpWAo7pSzCiA/mrWADjE58YLSeUXpJy3CFe2F4KAbPbeEMYC0KUy
Js+b1uHmwq5FsSpi1TWUaa1CFcAPorWHnoMNrB/I4MaMsM2W5B27I6DeY9hVxQgcKstvXxi10MQX
zOOCpdPGruo1XLVaBD+UDSorynkV5lx6GXhyBpSu/AgSsPiF6vpTVsM9Z46KocFSkuqYU2ab5M6R
Mu6IdKLEQ3Ey80/VMyNO3vgRSiysNFZwKPMLDeeDsN7qs4v7KAFophLTQ52zy4hmyUeqdOKq2qBi
hSfXnyUUbn6jAYLBzg72WJ06ftJCnENGtdUjeLXH+Jq8PVOGXY3jEuTCxtEDf7EXMXydYXduy1Hz
MZqanAp5ZmO9HUnKJDnjlZbSCcoG2DkL1gqhkk2B8mEz7PWJhQ+qe0xDytABMqjJOpfOWrvfZ33E
66Chn+svRH4pT9FhASmPRwXvnzJBDIUA/zysv3t32IGdx59VnbrToD/9OpPbMWoUZLsedQvLciII
UyBm+QaZVCGyvKWvyzzvMq9lRnL7xxquiWhRn/liFjjgpQw0H0Prxsr6ESh0qGgwYyayWoRLz1hd
ttPPXHTYqcg6IPpvzkFPH4WLleoGyAIyjFc2CnDWyJq97mjT3ooh57O61HClAIRytsE9mBsLkL1n
noIOpOkjHE4YDPvBei+XNu3vFkhISVB+nkcjCv+K3jA2MWwGIoTvn3PTV46KC9tZjB4RFyqxPD6O
idV3vU/upHyITr+bpR0fzufp070j/OfMwn4qd4XNbF6t6wUPi2NY8+XszRgoIL9V1qgJjEep5Bbt
esEtUvvZrcQRj45ARHZuuOP68R9QMfJkaL7ROTHzPpaKQhaMhjQZW94YSGXsz8go39P/HKfeNLv4
oOD9PxI6eAmxYyt9AayK55OsUVj2o6sGt8XG4/y4c27znMXPq2OMtLQZerE/NqmO8VhWbvyHJ8rB
Zdwa15BxpwNK+8+7z0Vht+vym/miiB2ykvQYA4Jx4xfY9pCb6ojvOdiXnbcOOdYbi3RA51C1ReVD
c+Mr7XLSV8fW3mYgQU3ia8U80czQ2H+c4zVCf+IbCWrbS4xsC74WOX3WaNs/vwmcDNeoRdl/2ogm
0hE1Y/RgUQopJXKEl+ZESckIrUKewQMwMZDLQDX/QITn6DFF5pAPVhAxSHl/2updmjnhcNMvsOYi
7X9qRWakrmWg89Q37U6C8HY2Vx5GYJlDMEXDYOtHva72bojv1fEmk9yGfdny6JQ7dTlMkLAzbcOU
0u4XhGWMM6BSomQYoJ8wZxg4fVAm/fbXypkyuvlAYizSbwDNyrMS4tm5UfxRotnd06YZ0uWxF+nJ
qj40JkAz3pW3KVrmptvUVjV5j25ZBJZEOILX7D1UR0ahzBQVz4podyNSh1P8G1P0fAiik+NxQIGb
LLIcAS4Eq6oKumIC25SEDeo7kcWUDPsdPl5sWj1kQoBvRQwn0NKO0UxTNLuKSbALd0wHVW8tk0Uh
mnOMPvca7NkF3HIiC0U5fqAHyz9li+OyYtbVtjuUnUI7j3ktBNVLtK8ZGk4uHHTEY/P4oxO8k8K7
6gu8UgwohhEhvdE1R4XcPO3ZJzh4mI/TQJWdCPo58JBXd1RztE3ISYj7OfeFWRr3zIQNk8nikASx
jZTlsRdpNMD1giHHt4b5sxy/UfADwdTIZrI/Mr+qxeRBd9SXDNnFBP0mKpCIC+xWUu287rzE9AtC
egyQPYLe3lSbotV2iawYSpiJhxyggRTE2TM2lm36eEFuFtHYzDxcFAfqJ5M9z8hk3ZDBJAmfFcKI
GXZZTrCr54a6HXI24sRqt2ugO+pQ8zdZesZUrSI+TvMgqJ+vyxWDpdiyablkU1hXB/t0kekv+JPo
sBhLgdG3AuDNUI7bVGX+GH9xRUF80sXloUCEKQV+Q1Y63lDNSHXZKzDHxSJHybc7jjkoLcsQiiaw
RtRdYD6SgzYUN1zWnnM+jB2l+MvKwA7Pv6orYLhDSbc4UdxoBKezwA52XnZz/8sCTGP+a5DCQAx5
tQLFQKi9b0MyLIk6PM9AHjcSH1Pn9aSMSm9wigh4Cgctw/LVF4bs8svxOgFfHP7QN9FVPeozynxH
5kqeXNqRbkR+APD5NpPtO//de6mItzKEoAm16yV1bmFnX7btXDNsPBUd60PemFZ2EtnBCYds16mS
jcJNabzCGCMfh/vk/V6BqiPBKA1UOJU5Hn2wJ3G+6+0iPuBjZkfJPtmlAiCN24oxZmBt7eha8RCq
el8Ep1+ZOFOklAwHyLo4DoVNhfFfScD5wFLOf5jECG+W5BpSjq7MEB2H8wjqack78tXJeLJtQNA0
2JfizgyUyl+NRAkqM+rQX0PTnh1i5hOIxCcFxnMW+GPS8resG8wzIvaSslIBdHyDYmuchh4vZFoX
nw1UxV6DGYF5oRQ8BzIvNp/Digp+XDERQ3ZNVLGVlmiNIz0ziFgw14nUwgjC+rNzFZA2VaDjeOjI
rrDcLfALvUmSAxl3o9KWAavBYjkeq3swKnvF5hzFuA5LJ5ngjh2+jQ28EDkAh1Q8VOXZhpMVhi8C
fhp1TnMlW8yLVwufW2b8NO5ACMGtP66W9KRxefr0CrLEMRt9aiuPPXTCC4vWcGOj9liTcPqFUicA
g958HtsmmPaYz6JWMtio4kKFDTfbJ2oCO2o3sOndNWp5zJvuhVbmC1JoTsKl5UWpmEA9RA7v0wCs
h+QtFolvN18ikVIYnETKT2a4YSIexx4Qj+iyhFfZLgnlivzbOb0btt4YnooH3BrPtD39nhAn0C9v
f3SuRV6kWo2uz7DidHg4ob3tgeixkQQhuorXJOvbacxIzeqImA3j78euKNVk2Mhubz/+ll5mwpzi
+jFYeYbp2r0CnMjlu4Ru64ISMCy9O6am6IWxE18iuOIufQxhBgGO5bGWwhNdH64esEcbqInyZOnk
gZGz2oC0saHBVKrX1f9vBdplimDF0Hdk078u1z1PdWC3CA4q3wmqbBiG9Mp+szVZWpaYSOhA4sNo
wm050ToC5WxGUYblqT5MSm//8IVjtXPAk/3VYUqCQYJPLyZF0H3XWrdRgZqZITc5gVMrb5duiaip
JvfJXRDs7UXrXjBtXD16n8249gmjIaZNoLXNxH77Ua1iCWSs6iM3pouNyg+cF2thihr1WOEW/PZP
2PbixxU+PGqrkZopyrJZGQ/t+hkdMPV5hPH/HVXiCAvuGckCo+/W9Mzeg0jiehkctqHdu/1uJwL+
hyFYOQbRCr9VJOU9om2oScK6kqVtbXeXT14mKW1zsdIGZoRSz+5NPPyrG8qZ12okMbLM9maDyB5b
3HAMKhmGuzgWeA39KErhWMyk2KHQkNwcn5R1Wa3/0sHY4hU0rvWuobbslE0MrxZ7xbJ0bAWgCTuq
ISMAcqpCtkqpIr36J8UMAj7uXzOYLMvEKZI40y8DxS5wyg0urRYjFXr97OQ3bc4wRNu1+PIodxPf
kthFpPDzn3xtfqK9FIWOIHoGlslQc5xVpwJQWDRWLOlDRVx6UVJbITdmDxSn9lzlBQcq6UrevbUy
VI+CrPohee0YzDm7XMcLjRQRanogkrY5mt1TydpsU6sF/9jw+ZoB/quHadLHjRYa7efXzQJtZSrb
BQkhjcwCwTQBZI6NUgVPwxEtp4FG+lUVaIUV53HMSgMBEaB21/gBL0yE/GtfxgUxNKo3HCP3sLjV
wt/rZNeSBEg7iIf3y97WnNgFHTGn3+JDywKYqgYJ9dRR9vfF4snXcYl0I1v+Rbbgrhr3i2z/+o6e
q9nxaykWbpVD/EUZezrGfuGwfqkWicZnvTf0teUAjcPGX6zYXXtBWqcA3MTMss22OKb75jIRwud3
ncxz80u+d+sg66fb0IL2mNDSkHYd7nlkb4UqHOO8EK4UkKHvuWG7nZ5U8J7h7BW6/yikaYei4op7
cqE5sI1ZsJ8TrESscnmWyxTTgJHrLPFIfnaW1elrz4CdVMEwzgfYXgKnabmGUeBkgZyb19PMD/yO
CVAizZhZ/zrl75Y7AFiRNeOxf9EUWrWjYV3Y6pNT2h0Fj1vyoxfGHpxRcm8soMFh70O8U0KsaQuA
2vzqY667lALMCEYeedr433cSb2q/6ul0Qz8wOfWQFIHgNYVvBB/ZiBUFMCExN+1YoRgwY4ZLMRH5
4qDXi+X0zN4VvZ1bL52IwUKmkrOUzoB1rBYZEDbOUZG8c7Bmmi9HSmrzRSSKvO1PyEWeYhw+Ppmx
Te/FBpk545X0IR4stlt5IanFlUYmqFlzcAwguI3fEVeYmnFgAXuoEz97T9NwZ2ZlVBD8JrPzbFn4
7r8/2GQCZ+ewb2ipao1fG/hV3NUNTvviPVGdtSRfi+gerSXrcMNfbouLid4bzOgXIzPrSST2omhR
xBDg74kYk3E9t0pDoEyRjWZ7z96tJDPuNBtvGXFwstMni4wpK0/FsYbTuKnofMT9423KPHVpibQg
HUBa3BrFkeH3sTlqNzinCQgfmKHZP2pemNov2Jqm7sFSyPMK8v+oErzA5dbLJghAGWo2iZiPdLVV
8mOOU1CzyTZrUWocbxdEY4TjG/HKr8gFN85GpvDwNmlLxcUi9E3XWxkYIQRkUGTsKB5zreyM3e5j
QkZXe/05N1uI+WIhRtDmwEoith+h6/idBi/dz0Li29nQamxc2BuVWRanCmhlM51u3GqW5uLNRvyy
G9o8hb8oIe3r1xsp1ahi+q0CbTUpiyLiADXl1YRMq4yJLqs0VP/qMdaN7vFZm1NNt0/7SF1AG2iA
HQENw1sVA2Y2i4mcOIgpWcO31GHo18gad+V8ezn+XmoHtb5fDPds+Tp3BY+k3mW4hZa2iTiNOtIT
ESItAC0kEGy5n/PwmVbvnSzN4VGvaeOiQEL/DiqwFqi2I+kC3jN2Q/WXChVIP4qXFrMUxipfHc5S
IZLaHgfwX2cAN1xjs2gDSLwdcjM3ATl0m+LCsJ9enIjSDcdXbyNGxtSHrQm+ukL7fDxrhelWolg0
xszeKeyeEj9ZPcjWpLdt5k0jP3pHP3BpSGjgItwnmtB0xBE52jtLuoB0vl0tqY3ZQasgiyvWq0rP
QNEZQxuqnLG17pROyNlg8y70UrpFWR6rIiqzpBwdHTA3gGM5n3y4DhLtkUcP23oQiWjKAkHXmZ/J
+Bcw3a5q9lc7Ym0qtO0kKGbS04mHxAGMUBI1BYLTZrLdMx7Hye52I2aVrd4zBw+cSh6wNaikLwSo
VThC7mW33OPBAJACcDBCM6i5LK/l0zaC/84SozbSSi76Kt0US+5sA+FTJpX3dXRh+qbkLGQF3R3I
X9UCeNLOkjbMnj2Oj7z7blrckMqqlyxN/Owv3pYZJxaAdJGzaPqZ/3K9nMobKvqcYfE/YvDxBDMx
thCPMviiku5hSAchMhv5n5fKUTzr8rJYk7D+um7b+PS+E3mTQMBITpOCeKV/BkzQRKyzT9TzfZ3I
kAZzSkTvgVDc/5KeMmCKpzM60shIVVRj8AGHyiO2qC8jR1Dh79Dj4DA9TpoOCCOBXj/Rsz9BVeWQ
sgFPnFmtOENMNywCtuSWPeqbwHQQRUwlyb7rn2uIA4raHT6gIqOcUKHQFEUsdXpjT9ga8lfgTl6S
pVwpvok5kayJMUQdUGHpsFdH8wcuXnY7tPaoJ0OqlYurx29dKIs2Zm0AC4L7iKysHlx9XuGkf99Z
9V3XqPHLO7Avad4yO2HYo7+Jk3aatFp02PY3WQdwn0DSoBkFuqFUWWjwHACZUvPz/CWkdVIGknIt
S5VSVwIm7BEO0VbBy7VzkZGKDQVgHV43oPbOJQmN5LBMag00/1Hs09etR1/eRxBkeHfwOvll3P5g
cnmFQf1vXfh+m6fbHcD2Wi6f11S+LqNod0mB+eG4lt+fDfOkIOdvQeOxugnDSltoAmvG3VMrUq0D
TGDhYKA+y8zbYowNm+Z40RVO8WP5VzIXs0Kkr2O/42RoBfI4pUcWtdZ+dJ1rNnNo4T4kfswiRZM2
Gd87GxMjqWKBAqmxWTdVrQ2p2GNShOHYPy4+1jWg1IC6OP48N6+5dVJM0o1xL0SrjdqqmzyAEq+E
6TkzEzMc9svfdYuCMQX28JKJFGwvL/1YE7M7wHQqNGBdeol/Zdm9rT5uWxs9Ri27vyIJUI17yIlZ
SdwPrtXLmo2RFqtMdLDD3odgy6DhgFu+7/H0+EqxTy3TUWSYwD6hdzi7RQI34Ko8kTMuzFu0r9bV
AV16fStvWUQwNLzrY6lgbJwyxjU0dG44zNC6hFihDVjBDygy7aIbvME9+6C01ixlodPEdJo8FOor
lcnqBnrjTWvllLGDPBYQbs5xj/XOTSECg9y6r/g4kvItHl1NIKHI8o0x7k8RjR/aEZ1wtqQhwq8X
CcPGmyTItIkGfxejYRL+WtpunrKSsiJhh0ImA8wLebCOVzc8YYw6407AIIjrZ9bAiEZbHQ1DwGuh
HnyxJ8TmCLGeRjF7KOVbV6eNGifi7mEpXLfeSaX72ebNP9ZZ1KOp8H/tKNjcrdMPGHGPaeE38OaK
TDO75iFV12kzoQr+uiATPn6CbpIhh8st+YedrigtvDGZ5l/ihN+XaIk8IanEFp4XXFJ0/R5S/TT4
LUeGduPG0DPACWtKPIzXHWCNPUn1Um9QJvRBiJZqSymrritDJ8nPtN/W6xdQC05GzfbFbxjRJ0lo
uOrJriZyduHWAqkIU4ViWGME9lIyvLHpx4ZiYl0ezUTw8C3zwuk5H0CflcBNrWMtIAI5m1qPzeux
bfFIAmTAHECaofwhjI/JNqoArzHRqeGKW+r/Gh08nLMCBV9y6Z3MH7fzr0LgxenaOUwbct5oW5s5
Q1dp7Sk6vvLwJ8/dbPIBbGiE+SRFTNYSVQTo9zlgdezNDi/g7pVXl1P/oEjPc1wxiaOqW/Z0nf+t
9cpnww5pDhaRjIlHVnu3ieo4MVAPYKMVqwNQoBemvoHBbZVjbYZky18a8OvoOPKEJovkcOW+b84V
vNncuT8eH30Zsa6ajBx2ueGO6yJOP/eXIoo65TpiNLmn1x9u9V00yHZEGjcGBaY9bH8WKE+oqsdP
uoGZYuzgQ8akWeSwx+d3R/uFNmnwQnN28NO6+z2USHdS9+zNh057DXgsNT12UlqF7raVoJpSB09F
vxiw0zhQg/t2u9pPUHEHJ/0PW9vd5Wt0ll2DoFxsmo71UHFKXrN1ZTn26V3cWwY30wzW9nd1LD2c
y/5MX0Mqn5Xk4t1gUrkOxJWEaHUv39xcaYjMUQWjUJBBguv8E5GGtnXlnYzwNZLdAyGpO3cBx8FS
1iCmLrU1o084gu8Oz6OTpES7BGGYIhX0sPeGkgDY9yjAuaYtRYK6cuzOFterNosPjLVurETY5S+N
63it2ee4iX1jKWvHR7f9WF48KkwZ+CrF5UPFY/q8V3x6AfQi9JdB1hjCXdl5DAaKiLkYjDXKIw28
wxyUE7HNIGBQ428WI4pMfYth0JHdxfhM8uMq2cELCIJAb8+PXy2ILIGKIE6QjfxfPCk78rq78F7Z
tqyXmWDIrDAanEbY7PEhVGoHA/DrBaH599y32m3VAp/PUG5Xa1qYMDPgoLY5w3xENpjZ/gXokiKC
TLAfprBt+OSJt+Pm/jARpW+zd/K/j2/rM45tsrt/ckAGDURMTSfwJw+1m4aN88J5gmleIGYh5/Sd
rwBYLJF1fYBmZ9aGGFtzlZm8v+EfeHHzMWYS91QB1RJTVutB10xS39tnySbX/5QBoWG4RXrjKG2/
UwN0MpUOVxLvnM91yJL3/jpB83btl7Uo3To1rfQGCUbSS/rQVa0bG79SGFBYTvRxGQRL2CRAuaW4
/zxBtivtmlUmUK+ceecew/+TD2XjFjl4ghGC+71QWJLg58WsCeiMa0NYsx5+shJnyBkVTDv2rCHV
Mc/4EZEay/1/PmlCDxejHrOJ4G4K+/8xHtvUMI7smJQ+lGxT1bTMzDoIPXz3Z+FOT3F3NcbjF/GV
forSutavIqM9izn+utjmUuvPDMMCfBFE289rwwJCifNzyXAyO87RWlafgTldqYYC7BY3BQUU3CvZ
yyEzoAPbwNdRYCOzRB6Wa1eD5LLeHpxTFKCSA3w6vL8kgqkfulPfWxK8NZ28zmOc2122FSt6niiw
vrKqbDYfIz/jwjsdhNWBTyZI/RD35Q5x9ccruNCMgK5QTaw3SE63yYtIgUw4AhNIilWmBB+tzjkF
jsdhM5F5FhmzCig4BkyPJUE7LMsKrXx8ceavpqxJOopVaPNMq91XkyiLxBkckOZlne3tqrzyfaBR
Oms5eo9T4mqIDW/FOGyMy9D2eULYLTFXPGH6dvdLB3+mjS+dmfM9DsKq/vq65Qp46IcFY1Lw10Hc
A3o8R7CfFzMOawtSTHTlnj0mVixMbdEBARd2O4nTgHQz/DBpyVa5KM83gHO6ZudjiuQtBrpqpFd4
zIm2n9wohFwOHsMonkJi2jcEwNnuL/rm+uXV+7CrZrh5NF6/AByQKoDn0zRdSYVXZh1miRTRNlv6
uud64ChO9tLUlmkLUR6tJ8RbGiQgha5uj9aOXsUJ0CSiUWv0Akk/anlS/rOhx5t8JTXBzLBMxgQ7
meZJ1Q29+as9eMRFl/wG2kPnbSBUqVxLeLgQ9yQ1Jj2hLOxpHlrlK+Frs2qs9UNXAjcNzO+VWg/P
2cYDmEFhajFkwjxfbY+22C2bknb9FM7U4hwQzan9ubmYKtLnGaOJSCkVcO6n66k284nieiD9bk1K
TTRLst6p5+mNQfYVvB7p0GbdxofjtVndFgCKJn8Hg70wKK+FOpD47vhfDD0j16aSc9G2CmjZ7tbV
vdMG00IwfBse1JOGPT53dgvPFtxh19Xggz2SGD0BF394rJAWJ8Px5dYC47CtZ4P5pnG09JKLr0RS
P0GipmHCPAI388j5El4Jbh3rcNO/oLcuQO6hv9RNcTSetxVMZUUTiHyWyzzMZGaSZIvNpHRQvRqd
fufgN7aFTGWXSwEq4+oDTvLb6MloC3sbWsKpje6yNLfsgSZG6Htqj2VZKE2hOa5VLifakurjqsBD
R+eWt9hG3nHuDBs9AS5cu+hh9/FgEEzoGkmMkAmQk8VUv2itiOma69wmruFC7rt+/8bpD1W2un7c
5TWKXnlXQlOPa5yEddBphp8Dlb/Ym6Bu+19aYZiZMUienUAFYwpzpMj09kEze+BBBAPRuQEM3AxP
p4DoMnZZ6zdQMaTNjTE0EfvJqn7eSaJQ7ABozbSfRFxqCgWYEm7ZFu+pGOO1XsmXda88hRLTiEl3
HffUZNywOy7m0F2Glr/25bUtS/K1ir2enub5OkqxML2ICxPH0psCunm22qmSuYscC6VVRsgJ/qc7
u6mjvJVdLc/b4sI7r8DZu+zWSyGb1cbU1aF1tatpm4g6clD3itkqJ3TP10Z5a4rZwhEQ6sW3dG2M
LP/2WiYhMAM4bzjtysj6cDXzlSTvrdJP8KP8G1YSsH8E9TZZAAJ59/cllWZ5zXSaJ9SvwjxLqqQ8
DPUi50CjTc668gb2GEOk4hbaFiCl7HEhT3HI7uQvWKJlxQ5QZJaSsYUapeM/Fn47vLIczcwlhUCB
7CKbFHLGneOSmnBUCvubHplke2QSU3Nf4w18+X94YlkwVTwD6suypdaDgRElyoeNaRGxwiyFzBgq
Pc4cv31hFxyug0/34jACK8lydE0LNhXPxmuMKx9HrmuJReUQO0SE+6UyX1FjzDlZMeQDF4iES9o7
B9sVrWN8m+CSvesRJJeaRfwEbPLo5q9vbbkSANWdpk5QQpAdxaoNpXLFQGUFitKD1akcwMxJH/P/
VJJNu95MOC6aq4OzMfjOOCSHd6jkot5mpe0ftwxfXc3ayYdOoIVNVQLCJBdSmjlrDbkjI9WWPXHS
uIv+7HEX/OaLTydxFhqP3NTelfsQM8Ulm54EVtzS21K5QFqkG1T6+HSJuh99gZj8VdynyAKgi3Dv
ki+dcTslWBNuJGE6aV86rM0cz+emObzFSDICA6KrRdqkzSLN58xg7eWvSV6vAv6Pjdg947SrTTh9
47CsA2Gp0G/T2rysZAr0ERmaWlz1WrkAF7gsRpWvYES8jbz/kIOlBXfrsqd5w/MZfQcJ4m6FDSid
fsUVZxBso3Qgd0ykNKfo+DiLc9lBw6TpBl/0zGnvG0Hzw+91BraDGdUEaRlq8LJuR7My3WO70ZKB
+nKo7ios6pLRmhdfusJMeIrOvbHBvsYG4+ls1gd1fPebeVDGqdEbh+j3EyklullBf2reUM9lwpJe
xPbpG+IOhwfMM1mlQb/ERyW0LXYuYjYwWHW/U+607n24lfcOr5OoT+n6ZwzXB8knHrzy6s+Ujm92
n5dIoJRqi1ntPyA4UVNgxNrgq31y8ZCf6mx2r85yoJLxRiCGxg+WUq/TYUtBD1zagEvWccVxLuDo
xQoLRoWcd2nXPUJGeU80JgshrJQSD4B+ZqvOYRdwetrxuthu0ogjEZovwEvDgNrcV6VbV6Gyg4cA
yPYq77xG9RKHHcqFXAy5RozQA15nf1NK71zhSl9/WPBQRPTynETVXW3h/PxlePtyM7bWIEDepyPd
9BAskHgHtiQOo3EygwJucjgRO7EpzkGBEpc8eGe88as6Wshpw6UjEWDXpzf7PT5wYB67RB87e+1u
K8usG6Mzp/9m7Tk2N5YjbhTBa7252l6LVD0EetkcyrhmO+dqZ38fqS0tNSk1Ew/fXYUpWCQk0B+K
zxU477pfQGECDcx4txEntChW2t5xB4gKXaXxUX2Bv/VahqvLzu4zXpk8FtHLL9BnHdgZ1TrZLnuZ
V6p9dSLaqPI+CnLL2jnlE5mvf9KE1B2ae8/CjJdpxsHFM303WWZUDsDggHczZR65zFjV4xFMTD7K
0hConIeMQ3qY+wfFh1rrgkHb69ojPOg5NnUwLAOmm9WMJPHrSJJJaK22/ZK/t9Faw7miJRkjPNwP
xBiPVNfAoAJizUGM2teu7rfLQaWetFhogsnoV32vpQZQN5jUDQBmzfq/jFHk4NG1dLAKOkz5K2NW
6jDepXzWfya5ES0AjA0QDZAAU1+3SqXEcXAbFLOlGb8OT443HrFnKUDLO/RibpiOz/7F9cqVA/8r
rKcRFoxyTmY5QlG1uH+Pv5tZSkqZSFq+u9EllDb7pZwxgGzthazQDqBOJzSN6fq/plhyq3ZsxGhd
xlhc2KoFZ/8ENYghLpD8B8NLgZvSQM0vv+UYHWkQQcQ2x3PggEbSJCUTwGGpDTvKPnGJdIxwF5UB
fCA1FUmcS67pBZz+QUvkCT4YyrLmkk12OYgMnTTJbc2TNJ63bBA/3t2GkGKuqNeC19QTXTk28TI7
WNExGP4wgYSD7YmxKEOWsC8JP/qMlWF3fSUXLp7Inbvb3P6VOuYuiEUe+DyH7MmJ+mEemJRJHtdF
vpoHhGAMlQVB5rP8J2y3T9zAzBuGRhO1/YABYomMbEawTf0NqW2oH9qc4s7KqedOdx8ClzRMKsZR
9/cd4M82eSj1jNBCg23VmtS8/RkVVtDwjC5BcTkVfuz/PgHZUqzfDt0fKCfurc0t3T+2uSgUCThv
YVx61uddXY8Sss7fQ/rDkfB05fUiGHw1HM8kJrAvIGal1ve1bhCKkFa+N9GCUP1hwAU+iLYquESo
x0jarfO3jqsxateaz5isEi3DUOBNzTkpAgNXjo8ce7B7F22FjoRDPBQBvzwq/d6p3DtKB17+UglJ
ioecGG4XsCda5R7E2iDDT0+rQnD8na2HXxVsOwbfC8VgvmuLA4qICsZI+HbPqj/CApEu+8lO3v/q
lMy5mhhlTppSSCjJixEm6M6GrmE8OGy3KmkXNTofXMlqcwQZDDuUcC9o+j/UpoBx9J+K7EJfZAZj
f6Er8CTaXRwytdagviLTJgq3Xl/YdfEpL15s/8ucVma6SJ+iFKyoUGek3bAGhQJHgwt9nq2Lbsp2
hBuS86Q/ttKE9IpvtS9ClwnkEx5q15Esx3EB95hO9tbwPK5V1DA3oDGPFhoNcRxnDHSfENF0KLS2
ahnl45+LSYLCciqWlb5GDcG6/cD53qO8IK9gOLNJysOiWD10cZ0wIo6XDGk+tmxe7LHQ0lBvRh7p
rZHASFHeQh3GnE8ZXIC9flBxBVkTPKAz8/UwSC3XKLIDRrcJ60ZG3tBq6ZRw/FZxPAnrhB4ir1ng
WbYkBMs1Jb/X3ThZmMbnygn9RgmvOaoBnEknvWILLdJTL9BwoB/jnI7wa9klsXp0lOKEhIJ0PuGV
MkM8ZIY6vvX+5jed5ADPrUxAM5HRz3MusLyuWeQMKprw2hsXgWD1Cun+J6/2uux9zi8JOkUFcTg/
I8yMEnlfkEsU36vvCcA+buo85sX30t2ZcJn70KAf7kueG31c+mGIakCzRc61/rdJL5Io80sNko27
0pbctRWk8gdTHjCXeeqFwRU+pcHtlm/JJGgl4SMxxHNCMFvoa5bEZBRcJzo4yF1e0z1oSwWHhSRX
PlSPBesPMg56TU8QVZPwGmvtYnnSVqbk74UNloR9OE2GgpAq2eqCx6diGzNEqYDUMMLiaITFGY4w
bFyZDiTfcB9daohtavFyugNAhOyVrHifnu8GJulGIE9GLXgJktTUEr3jkrJaMk/ibxND2oOdDBOF
+U+if3MYcTsZApejCSkX/gHxeciu3DoL7yhIqi6rX4a4UP+R6ciDHnlPLIdH+WOBKpHmnwbvQ/l2
5MCz3XpE5iAEUHvSUsAMGeGckaRqzi4HupmXObSVkIW3IzCsb99W/JnC8kNEWYsBKJ7S1DtR2eLs
0dS+6UKa1XXBq8h0Fpe/VAlH0ZoWUMHzrIdpO1IFMRegxrt2Kg8cfh/rv6nR+/PpGewk5OWfbex5
9fZtt+PSICq08mkuIdl7M2Xap1kFMzEcHgD9KFD/qd2dxjwCpcMU4370VKCD/QrFsAZFI6QXh7zd
hXjz/CE2N5t6KTMtuxHH9NmiN/OwBE2Zqrj7D+OTTSaR+busmqq5KepwSrgYVufRusOvmQC8oByZ
VaMqpwc2dTbeX7kC1yhJRpyLZHNzJIB5LGsi83ohOTlApLcIpMI49jiej+ChdTxXoxnXOHlJ/M1P
1HVjQy++6PDqchfmr6r91qnckDiH/1AKqM+RGINxwTU5SRzW/E7maYooNicxFmRqSGxC0cKidYAy
LA/pXe+f4Jmf3x7On2NBLdKYpMR1uZx4j4kFAKB+UB7/hcYhipNL0FWKyXOWAOiRTG6YBGABQJ8t
VOBqHlvrrlE/IVLbuolTmz8tkOk2MngYCbSXtYJTA630qBNXsVJOVjdbjDu9jvb6RpomTdkpy1fF
Fg2zsdghTgwQObopFf3SpPaLnX3qEmBy5e6+MlejO6VKCNOiyc8b+Yz5rFWVvQX4ldBvyJsgjcP+
lbgOzVkp3LOI2ew0ppNsm0FasKQvAwfFgkYIErYAnbzgl/xkOfTuN5+U7s4Pc+oBaz/psXAiGOEu
9IZyZWpaov9Sw0SLqJe6BuN4YWbKMgIibjxFktn69PcLmwKUzeesFVEMbKdkIK5Bb+bGvvLsSW8t
My6phWDvQCWwg5i3NXr8f4mMOnXL8p24dIAPj0d1fK5eKfm32MzzKM/AjohkoCS2od2YdpzCzcSb
RRnxynrfCZmSGg7CYGuLOnGRuvqa3NcMv7yfX1vs3fPg/ufsmt7Lk28Acx25f87piPJRfwpPvGdX
RJp0Eb47/PyFZ7VTyhz4/OH8tQ/mShJ/PTkgcgS+TSBFPk+3qRYJkiD8Y+GHA5fMgmB62+QYZh9/
yZh3GnFiFcQ5IDlaCeA2lvd3nD+4u6IZljAQmS8hJU+WEgZuo5OZTUguUvxZYmx9FoCOlxJBFNip
JH1h7AKbU0WDwpoQX89V5bRfrJhXcjUo0yYs39NMG0ClIz2w55U7LRd9bxD3zLVwdOBG6UJbFal9
1tpTN1woBAt1V+Z9xpZwx4tx3BZTR7tDe4tzTNLKt46zHUZhIM7txlx+Pwhuh0BhpSA91EBipFIB
4R0SMCYvcB1QP+bMuw0I5igOydis2t8YylmoFf6+Gdu9bHPOQjiU9bWUvYBaXM4ykd//o5W6nF+6
CfxXtoIBN1XtB1IeI6fXui22rMp9/Ejs6SNl/sJeedIiXthWsIhJhHVBzkLdajwBlZGBrgt1qSKf
ydHOIToYtepzRUVj06DsahCjYmrv4zhOfMym2CjsnzEAamOQFqWFA4zzdYE0TFa6Jv6RjqXTkUxb
b8juC8Gt2IliP/GvwaJEZ350nqSPbX86/NIHgahD/09bDDWadxlGKRV7D+qzWx7YARZla46S+glf
7YMouHnjTt2ttihal6FHp9fo2Rq/C4HfrQr8f3rjarVvLSp7EmAyBMEV5Q9BJLSDklXNLUMwWznN
L9jX9IXxnkc2S20jawiX9rXGi77jfiNRIJgc1kLlZA3NIpeDQ0gJS5wRXpqsUj5BMuPlrWvJFaZ+
rwJy7wnkNu53v75prXmo7uy4djEtunPYJrzRsmA5e6VdxbAOqQqfUAun9Vyw1sG/5zJC9vaw9lze
eOPOfP+WoLjJo5IHxHL4BEbDMYCDXmwySUdbCSp89yP0/iQPYsooIwLyuChAxyg7QCjYylMLOf0C
PkL2I+lXydnxcHJY7h1qWkocv6vxltFdanyCPgCm0vNJ4TSHlc5UtVbVOB4ggfSwkejRHKRbNBK9
Bq98R/3NvlrwoIGO0L662BUCjbGwa9svQpeMNy/Fg4wPwOE9Yp2+hJ/1pq66gcpLdOPSvlF37qmb
MaeohnsGiNRdawcXZqVxCqwOAWup0rdaxUvioZ8lJwaRjEp7VEb0pLAg3LUOJ9h0XrvvsTnn+MCg
CWe8cQRiMYaQcNgWi+bWBZ8HvfK81yOlIxAWPvaAK/YX2DRSXEV10tXsog4bnJIXXMXLfsNNIa6x
W9JKorGLtujXG8Mlhx/pxbIpkz3k5Fo5aLTpFe/XHKuubyhDUv8JfE83boFt0i/arLWrFsh8ID+e
tbPxba8exnrW2Bw1lUaMWHtlhsMyado9JJMeNUmbTqBJ/e1Lcm++BgpsrYnWj1F9g2wDPwD2+cZf
8sZ1MX9mvLkJzzD3pjnVTI3EIW+Br+6ucEKwEk5f1WeSdpyu8kXRVdAWZgiLBqDzp3xI9hziLIvU
3XOIo2bckWEuggGsd8wbj6uPPY1k6OOctBRI0ZpcXbIm6345uONqBoN+irwX4dzxq7X2OheKU+4k
A2Cch5gBAMosNJqHYCLv7V+xzP3qR3sYmJrW2k8JlVJ6Fv1IF0UCSu/QV4N/c2oDC1gJlaUnQRgi
EjNK55OOD3zRLWwHe8Cc5T/7xIQKDGAUPkrRKuhdfvugyAyTBXn5FQ3HUWErZRXoMjRJP9Eabbq0
Ha5nN/Ygc3hp7dBoJZExu4DIzKLqM2e1wn3YQf+2a3feR8lDB6gd/Cf462rTNKNHirt3B1GtnHPV
JeSKVw0PjultpnHJtkkrVunJvwOVEGJJ8XWRRHDiwW8yxWFbCvu4WaQ8mgSRtAsOEfYs1uw+/fuP
Jxo4uxqtg/496sAM1WDNhehyQSdOnVOAjRbYTv5t6Jq7jjMYx0wcPuSZJpZR4zqYXA7eR1GOFBE+
Jl/NPNjGGIlRBCIWfECN5q0gGx49CVcvnR0AYp1Vhx0CS7jx9LoA0LilJgDdQZ/CiAPNfKrIY5V1
rF8AZ3uRm/Vm3ZO8Siojm0657KnP90xJ5a+WAqy6gvpnUzs528nHq7dBdS54fUE41lyFjjkF9phU
QRAe4XlEqDWumz0UI8QQm9EC0COoaSmSrTEabWEW/K+7NpIYcirrJGd+67PowsULOZoAYASCWbcw
T1l2g/tV2C7buVwgFELXiJwF7RI/+Es8r1a7BBdX2EFVWdL6KqXfPjFxKSxYQQNh0OGkO3FUA/P1
yZE3zF5jFpegd/wZbyUJRLgXrHf/fGlA9iXtpfSb+Ttg3R0flJ9Hh4Sd6NUi8hO/GPD1/BT3seaF
1oPPdqF90xqk3Dvisi97wY5xVRtjhVJs8+ctdFgm8/rzVbTCW9+ECDgXTFHEGLQhdPwCZcf77ecS
EH8DprAH/IVmhAbblbG4w7mBHjgN9Ex0k9Ll7I4YqMIYGnQ4MJ2Vj+QQ4qvj+uCO1jw1ewGEgm/U
PtVuGQ8jKxj13aKFzke6NVRzu+Ko1Tj565kcC08j3/b2PV9HKFHH7K3kyxu8hYpnbC/NRTT1Yxm3
Rzv+WRVEQj5CMOzRhhpuUTrums5odd221UyP2nC4KHHn5nK+xd5s+6+wESBxadinOasXZkYCZUTI
xXZU0/F68MQ8k++PaaS7WhEDObhzmnI87/4wOyAgM1zdTi9eM0QveKmP0yR6Mh2Phaze039R8p9U
e5aJJu0uNjazaPHAcOmZH+7MhXwb9swcbuc79EbqeS/B9lqhpxZzuODAy7mBbz6UAH1grndX1c1d
VI/RpsrQWImhwz8w8GCMpwl6KLfpBkobuqMomg/N/BqNfWsrknzLfQsDwoBnTVU1ff9Ir4dYSQ7s
RvZw2lcr8j2Un/nj/pgPjlgvqNvSGg5i4v7S8Qi0RyHQeiZnT2kHrXkmJPE5PFUAZZcVwG59NCwW
KyPWC6ooETj8VmtVpUkSRZsVHIJb1eCFaiDr7Rt/XFsVwxwLDPYc6MwbU9+CWFCKVRlW2y+1ElMV
oS8zQOLL48OznG7tsU85FFCGyCK+0QlOdDJ4m4ST5oy5RMWIah7aiCcjIb7gMbPzjwYp3kAFOEDg
jvV+Nr7YKNDVE7EYcLHY7tpWgeWMpNfI369ZG1vh/oFB+x04pd7Ib8sB8B4MDd0CMuElIp55Ec/w
r0mF8X+VSgjSaAGX6MDVNEU9AQ0tEMxqNkwHPSCnPJCckk2yDp7pmxLXMWb0zKvwSZhOM3W9QBbq
Mi95vK/qqLeeZFKvJ5dBzPmkbAaVEn/HvMkWmfgyDpm1rCexsEnHGcgzl+1PUBI7l2+q7aOdTjYG
OS+Vn2MaOK1t8VdNChow8G1mtM5tmLfpu8I4TWstYzyCetx4vbtiOYAbM6s7iNDtERNH8DpiFmZ2
SkHiS7k4cocVWLFB9UDTyxk72a06CWap4qlHrR2nSdO++6bgy4hUmAo8xqXiJTccgX/BwsZMHHMQ
kShEFq159YYPVEA7Ud35CDcKdUkCniz4uA6p6zSO0+yw5dl4Kc4IZqxsm3hU5x18J7a9xhkvvfC0
N4hmHgzBufKCt23vxrIb+rwYZ9rtf3pm4lAiGCP+F9YOrcivx2xcpktt4b4rkhzvkT3K+dX2F2zU
PGgPU9/hJBqarY4CFmtGz2kyVSgGxjEQVhmxU5kFJyfmsrgemSttfv8qH6M2R7U/a4RCu7RQnUVB
MhZ2Vo50l0Ar9YSr7F4gs2bvFeM1mfPYYy+caegnJ/LxqhTZZjUO/LbmbOGR3RMErqMwJJFTN827
VvhFL/uITYmvNQZdWKRotutvPEtfPICw5ZoQu5BxObAIJrLjhEhkseqDSgxzRpwdVPaCuWo4MVyH
O7/7+oe2u8mieIEApZ7uk7Wd5p6KjWfVXIpv3U7SsqEdx6OGvOha/xR0HQ5L16s4LU4LQiTueX+F
h+8Mi2fjfLUpA/Srf3FrAKjOf8Vv3CmLK1bMtmtFRvjAZT6ZoXmpjzMDVCZoM5l3hzCkiCsv1KNJ
5kRy9zkMsAV4R3VG+5SNeSadTJrAIYa02Ayq2ZMvh9Q85U0sEBEEzZ5impMxiPuCcYOZ184vzNCW
zHBHKGn5bHzJV/oriaeIWCptLEOyJXeLa6RsookUG155dvX0idCvBJhvu/x076CtoJD6SBNSSBwY
pswGUpRz5DEah9gXdG79q+bXVJIax4KjuQUyQYRpW+m6IvlNiSdcRMUiLHrYqSYv+YpQHfNrS/de
jt/jpToPbUzI7xonn1F1X0Q+Te36BlGATuGuP4azXmOQNpwvH8/+6TjGsNCLTyKIX7f9KAjqHck6
npolkTYTcZjxPGATbRYm7nVlHjqeMOGBIV1AX38GnhRERjNtpH114N2+8LcPnrvkOcKsa2w6CzhT
S20vHZ6Nb3PCAN1oMnjdjqSi98ef2Q3SeVNV1IANy9aks3OBOUBPM8EHWKz2A0D+xpBVaTvmsfHf
QmOV3xM3kzEwcArH6YiJxV9XzmLfArmyixsrRhOH38y/ZbFD9lHWegLHK7bS0LvReFvtQ8TT2ECv
XwmqhP5lyNxHc3SDBx4Sh9vlnMl28ps7AEO5lYRkMsoYI1bLbZ0ohHRWfSSLJCEcH1pr7gXm6u17
HGu8FnX8Zb4tckpBNHVebQnCh5G+3GWJ23kwSDX66yShvVWHGHnWu1vqwk6udc9bKwovXEiL6gMX
poOSyDaAhqbOGgsvAqYO8PVLCdiXC1d2xvoZuBlIDpTcXE//c8rKFihqUTR2qB5BWuv3RIEHV3vk
mcOcHieulga3O/qI9p2jqSiXN44Gytyu9A35rFOQEpOTZjU+jcGxa0Kn/qqao1JM3naC3UDQG70l
DkS1PMmAPWL4HzZplSzJLmMaQxFtW6qQ7nU0skoLHCVlG9KoYyxaFaur+YcePhmModldGrNz18vo
JOxBwPCI0NCu83/QJ8zRL7uOv1gdlh/f7G59oGQMmgzNUjJ6qKZ3lGHmgj7tTbpHYtFr2XfQxRAB
9WCaRKZCLrlwQKKo0AsiIQ+ehmeKLt7Rt/jkU09btJg1ERMrE8MT+qSyjXoikh4gajyIi2LHmQwh
cEAcO5keE/aWDv4PyqXEA9bCrDNCfm+FenBko04f6A95cli+bLbwBDu08TbKZImkRtLPrtleX2cB
GYutG6DjDB8SMYUlnQVYmVk169mCarOUGb0b0uBbwDkmMqZ9hT+7CIeSaGMLjYCh+9+xFOrWlN2Q
zcDdqH16wdA0g6fsz2xWHLT5Jk2Qr/ZFvIcAOnke1AKj5IUsPGs+S4yDTj+B2+6CEMiHKVlTh1dE
/Kbe5+5ZaIm6tACbynIIXavwVESNF70RdIF9KXQR8ip8JvIe9BNrpHogk+PtmTlyYZimg3MlU1Ye
fTcTAK79kPQCGruBAMZCG00YSRWk6eOT8/y5Flz2207CrsnoFarVsa7w0Nca1K0327S0pjBxMI1b
0qIwHkur3g5AMH3OZHxsSkT706n5wCU6e4+EqSwS1rVjLepiJkcghEEYu+0ZzKsWPnO1Swl0kl48
ZWlXxepHID2FYL7mFTcca2YNH0hHhwpMPeg5JpLT2zVScm0zZlRiSa/UJ8/DKAChrVQErAkojD9w
Unyxr1UWkh3BON2PErQW5bu4nRp/ZaHTp9Y+4kuqmiVb3TAnWHF7U/G+Vgm7OW0IyffUlKzIc1+1
lW/QEqL8v5FScu2ZBkP4fiA6GNL52SAkKZ3dV+f/lKjvgUdz+Z0mcIuhClI7k9pIr4cUg52v3at9
PApBrOhIFLEAgqDGz0b4ZXoxO0qF1DzHSbjwnvaau0Jz09huixP2hBSwk7CAH/5R3ciABtfM5LOu
XF7t/AHvuyRVrHvuBw2jZUwlnn9f5DBL7Cut8ATFpYBxNWP3sWuqJdpfSLbQ99Cxx2adb5lPb1Ug
ftgjX64thbog+a+htQlvAwWi3m1wggArVJ4iGVSsynDNaqpyjCdP9uhxl1wCwomhpAIvM40K8CCA
ITJ8GYGH9gcgp4b5J68F+FCTwGkK8fwVxsGy3uJkO0tkJygpZ5WBhj+BMElVnub4LAY/clqvR+5+
BnRSbeCAWEqikKAGMb2qiMoonmputB7EyV1Ea7Qys+ITgTOQNgDt4s4TcNvdeyG8URNoF+cs4pB7
Jg2gUQrKaFYteVMBDMCvfR5G4IZRlkk3DApH8U4dw/sLLQeHzvG/vME9k1YbQcvIEFpEKcf3SugO
CVFpn2vgKb73JLSpul33g+nhRzBLQXP1RVpiw4bdPLdqjWcBAh/H9C+ZAWwIHpyTohOdVJT0OHQU
C9sabP0kOn7ww9Rj1TUNM7U8mjpIunA+UATatVeEH5WIPrW2di8CQjj7E6F/eWUk3Types0nEBZW
JV39LppEw1VBxbbCoOHAHLBktJm8BWMurX1TXaFFHb4hra7DITucYtBs7FT4a9ZOgugnSRjLyR8C
WpDnbBbtSdNXqCWdxdge4/WP0JxNv5v599mCX2BzGqxGPjGbzd7TrkL1QDgO1J7LwOk7rI8zeaQy
867djdJiI1g/1OFzoQ7mIjJDp+k+OScFcNOsohL8LfjGj9QlRjLsiUd4aljMyX560bJXbuXCTTM3
JLPW1BlH/vo9xrMGnxgZcIqDA3cCBeMVSzYFUvsFp6XEGAmpGD2vZO9Nu3y/BSmkyYHRITrWfd9k
0cwf5gYVh9qSw1x2xAQNp/VWHgzkr3mx3NRApD2tnMmxH0LefNlZCwE7GoF2sEXvuvXatHuho6xb
Yv6dG8jwJXfyELh0MRD5XqwB7rjoZQEqm0pJRfqp4+EI67qTOWdPwW72Ges/b2R6mHcMT9nVG600
IYCB57TZv/OjPvq/ASwLE9/Tc3E/+ds8MwDW/lHa497hBTiLkJgyNagh/g5L5Xw0/2cpGMNTCfNT
dzenQqv2AsbupRYRyEcAShFMHeyUv4lGw8vMB4zZk7dXWwnLRGModv6JK2o3ClXutOfQY5n2mlzc
RxL0Im/3FPEQ+a1yUClvECuHcwjgT8nSHFP5Dl0RyPixR6OkpOEKcY8Lc4GlzKygXtXPWvOU7zCi
2iflIqqAusBOqKAvrA+uJhg3KK9Jbwwa1DKj6aehdHgWzILmQQb+G+Rb0zP0S2RavVpDLXIIEJfT
JOL1ka2dJD+7iPZHWYEn84sbWBzfVMbirsiZ4PnhVmVGuNk5ES77ljbxe3YJEpI2j7FimI1I97rR
9Bhq2RkNUboI7qo1JJwzosLQ7rJ7Xja6LTeXBivOW0eXuWO3NbHnxetl1F4+AH0Q6AZPpDoYLq4e
42wE6M9XX1YAQkQjdZZkZ/KL3Yc81IPl8Wpz9V9BJ8UhySmtGFIiaTdQ2uMikG/DAV1d09S4YgvT
5F/7K7YJL+rp3CMAgTUjq1uW2JB6oewBjDMbLkwdOTJY1xJwLViYKzdtnCbdsDUpoFijLzMGTZw0
8Jmpn2xpbGugx9jeIW9mqS7DCpSg0vC0AuYQEtyeVrdEsiPPyUS2of7Po4UCkeuSt5CpXQTiyuzU
b4ncyfUKyrkZvzGazINO9/ZVRGl0nDJpbyRmICozzNB3wYZhycxeZ3RUWRt6QZBmUHOzSGvJVOYu
HuKOb+lzStSHAP8MYNms/grKLjPNbDjRCysX+/ZJ91kjxn8EmqXfW4K/v2SLnw2lqruat7gUI1dR
HTxbKQw6qevhdGIzWTwPl/ZzJ4v6xzi1+2bG/RBSy7jT36oirmKlOPg7LgLpCZxwKTSkgzlAfgNB
ANmRh4rlgyo0sh116WespnJhoLSEQsbM5Ku7R/pvzIgS6e9rFYXF0bPFLuYF5SrJ6sog12zzZ94g
8SOjWRv1+KUEL3HzUvLZ0B15cBrmkHtEdOYSpdMhkaeeGlqLPX8kBDi/z2N9U5q9jMS0nHUYT/K5
dGUD8mlQc0MKqZr7+nllkOi0Vq7MHGhTlpys1usTklBmvCW2Wzw3+prrS1ziAX1pBtCc14INATWF
/+myOo5nXF9tx8q7MfLreZJNzT9qOsowYv2rZmQBTXvhUjIV4ujjdwwFSEqcmNXZcpofaERPmF1p
+OTJ9M3Vjz9rx2IGgBrgwlTDeNjpTT4E1cycfZWEFrdB/w8OcdKj6+wUBSvnjlNahi1SEcvJ0e8t
yGibmicbgDe7JAKd5PHm+0xltyokx7u+k6r6dcXECPafk4V3OmNkWSrhjqAo3zNmsVCTs/gAXQsW
fO07q9XJG2R4vhKY2QK4xylG+pw1ulk4J2n4EYJBK0dpLUlEd+zu2Vybuxufei2iIDqc7TKPYyyD
d6bbagJELSTn2Be1yGvq3xmKvgIa11FmTxbi+PYKeW8gIXmFl72hls+Ik/w2wHv/0pJdFL28HIGE
ZGx3ogwCNtmyxTgcXhqDPoyRgzxr0CQsibPw9e5L537+z0caH/VUSZGEiUfpg7O0Fkm1dOGgp7nl
UidheZJpk4Iah45/VATNM9tOfxRCbVurLw43EYOc0LGBjNB8rtFbS+0I5SPU06SXhnXqahh45Xso
kqODZ1RM1HP4YDQqT7HyFAmyblkc5KNooJQOOFM3BqmGVITfHVA7vvqn5rz/WGIlK71siz7qiV5i
qdFa6E2oSTQB2Yhhm51ZQmxzk17P0TmYDJfdFx0YSZukFUqOU+n05UwG6NAo5m06HJubIXEpR28A
GbOeKbAdDqVuMYDTsWqAsL19vXEqnI/wo0Re1nPHVio2DFa30eVSbizq+SRt2VrSd+9/2hi2/zl0
ou0JEtK/NOP74p5Q6BcFjuDW3xdtigB3UU0oLNBYlKmlsGa6FI5nVZOouigZzHcDBL1zhMSjrlN6
x7W3YbGu6GMwo3Xf1DkoRHhEyvemUA+8CBzdQIUTkm59SKT4ao9ulwIPXegwHC+V2IqF6lbbxgNZ
oUO0RiDEDkA0Qb2BudqB2SlfM58TVl8RtTfLMDUJJn4K+DaryyIa8P0G8psnFm2zDCYtfx1b4MSQ
6SzSYyR3ebjcG05kX/CJoMncnfjWCAYZp2ZUhHZ4IjDp9JMwID1Pks5XemrUdg/emG2OvzG8y+PP
+iu8GBc6t1WIGL+D9vJr5tvtPx3xPkQXewXqknJutjSbTTdusvPzVG7xaqhqc1u6pWikV9K1fuiQ
wy/rgYpGenCSYRetrv7f+drGnnRox0UxKNVn30MA9p11GC0q+kBmFnHApLMzlElKM5Low6Qv0Fyq
0f4B4+TPgpp26+bATn0iZVfpqk+Ko7ZnAhZr3bTEQUnxbFfFaKx9F1kxosLvRrcQO5Tpln8ke2eA
sgYqXRyUSTzG0EFoo+K6PHBg69eWXCNAv68ezxpuog9miCfivMSenO+aeMEzJViZQtvteIi3qAK5
u6+XfLnmjpmXYT7ru6siNkSPGayC5WyE9zcVbe32FirdF7p7sQMNWNyWJYSTfdLXWk6TvKrI/dYp
6rZ0hLZ7O6O44nXM5H8bsEF74XFtgjvjbWiyhn+5b0HxEekzzfIBMYdQDPHugYs05kRHcVdVm82e
fqA4x/8eDrIB7O+qajgQzkdVSxghQOoKwv6T0gUlF4tR1eZ4tqrtkhV0ZHt9dWrtFWICZ02vyJ/0
x/zpZ0VYvPZbT5YtQ8d36T/izFZ+95ls4TioWyYje4pn9lFtl10K2XWON399vN+DcrbvwrkCmGK5
uGx+0chnOF7IxeOZkWWJKYyZqTlAdKgAIQikFGr78GzTGGygkw1egVJC8wEuf+ns8cRpcWN1cdHp
TEaMbraN6t+qgCl20DM3BZVF6FDMyL8tJVB8X6/eYuAQ6qWKmuf1437OG4bt7pkhNKm1bO5BIi9l
9pYXKHbEfoU8arX7Khd3FzhVmOrPNm6vYko1KT2teliXnBr4YAjxihXRxQzsVuy92HUrXpJyM+VW
HBSDxBx9Yn8s2dQDA5hy/ZR+gf3i1tfqCB59tx6fU1S0HtjIh9G6AIyzWkZSIiLwF+vIEVtRjmB/
CiIUyo9aP2J3gPLooktHzMsOWB9lYFbKwrClwkAjiNkpZq/QYMHqRQIv5RjksMPIosC3IJc5d/Cf
FnIJHFdnYGzy91UJiMBlR/OILnR8YYynnV+rf4cgmvhA/JVj55wwMn8fj+UHkfuAoNm4YEE6evCZ
p5/pWMBOrKbptoDLXXjPnK6EEH3Q08GNUcGYEBgMLgJPTBUUDr6Cf+6Qo0pMZn82770hbpPHGXXp
VxqdNgUUboPVrw+OyhkZUeY2qIUmPIUIxJial0SL6bqnvtxhp6KvhrGzLUN72E9KfvkXMbva5RmI
qRD22fnA9nPlBg9YoEX1H3ajKkg4OCf/G0g0U+O8wllSYcDphEBmr07Gxr7PI2/0LTqUirW82QSO
Y+lC//wmWnH199DuI5BcOXkwrEoGr/7eWWzFJHlu59qN8XpNejCKCkO+Enzzvr+s0SevrEXYJUaT
vU9ODLNnSMwlOFCcQdC6uFSr2zt1tL7B51ouuaQEaJq7X+oMSLjoBUj/3SvXEF1VS0W9NVLO3Wsv
3WeagwAKYwzgaxwR9/nwC4MMAMFLx9KxvKQHv1BE6LtVWyVBe4MM8aqTuZ8BOOKnlayKvS5wHCdq
MUt5HjSM4CSOcPXVYm0iLujfg0c5nmK5sK5t8f4ceHQIyJS9PBncmgJRowLO3EmF30p7rMZqbyve
1JrmIuyfagiLnq80bYiGgv8tKVfkNdhelnkM/SepWYEr2DLgK9NWEhDaZdYr4UrSxDLeFKSrJeQ4
o3FnG1Xv4P0ovWeEZMa5Uiay2VCUS0ZjDC2NTk0hTAeBPP+2/+CoH1OlIfDY7i447/gC7eYOxGXC
m3Wpe1gAZ3xaCLiQDAuKYIr+DcyPr321RBGX0Vp7O5J+zW0C6gUcILiE5jBrBnWmu3BoryeRhrja
BqVF240tK8JpgYuvBaka0fharb46E/c8Fd7eqixNSlLWshiKQBTAgTSjayDHNy6iWVFoldq49Q/0
e2m5I2y8PapIhuPXwfqpcgZl3VwpHB3LxbKSUjZo4kd2XTY4PMsVgTUdSmDkxVkZIa1HhRYwZHpq
JdXyyazgSFBLZ7bSA0DL3pYTx+KYx2ijysTxST0SjLPkAU96+zhB4osgAaKVvdm98rqzSiJpu2qn
LMa7JjVmYzLS2X4ahj2lOVTiIpPgcYIoryGMVYKqOKNJ7Z3SL4IWvl+NDpie0Wq1bXExud3rU1W4
s51bBdoBiSacbLex2b/qgOZ+UTApoUeh2lXyTZxwinH/bCxOGljMzsZtaQ1ZNeKgdRV57nYbuqyU
2LhppYYWVV3pBSTi9dL8PXa34arNUO1yuekmPOke4KRHzqkgtH5mg+iP8iTzZm9okHjwHrUU5KBJ
1tOkqJxfCmDSpo8dBN4dTzFCA5qDo+QwsSCxDbicTCiA2hY7erUdYH6QvpBxrNTInNRe+gRQoBuy
6SXkR8dR/yg1kYPNfGNd+bJptwAgeRVSJrDpGnxte8fFv2npIc6cCM/yrU7GRUi4J211cSJLqBdx
CMfVIJ6BhVe5qNwtYVRFe17gCfoY1Pt4FiBxQDaTt32mJQ1zfWDX38FJpRFsyfdneGLWzx29ojyy
GQFm9Yn9Fy2Sr2mRmNLpHUhopET4Z41Fn018/m8xfSAFjoo4uOTiDUl/si7PHqO4DLW22NUbsTgy
KN6oBm9ZyffxwYR9BTvWFyOn+3I9UceAz9lXBbSX5KC9uhl90BzSuermnNpZrqggF5sdB5r1mWOj
/fNSWYW4T3gY0LmqPOBT3olqbTbWTtEZPBSrNHsipF6vWC2Oh9rQKqqLA6ELWirrw4yN9gTzf1dJ
u/+134TXf9ezsSAe+O4XFBUkS8yy3ITd54mtk1FfXLTAXc2ETq/pbcjWUHv8K9o2Ca0HdJVsxteo
Euc/C0IsP2KkZR1ZKlKb6RpT2+nv0OtrbaeHh1XwKOrINE9Szh25tixWbCWBQ8KEC2LJXKTf/3xe
joN5keUHZmPHSSF7yeKSNkMZmdsWomJcmGYUqBYzt83m6QOP5J/rOJ5Uxy79yplZ5DQ4a2Xd9jLU
TRK8s92ogSx+5feJfxf0rjH/uYhpCXbtUqVrRb9mf9uKU2HZtCyWq1sz3Lk7dxNUrrEsmXqPzJSf
lVRcKivenRCRsuVd7KLR52GJDJO9QoorjEl6ptJv0HpvrvzEbrAJEGq9S7PQMARXpWA63MDuQ512
bVIPMphe5O/s6/C2gu6N2eR5UZ6FkoPChuljB+MLrCMkEDx5SNdqYYOn6Khy8K15eYjFCBJYgsYT
FZz6TEVI1W4Gy2E/mmScaZusbOkLFl8Ob77PYKRlS85ATJrj3FGWLx7cl9KJt16RGPW4rhhRPAit
W4pXCjVSyx+AVT/l1SAv4XU/dK+Olg1/o/1PluCEZlIPAGmTwrcFJ7Ig8Ed1sIU5yI1Yoe4CptSH
umh5GRSVzhZlst4x8jLk5ZgbAfP6907vYvdTqJIf4+Sj+YtVmqlyioWWNsY0wZBigsRhk/WpudUC
vvM3DOVaKnWtGZAZSB7L07T2ORci87garg9tp+uM9ZFlYszfqSjLpPdMdJOcBVaqsirGAdn5cQdh
Np5DGk1kvfVGhdmyJHHVP+AkREjDToF0c0HYj7SLoI1MIplUHuXxjco87mX5mKezj5vMeNOh4SbN
4ZfQZbctMhJuIoPmJ5MsCX+L3HeUwoVlwX9L7D+8CNRPhLs3FtibffPDCCZuQR+hpKzlwHBZ/mCv
UhRzhyFeUk1ABxFB/yNz+8ueYYW0BuXkGRBNJ0QxTZhuzwEBzPxWGClwP8Whu0T8GG6i2bxhbitJ
oly5I6o4bbDyb4aTQ79I+tiGhlBTMRkpf4fcHUWXDHEP2S71EdQbGJToQtuPXyfzWzAtIBtpEP+H
LWaKG5Yp3VB029K3dmXViA7ZrkzWyjxvol2Ojc+Uz1GMD6M+jtj4m+KzwUiQdG+nveSWT782pnYm
1R+6YmNVaRBnopso0OHGdjern7Nzf2onC4Ivmmrv5W1opf5vAPDEZfegz5NuB3G3NAsWg3aFLzH3
AGbGt+ZJ9nTGDaG+tKIqBS1ixMN2144h6gkHxTeHe9q1gd8oNB7noUlqO49uNauMzh1GmbKy0wB9
wq3H9QwD9Ntaxj19CSwN3oMwZNiasD6+hBy9WpSbV5TCEvQTPL06AycRbqfDcyT/shtUbfAR1WAp
aFLltlGbSkFnYiRezuS8uaPH6LOs7N5/S5o5BUVnW9RDVyqlaJ7FJfCH/eDfNGtsdrHCsK9+uvah
CRj0z2VK/2+PgtfBqZ596rJJsCnQj43m7QGWT7u3/Uh0ijJUPhkUx9Mk4YEPsH5h9ztJV2u2wZzT
bX9iNX84yZk1prYKC7jWWAMXEXYPxk0GRjy002hSUEJ2RDv4E8KWbna8j70VZlU65JjM3pnhTFCt
aKRtK49Pf3N/97P8x3AnktJ9y8r+23e8S6ezcdOnnyq8L+5eABdJmlCkoxLXBGZYjM7Zzkwpze61
mLJ8WJ+OX6bNjt1FMvgg+LQw6J+M47trWl9N1RyouH7sZywKk9dF8ykKJP/kvYnWz3GwKgmfFjHa
dUvV1SFKYsbbd02KkS6IisG12d28WPNz87beR1TtwFmGvJoPb58r3msZSFSANHIxLTn+ebH+y7td
aIFXkLIlOlihiBsP0q78yfKx6XRpmDtsURqyJdY5dDLO1Nq+N7n2Og5wlXfy12CJ/pqJrXYPxDM9
mrSU/5mcqGRWcU1H6ESvmEUEXFcehkpv0Z0mf2Fx9XmoU1aiaenD0hWrmlqPkR8JRGgLvdljZapU
7/GvJbjiBxekb+lhOgFoghxSEta+IJUqeoByn4G+SNzNrO1E83Bxu0bo566o/8+5H5aF6yRBe5xC
av3ykdE1buj10XmryqEAiO92QmwrpClBhZk50Wh/yN4W/45zsYpndIv7FNh/IA0BjYPaRDlWoAkz
GXs+jxxlEPeWT1/+ExJ82nHtTXZE+Ai3LMLnVr6Pq6Us7viz+CGPcnp7IyB5EmdCs+hCfadOcvaH
9wZiA/DpLFwC6mE4y5pOtpyqC75hrUzzSM+CxS9sgibYCgomkvjY6YUHKiawvZ9ittrRuDUgkHUy
uRBOCeg2CIsRcLRsRwJz+iMWrhFyLDqxgasjhiWcegYTAJBJyZtasbtsU3J4azq/PNP146pvkB0X
34iw51VowmRANaiJFEnzb6S8xd/3tOdZhg5Oe3zOgtxCHFg72Uv7jPz37BqxMiIsDSc36UlFPmMq
iQqMTkhn1B9Dv2P6ZLKQdksqcZqE3KcsgrFibpDCzPn0SlKxEH+CimkfL+pFYINgJrhpUMa7eu2A
pfzJWD17FuFk0GJ/I4HILQ71hAJ9B2/fzc9+R1t1L/FEIvPx6hwWpyYunDz+jGi4NlzwxbjbC/FQ
3JEmT87bG4zwOeuUA33cDbCeQ3GjYSHH51WgAH9osy893bRAjmab/LHSZzwHGARY4OruNK0WMelf
bS/joZhTn9lubhUJbS+83RwiAlDAh3mru2glRg0hcPW6VWk2bIvIUdi1cQQ4T89AWfGZxc74hzrG
s4gPFbdEKXazGQBRmpSmrTUvZcKNpxbwyq6RW9NW//Jq9ULZGFV8O89bRkh4K74RFnPhulm52FkX
pUwYve1nIW2ep4Xj2bzfvZclw9Rwl0g+rDQkktHwFyCp6h4XTiGIoWDNMvZE9qKFab6qrxAWpuiR
kF454dBHvG9L4CwKl91We2nKWO7FATqLth4QqLjALt5F4NUHW4tXqpkaf8/9gZ9WUHqPS6EbD6xz
YgwU0KCCNAvbcD30IrAhMV9AgLwhZ+8OKII+YDmX4tZxGRxwjV2yo8eNFqxaVdxFkMC6BRtR6hnd
vHXP64c7+0aOVOT0mJDuK5VHZ5BC3mdXiM03b2Fwl9IjL/gYKQKu0J4w0hoWYOUYHth3uqC21hS1
DO2E5B9Ru8CVQe1ZV9E+Hd0vAlLeKqrpctJGT6U2f8vjZFYLNG8owM0J+wjnwOy9U3anseS50VwN
IWjBDTJwBgitTLcOMpg056K0Kei/BGmhV5qOGFf4knNFqxcFAihsd2P+Icb2cbH2bmefocmNKO2V
3BTo1QiQK8IOz4LIArjkmnehZlOb9QpD+dRz/9YRH6E4ufcE2VHHhD5CbeknfrvXWhlSu/VqJtdg
cCUUJpNMxv7izhuPQsbR/QlT8xY3iQHN+dpqX5JPRbfjfRui7i3az/0/m0HAAVHoXVw8scR5gy6p
fAYCV08Yso7IfCq++A56YNvfBYqFGBFIgYG/dVEatzlOS/WykOXsqcgflxNIAkvUVxcavn2cdEcQ
ArF+EMPmcIfmrS5TOlNOdhOvi03hD5a59DBEcpXWxwK8MGWtQoAPRUvZKrJn1hHRvw16+wmasDIB
55iX7nWWZ1QDlLDu/V03Czegpp6iX4kpuc2ghP40O7hCrVOi9KivZFU2NHvD6pqh1gN57XtOhU6s
2HF9Qb71GXAodj8H64BucVRnlImYwxE5Sesl4AUsRucLEljyjGF4h+MCEWpmO9dGkA+w/0q+W0uR
840hgi6swLNVi4F9xR+B5NTbcdQ5TYNpVSDNRVZv/F4FlPe8EBFsy8oTJTTpZofPNgCUQmt4gX71
Oi70JoFmRGJNnAxuAg/JnCNlMYlq5d6NGrSiSuIdiPL5ef64ad0hprN6XgLGyxA6dXyd4my6LG08
/7ecWJRQuRZcmRu6B1uJp1a0I9cPsngMb3zCXLg/X09IG4YCu8cj/Hlfv6EUP6GpAwX9WV8xQw+v
RhO4AKS3aPJJ/Ta2rxk7flZ4s4XIlpiuNcH/3WxYaWzt051GCt17jZtZ/Ehp6qKylQTKJoZ8hYrj
UyxjV4U1MU/b+OEE00g4Jyv9VgbLljTZh7p+CfN9AdzA+sIvWKeCSxqJYQ/lehvij9LJedxd3rlE
OXbJQm6oKXlc0Kmboe9N+3RYoMoSXs9a3wMrCi2Vb3DegJgvNETLuETiVEgnjMggk8b0CZykIpoD
r4y+sIdtknsBtvuzXISkoXdXYNpMubPff03oHXPSm3iEUQdHJ0AggbDDN7skK4iHNqiurEaHI2E7
lbSM37oJw1fRuNybmvZ5R0yR2/JTb5unUBi9xtDahuCI3gCwsstJSSs1LHxSNvdWj4ytMTZGhsDL
fQ46m5+guYc6BgbBgItH8fKj03KA+IBH/FwS5nExGseyg8e7YxZLfI+eo44F+knJ7rLXn3oTbqpC
4ItRhiXb5f4JSHtPcupJRIh+z9gZBORqi0L8yHamLwAOwCMuJoISVs2SnjkdnUZqG+4JjIv7vsR4
K9A+n+kIiYuYaHqDSp+exhOQS1Py6wfxJKkB1YsuFgVSrMVTwkuZC7R/ZF5uGB2MDgxzQ4WcWEX5
hvh5BXxilMSJbxOs425/e87TL5s/JMmTEPDWrLPAOQzwt10Sjv9MjCXHl+TuDWlsQPVDh12G7OYD
x1uXgMZ5+VyUgVW7SRun5qJk0wV6PG/iZCPv4Tq2jb7+/RTl8BmgOnF6ne6nVNl36GIMbSmOOxlH
/9Hj8CQ2gQtNYaCSrbAlahuwCSN+pvKpBwV1RdnVDGTFAWvddQlo5tAb0+VCeGXM+DFacOTwnsb8
kINoKRs5BBOTXuel8v8SgpDK1glMkIcLnpB85oFTiLvVjON1m1K4m6+LUNroWr0QgxjUnOs0gvGF
LO32v5kfYpPOcoeA/lOoivY2rmjBS1x7U36iH0DJVYCDowYt2Z7br6VqBgAdgXu4M5/Sh7iUglgY
fDuQd25OCj+wh0nUWp0nrfzYgrS0LI8lc+POHgRQHCcQY9XVqZYS4t1mYeOkHBj0GTooDmZ8INsf
uRJKSCJrU84iybHzWbXfUS+NnnTvtqLk3wRNPP3srH6XbwBcjtSbSh8x+kePRW5pWzRID+Rza5hF
3V7220Exv5MImihDxT7XU3NW5DomBIy/5t9lKV04cKA8lCD2p1LAw0f5hPVCCBFuqRhcZm2d6Pci
lbPhCnMEavnicSj5VSx5QYEqgUqi1CENa0ELtJ3wIv/jbgrdFPmnC8yl54NJKoLMPdVuim8vtTzN
pESow6pIqTFda2iMOz9rno0l7MrQBUz5FK3pHbrn85eG5so+IJvVTOsfT8IPXBepFqFuy4uZFXCm
f9Vs/V4y9BjoixZZ7puxqEoo7eBNoxqhz6rvtUJvSBV92wWud73a4Rc0jJyALVngFZ/Q7qbusILm
O/+cZMsJXNsqUruaKooz0QwGpFvn4rZqrWjtn/phtFgg8dHfK8g8Z7SbROBBY8k9bs4X4mJDem7Z
oVjJYDRFrZI//Ir1FaIljxBqU9Usk4cXfxE6YAq1iBgkHagmW6fFoC/CElRLu19lCTBWqMzp0A5G
FDNO1orIsTlG/C3P9brnasSyMHuoJ7Dbq4VVDimTWhRglbAZHNGkGOnF4p+iF/WBq0xtheBHUBqI
qNdivc35rbr1uLMil9kLaJtq0aAr2a9oGifjYtJeDrzJ74qEb/qusUBaNMS8aR98S3SeROizX4R5
8vEKs2N2VxJhnOkA+9MIzZNgVzFeCQOfG2jwZm7AYTmE8ysf0iFKdD85d0T28lR2TrpcmE/RTqHu
SF4+unXqjBfzG2hxi3JZ8PJVsqukz6wy4+bF5iD/1j3xfWA99RA6zivyH+n14I6gzsLvhTyVB4uE
SPvb6kKx+elVhonBMxUda218ox7QjgRXFOltFO0qOhLbfqxywGMGlWarz+VBPvyaWjFk+3I4zJ6n
r6i1Euf9RMM04nBV6ykjXKfkuGhJ3nPNLO22RBG6DSG5I+/9/KYEJQ9DtrBzASk+eOjzhbqjhK5u
aPyUhtpe0cz5Rq2kmzxrqTcRCh+tMIX+fNOtbd8aP1zmWB0PRRhaAoTF8Ot7DOj8yjXYlHFmVY/0
vrCENqzxLtgqAu3dvMfMHpH8kkk7XeoE0RiuSvF7/KGqMGvPu7jkbB8PJQmb5pJups9WuUHG5Ky1
U3mMpwcyjaI7o+kIZ7/YsoADR4ghpBhwC8YYyPQ2XXFtgEjtpMNMWKhuMGfkgO7x0saeZp/XHZFJ
lakrwiMpgWs5nsvkLKXqArYPKJ55eiPtF7/ZUQsNZbBT/itg50Wou5lnHrPm+wWwkhyk8XJkYLQB
PbXzRQhy0pdsR7eDFzdLVQSpzKAIN0xkTVajN6oUuBqMf5qSUepFleq+dxhdu39aGiWYXXx1PsHJ
KaMaDnWnRzBMha3R8UEaK0U+jgzytVI8ylWkOl6xGy6EItynrREDxioTJLjzUPdtg3WiwbvZhT/D
zPAxoGI+8uptPjFQTkqN6MNkEqUe+gpXTTLbgXPfzAGztzr3Shi33YFwtC6+S+s8SIOgKQR/r+Ws
ZI1RZieZka3xdP4FRicrKj/v1EUAtJZ2EqlKcHZxOxwTsSj+FCMhwmqAVYTtO0bHoeIC+ltt3RBt
Z+sWGHVP92fmhA0xEIwmyKHIXUwpxPvDcAqSyTKDewX9edp6fC1SwVC56W1M3FPLP6WisEBvhhVj
UMAkZyPHaOu9mw89fwY+XZkDK4SQlp36jxXZEnJY0TxdG9zG1k3g0Q/PjoE915pxDA7r9lSALnJ5
wQOkaHRQkrtGgbi1wGx25s3GtgSocnXiZVQMn+Ox8rDx1IjGIBg5ydv7TbPp5qnUEozusxBOkEhN
rPFEJNFQ70GL8MSiM4OEAxRpYZfgOyu2/yYsJWVJuYV/OvnS7owlL8eN+OJRGDUmfcNTSS4irAZp
fwVwgmNn1CpQANfFqR8KGewxVKulQEU2UIBMK9bydokh7+jiBWmKR3DoIUi8IRs5yc7D/1JuXKwF
w7lHsj4FQds1PMlktMIYMwL8yXijodl3a3WoTFGSyt73w/j7nfHlWfePBvnQqumKjBV/xDJhVoYi
46u7AcjYq4Sg+Oseqg0eKFmeITMI/BWCHshnqU56Ra5FkxIT7YOtPVPsKoCiJFfAmM9U/RDN+/nJ
WapAvcVH0woFNpMWGd7yAC1CBwAtg6jgyqz1FAFgwkFQD3VNi/elX+LulHuC03BSiKlxvuegTrQ2
NQIbanOtGs/V/2HyKoWWHRCkv3B+FAyLe5AbEMAPbBk+JhUd41MW3bYvOPnhqlBpTRTwHJHKblbY
2uKkcT2QeXbkwtLCpfOWrdROSclJIiL0dE6S7wzXvy8h+xb/wKU6En/dCbY69F3QO50TYzF0X1uq
L0HUzi/g/Si2R1OMX0T1SWvCMIFIA2dKzEzkBFnAx+lFcHRQX9A9v/1lDopmR+px3U6efbW1IqMZ
7dW/MBStPr5LZEAHJ5VwlASt9IXUbJxKZSozQqJUy3Z9O7iNbxF9FVYDP0BzPCgpR0bovkCPa7g7
prAKa03wBb7cwC7zBbJyahwtJz/+xAT0sAFZGZi9RKGO4rF/Af/+guDMtRo4K/vivw0P+vjci8kA
qpcUxaUGQaH2qqbWhBQJEFad4ZrAkO5PkuQMALX1QhMlNQFbChizOjs5kRT+gowHc556f0d6HSkR
c5VbO6FHjnlHmpNOrT2JxGFZjIi4NVlfvjfpZhlymYZHszrybKrmoECFJCwAizoOmATlA4orzKV1
AK8WK8JaUOic27C9k/Tg30S97eMXdgCaQmHtHldDZubKwzue53E6RWMamLgnsb1y6IXX0JKA3e1A
X5YIcbRk8+vbqAWudo34a0aaK0F3fRC968J5V73VcZ5bsulSpwtju+zExbYPb/t6PUsH9bTok8tj
pcQ24kQLgW5WzLGluhU4qO6hKcHdm51rmUVQA0XAadB7NTmEcldMvmEJ+gub2kLtLwjWcYMTI66f
nP4lSfthMlKQtA6CiqRF3P7MdkKY7icjIb5F5euXG3n2csZSWmL4c7/k2Oi/6qoFEsIKqj5G2Ri1
2/sEsi8nl5/Wz4cmCSW+/VXusNXAK8DipCl5VrI3j9TDzU1GdwDxuLSTPjDliHL/APQ7YzKzZpNu
NOLBKq1XGvBIphWQRMyIXOUadHddNYxGrK6xlfB2ShztdComu9HpiPjbaxG6XDOSRH91gozE2v//
QcYS09LucYaQcTRp9WWbZkjor7k4wPamEtu4sKIccDLwqWMT+0oWp97bTSBJ/t5xNmTuwFXHr+Yl
u9uwStI1GimkgzPk1R/pAJZqa/t7XHN919T7vDGGLDCVhSQ55XVxXNj/D+q+6+gX6TbPjSk0mOeZ
3SOFheknZbR+eoKAKoqqtYSRYO1a/PuEoHUU4TXXAj6Ex9ZiOb800nnXx0Xg9XuDvwjD6Gi1rT9E
w3JMlCSFGizbk7OmPjO7w9xt175UNhjSR/4mFi4vInkZQn9aYKE8Cargk7gms1tnyeTayWANhroZ
iovqjHitnC2SPd/dPTu+mQfAI6gazzE+846YL35I9ITLZqgqOQvnSGu1zLGcklf4rJATduD1dd8V
5IBfHcD4KJFzLuMUOjNAcPOuIVU417QRpDuvxeiaEkA+bosHtF6cGrYc8fnW2I4EFD3RQnxdDgSy
Ktl/KkGKlABTZ1DYzLUJQnSXKP31/hvwLwl/9YW4vXtpKz+vNFuTsu+aJdJ6BHm0bLAifspp+xDn
LqTgob3jMdrK8lPXS/MfrH+LmKgYM+ndo9Y9UygrI7sZ5+clKFOyWIFGz+9dyMt6QHCWcxPP3wCy
u22BmWuxm0FjhhN6FzwRL3F2Q6zVUGPxOH8T4gnCWb4QECWbq4uoI9eeHATf7k1x568AiQB3Lfjv
Ydrxtg/Be9bll8/a+ciy/Z6AfqW53lyd4MHl5QwvxJHAafcaRczIQ9NtEsbvqWOVe9gO3TkAAfcB
IGRrRxdmErxDmMPbaeaDfITIacn2ldBt2C/rH7UMRzK0GIdEjDOMDuRNz57M7cThvhGQ/iGA9ljQ
vT6laOC+qKrJEHur7VnDiUB8/LSRcMKJVGeuhTCHVbg58Ge5nk9XZJg6xdQj1j7jxwRp0NNGbkbT
Purwy9LNidUU+yLsO7oZyFnoKo3SBgXzs4qlIwmiuSiiyVzuBi3MHcrK9msxRmP+2AcX8ZLSHIPi
7Vvr4tQkx94lzmcK3ThTzjnogDtn3YGWW2a4P7RG4qaVhtDL/jWbsp+3qmg/ee7dil3AMTcAyyfA
3AS3grArLWa+0Y5TcMfla+MQwnSWtHtKkKrBvyOxICaUc7OR3AbRecXR4CqlS+4DwglRyG+fNCUv
1VANO6ZD5BSqGRTGhAlaNUZ2j78lBGWRfcRg5kZkOmAlt1hkVhKaHQkyuh31GmolnCWK1j3/pClr
hfuxVHAYGVQV1hY/pOX2upWwxLV8xwY1cs6PKj/MuG9PIHICUOpyfADZbtn2EhDjB7gPGfJRUxrU
c6FkUnkaeWYr4tWEEjWaw2Dv1zrzDod994MgO7qLQq6YwolE62JAZoCKAo15IZWLJOa2v029b+19
a7ALcMO/VmAvYo3hXk/HfKhiaPfiCxo5TMLuAd+oQHJL5iM/ssgTAXAguGv4sNFTtGg7SWGXPwMu
9U49jdP/kg+l3vxv7MaXvKifKqE4iv7/Hx8GkTrUvraAAMatQQMzwnwndkKvV2HOGrtWDP6b+aP+
YBSIUXFObTKP0A0QTp+nmYKK8IIz5nVJ2wTGEs6Rv8wchjWdikPwcdWepcg7xe1QcUvhfEcj0FT1
RrAjvxDclw1Q5Z7nlBl8LnQPWgMeB4xCMlg7DffJoh5Sq1MhKr2cHLm2d34K/Z9gWqFHZcni8gQQ
cCUSMqFT6lp8J/KomYxb7qL8VCouhvIqM9xPbs+fU7PrFOrGeZzvHctTPFxdmbH+I21cRYN+55Y+
KJ4Z5Izbo6Dh4dxjJbtBVG+J/NV6ALdtiFpCn6cSMrZxWttDjdJXjnFZRCUZa3RFPfDmDS16BzBw
nCU6EvP53QVHe+Y8o8K9MdJ6V+6FKkbUhYHke8HXNtXXMXfrvIoNwpZEWYSZdJNxwF02MIrK6pQ4
/NaSw7cFT50eI5kDzfBydAWBE74pJQZSEz67cLDmIs00u2JlqTugEZJy23ZLSuLSpbwnXa80c1PX
hxpcWjYUggwj7QIvNynI6iKFjHGVDLIhb3NsMbzL7O74l7j2EOKsGMk1aCDgXjNOSm25rqTLTqCz
jc3FWkQJ3umaYd8EZ3ZmEmscxb1fGIQNC/2HJjDnoqT/zGPiQt2YhzIl+RSeZRdfV6D0R2zDzmYb
v8awUlAGasi+78MyfQzlMFYsYF8lU9JUxf/MwEvP8a15Hdb3nTbk9aCxuIzT8lNOMKRB28lVJHZ8
lg5GzVGZaoRN7lX9b4eYwkYW36Aca1XodR9N5h9KOTxTV3nSDPilbFIE3Gt3TbK6VpdcVvaEUdoq
WgLXx6CjL5X576tSaW9LdlyzQXkhiUnHd34VbgTLh+9d8RRyt4z3ICkvRzJPjf/LM2q7Vxn64AeQ
EH8kgRxVWD16orhERACOqUrTfWPYF9+5LgMZg8N1nrkqim7e9xNXmcNkruqX1+zpsqimIW9PtGu5
zj7JaqI9Yx75XN/VCthLlHR1lLhSfBa6qIQwbyo5J03TJYsgRkRkCoGwm9ls+SpS7VIMX3q9g4eg
CenEA+t4OWQNyMN/3XpQIfK+AmkVRKuwMdd5Sqr0qIlv4UqhVhzfNiM1aEqaJqKWURnFK6tQ7rc4
t8LE0cNBA6qzHwubdkUK2mOrSVVExKu0WbBDOc3N4GLBqFXGVhmUKJ7Qoj393a55dSImPfFmjA2C
mmGNgCIIn3jACvXLOWbsC6NoCwmPJ0YQd1S3G8goWN6Y30cjpMA95Jr8e1LF4BadtFgcDmP/niMO
/mknGU+3BCKHnteiTJvVytRQ6U+biPlJlxUuUWdegeKsw0/ZeS+ZHgxCQyUjtwlesJNLKeD8yJsl
DQ2kIrEAvudqEtViC3DdkkY7YqUZV1i3Az87is8fTqFhA3JjMpUK8AdPSqS53GQahEoUywlbpxoE
DASgVKRhR3+Kw3tHrawDqZUcr2UDwTJsEEGMLeqmmZ0m3Ac0wLNNz6horIZHV8kmrj/XkXtMT+x9
gExF/5LfPMDmI4Agt18QkF/flyh/Oa9R5Os4cAAMj/PU+N7ktOllyPafJvKZVS03JlIoL3OsrJXC
Yz6039y7DanoSYua8vsOBuT6hcP7LS9+VMkCtwjSxmON98XwfuyYC7tutb5gECseKAS9WMde3LLZ
NJh7goZqsurizyUx3pwQDPmwUyMYtYWE6VcyWSSB77wyuDBijGibha4gJF3flh9oeEHZITlrhPuK
B2zjYI1DkYRYTMjWP5Z/2kDb1Ma5N8xD2RF7MAAMwjL1MrO9pEd55Icey5gTBd6BhZ7z+eyDsIER
db9HWTnP4Edx8RIEPa0HJbNozNn5oHnTKfEhV+UIBvZIn8vJwV5JtVbkwvQz500kkHNsoG58tmKg
xIXtXEDMLoHZXJOmNBdQt7e8WOErkNv6nu4rBZZoXbkEd1FXg8dxREpVWC5kUGAythTF2Voi84Kb
COjaMUcGYABe60ks0TYRQKXiXZ5psjfpdxP1bE6Rq08qJTRFHzT7xXxY8GFVN0De6ApI9gdPAP3G
DdITdTA3KRqMIRkflF3XaXGrS/RUc55NXhm4hA4be3r+wDsocEf7KMjrhvrH0hYiIMFw5T7m1EnR
MyJteaLnLwrTKOKDE4eMVsGl2ZKZ6F+CMLK0B/yhSZ4+wSbv4l8FQQCc0Lr4yJ28dqaI2iUWMoL2
4jreK+CTDF+ajPX2GZUWtydTlrjWsRDyfSJcm6Siy2LWZNfN5sersDKZOus7xfGHy6rahIATenaM
CzLisPzdpsCUWIiokXCmvVn72OvM1wyA6//DWwx7cw9s/jIdKH6zDdGWx6BzxJvE3kT46EMCfz6K
210LlH1PTOi03N7HAbWI94sOMiB39Pi33d4YNv4YVCHM1L9VtwW3FhW66olx0U/kgjpADZwXSSgr
aeouH+R0Whru912b031s7Ao68h+jRuE/vmDzRwZshsurhlqkPb309Lths7UZB+WFzGlRP1Uf/JKA
6MHY6EFCtOENcNiP2QiHDGWLIk9V75FA/zsKpSQO3WDlu8y94LJ9/BjVQIpd4eNLrv1TQfvOpqaZ
C6ZGT35HcuOa1BfFnWOz9l3WeSxrlCwuHb6kQ69yLBx6HDjhEc8kIAWMX5Co6lQNRzJqS3Z+SXsF
Nl1DeVgQNy4Qfye1N2eessZU6MGVXveB3NLFBQ89AlObvV30A3TSXgI+f7NSGZ/aC/ryEVPcwyQ1
pzNzvAUCgPgcUIanqb694E94SeAJPI7UnEjUk6b2JtImB1IQVQkxtsepk3VrHB2TjnYC3erVRBLu
8/YjG3Y2WluTfu6P2cCVmbiIkaYMhkLgqoHdozOVbxP9P3n/u3JQ1FX8zcTcTsAa0HzZci9918Y1
8MZ4p0Phfw4UCpOVgtq7dDBO/rYSv15T+vrRU1RlyjtinFw5QCUa+9cAb2Jy26ma66Fd7tgTJH6g
CSdye8MbApXFYOvL3+E4n0rrXBSTW5f5gw6dCAAxBsss1pbfBYJTL9CYQwjPamWa26jSAuIDplRw
wU85Sc049n47g4rygQy2VZMAvOBcUhA8s7W+DCZ1zCnP1xtidZJ+f0Dw8/11w38M1pCAId4e4xsX
xM51xySdluqEdzH3ZIlcMaesAEWMpJxVgcbH3tmHeuWSuoOOXd1S8dDpWvgSfV0Wdi3falN9A+kx
xG+x2HHEgdW2ISnNUEY5pwlC7N0Kxb0AikJSBBxo5UBgJ+r2gwh/VwwJiO1C7gjdCOosUzRuLTz0
w53/PYgs+WB1fTPfchgBkBuXAqQgYrZGO32ot+aLZZfpJKbK4Co6Hle7wnKMECRFaTaI7QnNr3tM
acFgXFWhJkpg/c6N74LsQBCm10/8pWkZfkwvUHjFrqOaS7984Xco159bccy1/sYqLhDp32+CZf4M
+2aGF7O3zHLsgn13cp1yk4J+dFgs2EdzZcpPOEXhiEEEFC1POsPr8bJgvhZ23fQ9uJ9N5qPTmjaR
EVgJXzbTqOGPkJMpZuoO9lXIPUiM7xsh/9dONoLL9nxafwbnopTFemKAndooPMMXYBEXnGohloQB
z968lxDWHP7V1bXI6GT2uh0keN9KeHlLjZITr8hyGD4M+YoG4wfkj9M9EEC+2UpcZrnjOukuNi0n
MZIksKGPIBVAZPY5JXJJsd5KebXvzfm9wmqKTEuCFK6psczVxn3obI+5ySjSGyp8E9EI/TnLOq3d
9Dn18g+RKWS7y2QIiYW9ipUYwZpwmtsFgMFSbGkJ4HpyQEZ1O3x7/CxgxZzH3tuL2FDhti1zuy56
zkhbjjEQXNV44SGRb9gqXdX0SGnnXRgKECq7gpxYctBPiFm35BgCp3tH56SoRx43vbkJvas0eI+G
AtdVfWrqNXr49Ojm9I9XNTYdY48WIWx4HFyKXzQelFt9Z5mZSIqNrbHLVD0XAFLhSo4eDdn68QKk
hA0CyjRZj5A1S/3NdOAi9rWCW5IPmekVOk8Y0e6Zh/IAOl9H4VoWWW4UM6JZSdtmWm9HglMFM4vU
jt4Fz25rbAsKU6iwsymi8FapFlzJlY6Z5FAu7Y+PyKYO//31XAEEKEYtl5NWX+4h3Mzf1SQPOAyn
M92YNt6lQExNY5caq68dQX8+qFgjdvXg3CNHbkO5kyMExKA0PKDHRNOdBq9lk2BYMbU+J2SxCI5I
vD516EknTnLmsLn31YS+WHeG/2upGTrqn9vkF4k1k7wGiOJZaU/yV/2aunrKYpOibaq7lAiEzj0Q
Aww2R08BiftEE7GIrsLF3OZHrjFdiWkxu1zZ3e/4xvNEvgqPc4oeFmCcp6Y7O6p7Aqv0c+guziMc
PXdGXAI26rPh04m46uYUgw5Nc5jvMQF8DlCqBaQ56rhjiNIW6PwZPOkSs0ICyLTWccw3Uq4t7Kqq
+I2Hm2ljDfinyJpX/ajhjtBCxlstXr20NGi3aJPyfFfVZfRE/U9kgYt536pqHoXYkPcK57HsHGlK
qWLE9K3QILFw8xNBN0rnjUJdt9U9J6pu1XkWsQshkXf/3eJYl8DEH4VgNTMYBMi7H5MW+T8Oplzb
nKH718+ZRcLQrA2wdQPu7pf/MchwRcJ410CqdzvDVuBcRoePng0f+jplO3/NHDSNP98wxYYBm11j
DUQ7PFFfpEEdkxOcKVp3K01FOy3TKb3iXpixXXpxwqBVMp9+QjKRWn1tZXdsUaBowl9r0fQ5UHnt
Oy4sEIFSr3OWI8dQuiSSE9gJZY1sG9uM89pIy6WfX7qj8ziFtyS9KaPXE08pFEyBcyB7zs4nfa++
vwTXAvFu/fbQZ3HUeGCQsdECPBSvqYPYAu6WrJRN98D9PfwkQarWnuiLG9HzH1XWKOIeie677Ga2
XKb7QnAXHOWnFL/hfta9Y5pn9MXZD8juTpUe+wOgxv3warjNTpfOozFwN09bPBZoSC18iquZ0Yxy
AZoXayt8N/3y4C/YIvGJlyj8Q2NJOOCTvI2zVslkZl8Jocs5NVBKZjFPmlRo1m3d6dPseEQNSt8m
EtWHMxx7mdJbzjTGPxbUEHxZdE8K0htabb1vS2xj1p4QQPKGK+NEk4Msf+6vewCVL118BPdxdKef
sH3NbKkOOnm9p7J0ilvnLowEsAyw/bu4jgbxwZvD4hkt+nKPcQGM209zISe6xzL5eswOy5B+6fK4
eN/pWO/5ouNIRL6WHyKk8kb7t6Ebl43Q0liY752JhSVl4JcaehXTM4aaLyuuT32EUNUOcMVFusN+
+od4rxfOsmJHaLL5lFXk5ZZtWkCVaPPPkD3Doqx6tyqWYAgK+3uwVtyJqeXPYEiTowcQp0gmqIG0
ZWcF80MEPtdV17hYxQrqMEdiNcaV56XcTFH2QBavtlGv+HTU2BgNsvyHg/Deb//PaR1gCHzv8+TK
jojO0dFR2E769wnsy+ziTVDYQ4rL5oYxyhPvOps8Xd8KI64Z5db0yHb4C6cVaB2JXyO7RMg5Ar3j
MMHBkfkyeveXUud2VxyqCAqsSCgrjb+ljb3CG4HlnBnC+zvJzBeWPTF8ZvcF7FLcMCuAJN+ZIs97
CJtH4SeAfXHcK28xrR00r2jhIhjO+T3QdHm3wRS6QkLxglD9N5nCjAasvbQC8n7ML5CPHByYtFeV
p/rV8KETLbkfnCcLTUulec/mu/An7Tu+PVBgxT7spzFSscxWypxy78bqXqTGVEJdoWAvbfTSQr9H
6KHUd6G1O740+X6wI9iRB1DOqRV776kP0LbAiFgdQAYWInFHRN1jsx/ki7zbnopquWUvsA7dJfIl
ZRxcJjZ8G4gsZWpZ2DDA1vwstshaOHwq6/3HpWrBfUkK6JUCUmDEIVJ+NEMrST23EUnMqbMS3jt7
T6VPyUUIGec/3tGYJav3a/uSFXnzUwgw0ygbIRSR/t9udvI6T8sMtTMLt7HS3nvws+pURrCK75Hn
H2tRGuU1dQDt3ieVhL4AMkVmGnrFYEAkKkmS6H9IeucWqluaA1VqrjwldmCFffqozybtN9AAE2Fi
avOK2i10CqfyP50E6+ra6qZjfcUshF/JjTAYeijIq/8Q//mbhtrOtdUsUfXsfAbgU6PIWBJq1Biv
1wUQ+ASDDekpqZfIv8LlucGK2urJg8ckaPQ9y+HujNZ2LeI+X3fESYy7Q8sU0hXsJjCTOjctW5jB
87prNIOkIYkwjAKwe95niirzpN33NcSP3PG6i+Lkdo+N1jYSO9IvlKjw1wel+OLGW+hRErtcwLCP
OHI8UdLX0G4gyrdF9JXi34uO6U59x3GyYX1dzPzyCCroT45I+ZdHHg7AufeeU057iUCWPcArWqKh
LMT25WPLTs2UiugeyB8lNtRSfvNQnQHhKPeYWcd02awsCHgwZucyqFtf6QGBOpIFKGAyuyyyJgDz
Sr9uuZU7euai4bH8xggisple/xzEtJcO6lqy8AwTkaW2/kWj6CXAvgAZ3U2SM/LTTRw4KUjY5pqV
PcTsOX6acSRqkB1wfwJtjH3/D53hFpQPNT4TtZ0cwcS2xu3T3HHC9fDHfL7WQ/bELUvJKPJQF3NR
5sywATfQXMTGNj49Wd0vanL75Ys29F15weq2thzjhADTbRCi5DgBzEUbqpWpkpRHnJA3TuRpmCn+
GvC3s0ehxUeaAjcEs9m3RxeNU2a9WzCXFuNJgDgnFIjzL9SAN9BTQPZ6oKb6FpKGbaysppEZvjyV
RO1Vsof727oZn1HvDSTlr4Mqm28t4IIjrlkJWsAor6kPt2Kp8EDsInmFsslf7lSJrZx8FDuCeKHH
mPer/GRmlh0QpGzWCBE8hpx+LmStgiR/aTq8K4LKnRl67i64kIyF0STMzMk2TBnpJOPGL34dN3Rr
uPCmVG3DcGOKESq6jBeID8lygowSTkIUj0ngfhDZ77P+Pj++UGIdU9Y6tv9T3H2sWmvl6zXrHS33
5zecv0wL870/YcfRFdlGHklK94uSCgYXVETevAKJPpuKp4RMmv6u+JVdKRvSmxUVWEzap8MF2GtO
LynIO9Ya0C8chQwFunpMe1FW/VSftmcsYj5l/SdSVrPSZxMeS7PCN5VJ+Hhfdl/KjniSd0S155nC
r2hh/qG7VHWZk7CCHWqXHA3SWYUGbJ91itxUMa5dUHzK7eC+DXKHVcXGn6319FBNi2yESUrx0cQ/
NTweCnBUc9L7O2xHxuoVT2wy6z/cCxbx+VcxZxKIEH+cSrIa+6NTmHbLe+/yjKGc3BwTuiweCKW/
9b/kBa7yzPA1EgXEsWHJzmDr0+t5UKp3j7Rl2RhuRMEMcQtepBxbGwLekLDnwxmSx6DJjuJIFdcB
bW9JuNsv/5GHGPZyOaollocGQvtD5OuM69lLgzkzIuGjmyRNvHKKtJlwCelQ5xIQqlmF4rs5EHiP
dgoavcGLEoJkUUjqPlO2zc0uQ4UaaApBgr1cBSTZFHpbHMK/+hgZepV4OijM2RTuZ/m3NZD5DnNL
xqThTuSD6iSskW9gYTTLk/mNIKwdKhNJ8xx0MhCbSONjXR2JH9/S9jouILAhIge7C105dZgiHNqO
tRNq95ZYhCsUQOKAV2wECcW71k38NVSNEj6e72nDAlcZ/i/cAmibhfpGd4NBTnS6jlpr53V1iH3o
TEdP1CFv36FVAg49HixHS6RlFoKKSxpOBHSRq30uhxTb+Lh7QmOT3hyollDxWLupVC9fl8dexMFW
JP9AlsFbgnSp5vmS8z2i3Lr72J0Wb1FZPpghXaYc0KsrnNE/QXU5sabPVjEmXt8PvdRpoVrY+p6b
H9atRKcPULSGwpbwSzKwCrE2YLqQ7FbuAW0j6KBvqJnuqjPKfKS7MhlkYlgMzsDdz9Yk81TiWqH1
2DYDKp+WAlhhwKZsUFPLvaJE97Pq0IjvnZUweMUo45/EU9f1kSs9FS/wA7viH+x3ShXXIUvFrP3o
8EoSCY1CBxSTeCGHjmmgdA4NWSE530bbtLRiGTzeJ9YmY0PsgOu0hA8t2ikwhQPpzJpvMwARAcyM
imcwyWuYbQShoSplIB4k+rp9TM49LeADWmbwQ9fZaaQ5k3RNzMH/LNh4iHPMhdc5wvhpFMx88QB5
nc18m15Tx55uEawuxAtNvZKLDawomWbReFdTgXYOfsDVvZVzrdOTL266Igf8HKlYc6ny9sHR7HbB
KthPfOjiUDNQy0Gj2N9oLV1UeZtG9GdQHuF6bXmh3H3N0Mm+N/wuULbxKOerWfebWrElY4JIUAYI
oaLc5b9q4nQLoe3ycJPsBy/GkdEXUgwHT78Mv4N0S91LXx3Or1/HdfOZJ/l6WwSnIxdlld6T+4ZL
s/fFRDMud8e0nkrP1Zp8XFXo1JakVRCmky1bYhZ0oJ7zsxB3v46k9tPCtNPJr5lSxSsjVVDbcLae
NNUKr2QVqcVdRaR9J8Vxzd0U16tCEzO7dBpMp+O+ICJPgfTr5WWa8Yyi8IeUd23uTQqfMcXobZ/b
8lJN3Su+ICkGeJXTFvvJbnM71wJlgbfMTfJJJb2Y+4IM5SUjNuk3aLOOgcOtEAqFRXbRPIqUAWXO
Gv1TWh1xDRibgrmfArBa1BOa1j/PxdFA5ufdtB/DIUCV+BfRbIUgxeNF0vkWyLW8H40cdgdfPZmB
2S52bN4gL9iq2Vh6Zzw/HEhvM4ZnMiwruskr4H/DPOG9JVrwWWLtp9P2FRkTIGZmsTbHQ7FBaNaJ
Pev4nPOAzCiAwef9dtSiGop/6kBr+XPiGNEGYJuIZGtgdyavuwfaqlJoox52g29KerOPlK6ua6dy
9GjDHviQtu+b1z+zlpNGBnh+GC8m6h+dbu1bltCHFOEn9UXK/D2PEzVTS4LI20z65J0NIuEHCVtz
BITdA1Ks89kWJDpBCrAdofxpmM9kyO2RcPwwiTe8LfoUHAiURIlhTAsT/hc4Maxo9snVrAKFVYsy
HsxYa12IA+EBEn8QBIRr6yhEqMqL81XckwIYpcvc8oMDARybkzbomdfaH7J3i4IkkkPBYKMSsmUV
+NJccIk0nf/CY35wrT1cvabb6TWThsZGXBV/v6/HMYkbkl/w66E9wHMLB7uJlu474Am7F3ZeXh+J
Vgw+e0bydVpvg3mR95Vyas1TuEelgWKFkBqYeTRcZVK9/gCTyTuKKS+MhKCLCTyYUkG6zqVl74HX
pvxD75bMnxh6Ga7QG6m5XUNl3SE/Z+H0aSGOLrPMQpDrS+vjV4M2TnGHxTyt/NLDff/78O4B7uYl
okDgDg77OjtXJUDjOplOu+bWsTipTFSrAhriw451UdVaS1lK15z/5JD4P78GDYVG5vOz+bYnKtZG
8L16mnPqpRGoJmf+PmfDvGiYB+685pGJw6wdZfNSH/NlpHzXT/RZAQrDFoA3z0LUN5fn+V5bLYij
KkIJ8ZIMmfkYIqoLn9x+69bvbZ7gmBJY8g6f/3Q0EXOPa6POz5o0HYkMsNbOmAa1+zSo2IG7Bz8G
TFy02YoGHy95TJyxsJqGXhLUtqJE3rGmWXqwo1ChYT2cP9x6J7cvGrzyihUIE6q1jyoGBWcofiVR
MXRXB2QNA8csQ7aNCyz/DRY1onyMn/nKJntft8Ql4OqKRHUZ7tiePyFib9YNCHEGAu/mddDrStlH
Oo+hww8nhzOUsKTnC3bJrveyv0lgD293jDUIXbi/30VrG+F+gH5lykrR0zyvztEvRwWqkm6+bO0U
6Z5J6inlA9ZY8w9jIGgpOT3fVDm0s2p0F1Ht5xuWklGYmhjskEQcXkUgz1nZ+as9uRnJBgavytSO
rlW0THqq2mp3kL+sjYDekmn/XtvnFyjm8IaJOeEmD3zntRL82XHlfzpITUM16Ulyr7PpVfxMGTqO
LWpbEdxFBiHRYFufl+PHwYURaN40/tbrF9YDi3+nt++C3o4VNnEr8GzdtdVmzai9YHAC8D8vwP7e
PWHGJ6NHgvJqko3jyJkHyOl2l39PBiQ1BoPZY9JdbqzcI3CrAstPT/43y8xTYAJLXfev/blFYBlx
4SXkhQRXUId+P60YFA4hVzc9N7ictoL63EdOgwkSaRYsak47tIvelVv5dE+NukvKXgTJexjMlFQY
N0lBlH4kZsSK4sMEovBFHMVPN4076rkjx1kDKqMo3gA7hocABqIFKKl/wwic16zOGrff/AYPEJXd
Ll0ydF12XcCI0QNF+fxFj8dkJ9D/YkjDl3YAk2psB3YfpZjhdtUvQpILHCU1/N2QIyD+VlvvmTTN
2Br8UkhSIaAPaqYPqkU8B6aeVlCRM0bHK9jrmw06T6OIENOGNdSHMJqgd+6w2wRRBYfOucSUDtMW
Gms4hQQwcbWNsWQ7v32iFQQ6j1Q7nG1eNakRcCQ15rbr8TgIvhUfO7jJcFbtSgkTs4G6w9Wi6ZPj
Oc29Rx1q4ZRB0SfHAhSGFQJPURNd1+Hsc8LEbfvy5+swavTOHT0FCZpzUrMS4cEeFDF+KAAU0DUX
ARAvhIrJMGpN/Ta9HP2Za39K7N2/Eyk2Yw/oZ1secfyI4UvORSj/KTdclfhYvpszl2z+FnyqgnKP
P7mC0wBXTkJSbwOcSUqEU40Q0cDpI25AW0yiegnwrWLuFfU+deUDj4F6Afv3xwfyDnyApPLai5MX
FXxq/9z7m7v4ER775uZNzOl96gUQN87/Si0SIh0gjLsbEv8UzUhIjMmhloyLbTkbD/G4H6LlxsHI
RmBDQeluqnDvNIP04FtAXB9eaCRovwvXZzTpuQ9AXDvGZPNq8PlbEob3zfD42/0Ra5hjpdgPE02r
IIL9cD8DzV+rr/fgOfrdtMaogopCH2Jfpg61CkSZ7JY61b3uryyTq/t/iHQR6ON3LkSAOUSqV2Sz
vkrYuTlvruzwoxWYdmnDRTFZmPmOMCANt7lPP1eN5uFVoTDLs2d/h5uEG1ANDU38OFyWix98uncK
BfaF1JuYtcD620cqGWLnJh3LYUNV6DbUfPGJpnUEuAs5bT9SKPvfN9WMF+yN4aDPR8G0wtveToDQ
EWbQZ/KTHnhsbDpFK8ObAvjo9GRzjJcVgi5rqGX9aZH1bXG2GChR2ltnf4Fg6Iw1lft39Vmvy6EL
DsJbPF3k6tk89mEWvD89XwMWtOoPPRfCgHnQTsFU4pxqMs7fhxZMJT0TmaYPHJpGyS2KKpvlxJU7
3pgl7gwrYQIcuaVeRgsJz/dJnwDgc4u2nt3g2Y7a7JKCgixjP8T91ZOmfU3FVAV5QBkC47qbx6QG
a6xHEFEOiMAoC5hblAT9XppylHYi+9O3th0r6LYpI+MpL4UQlGLw244m/tOb+FJ+m6ppOat11klo
BxszzCMFfKSi4VQ+uG2AKWU+qSpUBGCI7Y2NtdrfarXUiSoi3K83LA6g1tOuPBEeAa9z0dAQIFee
KbQ5H1sBmL71z7EYQEZXBo3BefqXjRiIc++H0uF80X7A1hzTm6vPo1xmM+/Td4iIUu2B17OXFdBG
xBOp8lWO/eib/5wjGUYdTxdg0dviTjxKdakjYsYuDAWe5uM0D4fyDL4l7ic0mOArmW0I/uA5Skfc
ea9otUdKaZqgioG7crx0J2jBfmJl3OzLl0CKTOqmhQdPnt3X8hlQnB/Uc2fZaetx++e06SeMoH2L
D42CMmSKyuBFohtZVjGonNPRdF3AahbZyBV8gtpYrkFGwwQv+asqGkmweTayPCHtzTzH1sDjaoVZ
OQ3SzKEguLjEV4C4yl5OixjiDZgYVXovbpP3oD8mxdNUNlUPfDkf6PeanRTnp1mOkruNisIjYnPU
Jdd+Iyt9DjQXenongTrbSQqXbQOL/Rv19Zii/a6hqCNo5nLWNWp4Eaxn4Tunp9TyKZSN7QIa8g0Z
8RB/biXqxRuY1JBZc0aIvbhMJzhskOq1JHz1Al4Nq9q4VfomvkxD9nTdQc/q3CuFg98OjvUOVmsc
qZGAfyhv+XdW9QCjdn2ERc8g7dYt2ragCTqFTxdHU66qTm7IT3l6W5eLHOVbrfrGS1nq3UXtVPkR
00Kahmkn749Lzf4t0gDFt35cGAg4besyuYFyfqW2PBoCjGX/n+uUt2hpSUCUd0XQ5srSChgJxcWj
USXo4V+XK+NcqsPjSHsZ4W5XSz9JKpiUB0SKTs0IRWBX72dmg5AKQucitZP9E7QfSYYE+/hfDNy5
zLni62jr+jVf3wRCnbQP9WjWAsq2e9d47QoyGDNvnGeHd3HQS5O66eepOt25zIEcf9yF/AQuwSu5
/WMPsFupDSCUzJsk3ffrMS+pQvT170VZ5s36CAJ1mbiwA0znwIIvZST/3gwLeTNGkdEL869aT60g
WBuKHU4Q/jSCM3K/MkdQvfo8zcELxtoqN6nfko8f4swLApRFlTjhFY9acn+Hx7mwf5/kBTcbssaY
srHTYLQlUyY7DPyBf57T8ur/OukcIvqj0Jxd7IB55Z+D9MU1becFI1biKUugpjZ6cW3+l/S6wDaw
HkTpCRojUs9uUI4uLQWijpQlPaQe0LjviH1km8Q8qoTwNBjzp/U2fp37+XKlu3jJOYk3zaWp3IpC
52berQz8QeubiTOUHxrJlfq9iQomTl/xvKgVktrcPyaB6TroLOOr6oUXUlkY+Uw06nzSne1llZHf
vfY3c3cx1j3Xm/LcJQGyB3vBTEVLS9xaP/mEQBI9wBZ82dbOrktrg9sL2QT5GaV8o5lAOc7zpeIz
kgFG5Um7Uln4Jt3bwApJy19lzmsbLdr6vbhl+92pEGAcUZ2UohNBsIvOC/1Cwp/N8ZwY3RZAQ6VW
zjL98aN+nPOaQavCxq94RYJRZzSV6SlYAD/c3ThKvrSEW1bKettOsg2P0ribxVge0c2AETGvNTKs
EBiYcM/z5U0Uw9BYVVFi8UrLtL9Lh45JnAGdDki03xYMs5Cftze+JYBgv3P8HXq6fOIrcK2BVM02
FdERyGxS68tqS385X9KOSggdcIp323VvwaTldM9lcQWKk5hVeWWmI98EE/10fp0a9yqK136X4OOg
vhbTrqtkTMHvRyt5ZfUdoKpo8V1gb4Fn6RAEsRjZwQaYasbDkTkQaJt2DMR8TNhogOizMrXJ8BOD
LSpqSd9lIHN2yiuY6mBs8AhLQFqHzAUZx6Qx2F64hfgxP/llTdLQxwo5xZHCHVNoXl7mk1wXnsGC
BdLpGj0QwQ+HX3y4gOx3fenXM+4bpv0su/zRG5+YO7W6dbMDzsrWVcX+3jNP+heWesJRRdsItRF7
fh2+iNwfvg+ejONKM+OXKKhjxEcClH43G4tOP+oTuKhm5fYwiZ18jwiNcklGyvu0UIun0hp2RHvX
olFPAMpFuhuhvSD+IJAWY2p4ocUN0/BQ5KIARiVn8Jtg647PloUBujRi/p31pJcoKN2UJjZeGE4C
uKkHsCFjtSFncfk1SQnfVROuleZ5hRnqMsLLF5JNzmFfCX2GWLy8zl6lsh+zciqCmj/MXvvE7Mhz
g3Wm8NFl8fMeLcCreRbh5G4NNeI6v/kGlpGpcXhWTDIYUtfAFWDXuSUyLWkpk1y2m3ERhi2Dqx4h
DwUBxQnfBQLjlKQHuCnHjt8OI+CW84ND3vCmgvFV41Rw4e976gWsVItNsrH3Sf+73dBx7ypOcvSY
l5ABxx9Xscs+9FBNv1JUjacuRlSSHCwkNCYtP4je8e/uqR6YkylbVS+GEuj13fQOy9fKzwYiJqsW
ABoW1sIJ2ss9Lv8wDFai1QgK+p1PfzQxoVGGOD+bgvR3R0drRPdxDfUTRB/O5bId2w9pCX6EDJQ9
hd1xduXht3GApZHc6hZalFZjM+8nx7o89P5kIgxo8xghgXM77VGTvEqe6oqhxJ7ba4PTDmuZ2eIY
CNseM6kEOaITcgk6xnmnNxORdrVccEi63GO0+FBOP2sSDmxUfhnN9/KyVZkzWZkzDYNd+DnT5hny
F1cG+d6KCUSFANMUkIbSLe2P/liVitDDr2A8NoH0icF3QE55O0MJAmeGJMLUBUL6wZ7a+FWexUJG
3AZamxdgnRkBCBurU11FkPqebUzj+IhBYu+f9na1hJJ8SUhpHqibJECjbbYwDZbS7/fyNngVq4zc
OW1+/etOmeEb8klaGRw8YGwXlG4D6bQzeJjfSwNN2nQzO6YGPhtJ97HUvuWBAC9dNjQYpM2awwAG
qSS4WvTFJVX4TE1+Tnx1PLjSsE1LeBc5jxReLkpjunwMe3PX2dCY009r0U3g3CiTISheFjXspSsN
4O2IM1bvsw8IfK7szxq2bWbwzqEikw0GlDdj9k0y+GbnXYxTeGWWe5D/GAQK78//8ijpymm6o5ol
GrU6uxbrwXy0X+TE1ZcXkU/LhUTEs4xOyx2EpLlFBNpUdI9M6eisgqQVxeMoAVoMQ5DpUczlSt+U
afzikLwqv84gPWijMlj/GwD2fdGBzM5sY1J8lD0/r+uV0srPUE7feytotzOI4HQhfWty+A2igtas
9vv1JV54+upFRdcTNvi6A2onmBuF6XmdexUyhgUcEXuTDPa8awLR7p8CtDJMatk+396M+Yq36Vhx
YZPTOYTjT7uMuHdAsnCsUmp2vBTA3nE1WQoa9wTCbychuMbmf40zRr1kMQ04OWbcJ4UL1wDLFjtn
QdAVCvFgBDVTlY3IrO7uy8k9HosE0F3pzaWVuV/djuxfJQ1QUvRnkYTvbTsrWshutQvkKGMVQrnD
vHhLsWA09kQ6FzEtcv5rUnv8guA3G681bxgCk8T+MzaONe6mzVNK8SwjTCV+Q8sf+2RjnrjHRSgZ
P5MysLc9794GtLUCK1MZ3kWKZM5OLcMVpn56DxKrivuKSbmJwIjlT1hht7K6fY8CWIh9Qxzc6KMK
G6U9SVyv1N5QB+oFZK9JRfaMwFh0FRWzhgMacTLFy7RKHphHp4L0qBVGAo+Pxux+92uBeL+pj3Qm
GYm1iQ9ZKyYowuYBj4Zh5+hm+tla94Oq11hiPgi7gl2eAgIR76H1iP251Zr3jzRCwdNolnRHz/Vg
0WawsCMl2spDhe7VbmB6vHAHexIEV2dk47u24H33E0Xe2yuS4PE1o461qEMb/RVk99DlHRJ6PbaT
9DqnKJqOVotxWZZyjnKvTvtzCUXZDwEJRcHpiPkai7WYzuPONeCpiTQu5d1VuZuVKDKweUjOXWtX
A1ZA5XXsuWW4GoTsWDzB8uQKDFbCp0DZgppvvIwTHp38wpGNuVwtyQ52A+rGs1DB4vgpCoFyK9vB
KJA4LJHZ/zi88UNHJPnH0cyL+uzOWydqeGA0BnU/WhThw/OC/tFMEuDelUHDNO8GEELYfitzLxiy
ra8d9Y/JOHNvdmfPYLcAEbMvrdS3MDlXMmQfisb3M/SEksBkoUrLaCNhqaIDTytHgaBFBQ+6eJD+
VVbO+VqwhfNlPFuYhp9wI9zLh0ZXrbyIntpiKVXRC6nfYnoHEcV/RHPhsn8pJeM8JuBUtGHcioJ0
lN74z0rH+PmEWAnW0qrxqZfyJxW2YmYKBuvhy3BFw2rWUhj4Rr/8NU61OmbqDYAC6RVQRlKAfnJF
HfT88gTXU3mou3v0UAhI0FAbfneUoJDn9QWFCvMrb5tuiAbqZP1IioEoeDy34Q1WscFqDtHGS9Us
g5FHUE43tNTbikinP8nwWKySJsOhljF+vUqOqPObAMjAUziSktZFvGkF8MDVtMXitGeoeMOZfk2f
Qt88mKSV9G51Y1hUS0eLfmE+X2qIthuGbnmO7sDOAUg9Lj5RFTqiarrndxkEjsC541MOojMfJhPx
8cH0ybAoiX+KATIFn/unt8O292ctiFiyj+A/umj7ZIVxdJfwK811+1O1l0g6mu3ukaosyapUf9mn
rDXDN5yYJ1L0d+/M0/3uDlcFDGoD74aj+bqqcL55yENy7joLX1k6oTSYGYFeVkwjGik0T8fFpJGV
wboPsiOEpgbeQeyKuLSDaBC7AiNL05qXHgw/1gdxKvhm8eaLCG7XO4VdebE+yhUdhHdmex1I6atX
9+3Gu5zver4RpxF3tydDfDB96b8JI+mylydrrKY5ji53d8IE3cUt1ABRygqNh+R7JkKZD6K46XOq
j2ugW6JsIFGtpmpNHlb3pP8lqzI0779eQoUUg0ZensN5LwLFJy50SUBGouzo3w5HenR3v67WPRpR
SW2F6RKUv6+6uXSBlxWth43nWrQHmCxqRK5w+UYQhOuaTVK9V8ZESK4tsm9gR4u+SzqnKD3ChndS
unrxHI0f/j0DMxEWboeGt5HlS0MmjbVOqzkY/X9lwlJ+IBnOWh/uqbymRPuYFw74EnxUaE2Zt5BV
xcqxKnfuhLIDFEMKskv3LMoIM5xxqJAf426KgQ0ANzN+IAnMOONGWf9T5jiMdq7BLD+PWd/3if4j
sQqQF6s9QWQ+6PuqSeriJrYtbA8HKWBVf1pYWL2qTvZ2/wKam/pCOKg4jS+kXCOZg8tYHxmv6Wgy
xLz8k05J8JZJ51CokbUQg1GII/GXcAr5C3/aqyJaQwYuZsDSBHMJ0JP2wRXtePxsTcQzApe6mWCg
T7t5Qs/wptx66H6R5FXfO2drvPImSGnJLcqoEg78WLFfItPuzUcAQtS0hdMV0HRL6EvkP5Az78tG
KJ3SvIe/db9XkzN5zBIEauR525qIMxQbr+lQV4DmiVcExxZPG0nAMi5PH8aXYsmwnZRyVZwaM5ka
XA7BZWzMRmTkQNPxw75X3Kimbc03+8UtrvhQlF+ILZQLsFDWAuVPiYm3uPU5dQaTmxe5wToe/epH
3yFUaN+0XNsNqyUsfchLjAObaOQxnJl6sgCXM5YH+fxjWxYhk1lgm6LuPWK+8iprbtJgugGStFtJ
qWQrwoCQLq7BeDYlJh85fauhCOmNTuuTZqJJ0p847heAY28FPUraQZtG7nTWA2WmZKe/YU0gh+dy
si5fmAsoDS2ZKdnOrS6qFFBmFBG4ZkSGD4NFTBQ6HXVEY60rI9oL5BCo6gNS238x28mvMnfCsUp1
eLcHCudOvn4312edOZeCKrBAHloZMLSCzp4SO0Fi8+sPn+SYneIZzI1JY090NE9kPG9CiwRKt9JM
K976zUzL3xWvkNrhyg6hb6Xe94YDNXsdSkqkFEdtIR6L8Wk/ZzcWMrWS7Roi2ZaliHLMEhwDZ4do
tM17TH/KQMSD9f53jlWYsO4YfSn5vZ1J5LhHKUphFn4T75UJZUXsOXGqGk2EIAzpMmaNdPX6j5ns
0XjbMNhI0OISQf6wYOxm7LCcfkrT05jz9ahkUxw826oaZ6iKfz7w/eIpx2H+b1Ff90BB/itCdtHs
oCS0sWBma/FF17QV74oY0PKAWjQJM4Q5oSzL+eiZHxgv1l2lnKXHHwMTtx/by/84NnUx/UNIm0a3
tV8p4o8eN6KqhxNL2y1odaHRR1Nf8wnpCpE3Ela4+VDXOWdNCE+THG03sMHWoluwhxV/+tDPl82v
swmG6jpU6hl93HHXJ0Ot7ple0/9WZmnWEkQarAZwrNeaHW+GoroBBLfEOANEckKZCM4NGeZ2JV2V
QdNt1AHykzs/g0JbAC+la+Sy6pkFR55Ce/ytjXemtRIw69PJIi80rOicPpFvJRRe4Qrys9IKeGTc
rnz9FzM/+tXsqNf3Dyj4XskP76EHPujIihwFNLT2Ze7gvvlvYfE7uaqpd8axK+viKZMSyf+tYTqs
YXt+XbObghTv5O+Xnr/tKiMxlrD3hK/7cvlCXIhi0aZFAl9U02Xyg8IkySHWIJ/XNJgyPu+nMlSS
QV80dow9PedHA0BUfg8etPS9+9qx1SKkEDZJeE9KBD5NZZ690H9HJMFikd44K/Z3ZVMk8E6vjwk0
43tKvmEs1ozh6dOsVFlFTbdhi8wCi6l1PYLRg0AC0D8FXmcnzT2u54pjJed9h5w4vqbCp/Z4h4tK
qhzvNts4qdfIiSkmnqM8o9Cr37N9WyKJLs3vcRP+4pvdGdZtqsvI2kT4KlSwod/QLz+KWTptbZNH
ggpdnjY63ckv6SR6UuqNtHGIky7qfYN08FUYloYuZgp0bPvlK48laIl7vK901ES3qGNlUDMlBy4o
RwIR1L5Jdfzu7SUWK0p1RHBveUU/SqC+mQO75Vcip1lXtoBqOAkWs7AMa/zfJDuv2x2tHEUNude+
pFhqEMkfibJLADa/0SKtZ9nAy2xX8BX5kSirzPcUikf+/2QQWQV5sOiIUzqx1pIlWU4ahVrxMY0B
hrUultLbD5A4pi3rX57srIzfnSbCkIhBAO9rkgJXyArrtJ+24bWSLQRRAhuAqeowJijPfCMgazoe
CcNChOfNJbN4k1jUTOmwnLuVuz6Tm6O8HzPe7IEvMR2FgmB4eXAs9BKJQWW5EGBgiIo7Pu1530iC
gK2SEjHuoXYV3RoSqD0MwIBIyqLPqdtIWo7VasUkF2+eZ5jA5zx2CKxBULqVY1ypB2uvPIs3pnHb
AfOddEtvf09ojni7heDbFlRd302S57BJURJvuB7fmaW2p2yyEyWqPXeAXmW09zgvIduZ9dMl8C0w
5rXcX4oXbQ2Y0nji5KPIfJDJ2p9rS+/Q1yCt4Adex70D2dcngA3tbOY4rDOs6FwFWts0+aFZr1f3
wh3CiF3VexOAA9LBaARZn39YkEPTlE/40X9ulm9G5QHJsKxVIz97aiPvTGZUcF5ALCh008wpuMhO
xUZVTFcw3KqtySc9IL94EYfBRdAIXCv3f1At+Rt8zGZv0ugeu/nhoQhAHMAnGECDMuA934amM/oZ
esAEx+yLKQWB4/Qyx25T/pjDiD9olOjqcni4xXfadTvw/bsbPzE+CunpECxtU8ZHVivx10vnwN7q
np+uPvBUTJvnIRtl57TUmiAjWt+/XI/Ji8WOK5PIPy7fqpK3ofFdt3RvZGIuVxArX9TLlen7iD2G
z21xIylWYBGBFDOUBOEzCrciTAoo+/7tET/f5rcHngoBsDZIufecrvttLTgF8KUkSQ3xhXMVuxrz
EvZE2m662idVac2s6+k5yj9i5O8yJGB1LoSeDOJopLx5QXXdhkLyMqEaZM/v8BM1ipBb/SIJAtQs
bHLUpnbPnL11wX4hSpTleATnVYRzM0uVjRJqBk8V/mKuehmVf93j1hJZJrMtvwEq4nF8lh47P6EU
yxnUIty6l28ejkfkU/eiTvDZsESysT+3H1slUUrRmLZqhmDEmBSw7ftcGEVlzehX7FmGSxGGqI0Z
UlXoM21ITz4glCBCfmVVYqKxdM1eCpnEIvkMrEDN7xQFYen0drJ65Q+HWXmrMnYUO35jxThhMy6q
D9SdAXuqyFcBYjYLLy4pfF+iTl2ghYN5Gx8ufSl+7UB9DphM/OXzMZHTOgN/wukcLVLWql2dIVWW
RracyAEiQq2AFxX4n0PCTbk3wiwAVRqEIBVrRk9wUXQP4w4w4wnQYwIxxLL0yffvDvcFCTa+Zh9K
QF5JCXlJIo6S4hbB+HHYsv3iFX1Wgi5D+z0n5DFsMhK+FjpU9IiGDn+KbOkcty9znYnjS+noJrM/
wGOexZbEskdLSZvgt/Oa44Pdp0KY42G+Cxb3NEbb0Qi3VKGJChAMBDWkBb8tfJ9wluMuO2cQdTI0
jdZLm+fx2tYvKdWqRRprMDHUhPzvV4trFMoMjMrDWQsPj+fRbaz5pLO4civ/U+UvHVPUdc0tFl1k
GMFuid68tn+/5/Ncx/ddURUkInGxDf1/cWEPzwDGkmaMqo7S6Qa9voAVHs4yi3Ctr39sdhe5nwEG
Rp9cAkGIaROqy7OLannLot1oV8Jwfy2NGrXBU40Wl+oa8dqHNlfqpyd2nr/F3mPYjYhZqqlwhBj6
sKQnacyCa6ofdMi0xGwX8QMX9tOVNL3J4SL0OJmbVN6kFSpInLpG2cW3t+JxlUIb5ZYnpAx8KtCe
vl2f5ocGEKvw2LTyFPALgXRUUTKoWMnpEJ12Ay+2W6b1mU4/Z+2Y7Tx++bC3STYkBVYbvPJyzVIc
uhadqV3qug8N4TPQGmKpzWFywie801lTqjpvFoUxOY9IQo/Q5SnTNa7HYHKZhHhHamHPFog4xxm4
KzMSD6iE1L7HqJ4BJpTOXoOuiqmL+86P7OLnRT9TlCqh4hM2qeK5rmct9JJYIIcNqx0f5rvZBMoL
j0xWAviED+ffkCACCnA3gzVhWnZhCFswZ7env7Cuo3KsEzZwU4rzomV55CV1sQzqesCWD9YV4yEK
ULr/g35ddN/ypjAV/n9ahvMB76SB6pAgCb38Q7bsa8+VRjPc5VevAzTwyoP0b8iNSOLe+BY2e1Pq
iwxrrDLw4i+Eh2+sGo9G9fa8mNdbwcrbgb3bgqc1mUdvCscLztLhz/9LhMWrOOSjhAtWxPaHQDwQ
dfBOyWfOzfebX4hMT7Zt9RfL3mgy5dnZAgUN6qjVrllnN2vK0EwhpRSTOBS5FKKOKsBtlxPzUjJu
QHhHDRhjvQA9hL+9K2lzqpbIyD9K8P745WW3GmGFOdJ2jQ4EoRHhm3yJ2d66KStqt2KBKZb4NQXO
IjHLCnT3ODcL7BRYPO0qHKsAlA+2OwVBjiCccsOQvCYWJN1bl0nXQzQoNUopmnpSJLiOwD4Sxr5A
6S40zn5oD/b9T98/vPbJJ0BZwwM0FRBzw+Zq0nu6STo8XdZgbj22u94xaGxpIWjzK8uxtFYLp0Qx
jt4g6H/CVOJgPBIZeu50WoMkCcIg5cOAmgZBRVYGoIdLO87EVH6WGa/KNZOwwjIQoaxfmc570Uyv
U6NEKx42LaTQfcb8Jba9dLtliW9mV48pNmnDAIJGII7Nbpx0GytNyqG33T1srcM2gmPXJJ+6KF6T
kTvspkKsLm3p1TPr+O24DZ/7ue+V4lHe+DzXf094Apr6BNTML+fXtIijnXkhtu+KqaeebNy537Rq
97GnfoVHF40RBMQOdtICc2fnscIJ69fMKpN0otQAol0VJwQPDHczz1tfB7LLrlKLx1dGx0yPhk/F
1wxjdTzoC7E5/ELVx7soLS8NECpAdTgVe7A4K/dyrcFFy/WEUWb2HQ/cB2aA1OgOhOTWozda4uYt
Jbhngo88txZktCNHomOAjlTGynGxRbRArlgmheNclFWxdZSGgElsBS+d5RPeDH5yEfqzR3sfil0k
fYsb8u44Momndriev7Rhs2qnSngrjXks6iASCK1VKpbcJAkqkCQTzyJ7Tj7K7KVJ92jXijxJ7dQL
8ja6fsnq4tngVYjzWGHBQU9XfDwx/mC2URmYVdf/pbTppC/ZIDJFIPN9f3xSkJDU14Ytuq4gn2SW
nfEh8Q0dk45YPoiUOTQy+uJJSWqwsDFlDmPat0f9xvaZ5cUTNQOPHq5BtY2z7hmYktg8Kg2qPucg
uiBp29u018/D2lxGK/Pem2l5HhTE/OjmT+7y2SsJIb35/xYf3u30Ee+AHEabtHtwe0MrumA1m7BR
FtnAKpaJUJPvFo47GvyBkoyuZTk4G6tFZfN3vwMD8RUYR0Ou10ejmpNa/ZmsF5IgthJcVYe58U+B
dWTMi+sbwDnhP8ZRIJ1V7MZqpqikKPEJcekqC18ygbqGYAF67bxfxWnLNps47RFEhgEad1jX5Xr2
R8EbHsk6txm5HXPPJXzGkFGZNL2VjErg2Vz56/Y5mPM0yemUMDv4njqD3H14tOWhAPmDrffTtTxB
faqGU5spTAiXA5aHmsCLuN8/cUMSyyxVxsf9zkAX9MFzGBaEyXzD3ZkJH1KQEbO7DXAJIeDMrDuz
c2voHIkUKuA50DYaUYlu1vwQzzfN+i5fs+THQmWmVsQ+zrJAK4L4la0MaENuLIlG37Pk1gs8KDvb
0Zuh2x6z3ji508axpJOTs730v1BQ7CSySr7/pfr9utkkRShSv0aMKXSRqLrCEQLHKULusM466w8O
a4JitltnqRjlBMoDoOaoL2oZgccmvpf3wUl/pZ7LN+KE3zEa6CTRhhyF1+y8KoL0+645OgnEFjUJ
RkLjFAFRiq7iCWHIZ5ueJ0SnvVPRpDgRbJR4NpwUArh29xxiCIYVBh8gV9hsjJzTTJ9DpVFaX/sf
NB6xSDyZ6/8wmazSPFUj3ih5hldPXo+eBAdnN3p+UUg/sYqxcCndwAxx3bdbDWmLiaMmWHXyEdOp
wXZ/Kj7PfwVLv03uYJIcGg+Uwp2McIhew0KaTqaeJSVM/jESX6/nMRakWfm2mL231e/QVeZ6w67I
/SPXETbo/+Vi7jXOB5X9TQkCzuFBHZOwKhjfj4lC1dzAdWUuSjWKgzfi6Br0c9omguwoGUMo69tj
ruG2oWDusL5ZYyMNWYtUThBhj+7N4qBhwrofKr0++VnmAqxsQ0tfRn4Nf9YwpEgr9Jps3gnu9ZtA
l4TKVrfQ2N1OecBHOOQA4ZYhzQBU48UzXZjVTYObuk4nSgyR9GrlDtt4MAHerx3pqHsQzfngYcsi
OLon8NYG18hvzeryGWPaUAif3uxNOSH+KeaBgxOjahYPwkzzZTqumNxokbNVUCd2Ls6bwLFvea+J
p0OIsEyi97Sg03NtYcsmI1LveOY/hfon5stOiLDJvajK1O7peJBAiLXXGaDbGM/+r9mGhlHnDlBV
iEL676Wg7TirMojqrH5sfs5lcKZwy4q4w2vcWYXBueeWrkiAl1g233vIZ4BxbMPTZygdOU3n0w5Z
Dm1sY8YPca/4dUtfYZd8RXh0SnoTyhPpzceXxGfA99vvEQrY4vNDCUXbd2KWGcHGTJlhNUn4zwmU
zq66ZJBAC7+ZrAaCCfsmPdT9usOVH1TrzHQfm8ojcvfriHGE3wnho8baESFj9lyuvb8pQeBwCCDw
Qvsoq0di/HLmgbCiybQUNYsvyR3Kfmw3imnE0hWfyAzd2/FRl91V3sIw5a1ARmTut14TvG8wTmKi
iyf6wOXxoQJZNtUQEUie2x9+1VtSHGNGZZ5FhlgQb3vtgyhu6QW6Vn6b2ZMI7lji0TLMhQ6/kB2b
8Vu6wsz608C5DRL+xwJ4i7Ji3vo/pStw/ZzT/AnaKwFRn/QI5v3R4BeRAH1aNuBDwdmRhgBv6dg0
/AZRNWiNNTJh3MwkMP3H3pOVZWfyZXEaNzlf2Fw3DdCqkUE3AgrTN9BOXMS4quBgtcPcAWYayjGz
jc8swV6sBqo7DTHOw+AWnkLy1bHZW3rKpUbJXD3NhyOXYSULngl+36/ICX6ze3Vr0C064GphOA+/
a0U2U/h1vNGZnIgacS1utVTHD3MzzqHS9FpeQRgkuzuz43c4U1cyk2wI8HD6dO1n2VkF71A+mVKL
HmsiRGBMIpB+/RsEYAtGcdQfnqcX0uxBHKhyXWYvty74DAQaL11xESZt1OxQNks0X1SZo6M5VvHH
Ba5N+bLvkIn5oLZ+FSXwq5v5BVOJpTA8/YAzyEu5YKxZw3xxncFk21N1BcDXrfiMkghm+2URLaYL
1simRnZ1h5mhff+FHghweAiRLRZ8Zj2KX0uJE8GkjjCnMGuq/G1IGp25wU0Xfy+px/LmdikuS6Dh
a36NGohx/nzuy4zIKa4IaeiZnpJGJqgzIsifDqLVwxCWPsKaIkQ7/HJJUjqZ6HYWdMw/YJvdWkUL
UPGClFepK6d8qnwSAaOiOf6ZOoCwk4fRvDoxmJxPrAs0e+EiFLFwa08Ep9VajGHXDJnl7IOcE0wV
+vy6ju+uTam+kAOMxALPWWH/1PUZCVshG46oD4vwWYizKmZ+Up3tKVW+L5e2evqgIIg0SFtkXtAw
BSDlL/rG8nctTFdHoAtyPpHIFJfia9ODb014jTalT9O/whvTN+rTtfMQVlz3ScNXXm5ft7quAeuA
KICK2DUF1F9+3i/AK6lSAJyIkPqm2tyK7DbPIdBpL/3WVkygbnOgyBMU9WYzZv7jf0sAPWyer4FY
H5IoNyeCOjStmkHiIhjxNRJQ0SGkjJtyWgoRbjxX1DVol148zUAaUw7EFn7AxxPfEEZ5tud0gFc4
g5vcMq9zUpdwMeTrPb33u2Fg+LEJqX+Nl9Wivbroj1UOygenpj6MezXvSPKALXFr4p4I/jEPjiR4
Qkq/SDJSYHrUYahd+dt0eRGYvNhhWX5O6HcCnCqjIq+mZ+YNATmVIywDIuVkx+UbUAzbFoYdAGy4
54pW8RBzWWX9sKPInbJX9vE7VTsAomsCjFSSwdKGi0MhWKDbauPIBVX1QEHHZaFR9V5zHK2OZja9
1ZIVWd1SBcb6NxabGcvgTrBkwH2j6o0//Uog+KOLfIcXtNo36FfAS1Mjc4TorrWf8K+Krk6aBm4N
/YjcYVaO6J7PZ1G9LKP9r7RRCb9P5U9+Tcy2OIL2+WWsikkdwKonUQgqd1Kki32KSbz4aFJr+rci
o1LTaNEVtq8n7L1ICf9RqpEP+p2Ui2w+1xcRLslzHvgqZFxvgDLlPGNu+oSpLZ38riDct+Sc3H+G
eKfSPOBCyRXcl50ha9eJVRLAy5tOU8/mEiFX3p/Z4+VPZTdyWdDKQivkm5eh03QgiRUjJoPA+1lu
lLaeEMuSs2vQoKPwbh+LojqjRjvdtZVL3Zkv90jusDjE34YdHZ+6OXSU18011/0mkwfjN4ZbkAoC
0J/nxFNGesKCSHWvI5Poh4hopPZwB1U7vHWACrYoektFrRTBOjeBiiy9pcysw5L9h+sD24d1L2/j
nSepHAeVwONxzTORw9dhkL9XuyTjefCwckT5gHLed50Kz+g6TpysRA5rd6I/QbFun5aRc+Ve5Aal
4jbDnDcGKFuMTSv4w6zU3iLzCRFop/ACzLF+sTdQQoumrN8thJq/8OGvtVTC38zsoh326fLMHADK
qjL6iQBJrrHB3NiC/+WX8Tkqo3yKMB9wANPqYAwzsSYomuaL981mNK6GKQlL8kTJmiqC5kSSkF0h
uVeJE1w/lgMiuGallM8p+WoiTUXUMNxDt1PkM4Ifg65wO/yePaTnTyHQ82znPjPBcReCzNDHd4TQ
DS3koODHNLnAaSM72rhFOYTlHw6LS3/TS9nD8N8llFcGZ9+0VSwB+v8Kg9F31RDHJ40FBE1/06JT
LXYyDUeXoioZ4EpMqRariFpdo4EjtrBHIjfTlrzJ7arV+NLQFsxreo2Fb4JPkqP+/D8Z1BccA9GQ
5s8iBuZiZJz3avjk/6fHRdxRY9lNGhjI0h2/Rq2umyc7EaMmqFBUCP0sqngbzQywzE8dyfBrNhw2
Mxk9xKSmLvSqUvDdjW/esBsDVOPUBcn0kfQ7sU9fwdvVgVB9Wyq1MkMwDrZg6xqTuVUZHzm7Nmkd
PcLEDIfVR2kiiaF51UaV9KKkNfMlUDbxnb4Nf3iIOgOwoPISskCtv/AdrEvzLu8dyERs8+fMbdj+
zOI85msHk6FP1DBgaiiKTrnKVEqec5B+8bDOsnN3xoJJiq6pTONOzX84L8ksg/zrYhvsJD4osbQH
/rHiBVchhD8OOIoBu56Eh8jpxSpmYiiWtt787QXJFJkT7GB2IzvLR0kFYm+ZU/naM7bEjOmtw8BU
2k5vo2yldm1jXTdW2kefVTgvJcWCh8Dk9btXbGBYX9S6i8ZdNKGCkqH4R1R/LtAAyPchdmC35r81
LnjYgIhQcAnrS8XklvAco8M135kw4ZFBqpMZLdtWfb979+kjZfjravB1xqDna6NNKM89f5zdd44L
gW8lYdInJWXV6q70/du5SxBQ5z1wNuwTDeX0B340yj6rMb5g6igwz8Lr12mb81OMluoaDbm8kcAf
VUDQeoyQqXFGpXJ9xfeskyV8TYPOpMSEM5qlfPtwjnckmnebW2vtU7I9EEHYRix80oMnBSbMKhuI
VnK4jYZtrcD2w9e50Ut9EXLKXvCA//hB+ZZbUZpjiM5T0YDV62rlPIhfaZidbIVlpOf5adWpzLk+
27KUHYCKcZPAA9e4oMt8THFYkco3O0mftCGn8LJspdAQN3GCfd4WIwR3DqT/JR6xyC8+jXh+ALrG
42itud/4b6iz1vV5NwVC+wJmVa4/NGOYLsqrWDnHQdVgofAmgbX/xx19zVZozL42LFQXFYEwu3PW
Ol4u8+7hKovUXzQNHE4m2JlLeINi4rj1sE0PDh4t4Q+HJSKdur1FCe1OUrfX+U+u9QsuVvQa1LgP
bVNYusnBzPOgUA4qthNANtK1AYzUrPjQge04QJm2ttTHxm6dfIqT8hsMOwaZtnn/rE1b8CFCYX3N
lgP7krI0Yb0eGCF5mpna4BGiWkJzdsOeAccdt/Mdcw/GVb0HdM5vpicai2ereigF0Se2uV0yEfWa
BZ3Kk2uTdDjeQiRsYL+HSqy1VkqhsnPRMdV8cCIVXpaTfvl0LbhSHlpHsGQtO4yH/c+ucBV617C2
2Ed+9obXYuUwP+sDJO14aymANfy+29N+Sj4yhHcuLywJdmgPgvknftLelVQQnibN3lMG30ZTa5Z4
4cHyvioSMzXtbVJu0uAwMpxlxYwKqYbkT5ZZOp/5nk3SvSMM0nQdYDhXNn+DnO6y3jy6uPvoMqCC
bQkDY1K+Ol/m9YPtUcSkJDQYgMNSWQ9BuaQAzyaj97xeJRob+HnUk1fdaUYlHaySCZak2Acj083s
G2DDw/BJ0sm9jAwPwfHiaNAfdLe0F5mjPR2bb/WB8vpjIfgvlGrZajE+tkrjfsa/ENTP/uDCKWgr
YMHBbPZ1rEYLp/T0IbWkoZwksQ0AZcRFPn2evq9NhQNkf1raoeFlYweC6UQQDfnfUY6cpy8G4njs
Z3c+QcaZaGhtT+OT5j9Uzy/Am37O7oj5d4M3qfHMXt5KjrCiTZQ+shHRsbS4WlpASg4il+qgTYOM
/suD3qbJ7oG4E8W+lFVVdRgpQz2xJMPMokHrV7JfqawCBRnr6ckPaUQghMD3wkfRFenTUDbuX/0C
Cmbbc5F6zOtsvoNuL3ZHpc3nDvwWVEZ7OSnjwUrvGtfZUc47Lf/6qVPUtA4AeiAPlUhseoClTVgT
Zc6nEFCQIC4E1o5T0hhDhCGqZOsBJgzAx/CULovEiiSOt5T8OXX4y8LPcUvpg5vhz9LmlUp4/CO/
x6CXmyQ79swmRi3OCzbSoGB/ngvpBl5wiW1VkFctphrxEXQOBKUr75zT6qJ/SeZEzpD/Z5+5+Snl
Tv4iE+l3V7XlKJcWbwTp9ycM8QEKUJNfr256F7wmJZ+CPyw9RTTXxiaYpfp65PGBfNnm8aAzjXBW
gWQhehaM6sDVwPsYa2TFcGPfkSn3UHJDQzEsuioKL/xndHpa6S9QPDy/EBqlamo16WQj/qIUBObu
TrOPojaw3FBc8c29b2/305ewAEsFDGJ8n3oQF1EGnBprSR7X7gGpb2tcDpOcrKKRtPHqZrNRJ0Ss
28bKXfIZd2d3PiOoqmJdTnOIYa6GHg1jW88/HD9kFssOrc196Zngpg7yNQiIZqJxJ8oqNGEBa6EH
E2Vfpg+qHQUUdv1h6s6ckAE29+33JhXxcREIDStPzHMMiJir48E3DkLIOKLsnFD9tDcuqss4KK5X
xa2d9ZGMs+6g04F8gXfxvAylHxtNsZdJHoxbcziWmFXVHa5FZcPMpP5WV961BCMMPP3OsGPF8mFx
BPynCYBs9WCpBKzt8tdgUODBxv79CeKAQSywme50cEjVy1CNgUqUXMqGhlIQgRdzXF/6kZlve1Bb
nRR2aZiX3XVb9Wx2NoQ51lC0dgI8j7lSLASSHKx1keSWLA192EnaDm+xh99y5Y9pgedcRZZODBqc
gSZ/AYBfJbVeK8wEedT4Upc4SsppdpiHX7nZ36HYvB5UHKX0TAQ/+KdsqIQ5T/5l5FoOeszy+3r3
aEfzmCnFjv5QgrDUoeQnJZ+VK7saJ21kGY0bVoR+dA0Esuw9Fs1m30U+4pjd7RiiHV+5Zg6cjooz
c3rHkdlGXLVpwD+wR5XHpsBUyS8kMwOiucg8Go3MIxiDP96JsGX7NvJc2BarR28r5C8+pmhFbsSL
PC/BzCykYfPToT6vkh2n13DopM57/WPp8kIk0//M560Mni8Ce+dJVvgFuIPWK1qhLqlHe6b20q56
5hkSE+pPFt6zxQ4/uqQe1Wc5Wa4IHNpw4i2qjU+N3J26mVONxUiNruNJM8no2e/CmjKk2iinp8Kn
o8d07mmLmLbKdDCpU7li8aSQW+F2GYQP3l4dhU84PVarOJIdOaRtwlfMGrukTLFs/o/1QZekUpEZ
43jtQ6fJ8eT4qJ2eEtZQIDvdHv3OLu/mbe2/k9YIy264DlHPRdy5k/XE3aoqN7Xg5IN+YJhyA7i5
qRne9sxJg5cciQoJ3jHSrQb7IpbjuWs0XwAAkLgvLA/T42thbUCBr4LurX4o+E4HNyY8px6ZWvvl
qOHCkHcV04KqVAjRCB5JYgVAmSClZ5bvtowR1UzGQirmfLyiYWbuKJa1AC66YsNPG86hrAwzHqDI
jkdEkyvZKiLcuP3mny4LqoJq03az4Vbzcpyzrx68BzhNvd6FTcy6ruTgB6gskHayEo25LBccssiY
5iqWuQmXSc7R9lICyCgwDa8wcXAM4Bt6GAfiqxkqPNfS2PdFMqe0QTtDJkRZgIz+1f3m/TZCpg23
QRcDNluMzEL1EUVJVFhGMWEaM0PC5ZxLmmJdvRuehU1prQjiwQrLemQS9EH7evqweYp4lXPYwzl9
BEeS5RAtCIl0vsjkUyu43tViU0CWAk++Akcx9FlW7aZTCkAbhltDhsMgnBbVnmMQeJUZ4/1V0YTl
rFfgmCg6qq6tKKeWVB5U4cIMdMJeiOCVW35G7RPWkNpcj3uAup8opJLeQkpWJO6UmQvP17UxBJq8
yYxY/A8S03OSybUWuTzCBwGcu/Awrod2xett7Wgz3ie5nb8ACSJG6JuDeBTnRYQ07TSd0mxIT6zC
o6SPAeMiFp4UI4GxMhGs0RXd30qvBb0V1rvlrsQKgRsVs1p0Ajpz3TnxOOq6+oyITgHblYAt17N8
8O+NETYXNCvmlXQEWjL2jTxb0B1oX9AmAdo9QD18FpqfceLB434uM5cFp2fqhG8TUnQn4zDXvezx
KL9qk7WKGFApHWu+7kdPdZG58yQzxUmpSh5Jf8mB76jm79gV/XTGJBR9pArUKXAmbacJxCiOf1oW
aCAyw++Mw9J72m0vDP66rJasEvCD2dlXAqZirdAYQyc0tocQrXdsDbBNPaZh4MJcvj6vEhIXKvo2
nHrNZTH2SimuYhRUZDuAuoU+1qCzuRqb/+4H3/8oh47kNPmUAtUl9sjlV0IAC7rK3U97XlLWpmpY
szfuTcEqKP2T/9KtWxnm7INzcpuxmP8gBVPcsYZ/6ZEnfEQbDxFKbONRevOsebIToQs6f4o+ekYI
YBXX9otqcB1MeBez2NmkLit12zjptusecMlYkasvEG7YA5ZteNlAsyTqW84/VTQxb2R+Rn3gyiaV
h5tzCMQKEpLQzK3NQvh2mhw5qmm6T7gqozU9gMjfiF46Hp/aYGVjKoklAaTvSHA59I45jKSC8TRz
ymzLeFYZ9UisLk49J/IzO78kJDZS4Nu2iAo1KKHRUvfqPcMt5ZIVNhjhwIDTfLo94r2WpXDxrSSm
7PqGliSEClz6tJ0Pax+49eLbM1D53VL4ypDn7dydPT1cG8FLevN3J6+sE92T9jM4PAmlSnqVROOO
k0OoW0xY5+XmmScEXGpUd0JIWuLapZvMswSO7blWy1BZD6P33k2qOfqP33somK8YLjQRCY9g+a54
34fkurPxxMxf2Dd4Zt4/TnJFqQVTHxHOApOZX6KJJANx+uINQ2jJS1xhZyW3CCnKTMyWC15iv3Tm
/AtrQp7EM64ThkNy6knwFsT/G9+SSbpaNPGtvtLg1I4T+Sr/MwLaA7FHIaoS59AudZkbMXyODukF
Sflm85Hxwm4ILzQfmtLZ7uVPzcGF6nkuCcKRlXQGEe6eo9IGz3aEUtI5YNQQcikVF001rHEUaHc3
1GpdLP6KXCXsyJ7NH22DPoNlCrbng2VIdxRykcO9bY6nUdgY7vrDZb2eCOxKx4GHLXI/gUgxIzMt
8cnsaBjIzFOSkwEtcBPPMCfvbx/OB6hypQxSIJbVPVaDpPUMH+e99DpnNFc8gg1t8BRR8575ZXi9
zYgyjNj/MbmT3pBe3UyzXwhOwfaFJFDNm0Uq9SdPdrVwJoQJL5uYlxfAdWO/pgk3ppUL8bp6Iadj
+0ZHTqPaV0uax0Iq5M3n6z4YZ0xus+2N/MqF14LgoTuPs2rQOyaNivA7PU/aei6gSwHa+UgzpRjV
sa+LZpEj59DmJLSTteuuY/6yckiMA5h/mxnUei0/J/Vx8SGOOASU1zGNc4jWA3jIqblH2WUuIGBU
gtYcxe4ytRQ/bMFejmpYwAEL0/yNEpHAAGOpbaG7/z4snInpPOxyb12He0wH0rdbxlExGtt28+p3
B15/VVwlf3DCCVZXnspxNKmEpGKQiotEoEyY9eZ/DCxncc15iCsAgE9m882ntfXHr513zRPcnLCl
PTV5E/K446Dht28uOvkRmAdpn1Dn8SKPe6RtkfICA/xXFNAjX8eSXy+JDUEv+s25V/q/PIJ7cC6o
ABTzuzsdUPXNrPsG8JmyoEb+gn+AkkGT6DdkTWk1N7vTcLL9pUnSD1UNOkHxLmTH1YEEHpCJdQio
T9Ks9iImWGyMlSoLFJ1hlg9ZEuK3Wjg3/ujzh2qVcX/PWTL0KLiHuD7pXC4cJZq+Rmne6K8NB0FC
PohV7DG7C+hmjwLxvcZuIpuzrzo9l8md+/XNt9Ro73kYMt6/YXRFaV2c9GDheBQynTbRxcHqjfdJ
dN6nGlTEleyphUQXZNmEPtnehsxej5qRamMgzs1yI/0ZOvXX2E8N4EiUkMk/8S/ZLcZ18joRcErY
Su7O8z7zawrBMOp/APPmoIXLULm9XpYw7EUIsElqHuXhYrFqpYoXfeLaLbLgQ6AEsHawmT4jAf8M
e0gt+y0qbfhuoBdQD9r25XQqpLcNgPK33lZlbbvMePZqq50YhqF8ofJDLixnCoq/P5GwkxfiZZQd
bTqOpEqL7dfcwtjHbCoWWSIZi4Yv850f9Z4NrKH3ffGdNQweV6X0mxVZ274se33uwht9PwwuE05g
yJ+n8aab1yE5Rci0Z2G9etJU12RLqZ+ihqyyHdok3u3J0ighIfqamWDczFf0mqfi5EEbb4eNWfN+
FhJNH+swfPBMxMuQz7LgDHw3NHUqiIEY/6RLlHckmYGd0EGudhu2uM0d/3KeHXPgFGasSJo9zQ7e
Y6qofDWkXLhj1pwR2iz3mr74tpZ0x9RWp7kmK6MDElwOYtrS0gCF5Zw/3uoNKqsN6GDE/uewo2J1
0yReZbmc/+cK6jOqL49GwIeTPXws7wqng/AgsfOSIveL1dtt2pY2Xbvs+r7xPPB2IwS7ownZZ2Q3
f+urnZLZI8LV04q9NBZUmLLKTrYG4RCl8Qoqq/08VUUfhkEVpnKY5q4VB1oO2s9Srm+GJZr9bTr1
Kzg5G8vtIi3fBDA6mdpD2oPr8mdYNZAFOmkO5b6bjtMQyn0QTBP4xAYPMATeJ1DGyrXcLJiDkP46
77hZWYhTmFaB3AQ12WOqpYRBvmK78dJcx78/VeQJo3WuxmpZ63FQOJR6u7IJiI5/DWixSpn2r9zK
t3v9D5GwAFDZMwed1ksHVmdPHts8Kvix7GmH56N6oDWvfc76v5O5YadGyVfw0muMhWy1qzYnAEWV
YkICurINOdvme75/uDzluukdMlP1Z/zsTr6s3OeQ4c+eb+G7us8IcfZAQYI819F6uw3THgk1wsal
vG+G+miipdve/lWOp4ejhxuyYj/ZlUcjI1faScU3GYwhmKUfh33v8HpMOCPs8ZckNSHkWjvYZQXw
Rhe30ELCKGIvJEXXBPxmzmPRGe/eQhlIfdCf2Mol+maOe4LZ+6CrBURRlYeSx4CiWJPCPL0tKWDH
4EvDE1lvSGtwVzJunsZ5DIC08MtQOkfTWfSVN5YltQ3kDWqP/6Nc5v5CTxtEAoO2qrsdRck4r4Uy
TUPn9pwBynj/YLZnUrEPSDdWI0bYrUvBaObn+WEw1evbmpURbpSbK0tMk/KJfNepKxfrq49/gG1s
ffSMtWe/fkr4yxlaElBEEngWpN5F3OwjyaW+zlKvf/NOr/EKlijwU80oXCeKQQ/k8AalMTo3qnzl
kxFF7Gljp7/hbXUBqu9S5JZ85Hq4x61Dp5O2cyAkhuirvkSHE4Oa1waNQ6n9lJ0aB5IeDiNRR0be
M2nDH3UAIWCI7ZzqGNG3JqTTXFVi9XK69m+uuUS/VaUeKKNcJ+371LUA9J4bCwbG/ekIgcGESzF7
1PGp5E6wWupQwTTeNsHlDhojuJJqYYjKmuWhLlglGU/9x832XaMPQv7vBKbD0Fw7iSSOK108Kyj0
3ooZVmtTh41SjrMFdGPIUFQvAdtFdeQsHMiB1amdIeFlKWXsVbSPv2s2sFFsk37No2tkkYyLlf8m
Lfp/B6jDeigusETO7L+As83VI+R8RqZY5MukOLyBOvIBgg4d6Qtn4WFAfgetG+65KNRxGdoyIqsN
ZXMYh/9RLB9CwVPEIdlmO9/3+XmtrNg2BT2yNAVFRYwEsZhi/18Px/QHA9RRdlNNOE4mIKbIrbeX
uMANv9rVtxmRj+qaWvEB+XnF1e4KPorXjluHG44014Zof1Y5eqn/ehLghjzfbhpPXemWYvMssg3p
2hy8nPuWZp/ZKzrPBdAsE4QFzGODBxgkfHjsMsOjfkMzBdZn0Rvc4OBV7T5FlhsF8bqeXzrFNpB0
sxgDnUVoOoeRxT0hWCiaU6pefLyDJx05nXTyJxZTNEHbs5PcLAHJg0PTCowucpqVx43HI4MfwO4F
bstoJUcTp5SK6ZHBFsHt4/L+aeU+NFqioaA6zhx/GTop7A5Dz4kqY6OT5puo/TQQEvhxJtVX3TVx
c5Xhyy9uLqBR/XwJEiShdZps/P0FBDPaTsOYPGEPV5WJhp1lzu0lt90vH/U00QesjOQpYBcNgWOk
ET4UUpYV7ZekNBr9JJFRUID+lz9VpRoxQuj0VoRIBJu4difpblKz+0Z5F49esxhK6Q+KbYDOrcWS
t27yVk+JKwgqOP27mEOyWfvhBeLCV+tTLcoqQpsspmW78KTGRWXfH0JOEAwSDjdAxG/FwOClFCCB
0hneBdrU5B5ruwHyfbCr2cEtscUO6948ys83QqLXaTysl5h1YNKlpK4AQuwfkGPT/sHRjwjfwW6v
mG5TS7NUOEyiQ0srmjLYuxq2QXRFv8lhXG9/4JMtylsplaHRC+ikI+8kB6CGgQs1dEqj7lEwmcxP
BBg/TmwY4bYoVIOX5sj00l9YQvBlIqOmFTto8Ycv39C7tEemn4k8QR/FyNqOnflbE7hZoGZb1ss/
kgfnVxn2ve8217YnrHruFl+/s2itK3jdbq4PZGCdelO1RPXu5/hgugOg2fAbbWJPk0/rXtpmSgCX
SwxMs0CVg0zDdR57Uqkng50+QeF3ss9RNPRhpqN8oai0uaBYeme7Uh5N+X9o4fKx99/gIsiKkEe2
oWK0CXxdGPh8hoQz/vTioih0FhbZx7W/P0GcAkCgUBQso2e3nKEKS50eOZbBn8xKe4iijALh5R3w
HUlmIXhwn5SoYXw2b4/xvF1Ty173RmID6Ozc2esVxpMAy4TN6rGkB3YkM0ppOJz5LDzBfq8BpqBO
SR2yQWCYw3N6YEdyxQBGMf+BlWD0Pwxo9ukSFdpGD8J0w+Y91cK9SySHcZ+VysCyoBPIIKhEpn9c
AcBkW0Rqso/7Z87YSeZZdL6KYiTG6rTj4hnw/9kd11xUlss79wPOBNcLxLBKH0ANShI51Swc13WW
eMqKIm0jh8cTRx64UpU7ai5PDzp59Tzqo6dgbLoO7bUdiwOtZxxhyTDMYn1+CZbK+4zYqoX//Cfa
FVms3gT4EVJSBXMtIEKXV3ctCGTuqClU0S93gMg61/n35SQh14qapdkGmdYsqnyIop3tt55IuBSO
4pgslJURWuHJFEQ2kOAvTjuDHC37b4EmRjSBLd8/WGMDrddOL/l2lfCi1KltSczNZkeqlyDQYi8z
XH3eUvArm1QL98QERSyTpHVLJGVkWyZJMPutHAoxxHPQ5Giv0xoCrGlNKaz8VHmB/wv+z+70AXhd
7ehE+qIqGA/BbS9VxbJPRh25ZHJvnBFTxp1Y7TGHO24LDtRGGrqArIdJ2BZjpJwSxRkc11Dzge0+
SyYYWDHkEnXMtBn+N1N5NhOfKZTWy5ucqfiy8mhP56Ov+suBi9cqvjMrnb1ILSZTwjOJRQNL1Edt
bXkH1Q0r6rn81M/GcLKWiXqn7R74tOFnV3o5ERmxJN8RJV8Ny2jQ1XG8E6i8UnaMURQaR6eVB8Vx
eLHpuHeC/sWFo9NfcR+xOKeVBpKmVLUfJEv0jNBlfbjj6cXixwnTFp5YWU/iHwXCXxQegwaOgNd1
Tci14GOKdlgGvVhu2bplUUMsxQEcs/qbAqBV1Pnx53AybyUa8oMqK9s4vaFSmvENABU/vDgY/dIi
u5eOoCsTwvXYkePfJvS3bmcJK+qgSSTn2/7dF21dA173WRvZ91eMwA2dSx6VDcpceUAvpysfP8Kq
Hb3xlKvsIBIgUTRQm2tg3osqRSvf1n86lH/GHYMm3JJZEqBojDLF3WZivmHs2kCjfWdLbnj/DIxY
e0mEErNDD84sC/Ijq/zVwg/+ctBm13KyXYQnpzY9HCVdz8krAVPY1b8vZREtb4w05rfKkKBQT0yi
84Nywk/FMJ39SecvqqApN16OuG5U79HOjo4YmEkZ9T9A75+4ihJ66+mqeU1dr5JYGYEAig+jrDKG
9O7bM6MEh7XRel47DI2eD/fbDfBF0EIamHGJXrY0wGQMKOKSQV8mZCRXdUAbX2MYXAI+IPUquA4P
T3tNP/ySiZSS93iXjYhX3hIkZfgMTQQ+56U4+PCj2Y+o7hPIShw4hRc0IYzZZzlagaBKt7fMKuAO
Sv4GUBtCX6U2PGK+3RdKExzdJ5QrKO4V0xONJL8VAcc92E1wPeL96B2B+t+XwmbJBbOEpEDXx1uq
Y8JLDHiF0KTVpEoLCI8CO1oxA3QvK3FIAeRvfbx4HbV8CLo/Knaojm84XywhlDE7Ay/LgvXvMJ98
a6yGjgZLK3/xpccqX8zeVbJXJVlnTQaUiDpKP8lRDvfbGOtWjZPVPNrMXGpkFwveT6Fetj3iH8Sb
7WtUQDIxzx6hir5PbSlR6Yy6cBKBwY5/hyFRZGsJ5bk2OXUgtM45pHCRQgiMVs8NBO6BKnGp7QlE
e4x4hKKjAKmfNIoBrqYkYPQodPI2wkqeIdUVGVMq1I/BP4bQ4So33fqPpdgQhQy1MRQ8DDxzrM/J
K3H7y7OcRKSknwzgYGtJXPzVS737cZNqIyZdK/WqhlbVh78GcK8dQRJQGO/XbhqguHeTDPmIxSxs
Kw/zw4t34vB7aJea9NyXVUc7nVyJB4duf9mCmoR09wMcG/5VbRvzwJs0adkyMg3GSmjvjXqbWYA1
DBnMNnHmNCErr1QYbzssvMIYgtwWpEcT5CLcdwAG7z7cU+B3XZ2+eCkF16viXz8TJ2MuDbA8RgtK
zuRZ7MYEI/NCWXnrpFRrA2TQ7mg+7WlPTlmb54hpP2uH1AOVef+2bZ/mIABX91SMHxYA/VK/mFdn
V4XyQzUbh+oV0pWddPwCZ1J760v+qbzHvkHhi+6pBELPgLQ29tbs76Llcwpk0ko1u5GTxC73rlgg
1iOf5Y4iuYSGWlUWcDHV0ZVb5qqV9chsqT0Jtu/Ri+n4BmrTAAq8RrAXlMNPYBFfdH5ZBQoxoBPc
bht6eDSMQ6DnSWE1c4j/8e/CPAv+cTg+RvDHMCbLvHZ82OSAy+GSIgumJcjUspa3Rdtxze16ozit
MKrjazngg3NI9XQGEl6hkaRi9K9SdPrChJ3q+DEnIOmRa9z02UqtJgUhbHhRZAVXJ922NqWRopOC
3cQJjfQTJYzhey7n9YWeX3PYI68nN6wiIj6OOhX5lo15br9UZfiAGhC8iwq/3FPTXbEg66As09A9
2bOopOOsNumuD07XLdF0tMk3zNBnbWOssHhRfeLoyytAzV+GHk0mQ4xi4Sh9LmTw7as3fjEMIjlW
reIzuyZpc2w0Slg+nRBvbNQLtn2PXvuULo1lMpDWQZyxVWmOcxxP83Q/4lL9V5BEEaWmUxfF5WeI
53cXt8LSZ+d8L7Yn5wyVHkZ7B+V2CcKuIOiZ0+G+XQ1iSYd5si0BV9mWYA9HjPC/n+L88WSfXL/9
+HvLh1tCalk8psVRwPE/VbhD9LJbvgAoWnG3yBj/ZsIRtlaQ6Xo60wVMnxj2yEJaSLbYDkRi8So7
XztAh/l+/tZupxJtGXk8rPvOs09HFx6dW3IHHQAPrwwOzGwEnZj0bvyMHvVIYanTeQtCpsXDR6AT
LAuEe1laQV08wC3AgJlPQ7cL2MzhkOnk5Dr97655k9uMzSitzh1BylHAnwok4ZuAzSvbC1DBoNLd
VSsZ1seXc4E8TD/7m/mXCpKvAlXlLVpmf0Xk5Ctj3BeTeuiA8Ir8qlP11Nqq/vhQ7C/pbmoBoM8I
SDvPAyZcXGcT4uyayKiEdZKzyQaJjFtlFY6DErQWqIHwKz3JUGWAXVpuXF3F4pU2ITDyB3Mvw0cs
jM+fiDFZHY56eF5y8cUMuTMXn64Xkk8i8OPMqAWvhFjt+oJWeWC8CRUJVS2hnNvK7oJbwDq6ielD
slXRpWwOcAFSsFRqEIe75lBKBlbxyfo14bbAbPKu67WVY+i0fcB4qmeSGfxns/m0NHRFB5vmYoZP
A5XXOb9Trj4PgCDAIfdwsBONJ5oNw+xKXeOvLiYISnr725mvROLblmQm0mpuaEgqwpGG2J/IRakt
mi5k1U5gyV3L4SG83JUPpRhTd7l+9uwvUHd1PBYrzYXnqO4s+cs4Ux+ZqlFJFIDvtWrH5uG/+YB2
fEhzklTPsNmq2JR5kI7+72dNP7C43qTEp371nNtZrAspHNnBnk8o4CpIgST3ZMST9eNMR0Zq8BTp
v++MNLetTy+Id8/gratUPhBT2CStyuYWcve8hFeMu1r3fxsU9S9EGbQOtM7ADH9mQc52jLSRmF+7
c1H6CGMmdtgcFfdN1/tQo898sS2KH3P6SIM8Ibku5XHQ6invhfEllzQd8GSpYeLtHJS278zLW1b8
0yf9wwMXmMmYWgj9i0j8rA3XxpGHHZvMQ0WsQE6TfcNz9x4T/KhlrBYnZOYCok9q6Y/g9oEDLKgD
xEbt0zeMujHRDmraXOgxpsiUtZpPHcEsNz5MJI4PG88PiBQ8FPCN5ivLhI8eOM0oxXHOAN+nQiw4
kWNwdRgOxmdauNHYKiIXtzau48t66SyS/X0ey4vUHnOfGr8uQsqxzGS+2jR2o74cNqKwcdepVmYv
XDRl78Qg52/VRAVppdaHcZ/OZ7uGORLygSW4C9UkTta62f8bJKTXSI8jBMjmGgMEBL/JX05E1ltY
F33zsarJy8vVczaKcbfzNScMkNgD85etNZtynaag+tBxfgl5G1MJc56QSWyKpGrxSHf0meSuEZLR
KZc7SEt1/kCaTUvKOQYXRGIjht1Oza3KDIThamEsU61KhXWrx/AiwW+zXWRT4KJbeEnnDLAek65/
oAbw1gdoNcl0fX8G5+Af/k1JXuwzf3T3sW0QfDaNSC2Ur1tpoRRd+ZqnYHEntriJpzcCkZsZuJhh
LiYzRrl4ySnUo6blKSv/wHP0M6iIxB5CIHDX4IRLZF4ixzI82a+qFNIK6W7p3jskAhgFknhjIR/P
LD7kPXhpl1lBB8YGwNkTbTlknt2u8EZBaA0wMcIIoNvNfytvnl9XtafgfAn5dHEPefrXeyQz1mAi
EdZ1uxGq8JvPISZpvOml83UkzJJLe/xFXxG1dxUc+tho9nOd7wvz+0gjBLgoTOLIsW5FCQVcjv0s
tCBzjJ17G95VK5sGrRUAWKXtIiVtFgtDlwXeLvXLK/7LUDAfXApOevQaZK1EFOdTwZAcp7PN4rGF
BrqzggVgZ+SfVupeBj8hctruzgUSMjH6gZszCJFiaLLSsfMfPsisbzkwl1+46M+uP9juZCqoRFyE
hMIW3mWYn+UKa3tJP+oQm5iXmpO+g0dntpJ28byD05eoUaQ6YxPe+4get7dqH5x/qx95P2zM2XKT
2ArmHV5Am1jEfngrWdxdAiaAnVBekkch2gTA4eYqcFqx9DzgHa/Y5E2YTnAG2MqN+7Y6EDLlhUc1
2VQHPlYtyyy0nhowAGXL6fqaiub8mMU2sV9x/b6ENgRUC5lsGjcIEE+Jc/GJSvKytgoLq9hO1z2k
qgeH6aTgw6/lvL3VVwv3HM2Xi0sA4dWCyQOkoPA3eziTXBv0A1rdfQf+lqQyhaeI/4aARZc47AIm
bFjbEm1r5bGghKhvF0fqLLsBGCK1gSZvGs+448RD/muiU7BJjc92mNUn1eP+uNeEj/ko3qwO3zAF
Fiq+d7y+Q1GdWpKpxhKzURBK8NtkzkwBbDbuVP6tGXjRFDCC0Lt7gcnP5MptEcpxNn9llLXnAaMn
nb42HIx+FKn0IWxn/XVtS+9PC3QrRuS+msu4+gWTfF3nf3cEhkRPnA5CWwB00oQig4KvUWsrPwWy
XD0W/Qi1E/5VTI//a+7HO+5ONsJCWmTPB5RZdpwlt+EWD95oHxPuJkhpgUEW1RT7m7pB6WtHjzzw
avVyrTUbA4F6rezsAFArPpHVO4jgbv3WDrq1UScHyXW5EmVj9CAEw7zVuYNwomhJLzlD3XkLIbez
B/5Pcza5qG8P6b30ejr8hPiw29Lelxe9oDfrkICjTVD35swRqL0Lb8qIW+731a9N92KLlv+VT+hc
5LmvFZZXNAYlwhv6aE/XyL77pcZ+v4fkaAPlPdFPAXhA/mkTAFfsEn9d9mu6Xl1U/OsTteTaEpTq
UzGamU3cz6H4/rhQ3M9MOo4GfSHMP9FAAhNOZ/dG9fpFII1zBf7cy9hjSt2W4u+BHqY5tRxlPJbx
cDm3WMoK2mB6x3R/lOm3ACY9JKpcJsRanwD35ksUsKQBFGhX/3cATEZyUpSFmU4pbVqeMYEX23uL
kb9d8ub1ebj0bl4O/txCl8FNda7lI9hCenGtb+/s3qMUCk8xwWvHYlQJHdxOunC//E78ODFqreFl
PD6Rnsmx39gyvRQdRlJdcZDZLnNshRjVk+KQTdrt/JwYd5g+cXSV6y/1uAGv24qTTVnwGNGd0GIb
pR9U314p94G6h12Gb2bq6tfqPRvuyUUF65C8yElCGVdeKMZCHAo44oRU9NOEqi9I+RJD5JFx7WCR
5zxnzVuC12ezwtfjfnKuMnolHhG5QJrc39OLmK7zyud/EeixKWIZ+6zUU5/O2orFYc3mmjvAZRIk
E343pJO/tuiotEqGpI4cKgXeBP8Lvq3moFagO9K3kTrTFAB2ciKA40RRc7raN9NSZWpaPlJJYpPL
ZTmd/TjzZVHyBgFBbTNIAeQpc56XFl7AoyuPwnFn7A+bXxpKTeCHmc+gb7jpcKE9+YID0qnTbXAr
AkIfy2AXlFAMbB5dPaw71ZOcL4oIH9nxuY1HKzbqWYtZ7hykPqQKOU1CqJVsuJ4nwCScPt7oK4AX
BzlpCQt3ksaxMQGiDbwYaohI7OEzOIoagfQylfhQZZiY+wO+wEpzeTuC++TZcwgJSDIv65ghzwaA
C7senAo2aB1Imc0uqDwr6figRpvL8BEgKVWOr1W7dZWmooLQrhaGNQjgkdIOXYrXj//IkkVjrk2d
PNMBnetcHeFqNBBYE+kLl4fMB3i2ZDgTRno2E63lL9Ll3U1DoYZzhuoxRBalrOCdSUV15cI4nR0G
PZQzffnTj04iN92wgkjcDGXSrdCrwdAwbuAJmoS7ui7JdoXTAlfd7NVNEJMRlFiZkwjn5wvnNcws
KWQNePhas+hQ6LQ9UBVU0fatvJIFLOgLCAxrJZlFJEYJkqaYXzA4jaGX1uGyBOxgk4iPuqlk58DD
cEdQGF5uS7KeYd3MK92+fdP6nPEr3JMESWpyeRRamQ/sVZbwrLVj7YJ95gDDSGKy/I+AD15eshbb
TtosYv/EgyIQDvTPx/J21f0SPRptfWSBtQgtmeqPbSpiggrnOiWz0x2t5Y9HpRUAUpvow3QNCRtq
3rsrzYjMFKfCY60k+tuiw2i8P+/KdGP5PVWUxj+5qR70EUdrFUA6AakcpNP8p2acx3DpM/VQfIjH
XMY38wDON1GAtclLTaAoINh39abbdtYJt94fT7Zu1ZMnGLOu1gpJ9o2uZ0i6BCCEj+F6a5OLpGoa
KD3mAqOLxmuQpXU+2rntSVV5YZZL4fO2po/CqbssSM1eCmtnYYk5pOMHnCCX2koL4Ysiou6rwSPx
shnv850Cr1orZqzTF1w8lFMaAO+h/sSOBqcDwzl4TsmoSqeofHhm/OpHiFa7AOVUgNokLvR+AlxW
Juc0vK4sXrgl+4fBjdk/xL+bjNIv0w5VVuJx57sHJXDZ8URANT9Rs0Q8ofo3yOzMHP25cbsaCifN
pToL48jR60GrB7fsZHN8TjE274X0OAiXd4JOMmHiIVpaT0bOd6aJ4D8yrjsPp8Zp89v805ay8syt
VL8XU7rbYKbR+DAobbICBCoF4fT0iQ8F3rAbwtZu2uvHWG8TO8EXUCOkvLZg6OcMpDHskVqbvrPe
ebWgwYxunEvasOlkUINw4E4GKzxpveMN3mig35w1Da8l+JSHu6aoTifeEffkDkMCMPd+yh6cmcmk
u6KCtP2zaS9MDoBoE4lw4EovOZQuiYczn/UoHc/nNCmQVutJsxTRX2e7ExkcNVQ+Am8H4nLmFgJp
cdn+tHOyNfkXv9Z13qsNYN34n92PdshQzDe4vGO+MCCtM7KtHjNTBi4yo22WX2kvNijkJ3CR2gtQ
xyHcTLUXmKZOE7qav/2eqO8rbNxLqa+bV0oQGtskUqNLMMqnX9lYrfwWWSKvHxWKSUB2z7S84wDq
ZeC0DJmdSED33nr4mGTCDTrE1dqRV7IWXjUSKQqmPTAKsdAZ8IInMEJ8trv/swe/343vyUdE0PR7
9tars79+efUKWvmVgRTgy5I9yc0leCEqMvk5yGbwvvB32AXriOsVMOuCmXqiEqR/S9SUZ1+4jiwn
z0GKk0hKPjIW6MBHmixlGmQ7cJxDJVoAy/MD+dl/U79eeTX6BqrKfWUV52PQnMWS+DBBuYzx+lyZ
tqpZJjmC8TvqKSG3NKGh2ZCY7kRIk4wGhp1KAfSY5hrGtiMfwFaQLPM9e0K9rPFL9cQPorUzrDoV
9DTVeV5/PhIhdiFPw+TDXb3X0YinBRpgJMoLewkhK67+5a/JCuXVPo9TCMw1ozJ+SUpedAOXlPEi
WjmGhko/4+QwXAu32hdF4IcpiKBfQrjlwxa15hH+wgZbcaPR0jA02BV/oNGLG8ElU7dbvYo40GHF
d1uOVZMSJuLlCzu6u+J/eX7fiQ6ShlMHBmX2FcvDTpsKDpx5FlVEvZaBlP/AgCm1JNJJT8vx/Nhk
zRDZZRcoghbIhAqKptqNQN7h1W8ZuATdI4tqIAWH5OJ5Ul4nzNIUGFd78JwWWUoY7nseD74nzvlN
aNt0kcL5qRonoiDeYl1RQgfmECyqXVZV+1do+UaJSP4hm73nx0Bi913x7LEhiSe+B5uINBNORc48
GBY4/uxxXE9/WTQBbglRtkQhKmsj/LP/92764MLW0f+MS+ndKzW+EA01Tlg6rsvb9ouauRGdTFKb
OA8zNWSMQdd9dckYUJfSXxSrjdR4b18H/NQaX7yec6tTKssZcdiXou3R1kpVS5ncr38gfGW8zwmN
5rmc75NWMZYj1bxKsM3YNhUD/8XW0jvNnJn8p6eeybDv8wcBOctGnp/uUZ972D1BQHZO3Ufcs0nA
hPrRZQ0mIvwlh7vvF9JIUTKSKoHhiq5+FOc5+c8d64hmvzBPuKniOMZNXcE5ExvUZnI9Y08mtx43
RL2D1Erprv1P8TtQlOWg+KZRhDWGO2al/hcptL7Ivdrc1JijtruH3vdzeZKgQ5PyM6aQyhNaRjrK
kWW7tbo+KFt6kvD1JxKh60sWu4aGjjKBe2Z0EsJN71wFJwdzjzTbo7Xt1GG1adpr/6F33OGCBXz9
V/s0UdRVvc8wWY79W54HXV7qlWKBUDlREnGmAFocU1Oq10GNJvd0kLR1wReKsK5SsdfE1Advjeg4
qnHeMQ/q4Ei9odEPevQ+SSF1OpE2F3r7bPbKnxPfZQl9FS4vfWhj43oSevKuHR9IBnpq7p3J4URH
vszGyUl7/yjyZTpo50vLxwZqeWy6KtwS+sR4oucKJFjiKiQyfhCAvGf+57lceQiJ2pCOdRnnFOch
FpD0K22K2RXJBRpFl89eNLjugj9aLOYs9JGQWoDntTT+BbYMiZF/b51r0J2OBXGgWFYWk1M9vZV7
JvZrzxksesep0A0wTIbuC1qIMt8+6fPfaFM7GYsiCLqtCsTe2jlaItm2R+RVtUK7dGFN4bK6sHiJ
r+0c5YLZsvyjskcLcDwMbgV7u+wkMVlG1YexEBA3fwS5jEUD3xXueoFxkNGWIZOZM8uXKbTCoGpS
uGFm/ToqL4GV0xa8oDkoglhPQyctVcJa+uBeP7HyWuPucmgBz3fi5VgEGM59bQ631O42VzoDzQ89
rhwrdY8zeyY2BOfuCer49CMG//Ued6fBLnKoG5iZOHw6Toy1VfR4BuGIiP0o+Ct7WIo0jeBa3TsD
3D2wBDBB/lR8uyqmIE81qUF1QzMC1chDG2MfDzThE6tkEDfoeOvnFFdME64JRz/CR/N77DWqo0my
+0Hk0hObrFycgsPUODSjz2fDBdMRL4qzNYg4DpaGMqrGWEa4RYc7se/sBw2qgQrRCtCYIpm2C1wE
J1nCGfPk359+dKYCBAY1tMJgdmUlvUSdmWs4ZE9X4l2CUHC5BEun5GnPwbi5YNnL/6nlhN0RlD4O
AnA4z+kHs5EtjsK+OZYWA8nHY1xwvOceAoaueMCdpazM9m1syr012SyNfckfZzJNHy5OvGqxBxoD
iPJGsGHlLjg1EkumRubY1WjW0nF7v4Y/1IvHnkmh5YgWbeZgV2a29IvFAoEYhvNn8KrK5ISpBCzA
YgX9S88THIUYx9FbSFcmscxND+J8WGXOHLNFtvVxxvoKhydUcFkzKpKO0rV8vjC3nvp3yUfO+yLI
0rbqgOGqxZOw8xAHu+d1n10JznMgMb6vYXGIMmBlE3fx8cWIhMTWup/3mIjQxskawSBVWHVlzKOB
mm1K3n2KttvFf4Vr88lxVIF0mP9PFs0mOdcO7cto1f8UQuUVxIbyVF0L73k/U4ev/ENJyx7Pnb5h
Nl8qTNgwqgBLYx/EDXEtSG9a6Y4QUMDLVbIKLX8vzu8I5R2IWoj6RkJM6O6b3UvA2B6uyjkOcbRx
ypSJBfGISNWyete5eRJKHaaWY2/BjilnuHpwnBt1LgNJ9MXoktOPonbm1w/AMiI7abuhMjDNcmK7
p7Br2qPMkS69kxt0QsLl/UsjuKvrAdHUin55iU+v1sz9Xw7ey7yVlDivLh5pkMFF8GSGPjIo47v6
xBdqAyJrY2GJkqAoQ161dbMPGHxVZprF6+zjcOlvLX17hkXyhqGLjw9oFLsQ/BEwqPqHaB1y3Gl3
RY6QpmTXTW4BglE9H3wR/HZ+8lbEsdYQ+j7VIY3wI9aOi5t7uBKMPLUyQqDOm79mojhCfYfq1K9o
pRv8how3SVSSDujNE4TRqb1D12SMHQ1ysEkiCZbtPnRw/WFKQf8cN+HYxqEIeTKv3+G455wsfOFe
NVxC4Bat6gUDyZW0yeBLx2pYUvkra8MXCdbURf/iilzZGRv1LUDXJpdso2imbJB8W50ziqpYBfQU
u7BToi8lBUPnlGNpVm6xmK85HMMNfEEDF5UHwrTwymhfxxebxSz8HYQIjNlUbpPJ9ubBddx6nfti
UhzoB1wVtaAdBVBbuG1rbVXMbqyIeYoQfLAWULqPMUvNuy7N3Ql5YG807fMft+yqZGpUl3FmNfTh
BAT6wK6qFyj9MuINJPAFoxFTqocFkVRm/0Yr46hgT7Cz1Uew2958UznktCgmMzH8ZhdfSEPUHcRs
box3S36lWaHAFE5nPkoCaXVeCJjMQq/rlfXo7ZzS57ra2f5Y8SPTNXUHNs5Fa+nAGrHSSOZ8eJSL
pZRLKxxP9XxUbi4YFMhpIWYrwbwXg7vEitigv0MFZOiJT18WfJnkjMVxvs5DwCJFd+HAb03fx1FA
J9IJX9AY9JuAbgLiIf6KFNolB46e/w/AG0sSHK0rPGPFXx+77EAFFJ2jFm+CN6XY1gW6U4C+4n+C
YbDJ9rYI+NTgzKN9EFljnfwFMaSAhPIaCxU7ckx31r0FORkDnULo7NThQPwFgwbStBZSE8hfVvH1
n22NdHNq2pZNRCBWa+7taC8ima6CmkqW3uNyfqi4H+/QbcSXkRZuY8Dy1tTKHavySk6RvbT05tuk
U144FIuhm9reS+0s+dpNqGtaEqKrTBfEj6zATtHMCRX6l0MW8o6gyGkci1eHl1vj+OwWcxbFCcid
ukjAWK9h+ZRRCHJJagnSz0yrIWp0BNUVDEsqi+RMEIrOPvR5MPn5JTTAY+5G4qcN3kRZuAaVY1Gc
iFLU/W1Divy9wKn7KRWEs+dRxLfshphZmiL6EK3MWYihktAjIGc4zxc6SxEDvgQn+MdTGbKyNbkJ
GOBeXCPn69HZvVutuKX0VPf1bK5GEp2YNGdZDDuyCjKvSEZiI1/sCvR4vSlxrgwNBBnc87RA5xXR
Hi0KY2PsP61xCL7hxD7XaNeEGhvqjTnKqvxxbU5CsIARCF8j6nsKr7eROhSPmFhffKGnuFrtvxOL
I99nyVRN2GPImWUTL9urgQ0lmtkEExCRS9O1AgYBQrjDAohtLUn6+JczO3VxIxj6LRdSIw4zjZJV
lf2bmPjYHGnL4V/NTcBaVMv1/MTGsTOyDrEVYMylR0vsZjbHdPBtpD2syyI7npmxzkXJQOIkZ+cf
TTHueQJBOwyj4rh1qUVUcM5sS0aVmxBkOhb5Bb+CujuLC2LM50vyW92izdj3wccyl+wrtXcFBSbI
OOPLKp/1uZgg++Jy7DCVl0OrWhPD6pG9FfbHKX7GdtkHnVvS+bM7XPZklwRix61Kx0BaDWyPRRYc
r5CkidB6KZnMLl+4Yb9Y+iQvTeds+J7UQY8opufYQJDKP/Wmaa/vCngbx1YEpNf/b0D4dIhwiVLC
la6RCjvxF/3keUZKYXmOSkNlXx4Q1R0Cw4AiqWKafd5/Xs67ALIUp6egpYSW991LsgblIUG1Pich
f2zgJotE++aJKGkHlfcs0kR057CyJDQP/UdlWZ2zaLzMsbI1N7P4vOQJ8VJyjPekgneunvBoDRyL
Qku5hL6IqG3VEl9aXnXsfHWL8pYgwAYvRXmXVszGsthUkjvNpN+x8LRNQn18yMvnaYo2OMMtri7K
ow73r1cvGBNGyBSEeQpCIZKBEwmEO5HZDBL8v+R9dPEHvf6nHbMzRtC6pPpD8RLCFPGUfLpH1va9
X7sY/ttEckQG6Vri8Eck+7zqKTUTWK/7CIS9abpWLml//SHOL3e8SQdQUUCYOvbFsOHh1iFMctq3
MSZdxrIZhDEkLg/viF7xcaN/bDzx9gMgUcM/rM01E4ZyxvTbWdPJ0/4skcd+bMp2dXXtqE2TFe+a
GWF6jO13pb0Wz7rz8P2hIJPnFeZ77MZj+rCZnRXPptb2qtMJ/zY315BVEHCSBSw45+8I+Bz8d7fK
tH4oOhNnpaCkNL9HjLqTY84s5gA0ABfW8t+rWIm+PBHLiiP+A+nxCWAsAOo1tDrAW8hNEidYhBUk
6UEW71K8l1ROl6+NWyzuZev58pwp6wM20jbwxfpamzsKKNfJmAnYCesLuC1j6TLfjuJIGjXbc7xe
F4ToE+oGN7vV0Ld81rdAkRV9UwqURIe/+wzpqPyyIEBD6CLNvHIWNPQVrtMF3/6QLeayhEfigClg
LoIU0zMPBNK4ojNuYPnpjtf+ZwQv+s+y2/1DcDlla8v/4J+5JG2IGMGSsRRu8NvomQD8acPzWBbF
3HaRPkmnb48h+mpVRcWnjvnqQnxaJVIrg98MYIDx3OxPt2SRqBVObhAlP646/745OC3S9YpfsmsJ
/KnEJ8CZkkmweJrvJ2X3TXRZlrzJkcDbnb/ABcWT86zwqO9+eotl2XxybE0UJP5Dikq6f1PA8MI+
TTXoBxSFvoLpRCS72GTaUJwX1A8UwAexUZMJVh6l9S+HQI8JnaM8ezAgfAJqWZSL/vELCx1OTslk
VeiSyJwqZ37c1tYxsg0R0GBkOMF7qAioIwM+PdwcWsRvCaVcF2BQvhpQaKSvQkIHZYH/RZMKrOOv
Nw5cnTdgh7joQPcbchGiaoI90yrU03KS3zW3y52XD0BWOdYwW10pt4jqYrQjqCIGA5+NNDPsSRiI
+cEblmvmdBstdowvxqsxpho5jaVxegzsmldIZdqqmqCW9+8fTy8oZJMXAZ53r+KNA/gSyjv5QyHH
xOsGrS+DHyZcoT3kx4urBeInqjKBrKzGPwnQ1xp+wgmK18ijmmZqk8XJS23VRzKhCfXQEjO3dlK1
90uArW0N+G7XGhgoBKao2Gv6miPT+DMBwihQ2/nC4+KJv3bdQBl38O6sn7qqbO1matqTeaYTtAle
52+2dny+1jK0rBwIopqwyac9Rri+wfaJ4q5xl1S6ewVckFZmzlst8mVPLm2o1hgPlDTM99fdn12P
4anMmfi6Y0CbsH0fsARo7GG9F5KGKNobC9MAG+rZ7+bK6csx+OWK5VFTbg/DhetvBYsrX+tP7NDq
3vt1kA4Dg6LlJsgV5blTITrZ3hyEkA5gz+SLU37ObfqRrseDYIRDbHWvxDrIdTOkjH8fB3kqj22q
RKidEIkyiHC9BQQbEFjCMq+ZUofTIn+I9nF1UkrtXssrmYgLbmTrh1U0LpNbscfuSkmUCzWumuJI
rfRfMcuLFQ+gUEMHNQ3OnUPqHZv5K9J2BCBVpzkp8N1XyJWhYKaQJHXpdhjjjVxgnsVwVPR5kPbX
+BMqEBSgKYnolzXZNdrdEbfO8h4HehGQLg3QeeOhj9EQlfa0Du1GZjBQln8BJMlANUTme1kV8dzJ
rT7L2ktiVhtFIzqrGMTrOU1K3/mK/Uh8PH2e1lhsY1war+Q2Zq2SHX1lNmOXR+eHFDCf4Rxult7M
PUk6EuNH/womGYLurgkdo8mz02KaEXFVBD8P5Y0AXgmx5PpVGkoBzKSOgyaV6WWQZ6ihqYCX0yQx
zdWSLONARb+23Dl7ULfBrTF+Fb3CWjDvxoUi3fFbkA6lypAX+RZX2OcPTTdHMEsEVVles8TUSlSg
xVpZRP0AFyZ+on23p4WK2/Iab48zXTlE/YXW+Tg5eRvf54aquNd3be9N9tmaQZy82miGDV7Srvvo
mfopdJRA7TovQYmwaOn4fmaAZa4hg7iMrKQ6T8VJL+Yvn4yn68jCcrByOuW8h+qmoCvuX2GN6VwJ
q/j4g1KMwl0a/cyJBfSsAompidld0cReAaTpbuzC9nZV6cLZEVIaZ4ufBuvJPSE+IsAZoNNMuXaR
Fa+Yd+98pe5B4POZ+HdRmuk3Jgq7I+pyugNv/9iJar7LZ5B0/IjIOB7e4e2oKuyYg2TSnw1aIzsa
Sp/cRnyJEtZ2Pb3DRADYb55zvaL0qw6yjFYZ5TuWUHPHZHozuFdLa0BGpuJ0ypUwy0ngGfxvzObI
HZ6rM8OixRSCtwfXc7g/5f0PohAVaIwFSKifaJqrHJq+4mvh3kh/NvVLNj8BbgHN5SNB9pwof6Cz
dUAsVxyJAmj852ok6HSRAztaQozYAuE+nRg2iZzxuQXoDRqy8z9s5EAD63AgS2YT5YGuwc/5GVeE
x354CYP0r+4xyJirusm7kH1gydvgvug0v/3JblhnTuBuMXg0fTAncNtfiHkypjbzANHFoz3Sa4KG
QozS74Q6evwOx/cxXG6bE3ib3LQQ8us9fw8fUQCghGhfkdqzLES4UQEKMush0m6bsxne8r8jFPm1
W6LIDjpHHePFEA8S2kFe0GQ+Pe2LBSmMwJ8mMqGFchNOdTs6cpygmA+foBSRw7hUyPBd/5iESTxz
xZ8nLcV4Hxkqif9Q8G8iTSXh7KncUZHykuca+UtlNU5La2p8/pQR26L7Q5dgpemC5KNcdaDDF7mM
kvhxXoD6kwMxLtl1ZB2G+YsgVlBh9rEJ8PfZZePYlgO4aAVuO3GuVVQEcO1EhIDH5vlA+UDMMdFH
GIvcIrs2afbqKFeofOGrIWb28JXhuSF5VprHrYRWfL3vTs6+gKk66YuJpay/Wb33zktj5ywGjUen
BUg1OIP0GfMsSZS+uU+VpzrO1fyD7lg5+Q6OxtQaGd0d/+wdQE7hmFrClXQuSZ5Hw+QOMBSFN5lV
YYDtuopq4JjUbhDiy+zM3bEwSS9NqkAHUaxKkVRMsjjO/6CujauUR5Rey7Q+bzfBd4iuTXkPB2Dr
WWvQ3yClMsb+SdMa650CGSZ+zF7322qUAlS2mafioK2IADkVOfRz2a5eTsHQFnKqDdrpEnsUv12j
7MIAo3inhCqT4wYCiS0kVU/BvriZigTlBMgn+S8OJYGCwHv8z8qlcS8J/+GyBUtx9+dKS1OPZrkq
Rgm7ylEi2MsPqMnlwn9pzfzbkCLxbDgsQTN6vhyEjeGdDSzg6h/vzelCF5XyQmH56971Vff7gkML
dntuFKjHJkuM3ngXsNW0S976grQuwyKeDdg2jDH70Rqy0pCHRvEkxP556GqkkztTzDHnNm7n9avP
zMBhfR645yt/l7cXucia1U4oYeiTwxmQ0vgR+kN7+Gt8Hurgz8ysLIruzz8DjHHoKfjm4jTYyI9I
X7zzTv51zsfTffC36bTUDh0WeLwgEsTAhdABg+qun7J4a+6JpBEzG9737Mjtbv24AJlBi3mXYdUC
X3vbZGDt/IbNEBD3mqOTqXRP+tsmOv7NTwUda6uU+Kq/Jwhri7WBUz+XZlX4fM6tpKdLVq/TXRbQ
F8PZ3ic+XK4ZDoQpl0EBYu/ZE4u19agHMPDpYvudgTDygVf7MtAUR8gR7UvitavOiVmP/us8rbaz
xmP3nHnN3MbPGGLITFilPbVzJUdKa13MEga8mxkamyoKxAwy01yUdzqDqJPe24M46syCfh/cBevt
N9E6kz6n8cuvh5rnaY2L2q15st7kdEhjdtpjHCK7YiPVcsI7bwi7Yh17iK2TVJ6Hv1xLy4sMJIB5
leNohqu99hMx7Ilv+G5VFHxriXZAJnWodmKUGrwNTJ+o5glFKL+LPzF4SBXiB4IByiCM3mzSeIXb
S6O7XNCDPyXFvMHBDr53F0dbR04/xqvx3mQbwH7Orj0LAuQHaaLBqi8V8G0c1kp5nnmr0fq+jxMR
//xLI32emL4YYch9pjDyMQN4rbKNv/+27h7zLjA/G7LoGzJo1uKG/77bTRRVtRfQP/42D+Fwr8+b
TSBhPDGFWiKqaLyEK3Q7O6dhIoRnxnuykNFzPogo7cSEmo8GHEJBTSbl9rDm/gdDS16oLwC/z5FZ
cUxgSC/7i6VzyEZavO7gUlHFmJ5rk0acLdp5m8/h1TkvVT4QclZ6m/Zkg5oT9IY5YbnmGiPj/aSm
9mk/fgnuPm71tCrcKSyw318fWFrOHQmbH+18fjBF89GXP4OGG7QkKx8u05iC37TNXiONf2L3DHrc
QA3f8pCGETNfOHN6u1fTNqXn91M3WCLqNwdEASTcovigQR8fipKEFjVmgmVrFK3oJfAmS7BADq/v
BrViKpQN6zV4Ves3i97U9ico9dJ6Rpteh2+5GAN10LFE3gBGupe2PJR7BUvpEnlpv7pW/JO9D+P7
KF4CcGDC5E8YlMJEX5l7hS+dCCHxAv3n63DaHmyMiH05xeZWI5WxHH4jS8RBxWNesWhqn42GVH5k
Om35p/vakFcLpcH7133NwE4IcU8rtJLpOp/uVFmr0HmzcDKRetaIYSIIZ6eMobDE62yXE2JuaOcz
TVnYDkNWA2SAMM6b1bKgGqSs5G8LrEL/XSGKW0Kj+tQjXNHV6z1/CpRWn3vSjeVqe/Ol8HSt87R/
S9+Qz1hEjnSRn8H3fGSxGGrsOJp0JhSjhG75+M/Qk/E8p9/K+id444lCCcnx2uoT89p9rBnT27+7
T+tSehG1Hh6UEB+dm6KOl7GXkF8ip7x1nOywVIl8uUTqeYaRrD0YoKkKUaopg8H7207oB/1BK9/0
+tB2BlwzTbE3iYB1+AD/mV7qAY0kNVTu7elB2ILdgj94qy8nHzBx7KzRTjWnDf9lfjv5osh6fGdn
O4Hm436p2OGXeqj03ONFZzIsL6e2scy5hITIlcv7cnfBPlH9YLV5QUt1jOnSlKnIk4VV7gFv5LYc
EJk3wQ7D/15iOqA7fl8pq6jWYhKIvCeGAfshymg0HEaZe45evRxlp3nSH4ywLTbwCcy3q/XcCc1i
7KJZUauNLaCbc0syVqKhanZUZ6wCz/U6ZctVYf1B3tSux5J+df3taExztJmNgbZk/A85kSddv8sm
I3/7x0JxiRBIDOU6iXPrjmPXyK44QN7VuNTx9NKO+dGd3rgtY7/VZaG4aq5Pf40UUwh1YBlHBL/O
+0lpW6koHNAynsrTOb9gqy7H0zp8wKq4KJYOBmlHOyGNwx54VO1UDlDaGG2Yb7zHdfSzYMOvrXqc
aDzwPYbrTSM0vfGsF8xMgMzUrqfkKZuEui4RH+u7cCBuO0rND6QEwio5pZdcys/A47lO6QNfQGNd
3ETMODo5jufYr/HDL8nvFutTbooulH51v3FpEifHsOHqLGUAjDLJhFmJ9ivDqIevjblN1QmyB3lP
V6kxi9jZJ3NOkZDbbD6dtq+d4WlEHpSKkX7ho9QPOHogFinfI/rlDXiytEBXY7/J7MHN5J6oL33F
GNpmHaRBhrfLcjwhXsTB2Tcyk80zf0etEv6s1uaJaMD/21LZRP6XcHWjLGSRSJ5DGXsQA7sbtVrM
LoijGXIUG1injAvZCXxxqgo7wG73zp0dz0D3336CPeOfPwRt5gfw+h2RtzJ3TwCJwZvdQe6NZpod
XZnRc4xXAjAb5WBzJUrzGCI/i/wnxez9QS7aXvnx8OKuhKoW5s/h+44h1wedxg3COi6+R+UYLQkH
RBXA7bUctsGT04IONduTnrpmJ7PQM5w1WfoTqUBuv8tg36SipYlC8Rah/iqapiFT3P1ZGMrh++gV
+sRhIrOOGjSlVMScDhTCz8GqPBisV7cSFfgbqB3SYiklW5DW0DjbcsLHyGVKalp1OHY6/y6KSitk
rHbcrq3KtZVHAe1hfNmD/rXApAXlcVO54Gz4UbZjgvaf0zWo9FfAFtmvZ2mx46MZu4B3CQ/7bNl1
XkMf14fi3tVCr40N/TikvF7CXUsaBT9fPlY51AJT2ZxwEk11nNfjxXPQ2BTGC7SrW3nys316duNe
5iCSJWzLIL7S8KkpK7aEoDqPkfhdcapPpZaHIV5KKoPqgTIgbcxcTs0VkcEhAibeSmgFgYDTV9jD
r7H9eR0EM/djOKyeO9jS08GzNulPvsGB3N8CH8Zmwp9+UKE2YevxciLW38sPKUiSu9MUx1wkQp7e
OOKl4oCnoueT/PQTrPW8hW36vy0GkkWvZK35cMBQ9paggOkc1v9FK/I1sVUEenPFIkqsRJcXIm6E
jLSiUiGTpK/1voVl8ArP8OttbP+7hi8At72RVETCn3NHL5kSoRMsiCoIEvU+4SwuZhPbmMsZuNOC
PjvaIIwuc6LI6qT5uQ8VQdK0U1oevWQHz1dFANjc6V6fGJPmGlyX6eQpEGrBnKI/9ygXEJho5Iqg
dfE+7/zs28jkguLJ9Vf98gnwEWWOHCs69MbcCjfQww9Az5Y54sQPx7E/xkI2TpSJ8RKVwtSE8SYJ
/HX9qd8z/jRYOPrbmDdBbtPlVl+iAuD6zc6cOtmv76dc4ja+BDebUUQwgFNCdJt6SMGdnndTQ9Jy
lkq7cKdjeA2aQOhGHvFr1O1WBFxOGApdI391L4b292lIlXeT5SNXzfo8JqpSGGsvdmkoMgjMcRvp
jWlaLmXDcZvgaeZJ/BtuHDbrrviLEWhsGfgrAauJRMAITuB/xavpEiWdmoEF4Lu2zQoQR4mIMCGS
mjgAIT0dkBvg3zuVwqveHt/ftshj7JnGfb+IWdtiaJy+0m3wwQyFI0guWHzeUmbs97MJrVTX1F3a
rm9jmLkTGpzEnnVn8hhBsfuj5djKMWdGdoZeZemy0suVFFQKpxS+8u4CmWG03ilBWaywRDJ+xrOy
yvMpQsXdDlTPtyRWYT5JZvPwGfMlhhcT+MWd/EQZwKFfF9Kb+gEBEgidb6LSuSHrh5R1uxaT6vDc
gV2IQZ5mio6c0jqNFNCJjOwE72l/VZnT9Ibl7aVp9Bdd3J2dCOdwWGbzcqG0NEu/SxMGPlPHple5
836aJgfDqs/00gJfHPxVa1NdbCxi6YNZHmYw8L2SFT2/E5ao496dkSX0SJcyO6IX4ONp8IizLiho
ROjobU/tHpwg2x+7UYl9t9sviI3HMhtL6JsVDnPVfMn7jyip6PlRSnt9e6UkdDmH3cW3YHdeNcOF
5LjXNsn4uHiwrShnMbmGKJvgLcZBCcaXjjHmGJtd0KGqxV7rvpMeNGcmHnEpopHdZ+/AWkyb4yfV
AVVY2oNQ8qEEp6FgnEAYn7vM1Vh1TzOMI3270SIeKRnIWA60grAg8H5mWZzam/j4BfD70PH1jZ4l
Q9t8dKqeDtfrW7XRSjfffPGBT1Wr8bf0lEm1gRkUPc6GCSrxgDBxFlarEtvddR+KFePdzYiXYtJQ
kALPWP/i86RH4uA3YzYc/0tm9axGDwWDhe47VW4JEL+5WNj0zSaYbRKrLgpkPGFTFgIsWo6K5eAm
WOPT1yKkFQ0O8zoxC54N21PkxqbM+cUEUm6IMT5kYUgxHMwX6YQ8EVHqsVoOEZ1EbRHKPylrl/Qz
dp/3W22rWVI88P4qlcbSmZhWgHH3VDH2WqSVvnb7jfgV7QPURsn/O65fhniNUR7HJqdA5UKwz2da
90DPReGjP1XXn4Oicsqpjz7BeRaRLzoODO1EyqkNPslvX7aSTqs/WsiWen7WnjJDOeEAt5OrzuX/
eSnQZ/IiLEIDrA66W1Dtay5tfOYfdECh7e6cRRznp6QrCeVC1D9kr1Y2Q1761oKGztOquBibWZy2
fJCUfbHITsRLCWg7GWMvSDz4YeB6Ua3/UCSyShPgEO66DqNCmuRpsBZEgaD+I1qzE1vJReewVVOM
RmaSNPiN7CjMiiZYgq0C+N4ETnn/bT40jkSAZ8S0NET0bBx4EBiKaUQUbpQOjq7pVx8KPPyEx9Rd
jHSGP1D3jF0SoF0byBHtGu9wNSa/vcP7xg1Y2s4olPL/xCD08sI99ChgvlBQNKchCTcV7JapXIQy
R7oB7zqIS4cB65UPRm4L/8Gl4dzwafOk1sd+GKWxzBg5EmVBPLHP7rsZ8tgOTJlyk/fskk8abYN+
dIJJgvKZkDAvhmHFaGQsj9n3Wuh+aK/VfwvtMdGH49ggvUjQR7JoO1L4CuZQA6QJ/G2XTCl2s8ia
riR92dSOxEWH8GryHpHDCB6NWLVQ7hvJhQ2vr6+jDmKB/4NbKtlziFBJ5w5Ec42susRS9MslPk7T
7L/b3hb5mHIGS61F3ivAUz8rKi9ehdI2RUxt+Ii4kzwZDLNL4XlLLQzle37eWMTeHFXCb3sRQ89l
ooHU3So0z/OAPDAyNVl551JAceG6e+xdPTYhQZ9U6JYTpRBjCFPTcyS/p5LX8smxaKxHkuwqVQii
n7fq/EIbhO1iy/Je4GA2Tbb1yE6aCWJs5Ma9u4THsjYm8XrPPbo94dWwrcNmOPZ4NixuDLzYqrty
YX/qy3RN5Z4ceywJ+ss7xoeDf7y/ugQfhEYCbMqtJSLrIauwri+NIlH3YqDTWvAFH6WlBj8/IE5y
hHWUX7hL75gegNt1BxPVUmmiM7nu+eM+ojvfl+aFClFy0hGanoCYsQuAoKt375/Tq55ITtuTvhps
mpVzkjQmOlttY7K7wKzqm6RcPXpVdeAFE7rJEaca57EwcTDDMm+JfTBn4eJbBK0bNnoo7nC9eEkP
jl7GMm5hJ1aajROSrGLtk5VZ84Fei7UOowdmeTFPrA8kBJOU3wQLGkHgyQ/46iMyP0sXxQCIxe3M
RjtuLpwWtB2K1P1pLq86H610yqp1R3PcNj7aOLxEyJSbVQ+FIoSaE+wRLMOYLYGsIEMZAmD2ijmO
fxF/X8ZsR319i2CdvMlzNp7qXvzbWkXwzcZ7lsF/cxoU84MjUxGap5phG8KGTwTY7KIpsHiTaPIi
4nihkEd29GayQMWj9FCkAs5qqnPtxHK5t+K8RGcprYalRlFzChtd9qppi3tPZV1N6+hKs1egZqyk
W2no/xyDhDubA8IRdGX8XBbZTek9xLTbZY0vWqFab7T9mBSNojyX2GgqQ2zhhAHvVSBqBDDO8nrt
VER3LIqel9n8u2iu+wYtNlzxV0JWZCC1Z6a2LkvMy0mx3Pq1cOBF+M2r76+3WhtCM5Fl6TAsAIvU
4oa9OH6Xy34oGBxRy59k9L/k8BZq+H5YSEq8y691ZfEtojto+kOXjT5IKo9s84s4U2cg52kgTFrg
XJFNlbd61DnnklHN4tkur8ddShJ/Hi5fKUaKHw2P4c0rRcMqemJatl/V8cKrA4riuDrIohQy+zZc
UPqb9touMzbntgyQwrYAV67N7lq8Knv5IO4F0t0Lh+M0Uor9dk32qMH0rLO11d65v4qVO50WyGs8
mv7Cy1ukvRfV0Kowxaw1vavOaFmawK4sYovYebF/fDip8u7kQcIVB0zTiOgHd1mM/prTZrnFt1r8
QOKbEiZwBcuEEeSv8MfpVGLteriIY3LeiZBEx9pqqQrMLFQLxXLGtdRYL8C6KHtJsmJG+LlP33p4
qzxxYDn+zUDMj4EXdmULWBz4y72b9JMbS+CWMD98Dqm0yEgAD3hsiEifIrIidLfydcdfpNiS42ZW
j/iMP04ktCoExOZBtZ0ynPpXH/f9mIIFK07C9mqOsfK4BvygnuNx30Uahbzoylye0+/gfwZP9MXQ
6Ro6InkZCUpha2YuDmDfLLry22Zp/IlshWHA/cnnsB0B6RcMA6C3IjzdnQ3OUPTC10WXQKYy8Fmi
AZb3TN0pCzn4HxFce/kEcd/0xKoGRSfZWIUI3RCci7DNDSUtvOvKw0i+OXL1TV8pkWfe+5Yy0fBq
1dKJhWus6akOjn+c/aKQxvbADs2zmFkmKtIQpwTEJw0vgqRRFsbf0fJSJS8mAiFt9R5r/nV81ctX
JvexjYg2bzbl5iZrT+BNIEOzmC3tYBqPdOlVc156XIg9/g3TP1hAG2M202aDXOkTQwRRQrHyOI9f
opxCbq4mWprKwSlSLCD0/BkSi2+1czhmqbR0h8LJm5kaMhgeVeGVunIkADFwb5x2O5w/m3phQpzN
HssU/qVnqMVX43pfYRtdUMgn1lzbPv+vy03Dogx1kyoy2YpGXbaia7qs7qdER/Byct5sw20XEG75
rCBCCWp/usqO/tiSIr6tvnovdfR51we2HMQeQd2MgIUUwU2fNo8ab6K/LALLrPmG8YQyFmcVJUWr
xhY+jwuwULSBcQ6re1XkfQio0kM8me7LaSP5d4fWlS2pP4TzJPM8x5XLvKkgMsHGrPv6ZsVXxpCw
QZDheBfxDmTmn8ht/h4EEUgHkaBOOoVnVuUO4479VHRMV4crXMfqWQ1zgG1cL7cWEE6XM2C/KUh5
+II2d2Q8aYMWpRJeGeNKNWkAKswW4IhB45RsKH3OZa9RW1wuaPm9Uu+ty0j9R8xweZA3uKtnDELe
Uy6YAtH7eHkWPYdRD1xGiCLIvPUuEyILZNhgQnQTYdKcsoE8I13Nsg11XOmstMIddzFSU2jfl6zD
gLalCrOO9DcKqQnEXGY9oJ8P1b+Lv194V+rXBJk3Hc1S/SMzfbsGCUqPUYPhfkKbZ/ZQGtazKSYP
wp9WcZSsMPcrdBnVL3dcTnbw1by3noNs9raxMfmrftAEysJFfwU5U7PIs5s0fRjfneIzQJlxV++H
YZySURXgI+S4sV0H6Df+W4FeK8+YKOH770LR2rzYKXK116S49mv6n2tD1nvesW1OJ68FB59unNgv
2T+Del1LgxPoTbyrbrkAFguaI8W5Am13VNDZG1hEtp/DTdR9OnrR2CzRAfrUQ1GIjz3ECxhGVrGU
0Ls4+/tEF2SqdjsVC+ovb/HpjY6aJX2DqRlZD3VIWw3XM8LLQcdvujN7/n9abQ/uJROUzyRU6I5T
Ca9kXaCwTn8p2ROWdaOPMIMxPHGqpLnPdFEBA5tJx4QpjEZ22n6zUTI1uX2cnoxo2++BIfsxwS1v
jWygryEJWPYe53kOCBYm5tBnN3yp3W37PA0FKw+6Tj5+Uzt7rdgav9I0iYLnBVWZJ2N2YuBk+EcR
VjrP396Y9VBLz6SZKcUKzAaADqoMRiSO0Llejec62yi5m8IfJui2qB784OGss23CeX6ZDlyxGcZb
nN5R6yNUdV6cpMUXAEHFeEBxUmPEFud7fHyMGfn4NjZ48EM9Pqhoek7EeOkYmEl1Q1RcTzc+iZeC
bR24QVK7unfOXOrYMGUmnr7CbcQTyg48ZmN158n0d2qbaywya/nxubyUdxzbRnZJAYpS0qcOv/NI
E9jdJMwv5EzPUkYi/PKcrgVsj4UeHJHm4Xdmlh2ZASGH2OwMf1Bk5/vas86CGzXamAOxaiSrrTEu
0fa3bIrJtKH4i67RMmw6s3rSuNbs4j2vkJfgcBc/RTByB/fEpqtXJln9mwKKXEkxfKd/TiLKKXIY
iR9lPVIODDXNGI7Z7DhKImshOZoRnRk2qytsKDNeqX2np2hziP9rFZg5Gj7T4CjVm98ns2QGJQ/K
kvJrQZpsReeRIFAo1YDskvZZaNfCguBVJXYmyByqH6qAVuGbxUuG+64rI5zJ63nxoyjU2dnEu2Z2
m5CwcZ6O1/IhF0jGnYZ8bhapeUJdJ4T999bkJKigeF48RbLox40sBiRloJfdVqYN8OHBvnL02GE6
mHQWwuJYBCG4aB5hBNeqlAwxEisjAwbab2ZVmXJOiOSOHNkBC+gnCFBeFopKEXtITglf0VsjTcvZ
xYpZskn4EG/b43o7uJymIoQb9ikPY2d+FW8DlRQI1WEwLQjJA01/L9kyaQaY+AEW35DYUMwv19fZ
8g/tDD+lCy6mBIqDE5nsM7gCyLXGbzjQZhN/TuRb5WCVayhuX525Dx/N2DuHffktU9nz5VwRHC/v
i1ICbW9PclT741YrmdUVm2yb9MCLYQ39LDtaOptyBuVRAlq7FcUPQhZx1h7V1TLV0fEDRiettgT+
WGNvKJ9+fLKn7qPvcPotsQgV87UoumXH+GY5Dgjrf7xnEh38L8YsiStylG4LDDBkd4WzeGf7+UGz
+clwotm9/mx5QIXcItUFHpk2iJlKL3EDA5ag13Y1HmaPmmJD1XECrifWx75+XgZTie5pWPaGx4n3
KX+Yj5Ssli1FrNzE+iovG6fAYHPThya+kW7Uojmw0uVZTPoSFyiIxBqPUaZmh0IeodcdBNSrBXU+
qUmY11zeozuoEkw6AB3IqJ68+3s6zvfwzh+ydZAPNrZtoh5rU4Nj7Qul4wCezv9IC5LdK+lbDJ7S
shn2GQ6vLwbH73JLk+AW7u1uQFdePkj2nUHj+jJpGiVXfhkfHret9jnMKCP0EwvXxJlsEmeVowgQ
ppZICuUJUvpkC2algEWRgEaW00MGkxBogpFbYr4BYuISbJe39X/klzQm/kWrOYMOpejU2gbX185F
1zTiCZH7aVSDyCl+W+BQVvsI2Cv/BWu3/SosAt5RnLhVW/1F4Qlk+HjAf5Q5pBwQZRUGJXGNQ+kn
U37uSz3UpiCopRBnihwcpOpbSBpXWepse3KNG5idfQTs8zt7bMhDIRWgCgR/zh90F+36hMRypDd/
xAPcRx5PKo4o6kNAa/yaQHebryMEqdjHl0T1n1z57Dbk7ArStFylaakG4xg5mGMDNHGxI5ti65RL
lbMiAmAe5gHBximUNX2HnPtWM6zEUvCOFoDu8TRfzgF1MtO3sEX7jDUIyBVRkZjXVyixAa387EMv
f7uInpKZp3v4xVlnbSWxeX/6gsQpHZPrCscod5vlNuiZ9C+UsX/GkuyOJvlVjX7umjp7FkewkJba
gNVq+MkvJZzh3BoT+O4+XdA7Rncfr+3LN2G1aHWLCKNvTWAZhcvA9JjTZTjfWo264srbfeLvt4+V
4Byc0QaFCuwT9WElBQpy8AAue/2BKTEq/aNVcDK1yQxMnimGU88suAjllwX0CfDoDytElwIx3d+M
ObCpShHsVrxlq1bmcjnLyogIMwFesVaO/J8OqvgL2TaTcz28Txi/QRA4yb6p63i94zB8c6QfdF4J
QO6mrOzZd/A2jeBeX2PwaCXZpDnN1n/4nt0sc1Lf8vZ5U3ujM0+g4YIvmD+UWql9MW0NezYUv1rq
Kvr0M7PsBcfrtOmG1fk/5QeLNgdNsS+NLcTZwtL8N9Tka7O1uazI0w7wBieHB5kbFs2QMMPNAtdq
PfniASOJF5GnVtsDO2KaymdEw52DdepizpTgS8X4PBSTPdkDRXiFWBdZLcJgScNHOzutVDJJp0sR
WXJGu2kURLUGqzZlIvg9DvChEDZKiBgID4P3Tz33Q7ExApI/7AqwMxbPkIQ9trbCFVJcFgT9fIIt
rujXv6QNF9F2pAnVdMzCKaBOmZYCkElYOG6rZs2vSIcf8jp5XNi1nMtUAThUAAuW3hR+QcGXLAAU
vsT8ktLfIOZpeDoQKqQgSMf+ZYvNMcG7BXnOOKPXDYtDIyL4Se24O1C2/1Y2Q49M2Dt0m/5mWVbN
a/AZiWtEyiCq0mAsJ0WU4Vim9bykQVh1pcMCBgv4junL45LCMYK6XC9i85X7optbqqAIGrYl1yLz
3HFZmVD6sqtN73P1VZ8LjqtmT8nRhod8us8gP9VVUPLOG5/pG8cJ0gp+SLuja7kkoHWJrt5mEonl
qnxgypWpOduk41/EBXZGRI2jA/mVXDZlhCAyoPcDtEjE/0bBWDxnQGsxKzoQSSbP5vwxDsYVJDtU
1ZzK0WLsD+mBtYVJmjD9zRIt8TO8UrGS9C+oJv6nbG+u/YqttJiwMPfZ+z9eu6becZ5q22E0y3dg
BQZeByp1mt9feBsjPTpQAHtuRNlaVQ4v3+IeLP9XZAyD+bhgeVpY+sS3/QnnAmboEStivf5tBY2G
TKYUctEMyyxouBw+lUlFwHBSU3nKHZ0QTAfefm8FooHOBvkALMgmVHrRZ2yd+CCd+HzgKPovxpvw
Y3HuEW+ijq+CQbgv024kKNLdn8wmitLkA0eWF2Rr20RU76Fh9o/Xwua5FeAczGPlA9jfMpc3HHmk
0ucJhWhT7byCkTfDBoanuwfjgulNF74YMxUn+gpHGZW9NsD5fEP/XP808n6Vv/iskJSA/EZuJWIs
yZTqrfYZ6IFIZSm2ugH6m5Vd26djE/AcYu0I0mArnWfGcs+Ib4e24tpS81u5hFHMqIe3WHWSHVvg
yKB/ouRUa1qIv5qZtu43QF5pvs/xmj2cakI0rMIyXb0ngzVe7ii2ZE5n9AsNQrfjUtQKL7Iz6Wga
PVQPcSu3DEfVcoSG6WAeEZpWqqRqQA44YID6KbA7Q+5IjYOE7FS3RuJLuoHsXCfOXKrHp4JuqQ0Q
c5Fp53mihcWfNv+IXHELmSbI7CwHYfLwaaRBCkzyPtOhUT+hS8cObeFYWViMr+3RQnZOiiWw21g9
Lii0irRWb4010//V8NeJIl3U6nHlDlaug46UOz6rjO4an615d/Ls4UloBBzFbIO1PK5RgmiEJTZg
92wvAuW5gxRccZzh2Y3QTGlDLe2Iw95J7YfmfYP/P7NUF4I90/lt/9di7yVk4BTvAHh49VUMbRR+
RI/LNbtXtUKxfLU4P5syYJPHIWOVsHdeUu5BGIaSgqet+cNTEjEIhSNg2NhEsHNLMSQOd98l7rMt
45eTB07PnuQlETV1tWiUtfonlhQ1PvYaJnkKgYtlqiSTYWS8U8DUo2j/0mqVotJrVhOnsuEfMhTy
imzMaPrw3+NpeoT8Spy65d84sTLB3FJZFAT1kAPtM3LwGtH+VEtq86RL0brPzerddcbyH8S4UKqw
rWxyVA7brUqa4UjecsfygLUTDCz/l5pk7a+gvulmRzvnltiNtmofQv+debiBCB5SyThYt5D5zxu4
mx3QxgUgFuqCRDq2gwR8f4G2kwedE+pmSoAr8yZ7YOm0LOQ4uSbvACJ/ghaYwz9RtUWSGvddNxSH
UEwMoquhm9hrpvDu4XNFhpQ6M1rK91GRtY4p5pyFsoSyNaZZPk5C9i//4WCmR2cxkJWrMmh8E7hY
eGgaxqMvYad8LCBTfwJFd91w6iFopCz2iaR+kZNqB4NaFq+JMEE9UYuOZMVuFrsXtWWeI368RLP7
M4KQXlNyVumRVz/Xkauy26Zsm0+v9V1xq1frzF2zTmpEM7rXH33/NXv4OyjeEOffu/M1H12mW3Ci
14AraoW6UX0RXCAL0xgycs3uhknn6pekkFJs3khvk3Uw4nShRYLxRvZM7hxMLtBl0dsmRnA2h1ii
SNXW+++sUBD+2rVWJDCkMZbFH4rGLSAlLkdB7igXlbmphUgjomFhnH+ozCqTBLLemcN1TrciXVSN
XWC/NxKJ34XHNlEiKalniA6BkgJLslWyF2ddzla85fNhWw3o6cLLUMAyjutQJOn6OqCOP1ocPPGT
xmhEZ78b1poXkDgyd0TbaiJFPQ3xScQjuVoaCWwcO2oQTS7GcPf8dGpwMwwkON7jumYscMY1goLd
9c5u1ZLNZxCnGexJN0ekeBXKhW39D9qfnP6AuXqWMVjS8EX70xUAkFUjeYlf0oUTBggyvEb1Kvhe
TVBwoHN0PEYy6T+/E1RutLAGaSZrC2TqICXG2Bq5tZqmkafRgrYbMiPVmYireAwhP53o7Q7cTWZ8
52ppAVs00/s1S4y1ZZNctV+0H0Qk1RiMDRe/qNx0kS/irvgCxz62tYHNRF4NVEwo0U5UHwGJtg59
OQPYi0zk+/KBC6qVcA4Bw4JOMGHL/dxLlwe5TcyHKESUXj0YJwN6cGSW06uz62/ELD5vUyPKxAx9
3T+dJZa05tluwLuiIFGEQcGj+00ALthTPSVHKkO6KWejxDcSCHo0RZPYBleLcraDbf9sboIBFfi7
9N35/PPquQl3D4QNf/fVbNAoVE9Ce7ipsclfYQdQ2agIShtseHgWl/xMMGLY0or/NVIsl+Dx0XGx
GXHVkQjvqYonE4lT1MQJC2dfaJCnnjNX4pqScrYOBzHbhlxZl+Wdo3D6i741PGTM3i1Hx6zNYTlf
voFyumNlxxLF6cvwY6rGk6xxTc81HbtCXbp2m0VyM2HbzPQ6nAHr1I2Lfe7zjt21Pmb1VtJjRlaC
KCud5R4ibKHqRSjE4ZcZ932Jow9o+I3EO32pOYgcPjJLORZEA+QxufOUY85Lfedo4ScMTBwCsBwv
zAofw822y2QF+C/T2s244x9dI6giNF6gKBdm4eZRX0eouGD0BNltTkrsRD3xJOYNailzyTJ0XjQw
Wa/Bzk2Ee1qA3beR2IRRaCpIXx3Chlm5lVXI9oOLRDCftAzS6xQbInarwwpZdK7WwrJZfpdigWRJ
RhJDl9AENUGq4zD3rHB/ovtKgyz4hlZKWVbiiLrI/O4EuE5YGt2J7m39OnFSNjIGLxZuzWqc+j71
lFwjBLtSEBfcplkuJsUmU0AXMOYUSBUrwLnUDGN7HiCVplz1ixVLz8Cr9KAVEOWUvkdSQc6lZeeS
SolJVetvJFWa7ycRlHaDuTaqFLD6bILu7JmexWvfBgIItz70mvJ+MstfIUSCPQj8V6tNNSOffyVo
efsFCuaNc6kmNDBRiyIbGein+CAR+5Xrrc0qQOoY9PnPCg89P3yz66/+WusacZAnu8xrfrD33UIa
idopf1NOYi2FFgghc0NTTp3iGNWuTuqXWDsclBSaVtT4VWTT3wbNMFn7UVKqSmEjUEHhyWoRZQCi
o+ecEu14nvwq8Fh0fgFqA5Q/PH+Y8QIKTt+aURph8KRm9Bdw7CbHhGcIMiU0cZVBuXcyhk3TTjx9
QpDersojhh1Qe6UpfiZ+GmQgOs+lmPJjD7Oa6sHuAE/+VuDE3nvAhTr6oSnbBw89w6rH4Tdzvatr
xjom2bemzoIQu3dEuOo0QtGlum3QiM9nXBeZnpUGdeqUAOWYsMI8FHUHJIOvSnvc5cN+WvMVRSJh
iN7p28kDSfaiRa+wpqTxTquYo47h+pv6wEFWRy2DL16MZpxegxIekoVPOm1MylceoY7ExCgfH0bn
VCO1C4/DdWnSlA7EXfK6VjCuDS2dGXGqW08+qiyn4pXRRNgwOlEyGl4jFj3LG/FecU8LXA6K9sy1
+Y6Fgo0y+TJTakUTNyYeYCGmI0qhO7axnRiLd7RWhvfAwbhvfxxvo0uTcFt91TdTBXRf2Ts/pZZy
nSSVgNVAthvrvaFZZhnaEWhkNVPq9DDcxQke7XD5kwrLfM/TXnELmEnbQ6jDGcUGjk+syVXA7b0Z
8YhxIfX1ID9F39LoQULUlCwGu9GiQsQPQ8O1uO+Y8ruyInV0XPz8bq/SobBJDu6MThXVppcpCO30
Fexsrb/+sKCMT5My2gRf0hllqemEaKfJZVDceieEzs64s1lpIOR8Np0QHmb+KZ8SgqfCGE0JiD2k
/noRKt6pTZj3NmHUy9Mek+V1C/xUz6I4bOhgK1Liz0TCC5eXlts63uLmhifQH7Q+M5TyzvQAHhJw
q6JsT1ezn/ODlhrO5z8TFGy8NKU1gMzV8/H9Hayqj4l85sYp2NmGeAOyhCELjP3/Yh28rfwgwLbm
SBRgovyeWaAVYlOAlPu0IlGiC7top0KnzQL6Vkqb2RKxQ6V8zsGFZAZ59FXeAuVMmetcNLWq05EG
aD0flr0+LIaQYYolObDmwPkbYhD12DI9/fzrQIOWKszSBSeHSTuvv366i9S9v4bjOg1ca0VwihKy
9TbSD1xWBEYdGFFoWtQxeClzWbAt05jpxtSiU3BllzZnpC3Gjlnh4yVpgXlXwsnZriu4XDqlz+eB
ZUcvTNsr2U9E5bIy+hsYrQpiO8HenbsjOy3tFxdT0MlWso+56NBBCtnk8OFtQjuKZf/sCQWOxUDB
6pxj6Mmnt88/WsmYPWqtcpGaRBCjtq3ivxr1URrmQchUX+/dU7WdbBRzU6YZH4y4VETzy9B4TIX4
0xnngkUZthuYIFMlXWsMFBsxW2KLcH1f3eJgzCOoBZ1Z2XgCdhH2Br2uEGjWh8QyF7EVJZf9lRj6
atdeW3y4wDQyhORPrpRQ8Gez+lVqnnytEE3bFKj1Y3IFI4Z7wuDJlGrlcg04iCFetq6yyoIrJqGM
rQqB4HKyUd4RzojpZXMSxXqQsr1rFhUni+2UcLkLG4P/YurTGx9F/VScPFNzueTtuzWhqe6qG97k
hZn98nHtbPm2QTnRypmoawnJxzlSppUrO2+w9Eoe0OyKL2E12ehaZoUr0gHH/tpUk6sZeE07EddF
cGy/WNr/ECDVOBi4tZCSFNrImY7oTAwJxNPKkXAnaltY5b6EZ8CYygBp6zbi/CZTNr+bWJQkGMla
AX0XmB9EwyByYtI2qcw915u68wCHjs0elzSPWu3kLfMCyCT5i8iJdfWY7F9UQfIbOxJLeM/EsaJR
/bgY+vJwhfkO7HlO9AyStkzwgPzoRh04jHFUGGXBPmozj0Lbd4JGH3cSFcUEyDUVQo5DvW7GT7N2
FW4NVFP25QiRD//KZakvADH7JBV22vRZejp7BvYLIeyTb50xWsARAoaTYM/vHo3uYM673Cue16Bq
8Ls8xk/r3hqzW0if2fb279RQ14716UyE7I1zqZEygGWshplwK/eWMx/rUOBLpDO94lf9eSSEg+n6
jOSXPm8UGLQA/mYPdyvZG0M4kwgLL/+Uncfl37/N7HYLw32ep89VYa88+A0jQ8YwpL/WTRD7obAn
p4436Qbasg1pcvpUiO15k/8zJXFTjZ6BHLF9klL/m7OZjALopiyvSr5YEONp2TY3YEzPRostHj4f
K05TJbezt8pDyEgzavKz9R7JskeqkBx7FplO5/dZTd8qxaJ6ekiO8ACtn2MfdTP+6nVC501uhLQ+
4DC6gZZ52Tv01sxmqVe1G6WQMvsYoo3Nu8gk98Gn9AC07FoTuK0cYkQ/HDffxmun+V1Y16dFUpeB
ZlNriWsmFVaIvqFpM36oUyMEVeHRQpLGSPRXtNZCpXn96nldunoB6LU28a8ho7Yrhyym2EIf32M1
IbQpke5w2ZESh0oMLj02coA015XRnXgY9OgtmnnTcSuOgBuCN/rnVrUS5xSo1QGQgaeoAF9e6Kxk
f/YhYfIeg4UZtC8EXOrUVA4zogAEkjsERIU+xlhDUtnZijE37MYb/E5wmlrC5EM5vBdij0VzceZJ
k2/wioN8JoczSxBLoQU82slu8fC0mUu/sMVJ9PaD0HWwYrCndG8qYMUlPUnmo6fRMb5x2b1pmstI
NtkcGnZ56FXU6AViygbg141upmV63xHyRwX7rdZ/sb+PZfyMsEYLmrIDb87J3o58fabKZdq3KPYh
c+Emiqv17rhY9QKKuV3gkE8VoH72PWqQiDJnf1qCCwOf2+ixOdI1NgVPtUCQNMjOmvqAlm/FVMRS
OcogcQFktCLst/EMhQ+D3RVqdOkunIaAYak9/bddOLwxz+tUngxiR3nK5gV3h3yanOjKP7wwMR8l
pEFj0RCbLSMXHx//xk9a1JlYivv+M3b0VUhzRaSoO41dpBhNaRDYU+AoEwJQdwZ/ptiUm8WxlXcH
rrvCfRG/AmDkFsicmjGOXyPb2JGw9NR3KWlURO0oHPNM0Oj36HgaK9bZsdN84wd4pytXGNjjhNnP
t9ir2zMmFwXEFQ6F1H+fYxkfP4MkXVh0lty4bKCDDd3nMvHVJ04X9izFK5Oz4c0ty1DrnaJ5JB7F
3lFH04Ft34dU/QMMkvCF1Kysvj22JyK3gem6KqYTXvYvnumYVkmV9ROJNn4aD6bVao7h9wz+kSC2
6O+glVeUxOa6wRMcOa9SV23bIc81OsnVUJjw6P5FkAZIcE87pub2LImw81KsISyZy0TM8NKKM3h3
VCCcaXiWj/UUG/FzW7oMERci0GGtORWhmCsCOLuXN0xgQVyYG4BUo8eC/3SWg+r9VTdORP+w3rx5
XJM2R/POTCuzHpTyMGMgbHyDtBhIlB2CWxZotIe7yhr+WXPZDCTX5N4138O8l2+DouGkPEKRgVz2
mTcz+fsEg/SwVV+1QapVnYoqA9jsqad3aOZQzvMQfuImCJeD/fxN7anPvgDoUoyGowNqrtlkIi9I
GgbWbkg5wIJv8eJnjP/xFRHkIVA8jgKgH409OrLmuGaeWyXuNHuBQXIQbjpcrk8OWAwulwT+oTnc
Ys5/nqrinTCZHErVTqgm8CBeV3CYstnMGwl+ih0fzfOCumSafbGwEgwjUkVUszwft1RnHBDNLfKj
BCzFERqwbiVAzAC9N9mfOGXA1nYHsGyzBR49lS2A8/DfwheJquuk+kwyoY+OCNX5xa+fbNyvWDjm
CKb+4C1ldZyGM5Yc/vhn+DCr3EzzfPiiFCa/zxzKj/7RGqJkzvYwo3h8HV8ODni0UIbbekGEDw2s
RShvZLxca6gwZ+hsYR4ELlqcen4k6CqzaQEEVEJgyt/T9CZFW7r6BcjjgzetaJtJJFtvc+zKjT0E
0/dzM/YyaaBU74mfPi5m2YVnFVuc99tDYWG+MRZliL0ZO0P3H5iQgQtD6s5BXYKIVGE70nNgjeHF
aCDY7nr3x0gdiiMtUCRfnq6pUITHHzkGk/ggOg4wtdJ+RqcMYRJ0JUifO0TCD0DRE5hgj4alGUAd
QnsAMIwhcjpf/n/lyrcK+gnXmEDF/l7gtFo+KoafgmnVby0wsurOPi87/GqgqriSwLlkDbJeCLhy
y0PnKotJ6dMVBe6DTg632KFBP+gES5GnrDtIFqeXpEc2Uw0okGLKFwVgmAKGLt7UN1JkaFS3JqYe
AZnqCgs9ukeaV8/1MKt8rAKGnz8l3B1Gmsi3u5hgig9DKyaccO4iisVmE/itRnE31Y7XR8cwltYO
p6caKCmGpbYQbtUwVRQbV1/K0MYWa3JrKvsn/HGwpuPdkLIwMay5l61R1NgL0+5wzk+T1DzymyfD
sXDga677HvkskkIWm4b7FOOIGCOMvKZ5YjcDNgxvlK/8HOB5iEbdOJ9O+TtFTIv7nQKfS0S4sB60
o6gJAd6jHXPPoxXdnYxv/x+wO/+B1E1WxHkyENyZ/RkEhYmkn3GgbNQXOpwpmxIbJQhhE5H5R9Ai
PE8wEDatFwuigcLCE04zvk34N+k7EL09/2X1VEKeAHyPhTbWcd0LLzrF3pVxW+ErLnCnHfqa8wYz
ALSZBSm5VpMCGc7aQpOoKCV60QBV5h0iAXB3Y66QCZbftDUl/qvSIFrtvucZVYDkoU7UiHKXzdid
XxTnP3Bbya4MCR10bxsTdOLlWP/dFZh9+WnkbcMjzKcgO5q7McjbnX6dtea0YIbjDhXybKVi7rHf
CGg9oKiEmHdH/nqpEVUpuDKRgFSWdetIYMC797GrUImmRyM6tqCpXWblYqvrOytg9J4sBd1v8sZJ
D2++fv8M95YFZNIvrcpbIbiRxxMEt5rb9MqlCTd3xmCTMQ8jTJdpxqE4dWsNFJLMDg/ZOUkNfwZs
SQzoVDC0tdnY/3FE9dVtZLFKJOo0SYyQiiXM62Js3sJu3OPNOjAWulndGCAipV2dSnEon2t/ETfO
5uCaUzLKfYpMKD5uoIxMovD+siSk5BR5h75zG1vPjaJWUnH/5ZbEh2QqFgVbdZ71wKOMicHv8mh8
N/DZyWQ7xvCwgRFeom4TtwFdrMumGUz5fbwECbF/FEQ0yFqCLuMmRn0LOsIoj3vWSBL6sE9TGgDA
B8xYYpk5ET5OL7JqvtXhLxNQX5UTFkqbAVpbpcAU0tUS/DIesqcb77cPrDYj6ZSXbDDbWeVEop3I
AW1R6j5XsYNlixpF2yqvZe3DK+WC7EBQJ0fsaN3BdIVOflaDGg/ILaQJxQZ9I4mP6OHTmahponWg
ClKMiGtRV4RYQT/ZL+F7oeW+7kCmEqFVmrQmiwANg0lWxmxN6J2DrtqRRo8/cMr6Pu5qR5UHh+eU
y1LDXhaIZw3TJ7raxrSBBZ8tq0Sriwmfq0TyxnCLJPvcUW0PL+CcqKua9cTmqNL6Xw4zMhPG+HLh
8Xy3bf5474nf6LL7nqzq3Ga8iy+z+GrQ9nmRiodmNojnabxJhv53cZWbrxvhXCt/ND3vJP7I0bbq
r9UBKVgID6ykOrJyMwdxskj0nQPpE02gQdSrMzQffnXz/Qedgy5BNzU+WEFufpTVKzwKkWhSeqaq
9GQ+tp8uvA+VwfnDPNrGIK0HNL4Z0CnRv6rszpMeQlI/feOYIGElCKyTcJA8ooTUBoLAdR31KL+I
mzLHuufx5ddjLPq6TyyfrLQpj1CZ+J9I8Kco/8LB60fz/rXzo9ayWl+bvpNwAiTwAJaaw37e+RPV
ruPIJWzUHFZEo6vrxs9H03BjZ/sMTSMYTf1GOl6ELRGGDUnJTCQjUWG1VaqDr41p6LPmXgAwrFi0
XWPBf7rsKmgYf/GWfeahyNOigiZ+a0I8xeARvf9ywsKxgDFSlJQhvTINZEG3E25dP5qmD0TCdWNp
LMAygtWomSKCWySWCYn6T3DvSwvbyy9padtlYB3u/8r5bmBHK6sFurMihmKRJc9SaBcv/eVwuwzR
Q0zKWAsKQ4M6f8YXE+nllEQpsCswkvlZkJ9T38OucajSw4ASJL50i+jPjLfPXWzhHKg7cfGXl3bo
4rYROvFS3l0toNHewIJVfaYLslUeZdLEIVZDfojSPXDpVgPiqyFqLRexp9jOfRw/E/NeE3/lcH4V
CAl88fsRLU+bnFEjNXkKBmOBzMLmPThpFlz7GHeP9vIWi9jJl+ynBZEV8VYBYsJuXb7yzXtdXSKV
D67JuOk/TZSJuh+UsNjsXEldMOIalQigfFLtGhLv2DeNi+sYP2pxDo2fK9uQPJCneoDhKjTDLGLz
JrnoCAhZJkxb1V+rmJjSH5EFD+Ey0c8UtLd5GHeghpVDr0xyDmp4dXPfMChcwfZPwCZx0riyyKIr
vjwrvjTOpNpiwlAHa/wL6vJw7jPK8NtyekIM+BWV3nhmKMMzMl9xV155YQFLKqiB9PTXjYX+Llad
g02MrJoU9vwnSU/32ywdGHKb2bNHg3g3H4Ht1POjKq18/M3hulaJQwZCTU2Oios5UvI4KNWFq9up
UKEsgy+WwhLvcXgAyTNY0e5rJi7frq68UwmBSbP/0w8g0ry0D6mDwramHxuGdeoqnXDgmkplaZUh
rb1CvAzDMlxGLUvm3JeSBk66+CITjqArDs7r8zC6gQ6hMFoZL0mGdApCmFBW0OjvP4rwKuJNtpnJ
RdSfFJewy6HH64oEzrqvgC89a7WQhCgAHTvFegDmHfMl3AzdxPi8pe4xR5Z0HNopzDUQcVVw+ivF
2xNJ2UMY3JVS4bevLXN/gLFrDrbZCRo0VEKP01m/VpWLx4vyprj3Q9S7s6/WOmeenYrNgVIASCiW
160uaSWDv0futZBsaucK5cjS8SWDBAlSq/O/yZJeWs2H9u/nWENjXfzAU1+bS4qdRo+xzigvQduR
9X31sW/woSbkpIGI28KpzD08fH8SKqBFKkATKr+WXhkNmP/a6CPro05LieJnQNUlaHE3Lk54M+4Q
48pEfTxL6FAgUbW/GG1ZgCUIeiHK47U3eiPtDgSqDh1dHAgVWsvUM8Kcp6Coj1EVz3MA+17hsrtE
LZ7MC5SDcfoPzoSkRjNwkHQnsE3qllKcB1LvY4jOP4PkpNPaMfQzO44+6IN3pZ0SlW3LVLD2Drz4
tYwLdeSCvuLRPkZKeo53Gil0Y7s7SClqgWh+CfKQacAcj+engtkukrFjahLY4ToqaxPpKOKtbDCm
hNFkXC8nyXq9MoBGD6jhXwoUCb0YYvrK2ooBlPgk1642z9MiZXxmTFK9DQUO9C6ByVjzWD+9mX6e
OXWIgTotsbrYQiGasSGRb/M2s3mqa379csUXQ7UNr85tWXYdckcfhNVdTULyZ/ycH+QGd+ih8Nh6
LBqED+tw9t+xsX0ncC9+e6nyYFiDWEwRzKwIvtT17AKm3Bl0wASgbkBN+ZWswPs0TLs1K1AGoETH
UNL7JoVIJt00XG4oRWIbRZ+qS8xNIgXoQ06fBOuFgpqvycrUXtAQsU7/WD2e9amtvOzU01m66XiR
Lt4x82G/tf8MnPgVdbskAL4BkS2zV1BducEF5g/1L7WgvDbGKY5kSNApcoqKSEI1I5IMn/WyOBJg
1teOulFvnhtiO+R+V73DTufRFE67s8/Nly/jgi8vQaVkKVdX061gJySIzhgIsnE7++3Jsur669OW
Wq2JbyhYj2OX48woDVRiRq8vW8PiHLkvRbSb3LUtnJdVxHCVJlIo4bNlSArB0oI1JQZY0YzonKNR
+ZgRaMg7jhJ2x9ou7vC4XzaWOLuRUy59ed8y6tJP03b7llYym4QYdxavDn0E3T+/y9B5tyTkOh+U
3c0ydBxlYkehNkfR9ZUZww9PCGtFCKfjj1xWA1zHm3kiFFdpYJKOpKn7DBX0xDP2Ib4b9+hyhd6R
HWa/zDpNYuIMDO+FXYIJk8BQhQEQdX1P0cLs3HMlJ9zWS8qwaZJ9cq4xPHY8aBy54Pp90X4wmHSl
91DfJacNE/FWyscvxCCOtZdTtK8vM2u+lArEiwpY4+KQVpOBMNn5oFe9T8FumYaYmKhTrNTK/Ub9
HzYZOA61uUxKlE2R0jLav9RsL+I98M9ZsaCi6hUHm1tulgSCpKRntaZD4KZdqSs4Emza4Zcqr5MA
kPqVYtgq0JIzdPEGlAcbTG+XHjpM42UXLRcOk9XKfIG0RCwGnRqPDHXw7TTFpiOR3dYXdaJVpjcC
5Lw4kcPQAGuPcRbmOkNvugBtcmF3vW02+v2+pEqHN0s6VoT4oZmDXK5Ivn05udOEjI1qdaKZpTVH
XPnbyW2ck8LhpL7ypmctsBme3WeSJ/HtdmxB7qQAXXUHeRvbS5l1nsUFq1HTqVy1Bh/bf75x+Fm7
UbS3VWqFpDFuTe1m0FmswTr73VTFLy0ZW3zWsc0oNj0UpWzNDcbhppQza0A1Rlr1UxMG5/uKNCDR
ovfkvt2fsEJ1ctdyQTyQxMjee8AUpGXzQKrdVRP3lTt5TRC7JYXP7M3/mX/SJ/J3Iw27mg1FhUQn
Digh/7hBSK4+R3udHBthEsqxIBGOSOWQ985flmTrTD2nRnNhuvGe27rLyo9L2Q6kQ2tcv0pVvEG3
iTz2O3Z51XWTSBVPGxczKPZHQifCccoqvN3n/v/x7f6BwRI43yNfC9xbK9fV+ZDL8flihUS8mBKf
SFkXV3rzB3YpUq3pM9WMbnxs7MfvxEaAJ9J64jMq9FOubwvyAXa8CsWC0QlLqUNU4adCr+gwp9te
qduiY00TMvJVY+2mo2eGMOBurPGnYnuK14LXwM/iouYDoMNlxY30BMQ1CsMI/8FskA667CN+bwQD
UBl1mecaXCS/MMJK//v7DnmBoB7qEC2mTZNHA6vEVj1mWLC1W6cbnz6xsOqSX+AwjIWDl55HfED3
vH01sItvGjkDxJXXLXscLFiqPVCNi/kC22+hlDksYM9FIgmCAdhCKg/PGJCePEdNuyaCTSaXjz/p
g5etqPhtFCHMHDMMh34Ju6BXyUampq282+olFYNOyot0J2dFRDVfN/2uPYWB9F0en1LFLhslEU39
RduyaS42HYAIWxQgL5/f7qnrBkVBr32pm8RW/57VjjpyUG0yCvTmBpz7ZCxcAJeWKQu+yG6VAFBV
LDCGYLH1pdb+IMuS4ON08oRt25ysJEVOu/Pm3ae1cBJ+G2z7VOXivQ1nmyUbhLlLbKz1Hwng2LB+
mQbhmSpa4tJ1//4B/X4KJuk8KIXRjRLqQxZmPBH6erTDkqSjr5ZmAEqo8dL2fHzaYhDxCaK0HVuJ
wurynht7+eQ5ric6PiaKbuyooerca8jp3crLu+6Spw35X18dGyHZ/nSy7PP24XqB/yYUuVgD/5Ku
vLyww3zmzuELAKMfVh5fuT4+L13CY97du9Evx9pLsEY6RA6em1IqRx8NJ42zWGxszxaVQWIwnMrw
OMOZHQbkD7t09KrCvsmlucCsMioZBU3La/srT7axrv7jNbouu002xW5A+YTlMsxBvPs1XTPdj+8v
N9aWdgrlNhDZ5zdVrJQ2kRZhmffvpMEsu6UJLbXiaW55rh9IrU1hWfgcX/7TPn0BG0cUy7oub0gG
x2fUkA/rl84vfpOzvuHymALdLzub9NvJubY78OybTrI/TNCqAaWUZ1OWPCX4sASLPClwVSAFAPss
6ivxNZDYPRMDjIPeK+S0JOtNQchYlpJOkOR5GE6YYF5zakbsbRFg8736R7rAQhvzrGsAbyxfnMbK
voK5tx07hpL86WEzc2WWIrJSV7spQMMPTLUaWxSQPZzrRL6Qry/6GwB3fmsh9UlczJUQ4r6LJ7pZ
UBCZrdvBPnf6lZyE5zpaUrD7n6JPmxQtRCp1CRvkH2hDvT2ailNkeGltEV6jIWW1DNrlJMeoFpOn
mb9ivQeU/Z2XSTFilTRqE3wuJ65fc3kcxC82/g14cjZpNhzMpEnzpbpy9ihbHlU6cpYKmn6qU/M0
fiz/w/BoCc3BHjsmInyH9+biBXyNH8d4l+116uFU8ywtl/ClGzbGDExWcyXBTx5JymKxH9vXox0r
El8sfF/D7YyIzyN980YqqBYhc5IvRoCaef+wrY66HwA5GDpzaFbSindeDFKv7wHRepbuW23nqRaA
mY+yD1O/K2KERieMBDRO74UMdVWjwa5yRJ1Sq/eNJSeBnaCS87/VgQQJPSTfT2lXszqfzUV1Z8KY
NHRT2PPMLUWMqXmSOwcFKGWQ3fCmapc7KbolTXfH5+8Cj2lbHhyxnRCXDnsGlVlsXApS7fliD9/Q
SB5qbdQdiSnTUP/xKdmvzn2J4b+U7vwGBqMNd7csNctXT28x9HRiNCNRjoh+DsYCjQimrOdQzKCA
19LR6ptL6/FCa+Xq31XabG/PpWNNyYsITkw7mcqMXY3KAirkcPAAMExG27n6RT/rarAUS2SQn1CJ
2VmDhboJ+HSLQDQvUXGbf+1NN85sp1Q9fXTz0w6Y7vHyfktmCR0GPH1SY20evzlOFkxKvN6gfBIR
iC2qqx35fcVLq/DX8PgrydnvWNyr7tnReujbOr95AQo4TSp1tHS6nlcHTnQOQsvY+xWdb5No/wU/
0/Ntn9dLBLbFMJuwOtIYrb28mWuMoOglAGWZmhASQ9UoPqaXd+OGqieQu9aPA75c6NBiFKtYv0In
gYvimk2PB2X+8//OPuhxw1hp+qfdXSyyJ8aL7xCA2rtn5McMDhOW09/WyHj1Talcc7aDZkzx9AIz
QQxu/weKxIoXtL6qSWZ/ehoFGM28OPfCAK1BRUxlNVQNsLjktl+BF8z2mBiuu/rT2pm747d1gB6b
QtG5dMxX1RmhqGGjDWQffuogxV+uRixZUt9/o3SwiwB+RhfoJya18swtBXlWwsugd/1ZJsim3JHG
Pb6I1DvUULqhoW+mdwNUdexJx7QBjl670agybla1IxbagkIsKGzBNf9eTJyeIgnGqVfEXxp+2Fwk
jQLaadqb5POwtGBnUFJGY/SsMrPJ/Oty22HIhi4LHDAh8iAEI6VLYVjTsm9GgFCNEXqp9TZUUSfc
yrjInKBNH3Bt52F20qkrtdp5kp6iGbCc1bM9lDXfD055tdkw2S/07pVodpPtu4cDcoq+X8kRasKm
NDwAnKNZ6I12nseerbES2FUudXDoWmqYwm8t61+S0Fin0UtU8NXEJivi++WBuBPpEK+sdnI2wskT
oHTN5+fysJgjFgsDFcBbXDCGG50HA3UTdYM2t5rcITexsLYdos87nKN7ZV+X0zI3zCl9z/bLgPgF
nY8yiSfZ7py7QU/9d2lkSKeIBb8qlCFC4PLUUcZzQNP/yzv0+GMeYhDPgAOzhvUdbV0hP0g2woHP
9PIsdZbhG0S9FoQogEOQJuVLLbNNfUcSo0sDiUQBjBSw6X9Y1ah3mbzFCOHPhOpoB3A19M/9ZJ6W
YN8ZfJehezk+sS9OkoIRhEOC8hDYA4yRpvvqP7HSbXb0hfXRIb5b1oggIdB57K/bXmDPlOHQFU7G
dRKWRxB4nc6nZqR0a8gOX9C1DUbBbyxF4j4K+qycDXcdUU8mDHgzlpwgKDA+TgQBQnHWTb/vUjP0
J5d48y3m0PqP1DUnbtQjcyEM7BbUZv4cHUGzmvSzOj3GnMVo4UaCIPfSPaLjdaxbvolgj5SDxmtR
Rg+sz5L2etwsjhxWtR2OCL/KhD83bivoDiX/8LchC5DzrnExojcBOGmlvKTek/fAxNgMTFPn9Va5
RDHAfrrh0LssIrNm43aDRSYgY5SXLYwquhn4opp9HOM+F7DBLis4iyxzw/Pnnua4A37jxmwNAmFL
WKjA4+rlasxw4dH0rxgM+VUN5aef95X1qRaCWJrxd49gwqkyDvTXpitVB7xQv6BT/FFjvpQnvXZr
Df7MeV7BBRo8oMYOoj0S/RxrWf+t3FTIZynBllo59C9pIrFcvH79PyqpSQ7HUy5GyH6dB8IZnPNE
5Nj0i+NhCq9DL+Eh1bZKfcWDBZF6ycXcqx2/qM5L3tHNKjF4x1kdp6mfUP9HYL/Kao9Jm9vrQIhi
xGBVbcAHGBRq7EzTddNY1p5tZy4rLgg0amaISOOTPadx+hJZSasI2r6gAc/jEk07mPu/vRrp18k0
n5q0+wBixQ545H0NIV8UMHaJ2EzMsQFvcj+ruBuuFjvKubyXWvozpMzGUfbak7DWRisDh6VdeD85
j5m0DmEzxRuaLuHzrLkxJRwDqe9nLozOAjA+EsycZZ8kbLbHCcI1B77LWo7PfHzUMLmEghcC3qsZ
GMFv88o11TKgqKOWLbK6UkOIgzSP0V6imbKe3+ioigZNZei/dknC36zg4OoFHSqkQtRM6dmbWvIZ
RXzrleJSLslM2onijHf3tV1SW0lIOQa5PFKV4bvddrfT1Xku2as8wcXTXcbR5qY9CSYeUsNXVu/C
mcRGr7hhJGYkTecbI4J8e7nL25wcVEnWbCZyXhR888SmSKHiYLzsi3kkwus9g80rup8DTa6aL3ZD
vskJaX36RtchExFD1JFlhMeS9C4I+HBsukaAkTM7uI0WaW03mbozWgPazGCTaOWEtEmOkSPNDnKg
sFnp1IlubbrA4bPVyMmsfCdshpZdES7fXjZbkuGtfMBUtZbwSzz3qPMbEPKQiEUwJtMZ3ksHjyd6
vgV3VIIjt2hJXv1A01Ecu5ml2GPviQ544wWvn3m6y52KnhVBKY5kGrDN4t55DE5oWkPkUShyihzD
MiO3Um85jABhlynt8chkD0ELe9LiYcG00XXZI/FS+L3KB5/lpUhtLVu9Y2/9E4nuM/3TIONwt6C6
5tE4boWSwKhBpLpTXIXktPmLmDyUBBj8uGaSywreecaPpqmzKTipFb/R41y74eHwtZnFV41AJqrG
FKbQIKnqczHyguJPE3Pl20ohVZHbp0hX0A/exnG5yKJWbb58eDSknrVfSoBszScS6vBChDZQhckb
pInSnnWSvvpMMzeNZwixTjRmFGUc3f3iQBP5aZ2bBharrKu7kY5O6+4yruRC+MmRvjWpqeuRDASy
STNeYxXNtsapMfXEgjWKv1VPw2NnHiIyURnNQXaDRx26QcgaxOexPxSHOgGDtmC4hAdCfxmaHLSq
wNcDlu5FDj7pV964n6y01TiTlPDUb3atZmQqynu3Ftl3eSP02VYv0wVYgJZlGwhN9I7uEa/YsuqD
kBkhh8rkW8z1AUQg0YJ5QGbZc6LSw8H+25QrrgezLmJLOZLynQ+MLlDVvvJXaXzgs4Y6fzlwKmME
N2Io0eyEkT3qWBpIwwb3iF7oZkxp4jbadwXWyfUOkgj2/VziVTx+8uvzZCAo681HrCmxACWg26P1
sxWM3zkWr6Ji9uHRgTzHVVTvw2OUyNckORnXlz9HNwOtshQXmxZkhicUx9NRa3CgtvcGxadS5p1c
F6aDjGfEnUnKUKIvv94Db8bOFcqWi5CzJXfTigaoK4j1zGfZllDUlGBZtZ+Ta1YcxZQ1YDd/LS7S
g9vi72ZMkdUD/5fqTonvoKubPy37v88bUOB2CJ25zx0h70g2N9D/FM1mQPKWf4BZnTiDLOUf8m7a
TBo7WWF5XUr+oOULbuuxcjUIDArJJkDt6TdIpHSlfoRJ7J17y1YMYbAGW6KS9YnSXoxybF57xQMa
SHlqVSMbW8WEDT1rd/k5h+ImBI5T3iVEu0F61blOCJ8CsTbKZlIylsuOORFrAfcBlQlLaKLWgT6p
wlXLOoa4khxQqg1C8/oUvxwZWT1HtqMjnYfthnN/8Yq6+c8cuaJSO+Gf4PutqderkBT014InDiRf
Sy/gkJy2XBb8a2yLUg/vzRMI9hnOfN90S/HELjefO3vhcBGErFybDG4bCYxqQ2BoKBQNEdTxnPDh
yBYcBYBtWuovNB5TGMVh5Mvu/1ASHcbr9kwD4Fw1+Ur6dRe6BpOiTp1Km+mu9h8A1Ufj/pInNcSQ
EG7tNRpY5PdtNefF8jMyzdQ17stTUvoARv3eXJPNT/kjOZdJI2sN89t3tzOW5ydtqEVXGRfYJu4P
CN+/5XpDmph8xzmQ++LCg+JuarxYjkqoj+4OuWGuCYfpgRmgQA8o/zHplMXMp2Dw7+wnc7uzeArZ
fFv3e7EdFBveDvz8e2ahOAV2aOHV5PZnyT6HYQrm+2X2nWgLS1cyN3a0HONJjzYE1U/dmCMGOLoE
rqF1iRJW802mvFhpJZZhXR9DPOHiBF/nE8L+jzCrUwCwXjXfmFaSZIb25ghTok/0m2gA/MzghOgm
5XIIyNAV+L+nnnClm80eRBHppKY2OT6GsUTS5njzPvjWullBx6ZLasYXt9He++cnkY5CP+EwUSou
dNxsB1O20ay3orFbknKivEdiJOgh4nf7DnDhM3SNXzLeLPcW25bdZamTT3YtSZ6lKRcBI3jZFGF2
M8vWWX7MyxF8C4T4+dIBQ3b9Pwp7vGBkaHFKVomBiP27jEG9uAAXgJK9JRoENY/ialqyYbItTPuh
1Yr8pbCLYTmrF/X/gUaP0PcYWyvcaewKIUhTQDbqgb51UtUKTcuh40Mnnmzybz7LKz4NOuq0b+xp
SKmA7xKi97HSu6eSw8xmtpNrhi1eS3cd/OzkXr9uhOR53Sb69TCMGIxYdmYRTlgaiUU0hE2bY97d
AXFnv7ETBw0hKjUnQjhSxEj8pj7mwXs+S68P9dSxnZbRDe5L/rgTLlg2/xiRk06rvRVkz7R7EXIh
yPyLtCv5MWbJGdjepB/+HLQ1Ci91IR4XQbd/tc2EsuWJ+DS50LHwV3G2GpolrK4B4osH0m7OI42M
d7iXrzRPhTyHXzA7hIcIT9bcA+o3KU2OmlkYTgd7G1XhhqpzYc7bj/V1irCLyzUIhFuKk9wRcgCh
vak8d9+MVw3eMJ+RZNL3j2S14UnohqO4qoR63om0bO4nLwbaBQ2IjZx1XxUm9tYTYLRR+V0tUzPI
hZLxnHQCWtq8yLepetKjwsR1Ue/+g5eVubJ/kV2o68hmS1cyYrum8fljbA6KPUwUUrCr0wVVuE3P
e86JPWoTGZUO8YWTjpcMxfYHblS+JQcIeuOukDci3herkQPpCmmKhMcfqLEXPYCeq5Hhtr+MlaMs
kK8qdxhJpsw5SW0kZ81+B/JctiF7JCyMf7SiLKHWnZSz6ao31YB7/R52agu9mZtVPyRPRKf4K/Gf
OzJvbEcxOVtPVFbv3qHDqBF8q3b8M+wK14RFp+utdPRr2OwJOc555ZdUqOSh+RCyNmfZwc1ipK2U
uBX9pvF8KzxjEFp8yCr/FNfpW/Q1+3QZ3CgXHGTAkqMHlPD9+Zi1DrfFiXUOuTJ6yndMrG8ozfbl
dtvK7MgSqQKGwMVZMZ7YcvnlrvWo9+geMiYW+9a7QG4NfKRm/KDwkSVeYTC0dYEh74FBFv/g4+9O
rwcfppVqRqA0LbspYzoybBhByyLIy7qIakcpPTrHdg2bWVPDeaR6BpEWUia8jT45te7IXzsYfT8F
9ZNDomUhwIEf3l4SV67fKghOB9f12BI7tUdTmNxftu83UmOUh+PcWo8lMWFrkd8b+BP50aoQNO73
YtVRdfRioJ5gHCZPyZys7b27emnXI1cJpaFkRBUuS7AraqrRWQOmFqgqudPIX6SoFXh3yzBxaD4P
iTWjMPnTiSIX6mT4yscOCtj51TLy5ERmKZToEGtGVBqkJl8DrAblJ4eu+S5jQLMlsz1rGLjMWz6n
Zio1KZKjdvLd8CQyJh76ht+UH7EqQoG8kGONACsqlNV3loDroI1J+8xj+Y3UPk0yalc2o7w2GG+j
1kWYIVlX8IMDGCuoWgbcwphN2BzJgZw6N/ECenM7b/GL/V/xUMjipURqNbt6j4F1d9Z65c3Gy4Ly
csNjK+U5gTDcd5g0bXFUEksBObfF1qnOgdcOKoietbc4T/ueK/htNOoczuUsMCsSZnGcaTEB9bTS
w6QIDCqXUxzlP149sNEIPmf+VR033Ye4nqMYCZou9Uv0phC4Ga69lpvU+Dyqkcd88gkVE7zZBjWA
ng5gbXQsNNa8cRC1kY8ThGqTdSECORm8POTZXnMSk4L27plF0X3H7Y2WCyRMG5DtPA2+E3c6RDDr
btxGG+tXxan1TdPGpvGGSLLWyRTjDs26HzZKghrxSmBAFKw85/xc6eWW0D4lCViKMaTSRQnR9Cx7
BfrZXRvpfxI3Eo5zYQed3Wh9MMClb8NQln+bxNOgdBOoD2xAcVqv5pEwNOnB5mY11lJkolmTEdcV
aH8lrgwu8oPf4off304B564+NSbA9j5TiI7HU5Azintkm3XjcrVxjHF5Ac6xCyXmIDak/zYF6+F1
AYE9L278VDN66hsSu2XugTdYVcX0SqUJ73jz06V4LjjOuyLcha/ZUYl7heDW+zAWmkknBVSuPHwm
wQptJXkXcZ1H2Xxu66XCwghtsph9Yr8gglfQI4HTRmZlbl2w6ewJk4x3FqfWETMRiCMiGpLe6rwE
DGHzI1ccJDT88uVzh8/yllFoU3zozdVjGouqQhfeuYIqZjaND+k+cyhvNbzXq4OIYqFnLaA5DuiU
HBcABfrMRfOxaXZ9sCNueSobJWubrjKD8dfyOaLWhBFuAVY0jLxkU4EWsz9K7NvLZkT8KKTr44K/
zaG59PuzKqkQwODZdOyIwJjZDArTy8AaJmpv84bX/QYPNdWrhOfV7ID2Pr9cCtstFqyDlYk7KkjU
osS4EHtYo3IEXb4T6BanzxtTNiELZLxDNOYm7bjgCrc/jg2LbJBH51cECWt7KufMPOHxu0s7QURp
5r+X4U20EoT/Z4eAw0pGxD51ymt6Ff8hOjgNM0ocJUEICMnUkbQoyQL8rN1XQvFdozGuo+Fkq1uv
hJlIKl97tEzQtr1GPpm9ZhukG+vp9n57kUxoHkrUkW4P8s3PbJbe1qBMOdg2d51n8JvkImaca1jl
FZQX3r4WUhUJxLMChmt1HxREGKNEbvd4wgKhsoS8Qdlse1N5OakdWfB88PO+E7+PWf31gducBu91
isRIag5GKjtKIGmhx0porNwauDNiJOU+zLAwOEcbha2G5i4uIU6nKXkwyEwFr6YkaUYpmpiyK7Wk
b08YR3BwaMDhvBU1apm1kRrr1cgTbFfob9d6598Ad9J6EF8ykuhM33uluB7OxeU9rtk9sGKDd434
d0dV4SzVXTFaJFnKuXMQX4jMyI4Ct9xPHshbU3kAuWKjg2YUyPuvuLIABkBX0w9kvB/GLTRRSWTT
838/AIzLvOynAF9T9b6WoFVGMsrMp8IGxgG3aYiJoiRiP6ep+nKTAnS4bph9iaLqdK9vAIRg4OuK
rpqvmKoKJj6YJeXKmre9xQ49QqyFWcCEZynRFgeQzxleiAS96VvGEF/EQNk6VUsLWWs21TAkQWlC
Zt27o3SwOvK/eDfOEePOYn8bDUJz8QH5K8fd5rI1Pg+WtHdcDGCeD3DgioS4hLpSLUFRgXTBQKAp
1KvjFmL8DiuyseERzFqACH4cBWBnuTkNKBB7gMAvj5c+ZHCI5a7iEd4YD1TY0qlqASb9Tv5BIg82
fxtCcFrd6syhD1wQZUaCqBNbHgu3R1gcVy/gpbSuTtZI2Io1N7ZAQds0H0mq5NQTFeVGQ7OBoGcw
ypamlEfnVRBGokEBOxdw6vnxRs0EHu8/HTw3cA3NFu4rKXNfOLI/cLUeisRClWx5bFwGDMvEG1wE
GnogJl1vcb3vxgdRBTBOEyc9cJiBKZcBYnycZyMgrDDw0hB7ENRPWgWoFXAklyXUoD++ktydT84h
FTMs68THHYg7xmi2WTyt8g6+tIurpT01n6pM/P1rb/+SDd0R4hDvb/zL010G5Ll7UslxyKOnbtBF
1B1k/Mcz7QxLj66gCwM7z9AgFon9iHG3uCojup2Xitfh5nbnuMG+sILQxCY2nb0b+q4SPQF+BHeS
iK9u+DDpyjnbG6qJQaXeR/nF7uHDxGJRnnDwjbrMNBuYO9oCCRgE1EwWyXyg3lcQTIKKrChlXNKD
OLm1CJAN+NThA9EVPsA/ZEh5jVXp1DrcxaaWficXxIpbAQnOq6TQNllWP7epdh56eGeHoMrxeVem
M51F8Mh9oQw6urosgDYupcidbfyTyX+ny3+pjT9ZX1L9XUl6I8M22/tjbJuwFipwIm1dFE8/NiM2
zVsJmA0liaZavjyOIh5AbxWTZYAKxCf2JKlaIaDS0IueSN6OBMt7GRchsNpX5LqZGuRx0oBokl4s
CLh23vmmmnYT0cYRdZ71gpxbxZ/8ZtfiXX+YV0b89gnW10H8aDTF6pz8wW4VUiHELpNubXtBrPiy
7W98j2Z7bD1LLZ5+s2DYDp5P94Jh/+7ogyxIOg7tGrPrTGQKLqGPjoTxezjQSvXJLB9AK6SouM90
yNA3hE9ULpu9PTE/VJavEf1vL2XWmHBWC78uZxdgR69upPS6/gpR+hwdJdHbYEdeHFhCL47zcZmR
GQqlxel6qX8QULRFgYzf8clj/nBWYz8Fj+tMl0OygytMV5NYlK2E38mUi0E9W9zEPjsyT+2XGEqK
UKHYnVN8wxTuPU4J9cnlfyf1LfgGoO1d13TqUdQZFPbpA9f2vpHYuR1eednWJx8eI/tBDSSGDhHT
pRQZrRj5xYraT4C784bpCO2Q8zOSSsl7kqn9WaZH79GtlpL+p5ijDfyquXJDzGuvN71MBr29ZbME
XHeeYEolgigWJ74KoTgpxushPa30jqjZefxKAScffBeb3NNFxDHqr/ETOnhb6r3ZVWWVyp+GEzGI
ezq0GZ0DT9u42bKBq4xiRUzfbaysSufQqUbtqgPm+qAiYqKAYHI2wwBSWZbkp3sJRdVgBKKLRCik
KqU8Flnj1TLD84DQiSV/I7SrlstHfb2HKhSF9N/h9OsJ6HoiEpGKDlDYTRF/EXKnLQ3YapZ7rwQt
ulLMmVMjWwnqj+2roGNdAoCdruMTSqFQHkVNBLIuGka8YuMoxIKT8o/7O+oHaKlAJbg6RSI/83iq
U1UjD1A3I+LkxdhxyosKk8JIHMVwyjz6G7HwIerWfLlExBPu98Vrzbhpfg+YIwgPn5guxKRhCcfo
x4Y49BdWQ4K3bIOKL/emf1QcFYKS4TnGO+mxSO/Cd9+7yjya8zbqRDkOkdiltLQ39D1ID4CIZwue
JHuG8dAL9LZoGC9k7fxWvXsRG999GpH7fOhj51cI2KUyS6b+TkDUlRtz4djPjGbUGlO/PfJNMpoF
HhGx3oAWd9wG4ftjEzEbR0t5mf5ZJk+fnJuijc7OMRwDHWwM3lrSkPLPQkJZszGEp3ilGsk19RPn
PykurP1qEO9PEYZdvVCmmgvy5SO+PgXyHmwulAkKr2P74uGpNkcXOXfpBN407zBZT/FY2dS4oBML
4feZNsoSAkCHlsGpVxkzA0EA0I+GBZcOCAzeB1wwhfiMc+VLQeYG8Bk72ulOjtFm+SpB8NMpi4Wd
6emNbZTi4aWjW9jS/shOz2H+8gziyTbC4Uw5qwi4yt3Z7Bu6NuL1Xzg3XXZHUif/riZcVxhajgi7
oKPmt3j9OhQ4RosUuSkkBrga4F2kIvxRrc4/tQ1b0AzV1RxdMbk/IXgw4ZBcXEgxrsOULTD1fTdY
P3cOEEXV+K/MaKExGqjXC09fE8cYoa+s/MM5xjxdj4xALmA6zghS4JfDOTk7LAzhh/hGcOOH9lo+
P9Z+M5+9AEmhSDlFZuhJvXA+hwArGdDitRHVqDXM+xm4Q6yTh76ML7fIYZd3eUA+sX+cmWuY28Gz
1rQz2RSEEbNfhPC5zsAxHIuKcCUINKqU19Ukg6607taQQaFgN4YhUQyxIkIvrMW1+53Cu9vErxKV
Dx77XFBL1rABIaYgdGRhkwgmf5krEQqqb5u7Mdoakhee8h719VargZwuEaEXnJJfRKmKjsqu7GdW
wMebo3D+XPihoApm8T4JSy+R2HfD2gEb+T8uSH9hEW9tsYAUu+37crmIbVOTuw3DlwlnfQgdKDJo
l9LhE7SYRQS63tMVxE89FVsnMcqVTRDfks4Rur1zClc65GcUVJQ3t2e2oa8QOLSCKw3HfpjdacJp
+v9ZikOqxgG4GDd+CPRLP0sOlq7QgAX9RchA5pC6H8ZiR0iRKoCyF6q0APIlUUBQ4pig/LwKUKO0
j5upApTfIwxSzgMz0N8y4PpeREskOFbr+OGQoX4KYkxvg69h44fOZTaRDq2HMmC1vjSMDczqOU/8
c/vxlug0mL2R1Yah657F6V8hS3bGyO0I27In+QtxjGLzfR4yIy2yyZ1pAPRGNOW5zpgo3l3n0EvP
FcWuox6BT4OTKg+79OoaT5IGn/qP5F9GjlA6VPDcG3KIY3DdKVkJlQwNJiazu3VsOEbybigIqAZR
L55uTBK/YWIXCdUtRVy4IjoZ2aRUyqrREkaiYfXECivlQTsKu5x8z8z812zl1DSg6QFU4zrBZpZ7
9rjiiWMW6G7z0B1EHBcRLccHKMQPkrn2WrxwzlIa5YqWFbzF25A5OMUAPcUjEHUVlwB29F/mNHRk
k56dS7EQylW8gHOPKTO/oP7JD4+Zly0M1Xyw4RZhjMol7anBlFt0u97e0BTJvRif5BYLClO2hnug
1iElP5t4NXAk5MH/SmD9n9eHIHEkkPnNk04twnWdHi3OmDFy09urnq9Xn4iraX9aJz10OEIhD3r+
tZefCU9gookJVXB/BmXnijsprH0LyJSr76oxSv14NmSzQtRISSirYDUfpJk4kSylUamodlYsUqI4
jeAGESgyl8aqOwA9qNXMKbppeSZaECL/dWP1Vj8cZu1UDtB02smd2X/mCE3vJWlSvT9KGTaLzbV0
1TS9OVcrb/BRM1ccALsUX2uPXDG1Pg2WLXJqpr/WO94vYMvTMKyxby9lroMPJCTA10grnqvuewGq
gV9zV1aAhSM0lVj6uMGEP31LhSR6wRHBBclz6eAa/JcbHRkrgShYXAFjL38pLMWeoC9Pzx6tWa0E
5o8IhIsNInNuYEI63w5hAsmmCBtx2tXW5C5/qM/E8WwW6ttJlOHomXSGHr3uYD/GhmZLEilJnfvj
W8x2HtkfOSDJx4sORhfSfJL0uSLD941eKX0MtZkKSmu3kj5QYswZJ8FQwcVDCS6tlfNs6O1cvK4p
5GuHLLj1sL0CGAnG9jPGMnQ/yjPq8WdoRUhJS2W/4e8+pjAW0Gsnqr/FT637uTJzaKaPm8Od9o52
SGlWDI6hOIqGBB+ATi1Lf/E3HAxrnH+1qza3fjNcfmrA0Zg6PVgkm1P+Mp3FqO7ZAOXnJ+YBCrQ/
32z24jeKjtLDC5zHrKt636KijWaau3SPpRrtnY448rvqCqXzGSVcDlZN/Oz8cho/I3DOS9P+DfVo
EPT/BUzao5d59NTpg2HLnv34pvcB0e2crvWkyChGRJRVk0k+g5AacKFuN5nxQ0RHKZVVG3f+2dq8
MhXAaci86WdCnqTBOJ0zz1MjjxeVkdvcduZqJFaNmozH17GIZjex4YTRDC9mTvW2mo/oDSoRW6TH
hy8EefATIzLR6gHx2gnBgeYVrp0kGgJ4nD2XaPDY29dNViYHvYSa7vM6FLdLlosOIDNyMTSB1xOz
v9910AGVu2gnmGraVjQsH5nI3LY+O4tLjvB/Km3MaKRss3s5rfZf75ejDQRexRfmeQuCdb2eTu82
K93Q3kxJvInJ+hQNEoFpgjqPNUrqRr/oexQHNriTXmJ34YmRZrIQqwv7ScfKH+EHOB48pv1YiEPd
YJeWApyYrVhGRiT0hhqK8y5NCKtA5+kb3BEOcJMUSeFjJfceFc5PqrvwoCnMjqfW16woVOk3D0V5
jSoAuB6OoZQaUAkWFlmgAduEVqufdfK4b9rEk3iwkWKYV2f5XoQqYyrWG8IRoBpfVb/eRqixXww3
KqVsNFwegtTsNgFeYOeg7/zBRS5Hud3ifxvAh4UTmZJVQg4Yvfloodw3NDl90VQ+29gv2UGK++Xz
muDcBdTra49ivF8QuhBSHZoN9eKnUn3cPy6Xq7Fgeox/8Rk1WvYIEdivn3E3yJBUXFUtg565NU9x
ARQ/ypPKRBagZTHYI3Yh9Iafk6EDR6rGbmvc9HDE+kLkuLXb8Mo7ElAVbXQgeovCyP5jY00Et8KI
fKSSPUZK6hPHmxFhUQj1PKv7Ls1a5eJaG86DaGCzwuks9XpPrcvT7KfuclLIy8UqhpFPot400IDA
Dl6oIH6jIl6MHbGr+Hr3Lp0+Jn8Sny5uReDWA2SFJYHoKuVUUaDvbXgLgrKhgblFkF/RR8WCAX1Q
wy5vI8VfPSZOhhtlsMGk/YUS2k89k0SSasSuUHoaR66tbqHnlLnQLWc51OXHBNl4Oxrw0xEJHPwC
C3keX2hCDD/EyvF5yV+KaTUrmF/gbgP75LXeOM4jBFO9jj1nyF/RkiGrp4Pv+Fj1JhYmKDt5ulAf
Sh07VXNahs2Q25hcOukZ4C/UrpLWIuGC8MnZjR5tnrbPtdSvfA1fsU8wsgeeWvpIP93zrNdtLVzc
L0vmVe1yLx9NAQiPdLIFSFQPv2k+nVxQF+AVckhQpRmLdDfCCzPkXnmK4BWvHQWGwlM0UAyXS0PL
ODmoZf3r9m/21WJC1vGFCVuHiliJMuyIBaNRH8X5bxIeoisKUMZ/h90gcKpPtG7QiBP9lcyqwD42
Ri+piBPMqhB1QSGCYPB03WUB3Lyxf/rt92hRH0SAfGMKJGRQrDX9RqicffZeLS/eLJQl+bJnb4kw
rb3BS+hUzsfOgxjqlKxmp8zwxRoxXZ3xwGC1qv/K2Ga6fIoCwNTOqjbjSR0xfX9X8dgsX6dwL+F3
kp4+j5eczXFS6PaEQUpH6NBZcSgPrkQhhpbYa9Oo+ri5gNiWMPvPkXGIL99yY7vsVkRscoyYVuJg
GxDFIrfx04kTGo2ZmzpyIAXuwK/PhxFzajZfMaOqJS30veYM6qOBzO5aIW/9OjH8VwTBEudy98j5
yiJ18PG0mRktVJPRe/Py2udwpDo55iDKpTCj6Mv3JvHW1+Zjj5Mwptnp2/0U+6fB0d9DJuMGchGu
au0MZa6kkEDK/fgtXTFiSkOjtrNvZOC8JLAtu4Rtsc+C9GKJMl+7Yms+RN0Qk0IHDFboLe8o3cug
MU3pKKNR+8G7AdEEcYrBUET2eYtE6xtv1/wYb5bVIW4pN37qE3Xz8TcDDU+GKmaW1rH6wsrlyo2s
PFLpySxnhygZFxtkfAV7X3u1KrlRraho16ZVSFXqHJu1oVdH3RiL/RQgTArn+k+UZ/IyUTOddD7F
IhhyMEBuWtvFR33/mapRUDTF8bTN3tvB9O5SJagP+cU0gP3kwdLP/1/AprzSt1vca9J3IxlicntY
sbB9qt92ZbmOF6t/1G79CthZqFyBSUA9nPc9c2HaloutyjaJDrIsNi9Friyy/pnB+Kublu72MQRV
5AYoN+ockd1B5IqcS78hYqawYtS12yhJB+Elr1hqupRvfqt65dEQIBVZUrPwk/DYabr3DU4P/o4g
XY/n3RRqh1a5Z5eg6+u1h+RLrAKngW7sk1pYX9keII9xHnLUClB6D9jjZ5+fbyPYMMd3XBoCeUy5
wlRXvSb3Y6gWRUV/K+VneY0bXSrbQAyttD6XPjAz+6SAVsCuXeYGc/wPHBGgsXvcA/9KlhH5HMvn
t7PLkoUsJNjMl/T3JEGMzCezyV9LcIXW3/BeAuz7zRIChUVBawBEtu7krU1LIJMwRte27Wg9kay5
gCAEY87bRoYfdWqV2a9u2lD/vDfN9mAzv92Erox6A+R6LVGn2MYvKIciaMr97cJeZN06tMFTV/EG
1zTilndCLgIR/VuNMpIZM9MLV4zA4FyRIZDAscZnU1XeHPZVPFR54YmWi4YmRGxpRuViIrElbOSb
j0tTRuDo3KfesYCzZUFu/exKJZPmRQkS8n9JqfkdbzGRNJsswHRnuw4PRWQAoEug6D7gbcA4ADUR
9xseAp+3uBx6M1Jlet9F/AZWYSviq8nDCrrtL04v4+jcTn181Jb7DFBjil2yjXwghIwCvmGIZUNp
YLDP3m2f5ySdjG0DTOwVKKAffjWQXBdoa4TD/+z0i9pGpyFzW2bb02vI2B4N9+jWXjmR9g9yz1y2
6JiTYNRrV8juhRIMUbJogqij74drRav3Js8HSve+mE4BKIq+9iCyyk3C+ByHLSIRIpCe5Ub7H1pR
cQvwytlsL/MnLsYammN4PqQ0zcgv/m0M6y8bHuxDKKQKl5Ij5gDy8j0YKH/GAaBpBqyxOrubKvXC
g/N6NplWjxoUQYcyxgH9I7dUIBTqlUlyYQ4eFuxF9Fo0F6Uk4bqIAO+1PquxvCKVztKRvaS43HC0
GKDV+QkHfFIP8qvDmbMmqgeX7TJ4IVYNc6rL/Pkj8XO2RXaqQXVkKdS+MlBm8ZILfg2uOP3/KYRR
S3ptB6uQ7r1N//riaPfJUZsXPBqPkXSF4nFeq/Xr1tCcl2q6yh895AsTley785bJY27RHMwv6yO8
ecQ4wYHTyhgM9aWyejfFOx5oM9Quu+oZP3j8ww7RmkWDBn/0lo8E95+l9nnHrOaUH9Iew2h2wtbq
Wfjpg/BnVWtHRVvTIhPTkgd8gaUkx1XnsSoGlBnwYHH/yL7rmOBWFdXKDpMYkiXG4KxVOopNOhfD
YTmZ+znswAbLpZ7SPfkKSExzZP8SmJiwyOI0GVtavYzsOfVEoVVk7mQ8tid6pMOXgTrrZnVJ9XIo
5EpivdNpgaifxqKEtwZsFkbxH/8M/bk1pGKYSraTpggZREe5J6qK75MjtZkgG2ZERzCCy1SjKZRe
ZRiRu+iL266Rgx1pD8FvBHCR5a0EME51zKuwjkrSPeQ4wTlhMLvpOWQEyi+9O6e70S1t8eFf7rHr
v7nfMwRj7vFCIPnH3gmIPREj977fztej2nmbcjHI7BSdvWRn5nUQIJkOOwOwuUs7y+6aE+hZodBY
OzlUJvryAaADC/1SDDFr8hCwdEV6xKJzeLmlOUS5iz+3DmeF8dGo6jOYuK1AEhVBeW3BHsKRRiUa
5aTpld25TzJ9lH0Qs+59eMcA+LtMJT3PJrO8/2F6LqUUKMt2F3z7Nu/eNVC3LidRGQaexB0gYo0g
CPisC6ErHkn2DAlOgYpPELqT+xWLUfOH9/hMKEE6AbOPF/Yf2pzySNMZzjrC3/HANp5cf1l9icrC
I3ldj7d53AhrsazL0m2uVylJlv172EK6+mQuyQWdVWXpoVqMqMHev2pCG80mDEFFPWHp5YOY+L3p
EfcnOY2I8lA39N4z7kuD2HbleFrMp4U8VVE9pqgdPNfWqSwqKkkZlihP90L+Z2Wia1sRNrKfQIn6
Adyvg3e19kTMfq1oAlIUA2WfcY9XslmO7qHxDr+qzl7RxlbX81pinVPGGTc7veH4sGReYxLUy80b
TCLpa/f4U7HDJbMOlOCYTxJ2lJY1RLxxD7BdDTIGom+x3U3nOIJCSVsSYBOFakty2UYodxEiwXxn
5xo2Ygm8IzPhcpRSKKHC4UnxP6P45DYxkFb1nnpFZcaUDRKpKZblp0RGoMq5KpfhtXlKOdaTa+Rz
MFAwYw6WIJKJ1dI4Q88PDO4U3vXPDXPbzlbCS0EiwEa/wOOxZ5CmlpDzp0mwqB6maBWijtmZ+KF0
tam/pbkaQjxy30ctilM7RxRSMqOSjgPDQ+gEttfC7DtFeavc9U147MLfJmEWAv7WVo3qEYb9m3s0
YgUEtktype7KDW5aQfiemNiB2GXR/HqJwMS06wm6nZCVv274/fyBinhjwcsNJmKji3oWk7/VjWNA
97uO7Slk+aGrRChf9iC8ZjNUtl+Ls+FHYedBLZuEu+DV/FfTc58TW2VueEguPf1P5pNpvtigX00h
fE/1JvMq6KsE9LHZFhxJJJOBPkpsvpcDfO9d4ZgHCQplyKGOfnZxGokknASr+8k/u/CRodHD0BuA
RZrvTODz7jz9lufYYBUPAPI2PTHyukhqfEri2ssTNC/CWAohsfqWhHaO0T7FdUIiUIefMOf72noE
OYvlkokmD2EQBy2l94abng02HnOgpGCZDWSXLrEDq/yziQSObHp2VK0tz1sqkDubUWDfTbFu+dA9
19K0cOPD56pZ9bf5LludSOzF4iCYPmLJyJA8aiNQ2ZZOO3diCj1v6+m3q6rh0jVpT5as/bJ7yLAu
H0QQeLlFD+wvK4hWr26QYUXig3rhLRIq/X9W8sUvtUlXUAbIJK/Ep+6yF9PsMta8ipD0YNutMBHe
MRxnKeKgPhIuh5s+qBSfZ6ljgsKKXeXObljguby/XyHn5MxawJbycU5ZPxxz0KZB8YuOg0CYpl8m
MtkZMYdOGggKsM1sPl0zvadVtWL63Gb4hvOOXJjBbcu06CAyW0ngMLz71iKzI+dLETQeoC86wSkr
b1zouLBV77fmNDjq6DuzlcgqUrwM8FR8oJ+p02gegqz+I3dT/9m7eEIEz/i/8xSvW9KPPA/KskCL
I6ofsADUG/880/Y+uAx1pqBgwK9KQLlej30PYHeyFWqCUHhaadxXkuM2xcEZE9D53Xxa4iPeIDac
CUlCVkT0FKnU+FHUWRgwG46nmtp1Z+DVdGBBsv5QEhWkQQCx3a3TMnsvFljL3TqtvwMH7FFFP7W0
/JVp0fp0h0oAhyXedGBPbKnAgn+P41NLKq3ossaRtuqoARZ4I88OFXUck+PRE4E+sV2ERILOYS51
+H+0ylCd5XNgas+BxUO9OosMKevsWufaEZZYUAaO83I2GA+7x7AvJPRswPlsiC7XpdkA0siCtPoc
sCbq0mlL9NM6ZMyU7t5KYbJ5nOEdqBZLvujnZG6JPN4yPnnRJRowZZ19rIpIMOHjRZZcV3sWkdaP
QqIr/wVcLTcRLADk+qJMC7+duiy3R9+UejLSUrNMyqBxiIHNguQdCmxMCyjEpbW7oPnX4Bp8/hQk
A6OShDT78Y3vNxMU/rzVPZKNLWPfRcNLabqRHU056Ph32tTNzPmTfblmI94PEECOoWVeN1cuhB8Y
CGEWFbCGa+M5ul5Z2Cdey2zilW8q2lvwEEjFzRT2qFVWqmuL547midglHucYWbOXsP8scdFS2QvW
euJ9x6SdRSnj/ZNYcSIZ33ELnX0M9nC1GDMmzeYy9rh8uTbSJPnI1MqWSuQbyIubcDkNUxpvs4p4
lZScbiNEx2L8FTA2O2WuOQoL1jX1BA1hA9ZIEQZPL75l1/YTVFO4knct6LMrA+sl6IkCljdVd6yc
kXCxe3hVwNmt0o3AURZ5EmVe/SgQUbrQnJcgGoSL/8unSzH1c82UOPkpMLBOgQQF7TPnvTnoJ0oi
w4MW7aTu6jx8xxR36QvYGzeV0YuacbgvT5ZY6n70f7Pxd7gq2QcUuXvm8R0wqjsY7U8mexfOsBGZ
qHNJzDfKlfnKsPCEgQUswW34263HPKwYC1wZp/+2NkGkcvLaF5DxRA1u8yhspKs56Wyy4XIh/pN/
bLInZbRWUSsIqLzdWdAsrUKPkduRiTJhcw0rP6GlO5T+VDeyub4MZdPeqY8yHdaXh1lguDz9bW6T
kw+yAUskOmMnl6gLN+stczC+AQo1k/GTV0fYI/4EnRBKgfoWTLJ9BM8aJ0HHnTr8t/IQ2WEUa+zb
7IVQPdi/tfQ4Yh4fuCOZR7mAa9tQyEGOeRERwxO7pcDghGdr2vvqThb98SCp6RCMOOdJM0Km9m0R
ATD+5M2fG2VxY9AcWFeXhDpbYYC6Hy85/11Aihmuy1jSus6SKIQUK04vBZoNJPuK9EYBDkcnOQ2P
dK7oZsaQh9NrpCjxMVpyHx98NVMeXwVTVcvsHv/cOyUxAb30h+GEHhohjRhJG6Nwv+lWhnOnSGwr
23tG9w+StE3jEkPENY/4udNqUO87Twxm9zsGnN/8r5Ylt7jfXQxJ26TOrZBtZXAhdYdI6VYZgHx+
QwR4kdi4yHFeVUT7I6g/VnjwDq1cW2ATo+3pJsokqzbljdy8BcRJpBK1cq2umUlYDMcPRRfXTiTm
wreBNLKMCFQNP2bHTnzeLAWgxpvP8arLmdVcJWmcP7VLXQocMWB1kRSDQHz5g7Tnq/Nns/EOfnOV
R8qyQWdyJpORKqztQWxt/Fk9rKii50XW22TDGAX0khEpVAJX62jeh5Vcj19XmGkDnquyxQ2LWT31
YH2w/pDCOZSN+BAIEkYQMoWgfvWq+2PlpquLfcwkR1UOSVadu8tfXkK5/TpI+pys712CvxO4dtkv
9QhHnPJw/kn6shcftsecjuWWiuxUTdinisemZot9QuYkWBeWlmeqH6ykoV8rePZplgHheT4+L65P
EQiPfRFbje7DN7uIRBnPT2HIKwzuFlSoGE5X93zMG0A/6JvD/NWo6ji+qqNNsi804BhznTAXCdUh
m4ySOvFTca/uelfcIlIwOc/+a78EJ6e/GLzUV4JiU7dKt+ThL9yYUIHoIac3X2g0X2kKeiXttrYF
NggZq0ue3oV0xTG9Iv1iwbIRgwm+DXFvipgB/vvJpxl9qpY9hxg9UT46rMbtp+eIiwThyf0vJYS5
VfhrrxO512NBhLvmPdxahM9YLMhR8vaLT1DnKtXLvvsJ0qZvc+ahJUA9XCy3nE6dFnj50ELIieLK
RuiacZf7ll4qD0Q7/E99fCq9VswsaabK02E9Ukwyt736muons/rUe+7y0D2KD9rJUEUvw6bzcl/v
MBlFjyVacNuj98HJ4bu7/FOWUbcCw8BggwP+E1Eq6A6uIPDVcWCPX0cdu/nK37/3O39hT1rEbpco
uvkbswN/XnCu3r7/9b+aDlka3LUvPFFO6+3/TaHc4SRlP8QGuid+uDetAI8weC8eHE0jvAmlzUre
wzD6Pq6KSYDobOrYHPA0d9VOf66Ttdpkbp9BVZQFBv9RzxInVnhP5Kta7qTWMi53I24vh9fyWmGm
t9gXcVfoTfs0z4BHduVGaxIRsgRfQrqMu4RrAoww6OL7VD4cj3AYeZjzgbucsOzLCjZUlP9DlVw2
F0ht0irN2K3F0JZJOb1yUykC19+/hWxl7Qk6VR4YOojjoaQwD5Y1wVdRfSb8AQJosdqeGS1TvJnt
vEp2m1a9RSODsj68sucRo6FKUgsl1GCmQNMePJe8UgwfnEeixqQeGTlRRU4/ulT2Fq4APDQ5QFAL
mHVHRtJPcBZQwzckcrT22XU2XzToLaZccdqXTmSzE/Hj8StV3n9CFekikRQIM8T5vUKky9N002Sc
A33HHqTF8R0NYXMJJZAFSBHtVURWfsixoQTRIdO5hQa9G1xfYCUDFVlkGGslWI86zR0YAHiIw71Y
yOMhKTAMDHNnQwKZnN1N6c2/BAFm6TQCIaQ876HOYKLCd8RU/bYcZn6SYwhMImQf+Mh+UNCMCiB9
ydWN163EyKWZFbYfWi9z1w4agT5a7jKjw8Hoyacx6duuqjhDvxDVlZB8fmtS8HKYGbGGZ4/I7k1u
XKyoFoCIMp9tRh4yl0DWhcVpoUglZVkv91nTqW6xJjxrAxBJFhwVDvPIsVyZL5RtWg3bicwdNDMY
DQeqAWZiasXIdTtZOUQlUixAd14TK7kgq+m3J00RgUrYVtZWDQ1FJaS3VHlzalQsnuDHB3OA2l9R
sXG3TAMtlo8wsI+S4gk1zpbrvb93bV/Fw2kvnyN35BbTbcTewAY9Oq5AUPwGWRr77TLWmWdiJYo6
kwCRmbppUj1xhVpSsj7z73w9Zrm7ji0PDbXla5iy+BloRsIeqsMPPjuPEgRH6RLJOSf17h88XXnw
FGOMDZwaIJNSofRfU9GwRDbqBDmcVFMa9mMWuj9i5LQBiICK1vEL/3I/waWnNRTTEYARQzKe1nB7
dS7O+vbvb9RL6h9epxHEgJmllktE1X2f04WEzrwbL7/2rMR2fccXXBSulhYY7DqqTFX0+uwPR8s9
ZMMV6X/IoEI9tSofCDGV61YPGDcL2a2WmnslDeEXpUpKVG4vY03vHHq/CMhiyCWvZvmgumyoKBCC
FHEhBHf+e2F04aRj0iF286HwrFETRWmwHT6L4kJedOkJCqjZ0qZrZVL0tY0oDHS0jSZkr06oNhFC
rbPGjey+vo2bhLsa7m1K8uVJm5syMW8OVWSLGexDCOBzjGKOF7rLtNLhvqAZDWXgr3FbKpIbyU2Q
tcqyvYDYjjO/PruJ3ueDw7rykWggWvcq7l09Q6tE5ymxteLIIQDxfDmsjGG54uEPUTU8JpuI1kjV
AUTNBJckndkppuMiG0cA+f2HWoMoLurBGnCbBJ6Z6G5rgTaT213YG5tX0MA5qnyfzjpOIj0KW9cV
LNMzk3NKsPjI4YFanPWvHQuGFR6JqoAgi6NusgdNRc1FFi0FgAyKHwSFeWuWXfxr2hWLxz410Wrf
CT+O80+NlgbHQgZqNws4UEG0lYeV4gYOobPd3C35TrpNrLcLa37RT2FumQ5LqNQnXEyY2HbsygrD
U0eNcxAL5IgjcjGugO4r7m0fqM8db2nBbyZyCK8445b/f4aHS/CfEdKyhRr0rNG5lkjubHAgcgvl
D87BqLofwbSYTspUZx4cMPNhHu8Iy/5hXiN6tpHM+rvWgQVbklF0jw+hVmPp/sSeyAjonzAaZFID
RP9YpjiFmtcxHDwHrk3q2XGYfne2gnfcdXhlZsHafPQqroB521bjFI3AZle6TyDUzfsOMxn8AEzm
l61y2btkEe4JGTj6ez8UJmi8aYa94DMJESfGqK4HnGbJRBu6L2JWcsOpJbL91wPZundrY5g+Sw0u
awHszQFaHWLErlvue+rClU4DMkZNrxdwehybvrE/O1bhEo6nDoV7PuZglAHg488L5Jn8l9y6bwIg
qohkgTT9XeiQXWMOfD/ox5cWL6itjYggqo/FxTbYbYn5qGjh7vNh7rtPrx+naymaoez8ayp8pg1u
D4tmlw9OGtPaQoS07FrwxOsf3/xufg7LqS+YLnKRCRYWLvVR+j8FMXhkA4eofjlEjFJLOgDKI54i
6MH9VQTl1vY8wKfol7WP5ZsOKVNPLI1SfoXhytB+JWSHJFQWZSxg5WBlt0Zp+ZFTSiHO7Aqb5cbI
FBnMEYuOBZ2QTTMbWOb8brLa9ZqoCHfWxbPmGT6cZWm9H1pwVhCtHGJPBMaZGczT+ZbTNdzGS83Y
L9LmHqZgR5ek6Ia8ztK2P5CiNPRsgxqAK7W4bKC4NP5juUdoIGakqmkEg9efWQi+G+QkE6Pw4Smb
Lmq8CeUvRf3Qa4SsApCQ/wULOsO97EYTw+Nr3PJb/BnVckeNZ8IgDcrTBtZ2rbZJNkcqQvUuDzpx
UWt59vgbZ72joJmGHyroXzraGci+26dv6xwCVJYyTfIVOJc7V6yzHgMO89y0XKXjvKy/rX2Sugnr
dHBEu9/fCOfIY03NbIcQaBJu+VEiKhXWWMW/P/m5k5ZAMzvu314cAkiZOKU9BnVrqMbpVkH3Mmfs
ScY4nslp78wRMn2OsGh58wd9gyDdcQKpbtpKv7FV6dq1ho6hbuNtORZOigqwhpwguG6A48w0wJQA
Zb9IqCdZuLjOf6wGWnU9exzTjx66V1Qzz/6wtWjW4TWLupIKzwpPmVWvGseRwCeSBF49B6wO5d4+
9SYY3osoxZHgiX0TFs4jf0qpHCkaOg0PykUvDCnDG5UqAuITsOdqbbmoV36Ge8pv+vxQxtRmOlI/
MOT/NNuolW/kB5yQcBBqa3pbcXLvUDgf4ZC7JB6/ESTk0vU7I4IY2rdmNgkZpbsDqTuSXrVJgG0r
E7GRXonh8zAE1jo2hvgh3OeU6VlKL0fuMkXEvMk24eG7PDZPJoVM3BJSY31O7vwHcuF8iKisK0BN
4GEPmBhHZVxaxGfSvrnsH75gmvmvMPahQotI6vGiZ/ay2DIXbC2zMBt2Uj2F1U2Tn4W+tW4JY9ke
FhnJ1D+aaKD/ZiVYcexmp9cDjbWfOcZTGG4rO2tptefbDMjfhGRSPeVfFg6wbJHgQBcoYSSV4L2s
U/vWDAryc7CJ+4q8wpi1hbV4pf61nDJTyxDcFOrKmjMEZ31v+mH2tcWgRaXMbhe1/CAAzGOH1PCA
1/cEqxesa53ZcxiYopwiUs76LDzqeKO8pdg5UfuQO1tpL4+8x6Xse5IZZ1t63M0tnmp/H/atop2Y
aSAhEjXfHqbmBKYKtg+k6/9ovfXbRWIqUBefsA7CHnDXdQqhQwOe2XzZAIpEd88GHrALap6OCGyh
6BDuP4FfiKOK8h1yq7x9N0X3xwK8c8yFjg8oO2E9xON8e4wl/h3ZbZ4NMtQiCKNi9THw4+YTdAmg
TI3fKlYbZl77gU2Ny6b19N2L9VVDKjQTOQa2SE/GsHAqmd7Jh1MACyRS/fXepvZu7UJXaVl8TsgI
FPOPcAQ9LfkZt7suj0/coqeK1JFwflFvpr1fJoLSOkyY/cMfJNrS/vQrJ9HZlXNS7RPevNTKMQxQ
lsERinXTtvmnQCwsdB6tIo1H+H4GbaEW/E+z0oKAYBHf6GnBIvMkfL0LmJDWCCERLb8ot+CEY9GM
H7UeJSCaaxX4FZHi5L3zYTQSXRDUs8YZzXvoqgZ+YWIfxhSBhBRuvqCne8IGqraK7yFbLNjddY7X
0zM0uhurDaViiWOvbY45yXFF0D3whzGt6wt7Jr0I7fcwa17seXPXQCJLFZwbkxLkFsNR1nTxBWdb
iQbChzNdx6jbNvLQ03Zc/xP9x0EKAe7/iSpzpfeqDe7KlYpL9dFeLQRXZDODVwjv+zAD+mXPOVhy
HpsXe2MHpgLsgM2Rn+pPJFJ+yjOUgl/6Iu9uuGTa/vQsK9Rgrg6AjPt7jmLVh+jeYhV9qhyLQ6zF
OWpAMzlgSVQAG5Cl2Q7dCMsVPJD5PU01WXsCLqgn9XYHeIlfbBRdhCsbmCeGdgVggucCwE30NC4B
q4fvTWwebEIC/Y3OyKGFzYVX/H+YSDIcxdPOOdFHqdj1U2UiygscXgCValob/vFNrJg+OMrMQggp
6f1JWqJT68XZOnU+TBtLcZwXmtkk2E5CQaKVB6PzSWK+JUyAPsqMOkuBNm5vgHfoqmhqK9K0sfQN
6Pf0mxxXcwYk6j4RgvNBZ+JxaeOQgbZ1NED4p3w5NnE48D44kBQLznQKtigjq2AHoais9MM/OzAP
XfbbOAeSey0/Q+sEJkWAG2LF4lICTe8psu2kdmhVOe2RtgTeQwVfC1K51Xb5MVTXeKkCauvuNEOE
7naU7yOlylV3S4cNgpejRZGZrEJpl0TmvPGbjhjktg+H0waRoJ8eXeZkObZkkdNWXq+jVgaBRJJN
C/q4k9UieLCyBkCLBrHjEyT24T6KwSQKaqU/YM2Lg6k5ikQWBP35oFJwlxV60dux7ySKw/7H/sFI
GfOXPiH81Yvs/cPZ4Lv679xxrVKWg0a5fzblq7xwVVyU+HexkC+BEu5InFPzXJBlUEgTVAdmUes7
FXOvDoXZRWIunnNvgP0iWQEZPpDItrFS7qJZ3SFEyVB3Cv4gSELXI3tdfPTa+wctsF8l30+cPcg2
CDsB11HHzq2cDvF7XnPjFtBs6AFTlmCZeM+Bsm+Yd9mDvthluAKtNP2WXxUkNzalemecBwmZUA1S
BN17SYIJbGTfKI1ExpypzfygX/dpc8lkY0BmSb720/3pXaIwKSO1yP7GJa9R5z9GQucslmSHiL6L
82EOHNSQFNOIzy+ZSwnFnQCtHSWz4xgC63XVpjST6Zjb2k4QjdwFFiXHUjB54v02EviopTCIybMc
37wzYrc1kAX6iha+wWsH4KEP6AKiJmBVVC87Mnw9ZwCJyZdmA4mGdZV6CnMfWTAlQ9+ppzqGK/di
UBTjKyvcHnmSJ1oZP6IRzejEh9DJjFvFlualoGzVZtpIb+xodC4xTll8gVK9MqxnQx/53yFRcutM
XdN4T5bNAXZyGHrZCG1EV/yZ4/urDQXvoDXWXsWE8gG6IJFwNzIExCyLgzCiXJDoZZKYSn9GWgRD
d0rShtTGBaqw0uCs7DQQGv3yxAMfZzzbUPk9EcFuPHmZBJlCBJ0rEA0qAQYG4R4DHASwquWT//P5
/FtUIvbelxooiXLGCTBdZRm8HSM9N6QXC8voUhqDyuppstiN8lTHafb8NbEoaCS3FZjDNTaVQA+t
D1rs0lWBnpN5oKSfqtZkQPQIbah363AFWxk9UtxhR1+G0T47GNgNUZq+pDmByTpURf6a7YjW6yYQ
RlyDn5He//AUdT5r258UruXxY9a4RhsauJrrh26m4ouvRwbZ1dH3qHkrceNwPFGIqH6NQCv7MpuY
sAijGPP2JpchKDTHDO7X4RzzX4aSc8Ao/wZ+/FLSmKWLjLt0cBuj2hcCwKjumv8DhOs8LrUPw9xe
QpoH5hsvu5x7y0D5wXPcwGnQj5UaR9UGxgcEkD96IUilGs3X4ljbpTLPDhbWSdbW5JftNgBFWz0D
6bQ8dV4NReb/ynxydsf6ANVg3MP/IdsbYRr0ej3xzeLzjXYhwo1hm4b5r5TBiqsCVpScc6utaC07
vVHNWwlHGTIeCh+xkp/EFt93TgVGeIsKNvQ0aJpLmhOVbxNwDcVAV0O65BSqik4bty21XfawY0ET
DvBsHI/wAaZTWMxSzJXcDc50mx3K55HJZGORqFOvuuizvddXWwLNS7FZo8yGF4XsN6yHHBiHLAKF
GKFbHb/KJSr70xErqsawIVLLTU6s6obFQ8KMKPPmeX1auRDSHOrO/PZJKWPMT+M4FBbh9J91J2Mw
73SrTD/wkLon0fkFxy0ZJ70213IeZqgOAAuv9rl8KawcpnZC3XYWbj+1pyfDctnKkMCJUCmgdlkw
7UdjXToDrbJ0XcX/VMFSdjqrQp6o+c0XKyrEM1UgLkVYPK7ogWOeHwKIFbdkXh9eeVLIa3Fu+v4X
pgjz/yqTj94nxyGo00ACbex5ehXlyEZZWTFHSyj4/Znbm/JAj3x/4Zv/U1PZXpKuaO8CcRlcfyFX
jHgGVYgpbggKQifoiy7BWmoC9F7FJGae86ANrHe4S8lWrSxbXd2LWx/0qtX63d6KR07YVUPrPPMj
xTGtod2e7JMGpynwZxN8u77HzlLFQ5JPrm556IP8iPSFva0sFpmtgm5KoY0XE/iTR4Giz8BEfOCh
iLQgPa7ykhoKPejIeGYRSNBVFuPcqwX5KG52ebZG9WugCz6kNA3qCIUT98IVCKappYsQvWTTzOUo
4wu+h8GloQjEl/L6FCbj7P+PttoJOHRM2r5xAZvYL6ss+oMtieTKxGv8ilO79E5//w/3oE+FF4nW
5MNADeujPHUcF3dH8igeVbKqIoOVDG7nNBz7G55Y+sfnpQNQw8IARcggVdZd5G0p2FiLQGdbnN9b
uMP4IahKmMri/Yz7IN/LON8lpL+YCAw4vQ34vq9Pv+ZO6AeTT+7tNvhkVZ1bhEZJwIwVZUB7JHJE
oClBswjz0i9IMDtYaTmHnNwQoqqc7T/RjkKeH7qf3BZJqUuTDmeI25QTIrxZYndIGQrImfLO3yGF
5qO0dnvd5vG8EBQUV1WRVMMCEf4KAz7Cz3t5pkNXyWZYNnhgMPotYvprRljs7xDN3GwB7Vi9IbvA
QUWx1OsMDyUIBEDUjePxRR6zE4SCJm5235Yw0PSln7XpbIGssGhyBP3Uqg+jGpkQXFSJsdJVYENI
IchiJW+kIDw+dRWZPWT9SfAU5xrIl3EUoAoRbraUN2npWJ8DiloSg+aQbZtRcNt+um9vN/uqrrrC
o7OzLjJVNhLbn21eTadmSLgnGZV6NBIa7KHg+Xv0wRfKzDHu5jbKnEneIg/RB9QMqVWBqdgVLA2N
IU+t9Yde5UwkXefvDLYtdVmKO7NigkVkhTtCbJFTmheJLv7kgbzI9cpocIJaZ376YqWZ3MS49kdJ
UyyZgNw08m7dsN80vn/8ga4ZPZpqjDIKQ9mMkD8fJziixggq9uKGP3yxohozgDqGpeGOIBXtoXhb
IAbz1rx+pMDTj94PiVdvShdrECtbVorJQ4dRqFPHVYupzJfQj5i5bKzZ7TXO5ePh/uHKxXgeOZNF
FxHOb6UqJscjAM2Lg9G0ArGzBtUdVdOWSB01C2YFkuCeeZIzpJJComJPKZwqZgT20aNqynWokf4S
1DJ/USqaZojkuBxYyMFmnmVkJwr+EWo0fCHJqcDmmQj2M9zjcWvu1nWMrDUZisyH4bXqeK//Ttwk
wjVoBJi28hy/GOWFq7JtnaZRfOlrJ5JwHmgTw3XiYd70KnkDgU07ImOGKKxKE7G7awE+aIA7J2Wp
iAAfUrD6UqGvC3bXKToWrfT1n1SM6uFqioInPpadcTdpw9EtQMTFJtrvrUA27MnPaQNUbXoKKiOG
o3pxLxNT2TJI6xjpGhutQKt6H1F1Pd/+FG/wu40C0sIluu5mHDmg2X1diuwzfn4kKr3pki2Qhg4U
+pIyR6uaCdFFolr3SIOPe97wfZH14Q605XDnK5bcv8k5rqZN2orF2cJ9L/JUv/1i56RuIIFHue6j
h5TVOKPOpl6t6++1iBlxSxaR3SKhyStjv6My1u8remJ75QrBktKD50Ag3T3D8gL4mSVRu3saDVDg
/S4AOUAYNoK59+0zHYmSMYxkm1Q7emLiCTbkH5IW2iAeW+ZEcWK8QuWPdR4E4jIvBx/2jbTAm/af
MpkOo1o7R4T8SHBSPeWhPpBuwn1Ac7VzayAAawZKYusy1TH8JYnP0H8Bo5Uj/BEkwkAjH8LLm88H
bbGy1ertZBlU5Xq68CvPmf3MDcwwgn+yaobEwTzepI4Mzyvle9f6gkZAZXmeFF0BxT/EEGwnNp+M
EhVYaYFJ29CEUM4b9/pJp0dxmvFl7FnL9VmrzNlIcHmgu/5fYl7nnkxIJRb5/UMgqCIPiMAOEnGs
nWfaFvZyuBEDN9j409NST/BeSBGhdTGSzTxZFs4dyyTem73ZwZ2IxMPdnVpsV4kmzvEHV+Yh12Ly
/LrO/Y/yVuxMczGytMJZ69w47P6TXUqlmj018vPw5YF7yj0Hvbz+DbrYi1pAnLWQjPOMpVStwSx0
PJdikgucClWnZo8tsEXu1X7sTrNm/dbCM9rqfekdtrMMOVlbg1/XBZP6ik+bMOpDtnFxIdW0f3qo
opUPMuW4az678ti3qfsA70uvBhTpI56TaZjaVTJrT3Jl+cVYWmQrFJ6+zDF4BffAWgpWAxt43Bod
p9pvb0qwwt96kG9k0qdZamQ41PAuTzmaBZrm/tyl6KLHf8Y4V+/as7go9xHioXtvSVoJKrT+4u7R
h/ToORDpgZoiWQBiaB78dvcmiXYf/AJ+qOPlrC3RkxXchlPr0NeDGx1ccaLJT2NEV9nBMGopx/PV
p1YIfRGPQ+cEXWFp+VaTFC8qCHcmk3HY5HzflGMYcUAZUH9NOezqSaYMMdDxLkFYcjhojZH8n5lq
5iFUHO8PBqOg9hiGH0IIZo2KGj0wVtVi33dkq/9XjBvKvhd0VyTxZdUJP1GdbpyqR2JXgSO5Uyyu
N/+R5SWzarPpGohp0yXqMFQzwrBWuoUIfohTHALgAUCy+w+IEV4eJv5cKQVQilDyRQkyY6N5XCjs
PoQkB1O705ye71q7F5WzRUqRkq2bG3298P+lqsJiXgB5l9zUsItR7b63h65kcSNJfhX8dWSbLzL7
xMnnnW/SiyizQvXsWVvxWjBHFwmi39B7rRds9iqK6e8TJL7IdK6AXQk9JGZLDADmo1u7Bmj9lhg+
gjsm+5WqS1xR/4b7CFwuNIF8wq1jGDkiarILxgrJqSd+8Hlgzte++mPodaZqHsv5eS9+4VvXBj87
8Ez5cAAsMx0DO1zOz+dAowFwVvQV7oVzeRU7vaAB671YC2X7chMvWQ6iqrK/3uyqEPTj+p5GIj8q
Lfm9EnByN0Hu740ezzJXRkkhC5Q0pzG/6yjBPCKRb92EPUSC5Q7cpfNmNBozdXjh6JqFw5l2y7iC
kC6b6u7kHaCnPxnGq1vxZ53ncTxHzuj4RW8T3fLMPavX87KTYm3QtPE51fkv/Cyo4E/M7cStfR8r
QhVf6NuORVj00fIgCIEUEqnf3PJrZWKqCmpxrupRHU8m4Uiv3QB7sZMnEyoTWa4RYxO6iklkPHgU
dnulZRb3+B70j2lJ0ON0ZFuUOMdUVzkj1j4YZaGlef+GtD1DMPHDlyGEZtgmcmfxxUYzWMbCBqaS
KDzUeCcHsPvCvQj3AeW/9wTD/qCAwRdUygT5i1IAgNRD7HoTHpogYIIikHYqAjWlAPg+kLM7/NFP
qmY6L2ExOEKhKPcBWO3Vs/XeqIVnaMBlVJoxy3skCzeNMOle0Kq49tnL9bI26U1dP7G/RT6KrjBA
0i8kY4L3Um1MYeWXze5UrxawVbY4AMMqtcdJZy10LULzejAp8xIzOyZ9C0SNv/8dz+5RrZLxrwOn
bV9DENZFYT1qYUYEF4Y9P6cEmCgG2MRZQ19jpYyCjV2s0Hm2659Jx9TqjJvU1gXiEv06b+szAkDC
/lfT9fYxWKs2/qT8nkL3z/A6UGdjX1xEJIyX3zJ74NqtiEqJvk5Qnd6GGb0wE8eW8lw89jeXCyy+
knbfD6Hn6XjNVsxH/FVMoUB+Vn02qEhLisEHCMfkfdQ+JovtGFmMTlHK0AMNe36a627y+wNPGi/G
S1yoCJdiKdZWYfYBXWLVVZDM8V/nykhRIUUdoPkGoTFABp/0ReMSWlXhqgYXcX9rYWjmwK2nkPtm
db6OhLufZqnRKS+XLokk/O0nINc6ItorgCE4bDCrBf2C3+a7daDCUjfd7i70NhjpFcTIkZcSpLsh
FGErm6mn/DXz2okhLk/HrghXSi69LLJ+6EFNz8yphdJMN4Si/o1Qhacz7uORj2z5EH09zoy63Bp9
cEqNkHr/kSBYuYL/sPUb8AiTtGurYICgY2Bk2jzHe9wkDyYp2cIrvBoUy6X8czJPpE0PV1Nki0dn
VcGs0VHZZVovkMykjl6zht5a+wF0gkBjNbMTIZ3HJsBmrpXnwFzpxQRCGRyGsLnRnEnbI8NFg7ou
UC1pFTupbXcnY8KmPzUPEByKxA8fWkspQgt4Wq0tnJEgNaxy7fWo/MfeBIFv37KkeFZWPTrMxMAH
i9a+ulOmhcxey5ZXQ7BsR7Xl/5oxuOKoNlyQGkEUCiq4s+PNVWMkGjUBM1ZG1ccmI4Mymkzc2z/y
UzEb7MRgq+3Db7BxmVla4cVlg57xohgyXrMMo8VTO0IX0xMcphJ8khts1gg7N7NJz89GGzV8PTqR
x4MoHiR0P1+ZRgMr/6YpQE6MIkoNfHefZGV0+yniOk1qKBnQB10nlmxB2zZIGC+dZcMII+Yq1U1n
JZNu/ZZmuKKWsUwna8WIoVpVNEjMwTchZqLmdLjMaOLsSAtGEy15Ho/xd0KlbgvCumJlxSEjIWu9
gJb0YaaIlVvdnEWkNCQLhQJeTEJ60Wc8dhzWvi8qb5gFYw+ZsyYrHvVnWVLfm8Thx4XbXuOTFI/A
0so8bS/BQRKr3wtHzDSWDQriTTQTJuR+cUXEmskDlXX7lNaPlQJjLKuG2eSJqoaq67tpc9YKMYMF
qW0FepbHGmifJufqbvv8MMUpCtTXs7YPwIxHPf/8NXfELV33ih/1HntrK16afgLKFASTX0RSq6Kb
OaMX8m5bGrMnMbLedPJFqph6qgoLDktoBvGolsjN0XI0mGdZDJx0J9+j375deIOnW5CDDVGad5el
GUyljA8m8BYBQSVoHHOdMAexx6P8z+aDw3PsbQLOz12okfGVPUBpHmd9JA0zT8Ebkz5dhpg8P77p
W2sgRM/D5bKHFXJ+5bm7hjkgZuFUBaeYEFuyizFRe2CjnjQbbBz6Pb1rvWuJjyWTevzo0MBseOaI
4Pwz3pR2T9nkFrnvPKnxSmZygxXyjoxvFr566aAYRtga4RAj4E3Z4WyhifQjipaL70wmJgzR5xp9
n/4uOdC6vOzfgfsvrqo0/krvbTKmEzeboSe/Rsg48mce+/Fqa2nUA9OfHXeBRBR/XZ0FjnmOuMit
q36HrswR5FT4yjnSobC3ZsqsLvenMfawvWrTiyEzdqwO8ZLsoO9kRB6NpLG9mRil9Z/zHXRrLWLH
bCiwtkwhUEIoY4ltBbDNr25/OcUF5L+R2CoJgabVwoEMvVoWeNpSwLSPbuerkssfLzcgkyot9PvK
FNAsqCRKd0bht8ScoQax2q3c84uivcr3lp5kzTFJYSyxQsxRTUV6Zo338P24dEBqDn8/B6Rjdsad
b8FNiGWGapTKDbsMmMMd5Y9JFiab5idh/xNnnq2cQDvNYLdtjGZgYKcayVJkYdN8R1yfAo/moS4m
w9tDo4FCoqi4dca3A2HmZM1VS0MT4UR6Hb8R14W6glrYqexbWFY5IwKCuixin88CsQa3yxYYEmHS
humh3TEEbxgTsTUmuPEj8e6vU8FJ7SIrCu96GQC86m/js6HhBZImCfK1PclS7PURjdDfaYapD9id
bUn5c5MlEJZwMVDKXYxso3paKM/pH7qNcHGGxcdqkVpMeN5ml3nxh23NHzKZTMDbjt7RWgblpIzk
pt8sQjCEI7lburNWwqnn1tMsKN8pwupZvPthEyNSxVHH37RCopGlmWUn3TjMsv6Lw2UbZ1jmwK7J
LHgo5eSaYxmw8WURDKobDnjm1W6dQYB9N9txrTlpgM54NoiGx0zAEQc7b8+YRSsYrfPCcGX2IvV3
yTiy0pKqhqA2vzXJgmlJtS81r4jOwsWZmrNIB83g7i+uWgTzg2bJfui2xzZsg/soneKzFp6KO4Oo
0z9Do6/yZPc903KcL86x9ZEaukA4LvynmmkM4Yztaw94wwvhN4zjZxbKRblgSyeVkEAFep5emRgU
2HY9qEwcJg11McBr2a15WyNOeV4ROHvYpocBwexgaXclWl/roYcNQQQT1JALA8uU6koQhCfVbTLm
weZGOQMJmpBr+74F0ecCwTwmXx8GyuozRZozjaEjFA4hdS9CDbcdxyBEg3b/RFPVIb4FFOSMptq/
xAGJCg7R3sEe70tNCM24G6ZTwPpauooEh+T/eO+LZgpb/SfFv1GB0IDhv/WD07tSwp3b9WpUJXLe
8uZkh1jfqg7UPM693w00XQ88cb17vz1/+O0pBi4WCM/erra9CVzCA9NtHIh7MJmXSnHWdEzItKo6
RkTzoBR3mhmlwGDMQNdF4ZYEnzM9+Onz3h9fepPKRmWMfdEWLZ4NdVxQfRxDEJ8oBJDgwSi0NbMs
aPfsVFe8i/Et7BB86Of3lIR5zOQ39gudW/rx5aDbsboWH2MZjhHcT9TH7BiQNdu0NTyi28jrCNs8
fYQuO2v9RW23LcsgoLOI3xB9u9EeThKHpZ0RatoR/4OsaeOQFCnCDTSrnJcqKEPr0O2oBhx14UAU
L+zg4moSNkfKGFTfWG7cuwFXc0EUVMf1H2OvRWZm42T2o6+hUDrqFXSOB4+MG8lWYY3JvIBUTdeg
lu4MVWAwMJRpxQ2I8h6Scp0tVRpFnsQL1bcBDy7TZr5FDTk24vXy9FxHheUGKLuoM6oD7xv8iL7w
Mb7T2y/wngT2COXsJecFfsT5HtdPhhSs+KU8N2Fq/QSV7hGmJupatLI+lipSp0Va6hIwifGO22AE
+mwA2jTO1iB3oSJTpj3zEUWGYLDEi3fyxALQA/bRFfE2Iy4992Y3fN1zLWWWoj4eHHxyhXdpwPwX
OtDRVb6mCdHRl7IXduR/UajMZ19aV2WrNG50CiA7vMnqU0ZtRe80gJ9ED7HWg4JBvCC0t96Hr3iw
2VkxZVcmVt4w6piQJa4hSgjxpJ0QzEibbPDngllUzrCjpEfyf91AOzrx6I+TJe5DihuOYf7aHqWZ
ImL3ufXDhvAtCc6kPOpVXb3xV9zVjd4CTkeAj1yi9nrwsHhUGzS73MmSp19tR0CF5uRfU3xQPVAk
eoUCdVCzEX10D9nLhM3ZfDRx8Bya7uvpKjwHxsDMm7vlyDyhcy0383E0qJJcElmF7dZDMTxsk7Vu
jD6sjRvdV7lAIEDrHQOd2UN0SO7kBHhFna48G3fBDATB2SE5xCSo9g7tGcZx9cEDGUlk99ckJNAH
w5X8fikHQPFMQaPPp/v0uyppW5ONB0Q427kcfxjiKpTTYrYra9woc3WqkO2cTYM1w7TcW0SHeuBo
6dB//Vp6/jHci4HLiV86/Fc5MgBVZQWnJGZ5DfJ9X69NJjabjxFN2tdBGAVjLqqSM7Bb7L3WiVsN
o8v19SZwO+xAvX3EBkNRFnQ3bwj83baXOuCiBrmk1v7mkx6qjkjSC3bXeldAP+o0IzcfK7VL5soo
9oF+yVgcopVrjgS2+JRQcAKU6HM7IOUWAlCqwKd9fCK8v9fx3OiQW5+Yh+21egkIdURv41WCR9y4
HIhxhm+6vCoMHE8XtkhRu9X0tzukZmZJ3n42aKEXDOdEgNn/KSb9++wKm1TpgBrzoXVGMhc/awuO
7AuceK56Al7ESABdxftkfwhz89j7fyqGbHFAz+0ULPSz2oBAhiD80Sp/UTYo9T2CYoGuj8+xo1Sn
EfUseZf+Lwoj8Hs01C+bi2PE8pC9+3a7vrXJv6krl7li+uCnego+Qu62G/bn6SpNgr3IDdsN/mPm
iFork6bmfaQvORsMOzEmYiaA69w3updqT721lOOJODOBnzHYVRdaPJn2YZm4yE6lO+2VXkfoHf7O
T/H+JFAYOXDMDvHxr3q8qEfSOO55biDki1no+a0850hJ9oCA0JUqb0tiUwmrn362EOW91YX0zR1+
ey/C7neDRwXY1tlO1bdPEp+x0pIR36dd5oUk5MzaJq1rd1cfb9nZVHFw52P4i/mLrZRloOCdnKxR
4EuEGvuRPPvsq4VntEGNOJ6xTNDElXuEqB9h52RIDJM8l2NRZjdHc6JHT4XV3iX9GeA/K6ngXA14
22ja5147G9ABKlzeGRWBCl6oA7VFMEaXBYYNV/C/dV1Q0I5uTpAKONYtxmJODGUjWtZFPV4ZjeF4
yCSLGhsHajtjo0RY8GuuuJBe3kdCpWcP4HGhs10dDMI7C4CtdnFrBEyCQ94ETiPGGdzsniqXIYsd
hJ6PRl3DOkRILkE0OUi5JZXp0XCgHVXTt45+ZphYyBYw47zSerqvK/Msju/miAA164YbOzcX3Tjx
WoJLVlzEDZXxlByqQl8gmTESRPGOfnAzvRUP2m6NnXJydOE/GzGVWwck1c9jeKoHsfB0OPXuRsm4
TaMUh5h5uR25jqXMnFNvhZS+qEshlDCMdqtpzUGLkFDEQZsWa/Lviz0NcVox2A46EkfHUrnngBCW
DbmFCD2UtiMEJtcQP18RZ/ryEz9iK0UX7Q4FY8TxR87hgJp9TqHnhSyR05Q92jl7BKl1ZLEvUA6h
h6tPhxRyESINg1uvSxtddyXwH+OUpIAqRJGrdCFSZKoG6N2aXOZNTO8oQ2WWf3hcFKR2Q9UT30ki
IyIQyg9nDSapilN3x5O3vtIJ/Kbx9xSRauOmwTgROS/QtsIHLRofZHmn/SFkQJ0f1+vbhMuRx+XY
vwOtqKTEWs6fWrGcOZwpH+GiI0LHZjEuZ60ZIaTHnQu1fNg5Czo1o/RdM/D4Ve6a9fMXYjQ/czrH
b/NvsjoFuQM6uiZCXunwum1CdtivuS6Eg39NXHxf+91Qjm2mCaSCxT3dftSX10Ezx8NHAsDivdsv
YXJMn8E4OetyqVEKR7RgI2j55D2Uw+zUgpyzwhxev4wafryMAAjEXpbNYJOgwc8LNheoyFlyZh2m
eBPs7lMa8MrDDvvg3w+aqio9XB8DDc4ezcVJ2Qdi7w50BpVY11lcrCN17ZE3mBNtCmqPxM1bMuM8
YlmBkqGUel+oyRNgryUHW8V5X2ssrGjDMoclkApUU5zoM5e030BaTaDOHtB9snhRNn1nd0MBa/+0
fJ9uDY/YW902h8YNrIxbuof41Eg+qKg6zlCfe/S7NF9LFUTN7bM6BId0XIlPBXAqggQcggmSgbaX
kF8tqlJRW2rpIM6EK3ocIkbRe4u1IoYgNWY2dIWJApYhbyV2T0VEjj9gfwhYyim2sx+CoG6O7tkX
a3LyH4q449ghVrKcoWXetGdjleCW5qqgsv7NhriCB/VeYNmJtqCm+rqsCQ7mgQ4mR8zHh+HxUq9Z
dmqECyIYhhHZJF8kN8MPjZYrSTBKDeIv1CyP6fwxgdZLIpETLabYnUwLOPpDbAXBuApHl9b0Ooki
EmCW9f7/MlQHR8jNpoYVAQmqT2inOaGZc9o6DTZg2TzLhuPl8jjFAqt6fGN/HzwlhO4JdM3Jn3b/
6om13keflPEsU07XZfotVxOT6Azg0LTSKg73lXrwl6WhKnorQ76hb77M3+6eJeMyCIjMuIyWxDIf
WvNlzpxvjRNccWyd3DO3G50/D78YlP062WNn4zgpf8cU0p3wAzj03vxBxPvh3qRbpRSi+Pg+93W4
a8hLwgAbph8Hut8yI8nJNV0iF3bjqEfHtesSVPbdYTqAZOzIfYgSG3r5Y7o+lDxSMv2TV7dg6rPM
9VOVqGFL97tpMuA1O40kixvZOKeSscHKSZ3ISbXd9yUjMPYW3omPXg7jKgQL5Dorp2CjBhP+6h3/
ZzYHZKU4JQlrdvnr4akmco0kAJWnY/S7vWkDevq4Ofexd+sSPCqZf2Mr47sj7mXt9YfkSJXT4j3E
L+u78l2J9GxgNsDFf+G5j7UDPcpEkM/mK0lSNLiuYw7RqT8vdORenRYI4jErNu1xzEhjOANqgAWD
unsK1Ox2cONKbifhxPlp0a4jVG92h78O4R3M158vFGAI+l54d88g5laLY35Ap8ZtUQMEkTBREYOv
W4MLnba/2VP91I6cJd6Qqz7qA2zeoZvtD2vGWQ9usbw3VuwTTDwIkl44bBfjVCAdpWzpFChd0In+
OEUSerkahoPqZlqUzaBrlmhD0EyCdJpv32rFK6RozZermXBtHrciD3fayLkb4PooktSdWsVrD7se
RdajDi78OIwdv/sjnk4yxvgW3YAVH1lxtY/pFXUlz4egis5W/hucNfbtkzYHc6DsrT+W1dg5hiGp
bfVYtry7rs/NbBqF7trHwRqyEd+mkARvX1EP27u5ZE6torM2yOq9wHduDWvfHeKq/epnhkSMtkeC
Ava5VIuy3l5AE2u7GHqB5Ru3CdVLBGafh497jWJKh9l3RMroAwpAsYxMG3FYRL+dSYH2UI6viEgP
dg6ZsBmpBs4sx3dGWCAyEgYiWBs73UXVEmUgzRGKubDJCG4fs2UJRLC70UNG4rJNM+BmAfgtAL+I
hTvV6gh1bfbzrghgEE5Jaj8pmPboh0f2aAivTSlmmlMbk2decD2GbYpXlDfrtOJ+2/NGFAcobX/A
9KP+u+EOtThSczjKAu9iCdc07Ytup/DhuA6eMxAzFWRpHCctNmnexqufWQpoFJX330/BtLIXVEgl
U+iS/E+rye/gRevLSb4MVkpshMc6N3DIheYJctW0/v25Ph7DRuq6b4l8GPZbYeV8Abc9/wytI0/O
gQRL1iiVJOVT8r1froXIkc3WHRnSsJRfb3UQSV1kMfjno+X0BnFG6l+sFFGNzfHtVEjOF+1KUpui
PfP3ltFTDHf5fqKxZVfOHzrBnb2xQ+VgGzZWcofGGJX6BgjpzQ8EOJ9sFxJP66H3dzMzTPJV8X5W
u5zRC16w5sVzNcBD/hwIs0IMmPICS6MdVUfjKo0iJihNcRs51OIBW3dsQkTKX1ufZEdN1WSzjhpz
QMFRvJdggfvdUaPg+zb2w3hH4Sf2bCP5+AAX7HCXamc7UgxeljPokYe4buRynGx8FM/ROyYHNWEo
zREEqKQ6NrQjOSbgZRSPzXdEvDm6syR6A4hEINhdcpL7Fgl7ImJtlc5UqDntmQapNJmHIHF/dkqx
h+NWyAqWb5hMpuOhtvamFakngVFQyc8Ihyzf93Fa7RePQOb1zOQJIW2m+eTdFdprLRr3Lw6vKJng
thoGnIY+3p6CyQoJLGbX1UflVn3DlPFg159QNG2yo+er9MHqhcW9OBrYCggSlQx1AdDnmDugNgs5
X5vz5awZxQWr4Tva/9ILWbbUKVee4pmRpkKBnlCX1gVy+1bnbUOFILAci4dl3ilQRN00HsSXuXG1
VFJmQnFn493q8EolzZbkgiOyi4JeI//qfzhOr9XsbhHYEvwHCUqvZeh7+IMbqgtXCC9D0xmh/7U7
QMO18oEHohKV71gHLwltVPJCS2Pb/VVEYNwC/9143IED3ZMJYnJkTYZqjkciYrrRhahfRbCpyhhG
b+aCvYwvUMjYy6qcy94NCL62drs+fJfE2vYom1jFuyUMSs4/9TiIMqO1aJxc6rBn6Taa9+3IpxlE
eQWjRculUGY4Rdd1kdFh37t35EHWw9iz6MMaos+SAUEbEyLrbcQfTAKABo34EalQxvM+qTHIklZl
OgwIC8jVcj4tx8fIjiAzETSPP/A0cpWEvHy0OCAMZLICHeoydXaUV9fYV+1RE1cbJzz9Mkcxj61M
+rbnCRhq8kB9OxhI3JE0vJN314rpdGjIen9k7L/GuKqiKQgC6ubIojuqdAu4b45tRQurG2cif+X9
6CTk/NVpMRJ17wZtwKx+46XBFBjL3eQah8fUDC3KHCPreAQdqlaR7MmNx/g8Ai+paVUWbsI4421G
vWSpeh/6ahttW1MWZUIheNjRjAsIrsY+cQHauMgYBD51m3hTOkfzwQ5Pgl9KhqcjtUea/5Wbw5Zw
4ZVzl8LqQy14SVnAvEKSdF5zFQQrxvErsOZEzt6i8BZpp0Cf16JTfaG8IWbUF+lrklNaCYUq26GL
QSQIojWsgwdwav23FwWHxgXKCNHb0GnQXtlTo+NQ6ScttDtsu5usgb3VIcRzLNKD0F2qAAgM+pp1
Q9A3CpT/kDpJwsMwDdmrA++FQ38q9Py72QYfmJJnBZUwQEs6MHlA4V1+jnws/8mX+lsgaYBsgMfB
GQYMPeswlKsNlo9q5unqo3p5ogGF15VR0kEJSpO5RCOunTBBkQKDRZMQVrUeujOJVriGLK46hmpe
EsAQ47WMqws9mg9t7d08BnnciRdBXFZG26+Fd9gGJ2+utRNv91asuQyroQpzMOJRU4g4oP62Az7R
YAMPSnpLuB6hb15Wi8KU0E4OwOuLBsc50BTSjmj9jT83jldZoJt3q0JKvKLgVYE7Qtl3yBuwthae
Iq7xU903EbykgrtGxMROPsxw33Jj5NMjX3nGTXeFzoQSB6xrBLg5WP2HzU3G+TXDq4hjyMTuBuBO
K/h2DW1S5XF97SWiCOSDRhwxfNkfbK9rjW0C0EqMkI/PHIwFhCHpmuJQ+egziSJB9B8roGQ5xMS+
Q2iCRTMj9MnB+nHnM2pyzCk4BrU8D16G0hW94X3yaJ6Xm7F0UliPgbC+KuLP2C7L9UYe8SADf8L1
VI7paL7ERjUx+5VKqhdKcXu2aOn3um6aDDFqobHGn+UnEd379BwYY1YrVamS+sBxb4O28qlKMEZx
0m3yZny9UQomju1e6dm1FLQXgyFPdp+OZbGh5M5IaocwcPMzVx0qkmBqLvWm1FLI3FHAHO/jtgsZ
J04apU+7sRNIeFn8UFwl+tvYAB4U5+khk36u7iN6+K0AHEY8yL4z0uFLE1eRNtubuXq8k2ZfVVf3
HGLThJuT4B72AvCPVV571kd80fbMLl9r8YsdIrNOFWCzHVscA4oU3Pq5KtiInOGLD4R71I1RIpOW
HhOGRe1upHtzabsE2XCZ7qyTJ33x/YlbPZh5vPMbwGcPGzjhWxlHrNph57iO08/1NUT1tm5TreGh
ll3wK7C7XKAAv7MHeqWUzXXkuNABDUmcGaJ5u87p7BprH3/l565is4UKAsn2Fm5lnn4bNM7hHnt+
ttHnLMxl2G1eiOpdojZNu8H56KJm0SChK8RkVSSGHhPr/6t3UzuJxHf7I41fTnGKAcYr6XimcP4C
VLCZ+xKmo0Yz8DfmE+Z3QNLMgXR9HnVcROV0KbHsphHPzFstmvU03zhFxiS0xzbfmbwFzRcILPvO
qw3XSRf4bk74cZ5D7uzBBnDGhxm+T1wf0fdsaGGEXmOCZ1oaTW6YEzLrROHyYChwPdax3IJ/yvhW
5ioPJSfCByZS0Dn+TSOB+uVUF2BCaJ36oFs/ByAgqX44HTbL9GH4T34LR1eT4tm3HaCFF8CRtvq1
JrRMBSGSQPg1F7x1tazK7KJXlJ+ZaRlZd9v2knzBM8SPZ3BBi7vfJagOmHhQXguK2xXOedRKXAVz
RedXAVyeaOlf7e55sP8/RbkZfF56YaAjEcn+s5u9ePTl+Rp+3mFmE7rVfI8/Utvf3LboeEnzO8yi
fEcjSaoacBStVi6EtTPN98KnVZ/4QDxxXuE7n+EZCWdrN8d2EwmvcwZXJmZ5JE4nRBVAiMqWqIrS
66GEkHHovGD6HT+9xD/oL+MFByapboPeb2mOeBYnePDqR3wLwgkwy1/DsLDi89cY3DqlaHVhCntU
99XXpEf43I+Zbykip2C3pgCCjex86JWLZuLobp0MsodlDm7C8iqIUkjhgujb99Tvkgm0sfBbuBHI
Sbg26e7U+YD4G7tVMqpOu2UFin62Q1xxm4VGK17B1VVztj1MObtiw2qbzS8DOy2YnqaQIsm0F0xV
9WaUD5PbsKZUS4EsNMnQigh9SmlTcRETP2KTLiaSwSY3wiy2aLemmXSDz2TuQpToDNa8YpHMJW7b
U1njYQSPP41s/l+LV20zx0rq9nSRw2R6i704uHWQVVeOfGpn+F2ytnCbIv5KBddZuzSX+00qTmoh
jAtZK5aFaOxL1GTNemnj39yIDT9fEhjvKd1LIuOtr8evLdG+JVPY17urfpH+E5hxPOeW25kiCYAE
l4IPwFydBMNAMR4qkJZejlaKuBTNOMN/a6+gTCPJOBPh4NPEGAkiNhG4tk4P3tkIweUUtFHlhIbh
abD5/xr4tJOInAUpZLzcylJpFc3sBshmfCRvfV/Jhc0g+gyJr81DIrl0BmL5pjA+LbwXT+bmaZ0q
vut6kxQHp9eLLcEMhJXLQYvorRhZaFQRG8xY64GFHLFeAiRnF7Qu1ceY2e0Tee0Lq01G8tlEEO2N
VaTB2FAkuD9KiBaZoAJ/YsssSBJ8wg91quqWjeX3OhFEpVc2Kn5o92kY/nZUhUvn6M/s+aTyONuA
PJoQpnfkicKeMIbS0ErklzBZPEBfPiNlax8EnM8vO/0ujCsv+ylU5ffacdKlZZOUi0/P3BLoe227
GqBTgWtCvibZVH6a9r/Ymwq92ejJx2fWsovbnwjjxW+X59TmNhWkSvzB2dufdfg2pKRdlj+YnRUu
lYAfi5hwgshHX7Y3SBoE2j9JwB330Id1j6yoxVoFgOycqmh+bjWlaPEdH+2T+/6QkOjRVoFrWlH5
xSbBz4uZhnjTqb8BLDSuPJrBpK3oH7P76nlFVZ8MVWGU+l+jsPJliMzJHUn8WUrLhIq+3ZAp/r5v
zbkz3aQJ7N6aOhPFnLM/YA5z2uoJcxCpFmeAX/kLdlRZ2lNz0ak3sd2AjOF93DFVt0DncmbbX8B/
+EO5/8xD7cV4IBQnXikCpVR9FofnoUNo9vcdG9xqB1FSENMvrRmCkCh3a2ExgLAgSLp2rhaYmH9W
pxI42cho4qHHbSuQcsV8zoPlXSpldK7WwTPfvdawiVz9r/n0zJ33yok5tjiZfhRalmBUeJUseV+R
VZCZvJ/TYjfGCL03wpuTS9gZ2vZK5kQ48Wsf9m28LKnR3PXQ6s+BCjhYH/trJEqH85ue8GaT+4WK
kUFSD4kHb1y5dMpqUTfaAjb/ziQTOLNs7GzsTDFjYUDxEllzBNVVEcJlQHN2KK9TnjzDU4zW4YJJ
19xZBDrog8gfYCoa7ep0tOiq/Th4uXZDpUPdUe7Sh3hLrMAXRSQUcKpiaQwPq8MEVImVRkJdZNi4
jR/XaLLbd/xkrKSKcy9pyMaTqi62XRyCloiGWrB5bIFkMsLI0H04cfSH2QRfYuy3zoCXButjaE98
ajigMIlKt+ljhDYivpaCPSMK/ZjnwFAsTR3rEO/EDCM3oEAqCKL9hxa2BO3CvIuptLqHXQCBJaLP
uTrFaG6bjI28uKRQzmCWIdOsqS/9hhJoxeNkTq5rsNU8BVjQzP/zPBsQN/M3CR2uULuO/EH8aNNt
dH1/RGayHkuY7wR9ykugLSQoPnSpw77kLlo7sFewcTSRoIGgM1+i9CC9+pifbgN6CTs4wB947AIN
s1iZE3egLlv2qYtbs+1bf6CKWIURSxsrszshBORo5wRVSSntS76by1GglhEQP/wPN2msvQRN0nrf
l9SFDPt6fnkJp82AD20746L7qSK9hLTJHxDtv2qNMBTEKhpJUzGAZ3JLuKjJ5g7hFkWox5hsf6lM
LQa0McQIgMMPDTk8uYlVxXfEoaeMF9vvE0y++akTBCnQnDsqzu1MKpt+LDhk7HiZLhdbiBY4qZod
8e5NxmxPFJmsOtkkeIDJktefQLv8WzU06JS5I5w5SW2osQDM2BeH6qAIf/ZK4yzRet3XROTdZKXC
zjYfg+pWvzAzWo+Vxa5kFzb01r2pox7AXSQwZg2GqbcNna7uYxEIHntYO45mXgG+AmG+8Y2scaxb
2W2qgIS+7baQwmlQ9bImedhHwvoBJzSsxUqggXZ8w0JqffsdNCC8vy37zxQekEFcMOk4RVJOIs0r
Pt7wvyKAN/8CO6qF8RtyBHBcKXnb4YOO7K5dR+IZR48Vw3oWboDTg5vpGfiiTvkJN4SmgtLcFAWk
6FBQtluHiy+D931HEg1b5CY+6bkESEgIh7QDidyKtSSR0ol6WS1xBzpqTtFd1uTv/FLj4lC1WdoK
kMdx642g9Rwn404FtD0FGzOLcawpJHhgW2sHq6mjcCzybDx0CWPKnrY9QfCfHVdrL03U7dAX1947
59Aqv3QZyZQ/jH4R07QthP4Shxj70nkQYW2uOIuBfx/lZ7Dmc2rpVQfk0Wx0m+GK141eRduHBVaW
xZOrLwbXb7QihWsg7jYj/WJw3kPeOuco00qtaMyhb+Qy/rX23P+9YcrR+5XgnLrJukUZZ3DN3MUt
0aTam1vvj9LMxcQ8BFmTI4dng8ogYARYnwwLF/m+6l2qeQiGsg4LD9ObW6aOam3O7cDCGMFe3CQh
FQfYuTAtE5QaOS2IHuboEQlOeyeQcIYagx3ACbFSJvKGp3cPLBpsqeW2DKg27JZrwmn3oqef19P7
aLfXSh73qo91JPLsvBgmsbvvFBMunFQC8n0s8rwBo3IOtJWDWFGh0E/lLH7Dw5g99qL9PVCkJMJn
TB8+DNdnR2hog9db5r7Y2JsYctAlej2NXBoJaF/OS3hNQu5ge17ItAy///EeJv+U2EULuvaRnx3P
fjt+IZwtz5FyAfJWY+FSJZxUcUGCPRiz9if2klx1YYXFKjVm+TJ4A/gB4/14dadyT4rktTdsKuHn
IX/OB/QXDwH+e8cAG0cCJlWRUkMVojF8No58LEuies1zQJvTP1uwVd8+NaQ/Wkl6LjUhDj9iOcxJ
uwo8CgJKATeFHPpgChV/CikP2Xzb9z5gab51b8BcM075xnrtodOtc9FW8Efke9sIlwwlXitFypMu
ot9PHdYdU40QamZ1TN9I8ei15VzP5IAJd+Z4T9vOq99Wn5veP4LZsx2leSze8/wNd+CbvOO8eL48
A1ctTUCuw3kihcxD/ya0YkhFQIx5IpkAwoHNrhYtAZIZ9AlZ8qEbzaus6pQA7QgxhYyX+uZOY//d
aoZRxTfQ6wbUYAuyaAjn1C/TD5yFGcJniWMxnZtVIwbPzhSSO0lOkKTXE66zoUNvBpFXQx77dL3u
2CkwB4UETa8xsKYag8XDQEZaXHKd433xN03QgFuns23msBDYwk8kyiFR4tYY98SlZocKbxi+0Itz
+0lPL9chkg2M1u41zmlOmTu3IGH3wOXhr8JYfcm+IZDUa8RaHbtlP9XdhG+TlMcsib+dBwGau8d5
sp0/AaGF9kztwbIBWDxqR9mepb6JZSBeUZOhjc++WeeGaU5KaQJDxQBALG+zZU7etTP5i1vJ05Ro
MKpSz18Yh2lRO5QyL+y8TneAmGju+8oTUHLPNcQCr1gmxOyBqsi5YTheNOhpD77UHAjLpyGfO1Hh
/f/3LaQ7mIhMuQNd6UpLYqNoeDFq34QTmfji2PMPFAd0/6zRRwInVo7iRMP3U/xEbMIpMEE4HtuQ
L2vSm1MeURktUx9w976ai1upv+vm6P1wCevRiocXB9MImNCnYTcwKA8mdtXkNyTFhnqr+5z29f/4
hSuWmC3iPXxq9VvYeWT55310YhZ7qc6NI4u98SDSeKHviAx/8i3fKKVaCvgKBTuCzzQixiXvaqJB
4l5Kp3Fc0HldxcxUeqmkVvYp9CR8sWEoRhdqbJ/NU9lrsgo38QlPNQEinQ03MCFSG/0qJk94iO8P
mc5gjfj3kL+4nofNuFTlrP73sSocz7nHqHOC9NT5gvOaQAO96laqnqal9AfaW+BCMEZ1hVox1IL0
z+IaOf11QelCXOyKcsIVu24HiPIhabinyMYhUjgoAzCnsEZuctcB5wOPkUGATdWiC1OTUzA6k0CK
ER4z6fozyW39JzzNA41eyL3ip90QKGWtztp6+kFb/ceUHI8y41MsHZQwbJi4dwST3OZtFUOJwfb/
rlRnwDRedGgUPrb5Emg1xsfQPACiwZfJAVd2+T1c/rvu5tgDGF5g/6D6Xg5LmOIz4bDOLroggPn7
qQYZvxjso118ImQVPJtrPl6dPG7RQDIzk9VLcv20/aooAiBiRLek0LwErZW3LSXOugGyGU4EJifD
3ZLFR/crAIAuMy/MeO3Wf6FwRZ2tHrdPo6T/tx81Afkbb+AJt+cX4FaImPbTHJCAFU9EQIgGxsXa
fCCSDvFra+YctyS4ctLJqs2WS8qS0dR1hyengk2lIPz7kUO1YMwpzZRTMFK3ckZoEem5bVSSyauO
LbtMBgkLP6tGp9zSpssi6c+8nsgUJfx2uNPdpOGTJgHW3OO9wVQiHNtVlFtJEtobf9RZgVSTl+qM
okztwMi/+zGOovS6pt7XjzTtuH8MOtZCmzfcX18JMKgRvQ07Isbjj1gVcPq3OKWG8nwIq5ApjS5a
NJLAjKkxAW0XPesU/6P6vKd8vQB8+/9kXSUrcnpkfPTrGg1s/+M3KJBTp9nwRf2DZQpq7FdQcD/G
7b+LKQJLbiuv+Qi8N9jt+4764X0/beIEgbvYr/EZwUb8a1uvMpvm4LhbrwZG+BIq34wN9zqU0Ean
QrTKmehyFFSD8vpEhPcHRzDL5jkEh5C3t2WF238p1DuCyDw2ytna6RcuEqjw5Go4tR6OC+wbAQeo
Vw/1fe6QX/x+/oE1ZDShxLlvOssnvof/ip6Jwu8u/mT98Y+KI0y2qsKazMYueV/cf8R3ELkzKPm9
Pn+u7eQ8dAFHUswB7YXnWuv8kLuUXXOlXdPYI0BKPXUmhtuZ7XGmUrEFNuvxAA+2WsMjRid7zmbc
GiKMUoWUu8QbNUfFGFafXO+LmU5gNKi07GE0buxfapeNYbBhvOy/1R/gTQNz7IyxXmf5ANdykYo5
BUeC9scS4Dbg3ZFmlk7hby8ZUx2umhPQtRluNvfPvRHdQ59mqkctEtGSaMeVevLKHOlGM3Xh8eJ+
XK6gfrxk/7tKaEnKleQ5EiOKX4AU9W4BCfe3rWyz0irrzkveWKMGsxGbAp2wzucd9m3o1GDBXWRo
JPuhYEafqdm30j4ZU3meKuv4+ZoBvtKwzjCapkmhCBFhA58CTV9Mr7nFRYUsRwTm9Xolnnc/wOKs
G3ngcZdW9TLRtdIeoL4XUkzi0ccOw4i39jwUAMoqQ/boBY21u6iCuK/BDu27iLOJ9oFS7d7S5szE
KGWH2gCeVAVkNTk2sXE4psY1jvYEfSFPlsq+NS2Cdryqr20tMwGrjGMRxQP1ZoF39WkdqpE3Y9v6
gd8XgpPT7+Z/N2aCWuql/EV3EXGpLCYfkfJXR1aHpsj3Cq7UGGDbKDtLjdDY5C4JbQH2GUYI6d2e
Om8HRuOJSQCerTWFtS86nqvbu9jb8dleGSMP4OUgCZ/+MQ3yOVOfZVO5lbdNIqscfqDHf4f7Zw+/
QqvjWWn5wS1T1poVhFkoLNK65snFm6xVq5Ug1Z1VyhJPluhGDxfZAj9TbqmrLy1fdMuMBjhEJWYg
5ujat76lvBzi4SOduOyoSPgENDstCUWAwEitthEdNmODJadspyWUxjfaV+InH7ZM82zSxA+Y0XON
AYMuBnoNtK/jpjDqjoPm8q9FErb2+Q7mTUhEfMjttdnICe4nWdmXLqDsSpRtPPkOa/u+3NadUJX9
3xnhubRjPSZcCLYBMmkRaqufJAOkebzLMh3NkDCX9w6VWwJqXaazWUmq4xZpO6zt/Sm1T5iq6FFp
LfgXSLOT/uPWSrpq0Fw9Xlx/rntdrWiYTHy91lIPbNzuizBv+yIOsqKv8pGzD4vSb4IG92bCV6cg
GwR60b0EueiNW3k1dXXLMzcEXV6/3Sbu6q5AXGRtEqad3Ce1mNy7QrfnY3+01p30/7SI4njMGZs9
c1nwLGJ3n8lbeH+ue1+LVgAHeZbCkK7sP2TdyA2sp6a6iW5KgHYqFvheDG0+eZ10NUcGmg63QvvX
fI4KEg8mHFYu9D8GXjHAfM1d4L2mVU8Isc0KESPPyCdiKCH1aQTXUMIo7oFaBt6+yaUek3M2UahX
cM290yCSfR9lpTMvvVn5zVIoNjrQt2pxlak1B+HJE2BiEzp3phy3foGeWyN+tDKimjRY5niHD+2q
syNP82WS71p2o3lJnC6v2BCXZsd432hv+s2fCa2+p55fRisKGR2F4zApH2j1jE3+qd/97Whlfvw2
38Sr2dBk3gKDRMqW0SRGaCLaldMKXlrCsABI1gRhvSrikAisK7Otw1N7WgGYFUuwZyD0kJtLutDJ
rRpUD2e2qsfyAtdiJVm4RXeAzo2H4gV9Ss3MPWlxnplbfF6lwNyUC2315WNhj4STSs/R7TRJMe0G
y+ti4qL4zh44sqLBzx3O4UI5okILdsnk5tI8HGVCp2kg17h6fRCmi3rTZ45qu2ECSJjKfFQdXwRl
zp9LXGKpzkHC/EZxrfvDIERJGyKvIgcL+HfdrQwPU37rE3IJueuExwpuQZg+YYMZA7Sqz0IN3zI/
2IiOBaoKttv4AGtEGdST9N9xIvuKDIqWua++51bZ1dltBW3ctcnM9MfX7+Cz5TpmyD7suyvYuK15
yaM5tTXN1SB4LIgqtUYruDXQKINYbQWTUnjk7zaslWXs/5BKhW7hC2NVI+M9ghheZH5R46+9nmfT
oBCHVUYKEXRg8tFJCGNrxa1gOrhRdgh9qmJzyr6TcWoxhc4sDtlDEiIF0nTWSPYsKa37HCudhwl/
8yOhk7pbvqiEZJhZcpKYPfdPcpN89qS++ImJFVJN78+GfdyNHJaUPyN22wy0PlJtcxW7iLXyOso7
e6Vl4q7YQT6puDHD7Xu6v1fiNcDG8yO/Wp4K5p42nM5lebkICKHvZ4TvY5gXEk1ajEQyLPeItLbU
qaozeYbI/A39W3eeTAFYkrIlyemHsShHXC9zYveU5NnttSyBhttFR4XudeJIacwiuG22A+y1EFde
HWFFlCVmmOj/5GRCAeQV94S0tzh9RYagmCuVu49nVAUXJlAMgoHlTj6H/Ijmbw4oKaS5cBDP04N9
C8AUcq2W2GHGmwpfMVDBY0VJITssdUIT+s4Mlq/3vCj1dbljz4aTxaPDk6XRt/WysOSClG/t1RDI
kkzjWmOJ7Gb4+GsaEE6F8llNrZWZ/H9RRNGeVFtbwxXXqaOaZU65L7v31HjUsYzy5D4ow/hUD8ua
RQXvb0FmOpbaF6s5YZLWxdQnePp9ZuGOzfl47QIU1lvuU3i1T7XbVS6GWtWCjEjXK5ekL72t2N3s
cjwfl3oXP3HDOUrcnRw+KCiOapAkh9vqbXvaZR0jhWPFln+cC0luuTwUxprWQQSG33o0QRgABP2J
oZO5KJFNhwSXElhuYlMO6MjQrHqSoddt6+OhaZLlxXYdoU8tn5+kUN9zAC5wn/61DiHkha+ma/UJ
9q3Jm6GMhfRHgb9lvFDmMRpG+2i/2n+Zf5S6ELwUj1UzIHTbebd+HaoYwMAChy/yqW+VmKc8cvzB
iD1NCDXwOjjCQZVl91d86iPN7HCPHRYz4nS4WrBm+aYvtywY4pVD2/30kgp8F4oQ+g/Lj1rz5x7R
FifToJ4lEZkfTTGOUMDyHW4y1MkvUwaJTOyRpbzp92gXimKi7bWHGJ+7Ydwqt6meh79jSRY8JLwP
VVWHQRJjRxlekWUqmGhAgUuK335avgSHX03VakBaurm2iTZmgIvpNfT4ah09kIa7gNgFllibOHYL
u/uLNuxa6AqkLqIa9G4XlOC/7R+huD8V25RkK9a06I3wlQ9z8V17kGie6X/EeH1RJCzt+j0tw92x
MUyPjM8lG2IUqaarEae0I1n9bGa2Zzpezdy2ExnVAQ9b/ZOHETBqZSfSYKW5XU5ofGKTK2mt/XsO
hKBNbbQmh3R5HlNSf6ZohqunWi3WKUVudIpZmMr0JlclTXAPO0gWyvYmFWLGeNqobbOzT3TWLl4P
HDN8KVn/kBeFMV6MhoruYJHAyl+E5pXm9Gkt4hTv9qLsdP3lMGiT9rzeVt2scma4sbtQsUTXvQ8v
IXFmp1+si7Sy0Bl5JYD6DBGlysAuTfmhHW+TXbI7k40MNIifDjywDnvgU6gaQiHZI5Tw5OV/IoV6
0vlQAqN2jLLxu5QdAu0p26tcI0iRuTuF3ULC5r97MTvHWDpn6P6sh2rRUCq5YKfRjaxammThgp1d
puf+dP1Z1ENXGMqcF/lylNLv+qseqXqmraXdbTHjAE1UEGlZadJA0BarCkkX9e7kevyAedhg3Lla
U73dng3LezQrYuzMk7esELFU0E5nB0NXCNluith/Suq9BH79cdp/bbA49raTyO4/WmOgFee85+1+
7X8Ausz6uwkiKqGVvAi1XEuXzvliikoTm9jxX1VVThcUSt96UQFfq+aPdWM3Ez4oQ/QgIEz95Jay
0TJj0L8mLkuJiIk2awriHOVdICbVWRBqdJBbAA6CXq5GgAoJMSZCkhGRyGcqvCpR+tHbF3+y9gNu
pk+spmCG3hFEOGaB57ZtpvCx63wBt2Axa0LyCaKpM3kz1tcWPq/gJICtWP//H0Lz5B68a4BClHYV
8WOw8O1T80zLeBDbaMF0dDiqfAZbQhgbDwRCYUQMdQlgvrmHZzXIXylrvxRDTQ23HptLi72nI1vq
h2zQEZGa59ebLbwtSeaagRt/bgY0zGMSEP1u02n65LIgh8aiXoOZbrwhG5LJSnI4JfMHewiyus2N
EwFlDTvBxgs5C68coWhVNMOEBdbedj/ZLJetdj/nLNCJOH82gL+oilYGR+tnH6uzW+Ao7gWpw4iC
P/nJxVkrkOnc2c5hnj6W2sfwpO4vd1BpMCSQcWannBDuRqTddOctaMBvbsmzLiKKbBeuqogDIA8g
jEEcjmYMLwRarrHaGL4JqAiyzaayS7KYzRtskfAR3RvKZrfIOZM+6jk9OeyXHbgJTjQgYwMCa2yq
dZ4uM4PhbFcnDuudye2zNNEI5ovGwODuaF+Nuzdmsm65XcyymO3xOcnMQjpgz4J7Gh6VdwymTywe
UPb47tnh6w3dY3a4OO2O/yKnwomhPbfkZUeVUpCU3hehJrNvYHEiJiUEPOitqHt0zG8yoC1wyLyy
zcHuKufpHvmEVmUBAX9lJxqzgglgKjTqGe9+c7JDsiwKCpMNh6YaGvLltIN9hWcC4ryzLq/K2Gde
oOr0i/CmegKMuBTyoOnk2qGnr9vyRotUKPTyMlbarTUklAtDQ0hvZY878cy98vIprIxnRjBA3i8V
TZrKxsOUlf0sP/Li3/cVfWMAYEL5n02YwmkJePuZR+8c+Hyv9ooA/PzvUcbJCefRj5wumHe/CpR1
mWpmi9EOH9uP6lZ3swEro+7eP/cLrYtDfLLahLkwmkfJWF4wPZJF2ne5xJsElY+AP2mJa9nv0MlL
OFWTCAl+RDPCBbhY7wPOsCE38i03Ja2j50lO/l7tJR8AAFXMUlMNM+I/ahc3lVbAF6GDG3I6eZoe
p4jl9F/qhas/ZijBtKNmMn8a3xeBjH8bTzTNsYrBBa785M1+gd3DotKgGKIombHz8x8fJeQtlia6
QanUwAWCg2An1rT3tGyRqRFqrzFmd7SKriuiC/BkeiyZu9dvT6AQQW8E6t7UiFEZ91cAO098xo4x
uEVvMvVf8IlYQrn4GGOM7CogUUynlB3WjpCiBEWCOyNMklrBtr9AXRusSUnvOGo76Z418Sb7veNZ
1NK2WttfH4KSZ+hOUpCi9DzB49Euh08WSfvOhbwUDvDy7gGzhj0DC6QfrlTUgdFOlrtL+BmP1oZl
c5IpURXJADJPEmaSFyRn37MV81K83V0f5Z5rsmyqZlzGIztBbORAMlpff97PCr3fWExivdkH1eHV
GsLA+Q8xPUvsV6X4tQ+U1f0rgw12SGWwfQ1BqYfObwodnpuml0AsPSX1IohBYz30eRAXdv9g97Pt
SjDe4oG0X3kCEfmSJJcdJB4rJS2rGGGc3j16qdIM8cE6NMHRURogAMeFtaXVZjaIsJTQ9Nc36PeT
kpt4bd8/th1gKP72c2CDXO73CTb1CSioxT+giK/qwTwnz9EzeYHny6ze2188KCzq0ItSHOSZbr1B
vaROh5sPovz0SpXbjlL3KIJTVU7huWMnydktHCA3NZhdkhQJruIzeDInmvJ2F34rvvWZW035Puf2
isE34u3oNXi+5aCmQBDuYTuXPBmCXUqc9/UGFIqss6riJ2ByUvb8w7Bnm30Zin8KP2yJmCiSn5oX
eNkI0FiFUWLbT95+f69If9eREBuuRTIJWZHTxLPrdpV25Eg40Mixy+PtCX2idf6XhYQSx7bj1hAc
ERoNFhTR9PCHqooQPD2MzxZxkRHxIRdwexCg5L7dgeOdV5MhbnoQyqJ+/m4PSmddQj1WPV8eGeqP
xj24oHBIZSqoaQUOXP0ohROmB0Ye6IHwBObBgEAxv53YovrjlH7EcsPjLluBVyprWQbhjmVwCiYM
iRUOd3wi1aCNw91UFN9EJZ6bDnU4ZhjOYUD9XO5nmfZ4WLCUOKJPOFVXXMP+UTECGnLuxDAvuuu1
utrIeV7Yy/QvqDlYT6La5DSjsWTXQnf8MrXH5K2oHGTjan7DR7ZkwSJcB7ynuEpqc11WWnhHrNpx
aNxZXpyPy2fyVNPa6lBPX7QxEjCqiOJGDmfjx9GmHwSb1Uyhz9kIKP27kCtrSyYO0IfIAepzHjb1
MCzju9v9NIV3eGgWIwvCMjuWQm6XPGdXcWw1vDXrEIAvRdDdGAQfrI1k914RO5UV0xXRcvLUqstZ
CDD5BnPKtEt5Z/E1+er4+k46OC4F/UZSK8nvHCgunLuQgipq6h2Ltm3VzkwvJUoXQp/MJbT2BGvQ
lQ9ZRTMDQ+CBrGicDIkaBXWvMK72Xe/YT3U4phrCmkq+qbrD0PxK/5xJOrx1yCU4SnW3tjezO9Z9
tfx1/h5gBhmCfEbJKBO2di147t9+Jf3RnJIqtvMCMjJJ1kOe629jpZ94IsK2NOx8v/PIeEugR3y+
FruuHZGjAI/Cq7WIOuyblbQ231Wq3kN6w0P0qCC0LIf+VN37LmFakI0HbuLFV6wnof0sW7lmO5Vr
NKF9Szf/D4xZGg7RX1I1koc2nySWejR4qHn+W1ZzTBZXNTQZ4Y2XG+aga30JDVEqeKvJib4KXZiX
1Ck2rgU61kxN3j9z4zZJ/u8hWxNEJsJDMNHgNtpGp2a9EW79mzL3YGn8j4a2i19X4mOyvpwmU/J8
sUsSfwl+WItDHfpHd8O4YcRHCiMvw4TLsrfDmofpokF+qvgbCQQXrO0OhDjxKZZMikihjeZWGc3Z
39WrcAwjDmqp49S8jNXueL9zDGtG6USh4cyJ4//+wx1d2uTYcQqPAs0a2+j/H3ixIf761mGlXCxY
ZuwI4mMteO+AZTF1/r6gUZs9LQwFEtPyVKUMTJzj+GPcASo81TmV8qSbckGVml0aMYgM9FGChpx2
tN4pO/ec08jvv6BsKVqFj+5Loqmqwe9dBQ0YkeLvrILfE/RNhWbd45lQPBXysve5dlMkXO5vxWOW
5TDTA5AK0SB0QfV0qQeYGYI/FsoqLCzoqCsQJqtq9w/i77tv7JB1I8mJwCOvHsBbom56E+S4dmv+
NxAAO678Ae3EuEHoOFY3i0Ij/xyXur9SDIBFCPI9QfUuEuYNvS7uhoonpWm3QqfmEIiEHd1DsD2+
Raz15EJd5Zs1MOjwX41f20zvGqkPe7txqInviXbWIbc4KW96UgDJs5CZ8Le0knDkHr/dTASadAu9
8xJYu5ogP7BL/Pi9Y6xSLOKb/DBh9gG/OBHppnbrxzr6hIwjg6dtgS5y5tQ1foH8T0pLcY0FFiNg
y0wb5fRjsdoEpWMXqeV2V84PjAzbIR9A9ILaCJeFP8QsiziFrhpVMwo8BFWxi2rTZpSBFWSKpa3u
AKvDeGqHFhIBBQxPWvydRuz2LHzZR2608ElG3HXSC1XMg7zNNUmaMfiFnEOjQso6NUYNoYtD5r5o
hIU68oSobUlHM3DztBXPpsgagzxO1q4bqMsrsaliCCdLMDHqDNJNphheO1aRupynDyxlz8yG1GBS
O1Nd4pupvSDXw+D8rDLBEimMNLM9g+EhMGV8jZwWNBE3nz8NF+Q1KcE5EdbdhrAeIGnahr94Po07
KwewF+jj0Wq7H9F0eor5bjzwv3Gbev3zV5bIAWN/QdXqTaTZiJ0GFywwAsY8AD5426lpJkNDeG6E
FkVJ6VKGe8eLiuLk2Fwhiz2NftCEK8xGIEWfSIrD9t0XPtY9+B+8TDNfaArZNXhJX91SoxN7oHDO
XlwmqOr6CiwK4aylMCcu+lrmHWiDy4ZJyvV39RYrEvIRn3WOe8LNiuabO2ZWdBGZ18yr3NLwqqxH
3fEXCWd+7Og11/8AogxZhj8rY0+h/Gh3s2ysngYpcC7K73YIaY4zswocwP6k8OeNBue4XLkSKQPS
PSMGYYxmA3nWVyJznK4sI4QxdUhKFcDmmUKWVCk6mP9BumpYgxVisItdIWnpH6/tL7gfiO2LxvVt
gs+AXmwbAf9eGG4mpBsGnKJQApNFpIh+UXcMO0SRhIYCwVjjCiJ+wbnAA+OPj4o43cYKaiH5ecyS
vBz4geXg6JNBwOMSiJzgfc2g4+NcJ9qeJx/ulijDyHG6TDBEICAEmpPOtx7XNHG70X0qPCmWQHAS
47ryVWBKr6i7ubuFeY11jWndnYXvnsZ+ONt/oqk+hLoiFHlPFiMwfBoJwF+Y7OXNYKMWmiy90Oi2
SNXY671nLzY9qkX2aLVHUoVGP1GshEU3Mw0AusOVG+3AQDPFs+zh019BRupW6NI6jKG4HbwSbSH8
pkq1z4W9/hnkp9kjJKDaBfmVyBo8TYZlzuyLlmP2NLSGOh7biUbuFmuV7KJvnnvFkAoeUI0dFaXO
KHIlUJCqt2G+8UnBCS/ZxnyBk+VCJRNxcDeOSqn4R+FbduPItjABPZoacCdSfq8OkZPhjJIbCCwr
xJ964c8XIEyz4xdXLb3nneOoShMMS49hC3XfC/Kf/wxXx2nEfMmXfL6uAK7t0hh+zZsqSMcT+CpG
S8l/bMY4izKn6/iuVhIpOQtC851uoByJocw0QVRgDNMFY6aL6bN23vpuZoDyBtWqXmFFIf0cwmwj
43olQKQ7vGHbBriaBtrqgnbCsYWiNcTlEcn8jewHfllwCJxot29IxNVUhkbo1z/kqssHwSIHdfba
XvrmXv4caTRHOkv8h9uYUEm+Y/sSX8kfgqPiR9lZk16a/KjTFTS5/qR0pByhXn0b+nCOGDDlY1tJ
Yzt2RcsHXBDUtmnvk2kt7wjfX90zycUTu9Q4EJiMLqzu8IJXE3qI9CS0sRaNT/aYb3ZjjNYFdUyW
xFMF1UMWxmN0Es2DtmMmfKK+Wng0IC+edyArRI07M6+GQWsqin2gc0hMwQ9g6RDfwetg7nfP2cgZ
GYbuypun8cBTTldhqbZWB/rbcsQkcb4XqxPt9C8DyD3vGxrDPIpgNV/yI6TiimvDUsf9eWiWuFjE
Xq9fl6dDeBslMXcw6Y5lSxLzrJYwvxBVVzHR4E4il8ZWdmefBuZ6H6uPTOp1H79D1tAo5Y9+WzRW
AXpoltQIVrd182Mm8RSeYYG1JPZAAvk8ZL2/BRz3LoD9Iy3sMEwGm/Qz0aNNfljSPwLUCeyh3CPn
2o0pd9DsRcco+eNgqa5Y6IQJQUxejJNdk3r6wScDkvqKSX2VXrAiJOgU1pz0MzSS7DrHNyxGdNqD
WnmhjiaSs8oer/5S7QJAUL25Og5uKmdUfh4YxoYe/aO7j7lXEy5lFCl1/xIWkcjRmRSm3pt0u5G8
Ps5FdrDb/GHf9QYpJrWkFlSl3+Kppy7rlHFHUGk4gNiKKX+BW9Md9bo7CKEkhwiuc3xYKSi1xErj
SQVRfn0HH0qZoBPtqKlpdWQa8tViHVrKbQPTgDxxLM/YJf+y0EPm1dR4kCqLi8LdsBQp8kRJuWoC
fkP/GiwR1XRCxqd412l2djVc+VG1Q3m/M1+k1+IIXXNiUTv6OcaWhaCmSwMns/cKlbjyOQ0JbjJw
aqlqvspQysUcJTmb4dP68um/MiwgazHSUq5JwjYiZVAEBmBGNRkXp9+sDJAAalioRG/5CRMEvO8U
qiarneKiao3WbS3LqDE5ILtgU2sUI2ruqBxdJrJgxEezyi7qseDc7ptYcZr87P7oIP4psA0hZXGe
/A+4RrIj9Tjp2O9IZmzCyj6ifdutg18l5vPQKv8G55Hihrcs7/RmBJidbAgBRR7hzRbIcYVOilrn
DGljPL4pEPlBpnbppk7OHvakXHKs2KMOdBdtqlTsUVZNsvOOaD16vBBakkkNjMOnmukr/BUf2Qul
417tKU3tI9ZCLsl0NijHQFc2usypFPWBlYXEMBI+YsmF5QdEcS/EMGouX926+czxTmSwM5IVPadr
ZUDTBW5NGRpaYtyg8xjuiMBIPh8X2wVEdNrM/AE5oG1cnya6G6hyiTUoyd8U4ozm28P4B/SCD8yC
TV1KGH6lRk5+pwBI6S/FHA8qxjN4QdruJReBhXyyEPiunGm8uyGPITnYO01mZFb8qCe/ZHoY8/j9
XP7lvdAOox2mhK1irzNnrXDWcWJo/aFh84om9XVe4+M3zXQpj7BIUlmM+1Vw+lFr+p7niE6Yd+/9
usXinvfi9gsrhHPP/6UAZ/iBsUxLShXo+rBNBFZG/7WfoK6mfW2imrnq6+n7LYfOT1Z3u3ive9rJ
+Ip1pElvUOwxKKBopRlDtGsAQt86MCdzuEo4sPVPNLRz/IG9LD1IkBsPn+WK2EuTAWC1zlhB72V5
F5NJO6G1YvblsG5tY6fyB+g7SWoobyMfeX/jsYBLi9HPs7ChWHqU00gJbghUpH7BRqmvDLfsRjoB
Ku+BXyYIJYJMwSxjIH+yiXvvMJ43RF3h+z2C/GUc11EGxzK5gq1hMtmEA5ezsioy0tN/iU6YGBA4
tEhzxos1+6eaBRwt5Xp+xgrjVa+ZZfTBoArpAKxrczC2EUKaUVDzYnGlosyVKyosBrojfWCDEuhf
ZUbCY5xLXN3PY0JC6MhQ6GQJcEo9iUketQjbH3cp8ezLgCf2RvinCzaD3FMQszAnUxFMGPehNK39
cLSCpQLR1xvFXRNGcK+UZsKRTK7jb/+ZONsCu0jWD59gdFZFVBUCGhPwKakrPIwBRmyHkjnjCNtY
v1///jzv8+N+0vPCOHQzKt1jL0xIyMdNm1OAJZREYrSmFGZlM+AGYcuGa7yvbMMkSIoCAIQ+qnnU
1VgPlrjYrp+zoUpQhBw1Y4MAYpLiltm6V2KobtyIttnI1uPgPLG0onKzzqcM+oYNu5GZE5XHLaNO
xsGtiUMAT9s3JwxgRFTeyeOZbUMKVt3yUhrtwIA8Kc74oMvJgLqom+WDJpViBO7FVGU6k6Ts6BiK
kgJwtzSwrCbMTS6tQWOFu3XxJGdsh1dyTMY3c6+IuarrltIr0ujy6qiy3yDPx16vh/E61+qaeVkP
GIkTMiaTWw0bLAqPuzSaa+GVizRxwCMC/zAtSicBOKH7CV/eVCUU73ixXhKsuER1LTfhkQNgJnp1
rbpv2SgQa4p1XOsrudlG+0d0mQ2TIDoDwoH7bBhVglxsgH5Oz7UOkPGkCb/rN4p0q7lRxOGdumVQ
GODcaU7DVlB6tpLqcGHkyVCXzf0k0a5gmLpJ0CpqiLZ8d3w+AnEniBXG63OWl9vLhKFJsrWwWnp3
XK8AJTf2E9N1+Yxv03H4Jxm2oyfyKHcR1876OcvjxmdA+MnpDIE/gD8eZy8GnnRE1dPpyTUKv+lh
5MAG24uoNm1QXp6bKlo9A8xN8JBgF0Y+PGbGhVnfmPhdxZa2bCBLFflXfzhzDQmD/p78GqcaWxAf
MyhOputmrHfylg0MYpm+sORNP8L2FjSgXhYlkMk3cmIxBqIP/QYDhlJX9NgN0q5BFe6B6ixz99rd
dT3HUWAbAO15xn3IwLaF2IrwCJ+u9SdlFrxNjWcxpXe50kcQ5R73pG/hlWEjWT/gi5ZoL0EoL4VN
grEMn65j8UcPGtP7rZQteD0vWW5Vqk6/H7e4kGCxOF8Mco5/7O9MOEZn9Kkd7hvzGAIOodoqJ5jf
90xuBojQqEBnwS1ZX0MlvSkJNXa9wl44wAMEQhzWnb4v2uKXWOS8FoRSWirHJybb7Mq4rZSEyQTs
4zu37+LLjMW2hbvTAy+lVvp1pkl7s9Eg0S26fyQ8zq7wwp8sjZ/rzwwe0HBDluD/8gSn2YRe/M2l
u6zcqv4jPbIH4DR40qPe2YWUgKXGokwALb+uZF4jTyOgdnX5Cedn2VQ3JQd+Kooq4MkWRvRjhUtv
dl117fiGZHGorWWupkhVyRK1p5tfM3tX0oxGSmqdN65pds4LBDp3HBnGkgo9BNI8ZoVmptSazE7b
RCkOuOw26bt4xdUAVZuWYN0060iAL5a6hawy+0qYNSrDrTOiJ4FekZaRAc+up8POLpvYFGUc1EBW
5WF0MB/JW0PvzLT2kjcNjJ7nC1UUiR8iIOmsSbDEMi3wq34+dzE2KUQKToYM8Kp/kSqRstbzQLP9
/7GzVUhAsMwtcAqhX2mg3pAyqzuDIg3TBLUDsuPV7KBH6UAmIZnhyStPPKbfaMrQ4kMPOZMJdrOy
T2LMRDBArxYvVKVlZ0WFZx8xTV3gmRRaK7IYeGMsBDfTAhxf6OE+k3tRZYahsMFHOdkp4qs2+0Gg
PTo6WToBAYTxTfC9wbURIGy1dof/5JoI9XSF5C+axs0w23Lfar/0l15V3b9vVGjl03AZlOTugtF2
ubcx9LYxW1fFmcDy7urvBDYK9ANiQk+3pt0zdmUs9+nWa35p136nspHSuyuuO+f1dWMHG/AakeJT
FRYYgruaYmu+A0SJqmzBlLtQvGQMb2+COHAyz2whISyT1uNiccSJ/hC94MTwk9QKcqAEu8LMn1WB
rtHFZANOxTQEUnZauvOfJKNekGArYjaYUcA6QfuZdPSKFB6sZMYljZ8qtYL52wuBlqC23CeILTbg
K9/MmgIcdOn1Wh4M25SeMtsngJz6S3hpjmxZiZ8M1JGp7PMPkfBQyh64ke3YR61OVPEO+hANCMql
DQvbjNkUTGnF4HXWW37dgpF5NgWhyuNLnHO/fLhRaD5+jx3uR2WBkJT9nHWHZbluse+XlQ2+s9UT
Y5958VXu68rl2tQXPBpre85MaYDHzGg24A7ycSxZdCQZeBi+ykHoSbPGgUtuohUG4G0IWQgnCVyH
13PnUPGG9aG/tM/iaT+4m73gU9FA2mhJVLcFyi21maSXZ8YhqrRlEaOm3ItY8wTNoVBgBLOXoiBW
JuefO4ey863YSOe2Hm/JKHlFfsqrcVTOuL4mdamPCumYMzsjzjRQZqBlk5oBkdWDINaKoRM7qzfT
t5CmaTi14kduLj6pcEo9pKnhHQlzwb/5BAiYR030Xfn1EKT4a+wfqSMHXSik/N0v3EupWAFMgwom
8VHe7slxX8hJbZ3rHahNjsNObFsyBmxSypvA02BjdBvsfxqc3pqwRrwFbGZxtdYQG8NfKJfWB9TP
FV8mDghXE8u2uebUGBE0KtjeSQ8G4+TRrGvImzS8WpUfUC7N/C0OOOM5xaiKdZ1sm1zA8OSWQv+f
6DW+mBBS4en3pB+mcE/Z32KeaVGmcFlHWfE2YUzGrhtwzoAmMGi0iY/aL1Co7v5G/shC40wonQFF
QZuc7+BinrxFudY1GYbu/mswk+qsCnNQj6Jg7rttvCZ0Sq/2KzcxkSloMF9Zy74laOwQxsEEm2N8
Y7qu9oYdXLIaQsmhc5dvtLnCWmqCBtFjp2vM2NvSzx6fmCX9eoN1DU8VqN0UoP/gbuotDgsQhxzr
O1m/4icBjqd/SWb8WvpJk+RUyZ4hLA/rDEUZt98Z22EoLHeeoVFbg5pomzLdD9fYkSmAYcvl+LR4
4od6zFnihdJqAbVLjelj7HZT1nLswKp3Eu2yqOlq4uG2/21ldH47rg+mE8nBgdR5SaN1YcdvKSnT
FIoTd1M2+ZqufOkKJaSr1s6hv6zPi53D7/tQzZDTuvzkHOMHr96qmWmi93O3y1HFU5d+kLZJZXq2
7fN5WZPNyRSE/97hQR0TgQ8kHGJAsXUfSky9aH3i5kFJrUOVnbLiy6nPoKy97bZvHpWlyHcxYJji
o+JwEMAziZgvgLaG2YPEH/MDEonbuCWmVp3Wqc2/UfXi6nSy82SeBYTo0DbFWx0GKOVnevHB5tcX
essugDGjtHxs/W7SyFdxbiAFUBEC2Ff+dMrJss50sddfagDvptuVgBGhNjhqjIiiPWKXGdYKYv0O
16Cf68jYmsQdIINN9+H1tmmTaSGtNQM5aKZX7fqJtqFaGbS3BvNn6AiNrwFhoby6KJsEpDrXmsPO
K3QETd+4h9AtfPd870Hg8FIgZk3LHfZlYziuem+U9LB1dRzExUP7vztQ71ycO0darN6ExYevwyzu
NzUw9iSM5gZMiSXmOSceR71LBn3rX1wkS05SRWZ0Qj8ywpJqzdrvaTIKOMdyxN6vsHnurr4NonaA
uBpmxWVqNSy08VArFq+1WXcO76yXHY3kcP3RJCoi2W5i02b1+WnT8Bjoy8VqRNT2QmkfZdl6Eamr
kGPoO5paA9i+zto1X/hz3olK5dmHsk7LmCPHoCK9VfCnZblDCyplnbITKKzR+OfdJ/W3WOIGD0fr
OujP7MTYs/IOYycmr+3IBqmnoVmV/1MYyXeFDN+uz8JtHmZaQrpEQVkVTIgElSuuzVwGlIDwCP1+
qNBzMZ0Ho1ZCUC1SKBjtvsa3Tecs61PkPEF85AiMbH/CgUJv0iMrb2YuREBo9USdUkgYmJwL/Zto
23AEvg6AV6DQc7zpDfgi0vwb69ns8LVto87HCSguy4R6R4QuFyxCMxL73GBkiKacHBC6X1w5+qIT
Qu79L7L1r79VT02svmgnXhrDMN+KD8sJ0G+lnJzta0cD3e1YZkiaQy5AjOvpXQDnwB0ESLt3IKXM
+WGZ0GCAWE/CEST+2H84dHT9mFQfCIOuu5TReDeHGav321IylvzLLst9A2t1VJBH2Yr4A5NbHL0/
zrAFE+z5CQrRd9Zyoh2OVd9ydxydkxsd5jprm72OhN7Cht13QN+I6+NS5REQ11NDbqI6pulUHiYR
UUIqRBXe63Yf7hLxLNiuZ8LPbmlp9g84BEpYcJLhwBa4vzgr3Be2VuqwDWDVGOzrtA3wr1r05u8B
+Pin174iIW1xoRT5HzN86LWq4qqCOMc9k7pYObokK2xOnhDYeGyHkhQoz56Ply8Wfj3BAU6pMHYi
D9NLIVUaf+EzvF2Suf9MiUTeT/m7HvbGNYWvPtNV6IZFBn7vj9RWd8eFQ6ncDrtW6eXAX5t7YdI5
7G2GgF5zm/BemtBXVV25sExP8qPjuB6vACOf0ZT1K/6YIAX7rm8dID6p3/1BDYCwFq/7iueYmHz7
Yjlzzsq+Z6TQjAmi9Dj6wh9gNtNdDVN3A8SXaSq1KghfUjju7Yf7dcqk4rR12PS0A668zEpnXi6o
KqyrWIKBeN/5CRtTSFGS7lltJ0ryXDByJkVwNj1rFgmO0sHDdJBMq9djrVIqlaOfeErq9s3fFQzy
mX1bQWduntzO3+rknslN6/TX+WoalNe2hU5GQuW0oPO2ji49tX9ae5MCIht3BpHl74BSbm9X4x9J
qvaAfwvURSSn9iZYt4miIn0gZH0Jim2cvZnY51eKoCi/8hhtw50HDpYgehsLsxKrC2cKhpCin4+y
x4x4fMTTI8vSxbAW1Hmklqc+QHLOrs7HD1y2b9MP6+Dp2+2hpQ70E9gc2YN4lZN5jlPr9ctDx50j
wj7MiUk2hCLvbBbmNBI+30lEWQiphlEbcMhdsXaZxeD4jz7oPLittDMEGJm58cKABE4E1g4Rtltg
wFC0oQXa86Tm4Fm69Txek4SpgxWKBRKgCLAIRyBcRhgD+XLfvDVGymmwPtjv1oi3B+3WxnXyxGpf
jupQ5x281bLFi9QPMXGzHy61Ggl8M9VPo+5fPed2Wu9EXr2sCnAwtB7XRDoHtrgeCrcZgZmy6O43
Iowi+ACYn+64Byy8IzW/K5wzx1aHf7VwhrR0LfFTUK2TamCan/tkCtjZAfN7lKdpMkFFyOBmhg/Y
SHzSjNuU7H+yCxYGP/oIz+00JuYSNzdsiwRJ9k5CBAnXgSBIjcVZIhIj+MhMY3/EYhiSX3uYpa+h
RAqtC3RKTbc62F6nobLvkeJ27foyJN6c4+dsv1rQMTXjjYar67McZQ/yH841Dd7dYPT6wihHWeb9
CCvlZI9aWQVvPHRc+F0igj7hFgjpb87B354V4a5q2zMHOKEF01sEOHe3nrZuo9etiMUKBORCpeHp
RQjAQV++mdWiEBRFUrYgTs8jO3q2i5qtPbnfREPNBOETKeS5+zg1HCFS8//tAmCw59Z1tRzup7+K
e5YidNHetJc+ikplv98AQd5428pc+ZnetoJpmTLUHEzJCkovvMbX5xh0r3ZHXdID50Rwl3Ux6GTh
6XiqDL2/3eH3Ho6gsiYfNUPLwI98fPk5Y7mC7FjcoxG2jwpFq29FV8DXZ+2+LJLXm4AK5NXEPaRk
a7HeOe/O8TzNVzNqHLxzWPL2EnBKkFR89BrsUnsw3rcSzQn+IfOGUd0tSRBNQNDHN2Hq7hRlBR3d
t3njmMqnBW6w7V7tlGhpVVSiKQsF/NbVJbADsZFVHKetoMi2Hs37jaszKMCk1b7Y6yrr9jy+YL0Y
Q3nKzVXfEy9qPTq6sIQ14+1wFhGFPOXtZ/chKutH8jMG998sI9rTrtZU4vK8U+d1/N3AfK2YLgpC
9mhF8oB4qhB3VXcBmjdo3jkIya/LmOr1Lj0iXarHyGSqGaUarAGMcc1aJYpunMS/r1MKGX9d7xcV
KrAy5d3umyJmaUwYRIxeup/aDdDYI82eQAjBZDRG4pH3rgEZEDjE0zv3fuJ2h9nrIy4Tva8J8hI7
VzRnD/PJU6gAmWuMfFEtwhPbnXezfaMuMd/B6xCYqiAJbVdx8F6gOqMNJ2mUXkZCm/rWZrYMcS6p
Rfvl0d8bit6vaFTwePJd0CdKvJJ4AV4gXpMhhs2P8GXHYzzqn8MElgWqlrbBgjudTRVkWwtfl610
dLRrRMDZMhsYBM5IM9Cd//DetG60Wu+BkeO+sU3Xo7uktoYdjp96Spb5+bxduDe6QDBDryk85mqi
MhV4k3UFED5CWWIFjIRespMChh/+ULvFAYuPs17CeZI8+XDr+Ylm6onNzn614FBPJ5lYqV5Vk4MK
8xqgucfeYdr0YE74ImUbz7Qctz3CA+uvcSErjmhQBkeIeZxbFIsVImvG8sMztgscLwCwReJfEL0n
3rLJBTdzRBq8NvG5jFv7L4a0E5gyDXL5FhAWoWz3AkbeiWWw0bCA6b+xrvPqrogMz+nL8865/teU
yc6EQANQBP4OjZEnqQ1tjzSXwSMirszjUXtTYJ/FYFd4hoH0Dbqkm3Z4M2E8YQY94ah4YrVPNI6j
1eKDPXLQwoNElRzG6UurVTCTp/390YJOpltsUCoD81XlsQXMb7SgfZ2eb4b8A2mxURuMrzefBQ1y
l2549sa5pNxln+gc2ZKROVx/QH6+V2zzmtoFBjzfb8ouNUoJbiUzPGFb3ezq+Z3bXlyYwejPGPAT
kCn8Hh+pP8PvzdRBnBiw2etsX5C1bxDDl7uZd67AfA/+rWeVPMssRfjokKWio/lPlQqb6vovtUXx
oMArj7LvCN8WcJpY+0PLUBXkZdLfj+fSaHb7kvCRbv2xspqdhnBqlKNlnJEEInQdUv542hF7l9oL
3dbZsPzccr9kdm1YsLmL8tXIFNrSquUyGtV48XRRD6Pqw8P2fg0bOM8Gpaq7tlPuhhI8UAuIX1pu
t8v3Lg+1AImlxRMB9WdLl6+6A5rPMBg+zR79fZEcePyPt9/acqnMb55YOFGsRyVAM5YY17n44qmO
fE/R3nVy447U2tE4GUFMhSBCKMeacDng2i+pSGaciOworkoJ6Y+ctg9gzHWYw/bQnUh+7ZEv8phQ
J5xm//6mpCae2dy5Df1ogu1AHBpH66TFVj/t4PqhYfhahHEWVJPicMqFKGzeP320zPVXyTgpgqRy
60YyfYf7MUbX8zXT/BfDgBJDCCPeTJ8sjJw2D6hf/g+MfEpqJIFp7ncnJHdIP5hTsvIpkPqkTqnq
OzTIG4vorTpcYvs3ZgHjtXXq1vbo3hS8S3ibUoTenF7INPf8KisG0RJmQZzINGE9vnTROBpADZ3N
/lzeTLaxtJg/Pxxq4d/04FgD2GNzuK+x23YFirfvR5NprOaXeiDVPQ5Eg+Z3TZJZmEYzfDdeUzkL
zAMB2AB1Zd2+/02ROLFRxhE3Le/46ZpAXys90upT1vy7e1pdvofxVe6oINkHQZ7JvwcCBlTVEfzW
rAByj7p4qfmazWOjK/QmGZ9UK53ITcoiol/4K5l47xdsmocrqIe46Ovi5LtemXYm2HbaclxzWJF0
Jpk4c1cjVNDrj5OdlBSTMsxLb+tnzcLAFHPGgGPl/PtVFrfHks4HeRWrYpcYZb3mB2E5aygY+Sf7
Fus80mw2tVvgV81rtB4/f48rbb5yYQIF+W5HAkD+HhzoPihSRTBTs1/ggKlM7G/uOA6NIKEuU1r/
l5IkRYl532sJbILUpzr5HPMQqfw3lVETi4qT08zsi+OA98HngFml/l5vTD4N+4Gn+r2dQzYrAQXG
gWsafvD6JbtmV8gr80Mm09v7qjkM4j1jxhL7yzzlPNJOF50kujWsvQQ7a20h/E+uSYth8NOHhn9L
8aUfKvJ25wQo6sYmh4W/6wF+hCridw5SmdfdEt5wT9dXSuC+rqKse+2sEx195zlfv616JTXQgJg2
hVu9YZpb3Ii+SdfZwmlsITA3r5BHP0MADcVDv1kkJLtyge7vM6tPyxAM97wzLh48HFyU/SFEZVnv
zyygEfRMatvr/J/8obhpXbjIMTZVsIfs1Hs3MGX/fEb2Ecg86c77sJCp6vpESkIED+zMwnUnE9Y6
YKDgkAxxKwLX985Q4x98gtUsngnjI5aswCBYF9F1uYRhEyVtvcyZqXVSjI9KC4S17eiHR2fLSqD6
jx11lmJHruahkqlMcgEvil5vjPiPCef4f3QjhuRgih5EXEDUujYQQgCPY4kRQ7OL4qd0BPreczxa
2ZVPlwNYGRm48WCJg5XLdB2jflqb3I/yerIBWLP5ZsATvLx8aBB5ewtxKeKIM1bCRzaGRZuu7A55
8L6aEMtSXMlad1UQhRIFIq+4iuIPLWk2l8EVkHGLY/tFJvE9l7kir1YP53zHnmUMPSUK6P34cyR0
lfJvgNbk1yEG/29BFZgZcu9s8SdZNZjTpnvhU4V854c8iRintJ2G7HHW6OA5jWvM1okUJ1Ox4a0x
roBYZAIaOhGFXAvjFeI/4wNPXUKb317+qesrEcAFgwX9UjbpjPfF/xcyfVs4HVsMsCBRFm/Y1vYq
yGDJTUhtUdc0clC5szVPWlpTF1W7CGj+C4W1FtrrzkBeYFab0/6bN6cVUz7wBl0PpE71rZ4+N4jj
7Zhb+DQOhDwq/pEezR0YBWeJEm8kjPTZIzKHmTnSOON1a4fzcUtaunBw+z1mNw55PktQ20McobHQ
rYkxVzL5I1JvpgEe0R8MXQzgs6VafMrfyei++CtRv95L590QTdc+lf176lYJ4tt2yzX+mudt3hoW
4hmnJzG3yZswchS/4MQPGzBaxKrLgPoLvZzCyx6HJKwdjTbKjf2HCZl6dqKewc+HTFZ21+DX1eZe
6WvX7mRPKYlRCP+ID4RCVZAyt8W06Cmk0aLi7LjtkTNlrwTU3zan1jKxnXaTcaTFqkxmB0H68wPK
rYfHeLzUoZ9XdB9DBUIHZQMAN5sa0AJMERJuttIJlj1ciWEOD4YCPN1Tb5wOaW+fpySr0Wo3BVSw
6H0qgPwds7fiSdjjFzboUX6kDAoqUqab7Q3d1Tn7oM9Hgq4h6slBHSx7dNDS4q0iFJV5a1EU5nNE
/hbWXmXRklf5l4sw2daC+RYXcoc/lIwp1wczmnqp7tDths6iUxDi7lT5WdIBAFznLICfHWx4vJsj
oANWc3fXvseEdpW9kwbF3Fgfeu9erDgr3WmykYYMzRSbrgihBnOGUSb+0b6sxLJZFzOMctsxA/5z
Hj+VdIEkc4Tw97s+MIActtwiHjizn6qvraeiEl5DXRlRmTBxXXgyyTEZZwtDcDyLyRyx9Q38xbCf
Q7QsTkawoONC9hmtEWtPdxqLrgEpPX0nvRoUI2G0DtPhTZYfFzUT5FA93QRdGPWfWeuTWEabG0YU
sEGAFz+5zFKRftkaI5SsyXousXGVGI2LDH4bf2u57pPhdJajYwc4PVLvqyvRUatMhRJtzDNpPuzf
LJAbyBR8ztaAqQx4Cp4RJx0UgSeoBLXHIhhfcn0NbncUgYjmWuagU3oHHOgBuAfuTvlp4izohCha
1/JHP5S+P8NvMrhZ3lV3W0TagPqA2z1OT4qVHYq4pzaLBhbaKs1luaGD7bS4KCEAgCz+/9MVfvH/
bG+LnSVAjbZTN8osJH7ik14+s8soclpDgzoMes2deok4XNSJg1XBr6jzaxcE0EEi47EYeKVmAdTW
Z4nySps0Y1edV+ds5tTQONO5DUcpYHbiu4sGCCVji/9XYf2FVFGbIsrFvd7RLEzh0WyGXfuHiLvq
8z9rcGuEuOBzNRURtregPrmQ+WG66QNr33VzAWmwCi9NL96V49eUYYgKuVPT35zF6FqFrqTfEZmF
wuyvhd4hyEjebZHAD3iiXub5M1WEHrTX4Nd40suvdFIWXYyA6QuhG/n8Y3ZI5HAgTUWH4JzVuvh+
Z2DQEJDm37+PzSQC0lWwYaHGiLfn7ttr+iFYw2jV0YxWGmVqbzM/N8AqYYZL4EOru+ccvRYQOp5X
hGpfG7CznowwGlAzctuGOYdi6YBZkAwfVVhF+rChac31uGY6n34r9U2Nm6gLt2v5XAmqT65m98Qx
pZkBmF33jXX5QWyNHkhf2EmHRTk5U5u48VNIhefV4VlPQFMcCww8RWO9zp1BvzuzN9DEZR2b9PW+
j5pu54ytAF76xutTUf4ZUzX5lYjaPIMfMMWUtGh0hrvowRY0V7pW1D+4ogH/XJ3tirVpfW2yvN//
dT0f2HUYCHb0iJPZ0+Ic1HEzTgwLCCv5mXMOOUTzB6d4q2w3uCtjB0eP+5sU/n+eSbSKt0cVnZMi
KBix0SZxsck2RnffaV+uDlKRqubd62uy/BMRBZ9zJOVpkRaVU/XErxUfqEqFAtKUXuvyX9CVKavv
1odWmu/kN34Jro9ldTnFc+0+Q9ARsgnkdjsOEMMxxAsjsfBOdoHd4Ck0tfkHsb4ol0+NvMuleiff
9KIUffqFRo4tyY6bnko5AXiJFnVlO110YVGY1TDtUj8+Qh/BU8sznZJVAJc/pwSLKtWNmH2CSHQf
D3FBlFasddukqtfs6hM1xc1cd+ICD0CJjQhjhWdakCk8m2XTvgcXFqZWxNr8/1CamAnQoByDFrtK
8ftbFVuAyjJT5mcI3lBxQ9u9o1xuPdLk96bnkmP3DKf8aqJheUQxyQcMLUrdKnHIkeFj6UVSMy7E
bfdg7jH13J/7WJH8Bdsuj/Bx4jdAms7W4uLFoJ/8O897EHDriifvi7rgyaBk1zzmtU5ptmVwdoFF
RLJ34Uu+XYn9pasIqZLY6k/56RUIp7DiIyndVvvbnDrtpAJmp3/B3Mi0TzKEyfoXyJVUw+kAFsSM
8pIocNIN6FveBO6X3pjbO7RhqEevpZdpA5pk0UTsK7gHXZ7iK7fDwYCGTGYxSYKHfMKMpuej0RV5
V3BiRlsqXNQ/S/WEpLPBKmAqQqk8AaaOQCuSJRKg3eRkbmfXwLfEFaGZJ5YUzAYKDterBnHpSiv1
c5iHTOe9cTdJJjiY6dRcqG9QERR/uqlTKSU+SQ/lc1GcWTX401zX7eGXvptARAnjhbrBz1BNOzGm
vgaar1DDyuCl7wSgQA8DnVYH6ysZlPJUgLhv2KaviWX33CCPRA8vXthnK+dCcUCjHHD3vtIz5Lj9
G+8Rc5xGWPxiamM92iYQFjgH8xQsZSYEshqBuP5fpZjY0IS22JpvTm/muR+He/jABdWiOtt9aq7q
7pS3L/7OlVrzRKtH7iJDkzR3zBufxtd7qrvNLG/4x12oHfxj+wmk/qCn0DPN1vLpG7HqcpP3d1QM
8DiGSB6qy8HYAbR5KYEugI5gTVKo6hwGKWLZ67M4R+t6J/tMI9fHBsBwfEnehMLurWZml2xnOogW
RQfqmUbV4LWT3M1UnwZcJ7GUSfO5F13yoXTbSfdTMRccOgWUG2ctgzzdndRzPt+GweDBziqD2eGR
Xjz8UNkbL6b18Gb7YCpNW4rQjQFdVAOd6lYKsfmrzdUfUcvaGoiZCzXSJfrfL5qXQSMTCwlymjr9
QxUahxxVSOvRfiqHSEUQv8RlM/z/7Pyy0Amq1Oh3WBpzpSnhMqNXJi7sDQO7VPWItq0zkX9NjPKv
jR33bTr4QGq4Zee7Z5u0SnYXJEPDrONncTLIJW9/HfitrEvGyd7iKK8PEnVDudaOhQNGt0Ke4PU7
yvnvL1enq5kJLB21R4UNPUs/QBDNqAkuYnQ+XKbp+RP2tZzzQR5k4W4smhJjg6kZwT7brlWZupnA
HIN4tlSD4MrFM6c8W1hSWYEshE0kLshVhFYRX0RCfhT7aNNZ2sx2LncdU10a2NMr1wIN49+LFYT/
Ju5M0JN1nXi00UFNwujpUe0Dm9VxMMMrobGojZK8Z/p637cK3psfFIh6vITe0pCtCFavL39doRmW
vgNA8OiRZwEXBEE9yL8BbxvCyciZMP/Kjgtvg+Drwpu8GjaC7KkXOLYyQbV/H2YuSqa5YFCc5fF/
tGEeTR82B8TUD0sHsR/NH394XAzL1l4MnyQhTjQzQv0cK9VjkESRBm5ngjZxTnFG6Txqdp5F0vUu
Zea+aBqREt0soPZCA2Z3/QCxly+GaUPXFLKAL9Tki7/6fsA6nRlssPrgZM0D9z3ni+ma3/WPrgxL
BT/KupbjHTIO16e4BgARU7I7XeM7OhLLGB5z4b79WYWaw9BolJI7dNVBOXDxztzZgyQ1AEcyduh6
oK/I/ylHcFMbHdWc3haTI/3+NL3PmeS3MPSGBdIx7j2k66SanIIadqnoR6DDEkLPXrsRmU5/X84m
1LwdP5wmOI5avZqlVmR+URikXO8nbLrVSfV2rVfk5MbLj6ZzZHqCOpcNXXqrrpm64yrVZ551+PJM
ZnIjdBjt7mpUNQxxURsVvHMmSH3MZnkJHDD6PotFJzMxPCWiGK/EvypYaHjdlN1GAHqrVAdeAAZa
+6DZ0td9m6kTzbq+5Wj9+BxycMb7rkNq60g/ZNGBKUcmKyu7kwzFCPTmWkKbJtLfyToKownoAGix
1IPncliGNvROVS1k4eesGdXmUdeez6gFjpRZfaxG5FXGFPv7JXjI1RzXCpy0qDdsM8/8mAwQ9K8Y
UgDyAPff6m6ERm81SqvaaNE5mv5xNsrNnjLffDERBQ6/Wucuz7ij1EYl+c+HjHSmr05FiJmUW6Dm
fUvmfyPWHvirxtPK7SguHk3Ns+WiEuWm0+3BfaXruykpYFDaP6fNG6+UvyWSeC0qIw4plU73h2yd
2M4dVYqStHmX6cSU538CzRtyxqsELzaV05RSfXAci2GpxdJUfTWg3c6fTchwjrjFVTCgrDJMF7zJ
7JTqOI+LgqRTFSPBOxBKtGT26COcvxASGf30VqFgfRZIYIhoL2+FFp0UFPsIcvH1B2rM34qTfNu/
k9WDlPFSngTgrS8ml0vXyGzHiMYNwfG+9fFg/9dcihrI1rGgMSwN5TekluQMNwhYgHnVL5PFRkkV
jgKBKH9SWtxAfeXFdXZvjm2TjlJFNMwFNvr9FvPz5Z1gByTo5fEIX1JBJb70eP18c0Zl5uaYvt7i
2/JKtVLZjLLzW+TQ+I24VRkynNTLdk6D61IRto5Q8ImDlCsZoq3MiPeKApSabxg66ffkYEnKNdP6
HvfLGJIkohE2puCbwOSgNTvHsKY/Cd9/WRZ/yoG5pTzLa1w7pj6d3EMjSAq7OIpiS72nni4bV3eP
vDAwAN4fWhlrGR3iBiy4fcf3VJfRnDJpqT+hoTTmdFdcokwCsEqjTN0e9uxpXh2MGMZsDXqnqgVo
47KzLqGKjF+V8LwSfENQW56DQjSNmpQ+lEH6mNczirZKC5ugYFGT5xG1Wxq3jl5KK6m4y/bXMdDA
LJCuVGzdeJuhMcAN9Khk/+dsqaoYDJjKkQgxDZWIJ87iYWckZCIMJn0WijpKj2uy/JRTYb0/knDQ
9Rc82BlPEmMrhu16rhlicXxxi3qwmhBSyLuTwfqXaefVvV7NSqMJQn0ZMolIvMwfC9vglXn50G92
RNiiDcacQukEVIEN5tVQqzfLFTXldhhoGE9HpeuIcDYh1AtGKzY3y3sVQAgwnt9nJYtSZ3oWSJIH
KjirBadBJjPt1lH+zib++z74cpTXSwABdpNF0effxIToXd2xXZdDQYzq47JgOffeAyUcYDOokHVG
lkLjCZlliCLFcfNZeBRv3Gsbn/0ghuJdilbCpgSGu4OnY3e4yrYL7TWoenrThUEisF8uS1wxt+h5
iZDdx9uJ2mEzbUJ4XAgxYf3ASGyPr07J5b/ArvOJ0cpWoO74lK2QICDW07HFdqZNUyszskW9AylA
6wrx8f1i0C2o6nv9ZuAGGvAcpj22vuraC80+4Im1goRdVDuRwpAjZl/rZGzcLI4pqbaxUbSdgXMQ
sKPEGj4/KofckSB7pbnmSuWAzusZ4cXGEoQKYyAlXn0R0wikSb9ffKJqBMhMcNduSP9HRvn157lQ
R9u6nzrbM59k/WxO1m6M1yRcM7vbWKR4bj4ukEN6sjlkMJdCLnV1f+6IfK1BkioCUlAJywvjnBo1
VjNWzeLD/7T2qtB2XGJBsGZW11Duj8vgcDeeNUZdvlIpXQSIUk+KLN98Wv/4ZvTBfysgaN7/cJlp
Lp/by4bH+wKdzlvnyDO4t9ehPkT89N71m2C8qiNBNRNk+oDTXCeR9pjQqIqyEyLokeEsUCXr5k7Z
IZ6NWuTkKfwblCnnkcX3rvGqy6b+SMWzIlq0xvzmtPm1TLOXwXl55h6RKhVMzT8lprR1qtPlFfFj
dgso6/hRG7fMhjY46u8xBv7GhHOdF5f6aNN5uMa5jwVZ+MoWWfLSOQIf28DMcAyRReBlU+sh3c9X
RHnq+4fxb4BRaqCnem0YyqkzbfHoGD2+tNgsWoXB9eTcKMqkX3FOLfF5OyePZbtHvqy8bdoIzPXO
A+Yun1kuaEAP8bC5sqyB/eq8iI/S1hfQYWFJcdfM315mpVsp8elnZHYZxhRUSPgz2aGC1Fl6o10+
FbfX/UTTX12XwyoUjwMWi7rYCFMFC9uNzu+AwVZNRV6cluiW5A6uOgSbqVcdflNyIdfoXoyLyi4Z
rhW097D7MHop3KkCm+QV4BPcHfdSxTFyj1Lngzgi+AJTp5L+j3VSbQwnpgp7NXfBn+TmUxfmnc6v
NfrBxKKevbAlUJgCS70xLq7+4ytNw5Zf8CiK9UdAWukW8FxZ4JMjxPoRWY7gVjaVCBveFmg4D0Tu
ek9s4WUaBHL1bu+c7zl6dq09rxDtmV+q7WeEfIKa+r5YzhoJ2zMv4ZBx9xq8WomfWGjFWtlJ5AAF
YCWl50Frrh9y3HnguRlOS6ImhzKwUvvYvbyJXri/mdsft9unBl3k+oCHavAVIgC5JsWOewPP4JxM
J76Cc5qYbzZTZRnYKTtnFluObLGZ6TTbCag/S0ShzOPaFJ9BNjHRMFOgWpimE4tMxjiyUYPV+WsA
U0AkUq8E3PzejjMM3wytBnuAAMNEVH4Ab3qwou+HuWm7NHnN15wX2a8VT9VyQwRY+9zvhHcsnkOs
h605047EL+boBCBHrzfTMW1KBg3IoFauN5U3foG7FRGZwMgOQY9vphYLWc7bpab3dOpEn+zYLYWR
F6XqUeFdyYYu6jsq26fbfpWlpx0TEQo2NyhsZL79f2CbqKVYl2orUG5ZWXagIzmHW/eq/x2Nf6Nl
mI26sFE5r8rYu56Ic0AHy48BPdCKundUtckEfNNeda/G4+K0HJuqWZA4lFPjP50sGH9gVD9rHPeN
zW3d3nKutG1yclsc41cI+CKnAPPoSKO56LELM17jMkHk5Uam7Lq/M3+xW90Cwj/nz5PdCA2PnZis
yujqmd0IHr84u11nOY5KJmVFDMz1J+T/CO0eE9gu1Px4VFA56poCkaeARmclrcgZloYai1Z1VY3L
jKPIxHvzfVmR8dMuS7uZD+Gh4+gBPSRzyWuHQgjMZLxBHwal0zFsDHRlyPQEwegaV+YMIl6PEfuI
p0SUj0fWckLboBNh90foDwho0/FsJ2LOJJsoJJmSOVR2KXXyfKOzOSZp78XXvf+BLJlHuqleAOfM
oN3y3w/yh6BPgcoA6eCGZiutIS++/Dm0ToYguLrJFScZ1UdKhUi/EBkS4nKli+kCL1o9qJtsPwKr
gN0t1T34sdlmL3QUgd9gJrapsRvIhmWRJNQyCZCinyw3jiaE2jiyTFYXUPECAfThuaFsrjz2XmfK
kzmnNGTp4XFXNzoZzl2sjSRzYWN9wU3WbOj5xdh8K24UhnehserISD/N6fbl4PT6RweO+lQutq17
MS6t6FdfZlSFvcqbvJ9owQhuV9pLkeerrL6iBWd/8EMaj66Eo5lsx+Kpp9B63cL/AbdfJeCyfbMF
g0423HXGstnHlILD7QaIhw75xRqi+78Pt7KB0FDoR5jdK3ZBjpfARWvcElgb3PTHjqTJPLaDnjYQ
ua4jMCPS+hlrvHvybd9xBEmtRlQ1yqJ/taiw0eYGkG00Fb4ZTV4vj10UhI4jP0aM7EBWpVxj5XcS
vMPi2O7BTDCWOa/FLx6JOPzddjUx19telEJ5hHCFQPkJMN4+5y85vfKE0+dxIltzkePfLzNzGpRi
Ux7ursQ0UqoRNIRo/iwA8COCx8hOQ8hvymeibsrdkqVY9PsEfK5A7A0W1nc/MVvE3Xx7lBN28N4z
gCldFaYFZXryHdDYHXz6/e2CZUsqLCZ0ng01nHhpE6qlDqi3Ur1qZZb+l9dDrXfFbNTbNdNPNTYk
yl3j8qnO5wQKLu4o/UvdeakVCoDpjwHz5sDjZTKao81k834iQ9GRFsottbdy/crcD5D/tcXSo2MM
v1Mdd0V8/tYxGmvmqaU3vOuib8b65wdY4ukDeXp8fbku4TEMPHmjO7yAdPffPz4HAxb2Xf9J106y
UjAGHVdlEDAHQkILnEonpRYTJRn/OMpSM9YiiRZdy6CnkxD2txuCtRQPam/wftcieWBFf1FoOlDM
zUaVmLGidWP1dmKeQQBYKCoHsHOGugqNiywtBT19if/LYpsHj+uTjX3Y5UnI/T0dhrkBW1Vtkiw+
rOuubV4pcH9Js8ixBoLy9dW/60qOB8WMlwEfne3OL9JXSV9SygQFV/8RGGW5obUAVJS5QGZQ+mNv
karzbTs8AhS9npdYfTwR76H+nOalyjyokY9CjnsYQ6mQ9qLRrLWiiqOymWcRmasj9jPKMhA0Lzyv
cT3Mc1FlygPg3hqiC4Fqa6jebPLuMGoGD1jxOtQk6Vf6xUC1LK/4ymHWpNGI5BYQ0OaXFnYrBHZn
UhceRaK1KHY1VdkB6OV+MLo18bQdKK/zqhFhAxO8ZS3JZ26vNqRfCaOhRL0W1kYyYaubTAo5czuW
JFtIT4JQoMGkZPLSebEtJaoErlVO+GUE4UxI7vhlJuqtDq7aV60l/No01VdBG3+UvN3p2TEPHIkU
UqrT3gTBm7wQMwpX/IZSKtyjM5HRqxmcOquf0ynKy2XOizJnaxFUDUY2gqlBHO4PEZrU39VmEHWF
mwA87yY1dT3pUZhY6rnPNOPTFkBpTovdjA75UbU+l/E8nk+2K8wDnuIcLZP+JMe4n0DDfw3gwFZE
QXNV2YOiNUk17zZg+L6CVMJsMFutJws43gS+E/PdkIfnDsoY7Uf1BdRwkXs6abvmsDjw5WeQtcSg
uc/jHiIDeQ1dvm1Z8w84+Owrxf73wECJXTgA6hMn0dmQBvpNNId39mE6kq25mSgHVx9w9cqmDmYh
XKhFtTrhu+mth0zUNbDnlwWGWxDKiSH6unp9AjTZV35oEkvY6VKF+YF/tFJpJfAwsJRKZc9t9qcZ
0fqAYc3uFPwvm3oF9cM6dLf1vYa1qcuPYyIdzN7mvikcGBWYJgixQSb7yjoj6JzWx8TKcbsiP83O
tMJ6BdSiVMs2mVe1KRvGaaQfeOmtUCTMyWl9Y6kWBLU8b3vafMdAQaIWeqzeTJMIPxT2q6fdxZgz
c/IgZD+zMKZnBS1hKfcXZLuqX8lSvzuvDDnSbIutr/pT1IYfJzcBXrqMNInj6HmwScJPNjt6u68q
Ze3N+kFoyWj1fUpV3BBd68alCWG2+7hjvlMHdrDcm1k7HN5cdJtj8r9nCckS9xmoBgxgQQ2xnikY
Afdo1HDbKHBDUiTdZPyQoIyyaJpNSCR4AJKIxau52w+iTB86clx0qE/qxbgf8ZXa4RpG95/8uwjf
N9bAizo0Nr2M5X6dgUQhVCl9e4tvWToZ0lwftQ2+3ms5X0lgBHggR9CLmdTgkNYj4Geb73oHdnGk
SJLO7q39TtwhVuDgJFLML9L5VKw1VOzirFOWonEy9L2FC3/1JiwN6bU6hAOerjKj37bgYus8165P
Yr0okLx/JnMCye6RAaQlcwclSO2/xbVO/PgddPyphl+pWkwuawPZ57aMAEPVcT0nJVD1X9CsjYNd
0HNCDKJ7V1TMOorwRX5DJbalgm+XZT8MW8AZxTs7rrjEoznKZwckVzCjU8UZFS1PmxQ47j5shVhq
cKnYiEEkPo0gQ4urXakT6T46ZxC8Hdy8Vhrk+fLcRIIuxJ5eTqlJT+eCb82cPmpFcq5IJnNqvZRT
XrWtVMBN5CiQFOoGzbjB+cVyHYq7xr14bOFWw5H/MrpABBZhHh7XuyEOCahWlN2B6yutMeo+P5Ue
SCXXFAO9w91pIaawn53BCYg8ZvG7j6N1WG6gYiAsEYXyRcI8PurhXJLSO7Tfsm5LpPm6a+HJcN7i
Kr+OdVhRQzdBQsmqSZW9OP6fz1ktnLBVCfQ9T96YyR3N9Mc2KZ+79XYks1mItF9byvMhiGAgxBom
DZY9TiwmwffZXRtl45zTeMLF3SrU3/qndBUwhhfe80t66R1KXMVg+2hk2Ic/XSRnNAHQ8Ons5/cE
B9AbgGrf6371/5/HxfdMtgMoQV1/OpcS12RXWr4c965obhirZ95aS53Xz40H73VaqmcgFtrd3b3n
G/UuGHRYf/4S2Hd487p3LATX6RqivxGblhOYdMy4NliOpBCfoftV73sSXgI3ZuB9Gpx6nmRYIQKz
9T+Sf8n/WUPJmpB8x6ih/yyWGM3F5Mlv7rkIX3X4lgKvXiYq2rHwhu90HALRyRO6wjDxKKGhqeM9
OUyUna45kIRmZl4QeXzTJo9qfAHflG9UGxoWz3QsXTUuIBYksTcLfq48wCE8pANg+PGNvoKXdxIP
1EqiLOQUpfYEulqhetCmUcVK+FmEyP/bdYbh8aZpybJBD3FlhIKbk4GJqFUsCPmwzng8eL4CFDhF
GjvFCO8oq9aGCvNsJGoz/IM89vOTymoOHHBR1Bkp4XuztlP1kdsby0BeB0OAHMnXNdOArKo2RfvP
v0WHXVXRfeLoe2f0LFTFC4poBTA07Q8SPwxA6PWwBWwMY7iAxthHulLTZ8TzD49vDtzM3jg67dN+
j+1n0y9a1PhYG46ZiEAxMoljG+StemOXcWBEro1CDx6R5O3MRX94Eyzq8NavOZRaIZfKmvYcI8bu
raSveUzT0hoY4lRh+RnmPy/yBGKwBdgFrBZUsDngNnZA0kY+9fBS3xJIFjRMpiyAjShzUQ6NpHrC
Mtq/IsJp4ppNonJHttv9DnGdfnHXlSMWIgp+RV6dQJMoIp6wEcd/ovNEVG1oSo70+P/o3EB6+TE5
qv0uWS1CMnvG5ZGp7x2HRdgGcTzhe/N6hee5+5Hdw3soLxHilfioXDKb/WnodWRBgqXoEJ/ELu/6
jyUWzq0lm2Yi5cCYzsZkkYgHRXN5w8+WbC0VKvmVt5PVIaLxEno3AW8sKDr4SJzIFt6aH8Gmxo0H
eYdCEGXeiXUy+rloeZQ4JRZC3FUOThE1VXAWVekEXw60HXhvWqFWvkhJo9861t0TWYjzC27Q7L9A
7qMQGGnxYGb29l7ACm4B8GCuzL0hgWl6RfoZTEXujVdC+ZcCY0b/QRH19h6dEBMCAo0qWlx9ptfV
powSii5X3THcX26vbhPi0nxMDEXLhGUPv5eOowTI/jOU15gW3zs2GxxNrM1EnttFS0RkEUYQaLRZ
9pnWJSPG4CCGAXrC5kIRWIxLSI3uBQhksPuMlY7mLVtCXKs+lvZGKKKfmquy0Rp4zJJwVDcD4hLI
YSWH7S/l5/GA0Xwz5bqU20JxJcCTMNC3dPwnK22lG0hCBGBSo85WxoFgQV6awHfbEe24qfEaAV7o
q8cogtnm87yXJHoFMJevCFICLG0RCKSjqskGHSlDLfRmkvkJPL9IMA+v+FrrmaItyyxyleQM5Eo9
0yiztZ44+v41ghGhPcNWhCJWWEcwrbzVt3pMYPURse7qwB70vSl2FjiJ2s1HLKCj+66wywMe3n8I
VIFhZc0JWQeFS/Z56BimCWv4xMsPcDGF+90TM8nRAP0jod64iZkU/6HiUYQX3CRjEIyHknqGWyCB
McSvTauSXxhGVSZEo94QKJANRspNpsdPJyziscSDd53nO0qGa8zsH90szNjhdMsrEKkmHTgzdgOP
QOwdznIZ2goHL7YO1XeliloY2yXyDMfELDQWKfshfwQLIu5mf8tcmUU/4kLf60VqIGSCahMU2++F
e40tZQvY6xowiX+3W2RJovjIJ1kPffkvvcEtE7SLFyRchyKnM/i1E5tI5swqBlMEnPkzLVJISTf3
BrNshyQwg3MvhgiYVJuzGztZ9TXu2XpBlpnC/KzC3wHUvLt0zwVAFjf5XceopziYenQRZbOlCB/j
IqWfUEl4WYFuSTBU0oGVl70ezq8Csoicubpw0xzRYcwXM1bbD5Zgxbs7ghcDO+jUMQmw2hhHJ0RS
arOK4CGSqUWEsRyL7gXc0c9WPnv9rYCbXQWbF2D46p+TmHE7RpUEMLh/JhFmxi7u6i1hrheSOOy+
If8TS9p2WavZU6NWAdQ1o/EE23eVc5VkP4yVCjuLLf1JaLFPpob0Txc3oPgPaAkhnxelrmFNhM5R
Kz2QQZ73wSZsrHC132zIN7d07ktDkJ2KI/HKYNq4R1xVO+NoRyF6ARAsd0rEiZQ1SnB3q/GSGtxe
PLl68Dl9CXtWCmfIb4WMPA10LXPuzksv8h5AcCdcMaCtHWeXCEYRN3x6SFOBv3i2MCgTpVYtGc7D
cZVn4EvFC4p3QsaZm0EsToiUnb1Gt6NHXBDf+qeoozbfj0fMYtbWXa5uX2tAg8uIFaceIxs0Cx5w
YHgWwVHhUUhH0bUKLezLfvN8/OxXepaRWWETamUrqymQHK97AJh3sTe/dG0b2eAhMqAj2yja05EV
vW2wIebwwYLexdlkPqbO+QVHhEjK7cGfW11lZwgE33MrQGrgwJnIRc3iX3BWuIKuoUzfnBfzMZrG
NvYfDglpDZYGNCjVI7nLedyCraXdvrwFcitWASwi0JUqMD56QA6jhvG0o6Uc+7uqrG++rrdhqHWi
8T43M5GS8uFn81MN6eeHUX+htijHKHTmT+YtqU0Hcbszpv0UgiuLsE3+uAP6ttkRUxdx+AtIOydl
EUy/TbXOzdYToJ5wN/xjrX8syXjcuL9Xq6dNuRZQV2rMSTDnzSvbvpzMTneeiKq8aQ4L2UL1mhOs
ILH6Knnl77U3+kTCFK1uFTM1NGeJ+I5ADKWj3XdFuiOJ6iiB/zGQnZBXBn2nbmLIFBx2Rqxl+e3L
c9ZSNavslKM04q1zDe8l8HaVvnv2pwtoe2wDtPArf6XB0lQVVzDw5w8sCFymPSQFK3cY2PEJ8Qgs
9t6Rq7dvJsHGiH9LMAYui+Yb/y5/yi67yb/jIvLNM30jn9LWSsa8Oi6p5ZEBGVxbmeIwccmrS0AZ
iAJ9xhtBIMOM8baUY77J7P7rjv31vrHhSCKxsUGfvqO45ofkYAQ1nvHT5ms6cTGs8FvbOOTJTENm
4ErcoxzuhJnLWEkWtZUmBtrviEZYMQxr1LSQtkZARtDjE83MMAOuwpfhMkapn9j17Q19hwmQhP95
4RppN5wZ4gTXQNCkx/bksYQejJe0itjgZ7wgQw0aE5OH5LU/iEefXiNwDNAuSMT1KtvV13QiR6+y
dHCk/5hkVp6WadI2bcWlswk59DK6PZERtdWc42iMCIMInti4Cvd6TpmegKMBFeHfqb+Ma/ouSSF4
qoraHbKgWhw0iBg+RRCvLsdv5f6OvZowi9msfYXpP/PfiBhoPIhR23J2D7Fv96tf9qdvbCVQTHc0
RmRVGTnk6wE+59/rcGFJ2RWzIds8innRYI1E1RspYqkygvMvs2UCmwL4AmIqaC9R/n9mPu4b0+IC
MNbKFcX5SNFIIFplRiPn6oMpVCK/NHX4IYN1S8cMDmBcaKQBiwy+FmpjE8Lx5je1gV46zV01I5Qv
sbW0T7sOMXPwrPrP7dtrVjgW01aC3h48Ga6nKAfIy+mUYvQyHfIGDKZtay1JqhtzxAXb6W1RTi23
mL0QZ6m5c2LDFrk9mCedjZMIHls27++Qp23Q9nrSZSn5UOuywY3ENLOxWnVM3JsPWT+LlFlflU8Y
+InduZUvOi/KhF8bMP67oescqdswWVy7AZccv3RuxfqARKIHoeIg1WAGucb/QHYYaVgMX8DnB6HS
+PAnGwbDdZR4NBvAjo8k/SZs37xGVEaydrnpUXP69Us6e7twtEJIgSd2bxElRlBeVMewZ0ZVkjQh
FQPkPyBuDqE8MlWMm2Vv9qntZo0CaA8GoZlA9GsY70tV82A2sJ7uw8G2OItxMqSyWat65sTNqbYH
jGsNAwAn/eAYr/5Hh50WmbjnVHwSWjt34paBDSNbW8Wc4/9Z4g0ENapRMpFMzua4Ijsyw3ZsfPrt
RVfM7sM0jW4LE8yQSpoeo9fiUnBPjtJlqTLczugJIc1YPMwp+6HMtesCvMRSSfbA+0yDr02Xcx26
7yhQraEViL3oi743s5Jlm08Vpl4n5esreNfFfGm3brHoVeBovPR5qk3nOUW2RSM6rsC3yqQ2C2tl
nkAimjNkj50RMLti5XRzYzegnGxTxuKXTkvmXjZkBneQutn8U2N6p635i6Cp1OKffc2LUzoRy9Wx
Ds/wjEru4/uNVRPJtvjuGY5x+CpuYuTpyZjgruNQac5U+xt05HFaXvJIRZaGlbs+pGhtyLRnyJyj
KjMcSifi0NALJ6tphQfJtZgqUeFVnMs6Pfmjwdb4MnpW7gwY6AaQLW6yNND/eScxt/8p8XH4VYOo
xjua15JwDN6GY8yrJWPKFAJb02JvMNzeIQHeeifsZirCNCcje5QkkbZYNzdjd6PzWT+C2BuvIyzw
S55tep1+Il2u7gQ54om26EfPNwF2nVZ9HoHnkTzNr95HkalkIansEDtIfdqnVdrph80P60hMUBD+
Yiw8GwY7YpNO7Hldz9VYsSyO5Q5bIDhjnfuBRbSr8IwxQfI51a3khv3tc4ivCRX+u5rVm7pREjMm
xkt4mhItAJcC5Z6bqzS+pQLNgYDF4phW2AnGMpRp5z3UUuqmWsnRSVJqGFUyEkMHf46qXa2wmPYN
JgpsUAdy9bvPyDexpxxa2mhLbhhbmIfOuF5qD01Rt+fXu9Z38WmygO34lAn3Lf8jr8ClhemlOthc
UOXZWs4vH14AQVofXKJKrSYWzGCJdYgXIckXfTQdZPDHFPe8YIlmCI8WY3sOCV0FifWZkMC9ueD2
jUMPZE/7mf3EqYcG7jjTTnsQt4rdY//7vr3Mb3Tqy+rbiUxM496i+hGolh+/krOPj/l2M3VMupV8
9OoiRoYZuf0zJzZl5pFfXqpKN1qpaTsqeUPIC3znS+SNijzLKkFLpdg6yfZsV18urJXEd96kM8Zn
/81dKDWCWvH/j0Wv3KkBlkxviBu5JoXMjm0ax+B9+Z95UMiMKVEotpEikUGytWkDzdKZElbSbx5H
yJOOXPsEwYTce/pc4rrXLcj/LnXLySY9Tmh7dKE+XDLm6FZ1VcrYycaR5AQe6cDfQUfVW5Vi03TE
X6SPMp0ebDiC7e+4gMWQocrQTRTMoagUUH+bhmgHt3yBnr82cHa5reVBjg2/6m7e5X7JL5rflQjT
LJbKwd654YxIUPW8yOUknHvtjWYdCk2rsVBArqu3WjyaSRRev7Zuwez5fOIFuvRG1JOAns3VvLFf
Ml0JmOfsCNXDUbZmpP+Xs5bytNSXV8dlC90qCVzbAsd6EHjGSI3JyLI4daHXA5saQ/8I3BTFxcqY
u01PGw6uFzBx0QtLc/7QtapEQj3kjgAUejIay2GvS4lnACy4GYcOcvv65W1x9cXhv+OU5up/4Vxp
II0cgrJaFZZ7+WE2q4m9Lm1bbI5Yf3/Vc7CoM7As3qDf8oe1vzJ4AmyiEcBqVhzpE3sKLHEn35Rx
f/dT3ATc1x3C6FVVQEOg9/2fO8Xp4OqhYRSYbAzjNr4f6N/l6AeASh97g7ZXALThORw3VHjKPiUn
/E9zLwU/TlKvs00DD5lQBx24RamoGKSq5+XdJLUM0fbaHkf7IX357cgER0O49VOHff/OQf37byhG
kk/EhTb9+Tc0ZfGpYiedfNjcvZ9RrDaALrNMC09sS5pFclsMQqD2vyVX+6k8TvP4TjFz5s0WbxZ/
25mcqJtYPNvL9SxHmCu+0nxf2Sv8wh56OH6YPxHj0ZqeazwtKWxw7l/35H7Fudiu6K+Bxf0XRqJb
zgFaqcOVIz0RMnnC+dHlKTnGBiAqIGifSBtoudE6X1AkvQqNTVIDyXqWNLXXayNKtHnze3ISg9rb
pT7lJp2rmxD0hWFtlvlBWu+NGFoeN0usEzVR0JWsCOa9dFBLC8ft+2wsx4uei/G0V+O8O29rE7Iv
kWWrkztFbRVjQ4TZ83DQ/altatIyLErMr4EOqGVPX2Gq/RdyW+NuuVlgCSY2WjAxrrXbkwUcYH7h
HVasZVFIM+l87kFfPPWd6HGBzmgJ8c7Sl5mSmsZjihe0GuqDIyJEixGOMG0nbad0uuuEXh5I8V9e
woKxjV50eOepVqg1jZvzhnHafVzw23HGDwXr7alX5W9B9hlN/MotDzDouc+AU96gBIkMYk+VWLdJ
LmE/iqUBtC9EVFpsqCnl3yt1EFHF0d5mNzxyYhH2Y/TQEKGoSr5Zy5fRxAXYBYlu3gb1FG/GGcIq
lMxoLhGfhN1qkg/TutkeLNjiVDvdgZ1x2HoDJdh+3kfmyZjFHJjqnNaWcHnfuI+6p+p35wTknu+y
eSrC/BFuq719tgMRGy1cvKLd7WqyRYkFNyfzMByrekcqXlcbfJyc/nBt8My3oHcPqk1bH/Hd3MkU
G6zvYcXSWcRtbxHTXa1NKfwcIAm3WrxFpH+MEU6GKNBbxIcoXXvUMhXDYp48pcqSJ65lmra6+p0l
3xMzRvGCcImRiBg96vSRCn5T/pdh4+u7KZ03U45cd1H/Hzr2S0IujbEJb4/YkXWaMwE/x21NtZ24
D6j5paUt43jP3TY+xs4+qfLQI8yNv+3CFiAp7xZjsObJwKNWV8WxoaGLsugZFwv53+ti7LiLovh3
P04rrjEuH4m+3xMR2w9alv4c/dOhhWkey4oFVeOUCkwFuDiC0LiNm2w2mHIfoi21hBcs+322j0KY
q3kB14n8h/dNvrTKtZ6FiC6MUZYUPJT3oexbU47UWnn3qQhDq/9NFhFrhAo9nAzO5pTqW/FyRyS1
RPGS6exzPdn8FWXEClP0ZFmtLZlJDDB4xvHXPnOjn4ZJp/KIkCCKZcWezTUdoDyLNzqRua6UwD04
lAywRW/poO/SEk1ybuZkqlkpep1NFy5mHCG22StjsXpAxNbpGLLCZ7+DXjRBQbcDOkaUkYf7mpEm
n//E++WJL1TBRrx7N5fZ0/o2QVFTwFs6hpf8SNm3Vt6i67OEmPv878fe1kf+eud1k8Eeb25yQpZk
FcXj8+g4j1EJYmLA8N8qIlm5t1JknhzNf86FomoUrXr71GZH/rbkWmNfWqPahKMgQBOpb10vYdev
OYwMKOUIbegrwG4pc/PtRfbb08KnnvSzaMjcPMboxr4nO404ew/WBTlTyqbQIssWGbrX+68hqWmR
/OiX1+pvJBWyxLJaDI97wWSRepovYw+OSzu+1TI9z6vAgPu28RDMVklngENWpO9Y7jkn8K3vcrC4
jP1LUsOamJBwCxGORNtdu7YgpkgrH+Ribnxmwo7cw1XiRWH9GzW38v7VxWSdCRengCAqrgLHk5iI
WoRmal8obPDe7KIYVkeYTMKT17RbH++gM0PZzufA4plj9ApQoL9GcHP1uqgqtovHBq8Up4BEBS0C
IUTnqfjr93Qxu0Pvd8aVtW6IRgYtC2rNPv6USOSp+hY7Pfh1jTwDwOoFZdoqC4v66HR7YVScqPeI
i4Pg8MR/YtbAgCiDn7Eq7DT1wGzPvUQdHx9U7+ZVbvc4C7X6hOIDUZaeftOEgE1FZmi6HZ2I0Uma
SFWdbOANliywdPxKoujCj+PzwZkx9o2xKDKQeZChFWQIaoqOeACfvbx5TfgZDfTLcL2iaa9waYM9
1pp4Atnek5Y0zgbmPXO74TIMcHD4DRi7/O/zkblFsJKL36LxrXznrtkA36b/hEchNngAKrArKT4O
AROnQNrLx/zQcVabgb6WNYKDcvoG5sNvOf0g1KT7I8lW+eTyEndN3JNPicmA2GqPY0XSqgvJEndi
YVyq8Tm0PVuO/QdIDnRRR8q57rCkNjeZAMDRbyXviKjaoFrypI2EAmPkz0V9NECvT6cpab9nagw+
BBpRvM2kVg8L6CcIa7OSsXy7yqlhux1Pdl4j8kPWDo8z8wBXij/RecJsCwciOBQFt86lQ5FsU0NY
G1C5Kpp77ah9zi/oSdhK45dAZJ8NOWJeEU5xcS+UXdOjSyGKd3VjQcpkmR1cWQmdT6U1xBthqJif
fA96bjHFOyUZAWFzEm05TXMsvbdDRNy5Wnk7XC8B23wfS/CZ9aLhUxew6wNVXpxTj3fjKPAurCzA
lsRM+3cx96WJVtFd1WFO9rOyySPJYEQuVyJkviRnFb5bkV7O7qizKiqjJF5gjIp1vL8O//8pEnk3
AsqB2HSSI/1ZooR6tnDrU51B1qJPBpNG/fsi7d8bKouzkYw+KYTpleqtc6F8ssiC/VOqz31EqsEq
tbr9Uc6IcSS/GDAr7bLd/dtbIiFdTIK8xGanjMdtcAOltdLvmIvb8KrYYjaSNA44te0kpPrDzKOR
9Qd+i4501bN52n1F5bF/9lrAfsRwa8EtH7OM5C+pk7zd5p/1FymsnV4txqOV4jhKrD3oc/09/Lh+
YXUO2WYvjQLqskmxWUmOZhGbqg39pL+mcY2760ojQo6Xx5z19STclScoBZ9d9W29iGvBA1c9C8td
xHw5OvDUcwH/JzA3vgSRt8vFdvYR3ThHDdGaWaMZfy5X9UOo+jbQ3tqFsKVdLdsnR6niWW/du9P7
qSCxefrHn9QA79IAoetB2G465skEgWDtYEKccobJya9jszwJcHSOk6NRIJoWCXr3sO2jUhD8LHA2
5/KtNhTdXyKIqkF6MGSC6pHVavyY+LMLfCcgFdgz4gzw/zGMRi5H46Z189MLUlQqdu0Wqhc6DpQs
eCj6mkNcahAxu7xBW+ZADP2lC3LXRou+I5ZakHQXxC1SnH4OVe0plmQX4vNXzaBn4FeqHRqvt1je
DCx5UK9rxBlBE/os6BJBd6XpVZSfJP48SifgnokYG8I4keuVW1yYhizIGqLd04EgjITVWdz0OJYX
u4h/wg2JA1dxwv+dcdbLLmSdvFBUdNgKAcRGq9u7aLIt24XWcGBPO7R+eIgAIbMgnu9hAazhKlYs
UzRY0KGlRS3Xl/Xt2bSfF1tYjwv91E5NPdv6gh6UGNfPetKy0o/I6vweiG+2su+zE0uK/9zpuhSv
0zffgkp3nwcBBzn8ceyeIYGOwK5J0vPBoZ6fWtp4+g1tazv54PspAlpJ6S6ALBiiHL2pvUM4ZU8O
gh1aDVEivVvWm/B0U+PRfXZL9OHoclcO1+0hLg01qLbpJkxUY13jrrpqBJ23eBLzVQyzRszgvi/W
WMsZ26506f+NHJuABp2svNLN7Ec+7FdvYwhOm+TeMKo5Z1cKPShRQW9dqGYgekyxGdgdSgXDcX85
0nDTaUf6E0X9cYOA8hs7hCvStjWsC6zwMK+Gd11cJVfUykrbuaL+oiZikF3dKn0QCTKMEXx057R0
ZBa8UREtXaSBMhZZG+NpVjo2EMHXOv4w8GxIFoo1szDD1jw7UBapk5y4egpW0gbYOjgiaMcr869k
bfcYxAl+KMPvk6JjpN0SVpByc2YbZ9Q676VB/A0hh36SRZpwycNkMjfznfIWg9Lp0TpzPr5DkVFU
X6jSzdEgBWPdDEozijk20YZTCQ4OHfLdGBW8oE01GEhwiphMLCNlb9mzHqvxHx9wum8tN6AUu6q1
uaVTXY9H4MzHrQrteBUiuge+A4zrEv8yj8mddsFDgIxvbfDEpPf7F8yzIYkI58u0gTZKwmpXgb8i
CCM7zCYqOYSPjk8Jy+XdQWXpDb5XV0S9I6HdMBSBUiTG/MvWNKlfizmfYaT3BEqJcOzl17QpptJC
BUdXiqXxLeLZZ95TKdNT2SVdrUb2cGCelMX1uE3WuV/QK+h9I+5QlPZ9RgiUc1ruNzwPnXKRCIhg
s1yoMOMztottxN3JbDr7EafeWVprOOhev7Y5pcrMYnWxgoC3T2vgOzYJjZiFt5fkbAIGtnzyn33Z
b2JXuSIivquB5r4sJ5CQFr4F5MSmz9waRBbyChz/qI+uFG9H88ZI1Y3ncHg+atafBIf7cV5U+eEp
xs8n1rwfCvfKvSoMxxg92qbKjwm45PERrE4Z8Zkkel7J6U9ShAEbvcZVN+k6/It7Kjhx2g4d+MEf
oeONhLPtW4RnD0/ZP8Yyn71UqSuzMbeJ7ULUpRAJezG77tt0n1tbhvy1iHxVrPnDXxNe4Dck58Rk
fGP84meApNpLfRQzLG7noT3hAwiQVzb+bk1WmTENwGFdnLxQCm+ZxRPhkP8h43UMGjaa5YAdesEP
bBBqlqmCKSnWigKPAfQQtAR1Tlem2WOdMW4v47MiKwUpzT63BeWGePyY9r57OcQFfgryncOgBi0p
5o913C07TQxuTZOPTRw7eDqZ1GiSn70adf7tAo8rXOCIyJzyg5jjIqPyjn4HZo8vUQUvVMVTGZAs
KFpyGrHzneVWTwdx9tUnB3alCQ+hkdl6gI7Unxa16e7cfRIeo4hDrHyd09gqVZdXMU1j2DYM98jg
Dx2YRHLQBReDfjoBPeoqJO+Nl4LRe44x7xE6ckkogC3DDTBhAc8gITJx6ZYS3QOeLnMqcl4cSdq8
hHtJ5Ra/aIQFflZzDfAXxgDhTEH21WTfmHCe6fB0s7/0Mt89PaElxPe+W5XJks4mI2FrqfFKNeMI
Y1zftL19lsXNB7RO0hu0kGpMPNeTyDJ7DyItVvKYXy/5V6LNcFoMQFdkxiPDERsPntWvYEuEGY1Y
MCn4t3alNvdv8funaaNqG2nO9UtG4pNaLN5GG7FUZTJxfH1Q1ddyAZndd2IPl8uVeluGAd73j3CJ
T9YehSCKOEc4lalTgpyQ5YTS4twrev88jh/FqDPos3gjHASw9q+ALW3KNyMcAYn/KGaEun7aekl0
R3V6wbiH3IbRHDIDMK3hzDriApfjTmJQs7+ZRS3Ax8tMH5E/9oqvJiCIBn6kCTiztF8DO40uXhSn
pgTHPIotG7fmElSC6MrRkPjB79K1dnI0+CkjU0t9vjsTcD/SvVijl6aMbtPuRKqT8YJN9O/h7LUM
2K6RPlOXRx9k9Ae5nxQ2IKIxNZ9noImCrlQqXIG1skLbFDSYdTq0KVvMb7aIaUR4TFF4F8XMwuKE
UfrLiCknO2c/XMdedKnx3B9mhXkWX3jD+2ccm5uI/PJrt98RNpGttAZXFeHACK3Ss5jTPeo7ZcO6
bwuHaUKmocjKaIU4mSfwA1E5NMb+zGwkAQNs6HgwA0/2rfrBDInzk8Ho4WAt+kH6qHLbbx6A8Fe0
ls/M5X00mHgT3P4S9qJifEAmegMDQqyomz8JXKhmElNy0ZmSMUfrz81wYBCGFj7VaD8Li53n95i1
nhfBHxcq31UeCs89OQcfXQEsS6VEdkZmqWh8Hkfj3DKfmTlXQw9oqKMc4Q6OWsd/7UQb3kPwlGZf
z8JXyrui2ST3pZfzn1fq+QH8J2Nc19rAWTuH86I1lOIJXAQxTjxmgq8QfOb7slpfWxRzTlJWE8Xe
rOdp26e3fMekEhOeceznHNFwTV1epEEeK/WxUJh/H//uanlIbUc4eLBi7zyuovHC+TslJup5WXxb
wy2ijUIS1cPviT+Qbq1mTMt4JT6p9tcPoHoFYfVFWVrEAgKaToTrKtMSSt00ceZXEiF3suUSZu7z
lI4ge/lPEdDp0Hlkp6M1dRsopzXl6GYtjOAkza9asLuPl7YjEff4DfgvrErOo3+7EUw4JaqJZg5W
vcMi0Tj0oI3iiGJd6SLDkDkpKUSFl3INUsTg8A+h1fIjkBQzeBzuZAku+P3OyiRaG5mXdBg2qyK+
BJZ49ZCQ365rkENterV3x3e6JeF7rlaxcHm7OSvDRPn3fhaNRthDuXFLQM94wHFU7FyOLGV1FYnw
mTttppo0e7+kY5l3eVEhQ9r0LqlMZN64ary4t+RmZTZnJMArDe1WsollT2Q2tLHTSUb3uIt2YD9C
jbcfoTRnemvVbs+XadFHPtcgcbDVaTPZr/zkjIqTn6Wb8mfQfdFbDu2oMl5YnhyHwrhZrCPyAMd5
4ysQDagII+sSR1IjkAhhyiy0YQJx96Y8GawHt4+OQIEOhVANu6833vO3yl4gnFO0pPMlX/0+JLRF
yTZHdFkodXP6X4dgZYLIIWlRQGAQu5M3tb+NY1rWIqIvX2br4ZgWX9m5JdIh2bViUWUYH/MT6QIF
qIcBJhzlWEuN3msww2NXmGwxVWEgTFr5oBvGPK+DDiqIEiqXQiiqrpjZyDBBXunDtQ+MWfI6Dx1t
ujgF4QFSysaxezwrSGx+3UA9UIedb5HOC3Oj5Q5Z8unGdqOAPUCEtXwfZfvm10Jx7WluwaEOWNLs
DsYHuyyohtOX1tl/hdtncF2tr06lS0dFQ8MD0cNYcI7rHJmloFln0O5/PNKc8EMzEBlPkG36SKjL
LGQELrOovx8l2p6RVWnBrCBXykV9NAZUHAXKea3hA/L5K+0cwoJDNfWt07/XzMpgpMaDtLfTiTc8
HMmUwz+de1nlycYbuLACqMKOQP8cRDldmslRlLm5lLT1pByxIRSOYiVuLCX7rLB38T04cLunVnxL
nS3MdrybT90NQhzFWxVk3Q1CbCTkRgMfD6gPWZ+8i1Gvi7m7DM51PfEHtV/0XJVU5ZTkK22bqVzX
MzX1WEPwYQvAg0NxeFKTAj2ED5w5/Mo0E44ISY9Q3jy6nBAq6Mq7O5rKad+kAy7sszN6Cf/MHjJm
5bkFDkPRve7OVY6KSlyYUe9FOZQO/LKrttONTFrEPRR/474nlk3zriYCaV4v2DFBn8JN1Iph/CZQ
6Zk3oDFPT3UNu30PUQjlNnY4RuvC5fh27CgZGLcxQVRFk7m3Td07jgISNnvcv96Gi5gkyieaR4KM
TWK7Y/e2IQrOzzJCGC19GA9JKo39yCYE+Tdj6Ax95lDMLOg+Xvb1ZUUPGsZEbXWIH65wencwhZsp
3cT+jE+e90yOLwlvFNTTDtWt1mEuNj/x80eZdPeYK3pKBJUQJuHn8NwcdfE3U45HfLzeOUw9+ka8
p3Iw7jikEidvReVwx3gYEB/IslkFjHz39awfzHDpZ90Kn9MNdfaJvmlbrLH3rJ1jlebO3BWgxvPg
YXtVNl8wiKayGlCTOFDzGzfBMaxk8axso7y2XqVxB2C3aieb8KILktXiM03O2gyPO4Ipk6hGue9R
2qlQZ8jOqUI+VXyu2BOFVcLs8WoCR2ESYq8bNNB/9nJKW0xgHZJpWjFjWpwBIHT4zQ+QwfUZrQAo
N0+YleBtfL/cRuuPaooKpwc/lbuBOa/F3mRm10yjCSqcqLUw6XKvEexJTzC2ueM6A7amGH5u6b6X
SdkY3KCv3rN60mAqLmQccGWCI7RxPG2ueQN/IiWu/dRnl8uqS2tmUfli4fgHSnhlhHkrecDQnPXV
/ufeX0y433XOZx8Nrvble2dWAOTKq/6COVu3WUkkBy4igu/B2JMp4xjsZ1uafNgHAAj3N3AMIIvl
XsFlCCFU+RN0pZuRC4td3hmESRF8+EqM+alVo14cpY/KFxRBnBGb5a19S2gdzq44VENu152YU30k
Jfk/lJSvAvUBl1sSQ3sg7kL1cAy/h7sua3Pfp6XlwJ5fWm6BVkS1sf+KZt1feaUrJVW3BcF1zoS+
zpb64ZUn2DkgSYRvGd5WlOYDnuVIVvj4ihp03m6soHBcRBHinY8Vka3sV+j1LmDKL0qQAOVC81oi
VlNoOmTa5SNuMmXAXJKBg5IEPvqkwao+YHlSuOJXbRmYGnGevTeZvdk7Ms7lR88wnPLDk2v/rVh/
5SD8rLqXjaOgjjikxrFWJunY0tx3oSwzo+la1S+30pmdoz9NASoI8e2Qe+s4qRbamz07+i3kJ5Nl
5I7CM7u+BxAuzeN4T4zujXvxWF7U9L+47BfLLwogKNMJ/cDpK69hS7HCfOS1ZqGV6LHkHzwlWVJW
aFh+aTMFT6EnEsQhkiH83hSapAhozxrYNBhx8Y4YVQ/sFsLFkb2de79zzW4Ap9y0YyYbQVI1p5MB
rVUDtIbsjSnEzMm+44jpbuupaiX5tstnTMeSjVvjsprxwmY/jwjnRdKW4c66YDDEMLolsSTwCKFf
r/M1Oq1x1yPl6VwiE95wdu6ermxaexK2rr0PUUIqCAbNIf8FjlsuY4QUaVWfYmewKxESh1+NTuQR
zcCrktn/BfW9p6WAQ+QWqFUtfSt2l369zxgCyaZz7cI5aaLIbEvsRJ9hEYSuf62i93B+HrxQ54cp
vKxfLJB09oFuNc2x8Rfp2PQ0i/wXsNN98pTZfYzaHt+/lXN3hAwnZMjr7f6eXSVtXQxhGlooclVy
9+9pNL08BF/Qdha4Off+ac8V1Zr09tJ719UU2UmIaAls9M3LAdHD56E1q32INt2/+p61a6KwU80u
v8yF60R48nQfbmyZYRRV5rwZfv7rkCGhZKQ3qhSdKxTOt83HqWvlib4QnBzLV8cTVEenRpF8fbGa
cXXZPUcpPXESqBjYM8DqxIXbNxl9lG+/c6vJ6UGx+G9na/p0EEaSLnNSXWegcxGsyoXruZqXDUwW
jjfiJL6ohtIwYBvS/mp0OqA0VsyRu/1rHT11xIUX95lJhTo/VHSVF+RM8CjlkbaBYtnkCYvZgeZa
FTPs2cGpLZsUIuCf5ShWMXhgCMIr+lqJofGWOxxzL73dGpqB6kTT4glYcT4fYhR0fTccq4d7Cp0v
diY3Na21xE1CbJCGuZE2ok1yGegetUcSXjEKg3gKQlV4qsHUH68TGtgWWfaZ0yUQLfp5/C0XCx7I
974j6N3FmDeIAumysheWQOllvqnbul3eCSPG1XUK60DepCsbj+my9ZorKij73Zk7YjOMeXdOyadV
pYsZdO7Zvp/JzaeALu738cP2Na7RutIMndcsXuMpAT4VnJzt1r8vH9ydqxbaavHbqaDX/kG0avOx
Y/y2GklmNReCUzxGxKZGq/+bSFaLT11d27gmyibn4xt67ow7qJkJa6NuCML5GJm1SvLimfqnCTJo
wp5GlBYh1kNMxODaugwEDsPS/80oEWDJXcl1ErEctEm5RplSLVhmI1FQa4Ay5JyBjcTLPNZ6gbjz
xbFbU3CgjZMYWVd7wOIWN+RGu4YJb9nebrEeVOJgPOkPjmsVcjenLnIPafupgULgtZtlh1DlFcDy
CLDXT0Urx46fHYqncRtlOtnIU5QDEUzDJQ7C9jpEzbueq7Zqt06R9s9/G/J1/QeS4gyZEXqsd182
TxcIf4OceaPxyIyWFiLQOY94wswusz2txWIE/ppu6Y/nvxjZeJISmJ8LTt8nIu8YwB+bst2H050n
STa3lCIElg5NXs/YxVvVGXlNlZ9K8bMHJH/Pn4TvNMIF6hVFJQwQI7o+H5zxg2uIlzfpn/TmUR8m
Y0j+fDAN8VCm3lazw40+FqYwWWWqB9KziQaQBNfSn0myiNjnHRYuCP9iRdG/Eu3XmC3iVHRFIhl0
oTtx9b+Te5r+k8nCDVe7qu+5IzznvGFvko7QzvPl8ILKUXJ/CF7LOL3VY5DRnln00EawviMde6sR
tWpXXh2xW6GqnfNUt2FWtH/CoiUKI1eboGDWDmWTBa4ZopCYkCdJmrFtu8zTCpkUjcMwI37KF2Ds
lHIbZba2ckGxNEIEtkWmUW3FvhDYG+TbXs3P3WHIsoK/usL6CBKiVYHePKnGx/g6kSWvj7SYX9Hl
s5unX4kvYvx5c61I54UazLIQUA9Uy1YVqODP+RRD8ijvdc50E4zs9qgNwoevWzEI0qd7rH+eWJdZ
TvHkVue3Tycepr+kz2t5jEU/IktDLoRr0P80Sd2hlvtnXmquCASyUgZuT+MqyeQ4coOR4mg5ddwo
K+Siuspf2CTSDsUDoavf02e3cfXnf010Lx2pFgNAAsOk4vL+Clsb1caeSxxAo7+L6TZ9UZNHWgOY
uIk6O0HXBzPILRksvJjrYFuAoSEL+a++714/zHo0mp4P3hzXdydCYEAfFuTr+l7W5G1082J2rVKZ
7selZR86bpyAGPWTb+B3B7dNAjiGFoUfyhOkzVUDI4pXJdt8wUMdH/z0MT9y4nO8XvG12AXpfiBV
sVd/lXvkMKkj+dpwfCnDCdFV1pd0G0mDMuGPUNW6XSzkCC/Ls1Fo7ozjLFOT7/uoOFi8fDPte/6v
WTlff0mLYrIrJatBujSi7Z2iHBhKqpFFFw31wvU+seIYiFYguo0zVoviUDNNYPDnzHbvnzEqtCfn
A58dUJTCFHVSF3ktb2MMSOqk89xq+YCIPKdSohacFV+VsjZqhWAjlbfuaVUDNGP0hmJKX6ebStMB
zJRtp0SNaX7C59OdbKAQjAkHd1Z4PtL0FAjg9zPAtiJQ8xnlDaL60vxHHxfqACeZEneTofFQldzi
XLuzUipnoC+6vdC2PkIo0sLiER1/fA8HzHXU3RkkxCjSLcj041UsY1MEKUzl5xIQoC2ZjNS+qUwR
L9wCq8iO7GWmhwhytbwsNtgDby7+qxKU/PAifIz/VUoIkC/6Hp+SlkoekcgZbyoCm+wMrPq2VWQj
VmcEquFqdy+wmaTkiAo/muSpr3bT+a+3kzWMGHNCySh5byuKU909h6QtF1jlsV7pPml/zz0GdrKS
VVZXVkgElpaqVEa9eKQAs2CL+6UVu8gFmBiljdZOoUvB7sJEu4ck5DgFyHr/gEEC5f1S8B7kMMBB
e9/jMGNvMh1j6QT/LHPNOAfV89VNGFdOQecporFmj+rsrEF+Kc+EwHliQ5okrBPwrOGSduBeU4v6
HcYEiiOjRd07WrYLh2XHo1RiOGTu49CI8PQcpcdnQVbJiZOARsWL/9ZE5oMu9WtAupsxl0foE8t2
uHdDU6C4bBNbjEavpBG3bPS5Wr/e0RzZs0Bb2GMKoZ/KSTHpzz2GhZlEomd8R7waseUIRGOqByn4
2s4ClkLmeGkg3o470Ke0uuWFd6WvRI013uAoW6OTw7bW+D6qNd6MFfEV2J4P/pnz+7XTIpawov/8
P0A0CzWiTF4uCliLUIu5AebK1V13zvNWOWs79t+eAgQrvMWXvJxk2uQ6nyAZskHbu8O8aRVTwsUa
K7FBb+Y36TJuIsclCUlJwXmuf8QvhdEMOEcowp2k0THvS1VWfIqaDN3hXJcKLH80YFlI+2snJ2c9
M61mlRJWe7gYC9uhtSz9Za0yHf1lgimzTC5rDg7m0o60BN8qDQHgjSTLlXW6UKpEneG+RkZYEByJ
E8rVK8D+Smc2jMawePg8oN9SSzAcJwWsHSyc7bMsuioBVU40go/cq0IHITUw6Wacex5QVoGRpikV
RGKBBPcWXtRfXQohEvCs2QWFfdtfOyq9rwHvlRen9dAe+evZHMW/RndzKTPHhgvZQBFSOx6OP84i
ObOt3rLuf3DP2rKGyFvaBTzAN/ZsOTSff8w4fRTqf4wLqhTIF8OtlHjO+ns2VhcwnVjGHTqZjtqk
0vhewN7VXFCmB/+Z+RCWzoSWLi5OeeXuROPp4QYC05tyCsQUTB73FJOFX5BYrIZVwGL+vVjpzyQn
q0/fNWSogu8a72EtjBin5gG+0Yvti3l7k2uNenzOoJ8G09MHHxjHzpQzqtoHnLDNwwZEzZ2JL5uI
SLSI0QXZJm9GYZ1rwiGcF2xcW3PUOGPBtyr12DgT03/9plskttx9XPTrTPi0uxaTJzm4NCPmCduF
8bElhPIuKB4LgJBmWT5rah6dL/oVVY5oUtdd6mWB6BN0c8EAUYWuaIamhg4Mz1RzSEBrntKXmVJp
TDLbbVsajebH0fAE1XdJhlbciR74zaCV+uflqdVYJ+TQRiGDe/U9fc0pFKBFsQWpSezkr5e/+u8l
S+tdeELuE0Mt8OWv5RXHzx073lVGNonbxyiy0LWebMpeviHGsel3mgVQ1NS0wj2jtk8oj64nK7yU
oRSOkTBRZ81/+SpN0EuqUoZW0Hgc+F5/K1FGicZAF1dz4/mh+LaoDdQcs2vxMfrgdsFjwQwP1xjN
9C+WCsDvtAENdxEQ6nx4cd5+memgai7v3Y8oNJrsRmW1coq+Mjemsvt6Gt6h/0WWjuqgAIkxMgSc
3VZ4MdeF45MvrclNEMKEPdLS2QIGruuc3OXXc1ZST1bMnUhfnZIjIrgnB2vbV2JSiaTp+4U2QbnP
SdumgjyzoqKxKlqtdqNNgzFDO1WQaVLdcR6mYEplRX2fWtGbq56Y6OiNu36LOi+RS6SCRnqOo3+M
sS4mS4/LyOuQRbPzsxeSr18oqJFCJDIYvP2Dw3V+MYUZs+qqVGA6NKJiiVjaGf0TXzDVnsg0MiXn
x93MyAa3+6SwtpAGwbF5hPatnH4oZ8dZ5z3NumSmwYXxFv2YVXPtAZzlf+NBns6/As2+WR18IHkb
G9xzPLUSmzQ2trLGl2RiXQgJlzZyJFJoXFtAYFU/stpR/9ro5A/h2eIYcmQArcqjHgc74bZbX8D9
ZqUiuUCdf7Ct6tm4/O8o3EgdhdYwf91/GYvAl+gZa3u1yBeTl2X0hzu8vJs56COkhCdL83mNa+rG
Wc0uAEttvfKBbofbmrwNm/Tok9HUJjOxAReaxWzQkB+Xdn2JqSBDoHCJihcTOOjIU+p4oHGveiqB
MhfOPa50pTu6KB8WTWULI+AI/cB5EfJa+cdDUj2wc6bAEqmry0RWR/S9U+JbBvYg4g2PFXcTIlRm
T5V3IMIsyx0Yr5eJZcdwYlk+uAj29RGPqmccz8+AzSueKluXdLbugctMJCtuTZIVVFJZSptwfFwt
PHUgCMk4k+1+UfQbCRJfgxf9nD2FLYUai2LY7z3i33J6bSYs95fo62JBtBapMe2kFermC5fdvB3/
l5TG1nwMlj240F+hym+EPvCXnzRGyzexcEaBd+aA8BXbefOSMlt4sl5M7wjMx/RNqoCGxeRf7TuX
XgycTK5Trp6widabmAmcO0Zkxoo3X8UcqDVwxlfZ2ZknAftaFP8cZ9l36zjIj4NWhy8Fy4qeqVeS
3TioLhzL1FoSl+XvcT/lEtA+FHE5ZIX4wgvTqRU2sTrO+gWpwdQWL30TargQg2pIp69pNqQSQHto
OeseeUXqvP/oKK3WXk/iIDHHF0HzNe7Iy7EE3cFNYG8ukpDr9GKpZYP/n/20vguoUb+1XpfFLzX8
e/p2RvUAEe7iZnqPQBySyeXdDGasJkNj+U2sNcchHXfHLXqhUgRtpCrkoqOjul8wRcXJztB6jjj/
M0Yd2D2h5o+PWWJqL9uU+o5Dk4uvKma+Pv39lde0hRKmLPveaJrHfi8tYc4YACp2rIYNDnkw1eL2
Iaf8NhzpTXhvGwYMyPMzjaA0+0sfErnX4b2nGdrf5fNnSCYbm7NvrEII9fithy2w2MWyODArp96Q
n9939kATcBiJ+NZzWZD1FzaRQ5JdG7eEgVwKQCpqcGw4KNL2I5hajjSlMY5fi8rjpTvsjg96Aqjn
dtjOdsLBdWQ0EQT9T5tub5K1x/63Bt8U/BQFatmqIQPSxRAu6Wt3THB/0mUVMDYpe0vEfTbGEFiN
YKUiQIE86t3v1WNeICr2Ozl0Njt8TfjCpBAJt7HpfylV1/Z4EdLxWO5ho9XOy6iHbKwT5cFlgf39
SKK7zbRny/MmMeq6fRJfozY/Gk/VinKlh4pEi6P+9B1uo96katc5+nWXiQ/dMtuFJY1+K7Lmxs28
wPZ+H8l4eqazC3U+5hhkpY8FfD019dAiiBGYN6QrKU0m+xgPFIOldnhLAKsRVy/vU2Aq084pFgj7
/d7d2jqJjlj6pW48rKIXms21el0cgqa24GXV+AJhn7uKtLnH7q+LvFz7VsAE+4tz3cELUOBvly2q
A2F+4EbDaCp3oYOElrlPtVhNPOu+lBr1KhzguFNLqwsFFL5HwyZOIyt/4wQwM+vcoLFXnic2iMho
3GJ7G6bPi4Co0Zu2Q/8Sg2Qgag4I2VHsvfO2Z9mJiItgIDreKB1fCtIelX590kMJsGjjYLO2nfIQ
hNsH+AJ0HQ/j5wFh7bderoYg51e0JlnZ2H2K1fX6vbS2gK4oR3n4LW2xtxkp5yt6QsRMqyZW0ygl
+c+6IbWTbO1JGjMkTSmJdxtgPBVEe2LOKvpkx4Alz/xAw246Ane3SXzpa7ZtayonoLJZSA0jBKUT
xo9notjk6LyKaZu+1W+5EH6poVd4jGzgtO+PXsdijFrUlTnYWLVocw9fr9+Roc948RJ44O38NnY4
k6DgzkjlkP2HuzaYEGWEwMdSRrtrrD8BzkAVnFYVrI8gorggj07SnXMJ40cSIDs7si8RGQWhP1A/
GMHX7TSQaWw7ZZdsZ4Blqu1ZtGYxQEPBN7c8E8ioZH2MSqayhjaxx7YJNZRgMZgF0COyYhDfLH8V
uY75smZdBi7HJeACoQapmQD70Cn6xn7jqb9NBWxP6JUN6rRmuJTCKziHUhWiPlMy09tKiW2WoDST
/bOo86uYnTrjCzFjkqEz2Os/4RBBYx9kRgsN5h9FF8+0TRGEGh9Gknh3eaqmsf4kKu2f1iGcnULw
BmgvgWlyvnqsAcx7PAYySk6h980iNW+Zg1zv3wVvAiegPSweGwrwnqoaqsZeg8E2VTRvGT0oeN9T
FK8oH+7rFNeyzsQ22MKth2hsH5K0pS5cE+eeB+/UsaiJvWqTgbOuxqQhcslvjvWJYZHOB8aQkOw5
hkt4akV+L3FdKxH+vW+w7FGKQIlTzJMe9+xF/Wh1fKi972d8jrSs6H0e2Y7t5gfUsjnNZjZx/jpR
uHuyd7rjgpQ3SSiPZrBxKD4p4vRP5DzCWgBX2DGo5K14NpfbimKF4SnQgslGtk9osG8LxeQ5Qv/F
4AKFibd1O1rVbFKvTCYN1NCQCn116+EfeKHC7dLFYTzJIhMT9PqAbikDn3A6aIFxhH1k567wxhuI
wkMzBVHcrBvy80OI+cT+XXWSapsyWjuwQ28I3JcsdlX0uzI4kB/mbFTIcGo1sWu61Y7wPGayFA5I
lj9uSj0SbOxjVZ7B454Uqz06RUf6relWrKv9YpaI89MUC8Uf6Albx5morrRNSKn3T3CR5i0Y1Avu
teCZQ+zpJBBIImrCWFa3nlPnZQk9vOTN1I5LFpwjz56LoV4gLegUAe4jkMbZT4S3WriEwUQWy1Fz
HboGkWq17FRbpUkqnOOxvVYO1K7bfLOTboTkhNp8LB7Ytn+1LlG2pvLqjjoe2vpC/Nbq/EoN1S8W
ShqL8yYBKbYYWKhdd8/FtfqxNabVoznXi15fKieEuDDkru2B64mivI8MKNlr4csxD7fU5lr5NiWq
JnULOqZDjXI+S/a9Pz6ngQkwuLLJUQ7sgJShQUIXshiI8jgmYUw47RoPPbdYHanh6NxXfsGl08xS
2uYW8Jt9XkrgwFh3WO+CjaqLASxI8WGX0GsgIImJgiBpu8qe6SEIYJPNl1MI6P4DTr/4DpeOUSCN
zqHN9RBPjRJ5LtGSMwJHAr2JUI2lxfuF6TH7yZMWhk2eUSov/Q2OEDWiHk4gGKmM0ft31AUf9nGB
cW5LQWFvoGbUuOiMF2EuUFkGxYrgeIW4hU8BN08TnVIlE10RhUIhgsEOIhSDsSV8muj5rTI0kc+O
rjtG7XLg+Y4WkDWuiOtTX5GKd0876xMtECzytb6X/HrcHL2SqATd/CaOetKrGNetFz31dRRamawL
IHHf3G6rJ2b1HdxNyg2GP5uNRLs0b4557ZM6r7BXsrcyZXkiquyjYOgcFD4jh0bhLzGb7zeWk3uE
PmLx4TWeyDH3CpB9d+yx8RbYDL+Nag3Y2bWGi7Ah5ChE0SAi8qp9peHPDt7oilr0rUOI9UZXNQvN
9PjpvIKkZ7dEjphBEHd91BFlh8mq/UbMl8H+AHjeOEXQyIgEsG50Z7blauKTEuAKb/kuIg5DhLkC
r5fsI6aSxVUvtJNDSWWybiSHmu7oCxm1EUnyALidP+55rC/Jr8a1NaKxjKd7/he1dr1uQzOLgb5U
XSBVZF+2Z5+Z/a1sHV8ZQiQPbSf+amiRDLkKyARY5knkN8kI/fm7i3zesjRJI4WE2gKNZQoLyRF/
LIlBM2TibnNKho7oHSOcjIHgmnDb/Sy2f9fUhZPkDNcPMH5RYJ2AvERbi/gEfQ+ug6egn2Yz6XSe
1nPC1mVzuXQSgfwGrXlv0gKdH9eXIhKwY/WceNKlVNtQGAx9YVsAM/e4jMk2Zu1bnrEFE4D7wOV2
ymNn1ec84EvFZs5Ycjs59rjRvaAXfyytigI3ncfgHe/9tQ29ry4lyWXNCrEU3HUAOt5laRvksL5w
twAMsYf1lrLoP0TYzjyrVDy8qmaJh3jKxz1G1GRVKqoyrC5sU+973Hzj9PJh8cJ0bm4W9KVvbLSJ
O7m43d2tFSoBMHzDYIqVh8lo+ZO/7+VREHQADe/5qVPhvHAeVX12okuGN09fbYNn6ZrbTirPFvcm
UUYuOGrjdHxh48cYVL0HJVSPsJSCZ4HY8eedQvhL/3LS4nUQbiV/PhE/PSwSie0MzNNiIf6aiQtD
00WtkrUyDKxihy/BaSPK1JPJixPLNbUuMZf935jDxMkSIbgkIYr2xTrtMwWlpND9TXtU2j0svka/
4VXJ4RuNs25wMYZKj7nK5vwEZDa/qlwL4pEHYxU7Xrh6fjWSIE1f0m+mxx/99yJWczQ9Q1f90ZNZ
QOyFSdBb31ctglbLunNAJWttOp4QAJrAdyEmsClHS7UCbFLHVn/GFlI/KH65+M2OnCfbV1wC36l2
HLL2qV5lRWn/CUIC7vT1vvpNANkt3JWzmzq6Vbhh6Orq6sOf6WsBnj1RhFyYYyi5VRm/eyuklSFc
CHMCmGIYZFWFP6Tah61scZZqK3mNAp1k7MZPdbzmZZ85pdpWV5bafICErART35DcaklDDPpI7D4f
KDqO7a329/e6dpE81WuarQYANmNTp9PFOcqWxYKIzs+kS6ZsgjtME4BRvCM81QSjJllnl5AvUhJx
PxbVP0HABMWvOMP6Y8m9FRjByByAvEvKhUS7oyi+O2oUf8mtiKPW+YojJlPuWt0z2xN28OYJNK7M
l/hGei3Qhdki2z8y9dQisshFCHATrZynyCJ7f0X8xjxucsZZo4MFriTTTc2kjAou2rW2Od7b3mYa
lEFVeXzmT9wx0Ibaf4vTv0elTNqq4rHa9pJ7yKWZ2TzXDG5F1gV9ec6n8fQBi4Nkg3AB1v7rFDxJ
Mur6EGWqaqXlw7oTU9o5m/K/3rbQ2Z7qzXLBOjtnMgH65fosZ7++2Lensh1N2V7WrZ9onQQ/3jGw
M2Bw/1sAZav0kbcc7JRKcdIuasImg8lcIdAqb8KgIM8dfnbugbKAqwztXTeaaqackbmzBaPb0xEU
Z4twVim/43Laxhmww7ERsDhnmcK/kCA064bQQ2pzRY+1IohEBBKa/GlwMCtdp+EFkCWD6QPSajoC
AHCQkHJYE8Q9gykbgU6LKhRmUGSxro4vUGDDzlFuKxsH9rJJ4+7GKT8aRnaX1aa1iS6L9UqmDfLm
I9Op7iVDdRYButZwMODdbK0CMXjuKD0ORBRjqSMFc0KlWGTU8S3Qi5nQcWrkInqH239P6l7ASlJN
n7vGB/PamREJo6mjQUObmY/JIGJ8TUJBFjDeArdqL1Hp7gq0IsHOxdUQMGljZDCk/gescskLzIRb
opQt8oDR28RxjVed7wTBJTqp16c3fBo8eGMwGFXk41GeuN/0QCT6QZh4hSY6pfANdq6vnj6PAfZ4
3Fxq8GDwq/lY98hgfPuOGihzBxufDZKXNUgNQmvZ2iXUFcPZ4ZnvnU4ARiP3RJh8bdQ3u8W2kWF4
QypRECQrkTREaGl3865SJ3pSKuFTFQax1Kc7NBp6Ll55Z/f+hGnQ+1rKxcCrUXsMfJxpKnvSh+76
ZYBhMdgE0jlEufY4RrIn8yxIg6jqhG3i3uhrniFzgYV18+N0hC9LtCCUncvzoGeYRUJ0yhSu3UzH
EhLpxc5n3JFNIEiBxmIlS7H2mUwz/NVrrFwIffc8cLNOsLX8oTGiWQwGd3pvGitM2Fr2kH71DEBV
uxErwpXi+aa2oYqr72JNMScLNnKmg6xPz3UT8YDeoYy4pCZso+qWDw8oS6rM17+dW1IXgdcfBJIJ
H9ldHN7m6XLaltvcmDYojHUlSGC/v1v3f0jUMTqWW/uTH0QoY9P2vlMEZk7ElJj3ItXkDeBTYjTT
nNzrEMDcH8y55CaVTSNbtmc/u3thI8EcYja9Ah7HfV1a/+SZM4XvtPYRLx4FGURU7ljOTJrlUOSp
HXJbIBPSN6SvKuDALZIRX9DbJFtNauutcAE4yGnagurzvgJL6ZspSYKs1Mxhvh/B2cY6822n7keo
jVD0kF/XqocMsf9luH02RIW24+rgF9miIQTkxFtcIUz2//kbdCXPp9r89/cVdLszlyUVqrAtDNB4
aNjs387A//LhXdEmpcpgBPm9SghrgTUbFZoQvpjiEZhgZIEpuOyQvgZG7Fog2Y5Xi04RXrObEG2I
mG3vazErFyO0Zm/z8C0pjXgMMZdwW/ngIWETK+nxx25FagKd/NksXxNUF8ZV3WCj7H0OkwUC1Ml2
5Dk7oW7mvs/W9wPkR3mgDFvUALP+DJ7nHOb382v21qdJ+NxdX4qalE02iRj5+LiCLKfYJFl2/f0h
e5C9bnssWyeuWgjs4b3BkubzUrru1/oMwdV/KfgEgYQhZRCV3e/zAMWDBHaFOudYakK7DAw/TQEl
IEuZBlSVMsqVnEhyOiS+H4KkQFKcnkJ0fVyN+SISDVyawgIDu6SSC6PVSPK9PF+CuZ1QM6MhmPaG
9OqJUMOAOvK5DJ33WvQgFyme+Hh9lH3DRoiNsI4Xg/2yHpdzx7dELtZh23374kYtSHH10GGrUPGb
YX9WIen/LD9ZObnYEz84KmxC7Icsuyq8spXV2JJhcHM/FAAAhepBX0uKcdjcXVLj3+gtAIoaA7IM
5gCbol0XmGd95hUzbyvmniD0/pnb6AQknkFy4xBcr9g4+3Y8IwnUxL0pClOhwiajH0JjrcdonLfk
/+gbj8kzDxQQ+TxszpLPcm5mw6g+6n4goGOFa4VAA58/Z735+2AHQt8S87yEnBM1Y/oVVjhfE/SL
DZMDQzgtR9VALVWmj9pcyMpEjpFnVUc2ah+FOTNCPFGA6i7LJ61HewlWHR8a6bkpL3dKoIfI0Xaj
4zzl9HFHPlCY3CoT1Hb941/PqWEMKjiSjL4M+tOZIMkuvKp4bgk19d2PGa7wf5rZ8vrFcxZTFaOI
MeRRT15vtEv8QZCSwB3xDQIWiFD12tqhoz0pUDA8Ti6wHbXeWLbGiCp7/xgDRZ2I3HkIk8cr4lrn
RDOp87fhwBvQjX8CiFOF+cQjc5HxM/8SD8KWPjl59NhLH7mShN5vUrxr9HTW1EIdNgO92SUDDafU
gsQo5FRe1f4AQX++odU5IWLyHadLVKvCHfkcZsv7PH/he9Gf+eFWI22ymrgjLD2Cy+KI9K5cgpKK
IndvJuhDUOpI4K/3f0UrgCXzlQ6un9xA5ZzSFvcjxwSUNSTvUsCZBgaZw5xW/8HPdgwmzzZE10tI
7+EQSsnRqjCGtr0e1Qtfg1bGQXkkwas8e0GppXNQrf6oXjWwXJtAb2a6EHzOv/bx1gs5jAW2xTE2
QobVIxIRId+Sryz1a7WPA80/EkVhf1kyPnqZA89tLZEUdAofoPHEcj5xYtaQQYLF46+GctujfBLL
KHkNRy0lNrV//dhzYr4ds2tL8r3TpjsNZwM/duTh/oQtlKOaDFxVOdj9f/zCPV7Utw5sorR2K0uT
COFYztaFUd1wyHglW6xl1k86ORswIQgwhIhVEDv0d9o95o929tFqNFVUniFSF7zxjAtCKBRl9rWc
QBQ4Au7rZcR7wj9Y/2hjDuP3MtqX4EIBSRU52DZcjrdcqG+ZLuY9SAF2RmoWi0Dqqz9dOG62/9gM
SflSFreN7njUHBOG5jQm9235YyizajF4EdEJuGwfVp8yskwhOuOiaF8TpNNH8uNYH3QskQtGbLZj
jVQisMX8Ojs7T/fM4RTHNuILHqyPFajAZHI0G+Jpsvd824baL9C4Zc3Qnr/bxyXGDwKjJ4Cu/Awv
U3tFtmb4feRYP33iss6EicuaKVTn7f02XWfwllixuJ6LW91vmpnFaiXLnZaUWAqo6Am/d0r3lPB1
/GxhFH31K1ww6Nd41kPwNf+sh95SQcOE0FOT2WgvTmfcgIFRkSmI/nMuq3zZdUfcXvqptSdQJp3S
Q4BqiBht7FYT06X6s3lYKHSZmlf9ICC7YfyrRhb1NnO76vJJxRlBxoxeyCl+U1s5b63vOkh3zymX
kijiijpS47tS3W/uZb/L9cfx4wSMkmoC2e/LQck80Ofy4zYM7EFIdzKQQ+dnrvGzE4nCMOjhAGru
3ODAVd986y59r6YM30CagR79fY/45OBKJJyplG3qvWyMz8vtxhJ9fXS1QMG9hTnZh3TRuJVZri3+
kBX3f8T3HerowCxLaFBwIKYBiOLCDt8bynevV9hmWmKjdI8YS4vwbVlq/RVI5F8WU8xI8+k5eSOd
eEdOEGy66WD/b5xCB5xBMlwIiWsH0gre37LS8DXwGJk5H65AfSM/y0AOznedLDJGM6NJ72/+i0wY
6h2a13aw0QI2dzhMUR0OYI/DLJuy6iIBUx3uC7LZg48/huT449a8g6UUrOuU85qOqeoa5zoFkkh4
mP1cruTLkxlH+pEkAmGRj6vNUxkVDMKmlJLrfRdaLTWrxDisPQT2Jcz3m+5+oa3x7m292rI5Sysz
VxrqegdqdEPMjuGM4fwc//Dx1DV4brmjbXTdj4h7+D46YSfFrbVHYEZSwheoN0djbIAa//sKRGZ3
eVJAEljMOAJpE7K8F3kD27W1kV2Qy+CEe1LMGp2ZR1iHT7rVkky7x9rmBgw/uOcDiKWFCgsIMA+Y
/o0GEQCShotBpeB+aQ6j8BM6QBR4XzugrtiokDO60ZXZNFHtajTcXmpg3EGCDX5mdASoJNNG2A6i
xcodHG6gkbYmg1DsD66GcRQxXk1KP4YE7AFO4a4yxjIjbAhv5Zig2vGzaP+zOOHeBVtEutT9FNkT
72Im3cNTU0z0vyfZwgtSOnpLeSalda4gM0lEotDxgseB9Qd/NN/wp7m4XV5xc24IZP3WOlqAg8x2
5yNs/sfjon+OssuaJYcACqMFZsTw0Y3/XoPG9dr0IMpqAt//qZF/wegZK98BKAA5oNZVi5FveUqQ
uGVqHFzb89rWsWKjiZgbqQxc/0obbJpezd+KtE75bWDsC1F5XNIuW+qkmtm95Qjt6Y2p7W6MfvNU
npAKG9ABWnhq0j3LESCIGhM8gphPKqb51TPT5290nt8uK/AOoQ2Q7InlfvcP7QhakF12zksnFS0N
IzOCgfBbkw+apceLWEDsQTbmMFL2VSCyJVPAlqFZPW+QaxqLSRrYBCHbE95DDtMeuMxoef4FwQUs
xCB6+ZaLVruuGJ2o15WcA7uXMYNbnennW0x2qyMY6JbHhfGuo0HfRjmk95dNwUU83xyY369EorqH
6Q8jV7NsGUXu8qy4AbzahWPCCZIzbRbT/ppzEXF79DTdRO6AnnCWuiUtha0Rhwej275+Al1jHe2u
RPZB93kZg8BUwWy1/Jjx9kotOHFS+P3bsOtGaJO5MJbQunItPFLYkzKTx/eLRJoFCt1sdet+57nw
E1eN6Qj1jk9Ws3H2JmiSh3yiQLkAnNRrmkiLQDvKOUEeMLmDn/rq5bDtSORKHZBsYfbKV9R9ERd6
oOsqye3CNVumfiGHM3Dx98hbKJqAu6aggD3Ww8Qq8aXDYV+9UkXSc+T2R61mvDS0275xO6yBOLlZ
7O57vaQ9KybYWhxT0vsKdV2kmudPmEAJZqECmfH1VqawQgT+pym/xA67Y0fMXfnoEkAfjeUw1qpo
Y1oSIfKSeA50UKuoxLBRfy03YmF2fhvHiC05Kpy6bbDZm0wYg6AkoEt0aHnEqunWZJCRjQ5OUKAw
hswnuzT9FFVbKddbXBTCcDdQ01uPntRBgwTXSjIN4695/Pwd8Q/ilK8qnYzWd1+2m3ZRvqxBRVFG
Wg2pyKTE0xU9d3JVZL8z6EHQN57RAhBk7bEYN0uoCSoNU4cfIhUIK12Zo0/u5iFF/pUm7Ap+Dq6x
ZZeYNaTNO8+jgVfj28P4je5hZQWbky0k7NLHudgfs9/pgUhNdo8sYv3T2gk5Yxb4baFX4sYylD2H
iOprkcaQylZbqPyYtxJuRW2F3xMrCVF4yDItSAm0yJhATXYSsk5EW84IAXkoDNcjk6Fh+YfrqLfT
shiJ5LD4RsV32o11zaxhrWFOtFGs9dtayGeCRKgb/OrjiqL0XHn0DHOGTfW16DAtJXan2Mjbp5OS
jTjnxVAcMmVMzbWuL5UByFEc44zTDSha/kKeE71qUOTAYHQIns5bC1CzkjIgO/2UTyO7Q5wqZXIA
LPfydH6/ZRgSAZXc26N69ec5B9dMmAphNfYP8leV/lmH8GECiVZy6kBR/zQHsoK4RotmqBPuHvgD
BNQ6N/lxrRKQ7W0G/w8O5aV7M28lwVl9EG03MFQcragMvwHllRH+ifkIEwfwKkElLmJU1QCxYJnR
5wwKLQ3NgtKhoqsV8K7pvROst2c33wUeN/XoQmrXoWq1ng1XvJMrmmQzpNsvI34/n40azQvLARup
0r3x3vfZA/Av3favIAblYc4tu+aja0yuLsuPLIZRu6Z3h2hKOefu6prp334xJXeLEU+rp/qZ4QAt
OH5C5ZZNuWgR2KJBgSUjFc9k95u0HL2Di0jH6F2OjzWKYDZ0se/KCGKPRjFafqjUJMNX5vToEI6d
0gf0bdsn2WzoqTmFKf1U2DAfuNsKl0wEjJ4tQSc97i3p1eh8sxIfYE8o0u4+Z9wpWw/2gLQR9leH
VIu2sPb9nTtq+H+6zVGQk/I1a1Z27SNV6GHZem2kdtehD3m9AnlwmOjvI1H9mBJxykl8sfGJhLN0
5jsJ/SHtU+Y1rCJ5iQbTuDm6DNRKq70uCWnnsrIWov2aDnU6yR7wfC0hCb3WOndOF9AunDi5rpJh
trstNtdiKqlkUHznTPaDfrMGa0aPs509v1zi6nPa3zVT4bciFrTIPgul49AX7qpkNPYety5gM7jk
r5CCV2Vfw37laqHprWYZ5Ync1+39ZqLa2UqWrGVUPv6BjOf/e/BqGVmFAyKeAVRoMnZkP4IMkt/l
5iDGivgSAblRX6rj8FpDNxGGo4RAWiRPW8DmIcuxcu18Xt+9KVyRhO5F2NI90xckLoYia0tHLZjs
C5kywtD5KFyFwpec8bqQwUcLScgTk7yT6HJwIV/z7Sv05i3tqCXseI+sl7D2yUuYVH4GoQ3peeuu
hPjKNGdph70bsN4n9psI8oZADa+ZThM6vz7zkqKqLNao+vGujZGa2etBL8J/1aFMr0ZKKpE+n74D
mujXq5/AwfkoZgErDja/bkvZFMcKGPiMKAgtteCUdO0Xz5CZYm2T/BgOpdPfLb/Pa1HdpdUaLvEi
YYTdRG7KNJbygaJtoAtuZX4fmtb2okAeGlk878RbUZ09CSufkiDByBWDOfJo1gEeFBSmHkDLpIfA
FHCbymPHzzqvKfp8AnvA6ftL0MdbWVTOTQ/6RaY7qRx1yLAZQ6ZhaLlgRsqoaCobx/PrIWg2eIeN
QNbw3eINpfqpYBNtNAAr5A0J8SOMJjzPL7lq1T/sy+dbvFRCGFDiLgH/pijToIwx0tzKpX2gJLIG
2w0SsbP649qkjfWeElgWSvZ4WuFu2Ve4FitaJ2gr+5NW7a0ZTT9/5nw5OkhLfWXpHBP5i4qOVvW/
XCoVKTwaA42KUGkoyyMWLGxx8n3kGWfrYNDL8lThM36/96iNemhkcsJYvhrhyk0KAfinxUcx6MYa
piP3bOKyk7YdiPVIZd5iP4pvCvqe3zGt+1m1sPst6zyubosmUXbgnytt9mIVwZfw2Az4gAD9NsHL
V3rPOTG3EUpYdygH9lumtUkSMavDEQb+j2m2d832DNxTgGDzgQy1MCgNpNm/eU3bcqH8Bniv9xc6
BLYoRZe60JvmsH1qK4jedwJN52UqgKRE6YhppuUHbctTcvc+z5pY0EItTUUb73x1XqRhwT5Can18
7JBAd+SnVb88ZUIwYtbqYjJQ1rPZhZwQaDMticcgI1+IbsI1eXSt7uHi332gWJyW48SNcsQHJANh
MT1agHT78oiph2OzNflpkRAUxVMvcEgb8gr3peV/7XVUAQ2IIlGI0D63DZzZD8etQTaQ0hHm8i89
QYgesWvNIVAdnb9Ds+6aqToA44imFfNtXXSpW0XChTPd1d4JP/3hSKjklqSSSitVfcuHTyEe/I28
EuobheIlI+ujY3NAj8yUxMJzrs8NlA5s1dkAIFWsuZoJy3cg4nXI8GBGXOqJW9/ZRE6odIxMW+bH
moCYiV4mGwGuRoieHV8VPpbzOskuoZ/ETUrC8mTzaTZ8NIacBK5HiYIA+L5BfzO0xN0Of598zrpm
bivv/2KnAaMsMmndtHsjDtCecaJRAVwSVe7yLlLuI8RQCnpyHiek7KDcY9DTLPKkJfOLDw3jotxZ
63LaLcMGo2IMtc+97TwzltnYBc3COKYDl+BqY2RuFlgVzY64zo/7ymqAYwQVga11mAXLZhLytPi0
ldG43bATG9mNNCxcMPZHbjxYzTfBeQV/XGm7kC3dNHfBRXMYXEpFISw7cVuQ+iqE8kOPTpSW1Sus
tsiHf7qtiTfRnbNGZsTs5dz9IewSzfiM3vNRvxlweKpst51Mam3AyJ9m9fDmkfJ8rs8ytDlsw4Ca
qk2Sn890axfK44C2rA8SvdsINPUw7vA0fyH9z0HQJF1IEoRR9pCdFB4V1/InquJAt0FF5Iy8mIx+
2gQPiWgZ3eM+4ybexMHuhcRVikOJKpx5mN2Ap/nHuI1ZLPfFF+QV0dEV8ZrXUj5y4TLCF7hiIlnS
H1R/hUj1ptuU0RSYq5TnHp1GtFG1A9D5A70RDuWcjj1LSHFKzwk4ubRQxp5tpSDJhmRVJUCfybJA
oNPwRmJNwwufsT7ye6uZ1H5eZPbbRcTbh0dVJwCn+Eb7H87SM0H8O/0hPelktPZE3uvuv/Zk+KKT
BEVBg0/ssEA8988m33aLFmwrAA9r8w7Zy0AWtuPIny9L20U1PoaVUOhyCc1cKuo/l882CibtV+YJ
DcgdfgtW0jqJk2E2qDI3531hBb6dFRygJStxgtzAkCZ6yd3rPapNoEknp6t+tEtVMb91lt4swQju
R1HcrZHb3QScb11dk+fdyR1Az7KLj0EfVVuhXetpya3z1KgsgyAshImGhLqW5sGsNpZqa+o/dIM8
WFcuTh+vgpofnUYvuGEAu9SgzyOxVEHjZZf4rUiq6hOZaf2MA+OoohAUqYdg7d6RxFHhxhzJrV+d
2I8ymLljUddF7r7Q2rmLiwRpcCfPtO6gOyDRHKm7RYyurM0yLUzwvgOon+Uwrk4g24gUC1W0GEcY
jzAzLD4Uv64JLBqC32jFMLHGF/oDOVwwo23dIoyQFAvPj8Jlis6uWF8gkVzQrg4uFMRt2cCjWzXi
8jqSVXNLpoCE4TVMr5I6Nmu/W/AKlWgj2dcnoLiNMBbvscdJkYQxJZH26OTc1On6acRAUk6dZdMr
KcIXcxhq2Rkx/OIHi10GHIggAq7smLmrC5Qxyxaao/NrGmVPH0+CUG0VE9xv2heFOoM3S4wQCuFK
vhajqMqKT24vUIL57QQadj1ZjON1XyDWnlM/lQcndX6puILeP5IJGBVzxjbOvtV0yvo0sr+SlzYy
Z3cWdJBBREHId6CNmIW+HSO1jfT9M8Z/F7WIdIZKOYVgPeAjUjS7nGm+RWrQ8urKNNvb3sEXgfT8
io9uIfhofXv18icAQdpH99lBg5/q7f/9VyRdEaisi1KQq2UqZag/dDbo6pDFHrnhUxAcXfCzxK1I
yYfuw3SVEm8aKFxzq9PFz8VzV6HsjWo+jikh8PC/xXske7hRAmv/r2ZdoZ6OCfYzYwv+3EEJn16V
zbdLVaA/yX/V31IgzHx4QJi6y0Q92/3k03Qwjud8U6NUBcp78zg/rgZ5daG7zgvNVIHLZi9Rdp0O
bt730WyZ5qUqC4HVQEgTPYM/0Hl0e7BJAqxShOgSUhJn+XrH4f8lp6l/uXudrHlETGMTFfs12rHk
5uKU7tstwDZAx9+wLm6OKyOMbptt2LOIQSxwZyGFpII7kTrvOZQZ/kTsYNyVvevVjp5n/61uxzyx
jnNSq+nfY85Xvz3w+EK6oixAguvlQkilM4kMjdEDDo9Aq5l8EhLVEhM4hUQLdAPXBkE8hcTXOnNM
EsvmtnSkirfJ/EpifbtZaXQMmN3bpBRcT/H0j+GKZeGm5aYTbRwwmJBV2vc6/69w+uzLbyWgDmuq
hI71KRwY8fULmR8/Q3SDCNdGwfuIsZZ+lzsz38hoMNhd2OqVV0Mb8dXpcIHgh+A/2XRYuSt2qUKt
rGpRJ+V/cjMHgXPBELDdv3XA2QCdv1BecIQdd6aYfVif/ku0ZzqpWGfovSTgyUshcOqrmU3qAYUl
/GNdApuOQBfmfwI2x4a8ISsFnZ7+KsqEwXUAQaWREMJA2w/jdpoQoOAbFoKDytzYXkgxT8t9OZTP
u6IfcUJBfh5TmtEuhSjlLAFe0+Hzq/lI6Vg3B0BbNA+CJP05OaotmX8J5AvU2XUxgBRvR47IPD02
VpQE4bt34VJ1LiMkLt8cRP99VfTVCvXeoLkdQYUaUVW58BroQUPdLk5CuezViikttDOLeNdVcuxY
eVAZBYErGQ4be9uOJ3q1s2e4e7P++2X6G8wgMX/Cy1Xffo36FcSu3pYoHA47mSBd1OIhWj1PHxyI
I6VuTLcqLoQ1dyC1BjTYRFEayNc7Zp4cDSsKP/K04VONhcjZ4xMuCx26Pm7JEx/nvxJ2oElLMbJh
O6pvvxMTGZkrc03okR6jChdQ7Sg/hgFVn2B9vXyc18/GxF2+YFJFsEYzZnBP5wVBZbMuhdg9RA9Q
uYh1zXlvUJkAB6Srq3S5yggInY89Qeg2OTpfFRYkbfzdrvJ6OtrZJs1GAXkpTg63B4u44R6iWzV8
ts9WWfChw67lHGoh3X88PFAsIzeiXCBZONbyPjagn4MBw5jD6K/UU0+cpoBA3ZSH9CC3TKbf1kNM
JrDT/ZAFczTs0SLz45MKJhY2RVoD5sH1cciLwONLVQ4+gK+jbIXSZA5/sKwlLd9AB+xWBdodXmUA
kq4OLzL5TCmIqFLVY9+BG4Tux5zMQZw8EZ0VHuFowVK2iHglVZgXq4NU4K4+bzTWklJqAm/12+kO
53xSEKoHaNeLZL6tHuXrqPYfogD5XPo9D5nd/xSe2/9f2Y3AA45ppFj1Qx13xaIaQl0QZGhfpFEI
n7mfIl+krRUQJGLcOqFLWBj2hTkxwIPHSfX2JZzFXYpJiA67i004OZ2bZ23dPiB/RF+abuOaepMM
XO8Cu0YMmezREgXdCStYeE7ecRwASSaWWFcBfWLZ3Y1EkWl3yKx4PSt3IkzJFvANn0enuF/G+pEn
j2WRDkImRXxyiinKY+HHLDkzuQOjPoaYPvf90o3ycj/d0CcnO3t6x4GylnaRitfoQP8D5tpP/ihi
BorGDEBzlx05TXtBmPbJwjeRwCuoZozX/Q08R2N7wmNy6W+zKnBnR6s0evoXitWJd5/oDkHqBUD0
QAi9xC4klXq/akunJSsJm9KR5RVEHC4JERMXi0GNJVCBCboFLdae4TeswHCcsONfz7JsndWi+cIz
k/SwtHePrXc/G0y61Vi7beWkX8nmaukr/Wy+TMCO75r9wznpPrdAyMnXbyjHRJPiX9SCPklzgY6Y
/u6TE4cCJvwSNArjJ+nINUIXMyyxed4P8ao4PrcxSPc1P3IRu9oWTn0u3hHcnfGM6XQfJxT6UGgI
kG6fZjoHGzqqDwoDefhE3j5pEkjJy4/A9vgBRVw9gUm0jF5MmwELwwLpRjRiqsIa8CF+bGv+/7iv
vIOr9iWDR+4+MeSnhLId1hkc+GEjIWXT1G0UVkDIPEf20JRa7QgFyp7G3RgORQgvG/aqNOtdUNRn
C6ScgmLKyNd2Ptw8UlsS1VByMigSzm+5gpObxfjgQp1j2loWv3QmCA9l3vMg7LCBc+jXFFe6YunE
KeFDJl8j8HqWrMDJWd1Iys9Fr48PU+5dQtKKNfFAQT2RaZt85DWMqXID0OiptakCCJuBlBOIPvGE
0oOfX/QTagGryZxKXFRMHCp6TEPdVkYQbLk2uXkCTho4rPH7HIFaqBQl99NZRm4plJSV+hBQyIiN
eH50nux0boKh9INFoRle7XcOlUI3lp0qHNoVCezT2U3PfJRdvbTHEabzV/ok7XzLs3lCfyMWfw2L
z3kmCDMgzMcKvlnESpTLV/nS2L219kOYQqwXdNMuM1a6JOTFI6cRaEIhR2TunjbEebbwkscckEGz
W+p+AUNKweF9f4lx1dyvM1MI/4Z4UC8kxEvDazVwGtJ0aH2DbIybzxANQacVBTbDefJVI6+8HzQ0
gwGrRIMvn5WvLlff/i2pwtE3Q+Dhm64CAJYt+KT+gMVEOymbVDpZoU+YakpHaaSFJ++iOjLXurWk
7Iva2faSNcui9m8Wyi37nKDPxtMV+hTXQRP8JLDu8DYOqbSAoyTCEkwFjHlV/u5yRNr9k3LoGJt5
aKtFY3obp6Krzw0Ue+8jMdCOZRzJByRZCo1Fy1ADkK0zcUB8vPf6iQkx3E/KAYhUaIsTG6u7exA3
NqzmJDycIJSKojmVfdoIWh2EUcKGnd8GQpE25n443dKC71y3C7TqVYnsr0R5RyZ02UIj+SSbIrC5
uuTPQEognlIQswxhLcVNzmE5yOnAmjGb+spMIeld0/pSrrX3zs9sisl08UJ4slRfov0CE0giKwn9
PSjeDX7QP7RQkNlSE7naPCkH0ZvRbV/dISr5oozxkkfC7Ex6O8yRqjpxtfEL776jCnWUGDCQ7m0p
qJxlyKWYcsJCKK9nP93P4dUGvIFmSCdJ7NTD+F5qkH/RcSkjFKmO3k9TqTGtWmewGcHOy3oqElDQ
QyM3MBQ1t4UpJqntfUnxMMCSqFpxAaAymWbFyufp2mvgF6+dcLi1n7Te3Bt2Y7rBfYrXl9jfxHwl
BFrfNO9Vaalvsh3Aegbu3iZbhIcYJb3Bh3YOlt5t1EFHVyIrNOtYQX+YN/9aWGxONEOmCJuzvthY
AqKBCYRKnKHPLX71OomuPyvYaE5ZXKN4hXlsn0hjASuBXttNiDtK9JjXzK0NxJESSTHF5EBK6GyP
VmwXSdp79HFFmc2G8csutKKNKeZBPO7N2g49h0zohc/B/sfklb9NICgudnXnXjvwuaJi7ZTRP0kB
PIzfhQtveK1rCwHMOduZ4jxEYdZf9QecOLRG2DiX2dAdvOZRYHEMVwF+/zhDu54CHdCuNVJo5kYY
nHMmCotvRd+BZcJ3c+GqIy9wK0WohDeT4Xz39khzul/ImlqP0Hh1l9TA/O8m/N+sHxt2txcNpkX5
8ezoYIc7gpwmheo6xzX5pu1EB9dT1MoCx9dWK35Al02NyETsbEbzGHEnx++nr1zRT6EZlGgEEli7
CnY69chxqyxouG/4ahIQ4mBJHsKK1c+gd4b+1qRHqZ2PVotYIRovhw5hQLGddG2Ca5eW285qsy/X
SbqrPyPhnKkpjBbesu3hBEI1+ItU2kGdC28IOWRwLdTzBpkXfuLNwNxKsusWOdgCeTzqBMJMpkOQ
R005qA9rj3TxxO+felAmJWT6y06U4wqu4CiFvw0yp/5UvWpoTpD27gZr58T0Q3QK40vBzUCKZaHF
hytWDL8GCfLMY5L24ueduuHukw5+eSgdpb73Zw0vH72SAbCciEOeWiLKRtL83Zm08Y9FKD7jr2E0
yG26kDZI4QAZ6HaQ31Ow5gXqphvf3tN2+fDn/yakSTug9Bw9FhoT62/lZ98qq/3z2L+VOZs3K6YM
ZQ5nF6oqPb4h48iJaW6UpZoBaUxgCxUGN+AEsSvYIP3+zIpVcCdcA2iYp9aFBDYwnXtxKrw9Jm2o
RWiR/CQCwsvKymdWHm2iVNPjcSBS2t4hIKZ9TsJpodXNMiu+TSy/AR8IYwV+vzRVK/rDSu+iHG/l
m15UZ9ifz9zeq3haKSKxRiFwWbv8rJu8isXTdwKXKmp1VfCEfHDaKqolW7GQDjwVD6mjfRKz0Q7j
s4GaQZD0JUTh9u6QaqhMnRQU6vSEluuFBRpspyKwvjl136cVar/r/QdO+26l2H3n+2dcG2fyi5iM
ecP1oVNIgiSu9D392cLpxhiIt6RuBOoNlNuS9oEbspbow1pPa+HEGqw6WWFTtTOLHsHBxUmjVvmG
5BzXQI4J4RmX23iJUAz9vCcs++vvGnPBSo2dPsBZCUPghzQo2hsv6jwki3ttYmGiLalw0n7JVqiH
K9Av2h41/jTsE+7dufFKon2PqYT/cwPiBlOlWnlkp9sVhfPAHswflcLI48n9cVCnNryk1dmG/e6m
B33Y7L6vPUbjQTmyQnrL7ZxHrt4I3BB92e4LQAKcR5ms+/gGwWBhfojh3mLCzyewOE4M/U737j86
LuGiH8T8Fs9D/voRQs4HaSHAocz3/W1lPMkZ1bt7MRvGlCFNxmNMlB8sciAJv4wdqLyP9+XNUiiO
OogYrbcxDStALHCnf7lsQ0LtUzrHWA7I+V/Wp5JKgyQGmsw7wcMOwI30uGvbQ2Sn6XB75BMQu8ja
/JxnLEVyYyKyKaW0SDmO00NJjxTdzMtuS+LGz8xl0qlUxkDLyQtt9TkbXNb1LqBdcRxBl0O4WEe8
Py73UGEL6FDLgTTZIp99UiMTjIMIfhDk252cKW9xSW2RUz1+MPbVxCsyACfvMvCgNU3UaYuAfUW/
6LgdfHzzzO9u07jtO0L0ZbQeL/LfStBgRTncdabkT0bgtKe8IIsPkZKTs3TyTfuUW74wTTZchklI
EfiYZLkTGfiRt3LH8upLStuaKW73vo2JUGsCtzwV23Qz6mPyKOvgwkS3e/cOoPr9oPcPbeeCz5Yi
I8pYhbF7X7W2NVf0xf81kEqLibZ4IoCKGWtKysSuoYWuD1AOS39DzUj8PsU0VIrYpRtB8iePj2G8
wEFzEr6DwDmHT9ervIzTFRZDKYUYjFiNywCvF9+YG+6P31Abrduj6hcXYpGpaPCy+02+xz0CSoru
a3W6xr67u+apHci9cp6sNlCRngxfdFC0hDpmaUVUqi52E8sVv0RsDCVVeS3zqkgxADiuMQltWTjj
Jbg8BxnbU11GT1MSwD2GBkrBWanQxVyHjynq6ntmxL2E/rECZIK6blBEBMLtJNqKfRRZ9Z7e4FAr
kq8AUv5opL4gRXFVY6kVPsZWCVIyZBg/rs/gJtRNdrz7DtbbDbgn1cNefIh0Qie4kkIb0W2INlp5
NEAgLHKlM+lUITTPMhTFh4HSZLvpVzonSYWLN5xFcGd9GlKrvlezyNreQNxREDfmt9yFKZPaPjFG
ls+KVC7N1reArQKAt+8sgWFtkOeNTf+2MbwFMAGPvQ2n8PiyLqYoOpWBwO3GdnzCfqrktJQaieWR
IHw/I/yFOr94lne3/P2IjekMteN0/uH6WG+J0pEkXDkbuPyKhgGDccbqg9WDHGu/vb/JhrvIgnpM
4yppSxbQTwOZ9yGy52ctTPAUqAR8YHJtDIJsaB+SLhvGuw8HBPBIGm85tFTkAEG3kQ0F4PVMO7Pc
1pE+1wjTE8L5BJlSMErN5RN23Tms7LcqN0udYApQl2L84vanD9qFkD4WLJSs/AHawFzcZjWUe9q+
kRSryLIVtMbOfRG6B4fCd6enkoF9326y+If/f957EwtJUa6EPVYveCqBxpa8Ys0Gj9r2zy6rDRzf
TtHtiF4fBTdyeIj+KiK7MqC+F/jkb0VYktK37SjSVKP/iP4FlnjI4dqxG9JQZTClp0m9NX+4vU1E
fs7sCUIT73IRMJlCth4Nl7XQtSETS9ZbYT+CaTaD/dZtVzarKVGIvDH87H8iXDCY/T6byBc9FNfd
DBObqGeJpU76ugJFjlaIUCU52nfVKK9BiUvH0VWrw00iA7tMP8dPVo+wWkjzP3t8QsWnMRsO49iA
whICFO8N39Y2aFrtVSJrpkJrG8z5sxe2iCKjX5lvwo/Ozcjp7uF0Mzh4m0NXc4E0rjT4Rh/SXNFk
DnTFMinC77P33ISwUvr1E6b959KgLLVdYDC0S5cEusJyU0OA9EIXk5Ry50Tag1ca+oAceZSXo7C2
vjYlbdg/sxuz/UBM8eUppGXmXTOklo3qyagFRfP009PBpS9VF0Ro4zkTSwHoIsiGWpzS6LUb9RNl
cTZLEz2mpDsRhunFoR8BIDbKHo4AFayt4B3Tu50oxLJv1gRnByvINFndGiyz+C0tFs0OGegb5AUI
LzqI29GHjRDW6sF4lfkg3/vc0feW00GGCr4iI9L9P5pCS8Z4CYDFlR6tV7BdIIVKz4g0aWBB2S8R
g1abCVXnV3kVAozkw08Ao7SKDW9oaQi6HWbRSdFtWd1tzJxgfRt5F1arnaydTYMFU/yGAae4aoPc
eQcoTnwndTaJX0IRawHNOqy9ojo/M9YBUhyiuc1vRvufRtjxGaWD5kQv987lYNJmt9bxBxqgilg9
8h9COKKeb6qZr+2f0xO4qQKL4lN1woZIX3cYqSVG+XdS1hXlPZejuH1FRgxclYrQI8budVe9fWWM
ceW5mgG21xzeEizbY1PRy/n6kp7qcdGN2N1HXAoXt9Y7mxrHOwj9IxvrkU51QVmN+AQwjD23ZwQC
9loEI/lMAy66ah9xAAjmEXfDurfwCKN8oreppVfmyEv+FZNNP835kLBB58xdZR419CmfkGHdc0ri
fgpPkRA98Zdgpvp3JkKdCeCpHCHPuWzxraYBzQjs27NCaOpPPAxZHzLbHGCQ++WiMrTdG3uJHt+I
pO8D71iCzGMNpSWZ3L6dnDvd7O/4cjZO4dM/c8KyPXFyfI9eeXUCkA1hIA9G0o0a/Vv0p2wu2QCi
UR0i7T9R/M3pdRP8GbAbXjcvhmgaZs+6j8alsq1udF81bLqob5ASACFZ4BfdrBhHZI9inBXsrGzC
Lrfdlm9HMl1Pp7ouyMKBGW3pJzO76IDGEO7jD8XJNcCzJI7M6sfHNBVEEtYmrb8xDlp5zomZayYr
kslx1LvBDI+ntP2n7SoVbTFDDIRZ3ZSnuXnKcf0sWbUUFJdw8Q0kIBN0BzgJpvVsB5Si/RZpOpKH
S9JVklyz8RWuwkRESg8oVjVOPILmdGa/JXs1Yu03i2/F26sjccljWmaclyCIII6MY/lcxVA8zifY
ouLHpCjQBFOdvdIiC6AzWYZKwBzIbgtGkUgV6sWJKTxsGHPw+Oy8PfegwfVT3nUS2Crusc0fXuzt
HHMB8oZFB70xWPoRallVKgZdj4707I3+OrkhPfnQEOVQqBT8J2WpiRbGX3hrOmCkURTosO40QikM
3E4YnojOQ5/1Lf+kIWVeaF9zn3ErEyMw/FPCGc7Hh9RUvDH+PCP5RLjXfjY+6eLDgr6pZ0er6yud
TChS7fpTIXPIHueJekTuA5zdgkVJ5KptWaJ92Re12O1nyie11h5SLOHXZ71BLXY3DQllOeUGoCyR
qPzcll56kyd0qiv+Iw29QC0QnEWQsd8IYQjfJdxxG/FYSri3NWVbx/tDPBSIe4sNXSNuTtayjZKh
J7wU1WX5xANmJkVTSiELru0Io88CS/ud28XsvFbDvgi2qVjxfH2futrl+D1obIALTx4Gob9lIA+t
3JF882V9OccdMOqWcAifv9E9SQVaIteQIdPv7JGY9WyYUHg9HWy5IEmaW0SmG/TgFmFpULKbcBUR
ROBAvz5EqCL5vjGvM0FTJro7A1XyZD/mFzsgpvSG8ArMmzX4fPjEb4uJdk46mMbxLB/9z7Jvakeq
5YbTVeI9jaK1tWlTjYB6pnD+YG2rFLX3WgZxAuhUFqsBwIBgLnxFDmWOuZFPnlsu+MNKWP8VMZ5X
kD6iim1QWwDiceEW24pvbObmyRUDlV4Zxy7Cfpzn3wixB6w8GotHSNkX7PDJwRmFgBZ1YFdzbRkW
o7Dbziw29F0HxLOug09c9Z3AkPDNdi0Jl4wE1Xps9SHV+8XYZyueccocrCwI0pJN3oll3zPbwSca
I8CjXrbeN+BvN1aWhv3ydcaxgXieT+7vX7XmwQHkitxVr8x7p3yrNe/hwvI8zVGG/7Yg1mJdZRff
GSCMEFbnwu76M8PV+KZF5Y5Winob/XmnWS9XS1rNOZCjchyZKy8mPriUYug+F2MhvUZskfw3JpxK
0nhpoRQiJ8LbGkApg2BB70nS4N7YXSsLIVORO9u5nUpS6sWYWUtz5Hun5gN4BnyNCWX/SsVLdNjT
BQ/ChCr/gJY5ppq4Lj3mIBJAtkCh55m6b62/42q+pz1T6ZBTLplDDK3HC4Ny73E3+HWH6KQYcMgj
dthmVukVQRGZ3Ymg8HXBeA/4pA7k2pyet1OBnS7+pdq8zmgZS29NMmvw9ZPQHB/Y2wDXbKcRh9/A
+2eHSgLR78HziG8pyw4kY50I0dTzx7w05PRK4a51aZQlr1cOcMCtLuvd7xHjHLqG8E+T3KXcF7PP
2PtHn19ElDwqaE9nMAYPe+CrKeMBdjAFgrli1prJroOP1BxWHJotqITb0IDRgVnL+9czfV76G9HN
DN5PBx+hDxrCxHI3G6mdjFMFrLPOiJNVaBmhtDzd8oX9ANiBKIIFo6Zh+jvhilQGkmIuWGJrEbym
2cDoe1OwY5HE+REEHAWrR1iBNeJOSCB2oII98uWETJEzxNBcw87ksVhvq5Omyw22e7AWtGhgB/8z
aTgldNnR9TuUqorPETCge61HDmyMkUIXcOLhfkkLwnwrCflxRSxo5kW7qkSUofB1u+gQO7QeL9gq
jWILccohlwCmATO8MdPK+vWwR/eVXZfYNj53oRs8pDsp4li0+EqXRkumOxfNxV0qz2klqk4RDBac
lOEQYMbf/uLXM2VEs+L/uUUXzylo9FUkJ9dNn3EG1PulBnpEGfLwyTc7J+oUMPaqjYa+YDxWoOO6
quufagy5bxtBuR04CfokMVktoh8cJKPLvZFVFyk/Lo6ubhYe08hH2IkTkRkJNKFeVWbacl+fmWTW
mbiRAV9SpvOsXRA8vruqKOmhxbgPTi4Bh9Y2RE3IB0sf8wnyu5LGgAvlYATs9clHPKtp02BxBu5r
PEbFw23torK8HCwyyl04XBLzIRsh5dIPZJjrbWcWl6af8leul9xCYJuo+YC1PNxojyXmedFUIxv7
/iTQ1aCyuwI8uXkD4Ut+B3f07DqycXmacLZ6hcw/mjjXX3Y7VqcUHFsg1vlPACfbwdAkwCl04y+y
YMiwesnNYCs5gtP93kzYT7weec2wPILP2MfL/GQx6ckPjtpcoGxA2evsRsIfkYJ7WDwoDqZCyluZ
UiF4IYoEu2mHFxhzs4PtnQai+ilglo7vNy0Ka7S07UGnosQ79AltC3GAdwxi0Jx+psX9o7ibo53x
8LpKqxz/Yyds+d3OxqAhTexeLJA7XLxnPMftR8iNM8iqbGS4CtyuPOdyy6DHoPZeROrrdiRbH1aG
4T1ZTq9Il4e6sBzYIuDSkLB5wXK3v57GKAjcjL3nL4GnSSME0hQo4dGbf9c5NoLJxucBB7dji25R
mfqYqAmhRZy+9dBi36qEFR0LDFMDKx1kf47a0hiBhrpppr8Xgh+nC91NAVQmy2+65Dxyb/mIkN9i
8GkSBStd1SNvlYmK6HHE9KyIIiHtbQujT0LYKhegi/cbfNVuNSq38+usycfCCQSThggPIU2zkoS9
BG9zD0zwpFEi5apPP/U/PL+G0FXiU0aw2hBDudjQGnGNDYiVqqkONfJnNRfT0Tyd1JTd0Ko2uBY8
QIBO06gXKOR8sPrAI9HLgY+vnwbPslwSIcDe7JIehGaXqwlTNHNNskF9VxEWwu4OIH6YDYiYTVVr
QHtvsHqlm0lcGIUgDWtc7U55Mipz+oAyubXuVns4JdW8bnO17NK9TuPNHU/WdB10bJOoCDpL5pSU
XPG/dP/yUgMn/5kLlfieaQMKevKssO53d+8nAUbjMMP2MVhtAQ8ClcthLLY1MjjlFsLuT5p//yQo
6qt9rTsfU6iG3/HRg1TXBgg3lhaXAemHx4BmGNQqcS1anfBcgSGwXPPbY7Ko9glqShcvgcNS5KOT
a+0tV1dtkRRcFB8wGugYfhZhf7fdR+ecdks+QUi0EgPREyNu8wcS3Qh8qN4rgh2tpIieBd4N+Ref
pEkZqX0B76DpCrcKH+UEfvWiHYFUwpBFRdBg2/T4O7DdHtxGIFZflmhOaCTije8YA1Qzh/bHzffg
itTVmDJfahE9IAn3gWhjF8IW9/rEEIC6CN5XMzXCKjP6C12EkJIBqHwof+ZYi8T1k5FAD2cLmRe1
fEnVGXaGfG/JhUux9znph+2z3cjvLf5DbILKYIqji9z/315mbSBnThctyv4VIdSeDkk/ETU9ihzg
nBncWHKRwYldAAkSxHjZ9jihtP7bs1SOAvjWxykZPDojatqLiHSKEOFCTpBZNOXW+5SpgSFGJM2l
bHKa4QozxJ6FCXCEy+axFxWOPrPAf3Ho2UBKydJ2D/26c+4HEHagELvPvj99mE/Qwzi0fAmLDvo6
DTnQeZd0XLUQZnMb9qGjL1zSiYxZJM1yGeLJU2ryr/iBSDuVj4ltf+A7EYxf9aIheA8M3G4GXwZE
w2xhpekm054q7kFSzmhwyRgrxXZIg5jEvHSCEW1QZR3qPLFE1Om6r6zHTi1WOs5HKTTROF8kjzrR
TkAuv5P8NdazNny80fxQ8ChmFu7cLT8s0cBpaKd5VfC7zjMrWymlNu/HQPDalzraI93lroF3rvfD
LdXIvAZlPtSidjO4hqCBiiiuwyZY+t01bYqFUr2m4r2Etr0FzfOOas756q6f5EehYV1ZfP8PB4mc
7M24ZAz2Lxl/aQGAZG8I4W6lxW3VbRoZCc6hBrK17Vg0d1HZAoL3PJWQvHN1xNGJFNd28kwOweVa
gzK2/QSzmG5EpVyREggI1VKNnhKa7oOSR1lcMJGE4tgOzy3C83xfV4Y7TtrOWRUAzlVP2SFsRNl4
LSseUe06s+GYbrpEPbvyhlQK5+uUS65PrfLgkwlKN/70Nt/3Mrveg8oRjGALA2Cilbi6RDn8xRlk
tChpiRvxd/IiBayLn3CCi3zQ0yWA7hOoVW0xZuBx/+MfnYbPalCkGckWrMWlmYdmhAsWhMVJJa0Z
dBewTm5k9ArgMNBjg/VKvm2EamUAAxVMr+Yofw9Ooab3ccaRmqSE+v+Hiya0j5DFNawBtWeX/PY/
NHYGDL4VHv0UZYDMvkUnWNRFNS4TUbCYHpJvCfQUlyVv7ELHv+eMJJFXpRsyjRZ684Ys/fUJajBm
0rGc7ilFrOiaHUEAFBh2GOWur+IVbxidYX2Qejcg298lRiNCZl5fcxFN1wfxFrHj39rmLVOGhaIv
orR0m4gl+yfJGR1AkYzZeJ29lGKU9np9rTCRG5i6n/OuMsG6KDLB9A1BWEwqdD24CAelwUUKYDRZ
9pUhHCDbULHVn4NWxXE4UOhYilWe4qDrN5ShzwJZvi2vJUHNI/EnczZiEzZWbj4Hnux2JgfvB8B/
PXcSXu0kavZwL6E/pAv8wed+abaj0jFWz/aiNM+9w/D8YyQ0q27b//zG5C9L1bQpqefjQJ3hFlMe
9+2Ep2EQxBDHxknWNCz3CkmeSAR2e06hboamBwERr0IKt9cYMROH4AthaXIPFTML+E7Z2IFWIfoe
fcVeklnhS9yZPNxHMRRFc9uSRkhmgp6FkWidIUan4RVx6OPZ8txMVVstpXmdf6iUHtSZluOY4xDe
inHkn9QIBM0Hgf7KPP1PkwBwICm6svA4ZPc9ARVFbW78hS9VRegGfkF2BO1UKJ35Miw5GGyK3kLm
fPY1ucnm5ehxBxzSNU2U3ovnxQjn7w5r8KVmOnn7mzv5V6Ij39oG1JZ0VoMu1T6IMEzw6pEbBAYn
2jO3mYYIngFxELfIeEQHYL95yLFYuH7LYd3us8CSBlPljUP+K5yIQSlJAPP6Bw4A+ja95YwiVnuY
YrbLqH+Rx1pZkOTHJoWYJYl8ZUfL/6hhx/EQrfbS3aslOskpRJ3fvhVREckajizu8OfWefLaNwAD
nX2S3pV7waz3OxWvOH6QaKzVPTlFzYCFbXFvhzivXjmGLiJTznyflcyU+hYYvWoKVoYq5D6cmSdY
caRSzq5lYKhVRyaT32cZ/cpg0pT+oQsZ1OPrL+us6E3iM8B6uPAEbCkDltFdVuvgMxt4yxBKBnu5
X6OQAHr9C0KhfuO5KsqhxRXCy3zwAfL+S/8YWMsnjTV//3JoLufcehiEnxn0ORr/GhqfSUkuGIjW
jVUD9VaJwiOIemabgWaII4F3USOreJQqgY3iwjrRrTc9IOh05mRieZth+y0Ahy2pQr+NLQKHPcTX
V1roc0ks4ap8ue5Oz03GKU7J+/JadiJ6VqGzRhBITRZawn74EnB5yfLFQzX8Agf8uxk1PIhY3YG9
zVsEgOgIcxao0Tkqu1nd90IE3+05TJZJXbhPiyW2yTOe4UW9gRNrf4L7UCMMcVnc/pQnFm/4oMq0
msONXJ6kiQQPEIrmeHR/nMHksjWEISkpEXGcYvA+q9FuQfgMy/5n7uUqMZv/Ve4yr6DhcJCBFb+E
mwTV41TvdFMnMedMzD4OLBKzuLaYOjEYm+gdAIDTvpO0MHkavaQyJHi6pgNbS1uq/tE+oRFZqCp3
X3R5fSmbPp1Exb2uXmmVF7Xd2UgoIYQudp/43bkK0chUwhXhPBy5HcHyvsYmmVPzzMS9IqD1lUxr
rB8DAjyzr3e5HX2FuT1F+9n3uuVa5BlsTGIVgAkAmDNzldAb1Bfn4QTqYXK3xuXWQyRmC8Fhgsye
ak8oYJyxCDVggqtMBGz+KROk/VQvGe+kC0juuegwZnbwgIwJllWhWyi7jw4Iv6Zl4QtuVjkYzpnM
CLplmUyN8BBv6x8zFBrXQkH8o3bI8LArLSd+hb8JP35/XcpKg+aur68ZIUJePDLOwrbkW7DZtH1H
d0pomxCis043dDKyRTxv0g2TcqEbrkUR4fDvwdq23oc5s4uW/FfCUmFy29OKwK84RmfwnEcQji6Z
gwrp8TTxSoXrIYKPvZmH3ehEfPe06LF5y6457L/B2FvYRh36bBKuq9UgqsoJE2GSXlQJKdS3pKbt
topGnic7D6PYLqvKipn447qprT53ZF9s+wwSCxo9I5XKU28Emciewlxu5q/HhxTu+CyLidL7D5Dz
AvUBioGmMIwXmCsqIKHFPoL3RvoSEpX0prd9V9Q1gMDciMEyZkTpW1AZuNQ5wfQ+qM7y0enddL5c
KyT1oVT20ACynVixxZ5TyzZCnCOzWF7eo4VRmvIJRBNHBUre8BgnhjKy9yClBWFeMvUqUy/Vxavq
bhjqC1CvoD05qYiZ306T3jaLE463DtxFzudYv9Z7PujUO6yXA0cJOWIiRcSNqfoUq1BB7wHYT0fV
doweK5EuIeQwI2rWT4lC5EE7CatBKv4FpEJkySnP4jyUlHD17WGZxzeYhob7c/+pfbcNU9DjcDm1
/qcfmaybq2RIhyN/fJUpE/ziIfvK5YPBTlTgWT7OIMY2zWRSE6sJJBFNYuPT0Bb1ZU8lihRPYof5
1byava2xzpTT/irBT7zswe9Uhb6Setl5hTQnWJFEquyq4o1HHyHV4MAw8pOHLmKLLZaWqTTjbh3J
XUOwQoTkfuIOOQB9BBNfFHb+233g7qHN7y3NJetSCWBK+ZdZwhmLpuQ4wmOsiR8pbpc1SZ/NtSJe
hBV0lo5CekRHme3BafG+6BGRxBPhI0QNdWtVzwYcFd1ckMm56ogs67LR8/OpiCbOEDmU7H3obR4d
+2X5qFtt0mRb2rzkaYfi6YLESemn1aaXCYJnws0aGNs6oC+RFwf0BznbSCS0+bYK4sbrr0iN4V1d
13LyGhF3hEVWEHZDwymwDThcW9254p7qIskkccGDZcQNlI4zara5MdHiQy83Ld82nxsYplQkgqAP
asX7qg2z85dCgGz9rbCy+HksxEngrn3ffa+/elP8bOrWfmH+WhA4BgjIQDDrZoUMNvzcCGilvbzA
Hpzbl5+gqzTIj83u/ONFiZNZNMMwTO/1ByKUpnhQmzXqCBcDdZZ01iedD6fYhmCv4TUiq8l0xNvx
OMrjgoFWB6b6IVZj0s+brLr5278IxD72gFPbAmrDjGopMhbDkEBnaa3CMaaWV63ZIpyo4m+vlAfN
qgjkPcV98ea6kePLthe30gc9Z8oiGsfFT3xMwppj0jefC/HAXglQAr/+VAEYZWqhpv4/WGR2GQsD
qvc7QnlyDzW+DhJgIQtYb+uinK2wER+Txv4gTkoQev9FtZiUxwsPa9eXFpdDNSAmp0sTmqsCakaQ
X0gcuo1Ugvj4x5eMJvMmV7oz2AQP45TZPwP3K7Cv14y1FQWhCf4TyY64r5GxmvlZmCfnhQxN0RXk
bfd+yBcEXqv5KBU+1OACKUK2QMf2KmLvqFIInERwtCRpbouAcsMB8mqDiAYDr0uLFMmpGCXuM4zj
yO0jspj9YUg32EiMvPK1hc7HgroxN6+5x5DvtBQMh0/+3i58fwAaz0mFj1se3M0FQkF7uL8mKV9k
0ZF2tqzNxQTgZMMGvryEYZz4mVZp2CqNDEUH173dhstnkr3vpWeNukHLVwPh3iY5u4fKvxjrs9/d
jBV8Wl6ptZjgTLz0h1vxc6UTI4SgHu4CZo8cotNAtDG9hLUJ5ZeauHQdmMZoWYGN1izbi02uTAvV
9ZLExdKrzQtL7upwoCbUwYKn4qR8NP46SJhhhRivND99ouzta2uWyIAWAXZLseJrtjfIithm90AU
PDkzB/fuRg3SXWGvxnSwcQgmCjEkF2Yvhqtw82K8CkYB2kaiB2eEo7nV8d2YIcfjjOhqSZDu1Qo3
CoDcuhm4NuFlj6F2ArB49AnVbjbmyDxW3l/o+NQX9lFPzWB5oUkdIY9/lZ8qFGgXN388/whVEtR8
iCOpj8vKd00z8e3EES0dKEFAOjScPPLxVDFsa3PApvI6H10FMBa6GoLv/obDvfWXzEDY94YYQWNA
XcXJaU0thd4ekgavxsaGV9iF0TpTEIXVbD8RH3CE+ZcfMsMDMawOTifV13GmEFNa3tpCC+oewuAj
lqZOwt0eDb9USiS5zrmDQWhHIZj2c36/fatYaML0P/3kzcOj2k+TZVDq+/CoknZOuQkISw+XUHYp
Bu1B88lrZPnmU/jRTEB0GD2xiC/G32FxRUoTygHqZ895TIjVfapgK1WS29FnY53jrg6Tk1CoQF2c
uSMGoUSQo6aYcRtGL5AivCnTu5kV3nI0/jpLlHz0dLYerwgAycRzq3uNS5RIjLe39sO4fM5dY9bC
SEK8du8S7qMEF0CstZl6PJr+TpdeaIiAF2u0WTwvRMnifPkGnmV0mPKLqR1f0cBg8Q4EYPXBSp4J
dHEbiFNLLFEKreMjvg8IbIqzUiswxgonXMu6GMeVC/d4SHEarkc55dKzSdiksr38kCjV2qXIq9yc
GUIDptRSXp9dsreDbpDkRcxck56NcGv30O7CENdKiPKgpVPA6+fbkKEOOpf/f+Izr9ghuCQTVyLx
zhMHCOnAWEvm5v0i9poZ1rmQ3+U6d1rA+69IQ71QY0rx+j0PjwK1Oa1ryGJqZ7z/6BfJzIbIv4rj
v4fas1mqAob09XLbmHJh6sYN0nfqqLMKkLhVxVRt/JdHDprdF6Uy+N3YUy+LDNXaD/uhV4Zx7n92
k82ZkSC3Bi7TJbObfncJfVZLokb+waHlrp02fMAU3k6bYl8yp6VuGKCAwESUFZTFQQYE3nQJXMeR
FyL/WOqGRRW0/YqhU0kTFDbf+hlJJQQOKVXO7lmVU/E4OS76gxIuil60ifwJbVTBsaplOImWZ0Vm
YXUy5JXBNBLIhRia/NBUxsKN1FiHVV28B19zxFrHSeYz07AMt1gddug6ondGA2n7vjpt17dkxinO
rNU/UhblPcyn0yMwg1ppRJxHAvnPc/2azX9L9FhjxKrKea9VUUbsGXpAFb7ZBTMCXSRYia42eL4P
FnAreVm469Bn/lpzBY11N8PW+C3umKAnMFAUStecagAs1O2XcYgUPPkl79Ox8dtg2gIj9LGEOhI2
IioLbVI7ghPbUQQ1HoauX3d1l9Vfi0K8ZTcidlSbsqX1GRpUf0Ax94EQWFMNbJZ5gxt/pDVOop8p
OkHoqxvfwFemoTJ1oMs+9sskPRiDiggKwAer8C/WF3s2pJFpzt3P1MNS6dtDjz2QIVrnE6UR0erI
HMt6rSRv7HzEbAnGgp50wwZGNHVLdnX7AE4hdqnxmtEimQmaL34Dx3GhItRFap+0uN5SkLCorydp
DvLKlAlUyXn9ZFT0q4XuxlARL8pVXrzgebkevY0qiNx3+5kbiH3QFpTm+MEWT284OflaUXAhL90N
3hd8FSiG+qfUT4xR0qOgsKxts4mplVxgn2PMXZR0v9kq+egMslS39J/OHVfxdMklkVTh4lru83gZ
CNVJkjKBmsPnVA0PVyeB9c/jRammo7j+olerZuh+FS2m8vT7YhOTg3eTQH6tkFJ37S9KWn8uroOK
CcVpHWL281JUnZK5iRE+KVdq5ckTCLaJw0s3Dh/5ShHyDdC4v65cRrabt8sg33ETCWZKV0oU6t36
D+2/PgeBpoQLN/x/+BCa4iuvC+uC7mj9RRuEfb/kENbpY6pgbh8ClKN4JmL15Rg9ClIT6tqhfvUx
+INn1e1n+bqwyf2BMnXqxrTwFMhR7PSLVoBqJFW2RGNqV4occ7BsONn2GCgjuNKJz/lmkrXZ/9sl
pBZtHNN1/BW4IBBs8QdBsYng9XX8QT3fc0lqb7GMp3zqcLh2c7DLO71issRWJvVQAsgpFtVMeSEA
ZVLrY9Gv0OXqQBeN00Jq8DVmOBREWWUIgBmszjvzRsMe940d0FksUz/r/URRbbop0VGESu0qjoxs
7mEW+jbQsGwvWs8xC2aKjEoTAiDGKxAx7Rej3Ifr2r4a+/3/F7HUQ1zLfCI75RYvvdlf6K7dsyLE
ClH8mMJD5kWbw/ev9kdeROQJMDlkhyM2wEvwtBjvgEn1QH72JjWHv3BN+TDL54pEm2YnDfMLehfA
bNTdNbVm3iCIInlwF2Rr34v/f82sjTpLMoIVW/vQeEuSLTuRWO7NutxXCnXr6R6iJHNndCoMaQJS
JNP60cDcW0ripT+/A2VKQI821cR42VfTwkk0TC8iBtA9sfCvAufAHT0X9b2KS6F2vlKx8Djdp/qE
P297BK9hWvqvnPgtAt2VyTZgtjkDBeiYOb2hT2XkbL+b3FbyAJGhIssH1bu3MuOQSssF7eTamRpB
UpkfPQ5mGAC5WlfQEUCKDHXlpVHEuskYgY2h2AuTKEOKrSvQCe8Ho40Yn1HoTdNb0WriHsiNXycD
J1iYUsbRk/JIBpOD8thnQFJW5QhyJ2y1/0w7ETCoG9ruavV3gTzPYtQ+zAEGWGpPeE9NPoOdEe/S
MCZT8ILVX+v4zLbjKvTN+4zBop4yz+Odw63f1GZ5Z3BS3juNyGruQb5JiSzGzLq9FkSvOqYLxzsS
nasKNruII7DK5gwb1V+CtVQYnmgprmu5g4xMVsQWo1X54R8rpHkKKfiKbW2DRLuFQ8sUAJzI/EIf
BEg/p6/+XM3Thu4kYSfK8The6DIWJnnyZmPG2W3/5ZhT29yBuXeZbIZAbHtdMG4TqlWYod1lmqXL
2+ME/EiveCicIi87PRctxwlzKonLxaju7Lx04ctpBtl57aZDnB429IfGwGwXcLOYi8DYXMnj0eO2
VCzVJqeXMilijfz2km130IC7SmDzXAEVJa6ZJUdvXGj/pahNn6vMh6JSLCSyuQJsW1slENhNQcOK
LiWGSA+ksYL109+iph4m+8zIAWGOXmZsNZrZuPDtY7/K5ceb4SW81muXLgcFAWof5uzm4VnwWmr5
Oocw8oS/hYfFARV6gkPUglP52R73rraPqd+qQx1Sdv72tuWVvXtVj+ziLk5MHvaQZdUlV5BwAFE6
osV+4T28ObBD2p3gwcrNKrOkiRBH8JD0cIu9VCJrdhcO6OooofMZVVWHSokVwIfqChWLi94Z92Un
bZwN6Hd4xawj6UXk5h8YjQ2Ku2y4lmImvHRiQXjWYra+YxPpm2gVuMCBR8ykRdK+p2thr4VFvu8r
It+p7THwS48/xAcBbAiFW2yfoQsFL0pPxH2DNHJ1888iTm1pBGr66rfaZChbgd6okb9biCXynPeH
Zd43oFlZOSRNZWkKfBaphxPq3d0FysoyZWKbpe0TVQtWN0mCYJdfjKIWpwleLIDUrgrA+YZsUI7B
LVkTGvGOLpurlDgXzwMy2+BbhiyRsKFrftOmm05y2je1eArjEgpr2O79STneUjQE5bIbuv8ZW3/4
04rY1cj3gv6C8iV5mVfkFQCfW7TfbfZUzIE7RmthoUz/c3jXA6mEIHDeA+SUPcTk7VgQeVkJnLm0
CiMHzwqdk0N3OlAq7LRNyDwfvQo/AFrGNq2nWtTiBD69rxOyLvCO6IGEq2n2CsOjVZO1nOgpL2mF
1Hl5wE1VhnE0TNEYpv7iKBJCZij/WG+Bt+jJDHDkmqSfMhz62hOIaZcS085a+V2e8w6b6vf6EKpG
XHNv9j5w7kDW+HdQ7AbnrpaU/15TJiBxfxaQrGnikyApjuJZkjo0dzHQz+XbDfbcBKMEn69FmH5x
EKcs1Lr7PwbZRNru1UYO9W0oEEYrmqwifAkzx25PyYNp0V4KrRZqa/hfDS+33uZPGLZc9hWoH8+o
Avx/joxtt0eYDodoDzIE8vM3DzO/46qwkFXjSUKaxKZwitC4wBhBHktIYr4atYC6SZbJxdr8Kqwy
NWsQnhVbWcW9A5D09aZGeYMNNMqiwQ4pL/ojUIXMsnWgOp2yCWdPys09OeX6//K7/FSOflJSAmx0
QQJWobF44T6fY7addeFlbaSthAfohceySGeTFO8QEtapeqOk5nxteDPiyk+emf/9OamC+kwD187V
9rzEVEcUWEm0TbFDisT2j779z7bjAWlxm0BriJr+U/8PmwDApZ57oWCacCJL7F60YXXf8RhiLxca
MtUo+Vy/PnHTSCf1inRLFHTEteQcjl+KW1UqZQBA82C9DeeCKdQjiZCFp3EasGNTB9hlmdhi1RTM
cQ89CNTg/S97HMXwL9fQjYeiOCgMIA9kiZ8NIQoMW48hmy6sDK9uX2mPCr6V/qtEFBlLZWT/1TvC
UG0IhdBnsGEV55Ncaf2dRWRRdw3AtoMfqNDbxJ13pHhnhxAwODBxPzEdu7ZQacAH3ipCZfVdNuSo
2jiCOLTumIczwysS2+YcqFFaUbQdnRUiipTRbYKP+pt0bmqPvLIcGE3kUgXFNswNvASZOti4vpYd
bx3GqLVcgvrPZMBQOXjZOT19jHIp/uaylm5X1TIDsvbTO/4XTdUyyJBbfLBoYjcHchHKO2CQor5w
ThQyXZtf47VfGUZdIERHS3IOAgIqXDabwuXuqaWD/UWDppZ7VgQ4st86wk7LBjPeaIZFr8VqALd3
eplLO/XVcCSJsI2X5LBiTXAxMr0v4hp5LhSlMdxY559YDT96lF/Bvz+GMEj41p7TbXtnOYWT1U4x
gvBkkqlYegP5uH6LBLTU++ej4caLw3GKXs4g6kC78uvAxiQ1/pdqQMms/fDUeB979CnwNumu0UMD
Cp4uBM8HgSRdTGu/8mj/pNR5+VbC8hkmGNhoxtpSmC3dQwG7pMQ3D/QpwqXm/h9UDOfxShFpKssD
fLizLp/MOrlHGj7COxJtR8PVy7aVsJj1d0Zdc1pmfC7R+LDwATWQ1v09WVdodrfRK5FEjEAJmksB
9+reHbAIdCLRnlHWJtcnnTbDX1HykXk/G+2GnW0s//+TIcf+yiKGYGp1jEzRaOGivkpP0tJLSwKl
i2fDzZZyBOOg8eSpTqeiFbKFcsLV1a94GJFC+yeR/I07dr+26h1Iz5h5eBgiqQWfw9MokBA6ngoC
Aa8pJWX3PR5Ep8ASIIwOkqKVYYuX0s6y4GLClf2s6IlllEj6H1nOiHteagwobk/H+5/R8gdBOnXh
O1FF3Alhfv2ubwNLs1PnkgQ5S82cedATkAPvSx5XOw8sdqMNie1steMZif7lxxfj7mJePnU9pJWx
K3I/yDNQ4l3S0ehKD6DIU7UzYMDtkA/0yO2t7tnRUQ+3Bzuensgfz7fdyv6nXLX4Zv4xYj+RCekd
Mev8gTCGq7cmJRO+TqFyg3ibF5CEI9SWwTS/l0ypqzeMbmxL4iKFqcv9FlvZys59TbOHyiKlXG6d
tp80ZuBgZmq2lIvOEQZ0sAfED1YiSILh6a6SXqC0Vm+OH9AF+NEdjsX8fTW4ybMRARc5SnQknIq+
LvyndTXxjYYmvPJ4zD6iBMjft4NU525gm8K/Vuqp+mQZ2hxWPPz/CoKzTBGP3vZOjjKo1ySgW4KY
L5WIWwi7J83X2IVCuUO7Bj2Je1qx6o8BXeoNeyJkWZzo+W4jIv0TI/R5UyN1DioMUxWQgTuYIXyp
JAokSkFmVUUoWlwbul2bUpi7frLxctZMCYe6mA+1wmEWn1/v/3EbFkjfaadXeAIVYjrKd0GFT2Ck
oVSZkMnHhgSW6IUyhMi4RqtuoblhK8ljysCOd7PON48banWnHkSRu9SFBOW0kzkGLGJB8NwEnK1F
JEkeBYEh1q4FJgEQpgfyTtgB9jEJw32qVXhvIOE7mqq/d/P8IKZYQYB80+CgxMAPUwXwTUHju6tk
m+C7N1aA99yTSw4YizvJT/g0/TjBNrFAfjh8OgmJVQETIpGil93PONU+14OZTeadoUcTnTx9KXwI
HKAbDDIb/jF1Gun43jNvsG111ZdXYbmhVYV3Iw9aYD613NjU6eHY/e5J6ECEW7FqHjdHE1rxbI7B
DsFGHV2bzhqshLo+SoKO6QmbrpzZL8n7URPRvdZuj98ZSUhruSg/F/8TedKHKBeL9tgiLhbU21yO
CVDXj+qQ5+XrlxvQ9eeKFVlYCYoJfroQehJXv6NKEZdlZm6gxqxXi4qbG0OtclhL1Pe6iTmo9nGL
SYj+B8fTzJM2apT704qbSjEC4HR4pOpRwj/rCnk1089lit8Tv5UbGAR3XEl4kUzqJ5UXdEWR5u50
X8Z9yc1OYtES+rDKzIwwq1bM71HGuWmfj70sll++aklR1j57m27R4a/yasEYQmO+iDmQif6VnRsf
NCiWHBMzpFBki2G7o+MN1qKPz8S04fZbBDx53rAOYh0bPm5UnNzBdIjVJptfdyY2OgxFhvEo2nTd
ilzfdT/37P35uJIDiyToyYQYRsrJw6bUkeFC3a8rqSpUuxa0UYxpL5sbibUVXkZ4SJly2hWqqnFO
3XQ1dexwwTy/cBJRyWCigZ7q1FIppj6ZDqjSDv9tmXWiatqqj7U8cAYv3yFyRcEfQ5gOhnfyu3Rj
uoMH7+39AElViWEzaGR8o81cm9Uq2WPzlSbwT3BziVbI/PF5pgg+NJUoUsKJpW7JySMtIwGhZqSx
uGrj729gMfDINtWfU2GwDKM3+AZvklaj+hW/aNZcUxPYGDtFgaFLOhVgZ+GWhnHOFJzCNZ9InEvJ
cGKsMcS62FY256UGQAfwOJBbmA2wvxP9PlMvQevYqzlD6VhY9i73B7cNzPcArTFbUnstuJdqdE54
HZ/T5ikvVw36BMbArB1NJBAnQr1qAlU+nQe2hKqI0q3KdlW16MaWkUJhWpi57mUgG5EVG7duen/o
p05/KGIHuGD7SUs0Ifw1+u3d7HtVw0tfdGYfYsOBVT8dqszqgt+eWzIiCpwf4dvjrmc4mXCDpMLx
x9a4isWtR8YhHCD7jG4PSrdlkPCsMFQ3pf8qykAzpTNpxFb2nA/RCU23niwRsu5VsbBHnjwkGq1k
3EWzURe9VK2U3sZfehwJVHNCKnfczdZ9VAfWXAhB6M6O5xnCNN+8+eqmOXrSgyAU/e9Oid99ZL54
eUZ4qlHajHwvL1kuP6e1NutQVFOUIvDIKQEgAOeW6va5xaSrQs4rBfEbR61a3QyMUZFuoa8dz9aA
KaffMo4ABIr/isw4WNNmTSBoOOkXzCPnmdBvXCDOQ0L6ueWfcvBzEwSY+6InVK348OAba5MR/Oqq
ThHzjS8enw3Ft2giJ46SjTLu0hnbXlx7ti1K1DZ69tUbTzGJpn7WK//M1wJacyIT/K7IbIfaBZci
vYGhiFSp3yzN/Fo8K4djH1nuG47L7Pidtg86/BjmM/ZOp1igCaO0XRCb1B6JTyib4qGN+SwNv+ym
z2F5xZlgPzcMzLM1DBC/6r/tO7aNMfYzDxV8FAbegGO/EEy9MZiu/FwOZg0DxS9DpE7dHHuAhSoL
khS47vYySK9hw56po26P5u0/ObjdERbOWWYoOgIyrRE2IOVQ5pJP0XKNOyGiLwnGrWfLW6ZOtqei
yuhGcwLjjnS6Me2/aaiD0FFfZvrLHv4KvPlQ7N5GmndsEJ4terXFkLYMkDxXC/T3B03eZ145my3I
FEibUmvp6YcBk5F49tQ2VOASFEHushoulBqzwD8OJ57836/SbpgXaaGbZSigrnvCM8EdlmIf+MR/
glzSyOyjd7xRSYt3MCMNXuQtysnY8kncT6FnUBAWKbQOpuXFc3pRT+qZK/LqnkidmiWqpu6IwQKR
0IuJsknkL7FR2pDkjn3qdob1EqVN5aX19F2HGj0ACnqlMyN47KNfpB+ykU9FgzjfLNdRlP4cdc5n
Z4PCD/CNs1of9J4tdai3uLcku+uTwsWxyopUxN0nLMN/qPbsGnwPqsYHydZUdcZgONfXpyJlmfqw
xKliIjQFOpXTfeoSwTAqU+i/L5cM0Y39nc8hIYTcD7dpNjXkn+D7Z40uJcts+ffctA/S5d/jGuXN
Txyjyzd5EA6EJnZkiaiOlNgu83D0G8L6Y5zKCj/4VvJIyigT6UtDCjEA8CQOYX+IarXrXKityX5C
yfbbJGpXaUCwxGamG+Jm34Ef5RGelREUOcM3Td6HlDIxG5Iwrpml6VCa6AmMFOWVfxo/z5+/maBU
n0VOd0V1sZuSl3gIgKkxoiMb00LtmRzaanF3b3Rey7eBHs4S+b8hdRDzE0ePFzEN6txkZPkfOHm4
IvMJB7V9o8k08U+NGa4OWKdwbAaAVl5f3nS9JDWiTeO0cYu8PEQsASdC2XH8XJWUaQUKIdQl3/QZ
6FyK5p9GP64g6tnfejev1HjbvJqZtxAkC+NVepPipcRKwSf1enga2EwLQ2CgEyc69fXzjcTcKyTs
sh51eBnXmu8a6qhd1/BzYrKt9l3B961vVcvrTBKhClTQsaXo3unIgpSqJ0ikEsrqALU0zyiWXXr+
hsui4f/0BGZ162/0ijWvclxH5h2g7rgsrwwfuIozPoNGOlVnTB+wbCupcdcFp2wEw9vjw7PZ53aN
4C/HTEb07i5S8xcYQ9iR3cp6BtSkHtLqwxqU/L1Z/59W0zMBzhiB33f7cOY9u51rTKl8jEvEBg76
kWBciIs7M4OFZaQVstUtXnthzfFUatrCH3WH5x28jWDUFZ2jb2a2h6uC8NodywnyywI18UZsz8cC
J8eH5Q+IQw2e+yBBMIqKWCgC3sEJ1dhQ94AsdoU94Vw87gTi3wRfxunzfNIglPIYIOG3JUANFYXk
vz8sFo5zHsz7EaUzFBDNesaYW+aUkQKw4pWJcMMPyew+nkGV+zXXAInia/NncK8IG1lYR9mFMe8L
KWVMcYo8UOYFnGXyotYkk6IOjA0bu9fh7GPsGa8fBo4kVmHsyjwGf5nO2Ch5CbeGzUlKmNLJxGSh
VMaXyA+vMwa/jesXcuzfCjImEKX2/8aLc2u1LcdyCMqO2XWrm/LxRlKqurWY5+uME+TWZjmVmCyH
CziIQcQjxn944tiFuIl9k9aTS9xSOxPtt+wFXs5IuGkSgvWCZLpvcT+q1w082YKV0HMpYnyJnemp
Dq04AgPm8rig4bCpB+AN86m60rwSS0qOB0FDTI2lP41s4uJYytQwFb/4yMrGkhAP1SqP1kzBEb/g
gm7PFc0aNisCc5gcSrGS9/bVTSILQ+uE4YmsDdOJPJC2LIzRFY1fJNtv9MlMq1fDsHvf63JZvx23
RdhVDdf5Kh6N4UMflI89OBMBgaq4u0cqgcL72nJeUN+avXWEvzgesWoGAP1rouiJq2tnj8CGGIB8
0rlF8At7UjOfLy/jGX9selkXQz1S22pIopIsfLvRSMfLoJibaIqaABQwLLJPMDfp4MrKbxMwHePF
MhRSOMsh9A2I4qP0BHv/7SlszH17+kkXhWR9KSBgTDfSKrovp46xttsTkb6QRhbqCrFcHhrv5Xla
+nd4VkIi+cvxbn6cEh2t+MObruTsSrYeVtIvXiihp12+LoKyf1++VysrwVINtNEJa0uYPSH9s/i+
qRQk/xujs1LV7Jmjx+RI3ctriugvE3A5vC9Z4DNQzg5a2++qlgxZ8z87hRXpibJO+tWdGe+81sqA
LEvXKPvQysEi8uedNPmgwMx/TZJb13QQsdG5ir0FkHrb+XPp+aLFA/dxucLSrujnC+bRMtSxx4sk
Gwi/KvJ3tTqkktZUeTOwahPMlMDpV4ZBa5nU2CIJHjLVxHHdCSxEzv1nc1QgxGbNgL9P3zjgBsGT
AugO4rNjwk58tE1C+6yf29lXSK3gmnNigxJV2/cSzBDs3Y7mEp3t4/z4gs82Sb1QiJcNiLPIIxj8
yzTmafm7JdSqXh9v2pdZqHpOEeDkyjYZUk91V3e1Ujcw26aEGzd+14rh6+wY189UqZr69T/Gyyrx
3EePlGMFzQ4zU3eCp83r6n2UvltGb3u04Cx5+0j/qEga6UTuq1yf8f17cXrPpmaVVDQsnoRpYd00
W1RwkfQnDBqfp8y8b0mMMuhu5yEaiptV/MhXUtbCK/ltdL7FFiOiekQ8WlPAVMnS7w0ydtwGP9F1
XHJYoifenluhDuKveHyWFwyLQL/d1JOdUnVM1R4Tyo8hzKfJdB0w77obw/Kp5op2ys345ymne9Bw
fOqv7oPXdiqhKkLbCQ3sA6SKsSTJrrdQ/woaQDcgkNfyW7fUA+idloE0LqJ6iNMWJwYRhMauA4Dt
PTJitqKEQnzdFkaRyTX0dzTDbSfhULcEh+tcyZR06Qd/ySSsgcm/QoNW6tPxjrTAHumjrA/GPrT2
tD5w2ekIFZlei8gV5XITR+VSSM2Lqfk3CEkgCNyaQBQ63exV7BWG8M/ibFbGkY9atKHA99Jvibet
v6T7xLqVKdTI9eKcue3OBLwSeFKZJ+663vE8yYH/vQBmmhZAJdnDqXoIRf3QP1qa6bZ0+9JEukEY
tklOwJS0pLa/pva+KsBlRHjVWJ96XQ3NNyVZL7sTzAfB0lfkb+t4/MTxDNsXnMDQHWc1dh3XfPMO
bRj8n3YaKoQMrcUv5JKwNxT7oIOlRNRH+oVKVE4dYsVPjiF27Ko1pp+HCxOserwkT3Yje95bxmEx
6RQKA9uZ/NTf8DLuiMdKcQHWyDbZG5JNxtbjnPTyML7klCA/4jtiyMWEI/Vpo/zzv6Bd9YT7aRtT
/D3I9IJ6+plEk3WFLVPy8BdJ+v2HvuyfEGLH/Swd8rb598uVEtARYuhuvDsRkeXcuvc2CfTe2E2L
+Lotosj7D+O/zVkH8Xdvdg7NWpBymCON71Zcf//wl9X8ebHkYYzC39HcJbiq1hLTrBIIAGuBY0aG
Yf/XO42XcwOAVm5cCrSBjtJyyAbs4YX7LQUD5YiMZr0ShB55zoE3zQw4au4dbj6iyZ53JhzpH98k
dU/aERvr6VdA4o3B0yZE0xjpOOA4YKPMs2XP8GgDqDlBkPDXfpv/R6jpj9u4YFI3AH5lY1zC/AgI
Bu6vuMZuHoCECDe8kPtLK958NYarGKNv+rDJQnOFuiLrGQY3stAwfPpHr5duVE/O9wneRE/0Y5H3
ejQVlP0VTTSGCJV8aJSSJWq6MoDW6NdBtUUHDoVhjTsiWHBdNOsaulsEuAmS0f3CYEaGA5Fm3JKP
ID0ZMNLAtia1pDmx5T8oaS+WiSKckXpnP8QejMHqHcwlBceRTcaJiU8LfAlymLJKFNn/kV5X31Pg
SLA8kMW9t+wv+xgy4n6yrcBPvWnd0KUpITVTG6WTVK2T4Rdp+9mN/R1fQqPw+CtO8VUyWL23rZdY
VyhLTPpNlnOBi6yaiLmXESYfsL89Bxpx6qOrdUqxinWUob4tH5wZIpRJ3SiI+ACSALq8fCyBmtBw
JSUqLT2Fmk1g4Y/XhzKL05pRxqVLAHuGwVRdottBBi6aSjAT/zWylS0TKtFumNGpEpcRaxKHLudM
g38NAoJqZCChLfNhjhun2xgLmT/uzE18QtNDKC07LtaiEbkVHB6elwKg/zotBs2KHSBAC/tyKHBz
hD6Fyng0FKBkRUBE/phGzXMHeMHvMFaITczP/guStNG4T3QJnIdsooM+ExrgxWHnt4C5VUQ4DrFR
3R8i/Uo6tHz/Ums3sFiq8BKVHwcJOWisOGwmuVf06jCyfzvh1ZzyfDSbM3ZOqtkmGlsy3U1udKBO
eLfe38sNhsTDQCRkEjFXdZc78gNvinGskSeovk3W5mdRwsDhdK9vEKXVsjqnxIOFV0ttVYe3XR9H
GRH2gtuR4t8f1ZjWI9LNaXsqETRodklYdu0hWAbOMTBH1H4AObHoQf176Htjz048pCkMVm8Xz959
l/eTBg7zkVxEpAPzodZVDEmZCp4VGpCSvoVAYr1R91YZwN7tCvBOwCBVgFMzzfYUSEhMeeWWILhM
QiastrMCC+JRoG+qz8KiZGsMdE/W2KkxvTtEjT6OOCwQiL52l6o07jpnpdIIJ9l1hXS2cEn5L8Sv
YAzLvmOc6yAzjkae1R63QZfeTEOD/rRnEuEx2+6e+gfY3ONBykQsxFckKuSG1lhwEaGtyUyniKve
ZnRmUl0zFjwIOcYwQq6E4Gt3uYfOqoVdNpENslBPiuD8+Q2NzwOj44uk+OU8eqevcgL3PLNkoboR
9Qx8ArMPEEAQdnW/qcnT9T0HuB/VgreH0j7889DA4lmTiVQhrxQ/vLaRmgt/+q7L8WyrUgxjPFdv
QazrKa+7GM1G9wHs71wz9CFefxFMnTBZRB1+YfUf9ykP3WRbgYNHUzOtTfzeeZcSkIZO/sPf2uTd
3EzZ0WNo15PqlCzSsEZ4nm0PahWJPOJLcFL8afAYpqpggyX+4V3xvtI3e6EkdU1pJ37Lpd5Fxwid
/A2vZLSCcah4XuHOPtTstWKmwCZjN6aTHHp0rpAetfagzW1veFhHAaGVxMyQrDOI8ncoeqaTjaKj
w3VeqxTaYAvenHm/s0NoufKrjtKT7D6KoQeT2Lu/LOxZOmgwc/Vn+UAkx1zxSsCyBd7hsAyVKmNm
wiVGnvhwKzw/hvSmxAknVa/lnxCYqe3yWzqBNoMW8oD4u7F2VKahDOsfLptPot7T/4AkvnmfIkeK
xuZMvEz7szldxljXHvjOKioHS+4o8+FdIzyyG59Kjk0zvLc/+47RKyHDns/3ORSz/+tPUp4xflHE
ueQm9QfpxdGA40NanzZwFo0EB4NTaIV98QrFdDgQS0eVvK3GQAnxBl1yHTnu+kh9Du/d0/PRwQv6
ljpIg/9pbL36AGdjX/UvvZMoNkVto3+jB5LZtHNcg/YP5xM1DdMikS4hpqKSu+WeCVEsMaulUC74
TzeEmZLT9pMhliRDLRqK2veHq/lIyo8M6Zcic4aW+sgiuOHffblp92KlhAvHdohzwYnDGe4NO1HS
IeEOAGLVA3lSiGc0prbuGLTr5oRi3tLke/qHvmsKFzFLHBdtPAt7885l8YlLGOJcadQKlard1Ese
1EZ9VXXTyUdvyY28jeA6j7s+H0D1/Q9eBZHxPz1ysNo/FRuviMO/eUAx1YSycnc18doK+GtuollU
FZW7dt3Fo4mwC3ok4BaihQkXhcu608Wkyd6rRlJD6NLNjrpvMwJOV+K2yF9SzzOvT8RcgWM23Mt1
ea48y6+nCN45wCEZdKDF2DGr32QwWWVTUxwx61xHe+dgM7AJ6Fm3tC1XJeTH1xz1at/jzJ7w4vfV
GoMhXZvcLV86VZCg85nkyNBSQp4gehGrzH+nK2YFVtJwIeIMW29jgQh21TeN3+7JEV03KahP4zjN
1a2V1vLayzHZSS3T+hvDaBFEN+D1IfM26iXKwkDuXSgIBz+hpVKUKUWQtXzwoTyjzBgJM4qpsu6N
g7g/DDFQ3rcN8tnNr+4DjA1YkGyUWaHFc0bbibgQuauvmQC+yZqg+RUSGZ8wTe2rKzDyQIANLtcY
Tct6ONqlBCTlsTZjHRR8ibrM0+ttR5/B06HJfNpIfxtX+ygI0H9Krh4s9FDxh11ps313C6/YJ39H
h8CDOpnDsUAnvjxpvx5lrO//ZtgQAxplcu/D9Fq9meuZ/tWogyZcPZHrXicCBn8HixpuZvhyjwHj
S4hDPUkOUlpPC1ZgAKnCVBPAa5jrAALtjxUumf8h365K3+XdMx8SxStPNpAx/OHmDIxph+IUrbOo
TbguSJngem2gsrA644aEf1UUA+2McK4aA6u9LL5hKlRxiGzp5O/TXMm38d0PMXQ6WMlM3rFjcHLV
k5cInfaS4aVQhR2bn8GXQcxhYXpO/xLYOsGei1mRaulBOBst3NnM79cmaMu6o4MM4uFv0iCh5yyT
rKRgd9JXr3TRSTS+255WR8kkEIE9hJUlmy6zmkFLXj4LxLMkT/xd8pk8uoRWcxqM2YmJ2qTZ3OLU
QKLwnNec3JqYKatEiPqox1oaA6uBwLzUcQt+DOUIIp34YnFl3Fan3a3Ryx+lUscfIam5PW3+AYBL
B2l8EZC1eF9ntoZuL6RM/4Y23Wk8isa38LRk3XL+ht3N5ZTdjU77pyc9dVWxnW4pqVjhTEBph/KK
xJwoBcQhC9XEslKQG9AKXOttVl3LP84M5wjpilh0ktDEUSriUz2encpUj3nwddzVfwz5X8k7dyU2
2FuRLHHrkZgtQaXm3jXGgEG6L+Gb/27G+rOaEqHqTybwQmMiX3a6tsQZj6aHuZs42sh7WW207wuN
xw8BbTPrSyCSIwrxblSBNmsXesLF6To6NmFrqMFcvDsbHwktsyMnitoC+hDQ7c+hDwUjfiCITDTm
+5MBAgzCX+x7JGZswmN3y9uxhJ92A38gCisgnJlz20DYFwM6rA5JtD3qQL2tdWQVzSq7iwG8FTN0
TcsNl808g5p2zLsEfmvjjQh1f/ULHgzerkA1xnU7QHj26rMOI0lgmRnXJlWD3i2ZZbZkXuzmkXYR
yKk7ncqu+1pZ9CEzt+9tV26fB4NkWYcBe4yG2ABwFTKZHj8AcIK6xzUNgd2bW+dLYgBdAU4RDAs2
cdnlueeZFp9BxA2WMXvOhMpMpDRcvnQCnCFVSQiOCNbl97/C7tugoM92yW2F67nOiDYsGmP/JHBx
zaMhkS71NnySHW9fL5loiUvFcskLaAlplwShlYKJXRa4G1njUqZMaPXyAzZnU3S9JIRGuo0deGQY
GxpgX8voJC2oeS0s+N6OQwzpimW2ZSCPTFdpZi4AqVpkiV/3Fsqw2jOVzFcXn5Rfok2KvQ7QxQ2r
HM4wYH6ZzuOzVww5LwyPKDS9V0t/blEwt4XrioIa8p2htYPgT7bxbG0+l0HqIlIiq0r2zoellY6h
SPIvqrYLl7VFqCbqmUWpw2m6+Oq+c58cO1zEtoUSET9EsiEW7T1vjQdS/quJ3pKK+xHikVw+e4zP
7LgqjDEcZZCbBY4fJvGNdGUdpaapv8IZTb4jJbAXMDGI8Lwcqq5C9lEspCXRHSnyRrBkekggisxB
5JNNkZoOds3pLq5xuVBSA4oqhQDUWHV0KXFLkuAyTSQdTpNHYTlfgZxQxSNpeTjTHEoJZjyYCah3
5PTVfxhjOBnhNbL9gN+eEf8B0/jaPUHYdQg99xLmFPTnRoIyq40bvElVV9H/ooaOsgrVs0Mvsh8m
Stm0dEa/rIYhYNQ1mZHUJfUHc8dneFv2WBFOwGkaN56bId7YkzxjZGGeI6UCKFYdEev2bBWpDg7d
8CjDfWgjHo6aK2kQwbcJujGTLt/9dvh4s89x5tAYSD5V1y1maytnQRb0UoForFar2ibfMUiZD3Vn
D9T8eL0/mEdCB+FX+/pYA1uTiBuhRCPQfKdp6guMmZHn6wBQ0qNRg3RMiBImoRBjXxEbSWgKt76M
jqUkAdifWXrEqrFnBlDZ30BjhXjJo4WNvFSBoGb1vxLoR60DdzrYn1k6PTqXTyZ5lV0CWaiPGQXS
5TAZZMwvKBcfitAgUuo0oFxUWccuqilRZe6BrSi1y8dsn9adq3qo69OPorGDc2euVKUK/Jp7E+5J
wKhg9CRGd52rR8M4kS1Zhmm5z9JgengbI6/pYHFOWrnIPd/WnGaFhM/FMYl53QL9JGa0262gwWao
l5iMIyl0x8r5iLwvhzkAy23PFJr+6viY+BtlRNtxIBEr6KJ6x0UDOV4NFP4gKrVYagUCLy5DHbaL
lsafS1NqdA4y+/fYpYvtYEVRCdijNFAcgC19jXnFy3neOsPZUr0/tR22ADoVz9IrmOpx5U3WPVJL
dbbyaGuc5oqfxIngmaVWEXQx5lxaAV24gjWA2AFOtTBERS8GticlZyhEIwVK/E8GUE3nz8mtQW6B
5wqhDrxhWtzjybYs8xLEXnvwjYm1WKTI3dcni0a60gNB9WVT2ABKdgs8DJNrY8xdfspN7c21rAN/
wx8kBDDpK3g6U2nIB1zLAwRY8HFzpT7YgZxy+gJPz8T1N7C/Ca5PSLJkR+eZR0PM52sKSNmrPou+
FNTNqCRBl30aGuYqO6aTthAa8FofOVL/YOxLEdj8fBuwTqxV4gAC4RyEk5609+m/P/oD2kbsMT6P
TlUU27LQ2qNxx75endNEyM4Ns2IcJVbtDlyUdlFubhQ/3bzGj20YiHSQMHTjgwG6hUj/EYAMMrX/
7wLnpLmpvuFKDvY/cr52EBmRM9ndhpebprrTE+qrEGtCtB30yh7q1c69QjKGOzvoYiXPi1Ws/hLD
R56uMM5UlrNFVHDwF4LmLkAiXvgGQ2FEsvvDt9FDBf5Lc5ZLHHOIs6M2wlRuP/OMPYt4DcTq7kdu
r+RwbusyD3jYDUo6L5rT4FcKhoxfMcZAW2AISVmJA4LAOjcjZzukPrIEGSJg2P5qlcJPLGI2b6D5
pBQiT0+i3LXkvnUzZT67FDTo7GHVMcDKnOBjkg+PCoE99OC8wnsTbUvB+e1ipHCR5O2BMT95y/gQ
26lmqJmOFIfvqXqeHbJQW58EyjcoVdklmvOtIjrO5GIxky0cx2wJLMt1a9olxStuPd1wbgqFaoj2
Lo/C10/pgyuD3fxf4fMolP3H98g87LGA23fNAGjgXCGUDkVNz87vwmiutgIZiGmnNKBENR21BN7N
GWNBrABrEZLnqLapqbaMPgWr/2wQo32IzbiFEykkavW5RmgNFuWV3/z/9dXQLV6YHVrsWZayN7zk
jda1mh+NoLWqF6uPVBzqbPZE0NOux5sKd9Q7STnHK9NjYRS3pmz60Wnmh/Dkdsu+HG7bIZjoOic1
fTowoM2dOs+TwNRnzFqMTJPsUg6EppoFAX3Wovk7ba/WABz3L0fJeuzt1OmDlRYQdbVcR125/gn0
T/FZqkMIjCCV08M0Q78mnFm3/4eoNJgYsdosichiJRLxM6A3mP2gsViEaIrKjb02GDX+9HfTDvxK
XmzBymFyedg52vDbUkEpLqnl7um/qjg0pGpSwfb13quV6O41odWsb9IMROWMN0MVlj8jfdnrOPCf
Pj7DChzVYSakpWsiHtVdvrdcme8bSCx5aJyyVocXp0R5MHZBlj11MVXFoIJvhktMiaLrBPtvFAX+
lIH0znqMqp7d18Mh+rYy1V4QdYCgQ4bjzKEXDEqwBmD6lJmF069QorwC++gid1uEK8pcgkxNM2I4
sB+vRXUGXtY7BRGtfu/O69HeeywY/qeOE7h0UaCRG1k/chkSA/QADAttN1aoKvq5QT+M+Hgpw0Of
iYNzgXl5pEf7XWmSYNYIrXn1vYmODVMkR3y90C8IiVprZLKBeeAFXVCC3amfpkZtE7Q6k/HsPB6s
TJOuKTuOVff7dZf/DlqxgYeJscmMzOrfSP5eJuet7Y9OZVOE2ZQzj6E2HCSj4mXBXyn5ZAMkpRZk
BbPpazEi+LKK0AloVjxWYuMqXz5pQ4VGcmR/pmbCuYrmfDeqJIsHSKUA9yfP4BVka737sIhMZ0zK
v8gA1xWj27AhJautKe6FstyEFHHjLxnt10EwUHraLX9YxopdfAIwyywl6eccqehgTMyFRqxJVJUM
OFJJqvwGBDVhzHWGi/TMBYEFT9Ij0jKkKiM8w5g7hPMUrC5XufAggKG+BPLF9fgvI+5pul7DZ6eX
dDMZlq2mv90A528hzqhXOHAS5Lpr3jN22uzhkRvdkjQoT4eYr5493jD2bkBCHSyN/s5t2ZqWoRgG
BJN1a5caYnggBI+r7pzZ2VDG3SQ+0nG9FSdjOUBg8i6QcvRPZ+IKtMSOT2e/tZ0f3ERcGhJ7U0Nf
gTuB7m5sfflUPqvqXK4hB6Oygc4wqWsM6hrNEAE9Szjk7JxdpYDdIPuuiv29AJqr0dNlkcTtzALh
OGT8dZzn+0wciQ9s0JGBO2/83GYOTttdSUCasL7U/EynJCe2DJWzCkIg3Hr/yVQTLf1Kaf7m5QV4
J41jr3S6iIEwWeqw2Lq26VaQY9LIlNIEwwUkD6/h36yZ0UY2Uc3boKH22rELBKezQQic02+3wlj3
eFtZtyh0Lkh6Slbx5j0rn+CTz71bI2hZ3sTV/w8ff0nSNxMHZEU27mvKX9ChfhDH0ryDSmCw7lGu
JywWK6WFWTNK3ZXKM/X3HaNP3HFD4MMgtP6l/cJAt8Py3dZyIBX8LFWz5RHqOPqzQ0+BJ0MPSOMj
MnyoDdaPuM6ashmsFo7LZAFldgKIEaPKBgB2Dw2fftO3jekFzar+liKvCmedifTJXG4AhDAcdIUT
4aLYMAQTHubZ7S9+FlPfi/HkcGLtqtsVfmkbI/sW1BnXDeReEvCAX4mi0ZYpMX0db8hpDtHvgfx8
T8NYbUjm1X0ykHcXpSIBij47RWv/M0Hxo9QlUHdoLoB4rVxzlZaEkSpZhaYMN1QCacxoNJ5JAzyH
L4FrNXQrcLGAP5GSwZadUwOoEB8lv0B+wRYyPfjQ/NxeN7Obeec9keZYmn50jXFU3Ey65DOmQu+p
MxNyV9+BAk3SOsG7ilUjuEuVWrlawyNVQUGn5ZDrrlJ6jM9X813gjT2/D0+13xhFBbFcQ2BYYflU
zOseuvDJ0F4ME2jK7jPI8amJLLFIpQQ0hxzBIxb6sTRnBb3HZw20ZQ09h1r1ePUG4bCdKLpxvpxd
wJ3cc9/EwfEOSsG5W/tzMCKYinLvfc3xwqTLhaqfK+HS1ogC9q5F8/8m3e8vQbtv7Rzim+nJrDjT
3WV3uRcBkRocxqClgOnY3CcghHINWlIHmAPiR58xcLl4WMO19eRZlqwyVih+UseEh4le7S/D6kMt
pn8O6bSkaw3KQRRzhovogNHx738gXab351d8el1gJfN/ixw0Ngnuns0TlkB6MsyklLqcnz5h/WWI
s+FxNcVZKvTDPMHcri4fAjtSuN5ySgf9uEVOWQXhT+6YQVzGahkoRugpGjJ9FxyiMt5O/fZHCQim
y6sL1bTNB4KZ054ey29CIeEZz5z6JSzV48gZclHIpNLVu7z1cRwucOX2VDvPsI1dYY6wfMPmq0Cq
T3Ne8LG80h9agDH7ZUA4qa3m09rMl72ms1tcfKEDKspupe/auXE8iRGXFdvambuDosjqoG1mCIb/
maescq+w7WbyDSXmLGcy3F0pTk7GmTMaUuW75lGheBJv79LDW6/gh40pfSlc4lBi+arltLrLi5al
shmDHyqWYaBMieyMd29BfR7ajK2xYXEo61FkQ0i8OYrujThih8Je66xv8d1PBDJri9GMNgqgamgM
zVLFcTRkXOz+ZUvIsD0fkuyi80DAbAO5Z/VD6CO0OZ+ffRaTs1Rt1My2wX9GhvObDR6/5e+L8K/Z
6d+yjrQuLTyJOz2/zjukRqQ626Q2WHgaswjoiqnNi5VT8jxteqf08L6WNKaiuwB6kFEtqmeAAmXl
NkYe0YrtM7XyT+JoKgPR3QKOHBdHYCS08jYLmp5x2oPPYldZ+/0oUx+NNKgZbSxxxLDlBFYpGx6p
rXW6EsKoci04GIgCh5VLJEtPaRhJ5+nZP8OWxeL1SABtpptN2kILVd8PLbNXBDUEX7E6j4hXx65q
gMzpDp7P+EaVbyZe2ksvn+kfpju1gaG6Msx4yn6PdhfackuFuUANBbWJ8xZUlPAEnupqsIVTHkuW
CTullfPqXxb5BbhcTZpbcjCi9eYg5o/Ro+GjpKPuXxcsAauoq0CAoA9WnfTVBSNWbH69hLymOybY
xFsBDlgj14bIxRZg9HyiWi3YmLf/zd2QzgfEb5dY/1Y+/vGDjCDsCIeMym0wpjg+1lwDLjwga9f9
VlwBhDRNGWX3sUAJKlS9swIel7n8Z4D4RzvckUubgN3Ok3V0FyL29hLT468DAl6RYvsZVBs+ciga
ErkZayqSQbk2Ge+6jCfiPbUrCjGaoo/l54rPJkjGyRxU+RzHhM1u5//LCdiKD7wNVumgakGVxxaT
mRrrjdxvLUD6wb7nbPZxpeLOEt5FesR3Fq00U2by7w2M1ot0rfAuITVr15s594i9w1MLvRMRdUyF
bldcusFTZcd9TEKOGBWBRxoFLpata1fps4grt5G5FQSN5Q5qoZYXT5IDQ38vx3HbqKRbtIPEV1gv
7E3D0KQqPg/ubi5FUczXQs8BleJXGsD9pSEtjHG35jHx/utk7XKeJi/YiFe/ATD8cW2vmTErDzTi
yVkxg9ovf9whFxHW31qChO1Ztbti9Mb3XW+6bzJk69EuTcfsDIuNF1k42vgdyn275r5lRy+l20pL
WwBr4b9gP0kd2OoZvAhylv7HulmVTa+V7+PPzwTjlZ6LnyUKe9FWOoCpksMdUmbuu7D9uOnGugJL
6i1ciY3xznzFpRafxK92Z7egw09uxfvzobsk9gLjsNsHJc4uDA+slO4fhMvOTevIyN5uiXfME9LY
4YkqnOyZqNCUHVfnGXeMCXByQv3+NpmKEEaP7zva0sXvH0BEfhjqWuDWw85dXIWCDEBzOoKC5UHM
qRO3URJh5DtT0CHpmDzsi8urFS/BoJYeooqnIj/Be0uxddeU3yQCm82mxYs77FoDfRjpU8W4ezMr
ggxg3CIVEFMAQA0zdFglwbpYodjw49QOZ4YU3en5Thj9potBs0IX9cdjbbR8N6/bF5A5CstFJb4V
xZfKN34X+xmvSD8ZA4c+RwT1KVd9UZxTo2B5u192f9GRAkHHRYV9t/DU1pFsvBC9ILXGJJrYSrYn
/EMYthfTX4Hj2h+zihx9hDuLI4B9pXXWgYFU5vXxHBjVO9eRdD5Md3PnBrJYWsQ+rUXZ3PUYHK6t
X7XfCi+TwPE5onNBFSeEr8+xsBPSAjx3+bMK2od/Jz0ycGQlESiM47adryfV3dAqjm9LTV5GAudd
tjXI2A/BsvsxRXQyjmeZxn0sEcrsZnIouqJqlF4s4rIJocMCHPofKWd8mX8rqeqaeO2bOkY6iJI0
i2nZmYqPLVPj4JbC94q4JFlk7N/4kFq54ORK7LM4Eo/K6CT5nyTWs/iK0MeQ1v9G/3IIZW3JmnRm
OA8MUyFYlAVhohRir5ul00yy4GSqRS9Rc0hy6tGJoWLQ2VErxrNd3BsVtXdKrY4D0MvSqlq+MJ45
36WOREdr8u0I0lvUU5BYCeaItyIjA8oeEQu/xOpk9fP0xdTRjK0dW8TIDBy6Pkoqm4eKH6K76yrS
J1pNSTqsBMRNRB8cXz7nArPbk327x+WewUpIvFmr6QirEsmBt+TcoDDvKPiP6BBTikOa1VhZ+YOU
ryLTakBKjI3No496WvQeWIP7uJ7W5kuYhkHRp4X3hfu9s4HtQiONIAoL3LmBkckHIjK64gpgD9P7
lvVp111BN57+fF6gaTt8AcduN3a7hcJR34tl6waerKNXXdUXTALKAgdgJxhPHexZCEsufZGAB/Yc
nUM4Jn+B+9EtMsPoEuMuctqxlw1gCzc1uoCXFu6UCsOwQNQiaJ9MyzJoo2rEAAE7df/cL4AgW+qC
VZCJT9PEgLSasciBhewjAarJYDN6X5hJqdCvdCMIH+QLws5cW/P0rF85Z3WWIXA7yG7uNcut8CYn
9jpI/Amwbhdo7/B7wPUNlQBVF6vJP9whTe5p8yrCyoxyzVPsW8tIBmbrPrEu+XoQKGdE2pztlogF
fDzts9hlr2SgS4gfB6AGhAZADf+NafwEgd5w31lNVn+nAQNS54HUTZ+LEDsu4WK+Z4wLN4CrJK47
QJFI+djZCuDvv0JgKG9PJFLOYIip6fvsx0H1OpCjMu3rkwkcv86hXo6/SYbkrymgs00lgxvHrY8A
jgrMrKQeFPhx45CL1alQHbK1JP67qfXaWxebGRPF+3aQ0wj0+FkLKWkaWvNJVrjD87RyO4tO/GFQ
FKTJsLU4p5jy0EeXsdooNTGMV9yydLBnktrLt3XT3Gt4S94uCm6/cYkaqU5dS174PKTJG+WRIlfE
LC7R/xQ9G9MKZzieZLZ+9Dz7vX+47hM/rM1MIP3DsOR+nvsTpIUE6zpj+eNM03MBCymV0NJraekG
vHCDCLsxsk3jYNTtm/ZAYQVEPcSPgi/b1oW2orlxzsnGe5WZDIhz6Yh066J0X5IvC5zbXMz7wHfk
fWQ2v1E4hsslF4nQ/kfydtgvq1u8rLN1uEI2+j5Ly0XXI4zPtpwabaQrlSNshJNn8iGyW0J9YoXL
V+xwyZx5SbBo5Bu1dHBfAyQRmq+5/f8iIIbn3d7WnztkpRjCYEXJVosPshTnJF8TLviadRrai11U
taMnP/aulfbk5m7eg/DhmVe71v7aZtazRdK/ylGlQxZMEOVoyh+WVANGhRpNRfz3B1qWwyFTXtUP
BYLql+A4ZKy/VsDmRscah6L8LA+aWdLILVLvO8yiOMINqa5vr6IWOQsfSekRfO3RBmKQvLq3ei23
D3bcx92nur7y5T79PzcwpsmHv4SqXZj1U+4DO9FUHdENPDhuux14M8Fh6H97NM5TOuCBUSk03/oQ
ZTcuqAwLdXPD0c0R2jbImWkdtHvm0y48oUZk11OxfWpJvCU/SJQylZoZl8svhNsywVdQP2UH79k7
wTrlXk/EFVexM7+04I22xOfVtIKCx/9pQMcZbK6opr1vzwyZ4m3ewwdBvS9FoD8Uuy/PICBAKrzn
7E0VM99tNt0BbTAWyO4Q4e/AZu6x/Xo2hP9fjdUpWdTYWP04AaXVf6j5TqLZadxMexPkikxrHnK9
Gi5e6HC5LJMNe/J+WsvtgRG6GYzG2w7uILfnPmkF/lZWNqdHC1NhNXouov+meQMHib8kTl4m8bQL
HiEyHPWExo6co2Q7SnmdOAbEHC8JGBZ//dASzi+4cQFYevmTj3GxZLMYsWCc6sGE28juETsvmVpg
aruvhIe3IRafDVzW6E/pri9yk/ihfkZ2Pt7Vq/tGgfADcdDWGA2KuG65G3lpAPzNAiZA2g+oYL1V
wObJ6Nf8L9xdakBdp9P653dtEaTRRRGJW9ReLKhfHPKezC2nv+YpzAc4Fr1uUsmiHeCz7FB8aY6/
6iVOrQ/bacmO8pRMQvILffkbiSEHK1NTLQ+T7W43JSrrSpZh/jOcDgQJAoO4z9TU1ADBt6iuSZgW
jCr+U4m9nLT6vrRKghCA08AWYtUaIJwRkwOe5k4ei0jwEYy32SMnUmetShqyVDCMcBM3Co0L/mwr
KykliI0UxU/6B4TEuxqZKi3CIiPdO5WCXaBFfcXMR5DBHBt4GrK4sjFSohHFWSfQQG22szsgXoV6
TxJMvTEjFjECTdM7r5FnWPRDMquwNJ91uM0oEqanY8sSKUjF+s9oYiz5NEgR8XrmFLSMQ/h8aBtb
8n1sKcuHTeyCZmmOVE+hHAn4Brd3/+Y3sQ2a3H87Djkqv5ow97lQD0mj4pIOCJdTIpO2+8B2i9G9
4TvuKbl/Ltfvm4NqXUfAB7rjgvfn5fICS3zNv7T4QHOExnKu/7q1oFTCgcK9VfGaVAuhkG0N67FX
PeYZgO0mGvGcwLp1px0cJWvsnDG+AkkDzLJrqqHCzLNBvYc2HTojJXDV/6RlVFDr8SlsfTja5/Ze
4nW9FmDZ/dy7JafDRFvFolsTaT1wcoyV515uliXWg+eEhQTXw180aEDRRUJkYgHi3MORT0AV5YvJ
OaORQZ1+3uuOBy5EiaFexfq/JULnL3UTzVHHN592NP/pTe6qJnS2Kg+5bqn1jbdSPbkGIWKf4KdL
rljYb3125vy3i1SJxtGjo4FZguzFWJ7ut0hmExTM6fumuPO9a3G+TDA6qVb8ylgmXuBNRDOpU1ag
+JpQ+zRStrxVzVAuc6hixX/jLK1g3LtXUUiAnKSnqXDLISkRZVLEzh7XuZ1rL9DQh8UZ6kwLIxfG
zjvs3VnUnTv8M9bVeawiyF88zk3XV3/hccDcmWqUUpUkRv0sjMtnfZA1LQCWBrFM5oJJuxR3Vm8A
ax/OsHwT/by9/RruVzGG5Mkh72jpO/1jktZX3F5aATwXPRqrKaIPISdVL6ih5ltvfHVZLOB/bJOx
V1+pLwQ2ZFsKaWsXmH1bBz2nww9ZkcAo0iZrdOn9n2WvA4GxbBVq5RKIvUvptYWJj+ttvlw2B5Hn
14UQue0EmvxXOCrmm924U+vuqvZoc2hxFRNE6hCu6WKbnC6Qr5b3M3nKNHGEbcfyw4nHtguYRgKD
/h8ueV4O+6woRv9zpd3K6kgOjhOvCq2FlIvGkmIw9gWIgYNRumzdSYyEe/uZBJ8B8sUY6CqYtZrb
HeQ+RAJiZZqYR8PXA+BWay7pjGUAAsHzoGjQRWKflfS5znw+LoO4wRq6NstDPNK+MLK8yVNL0TNQ
QhMyBAmSailSJpJpQgKs6vbFL+FUx4bG+Xbmw6n9/6ghIv/8Um+qlnnc8liIpBVvp7aAFt3ULZKr
/hF5NuMi1RFVro9QJdUGqJcyvVr14Sx318Jb4Wo2qfu0C3zjTeIV8t8ryHonXFA+8v6gwsh0m9/8
6fXC2lelZwztdedoL9GmXloF+Y0G+fMX/5YBGC8mqsONXSDrp0+4fRuUpMiu1n5JxsFjf3fFhW41
BA6elJoPFkb2FbCF5oAWTskuGZFU/Xk57Whq8r2Z3BG2WCI0pzV3mVSMhOxPyiuWEkxnoXIrFBCw
b7CDp7zcuZmxaQ83RDbJknbF4Qzw3EieQIV6ERN3K3sRhAllGcNZwztyuvP3trekcOLHOLqocPzI
oWyTZrBS8GrgqzRVUBlD16W05gkKDkAzQxO/TwO4RiDODH/oxwz5mZVAs3syf0aqvahd221Rkafe
VR5laQT5f9X1u/HNnwQjoP9MIGIeuEt6/VColLljSClPrQiJjZqawEB9wLGG9odyyCxIf6PHT5rI
N5zIupE9swm12gM7yrG4/+AVX2xmYUp/aFeRt4G1aQQx3f9crzUT9GR3fnbkIFUKROj91+ap3njo
HgmvfmBrbcD8M92L9jgQbMpKG1AxZuCFxgk7a0N/znb++Pvl+Wd2ObbDsoVexv3/gc2jRILIzGel
+ksDJkduD9cGpM0FGwtGspqSqkujyL8C1h9rIjiNlrjPvM9KjsB/97zULF4cyNGMsmoTzcxXZdYD
SdRm03qEx2eP9qU9qoDaabrFxPj19L+84R0GsNF83LfVXc6kEuEceTo+tHTowtmAJ1kL99uQFZmf
EymRoeWLqPL3jAXs8vIkprKcvnCZL9Bt6n9Hwc9NVfeBFwrjrs7h4WvAUgz20LXQGKIQkWTqacYD
ED3XZBLzh3QKkAQbwZYJyX5zMIGX66mMEGRuk83ffSjC1X8tS6FVzHQmjfwZabyDMb178KCurkKt
yqWTBJX313woxJru07hxXLgkrkRNnkUwBk406qS5/HQU6VYfm78dpSY4ZplBRZ/SuOOBbhfKCCxa
kVUeM0nU/ANsDxYkD8Puoi/mQiy91Dfos477llFxJvxKzkJ4psnfDyYNh1QqoWMJRmxXY0fX16Bg
uZyAwevBgeofjLOE48XE6peSZRXG3P1VDcn8Rl7R6NGsvrt39RMhon2eWj51/FOQ7DLdE4rxlSV1
xJoCaHO3JBV3Rfb8cAC5lY7naiwMwRx34bO9MCWcG/UyG/omgK3mGIlB5GssnheGDwtIh//pAYh+
hpRM2UtLHJpw9NBK082LUkl9c2BjO4Fp0+moYWB9Ir8gnYlWQNTAs96LPPxCVKvPw3qvGyABDWGn
OfllWwDu7umPgVSzAAM+TBgkCid3DbLqV4yDccIGj5MknLdwhzRJ0o585U3C5j0ZbyH4CeuSatjy
z4El8djr8QbWCwJAk2CKJS7CbdxMMcu4TO66Mk0KMG3VmVwLTOwG1mJxFWf4SV8YwBrB0D1/0I60
FdB6YQNfMfYlmJsCEPQ/rJJXswOdajGYGxFEuQeoOFOemiw00SDL95Oeg5XnpqeVWgb+X57KSvAT
DiWy16aR0cO/HKY1HKmPyqg1XQuyizB5cKgPNMAeqDTlmuJpdd43JgyPLZE8JxIKANM4p5Hx21Tu
wyw6OJrTUkB7G6scsXFwsDQ/LBMZyr3sqGR7djoJ5BgtuaZiBsXMlE/rnDUCWitjGRYrjJHY1Lwc
F148x8awnZgRSi0IsTRBDwvqhT9VJcGaZB/rP360ukZxp3VDAjTQ23HnSJKUW3+62WNpVXIwO0RP
opf2VWX8R8StPo4TakQ/zjCdUuXwsY0oTT8JwXmj2mFRX7invWmrQ1nG+i7AKrLAvpdH/HCgRD20
a9UfXp7a1j4gpv/ziwTRoyITgxjRtR46tpX1Kl399gvCEU6gjjdLnDG/SMntbPdPryHCjhcvi4mK
Fh6vFzOmT4AdTj4LVJkM3SBUh7UUFmBnFY4BVk68rw5Q0osDGTPrd7ceI7+VvmAq30fZtLzaTlOF
zPs6DlmSBtUhuOy1uWK/sqpTZfoPRrTcyGXzSHOtNrI8KY7HYbnfx/FTAZ91sj4YBTdN7OQEEj1s
nuenYQXTfmRoqhw9JlqVh8E55A4Grj/Y9PUTov7NPUpzDbTXXLE4o8gYrBtYauqKvkK9gUq/r41n
PAe8aDfbdX092SwjWWhC+6voC9H3HUesK0GrL/fD8uC1ADX8HZ1GkZQJ1rPfehrGsivcLezZvv1l
b+4P5v8GJ7VIqHCGvVFmzBG9w8wsqEtPOweIVFWmyGbTshOYC5KSe0m3ikBTqBQzzHDVuTOBY5a6
otnBRlnXju+9Dzfa4kdLKAUcwxQDZLEMkF9N35iWVkpsh5bGFMoa8KYFX3DWlI00dGtkuFFhhI5b
IcUvaV42OoAZzJnfO6mxnaMWN8p6e/fg1MmwJnR46L0E522Z/BMpyo+8EvRatdFjXIe5i7MsQwCw
OEFT/BGEMVtxGUXRpK+ihuW6er8YKg+dqzH2YciaYdUN9jnTFALv7a50XFvEM4sJAeXeBqKTRue2
OrcZnlf8BVWurqn9L9z2hA8GKgrdD6RO80z50Wq71K6A8bFIPkOm4G20SzJ3H5O0uSXJycOZOn84
Ra0xxQmWHgiasQDxexikXW1filx8EHuXLAzqve4ACWRpzkCddw99g5Ed0bxYtxcdRpFcrbu/0kXM
3CM+GNK7Oj7zRUPn7ciC5dJtAfjzU+4407VdgySLYqzuRVYe20ntWOJUiSxJZjvgawjO1HvyQnoP
bR6ChrmwR/9rltY8L59CC/m6zME6untHOx2aqXfS/QzQW/buNer3rkGrT/ZxFh2aDQrrg29Duv/G
6+C+LgKDFhy96BRO2U9gi3QL+YBJbpe54Lgl6vRroWkiqUZy4/KL67w4QWKuKbINV23AJP9iTdVm
m6/XhQnNuR/gxee9gqHdTFO40al86ny+gTBJf+ghk9ZFqqjMQ93KIGWfpsjDjqURRMrfIBllPhg0
Dqi6noUQqlgrthkdds7bGdr1oqwre1rBkqBLfnZLfWi69q8vhvsLB2DQy4Avee5SGY3NyR1A9cWP
XsnKKzDZcBiz27pj/INjQtc8MkrIjqrAKO//wb+GQPqJ6ClXWGsh97XztK9GgiQ0FqACkZw330Hy
yHXD4/ePH/oQmpWevyht6D3esu/8NCZ4VlVYNHlFteNJiwhTxjKZPW6A3imbSF+PGDf8p3WNnbn7
P8or8xWYD6MJpaHDK7co0sZMiAcx7sgXtPc9RV9doE/BVOKcyFHcDHnBucFFLof/711GPwKdJx+5
lK6Guq6V1NnDmDHNcJ5398BO/wQFgZdplXUmW/GfVbn1xoLkQBWBQgFtPqraJPBit/qOamed9jyp
4N0/zMT7Wy7MCC9F4x8pHeoX1zSpWN8AtE0fh+kYc8yxO/IRapr2bw+6O+G6sttmudRDwBRugtnQ
/TGX5YBN2xeF6uW5/C8r0avynqSCa2kdLGalkHOn2WvIN3pIab+ekXvoByk4KiaHPhjBHpzUlqnT
jpi10UJ5rec024MHN2Dmf1trNrdWlZcNu81BhbvcZKidvPLMTZR6q1H8KELLPQI1zzay1eBI16re
0hChd0/tZh1I5MyEqZioHo/Jf7WnJNg3nOVOhh6eORbJ/obLXntQi6Ipp0zOQsTPJH+3+EuFvHtP
CyZTpVNsUoYz/fcI3ePrbGzirX19XUAsNRpGaCQI14rUb4vOJUHt40GskPqInYly/M25o2ConEiX
hz0D3InUycKdZjXLzs2YRN8BplZU4K0OtiB4QTYBuhZU3SYFb9wAlpprVzqbx8MeLT+eKqUw6u5t
yVJw56lo1ONdYlnP3I1V4ob44DWFZOzMNtEB5HcPolm0oBBxf0g9Z07lUytXc7MClGo6OD+aFkYy
WAo+Ts+XNxyCcN68n6QKllTz3GJpAztE+g//5kBbkJQbg4xGzh2LtXb472ruUXXm18WwIlrs4Vp4
tVlUed7ucPkH//eqdQ04YSF6EskYi3mfpS0Go2FOrSX8oEk7ERLVfQPxKK/dQB1ld/BcrFKQTb4+
a3U8jF9I3wOHva4BqmPpSMXPN4zelnPXb7BerNwlr4+mw2dPsf8ibblrCXZ2OVLLc/BSo7sKm92B
ELTv8KhCW22ANx38uv45fsLEmE5EYrDhWEZ2hslYAjqis0YYRQeaS8shhvKm/0ySzFbGDt06FL6+
yWaCnWmzCUj+Tr364j+v4Nt8IvZF/fNsle9gtrzCuB95z3LIW9LWKLRL2AM6eiGetc42iSSiDY6Z
YX4QitTFDgZjGa0dWIa2WRecVwah3EbvPvfBBbout4JqgtE8u5g6dZ2LvGbkjtv3Ak75yBE60AUA
jeBogengZNmx6wBlmPwfYV2ngC5KNAV9I/WRpK7MokVzKhDiMg5Yhw+KYpdCirbW6wcb/mmcYMI0
10BkmfQMaBGA3n3O7ptds7ajZWz8LRw/iSSQQIkpRHC8ndKZmcnG4gxUXQZUD/P3Uu9+yEjs0zJy
rQwgRYQGCIf/F3ZM7AAKzdXTxkZyg6XPQ3DtzdG9ewS3a/9kazCqJzvcjOdClYaXsOyibfkF/oYh
73CvlsF9TaZHKly7MbfFCxJ/B3XsxrtlvDXtGDRvA2ThTux8+JBylNzwlvbLm9LrwNGqvS+bbAf9
iXVcYQlz00AY+72Q581+kx6TSqqU0fdnlxOw6Uk4HGUEs3sYw9WEN7fKmH/MRc97g29toUGLUobg
ok1hY00Gf8VN0g2+89BQl8RjIOn4hmEPZ6asLIYbqrxqkfN/kmQHowrLW5ev9ssZkgxd4VD3Z0do
hoCiZjBgj97C2edUxvH0r88/3TXXYGB+sPPrF8CFVqXft4/UGZXMbjpB9FO5WbuIi+PHoRNfo/Eb
u5yqxJJCHLWjRPiJQwzI4o0JYYvOSVVhkjXUj33AqzAa5FCWyilwV2U3+Vph7TQbGWHmV+j6dKBW
/VMmVMOsSYBkUp0lsd4SuAbJMMeS/viNl9JadKlxQSwBekh1OAWeziAxIIIasgMs0MiVc2hMIhlK
XuaA+U1L67wWrBEj+B9SYUlXyVdiiX5I/yPn5Q/XYEDTLgrU6hVOfEYJzXiqTdA5EtEPSKwmwwr1
Aa3ifmwplNf2I5nCmBazEFGzKXcSC8z1dDPPKkJ6RUC7LhItwz/yThjNOC1i0CEtjcqGFTgm52h1
e3jUQ0p7KgxlgUmYSGmTaKAhuJTRXK2IfouIJAYtl+FKKrSEoRQzpTZL77jxTBwNmp1Apk/NYeme
zU95/DBMX/SN9W/929tPDg9jrAKLIpbLxYrLWnke0qKFk1xuWp/tDgSkFfw86g87gRU5E9thJ+dW
qbOFCCtL+WHLZq0lnT5mW8i16zE6FozcelP5TCWSsGCjdr6qbAYIVKOr3RSDVkRJjJJG/n3gr4pu
whxu4LBpeKEibK1nfRmJQtMuesCHtDnwwufO3hYm58ArQ+rfIFnIrkG6rGaV20/GI85ZoSKvT32O
KoexiEiSMwtEjrO0uZDhA2Cb40gejZhReSflbohWFIRXtqn3IU5MX5zn3OxZudqTHZ5U9BgXXS6K
dMEHPGr2M52TqyIKCMwo5JTcKefIMamT2gSUzCNvyzajZL782Aa0cJpm7Y09qwbxf9K2ismS5d9t
+wbRIM1TjWzqkdxkdMp9OeUJ+d7177S7/U/5LmbaRbuOJRjMU/+m3+Zl1Xq3xhk70V62k7b7B0Ys
1P7tdyWC+ZgSWSTjZ6wJBEyPtoAYelpwI65IxvxrNMwJV5pq/zDaBtXqEs7tHCkD6VKrqZziw87V
eNATwR9Q7wcAR8k1n9utrLNFektTe+NhNTugqQlVNrmV3+vwMB/Pbd3rHSyzWo7AHf7We4qZjtxC
EawUkuj+2Fa0DNMQFHa9Y9G1T9jWVwaatUoGSSwgrAhS85digtVhyQ5nph0R6/d36BooGriJl7O7
H1B6l1Dz0QF8GQHs2DgMaTSrHT91RRanoCyhAWD09tgR8b+OlfcxmLmbWOmcbLuthV0Ba+GsW/Yj
Wk9JGdIYguCSLQu4pqEDD9Er5pvVHp6i+S8mz1a5lUFOlilP19CSWJeYSoS6e2jIz/9ChH4pTw7J
D8ZeMK0VLpbJgsX62qIzEk1zAMgGzisu5B08YQchhIVSl2VR39c1QZqWlsXYZdam2bVh0FUr018Q
suD1LxzQc+1vOMwKR0RPIM5G+yXHjk/RckCYTaSPs5eURoCcxU7oJYmXIMXk9nQcKcc6hqv7qgfP
6Zhx+m/ALQcTYpVmevaa1NmIsyUwJeZN8ytMN4IEKRLEXklIGJdV6vO5LUHYWmPpFqHleO4WKJ1y
5BHwfGTJ1AxPcs4JOonaxwA6IAO/ZhOYrXhPWIH0sZtrIIyAiNWlGJKl9Qd+TNPrNKMwe6aORsfC
ydGIzipFQczGwVA2QiII0msWFnh7+HQGhxXIUwXBoXv8kmHvLQCFrx0jbDj/p2iQOdFl5eDyHby1
Jy5/wspuRn4BKeVoCMIGrkI2rIsIB9UwwaKqYimQ3pb9+SeaJF148LltLvQOJFfZBQhbbn3EkbAJ
x4ZoCcPxvXf1dkDoEA4ZET9hNWYx+D9fvXyMkRmoOlOycwMw48rpEEC3N26ThLAX8xYEMC3A23QL
H24z7FhxYCBlBo1QGifPq5k06K5ZuuxL96UaaEmURzmDgetFCF/nC+NR+k3rFUrOkLZ9Ew1P6THF
UUY3m+1oeLuT/qJmpXhNwWwAIEb/AdPq+X20tfEWR+kfMkjJdQjhU4rGCBUaVOaIzMujl4N1NsX/
HlRXEP9j6pW+nKm9Mkh8+wd6+m+kWKyU7pY1lc53lAEsoT6TSgSlixlVeKgRjou+sDtNagUt+oun
Nk506f3gqSGaRCkYIRmvd0P/nZcdG7H8Z+/dRZxf24BNVZQRyw8SpuztCLMnuxHy8/ZSAf+1fHr6
F2eF4n174KyLHxwrMf6Bz/e/RMW92z6Q32MKXOVMi4UEtSBMd37WFe1sWz8gGjm0AnN4xpmvbG+R
hTcaiJ3SCQh8GsbzK+DvykEuHz7rT+kTQoDOD3jqg/ipt/1rfWRlimKP3OUQOFU5lj3Iayx4auyM
+pYkH1unxuku1aZcaf+/VzfMNhnKwHwLZTecvXbsHXjYG+qMQEM409KvLUDRqG8oPDpUrT235Xqm
RgSYQJVB2CkpPzsebGBya9mX0J8T/JJYjIDGlebE8fvcGWxQrRRxYNORi9TSRRm+vZcO0EuwLU74
rnbhDw6UWcNbOxYgzmTaHiMWBg0sF1Cgcla6oPIoyZ6yPIT8dj3CSsVbytQa7tIrUyJcz2OrnYEa
1LrXZG5Zk3hp9/Ua79jtaFCBaigxux9jg+aDCAOksFzElkpZ6Qo7hL67AxR4757h8Ll2xGxaydLU
ulfHKPVK99e1vlNOVdBkebuemjNkS/kgRe+mp8mJxPRpVW/vsn3Q3BScgwtQHYfPMj4MY2JnpwpP
D/EEmOLgBQYBx6QxXyvcncWKYEomORFyRqoBWx+9UJ/p52C0C9f2V0i84W9Ck9ITabaOF2/mn1jX
+f9NqWPIAidMqQkzidInpoaNC+YRIDgBLyLt2NH89Y4lb3zJmbAZXPO48tqkPzBhliOZzJccjOue
ESklH78NnkUxmj/GS/RUVmR4nlhrHPlZMARaxti2pPyCPT54P4PAKI9c6N7CNqrwb6WLakyt5cIw
hdyHWoC1ug59gUz6gTSI+YSCvoAts1IL3LakTPmCxj7c3ByC57XYxMz1u00lXPVB+u211sXGlnkT
I0TK/VK4hIvC4sPferfzl0DXk/rr7VwIwu8uAymsQboN7EqqnhQjzhVBHdrrC4KnPc0MyGA6xuZw
yDgS2WC/tpKXPHo2xvqB7O/DJausXW7hH6rwLzqlSa+yxqFOc9bMpNVe9wRdSbClRJeTpR9HQvrz
qV4PPpsHiRkE3gRPO3b0AhcDWO9hDPrkiUfNHpb9RTT15klTyBe6wqh88waMzKCjav/Ri/ouJCaK
l0kgiiY2RYpu2QpvMHQwXRZKA1CGHKvlNBaOUx7zT1+4DFK28u9FF/foj06znWfPsRfjKsQ65wcg
8Dc4ufODhfxjKtOb6xSFYGSKGEChhXa/LgD+3bF9hlS6s2l4GZB23Us2N5MdYxSPhXR3TTnkSGej
+O2fNsCJDceBTSbw8dANmcUAwd7JKReo2sHUyiV5A0hIeQ0zYq96g3fbA2xfW87aNak3tVcPG6nj
FOiFz79/wBIZIlZe8jgqoK9KKDVVAaW0lJiIs2QOwGbdRblALsiEznub962i6GzYXN0wGep4GzRb
H90XOHNmoNDjN2/vnnY9tOwIzFi3C/+CZhF1Qyc/HouDHqPbNVhPqF+4n/ddQj2R/rzvTVOuFA3C
EJqiEbnpDO4eE6pQ9MRoJqPYEGQiNKceTYBftvZLVLGry4Gm4Iubgr5KYW41IsPLuy+mw5WKUws/
ZSHP9KOGejDRF4MBv9ycYE20UodXiC9wVzPI5KYZPsgl++kiFysF5kt6aY6xodQMHFHtnApXipDI
kySuXCa+/5JvZWNhhN9WaVVi64U9e/Ciulo+zg9Sv9HUSBVcTffxJDpWSC0rLV3rBHBaq3Fh1DhF
tqV1UIUM3yDzQXU4jSxMIIsUJ/7cxF4d+DJyJ7SqehIxWkwxNUf0RWFKO+th8+oG5RLkhF14iiDD
s0Igc75cD14S7lOG1w4qvXGSbpXpzBE7zGDDKBDOBMSPnTs8W9N+XWIifH+4gblwcXkrPJooJ/Yt
0Cpo0/NrPDG8KlRSU7Ju3h1w1J68C2OeDM6z9fSyCQwJLxFx+3GQ8LGoOpqZBd5fqq8SKVZPkRgr
/2yuD8z11JiqDDm8Gq7SoXPMaGSnr6YFZuVv9u/G8dGix1ltDPnlqkISPBQWoCHechoUQhDmWoCV
OQACY1e5LvQVL9t61JZXOfXxrDEfdTJwtcjhFywwK/WGqoExia9PEKtZt4KKtbMy+NgNS35G0gsv
RU8fEoYMOCcm/kXjM0MGLETeUq4H6uoF8XYwooeZKqTqdMnFfF7ovB54QOMSKSqpg2LYkIXdV3IP
QjNDAuQH0rpVOrP6qEXBQcYIfNPBXIlBdm8t0OZHdn3INevUwS0Fgkdv7Np+F3hT9zkPNN2p3O3D
CqmspNCmblvFYRCR7UMly4SFYkugANglk98gwJ35ArXz1yVlFccTv1v1L1IKLFlnK27QmxBUXfHS
RbYmMy9HgO8Y0on01r4Y4tVlfDxhOm9kNPet3GuYBME5VqTC2Kuxo8g79AxzqFMMnpgBvBYLdZoo
3xnOAfNGDnYPIen8erXcUsLjyLfoGK+dqWAGG6bg6cgYhDfzNXp+paeNuGbhbIYhWNrGfOAylmP8
tJNUUj4BdnCPJ3OEmuuZobdU75hby3STKWxFedOfrqHIlB9xJEb7WS4ul/zAtWJzPoZ4zWjCL5Cf
HFRextVKGv0nFWDw6Tj2mRw/LcH563qx15zoz5K6Bt6N7LbBEOcjjSm6Y5jnym1aLG66VCVmdJNe
dZ9T1cnGd9UOsHN5cs79kph92MYpUKQ0ub4xNVlVqdNmlk3HDlli+8oQK3Y/Hp3BK9R83qS0mEbc
Rqyf+97ZW9iNzIEEltNGliQgTkrKrQ2ghhK4BlQOObzWs4BjRmXPtYc7QQuau4K64hbxindyZfTM
SAwOb6c+mhryjOAMjaivxu49MkA98EP/LbFo6HZAtxJwGBfMsvqWFwQBnwfCcklKWpUufc6f5Ohw
Ghc1Quy0z8lyOT6kTYZ7pE61D1ozW09H5rGsqXkfNVf3YLxjtvlXlQKJN3M3x/fXSOUYyq5q1wdp
ifiF6gRahaFbY4pCI+9Z0fSucVpkuNKPphJM4ez25JItxfKcV7S9r/8Jnflc7cZOjeblFLcOxsjS
YxbPt0w+0zb7hiN9XgdzGB/SvW5rkm/z1BDpgr0xt64e31cqF9M+vjJl3BGqvX/Vh6isnYLNh27e
xpuPKWjM63dOOVSrxx3m6IKSrCjJ1M2JJ9yelreQNmXL6IfxEaDUSuc5S+iMPbivOzt6cxdVTOAj
nTiACtJecCrr7IpW8L9AxOwqPcYPAB3sNW/mrHbzHj/+UY402KreO3RGlFgCYEXQXbv8CsMhepuQ
nj3/MAgBro/IejR7DBO1eomJBR9i0m7WEJTEQ0DK0a6Vy+KfidE5JVGLiXUSuET/1BXB27ttEUez
bTwNqwUuw2Kx1nAMdFNH3XtqnKXLMBKm9xQ891N43vzQ8pFHWB/CflEeikwBoX1+FYg2u4lQJqG5
4TxNTwhOMkF3jeHJ80QAcncjVECBoX7EbO/bNgpA1P8QoHZOe8cAmMu6L7J93gISdz1dpjw9PBNQ
x4f6nzhsjJpYuqRJ70Ws1zcr/swo5JIhty4VsNSKf6HRRsopJjJSHgUI6wtzXuz2A2g69ORgEVIn
j04/6KzYpigfdMaC1WJY+dpJJuKdap9fDdTvPG3Ofb8l3PthU1rESkuF/1iLmRR7PEMnl6Thq7Q2
UlMaFLhpvQMddhKIMt2kUJN9dapU0Nj39e44XLetfE1mrVGm7Nccji86lSqybtnDkgyPpU7s6YVP
/N6RH8P+ke5T89z8VwSpu9ST+17U+AY3mKEY9MP7HXxvHCheEkKhpv9OjEzbthj0iyVcPWNmfcsg
qQSY3pRGMCkeDBT5T7KBcKofWOnYHVWsAyfZZahvwJF3YJUk1or1Jm4cqZuXNdLEAkLHUmAicaRH
8Sk8J3BuwZJudU0TQbzOK1UxdGouXgx4XMGkrzQD0PvLUV8r52iYRLRAhY7i1BgEGuTkzKnjIqlZ
Q0FP+Isv1kaiDZ5XKIc0/1sX/akPcxlAElAjfF/1fBPU4a0MhLhvZ/EDDq1Rci8wY/jYg7HRGT1I
twdheMnz0mso4hx50+slVYuluOlCkc9vJ1RKermkzVLouj7Cjbp0urgD+drfhIpULvGkZ7kPgi5E
7TNWIgm8WfJTapTcXBaHaF4inggQQMaggR4cHWBE5fYJ7i3Eaxud7o9A1HLh9uktVfhWH61pg0r9
Z3eVlEY15IjzDhvs6QEB5KBkYPEs7wFcITeW8tEZB163czF/kh3VAz2dVxMQxEAJq/dwYFmJmYXe
jD6p0eNprTX3YZ1K00k+9Ie2UKkbIok0dzYh6w64Xh+JNebiJJGr7zw8fGEV3r1A/Hp0RKXtxwsM
H0OVVBRxdDFmK3D6GlMJ3zWsWX84mTxnIL1EsiiFTOXtFjYrjXpmqLgxA804MH8gowFSY3/bmDR9
6RGS9Ms2P5wGe1x9Qe4/32ggV1NENkHvxUjSJ/zOrIn4VAnNpWk5rOiykohzt2mmI5TcblKWUi7M
aSiPUarAKRpVbDcDvv42lIg1X0kmq1xcJ005aNCNRm1kfqKaoZI8silxT3IkBWd24ll4Hv8Kg2xw
VEYGU2VAKfXhpZe7puIvLqgu93p95oUYrbdjTOZWWloJQ/hjvrpEQ91PtXavaaxxcd/k06XGFyZs
+nXZlsD2W8r/XZGc3opdBCt+xkxPUKRKSozVM3SqkU7SMS8hO166orCA3tv3hAqEqA0iuh/LI9iM
n6+GtKddxZFnnNCsXu9gfEN7JtqkzRvcfCdOjFuPq+au2ohzAMm9mAWjA0oEDfDPrXDnH+EAIZsY
nV3B7dEK6YbFW16JfVgM9LK3J2N9/2c4gItHynnYk5omUZ8nqmdg2jDPLoWUjJeS6+lilJukZpG3
spTPJ8kJbqPhqdaf40jZqfdqbhmRfnZLtrNLvK2Z3pMnYSJGXahp9q22M6mhdhcSnpFzyVHWHi3K
VeUOobpD/WrKymjqFWSLIOdnPYcc8tXS4Lf6eaydtLSXo371SfowuZ507aZVeNczlhF91fqoiJoL
jjH5cCNuqTipXu4nrLyhIM/cn8vYOM9n+T2iAtGuSSkRe8IhVE5nsYBu1a+8ms6R7ufvj14BTtkV
hzQCUCapGHBYCNRW9vuMCj1VBTgperPgfr+7ggPdTQ9SQy3rbuoFh2GgNyR2QojlV1QJbCbc8nUq
aTto8GxVqACV5EEf0cS1Q5LZsnonWkAjodTeKS4jgJWWWf01ugtdpAnwq4x+3Uc9PszoMJIhFInb
Qxldw8DIONOMj9xGHL3l/GXaFyKV2yRAdsHICe5899jTMWoZoZutHLuY1DP1VUYp8goyLl+lJAtH
JFI82uPwTcfGGuew/utPRtqKf9xrvosEAs6ORWVmso5f3sALa3jW7jQf6z38H69DbDH0YKm/Sbyn
DdUEMeLSVgQ80Q/YjxW5grS74ysPNh/kdV+HoxOT23a8V3MJUJ3n8CSvJbVD0YpX2BmbNTr784Yc
AUboAwyUkHnjzFpADj1n8nB05XZTqXr1DFVurXAPLPoZ9/+3djZCU3MwuBWp0H1U/jU/7v2Y3Jid
OInnbjyhVvhxhkfq/Kb7jTa2C229oKE9GfE4ibyfqe0V9A3T9ADzDGJs5YpPmbji6NXFYURwX2ML
EGEN35LEHZ5YMXgNrzF0aUc5dPV4XlJdSafkN+bjTNNTqHzOZ4wf9CfCpFKNqw0fLjGckrQ8CWjz
jtIm91hR+CE0eUxObCUf/suX9OcV62EwaTGXxuil8kjewDyLbo6z+cVBKlu+1ZedZpeukWFmr5mg
cEsCwwIAQ/ptOaFj9xkp5TD6kgIuMYO9czpFw7vJ/QSD1AY/0vQRKnW1//BWti8fEKuiAKedT8bI
3uPGGuGzBS8lLxwGssBmDlIAJoY79QGaE+WDQo/V4UzA9I+ZN7EKHZDAlLbnkHjUjBf+W3gapWGJ
tLgvzrSl53pSzBC6do1RnfKxLz2M3wyPnHAclt4iDGC+xhuMQ1S6Kb9UDwC5TpyWRbxA6Pc23j1D
aWnFy5NQPLsvJhNt1/JHDBmvHAmPjP2OuJldXJqMOCCmoPvPH/aySJYW74RWcafbJIgQVvfjv72X
cbwngzcLo/KmyzAl1OajHsLPLQbwafVHN+iqkEzIAMy9L71go5Mwwhh+M6cNATV4fmiCXUdIAZu0
smGWL5ItGCIDDQ0oepRcuYX+jPDRYB199dy8wHmLto7Thm/3/cCGIVbQFjwJcCNsE3OflQPxrv7L
VLXOpxqUTnitW/MMj2hlJMR3h/VCc/WfQRYgj9N9JhL7YZq3UMU0UFTSRvYanlz2m7CkG5fmaWhl
B+cdCg1dIpoEHbV7U99s7bP34tR8Dv5vpZAWzaqvY+9NTepDHp/9HBIEWfEbcDwfEJ23+1AnpYyq
suWvgZcYFZOcV+9tBUNMmgjaMUh87engvN4sqzc1hRZXwCWvAqS4IEsm1klIFMXwn4xPgigwwrig
5bb+WtjMwX2FCB91Yt6xm55Fah6qDSOeC9RhxlgBUoMRfxJMZ30Lp/vse/Bs5+o5WQ/3D9j+KrJZ
GZzbQ9FWLKPpQH8EqMPT6/MSaAuY+Aqg4vUojLoC1IKRbkzh6V4+J2+UwJY00bquH5zUI/Qpi8M3
rqBIuFwoG9jFClSdt6tP8mUL0QweUrfySVepgmJxBJB6u1NzaeEddsUIgDconG1f0GP0ntRD0AZ/
jTd4H7erBlJrb6/qt8uBbPTfQZemIZneC8KKWXHT+K9QAyfdrLK9OXiBpuyM5xwmXiWpsqIyOgD0
BgFeW8Ye5Ku+bTlU5NnFLI6DkTx/yB8nslBoRe+9ZyMuvmKrZDmFGK94Er2ekp85hx/5Kr9610NZ
lcAn5PATw/q8IC/4jPPVbBpTVWkLzUmHuiAvfmHBybIozpLFkjaj4cOPRGzsxuJ/M7eM62QigQsd
KVaFHyTTibbfM4UmENvRzQ9VE4UUj7LJfKYe3A+XZw61suYd+QEx4GqveBSkLgrEeNigbzzqm2JU
3Yl6HPoAAxcDeZ/jFV0YBgTqn0+fYbR+1lUGhMkY+d0XM9C6GiQTSMuqB8IZaeGSXr9oIK0y8BPV
TIX/IhZVxh7X9YcvU7roiWLB6x0vg9pMuPHKXY6XEQVDy/8mrJbXLSHwbLBVSF5W44OQtRgAjqCI
ck/GpxGeChvP5XU/Grx/8fXFJHC7V38KK/5ZJb7ByNCptZ4uc/SohfUg1llfKWQdvRIf+shH2Iow
HotsL4nywvznJyrEhkVPQ6E7KfF150DHpK/kZH0AMWX8PGX4t2+DLeL8A/+G5EzRs0cfyo/UMI5K
4yYh5XK+pxRqVhr+B6gb5ZtnMq/WQFVp5G53aQQ48mUtxIFDFHmbYlPY8Yc6ICEvkdVSwWKiRlkc
f48SjD74V64guU6qWzCJH9ImSBWWxH7pvET4i+ZD4gTWgnTwBrs0y3+h0Mqatmr0fmr6GKnFOGf/
Uy+uAbMUcV14ieuTZWYZR0bD2feWfWA94PYBclSGmPU8qcI1uoTgLcSea92CnK2hvPgw2O7vMA4V
Dj8HHayzvkSivOlhn6WwG0zdqgKRznjv84ApsI/b6aRpIBoy4pX2fSFcn4rbqhGDpyVqMTdQkYYo
usDWoBpodXYHPgCApfzLHfZUkG4vhKZtZAzlnnt337f3svrccHWAAB+rp7XEeHQcI56Gq+cecJmy
Uc3H6JXTs3W2h9kLCVRBVjDJ+cJwFzKDr7YN/4vHngdLOHad+NlpHzf8FDl+lzwIC6jgJM/lZ16v
S87fBb3o9i1iAOVUCntzGMAqail4eLNfwXveqGkEZ0TNzB7Xyqn11nrhaWqCBRSizY0FUF8Vdwoq
psBWyT9FBGcEyzxw+ijtNmShfmV9e384giBX0knfpVyaWlR/ES0+ntmTbuivFKafNcashE1PxF8w
MAVDfn4tmnk2KDefWeWTg2c7KLNMsHtaqHy+dUHx/Bvxpsn4GEvqaOCcjBM6X5I7q3rV8vlqOA8J
Jh3NC6uuQFamrdHP32UxZS1DgiAd4uCbP8xDt2QCvmIbwBAZN+pyM/7tsFaFsfUz5LvLU1paJpHV
ldWvi4IiWXKt7GVSBBlCX9C7lKjqpFdlXsjOOHPiqCtBs/x9AQsr55TGJnYQ5P7lseIs2RQ+1/gE
fLeV7ajAJ61nArm4eWG45+c6Ia93pmFB30MIXlQ8KBHQ5fiLhfLqjsZpU+ZTIFtiGgInkXp6gBPw
7Pqn26cwLRccOIF6nav9waQ6ptZpPZZwV9jQ2d0bRgVd24hfxgvghxJ8Qz1C4xpxWe6fDbAnU1Z5
b+GKgTvmOrxtOkwMIi7mQSTv+77u/R/HXbIdM6zoI+HsKTvj9uYJDIBBjsWE6LXFuM87fpek6kYP
6GgFEESN+yJqD+l5btCU411Hdh0CABR4VzOvrxK/RGu4JLLg6m9nuv7pjBpdvfCPUhpv8LQvIVgx
FZUm92nJcCJKxIwu8VXaz2imyw+HrO43GDLo3txswWpgyNFgdgy3N3IOOQa4oJY+NcIw8+5DnlvK
n5Bj0wvhYFwUEgMdKnKk7oPUrbxxFguiKKEh8mkpH87iB9eJmdiJFFLEB14iFb+Nod36rzBOn5Cq
PHawKCBS2xOUo8olxGAYCNzW+ydqde2osDoRCyaFbk24uoT8oLRdAb69G6VFogxnDpxxMeFZF5a7
aV9a04aQ4xbYVCFn2t+VVfOjXR+NYZB1ibteZP8jM73f5l5jqn3gQOqVhD0/SGelKLKsB1E5NqZu
54AWS2gCfGr66BLAf2IFybrNYDapu3Ilo7R9Ny1VaKPeqPcLhpls8lJeqvTFbJwLPP32rPj8ByJC
xYgNczN/i6pO3NxT1FTSIG165NYoZsNbjrG/5Tt8CFgemEzflRVlrTlF0gwcEd/fm74et+9rHFm0
2LHyeEU29rm7xh1KWO9fc1894Be8WX4Wby1Sjb7jgIJiuSDpWXO42CmtApqQomNZW/Cb5g1tz4dO
z1xFsDoMjBwxUTHasnKSHsbmHijXVlmzfE6VBz7C7hh7svvuph6R8tPD0bLJYmFCZERqJWNLM8dM
hkL7v7tQs1ePBRYcxMoEpbSqRr1atlLEMQmwMyj6MplR1tqjJwZD2FBLouA3J+b/sZTzmvLLdpP6
LUycAegu5CnrOqZOurQIbs2ts+cH+bMKDmbLeRCVJDn3Pe57kagzA71Gev5mDz7oC1BnzFPaIJZy
UCVUSFY4ImC2i7Ajs/B9vBdDN7xPkRWCPmKnzI1MpIPBEe9Qa4R1PehNLmrKuJZDaL5SaYVy4FUh
DRlZkSKjP8BxXu8pq09dy7wPFXftAOQwIc9JqjUBGmPoPUpvg+2GtRVqtMS+ku9pss5kpRjZxOXl
QSfu0RoV7TSeW5yv444o5zoC01wB/7rT4MdnOQtTH/WihZro31UyuG2ZlIPdUePSTDAIf+q5kOiX
IjxxU0GaU188XP0ydZPX7gX6agjeXhcXY9BLlapkuI7Iex8wtdhZQU9D67hW0N3G8Eytz+76KBMX
PJz48HsVErRoAhVbedZWTmRfldu9aTmLJfExxOWOYKQq1v/9jGKcbqOJdqiUXVkpaUqvHlWrCUqY
KAsFSp7CiIGKrAb8twYhzNyVBBHC07niX7Fxw4o45Kk8dOEd0Gl0Hk1lV0LnT5puzrQ+vb88RU7p
f5Pd2nfxvGvGmqfgBKW2tyToW1DzjdzBB+tHmoo8wBe1dpgamC+eJKCf0S+hxdbnALmSBOWc7PBJ
i01h/X0ga9pNxwgEcmE3ArjhcM7+B1T2NKnjDHivRkYE/MKobmBAxtWHYE5sY60JC4I/PtFYkATT
l4FvMr6QzveIPmSGrwTlUy6e4xtd0MyuHKMnT3Bm+pBeyH3fLzGfbzOfTglOmr6oSgCO/w21zLoX
sF4+n+spjr8XAfZ0sED9hzmbivbgxszSC0mq1db6kiHSmrIu8QtW2GLF0M1kUNFyltTlYk4ktygi
XVgn/e/t/7Us0wom09Xlv2M/nO/WopVAMfQc05OuASVMe+WdsmU9cgZNblDu5MkiXLWdQvdS0j/Y
9AycEbgYA9qjG7UOnlZI3ZPLvGLMbBzDaiOQVB1gpOFiSAuSwhDLaGLhAKXFsCcPS3WH5Pag1Y0k
Pn75BIcaKmjkXRbjfNYexn0s6f0UCuyyDTFmzAXrfZ79AVrJ2IgtFBWblevs3P7JSfhR6K84zGAc
TimBZxLq0WRvsjOXDQtHyDqXKdzUMhTc7c+8dlLiEQ0bJ/0tZzzjHh2m5M1Wm7ova7t9TjKcdIew
RTocC1s4tgP1RiX/ToHDOOlifmB2mJquJHYSrrIDF325Ps7tq0An2u+Ys95/Ep4bTwIG7PsJYjG4
680cEx7Rml0Sjf9mkDV4ANNszofFcT6IeRCzbeF/siuHUBzVid2kNTsbWC/LR83nfz0YKv67+aBY
VUvMi2ufR5fo10JWMR1FbDLsGOFy9hMijRxkONUvjGjaiPeEP1++Sma2izfOn+3w2RfNX+ukBOdu
xkTOhwU9k27RzKCKihtUzg6cbWWi0D1wmD0YMBbrWTkPX++AMrAk2UG3nlKlKWwZwGiQGmDBVaEv
Bxii/U4RkcjaKUHYZB4Hjaqsgn3FhEcVXIqJ46Zp/VJuWgHaL66vw0FRFJvUium3UgyunuWnL2qX
OsFmi1unPdA4G3vx+q/KpX9Edk4a1Vv5ccA2ecNMEq5YjLC2EgT8SHh8Z5FQMFXv2UIYnOxcrohc
tD1u2Jtew12neCt/DwYqLXaBlrQiKbbFNTLFTKRxfaFACorKCi0daSEm2z81kkFrO2LK76R54Smg
hHVlFv4ntaqatEC6ba8KqHmgCjZLoBECt747aS3C5l+FZw34FTRmssvdp+Fcl3x4AWC6b9FxM/LV
KWfEwcsC73OF1vGWooddL5+J+ZUJKFZ0VFKLHKHZaxAejreksBgInSRSjLlcpJADUUXLvYXiooWj
kyiLRY+Ly/ASngBAp0ol40vm3Efd0wRdmiEajV0+SOeFDBL2NBkv0ISJUAUDfhDcUX1gf+2UcWR0
MoOm/heFEm0m4BFz3cA2nacy1MKSuALxVHC+6IBzSzGPARNYNn8fxjkJwJHJBcfjg8iHYD1gmP9W
ZKXHGo5uKkUwGekrmrtz26YzF8iidyWeWyJepg1oPko1ZK2vFNumzkg6dmD/7NMKhTdgV+rNDQM8
5ZjTJen3Er/U48dhqvYGe6r06zt5GEjXHrpdIBokTxgH0ZHU+8V2mWXGemHqeh7cHAMyr2vd5G+d
0eYSbGHRKksZ1WiP+Z9FMxSydVpmvl3w2Um4JMAUDyIy4TZnOnjZ+Yo7TJmLWKmlhY8AltkMij9J
JYvlevddQ0R79VFDF9z43hBV4luSjdQDFM/7UkMehIK4zbKdnVZzSpxhiX9ixf7xPTTBpR9Zt1Fi
FaQsatW0iLS9M+X5J93K5oxEimJoMd54egQZe0yCvKMwYd20ZFI0JK4Kuztr/TZC+swRaZsEMkG8
7Hmvk2O7uosWnP2Ml8OJHJbSQTuZnOK/SeMvuAYS0ppuJRIFh1sigEWvGtuK4kDhv1IyHoMcxIZA
YTeefrNGd8RAyC/uOOUdtZEwnz7VtoA7T6gLdetb2wK+ARa8eQyGEVQ87Ddhg8XKfJhW7vplBhwX
tpHdI0N7ok8supH5LAt1COKr1c/mgIq2a0+qEeLi3HHt/NzRROvdLtPOmELt2tNWUcy6FaZ6PcHz
dBu3jhNLxv3Pk1c6jwJmD6fc9y7vIoBh0FP9lopmfhXzSL2TeEe23yhFMyilv+aJozGGIKL/8pBH
uTpXWOGSlEtOTghZfTgteL20hQ2QuGLim4+4czjkogNr/3zE1McHF1bwVd/oF/DZ+3UVsipoJUgr
QWvJOidFNAggfQpgG3FaM6T9nNSInfkKN7QCo7uv2RfvDjdNNqkePBoDW+ZIL8j+pbOfH6Pjwquf
mpJmmSe824iK+jKuffyIWuJCBSDF22FbNMVHraupTzJZrmPwYZqtu82ywfoxUdNGjJdCCEnLLIXD
fOlD05cN67FWuI+LVNF0AXp6rCaQWctvZErqFuMJWyhGXzdjlugwidLjae5S0rAF8uZdJm39ZOpw
6WFK/dfwPYa/hvjXJEaGwnVx2y4RohE0iE6i+tEpEeI9p0H5Sh2e3H5zvkEA42e4RlgVrK9FQHT7
5jEA6/SQWoLyCAP/Ua00UKIHHdMwQ0FqFAneA8udx9RCOft/yPp+mQFH+/vrOSDSETvrYrj5LwvP
ISlBSpmkpqMg1Caay0mYi3Kra9c3NZ0i0aPWd5MRQmP5ee3txhXvGjjhTIUKLhECVcSW82kLplKK
OtjT49erOq1spjUzG6eVwo/qJ5palYoiA/MOkcObyI4C+LafFFZCMVjib7HFZvjZrc4Xgq7xnBHk
STgXla/skZqpaGxHpTe14FLcf6Qy6iqKLdgZHiEV0m2TBR1nLszNETHgCXZoZhswd+Tp988vSSWR
WqVO7hszo3AnYuoezhv02qJq3u+XDliZytw3PRHbxFbnOVVqqTf7g0uXw3iM9IKTqrQeyJTnSrkQ
K3qA/xqfwQkAimdi3nWFBrKABhBVX3p78kh8rSl23VFwCCYicRKBsxdjLxAvi5QHJI/1uW+R+zrQ
o+Lol1XGlJ4OaiIwmlWyRt3pm13DqHgWAYSbSZ351o3OwrkDwwkfrvwLBdYu4pYLk0QfCk08nI+G
c/DBSXm0cH3Ld/WToSAkc6jrbyu7Nmo5jK+nIoSvcQRfy2EvSvN3tiGlBDjxlGbkljqffpaBlx2q
T1Q+G9OIBA/A0/wtNPCUtZkZKe76tNjugyTahomqfM1StIrsbikf37YQU0zL6Pfy/8Ls/5gsASXj
v3v6lEmraITIE20kYd2VPPiq27dsjazPibISnsnVmXSBmUyw/UpmGCMpP9qMCExgl9SLCRBBlmNO
HkEGEFq/Q/BsM25oe2Tg+6lb205M3gIkZqYfoGd4wLPspfB7Mp+avMfPHUmt70CPD94riU6fI/Zr
+3lro11Yua26YdDMnN3WA+mCtkCEqk5WoUL7c6nXDh849sNcUTvBc86sxdIvmGxpyyccOEEEgGr1
x+JJ10w/OVklcjfeQwvGxIKnNN2HBicLrnbvGNWXGRezQrpZf/zJl3HIR1npqs6Mxm5sEfm4x9eF
22IXEvGq9xQTjn5e8yR0aBu3LPQtAn7QnDqbZibk6PYAQSvcPM9JVO7qAw43Myv/lqp/r8WUPLWn
DLiYOZpjMRK8gDDXzkX3vCZwCT24pvqi0kpaNem9Zm8+v8LadWzSUNC5+JxOZ5K/BLcZGnL7F62p
n7hI4rB/VJ9Rd6KoZdQ4kkNQowC1HGorFPFwY4pMJTsCQY96688BixxDJfByr/jEbYF/wvmwaZ73
YEkQXqd8I1VSW7O5m4OO9Zump3uuwk0WB5yeFbqW7x1ReeZaFrLSXdVMm2CXYkGKE/12JlKwjLcO
UCflj+fx1b2mB0/KqEfUMOZjYHXikYF+ghP6pMIp2ePlAO00OH6uynMsgLSWiv6EJ2jar0c447RD
+OnXxD8x51N/fN/atS8N4pDpMuX0p0xGGmoJhDcrQ8dGTtzYncMyk79sHWlpzMOnolWZ+HxSPK2Q
iobSTcZwZgbbsQ7zBesebyK2OT28zWObqOCqS3Lms8X5FZci+OtLI+TQa5USrtrFzc0sVrpgLskH
D03SnIRf5WY8q74pPZ65FGrzSYL256Iedao1dUUokqxkvD6ES56MITkzisUCEmnsR+O+qesWiYLJ
FUyJzv0nN7iZAx6zq8DYqsn2HJuyi/t5Jq2bGHXXh7p+hjMkecKfu9zVY8VXQJuCLe3iogjEuSVS
jIm9YlodTYxMXodJ/CJF4SEt5tkotrYx0A+qLa/bGvxjJ2aTfrYBYwvDV+D3csQzwFzQizbP3suY
dvZ9GS41AmoDiWKiG3EX8wv86pUXI9Mzp09X4OxaGHV2ZxLvpD//VwN5WxvB+owVYV1+q2JCV41k
QdfmwHj4SKL5rf1LXqbvNgU6fa10pqNG5jisJH+ZAfqqYf04yLkf67VtyVr8xWcFIxiYWkyhUdc4
Oy0WjXbz3CN3AAPhdSvRLNzhXdiRk9ATs23EP/GUryL1b2RAt/8+irfu9tQMWAsBxnosScfRX8Bp
leWF1+s8O6d3HCdm87+p0yVayTVr2pLos2X2nKr0cXV4JOnU+Le8yT/VxV7qtHEWFaqw5HZLmPGr
bH6N6TGIqER0l2umvN+tiZo3pxBxnQbJEk7Vyqbh3IjV9UTn79PmfPV68cUB+MQ15mmKv9M/x0XA
ZLRWeYj4zByLLToGDW+DgXBi2yS2QCvk4l5p0dKTVWKtUnZsMLZCBvMR/r4MmKTbJLs1KPGeWyfV
IS3k5ezsaDbSrs/7PVoojKKF4yA/F7i42trYnCoH7Yq+ZL3OEHpZCpKg4gJEP1mOvVhnA3+yd3Ng
SG0h+NKywxWVHkYlbYAryUmEpWBUmot6snzgWjUmpr3cwk7sHypoj3hvxuEoQfIgFI+90wGT+cLs
/yClfL0nVRQh9oYy50FuHFxmwM3inAvlXb9Z553eddyGNo8QQmtixMFGnPNofrKOqNwek/jzV0Zv
HWg1ML32kFjxBF5wNE9/6AoYBx7hhc8S5AgIf9O/g3FehBTToIX97/PBLkvt0IjEBfOedVaqnr/s
mIMw1Y4Pnb9tmb3k6Xv1zPd1mPHAKiipV4fB32koz1306IiGrvQvK94jRrj8zdFgi75lMtB+OGi2
hEIhO+UE80Wajz738qxgSYtm5JRYtrfNYIKp92q6xkb0uuLLyuFfLeNgFCFol7x7KMnLYRGNvCoI
8nrg4zJEJq09nbhBSX7zVOqADShuecjJ3y4rjWWj2X+r4hKNgMOR1aDoc9ZtQg84VHLeWgVMI2TK
uxiLv9iqy4+mbso9qBSMsujOKhnxHdBkHHrPrWXUTxq9dDWVGvEkz9kbzJ4Q3U0nQpDCf5i142pz
BZ5LAbxvpeP3fVJPifsSWr0bcL11FPU/FpdnhqXEWSuxCp4FAU1PWaPgttpItV/bF/vFForIT/ou
MmK47+HKzHAnhex+ZFCrdgz4h1MtfFDn+NVid3J18bNdbdKLAq8xnS8RIpa2Dw9YW25JJN+L/hnY
eFICdrB6VcFp6AfP2KwOf0w2hI7gdegYCR9hscMWapbRa/qQbkGBfopxsjcAKvc0WR9na7bAdtQ0
06Os6GLkGTnmRSMyR4SF5aC6GBGTlMKvw9eTkDyky7scJgyjA0d6jLVglBzPLiPPPIf1wjrVjD32
LxJpUFl1eQuh4PkJ8gLDFdqFtXaaBVZNvB6jwNjOoSI6tdZSqn3ELugbSz9y1x8xNNTIKlYc47DT
TgJtXAcGm1RwON70TI6cVUBn+5XS3lm3T/Oqn9iQZsJtfaijQVTcUKUUxs8DM+g+MNZ4QMUsSi/L
jg5hQ27fJbN1hKkNaRMr9OEnKDuLdBbXgg+yVvUJXYfhnwK8HBwcPhY71Z044DvodcgJFbydpj1f
cPXL5EwFso4xSwF81EdeZTUl8wnGCT2GylHNGjY6GRhNaHEx/uQAWwfyAZfVfJFqZp4pcCZHnj2+
MZfTdl9PtOcY/Q5XB4kyVtEt0tuFAMyM/8zAZCUsXtAHH1AsDTyRf9gXs4tLDn207ZNuS2VDYDC7
dueqayn4T0ARA+YhNUMfeG8k2y3UZIRDYF12TZb7IVXG2GCp86Ztmy5eX5O9yDJj28A96WAHvIfc
TvN+FwAB/MGYxsIRPJRuyxk2ff2Nrbx3hz4FKa820gpej1QH+a0nNWSqjy5cnDp46716Oygki+lL
JSdi3U11uVIb/U7ozYkhpt7Nk3adVaQOUoFeIJ7zjfWM7tfJ7Obi5fU6LnaYqZRceOP0MoPywQnm
VD4PSjyRq+b1lgASTuvRh1yg/hiotU4HfwsGI9dUrgw+IXdcOE6HMyp41MgXFvV5C3wvs6oU52vd
omIcBNEEHUJj7ZqIkiQY9YASjqboQxa82ETAuGCpVxFd4/zxeugXgnsf58oAuxvr7VLHW4c1jj2/
KIoB0PzKBZaSjhadQ9GGGlk7CrL9vWPywqTucABa3IRKIWmkkRb/u9x1sKkCxH3/iCfvXUqKTygK
Am/YAtFdmK4Qs9aSJNcuSGZI2S6My8fO54GRTpDUKQn1Gy66e1xy6val8YGY1CBfIFPEdCvksCgL
qPPu4JHc08ZB1uVDltpxwUQjYGtDCzlcukrASUxvZKWVpaWIlkeLqxE/O+GyBqec9YboDqXkSY+8
M5neZ+keBFc79Eo4t7BN2BnmIBT55/i+TC0uDord9K27es2Aai4om85xcXcXi6zlEJsLVVrkzenw
4tRKqI/n2arNYFrSx/+QBbUgdAmly63TziDQQddTBpsYmQMBFvRITWyQxSij6j7cGpfhewRQDt2Y
6Dtf23X4bvACvAvtHCHf6QTEIpl+1nB/KD4q1cY4Hcwv3i8ubigC+3PKJ6wo1B47RO723XHwtqDP
QCY1EBg4+MgMse6jbBNmjztYLB71zSxuUQ9n1Qg9NWmySAkLBu5+FKFWGqfIX2fIYcmvqqfmOBLy
2Vx2ak8q65s7Fd7MCZemVmY6IfFPQV7rspnkyyLIZKU8poSfT1WegDxkVwxn3RM+azYOhqq2Zjzj
cqBbWef17+xUs+BIH3ggrUCGKxn303wi3i3bSuQHYucNUqAtqX36AKOGjuxR79oX3p/Tvn3ZZ1WO
QuJ6GogBVCzuZq9dpJ3QN8fQWE/dbiOwWy0BT4+053QquJqyoi9lTvCv4YSLUBRQN9dtz1R1Wpwe
j2Cx+6oigXSP9GXi8W9kmyFQywLnykASi0x5/MPauV7Jit36QefYLgqhsRrWHqxS/YileytjT9NL
I+pZV5Zwd7xLu04GyGr0lZGM6yYaWn87xeez4ajv62VlgBaKXagBHl/kBNmS0bIMf3w/QRQm9t7r
mfJ9hsTWN+i08h7rysZ7ImDbB9VdBlOvEUrpTz17i6+Yjbqxy1Cl3jPKB7YFOf6sKXbqpQxyvC5E
4lmJYAGTSuVJiPWA/Dnvyc6kd9msCCRBkTfjJbi77PnKAU+TeL2GAQnpNvhfsFB+MGifyqFJgUu2
gadeUIA19Mk+32oRD/NK40SyGayLlXi4clo803fc826iai5jz3NwQEfQsYv8uBjnekVOyGXjcqj8
vnZd82D+edYu1r4iWDZ50/TYkUxAXQrEtPmCpE5ho58naAq9pFVaeMjtKsC8ZS+9jrFNbHz24K8z
322LDHSfRGDakz50B2dl08v3AuUAMNsMAozY+OtOyygdZxN32Vn7PCceg53P5d6A6ZcXNgEVKahi
nyk1QMW2kpbilziyC8E3HZxjLYaF4RrGnKUjzNKBFJSuQJw/CNO5ueLCGAPFoiF2mX2zGzd6df7U
Q4yQu4PTUn6Ay7i/lKLjXRWY7lYcErDBCy7eUqgrXgpIkjq4vgT7DZVyoTYf4CjQxq9BNE/WOJev
3mbhhcXxg85QSba0Ce/hz+JcfTyhHjF098/9JtSIPBjlbNULausSor4ncUIoIwVkJHAh3bR62+gU
nLzUvJU2PxoYya/IpFTmb54RuzjoNOx6YrNAXRDNemk0MOE5wytwnKtAPKzqcin03g+ft66Y924k
ZVE3K9ff5VA9vqKcAweHhxBMG65S76fhWM/GAdoa3G3dE4NXifvkYDwjRHxAE1qWG+TyApB60jCe
JZQeAcAaZN4PpqciWWrE9+qxvIZlJZ+ZhLGKx5pTbD7onKKtLFJ3rqkTyCl1pQ+MiOnLdhSMeIgC
PlQm6EZHZ0zWNl3urAid4lyOUGIQC8Pgi/9NJFRLJRf3R1QjsLi54LH3IIjw7r139zK/P44aNXRI
gatybIkTXggVouH9Ut+0uuxQDVmhJ+o0fPbDIyeecQVl6yW7BORtN44Fx7xZTpb4gCiSVU9VHSDv
4VYEfet4ZhDiYbWo5sLtd0APjWs3cRGrvreQxs2EKqWy7DL/+fNh4PrlOqSzxnCTJA/xQI5Qzke4
skNeq/WeKoa2rshhdzUdgc3gCVsNhIRl8qa7gnFubNoAwWHufMrBpYNGHg8/lW28mHY8L8xx4kS/
uDaQOwRRxoA6UGXYJUEQ6hKqOjrr8+i+HNY1XIC9SlYXXdb3gWgdwXWgQLQDK+aklwqH4yUXQ6lN
+bSMmfPjkTQNB3Z18j6gpFs+pKpjqNNcBkP9TPmSqNlv218D8sG7LoAOceDV6R2a9F+xzJL+gqCz
/TVqswdK1Dk9m8kKH8vqQj38jVhwkdP/Ots6Sy3gFJ3xVjBkevPpfxW+an/avN9NHgkBOi++oenD
Wfg8ZWOoUKON1sDk7tOquxhvGKKlaBQq2h9oe5TvQAwrC8vrvNkPzutLbAMh377mm/KM92C7HdPa
wdadN2XyXgFt8rju/IQQlOTDpLWZL8B9k0c8e+bA5P1dygHIKz0ZF8pq1C9T09LaWtaR+O8wG9zX
lmkZa7gcLgzoN/bMayggPKHG3ShPjRNAPjwwj7h5YwsUdl/SgYJMLN1WR9qrLGBnHHzcQ9L51JUG
dpjEjNBzNwfrzD7Qt5RSwU7ahz0ZV8WzjJ44sI8v8EVXEDOlldIFuyRED8f/XcYEVrRpW1edu6q5
83IZwoal5hzUJyFi4qKfBlvsIFHGWgMxmrllLcIQtVxKHrCZaNU4cPZDQ97W2eNbePuCVHW1Ui5X
vIFeqyC6YSsva6CJwm70ZeQvo87x50EAoW/7fHFkldGU/iXuzRAEqo3relj5ax9F27TpsgF44jXO
fqPkZSfQdN8IeTr+K+zBFeV9SW4yENNSGi6dgrFpPguxfqKpZMJk4+G0JiTRgAHBQmlAGMtdVF7o
LpB1R1Rt7x466ueANG/1RQbRZ/JxYcIByEwGyaFAwY1aNA1DD7G60Jb7KOGIxb9/NELZG8XlebGY
l36vF5oGaAgVzxaumvXwT+nGaaUlJxyNe+nh/WOsI+xma9uXL+bg2fpYmfBoq3llrbpmEqPRGS6N
G7/aG9P4uBg2tjgXfHTAl0gc1kMJfX54eVTMj1GBQemJjT4UPpsc6rL75osF5wychPGt6jp3cryH
jRc6IKXs4F+Cj+WFyLpKZlCm/R4ejLGOmP3562ypYp5pZfZUTgHhA8reXL01ibIqPxE4BOkhJ1zd
EVML73qURolTjSvwMKd+R3L2+uncqDrxJhJWrPjakXE/3Mhc9B2sPO88qyRNC/palQESVdoWF2yz
1N09htOM8PDdIVOUetSDl0cjHhnP8SRSyldO1DQWmnG2EwawvqW78L6aqeYNNHFb+HphGGodoQD6
lXbU1TnlrMPNqrSF3D7rUrhyAaOkvjPBH+Pxw3YG6Fq4RZMsXkoN9qfe9wAMljA2A8Q6QXqMpW6B
ezjrLhN4VnObLcceZwSeM988eUP/ZycnaYKVnd0t8tZ3QuGm5eFInWa3ELPdZGEhpVxoQP0Lfd2A
Obf4PFIJlI9gZj623WHLI6RL/ORE5005KzKL4LNrgXBpYK03xD/2LbWw9242p6Bz53THM7kijpVJ
k/P3tHsNKZb0HsoOYCZbF4FBsHzx3HX7res23XyL97UDAAtFxe2HifkCt+1YijAIT4sEAxykJhKL
jz5gvgqPwlftVW0/xWa3cKrOAG8MwtI4hN/SjIYQncliqOZ1bwbedF39+BHAxv0e1Ye8MngHp80F
oKx1v4k8murqpJThECIIqr46XMgn9oZ2EXBt3YMZKzHqcUYxmXYvIhPxbwd1iiwwFEp3fIqCBHED
9ESj6MdFOPUwBYkrzk65vYB8Sod2dnbtKdYK1heDKowRDvv7L3zlY//+eEE1fSyc+MOD5M72DPip
gCZuKOMagjfABTebAFVvXU9g6jGXeuJwbhCF8IuSbN7ih+SBkbtMWYYn8NHkl/AB83ZFhcXB7UTW
Xso71YEEUN4mtfBVKexi+UveH1kTnTOoHTyEl4XYsVCbaDwKCILVE0tiQ2eSvTrdhr5DFVXT9fkd
HtPuuLjhmJkvnOFk15IqKvgWhef2VGAvpi2Ov5UH5JaOvBIR7bRTc2XhuE9cK5aOl4Pk/iwYJhwh
TDmgg/bFLSPEQOqFGe41Mx8VZrzfiBy0Xzp28t+AvJN0fgJjOS/kryzo0OIXBJqhKEpDMWP0P5K7
akE+ZU9l1E6QRj/d1amtul+gdJ/KOokeUXiHE/9RSOns9BLqRZNnIHxx7puobIRZoIx2DBH/0WGc
uPWm4+iqbZozh8AY3viJsLiAh5mn576kxp+adUaTml9i7mDSta8oy31UlupGLFSslL4YI34LU71m
2sVtrI/n2TzQnZ7uDEUPTvF5NJ6htPxUKLsFbK6CzBRRgkNw66Mr+xayQOMVEfawV+ipQ8+ntRmX
plN7XIj3FTsuNQpCFw9k+tMpsmyt6JllU46hq0bxYphsxCj5Vt8giXRfRmJEh1jWh4YsL0eEfgYR
i0MUsuPWGr9Rtjh4mfuX8fItWXR9XSw6ekZQYMci8z7c10kjrMxoB6uX7nT3IktAfrtGYS78v1dA
dx0PmqWtl+QQkC4GiW4teW+s+mdHI187kt2n4AqiQT0LzJnbksIRS+e6h6wKx9WcT8iwMuOgB/yk
Sp75sYT097EAolhIQKXgMlZ3z6ygvWeMuKKnkr0fAsWKdbo94w+BS7U1j5XrLjmVQqN2Mp9Nw2Ty
dGOGW6b60I6Mqy6BFfYlNOTIvIRj4zD6ThYCIGAkZDbbfyfSqh3aOsLu88yBMeol/1HIloPVZviw
Og39ZVUJqiTwwlVat+i22e5w499+2wex3f+AhnyE1D2SadE53uAHHoZqF8aK+mK3IjE+7TFvPw7s
fcig53QPPSJ4YQXN4pkZkJnU5BtCi0jMc70B/r+NqkumMPqbyvVg9jmoeNw/Zd0HZ0fn+KjlGEAd
ywbfzejknVm/pUEuiICRs52TpMZG7qIiKIFGyDgM3k5HT5iwV4fbwFy04AsVMql3aXpsVn0lzscB
ab4itsM+l1vt5aZvAyBszqEa4HBKfsx8lxITRgBjgajIi+JRLI0moNqDHdsafXwRLngCDvqAjd3i
xF5L1s08L75MtjQunR1I6MxUtdJFE0xUzarApYG5HFYRKKlsaJtkOAGkcfgGkQPBYmeW8YOQDltA
uhoeaD3fuX4bZpf5kAuSK3OqGWLvY79AGHZjw+tTVuctj+TwmMPlC2kN+KH/eXZtGFUfXR/9+MTd
DmFlvfUP5cz2JOuuQhVzdDaXclW3VZMYEBgZWVTuq+4t+eZg0k7E3mhgN4nPu/xvts+TGm3Y7vPy
C2MqICeQGl/WwhXGJnEwB2bTOumgc3VRPv6WDXA3epOywkj1PBCXGrQdUjX2f3gYj5fY97EFfew+
oidYMPEZZ9BwSUyVVaYlVbYkNAopzi06HcP2Ek1hG37No2LtMnZ3pUSGVc5llc4gntksukq/zAuR
fp7ZOfPFfhp3W7nLqy6ur5ZIxoDip4jHVr6LFsxeQaTIsqz5yAorxkJCoQ1PWe0pyzK7nPKTVAeM
MAsZPNSXQnRYuZHMv7MBl18/JUjynvSZmw7EUDpRRdi9SiS1jAU90vLnI/lhF+bggoE4ETHf2aXW
klQLwu/B+jfJKIxeFVdg8J0TshIiSvAHjvVzGPDey4khkWQkJtwmFaexr3v7avE04yrngjBIbcrH
GK7MyTVcNutD0Pwo5nbtt2XG7QNQQq9hdJgUoU8Tr6d0ZHQgwM02bl2YowkpYjs+O6cwLDTcGoRB
MGBf9abweonOLVdWwaqQYP+VSVfBxM3UcZHiNaBHviymBNDEXHqBHYS8nJEs56eBGhgilmQcbBRR
gZDNkNVo8u0ZwcUIGH5aAndLs5lm+omRjel/HLluULVvNGgnJ2Rd7ExXBIr8CBTRZnR+oyzgbwDH
VePbWCfe7/C5D5fxMVIrHhrvn9iS6lZHFNgH661clq1Jt0uYTQjYIPo8KPda2leLtchm38SkDTLO
M4yv9D/ElGY42l+6IUwJHggyfoAWd2mbooojPztAqIxxRhJD74rXxicH4aLNzRPSIzqiopmt9SrJ
moWgsq2qEvsHo86ziCuLKVvCArnXb9cNMypL5xSFVgdMxdoiA/ca2C64m/Sz/Pxer+Mwswzot9d0
fzHMTZKGnfvKlHlWPEXE1mWPoUl9UkyIxwjR1uZKuXadC8ZFGbMWy+1fdDmVry3frd6pcV2MtPew
mWsSFV3D23vPiWchQNV1HhJvsAFpUXItpa/qKbZfF2H8G6O7CyhbctEPRIhDrfA3PBd7rPfO+Vz7
L+psJynCutztwEy/KX+mxSrNQOBOC55IKr5usVXsKjBiFofHy09E0scwxAC+4XXax5WQ6w24jmVa
iT1bOZydaTfqKyAy1h/zBggFTcose0gCEW/xyLvtfDbNhB5EEavqDcDPx6XbijRUrXN3AvkqyTKW
/FeNxIRhlAJRIonhOdNeJ8BTB4qr0Fj1G+onaUq240tEtdu/l7LKNUG4i11H4a/q2wzieMf2YPoO
m/OzKMFt0NByvlrwMFeBoqvjKqiieH/Lv0T9Tc+CBs5vNMe9h1OrsCCsyatnTDD63LtzA7pZ4Cp8
3jwN4FJSuQr0aOcrSQnu3Wz4d+8iFoRueuz3emJdPpMFlNPAcdASa21TccZ+SXla9SQ++hWnfb+s
1v5414qLoEy+h1Nb57Va7yieZQJ1Dg8Jvwptt96iW1uBd7M7i0vWONCNpqTMIiyK9QsHVj+0U9ZR
bGLpFRRlvur8pW51pGz2EJ3wLdjII7KlqmXVBGhsWb/pvnsxl7y1mAoSw3/AK2F7GFM9cADlX1fA
o5RsIRQkTcT/jnA/SeRQpTjUahXa1EHfmEew91bk4D9vLbD1E+9nmxkcrEbUrwE7MlgwrCs1tEup
u1a8JH5YNdr+teF/RfoYsaYBisEdzPfHbtcyZRcE2pO4xovQjtsSY8GygjnEQ2IWQb5MbbLMj0+N
Ht34moShqt+8W6MFyTkaU1Ui8TiPodGENtS2hP8BHpvgHy5EWXHu8yE7PFZLZtRu6kftqrJuxsWS
oAJxGHMwLt77OHkg/Dg1O5VGB0ej7udTHo7sBqqaT5Q7wIw+hvJdQohzsc1Z7N98Ixgmo3lGiBe4
WxeShaPmL6zpJMdRwcuGsDSv406JkbptEvIZX+4n0XmWo7FeKpx5X/pabazgRI64EToG6ke0a3R7
So9SHKqTp2aVWqKpErVslFqgHGs+WpQ1l12v1nRuAgxWF7PMTAutjkb/ayXo5qnp/ZhZag71Ampw
Da+tufvDuigoRJ+vf4WXb17pFuHsbICOKT5NP1p//Ar+gpKQHHQlKTK+8qapEUkA5xJf+F5HzhrL
frI4Bf1dt87IPAgbMy6E3Jr3JgD8K6pUDDSC5nEmbsOurAwzRz0WWDaTBZxAQNBI869+mPYhNeot
C3VGti2o5P2cuchhBsUK6uDM0+PluJbtSPRVAu/XNmbE2Wu94YvJuoDGbIH+ykfcZRvfCwMBk5cL
7jLIUg5oego9CzcO85GJBrxX2HX8CqvPOu7O/7HJqbM+ZJqC7UmVADdSZ1F8ZZOqcFCBViUaLNCV
thfh9K0sIDfU1yj2rjk8oZPKfuqGOG2x4EdFLz8nQWiHtJyZ8D3qKd+zhjQ0o3oyfw14XFnZ6MAV
K/TIkYOg+/4IlpzF3zSRBM54kmiz28GhHl4GDIMXxiyzB1GOZWTaRrPQmGVibvKIvgOYQ/mb2/Mp
jo/zoQATSSAfZH0+uzRAOzyDClAvWiWQn9cJn/GcUnM1olTscNLTl2Pvsiz8n8SWTKd6++RjPvKw
0+WVFipxPhNVXKvz/IS7dlRjg76Ac7i6PG/tsicWlMarWOvGnXyNXW7F3eckOPQS6pkaiNny0E20
6c8J5XxzOaw/nft8zVOWKBey7RwlfN9Pw0yDDODCWz4jAFaffjWFJ1VRERc5SizXtNPZa2y+sogL
z2bW5+Zh7Peswu85Yai5VPXTvyKQsjVDjTO6LH+xX6WOILyaTwjfhn8H9vgJPbK+Mj+9UORtcnDC
1sOYrXHoOyvkflUZHQN+I/NCfWt4rxvzYJpHVE9J0m7y/jUNb/hAK9t+pApVVu8IObzmx7sryF+X
F+Jv+99inbSkmaoC84Zal3rlzOsxF5pYNVydT7Tz0YFCok1RQz3E6LVCReHFz2SmsZHkaUgZtDvC
VWSe+YyZcmLMlV0d0xSjwnp4BdLmUBVCt4cT2aTaHutaNPf0mTJxHXk5ZVEWExoOIfTgdrd2UXn6
67R2Diq8RLSCfFHo93A0BU+6jb2wpWyY6KeExFwypqXsC6jhzG1kx1JfHuSmavHbPiFu5zuSqdFU
jEiNGQugevsupyg03Oqk43Qo0hSHTDAlrklzhZY7Gn4Xzo0wjx1vSZMVqNwZfwy8Gkb8iPbw1zVS
5t9/l0L4j4JP29N6ot0TMhGVi/CTVOZowIporuZYmKmaJchG2A+16RYLpWjvs21KapKSPgPEjLaT
6C6XQbWMBaDCpHMgnUSc+a58WsWweZzaX1k8vInNcPXFpErnDAnJ+zueqPBrC8oZlyWbNwTPuejF
x5WmSC9ZcIUr366CLZMyhjFj01fycNpOqtzeX1JpJBusF4zj4iU+6sPmD/aUZusREuLQx983+EYJ
DOCsdzHdVgYn6yuhVvcsSv9G6jehLcTsv4DpYnmOu1IJEpTQMHPt/s32SNx4hQLBBSZhx4ostyj+
4FwFSFnbW7g3uyZE7dcmgkG7GmxATMAnpVDTt0e+jpn0XDnK0J7iOltfgw1xZy4Y9d3eZiXhhbEN
YYtZuuHTSZi9iDxdMvwI5MceYkvbuvXLKc2h3nD8o3P5J8f2R1qYYdh3ai7iRFWVNGVkrlNze2Do
5cmHxRKmywu6Q6tCnJ5f2iLyU13OwsPoETrjSm7iPuktPHq+1FZObMZzv30r+MMkNx7wRC6HMYIl
/MBgYJpBYMRZzrHhGT+UNAUOuLT/91WaAFWLnQqLxC8ir7FOYlfEu12o8TpCw57KWkpSpKmxXEUp
33FBbyZPBjVaehJzbFTonXqZJ945eBtIx9IJMxYnAuzG95xypt/vyugXkfyOpmjZTsKVQi4HxJA7
nqR49eKANISZ8RiaG3DtepfezDK3f2846U4AN37Hyv0W8UQKmXRLWu+dAalRfxnXTkNzLb8bAS1N
wqhvZT/TksaGjmvEbQi9aImoZLjQrRHgZgfi34Tdv7x2p+D1sShRRAfxVqDNy6JFl9u3bSXyRiG3
7+DxLhVK4Cowy6p2o1CSOAIodWA8jJga344+U9U6czi7N5yus6rBkVNMqBi9gC0NaCtRH/NuU7Qu
71l0vc5lQOGLmTVLSjsrVSvBPTs6nmBo79Tt+icAzkvUv2pehCIfaO5MAwDXTX3B6WBpsKuWGiJL
URljYwRP63+bDQ9GnWTm56Xqc8fWTYmDOU0oIDYQUB4n/pQqohwi1xvhD/EiYXY5PtALVbbaIjc8
JOkbg7GfPXE9eLWEqp12zWq6kg3Dv5xN5KoC3WYx2PtyNTEseBHK+dSVVDxQTQiLP0ARlapmgs4p
rsPHdIDknIyvYi0nJLLlVUBhxmShxq0IaQJm90yS96dQo4vK5bev+qrV7m8aYXhcyy3oaAOXYteT
kmtXg1BWWaRsXMNURY9QgR2mflci9HkCdK5LwLG5eioDlhgNRqaJDw5IqkU8clnHSXxNsKKbR4eh
3AtctRvfRewUuuOT9G05MOHGbc4A/slG4v9ldhlFag9u+saSiW57lOKzAerv0yUlzaAjZYHXGjLZ
tU9pG7oJFQwQK7Vmkhtcr1YfQEPRKd8qeX+vy5tsv6iELg8xLHx1SCd1+IQQQu88il6tL7OCG1uL
8zNWiOr9aiTNqbZNzht324uqEXE5kkjtd/H+nyq2vX2rbSl2iUnRtygxNa//0KFVDjJOIb/APPlY
QLv6AZpBgBBX0ySZ/E3yTw4IqHF2NCbqgeEPsVgmpNA3AJ5/Jv6bzQra1YJUf/6RvWbcyIyONCvI
2Md5p9msnuIBtTBLY2Non8/vlOCjOJ4KeHxTaboVfYvg+ddBWYTgFhCkTibbZ29TsFN0t7KkJQvo
Z1Rzabfw5wldNXDzVGyOMQApxdD/TUh36y+I6Vvmv3lfQ4gUakFDL6Fpfwd17v/q4ChFPwhqoM0a
4TTBpu1AD0dGhwAG3li24LUalR6QIHl2uJorvcw1ExulREK0VuX0mzLuE+dyc1LMJu0CW731dZVW
Beqct9ZVnKyRdyVmqFbaRqsOETy40JW70inT9aI2GfiKIwy88FERS2cdybQ+kEGbs/PPneSh2WV/
I8SpkaT3hkiYrkOoZBrFHFaF84TeObikth1VrFc23glzEan5Z+6yhxGhkUfoZYht+sJNw5B7R7q1
hCfnCL8KGXRnLNzNvLe81iq3FW6iM9GXa6EWhjE5M9jczT6it+2FL9u0ciJBO/De1TH+hELvAPF1
0CXzJHhrr7biwNuHmzqC+edTEA88Vb0AI3ul/qLA0uMB09cYImFLq1aqoRuv/MG3tfNjXt4E6/tY
IQUY4zy1wbSlNMknPOXcKqOWAO4irI1zDPawxFqDR4zYh/gTKGZa+WWsOuV0LTaTB1NhvyJqChda
zUZSA53DlT/e0byKnZimk8grUhlR+i7ikUXmKdyK8EOYiNYuDgJZYHyyqb20n9enK6bLsBhaRx9j
sBBRb9ouba415ZC06P6WjY1lyl5Skloy3BA3lGRmHjzesW53TeeHHkHLwnNRAqrpPWlum4hw7iIN
25KiopGSvAI8DmkZ9IUKK5FZ9u9rdWFpElM36SZ8nvYoLdOLYPdsU9ZV41reGZ4F13luouBvd2Dy
qHYy1LVsVPVeOJ8UiE6L5NuydKNVhRIP+GtM4040roM8B8QATbf1xGxLboJ5mPCbPbZnMN5nT+5z
xjcNWUHakb8Gtpr9BoY9WAukXroMJSVpNcK46cmtL7uYBuxWP00Yx819u3/F6YOtaiePRWKBqtb1
INURSOUohqFtA+7Y1HY2OQLXkEGqEMltoSpHlbqkIXM/aR66HclK0yuUrN+m5WAB2gh54+PfN6Kc
A9xHnRn3JQFtmIOrBvAaQ2YDAiiUw4cU+T+tLJ12ZvZ9+NkYg5aPsTbOf2ddQFSnq/Gjbf5vqeLi
xwfwJRPIey6LQpBFPEEhaYMm6qEyREBlxJkK0jwESLe35LgQxuWHchuLFn42jGBy90QlfR2r1YV8
gU4DdgkLSBlUmG78wyy8Gstew+h5/NCCNIR7SPY7Yu/GfWtYJfOh4/9Syy85n00Dy9rI5QKI/DBY
3VG04p4BalY3XEjI3/EYI188+7e9YJBPVnANLh6e79RNgjneW8+m+4pjxUrYmr+kvL6GHRcoFYiZ
HSrhAtwoa/BLF2EH03E8tplN2c/MPsJRH0IHNl79iTfr/t6wyhakLQ2thB2Gzt43xULsYlU+McnC
OffXfLs77ilcCD9ErIejVtokze//NbKTAf9+nmDS03MdWy2PpartdeAHjXz7Hmv1bfJ38NNjb1v+
dcu6c7k6iyEx0ZmONpRhRdnBgGE306Z3vDEw59kwAoaRlnLSBa9Ng0Cg7zpp9l/xnIkxQAUF71IB
apNZKDM0iz73Caj+IOwYEbM7xnsndxmOco5QWrtpgXnyR1/uh61Ss25/nRVG0VoOncK0wdWAk7Yz
QpHQXwnY9ywemZSwGBBlX4u2r+fr5LlG5XOP2PyyJXdOUl4fGDqF8+Shk5qnitwEwE9nCfZ/1LzB
sCHlNuSfDi0Izkz1/Tuq4BN8O9pdNnGjo4ar4rgCGMvxAq/oPlvXOW6IeW8AoueHqjytSNrd+7U2
SzcH4rv64iVG6vvucZYqdAi/qqRj4DR6VwDOT8vxcjrwn0qO7tiKEAFeQzjCneJsUPPLkI479Ntu
zi5XY/4ArD4mfVhv9I2fAynSHPMFLJbkn8PDO8HMPB9jDXEQvOWwK4+TMCoJrhazzVOvoTbBp1YK
nmvjs7ThYv01/c+mLSUniO1zJCbdSho+ai7xfUwfpYgARnj6q0s8jxQPnf49+1EjGGqOnrPCfKiF
vhZItOW01jVAFfFKyhnsWMCATHOMbTMfORzms8SQ64sybO+T9imfx3+aQCOAtIPRDjvzWqXL2zi/
XtSm49t7G8FpnCJQhJe/PH8MlFljTWfl9Efzqneozh6qqbzQRwCFYmYvZS1IKF3VYNl4qdewidjW
y+GcyKPIxEyA/6bX7PakNKRbfxblgV0qF6dYHdye9h+BRuwjpQ2j/WwhA2x618mUgLlrwd4uQy62
gQwiD6pgOfNv4HP+i39xT1Kzx9qss8teTTCEE0+CWl0qskGldAXbaYzXjUx6ogu0ArZRuyjyuZ2I
0UVNPmqQeTfhfx3Xw5UAKeXNrhEKPvd51JUO7SlIu0JjPPZ7KBB7WDaKW4bkjXRYeu63nekx/jf1
ZFkezLrgXQWKNRaiUvFFcvckEbKwfvlr06UwjguRUJDqWUVQCP6ravXlQbTBtZOoPNxn6Ge9LawL
JMIX1VbhvCfQ2+8kSohY0ZpirCvPjFGqftwlXYqAgrhytPF/Qbq+QLkjwW67AaS3zRFJXBHi74Kk
CYsHY4UPm/zwpYGE6yA+nL0U8bBKFLPNNMbZCFGz85KG9v6/RArG589uiUEktjL8Tp2QnxI6/Wfj
gAJBKZLCgGuQia329YRi//y+TQrfs6A0h03tjxqA/WOVIgFz/Tfs3dO5Ef1MYANOYZ6xC4SF7bBr
0v0N6ZjZ/Ce75HXk5TmWmWTxgOYY9hB8HFNUs4a2F7vffgWsVWtvqNoH3NowiyXkdBAATAFNVMq+
5ISYMH1a0cx4oF+BU0PuJsHeRhcDGPLEOyPdFZaoMPvuf/yE+bH0YisEQEYrY1hYoJlwsSb6SUdg
M0KHLw4Ht+LSmjyaxjGNvqMZ/Cc8C4swP2wcuM1KhrOIGBbkRH7B2tCgJw12c0BtOPDjQJKLXNtt
6FToDqhR6umG9D0nw94yGacZw9gZzbnRwzw+C2Xoen2zE7hXuVXukHNOEc5BQNXgK4ZpvwJ1hk9z
Q2PvG84MDWrKkeYuvDsbyH4h1xF5RvLvFmvLxgYlvTx51Tb2CrbhrGpMmPUpytf5NcAbsg+L+ZT0
Tg8rpzOEINnd63rvODqXZOAtj92/zcCCmRXDx9cEQoSgSxFMbx4m4Q5Cn71KIKequBG7lPog9yS4
3X0L5R4iy1HnUPnG8pj/MOcXOTHhBW/zgxgBeDxlzV6BziNw5LTY/F24xJ1fhShG6aELD5MVO2Ej
zchso/XAYTy8sudb0d1wbMFhG7JxoZbwpmUgsEWyalGZiQHKGrUdvtU8V+zr8FruzJAexdpzyHCJ
B6T/cIyxH6hfyo5d5/V1LddJV1XaHoAqaRrWYQVSinYu7dRtB6W34A5KWL+Peh2FrAahPl4OHdMg
ZCYOKhuhLxgonxvdD1AZsa50CXzZWOQ9f7wj9jbu0eqXKMNOSptmMRmiUTlyB+VL5+fHXBbzPECB
v5PUxXDHePTP3By2rCf7iV0wBcXVLk+KP10xYWuDgpALGFaVV9aE/9OnlQ6SKVjQVmLkm2BHn4Z1
5g2mIO2POw9FWJve+X8mV8lmqX8vpBYBptY+YB1cSruvB4fN6uLeQe6/1zMjgIFGPn4dTgvjiaCv
UZl/xrkCWAUyAZIF9hf2xtJwOf5+Aol4NgNuTSl7X7UACLV+gXF+EXNLX+SPJm6nyCU/S54ydfmn
6qI3pGNTnzTuqw9aPo5o5+j+gApEM2MPvZBcax4+nrKFXVvGRnPggyG5JEWsTs9xrxoSSwvzT3+x
Dvu6wvVfZ8pvkuzT+OS52w6FJ9rTGW9NrmvdN6atehkECuMMmZNSy7A2y9Ch9Eye/0GQ+WwaLxmQ
+VkucvLfOQ9w1pYKIAMYkCngGXW2MvRx5b7XbJzYRhEw9d12lreKMC+x35HGnP1AwbzKiVx8YOxL
8TiE2wbnhpWcK603wGgTZhELYVfb3OAzvc6hLrjOdEdKYIAQMe2O9xVOZgqJnFeyJDrrx82qqw6x
zu1efdartoJVl2U4zsnn/YDQOARsNGA8TfBIuDh8Q99JkQG3uEypzbVcFus8mq6E0ujLtUmohWMM
+098mdcAD3ilWnlfywuXeldEsHhXt5+lGWpi1zSQ26H0lLJst+3c2g78qBjLucFB7/yCycYS5c18
8RDE+xn5k7l1H71fTrqpE1bvV7cLakZcYjIiE+QuyO9YWhwM1fjpPTuJyr8bJLq47j+aAiRQkHXZ
50tuAQwYjJ8iijYJ5+8ay9Nnow8sgfN181fGogIHc3QW7HvvO/P+oSdTJ76Re7ZTVWVEzIVQNLTZ
JiNULUXuDMhe7cFl2CthVQdBsb8dKLvSblWBMMH8MpUB78tUiENYbXxylmFk5niAsb27CeXmlrMh
fkJblQCiAjCYr516PHHDkcozWAh/4HiqDch+hKCefItgsXA3lcA7p3/sMQG8SnbsUayBLuW11TC2
h1zt3VYbbI5D1HPuKUiKE0gYOMfXS0tZAGYG7G2L1Xm5Dx7QJlb0NhTxfk1j+61GTEjNIY61oMVD
Jxfme8Ins76bwzMYpPE8h+uF/XgxAk/crLOaK4hf5uNf6T/AdhpVwJMsl472O2SyaRiX4WTiMjQu
lYPXZJTdfbQ8OIQoyjtpsxr3VNU1MpYtNn0N48YNjvYtVUn4OMaRdWT6fkXTuhoFiF6rO+CMx2/x
nW4xt1mu/AZp1eOEpbM6rS5+g12Bp1NHap21EWuWeH5o8X3rHlX6OOlKlkiWviLM5gUkObfnVt0p
VKkX2hNuPK5o3MzCMBWhcAOF3QUG+H0DBb81H6OnhDdRG3+MvVJoRPqdyvS3BisysTAIbHZr9hjk
UlIIRYcpmNZVqDCO84ztYxhTJUG5K/xksWByiGnfaguifUUMF05PeoWojBMJ1Frtsu17VKLeMC0t
gM8eA70TB22I2UwZrotwNFq7Pw6kwb5FMvAatVndmsHzRYn/yo4ebbzYFNJwpqVEZGYwDKGnz5jH
QhhVRtFOffOznxDIoUiWQ8gxOY2+nH1zY7AEbCw3NoQrEjpYgaBGZx00a7O+gt6Ba7UMt6tPaUDk
npnqYFq57OiC7ER2iKz/2prXr7xrMIHPExsk5gshke+qseV3p8tjMhugGNhfKkoQ0K1w8E3PWi66
/ESpCjF1ce1BMdnqDw2b3gcGQ2Yc2hALUUIxStSw6HIJwVj+oFu8xaziTwV9n8dLDYf69cjpeJBu
bh1nfPuYlsGs0CC04dXFkzPo20SoEcY3g/NpBaeW3ROEYp2J+OokUKAjzNhTd961IP0G5ltvborM
GlP7PJf+XhqKDzCq/n/s6735zUERgjZ7QAqEI8Z/Gpxq/hex9Ilj7lFGV0+yPgB+X7Hm4eaV/GDk
XIEV0SJ15Cf95Xo7QS7S9mPdPxl7GV3A6W4ng5eO2C3RCZVMFjBjpYdaNXCJ5632yy5hkCyL4fTy
vZCuYK07onpPdqbsWH/WVNLZ7frFN197MvMteCvqOqZ2oFt0DO7yP2753+KYBs7VMmmD5hyxmM71
nBxVEw+YfGRrDx6f3XmLTtFwd5Vf6lxlXrcIdC3fz+F8oZT8KU03V0Zx9L0ywCD3QuSrtK1ZAKoP
jJOZ1r9fwYNVOGvSblfi0uXg79Yp8OqUoFDhkg3rVLFJMCekufIuAVaZthrb5I2tsoVySAGs5muJ
LWOBaL+N8EjRQ8YMZickPInkSjgD7jArMNpGJXz8qACwzG8b2p5rOzswwei7jEfw+jxiFRaxZffV
qidvC4uzq6cTvYx+dX0FvMtXrAZ+cUzKlLNO38V/Jg0o275Z9PgpAeIXxDVUixbhoLnoI7iALRjl
wsoBuwiCGzuVASA4/JMOMFqZIdEJe1oyR75NS2Pl0l45M0v5pHjvS9h3tatKGlDow0of8BqrgvRk
JGDIS2DG6qjI5OVYUYbteGlbiebriZyovucAwwpiBzeoREG9x4e6wt6DDIi/4wQijlSRvGIbSgfm
FNk8fzhI7MQzsD5hnKcbp0QgAsmwGq4snoKbeO1uu6LeUEu7HHcLdw0JEcvNAdYFHuiYlYQSomlq
l4bkHkk5889bor385auB801CgfOkt5VIQkxbZk8RD/0x5iR+e8SwtX14yZzwqMegvWYBfy8wSkmJ
ZjjTDgVf88bcGa4NqFc7wQNpKmvxCh7A/tDY4SOFY05Hawvdxhxl5lUjoO+ZEjuvn+o9/U/ca6iI
ZQpXdbgdHu+upx+vu0WANyJ+r/lwrVIJ0b8JzGtYF3NANE6m/oVk0Aw9GUC8znu4O+mGy7umhESm
RHILJQUzF40NgZz+xNtoBmZOgMf1SMezYN6vYxWXd2gDRu1FaH4v9ctkIeBDczsCSu6h1MKKo6AM
d3dBoSrlyy8jivDkfK7FN3AlKt6WIUqQCP9Ra+zDKH6DJ6kBnYlz/2Fwh1ZERlUk+mRKdT1/lIbR
gjN18rCuRTivcHlmxulOlj5mLI9B/KPiY8Rp5AtWB3VvSBGlkdRvyOjUm/vRRl6qengjnkrCQQvl
5NWFJsSQrCF1+xFmROdrKfG10i1vCRzjrAwkOIvVSvRPYa4VX2Y5xs9a0D49hYedsg5ROGtx+YVo
AU8LkJKwoLH/0zbA9sPFs1HPqGHohEGbSAloNinEnm6lDcUMXQ2hXXDc6RxLrppexH77rLxerRyr
DGa2+rz9Xdlbpi52EtIzAPC7pYvX4EDG5lK/Wsc86zLJiK3+EcfIkHMuszobiD/en+MObS1K6QCp
fqdNemTzpdHgpN42YyybcrVcu19XDsA8RqJ3tjuUfvA4Vj0H11wimjEwm/vpeZibCaqpGGLCN4tj
3nLr6QPt4BKBTZreXUkBQc3B4l4dgnOVZ8n+OZUPlwXMBJX39UlI9UreG5EppaOOpaYz3NjcnDJt
hlK+PyLQI7Xlc0NpZUJ3y8SsWnNyGGBng6f0c0aOpPpvmMiUOypspOpqfYIhtDzayAez/fqKMOHM
95de8/XwEaai3+uEnuViAzvwb8QuHkeZMcRdmVdjGDu2iDJGVfqtxv65vFI9WpzuJgPyOPxMFSMF
UnuLfQ5Kwh9oYKngWVaAqSB/JcNjUGkPwNf0dKmE3ZvFDD2lpKWPqYGl6HBuCpZNwp9Fi+QhB3eF
6cXWCE/c6jQMLfnz1dYknH8PwX5rNjCapN1p/6QJqA8JQB6rhO7Zr3DWL1rkb4OAKndr473sgB1Z
TXHaouLmip/BsHsYauzZ/wmCXpE4SwojKA+YiCKFZ7IVcVc3/7i4AMoUdBjptc+7VSQhUM7GCq+j
WMYcDlj1CLt+aut/3ZEnOoB8bndhWWaXbSnEiXiPqMmEavNol5gPbmtjFHtfzJead5lfy/lKChx3
93DKQXIeai/CfDa7odkkrlAgAX9cfm94+BpFjNzcfw+UNLZ2kjMPlXmBrcU+RVtU/xPSEIFhh/Nv
RyPrjjyNCwJJbgrYF0QcYpYdf/wNS+PsHDq1yykhxYduHE/l5cvy314Z37xmbUQ6z+1zB+UT/kbm
FDZFr+upo6ui0K9k/dfoCCJJ+ZN92NcCdFIzyCsfLmOZMYfRJnM9ZE7akVCN46Kaast1jkI9YWpz
N6ILCw9VEmyINveiSSdLrihLr5XnR3hWovcpQyI9r2RCinINX8Exi14/Xb/t1vkYYCwc1uTWswBF
INRYxJB8Oi99VNFHCBlq8FmDH+NeegYdvtmbePLe2lFCLRX6FDZLgAR9OzsvUXI3Z6+shdESWg9K
heTOX31+y7cJjhLZQfL0Jd+nchnNBX/YVX4WH+ESsEfZZSSm5Revsrl2YixYQobIKm82h8bVnXde
GnIqB31M3iQRGHIM4R+Kvme4D+JkBlVg7ztIbMWEkN3kLgr71EslOhPg1Bsck3wJw8/2rAUB9oy6
SRdqmHuZcZ1PtDQMBlBWU4VJ1iPN418SqmGEe3UCs/VQUglvxwotQMz0pqYOqu2FthdEi9N7vuMC
lNjKUcD/i1lpz9k5HIii81UMyjqFVNtsQ84fncEPx5UwB+QdgQQka1fL5a2iwh/uIEjIlSeEeFa/
wzjLrXfCLOCl7koRJ8F1bx9zgqK6mmdlqQUQCS/Gpm94b4vn9iE+FWPwdqRUb/i8uYk9tHgVsyCy
NKvoZavWLCptNWgg4wGXMnDhMYrtfm8q6ToYHTkaP5IU1re7C4d1NcaV+XB9wuuzhhQa9EhE/FY/
Vj78dSLQrjBJ6DU7hx8jqME0HTKAQYZ3KcZoBaoAvENNC6/iHen7ODv/7rcMZhSFm/1JqjYQSv7r
f5glmsO7LcHhpXnUaZ0kLbECvK2v757paHZnlOjzilSMjGtszwWEhDCLXBcA+ytXBjyjjDXZGzKK
sVnpWrwdylkDVP7piLFQeh3drKJKmHIiYxksHI3bjlsK8/sFr2gMJMiNUW0cG2IPWsEvdroQkla0
iXCNRXnRTKN6cDhYmQ8uBMqrcLiJH8Vj3gicoPvqPVpYkHB/KLFDxytGeKNhE1MtdATXJ0wyYaUF
beOKqlIqJaCL16sJ+Wx2wRNQ9jTlHwlJ5cGTYiT6gYJ+OMgKf28tMoVfd7vPoBe2ZUW34IQqb6Zt
imxRUMb/eHho7/Eqd7TK4i58MgyuJ+cmhMOIXqOBsOpbLF0BoMcJB4+R7IUgEswPFQ9bw48kB8iL
Q3QkG6X1qFMbrx4bYRhbsosl+kE7gKG5IfgrrZi/OO52zZ0oQVM20YBASyPKLGWyeALlwBEZrHXI
h4etMx0Od3XXqKJ1PbPxkXXmNgF71bEkROWQC7KVVqTxK5lS+I3E2z6dqc4p4gbcSViPYQh5/ohc
7WZR+fR14o3lJJFgLjTn3TvzozTBP7btIGBlfRAartC7c1xyU6UYwtJjQ+cx8r852kG1RgYwT9XW
ZAcJe/Oj3cXPBg2Gr2m4U9SVxTmngXYMJz+QhRtkgUY/QoZXxgWU+OOOIGPkEK1xw2fimuysbtrU
77vfbUwjAvbCHqXhlLxvnNt0Ov4e5qnR0B5XEbdQn4DPsfUYCNgsPsLiu3JZM23vs4MKvPTSp0xo
HALKn9uSiNjIFdTbGUy/IiFOYiSuXUPD8hlGhVIxnRzzlMhy92fcIfCOSA6cpw3u+YEKunCyEkT2
oNRFI4f8TJvQcXYFvN30tQhkcdpw5b1dWWujotmgaBfJmOHA353kbywkExNIpbtpxZFh2I8dcCxb
ht8l+85Jj418UyoQ9TXBfjYqj4gd3m6jVuf69bIhKW37KYIKS80aJau5DgxSTLJRMlkIv4gr40H6
3fJG8ZeJv3+mf83Jn9ayG5gHNE3AsN+F8uSlEYu38jQZLtt5/oWO3nHd2haxJXorQ/Oyv+m5iIhY
+RYi+HO4U4RYHBOU6nkKQStPQBnM0ub4P+5I/Ple0vAwH2I5SfEK6soBoyHuZJhQo0CWVjyOfygV
5S6dBfT6AfXOhJDXQlmjy9aXmwwcjJuKR4qnX5zOvV0SoVg1G7UxEEKf81PYu5bGMREepODp8+2w
9p/fZeTyUYamhIGhZid4ELH/MngNKPeXDvUZnaC+IM2J0jFLud4f59h25H+bPREHiE3u4hdpwoR+
gllhvyfutfJ3UM6y1ccFpNaN3mmDVhnSp6lqPziP0m+PdAA2bh+QZdWBv6LJpU0ITumiQuQXbala
MNNRBd+1rd75dnyC0pDPluJW+5MHm3MghnMifeoHOZKuPcrOtjEJzc2Kom2d8yw4iyg0uBvy5Euh
ps7cHyTSR2tQGZhJQ3/o5LtAf4P7vzsys/J2hb0oU04Cvhs86Cb5aj6Ht+ZznUZRI+7o1gb3y8Xv
LKyDtr+kxH6uFLUPChUoNtGn4x/2C4gMgXNExQ7c2iggrRHb4Q1O6vda+nHCmp2ov0T9S+qqqWft
cSS4o3R5Ytrd4FnwNEo5aNU/CIVoCsaoblW618Ct/Fi6ff4wjHK1vAHI5Py91rXNRq/R9GqCmf9+
blXBA+ub6eNZpnTf2zQk9aCJove2yIAZ5Z4FcCjqxqjOE+aLdh0hwRcFNUaCeayvqDSL31O9p9Mq
1QD+h2zfj5YRy/6cIZGpmzQmKRwcJgafwIGaieqyS0fDupR6P7TEBHwcoeSm3oiDQGrZFwleAV1g
BnH3/92vYBoUyeTQYgpOu+sFPcI2OA6NL+2Wc9QtFDxpITDWjQ4ur3uWmZE9gOK78DkSPvpsA6Ri
kuW4fPKZooIsGCA+J3BJs8lU5D989mYq74Rt6xWXoQh+F+YVT+W2J769DwPKSTR42fcOxPX+f/cJ
h7DFOsHUXSBSUa668z2jYL1MPnVtCH7japqu4ZXrefNrmGl1rpRViFj7zYEz0LLT2tQ1pkCgZV0f
bth2aFgX63TsKEPbh7P0lvp4DECIpnz7fds1maB2fLU3JdoMc7TIxJc1wE0ydRXI/VQHkMaNovHj
dh31K6FwPtdww7ac+A1ZH7N33P8rxHA1i00OzRtaR9FBo4s2qXSin1E23CDE3u93vPYpU093SQTr
qz+v7/+k0KAvm5q12mTbzrmZ3RBcAbnTRds3PWbonWRosekCZ1Ap0ULMCGEpsBPMf6Hm3NP7mNr+
ZzwW8dCd8h9x77j/E4/wGu/onaks/nfBCTNVBbb0p6IPhTlbz3a1bC7nPxqXr15ibXn5mBtrC2em
d2tThQnrhH2B5Etjqy/rrqBm/8lDJCla9ZKaBITM1GVUJxg+OMEZzD7JR28mLRKSxMv5P9/xuA9e
GNmZhGhcw2liPA0arGNOW9ykxC5W+0Sf3psBtUcR4XnRiLMmxRsJGelrUMT5YBX7sOUFmm4bH26Z
DGQ89T8JCtCwIMQSrxuKhXmhAf/a9os5jYBT9okhhoBRLjDX0caV2cIL4RAj0BHYw+Avy1Bvcbof
tkk9GWGq4ADxIFoAWKs1vOxckZjwGdHmj4qvVBVGUi5ly8H/+pc3leBlhIb1AKdmCt4/0YMzoDRr
C5AekTQnpd1KTv6X84hm44ORUYHlk7W1ibOTsR7iEpj2TY5HEu+1xvot6hjX26txbpLiWQs/5q2b
XTtwjITVOzQFKlXfHlAlnEMgxulo7m1cvIOARtoSQ9OCj77zGgBuaHG3SWALqBuMxyICLsNNXlcY
mrB2gdHGvywLS+OKWoduGorxkJEyfqndmBx1n8OrigqueErPwfz5bwkI+mvI8tTnKV9J6f+SDbdD
EcjOyJzHx800qiyakncM1hl3gnehT4FJcUpRGQfOyctyZWq5xq0+Za+/yYE7/mJw8adxxYwMAhJr
NwB1MMy2NF3wmH5gyA4FRTzPckB7QeO6/qnK3/fxrirus+7c29RMqiWqse0ixA3khgCY4Y4gY/lc
CLdHcW1bfwRPSdfLrRiez8leDNT/pANOkNZfV+POCz0rGJoqnEW0142aqLQFyo6BlLUfLE7+R7m+
ZYP+ZWHPJjYwOGofpfscht4HgxgBCa8KMvJi2RQ9486OIa4/Shif1PBOLRQAmOpRlgU68sHJaO6b
F8KZlkdq5cjtdkksdNK5im2d5mup6WHPKlni5kY5MgMrjMKxwQpOson2OeZz/l5aLKrRiYBEPHm3
x1WJE9ormKDSDFvu9p3J1vvX7oTZLne2AK37VXu7XhVK16Fn0cwyZ/I9FCaamN7Jfxwr8zGn00pp
ouwrtqcQlEBmlAgp3suuRS3dXuA2sSljZbVepUgAq6EZ2i+p6zUwv3Y7dLDw/TR3doYBGCAeQ3XP
ijj10AFFHZWQ8f/cZEWAtbfBGkQWPPhB97zVhCOENaeXFoeUkfevFskFKOege6D0WVchbtIQa6L/
mc2QRhs5vYazCWhl/wYpKWfGe3n6ogUUlEA9i3NxUe90yRkGhmMK40gz01VpZRodcoYqaJUZmfLf
bWkM4M2oeANGrgY9so464k7iyrsEH2m5mdpLnMn3QZtZ4QEXiuW8uSQnE8uLJqwuRnQ0jFgVNHu/
XyubUM4VXqYymtLDQvZ688QXIsxvJntDeIz7aI1w1LF3fkJdofqe1zq1QkGf8kbj2QMgQfsUHtc1
ffUENfON+k25c4vu6XKc2NWlybZ6X1amLEdcw/1jP5r9cbtIM2KpbuyymeYYSYmuC0/c514gAKK/
blCSXnEAQVBtZce4kh12n48h6Yly87pVmjk0/S0wOhdJzrD3a4y3zdSKqiddAcvjNiy05jvRr+rk
9lrmi0XCcUHTwGOyNCfsBKOCAXJLIhG4lQsxeS3HbsidIqbc3yddnT+Ze0k9RfyCY5FGRCYzOHZQ
GVVqw8fI0fLFku1wl97zuL8emVCsxuF/dS3VS7OkPl/eS104BgQWuP5Ga/UATcNKUEuqJ2hGrUPL
/fJ99Eqy1vnvu2TUrrP1MlxBXLR0+CzCj2h/4y2tobByRIFnQkRfbFL22O3J+T1790vfAi7OIi1L
/4GaJuHCHTL6pF7nHgrn+gqNKO3KZRzVylHQIiIcRCZLIPNX78V6JMLrUIrr1NlMV+/4ev3nfEC2
V5ACkabyhoyqbTe5SXWpIt/sjJus98KcRzvM8qF9omZMD/cCC1ZVqLd1NYCFMWc7yjIfAjW1XryU
oB7IUgDThroYXcIf5aby920i94jBwAJl5sWauHLl0b2dhMAv6tpzgpLuY+w28ozpQzn1OXsHUuKP
YK78l/rl7YouSDI0FCXRMH86xusBZZRqycbjIsJ+5EkPit3voAG3YN/95sPsjcHseLpZVWWVQ7X+
/l9O42R94+9Xdg+EmHoE+NfF+TjhBLIoNBxzpFWAsi1KBAciS6bbc9cz6Si1Slt+2o3z/YrxMVuV
1J7HF6Gq0qioOIng7mSaQ2hQPaEjGIg/1q854uuK0bYnRv4gzSAoLQktMT5dna+2ol/ioiNN+gM7
PjjjJOG2lxKx6hIH6N8jXT2GmYty2IEytoArleQ259oM7Zx3pTCYRL/ANStxOqqyM9Cexak0nnP4
QntqqLsKTXCvLMcYSk1I2TFj7SlAsEUnyWXN7Y3Y9zshqAt9lJc1TL6EFoo53RuHgN02YvbLzQgM
VOztzTtoRJWCqAdHiotGUwFyC3/4I0352qLuNm0I3TOkfLBADF9527L3iSvbOXjzJkm1s46F6fSb
1Tjn7Bao//ndensiupMg6OblXA60T0d/yTrRqLKgts1RPi1JpB7JFp6LQ3XpCCUQ5reNitq4AIAI
eBo5vf9xPZqmpPSnwrhgMuvatMoD20w2NctM9QBE7qqH4/2BH5qMhbuG7K1IzW/+bl6RHOrqT7ib
raJA1gRD7YpnPrRxXq4SviPMSTtPG4oxpuBVV64q3tLQMA9REu00egFEw01zVoO+WPgoiTKvabp6
yHEFwYSpDnd9mRG7+FDb3afGVsr7C4kBrB913FR2kzKYq1TJRc6T0Iwj9U+TfRMNyUtBxYIz3CUw
fB9/45qKzOfH2O9em9LlCFuoPkSNMTyLPAFLGaT8CASGRVkXuqBDjIF66uQjaTsM2aRcfDtxOt1c
1HuF/brGrtoPHObYdVar/2GsO6VLKAeXomwVvooS64tPGqjuVKzBze889anq16Uf4ykDLIF0ls+a
ehcuUNvpoODSo5oDQZzZ9V+0CnhqYcAlIRA4V6X7fp0z3TD9/WROn/9c9YzrnE97DUYOHwGZvhQ2
0cjhcWXnd0G71X3udnsp4Uw0uLkxmEUTGaGRm2ug++ETvxzWi7q1IJiSN3vCHTCi+lItU0MNMSCN
nemSLh6GJLTwSZs084azgHwH4esD31V2wtMkTv9LjyE+0Pj11JeaZnUYyWOYRGB7iXFRc8Jl4vPl
313k+II4u1f/KonHx6EC9PfV0Ys8mRARmP+0hAHolb8P2+aUVddGdMa/Ziob/nSAmCWKu6/k3Sd5
hzDziSBEL05s4/OWzS2QWilSLmFh5eCT/cKhfL5H9A1XCTbXGDbi+tD4foFXSz1/t6uZ1ISzJGnf
zd/md0dreh/t7+4jp7zohZs+sFT1KySMu1iJ00biFJ+7MxouicM/rfwStrvESqQsLCMgRmDBirs2
an2AZMv+rwKE33cO5TSIKkI0CPRrL9zYnSpr7OiMB2QEcVUF9lhgZbuiGkMaN4veXwOIGbO8VIVI
YGP/fMTcc3XKt8c6oxPR9r98Hj05AXF/sBr0eg5id/zDS9gx0kdFvNj2o6fziHiB+GrGnFcZJEtK
1/rrLlaT+KpjNxXmrD+FgcYq7bg+oQVbAOiJ6OZPNHBoO9KWdzzOTKOWc5dmC+aV9hWAZvEh+4F6
uUEZBHU1GSU3YO+gqkBK0Ol5mX8vCydDbtOs2iDSe36vrA3ahV4Br5oUhhw+aMkBxkVHdZx/00Jf
IbdbgDEbxVkqUnE8nMHF/1F6HZLS9F2pPpq9Rwy1LlrvMdw/RgkvJwOIK8Cwt9yWRlLMTEqhfCkp
6K5lZysVT7iD75NX86msgE+xpb9/WciTgPhmeeZOSGFEHT9/VaiiR0pKvT42iTQq6suvTwXjdg5m
xWnjk9Mrr9pPsMD1CAOeDFYqMeXJaqynT5RrOqiw8oZOrZfXgImr1uKfeyQ4d4QcS3WSrHCC4mEk
5vdW8PfSKMM897RfhGj1Nop+74XFHpIzTcOPpCxuFD8NkZxpXNXJn6sRZ3prSwrtqGFe4LF2vNdq
HmmMpXho/T2OPcaDxJPFWAo4xs6twHId0c0b0v1K9YUkgV/itsh84zhkzsIWtyOfTiLV01tAZTdk
2xH84DVgg4hT7/rgUWEeOl+LplvtReJH+nkloZXbp50gQKOHLOFdgFqjHFue6wPBErPHAfKefJ7b
34Lu3y7UguzXQ/sblBeizwC88SgYRXzNtlaY5y3wQJRuC61lyh7e2jHhoKv/j2N67Am9Wj5gSSwu
OTtiKNC5/ONmAOCsmhvyb9DMIcJDegybvYbS2uID8kpJlNwDczBjxzlwMfqm3T9g/o2nI2z48db+
UIdpki2J2PfZiRKQz4KdTyEb7m7tKGv08xSemC7wXXWLAMLKzel5z5jdo56iSE9At2aUotPRoaME
xLy96OK7GenB9FxENT3iCZoZcRnh1Cm05lVFOvft1x9zUANfBO47651I1y3oV1DssC7dlSG4NSn0
AoiiVYSY7xupBNGZmDhOw+ZEzKvmmZXJ1qjIXAGWbt0OnYZXXO/zXXk3ysSJOyCaBXUJ1MXLTb/C
MWInWNdGKD3pRWy5/P1Swt2I0NbEmkNetolaQ0WRHFhwCL2ZGwbVFzOt0o8Qz1hkwZP2A6W3Ywfd
TTlcuJHRZlAiHOF+/Xy/SDws7Wuq1+rceVzsTF5cUu/ixws+jv4611oJYowlH73+5yrii+XMiCMX
x7EoSi54np/RHjmnS7FvqzLpHDBbq3x5Vj3gMtX6LnKdPzaQ+EK2bn/R6gTd+nccTyXlEG1FCzyN
fgWhJsKsK3w425FdTsC7VdbO82eSFF/4xC0ofUiMk/IicsavOo6zFpkLrAN9NsSluYRUC9S+Jctl
59Hhw3ojsJuF5ISvjw6xEM6BIfm5yvCRbBSu+ze+BY5+eeGTI8+AneDCRYBANoNQKCuhaaaie6rP
iMRn9Ev/YZyyVDSVP2mqAVde0u2B64Qi0cIk07QP6NxrmZEgcc2x57fP2n2BC/TQIBTztPN8dHOi
/04w8ZRpm/CwTI6Wh/k3SLc4lnW4ZnSfE5zwUq8VT6dS808c/o7cp0OcV/SvliIIrL/byPPSpwqQ
Gv82WphIhCeqShJYBkCDMZHcptZskACnEKLYB1ix4/BTf7iZRgrIbdLp6w+noMTgFS3W4Xp5xVX+
WNU0xo/+/WkYjLmpcGFgaKBDsWStnJYB4AiUarbLqKtHIPjAAazea1j31zMGOzY3aoTY2lOU3ZBq
1GQP8kIvnBgXQ7R87iz9zPyb8fB15xyFpYIIb4CbpNTdgudK65Ix5BJcLaYmdsO0JGT0RTxukWcy
9pn0rqlJ90gOfhDx7ow04F3fy/ACiC5BlrtTt1PimsY4QvoeUAl4ODtUpZtd8jidXNlA0GoaYYW4
hUllqc2D4267Y3Mec858QXbEn1QOsMoDmIHUdwuaZs/mXpRXBzvXFKX1wG0ogC7/lyhw4cFYzX+T
NmLehNM1HEGzyppFNOdOohphCZvcEn7qjM84E2zqw14OYjG1XIQicbhsdGKaQWpaU01hWzIxEB/Q
287Qh8wvEAUWFV9bsuftHI9oN0vJZli2aCK1lS/jhjoXH2AoZ5FDRlc7w2zl0Vvww+C/GDLJeLJV
1Q0VkOqvOO5dW6Qw1BiBDPFYqy4AwrqIC+vQidcBjaiZWWOtWxFrNcqYor12NdJle6hs1LhoqH3g
kfkmdscpOLUFZhdhs+FmzEJb44mIETWUt0DYdqjOjcA1UdWQtuBX2iOs/+0N127UAzA3a/MduXPA
xy6prgJj453VDDWE7+TriceX2BKpfTk8UegC7FbomcLu8/jATswAjkLi5QJL34k5ovWA+y/YFVHQ
qLP3dkCp22TdFA7UA6hdvsfbgD0dywQES1ouWIpRKcmxUyxWzIUqgQnPjWs27cO6nq6RzlixdMdE
7sq3I7Fp30IM4nB8eR4oD2LBUtl6Atjiw8iHJWmzAau/RdZmr3hjvwrWMNLhB/69d/bqvZd6IFue
3Jx+pYltEPB0a+nO+lAhodPHY2/qcUu0VDt5OLz7Qd8JoXOO02QPFKdYVCQ+hUzdwFbg8C7/m39d
x/RzUFtFjC4//Ggpnez68BZUwm9wWoQI+LFMvK8948o6MioVB7RLlbToei8lIZ5tKDiF/igeXC9H
BKDVsKqKewmAlrxodqGaaNzJLRDyp5rf1QMc3pujsrMCiOshr3gngW0tKtUq1ZnvRzERZzRW2HU/
YrPntyleElnJz+s91fJizbm62AiZO+WoZPj0Hm2e4UOVLcvr5ZKROVXzBfrb3bW4IpzNBn3n3/kM
KWgJLimCk4EBwlv241DelKyqskDkyVzT8Leo8woUfJOyjvmgqziXw+3BGm91EeeM1ONiv+D7uQgs
lOlDtuDpJuO1e/wOUBudljtyWSv3UCe/3f/sjcICTmir4SYF68fpOHAZSGOq3BGSoeYVDnDor5O8
OxETtl6siWnTB9hRbZ1K/+hNByb0X9iFVzYxIGtiK3tXX3cElI1MNIQEh5NoKaHDFZUVze0gEN/2
ypqBByKR139WvhFLbZeMmJWxHf9zy/ZBK32R4m1QGGNEFuix3tIL9wngSjdc209aDYHZT8yJDBz+
KE7u2SR82QdrxsftOuRHE4N2xi0TU3v3j5YuMFIRDIU9aISJzTvTPuQHovbSFvqN7lt7UW4tTy6m
hbIiP59qB733QqTe4P/HBdtJ+wh24lOn0cAtNN0TEKMXB/zloP5Iy1KBPcYvx7TemNtgnSNONT7f
ffFVZG9kNGG4hKEbBNkcFT4ogbzgzpk4amMxCFbATwuwTn7QFDWOweuG5XZXsFSPaMpK0OxGtfwZ
qQcSErY/Pn/yThVXpjtxjm0YA2LImRNDYenGN3AkgjAqP7Gp6/+sM1UwpYQ8gNG0EAkRwkgrQGqa
DK6hx3x9qek2KO3IP72RFQ65pv0ToPRWr0NExW8mas50j/lYS2dRMCnfb6qF7xmYxQs6jn1D4yAl
z/LZxxKpWkKuxlYbX35cruv51Yw+nuQTU9fuUDYegbbkgGGqV+xTKYXONNgGH9djQ8licWcDXZf9
NWLTazb3occKkwHqJ5WI4H4z4E1QaO3DnbOuCOWBKNFjqpki2u+tvOVtOURRtuyl6OsAqBsFGpAT
FA9IZJ7g3nvyiKXCI4icpED5HgczEwBEJpuiacrbv63XLSpyDwuihMUejpFo9a+gOCZCaH2fNb6k
v1Sg885ezBhH5F8w9SjN+ZqQvgK3Z8sHiuwNd8wlnLK/Yy0tsDcqCB23UQgsRVsA6j5K+3Ey+8W3
GBki/OjZS0ASiP/8M5/j86MZz8mmAn9nKkQ3RG3+Xbxl+yUoUACgj8bRU7QDl6Utga14H2abnAm4
McJHbuDt7TvO+tr/WyNBiBSqu9veJHs2jX8KZqJoM6soqCrE34Pr6F8p2U2b4VZzCLtRBBZ1q1GX
IXJ6bXP1OvDVeWM//c/kgazo0ysusSKZpSSyHl2xLjizXbHp0s/+QjDA60Qt2sTMFtx3FoyklBk3
21TZTKHRxXfP45/c2oJXQ8e1bVKNVqnba6yMe48/yiOQ0bCQpHAL4huVv1Q7NWXhtL1aCFlmtohS
n61VwQs8ByFWdR3zMgwVQAK3hqVumneA/0BSxIH0K/8sE5A1hgiIxipjgZ5bhHDZhV68skp6LyYZ
f62aF/OrXn5K9ZFyieBuHTivg2TTcV99A1/Y0N7RatRVkkH7TGS1yySCx2Rufd6EbYBfs/mzl7Ea
anU5wKrdGppRXgJfEbaTDIqCyeTITEFkUB6OGuAE9Hw+58mDqXvxZbKU77WMtjTBr7ZkX+jWW0I0
93daN/7805X2hLE+ljxm1ZjB850HosLkNETyTVzPbhCE5AeTlhNFEAL8LNaUor8mSrnK+pvSQu6Z
H4BCnMXLPSIolT3HdCPqrarBubUpd/LuSWF8fJ+2stsNbYn8DtNimnguGFu6rBIajha8D3eH+/ME
hyMVrUCnjBedzhS3ia2O7f/f+uN3wFU0pjkhin8tx2UrDXp1q8WJeCs5EViPwNt7pQgtXRcfC5Iw
okZ4mx5xM06WQxWbqV+c8lHZygbrQ9A0wsrqe8/9S51FeLvwr1yIZzRx0tTWvjgtvW0INN/w7lBS
AUFBachOZMQsczAA39B+xHCrofqKgGb0x/hqCMcOXsnqCIqvQAzjTI+/sXeizN6NUobbLf8pvtLa
gGMrQ7JcWFqTu+I99NDEb+ZGk9PaKQVIzHVIl+vlpqSeudOTQ/S6NmG3tTmL+twyCxpyCvSGDzkB
yL8qz7Upq2HIZ1oCJAESz62gppufMHKBVc2fFwWISs7buo6ey784JmEn9/45GFeVBi7a1DvA8FeE
MZAcVTyfXF/7ExWPRhYpKQP7F8AitEEVNMu45DXRAi9t5ZDoSJK+45AnR3czbk9reJUwCtQtRwHW
uJ786zAFLMQV0zM9Q544SiS1o+l3P5Uc02bDWsD7K0QbIDE2LV7BAFzcfD2QkDdOykpoRMHXHyUQ
i+zUha/ukrXmwl0bGKkmnqh5vX8QpwYFqbWhK0ZnAcekR7RgpaY4pUlfiXpPR8Jmxtmu6V2X+lBK
h6EzJeWWNY9G5N/JFnw6vcp/LEgMSnUXuEgcADmHOMYvyNTju1cqFH2V+dXjz5UlHOTUMgLgee6x
BSy2tfL5YE6Mq5U2JK8jnaKb06CKO312b+uz+xB9b4zIBeFlzSFWgUJqA1HEy8U3XApwh9mFcbNe
b0I+MVegjYX3fa9vUE25LD9kV1a2tjzMF5mj/dvkR4qFV0L+wicXwOyiVCPbcvDDGOxs+uB5AxUG
tFsH+iidnKyxOYzv42y9QARnCiDzhX8om1YDJqYhMzYgzBHCou04hf+Glmo10ECs/59Bfk4yBVMn
gYDa8wMybKeYApJ0C9PA8p/LGKOaWutvJl7xu6HNe5Arp2W0YD2HRw1JhOVCUV1Kj04Fu9gPDEUu
dfEXechxoWaiBpqjPTy6TP89hhGitl64zmlXFTwR57e9IVNvubHxnTKvcmvZO44bgnbx0zf4yaEF
V0YVbv/a59UUCgqQfDBIR9lfb1EudOUgSrdf4M3tDg0hutnG5eP5w9Q1rUHpPfo0/88POj8OilGH
HcfhgZLYAqtKF9DQvEjqzFUdhGJwrh7qruU2CjxtfQvCg6ZqxrkghIqA5qETnNyppBL8+AWh+zqx
AvjTLFc+BaH5juxwRi0a4oEO2EhZFFkaiVr29vbKqhlHP4gP5j15XsQhyQqsGmK+5ciMJyV7jayu
QO1JkwipObc6aDn/IbMyqDxJXBfgYHDJ2YqTLXukxoJjBsS7QtIHgxHTKeZHdsPOhSTbISrhPJDI
Rmy7LsWJTz+v08z8y4fT4XcS6sYq51OK3ezuGc9Yid7igz0/UF4ptAQxDKfFsoTL8/elNZwU54ms
GQPLbWPPbVwJFrq5jspm8Oha7ScSAXh7wDCxhACT1d0VRNlp/FSJTttFPJEK+88fYEl6Hu2rzeOn
4argtc2PVKXlstr+XnuQmdrTCjv66iEJT5q+9ZwOC1WoDF9WFHP5KEkO900qgLFDKYfow5kf2ouK
OopKtTAACB5h/j+v2ALmq2v5mytZxtdiMfHoppJf2mLvzi9pBdJSYzupcrSSYwIc3mVerEo4CwOw
+6azzL55031NpcG4xMNorh84LoJQMVM/FTX8R3TXMUTfVRwnI2GZzbWsHXYIUibcewrKRRo6tboS
jDuJGZRUPkBlslBPG12uRVZPrlD8Hz3zc4lYcVvTtKVQES2Q1vsprnNZoTMHNXmV94NfstSjnBT0
LV9RVFd6Tc6HJrZ3KmmMaKh/GhKKDVYVAuu/cazg2RU37ff3VbXXO6JrJ5lJrU7vXqulM4dEEhRl
F0IkattuujRNiMq/NABbxyHT9+Pti+bs5+ipWm0mE+kMq3SVW84KvDM3T7JwGU/IlnosZ9KWjdrI
sXqxQi4ryqP7a9zVWZW5CAUOwE8KSB0IFiXGNaxjjGFuTn1ch/hWR5OSJPesXx8orBMj0qXuaYS8
VCi1JAuOz0QQ0KBEBwii+zPdIwiiMklOX6JmJt3m2VoIxUeZ1mM9s4bHigPeaXZ3EPVnUjR4hYyA
6FndkVc/RZJ8tzzH5BLXjj9b3w/eqRABX5Crdzz3l+n8xmUKVzzyYqhQKY+xJYnc9wd7Rmr3HRKC
YrfLnD2t1Y9YjABRJ1N4RnUYia1+AQIWx45GBegzbTvNYo0z8/rWcyVmQRDQ3dJeWzmqYPomeiU9
xBm9eRviTYVNbl+fCuWMFiExuiVTy0Omqw6S9dMFicHH4x1P8yC8K/6aHBMkmsI2hDgpEm1Cq/X3
hMuyuy3o0vqqnurDmP0sR99p3XFwC+PWteQ0G5GoxCdvAHc5Ian6Nh3CcFsra0QDINfmuiEoXhdc
qbdexxBEVXl8WfAedcWLK2KR/Tc0UsFDfNN0wL42xGWP5DzG4pyD2nvS3C4eXxiyYLjfdG4m8CN5
BqvdNFgAzjC6r7hJrvS3cw8ZqOs9K7Caspf/BAL4cIL2Se3UAlSd/BahS56egl3mljB77UPB9Cr+
Toz5K3u5E4L51UtcKM17Sg+nks3yLpqEdXE9eYEwofBZ/xgFfeLbKViGtGsXXW/3xfF2sYJqIFsf
n8XepfzPQEbNUcG5t1DtoI1Bg/DY5w7OnV2Pvz8g0X0cHUxvRIqAlB4wYrGi3wIMb2KBFVMMKkCP
QRcT+O9C/14unKuig2yvGcbSrTd5ITgwGMKIzKE7Zkn3/83b6/abcrhH40afAqyM94ZdmPNcsO8y
hhziTxzCQUWgz7VGoPvOr7nLo4cCytyHIR6SrCIybjE0OsdmjWVVQVljx1gMcNTyPnlWkZEFYzK7
u5Z9NdHISKW+Vf4lRTr2NRSavZXmozeR70zeAZ/RH7w+3sXkbD8KG7s8f5E/lWAd7S7MywuXYuYt
Tow2LOhHU1h7v8B6LPnCwsJ3ZolxoPRXlKt3hot/caprEnDLqaRMD1I7RTCeAEphDYur58doSLzq
GR4VVV6ThwigqUM0Qz1opS7VymHOLGXx569kKTw/Of4o8GB3YfpSwOoY14rO3nisAiDEj5UFk3MB
dQaIruj8ThjoOokrBusxmktrkGz0pbciegzJY4HnLFduQxr/tgO+U9OMuKtywPfmC6lR96Sca6ZL
WE8oxqXpZi6S3vtPmNUeT78ycdt0BcsJAheh4Bk/0lYxHnXTNZoC4Xl9nEt9jimQoFtvywfj5QRe
r9+NSbj9OLZnm1gm+vR+mQN93S4pry1EkA3Ttr2v90SkPkYYtLAUwLbXaPozDaFohTRVtXa7H9ie
Z1aA5t7e09i1EKuYb93VLXaQ/QdxLoky+gE1WWjdzj/SD6EGs9vas1Hnx4s1aNxpNCjWeRCn1xa4
Bh7QR6chPG+7oTf/uqvBB3Van4lelYaP9NjufRnv9IuvE37zKJpKPwGm5UfTG5RNpoLWCXRA1cIQ
zuav5e+SLahoKXp/XlreNET3fovGbLaZKx94TMmQw+2eHcJwx7B4Qe5cqfFDKL1TYYMBgvE9l8Pn
QyTX5SfMOUaNZxTncJkhXQwa0nB3bnxPQB2YfE7DUtXVTqt8XBx12X985FeUcr/NjZL6xH8CE/92
8/fQk2SyO6Y5Yb6TBpfX5sclPtcLiF788jL8rQurTgQ4djEK/NUX1CAXdxGeEbneDslBvOYKF/a6
fv68JmBs0hQ5GnRAJBoyjKWUE96Dw7zxWFSEyhepxEzGViNCxTu3o0yXWZQeQvQmjd4AgDuqFXjR
Ejm3en3Rz9wfv2L4peapw4T3JIIpsWfQ5TEfAjcO9TRoG2VKIbannQxnhYkBplV9VodjZ9rawEHY
fr2w8nyzdDrNjFUvY3D8JkxWfx6Cpkaa0NyMTEGtChvVAQd0l2VAhQqG+2EViNTOwsR6E9gpri5u
AdJ5oU8ZFup6hTLxYd2LLxYO9woiUeScuQDFq3ERq2kGPZOSE4YvG4GvCPHEeh+xaU+/zB2OYksx
nXLxV62aiNptrZE5tOa6lvEskz/e++hyvKNbbuELq3lvMh4ihmosLDJbt9Jo9fCPrVQSmil2PjZi
l45XG6BMQrw7L2vk0jfDRlcPV9WOj00T+EI73T8gKZMQEuygsjiHVhL9q3xvDpLrBLTIwu2A1V4S
vBTA31GTC7oNjNbbOZwwthuIkNvCHFBRNk0mlmMJB63ZYu5+jdJsHFwpMAQZLD850KlPh0Eeives
aHpecfu7X+rrIqURzoc7GckFxysqZRbTKnDWmFo0+EsCr98CSMx34qH2/rqPi2HVLPPu+EMI2iTS
I0G9IUEpVznkkVmRxHHAgZBCYNpfMlEAG4LSELSWvlDHGzSLoNW+EgYyzhKGGLDmNznA5WJuwZ6t
pbqIOzy1OcCGAx1SM+vtkU5rKS3OcESkoAyuwEiSfrxJsLE37PscVVH/nd5brHRf3qr39bJ8Jmqk
zZKB7NSq06M0Q4DYl9sXzAYiYimGIMtj5hBCR1/l76owWjrvc9G+zgpEWv/LDrPK6yK7yc8n1+Rl
Aw01lUYuHSTY+Pdw2T+kAXfDXJHceRxUaoG3ayjV0BbdONGMqZvYn7/LmwkzV2dx1euXA9RlxJb1
8KeYAb+ujpRzsJc5beyAUjcibTkjcU4xnGXoAhRSAxUbeShtty3s3xlAgMYoUDkf0FN8xM+eJCEj
Wbs+dwYiWs7ZynUajwt1cRgCBYSbAUpC3BjEcULrh+khKID1IUh7vKwRB05qyn26dx+DjXCi8wvS
kMqfypbF+joLKEJsPLJmlWbTdU8Y3lIVQF4RdjG3EFdBhTcfvTF0kCcEsQsKMfYynyj57t9mhryv
utL2gTa4npTu5PtOOEFXnG0zXku/Q36xFoHB0eW2L1uOrnIMF8uvWH2kETPbFDJgUdzUBkZBpytD
94Jo/o3oYT/VFfD5zKoqMN+f+LOIyqZA8ugZxxsm0ulF03Cz5PARNDsniYQCujWHtfz0ZWjf3HSI
72+KYhHhrhSaH9U9zLWxsqvgPEOQphVuKelflA6Sq/W1nmnZfJbsCcmwnxcdJWaYps/wzatlmhLv
LizJQ6bnmROSURzhwNOz8b9l0hMcoeqIefNsfVfHeOcevz+X35me/7Cw+UODaTb3WKHQsW33mtle
aZ1evcm2Wb51LoqCO7DylFfddcaoAS1qYKlXvY+yjVmwyeOWWPP+u3E7joBTwim5IXsLE+2m9ctv
g2xDhKhcFLkUmj1oAq6zhmoRRxsK1RHNxBTQiKUv5gqouWOpKn9PGJH7ob9K4gHXt4e08rpumnC0
1bqEXlScXrVs2IKLJ6wbhcdnVGRBGQYqTgZ19B2B+SrUJyYZW3wWmVC1yTKcfy3SJBnHANypcO/s
pvPfduUGvdbam8D6SoNh5LYz4d6CimGqMHdLJ7nh45FxqZO3q8bhqT88VeaEjKJiftCz6paLxn8N
yvCtI92xmMmJ76DDT26UndWrLa2ZoObnJHC2njQIe8Ryvw+HRpp06mMjoNDUld1P4l/NA6guK3m4
HdqYdSXyKB2mlIGh4kEd564jzLPpvN9C6zJL+Z4RN4NgKdfX5DfjMtTf/gW+SftXIZ506Wo20DVK
t4Oirjg7cMnUnBHuXsMb9UFj0SbXm1QtNanYrOFDmTxtTnJ7kQloFTD70uT+gF4wdcqPaECjHyEW
/XeXUJm7T6/ecqZ9vMw5tLVFCVNT0j+Geaa1ANvdl17v4kxlx0Lq0LOSP5vS7n2re+vPOv/ya/tm
3gJNPmb91g098w1/NnXVNErOTSg/qh6DtN7dqSgp4yBR2UUzZftSlGmlexVSkcGmGJINF3NEkSs8
xLzElzr0wctQr0GDpiK47MaS63KvafP+YeGhL4PP50acG2EbWnYje6BcNWux9LzfZmHMSjgpEaP3
FDo0hyiB3tb7QfPcTyiQNba4+qJ4eur6kmjNML9guU+TyzDE2DiqZhYaZrVEdKTQbie/1j6IQED4
JSzy8yuL1O91msDfydrzZG7F2hX6VCOF0hPfyhKr4+9sC6hQ6Yr9rZNypxpv0leTGupItitzYwBZ
NgUkpcWknWcxIMGE+5AKf5xEjdBfm1tHdCfO+vkg4ANXGgevyM06a0Vm3Ei9e/VIBGHSKxdMbLhs
uI32V01Rhpq5xKx2Zg0wOc6txxLKovd4YK5dghiFn0WZGhfb1X5/leFNHtr1BdIbhbxQlbo8ttCU
MFtEYCNhFHewhgzF+X9QzKRuqV9DC7yBNtp3hZewIh+YCOTXrOVnpVZtNukoHxaGYFtDsbToPaW+
c6m//ObsDnUFf86TWF0Hf3HZegeqWhLpjctzJCztzeXYs5PJkg0LGt2NVJsLCzP18M+Ka22omH8l
qeZc5LyZHpyniIBsJsqrLFpbXLzIT2BI94E2MT2XyFY5O6xpzcwtbU7eAGfcYpSuD0XCwx3qJlZr
efYIiGZlz9q1+TIb5nFZf02QXtD6VNRC7SIfL6OzSEzEUAFlbm94ajhPxI3+/rU6NZds2N1zEtVf
eJMGw0lsDxUKfHA8soUH0aHyTM3zb7ZRO9UhxRZnOTDN5+RbVwvM00xfpS1qKLVUw1rrBFoDt52k
DAGxucG5sE4fw8jn6yzfC8ALWlMAQrwRGO0zKC7iUlzS22kkQkwJmh/3MWQszFdhP3K5EiZ/itmy
C71iSL5eVVQVBrK02Idtq82+rfJmmfr+YHak6niB5duWyWkpU0tReHjghgp4ovZ0no0BXFDyAqxg
51S4B5PIeP86CoymSkg1fbE3dMhKkW7Th1noku1ut0dLgdrdRtfIM7XeP0C6ch9TCbAiKu69Kpka
8LD6AQ/8sE4W4qWBx6E5xDPY3DO/F5fGfWhRs5royC85YlhjaXBd7pjcQ4bRZ3bP3gjH461IaojM
z3oNe67j6+oEVNNznCINolSwDQ//SvJAth4ovlRQ4pjtGw7aHn05Tmh6V+To3TRXNHbJFRU24rg4
c2Mua9KpsWNAypaHRjWCx31tRvX66EhMqWlIBFjHaBgQvYuM+7caSvdugWHvFaZpAleYuaaBKvcz
ojEaVtwyaLGkWtx65MhjFlf5lxJ42orvBpL2NApHyggUm73ldScg+nKfFT8KMRY9vr1nxyZ3ElaR
Rm7397xx+viNbE7OQcq1Nx59TwAsruY+6dGc6Qx5SNQYgOUyLWe7et2JDqNNDokKUnMhPLlTI0ts
Fk077QPZOdjOAcgLBxuu4t30CMaXGA9RF5sFGKt3cR5U69rGx8IbU2HZ0RYMDfXWhPD/Rs7jxrr5
OwwZZa7wnWvJsXPLVCHnKUYRUH76dikMgzBBxKTsz5K0z5NwWouMjNp0FKoVRhOqGvzBWtGZziuw
lvQEUZW7870VNmBL9ZUNS9/QnLLpImTiaNj2qrsHB2FFsMdPk2L7UFUwvgmmz3fuA00ujTGX37Jw
M8YZ5nNHsb5wnumLWhfQlUW4PHrAfh/8WdQuDKq0/1y7+SFrE0/rYR1dLBXsMCuTFak5Nm5y34ld
q3XJOHWxsWeNAmJ2BoDoNi4nyf3IsAzzhfOu8wmmLRpNZvF9iY3zLNqLIJN/8C+5K0VBcnq33Dws
wT4TchiNzchWslRo1i5P9H4ymfrTeRqH1jZNoocNHeb8ttAuRkt5rE5quA/7HDq2HFy99IshxwnK
RYm7RhNmG2CgSnIfDBklZQwGlgtlGMRQRTrWy3l240uySf2iY/86P97Yghi8INBs5g5CNCR+biVq
7sJUsAMRoekt54G9Qt3BE/9Fh54ynBb3Yv87z2Os7w0VyIqnTd7i/rceiGFaJZD/UoQ9Y+INFMaK
dzHbleh9lEnqepw3lic9vfFhb43/FYss+8mreeaQBjKLUf0Y9bptZWH69rr+N+iPNLOQfj+N4Gzq
NyM88rn4P843wvXJMbO+Fj2N69gPDWrg7xiYSVUsN8pym99CSJq+XtIjxkacnLs9EFCsG83hhdwv
UcN10qNm7ndYVqKB4Lx+94io6ZYbzdNgQ+STtiqhYCIKXyl6BjbNQRC7csm12hKLY+2D2Qi33d1k
JOcxDNrvwY47mGfqXByP/BBbpKk8Rw9TgJ46qOBfggONzpfxcv7QouIlL3x5Ssxj6EdLSA5/XXiu
QSujW74n1GL8S9hLqEK0zOAPe+D8dJaawKXOZONAmusLjurPREVIhljAD8pvrvnq8Gcxu/+PXAn3
sPzuNsVGXj7WNkqqKf6sI5Ex47DQ6eJN+iOjm3MJ+kM1XHNiVASsrps+H9gubLuFwvmU5qDQ+RV1
YCvxOAQmmqOGsuCj98BcK0osTlBqGcfNfA9QV2wtsHTGx9QPSGlcoWJtj+V4yrC90iM5NltIsQkA
09YRKjUy3hhj8G5/3196bI2h1RmjnCc9dlaJSLWv47oPy70RaDazr4sLDRGBBuMV12zJk67/PUdg
w6F5IQTdHJ57QJDb+LA2TVchbJHlbXQDU3T1bzgkNJ2Ruh5MvfrFJL5+IjLXdabk7l0sU9pClg/d
1l3uzfAV+2ZaiI/PR7rh8frleP6bKst9TwWBaNEPHYzlenfm7bcA1JL0eplJZEccCcTE8DUjCV+q
7DX8+ZwEEcXlVtYmCtJf93jIePMlgs9Usw+Yb0xRCvAgyHV5SLrEDqYJ1KC1CcL3/UMD1FOcgSg0
4xNomRB87iAeFkn/a/Pe4McjwKVOVPnVNmf8LmBWL2vB+A163O02pnKnfOzALNbiFLqE2/4ZDs9B
y3jaNwKAx9nu9E7NSwhrFqFapQfKUpaJWsXheGLNETxNWOhJnSRQtjzQeG+wR+zeZ25dcfH6CPmB
ybOr4x/oSygS5WrfVA8BtqyQiqCxOiVVpnyJMYFK6R6x//fcC6GozUTtZaG6OZWdwstdfn1/faJo
216UtJ2r2ert60dFY1Bnx7phFwg/WGoQ588+bQFy/WAQ77lr3INaoFjcFB8g6ZMwbGWbBNf5mC3a
1sil++I/0S0g/D6sMpO6e66OgOlQbNnJbMUmA4mxYmqizB1jw1UwWMm8jMt/i0DA5ccprR91vDtl
mX8BF/3++s94uTEIMV6BkIqM07iLuEZkvwEaHmGNPc3K1MBGSlwiXNbpLREp7wFlnfmzFaY5l+LD
h7XPVFo9o/nvt4d8ENJUPCzjnhppbc3rXg60z3IfTFAz1ScBrh0vWvVWo9M33+zClJtvYpKNc2Zw
7AxIxe65BY2KYFeRc3w/MsWDYMQVY6ejDyT8hUdhznVo6ONVSAX7L6gDRnwa5bX47urARqsdkZ2w
nMiAWRlwBgVBoQT/cl9g7g2ZaF1AVDQK7SV84uOLlWeaUI4jHVx4SO7vGVVrVWo84F1tn3fAAG7p
fNTu504Iu7LAMZ8w9n9JY2aXiupK5HhXjCuNusG76nO3TIxCDZBtjGnN2QwQQkKO86btm6cTeEAf
j9LykH2bKiN7V+3ENvdc5cPR3lDWU94yFq04hNXEvDltBESri5iWHF2qwzLis8rHvwTC2XXsiaB4
ywVHxRgY4JK6/aNHomd7qydlhQsjSFrvyYWbi3QoYKwlbNo+xZb4S8tgNYvD80DopfAKesQZEjrC
vPvgHEJ20g9VH3pTY/dvIlnUFnaTCwpVsiOojOQoHy9uVyv6J6liHTnoqDPgveOsu3B3LV+f/rk2
gJ7Ar/+MIkjCEQ6pjT4lYvs4fEu7OKRsMX8XgCul3ykNPtpihW3+qPKWyo70hp9rP2lNaZrUR0Mq
rX6A9nsLoy7ilZoxFP1Qbi4XCDcDRwqc+vbd4Jm/KNS/XXAmXEcoUAcxKjUG7e92HBJQpEDf+geW
vpd5kFSyWv4Cb3uOiJzlQS0VMJEhqB0l7hSF8IHt8XTuFh/iFmmLC7gxeA7YYsqgYNROIyQ6lbqc
6updLY1q9G42qo+NSzR5FJjZ5Wpy4qJRwlhRencvs4pkpB9bW1wOtNYX1Do1+etBtO43FYiEil1S
CYeNdP4IZ+zwqsrtcd94C+Huyc7rRExXmIfhpMw7HpkgN4ZbD9yBMgcFfJi9nwYAPjEEEyuCpeUF
i9xsAFBavLS65BnKeKgjfTOD+k/bjRWW1DkpaMLRYbbspbSS+Vblq247x3ai0RWvcpEG7FrNcaQU
34nvjlYXxZCLm24oDku2O0mnif/ChPKZvFzcnjtsKG+GvsuXWwUzwdp4z7GVtylx56kE/+wNTxwV
mHPVDPLK/YWehJzvz+pSzrJ1zXxsKg3PhMFqYsnzfDrVl/dCUwUDKm48NYtD4MTR5m3DTba2uCd1
W9Pl2oAHWfryj8UgjKX5RcmF+niUWKo55Y6L9D0Sb6MGo7hkljNCVCw65iya2OxUns1EhgwPPswc
hSmxm47ycs6HZHywxqF0YowCtNOT2/t8DPYyL4vEU3qO7LyoE0ZDSROvIbjAHNiO8v727oEHgKGy
dnV179RQX01hjeJ9K6A+Wwq+B9Jwm1ofI8VvOzL5DboVufQIh07gO2lsIXErga/U5f/BelHkBGdC
HWiidZeRFCOljIOP6lG44KrH6zOupBLfFZy3pS2LwgpAVAfDxYI/tw5GMQyuzoIrZBBaIsxc6p6G
7poIG6b8InnEWRbwZN1lp4Ni7wgB2H0w57Xg3sKQ2H9Oi6i52GHDAeYukraP/OEpKINUraQOZuKg
xK/hfbwnCKPJGzpNuFg5mDicXSHn4gCGkQCdN4qLHOZnFs/FQC5I01EXp7Rs71uAbPbJ2HxMgmHA
43U3HMStn/XlkCLJ9Pfty6DXOMY2a1omwUx1mp2zD6R+F6eI/XPyQvvcTsFV08uh3Ta9y7itLnk7
dECWDMRU3YLirEwlEHBlC+kLqt7NsfNN/hivnzVJHLHSJTmtmBqebbSDCZtsSdHeRMtRmd0PFn/v
8UJZptIx/TgJV/dqnbhrlNT4kAKF+OqWD5EADa1yv7x65/wS+mdNjuBckgywvDzCuqthbajdW4Rt
LC81im4rY7SRXBDOS21SGmX+DEuikq5ysxOrNfofCB8x5IXXDOpOLfMamZcfrG3DubkY7Fot7UfW
0LQzLxau/7j66q2erpUI+Nx13uUnAN+mg3ik3QeVQTqwYzNrbdUxn9BOGCQUXo4KuFERT0M2vB2p
2uAMLI+qAJiLUHbnYPXnuWnMqCL1h1W3Hzllh16DeiKlZ+qQAUa7R5jtd4pW1AtwJM5Y1WbfK3HK
r9fDN2KQuzgiVghVdQ2gGjcZazZjw1n3YuJo5iBKVc0dwKZcRVMSNpvMNDdv5KQearaC4ustIyKq
TyO8BMo06xNXhpntic5mJe6yAZi7W7uekLjlNHQKVc31emEToXbKF9y2vcLgls/MMTgCKp0Bh8t5
DrHr8G893ULTvvb94NqfDi0aAJvrgGNCxm8xEkwlFpXX+bQCEY942VY2r17zQ/yCxdkGyCd6lIat
8yOq444YFpnaMFyx7f2vtc+uR8aEmvscxh91ufgHYdFpIiQUbFN3Bwi6mXrvpxGZ67YE684z2bra
K8q/NEskAb4jvGmnpZde7udLfM5EWn2OgnKxw4S/zHW6MsyWom/g/EQb4z6Z31umS8i7n8S9BN+o
CzOWXLV0+78ixi0CLJLILB5GLCN2rzjvLCHRiCQXzSv3QN/Uxe+rtLZ90jIreRaQk4vGZ1C2ySjj
xAxPtaZIIAPh5biPu5pSOxfF17qLHTNJTsuE2tcHeQuiVR4y0aUiwxepSkdCdNizwBYrDjO2RuzF
RptpaAfhIUEl/ijFsyrCMQfs7Jrgg65D5XgRWk0ieiPmiykqq7MhpWsU1M39/bp49UNvRgYs6LWI
3dNB3TEv8yQl2aQuJfNQqVFYUgW1zpp2Zc67DYVCiclfJQtrAgLgVpQiDS+Me8Q0fmRZPhFQ9+7M
shVygq6OsI5JVfDLdQ3aseAtgVfyHv+fS8CkEGLvWdpsPHtfL2OnOouRJGSw51vmb8T24excuEpH
kn9K9KzovHClNdzBQIF7J1KCOKXfhN+pHmpLR87jHCy2ongrO3A3w11fJj4XJzxCeH+AgScxmSAK
v9tL6qpVu/7xAYspTmgxM+vNxBFuW80uEj6eI4fCr5YuMdcsCgrYsIpZnFhO8vEB35lDdISimWgE
eA9SKHdijykFB4eTTIWhCIpQyiiSdd5MC4yZfQYDIVtOWHf6BBGgFc+ZQMhWbp9yXoqDwtdHtEgt
oRkAmm70iKHhYggn86foJoBRDvcXfbSf35m6njFyNaInvhdJxdK6CqpsaaRVN3TviKaC9DmDjZ7F
E+ObndNrl76edIVgG74QWiXAEGlcn7k5E1+tZwBxwFzj+CXdUa2sOuD+mvOVeJykw1lOq4BOcY4u
a2RIku85aA1t+KvZqmUBNxv/xlPC2X7BqspDOXZQ4ePgsilUEmWEBpvEwvHtA7NntiRqoFc7rHsX
526+MI1bg/1FpuzoSui3RZszAPhebl0J3XTVtdALDid0jZwMK6NWULJLXtaME46no/jWIIM/Olsu
Z6pEnQLPC9ouviVPMEbngJwNJIhamRNhzvUQ0LJH+eMTUXFSY5pysZqqd/FXjkyhlfCjkOT0bXs3
B6+1Fab7zd4qt4nMMeB0Ze5DJRLdzEcgwi7alUUg6h8Al1NRpUX19mk/2ZJz2gjp8axQJT2PHLFL
kMbSP3F/rg2OMqiDFtTjQruUCtyn0dxqk4ec7yvcr2GHgF+PI5ANr2lxwCuY1VuSXc0MXsO9SQSA
0//J/V1/Z9nB/UMxDNpkNTZ8kMVDT3EXwbsLcJmYff6cAUjQTie4neogYU1mRlz4j3UebfKbbRK8
7R00oeRUkGfhwAWG2uxR54vfOWF3Wr0Vjrjf9qf+psqiG+qnm/RlrUWRncIsAbTtFmPTzdftlcN+
WcBfrWf8zO16NIcaLj3AZYl2fJbbYeBd/BGuGdo52SL2axhX2LbhHqgZriBraz5lXbpTb3UdfRUm
yNmoieHrUSvbNZ1pyKzEYFvSlQHGszGBefmx+EjoL0+qv1eDoByml5WhNH4ikpLYPDh1bC82EIe1
KW1vD+GsIU18vzv8KLz3t3+flsPwahIwGwONZ8PSQ4Qx/s0JiHoTt7NHNvoAG0U67IZDqMIscASe
GBmaDlno01Sfquek0mhxHL8eNINX4bXk6C6h+rO3ggPHaa7N3ReD8YbZ/1l9uI83ekXDjpIKfnma
k0qAPVTFKD87SdPeNy4DgcqqsJeJw3wZmqHRRjKeuvh3AmoIZvVH+fTsdZybx/RrjMgoYIkUu6ui
ejrkkWPDsidLkRk1PF6qUfLCxTV+dvaoSDP4CgZKP8KuDv7KXTJ3CCFeyMIS1I/zLTfKeEgioQ2b
V2bmnwTtubVl1peUX41GIQE9x3fs5ydWx0p61/2qASd1yrihqMuQ7opAFFiHbDxGCrogPni93tPZ
dhoWu9koy4sXpEZb8KqTgDIoxGJd3NfvbUskJ6w24dLegjdPapk5/qlqK1GPt96MWwnX8zJDfPis
YfcClPlPXDB4VdpO9AYsy4Gp7cI/SyLShh2Li/i9I1uQx162mxCIfGbbAajdfwpmVP1HErC6dBlH
SRKuq70f2sTKMFQoPzjUCJIO3EtyfEh85Uns+pmt2QUa7prt1pnH4aLZAy0EHgiC7pUO5mdb+1mW
rLRTI3gLAVXITPt2jGkv+Z16AqetJCuIv3xb28T5Mzl4MYhIFojcZiKpec3gxOq1bxRThfsou7Ir
ma19YEduKeOqBQ3qtuOrLUNSkNEdFqY43eYSVlee5fNUpritEcfGmbeaM5zZDqTQjusv4ZfnUgyn
bd4B8wHvU2KoW1TDhbf5NfslzallW6devvlurOzE5Ma3RWKnUbc0MFba9tNBZ+3vBAjdcoNmc2K8
sU2O3MSKTlnkvt2vk/dlewewv0tr86pDgk1Wg7mS7TxXA14gMXsxkFY+zDPKF4w4v3JTbmZughWf
7MZse6h6zEM4mDqIhU1Jk1I7RXXoDVHbr/8Mj1p1WtndJ2yTJozC4UG/V+gQAY9/gkQen+MoVK11
L5GaKaQSlqFdALoawInXTbXllJqS75cUi4kO3hxGjeA+mPeyAA9qdkxXwRJMbcXhknjMQ2JzIfpp
zdXMqsY5IhWcobHs29aivwhArGxVavm2RaKkpu7/h4kkBbC6eHV8h4Qb+rmOFb17vl9c4tYNDe7p
WFuD4/MwgmkNrGmTrR3hYsiVzUP/uLveHjgSbGQkQM3OM+JJ2Kvs8pWKcYm+pKb8ooMT9xXsFO6t
dHjR/TGWlp9i8bX/yHSbt5v7GuA2VzqVCfXoKRQoy3gyvAFKwumdDAKZyQ9445GJpJhRyLi52PMe
LodAb9wf3RtfPDKt4DEgkXd87T9+zxpMggNYSy5hbtHsNCkvYWvd11wHRbZl1VvojJlNEVmDEmJi
FLOImDEAnISsCFNAfpTwBCsV31k88PYfne9jP/YMH0UruLaeDsNXJ8QfxV30eDp0HEJz4VdV7MU5
4BFkjLoeby03da3DOEgQygXRulKXQvPhI+Wp3bJUyUhrux5BhavrftRqmPmXSeSUCVH9V73xgqOB
5FDz2wzP7YmU952BTt/b0ZMpmTZub0B1g+Lq2sAp7CbBjElqZqrxYSbz7jFfGcTb5qrMyeHkVo/6
qaZ/LRvLlwz6dEGD37F36i3yw1t6qrbZZE/BsTTJiW4lBIeTbH1SCY2KDqOTPB8rW3Wm5odg36cS
ygOHVgHKo+h5rqEN3cAO80z+RBBeJhvc8+Zsha6yczFI3eHi9LUcB+bEZ7t81EoQ/0WXRPqQ5OdP
JNxAF4T6CGp+epdW+5wL6gdgHqSpVD3n/F64p8GZ9FlXi61QeFDA4DORryaryZWqfghXfF0fQddO
eEouJaYL7SiAz3vQFmr4CJV69QIRbVlNDALazTdIyjA6vcv6gUlqqYbkBcPc96QmLM8F5DwVjC23
HYEU3lx98aDlBjOIlsQ0jtFVL6B6Xu5Dixx3nEPZXAkWbgpZkLhWxo/xuX6pLmcvPPvX5JLm9CA2
gzVPPhEBxP/be4iOZM36Zcun1jHFr46QOZWFhI1/74/zxnxVCYerXuoUYrlDpZsA5XTc9UIMZ4c2
Q5VHSeWNxLpEFKPb4bONlhg9PKU5gzpKF3w6pGwjZigKoCzA411ZtdUr2gtHfdMTxbX+RPBPPGWa
oU/NeiS92jqsOXDR2ra8EYMemk6uAOObDE74i24bmxgNcpfFXmRT/NyarDIDfmPty58gtjvsYttv
FQYev2VzO5f1F8Avlq7nfKl65U+V97U5BK2OCbFrQZ30nSpmieAkFClOPSTH86ZxyRfUUJUFduSz
SFd3kRb1mjtTiQIPg31um6hRCA+XCYumEMYXWuB/ZNjXgreqqPdHM83EER6k5niOUN8e7vI02FXH
HGGVsT7P9RuqD+m9gnl6wvQoliPevGMYn+eeknTwQZL9Deq8VxCemejtxKCZRxMyhqtCQj3wdAOr
CMR7sz5eQQfI+9llyIzGDL3fpDwEXsteqxlzkH5cv+k5fxSmEgeX+lRcZ6Kx4VI7OFfpgcSHy3UB
SG0QZLbdBu+qiK7Yb+vUaWqyb3XjHLisH7BoQoIuykF4s3nMbLqY/8pzNAO28mlNtpPYayN6YRzy
/Vq4wbYogAvKiAEAr0GBefPnh93S9YveXPnFREjqQOleDs8GnNCq8+9VbXnC0r8mzW7OM4Q/ci0l
+71mOjOxUTTan9/qs0b0YQptxm0htPadlA32XdvhQw8HEzXfs0skubddPpLum6iD4JmIcEsQVfic
eZJ8I7nDQ+X2QQOuLiAUg/j/5bOn1PVn+DuhkQjXYik9+lWKVAagDdqA567WsV1BppxuBZJDOsJb
i+l14nUXHAVQaEv6ScDWD1esWxkP3X0fMW72odZjFkMOqWpsEdvVE/oojB+EbCC1NM+AIhhf9fn5
0xF6PTS1M7DmD3LUUxkTjEbs7E5m9mcs7UFn0RCZ7KJfgj2pGE6HlykdVGd0wXy0lqHyLwt8Ck03
q7vBSm15XXbAFmHHY1ryA3Syny01v3q7XaOHcvAIrFI8IUibICXQ5t7q6bhFlZS8D2Zmi+G7RNhr
ALCIde++KQuxZXQK4r9kzcKTIv7ZVPtRj4kbIzGuPSDFREZdnl9MXCFQKvNuCb1xNitawtqSoixl
hVI2GsMnM2La0UGsgwuj1md3VVIwmO5HkW51ChFnUZTXQ+uVr+jjwsN6ka7NZXALeKFR5cNFn+Fs
iUq8X7/DlwcqkKSgBov4UY4Jz74mZclZmUySKcq2Xs1C2AID6UJrNbcLYJ/VMcmE38JNCmNgQP/d
FTyxoWSfJjJp/WfZg3RCXXvlSZ9irNOJZjPpDgmojz0EbAbEbhUvYv/Q9i2MSpz9DwHVmM02G4wu
rQG5Z4Z2jg52r6xnQ0J6+xa2Ffrz4wNKQEh3iwJpJGAD99Zsc84YdodftBd3Ifzwnew+ybdKTcqJ
Oaj8BlW9HWVjfNIZt+JAOQmunpRLiFCkYzLLMmPCWp7s29BtKDcAaJhle9vvgNS3L1ifek7f5q9l
99gdFyAoiuC8HLef0U3akP4AF1vqjmaisz/JL5/27j0Xqwn1fRuxd/RufVmKLLR6nP20TIeO/nbz
uZuWHJERmD4HGpaG6QnDkm/iZGxp8IHUMyvcOkc0Jl6QnD4mQllXr0rlfS4+n4ZcSni3h4iF4NZw
130d/zJEt7AWN0UDbWkWe7Z/h3LTaZqDEgNcdwIVHXmFm09ihfSbnBxYWG6gu1AMh72JF6tv0iLG
BcYJo9OmQ4Vfoln293Gpk0zndj48RC+os+u6XF3aJTJr2yaRWxyXzTRyWKmyxHuY6t6gju/tRtTs
8pMiH45dtDaBBmXrocUUssxlUvFFtIZm5UBqTaXdAPsp1kMzCHvWA+WNs8sq2mVwTiBQ4J0kiK//
BUUVWhlZXgTjpJchNo8sQXfHO+gv/TOYdD4F8q86uzudsCpuOuNJ8KVAQHcnA0+F5eJ8tTv5PVNw
UJtpuPuQQEFoHIQ7WuFM/gpOPBp67rd0ZUAwsnXHaYXRe8Q9rON86+gqY8uuzlHtvS4ypuRXzzNA
7x4Pf+MWJqCYpTp9JmTViiVDlX9rZdHsHG79MY71b0JCzCVAIJKDGbwgvieHdP2yoOIqNgpr3Vmf
CPgb5GWd4Z7Qf585dcesiEBvGaTIJ34k5rEZlssTCv4Hms6DNCbP4qJtksEUZjfEiPk9qWQACuht
nAJep3mF5oLCyCDfB65WQyLZhXSNZh0diPfFN2qwUA8ffLELSUBfyQaxj0cwX9BZryzqYIfVQvPQ
D2zXZXm6T/QUmwJBLeGlU594kVwFdD41ST5u2dfQ20d0xl6mtOPesvYQU9XbB4tgoXCuzgs7Fdc3
QOJJ0LZ6D0/yFFXdRKhwrOSXxDm13S3W86OhLe2GtySQkiDIvjHI//mmZePQI+2qzsNw8Jw8827A
3rSENt3mMYx8tj/v7VR6+WRXhRET42X1BWpbIfQp/HlB0dRgJRwtpbr2slNFR/IiADARSqO85qaG
a+IxiPXe1t74WxYI+j0GjSEQ/BAUErTeqaT3VsLtwZ0TLImKucxsLmDBUOkaKwyP6pqEbT20cIfg
k+jJfnDdTfRFI8qS6Q2KNEC2TToiCOakhFW75OWhZYvbUeGXYQVD5zzqJaDRmAUNG+rdvdnAc5RZ
9o7aIPfR9Fkd93lZTezZuzQodU+2vo0GgP1tbeVczUzSZiGQ/bwhXK7LIPTVMJA2RMfW5ZtvF21c
JYKrmXqR96NCjYa4LrfW2hGqc0DrICIrIeDrT3uHfnarhuHi4hMVeZThiSHG4lm1cemdtYPuyv9Y
GkNrEQH8gPgpLaXCHI8lRtzF8RBzu9FUH2DpUqngy0gIRI+ZtGDA/2kbcD744bDw353nQdjq6iRe
O9yTDFhtzdXyudxwrIx5YWaEc9QbF2FsTmkHy46pbekPJo8h1fequEiv9g5ng517jD2LHp7WDua3
swjyfdV8Z5qddz2vojR1i1UWVUS64eslG9i6gfLUUVuxp46SA4fqjpoOCOvlFGV0RQTXnukCUfX3
vkzqrN4nSwrtXw6bDRcwgBzKeIcIOzqjoKZXtFnDoXk0OkdGizGfT3DnkkHGGY7WWEadQRIElKcr
vebjBv0NkooqpgXyJOLmBVsAdKDdCwD9qJc71BpO47gKLNvnziXmeExK5QoD94ROGY9sdGQ+1H0C
MzdDjhl1hU45vbVfk0R0VCrcrM5aPwBdpFK4OnZl9fm1eEF4ylif2MVXseRpijai4MW+EDEVXPdl
ciV+PJ5lahZtEyBJi9ZN8+LpVp5fIv96q0g+TScPNPyXtyhtx0gT3MWB5KIpgNUScfyPbbYDM2Nx
J+CNay4OJONDw6t44S67hcOYiOWTXo61gkptAEwc6g1Ux+xf28+OHaCkzOpLanYii1T3M5iON4BT
ePNBtgFNAnmyuEhUN/TA0xivF+OD+H+iG39BuWONCJbkDyT7zPyH9SH//jfvgtsNi/8rR9DsOiMi
Qfmv9uvMQXNer9NeNtu0kKD7JoUEFff5vjOwWsQ0+O4tLt/i7lf9Ja4GNOa4ygQCbQCI7eEgWvxM
y4wWoEn11Wu8n1vC904ljClI47pXRsEx8sbRUPMoklDsjj3XWc1jQFHO9eTmRZSdEG2iyDLxK+8T
LdyCt2K3Pe6lpIcYNo96gb1udjkfFUBUTZut7ujM9ldiWagvYMB5qGtHzxe4/gLtY31T3gWYtki9
/8d6ito1RLXiFPnp36d+S4CC3WWOL6b3Fwf7BmyvsDSZp+sIhs5B9pB3kM0xyL8Of7TGwUuKP0sH
YBQVGYUv44qxhSE+s3Wu1ef3Eyh/c/tam79gOtR2t5ifEvzQ6t3qh16J664YryiisUv77yR/pwh8
DZqxFDKPAKbsV+0t+g+AeJDRpo68gKyMkLA9urQsDQ4rReTZeQzMRNDvxmx9iUiFvKaxj1MsalKo
RqOGicft9g49628nl32KHwyg2cYDRO5PU7GNn4q1j4tMNCj2IPxNciSr9d1QhK2KfzMy7+QYJmQH
JQnLOZnJ9GcGadQ7jWIru/2DMA05Db/mrnp5lN/QNk26waCGRMuiJztFX0k6reMzK1buMfqo/Vc7
Ouj8G+mPmmmszUAoE86aRCl7qfd1V2Xgq1HFIkfG65ezkt0VWwI6hxIrSH1SrVib/4TicWGJ3IgY
42fMqrSlVCVLA1vbxc1r4/ROHDyqr0EqoVy/khsDcdeFuMI1BkceLhexwXCm45GxfqNyX5YTEzOh
YbqS+RgjIlPn1p7BDbDkkUhDzU6vcI9cZf9qRArb/2ENEO3JKyJDSbOlJmgrlww6h6MjF6BQX6zT
JBAMBcWcnyU/GsA9JlNlYrd/280uxmGAZMzDBAP7/LDJ2gjCnMR8rwotYzmaRWdxsJtbmPTYoYDg
Jt3CmwcsW1IDPd832Ls+PCNFja9D6YZPSUT/TXjy4ajjSeXWOX0Qk0SJGBjSqEoAb2992ObU8ChJ
sRhYZjiRrClVSNd0chelMyolhW8FCBBtzXTaSg5la3jDez1MxJ8jQOYZsh5XNv2jdFY3TLH4ZGRG
tTordh4t5/WosOXltY3GvtBUU8ovTPrKvwfiqC29zurHaWkCIuoDi6wDBJDt3PVItY02W6uC1DNH
FU26O0jcjbPucDf99qrg881yjieW7DLSW4m/dosZyuUB/lvkSfDSHa1z+N62kq+8kPo78dDCwVs9
xRpZ3TmY9Dp59FbUOv/LJfklhCgMShafb3SaOLVvQmTDfotBCxvXHpq9sPRX7vCK2jEN9U0oUcfe
rB39d2YKWeR0sU+v8IbhzSgTycAXgoZ0cn7UK2tX9VhZOXY82qEOjW1pnGKihxytG8XGnfgJcEvz
cAW3J3H4drnF4Pel0H6daQjSgYSw6pHfddixh/VLyPaBU+xfgsI5opyycHv4K3w2+vOgSNDz5iL0
bWI3GBY5IG/3dgTRU3C5rvGslyzHWD2vyObNeR0QbUh3a8mbEOpCg1W8SKg4mJ2YxfQXPWQDsEvq
GoWmdQ6eThjXlMYyxhMzWlTD26wQIJHsSnxHGdM27faobqZA8XU/aGRxtrlb7yJVxnhGhtlt+AWr
SbLqstCViqpzNHB1114oIovTBnMoetwgbwVohWAOKFbW8dsuzcofDDM8gPUgvqkgyZHTn+AI/OHv
HEvLz/2kplQj4hcwsWxRm6802ZRwus5uVCgKD++moO0B4niLX/a/FDHancLFrYveAiqq3SNTSv8r
S3PZEX7GWw4T5CcBK7HF8dAhLP+vWBe0vnIu/Uw4b1JHnCMMxUHclD0I4g0M+Qpliggr1CJZB/31
jbglWghp9cVaOS+cGLHjqjHBmoCM9YEUlC3NIuVN+tdtIZJLlCe4b2Kh/tfLYdMg5HT+36LRKtsy
wV+Ib7EKS7YUphaUuqnIcTIOO6NGZxovp9tFf91uf5XMUrCL2ifepykhOJVp+x975fn8iHzuf2CH
6DZegTScAq6FQD/zdQP5BbDz8FbFrREXuXrsmRhmIxcPo2EpP+ISUh8bmh7/F+5A/uZX3QHQe3G9
IOzHn7cSjp3bBSHRo24PLrAQRUF0G9wpJpD7lxvzPMykjRSthRQxPzLZTVahFR+drrgwreRUu0Iu
8N7oGuu7dEAZRKpLsEPs55zcvYmyZUuzAQj8u/FrWqfZ67cQ/+9eW57P1IznnxgyeAq5nj7wau4F
9M5KFjwIIuGhFwey6uSPMVw9t8GHnW+yD87eToOGKHchdumYEO+AEtxA+00xPYYGU/cDaA3vckOy
Lh5+o5ve24CYK2S9kT6UmoSfKsQocM6k7hvC3QqJgfcYUdDgS9wlUdeD5wXJiUPz0SGEXODFb/Rt
qTPWoHPZ3sydU+W1v9hP2uhAg6q5/vSE3Oaab6AYEWMtMjJCT69uuwtXENT05Sdp8OxEcejH/Cvm
QSuB2bCT1UB5kTNlDU03dqusxAiipPgbkYnJvPEM681ihryP9CKYAhHsRf2ibKyfyFUwpHSfdI7y
gP684uTrQmv5Ul8arTU71GHNr5AqsdvdOEcjWuO018JvDTTQIWhbzL/oeuN176rLoDIabB/5aPOr
7s9vfENwuXKEhArndUpsmtaLXce+POlDypAgnoMcfjyxpnla8o6RDdJ0xFEK7DKXDaXg7d95aQUj
Vu25pDfiytD1+jqUtutxFVUlz04cwna6KitpO44CbO0W2F/Fz4mkNYHsMVc5PLHsfWSuT0Uy4ysr
OtKQDplBZ72uWbTU7rKwvMug11Cq0AWvHvJtB6nNWqmdBb+PRE4ORgKdhvauIw0qwdnLe3jVktND
B5zExFbhAKK5AScglc7ie5j0W5mpcpcfRrI/OHfff3EoYAUijjfxwxWNa7eIJyN4lozgw30yLjSn
Aj2WI4IG45kUOcD6FkO/EmILtFQu+/LGDMFhvZYu2Nm+wdJUTYv6dDwPy8TuX3X1/nn9+LYOLCgm
d30hQC1bMFR7dvdqsYnCEXFLc0utme421tGjGZet9sKY6UwiTUI32SaA0PGXmZahEcWDvSj/88ST
EBKa9AolBgboRG+YEGi18M7HYg5zwoDQvBhKt8pZ3wgTqYFwnSh6Rf2alLdNN/BdSTx5pEqLnshs
x66mN9ehOCaAyvSj0dLmPHa3dA649YtrVVCNXcFWqIbDY1BRqgBbrD3G3CwSPjtKyRD/IAPryK2V
djvH768t9kgD6yhNSwrB1elXyJ9NYIbUtHVo7CAQuNBfr3ByBqPpvmzusAAnnBZvcfqSq7zJFyCQ
Xto2SUjXZjheCaW4FWwiFIWrCMgpVv4fLpibnFbiqQHt5U3wvEPJGqFmxCJQI+EtG9rwm3ZqfDP9
Jh2/O0rlAOEA5t6nyGg1aoUH0SuMQBf2kahAwvynevXUMZEGspAnoadV0MdENU1diotJUp6Xjzic
7KMAJotzrSSy2Mc0sSHro3mQdxXq7LRrg5wgH9K51yF3N+ufd2dH0pHL5l/nJGcn6p38/JfodVjC
8eXnhpqvRqCzZmToFugGmxW6STM3w5HD5f5R8non5ox0opobpRuCy8A4f4DN0Ebav4gjJ1bAwar9
c9xAeHx97lkzURUR/UkOZcRp7yN6KEo9MtFncMZ4LX60kgIqOf6csfDApWp9ugNM+rn/6xIoUj8f
O/Sh1sRsa2hgTBW9wPpN9sp1fJM8+EhUX2sv47qNUsgcKNtMZYDLuRr/l72YgEffhspvUG9wNqlk
KHTMt0i6u1I2S12d4rr3h9Txalj+f6nqjdvHOV4VX+lfPw+onx5e1eLq0u2wRtCk0PfRP5265eZx
AW2MIPscmCyZmkEdqknGtDf9Yw40b4zVGzMYZdlcUyqiEVnRvRVudKoCzavciJ8+5taxpRnw6L5C
78GBZznK3pouzOi8HKq4afYiQB4iB3VDIbLODN8tlmyE1ELSo/0ouKB3v2rH2jVnx/ervmNq+zEa
iwZY3NhtykveThkALeJZ8jJETALX9grUhkuwGdbeLYKscuoaDuO21DlbGWdYSELkO/EWYTrIjEoT
sNJhXtUBrLQzKm1/H2ujMZtHj+dGN+m8lEuxwcyfzfbwwI/ApxYzoAvsQuD6C8CzVNdPL1UMs8/7
fPPfWcF17P3nd0l0w6URhIBRJuKou3b9ydaNFCj+3q3WT/sCoYp7tQAbfQsOCOkCTaVEhveSJGLC
FBgepkqi8WNzkE6cIl8dVdrbhrjStQnUIX2l8v9wnHXxoq88XODHnwmNdiropSfnzeGKCmwttgge
J5sHhdU9ccFRSK9ARVYfbXgR+V2gmMP7vVg3HYhXSzxidpIqU+nPiQYdUfi1FuL1/hqz7hpKJ90Y
LogDxr16PfOqKPf/2q3z0xKl2+up63siAqb0fZVZl9YdIdlUk4++NbB2s8fINS4DqqT++SMMJG7q
jknH1V57ISnfVW2qYj0RTiA+Si3fpGulGVKT/LLQ8PnUbqBlSgltQi//GyUqb7CBMbl+9lyFxRKS
NlTbtDFeOVI4RObqf27jC8yXwkjzx2+ggt25Vny1gTBFc26odXNkb+qNbw1Q9HY6bI0qZMkBdy4v
n05nagGpD1ZFxJU7TIna/29tbyu/siT8ZrbMAW+B2z3qE31KlbOxaP8VAMAjonsEj7XbXc/DA4D1
hKRkwo6YjCWEwwn1Ot8DTD8H2WuV9OHc+ZM5pzgBPJ2x7H+pVJ/D0SYCHnI2hKemGRicaUmsS0d/
bxRDErq3Uoa+4JuSBK7I8JmqvnjpAekgUuquKr66IPtA9UavdX3m4PitG7ZYJP7SY1HO2SCifzY4
7/6R0ceenpY28tSbTymXwAt9/s+OXX5LSUwIfQu5sxzThFWKD4b8/JsCrvRNneTwl4TFAql4YYUE
VIkx96xdD1Tqay0hw1NTsv4eV4ps2kzPR8o6yFxWkE415dqlXXYVKsve6+lMmsjjZvpcnUNw4a5T
tN6SX0osmC3MEwXYdpRpVuQaTA3eSPl00THLnotSNYrAFXOFCfCcSOi36dBtlgPC1xnv8+NqhwBW
z0h57gFZG7v+IB1uNuqWNrO9nUqi+qfnh/LN7IWEtrmwNytNUyEYi8p30DYL54xK9IR0i9nyt94o
JgWwAUKe05GBdCsvFwCOIafmK+OZHTWaCPzpcMPOAaIOUi4VXQTYiJIDOdmjaPBaAWFckRQQJ4WA
xYyhjz1rjq3r4xwu3LROGd5+NNcBjWeDj5UK896QuHidR7LiIUxZ/bj3f/IQUjroOMd52lgb5Eo3
bxoTk+L9r8d3gpQTU8Dci761/JB8lt/fsgG8rIwotjOJDAzaQQlXycre0BeoV7sw6NO3UjLPwhvY
hE/FsJsqnigtg8TkjlgHf0t3+5wbB6puwIuKvXlLQEvsyvCnYApXvEIghHrODDVNkZws6AS9BzhE
2y/AjnR/JPK9+fepibiX7No82AgwJenvHgzL6InaXBomaaPZwSstfXcJEFr3xfT/vWk2ZYHp0Mx4
QwBWUD7EGQRiKwOwfL9mokvbvVHuQLXneo3jlUEByNNmXOJNs6PKkR7n4ikIXIIQdivuScW/HM+1
ey3k3WqJBI6w72ZL8TapPyyaISxTY9Ys896x9PrsRLLDjO7DpIMPS3B5Ov63uAWEhYERnhCIBNRz
RCIKPiPaljtFA8+t1VLzezN1tvDxNf2h4eH+xD8MISDP/lUn6pGe3KS4T383oFfz4NJ05/EfSLou
Qi/BieGpixqDPwZ4Hq4WliHHGAz/s79g+x7ZXtzGN/LJfIwix0AF5wAmreqQ1/gRNknB66U8LiBc
Absg6eXweiEq95rRAKajokHK9GRQkOhsH3zWAqNrP1Do/R1PcrvR6nq4pF0noQ9LaplzrCYkDJv1
qovRzsIF0+1XtQBTfEoJXVqiCgCiZ0got4iycDhuOOvdDMBfiGFHzTGTuQsuZCXP94/LyrzjSdHg
NMigUpZQew5TxLO6VmfmxQRwNMlyYnPJ8unit8ErId6f4CUN1ozNkGLHucc2Fh65E17EQDueNji+
pMV2VJrQ/37tOGjePoHacYqWX3BJftYridpPyhhY2zAgBpw/ppgZ05t4CzkdmEwy1NpLPHOGh8GC
g3iIF46h7xl3oFc7pDG36l8ekIFaKueAuePYyu+AAgSJX6Ubb/EroTCTflGTaxMSYfd2AEohu9ds
DZcgrIMaoAhD5/nS6sg3Rcwqj7E3ojeZRQD46KpUuKNR6x2MTylpUTMJQOzBZRY3Wxq7c2+AR01f
WvUGC1PNbDJU4xqXBkklpjzpVG13zqAUxTU6vgmVoA6qg0qw+Nh37ysEPX6Naq8crDydX9bUUxNq
4zXvkayBlqH2MzNS+RHqEtwbVPRdet5Au4f8v3g57c50hqCn6j1K63kWErkJSqlVANjljGxD8Ghq
Y/P3zDU1tpu42CHEub54VIrjxd7lp+QsU32m/WTNQWWpXVybpE4Wt92KSzX+S1fp1S7NfGg/lR1S
AdlfAfmp6DqnOYhzFn159pi1OfgZjj8mTvlrgDVyrbETcodWOmxJOQX5c3kxk5VvKTF18iu6nFks
PccEJOU0CXUjg+YwV0W9y4/6J3/qFop9k4kg6xdJFJRF/An4Vf5pwyAc0J24o5uXFwu1jWrk01v+
s2m0LFNNtdIprXsy8zkjzBRVc+rm6YzIReY/lVgHJjR8YJ6ZBYfsWNvKnLzcHEViSQ7K/2Sfxu9T
hKhsR+VHfJtvNJSBu4TJifj6BYCkp1+xsnyGUz/VXuDVLPXHB/HXbfm6/ioKncCCOjwRsMtERSQm
8RL0p6IgeKHjWMF5H4IWbZMFsCmoN0OpJdXsfrhM4xx5v5435AEwMKz2GZux0ERurvTwEj2eixI5
Oemhf0cJ3LITYiGArL97W0WE8U26L0Whx8TGjdQcS9lB2vYqeqoXb4aJS33Mjhh26HKnAtPbpdAH
UwTFsjaDDr4qATkoxmjDEbbH4zFSsqkS7wQAYLAvKt0XZnn25OhsFyg3eAheO4iNyyKH30Mq5lM8
JotsvOritllGca+q6pKgGqmFUK4o6qpjvkG8w6OLW2o38ueoJyJgC86BxXWQxyhevwqcquTihYgH
7KGxhinZPO3CIYG410h7/0eNAvzMAb8xlcxfhBDyE5UvQfvd7QzZvY0ezRVDllmcvC7D25AvkxiZ
dFTHIY0/lKhDm73ObiuL3pYMKfmqusNzfwW4zlwugK6dOdjPQ99ZiXzLHHqtlWAYaB65rq7kVqhM
Ih0ll4bPpGY2anfB3TdtrEqQT3hXie78jDq/6JKx1DguqoAC9sHex9xhQbIvdlh/jnEHTY5nXA2v
8rK+2Jnl++69yrIedP58E3RZZJPYxQ/K0W0MZnhjgwrQC+IkBouNL1JT9qSy2c5/oObAujTnm2eE
bx0AfEWtFc6yP7RMc0Aajkl4hQslSQcmyPll3BbYiRCNgqfMVMtDYFx/hodWFvWKAi+dgr/fLTxa
0b4ZMy36lKw3+AM9C2jIfOZ5/ilJeYQlyREf1SHsXqRJd8DBWmyCwJ0C1J+eeHhHCdCZ0q2/odAH
l+NgQF6IIk+Rs0TBWhwIvrqxdbx1c9H05+NnKN+FXYARadiKuDv8fTLff2JwrcMGjqPFp6q008v5
i2sYE0DmxfOI4mcJcZ2sAW+frO04B39pNfVIRsgltX2gZldnQn9EUMnDIfUtd0ejFz+AhW40ij9v
Zeyu9J6pW3/OkCQEmpxOR8IFithzwRNOGtoEELcS4iwQcsIt0sSqWxfDXXLBYIyY3MBLzz8hBN53
qSXubHQvUpFv3vPke6PqFd3CWAQ5IA3QxYExLYjQDvIMYPcGo7V2pkgeqUYL1wy8ahKQNy9jkcsF
Sfh61JiJO9Et/UmgbcKfykU9NlOuNLk/XXv2oGpuHrnSoICme+0zlViqrFjGvaxta4jo5A1JqlgA
zD2xRetN/Wjm1OrHY89mFKN5+8S8LWXAPSrdHY2odXOUXGaYEA4GSblMtOobaW4v0gY1F60rE5U9
Tz4miwHjvTeW45i34+qIfVE63hpHk8K+wOtb91kwbb6soBoZ89UYCH35BtXZ/HOrx31+7XDOgaNc
h30oG4cAq5k7bPud42mxrViH5ZGHAxGmbvTNc12lNP03MzZ0kdXoUCQFuS4vcP6Bg4n7ecrJjBoV
ZfT/vn77ZnXgXSql5G3PgDyiyNyAf2ageZ1PFRMv0q7CQvvRd3GSf6T5UlRuAQzatwhsa7Y8WfI/
m8HFCmpOUsARJxjoAbvkjTbA5DxMcrArDZIQRzh87qfs/fA2f4dzSIF+cW45FkGQ0hUBKfDIG8ou
9eN/u9qUBo0usQcGTpkunl3+k+8UVil4qDMfdb52FVuF8uAiBs/K8b0fSSYGsBoqUN7RPuDrIe54
z0fj35TwvTMy3N2YTbJFddNbh5hTDdi+ETjlgikrEzmF63re76q1uOuqWAEniViWRwBh0PemLM2m
LlII17842aXJZJ9f86ZXKCEewah9kVZhUPZQY+lpMMnXLvxe9pO5tbE36lUiMixSaYzD5vmDJ/0t
nO+MYSU6D8Xj68oRJlEsXl65TICYlwcqyl3koBRzZ9rZehbicWde3LmJqqrQhQ2KBm/YTnF1JydU
+RkB9Vcp13f1oDIFUCEFfHkT1jB7WpLqQV3x7oruOYeKYhrKOZeonA96iZZL5XUTuH11jdQnwW5M
lA2RdJ3szDn85P9azGR29ytuIrl37v0L4hhfcGsj/PW7YbCbnm2JG7uu8T6nPNnjXHnhzrDE+ZY7
SLlQSZcgVfiw+/oxOqom9UYsoApoffhpBYaCxrstU+rhg5H+IkjZyjPdKz5meE/RROcI3EVfH2dV
8GxayCyE6ObRFA8nL3g/ZpDJlYWmjW4VnkuZbGpYFKEi3Psg2gws8MhZM5vLOYxtDyY7DlqejVIp
qnOFCtc9VAtgZe6ZqzJck1qa+0iWIyGeVfwrHcHUVTZulSErylShYmD2fvrTkJFLTTj1ykcyE96O
rp96hOgPWC3tHm51pCc6VBXqi3kLmj6LymtFrKPeam8zEKD5EZDOHdOFkXVk1CgS6f3GZYUXQXBY
KsyhdILjDmPiGM0L9ib9dON5zHVcS6two2WKd1JD3yy3Hl5duxW62H986tvFuV8yYK/UPzsKstfw
hQsj8xlD2GUOyq1vqzr4VFDG3zpU8Km4WvQaDGNbsAOYHvtr93oCdJOz7xQvXgJydpCWzFZslq/f
1DJ+wwI9z2ZPHpG7o3phPpMC4mzz1VTV4K6cgokAQcV6jyTohKDnnnlFUD4xwjOXfH+lXmI4OLVN
ns8aChH0edPkcu/lX7KIHr/4oYQLKSCNAuN83xy5V68oJ3RxClAG8SSK4BNmY7PKUSIC150d6dpv
0kR2zrFeRVXE+r3Xgi6W3xBK7DcjYB5j5hEF6qz984tM3nx9lnqSv8+2R/7oPZBMjTGC5CMaENa2
yQ4US2zLhNpM98iAIpUZs05dFGyzflvBBIbZA0nWijeX7CCvhp6+1DEmw/qsJrnABVuhL9d/cGJL
aWVWQNIlJIp/52kBSuQjmYrz7vuN8SOMYH+fkQTjL0//jk2UrM4Cw6c75nNp58JDk1rxPdJu9LSW
Rg0MWsn96YFxg6YOr7d41Qm2X5XNm/KITTFCN0useGcOMtErT3BYVQB3e/y4SPGKOscTIfvX6z5M
HTOfD3HGwhYfYKx613m326OVBmrOdqE6g3F+B4R4oKt3vMuL3+u0RlMiZ/4piDGmE9k9XTZhhxEb
FNGw7tKyq7ifMDMVvU/DlYi2lLRxweBY/qw62yFxSfalMx5saOcp36VKWEUui88BMA4uDTHMuxF9
tbu4WRUuOqeeIbEUVEWQzNuoVJ+N9UchmFfZrKjI+h1olCYSqKZUgIiTnjXYizk/kIoyCNY5gqeG
9AKKSbNVBytvgFDyiSfYPDYInXXwkZzoQmBPkBxaBBQKgD3TbWZoeHiffZI2eimIx8fF8U+vrF6Q
092szkQJHvYdePOgMIhXDmPxRZD9OlvjFv0xrZ+VInH8pjzLBJsif+GHhkozDhxjUm4LdpTPbyx4
HcOrtyVo0wpSqw8jLTVo0cQldoZEZv/SbB+DtJPKp83AGbX0M1bbGIQ8T/rHn3azIz1le/rWGmwX
qNWgF+9ouGvHJ13UXpWHCs22A7ckIBFLgiUrCTVnT4FhJrqhQ+w1EQ5l7tP3PTL+G94PBLZOGrEe
pFrQJv7mf74hjDRSt6RJ/bkc/pbARqXpNibFTG0/HYoNxoJJTt3waNMUr+h3lCfqGuI8pvNUeHsD
a63unD7h4JKN8gIq56ucfVpFa3s8E5yh01Az//Cc63PLAtyd4eevmE9bcGccXDn0n5FIBmfE44s6
SukvokjvoGTxN4W98/QPJXQtjUoPn8gA5ovkGpmjKEtEtX/4ym7cUszY0jzBX9PmKjtOTiIBGrnz
sdQaMm1ip7XBqQLup0PZ2TojDy4WPzYghpcOuU6IR8pA9+AZ75Pqz6rM3jMjInaRyhZlPHpuDQ6r
7DNM0vBI40gPOgdVuNq2KCPbs3pJkjos24kpw7AZFGjqc9sWbMp1mSnaaDNS0LeWPfr2JXxn75yr
xLPBNu1RP8sFPsvvBdx9c9HItyXq0M3BiDQTB2e+71ZkQfEa+xxp0jEmEh+Oqu66hI/a66e46W6E
RsVt45sLsuZ2c4DNDQg9FkzLsuk9/fHUZ0u7xOFqrx1MuK1PJ0uodGI2eQA6rye8D0FxE581U7zi
pMeK92j5OVIXl3imVoeP8TylOIeohtNwmWaefr0WK5CAgHYGcRw/rpG/NOGD6xr9/mle1+Oe4r1R
JNQmCnnXgfyD9+Y1pQyKQU9S3PAuiapruoOp633QvKc1AS3opfZGrD5mB/A5gL9gjsF1ifc8pJmi
tgrobmrLhaFpDi3ZoQHRlT4zy4hlhbNE0EVgCc9JBmA4A9HS+EEdkAGJ9PI84fvd2eNt//JHQNsg
/7fVF8IQCMfwinaBPEc98FJ3+bEuyp1SO4XrelVcOpc/o8swJCTd3sBfY3XUDHRzsq48oYWlipcN
eRAdiokJQx+FQBUWa1/Wusav8XGY/u8qbBFmfz0cdHfP/dvZb909tqTUvisYSmCrOZyiLKngdrA1
aAeB+imvGmEO/jL5HiaD4BF+vaM25ydFDRsgPjAkkuB8tdNgilnVNOyqgRBJl/+B08P50dHwiQIc
SJwU+C0Z+NXxMNHXJ1/2Wv1H80sSk3miFHd+uYuYIuTnhMWgzbScYhB0MpxAyZ5SNjKU0rWYFBlQ
+c7W9L6CVZFIZz003++hTNR2IiwjPJflzQs122a4KbhclxUk4Wqnp/MGKJ4ACilPLKbTdsv30Ieq
yQPb4TOlagOA+71maM4rlrqhvtajhTROSWop1ogeS4gb59K4vRMmnvL9VufKrDGSnIurXmya/byG
ISO+R2sa6X72CcA5gKeF82v7HtSuP7aaOCbp43nQAN/dr66MEL3N9Xu7DXKhxZGTYnn7/J108tpj
M5Mi7fWAmCcb7PpstN5sjEtY2NZ+cVOnX4Wiuba/3gGw74I52YriInwzKl8YekZWCyrAAnJ93DCH
FWaM3pMg36lkhiG43mXW7Lo5FJHa8aBUay1r3edhj7ChFzilYJzY15muzoyB7uyVMIJvbUSY3hEC
iW7+gZJ8yDWAhMVpBo1i+vvr3Z0MXj/jRxJAt0lzPllgNymr8LtuP/A2ERwAcMtZvwE89AjUsrYh
45MN7nivhSw163/B3X1DUkXNvAS8EnTvbczZ2R8uHFEQ/k3gSPUVhCwTLtjJLzd1yGPRuz63iCl0
N8UQ/AX3DVIX1VYwRRkAEm0Hg9Em4bIAN7ox/+8AbJFIP+iWJoqHz4imuWeo361es+kn1n87YQ4t
PeJ5Tx/Jl1tSAz+aS1HTK/efOpE9WkuUvq/zwWYGI1DTVZfykHw6R2guVpmRv/ys++LOQKTwKz2a
c3R8vTovvCM3Y+bF3a7I0xT7NHptRpcWjX+HHQpKHE474H9RqonpLronC79vGiDeFnmA/Pjmbqrc
36ySspWEn5omr4n+uf3HHq0dt2XDimGftzNxEidvN3x6jmiH3BoTb5wApZpKG+hckmhABTsMhxOR
cCUsUkHjv8SsoApyRl12iOXfB0fnoaRuq3+crZsQ/aX3nYn++WScP0aHsGytJPzKoa8GuyzXwLkl
JSJ4pFSbrKzqmT+uZhOmgEvtLWG7qZay2FRJHMnmCrTHNzyHki7Zr4ZbLt0E9iCPpPwGjSkd/2vA
mTJBqCqQ699v+NdNYcMiGMIDwzkGaPYq+ksAHzFKWE1YhuYS5+qBGPw9wMd05bXGFUOHKprRkIf7
3JzQ2qb2he3mgNQWyYAQr0Bt9YsipuPXIgmdD8nj2dvVZX00u4/L78+9etoda1y0g8jmN0QTHBbc
m6zYa/fWmfk3beeXYPQEKTqW4gOTCjSuqiIuH59KpWLOeTyNjKH2YoXW0LD9Vczbt9xzZl365Ace
vgCfFWNAXv+jrIocfBB/7/L/Oz6MzYuEW3cl62z81TyWs8seueuCA9FtP3pFJV+f2HleVQKlp5LZ
jP5niKA4nV//FOVof3zP7aQusTiUaB+g/qMOXnztCjHh99BLgMgQPu+d1ctKXJwx4INBnqWPk9X7
BXmEJHUmrY4G46A8I2xJzzUbPj7Vr4XQazBZfMjvinS0grq+mhrwyfgyodRmakQ8V0sAp1brpU2x
m7gWq4MonJyrM2oEL5E27RtGT46OrJTrAlcqwXlM7J4bAPt+eMAzlBIuExgHVHe1A3uf4/m46Wvf
1qiGqrcbLaftJWovYTqK04E+ZceKRPbhPO5UFFFOThPvE4b3LTyK/cKxT8vQNHppnNEkrU8ywEWc
i3ZJ9z+sBcKA1QpsytjhuVmMKUqtSdNigfuedkS3Y0CmmhcEL1/OIKu8MCUeYxC8wTJx26WIT0Tz
TbI8rDVlQij7VFcHtyHV+C7Q3NdGckMHXS7D5rAIugD4wpn6iAmK9C8AuJP8lsTwroFrAJn0B2MA
jog3xWe4ty/Zsz3Pc2N3v7P3KiQaxcxouG9dDxBDQIOv+c6ZtHq18HXvFyAbZxQx6OF1XksWDj26
pXMsjjJLw6/hetEaNzj8ap8d2cWvgKmhsrr3QPrIMVJ6sQhc3nNmKhtdyq6oEOMKrqgbNbbiGfph
vgacX1HeeNhmGo1GSZCsR/uOSViP0WhLI0o0CoquXeDU9G6RP6OPXEFTyZSfU7H4qjU3PT9QfLXe
b1/4jryXUY6xlVPKnrJoFY2pWs+rSiCBkDV2AiukFXkTqnq9Pqb7TcK2GG7YB/Q4HQTYoMsPP5iw
x8LvEyshc9r7gEcO7ycsvXnkBQNvAZDKjtELZti4Ip0vPEFiszH98u86rMaMRfwhuivABo6FLm7P
lxXChYI8cf7AZNajt9DbQKIhX7Lu2+dbw0XS+xnZqT3mG/oA71Ukqh8jPUi0Fj2iBitUqhFvHlDI
wo3xyeKo/O6PyWjzAhfrTiHPOcr9nQYcyPfOqMWOnK/V5eeIRc3bvz87nJ6rhP4ers4rI7lRaEol
TQahdg7nefy4ruYRlsQ/VSZxlHqAWqZpnoXeFnDg2Q+7Dlm0S6zlULX9Fl9Zwrn6t5flt10j/Puf
KBHJAyc1kz7hlQAu43dY6FPGrqoJBn5JkJ/IoomFWRWTjE86NWn34RB7tJNrv+r/ztwoag/aUwrj
rtjUleNsh+NzWE9rg24rw4hTiM3szdVpl1HHC76XCp0vC3OdVz5wjZM8f037jL2IkLvqFCy1aGsq
6C59LarB/dpi3woT8ulTs1Kq4dDlbGiCTAl8XkVDkLfO/k611yKEBDn0dtAEnx6Yz833+yxNb5ub
Tmjn45oF3FyYTeoDVYx2lq+lINH/6uqOnqvVj2eflN7V0in2RhCPdZTvXOgwAp4ALccQoJcS/10w
KBvhUDrTGJ3Fl083M8LCAaf/Xcq0dVX6mK0J21Bh5Nmdr7VeCJohY0cz/erXKskHd609jOUKcX3P
DXLpXRxkKp+6VEOccoRSHbLIa92mwNI5n4oclDOh39Gs9Ll/yrTUca5Xpwww1Q5NOMIlq/FyanR/
3pdojja4IkJJVcNwPu4WF4DRbki2qDL+iN5/7p7rkta35NfiV7A5/o0IEN8q8cq3+S1PPDc0qiWf
4o31uX4StKB4sz5eN2eKH+fPxcA/j/o+FBsDcKioUz8A6UVipDoslfa6hOMSGjiL9sGoIlLZWh/I
Ov3bF8ZoYStsoebnDP5kttJCAO9B+ioJcf+I55RBkox/JctvZXUYejEdPZ6rkFXjVzuDtl0tPwfo
iqVr78tjyqFF5lTlkpk3+WG1GW2JuaaLWlT/MmA9Ci8nvIG7hhO8OSYwfe36hHlzqhp+MnwIZJAe
zv+B4wEtET8wFYV5ghuI+2QxY1PDROw/sPrxI9khmlVSCItPvoeJ8qzC2JTozWov1fYMoMOqk0Zd
KSIMBCkeK5Rt1mqT5MOHcdHDJNoyuC6cpo3QuvD5TfaxytxBKw7T9uO9QDzedX29Ds10a39jCgjl
jB/SwI8hpqFsFPlrJhTnGkeca24fJj+EZkQSMhlP0OrQCEX7AdwXp6AM+Z3Ci54irecrsAvcTR/J
RRJc2zXV8dgBxwx4HETfY8xN6a/xKhvHZ7/nasmVNgan4UUauRf/kfkObLLLoAoVIWFMEw6ejo5o
gXrPwmstkwnK9ZcppjH/Xemaear85C5TTRUlDcl96IPs4WvTlQNH4PB0sTdXXh/Z/lYHycedZkVD
HXuFvnlq3BCXbvQlYQ+rz5xaFL1fNnVnBuX1+UA6+uJSm033g+BpBJYTAi82vDh4ejj05uLbSmIT
NjUP3o/MfrF9whOvsq1qn5zJ8A/ddmihzoWnHwguMzWEHyiOoZBRfex4Z9CEQOAsrSWHjzavSys+
cNjhvXmfSmGvyi5X0S8esma/XTwQsAvrREEIJcKgyK0ZcvyyyaT9T72rXkmUSRGgYJ3vxkgLIncP
8dVsvGTWBM6UNN5fbE6wWuQw7gsusUvK9e1pXLAXVd53zgWVEY55pZXESlHB/lNVCpoSNQQItUg6
D5H1oNZPCdi15wA3MQMbOFKdU7SUsa4v/oJn0a96fQrABIh4ykrCD5mWWqar5WXg5W2d8hbmxaQS
fXf47tKKdOY4sfB41oju71/MJjBHjU/TbnFnsuI4mw6QzIu3yLEOHRhCS1emMVvxiOscEjxQ0lW0
npv9Aomleqm5loWwsCKK4H1O+F00VwUJ+okOijirJBXInPwUCySaZII9oc77JUk6aGG21t3kiVvY
s90MiDB3g842O/F7MYnk+cO7vrGDqmgMPrc3t874mtIg0kj5IJVpzDwpuLfHJGR51HWlGHPKB5hX
XG2kkp4plcZzVJ9j55TUesnZvB+UAAfnFi9vV4ou3vbKCvivEBh2yjZglbGLgJhwcIknb6MGYCWT
yPW+WgYh3BkWM2ExcCiYvXDhAPAxgdHYOaC3/KJvAO/G9ZeFYDUuaToXJK7IU6ipOewI+CKExLrc
tPzJa/ZwIpLWS3j9g/GSkZkxf7X9U2Dyz08O/VlZIBX8gVKAoizVIwZhdrD3ztSYXPjysTEdRDC8
gIxcMhIFvKoM3UJq0Sca9t8PKAnsP/VpTfsg+P2ebV9NCxHT65kBsOpkptFzvuGngARXsLpXzVZj
SzreZXSnBf6f86u9zzra+BoTqqoVLqqpHmWI+cCnHWbqiHSPXcdPJaaSbHDiT+cqq/uETc4YTOzZ
4Kg2nYFSOsfq1mFlJvol4Oa1ReIRbPfleUKcRVnX2Yfx656bZzgKPKMNipV808e5vyxLC91O/nfj
PoE+Z2m8alV9xZpJMMw3yc0dY1Q2RTx7bQr/s5tAfzXqm83JJr1ZEeP/AniAfsZqwBsQuPNJWQbR
0kO+fehUyKRSQncT22AtmjtHApwNVBfqStM/6r6qjg4jG2JhXY8Sd9BIZsJRU5ieE9pCKVjfnfEM
dtTuEtgVg8bKg22b5ApLod2KJC0EI4kQVmku+PzTZ3O3CJp8Ifpm1ro8m0Vn5sVBm4DQBUY8H3h2
clUa+a9AuuEdHXlFOIKJ2Tj9LJ1xfBY6/IhgqZ/tK480DCSM6dKA6+sprX7GXjuuL4YD7mioAihN
dbLSjNWALv8RT3im/PNIciR5eA/ZtsnWf840sc+mwbeRKqYnIWZRX16ysa+nfaNf+xqgyW2y4U31
GHA3tBFPO/FHpWMR5yMF0gSdqwGWVfrz6QVosTEgE0dsUnDafnPIOImdxEupZBVQWcRJszGfrbWH
ZYN1dODihOTrP/llBKvoIDwSM2C0/kkH+5YJrR9C7Uwzbh8mRhToE6e2xcuFOecAiljpn4zO5VMc
BAHYmG1e3alH5jYgMYoxmAMkhkpb8kMZ4MYAzOLUxfSXyvBZLVPdmyya1yqYgHL7Jc6DGVppX21k
WW8sOiGGrtfkljI7t7nDmXp0iLuegERnGG6UTVuqJKokxSPzyz4eLnrMYE/luqUYvvgrFTgJu5DS
Hh5nWCdMagJVOVyEvB9QK8edHaoo/j9DrHrIJKdnyY1YIqUMmopGzsbAH9NY1EpIZmdhhHX2H/s8
/tvaZ+f3+g/rqqGDMJcP53TFmi/k+7TzVF6yHm2mJqsaHcYkVjxqjRgR+qkjd5sEEIg65NZANAoq
1FMKAuMxiK6H5WdrlZhMpSzx8WWJPRJuxzB+WAABSdWo9He7+JYS2kSc8UKTuZ4Q8q+esElUqAWZ
WfwvQKZnS8CUY2ZKPRTi5bFjMPJ23Zf3Wb9uKtW6BrcBiJFcpmEYY6xsGs9EVl8v9SqP/7oHA5DK
hjLJM4ObEJdzq1D2gu7U6N1wvBtbJiMEH389IXN0SsxDyc5WZxa/1zTY3gyKRpQmx3PHvxCj7MwZ
6jQ49VrCdxofSBSf+L8M3ltEdtwJzNBtv9zubrVCalJekDyWfoVEgrV4Pc0HBy7Rncs/nJCB4AFZ
2LdIRgTgGgisO4k+SoNNBI9QiH8IEWNJ6MPemiR3wa3AzkNw0g/FHk1QdRsl9Svn+u9zTBEFPLsU
if3Y2m01Y+Hh0/ikkdmVTXGRhdnGbfCDKplDaH2rKMvIoi1J6Z1VmWI4D+k4+XFwQOGkAKZ8sPRi
I+TrQ3ZmEh+NYWgK49YHXdECZL3YnTDUA1ulzfwPyWdCQdzI7OVBYzYB3I7ZkbiOwQEwDOFobEm9
lsqixgj9atJTbS62m7PCEfCTvL3Ar3UgXc9SlZte/hSXfMQSnLw8VSJVij5GA1Wj7S5YBFojz/gP
g5awG3DCLyA0jvYfE4Yxeenr/NfKZyxPiks0ia538eOfjDWN3Ptwy2X09MbnmV8vABGGC5njx/Rd
yDbtUbHCchWoLmAR20ZeJIJNpBXMKwAaYgWP8TyXY24TWDPTGCMoc6yhecNyx2RwaHuWLo6356yi
NTSD5cTfa7TMlOpnSaUy6t3Pm2b7LokxT7aO+SS+Pd2tetAnI1fT0lKlq99KSVGz3gKxr6ra4pj3
eJiaD3DldBTyLH2uylsAFEywrkp62XFa6LZsfWCwFkV3Gb4JeaWuicJiPitXpN9j9sB2FN9GfAaf
I0Ye2khkFbtwevWnSOYilRh21UvO3Bi30pYvUbgxQwZt2cgdn4OysMOa780JxPcprLFmlNeha/Qd
AB0qStA2/xmF7n7pBDrIKVW5xRs9JMWb27LQ/JXcqNqO/TW6rsQfSQlr3hFFj0rLYUfisUh6yy3f
YD/ANJSkurrJBoTwzy3sD8xKkUlx/nf7+KKlCa3Bsx+ZkGkNu8ROH2f79VlGUnQ65oaPN4opbFCC
rw7IHJts4NK04Ffh/vYyxinozlIfYESZgjJahpbFU3g0Lw9a2YeztP3Ei9AB00vjaWQm77wMdbAn
2Qa0Ybtz3IfjdsBf4Pukt5nYH7cTv1V++VMYdJ/kz8MXcxOWUHjOF+TEH35R9/0GiLfFKkYzD0yo
wsdmzXgqX+7rHA905Q/BJ8M3MTl7YyZxysgIa9zbQ0b2pdevclCf2rERQjFIKpnm52oSmRvaygF1
VA9tQwmVv0+Jiw2CurqJ+Pat8k4fLNB9tamCyvkmAqeODgaG7VwXfy5h7f2O5Z9gL6JQ1ConsJqI
+nlMOfhcoQ6naGhphgKcBXL1+OMwlDpSQRQidmXXKGPKv5l/f4KSDTAz4C9X6ivc1MJmgM248xJf
UOLbKd4uKbKXfDzRqPiPtWe6spe5WljY7UZGLHOI2JKUY00ZtHJc4rLFRHJLpCdasEzl8Mmc3RjX
1N7kmxRppjEdPBnXR5M85gWyMk2o/adFxJ3lBftDttf54Es5hE2FLElFNe3qn6Sbadgegd4AUXIb
j5xpFJ/+eebyxONNNQ+xLHGNOSEKB18BWBeniOsZ4YXlzC/EMk2GbVdNItqEu+Cg0uaalV8nRnTa
xp55CsTYJXXE5xa1wScD6NxM3BHg+mLqXMBAmsj+d6drpsPzbExx2MR4Zu86GdGVEvkoQaCY5zx7
Kwm/uW0RtjEFkk1zN8OHBAfLHppZika/8R6Itr9UzV36HVG+BgS9qau6XUZvH50KszhyAnGcZIZp
iLYR+7quPsn6W1SpyhEZJmffBIzrFyfW/8xACXflxupUa8Xti1phxrGAhM2PRtNMY+IRKdgZioXs
f7sDvMVy7wi5kGIJ60rIAZCcS12C8LkaMYHxVWM/OjTSPKKgz/HolBZzt4SQ52re4nCpnypAIN9o
1Q5p01/JzcPXiFIStUtI+xuUai4vS+CpsTtbJind026cMb0s8oH8QsyUZUtuMw5B32OMPO+B14sv
yT69uzbCD6N4S42jiDrrSbl0KxpYHY9dfL30y4b9VImI6Bq8MdlIvBGwnlKKyRwB2T1kOEkH8/9k
5YHYSD9JI1tmJbeluGaHegnvXVNwKLel01voqZHcLB4hBKPEbLubbT99RXRGbinlWc/hHjD+4EuX
A2NnJu+5x1ZkcQJxSXTB28PIp4vqoQ8xyTM3oQqUUxOAmAZkYaLVDiTpjRJr4UD2MCBv7QmjCMHV
VLYXEvy2PL5I7hpRiFnjAv5nnuBYo4lNS+RMKb7oaiQcreqYejL/hVCunaIGDv9Xly2KryD7iwj7
03TecYfFFpmfrZ1n9zNMizxN5EnwsN/4XO7TRKhERYoyEjAY1DwnwZeSNN4Quw65PlNu6aR08fk/
6ompm07AUZdYgnaIiTsSqahjejyUgtQw18f78qdE/452YGCCiOOdVq7wnD/uyxW5AwH7xZ2TlDKX
frmD9LhtnTXJ6cx4GqAjhfOOuxkQ/vc4ErW/YGBm9Ne0utZh3AZL0ykVRCIJspijOoyRH2jG80Zs
6v4moXBg4S72fBh6KdVnNXMX0R//Ih6LHHus8FXAuMxDMRYm6ktithbMgGmOnE27m3C1l0QkK7Zj
IhzrpYpa25DN1UHNht/OAjxvhPROb+Dhd7QSVBXih75L8ROJNG1fZDKzY/NTU2JxT15P4BbV8iKj
2YDdHEsvTi8cHBGNGCAJOJqml1iGAcxlKJO+bXctAJhwf4SBVp5zNu3E/qEW8u1TgnCohCYTIQQi
JsfRkZAotehyC8gaPye0X991wEujtx8vVEZvJPIrLbjA3b47d0vjGc43qr3fWJz3CVjQiJFQZj5v
RoiX4x5sXaHjEA6/lsUnsTPe43GZbeaBflZpA18LaUDvBgSr5m1rYXXaIvEty0SA95zXt0HvCTLE
kBcxEJdI30Eic1YONVv7rOK5oKXR+0VaQubrHPMoflXP6+b05UfR1bPWQZ1lsYhAVy7c4Cy0R8qd
qA1F28XU822txf3CSyw3OsPy3Ozobqbs3Mc/GuCBnvmPGl9NmdOr+fHUUbvqKjRtQmfzK40TB/9C
bWVBWpQSt5wDGQlHcv1b1KEegzUHLmQSmED9LL5A0YzOdTzF/ALb4PVQZhLxPkDH3O5yjrNr1nyL
oGZ9N7dkwnb3DRzANimYWcIalBz5NvIt/46PcX+nAWzMv5PEQ+SsQprWiRHz022xB+iOJMbpnPlo
ImvW0/xLlXKqPm8TJRDOCfkR1ZYtQ+epyinAzZQbGKspZRTfh9az7tb8a5lBrBMZw5+7EFj9CJoM
TnnmDAkx35rLasDvQfl5EPIV+pMTNkYztuZANlJ6Ni065tGbgkctkcymPSl1XOdBKFqaUoqM5DSz
5jARMMr5fgjB9FHsaM74TReB0oMnMG5BDh3WMx+IySjtTxI/jb1jxqi8JIH/QMq06Yt+6VntZnTB
i1qisEOeEYbZvmieaxnqwyweTf4WhlhUCbPcIKeqwkm6T9+MlBJoWXXqgUhu0dwHknLbpuQHM0ZQ
eqcKr8frgnkBrIIEUobeCsszMC6BsExWGbinbnicMo9GUbQFqeXzQtskaEzV7BvR2kutFR5w09oe
NxbZ6J1ZbkeNMtrfVt/SqkKHpGgq5WEQrsiE+PCV2gLn3m/vQoONzOxJ2st8DvECw+vLLqs/Ox2t
UfUiPM4gQ38DMUrvc8sJ/FoQPXSST/BY69kaHkw2N8TXSCGKdhIkgXO+MBqntzsVR0EwaVig9d/J
ivG4RzFsZV6RVFT+G84OX032EAJmhdnW7Uh3zYTvYGX6p9QCb8PpUmtnjACjEL0Sgphlmx9zOkUP
jXAVllKcwJZJSZnGWPcTR/zPmIkcHx1FvM+Zla/TjH1kKBfrKH6as1jNYA9BWLvphJ+1jnrtTz7m
hpRQLVTi+qkwLvh0Sxx+zuF9g7X/AbbJAoWDc5wZviV6GoSQXzPdBrFlBX2XaLeKMt0a5W1DLuKd
9JhbD1TuWEfLz41T+fImwOtjzGfeSY7ctlkO3E6APvND5Z9Nv58YsMD5ebzs9ofhYfwfag3dlnNa
a67tjF1b/V+IuqioILhmiT2YIFsGRV0u3iu9P1lFhQkV2B6pVZ1ZsxXE3PyUghClE9i4SzVpn19y
1UcQyVNlSO7qsKrzrrCf/txyvgzMl6fo3azHWEnVSGXCq6A05WtSDXxGwVlTuoxF+m7uGWjNI5eR
lZGoiumZ3XL8Iyd/t1q8ELWVz0cG5XrQFD1gDJTPOCvJDIBme2Op63INgbW06meWsYj20R8uYs0z
z3YTNRR23hiMlZY8/ZH1A1ZMgFESOW62YZ8zmGR5uJT2bkHEvsLWXTnCCR1H7AKDybf8a+biP8Id
FUIsABXD7VXqzVdDUxHya2S4K0PUHC4ICPg3rWDj8bPKTXeCgzHNLtvJv0IKGYG/W1ySvHTEyb7k
H25ng4XE1WLrIfalQOcEwyTeC5qmQ50wEDuSVeXeOw2mqpUEFZMqLl7KjMFZ4cVeewxbtJjc+SF1
VDqNvq+EcdwNRGs5VpGykTEVdslLK5x6ZrG2TDrXYCmFNEnKAbtC7tjdl6gTbio8YllrmMU/eQjT
poMbD+SySaYeydQp9b646Rxf+gcapOZtnoX2VOgb6npW7cMwFZVm6xhUCpYXaCuj4VKXX490YLex
AucIzL0qoVTkQplzItkr9sj/tDbxpna/zVALQmO2T/S7tr60oXfqKBCOdQLuedgu5mk7px18rb6i
FjldXxHlPjSYObmWBzvVc6aByMNAnwy8u6n3ybr8IEd+FlCGL8OcdQ+jbR7557TRElaF5DvvoLVU
Mm6WXM1Fi9mVvZ9KXhZKB/lsvTh5ST0CqZRueo3O98tcM74vsLsKss0S03bFZD7j/MErTWh0WJ6Z
n+6dW+T4da4lg+6/H48pGd/sLBTWcIlwU7bY9erq2ySJSa4H7a/0cMWZ2d+ufGk5yeXxZmJYeWcB
qggdnsX74vBVmEbg9xrfZ43EWb8/ndCijtCoQBjVJCMF8TCutkQJgeUw1SPPwz98sZurwLY0iJgS
IvGXE/zaICYHaUtHim7oWoT3nsC6Q+n9hVtqK2XOvxCbuiAbKqRW5IlqfFjqWhkD8o3GVRYM/RDC
xD0VziMg81rHdyJDjmFDrMilqw78hvXtgG1hVf82pROUYleVhTvXT5hy/lBRpGHXS9FlMc1zyrek
bnvhXgMQSwbJ2jB24XPqoHjuln74tqcjnnsVlrVwwUUJxL3KFyz4uqG7uu3oWyd6QOP6mhAxxsaR
f7uQm0rtaWwuHxgXxMK/r8s9HdQMqPOXc0zOSWVOhx1duhSporvZNAMlreA8nwa7B0a4QUHwQTY4
6OHHfTLvTthAIqoBFTsKRnztNuOun7C7tXJFxgYVZ0iD5oZtANXGJ+wutcPjvxEhXNBogeG2y+/w
/V4W0zIOsbDgBFeqEXXGs1zaPibWSbaXZ+djTTEQF4KyAThVm6pHqk3kfqmL8T1Cj8lLAWWikcCW
tjow1ZuJOVeGnvThorl33It2UQ3e374ZyJSgL55kBfvl1jrQI/CW6cnr0GMHde1S0fEkmuR5u5dX
xAgWut/lEiq4un0m5csESQhB27MOl8NBIviyt/Rq2ngEcVoHYHmyWdNQb115j45s5W60umGS1r25
1RsMX+N06Py0W1UHOZv3B3RvMnXaZJJyvyrRIuKsPA2Y2HObiGYt+rLTtw1X5nvkpQyIHviNdcE2
9c33EvOxVhxTyEqyB9rSuVpdU7LpJ0Ulg1dBNGRdxNUDterLwSiCndsamAXScf9R/QZc2L1Y7bQu
oEG5RHQTlYLiz4wUH6lPx7SWmbbtFvtYKOBCXc4uX3WfIBKIl78rKjWGS4TvlhEAwSjiU4kjJkfs
gyM0O5apQEljjaUKOVsV//RSAiBUtYNr7heoUIw+lovrzahoyEmSaQKI3+L5L+f+6MkenSH/Utny
ecaI1kqJzuWGG+bR6Iebj/zf8Bfg9a2dIks+DuAMkcvqRoRS1n+hsQJliUKVPhR6czauop+Pijn2
XqBdhNMKGTBDMDfdJHByGJEcchw8Jzig8i8ThPBqyFfG0ymiq22ny5CawnstJc5ehLC4s5Pp3jkK
0GgMja8XaHaTDrhEcjfQmXglFJajVWQsKpPQef0yyCQZ5Ww+wZ/uQGxbxSzD+XGCVXtiLoxsFe0H
ngpPf4rhSaOI7dLQAJ6ClYh8AoJENaqzjiSL76JviDLZgKKzTca1M1T6BmmrflCHYY29vHNsKZDE
sRZecPW7S+pvyNwF0UzuBDgxIUT02mInZKHztsE1ERGFijeGajiyKce/mIeYC4wvskY1J3g988c4
PK5/fYb6PdfrK4kunfHnBbqu8ak011g7pc5ue1z+TzXAwRTHGlbBZ5MYrSmLMD2xNYAzN7yDhhVd
75YcmBC7/tNvQs1aR+HrszBJbtXK3PCp1K10DwfF2fFoueYwxyJ5BCKDfWHA7D14JhS5JymG1IOE
qeRAObt4K1fxub0w6XftvFJmGoBW/qg32rOTlp83qnswG0cmYDkCE1OYo8tGAM5SwU4G+hPhcz1L
U1CHGNgqfARvH/W1bqFMbkd1v+R5VCN4ZfGlK7P6sHNw62zcNNLESh1E96iV/HaHaf37SeJLEl2D
ssigzEen/TwEq8ZJ0Vz1Xvg5ij4u2b7ssRhNHWXtWgmKvJnqRBXS26uNAeYuk/UbTlkIm9TBT5es
IEBodzqbhgxhVo/xE4B8dKjmxX1Drr4hHMjYx+faXaw+YqdRWTaEiL9wuqV58wwhxrqX0ws93iWB
d/zqbmUHKrjwIuPGI7Sv0r5oXndLN2qZ8ryspv1/Yeolg14N7dIuI+aiK/D4YG0phTbA5iAnAdt3
4bnMdyDH+Gag2JXyZbqLVk3/QQJWSkPsRJp8By80q+Cqk3OQT8TF8B8+gKkmKUilI88/fMlgeuK3
no8J0IOaBG6q+JMhtjz7AX5FdLygcxX0lnaQv+3VOGK0P0XfTv6lbng3e7rCI1TXeWA11hMz09O/
ioagul6cla0eMCTtvzotwgbo58iWxZaaVamCbyxzZWZicA3/zTforZ4kJkgDBY/bX5KBekB7rqDL
KTPD9B8VwPiI+N1rkQA1c82frU3HM9G1W1GP96s5x/j/PTwBw6a5yCJg+z7P4fANXMVBU3LE3d7c
oXlqQ7HlHMK+MIgJdaU8tkq3np+p531dDKGe9TREmJNLOS8WrB/UH4gAQrcOtbBR48aoc6/aJr0Q
gkczmQGgAq79Ia8gjOTV2hxLMIpiiGLXYFQgysvd1vFFE6BEQEdo8lYp69r0ttTxFrnWQbyytMbP
VrINgpM7KRHXJnsdzmMNK02LVjRH/5CVE6PXLYWXKa0qGtXeRUpOYo8fDWXHOHjThZktK+vdDIkf
MU8PuHToZdsUpTyK25LAyOx3Ixp7OSdeqZsELfaI1GjdTcrSRFJVv9nHeJW+yox9aJeWvKXBwO0a
9rw1fnAQLCm+H85+BbEVjQbgXsVqMvtfG5rVJjlGPDOQqEj3Nwt6tdEzjFenE4PIxSiB+RrPqtga
PgHkdoy99TbhJI8Jpl6iaZtKe0QHy2OEOyRa4pij8Q3ZC8Ktmf4ywnPimvZwKxz5wByUJSi6/3A0
FZHlzGGsmJ85fcJcgrPOJz4c/0a5bAH81txGoveklaLqua8OIDHyNOKAolHt7IfoVK0e6n+qoJF7
0NqxlS3AaZEClNu2pm9U39bQOmvB/poAdkP1GBp3UZfI+DD0ZbK6hCCWPHePEdzEYTHi2TogaLB/
vkPE/QeXStsQ5YVKcz4KMf2nwdn5NiBrOWL6uIDSxSKO8G076nqiU5LnrsgVC3Ytt+r5P+ztwiuC
0yTJsj7ncvrwvGNZroQgYgQW9AT4Ar08jZKUa6b8Fwn/C7dfC9seq+Ldt3sMOLIevxpKVrju+s9y
iAL6l7PrxQO8rP6aSfwuuVvUmCx5aIhUeNV+I3LfBdfBCOXupbg7PfWKs7yAV0AH5M2VVfxJvYAx
VfruXA3dIZDzzN8oYNZcjJk3isLHSvIZA9mzEGBW7h30MZyXyR3gPsm5rlaqyUypvXZESF9kCiVl
x51RkcCk42NlpyIWJ+iYt/wrfsFQvJzUZ/wGR9ag+MEt6P5x8EPfwp1blmyfogFSpI0R7PGtO7nG
s+gpY7U5jSA0hbsr9ED6/BTYRpFl8w58AnwNeog6aP37QxH1z+DGIvPiOAL6hKlqbxB0rXkizqGV
IcECw9smcHPLhNsddyOPf38dP1bdYu/TfNA2eHKdWw9CxO9V0r4Tc88o3AI6BeGTkS52G7CCmv91
85HLuhQAk/vrpEUw7UcZ12SLALfB6DeMNHeiKz6QQ0ZX9JV6l8z1HGtmO/s4uCpqs/36LEr4eINM
uBGlzCxmZ/zx9Q6S6rhwjJwenF0boSzOL7wtLB3uG5JtxSmaHp6m2ILDRoMPbMncUM+m4y7s/UOI
XARcPFb5lUgjRqOrHGNYGUSjr9/VEbDmsYxBqgCY7+mlpURJBDNZxR2exsQc7xlZGwNkf+3Af8nl
D+zLoI7YgvX1L5/iFZNX2sXMMTHgD6vPce8Uexi51sxU7fsl034dsnrlBouBc+fVP4ZnWGFNs6IP
xb+0NQvpD45THPSqn7gvMgG49Ha/1I8RceWBApNiIS8fsA4S5eARNNA94QVu0dB6Rmkdgpp6tKS1
fdYQaY95B7f9xcphe85CHxpaRgQ19UTUXkQVpE8GidIb+n7BU9lCar/PbstoLBQapmlqfMA9BaDq
bonRONf7BJ0RE7b0um290BtIPD81K9dhy+bFrL8TzAJ994J+OthhwyIzppnAIXlQa5jVr0oakpEr
+KIpiTj6mkg1YOM5r39inRz1R+JugpNFvIGqP9ASqIjZCaCr/VM3M35BFseuT2XZ8Zp7W8kXq63x
uAbUAS1XkLuzSYV0tf6kTF2RcMK7sRJzoa7+VKLLOktgv8rNg7Df9KxXDIEFQDshjKVyeNIsNASo
3aWF6+IOpyoCvPkS9idkfwMI7tok+o/jf7aFLDKG8ZNp2a54AL6DY3DMe1Ihfr6L5zKYQKbNhThD
+rozdtwgOpr13+lu+4mLrvipAjMF1gc9sS2Pm/OCLsZCgBpp/ZiBWY3kNBazfoBPScQ1+7gmaiNm
RxsRQa+CzrYuPmq0g5P+OpJQOyZoeqqMHUvMmCEBLD8lL27ZhAsEvkIn8NttyNgrP/D8UFKYmNOG
bz7yRDX4+JotTvR/pAPdv8lqXFBKIo6Ogyuvh0VKb5/xUi9NYPPeTHdFkuoAyr5kv1abbT7iCmXD
jMoX+h/gTf0V305cHvGUjud4E8TPKk+jDRAlmUG4MPQXIkKzMCriMF32P2qG3kRbl38Ga3SQYBoH
Mu5vxOyS3OZQo3tveLpgf22hSWM6aZHVubI8IVRUXFcvQwaxidUtKp9EUesLb01qDNvqaMESgg72
PX1hu3BRfdnfMzi0isnrkSxBS1W18CNV25nESAxOvtJrJj4nGkAggUfNZCRUijvazGO+l1b9iOT6
5Ybp/umpQMJ/FnA+4Tp9KzQNpDJ8WE531luf9hi0baKpurIyBMNqUoi8wp33d50RbtFWriYciYww
3VkAnfoIR3b1KULAqy3qlDQ0JVGlZOU2V9GHkI6zmmP5JLJuy0t/M4UK65a9szMVprAQ8wRhRwi8
bL7VvC192SEeFt/BZo/5otwznf1/Hstfi5/YflWDtNjk46fej15yfk5ZEs0ihZxv962xwnH5giQv
u2bPJQMZ8rc3+c+HP6HwY3KPvjFoVHUe5dWQ8Klh4YOVYXb0g/k2xdrNvSpt/7Jp11hP5uBRDQkv
qsbgUtV0w43VfiM+LDa9NcMlrZgcYxI6CzSTQI8MQJOoBDgqv4JKPagSTW94Q1L1yX6QCPAMPyBe
fVEB8cCWBh/jl6FCaiqPjNWz5PGmtXcAI33ueNC1/B2/eZygy+e8z66T+hcLWTFeBsBrwstIJFzi
IYsclO1jm6x3TCyNLUIX4ZkPL3vR69/afbHL91CXpQ5OqEx9SGo2nHZFC9JKLbk1shBCpR95FsFH
rrokqBUbFTWh5uxapzpheTCbzWXmRFERul9gc6WICJ8NF+x8w0QEELpBXtnSUdmgmoD0oHLEJwLF
s8ArpPqsjTutHGgNPPhlhswapnIALO0bj96Dzwbg48nBsrvPkoHGsyWjfG57L34Y77ooKG693QLD
8fFJUguBHpGWuJObjslKWhwxTVuWcvFJTViFcZVgk/6msoci0v5NwH0jHO6I0YsP97+0X9kDzzRh
TIAJO02hUXEC4Jn5+uAZc3GFgXXGExdoUjO8UXxMkZuKEix+VBsJDJuOxHSUuW07+3tQKluF/R2/
BY5+IxQMvHqHXZcVaKsEAq6xhAozpU1YMDJn+mgwtURq+avyRyAa+G6mZlAY3kpPzaXBJ86cXbdr
Ji2Zo+W1dPaJIZk+pBwW1ZRuOQeh2aQO8pqXQ5NU6aU0uRiKS5NWtyMvC2PW+OuLEHuFAsqfGW+w
kkHasZca4/KttDKdx3ONRocZn0r9jWljYj4kAq6rzf0NWkP1J/NnZXL9+SNY0vQsnsf2Zx9Z7ppj
nCDFFuMyqU27Zwvc0+u/yOisgggQ0ib1w9nGFq1rhZjZRyESe+EN2Q8XORTJ+OG0HjUgHG8NHrsX
jb0bfm203DNE2upvpqhsmXBOqIYljNW/OM04vxWD+w5bZXUM10u7gUul9Ulni+wddMNQY3/y+F5U
SKaioupzu1AWqosVcAFbVdgSEgX/ube6Ytg9Stw5KankEs22QkX+of3cQp+fMmx2ZG5p1SM2eCKF
0HYChESgx3OtoZz8n4k8PJEjPnZZAQlwCFgrrqVbcqVvHK2fA7NOBUoAjWVAsNByt4fOvu0Xeuki
cBCyo5f3MZ0EncSmold/N/YrmjUMsCu9TFU7v4a2T8nwC38IXhvdeQlj1Cm3jZlR1LLZxiRu4NGe
26kG97wQAyTNZNo1ezTzDYY+P/JmsS3DPryOVDhhyLu0yioVhyXP1r7xYHPK2nqTnsewrmmP7mDa
zumy+0qaSCCgIWQxruhswjMDK7DgK4Z5ycW2jSbdn/y5y7vAN4ybWdzVOKxGovmWbMvifZ4SUy2t
NSoIKJj4qhW+PGBzFJFc2f6p+3mnbu7gTHgH9MCCGYSQ+BYD+Lf/MJD224uyVjrPjCGp7mqJzeqx
KoZQ0nnHFXr74qEsYa2ifbaaCyJavH4wgBWQhn8eEoylEkYf0fJ5DVRuXVGdrB55dx3yk+pr6sxd
JU5ZObYGl2dPUwKjjfd7XFpX2gmcf6cl+zgOPDrRzGmQ9TN5V2bzXKAAH3onL5PyUfm+NKRr+hUA
AJTy5xx7RRD85d12hGz7zNki69ggFw9lRilRXpwa0kZQd1cSSqJhM6khPqnc16aytV8wx8ehtTaY
fKN0cIWv5rv/qXnpMaGQJWzI1gnmrKc5EdGFt5bQwWFJaN/AoZHv9+2z+0GQMTkWeaotFmjSBCFx
cx9xwBjqqHOvjmYrUvoZ6OBpep2OC9TZS32aC1nTP2R+EdIN2lSUJB8GW14xKS4zmFnOfTo9O2cw
9A39cFqRSiy1m+RNsTdPZpbNnbyPMxjS5umehsYz3t5/uxkELfmk67SAULi1C/5a+yUtKcC5wnCx
S8/unBmOFaMMasRV3rCjCJmFUCxW07c8GeL3WKM7usB5XG2g1jWLu99y4rid+S2iudi/zic3ASmx
bPK4lXppb/IS8venawlFvhhWEODRUtf+n8kw1XiL5UgI29xssmnahFasNgLdkt1T0+1nTgHQYqKr
PlFOZPmijEwFKdnP+EDjYPmxoTxyqURNWTbBeNOcaLufWhRtzrZoRbPFIdZi+F7Ysust8v++HZhP
ksb+k0PKXKYZgXCY8LgG64JgYZkRb4+rtvM++4NigQhUP9OEejf8Pm6adFHo4Zkd/MhZjo6aLuHK
QDRjvlpFidHlR9I8JyAX+DE9Eux++Z4y/+hM5nDwUZTpBMrs4dV1+gjPdQ6V+AATmAVz26nAdXV+
lQLaYuRocR1JTnEJppyPWZFzLs2RSHKdy9vg27rI0eXDgVE+NzKsr7CPNkguASoPpBIgLdSJeah2
1soNnafXmDG2/UJqyufaww1kHQt/0nrWFRKXYKWFh9IAmwFlkwubz38Kc73rzmpWkykhZUD9KbsC
42U9/UUdvOhGlWlRjPSArq+dlZPEkQfz3JaEoXzT2h4lpiqz57FjXAXz0rONUjbCI6s7GoDm5nq3
vFcxNx8aEH8UfHjxBT/XQMYQ6d3gT5yuFBkvy6qp8v46CHQxCrf6hySK7nf9WpW2VqYCmpyD7Fw6
ekVDhxH0nDBg3d13H+ktl+UQsYXckcGKIVNw8edoBzhjnjUBBLrDf2gwDetZkBC3hTxBar5bBjYt
3RtNNj01Kn3IxDmQoRZ1FXo8PXA7+nnmid9wmiQF63qMSdE8dvhLQPcE8/dGYNdrWrcE2mkqTUhQ
mANrT44Dx1vaNr7BunRdn4uei6lFlOQT1vzj76tGygn4nhcWN1Zbxj7Yuj5wJJtv/54ZimNSGsjm
JCKqnkSHvNeMnTdpK6gkgpjjxoK0AXNor1YBgmB610vp5SCCgrLwVYg6pnLDC8eNXS0tzNA/b+vM
Sxk+O7PHF58jKIVIlyFLcboERnIbx5VPWt4/gT78lQgic6ZhSzv9It2mvVh29CBLc8R29o9GwrWp
oBJDvg6HlDAR/1+YLnHODc32Ggoh5skwsvEruKLGRv/8TiNH2HycFu/pBgDBAod7PRezsybACDqH
fnqDThjuIlK+3d/pT1RP2xEvwt2dJZXhGhYkhamGoB25DShvM0BUq1id8jFhchEL8HIrf11VmHII
8Hk4eQeFX1lRoLDAqb7ifsq5tVDtbN0huycoWPhAqdAPjaAwAK4eyi/ivCLUh6oxeMhOsOxAx9qa
5Pec4nCUPpNRof0MsnVUyAwQtREa5F3+z076rQxhVwoceOdZjommiY0ahQksmIwA/A+EbVQqLuuI
grn2KX8eUG9xsoKIOm7kw4QUH0dJzIzbadvzUhqtcV9vN/UhVBXJf1UXVRSwZRB8X/J7yP92USwh
VoV9lNME3uh5d1i1cwad++C4tGkB0RfhyxHW/gURL1zrZekXxlhBHMdye+ciA6CuPWmoHumIw3TH
JIgJeHoHYuymde/dvg4zYc8kG0eqVRklbA/y9f4PLSGvHQGErthKyw9a44gYOGeu3UF6J19Vd19g
jd5Rg8b+cTdYLhkay2LNdXJ2m6QrSX+6HunZ05sKXU78XPjlFAg7j68zDhp+bHRKpPTH9na9qHdJ
H7yaJDQVO0JB4W1vxucNe8s5fS61lo8ppt8kh5fpTzYrEhQ6ydmhm7//wfsW16LDpiQhHPRhzsdc
CnF7Gx4arip7TfrEo7/arr1NoIrtAac406LvI2+fBHqnN9REPbug1PBdg1SJMFXd+Yt5cX64KaT7
HbiQGCP+Iwo5SQHrXK4ra8FCbVl78Rva/r+JBaWYYM2HvOWISa+oT2UHq+E/rqXMOGyvha485LZd
6aQHFJ6cfxVHcofLdKxHDN1wu8t03C/ryn/BYhWM7fMwcv4yHdJA/llVuzuF2WLWeget3JJnbTyn
vma8Puhh5noRY1UjrtQm438vZqqfhWFoMn17y1Lffxpad3h7otjPnHuXNWaUIlI7w55xqGvHLSm+
Ak2RKEf0wJFTv7I64B9t5R2HunM+rdqc5NuAYPHvMfQzl8oFCE3Fab5zfNHfeiid3pUeieVMYMLr
y/b/wf4iE2oMCPH/nZu08V1PQ3gkB5cItjr8MIbWCZUK5QC8wA19bZzElblgOMa1wZv8lIWX91Gk
mKYXYiuCpyPMSNdUU3qD0v8u3N6S/5aG+JWYPbZyVl7H3+tfHjFgAc7Jysq0b29JfZDxzs6Q8XM7
7tumeeq0zREggRoViaRKnDqWq5YjtbZEImVsAcq9EWYuO486JwtYm3pCSN13EFSzm/FP76BFGOR5
jKNECw7lVh3U7Nc5NmR2JmO3Wwlsf+qkj6Esh204UxGcC76zWXcn89Z0pcArYcWTETmziSVgef+8
UxEV8UK8WHzHKr1zZio5jdEwRjNzPLuX+yr8o7YiWj8JDPp4RxrGyniXx7pw9csZQOO23LlIXDZW
bomTwXu8zmz+/LvUuOhLgjp2+bLG/Z7YcfnGSEDKn3i0H7zbzrW1icY5GcR/bvyHsAKzyy8gWis8
51HIe8x48L6WYHX/oVZjs0m1EnQJLW4m2CbSfxSLq6N+8gzqCsIjkHC3BbGqS3DNMPO1T3JUpuPK
1dbhy7CUATz/Df2kq/sPHumn97XnGTZecmj/EbpsLFxns8/3c/NM2S+FoC5XHYNBoiPkPZksPkmx
5KJunuPXffNsNZ8g3TZN+3OLKTbZx+kfWqj0HK1jc0y8SMYcvO1V+JcNi9dSHNYhE157HDGcRrOj
JiVRPUl6b9CfcfsTmFrJa3z9pedgul6WejrkGZlavtse6vCN+ly3freLw13rFHiQNkm82pH+Efcf
Rd2QmxBR4vl++d0zGKXaU4naoyaZqhNO2iIdjYNKSCXb0/rIJ7jeZUvLhHNL2r3nNHOZnH9XgTep
1icNigXq9pO5bvmKb9JVmrmtgz/HSNe4VZ0NNX/rnNA9Cw1vBVx3CpAgclo17QEAL8xr3IHlR837
TWzaNL7xQMpB2RpS5hXd/zQCgM3vplHtX5YVD7ZkDRa5WGt8EMpQNhjVf/BuHJZgX0mAH79Tijf9
uH7o+BgDBBA7cz6KsvuOOos9ocWfsuI49sGNLKtLTeEfbBGAdnclNgKNiDlnQF5yT8Mwg1e0YX61
DY4Nh01RZ3m/aLdjVye+IGlr5yR/i+nq8StYBclRMhTzMF8MT5eQ88sWxSexg3UQwlGoN2/tnytH
Ys5WXxDGwCVBiE6EblE8oDRQTPtQIpDXDxzvM8bMWDyYPVs2+6cLRvTKOd3M8Hjq4Rul70101aOq
9tIbigBkXkESa1kf+vAPPc253XGwlWq8SnEV/6fKHRE9l1i50zbE/0qYfWKLRSgKYdBpZzhKS669
VTekxGuDBp9rqxyX3WaHt/KRaEv14QJdZQW4oBJiiqKz693+KI5rlcQEkWRtRTuNL3Ma1LRN/kP+
Outi3a4+/MhLqMosWzqbyXnAS0JbL3zusAcT2ARj2yI1mHn5p6+jNv0jm1CbwRK1dsEVPFJdBEfD
jvK0Vt7E5yfOy8fUAPM1ZbWTf4hr88vAu1UfA5wczy0GEXr4zeYcrfDfpOjMs7VZITP+ldXVw6xn
XMkvCncFwjXrsWzNOSqa6rPAc46YAEcFiBvzRzR9v2SKCsUq23Am02nR6crhubjvngDaDaW0lASb
gT48VxskPSTW4BOsjRCKW3uhrGEAHTs4BBLa+3XTKqtx4TYmExCDJFYN//0nBRruPlNwq77XlctI
xJttznOEbz6oMV6mlW0o2MbztD8M3Xrg5f9JqNo9TyQXmQ0yBbxlqPMqo8AtfbT5lmkGqJX5G14e
BxwScSQ+zsapUD+wwjl6yeRGWPSNqtd2hf9skhK/6qEFmRaiIMsp+pv18K7Ljh/vh9We1QGPiora
3RXiPmtxmnGs6huiXygEWGQKi4sV0Mglb4O7c7sxnt1rYAb6iCq4aAkzDKZ8WdO9JxC6CzLv+eDc
R5y0Bf97LBGIBhF/gtLXQWIg6KEppj16lvsfvOG5ZhooQCyk4OfM48kv2JNJXJksF5lultXe4F+t
R7PZxwd/RidQt4GLHJYXVOodk48TsQvVz15Eck8O9YihOSbb7vu7i+U2L8W1QVyr3Z6EOwKi8mqZ
Q05jW/aaKDgc1OUT1Tx9wzYduL1AAnIvGlj+uAovWmMG6OAAmxKuRGChQpgDqNI3xigyYpEaFpJ9
uW49uagER1u9QJ4KV4pnJd9oDdHicbsMBPfFkuOnzzi3PxohsBRCz0fiasNZxsaGLamYmYWMSVFq
420/C0A7+bbm0fTmVAumqpdgoTnO/gtnHbEIETVt3arHWBgnsihxUgtO03QBcA+l4kxhfU3ibqPx
jh5x809001qD2dotRY8dtbhDiLcrcjxuXS0QGotoNyudc7YZD5vYJQvBJDpnt4tUsuDBVbH3vzSG
DEvbJIMx/BTnMm4s8a2NTj0AXbxSTEXfbke2KhNFeXQkxLdewW0CyTdMZ2nzkA3mmIN74dNRRgU7
9SMBuIV2mJepqNGc81kOa65XYDLi5llqiXoibKHmcWoP9y5DeBxHQsXPHBezRUYBXHUhy1lrbh2W
jZWwHyDiycK0Nz4whwsRC+0VxotO06v05XIuu0+GnEwEHHSn+lyvfb3G7nY5Zxu5X4luaO5QZf4U
yIQGm0/LgpR+hAuLHqFIs3rB+PPKwE4YXf3WBX3mbgc1H/e7BZsrlpbeB5NpiTBfAAGUccKVySmK
fE0Im80ouLO9iYhIiafjRNn1unvKXbRNV8NgZDUalWqAb5mThvxwM6vugqjFkmL+TM60bl8DWT3L
FqQSURbD5pD51rhmk5hDJApmomu8Mehvfv1/IA2Iz1yxdseR6EWgY/zAa1N1Ftlx+7KQWMYuATLy
/V9Gdc/OibPRsAmPY3wr/zhsJmvb1m2GFngEOCw0n2hNjNMjdXazzyfCa5qkGBnpy4KfaK5jog5G
XGVtNojXS8M/02M79HHuEwDVv0u+o44bOzOtP4KHkje14S50wSv+/O+iqXwE+0/glf05YTFTec7d
3caf+BV5AMpm18JhHoMNeuWi9Ue+uYX5+5cPU5o15wdIDy/GxxWAqCw3YcQJ1qO4pZkHd9YAZvB0
B8M2FEfz6lcNSCNZwOc56wMoeSPmCvyTaCL2E/5Cmxn1r9IkA/aFIUuPXztmDlvs5HqtC+IN+182
RS5VliUlwJNNHKBDzTEzdWCx1tb9nHSAAd51W+Iu0ReRviRCLHlEzcx111MW1yxKGNQxHt97UVZZ
SsOFBdgFawf0iH1/YtIQC2xkZr2A+W0ukg+Vzsq8/VtyhdHM/TUXVkFzPdOjy5ROIzxg1s758i3R
MHMv+SwhsYYKKbsm/KVs5a7iyKqAEnXRbaIv5I7FccCyTvxCH2VJuApXoBqBGcG4lAhUeDSdOHUx
b4/ywzXCi/76fcNm05ogIwZI7AfnxOmp87MZgVGK7U/NipPoE5tM6P9IIv8kIL95ECjvh6DDvxWk
ArSCO9fE9/Z10q7BDs2YuZufbI2J+HHJ7yJY4/kKnBfb9InwSG+RjOkdqoEinqrvrq34dfv1gj3Y
jmkSpStLzPeB4pperWOkKDdEqpkXvv6MgwUL7u88EMZzR9fUE/uq0fozv3zMEHz0JVsBzVpi9lCG
FE96AJmUV32i3ppN4auW8mvBwb8Hl+xq3jP0EEJoDjwWwoeZxq6dj0b4zX/pgcAxwU/nrPWOjRO4
KttdWi1hxYT+jE7yp5rc4biDBxd6qW81QI7q12hTA+ObhKpH3nT4p37po08PstBLMumZBIaTIeQf
8r28ZHKjdfZ+yQwcR78kfl99ipEtGXMnOlwrlZSqeiMczgtJ4hYkYUCYg7gRub4O1odtfDVlxLwx
fm8B1y39KVi829bYSEfesfLViFIKM/9bXN3vL3Ol2YLflEZdOV4Np0+8xLn1YATJ1JD6gYx0M1PO
rdvFyl1eOsNR3nkMKQe6Z8BtQwnmRWuLHIDAYccZr9bEJoWgrR2YVDkeDz+rx7US0O/UgrsjWRdv
B4aHZeiPkbORrNmtGzwFTl6UB7NAns+7Kv30gP62Y5x5Fhx5UXqPAZlYm52nP7j9wuzpLwf0unCd
YAiV2JvrIP8UIWBaKkzLxZSdU7HeH11sdwHpefRnvfqJXC64EJSGxm7r+YIt8uaTkfq7LyI0Zk4y
ampDcEGq+U3VV3HFA+3CLN502jZXn/JITN+Q6Bs18yk6j0gpbJXfAgmnX9mNHvtOYK99gduVQ8P/
JrNoLMR0hWeyVxB5foDzT10rt3gpPdXdjgMqLONXm7qj6tr19CgxlhU5eFvnNqCAs8ezG2z/OWjz
+lUOM4RJKxrkvUiSBdQHiH/Np0/cH9mtzBsB1zH6BEfgN/jeIvh1j1jWsawFzjYY+4UvYpPoLfh0
theBAoGDne/qL93Y313rOX/atoEZFZ3WdMKkXWji9vLWNyt6hkvjV3rwVoeUI+q9fEs2mjqzC3Az
L6sPCWpWMIjLEK1UO134VRGP+vMkUeAaVbdUfu1QbdhoHlMaZ2WISS1C0j39XvuRNg/dA5PKItcQ
axMmOBqVIolYJokBizytXYQhLe/+gFi6MR1mUqB6OGiDnV1+wOPa+N7kHVpygsNmwBqCv/2nKlZA
d56+KMezAVY5XL/yA30eIp6TvC1BBPv04y1OUiyg9dtE/vNtFR97tLAPVYLsLEXqPYgrJYmEeYDW
uyvxY7GtmPUr3Ae+zP7LbE6ddZK1996JKSSrizx89mQfJW6gA4F2KBd4Ar0zIjo433QSBZO6q9DW
Sf34N03KLnTdG6tReZObdhzJNyfZL8ZB6FlQIhFgv1TQ0VzFDy93Cys1zHwn9S/490uHhaHJ32Mg
L0JtUS9cs6sfaOSoqsosZEaGUjYpHxM1JfVKEqwkPFIB40jB6HKUdGeZ4+Zu8ClEvzWDLv8MJATy
09vekKD+YXlBQCWBOI3b94D4mJdr7tjOpY0ytG/djni/jlsUl1dlge6hcnnmv/XWy9QdlyuPvZO3
6IJtb28s3EI8I77u48XUZHuhkUR/bNwoyaKb66PNoW6YuV9kTdcviBWHVRZW70KzeDardyW54Bc9
STvWgCA/qkZiKMeaTKci19Lwxe5EiF8qv6PlCDBj0AlPVryu+I68P6GOkyyMTJm9nYS+mkhGGGSh
ONIeMno33PcUSwcdnfGiAoN+nYkOcLOBcdouMOTOhLwa+uKA16ZbHjGZC/9wm3yHYHhBPaXjHoyG
IST31wcPbZzP0+e2kE0dG4FowRYNpEtVAyTRnQfwg11Ds6CwBy9kUGPrEhBhzVOWUHCpi54L9nLT
+tHCujIj1dCNI+lQrsNqCbftc/Es7F9GXsYd8hBmMQqC/NzEzpLO7ql6aEbyJtO+9iz6fRtl/2gc
vKEnI2EdubHP2b6gaK8DGkrj7qS9sxksiHvIPbHneUZaWCdVs4ngKKgLgnL0BayozRd5UuI6fozn
RXTwoJcWJmqMePNM5vp642mnMthN9l1p+/0QBpLEASaRfkvf2lwovAMH+gosJmhGygdkOnjGkR38
9gzuyZl2sCbLbQhQt5IAw6FK1FBLJP3N+kQud+UjHtf3qEf6ilDXjv7IdrA2LuPbQB9LcsKHbTwo
TYI120zi2mIylMIOw+Izaii6d5XdyW2F4AMu4JK3Y4Fm7yZWq9sKLMgMvdmop94JL0zNLk71IGEO
ZRJDZPGplsGbpQhj7IUJcsfDacZWUYomYNB+lVBO4XuXT1xYtPD9gC4S1PP+FKMHQHTyULFiGHrR
3cA7V8zlcdo1BQ3x3GJDN1nfEjtA5leuVpYingEi3sJCmAMT5kqeMb6ITimFkWKUztzDlUZnTj+O
Mtymy2wH0JEWl9PU4HXcMm9XHN/2WtL2Ib7zWG8MWTppj1MjUczGK2LzL3PbkLiyKwBWBB+qqfur
lRiQV9WkMKvMH8YECYkBWIMlTxRBO2RoF9un8+SMlFi+WOYWPGJdBtXxvNWOHpR4dLsgZMCbBQV7
rbptvdsvWbjvBAgXYVHYdyAvNMhh+ziNBi5zOVITfd1+uPpLrFjKw67igCQiKZmfSm6qmIBcupua
PR+iOR1+7OlsbAqNXSqQtbmgWfDJdcauaDpgeK4majo84aOwddzpD7c5Rt++I+eKrr13W7si81Nu
/7oxHEVNbqIEhbgBHYYadEamr9y/Tvf/8SvWmX1Ast/1EOdt5vyovvVEH06rJ77OS7OU4Nmiruny
gDA25UlnGJvzUoPsNCk41Kyz8NPYyQLTiYtHlV65Y4O/ejw8GNZrN6BFKMSeWMzGDfhfnh+r72uT
DZKXDwMh4eIaGIHkSFNCu0zewp7TnGcSOKSDcMzsy2CbjGxIQjWClj69TdLN/aI913iKIXR+ffPN
+cSROa8rdSExc7nImqiiV82BeUk9qnENeQHbSTZZg7u9auKdgzKqp/yvQ7h/fOeHAoDcWrPPQKho
741RtixuV9k/UbhgLDCnhWflTw/Lzg43044T4rK2Zf6x+4wqY+8j09boc2kTCKiF5lJdVOOjmpEJ
VNvdUXYsKPN3YeCqY8rB7oz+pj9qWuQRm7kKljq1YpMqm6Q8DbAnn2C/QiNycy2cVD6DeY0bqbVh
m6YqdMfBlE0Bvk17mhaOz29te2JDe82LS3MReqcCkiumkXMBcTHz4e+iULlSaF/1OUy353X7fTpC
ldze5UwLVLOo0KcMJScKGbYDB8wc3gaz6SD0aQxuzCkUS2zDstt4atjhj+lF1Pl3NjpKXMbqZKkq
FW0oO9HRmzgte1HRTGHVHJeQVxMwpb8TkQnOcgbOcRsHeoIXK7KlTe0t6CT5HDO46hdLB3EVuxjt
uCJMostyR+REvQbqoFnfqeEy54qIQRtS3G3sHkO1zNZMx9A44aRY6r91OrCS9f9LTZ+6G/vcJWxx
NHnOZ9OWe26UcpTQp+WzGGyHpAlCBFG0JSwcUYX8hCSNBgi3UjyMnvxoqsOEdMn3I61zpqK/BEfo
Sx1bnOa4QHNPMpZqS1spvVuCJfqsVGAUzdcLo6PlkyAtWx5AUmndplyu/OFgGaRq3OUETxAX6SPA
J15QZt+i3uTPqxX2QTgqAL2mVHIohsY0xsumTfZdfAmHAkDJ5JX3o+GgO7QiDct5HkYOGc99JrzJ
HYDh1O50yHKg5K0Lar0EJ+jLIbJEcz2uk0MWjoXMWs97lwOwx7WwaWaI2pyUHPbjcy3JroJtOp17
fNty8hmCVLN14iX+NeJpZeBhv34GORUunpinTzBSn7jSr2e2d8dQQoG6is/NiDsKvytxVVaUSEIt
sRyC18Vmj+zli+PVfof5YRJIhtO7t6znska3z235wanLHuuVajVxQzgGQ5PtPzh0syGA+NqaBQVo
eIBZzxHiTKJFw9t9Yk4CRHgmvA6CFKJdxXnGI8CSBhdQUUHgLrdTKw2zp5VNdHx1SU8AV7cAvDuX
0MjfWDFl+p0Z4IlV0pQ6I7M4uaEgMqYmWjI2rLROWMjTVu21VIRgS7UThU4eZ3BbANS1Y06SQRV6
Hwew/rko9SHVKLRKnKzbbtEmLCcapM7dc0DhfHx2DWWY0lPTugWl2sswoG/hHqXc5qQxnYGYHK79
DMXgbe0D2/SdNZoxZ8Fe2pPf89DsOuFgoh7IVpbW9vqHM/PbG2xL49xYRLjid2T+ZS4HJWjf9zlU
N1cfdIE0wVpnLlGl5pqTrYYVoXvsik/SpaCCbF2w+YLCVS9o5cjh4gGt9nbDhrJf9bC4gBc+R1TS
sw90PQOjiZ385blR3pX9kjlpBTt/ynvrhhF5Mr8OoVQpEiLzUkEDLtP3a7vBL8eGHMXFSbtXgBUo
h2PkbZUeOaC6ZNeJBtTUE3gDcRhLKoni0iOEXh5WmZP5d4l3raBVsBdg7KUbXGzVPiMxLJ1r0BVy
EKcs/E/SKqCowBdVKV0sJS16bQegCeBAoU9lhIElLFhrt/M8+X5FpHrSGtBqsybTx//o1bjSg/KL
pmZhzHJ2niMeOTzRVd68wLDmiih9clnmNO3UkVRP9G7KXh2MbrXRJeGZ4+M7atkI5RtHxn7jTl+L
jYD9BUbNibV/gQlZXQqkGB7lNMDzZBXjKm0hCw0DSLi8a5rRDwS9YjdR8WQVozsi3JvSchuzwkOp
Au3tBMpR6Z7lqzrQ9K/hb89N4Cvu8gI6ispCrdeyoT6Wpt8IOtM2cmVWmiVQRR4VyRVStwXl9sMY
gcPdTzU3c/wDDsoJQt/FoitLhXB1CnzONtBGkoQjvacWNlXUhEtfb1Moa6JtE2A9NU0YWBGXtikB
nwKbxfMWBOJzIyZS+odNiREQ1VS/O/uKtLq5Gwf9jx8FvdZ8sWGXRoMUFMiy+pm270Ye79WjT0sP
H2KoR2mqYY5gMe0ePwAsWa+xKSbEFOQDcu6+KOioMXrqg3B95T2KcKQXRYgqmpF1lgDtHwbzCP91
HtCrcUq14Of0WjnAWMH1HJZDy//pmXMDFWDQbcnzcuL5FEhMFNmCpjZpBOBu/6KgBOFrwshCof5N
jlcAwmIgxdx9uDcIZT8+zntVQrr+Piomsz08kf3ElAYq0D5n7I6TNdB4Ana1TOjlDB27dYkwaYGs
ji0dJkZfPixP06dBx1xjmEk9sbDExCdCKAYjVhizmfKFCTxjABvquqSvhW3vk8tn/srWV9mmG7Ht
KPSZRZ9rqMIWzrCwJJ85oqRD3ijFgDE9WCDrl77ghry1smmj5RkGqyBPYQ0rOLmjlV0PvlQOPxAe
iwKLM71SI6r/IZefDNeaHCFzoHuiYPKw6/15UxwbiHjZ5R3sfhkkYuNrw8oK9M2CrV85u5zbFljb
f7x7COLck9ppoOM4GS26ZQrUIafnhR5KQUF7J3Cd3c7qps/B09S5cQxW5eER6wVIpLrZGZ75E6kc
EmpPa9PKcBLQZRM+vlbA/mqqM8B+JG7PfDnqQ17wwaVG/VLmvNMoByZsDVdkh23hsi4q52QQuenb
eQjWUgbM+xeC1CuR3t80wepf7+X+Gxqnbcn1idAot/RsyMvurmiTO2D80FE6VwiFKN4l5AfL3AIb
UIsbqyqhQ6v8kK1nF7DH9yuq21n7fAwd14JzHysdsaXtsBDPb2/PfJCBcV3+wPZXmYayhGUOQJvi
PSl6IZipgsybcK/eFVcikS3fOlgndlr3nB0HytCG3aln/Cl0ZtaRaqi7tGUG9CjrJ0EH9cBuelf+
kHDDchXgBnIhMnRZX8VZnGNKyJUO+jwI3ZCdbzqSm5/qr9kgWWAx1IG6PH+hdFwlmqv/kPKfOCtb
M5RUc3roGq3TRt0FUH+71ISscTIP11bS8soJ6Ycp7ScQI2Nf1mTw9lncit8XYBDKW3rXnq+kPel5
13jbc/1znC0pep+Db9DfpRIhdc4/NY8AV8VrncpNZF72KPnu51VyaUAZSf0j/riMRcKcLAYPI7xz
0SxKxlEAIPFfzStFWireo1QzTVyJgEJfHLHytRq/jqdwJ7VP2uroueMZyCho89+mU0StxUUEiEgc
OGtbqLbwPfudPEA1rC9NdXUSsozgInqW2D6ySRZaaK4c9PsLBFNB+PDS12AeZRuGkaH2WiYjWIDz
U96Ti774lAMjgIWIOPaN0fNMggaFS5QMsN/jcmWYFhntSQndQfsJ2mY2asYMOoBzq764Y0hhItKf
Ud4ub10xSqPrxmOCKtxN7uOYmTiuQUHu3Br8b4C+vqeLKRH+Jk72RcLOuaxxuxNl1zvBTx23eNXS
RLNAVKs49njUQIFc+satN0UZY0Z2FOLXvtVv7URxuEZ6ZbjnDsLeauOweTntWVxWAPJGlBhQJ1vp
upoDi2Ct7tw0nygyU4XAYmNuQqNsQbSU+eb4EEEeM1QUx5iXRohodhVh67YYs+r0yAwGhnx4glPS
sAo1cjQvNIb3yMUkMa43rp5gqQw8RwWIplpxRuk1vwQyG7C/tBIe+mEereJN/ABOA+hSi2DMgXT0
bFII7BP9iHEplBF2Fpe7lXdNlL4Fx1fKaon+kiv4ZPK2fUujAbt5BA9AdFFk1HwV3pmnZMpvgyOu
8eeZbA2CcNiOJJvv3NCGyg9K7EKt2LQzULDrOlkBgAk+8PaLE+KAaww3/krNLGF+ikTsuh6pZt8w
qnw2kGpx4RQ4vSV34LVlviwmFzR1vMudqfxij1COI/rlOMcHegHSwRdKl8kMNYAcFI2HLNGRQcBV
Npk+OGUktuUBDMO8Jv9+XJdwtE+IEODPwti4cUrrWOeAFycmgMjicPET8l3TDa+hhZU4mNNEaGX6
e4748hAOayIaa0PjLj7ofMHP6muSzGebluNLSolT7dWoyFmrrX9pvjbtENyrD7ei+LojPuBP31dg
iyX+qP42hJHWpcisvPNvd3hpj4qEDNyGg2NbI08S0bdNsB+mxNf9WsiGtMT7ePzQaMWuZNwIr3xC
Jfky3g7xL2XRARP2C6cANhIHLdE460B4w2B+tb/Q8N8b/hf1y5a+EPrD6JnihseAbCT8VzXaZEyD
3AtCdh5Ys35K8Owb2vWQgWSt/CeGvtBFgv1CtG9OlkAz6PhOwKyG67HN5ufo32mFXYJGHQpagUVA
uO4kFwFrkGDaQXuZLQzYe5xbMgTNe6Z2j3vLcKyitK+IoTxMvIVVwwQxP86oZxnkIKKgDm02X/iw
pxtLNwX3D1JM3Kw61Yy8WlhTV/+ulEVGRGTwrP7cNAWXksBVU+UVAB/z5oT5tMPdztbZYT5qx7p3
RWujNSlPURDyG4EcU9o/cMAAfNwtp7yX0cyQrN58YBIDAJCq2rHjzMsDiSTaSVUHSvU00pNn2wlB
39wnwVJhUgGYrAUoO3l30EUUGCpDKl0/29J9X0uezokAWRW3BbFBIS9/TE1+PZIpiQrk/bmxrkMM
0WzDj0XD6lUBVpjyfHMNIgYn2ZyAtLzU1xyOEbKvTJz8aN91OERI7x201BofxDq/TcyIDXCZ6Ico
0bSS5wtBzJQ3gp+hCiGAyi/FWaO5W8UDCxLBrDLUfAObEs896nGhoCAqLXfDdIfLxisGUu7BmtFB
CZLKv5JdmLBNIuNqnJ/a1243ZXnWW21Z54EiW1AYNJlzNqEC9shLSDYNmLti7hoPshv3oZWo3v/V
o8MBX5e6RTcQwtpCHWuurBesHDQ0wCn4i8hVPJyQ/4wHfOHPz6zyOOQP1P2NqwOMSp4v0jd9MgFQ
km4W8YPIUaTmxQMsZhwtGtEbFhiub4KB5NpAe8MqO/YwAysyuewTA8XI9JCkIxCtVZNO+tYusYkc
VG+cMwa04QkPW+JqWnLJrTnrRVRcajp600/rNa9vuk5GTMpR/8E0H/5VtsF0fzdIDzqEYVyUR3Ub
vUu3/RJa1oEPa/pb5ENU9siZjmbNklyPuO7t0oLGJ34ZNaqvGpI/v8/7ALuWuPT1vm9Crli+1Wpv
oFWC2FIKBO7RUAax9G6QVVowsJq3EOiP+2n8CPVMyuUiaVTZ94qrw7vpWUorCCAa8AVUy6SI9+jH
6c2unyY91lWMM02he50MzOQjrsybWwT6iwUW8Zd+S5F6zD3uObCQIzYFip2hMNnoaKKjin0vagZN
E3N78gO/ckCAasVpeUqvE7sAcET26AFs1z7L8PXJ9a+7jl1RS41I8AfY3b2Jb/J89KcSooDCTOOy
x4R1Vks6oSNA0Zs/e9kc1lW5sTZyCcfIrP3LMU4ofcC8D8VIAiCQO9GSIUgaNV6aSXBJU75JWBdi
kfXh8py9H1Yb5YuUrNXSOzLjvOnpkrOqiUZwTkA5KzGv7Rux54qYICyFmFImatSHiDSM27m0/I41
sH2q/trHtmLLh8aBS99kJdt+1B+AZZ1s2zBhBMpO8uZlNnAZrW1uexTx8SBz/AnjHbKQEgiGlcWp
rk63JUvffTZUmgki3qz11yZ++pghA/s4TS9rrxWYPWn6gQGEUred7of8khrYSm/H5XTN5caG10vE
pkDGsZb9asAFegQZzP/9BAOqXKcWiYgqLIN7G3Qt2K+6E0gKsTKoM/XIdqc2ntt15oK//SA47oHU
tewBayVzG5JxYMsYSxCfqGVp/hOFAq4xhLH82y4WXe/YmLVze0fLjPOtViE8zVwJcTUwFIdIDkLe
QrxNJbP33u2Hb6P8/zWi1lRcapOAPAEi2kLXhrVVIgm1jtKkah/9vId0B9lISSkekw4zcCMRt82P
Xhpnh8VYg8wEqZsfkrcTqvMfhhMOy3FXFvcuugwubV0QBYpXcXL4tFfqvqeeznFQJgfN9iki3zjj
wNJzJSWUoA8beisFOdapZ2hOSp3ubReiRvTQNFQUyAQUlkRoViKeHAIFdiyqDkcK7OnE0RCH1Pu2
BVCMjV27/eGxXqLMH2ckTceBsrVDzwmcfCJaSnzeLDoqnHRt1khHWpqmUrm17BUe/fy9+xGJucat
3zY7FJUmmHoHOHrxW1FDI3DJEij9tUPwDgVTxhKU14iSruiEU9umi/w8fL+ExzOyJUSIuASt+Egv
o9ufmirWyc+U9L2cSZ8rMZwXBHyLfdAO8dD2Iti1HDpDvA+EvhDRnUg3MNvXeqCRfZ5LKoWhK5EU
wxvPtAmkszzddkgzFbARymQpjzvPPm0vqt7gqi5haGosEMrvBB01+Nh3QFsQKfOpFbVRpPEcvgOb
IBw69KxnKg9nKrfi+4jFQ6Mk45gRIPB+1isPenAa0HK1lawanqqcDGSFqulGJhvkHKOGTj01FYeB
TOErMhFiGGQoHjtkS4ikyDQjwxrwuZR/obNvYk0+8y/nlGP0TdwyXAaUqGFUMAYIw44de88WhcT3
ivJajwzb36l353a+WJdqV+G2DtCNfP8MZPeH+iLkOPgDcxIYAAuqJEzp4VUdIQYHrEh/gyRmXIhl
GnCtmWHP0qjqEwd8h3TwOQqrM8/j5FRSIQ225nqy+HwrRlrrgXPBn23KVQyeyIuUgEKvAZ1yWEkL
TaDhuQabMh61orEojmMjOCQPwSJrxVZSkbrLN27/fzCx76fsfdVMUBGSUIy/KBCOg6GHS9YNv1MX
jYW1HigmNYYgqQIVyiPEaaJJ3jRW4WrcIH2MXQ6vYrivp6uaaSeTsjyUgYVoMNql7ZFeq2+Hz1UT
ofcyPlk1fHXDxs/ij++jrJOeWyz9TydYAf2LpkSCD8fa0X6a4AC6yu537VHDLng5hzBwHH1uLQJm
k0P9ozj4VsX/fXXbFw5xZZfJbvGekH3YxMaBWveSOM622w/X9oICifH1bDBcd+RiI0BAQjjmmvg4
5Fv7EeO0rJaQdE104mXKYmyJPYlwBbJnuupldWbbrPVGNIB2KNDq1UvEa5IR3Q3S42Yl/STQONpW
sFzu58RXf/tC1UcFnzq3+xDra3SK+NORFgVhziJS1lnZjiFneu0brkQdfQFfpu5nL7WYbyqafbID
hiikqXgZcgQikSblo41yUgCBqtZvgj2Jh2uSWSqzFyssSCJA+l9NrvX+CHsJJgym3x2DXM+cWfZU
bz3b13HF2XFVA4tyeUNxDVAoppfdqK0bDzGl14QOT36fFIyLHosKyCYRi5qkRr6TG2mMS3U8dXQ6
/HJJ7tzrnfHyxTgX8boPOylyLzhtiCIcn65RTL+EH4BYH2b65tLzFoP/wqoNVbGIcryvQVzRKOhn
PluHWZzdhEzP+SCaXk1GoVWuR32Dk/6TM9zDqrsdQs0HxHqR2wQFQE7Swo/heW6RgReOKTVDYMkK
FJ9cZTptBTYS4A4Deg2F+/zhjkfKg/nxqh1PUvuRhMTc6FWS9Y2AvSigSDyPG1uMNBCtbZJHufVP
mLTPkIsp6P+rg2KApaAfrkRWb5Zv9MNr60UIWX1P34hyYrqqqDatuiXNoeNiBwbwRdVd5wDPYq3F
eN3Y8e2JQQY+cfn3ZZMipOlArexorK1AH5KcNqtoT76D3jYTZ+5XXE40L9Y4S1DX8xUEnesK+CZN
sxdI7YFe990gZFO96gYMUEJ/Eg7OKIgFvt99MjRHTzKPDZc1Q/KuPFOaVF5+luXslsaPeEQUO3jY
t5MgMskAFEfujhJ854mcLXbzHfbQl94XKDBdgw53VeKPCNWFF4KxshvV4rJbUPYGgC0kFLNtu7kW
loN1w6WGRFlKCR4JPdJ0WKBudJALoNbLYvNiUbXkLW+umVYyYQEDiAWc/+W3srjQyIiwDfvj3CMp
vufuGyS6+AYg+Ml5wmiTkNfwxb6mQ2MbHieOEo+sJyMUb2Ykyi+WAvxXo247p6mOEU4Msmvb50ir
M1pIUWHD60QkaivI+Lkl3ifHkOuc8WiyVL4t/D3YvykPWL+Eka1w4swOzmKH7Mg40q6Z1Rb2JWhw
RLW3nuHGsql2d7fWCNq6wvMU+XgS66jQM5dNfz7aA8qtBAmGQNOP1npY8EmJA/rW2DoX36nzENxQ
GeSGiIrjSo59hFeKaQcmi/7cbgwNmbDHwpZ8/rrExyZ8DhYDzS5Y7TG1iM73ocv8rUaUCxkjLyJr
/LcBOSWmWf6BHgHag9tZu32XeYlAVKVGJaa9GboHDLrdpjsbaQ2lwDvjGulQMzcXllv368SgESgD
Gm2cvwcgr+9eYl4D8PFe4p+stlk4Ub+Vmq/vVLoKiCwxjqzyD2Hxwdhky/Vjv/n2i0+rclE3xepi
h3vGko/+NdVe90Adozohn04CmYsoGbvFquDDDBL6X2IFlt/lXJTyd6/GH5zWLl3wHd8+A0LEM8bf
52Mla27eaZ4h7ZGfenKWvHBnLS892ejxdgpCefNFaHNkheDaLJSEDhuwHQb7lNfHIkhE23dudB16
7zKUmB4+pnAcGTVDath0CV7eO7NAHtEf2SJxHsGfWQlf10nlWqwKHWWLpBJaLa0IrYuABj9IUNCI
VLqpJ9p4nEMYpeXqr8TobelIxRKtLM6wDE5PjHz+zMxGSvIlmJ5QqwlZ7AZKdbKqw1W0q1fGtaIw
eIUsgCA9NdrB8kH+rlKgumOjPflNMFDTB67nym1JIYcydw29zNMt9fpmX5sFX0SDx3cpOFVSbWUm
8LZkDjdYSAs9mdgpTT+VuJo84TSNoUvNkFdlaljD1oUsetT/ZDTZ3K4mphqEJ5L6YGISHrPP7rm+
vfAEq/XtA+47Nhy3rA0CMJYP+GUkr7ulv2zmR4E+Y500cjQHYC//sT/X8XW/vmiWAiGLmtlUj76R
F4X7sy/Kl1cgHSvebs/kKGjea9ee4vtcpyEwR3G0RKFj1TAxrDMN6OOPqJ8jVAdi1cpWVvxo5Fqr
msiu5KWFbkrpzug8D6lKSDym/H2u5Si4maneqzqFpVE2v1Pda9Yr3vJBWboYeVcIoVSQkGM8m418
5onx7Z0TG7DuhSuMAcGykQsU6UDIORWtHe0mNMyXSors5Vmr3gPYgyaxMuVUwOAVkV6hXGdiK2a5
J5ET0sMXgXJ2ObQkNniFsQeZVE0bhhvDcnn/MLje0HVxGYJ9p/jUU/xFEauL0U8X5s3TBdxc+1M7
vnHTOGXQxbzu88IgQo45L45yECrDV7OtZpNGaBtGfJcD2Iu2K9FU0HFIdslYii0KtCwfc1xwwE+z
qg91ov7+GJG8dRnlBZjpaacR5XEI4BJXuJstGTw2peVJmqTfgA8g+f1XZRJwr2Pyy+lY48Rkwfrr
4YlW1vISvhVXWajy896M+QT9Po6T4tBhP1WoXOvchAthueIL453vg9gYbEGafQZH2p0CRMunIqua
QyXdVdVk7kRRdraAX/RY9S2tlBnBO6L5cw/FcDWDgJVo7Ytu0PAn+lp0OrL9tsmmiacw5uAougST
qamTq2TvP//bQZIpKcWSuPIQF/kvMTYIc5Kw3Ch/RemJA6MbmUIcx7GtZVBlpqTR9OkW9r1GPd6x
nDBsog38V0+qUFCOByQXDDnOclf47nQcKRvYBvb79fRftIfIKIZTqoLg9mseUCk/GwuCFQnSQBpU
QLnzHoA7/dOgRT+hI5gT+ieZ4g1+l+yQND0jSrmpNDFp4yeK8dtn1ac9GsrnCChplglqy00dkRQr
+U3drDJC2WEqFQkt0sR2DO4Xs1bmvb5xrH3tGbLQX1UUofvw2cMtzYyYMVUwV5ALCeSGd7e16xA5
1l5tHwqGygk1ggsoJsVkpETyP6vfmdYFn8R6YpFcCSQUJ/ZkgCbI9h+hMUjQU0jehFNF9CB79DCo
zZcRCsFdjWkg8fqalvVEM3/B3bKX/wb9ql+fnjM5FShgr2X9XKi1N0BBKmDJGbywCu4nuP/6mm/e
so7YZ9pKgHKbw1bGMJfYtdMOikBzCTeMcjY8AfJFtBN2rFwn0AQ1zM0pNtuNpLC4+MkYg1fMvxgp
yqNiDzPmGqvncXdwCC5hBsCjJfHD6+5NO86dlpFE311F52uT+qDE9z+0LMb3pPFALjKOP9Chr5ue
c2og0t9HvQoayUxPpSk78on3tokRPsQ48HA9Z7Kp8Zxtqegh/4RnhX5yGrO39OvoQr9e0OqfYdsW
M2w+pnJIcE7gS/Brd74H7xIExG6MZpeqCcYIwzL8AgEWMnabBLm9bl68I+zkLK1F+YuUWLTFUv4b
CJKPRShS9z5bn8M1beDr4d7Yt+bqCvV6l4do7BMoIg5osux4RVs/9Cq1mNKyGrUFTQbv+k9iimEg
IfFhg/b6yLQyrYDoMZ6OI6+PfczXY73NJ++loJ+KodhzmSf1QDXWRmipBAH3wrv9evtXClIK9dxS
qywrJaouGBKBYkEPUu9RI3dg0Fu+RwwvJ26PP9Az/2bfk6m/5VP2YJE+pCzqHoAYwty+JD0+UH0M
IYb0OhA013juutEehOgF92q9t/5b0i1DPY4QC2d+IXhbMKBP7D3AEzIzd7L5rv0IKZLFhtmL4RQk
arkcKPwG//e79frKjnwx2CAjUBLsABdCLMg21hojn6qwnVuoC1Q3jnu/l7nrcy3JMvTZbUuOu0Yg
WyL3Fa/7jM7MqayRoTn7m8aTjM0GVIPJn+LazHfJ4mvos+viVvQPY/YBJ0Dd27BtDqQ3flLcyML0
nYZCnF2Q2OUN4LXtTCVV5l7WmtlyKyFjMFzNwBIJHIV36mgL1ZOxIWbufUyb0XFuNIrgEjJAX+zO
zO9W4Mj3yG1HNZCr+Z21nQgc1dPaex2qLG1Nhu2qDsUWMvNLrVCuL9bcpigj4Vu++Hv2zEebGuxh
sHdTIgmnexLqHP63/SJiP8/UHF21dMZ2aF4oyFcHXcAmZP4Nnoj81tyfSx4V1tga+9Qd7uFEqw5+
tlLFU2kg1s1ihoXP1RtG66hF1fgL4EeToAHtRCnRyt1ukG81/U1rS4qkMW7lzvzQQUj6AKpRn4Gl
VjtVMtjvHOEAoblXsp4yqWHlTosX0hzcftZ3H2Il9PGa1CcevBUuEGclHVWhOw4NIM0Pl9Mf9BAo
UgYAkwreRJ6CKQwtRoXrcqe9IQ3fAaLn+x69mbXxS9gct3Q+7vRbksB5/rVhLb4OLb4CoqlcH3jf
EEogqyK2hnMkO2CUcZ3FnBjIzkJV5TFAQSmIZOhAgsbCWP8kDkM5AG13yL5J6Ms3Z/mEIWWVJNMS
t704SzZDy/3lX/cKzvueswpcX1TXrEBlyg89CFk81gQuxu86eI4EUIm9c8IeXdGWpthgKFfns5kZ
I1PvLXSkPaKSDuZ+OloI3UIyoeDuF4FgOs7NU8yykyyP2gN1ZlwqkXdfBgzB3e9cAajOpBB5kgFq
DiQp1KRoCX97rCVRG08veoIADOY33wDyYtFj1nNRKg5l1gPQg39PtuKqXoXpAb1xqjh7ITXwvB4V
fLXRbIKGfiVgRPe6UacLb+/6Xy8KmXnPtT1Td+9PkPMTLXIPhCHofqBfCqJlnPWBJKzt2ELZUCfK
Ao7+uxYfvANCJSaGnr6PWRkTt7/14ohPyCykqUdiDCYUSzWV0Jkwf8zG/hz1A4KAihemxmjDZWDQ
uvaVKvANhtf53Jn8OFGr3ZIYDb9LUeuUUHrfsSD14HOCXEkh9Z1ZtNtEzC8bsQiNUu13/j2hMKQ7
mzhyVch8COpwJA1nDM6uPm3k4WI4ntAJ7fNanLY3ZRa4PgN4gd7OaQ3M0ep9KeVkUN0quk918quC
sKcRjm7lHHCZFL+kxqSLi68/KFvGAe5pjcqMS5bQe6gMduV1Nlua3CWoDTM7uLRVmVFIolTb8QD0
Dhl7pDAWtYoHbtpLtOglY1qQW0SLoB3EBNzCHNB4KvttwrQv0x+wG9pY5pTARlo3lSJJTnP2m8zC
Ppfp3DANaqxM2lothA6wclR5plW2rJX1TcPGITMsP3qLev+CUk87QYuC/x/kbQ4vRk953sZpiBm8
hpMUukdUw2eiEEJvuM76MOT3wNDKug3/iHMlWZgF/1/iagXauAwvzk70xQ1nzJlusacaS/rwMTli
uxLfOkGDnJ1H22X0xuGb7xJApsAUOvl7X/mCEr7/nBuZYwD6JGfiuoS4oqBAQQP4xVRDzQMw9PX/
K2HxIMU1RB6mqzyZPEkA1hWUG1rV8Rb0uamBTFyIYm30hJEjxN0kfbWaeAojQeEcPhbJRIWKg00a
//VEbkmc+ywGSqPJzOj+sIheWTT209vUB0UeeBwfjY8QXaa7a/Mr8FQvb8BlWLPvJyBrUD/4GI32
1GHnRvMSk5XjiSlg/ZNvIiLSW3uREqI6Wz8ZC6Gw8gaQwjD9PLfZmTcP74t3ypxLv9gJFnCyxR//
ypz9QOYJ0BYAavMoN3h1Xf20zxaqhpEIPVg6R3JVoT7OsicjdpgchfMCQddLKE3FE+M/O3ZTGpPS
1VmZThkKAsoBrsAco7gzHTRpd7p+HPnSusC+lz6aWdE55Dd9ttUUzrWAMwVyTFwsQwqmHrHkV1ed
BXyj49PJoz38oPx3Bm3/hbxIzoaQAxmGbRQQeRhNWCKHfaekA2CKWkWRdMGrp33uMBPXRpzOsZTC
86VCCxBY6Ysvh9qGh7aZMhMrf3NVDEBmwJ9CsJVGSh9sZK19/UrXnjuHT5vdOie+CM4q+votQrUz
2TlJblWtvrgTRco1jTPM6M0t1WSA86UEBElBpg3IT1pt0PcNPxMKxniNIJJ9la0L9iDQi3sE/jGh
btBRjKgg6W2FJ6VhvNeEk/3/NgeTiXzATWe6Y068wbPnmjjYM5pdb89kaypRqvNAhgZ/DbFQQMlP
f4px6B9k8QK3t2YOP8IK6px9Gvc6nPJtNHAuir4oeTjbD9VDy98dPMBIcn/fRoxQjpb0cv574lrz
4TL5kzZWBzWqW1Z9R6vtU6VEOanwRScmoe/f3HVlW8cLkLH7R12FhVyimv+1HpTorRNpIbHa6s/W
NLDMFW6dySXbbOPL++7rz6gc+Ht0tmH0cuOII7qh0FLBRm2MTun+C88FRb34qwTa3DQ0qlV+/dVc
IvQduilALQNHgLLxRnND4JoV0uNMcsGPgh7uv+CTKZA23TKt4N78ScHNTOlXi/7Uuhi1wu2m8Ad2
t0LsiRrnDr290r39P/RWvFvBpFh9zApaN80ObbDynCd6Twgt8wx4lvq4B6JkSg9+db7NboVa5e1h
m8iZkqViRzJ8b4yU11xb4xs5Bqz2iPqORbv/c3ZKf2VXVMiQ/rqHsqzZsk2yliOp6xBefpWXggrZ
intpqNra70L5eUf+xeNyp9WK3MS7FomG1Aaa4x3tY//G7hqnBRNrdYv8ImAuVTdUrTfJ55+eybKB
7Jos2cZ0kfepwpjqo+pZMr/xJ6QHSnlZTI3b012Xthah1ACoDMxzsWTCaeMT0uMUieQlWmmadVCG
U4mJOftiar/axudWgUy4kwRUSlZkW6uRAN4OS0POAEV1vBSQe/SOv6VqfU6WtvnUYDZdOqQ1qlgG
yeSYQI/RacVUHA+hXbvlHLn131r0tmwnCkmMqIkc8iWxYTbxiGcZLKvkIonZjGSAFOYVZpsav3CS
3+n1pi8HrSVyiJybv914NwFslewyRX0Est5WCKiVWZCQnPS9KJ0Q67fwYw+EYoBtwDpcysv3MtPU
tbrp3hENRi26CiJ1VsPG4dUr+GMkv0j//Yj/jcag4JBbqFCBx4jqPXFJ/CPkJH+NVLzOPNVCxNca
QWFeEK+q2wwXxVTfJfP7O8vMlwaXQEx8Ollf1eESMOwFfFoEPIEq6CkkbdRlBnbxLhTxma3expVX
D1NjR2P9I2/R0tPcopxpz/bto/XJeZxDI9KYgJrT/cjmwn4uq8Z+TBDYlWNnjVQv8NxrPWqP0Gsd
iCQYJRjwHzJ3Wgda58Xip9Qwj2LK1l1KG7zNta7U3LWlcV1i32ASq7RIkIPK76wtd4QhUiZOIjR/
gNW1LJsFCJZsu2Ckkns4Gvp6jPpcrsJf4gsV5oUrh45rwil64UTHWJDxfsmZXW9YES6yXQce9oOe
vcN+GXMXQZMAhQzKM2m1yy8ubL1jcT0DMsVr4He3hVkAcczlkWRtkyogCsc79R6LdtGQOTVbic0D
8D2574yB3S/zD4F9FCpUa1yPw75vEERyA+ZvaOD25hUNm4LYstwWr/4Vy6PNiIS6tbvS7B2sF7zw
YuzMUpL1v1+wkRQ1YssSOgDr0dJoEbLXgKlz9rN6tC7w15Ry+jkiUbYESO7IDvVWOLx6bKAKYCVx
aCd8CZEspsVCQ1JI2+4ur8D1fDrj1cwY4iPb+fa6ybf+btc9xdWDi/pzs5Xl2NvgelgF8IZJiNf9
CJkkwPcj4e4ur0W7gUIqIZu5QWthT5po0r4pLnBpibJ7shWKKrYAdxhsR4VU1jKzJMEYzhcfcsnT
mWROHdfZlh5L+Z5P40S2+H0JVHhNdsZvrlnjHAjWS+OM35wRXPKmvaLAeN/DdbSevZIc4FBRVOfX
v6A/XJC6Vko1UvjHbR3WYKGtgJropJRlr6lp0bU0HzQ8Yp81uzoRballi4FSAvM6pPcN20ZoiisL
v59wIWiO8uua6dv8GELYYmpf/j70sKPvTO5E3BW36EuDnpbsgd90N3JPiRJ0nxHrKg/VRtNF6mYB
JwyC6h0xZEpwCK6hcTpiI4Wpr8t/kAZa4F0MTO/yeCgEFLfwID4ckc2V0lvfxssdI8zyuMU5YcPO
wuj/JhauERPvcuDhk+hW+OOaZM8bO6DrgHXbvz4Dn8+S2jg3qHSc21UIhArC3PW61J0TiDP59nX7
TWgKWcnfDiJqvCHT1Ns0fneTEQn4LBCzAc4pIFqrCrXOZYMgCmcjtQSfM0JCirCdCPtnjAR847F6
OENzLUMKVBc3DE9M1hrr9G0200XELNkran1kHJg9Ael/ra9hJQ2EPTBJixrtbHojY3cI9kxWKwAg
taQplfPPAOA0cMaZ9UwACU5fYS1gm7Qgny9DQ/zwKUG3Z5890koArqOI4H+eers38YJDwOr+gYi1
SuT7AUneiZRn8aHAPUdIE0539fzAsqmoN/wxBrpPEJyrbDVlsM4vMBL42GjHjf+841aifE8PFF5K
axf17uBvY480rjskeNej2AXvm3bkf7gJiZ7ie4ZfGPHProDdWnxuCM2ukC66z4IQe2nFzn2edTNK
oCj3lqxm2Rny/7RRdEwbqviQG55Iunn45d3r8+v0YcbdTxnvRvGTE6xti7X4uhQ+j/LRWz14X7Lj
+OBNTmIg8lxnYGc2TE/YfUiyx6mWZM4GqG6RMbtkdGlYAK7RkpoGqJf0ejTNCyzMAkD2qrjySYjO
movjQrkeWjiWW1cEGUm4z4NwdZD12h7V5yl21HrYsb/bi8wrWIrH4K77CbvjQBUwpQnlOL5WZAHN
PZvy0i88ZO3gn1rVHjCi/1gyY8tL11npu3pRL+lOvQlHq5XT/VY+EWsfAwnP423kS/n2bnGBXPHD
hb6kwtXI3kZhePx6Of0a8mas7OCChoilXwOw8BmxLDvuy8oz4zmqki7R3peXz3PCI3vrAVoN8D+o
gMmeUVXBKKzYz0lz5KzoVE+Vo0NCbT1+U9YroAxjE3RiSld25X8TQ2ih7K9GRS5S9S3yNYXGMBKa
DwMASPjQ4GdOG0In1Yq4xaKm/9Zt707Yzi4l04sP6A2GlSbGEGpk7oiRpK2iPZAAyyzPEiek30hF
XBc/MYQLxBRyr1TJsSgjEKSfkVkTfX9P7kHdZ8LA4Vy7FVyZkzkZkCYtz5mnsc2cNvkdEyczzVpK
N4Gu47XrtcOZpSMwQw/PbWhwL8HhNma+zMA5eyQk5aD0wKM27ix21AnENqYd4RR12T9S+nc4/zn8
x3jrYwI4DdM8WojeLYsBHzbGVBnnv4x1T9Phaoq/hgRWE9lLWoK/rol3zecXkr2LB6bca+kke6lA
hXepne81PUZcziK+P00uAOGRKM5uJ8yh8uAA1YoxwOrK41Jw/AseAMI9beaZhqVbCfPJyVJcuUvf
BPZB0fWKfYqYuj7yS6mPQ1VwLKxp/O3nmJn7iMn1FpDMHN6A3W4YWu4jUPYzh2r51QE9BbDbgxpq
SAzCxx9AakTbY0+PxJlVHyh7J3W3Srfmry2KJPqcN2WKnpBlbfKOol6wx2SWq8rSkoPTRYB0uxbP
tXvXrS/602axpGQqSe+/mOIPj+QQGKzmJBqk+xPC2iLTrDaT7OZuXqTnyAnvs/kshzNWnLnj4hIF
A1OYB9bU3YfWdwLZ6usA7ocpTmt4378lh+0ZRFH6fpiGl+fDFG80H8S0DVwcxILT1p6zGxP52PNl
/UvWQOc8u7xFblnwohTu4R4gYui3LjeocFvvMzXJY/svUTbXXb3iuYVGieg3ockmelY8PDHkB4Ex
gr3C76znP2ue0Yz7LyYMct6C/fUbIu1KyvKqRooa1mfujotPiyvEoCrops8ZXiSGR5vgRAP+ouqW
2l5e/6oG03/UUTpkqXXY6oTSDdP/ArhOLjwd0cA6DJJtEUONAw5nCFXMxleJW44ZBtJl7xvwVa5U
gaupbOf4FL4CTmAXMQp2JuHJ38sSndEIvSeWTtX5Fnv5BeoBjpgshtu6QXtbpFODX+aqiQHKncN1
BQpkyLsn9omEVKH6MssiWF9M+7o7L3idyG5/JeYMhLnIuNHWPw6lyZWuweIsbVaglBCnOgJGnfWL
abyLHywFVTd+QWdqNa+fI41yTAauKB2e1q+KPWCUNpilVgmjIIQ6DHpUZZ5Gnrk5+Nvq2hXxTdF6
IrM1h6QcGKcYlxIXodve65gh3z6Ne1YDPH7UWxKRWs6oVB4KOdY7uRrGoYl3OLo9ez4oYrXrfcdV
Sg0XYBnUfaq1uptrf5m+uvsQthAkP+JiH4c9sunsmX4PQdid7JHzgiPueaHLo9ARTnhAQ0rP6Ing
4+nu0JbFWconLHLw+2tS259Nf4lsIj8lVehfFjsLEnEknW0+deyGMEPNq0GulHo3qJ6tZGfD3IqB
WplC66nkseHSmZjXauNvPGkbu6O5cg/TTmIWchtoKBzF2EqtWdvnnXYbh2cC94lzAUar2uk4as8x
1aKfJvifyyj1Ojq+S+C39a+jjEch01tdNHK72kBBMBzwoEBqjwbEjAmad4LLESXbvQCugX1ShhJy
CTUsyA5vz/tYXxZdqOfkMAbblzD+p/jWGnrtKWAIeCpPOEoRf0JYLUntN0FRn3+5DzhGxysAfhcx
92NGbqWZVlAtchE2izWADoezyyNGUlRTOo+XnA6Htl1UHbFfYOgmAStR/01Rb6qxFljiLTKqQrJb
VXJAqf6jmR2XXhumzuGP8f3YcKzP3bFV0hbgUHc21S2Idbie/982In/zTR9sPxVPFrFlEMJQ8KQl
AqEa4H7MI5AtwvE1rVTfhQIX4yYGLpKJNkcgOqbAVT/X7LJrBrXiEr1uz7fa8r5XMf50yPz+FMyB
chhLF41MyJN5WkWPwDX/GVKbUUBEDmNa9pKCVOySyrJNpOpSuAvKWZjL/1m3l8c8byZ0B39Aenr9
u/kqKhD3/unY80NyqdMiIs7zPqs3BYTNOkKdojkUg9QyLCOjqFOvkh2OtbqAv0a6TZ9lKNyX8UpF
dQK32YgMg+B/Qf+iwMLAhYm43U4NzOtvl2jM1JzYoE294RCqKDn97JEig+z85oFoXxqZLl4PNYjN
riyTKUGok9Q6D1tzBfHlJJd/OvuISfiWFf1wAUrIOFcy5J+WVyOhjAMM5Pbs6k887cZOlyVvnlyg
2KOEpu5P+RCLv1wtQEOPgV1Tl/kbgXz/1lbPaD3uFeMYtHcpVkrW+OZQ2ZYvRw5G4WejesIncTmW
KSioXZTxVbc+7olchZ4euJXNTk4mor2t8E9hBlCf69nljea8IUyDIsU/l7ejxpN+EanuG8Fhuwuv
7Re1XRWf0tY20BiI9H+rcYkoayEjzV/LH42x3uU61bJUYnm9ih+wgwfw9MP3YXkI6lxEXyhOwC69
fC7lM+YnvKd5rjiqLnlgoEKDtdMnuXiXnH908xe3bqdZp9MfM5LURWuijfGhA5PHAPwJyyLbpK0E
+mHnY2zlrdj9bRpLxkaQDmbWweIPjfDmaL/wFPo9oRou1qkWUFk+nVpTEiQNeE/doEFABV3LLoU/
X3I2g68rA4bfH3zry7oZW2yaT4014jrpGBYpfrCu7PxXx/MRdkvCCUextindA8ZxjeRfDOEseZJH
G9iSTghyZD8AiNOxuOALNQGpMNDSBE/R4iCC7UgG5RM7ZCjrF4ZegD8JFQNhJKwBZbXresLtk9by
CMrmLMpA3Ch1rPsEeoz4dzay5Mneo2TBPjKhP498SEAcx4eEYTokHGTWlqIwQorzZQnmIRHdKKOm
N7b9OYp+fRArckL4LO7Hr3vycrJeinAqugwDFiZgCVt+lZ+WOA/6M/Kv4Wo3AOXsnbAyQ/iz8Rjl
EymMh1mcJ3JgXr6ADdvv1SmqbxZRMPl7GtFcTM/qG+vxgyNKrWkxWeETK7d0T1CzIjFBEtdbFM+k
7ZSh4YV4vyIlWp4U0lwhBK4h9N/3Q+Vnr0UZx70sf1soSWb73sUPzjfw1kPCOsg1pu21TQ/pBz0S
REIOy6n8k72iXOBwiaCERwPtbA8pgyfI1mu7jhmsB56vXS1yggcSgcdaAVnduy0SpkboKSGjK33k
HiNONYvi7/1vldOTf4gFejV/koEA+j++7GaJ8375c9ANfZFefVIQmWNsi1vqxAZxZIhlinbCUIZE
7/DQdKJT1XAlLo9DCr14vMZjbNuxahlbtJyTvE+/sC67/Wibq7RVtAnI0CzNnZFX2+gmXVJP4tbn
3PIoy13JdAX/3lpcVafk8bMBiJvdQzo1SufgTIc9rmjLKs3BIu7A58Nc56bRxXZHJU82vY498Xyg
CVgj0Npd/TfVdzgFd3b8QJp32G3sG5jdzI645H7tRK23NMeDNMTGOSoJ4LnA1RH627qMz81nvyHw
AVDQVZtZja+VcKFrHV2uJTfxy3EWN0c9XIBlyGAlbtFlb+dprBLfGk4fT6+VfpOGrt2HesecKKK1
3BkMTzn2ozEeHoSF9oCFiip+UlX1f3wSK6LlNoQ44YXdEq+WvAPsnkHAjPeMXsPvA3mgdrRwQu7C
ys8OtUFOnnAvKOY3qQ7+T7dXSPEJ9ghWkIO56JUiFNBRPouS6KOEqYsY1/2OePzLCFsonH3tGXNj
VBecECSW2+kNqUq9Ej4ruJ0DwHrjUEmsDtvtjuOlMaTCtqZExOsDap0bLu6Xoc4a9p7kUgWNAlha
/K49BljsIO0M6gCwxDxsvIUNdVwZWwgmrrWpCmQQMQcV/9ms8kfeJ4ibLyMCeg9Qv8j+6CRuJjiH
D+DrezXf3kUC8Mk7ci7EHIbnV0AVVG82pDHnBMlQRAuXPY11TY6B3syVrr+foTEkD68LBpuA6i5y
Jw8qbzUkGwRO5rPPpofjDFgBWAfkW9bFxfyAiJoF1MVIZKf9CciRc72KwlQ1zHvpwL+PCULOM4Xq
g3C5daR4lS7hW9JCgzYxsnkyxqv0NW5O/AbwBMYFAmb+X4wxvZtOt8BhmcVghMyKzqbxLrD/iOlQ
euwbqLjF3rndsraoH1kIy200DAMB2t5m4n70QBrquKgv66+qarVzvnoNZnihZfAGXqeWdfRY2bba
oLZoT7AQeMkwtPYxxMBCpTbZ17ioPaEV47GmQyrhr+9/DcW9p+HdnKk8xljwcZy9EIM6n1uoLnzN
+0wq9BQ6ambHh+JxyHHGXTxe9pUHz/GGUTQp5wufcVsTzukVO4N8mqL3WORdv7ArG4MMLLk/453b
krE1fX+dQjWBax9Ou77hz8Lnr7c1Alf5yAtk2FZ5Yo9DEB79+pUDPboec1E6tuAc719acUmqG3Qz
pzn7syfUE2tjzivhLhTh/4fcIMpC7UzvPdrAFWs7xWwK4VdgmzpwLo5LDCfc9cPq+NdhZgTe8CW0
hPpoYzzxz9zt/ERT2NwMheGTGKv5SKGDj0V2bSWwempJHzSxVFMuzszJU5YlLqoEVvLK7HMRqVMB
UpPYzavTL/0Mb+g4UJsopBP9mYOZJpgTfSOL1x6Tpc4LA5lHa5y65DIWXqeTIq6iOZezfQvF84Qw
jscP8znjC8zez9cTpTjDztq5TiGd1xxEIXfD7ctLWcy9FRgZQG7OJUp4bZ0TLpwf92dD2nlgD1XO
/8fxLEys2gKiDwtSsp6Y2cf1fBZryks+zmuFvXb0YRCn94AJeILNvESqVdjcAScUdHsf/Bdrr2cZ
RijtRjCWKsdfh2l10qNfSYj7hbGxdDTpZbCYIWkVOOvcj65aH2krNdt/RfSwYpbc1ng9GtFYC2XX
QmWey67/r4l9klJatDkB9Kpo90f65pqyGCxIMESw18pXEDzDEb3ts4A4adp9gA8oG+QOyQ+m1PQ+
xQOMiBg+gYnjosVbqZRqoaJyiR4ocz3iHIn+8QDXeznXFT15W6vU2YZow0KNUE8Nx1w8kpoD4bFp
8ck+9xZT+wS6ITNN72hYwoNnMsGpMeboEBgX/kFVj0HD3PckiINo5CJitwE7Nj2EHQOjPfkcSIFO
Qtjrw2dPcJFhwtGate8Jmw9Q5Jg7CxcZ+H+fo22RWXT0VNqN1AoUDNNyzjVFIYkGt/3nhB+/ieki
8pal5YTgINevUerCzmkoNiALEdHq4Fp1rL1XnhyuoG9XxzdAKDIThmdw5DopEOjrkYJqr1DyMWtw
DsISaAMxx3Z9T45ODUbKzu/NMIWixUS16bh022EuVdiB6v2RFFR1ExjBLqa0zthAtsV9u0pLsb6T
7fUJ3+B66owHUlCIqTKkSoaiTbH84oPJmiB6zji8xy8OwLZd+F8UFwnNZyHSWZiKh+fBSbkyrQUt
Kolcl2Kdz7LIBApVzgVJPWlFfF4tQHboPprSvMKzg4A4GtaiJYHV4wqvPKkgfwt9BrGSxHh0iCG4
W4pVqIbvcsnkOqGwex7PuYo3mIVQmjV6kUjvh1Y70Xx6yhdbtIoktYXAPWtV3PcZTyB9woSQd7Jw
0KTbrxMeFk/fQTU5hwqRkNkClIbKGcwZNXylPaBPX2q1/i2lHk9iaRcxz0u1SnDQjtQwa1XjaAvJ
K8Bk3Uh0amdLEUl7q/eajI1U58OFlVxg28ItJPaXo15Pc0HgW6kFmYN7rHOt9RqMuwqN+SmJ2OzA
XaogP0LdmmQj4Ugiv7Wmt4kwfeBPMwTHT7AVrljwQWw/xLMHrTPN3XXplTrYVUfXbKrUSYKmRoFw
VNW21jkY/8U/kQFX04ieY0bhyl85DPt3fRH7TIOrVz1hdXjESynoLqkPqqhMUcElGgXDp260SIYN
E0yZREbWTvzDJPFfeQ7Xrs63wELEHq0X9P6S9agkQuVt+T/X0Zn3zSa8tmvZmPA85miHz0ZLFOt5
1GL6yK18el0qwh7hmQRUfbwKDxOSnN3UkwWem3RUpHf1H6jI8aDRXRYRAFu5AM+ORyegCOFoceVp
4SOknYSdNIz60Wg+bLdwAgZhMsqBlcZ9i6ROZfY+Dz5UQouXNfsGCUizea97xOx4LCcUdhuECNwt
xj2ZOKrXkAF4Tyf19vNvu3a1fzp22YeZFbnZoKrMGQYetBgSBYInyZlgqs+RQb+tM0qsWpWJMQm/
0xA8jgL5HhtOtTakvaDZm1s3Qf5IB8dmj2Kgobxlpj6zR+P7sZeEd5z8Txf1RXxK9TKaxASXIF44
3HEWC+mcFexMEIiRyEdxVjOzzdfzSblbYZhgaLMcuiwpNMt0KdexdJkXByTmR/47eZPhgFLuittq
iIpp2qnXSTUm1sraaEpJHUDZct5fkxFgUFU4rpHQs78DunURGqPfZLQACN5sQnK8kGTp/Twax6o9
nwAnvzcv7NIrRSG51f/GDCMwhAQPSM4SFQMOMbejBmygAaP62VN8CSOPexrGjRk7Fu8ujn8J9at7
oDg8aeVPgSU3er6jwNemRLWXXLk+nDfb4zrrU8Ir/Yl7ytlxcg51TImVHgEQgU9L+FQmK9lKx3Hp
fUqMX3bosLCYbz3560v80xxqaY0GrDfXTwLZUhs1n3VyFiPvCptt48U3CrsyYVwjChaBGJV8mMgU
CN3f9Yv7VrUnOLiKcUent7yIVjuFW5KQFUpm5BSVyj5mgYf2fWDgrz4HOheUTzwW6CqqhsUuDdqM
7Nhq2ytY83Hxx7a9rqH8kA9IqB0Xy7SihZbLnS4n2Sg/eQhgX43SRvmcJYiZRHZZm8SsUvz+z1jA
zt4mrvaFlTKahDWbzvlRxLzvy7liovPjGdN7CBRw0yU1o+UJCYYrvjCbs5x7vK1VgejJ0hSBp2RG
qePpq1mtylytrfdgrl6AGdeGfy0FaD03VolLmxIOc8pN3pwWl/+88bZYVDCLjTwnHl20eMj+g9Ld
Q8pXLgBKIPQ4f/I82iLm2BeowblxQb86zrFCPtOHp+SlqP+UbaKA3xEUTMrno7d+StoEBQNe2iVq
QHQbxmqeAn0bL22QN4GZN1mM07qQJTLE/R4l+cy3t4y1UUz1mu7EEB5dhhstEgb6usj/xu+K01cu
kNDjtHlbfICUGTaI9EuEYRc2ncAQrTBLjPiWqjeb07rCZwFvLaC+oYA4fGfQbjeQAYfIdRCyWfir
hYNOjYc0pBhKm3SmysordXp5U/Zv0jXY475mgVAhjF317fLu0u5Ym+x98WBwQ7O50zPXXAKbNQ9/
mVp2hkBA0462DGbvQX80JXG+TtCBsdr0JJn0WJkCTM4NkPGmzwLpCfMQARqCKDA2cQbwHX5GODeS
nDPldOm+5Q88D6Ji1z3RFXAG2/VWXRsEIEYX+5H/A3rCt76ayGKivO4ObdmxmvF3M/KeKm4UIpVl
3+5ARRbxpaR93ZzAUxWwiC/uL7U+QAk6A97dYWuQnWZgaDnrr+tWycQ+7nFZzsir5KCKWM3iekJP
9ygpKaI3bq57r7e/GU607g7NKUMbo/O12ihtKAyyDkoZ1pS+B5t50kTLAQeTlJlmSgYEbp3TpKzS
VU3k7BKO9uk4D2zxEKJrxWQ5etG1m6w8GP0Vr/q1QbblD/uVgNt4QH4+G/MY0iYwvlPVn57+V/6a
WdqzVxwXnWavrbbD2bNcmRynXHC/5/tbE1Foyxcdiy4/Xpj/ALysFfzuMQDgWpgTPB70R6VyoXeb
1P483Xw+/BY/Su3LdL2GouEN42Zx2BHw3SNdNQkX6gVsMGpROkDuxc0R6OLVYP8uJmTNhUeMx13a
0/Z4mlnrWOqt1BTPgNNW0wRVOtbT3uMplB/QqjHxKsIokjZ3lP914RISsrZJPgjHCll1sC3KBusx
Baoz9rvcGM7aoDFqXKirWwsOnRpPHuFgZyGqYAw9mvgyBL/aJu/qXQh8rSOa+R1/gBcVZv7z23i9
dwrsVhbX3iMGy2nAFf3jYDdkGC3nEJh8rDOVsmhWFSAxpMg0l3T+zfa+rlHVbaSwvs3EwujpNz6C
eDBX/55plpFXp8gKb+vYaPofFyTvcdT4aR4OHEJNrsD0J3JpTX8DID3p5oqydBkn2M/BCUgTnBHv
HZqy2D+5qDuOUKREcydeZcu9xON7hy5+aAMNwK852FcsnVXIycsCV95CKv1rujq/HNQUgX2thKjf
mTCyPTeY39T/Wd8iYoarf9VY0PCo08pZdYg4blQp4ObjPMFAkDx4fl1fptcenarzImrCbOCsyxsU
bd/tjI5GoZz/WsJ2zq6H/LADPzR1QOXrj5HCu0jzhnasCOWSrADFd+2JauxU+n0hng0POQxZBqcu
zGCM0VazF/4BVfxh1cN6TNLzjQ9fMnFKcjBlSmykgFaGR4gRjus/oiact/zLz0YfcUOCzAaBdAhH
7Q+Z+WBu29uBdYzkgfXb56JIBEtfAnL3lQ5VFXhKNskl5VVtUvTYGZWYiP+824A8S1igHm9KiA7Y
RC437tuj/2DfdhDrt7ygiy7vxGYiFng+8K6wuHiUharBN67Vy0aXOlRO34faJgeOEU+PCUp7kcZK
sY8TeaFfrwLN+nRuRIySK+5T81Xx2RvqyDWjrRMw/5HbVyTsFdtF867FjrSGGb7G46SYB/Fhy9mH
FeNr/Ie7mAZsLYz+cIMZi7pydwR9jz+WqYBTS5/aD9H2Ti2gtHCkrt+NRwY2k0m4bwLLghV2utdv
LBCD2yTdM3+Nr3Bk4Z9TvUa6jrCEFv6JfcwQlqmb/Rw2Zqqy7SsWZNn6dWsKx5RTBeY2yO/7RTYd
BwADU8wZRtRfHM81oImx+G3X9j6TEdJFM9efikBN2EDR9NpYUzaZclpS1agMnZQ8h/k6ueRmlw8a
fw77lNAROvsHjm7rEtTLA5HVd4jjH7oakOJqexCY8remU0voXg5t1diTvTTKME5OtZL9MDjqxxMu
3EbB0qD8x8ZD+lS/w+5EVUoVuZa6ClkPgdo5MLjSsRWe3ko+aCGkZNRZb1LFpVo6RQPG6sazoajD
PmZn3ecX14qc5r42yIC5N2vQm5RSUah8Dtpp58+XPkTOaMK5WbL4I2uDfQSL6KZvZRnqvvkQZFxf
8cBxkuZa03IIHTolQAQNPc9oTwHIAVHrS9hlLkfsAQNLq7bqGPSbF7nASlV0+bqeIKa2qYd/eRw2
9Kgz7juVLkA6U0CKzHxOtuybleH3wM1YwY1VjtEaTTYtf/SArbob/rB+GyNdOe+PxDUFC0avqTgz
GBJU6YkG85J3rWMQISTK2vbeWsjOHWco3FrDuGsm94Knp4AQq7uT5SPtqWkej4iBtmflA/zjMaNP
Ax5U+jIndOpKxFi07/vw40r68mhfDyfRcWxqPUPo7H7kdF/bU8POCbi0Wga3qPX8nRmSYJp4dS5M
Q0OwzGfC19dBLBdZYlaADbw+q85TwRP9pF1uLgRPptzQDkKITkFu8fOsAWqu5seJ0zOVocvUwlU4
bKpzB64OMYKAZVp0fYO6ctZX85wpYq26rIBzQPNVz0Oy+/9teYPfOebSGkFbbr/0TCDNWcvml4Lo
g1Y+mKdOr1+kAjy26AduPr3f6QlWwn26WPHLl7SUuePtuybFqS2lJTkAuh3HGbtxjwpaZCiJFv7N
Y40orPlYUpRJ4RkjyEyVSI3U0wnX7ZlbqxigNBIXr3/Q2+XOY0sM2LjN/68X2YpH1h4HHB4asJJ0
GKYsSNKhVV50mVlomvNTLnhZVez56PNwg/4r9OtwUs/P7ykgPod+r2dH5u0g0wFa4HYFuWEd4EDI
8UBhJhvQeqI4d6Q1hmpSoDZ298M71LFJrtbKeiO+2ikKsS1DPsmXtISB0v2dW5Y06TVJwRSXTDVN
Fq84fY/9SG44x98qWTZeilbaySGDoi7yimedVSXltHZKO0o3iC2jV9FWKoa2ybpeYTHRew26D1tz
b8O0iHZFHgWzyMAUMFLbnukAQUNjU4mzOxIK4wQ8KJK+LLHV34mxaW9fE/NyPBpPF59tKJs14jas
65U5qbPPZD5x9Fjnv0bny79FvFQoM11GLM2sl16MP0P45yLg3OckDWCtrsXVnQOSMBVDuToIcWzm
VXJbil3K3aVrPdXG95wmJ2vG9GNr50rAy9XHwdPuwxi/9ttR0YKWFpCY07sUybsB6KOI+ri7jQNl
yt0tZNQVpDBackXwaZlMYs6B7NEgJ5scPSMZC/Eb0MDYC8NmDZPA2DFh0bpAmqaFevgQRA15hgtH
wRau09v0Uv8y72GG/9VSmaa09/sHJAeHEdIcQenDDgYC8mxbw9NKHu2W3PDIirMowpW+edmG7SGW
DXSBzSpz95kgXSS5v9QT8NQRg2yQKL833lhI1WKQ0tCs4YwtpeWVyDuvlPG26gJ94gp0AM4T3iKK
Rvc39A2I/JgfokFxRaKnWwbl6iaU9BN2hMx7yZyhOicjiq+pMQ0KFGuQYcPMkWxYFhvuwxKwM+qZ
mfkqd7SUqin4TX632NKeUm5NLzJLpt0gv+tcKokMpAAQNvHKoTmYRCSSzjAH0BV6vDGisenELwA4
xefGzF0ZDwdLn0jPW2HFwLVFs33ktBXqdyWTIzfBloWpOTABTtW3IQ5rIO6ikl1Zsf5jHO5tZIEx
TL+Z6ewF5ObQH/MxYYfBF3KOTH39bTr8gduSVjEKx6buTeY9ig+lho7Dt0rjd5tDYzhUPSTcbYnf
eBPTeBrYlZ55dTR6Q3hJkRKQtFWOQibQIcC9d4FbcWP7tQgMfVBUE94Nf+mZI5GeQNnBtutLeRWk
gZeOWfce1O7jNT1M/4CSZ78cJSmsscRXSjSL1ODEryegTvVDpdPVRAArxkyGClvsxM+FwokhHscd
1EpezwdcxfzuV7oNRcvflrzDKq2mm/HVDUGi2+yaPeQi7YPv65r55Ccbt2fUWulmm5hs8d7yyxyC
IP0EThlO113fKE0jkmXO7+iD+WxqrSBzkUDzZYRwLTa6FZ1d8tfhLfCUr5IAhuLO+N21LmAJ/Wig
yym6C0JFwFtbV3Nws9lcxMMC6Oe3O3SQfe1WsMSgSl/JXZIctu8gJpd+PyWhzKAGZ0sGdk/ftFHJ
MRqNsW75+wblQxWzbNKG4llNq5sAG611ilbDxKXrkig735LPiq5rey/xg7By4HNWWcCJGUVfkcXb
UypowvctHlwoL6tdNMcsxlhDQ1GgV9OBbVMIIl/5oE3s6JTGwGmvxF0AwKNswZo9WIWQB0B5P2/b
AMFgitkUZ+V7t7Hf2rJZ7rc8TYAsL8KTFWY4H8efDkoGU8wm6/AbxIxFhBxALVDUhmGSVUfUOtzt
YmOvoYxMMbV4//GV3Ak1ppwyCi8vCsXfMNSm3lxY+1Cd4fxwguS8KYkh6BbVg5EP3GdHqZXjoT1x
r8smDZDq1PmCW7yNSS+oEy/ZSoyQHd8gFHuL0PQ/B+yH6zaVR40d9/UalrlS+DlOMAD2JGKaIXrB
DmOLrzbuQLMJgyAdvAj++qMUUW+6NDKKLpgaCZUfO0hqvr/UOSbCT2sDdQx6rE4KknV4CykUswdP
H7KrZjUH1DDSQ3fiduDq64TVGBhNatQU0OAYTF7w5H2sDUvZnjdlxZbzciRGclNUcYVI0kRVUyHX
oY4+y9LVhSz59n1rGd+9WgZM0HoICeYIsfIoX5gvDOYyugmXYQ02rKsLTdheKAIKRr3+wyyOwmG0
z2byW67PjihIBD/tFdxEZkIobGNv2aGj9fKrE+cGrCDjmHKpZPW3m9FK/WMIAy3oeJh4teaVxLxx
vP44u4J0wbK6o0uT3yLiJVhaiq2QlrQaFB9RfQkYTkFCtoVVzXNSOPf1khA1uH0fga/51zMjPP7j
I7rF+ilL0GW4ZUjxczizHFSpkvCRyNSIQb6ylWal0i/nQFRzyY1ry90re7kowJ8KZo8WCOzn2VBH
xfvSCPsWXWs9hXTUgIQfngbdlIMZKBfXRgmu89CwMRhmy1y4Zrbe1mUGCa8G4zI5EpjYnhLi/wS1
XJwLuDPl1gV0H/4KAY1xGcG/jAY2hlVMX9QTGmalhDRp4twUovQznN0tvHeenp6JtNcC9VsaDQLM
sOh/8aaMeu58q/fjlpogxRcQQWcFbUmBvgraF6Mgf+5X57lJYzCxC5DqV9K+Em0vWCKqxU19bYPc
qDyapJJx1zv61EoU81RP2DqzdN/uAX4zZLxDbCmxVQTTz4L5dBH4brQJYYP/VUUymKZvIXj6YaBd
t3sRex5Czq9l6V223HSGWxyhgAw6WZ+15p0htjTcdMWYQuch2jol4Ig357L4i+tXl8wU9jHkS/Vb
hgfdG0MbHUmB5XdSqsMpqv1y8+KQ8f/cLK40gMBvvOQ2Qx8hpJ6y0JBHx77JBAdo2tr/p6Muceg+
e83usCgfBi/rB4zeh8WamWsdaeKwqBoal3/qDHWUFHp5smrJKkoNmM5v61tH4+BU+mN8dr1tloNt
tDz5S3RDrudnb7TTXyFuMAs3GHifPrcPw5xqJDsQ+rGL32610MeRqoj5zXlkxbLQ4gcFmbNcCgdY
5P1Pa0RwweBCHDQAzlhIlF8jAASu0kbzb4z1eVKyzU3x9OK8jirFECyWTDbfLL5Rwsm+S/xL6kWA
Qy8i8Y2WKxLb5pAHJVRuG+wUdMv8ZnNYDgmWzLmSPBZpf5ZsUVuC6cFBWR7lLsW6ecjd0k8yN7MP
LQT/z678+P8Osx7OBSscK1P0hl+BYhtJx5u20f5Bz04ePcTlA8KwsoOIwB9m5fYM2FWL0h1/EJnM
LSe3seept737rXKyKlDH/b5HUtFHyiJisPx/oReKaxuVAIPVKpqIp+DiOw20US8T1q8Ph0bBsSaB
SpAUv85YR+COcH+NnF/Bl/iY7c8pGVqEFaxUFpFMW8p0H9bNHdPue9+eOt2yveVJy88Pj5NvbYzp
hc8Bcpo6MKPKG9j5MOGhKQXqvWTFKj0Kkek2jDLoelSW0QWkv85MDLakZ8IPaCZZ/s9Y+pEUXvx+
1tP2QTgrOnMcuEoZBnly3WoIeOH9DyexayFlT4fI/iE/u2BN7opyoLlIb+LuE+NNaQaGFmRL5VrM
xo7pb++UzjESsghdtsB9TnZo8Pp27/7pLgXckyzkPsC7DBhEIMpx2EjkF09h78o+uzQjJ1E/wAvy
oHZTDFHWKfWD7pjh/WA2fmZi2caI/pMi5CK3N0bhaMZOEyNtQhRO3o+XuZohZFNn+vUvfENQ04Na
bXkA+CHGuQUWdSjlnIlVGZgee6RknoIwlykq3kByuwYHfJiwhm/SkgA4oFLtz/B0Wmz/2XNu6Dlm
jXYoziX9p0VfJwdp+yT6hpV3RTK32lJlsCLWwCRdX7pReXF51abYgO4oP40JoNtnUsa4wmhNx59T
c8hiNESIdb/foiUa+h2CNWmiKtKzQ4FOPH4O3F/ffGzjqK4unWKRHFceFDrITmHYI9p46nYJ5EKl
DHYwI3uqqT3aaWncjbZAtjcMdOCGGqNWP21jH85cxvC0jeOUhSTtt+s1Kfd8wU3jju8Py859/YdA
3KiJgQOIvKGLbP0RtSSBg+eccYJT3LT7+zYdk+0D3T15nW87lxl8dyjIsS3CUykopyh0P2qwIHCr
dg1n9OFACZ9KO1V0PMDkCTW+JpNWvbQv2uMa/rJdLLJ+7tbTI8Hb/8e7nZseAD2br5qB/FFdeX9f
VdtO6Z8jyRDDB/OieimOqFBzTup0/qWM7hn9NtA9r+O3CCj8DXkVW8EzZ79DKRkwqnBXBSdwruv8
glZXPdxWw3FmrXa8gOJ4NhIzfJT747IjqKZg2E9stRKk9KWGoJCLHIapz1s+99pvSUfDrNL1asY9
OOPxva+swhvQAjl4mi1w0z0SX7nozXLZ43Nkd1szzo+wegt3c9P/xlHHUxRr6kXmigpPrtYGAPlM
AOKbEq/q6n1IHs3NBYrrduJtNKKTeKD9v28mr8mI330vXZt+oJw2XoCiaBAHt1lH9GR6IrKV8h/i
rTMnLSDySp1mOQMiHa6a3fB8fquUUuOm8lIAQcev75xv4mpNBenMIydZ8wbwajuYPybB7TVuFP9W
JeliGLr/AYSfNOXUiXnh+A8JgTP+z+YGs1IRqJocpizKe7Fea7Yfh7Rdc//6mEO5WsQvNehIgHCc
ncALND3Zo1M5vdCCgogWDU/LM3GsPPqxPAuY2oW8Wl3sIj2ZGg57tCxGum4CVnIPyGDsnIyXOb9I
XSFsrZ7pnk80CSCdIbFcmPKNK0a21jdXAA6nIXRYqaTVwpmEtnKSFHmCYKJEU5oh7RfimnQnU4wS
ItwUYjOPzIlLWhcjgAgKJOA+5VxEzaquv1Et5VPdgcN7byKgrLaZC/3feelaKR5E57TouaEFSlpB
IC0niSVbHv63liYWFV7lH6t6WTrV6TifvPWLJEQnS+8lt9/tCe75rCyJXq5eUoFV4RYCO+FV1Ytq
eFHKIHdJsar+xytj5WAElhQrHTdLb9bSbuOJY6Z1qxQoF2fNlCQoj2tFa7DoswRzlUH1V6scOgsr
mD3Yu30tjQusUB/QMlh5be1WxTjF0N/+U2jgMKZqbXEJK/B137/YOUHv2Me1tefwAHx0m+WqFNAz
j9AaapPFMHlAQcr3wLbnkFvlr9WOn5JoCnRdj9rUcPgX9L/dFgz6ewEblhvbEiCZsgZQvkgTyyjR
MjBOY6sjc51KgQWUT3AVqf69Kea1U3giuFOZwLNJ8rbx3g7bYTuMh7s6EEn4Oos2HXbuo1ckvhyL
aD9UERAcUwbLXMaamiJM3WKx69AIlAkx7wM1XhDcPWHgcl84uguJSnuTysIEcV/wopKFvi4+xVLg
ST9ThngkOZCaEWD2J66xVKWiG3IScfdCXkFFmDQx48qp8/LtKxI0JvuHSsbWzlaX9BPyk5TRC5eY
6KcqlTMixWDWO8x/Jar3LwdNb+LDfpPldF6HH/NEPLoUqOSb12c7Z/xwQX2sjiLoHDPldrSsQ8Km
fwer3R3dn0o/7vtGXN+kNQ+0iWYXZob6O+BZa+fe/PIyq+zQItK2Z422LRt9Y+xMgrz1RvV0+ZzF
BnAIwjDRnpRJKpTZ9t9xx1aGZmpQg4aa5FpRNynnHeuC3pMnzNEXZCesVyxRc5u10DgN1x7liQKJ
T3UW7LKDJnIzFqVzEdWafK3MgP20Xoa0yLfEUV2rfDN2VY5DhxyhGRu9oL9Ede1jY2CvXB1bhKGK
pWrK7aM5V8232y7PgD5SLvNOkeXfmriUS85+bw6M+wqVDYenunUN157Gc2Y46OFVEiV2r36bkdvS
eE+vR92yXrsdIMw3qTvaenqS62s+ODmtJzbDaaBdHOjXTctHvAMiIpJEw8XtRNzXj6hXgx24HeN7
U8MjWmrTMj5VNeAIQi9W+zIXGjySH9iobcLJDQxnz/lldu247/rctUxx0YEGFOt8pO0lBKrO1/xd
VRVYuH7MTrCd/fnPTt+T2JQgdH85K/7KZNBjVrRP35EJrVOi6Cbb0GBInqlMogRFO7Vz5KuyaIG8
42zdm5gpm7KZbX1CVbulSB9r/78EyWzKI77jd8FxL9PWjukuFVMH69VcQYP+p3FfiU9hvyCbWOdn
Te/jp2nSuizxXy4cw8gdL87a9Thzss7np7ROzegqKIdFiueGgyRy2Eyi9GnKVJVt0OgNRt8BExEq
DVzUgyuAN4CqPEn2dKfTJuK905qK41+MLP+2tXSL2HVgi5ZCaBZ9MoCZHHtRvbYF8Ybn7/069cDd
a08F7mZchdyOp3Iue8NnwFxk55svaAIQCYpZK1iYKr9HjO7rIpVbmFLak0r6ebyU7bVQlNP6XLgV
VyVzdVOK0ibhZK9TH+EYaAlpIw/5MApPkOBGI1T4WegMkhMLtivIqQWY+8nKmYK9wpuHaeSXLWiB
aewa8DA7nX1vqV9ZhLQCpi1KxUzNpmg68VpSb1UaTx5xMPPBCrICsIrqNbYqWp8+FuFZvCw3oVBF
VhnIjD+efvJODXj8PYClLyZGze6Kg4QVY8eByJZEgdXfW3vIcsIXkeRq/7egQ+dnDNqBRsnIFLPP
nWtuChar89mR6CQwiYHse5beUSw1iPpiQCzlgw8K/mZpRfv7oWmOTUbtVeiwUsIyvX5X/bKoVVWY
ECDvuJoae/kXq1b9bMiyamFAfrfZsn2z1OyjD7QRsw9mz+sT5c/pKRSNWOMFkyXTvWxHz2yDWtSq
RkYBA2qmaSf0MQtfZAs+5j399Tc9o3eIhFlgRWY1LG5I6l7AFZwTnNW9d05hWBFXmZhbToi4DreA
ViFLnSqQyWYzGyu25x25AbB2slygd7hO4ItJ/IoRRj0aq007FfgsW9QHgSF9BKpuAzCFrRaWB0XD
F+sUTime6jShFjDxmg3GV8r8/VnntUpvqP/dtbJLpbNjcCXdxaP/VLMg+v/zI4iS7tJUqyL60o5g
ggnWj+RfgdH3rb2F76cDSnXjVY5QW7rNqsSCNJdGhbK+ox5+kGtVkx3SWi4w81JFBozJgl7MzSvd
W70I5eVUbhkPyuwVGT7PbGNhOi1TXR++PyRpBIEijuPTGbuJ7cPXeUdOmpJDdBLRRlsFLh294BWa
BriBbKHvRYEtjCZsM6T8W69Cdz1ngnhGx165IiNBK1nHb4GJaBvTkfO3zZHgugFSTYWp0T/jL9gl
9zJHKEJD2Ju5R1LSeLCzqVPrrRYl08//zIjeubn/7FNYvzod1KhEUWq59ylb6D6kR9vmI+zgwOOa
yi+T5+stJ5pctv0+gWBtmwfpJwlNdYxzSB9dPa8AcM/LkOO1O8WbUtVJGJixFWCDvu9s/0yc3Q6r
nc05SXLmMlmwPjhbxn7QlGlKmn2AZ8p7QimKjsoaOu6zAxrdzDIDV+96BZj+URZU+ZRTZ+I52ko5
pFQLlC6MpFDuJ9OQ54kiZ//HQYUB6ShnzBdyr7ozeWerhCfHc5Jr/UjeNOk3sVoA7b+caBf3FAXr
VeriLWwpFKW1Nbn6w6TP84GJ1ezvxD/MIx+dmitrG2lMr9thKUD3F7VVotm5VSOZtjOS+1RlBd40
VI8Kpprj6mrLV31pA0qfo6KrBsyNP/TDkhM/bd/ZWyZ8jYOQZcSKqjIi8+uvKfNwv9Qe4ocQR6wX
JDAwsgnFo/5jHWtoY9+7gyycTmdbM5cvZvCazUzkeyKN6N1T17bQvIo8zXgONeKn+denem0KJOhf
yMk2Gi06V5A1nynZ5Td+hKMXNxi1CB06573kUIsDP5vd9KYRsr4UAFH7KKJW93V3R90yGXzWjo3U
EP0WNNSaOuRQPQGppCN2gQ2ZnzDj4O35c66ObC3Xa4TKYVifPjv22YSBRrqvo87RkQiP2BZeMv7A
MYCpr88bmcJXCWrQ2ysUvzQAOW87nKMHoC4ZFRByEIP24m8Nx40KjGS7Dhb9pQjiguPAgNweLYP3
trIfwticIXEM6jyCqhSc/HEu8NVIrbwrzi23CEreDIBgfUIluKdYoHNvWwoSW4TFCnOHv21Nwt3b
JUqUY19mxFjAVA+bA5PRjIAhii/3HB7Ei/wuvE7DTVItlb5k+Wt6rcztjkebgIDF0HW8rw+VTSG7
GdekoAr6CAnclFI3V28Fuwc706uuCXgpF62Fk/KAdpl6jzxUYOFZrsg/ImUOCqUQOEGlqkhY+UjY
17MaOhmd93DZnWl8fE1M0rlieFOAmtc2c67eBFM3A5cZ0nOAtd90fV4jccexUo2YMRjKxtJlpNLo
f7+9aDmm3ZuV8uUMecAwGmOYwlJUmM2BSjYfsbojFJ1YQCBYVGY08BbohzpJ/yMb2L1IG7rPw0SM
PZbJ+ta10tBQrW/2zP8BoJbifE9CYL8mahwXA7SfYYG6aRCc7t4+DFtHGyG4D6KtUPzLdN6bRx13
30loZlg9lMcWEYjiJfbV8QYlj5f51WcpWRAmzCa7PPeY8di6/LbFXHvL7pUmpP5k/1O7yzS6wKMq
N+F//C8wgKujabcKiMlusEaRE96pl4VN51eJN8wMn5FTd/eakq+KahYXA91Qkd0hy3HFQ2iKUzq/
fs+k/23+xyAQ3R8e8es4qK9BEqU1AOZi6as87mtnSEShF5XCzxsp323XvYVnC2Jgsth4BHq6gEpr
UwnwhMxaWWbDiRYZegJs62LHOfB+9Bic9PbrzmsYOzSrYXYXbgjm63O3n94saGYXVQnko3vFgCiF
vSkWFUe1FW2tUj/pDNIbBVe09owKfZOWYCsZgiu+78cGiqDb5tww3ISSs+LjP/nu8fv72oVJV69G
8vLTNq553OUUcL/1GiZdixwAE2u5TVaBRyngQFDV6RjAj7kO1tQ8mkUr7xwEdJklM5jWxk97iSAq
JNyRVgNrY3L1+qkV0bCBfSb2ytBZTjNvgJtRR72+J6DuHGZAwu5NqgdmSnnpBErQoOudg6Iata5K
uMDCWpxIVIWTOTrWnxlhuzGzitAnuCixaxoS1qPkFVwcMh6zdjcyJSr0WEGmni+JwBf/T8NwwL0x
a5v2cDQGSTV4Wr9bcsZb9NwVpbaE7AmZ8cPs3rWCmouWUtiXDPaZNjIjjqgUZSVpN3yIWbnFKEaJ
oFbJB/sSl+1eoueQpTTpYQ6G4sWRf2dLp7qZgppv1s5HaXJcuSzc4DmLvVjIfwnm53L5sbEPymYm
k5uTqjwheK2bokWJKDd0kEWZwhmTTPj+9Mva6wlIj8/XsfD0+WCTiAnWBWCfoHNU+QdHg+PcTRE5
X09EJMFybzY8r71iPrFdf3dLEipMj2AoQISksDaVa5TD0qQ3oH/kD5+ijoMXeJtuc/fL0vOLAG89
RktIbmKTtLC672i2DHRTxe0v96qe5mBHGJcLmzm6nUeMbSc8Fjl0MRsSrCJhxKCxMzAFd/lDYtZU
I/adpeQ1mKmaQO4ACA8cyBR5YxunjjmoVag2cgWe267IxgfG9cwR+mb94q1ifSjT2XOvzuwJs6+G
PxVLrDVoHvhgPTLjWOK75mJGtOjpZUDjm0JCB6yxadriHqBNE4KgrB97mruPDoIav/NhAX0Dmxsp
5y8M/OkC2lDEMio+oW2s6nUPoU745oCTHYlGQPQD2rkEzHimHRIJr8KqShSS9+30tWOVywRq0fBe
yQuvIDU3baWH17UHOaK96WjilLramXia9bim2yaIlfK1gIyQtlSToWIgpHnArLjsIb0G2+hDigYb
yDz8rsn2z2BjSaOEGNW2SItMtb7jnXo4w01q7dZYxjZk4YaPukja3hxjh2GjY0MoOg+bohpBJ7ZX
beePfJJZFGW38yih/JMnhUFDf9C05pj+MGirkbZPUleKtvvNHjt4EfKwfddrkdJrLyUfpAaUtL5G
4r4TdhG0o6hImrFrwZggUYcjGooQ9M5BxcSOsySt7ddlht7PybPeBttrIG3qRUWhAbCYQ7joD6El
19E9vEUxhEA+Lr1q3NcZ+Lloq+ejeLNVXsXSRikQLpmttJ+2i75Nu/rLD2w9eRkt9qjAHJQIHtLu
GwHndbW5VB7PmeOFWlPViJ8VB8AFASOSazarZIQx0W0isJ+aKfDdOs5BHYErfcfjxD/GTVKntXVT
X1JQ8Oth1H6NW2iazc0/mVlNM3eIebaYqW1MOqg2qQHPxZO9Pw3xTnSCFEmHB1PthIvFYhJADsGV
7opst5y3xvte/wVyHv+lPYgCrWfRVgeh1E3ux7wec7D3S6Nq3UcloTvY6yy974Pm8YghIQrS7fMZ
yEPW6NYpWoWanCWFsMPtlMWfXFmKzbgfZJQw4LapkvsbCZDqsTs7874xF/IrjS+ZOka10ESVQ1Mu
2r4BMnQokBonayXS+ut+C0ybCkxTd3/3stlm1e3q6h3ANubRVxPZpAAXONETuzhNScUetVForLxQ
GfXnBxSuUzhejk9U+GSAVvfPGqRnOO4a9+VEnPisoegUgUeTkTSj3uwnHttxppma/93xEiYUIGog
1YfmNxP35OD1G9fB2YXeRdb6Eg9/uKucCyvb3+xUHuIzyi4ubgVV3dVzkUyujbRcg83u5djEKlt2
urs9VRPBAT+hID0nGwXwnwEwlBbdN18rxm9N/ICRTxBJ3JZDSXdwq/b2urPFn2F6u/+VUDQb4T/g
OFzqAPmmXnMmtH96/Azmrf1Vl5EvDuU6Kqi2PSGqI1ZkDOiXacK2fkwsQ3ahwVZeGuvhFXi7RkF4
H3Vogv48zlMiwZCnX6GgTPMk9yauA19gSMzhsikHYOB52ldAoHKd38urFGi9nQ9I3t1GoaGl3S7l
FZcokndiiMkp64aPj+ZABMlxUCVPpY5un7+Of2dFEoYkO32rtALIDmD86O6vDc48DXZfaGPg57OE
Zd7h+phsUS2Lr55xyQfLN7T5OLwdEsTywbPBxXz64XDoW13FAZJfDexyxd1+cBEFkUxXpUysmSj5
7AwfRPCf/Icp8ywYap9N2j4Y9jA+Ud3p4kc1mZsG02xo28gt+wTVkJ0CU3eowTpw+1PDxccCjKXJ
YungM6w077VqMHp9cQZb4+xhNgpN/S31+nrNQV476XUVc9venTMRnh/KyDJh83pT4oVBzHoa5vt/
FZIIJtbgTPy/gzW5jGNVUbbOl+p8FChLiW2A1GxJhhjQEBPbNvb1ugTG0bUbncy2Xeq6/eLrE7u4
8MWdvqGCsd/BvRCStYaizoICZyWlrzhYrBkBLlC/GRywRB4z5Zd1Xv+AB74ZisOfSboWyDjC6eUk
xFKANUYsS8i5gIGapirxGllPE65yaJYqZyaexWs/FAPFFyiLLSfK4UvDK1vYWqe2YoTQaHlENIPc
MPz8Uxk1c72JklW+ZmiHh+npHdFFImhqBoawFX0qUOvzvoLvw9WzGKQf+EdOXvbzJ+oSMQWeqsJS
OE+E1ruHjJPmV09eauZmagYT/ObAKftzyjDEkvQu2/9o8ZXf94etTq3jWzeUbVkQz9U+SfMbMXg1
CRsstAK85oGa/BhsJfIbZP96gb+kKAv1cE1/6Nz/ME85zy0qMNI3kCkK5I70EHHwfsz4ON2GsHxf
j3vQs3RMt07+/mL1kdq54uiDV5nMnvKjMW2xhZLzvek2Kvsk1wCU16JzdxPG5oCQtG7AZLb/QIVl
tU3T3Z3k/BTQagabbPD4oDUvx5BtvFTD1SqVTjwZqUOClYC6hQcCSlLA8JilF7AtNr3WusruH2QA
KoM205DWjVAFSfLDs5e1eYstYqDZRyHo+rg1KtyLBvbAeeVs0MFDjd+dI6g0tS6mfb/zzLCXsK+e
QHVejgzcN9Mp6S70zz5U9W4fdk1sjh/j65qqjkq4+G7wvF+GZgDiOouJV+OJJwmWd/wLQchSZOSg
+T5wl38GXnsqhm+ZFz1iTuF+hsAL/xfVs8yOiu9EJTn/ih75MDBCAT7twlC7BYWRGYqph1ccVQCc
zQsBTa7ql1RtGeriMB4+2dUYSNv5sTb5onQRxazY8uTO9/4UlLR02GSY3tI8YxYXNLvjm2H+8U2C
r4ZdAonBj22AKVJiHdRutcdBV07kK6j+wCSbEgTfgJc1VRQ75e6eBCtU0Van94ikhbZg79YJ8Vzi
DlBTX6mg9NoRmgeQUozaOroVP0rRknH+t37bUp9rsYr6VIgZnENeSC9EWkwDdmJuuWO+iO8ACc3+
VvncsvSoVJZDN3M/rTjAXnCtHlHs8ZYrRB/l3GuOumJmcGKaaNtQ7sdLWZTI74MLmRA3lREwgIyS
qiA88hxqvSCrk2en3WKrKUPbnFdSdnhteZ8/NmO9QRlksy6gDJqZ9ERfqBVvLN6G/HGHVxz65EiE
9xbSMiaFYDAXIw7TISiqcr8YHnPJqBfHee6vXK1Fb6nZ0MoRC3srLGXRY+7etG3cXqtxDYcjAA9c
5LGSN5+ob4cjHaM0BzZDFWV1POHZwHqwWfgtxU2V5OsXhYHOIateRB3vOGuVYPNqcNxNEoaoP0vq
ktJ9UIh5KnVoJkKtoZhWvQwRdoDeX0Hq+JsRRbgZ1oGJQ+63kGtgeio9ZNduh4Vu+3JPLNYTv3Ce
/HXqZUR4aquj3AtxMVuzyJhupF0LIAXo1LjZvG8IvAAPFh0nSnWRulHj7gDsJkXbf45Fcc0saU3t
d4TMnAz67h3B5vsAZS/TvOr0egs76m3odoYWv+3UruAkLsNYIMQByOTBY2CJquLw1RtnWajswZEi
RKmPbrGnHilf8EHt56SFT3p15h9B2+iTKKs+qJA9HWcmJ7ypJUKFLBCCIztmJpwIoRoetLP+3KXi
VEU4CBldLO+pk1epoXpEJZdeT7zhhpfDoo983ByPtQM3CtwG9BaHv1ikmU1A27riQonToS3Hrk+6
wagmbZrNyoY9TzdeR4Cf+KFPq4p69i3vDCGPtKXLGy+/yn8qTEloUYDxim99FiudZCAEZGXTGLSw
DKL5qdDDVng+aYOjdT7ONPrVdXXZv74sTpGXEZXFSAbV9y661lYH4P1Z0VRfsXCK3kBwhYV8eZdn
Xes8DNf7GLOYdV7ksvT0iA7sESeBnO3EJdaIoxMozPygEGrUQcLOkXzWgSr12r0xDFUY/g4l/zch
bRuMNfu3VMPTBSi5klMBZO6uiSZiydOB1zRb6r/m3eOMla9mjsEXgWdQSrGt99pALo9Zwi1Rbmrw
9ol3JSVwgwVrLARm9ykBXO+o0BiLmPgbatDf967ZhX8gCa3Yt3+n62eQU1Zn/Kp8H6+qivoQMhJo
OCDwckopFe9Zmsgk4zmLcf6xM8sdUV/ixsLVy2WIc0LANMZfXbHqMDCIb8FlEO/w7qPYzpMzNhkz
vWRbW2C82PyLtury5nchmSM1+vmAWcHaDxyz58KYvZB/EKDQnIyrR2Mh8qwRpKheQl0Wl3e2HBUT
Ke5A3qhB0xHzTlRM/KghGrmGq0Yz6AvcT0SBQc99Ol/23P7Hw7Kx45ny5MGUcONzccz8evP7WVX4
iRD1S4Oits1QHESKRehhkSPC5m7WlAAmegIKz75JMs8qzcg6YJ/t9qFCz0NiOmdWiB9YfTEZ0Gnw
kp6FZvBMqBeDIrq07yciICEHdoAhpPypi5owxgvFcZNLFEFTSwVbZGuJPU5c359aoCb6uHxo6k1T
17AvCPsQBJA5PP/2VYmGmC+CioIjhYv4Pp7PzXOaoObgF+dpYC0QUTkx+fWlG/J2MMOfv40UACAk
Vmh1mtiwHXDraXE98/QcIj4vV6NCb/xgS/YL2BGYLjwKTQf71msJwqECRS6eaZfmhMnHYmBE4Mrg
+WB6wuD6Om8IKR8jeUTa6UsIlspB2psklaYgHyYEoAPQD2RTVDGW5EhpSY2phiT6UgJgCGpjXuTZ
sVTqjbGwy7leTxEg1IHA51Lz4snoCBAO7eUCwDUXZfqZK2MzqVPuU3F+FGQdE6Oog8I2xdDxBPts
DkVxHU77Tb4u3d+Qa4FMEJxlOg/AE0gX4vuxAja7AS6sbvJwKLCHJ8H6XlF/V6FvBLiwl330wX0t
6pu82yaOQY8eyJhVRwHa1D4rHaRTf1Lht4RymKpUa3PZFFgdQBn2fNUfcrljmeA8VWDT2y9vZ6zz
JcjSTBJ2PSwRgvyBwWfoGEy7/GdFBZ5ONi5/HgQdSY/sIf8pASFFz8Aey74wzWH8hZ5ThlUORp36
tU3ALsA2G1XQiCW+q2ur9XVHuU1IidVkaNhmJfEAAXITkwQM0xQQnj+mlrfGCOmvhIA+PnE1lPwj
NUMv6doCFiDT/oign9FkOCT4XhBP5p0/jG6VE6bEXpsCZra+cYZb7mmf8UphKS3HL+eeuXR401io
Bk5yjPpzy9EA87dn08ojllPeKFlZye+SSxA17DOGYpETY+sLpr03SBIcnqtU9WFhE8PbLsvjAMj3
9l5FzLfebUmYiwAy/f9tGcC0CJDeOUbOi+WwqJ1ExOURqqkGu7A8b5SlM9oAUXga9I9VxOMJb6s5
Va7J3zTdllr0j+K3YsPpal5LrrvmqFB/Lli6HPym3B7e3/N+KZ7AyOyBESqElr2rRl4Kxch54eYM
umshuh3XYwBY/MfJOHs+YMK7s0cXaKDJhIOIoOSgCCqwWaxfirWYD5qX5OQ1G8K5rtMAiogrEyn/
oj+veslS96Ace4tc9PYAQfp6aMPoyE1vloSI47ub+32vcBQy2OzAmz44qJdT3+GYM2a4NLbd5ZWI
mNT1UMfKFF+qfzEon/scKidNb4IP+/qTax96duJT8zt4JCm8e7NmXoE6HBI2CmXpPBtUO3He3fBF
j3XtqpYL9iQj3iDV1/smR/enm+z/k+mpOATJbKNybNVK5IK0WiRTAKQTqg5mvG7i5DOZ8XYNWMoP
c0xWaWgE9xBIiBPpciAlvRhpSKK7dubex8kiXFaKtxBExD0Eqj9aGGdIpiQMJceEJ1O7/twgrpSu
7GZhyvTU2yQvnXZoNvWIwH62j0KHux5541SHYnwOzAx2Y59GEJJu+s887haUgI/ojzwrD+QstMdT
9WT8QcFQiSoZNwEVNKRcAXgSI+okbygd1fg9NqPQAX8XoWGJTn8LqHfyNXkOG4o4v6kD3x5q69P/
1pvFJVyrLH/EIWXHoQdl4wN99jJZHJ/UMQvqG5FKLH66vka3WSkceJ6okKl/0JFMM7u4IXx/D1+V
wZWNB1us1crl+JOh0UjFda3HZEIM2sjLSCUT3xnfjpZueyvp+R+M0Rea1qnjRhdKLlo3k4l4S271
3hyNPM4jyfKFf7QlWYWI2cwTehaZakOV88K/UqTv1j9DM4TWZQb9PYfHHXtSvis997YunYH7Dnzk
E+BTfv3O8nRrUFCbqr8db0RZ32trGaRvt+2ipZno5wfOOKfwZFhSvDMI5PgtOybu031Ai7BHAm7g
atkrx7Mpb7xhWPls4PX+tiJSzICa8bTfqvIag8txyp/bpFm0HoUoQuc9Hip6DbBAfu5H8cgaxn43
NJG1nnR8Auckk/9OUkcafOdkfLZMeU/pIfwznAedh5hk27/fPPkGOKoIf2qZ5FUfaJZhDb0MkCm8
bozXlsC1qgv1kHSKpa8zPucobgmbQNP5Ic7Mx9RScKKT7NpTO83RK5mrqf4nMY/kou58ZB8L2gn+
WyLRikCoAdB/1nlhbX5w85kPnGfbjjXqaKkFGW1yLjTAZqznkSW3BvLPeVHzlk5a+rRdWhLa2tgs
+GyGKfPe+a7zTA2TDZLSZg9jR2SS2cUajAXf9aLT+7f1f4bv/GRiWzQe6la6sM5LIuAVZdOOgNVn
90cVqrC549psOS5FUb6U9gPlzZRW3TzW4NrWgprwTlQgPV5Jr1BxvcPUoIGig8hY6L2qutiAGTCb
4kYh15IZ+ggpXbGDxHU8rv9SxNAEBIvXUGSjplxVkKq81UR264FvBUamHENjh9j/H8x4Htiq5HpW
dA9H1989VrRdxZIl7wzOtw7Y2yGF0Gp7cQ7jyqdeyRudBR5stZEdaE5x3MLJsq6+glugWaHg39bz
+ANr0uzWjUUUDWgLw+g+deE/UHmrYrnrWyuQbJtkmv1d2Fxy7kLQqdnQoKNHdZooRGEkNGSQUPEB
HVjzpcqWF5x1c/WMiYhHWVNZQ0EKLpi0qL748e6NBfEFQQt1mUlY7SlI/pAgDdSsynSjGQPU7y67
I8tZvPX6h5lZ+9yJsxNPItzkYhhT8jDRLpiLlSr2gRYibJKIU4XoMPf7gCZlg2AI15P+4yWFUmA9
fkm7zEF2n46Of+xwL++ZjVzHtr2CbwsXEuM/k6wmDm5L660i5w+sRDCB5fEssOAkHa28SWsz+fas
li+9XrvDdfn+i++BydXwkYTHFKef+8GjL6NvjVPEuI80lYX9jCexEiFNFMA1NHBcA7t/tmGRUJly
/fq/kXa2y5xs6giL4NvjRkbo8O0XbLPsMqMXJX2AYMWwxBh1LbPEdiNjWJ/R8CZt7e/ODik82omx
Iew3uRskvyOVmiq4uDpdGuDc7YLEMhd2Hpi5JnzhItu8rb2k/+XCHwChLYgjO6Ee8KdztTCvXZSE
j0KlQ96iYsAVH2Vp6gp9e6CVdHCeObkxOzq1Om1zteuSpY/Z+EWdHrfd8mVhdBoeTgXibY8Twfrw
B0l/74Suu4N0H960DKQc48ZVpkronDUzsbFJtJa/rB5Yeafro2zEEeQUvARwtimQclN/GrwXnZ7P
49NbZe2E3KWhmLM0uVQtyE+POWMS78C9hQ7QkI0kxXnAunGpfK0I5lVvhOuqBmoIaqZtKXGroeZP
GhIWW5kX2uEiu6wLb9sHN0wiRhrBuaWMUMsRwDbbGx90fP1eT+rcZp2CVrQSrXEP5NY/epXwruxf
iJn7LCai0krASQNY9bUAHsvwfStRD7fZvTShMbC9oyvbiZt+TLsZww+k5l9/nkj9m0FsP9mDvX71
BHtgEK5Kfdxx/9+BjtP3coWHoEMAjQx0+u1xN0WWCaPJ4ehNzZ108LcQNawqPZl5JcGEXjMubT8C
phDYo1IKvwzQOGvWPK69ZC+WF88DUxxvuaHEqNwZ97VsRKBIiXGm8MlvY8LkAUGssYSTFZkvOfUG
wpOsV6q+7WT+AJf8jSgDaIXr6U7EM7KZQhvrafxnsUBv9B46ASaEcwVHeo4C4OdwUsJmCBLfYuLM
Xby2Q5aZoBBRc5pGjrSw6C3zUAxcIn6K5EznhtmXa/HGHXEcl8IRraA/oeuMnSy/37GFwD/C5WNr
3NDr1FF5hVifthlwWB1+TO/Fip9dbZlqpGfr78ZgCPhg9kWMSvBwR6HQqmZRX4dizi+b/uSZKeOz
RlKAj6vye7HjnxjG0MHCEC0kPeARTEU/bDY8VrfFfOSwQjR/+qnYQUdisVcqrYnM4a+zYUa9C08v
6yHJ2uSzQL0knZkHbCKMW/7lBfQY92nIaqIKF8HQJAOf/A2W3O+KjY2nqXUW8RsatpI4viGYlTEs
R1fjkrffN45b/UrhuVCEp/tKU2FjxLOaMvwC3laoq8GZWt5ofvZ7R+IOAP3T/cOT+2dkumamq2vE
1ot6gsGkB6+jShqwJwU0dY/C2/eq5bR0D9s/WK+3BolBEu178UbatjhFJedKp3imRTsGx6S6EgKf
FizuDsMunsn7yw61QAxA0koY9kgqYvFxulbMv3MyWCi3UAtJ8+W+bq6EpQ6rJC8m3yKPCc3T5hlu
3vEwYf15nwf4lkrGQxEYwbMNs59xdL4vt9nr8LU1NWKlCXhr0bwDeynxVh3JGch8qsXLRt0AMNYj
CufsLOOMxFMVWztgRDc3hUjHazQeHiNQ6dZVrlr+8SV1Flbli2qmJ/NzrVq3834J3dbenPu/Ftzn
7KHInMMK6aNLFxQ6LDEeKu6GpAz2Qj/O3oFaxbPLsbOz2v+kbl/PELXfjg5eP4lGsj4WCGINYtxj
JcQv8ZOCYVS8ywavFD1UJhsS7iyCjMiMVtKHGySYy73EYAlf3bwua94BFEw8JJmMEM4cVX9YHwaH
CEbcoOnpu3sNB6ezJbvSduA6g19ZNgx7wBp6cF0p7dJxLECr9/HSholgTCdHo3q7JyJU3J7NHkpj
VHm4yVSxebK5Vw8GssQMT0BJpRnbVjKpjrVAMPaMGCp9jiwS6relSEweZ6fyAK5T1dKd1L0XysuI
hLFJSuUpkPKzvNEDn6IWZxpB/mGJBTOBds9LkATZt6i65sw7vSBaKLMBHuGTNilA7Q+AnR8Q5Mw9
jjReQq+jVvJcYuzIzRH9WbVDYWECCXYiKa5PiZ8L6/t+/q7AkjP/JLwBXriblLw6DLQm6RP1eOKJ
+qPZIq1p3KIQq5ydqWwe3uj7O+/S6aPlB1ZiQy7cOUKHZ2XUTqeAfGwrN2s/sY5gUp9BDLgIpEno
syvDALu8Q4YmjxaPpJAN5uyGupSpMAOgsYiuPH4XAISW52hjnqm++pWH+C8hl4jPCrphVfCbKPWx
MeovT6lwfQowIWPa3xkVCBVaGF1fJzzkOQNOTTFywfyv5+IkFSJBUxT7kPAfHtLS7Fnd/rBOo3v4
A/SWf89kjlkO+K1RR/9e/2YEluiowob7kCEfDGWOWU2LQJ/1vi7OpcO75bIKHnug7XfpGBx8zouV
D89fOpr7FhBKOwW17bicvhnVrcBDPP3AxVYh3EdWKKQj0PQpOKILxvqMukstv+qAKUL6wsq/MC/J
pUBmV0K8yV8mBG50riWeYR+khBDtPaoPW2dGa6Qplpmh4k+6IQBy95ZWlDlWR2VW2JeKlJ4Ta0/4
d+Z+RldTkcuOEORaToQYlFIIGouHp63C/kXYbTJn1KOwCIkEZc24uz/V3EUZHuUNd7No1gomM3LQ
JDeTV4asOZnC950hu/2JnX4UpuMtzS9J+Qw4iIFxbwYCgvV9Wq+uEWipvXvJ4MzKYxJWOmqLXQpd
Ua1tzCuLOvL74q69KvAvnjW8yT2t0EI7qRE+lPJlHKueiE46BB6Hy84LBD9hqYpbCZtoDtYDfFLg
zp1fKRRiZtrF8bikbpQBX5qBSNabh/vk5tDLIcdlcscQ788qcY/+dZG3g3Spc5WJiMGmpKeQxs2v
CIydSGWa4j/bD5JejgZBxqXV6+VeAxT27/B5u0TQM8HuBxvMzA8c19rMrU3YXrL9/Q+Xbz5QlZr5
PhjC/q+BEQC2bjBqP5jU1Vr2YvD7gyhll00llBmyJg80/YPAVEqI8s1cDmU5rzd2Nqk7C8kXluom
GXZ5ljq3jskv1oLwI7cFlZ9q017OzMj7ADiQUUkgkBEHQ1MhcpVMI8Ug10mU13iIHqLS1r7JVdft
cbqt2x2Srhv9x9GrmRr1VrH5cYvX/FXSDF0l3qgwCB8H4NFLGDLB+9pseJ/BHbhAoiGNx+ZN29Uy
0oyvSOSxLYvuP6q7EE5pdXN5yynDFofmIyPQ2e3OJsQE/hQPauAvyG/wOVTwF5gPljJBQLPZxnzR
zoJ/gVY8Xm6IC1Qvuxv/A/b13duIAcK3HmsUE5YqIZxa7DAiZSuSz1jd7c7jewF/dcl6Q89nquXl
5lBRnxwqT8WWhmwDIpAXCG9N++OZldf7uP/sqjNhPr2FcuyfNI1PHACHrNXZV/m3NI/OBenTH4wR
mNXfinmpT2aN98cJ9UVjeCxbb8tsfyMzunhG5NMzf4CixX+xR77IW9sSMo0zj6ryPYIWi3dusAQ2
Vvo6C2joZjbhLnDfuU8xASPvSnGa/yneNO/L5uXYcS8SZW0j8qGXUS5JSMkA2CZcbW0tTzD01CGd
Rn2X4lR2XIFlvX9xJRAGnSTbiMbWqOh4ICmq/1EUWXKWuiJneMwwh/PKOzlJQjnDo36PFmiNDwyX
ZLdCLD+rqqNP9a0e8zj7N/FsgGEV3NZjzqlIiPEVA88tIUUFjDrI29y2gOmIxao37D/a4ILhQewa
46S1MMh5k3DzDHgPvJHvAWcAzYqgSjLPcJdPUNv8K7Y7P7Uz/XqOPHq80Eb+G4mvtR6g7BUtiQnM
W1Q+ySO9dHTfNkxfP82+b0FVnBegB889C79kn+3Wt0QUnNHxlihvN42m4DWybjx5K4rju1AVyVIV
esi9yER+QOxl8J1vT8GYPu73qV+haw9TuAC2L58aWI4QaMsFNf0qGjfWwdviFkgvZGLmWRzVNZxB
ys0kXa82sBVurPgdXqlkeXkicY1UwgQuJE6guvuPFu0+p2RtoMCgDYCNpRithsKhwoX57ROl3ANH
i2Cld63qalFyXoPUAvzyPVOpM55erRps/WxEgoJzt5ZAaz8xYMhgX2D4gSa2/WYHYEmld4mG7pq1
i0gVSnqbUiI1jmx8lN2vdUB4BylCmaqSdAj9fR9eb3M5SyH8LTbRavUA1A9olLI+Kt/gwCMFlUIr
C6N+BYcXbOANIW6GbW8rqx2p1QANM3FzEXvX4ehB7a0VolXvxryz5qH5x99sKW2fcDDt2Y0vibOd
52t9socJZfo+uWWbNTICVSni9ctB4wQPQvEyXM2i6IdeVzLVIpQgZ1TAnF1AFeLs5McANMJ7cxYi
mqdldzPrrIPjkFuX8l/XMOHCmtoIHlv9Ju6C/KJ/+RHPeUOOkpiqkMq0qg28NOiPXAxvhqig5uWU
GnzBMqGo6O3yF7+4HhtVxcN/1DNCFxkm+xv2FTQidnASD2NM5zl/3pPxJu9Mn2+H+g+0SeCHGC7a
dttW30yuuCVYe3Ml0i6JNI6+4kv8XhouairSUznjy/01l2qpw8guO7OcAsmROeQRzgdpm7NzRg+W
6GN6ffRYtKiL80ijyFu+9efdatq09zMHjQeKlJSzjFF9iL8jeS2jcuoHTRU6Ux5oJHZuu3hmO7tJ
mgaAHddgL8FTCn6JK+lLxCGbnLFN3XPrtQ1t5xDmZKVzLC+H2MGq02C9MGSC+Oh7olkuGSA90raK
G2Ap5/4KjWxQ07KWLBhXlSl/x9zgrC0nLuEKb2Rrq1zyQFmyVqpxRza6WOTUmhoxQUhJEXmoeQN9
e15VuvGWwUXMasyDGettG8bR1yRq32CjtPFjuMulBRqdFL6S7FwTvO/XblqB9rEEP4pY/kocDyfV
YP+hqs8oNrxl/nUYiASha1dgGGDmM0tzY2Loa4mEuxTngsutV7K7ccoPQxbTcvhtfXpyPACqvTlU
DVDh6ZKZJlVTHLHzlZ3Rsi+jXy/vfPKqKVdN4dXyiJS2XFCrpcSNR8nTOmfo9WYdeuz9XWyxtfFj
VBxtp4lvS48+nUQxAQBq/eqPBopYb6NBF8zTkevNHQVlrUntfqLZhf1fT3GphPyOP3FjIMCgwyNM
uPGPHYRm/99SQ1b2zXb1ek28MndXUftAnGuxd6jqxkE6vlTqH4/qm/D9VN7RRIeutm8o8ENEUhXV
nqjFChHJ/FCNnUnyLkdvTQHbh+ZySvzewS4yiLV/uwhqg454CJ9Kt3fLs/LclfFuylLNRxXK4Ave
T34imWGlud5ToYEg9myufO4eALkXxB+W0SNMbSd9QAevg0JYeGrI8wWxaLJi0oGlmWwXNRErVWgL
+L0Do3HoWdOKcMZ50r29/Ru6twlQUV5chQ1XicCBtKZ9wdhg6GAfk0w1550PJOQLFa4JL/IM+Z91
kysCSfNJMZ698EaNRAH/OVuWUepG4xMQ8kG6WtonaR6zYOYtiP8u3dUww50x2XYO4xUuMlnAgVpV
gEL1A6ML6tvShT8fy1VeSQFxWdF0/owVJufLCw6EffHW7A+64jr2ZghSAHCZe4DxYxbQBng84fMW
nkVNEtN+enBW5PAzyVsAVfGVo/qAcdRhWkUt6NBB1abuWKQso+vPUokpwzJNO6EDaA3J9vzLv9yZ
XE5v+xHCUTFtdx5QIaRFav7cAvzaNKXKkAveW1J5tBZiOCaSTTp59dXcJaDsxuFo6NjZy0/jrPYc
6duTZLNMr4XaR41dNbGvyDsqxlHsuzc+Ds8ZqeOLHziCN/BN8CqsChRveEMjR0lwWZPd7yyd5CYL
dVwweldQJk0Jt+1W5tJXv/ye3sb1ANc0EAuwxT60c3D1iuvN4m+DRIN3DAajUkkdcwun7PMLEZGw
QYjCSCFZoFLLJU3LKJ6E+v92LjuMAiJaq2OhrdmMVyJPPczXaTfFuoBDNVcexJsmhAbiZN2rB1dn
vaqyOE42haFFvCCeAoVbOFK+YEVO8qN1ukvXyovQ30FWW9F0EwXbWooYb2EUVRfZY3CBJziEu9LX
cesQBNrr+gru6UE66z6F2dGZ0TkhxtKtzHsjz1XsU5vTQrzbNsUivLZHQu0HwW/EGGT7rU5bHAzj
30c3kClEW4e1EJVYbbodWoYFl+0zwt89ugoVhLgzQEYSwgzgzljaGD61Jcc/3PmPNjcym135wVCB
Z58eoS1Bchp3gNVT3iExu43QyXs+6FB0n7G7SSEDJrFLWbYiRHCazppLSXKqruY1ccsliyU6DbdX
RhxnKmj3aIuF8a2l4vi82LN8NApf/vXazd2VpKBEQyDcU5QEwqmjoZeKrg0FvMQWqcDGk37dNSbX
BmFSVqZvX5jS0zahyCHocsy7EQHHkgtjfk8Xm5bYMFk/fRgbJ23nFX3yTo+srFcrEY536GQuaog0
nBtyiRf/xmwTLdewq1VYhHRbirVWQf3OWZCBdBCBbp7DDcHs/6vd50Nh8HvQtvvhSfZebK8KO1Tp
StbYcpHeOdR01eC9DWlJR1ifchPD1MWgQbhAM4L3Dx9qYJA7Srr3GIAj2WZRaoEDHu66yiSlOVI4
Jf6vNqE+O9B3CGqjDN8mLMxqSqVshBoUaPA5OWl7rL/AfMgtPw+T+AqCI5ZuaMLOJGjLoEhXI6H9
s6+/aK2b3Lbrle2N1PVjIV9vLfNU/IOZVt3G4afgBTVh6p7W8JLJyZjf7blu9hw5yuj3YlfmzglV
xH/5Q++vsGxTmeZaR20O6l6cjzNo4IZf4sqSnAguaoheGKENb+4YAbZDvp1PEZZ6jpjwmkTHBLJS
X5aLqjuVBWoTmAplhQA4Vc0aiWZ/pQx2cmhnBdjzCROvh7RymsgMrnlnRL00fk1obQlR2RCRGoar
3tsRSSsJkVZDU+2DYLVseZjCtoB6VNGnzCfJohzib/LLFvDGb3+NK+6eqRLKKNC27ZR7L29FlwB/
yWf/hiS/Ql1Uv8edyTqE8r65xs2fwNwMuoVslkyRA8ETwGcv8SL/sjPoN09+xRIB/paKYl9NBjw7
tkD6kRlAA+m698SZ2G3i7xG3vcxKjzNuiosiblgk0iikxPa1DmvTnrgNOE2mTy52StdTnGzZ4g2A
6Rg9it/LlR/pvz4wdJ5UfM1+Vi45KnWkv1tDfwSqQeFbXkhr31al9iN2Kv/oEWg3df9F5yg/UG3y
H49YFwNpVnXpib6p6cMKRfbErQStCKo29WvxgF1lDQ52ZFvjyY2loCX4hR4HIHMVhaVm/SQanzjF
aL9K6bY6YYjz6ClHvNpW1W/WxIYOoEaRwI5VFVZ6Lk6+6xWCw/yVHWI5jCSDvQqecH3SQ+/VbFwp
+34LMuPr8kkSTeAzwbZVaWQKXgqtu5dklIxLG6in5WTdWPdiR35SViOhITOo/CjdZ9p7dItFzWiz
+e16bhbrf2wmIa6f6TGlSrBjAhfdSVtMgxU6Dlnmh9CPNxGxy1YQLsb10oSd/Gy4s/UqpZjjWPCP
Lk78BAGyvqertS5HHCrNPOXEcyoUaOs1V35s5OCjVTooLgUAoUq68YNWupjl7cxaqz+ZT6H+dnyh
7wU9ZXvrtXTKfFLiSzIcvUF80oA+pUY492agiCTYC8wJP6QiKjNrlVsdMZuSgKcgKepK4u4OkSmp
Kw6jc8p0Q9YZZxaNHxqReMm0sMT/ZTrrRYh3LnL6MCMmhMgcvoKUJ/K6OZSMITCYIFm3zHw6vgJs
PSzkgU/c8shcsOZ3xlqvjIcE96NpOVk8taOWb76N128NGAA5uZVZE+6EXcUQzDJBUXDLM0UjrzJE
mVL3szEaughDilxE2j+hLOKHEn9BiwiQeSMuFt+mtlIsc0cUn0g77tSuTUNEbbGYOLs1zTVKI5Lb
LEAeY4o/3CxF7ZaY4hiKj1RopoYBPQV1E0fjnP5agVjs4ia7oWoJ8FvwHq9e7hAGWO/bzpLdL9PH
zFbjMXzbs4YB7+4JfGVqfR/2qMMun1I9oKud/ElHqhBpHG5+QjpnoXMn9R3R36RSX9hW2J27nnk1
G8c6DxH6aSoP3yPaDDcNjwSQRaTj70XIL3RsyEWjWp/jHabas2aYcnURAdlOtCThdsAmjDZd14Rs
+WUWWbomuGgaNWyE+wYfS1bY8OWKaY1cc7yGiBKlMKF3r0edTY8Zd8+3JTzL6524OwNEJpFV/LRM
HdcSlx0Amu9FM1gHGpM8rhtyMH4QyIzXBOQBGqyWZrFhXWda7O46QtSDjiptdL/Gpnzc0RNOFkk3
RgIQ2fmdzAXCQpcCrPJmMdopDJ8UcxGbhruCenzFvot11Myyzr/PYcpd7OxNp45Td+Xzdi2rTR9x
WjBfzS2vUGg1AxF790Ssbs8CRI0UxOWedsNZASp3HLe3HAhk+fqeMr+fEewlJSHUgiWs7ljWKmfR
ztGFk8qiB9m+HEhhMv9V0Y4WwxRmSi5Osie7uGVj2RqfG+IyU/aROr5RMwISAGi6YTVsS3IwYLEx
gpFCS36xwgAbx0JiiX/V9TsblzEn3MheCuzLodRvNqejsy9Gym9jAj4ks6dCADvCjidJ1KvI2kBI
XIdurC14ibYvl1sWgt2eVscAv8ehTWAA0As3FcYhf9QhS7sWTV2LlO+nbDmOBBRu1lNWNlPs2a5y
4zhswgscmJvVveCPak6UEQjv7vVmJJmcz3yfc4ZNIDnigNCDXMjpfB9cfdOah3/og/nOlLE8LWje
3COf2zNU9Sr/r8hjKLzzH8eNT9rEQeFNt8LVar1GfyJ4Z2Pq3n8MhEC+2Yh/d6MlsyFfJ/cc2zdC
ZzkoWfqukteZXjGX4HJh9/avuB/gqMYgB7/ksecwL1sieRDdNunfU2U0t/+qn+wWGroqoeJknfdO
/mCkd64X6QvPJGERupuDrwhsheYwjwCyilzarb8TaEo7w/LaKvJnvv0LCeZTAzpNBn7Z0cqlziTY
lwqSaog81sTIDTVToxpEP2O2ynt9GfOvHGgOgQx9p+UP63PxOg91fVTktgpc/yXrpuh+ev0CgG7e
Ou33WdZqfzhX/z3JT94yMws1XUs4AzDhM7G2RinKGxEkhSHsD7nT8RSqAeSDkrLhhnynFMfxOQBx
xh4ero0eL1fy6+hlsmzQuz6IGY3AZosQOgigyC24iLUyCZ5IkPxg0G+GoUmSVY5pp65w91xCjV8v
rf4d7pxdStIiVArqxNkPh6ON0+i2Yb0YZCCyR2C9KVWugs/uYmDAs3HQMfr+kmJ8sWrqA2SxwnM3
ZSelWT0hV0ebOSgjXa65ga2t65oF/YCQ6YxfCqBjwt90SKkczcqgTEXL+y/PyUk/hftPI+M7iQo9
gzTCfD0RDzxsSBH5Z3upodmk1FcKbt3qQhYeCfNm7eoDA/HI2g4BeFZk2XJQA5jU5piA6D0cZBBm
73NztJd97uipXEhfzwe5tFU2yUMVIp9SfHErF62GqONFDpzTYoCjVEkXmbdInL/8JVqjwTp38Qac
D5zGdw4YvNRhudL25AleMXoqVhcLC3aO45U1IUD+Od1vcsThAJPdz4kcmCAhnalYdYK0nEESdzmB
kgcbk/talTYvPl6yIWeKhPAC2OZGv+f98pxwyhe05I0QoNx3jWTwnJ6op/1rLHV1T5P3prlHl7VD
eeovewtKJLXut17ukFPnPappEE1EtwUKRLsIUbI444vQ9kwumkNC9oGvcX2IOddQ8zzaSui/JoAX
DeuerSXdO99CdIbp7TKSwmcCGXBiznEbGNCR/xKoAY1li4mNj1jhnYTfz9fMBZyEo3vFAxmVXBQL
mVSwQPu/723J0gIp7YBHYbNatoxhP5EVGrqLU/p5ZHB9YEnuq7s1YGEq5gvJgDdwGJA02f5saw/9
3tyd9i30TQIzPNNriWd/1ai5mDuhfI/N8FCxJ5f2u8Hqa7t3SZ+O1CAJyi23Zra85vcIF29fCCuH
h7qdDXBZpRo1CC5fkVALWnhU6mKsGh3gjV7zTINc7/O8G/G1EXg+GaFD8VSrFhWFUzxp90AJMdy4
elKpAp00xTJolkGXceZvwKTq3SG4cIb698xw8ExrmJyK+w24ynT/2QJ9Z6F6qZ/54qDt6nrX2MRb
X0EOwgKAv0uME9EdxmwHirTvbJjAjgJEdK3E9fDNjKGoXdG8Tlit9Pkh2UB9JbcVU+HB8ux57nSN
pClLYUShpMpKZijR1M7ndeGofmHHv5hysZvG+7QEBcc3cYGYbBJsTKrkj1V3jHVsxmuCYlonLdaR
q1Xhd+wF/01A9zLY6WXpnYrkvmar5x3255nk+pFyQfsuYwm9PVneh5mu2aS0DF7KW2SOjYJgyCBl
Ej8dIR0MNQrtLGrEbfkuS5DervimbgFD75HZwdXb8TNVXlmoQYziNZPJcB5dHLAIg9OQF465ulyh
Mgs1A5OJf+PRrrcjCNZHSpgQkjzB3nIIUQPBtZt6nDyw8z8ZDoUoFCQYDsCK+JAv4eoMqBUBwYwE
lOKXH7re3i/WArie5LKUiGP5R3Mmjq/qOSFKxzmWu8hXRnQF8+xMT0w8bKV38e6f2Vq/1S67jSZw
dpW3mL315FfzieCUiR0nnf7oLiXDS8b85xpdiX/jHHLsMpP8PZvxArvGvmABIQD9u0de/5cab+61
f1TDP3+Haf/pY9/Ub9RWRkl/Kk/tIG/GBVUSFyJbC8a3mdC4qGRoaZehu+3IHjsNssmyEe/T7Bkm
U2L7+zaLL5irO+/tRMAwDkX+CbnPqW7jHuHfoCyFBZQDSRiR6AUPvUVrbi+UsT79PziBXiz9SXAU
0fuh7Q7m1ptU3By5rKLd22ZEYc994VsVVRgwNhXxTtDwIuqDFiW6cd4wPXxPGbR/5Z2PiaXxSkaA
aklhRaT9g/upJ8vkA4e8mOSuAJF/Zo6pJ061oDJoLvH7rDZ0dMydebGyfGZY3UI1HaPf6cPgK4HT
dzujji2wOF8hfNHcKMw2BpANp7afQZMCvB4ZYEngGZS1USEtxRWjxaLhdbW724NhNndl2heBZvv4
WAO2z9alS3LIlru1b/GaKnMG13dNusLSJv1Mjasho5gqrRPnZ8nLERJJNNRaJAgbket/I2GO2ynp
8ZktoIwJB3qYV7p8pXqi2azvCRjZgAduJcFL/VkNIUR2f3e8PoUmAchrmoh5qBORImqrI4RA+UM4
22FKKcv/oq3WcEdXFwIFaV8+uH1i0vn6asDdUJin5riqkuqKH9R+NaSlzYNVkNot2uQs+KhOA4hI
O7+Q0OuJk6Wk2jpTGZ79SYcppK1sgWN2Z5uSIWFzIQrR2X02eqykXwEb/eyOeKZ7a59zUwabpKWI
22bOexyC4gMn1CRLKOgo6DW58oyLRhMNpSonKRmkBvXNFYSZTARpIzxoYRbm2SaXlY50Iaf0TdV9
jBIcUK6PyEKs6rR5BpMZxRYZsWvB2z802AwgFCIF7mECbNK+dxIu1ga58YdBpOmIzpXHyh++U+Id
lhuW9IMLMi4EfDKyUHU5k3ZM9IMTHQAfpeo/6066o73vyl+4CsWeXdZgTFRI8aPOO7JBt7B09mPj
ExqCwNX6tgpy0L8ZV4uRHMx4NDsWC9F5oefffioy5p7ZvZQD3T/+9KgNyTV59kHf3nl1duhSZjdi
9utjR7lPNlye+bUyugtwnpxqman2YrJVIdjfq6Nm9J+y52eKJN/dOTUUEbqq4sk2qcxfrvmEieAu
VdX8vPosrnJ61t0rFTgdZfypK0W8gIAICFPJpAeeZDEs/S+iwpUJb1guE9Sobc72XIZYd5uuRPNX
QrC+CJn/b0gU63h9ZgxtMpUZu+Zu0R6eyeFekvCD84B9XHMjQLpAzLMgPogc9bjUVSTvSUSFzbby
hQtZozQHKNVV88FuhPC2S0yk0+WM2VeTqcwFe0M7K5RrC6bWNpwcrCxCera+7F54O98U5XL0eUNB
27cpWEB6Hhh/Rj0QFvbKcXasdOlXtJyFVVF6+RRBgqSdp4ioVSqhNJ1l3GMcZLGD3p3AnP6iw3DK
Wex3dD8UifCtdyVP9sYjgjuU8j6yeswh7iHJd7/NpSDzU+C16hqWIU/gvASR5kjd0NsRSzelSTAi
CMwe6UbChkCCw/V6uMnTaejs3Wa6wmgFvmH+vi4bAR03V+BKourQjm3SxIgTtKuFxr29kjIi82iQ
uhIHD3XvewmC9lCPoEEDed8pRKS5Ega1+y8cKEL25KW3Rny9vatG3hS3CQ8zK6znvh4+0OEqlYKa
WY2Q+aNqg0a9DoFgigCK+VHKHnQVbE3QeUlVtjk/QpP3DYw6D1/EpF+mGDg6/3nWNlZWGnBd73P+
BFtYx+kBLSaqPaI5VmejVgZgn2f7kdqWeBmjcACWUwoVVvlaSZjqtCKS9WN6eQkk0yKsBoQASUxQ
i6N7csY0iiM37WOft1aRZ9wPKFIs/KDM3ztxWZKjUgai1kjryQNTsqFwOWBq7OyblfNJVszdCflW
aTtQEwXWg9mCE2mrzCWUjjW2flRGHggWigjgJ9dw1b1endO7ZcetOE3rrAcc/ZwxEPEU0KpckrBL
He6f48+xMSzfVUlMOjM0ZZrfRAQZ7hs7XTQbzUwA3ufJZzljmVy9H8SkWZp3U2G6wBizbKF2ncUP
LDIEZezFmIJAdb/jRqzRp0aA0Sro15w+t1jYVQ5kfBSyL6dTGDuv7F/IHdExjs38WnR8C3KGshS6
txsLCJkQVKj4Gg+K9Ha5OHWyG+W63NBau5FdXN+EzNkhssiLG/RHzTODy9gojaM+TBJqmsuLt7ty
srwxyckn4AR5FDAAXViCGyODHiutrQ1CiG5m8lKzrsxJgyDQwSJsuEdOZaUirnAVvdLtBKHyjZmR
DVDAgNrrpPDtxZJgs1sf8K2gXyI3lwb85kx9FenAdQy4Tv9ETSfK6pby5sI9ORCvtkF1/4FafucT
wrQVm7+43hvyFw/9RmBs9sXCasvWXatO7YyNfmoGocdet2jptWfdwGFIomvTysP1U49hFZMkE5FB
/Y15b+0ScoQD2Kd6zK74bBad7DjHU/RHeiFoqc6LztWB8a3+krfLxj8pIQ3K8Zky9035y9PJYn1u
cH7NNQwNVyKdOe0/3xL8p++XuDXj1AXCu4ut8AxTw95iozlYrRS1Yqwhu6ZWJdiVHj0bTDnI1QaN
7MlvzJO2pjgjKrkCYHxQspc/yQ2op+3KkP53L4tWdOklpEi7eAyY9Jnieu9dmaxkG+l3NzRAhjpQ
QEBSX/7/hISz9LnY2S48Doclm4XXGevGq4lG2lHwm7f3/y3yx0Z9IuhDzfz+6K817L812Rk/5nfQ
8dilXFwu1K70Hu70C8GJzB4v5ALA3LyhxPL2x+/FWOr5w/xWJBmoC6v/jlIr8esy1FSMnSRc4oPO
5pTBS1lS+n9gBuIYDlwfI0KvcUiIGLAjO6jc5tPeEOnkdmH9FH3tkD0F6SKWAC/kjr6EVhTAgpIC
qMnxA8bAGxqM/REt1HWAQvAdjk/y2GhTzV3+RC5ud9mcABgsbM/QLbz3veXpGWvDYf2gAJwce9+l
DakTfySh7WRBRuiBsP3hJYQamudY0tgkjqklQCZnozNCMBjzP75uK5h6A8BgVu7WiL+JL4FEU7yM
U2ZcJ5u1LR5Yx9AYpOjan91o3nv1DXAINq6pUSgDYm6hsO7C36UzHlRAflYLnRFK6bCcP+jsXe/2
y1EaB+HbMc9VNr5EyVrLaQxsEDTqfIfnbHiiiJcFFJTVhZgHJMI5BqZYlxuSsMFI7JpLrLon3p4e
v8rWHki+TwPp5eP7g5KTVQHEmUNjvYgTUoaY4EOgkm5pJOyLQ9Fpnppsltgrc7DnmvB91imEtkaV
TjhYbDNSfhSFFGql/TEHVh2y3n+izC+MtuDgpXqNZCJuz0X2hyqjKQxjeYxiU0hM92KfRMR2yrUC
oV7DxrZTYN7t1W+L23P0eJUph3qttf6cLsg83ROwgOqeMgKvLyMEHXlMOz4oNtGvvy0DM/1wK+6B
S5/Uy8/M6oQ0KzfrPgEnzR6LBXqhUVyGvnE0BfaALOxKOv2SuUq4Xzd3sM2MBDAZZo1y1Cbtgbbc
MpiWv7dSWKCqTFjfGRED7u4BLCWnoLMFWelOOuyQbpt9JEyZzH5S8GoygH3sp/9ZnY7INOCBXFum
53RELQY43ILnKTNAunR6h7NfToRiC81flrrQ+pZO5y7/zxssJ+I9VyJAWVUSbTSM3zFetQakfNO1
zE8vRlZaA/O8Ca9YnulNEkMfz2fz/VucKiCg8PfXDEoJlhgmRjwl6u3re3c2Ux8250qJLpghUzMx
ZMC+JK3c2VCzFJjPbZHWE9d2dnE+715ld+7XWz56q1x8OK/GHj7FeW7Ma2J/nUc8fjF6v/E5DZ5x
4GgmTzBKT+BXrcylVTBTzxAWeNQMGgO08keOKz3BqnNPw6Qi3zR0TF7ptUnGs1i0U9Qmh0xwHtHD
cBjpnaBo7tgKybF3K8k/dS0cFYeJxqfK8mT/fGrBN/wZ0PwIV7v7QJWjOsA629Ko/BqwqZLzlV7a
YCfL1vnL+RASZQRuUGW0MDjiXCuS+9HtyE5/XDvr7sD6KHcmrt6SZFj6cwJx8XcVudkMpG9Yy+YM
FM8EXp5uCmh4jUMN8upC0QurBi0bAWpYJiNwToLyBSq1rDWTL9oEu7K0t5A6i4+XZv+kpJGkMlcF
64aa5AoBIPUyZwoRLi+6FameisE8/T4uvt9Glc00f7ZHeejkwzO/4IPZZrsiDiqKftNJLc6dqr/e
YQkOMh12nl++pCakdmimYRP0SWwjbbI3fBp2RdrBezXrZEj9ldPkVTsdYjGoo3VL2ZDMVo3J3F5S
gbofuWuLzm37xkSM4QkDb+6mMP3ZvrKK76A4kKY3qvze9fHYTqW3Fgl910CsoCJVbGicF+klEDqe
9q+dy+GQJHXegLCfa49XHQRD7xpp1fCLhvVy7B2AoLAGZe8k/9AeK9VOyJuv3emGsFa/qT/DJzMp
0XbrgYT/f2NJLlZoVhpZfhYpMJD8zmzEGBJWdKnGVvPhIy+dRAZFnNogmz0MLM9PtAf5kX0YUDy8
Jt7r6+T6JsMOBpzyrLBKfH0MYt3yepvomr8O2SVY8qmzlce8v8Bqn+rjggY/UPAjq9yHDQmMZFVB
vdsH2YOiAjrnPe8YnAShzSWWZ4nLqmkZI+ThQtfewzaY6otmxJpCXYzMoJGrv2FZhPIKbCDnCniv
iIHt8+8U9gscR4kc3oYOV7JgwvptQJhDlfGkRH95d4vBaWRfKb24AzYcqxoLvn3CAN6M6LyII6Xi
G9QH/9WmcYihiVZ++qKDgKSA0r1n1jxAmLv47bbgCCqgDRwqY868nGYWZQtBE8w4IbSlRWTCpAvU
b3BU9Eh3Ip21e3Nxg2BrHXuAQaXmk7i77UDGQkgUKfXt0Q8UBxf5Ov6IwPUtCMz6WGl/HLzsn+Ku
BF8u2sHzIkHLvRliXfzrvBx9909bEvidg3xkLvxB0APyUomdR269t5aSsapfp7wo51x/NFokkCmP
O/gRhyCeKIXj34a7PkTDHnBOhFxeBNS2+MRR/HgFDERn9LMq7KHQE9xOxV/Y9kSRCuw2rnrEwnp3
sEbExRwNdW1DUIt/0mPAX5fQY4kP4WM2Lyb4floZ55QlKEX9jyV9LYHKThfWyPr/OUrGBN8qkbo0
gEjpeF0yz0v+StPYHHWbDGS7XZOwwT4tGCaddD/WB4tWINB6Tv6wFL/NvCUfXExi3vknAu8nGX+b
01MgEDtA8nqIRJ11IW18OrmzEVFLGj5IO4MkK9cLfnQaQGPHNXgNRWjjDHwU3JCDIIt4pjHE8mA6
lajt70AMZQ18ylJh1wJ6HfD/Y55yPZ5Ywj1atU+99kUEZMEsgVxPRrGiClol0BPbbd5VjY/jTiIt
RoYURifM60fEeEH5ZjbomsrD+WeQrYW8Wm2M/7oZrPO9KtOF70G8aJbVXRGu9tS5vEj+0G3UfFT9
ZlB9PS6SSYAR13srz2IM2YQ8oFjCOhfOVEftNstGgpumRACgq9gNG9FfRuaAsZ712ohXSdNQKQb1
6YeAjECePBkdOH/AbzKquinmqEPEPDv0DjczjhXacmVmTNYS4UPzhJTh8u2EB7TwLLN9nWIfnqyR
KCWuIC5gTEioxobj9hr9aaz3N52pR19weZfFxPIwmaaUor9OQzsAfePspNXyBnybvZV2+n1PRsmo
2pToeIhhlozLfd2nALHQPn87xI23KTMOWmHUDIDhfcWy/NhHfJ74OloQXM6JuGeMW+uXJ9ulWivC
eiRcjn9mkOngVCH4SepH6IIllE77h7WGdNbrDDG2Uad1NmGqlSqkhOaonhBub88J/0DwNKY8BD45
wToC8b6agIM62+EcLVI8OpX0t3qXQCe8usthDwvS3v9t9m22mr1fnjktpErK/mqYZR4HoHxssWMI
EtipgZ+gfKcSb2c9D0gExtIeHN1D7FxOKzGdUc+n2QIxJo3k2ZsI6k+gJAY4tVA0829j0Wot2a/b
9DjpbXai7K7SE3K+XBw003I+LdrZ/tgaRd/uG5eLumMFfzwFLZVgcTcLgIJLorxe3quhCn1MEKFt
uywM7Lkm6cFn9tPERyc0NUG1//wWeb1bLk4x/7cLFRe8uuLJAD0tLdCQsdz/7YXC9HnvL1IG6+LB
cFc3zBbnViTVFDorND8MrP1PUEVsFOpGl37wW9hFgmHZ+IfDpdYBJw/RXX8MxkhtuvQbO3WWr8eC
UKtUMm7ND/n+nsAoQTe1TMCpWe6WDoGJPL3HPqhNLXFmM2pzInI3IXq1cR6oz2S3rCzhU5tDRIzf
daabygtNWDOFdqolzXoVQfdt6yXJCB6NSoDdvjz9t/aZzgcQPobEohJhPl+vwYzvGEwvIZdQZyZ5
2epAy7edNBKxT5xn6ABCHSoSC+urI50iqYOSnRk7jHHiWI9IxSMCUQKgwFuwqR3a04W2GjV275ac
8iwVWEk/7os3gWR7LVawg51R/udOlT+C/qfRlLpYGE5mVKSVj9R/tEpqfRAarNUPjDrX1hUVz3s2
TPJMS/Hy9CHhdYw5FxUMENEUVsioXOO1ROk+M8woFJ6i2dThSaJoEc2QcagX7dqIe3L/4HN5vAQZ
i24LeZ4+Qn7u09vzO+NyergB6JutQAj8TnMszzQ6cLEaVz/JWMnQnA9HC3R4BXi6Kwk+uLdER3ZL
NaXIeBHuTQTdaSBm3pks7/wWmObH6tr7FHtM7Ae/246Jlqy457Icj4IkwkKNZN9IAbo2br2uwhFx
jPF1MR4apeq7ODcKsNzVOb/O8nD4bAAaKuo3xeheppzfFdwafun8zbyO45gAMtNg6BbdlVIdBn6j
8FPvivBgbr7EgSbFZkOMs+zIH10O0wjwIEDxHrLAZYq6EuqOEthXnFA6gnLDkaD9+ldt+R47FOsp
URXqaLJlDXEiPF7/IVSEDRcvfFYa2Y6VGRbftut3LD3XJrxfwdafDs4kSxKVqNpWAyXxqqikRTrP
Z14pEk13WHqVKsfg5ZV1s88Xm7MJU92u8wUIq7qS1dXutjXS6JpE0/Tqwgx0EB9uKRe0TwI3VUvJ
0QOkHoR/Xm/aTRG+58Qi8G2g/LMzafYb6GHmoY779rae7NfaecucfM2+KxCzQIdH5RAh0uLeCmzo
fcwccy51va+49+06ZncIHMVgTPKzDKZ0GGYaWfYahNQohuriZCHvrRJAq/RDkuYSAFDk4UHj9sbk
OrVXE3MTqF04B6sIG628F4T7YfvnwCsCvwwRSNypJYpTXZTH64UgXnpuF6v0+hTiaQC4GH3Q7TC7
MJ9BJ0RtDk8Sa3HBUjs8ii6qc4xwK7AgBnsEX+dU5OMLitWPC2kMXsgO4mLsvgRfYSzkPsWl4o3W
7p1+9SNC4PlrqZLU1RQqtVvkv5te26LYdAKiZI5+Sqp+4aGXAa6pyC9xnzDJN/3FvfpVZvlxtQZS
jQgWRjSrL+dPxYA2hgcK5VB7LniAvMkZgXjBHuqtQEDWfvlS3o96aaHtp7En7nmhlW5ehSKnZSyw
yFceI2HrPlvTNgmhm4GRo6CzN8DdKi+1wKpgWyPMheNhul45tBjZ8viq5S/fohXNhdk2LWz87aPN
zq9jFe+7lkNwKfciaZRPQ2fx8Dd0TEvanel/bIDcT3p+T/Sj+c82Qv/1z+3aZhhCqMVxVDQM0mUm
yDX8sWnWLGMA6aAgMRV11Q548D1XHGfU0RBQwRAH9AsWYBNxMytNmp6ipFTNkfUiuEUkmvCSlYDb
vmxXDFtvkWefovrVnFOXl0hUxsKXVomYNHuU0Ub2WwwlNlC1p8ZjUMkQQeLNvyHO3lMRBfgEuCd4
yFzzJoYXB4CzxhQloc98RazCihVRNkDHSkE+gsaIVYpjy1q7Lnsv4D3lbz+6aSfBc1nKh+EJsqoL
QcAp5I+FmC69Abtb4p6spsB11TPeuBBZKsNazbHxQSrfA2Y88MjY2UnJbghuRJDi4/c8xKr3wkj4
cJzRgA0lDM+v2+1quHTChZOnzP6IrBT5BC1LG3MdGNrkwv4+Y5a8IIQ8EYzCnTLGEoGMieKGzsSs
pbS+O9RAxb2x9Y0Zw32MNFC+v0xMnTqMWxeYTSHV5paflGnSPgQbzMrnBaQpEfvRcH/pAazUNhgN
PEVaSBPV60eZeIoU5QxMJr1lOi5kdiMKSM9g6DgJGE5RvO985e0ZIoW9MWbOe1eZhIjSBLeAM9nn
sZBGhb/r6LIVowIZxp6EVhbN2sBbJOqiYodafL9MyMsEQj0lQiPS7yPzy1gDJHItZw0nA0KxaD3r
vToFUNJ9EDwU22edGYfdTp0zFLD8tXkH2AcaE5LMqvynP9rF/F4qX6fDCgMDRKohxJsUIZ4PxY/Q
OEp603jNb+K9cwfzXKIlNKeUkxEBbZ7PibKcE3Drbu5N2mh9Ckq07Bx5xtaQIDwmSW7Gk7Y0DF9p
xh7OvUE9wMR6/i4RAd4nV4PgM0O+87FgVT0zC3f0kViFB9U7bWQRXTxzOaZNAVkZ+QcF4kaRLKBm
QaWxoPW61Dx7fOoKHZ/qis1vGJmHyvcb2uDCa8noYs1dm9wnltEErlEkPwStpePBDD5p8HTd3y9n
mvO7gAIJXWfvQ3o5VYu3QrsissB3I02XYBwlnk+384rZLVuoDilQPPRwoa40bzQMkF3qdylFSpHf
h/TOmj2xXb41L+CvRgYl2haL+CB40YNs0NkEoB5szmLj/I7nB7Ebiula8fcyrfD4tlCa1eFv2gWj
LZqOZBPwhRSUe4HWGRUmILWpn4NnV/OMGEB+SSALFASe4eIkaaUZ4SFOBt3kg/7hkxCsKugFTC64
yIClZW+xv88vlmuyxEdmYnkgKAnQ8CMNmTVflcS/b9oSC5EwvaDlMBmLGhsIU2lFvq964Bq+Hkef
7pL236F8gi2yGwmUaIobzM+97FM82ey2eLtPaEui+/CbaTenNVDAb0oC0sxO4AhAu7YAgEgThoj2
J66D8DS+lOLRA/EclQI5Q9BbwH448quGjb4QxXOZoFUAIMjS7FgJQsOZZzdLFlo1ewEZwUnRYZlR
bfawedIycGPVkhfK4NgjEPW9dQP0Loqs0uSjW+jIZlHWCgcpNyKyzonXcrPgvp25dhEJwuBRurIQ
Wqy4IT9IrtKsZTg0rtkGYdQTWrg2+bv9FnOd7VFdl03AwQm5Oir+zsDyVMgy2py/oUGSUEKtlF6B
MQlipLXE2eEMUFczJMW0m1p4BZvdBEYdhFY04iZrT/ukvJSSGfDlozNZ1SkFLNc17ylpU2XwLKYh
hp9YxSiYGtv8sELKu4GmR4mwVqE61ZsLWgmmqUKawIbK50zF4D9CH/sDKdclq9CW7sFK/X6bx/d2
4S+iMFg+iogO4okn6/ayg3REm0BMqSWxDbI/kWLLqLVhjddStKw18zk6YnfpdnVucXreLnrcA87E
Q9nbXArsR4vJjJCzODxz86bYmDyPKBNK2SkLIKuSLACdxbthi5YV8SKakZ1zO7zvR4YSY5pObf18
qOdAw+rSp9x1DgLMdncCpc7y/+/ElqVMl7oQAuIjeDxpPOIBbCgLTpY/4dLh2e6uI7UvsJVplnXg
XSFQBwMtfblT4Q1QUcvVd70SHvQ41Cyj4JmmyGLf2OYmS6e9JWIFIV+ZfP5kNRI0ckzs5wYv1yvF
JGxeeVOGgibDbkh4WWQjQY4UvjtxDK1IE8iiIK87X0pYPo3z+fVFX6/59ds6JOmWWaggaiPoSGJU
FfhmLWOXSAXtyNvRIE/Iz4CgTS/YQne7QTbOeumWjqGtW+mAgZJ5CYJVU53zVnn3jLnzDGYcN+hQ
oaO/gyYZWlnUXk7JymQGcol2aRESwWHBhSBh8t21C1eVvhp+rEEkQ4u3Tql0QXZWUhaFxLMJiddO
v4TNqNlbt+kDjQV3/WFDc6iLnpJ5RXO3jE49d3jzUaqjT73Ou528z5BCcEyTROdRZz4xkQioJ1bj
oKC9jOAIRnR0SkG8CB7sMgP/ZSMRFD1ACujqiQCQFMnYGfaJxO0hWdMaOT+d6JwDmnrq3Kwof6BE
t53MIyCOdSBxJSKmcuzMNH5r+SetJh/GkZ+KT79smXqb1OcRlhiXDA+fq47zUsgEOitoyp26DdO/
pwekYQqJ4sPw6Kv+g/sRQ0k2AjOol4ltq8f5P3kDAXdGr9LK8jyo1qYCCrdwANxDcMbXuiw4fC/U
On+rU+58lBRCNWost6PJsqIt4+UEpJLywx13vCY4A5M9/EfLsqH4lwgRzWew2pea7071bTZszN4h
wM80po0+qMpxrPEV9bCFfeV016iSwd2R0QCqUSzZOCFA50Ps/05Dy71s3u1Q+OatkNyfVsnwXs2e
3utyGLWTZD8t6tbkAnysJ3ytBe6FoD8pftI2b9dyiRbpDyAuOrcwe1olmO9VC4YwRbgDrjLq7+Ol
nHaWIwmmViI1oie5Jpz+Qku11i1LkKI73Vw70b9Y+fCkXZk4iSgCxs4NiV5RiJDZUhkY7pX5ujxz
bNpAwzFmLpGNe/DG6RrPTFE6cXzyEkHpfLoO9bIZRPcHUaYnB+/8un+DHJDqR/PsmJNIIUAb+b7O
mE7U7i6OVj8pKAKemcog5CPlXgMcRS+vgPeodDZuD3d0FD3crq5HTYqJpzYb7AkfdmXpcFBVsIJa
Ny5k26pma8/DLBLlo+7ruGax3xolKFOLRMAL7x8maOns4HKwmwleVW04+qRZ6Sun1YwzHN0T4mg5
VS32EZKrlB0gmdMrJuqCwbfzcIhxhVoTVRq/jxmPU/W+ZYhPHQZ4qyc58fc1D6pXjHdYPzQdX555
OUufV5No85QiyaIOIp6dDeGH1iI8JHV7WWX/zy8u2kHMG6LBzyWVFAKgjusij0vDfGTTYr3wFMtB
bzPUSLQ9qLWnc/VJnYzcPEcOnGqvyYy7TKbSlfZstxTpbVcndIoViYaqjZuZ9GVhBZzMstoJnqTE
qrtRP7WkbfHFBkleJzrMqbS3wVeyXH/lmilzvTLZH2IIk9i/Cx4QRZEdRdd5+Sl/k/sHhhaVlKJE
ykXKR5FoiYcJEaIRD2633lkkp/6gOxQscfnvneufRLCEVAEEk3Enb9zmFwKOzUtqZG77lckUpKVY
WZp4SM5pUZEAgD3c1c1i8kdq89qgtCO5MuQcrGacglbUI5CoEjlxjqMxn70pzenq/bLCb9n+r9dA
C/gjWLlLMIEGzKGf7mWvRPSZPp0Xnt518L3UaRNwUXGex1+gyXQuFTvEUg2W5mNM1aErBsZ8odfu
BkKwmFiLZ+xQfbq5Mt8kAgy7FfrQZoTXkNBEVZpCIpAEJQVAH1AAdFcPHCdNQHwhtJlQKsFodH8c
ex88xum2MwgEE6AmX+FZi46c8/TvZCZW64eoy4aT+woTZlq2ylsCJu+oxWXy20tWjMzTg3fvqQZR
Vjxz5Gt5FPtyo8nVK5+E3aH1r3PZZXLlydTOjj9eCQSkPlnYnuAiNr/g4uxRQIbFNQp9f+HB86W/
fZd3xz2rZ6uh3gM5DzkrnDwE5YgCyWfZhqAF489IcXLxXeSoHRM7LIveWKBKoerp2CfOOoUDWk5H
wugNertNtzv06viwcPCKGC4qLbwaVDtKe+8zSIdO9d5l1RgnYkNMum04g2YcJ9Cxlgw0jjQzYXsx
2FWGxCSh0JHyvlfBDd2h2LJwZsYsVIN27VBdn8I71epD5Ku6tvY2RcC0cHeB9lvAF6dAxbom55IV
9XiL+Hfl7MCc8PGVZE0UEZD7y4FwsvNlrTbGVvvr0XpBnqc2ik8mTCF957FubpbpUXINMjMECOKa
AoJmU2eow3lNTTxJMvLrPeQcNzdyaBUH8iJaBroHAtzE8bO1B4UPM16Xho7HbxMzgTEQQ610Y7i9
xWAEDGXG5fnDLNoGov2pORnnuciF0/8nUfC5kUPTYPdYa5Z5imIZy+uJyTZ7oymjiXVAx2qnudvQ
r7Opqms9sjgcZfQeGwAq3frrhr5e979aoWnm0qIgxfVfFwRtSvh/UN0Z5WoI3j+IpE1FtRY5nRik
GACNs4RGbEJA7OqUpzTDWGkGa5vIOCvBDRuFnnyBJzUvPS0dUhbU9dfpjKThWpn33KZnn9fZ+oEf
HeBEYaN5hBqyxfutXzKXr9PDuNKbMPuNP1obz/aED+bNKwFyM4UqdAt0tR3Q7QBbUi12sBRRmHed
RaOyiOe4UsXQDBLQgtlR1JNBXRhnOQr62Bt4oCpiqo5aK24OJ6XeNqvS7ixHEa1/1EToRS/K/+n8
WEBrwLyNuf+hO4MPt6hpsLRXs9KAelAyBKbL1SBZOJ/yR8zXnhhBhJJPInArW21nqqX+GQIeubzV
pN2QLg05TYR/8OO3FD2cYOZMyI77KzRfr/vXxFAh3/cshNKDP1FGHq/cQm0NpM4YL4doE532nC99
wZ+bY4WM1I2DV6F4Ex4MJur8vBe5zskQysxzXDwJoILDHvlSheSJoGVSxUhFuIVBA0WJN9fKX2JV
ZGmHmi+AF0umnfvqMokT0R1n1rMkJ7XROql0FjFyxo9CdqEAgzo5S0VPGVBewdSdYBYfq5n3ay4K
IsnUkPSTzp+/0XYK91ICYD52TsvR+3q6mok2nW0tXRMBJzLKyYBRBf+7Z1Fg5Ca08THRnJrfn7oz
LlHqJXeziRGW22QFgyJka01nHZwB+VFXqGzYF4y7ifXmlrl6N6sIS71yZULVN+3VX3Kp/qM3hJdO
umi/xnONHNO0EB4ud7S5ypc2PZbNXivRZk0BhwFHu92H9IlQi/RNGISEcMUyiquCQcjJJ60lP9sa
NbOFtI22jqzQQf/ExW2d0iqN4W92uHwGOg7p3wHugZXRUdhX/ZBEjEabJ27K511QZgSeVbW7/6cd
L7Qe7t64vuRKPWQNfNu6M90FPD/BxkuuedbGG2TrwUjT2uO8ojRbLP5IXMH2wbHnGy1i0YGtfP5Y
/GS42X2dguhsnRYHeoak0VBqWwFfyK9RcvME8qRuJx6ONVEtxt97159KDq+0Vg/gxOg1OD86BRui
pOKsOTPRu1WhEG+A1hWEohVWs5I8V+topQJIIjIPnNUBG7Raob4M+/guAAHGDW3nMOBN5uXpDLLu
eeTdCh2ZAIX51HHlf6dFhJhMXCQwR7ySojLpUVO3v+tRv4n24XvLLmc8fh0kYM5bCC6r02nABCjZ
r162nUHUagZ7gSI57uzI0Dwui7GOZkvMxDqOMvIfWjiInMiNn6BG/HTKaqznwUnOPKLjsdvfqqV3
S9xREvtfeCxeuNBXoVkKfliKCXV63n+Qyrf/4JT29c9mnWJHidkHOqZYCKRV8bNtm+NSnUIsO39S
MVtqIm5p5AO0uwTO3ZN+68mo9D3+b43BoQZgVAbEFx+8TY4qGcTq1L7LUiaBGtTTKTLW9TZTMunp
HfhV60VGua1JMvRto+AWkZCI8G96B3y4ndsSUHbsFECKZzfJ2APVrvTaxtiJxVnSXOx6JoaaqweJ
kg6wGyNLtLMzDkcoY3Fmu8KmVbIJtSAWq+fpQ/IuYAy9D11tAcU8VzXQjJf0Np8r5+Ohr7B7Fa/J
InXKFih640ZLQgoEVBSBLz2tNb+IFbl/rtnS46aB7atX7nJEQm/L2ZwWpwXj3TbiaOA3ztCx6XPz
6IgCcLmT+gF7VHAXBcy615Cb4An72jlx3v2CI4v1DIvcswdrL5hjEdsN0/dXL4wFAzRkLhhhEU7l
x/YqdaPYzKzzOFu1R+zL8LMglszX5ig3Tvek4CwXqn2l8OJzuQw4OmwKVjSrQxh3+HoLrwp/WrUO
I9/ru/+FBeGG0s2UvQo3DJGt+CeYaGuCarNgGUsROeqm8r5jILjRqcPVbKBmjNJill00QImdUCa4
O/WtoLd9PEuRaYCINMRWuzbxO/CuYlEQl84TV3raevY1yoTL4e72Qg/iZfwx7pwS18i99hMHXMxr
RL/s1Oqrp5kD/9C0MJtKtEPJ0E5H479IR725wKddBYuP+4BhRTmqMNwYdtkP9bJvtA+H23+SDD6L
fzWmH5QjhtGFNrcVO++HG7+XJw9mu9/aKIdzr8skplHHd2Q6XMz5pLejDkF9FNNZZMchjwOik6XA
UCY+0PX9Endb55m5CuSSAjWlAhrr85UMlZ+JgrvuAKH5dZpbTL5KrH/rSfqx1jysk1tR/0s2x9Km
XQp4lXN5IZZQaoeRsmMFLeQXeWXbXy3k0dvkx0zVi+Cr1IR2t67v+fuw2R/LHPwmTfPHEFwGVGWX
uUFJRLOUgmzdyfwB8HqGx6kz7R1mUpL9F3RNeYmzjmq403uGwzMwTQ4kqS9SgJSBTpF2Uh5BJmfD
e+wJmPCmZISF83ofau4OurOh8tB2msLg6Ihpp4eN8jfjIYoOg6kNxguQygHZ4XdL4y4iJ+vLSya4
YFtGjyQiON4XksCr6dD8DeXWKcZztpuVyaBnyb9YIizxRsQ5dv7NDPSO1JiB3GH1F6V/XCB1ZQOA
EwNTRHLqpGcJOPxWNsD7kZiBUZxyN5g9cwh+44RE6qKd5mkAihB4cNEgvgZ6O/x19nvAlr7Y1Gk3
7APAQrGOWhMbPhti0G5AknrECV23zZDmvgD+A4W4VSij4Ts+j/pD+S3r1SU18mPIZzNEnL2pKfZ6
7+Rzyhq613yArNeFJzIH1PwWoI9TsWs2z0BwbmEaEn87FVr+mmkooIXEPz921odQ9DuOaQ+UtdW4
R6cMdh+atuKj9wSJs1gzSQrx81iR92K8Q6xfFPA6ff/a1q8qW635nSLPx6AlQqw+ehQUfQPZ/7/i
gk+o7G98zvPoaNuGF/00rUOIlbqt/BpRcQ8Fkw2Tp2/PFLhuoBzCxG7rfjU8zGeMuSwD5n7wa45d
fhSnqxVxmVKKYjkAfKEwcShHbaQp9EPEZ9OrjenZ6bbICHyelaSYrdxg34Wk4LczXZ3DYTRtjWav
L51H34GbCUxo6oxnR9khBMk1ZIEGGcmfZ/DWou5mJF6S87yGPUflWiucQhEUSDxayYz3EZ5Vudk1
2PyH3v5ARKN5zgTWqNOnr7xCnBFFhr7Q5EBffOPbSV6N8zXYL0qiCx1mzMG/OxXD6O04LPC5sMCt
UPvGRRL6wwYp/gxZn3+kDarN39qDeIedCsCchlL6FrOofra31fZw8Be5PcKS9FN2AW/tpyJ4Gc7P
4ccyyZ0f5A7242ry89JCdTefFzeyBVUr8MrkvQiW1UiN90VYEsibdiSOT+LPJdfJ3nPrDCJcZRvU
kcjtlHue0BmN0sJ+kg2+J0LWQo96piu3Z5ixEwGfdRi7MrF8x685cF9nd6zeqOL7RtwJUllL9u+H
CFPEjuS87wiwwQ7aFhasZE1sbC1zMbLgwKS4BPeFo2lo23fT0BsKgU5w2jAJ8i2R5FPVuxu8vFwl
UsTQEn1phiW4ELkdzWVLfhkcrvqn3BD4BbAMUn6FxoIHdnFbfMOofjS4NtmNJsLjWU5U7AyZdNjW
XHzTtSDJMDdZ2/vFqWTDY6wFjMyA/olvHV9uW8K9i1d0oLGTNcLsoWnAFL61HotoxBl6SkDOcUne
Wl1Muai1dAXYItx5bIZ0JKIBedH/tv1CfNQQ+I4Kq5yV31AUWSEHPuJUd5SjTHqH3EY4ff0wl9H1
A/saEfFQw/919S8TQ13O662PZiE4L2QtCR2Oeoq7CIUxr0sCdasyCv6td9/pyZLbsF6iyjuIwB7J
GXmhJDOFb+RdB6UoK+S46z5Pm4GZohNO/pRtDjOjjqdAZW7yMG4MCwh9IB6oh5H8pwudCQLV0oxK
9RTSVef/L/bFQ9ONfktV4bxGeo9g3PqtYzxPQcN733hx8njSum1LfaKhQIR0FGHRKQm8oE/2i1U8
H+54RNQcY8E3wJPrtPdmGpm71Mr2hUDVpu76EPl1nQmGpsDVvPXZLzfZkT0gvBlD50jPB44P2qzK
7/EfyXHCu/rWfL5E1O0CDtidCMj8d7t6VIxbMoNr1Q6Fu+9u9KG9YavD343yUnEVBEFQJPHjF613
Czh73lPoTtGvk3nhIUqo4MGDrxHOH1NRtStuC7RosefV1Lald1W4wSkq9+GvLqCKCUO4brJC/Y1K
VFLWOWbC46BY8nVyuliHPN37itWvs8CIkrFPiXxRUqNfOeMcgRj48c5pD2sc6vc2on3Cq2Mt6+vn
3LxJ3dICBQ5ERr+iWWYpv+xTT0EY9NvJ0vVoAd5WXofHD8VWAw0PwJ/ctP6Ae6jTX3u2khHp5INa
R+Vm7NT+zJk1nkDHD1sEe+YmgXxBV9L0rDinTv6viUH1S09lpN0yqjAHcWPUui8rsk/vefh71j2S
h9qhYEqrBUibVeTJyvRodUeDIGRFlwoM/5BUGDZwe3+jFCLz5eUgA0DFGv5ej2wd/52fwycJjVdc
Xaw87pLpBKmzenYCLretcomWSmUMSVOScdNFEyW4Uu/p/6L7mqJQaYo93WAnBV1cQZmDQ0thlqvt
bupeSVqgP9gxGJPHq5pHdmivnqP2s21bQeoxzSZG4Ya5idDB0I2ObP7SCwbYj2H6grF5v3KNURSB
6c8HOd3fGfpyvF2Uwv+ZGEKsmyAZEDVUY4HCFc1J4aUGcLvWLcR2WCJXGYthxgTs2UX6Czfk9+H+
sG3j7BZll6dUZ2u5Gcp9lkqD4Rw/w/Jb+95X6RolXJxIqqeMwoduLuIvhNGXX9gN8BUfnabKco3v
HzEDw+bk6Uofd1Kc/dC/Xs40kVKzbXknDBjHlJfJKhjmmHMj5mcHiQb6zJTOAdD63EBVUgpUp3BJ
upHEiUOPJ3C8xhuKA9KfvL16ttboC9RrO4szdP/Kou5qyJMsSBy38H1XaKv5AE1jNQ7yhW8hxEhn
A0RHFfde49gSVSk/dpnlJQj4wh4Yot3QXVgsAtM0pps4f/zx2gTlD/5EUWEMU5Hs5XCR+80KtFxZ
avA/gILbrdWftMFwPZD+OmBYXLA6S6b0lY013/B//Y9o5xUhT2U6PVhsb1PxM2S3gF8Rlm0xNb5f
yu/WtxvN1iFx07gf40mADDlwmXjNqMDtL2Ql3NtB1bAukP8sNh1CD/GbzS/WHfxjLRdnq/x2M5Sa
4T5LYwODnUW9vNwFIL7H2WC946UJ2ESUJ7mQoWApR28Ho/wkLOCNqNckUErvFvvmkybq1vlUchOk
gJJgNiARhtm1ZUwbWn/JMO8NPIzKLmvmUaf+XmqB4LxTcKqtHfk6VMLESyJSS+kNb2hDrX2dCl38
vGvPtAocDd5cre4dRIl4mUEx0CK/DargmFV3nayYTSdS37DBBXqlqSjXkry79jK2e0qOcKkUyQdN
By1h4ulgyxrp354F3loBCZQJYdcF8z8Lh0OiWDr+U58DBmrTZoFliD3meNi9DatH0lE9a2F5rb07
6tebCA17GjBTZt1DrA1b/x2JGFmovSAbnWkS/dWMCAQgYkfn9hMcFsWieRFZzYm88poqb9xqYjhQ
daiCe5DlwrKu5pgDPGDki1N6uBsq70tuBuln7JYa7q6F+6FNziZ58buXLStaK/A1RTFY0lnd6zV3
jv2ZE2J0JbiktymjTsmyl78GIPdtaSZb0iTXaGmf0GyRl5BAACdQLZ9Qdwu5YDIJjE0EFH2seZus
WgPXqPjHwPHLnN1WD01HOhffsiUcinnGByRWpeJu5SahsNF5/W4bamMdroP1P5/wCPzynJajKeBd
FCBQ6JoYgleYOhQV3Gk3RVzSw/qpLb20OIjtrD4G8MWnKVX9WG22BUB26SDVbr2BiM4uuidVnMC6
/ldXRRPP9v2UGvJ6a1jg7xWu1Pm1n9N0BIqw3zaNqBG50gOSl6FRb6jWgiqQ+aPA2lb3fj/2CvE8
jWlPTTJeao3L24qlIE8BHvt+P0fwmnLPBHlOUS7DNzjAYOwEVMfszJ4hbgAvJ9SygM2bd14w0Mxo
TU8x1DMAgs72d6MghhltlTDd6WNCAAGU2ajtynE5zpGvTDjSyKn0p+2FMONycyFSNf8HTR5ctlqM
+UGePfE7Unvfu/nbAHFqGB25Di5HL1C1bTiNYZFa6C6PoiIiidQNcqKF7EguBPoMuQSeOItPoG4s
EAdyjszA8zOFPaHu1aPtrIVPNZbQkqfSSOzFOBdSqBuanS0+kRdhFhvBPCLGQXZNoAA0lo7vpQhL
fiUBaTWXnDlIqLkr30J4yQXoR01QqFHC244u+XJv6kp3mcCwm70FdAoQL2yZBLY5s2Y6LCmAUKlW
u40uJSSs9AmfmS5ZoIdTiaFDCPWGm9+XGh0BZMR8Q//GXaReXarxXPjwvlwWGaQUFc3Zfuc1hso2
hWqXMRNQXjy5y8ecfq7TraaKXkuRtwrfLXYfaN3p3WiQIAdj/vZ1M7udVL9d/nX7dwy0OKNxNFwm
4iZJX3DxvKub1hPAWTnvVBNJpo1BNvFsjWecfVYnRlGMFmipnR/rCJbjjS6L/V1WZ039nr/R9f6R
DlNTuNF1v/K5qRBmb/HEAhRDuw9ePEIDH5p0nK3sZxh2QG8ak3mwt2KUGLMVFXy1Rh1ODrY2AcVs
h2HBZhscyTobTpgFZedXjeeoPZ5WH7wqVtQhmwpAiPbo1NaGLGwaqltsF5FHMUGoyruE0cYOpgJ6
ang0latRluAZn6sXdYdB0uoJ1q/uUmBR903S/ipDwjPDTs2dx4ruri8QAcwA9Ux/g7A0iWs02uGX
fLeI2suT0QjN9xHKaJiTDTYV3DQXmfWycMFOQdq4tmqA3J4HAEoRNU00sbeSm4r+5+d1hz4yK2P0
WNTTcZriYNUbDTUn+DnBu67ICDhCz8cY1xXChoopqbJeuPNjKAQci5yBpksiA/PRiKDRtT7HCtV6
tyR5U+UeiMOika36DJuFabYGcg+/CMEVsZE5f0/9Aw04K+or9Ko1QKQxxWiB7C6FDgRpVmeDW2GB
EDCCYInUDbbzUVneolletUMGru4Wcf34DYZt3G+ZK3n4ZQa6yhVE8A+g829L76M+VRDD44N+VZeb
7O2N2DRc7gpek2FV318lZXAqKtKTb2ZIWA130qt47H8aej0itJV1skIqAPrMVJUBQe7HrKT7i28F
/6xkb+V1Cu917ddOyfgi3jlHo8JnwdM8kcc2fe2KM9Ci/GKzTQ6E0/7kSLg2StbgnHsJk3lfxNoi
JSSjAHHHASw96CIF8pBoLzRk9V7Gv144YS7DNYgbW4h1oW9PwNxuANeQjdk9vx18lqyujPGPnTHd
qtkudT5SUtGxAuC3sipoiPIKOhOJ+fy1QGfiU4io6tql+LODr7eo3+UCvOT2B8DPsOYcC/SdYPZW
I6zy517Be1z3llNbnhTe/6JCT5Df5jN35QTKsBTxzTpFPIDi1IjU4b8fklyLJnuGkhBx6B1yoZnN
t4vh8cfF/tR7Y7CtLvlhQAjfZs/NVm5Y7bJ+lqXhD+lcypkUzc5/WhMkRxpNvGK/FRQnhSEBgoZs
nzW5dl/5JQ14FEkazNNhnoOAMlq3wUX/BbBt1pJgNOcXBv/3ylzSzZ150DBzOPKnKFMykcudDNhu
DpLkwEUgd8qS+8Ug5MbFozkBSt682P8jlZSme+uHlfr+lUGT3dF2D6qtaOdBldKOOdBQVd6whT4X
hYUBpW5xP09bnBs3Xu8lbq6G5iy6DetR6x2YupGZHMpu73f5uwshEzpZeLVCeHk0ChJINX65dONv
DaPmN5hF1x/wi1Ry46lQI9oTMzoaKDnlBMsN9025HAhsiLxc7e5+IwojB0JvRlL0myU8uf6btv3s
vS3ESiOof8dwb7Y6qDZ45M30VYm+2AhXZWMKyhaNWA5Ul3N9QomNOshBtqANLHT6xFDg7D/t35E4
yt7f8vFEYggwea4cs671LCVMebpgTQtezzKaWTMoAwRDz8J99UHhYkvJ4XPFGAKDpqcbLMyhfgxq
HElWCw37uasqmE/8LEQcmx7RcImcUu+ZN2eeSyWq5erJ7utTykvpQiKUTSB7uWOWsp9me+q4b2Ul
+QgMwoRykbXdbU/rEwNWbD5ZInE38msBHXlPZyQbddSJ2ERynojjOot4AGuNBqPJ/BbFcINK3pAP
E7WON+h1Md3w65zftwtTihsJ4Fs/7oIhrZCiJvZHtz/+28hEWiZ9EA9sd68X/cu7cm7RU6SG0xwN
7ApeuzBZ2dqhW298BrL4pE3Dz1YRQo09E7KNr7tbivtxg2WBTfhxUfT6WaYOvD7J3qgtY8tH2j0m
EGQUjPyOGFWD0EObxAb3ixHQfZJ7+Sgg82tNHc4LHK0G7bcF2BqWhy4f5AifusTO6JTzkflmD265
WS8DGZ0OFxd1ns4q1g86RGCZO96MmdKV57PKdpDqC9/5RlbSRdlw5u12Z6IJRFyOp4oglYF6Np9/
VI2wkaZBSmzvLPKcbhteiR4bSow9RXlkIgLwnGeXt7vPQmR2s356ASpav3x/I5fH+cS8EXpvsKPw
ra+/kiPQL0Km2J5zq0yBY1dkizAnnj1yf2SUCQbkAPEgGWeoMmo5xPmiy31BQ2/dVNr2vXgtRX0h
HJcMblGnW+D92pAYGa7u3FoYn1nsBKISK/B+GaE7TWJL9C1jC6aK6uPpPH76/JLaw+stDU7WjKL1
jTxJ7tSrbmZ2aO9PVBe6mvXlJY93AKiQv6QKn0PT6mmZBuZiFc1l9bSKm2Lt6njUjLUKUMcZsw9s
GfIHnBv7EY711kxdlGJeWgW6Bn5ErwLG0LxlWAC5jwqPAX3zMg+iV02QxC23eFtMZfB6d7daADLZ
xWucLIZjRsPNrseVtxapLz5I62r3tFSJ2gIXi4OdpxHKpVr0kSnPmiXeyDMKVuC50ENeHkne8hb/
as4j5bbL8ecrKe2gJgkjBzwYWPzlZwSd4p0uLD4QwDIXZfzJ6mIyvLQX1h9by4toTt4sJg3yxvEI
OKSfNBrshnP7/imL8UL/Dy6qwy9xJwFJSv1NqeNE6iCO0cAK1HBm5tFLyq2aYb9l45T4sdT/iQnv
gdnkS4PtUhnGTwI0SyFq6u45r2msVqVpku6PRIcEKOCEX1+vxKowDeW+Hmtthzg5Zd4w2RlRag6z
2uCq3WLzflZnteuu4LSvoSqGDfjx6K7Jjanb3DKNJvXzgCB9nGKkHo/ySIE799gyURseE+N6T5av
lfIB9tCXfhh7jjzQEZYDYYLNnfCAiX4YIDbyMAbqihEYD/Ro0SpH0w53OH86tQgvEAy3Czw8ogkd
/B9ZHb6quWHoTXtIANIT7C+NN4E305NwphaI+sKLPFISypPVvx1vPMpGGYS5D6r1q2YeDpPLuHMS
W47Qqb1sa1ukrFwb2TXO7yGqwMOZLUGopNBi6auAWLtz9sxWc4yQ+F0Uh6t/frUvzRWq+8nukJp8
yBJENOGHqAf8PFhgc1hPJsOU5GQSB8GtcNFDYeYXxNlliUa6CVKi9g5QlLUdRXXhqZskkzl+b8RR
mehiATdQUZgSMLhh1dd0xIq7FHWCU3GMlTL7iF6ChuJIi3RfsRio+WbKee8EXjA+KgzGMv5irHjP
5FPmsldVkhB2SBouIQgmX+gu7y5wekukfFhDnnrBhipmCo3hZltlvEQp0rpk+InJP45CLkr8LP8Y
uP0Q1atphusHAP66OOs9pNxC/IHpvJfSRSNn0V3nF4BLvcKYAZvbYBUPD7/WOyW8gGudotV3vPOk
vO8Xc5AYhckWtCsu6EvaH787iiiwy2mAK3aQt8PaIirfzWB5SrpJW4N2oC/Q23Ufeb0d+tSGRcbY
8zyzfmWrV1sAE6RyZN5e2A+CMpJuFb/0/cP2Rc8IyX71/My90WbYLCfi++LbTXqNEz/BwUl00X/K
ruk7lIPAdZmvmN4QZ1sLBgDae/j2k7qPH/NFZeGmLvaZKbQ2rm55dEyCGtDtrCh2IOA0fDr/MrV5
p31NIiXDMptx4CYCkXfp11vVqN+caX48BInPaXpq7gmMv+N31qoodMB6tAi6AFeLFELDSc7r7cUa
V+8kKKwa33XPP3KXxtmHcsqlfH773RnDBdIS7knjfZcmncM95I04BEs/c0HdQOAIcZhFmeJTja7d
MDZ+MA+UKYNm2t+sgg54RTBAZP9tsFBoSUJLe4zNkcF5GbVYuuBuLzKgLbmKmQLLSNyFh/lHnHTP
c03LAzNCP2Jy0WiWd2lnUmZoG2EijPfX7z/XYzl+cG/VMVDDkm66t9Sks70puESR2396DuTkBq39
O2Onf8h1HIx0GIvjjURmTA8PRnCoXa1/7t5oGrXJeRDqXaLaYAAjvpsajfj/rbj9jZX541seEqLk
tZbtvFfL7twpVOgkhLVQH19zwBfInDQa1IQWZ2dN+3RPjvaVoD6viYSP+jfo/cN9vYj+vumPyIy3
MIQ/XJIZY15mryOywXITEQE140PHAemopQKpK5oljGvcMsilwVZsMjD/F1sXkHoHiu2o0qA8bOQB
k7aKHSO7c5mYXMhTDBnLP0GHUndn7R9AxbnpE+teZlk907RemJQbBVgIB82kvKagSSEcoArPGGi6
VK5oU9hZ913+tGvulAT4lwDvU3r8uzdw2Y5dP8/nS4jTx7ou96m73EiVZh8mxbtTeTQRswhhaO5G
8ZG0vTzFYXs+kdP9qOUd3dHcVUgZKWNGX0u3j88XyfuI9NDRQlKnKM/r0o3FPEZIpJYQgUhsYO3G
BEWzQQqPvzmWYmDg9FHrDgfJE63Hvdn3G61ildrcsEMm4HHdpa5sUWkL0XWX90sW3mcXoh3XDBJv
Msxv0tJcsZu2TNmgYrE40HhNKlZgJhYb/S57YuyxKGHWO+t1IcGtgfu7reZh4HRcMkhF3FV9nf8Z
lcEl8B0hp7upMqvMnkLOuBELfY4Aai/R9zzCqdsUZvv/WzFW8aLL88uQinod2yzCeF2BN8oPojaa
H+cj8BeoybHWM5/fgpcEqcRdLywEKqt+1BXezi9raxS0goKVtRKtpLJCGglHdBxMC3WPefWRsDGe
QEdHfVNbVfpMpNikmwhoYMSvDGSUHwpOsc/6nhUc1naym6DvFRrNvn7d3a58RHtjRSWuPonbq7Ka
H8pXq8k9aHe86Exa6UQhBxkiDrzptmxIgnTPcLMSREMlXIVZLRViayPZPWxzqYkLwWyjPTTENS7i
7k/HmdzbiELiuFmkpdqvj2KKoKjp0Er/Icc5r3+qPSr72x1Ax6zYl16qfssQtw+Xmx4gSoVJ1Dk/
pN+mrUuzXDMYd2guUQQDHlc1zwoaEbFsn7XtdZ3HelbLGMmbdzfJYHL1n2SWdYvfp1YjoPbAw4qm
a1mB2HuzS/NqZ1zZ3PJzuZBKHGyB83z7J94+isFbHZeCqwZNV7R7N9TxeAfdnTYgju6wf8EY412K
t0aO0r6urMH7G5oT6hMrOiRqLheRqKjDlCAgNaxCDzqLXIY9H5lNAvg/0j8JD/5HBYdfR2t04i7Y
rNchhwJH1mtrFVKyN9Q3GeIrKx3k1L98t/4JFnHvMU92xGtDW5vAnekUyIOtkHGYf3wir/mMUXtt
23ovzFSAqKXy2nJOqmt7DTyLRfnddtywXWBBdH8Dc/ov0LHxVqh4vJo4zYWZv0n3zgIp/CSx1xQ+
21kqkuv5EaZhZEM6y2J6a5D0p/QGGP+f3unH/kMz9LO7lt+4LOpQVnCIahPa4ygvMZqruNwv06cy
UEQEHL7Rg2J7yBB7x+g/CWAZ/Vh11yXf2XZha0BvUEGeBjYxlojBWXvlFFBb1kwAMRqm9aegQUqS
mRIZIHnACAH7C1Vo9zlUWAUtj+3kT2IdNb/y3r7clyQBKo6gQtgpA9WrDqrNrTJzpyG3jszt3gK+
LBj/AXVLNlvXh+qQ1RBZ/TmfgK7a/gd4RbWC6JdoxrfBgQh3a1RRDzxl8Y0eWPgIZ3cxKlaX8Z81
R8nEJlau0NsZ1C+x4qCWLQDufwDfZG3dTnNxMgxHWb0RxAiZBJe3/sOH1jOmENFZPBw1zxyKIvff
50TrMTzEdfgE4R1XAWQdweLmbnkzjWr6igrLYX5x151+rkI3lpRpEAGKdIwNmAR1sAczOdTX8g53
IyvH0bzM6ZFV2SbYX8Fcby6c5IhNCH2Y7oSNqhGYVBhVtBBPjWBJRaLnOkjdyBNcrPVTuOIfCTwm
VieDdIbkB1/tXfipBP+A68436WPYZ1enFfNM4Cyp9eqdMgnMG8qVurANhbluj7N8F9Tl6UVqcdeb
iuZVQ9JLu6JrkCC8dfECgHribVD46AcKosUBw1tXjl19HuyjuXWclg3vHWMq7/GnDLD5B0bsdEyP
88a8NYK8FGToytUhMRaXLnewHHDdht46s4X0wpDem2Nzbul/jP3xvhT4JPlnJdQH2oF5n8YgJPrG
8pp5UChvhjahPGnMJk55BQ8uAf14G+LL7UxHSk2WtilA33ypTZD4c5aD2kSSoB05U7a/+BM+hJl5
wOwTUNpESHPQB8qJFBWlqysG0R0SCXGHxSuoE2LcLUqVfvumI4UJsoyyS9pPgzGhY9SgcCscZfLX
fIY25v0O0nLCIC5R0sKNnKc6W000gU4ek1J/2BGeYVRE7jcl1z4rtZeH3SaqDHSt0wcHcbENxRH3
hXReS5iEynYQFjmeXSVBgiGC5+A6f1lVl5cLgtZBNskkq+azd8gD5Ub9S2JrKqarqjkBKjXNs468
iLNoqOAt1DqJXs+DmwbPF3IJe7QwBgk/buXusGbl5Fp2auHPJgi4F9tw/D2mwudiCFdbsrWZh6SV
JLqcyt7rXeXGyhwl0HdhhwiO5uuthDE3ro5C7wZzi7rt1/o4QVs9NyThlJ+sdwzPIh88fDxjqjSm
OoD6dwIxOKN/ZWbn/4Vtq6kKE5VNWPzF4KE9sI1jPguAF9mIE9KsU708satxGxTYuZQaGkBiNlT0
n6PwDdwpjBTnQExBQKv+gqiVn9qpjWBUEMRpiYQauI91UfUTk6yvpBH4yB2J8rwEi/qsmdHaG1Z+
Bd2MyBwmAb8+H52Sx+4sfM41vAGnPphgLGQIBn/EK+XzEvf5+A6zmi/93Tc186p8Gae8cw/YtoXm
oLguT55R0JdTiVpDfBfnloDYTvMmwuMWdciChLHT7Nut6p6N5LVbmzP1mCoZiVl4tSUZpy4olLOt
jMoKKi6Dm8eo0Glr4tZQodfrbF+CpnQgR7hC/I8gx6Y9QLdZ2siAD7di6tvip6Py+RiYmxq88w1P
YbTflF4OFEqrF5nrzeUQ/jg5BvvTAa9EqtBZYnGN7LlDHJjspH631mIYwiAnMr+74QjzZdkIS1SM
QhLZRX9pz6EhCAtReiwPfUT8650JE8fh/x21wvm+u5gOd6/ZIFfy7KqEJ6ZFJeQG6sbABX1UAjg+
9Tn5YFn+432LTMxSaUPqQn8eD6HzpGaGwOAEM5masn9Zh/9yH58s0YouM+ejEZA63LLxAFTISzM+
NNrZ72keLl+MziJxf7PfWGiQ/HoTEb70He52cBGSxs80bSK3koSa+N0GFG+mliTW5cYECZidt5tX
SclHoXtP5rpmoMJ93P/cWpWfHNwwi2bC+0YdNpfvvxgOybqdievqFh/9BkGQYLib5VwSres6A+sq
OgKllNRm2kOQ+qlP/6c1xIKxsYCQbnPowDjxNIJuuwiLjgyL5v8qwoz1YNv1QbNQIZxpUMc68Axp
JuD+kGiBek/tyaeM+qNJ8tLgRE1zhMR1/DBoEfO7AlNIf8WFuUoBcs8pDWhGIN/XGuv5zYjEtXJT
ojjTiuVQ5A/tr7rPFL3WZxcMzIZGQ/eCnt15V0D9Y6Ib17NX8yjJFeiW0h8ujUDxcxLjkrtUH6xa
vqlYV6yAPgnz4UY58eN5p7EFujrbOq5iXjEuX1BDLeesMnFk4EqR5L8PU20FZ9Ol5VlSieD49f2F
IJLjP7GEL2JavJDDQ2VOOWvxGAU5+o7dyVtY5UhQSU1SK5zLcYP1OBCYX7Qjhi8k3ivGB/z+8228
lo6AXZacjxJIQSEH4HuNsIMqMBwxXmu1cWZoojblxO989Z1IRZ5zIwxWoNLjG2WziPi1f2t+HVYG
DmTbAsghPD0MSjYXfNqNhZ5lBaXvvP+dqxdRtme2l96Th24dNhS6bd9OHU+eOppnLUeTuxkKQuJk
PhLtMfvRekR9SWNSDxXGt+0x40vMHa9C/6PTiGp220e7BBQwUql1eeGGl/kSaLBZAke+uihrvGWM
QzsJdXMk49DoIkBiLAYO8GxefWjvF3iVOx9Qo+AxfBf+i+ZsUBIPnPR0rlbbnSPTBr2xEf/Lywca
J6ivty5X099upv6fNvZuFarsUr/35QgcCKZmLM8CzBILQBPYlZnj4iuxGRZikSZejpwYWQjLZzGM
IyFQnAQjtmIHpNQKUGktz3baspulxH4irrvm+blVnMJigIZoxtSFkrvXrIjlYntHklHHDTiqc7ux
cV9ymuURudSS2jXIHsN062iFLBWQsPtPkAFb9lhfG9tIEXwNtnPP3ZO6CIoow4XW99GTQM1xFinF
HN8ZvmkfVvQFTH1X4AnUdoyHpD6xOw1PRlDqExEYd2lMGfwcI5mxM42NcBJl6zGEzpOVGE9eRWw6
OQpHxW0c9EhtPnODZ3pbe/mWL3sBP6dV2Dy51O4P2gyoagen63h3t8Z88Ywj+N0xh46AlOt/ScMv
rU1sI+tu81lnrtCeEsbDz/mRZL6XaveQ7sqjVYR/jkQKc61Rtm8mLk9/31luLAJCy2H7EBJA16pf
7D4T3/cxea+ZTE/jYqFKaEfF6IegZpeLVpgzafL+wsH5EHznsr+K/OjIPubn65nQg4Ohmsj3zmEx
nFu39891jNhr+e1/btAV4Hx7qiahKoOSaUyTTxaksn1aoIlAmQO9xz1xx8TvAP06jC13LTGXaMB6
nGstMUqcydpWsqNMUMwNUnGXo8XDDT6HH0Z4LpDo8qNe7Iymt6/F/vxJPVtoOGuamMRS1/bd8p12
uyv8BA79uUtrN0pci369sZlfFl3aFPxn3DiPSg6qSXaLKg6r3gHIIPQaWTsRHAkA5XJPuAVWEF0G
2ktMtON9icM6eRBw/+mvREVPXP9wKFxSEg1NCIc9QkIz8f3XRgjgU7PVynHK8MEGwqPvaNkVPW3o
EPYfOF4dnEFVauYA2KtJhc1yVNJnNz8WfuPFTgNhGjEDbr4z8tdeuiRIQIQEQPUvm3V8dGcjxgit
ZPSWA29OBFLklkvX1PTGClGl5JLHLyzjrpQ6dU1I2dPBxrOz3d5ch9Kyt/+w7qt+0i+X0TUWhC1g
kFVaVLcUNXteOFWx99aG5qNJiLycAr173g3zaCEBODkHkjKD43uLsl7pm35yNZGpaVP1u7j1SKyk
NpyV2aV8nHiaCUQzJKPLwTjhbftJKJmL8YkKwe4pCW70s5l51Hi4zBF46FGDLU2DQqgkqdWJpzAE
LmSC4U/Wi1GnV5II2p5VWeBqDIfUR+uGhvjMQaESWecnHuXhGDx1M/kpYOy4q5Xv35N3BrRH2CGt
Qic8/1dY3CZn+h90hJpUlu9DUsn7El824QiALkbYYQYOG5uEs71gDaVUI9Zr7BspFt2TcPIqoi/d
S6a112kKgByfyEgTmEt8rZhQyhg2i7QYKLNFhXWHaFtX4l5kCJ0nkSsQ810sJ2D95lDlnbiADZGQ
MWyarm4h3h+4EQaUehntsrAx/sj8bzBKVW+5OhoY0rJwyx4BYh9T94+oBBUDNDUs93WI3NRNwZin
FSLd9WfE5WFSaGqE14wahpbPpOgdTbMXA6tye6E6qtc325H9sdwsDYn84DhsxWRsMMoej+F5CQji
sW0w8vz0ZP6YwBazpM4EDGZYPPucz7OLyhZEnYyy7olqOk1c0nbe89M+4rr9bXchvvuWWzJWq0NB
S1dbnSowkC46835aYlFHi0uQbSQbdpJb8bCLk5kqZExt1IY5EXWaCzJVbVVlwhQAxpfB9nOZ+bQM
Gz+aU/yxqFbdcxWTY/O5EgEcwAuxqnhwheZ62O8JfcbJZ5Wzj3II9ZP7BlJ/mmmKl7YDCeUGB/kw
GTgstF+Ys4PHktiHomyjyTIWVry24YpbCSPH+znRDWiS7qHtKsolVXTkC35AQVQjDrU7H6XZflWd
hIjVAFBxyJkzdq27jGN7bZjWOEaAvPqdhDkFxsNrf4YqBhahBsciJDmXIksVMApP5t5rdQtGtQY1
CqtdrkPkDh7SlwEkZ7Xlvg3zF8G/lCSGW4Wdm+nJ5QntsQAbQmIwm/2BarovM9HbkNDhuuofkulL
X7ReSjprCGhGM4EGnQGIKhyWjSBGtsMo8OwfgHLhS1W0r9DDqaGNvC/xJqew6uuYSam1ZvrpHB9j
21qOinztP8NJvC0/60a4rU+3HqSKo/9ZxmPrKgelMicENsY+Y/VA9ZVunVGO2RaFn59Q0Y+viCeL
/vPCjDpHy7Rs6daIhrdv6jxhCaEHi4+0axE/KVUQJteHghp0ijgr+Cy8aISeRIcM/t5foLCz9mGr
PApmOSNjUgTkWyzYMM8PyXpvnGYcfiwf4i3aYlr5VepDlZkZm7Vgu2B0eY+GBXoBGFYcu20fOwQd
GSKrwPCTI+CuX4uALS5Nn4SxO/JynX217B+y7jSOokxPor12tjG7GIWKDbQjyqbEpeKsHNwjAtrE
ZaVBqhwMUOmsTkY79TSG+XNpCq8Efh0LyRgT03stuJkZrOHhlp0h5zai94bZY75O5ZbBRdh7aaRs
0227WjzjKKYTR5ugmnSxCE3AZdqQSBKjIVWt03u6A9zRfwtcg3NE5zyVYUfLjHSC2TE6gMHOAlu+
znHWfnJH0qGGaHVOjNxEAGIG7DUtTUCnfl3XBCXe8fKrcyUqarapZM3MVGSwbShw0KwSgv5vQtE1
G+CAxoQzP2hpaV32PLvKt+wZVLm06FxL42eJtTBuH/iqWU5hhOuuHZTViisAlFxm+BUYKi4LxtHL
D/np57qDFn6itTAZejlosUOWNc9r2/8n8XIsOd80Q6zXEiWVeL60VvU9j3eQYRThBkqstm1Q904h
COV9VOxgVI+d+s1UJ8hwEBYGDbd5nsUO4kqddfV6ISJZeTJBNrY0YSE5zrTSqLp/5xgkMYaIkEBz
Ge16ns4hjE3iIHidZ9jg0uzXMERytAAX9sbnXjKjDpFJJKAaTSi76X3gI8DuVC5IRo0L7pwnNPdy
SOKaHVf9G/gwR2fhzWz24GtBp/j7bH6E+hFHa92MVEUmA+2pf+u3fKc6q7QYz6xAib1v7c3qaVAk
zoFhvG+/V3yxD+d359yohQ5J7UBaGg8Kl06sM/K1AJRDLGi5kni0wZHcIdsshH8FwrVEzdByQiK0
goaLvSHTqJ1TCMhumLDsNKkEreOTLNrf3+hI76C088PTn0RXmeU+/F9SvEsRepTqxFhwWIxosPpS
LkX7vXSH6dnQ/dDDGTVYhxjT69LzlGqH7mksc44NzUzIyj9g+yMgEANNuEpCXaiPXQeHhCkuWprl
MvpAh8u09+KfaUAnMikZWAX68d6c7X10/Y/4mRST8DGHot3MdjmHbXEvIAfQxtog5nJWkiuYivRN
C5v7BF8XkYusID/dulBxE9cwAVMyw+9OdGJpHEEw43/LeJAQzx12SG8D/oe+Jc22+m1O3pZNuELG
eYfAYxO0UhJDm/kSIF+cXPcXYUV2p5KDCg7sFmvhqgzXoOUiFHCWofX3MgU1LyrNnNHAMC1bvALr
M6yfoWeRLEKlDzX+f1aN9AeqmbLCLpjcHxp1AXx1UeaXFiLCiUcv5SwOslD4IT4dvlSdAZgA0sfA
MHRiDn5+9yG1vb0u7O3YfF+dJo/JcVQf9XP+Y1qMPIpovKt9MFUEfDZfwK0X9E7PVLymCJK9ShNg
1YhyPCfS7ZLl5YTk+CReUVK+lLjyiNJ6Aj0fLvonNSks2CG8TnxKv57aQzQI+ZftuF6v9ON6YU3N
16OQqZi7Wy4wNMIqJGrllKshwr7UjEdVZeosoVXnmjd2urweLQ2L2K2L+0zja/DN6U3G/O7JSwGj
bB4KH+t1KTTd3OwGEQO2Ws+F2OoLxHJY31ndzf1lA5FAa4loUbx9CTTEamdcAw17AUok0rdwTACL
6+dYXsRRCwatw5CD+7ra4uZjSENSbzRfFRnYdRZblvF6oWoKWNZfcMZk0qWo+MFTH1eFkM2kiFx5
F8xPn2CJtt+qcuB30zM890TSR6/QklgMKnu7O7vVh6zzFla/IuT88L3N9e/zN6qhMwwESoP7F6bt
wFmzEtCJsuVEqWjmS/Bnal2NQQIGe1fRNUJUWnbXFadszrVF736xpSsxBXksCcw28U5nuzVIuzs1
z7cm8K0qHItjHotJPjutdI1OoJZDGlzf9ZrAS9hk23v9KCP0CTj2q4mVng7H1X3jO9oyPPOMryxn
N8M/XcX1ZegB2372fvpieGc/xbwKf6htD7uf32XP919KptYEa/XuIcrTiVAbcdra59h+I3pcgIPR
6Pr64e8gnsYTJjtI2lFfFn5VX/7WzW2hC2/Rw5iJoaY8B6QVDszEII+e4p8XZFDFP0S8ATOrWLdr
8tuMHPkS7WnJ3p8cWzY4Gf5WBektQurOe2NCQtyLQvk3fkpFMeIclrWwZ0lnLyjVg1qOYyVsG8Nk
/M1DDo8nmF3PeZ78W5K/wpB3y7W4KajyhMslh+oGWVBP9faKRLUSnx75SwbXRWqulXpNlqE97Hx2
OlxZSTieJWP//CdQskm4BJobZLbVWRQc8WbUGCh5bVt9IPzTyhqmE0Jp8of96wtUKWNhuW+DFpSi
O0uXGAmmfLNz/Z2DfuqVKTUKh6ElZgkQGGaJQsg2f28RlTR0JcwZYNNjU1gPVnp9n9s8q9QKceqx
tNFsvnycIZQmthvUz0mnl+SPe+HyEsClcO3AXO/qmAOH2retstVHD01ky/tNrN9xBEDWztOeukLe
0yLsuCQhyh+S76vvhzCdhWgjqiZs6d4MR1/d++UqK5qeguYDW9BKAmwk2UA2L4SXrtS3gavbANMo
/b8sVz+4RqoHse+w2jsdqWHlnga6ZTozSjf5HUCbnbh0X81rjqYvrcwwb/Cp9pEBPalewkAqzfaW
kxAwHhKBXbbGWMivu5CVPy2YQT9WXRxnUp5oruHLcp2qAHRaGLjNFNig1/Az/iteZduz0PyrRALb
otKocxlzhncCeOC8sIzRoyeac33jqBQ491hol5P0EFazaMQ+CXD6YrhOpEGuvuTYsxAPBmt8Ju45
Xdf2tfzVm1LkZ5obYuf/qc/GEJHe5mx8GId6fkQZX8KxijNEQfSHnfliNri3z+77ii6tCHnKRSoR
S9cKfGjntdkCewUszBGHdVdZTqhHBjLWoK2Ws/+v8anox6lTQfWUNGG3+aGIPfJ2E7KDm0QrzIQf
U+6xj73xx6Grq2XqUM7jMZEysH3rKY78oVt9fgb300Vry2BvI0FsiBjnfzq55NY8QYDA9K7QUJk1
IBycmvnkwaE4X/CAJrlQxp2b/dFv6ftd3FBf4zL53GJ1D6s9qhhfo6C+ZMPm6c454sfc5FpPBtDO
Hun9d48PLobuJ6HEufOB2FffrU6zEDr8ROqNq2WQvjSxTJ7nXXPtSBxst8r4Y1vkzv4RB0F0OTCj
GfXjXDAdsABiIfFm73IdRw8a3lxOg2VtM0cD1QpPuTtmscsVO6cviAzESjURQYDTlKveXQ+Jeugm
sD1Xstesf4gNFZVVzN5oJYIR1+kyHKUKk5v0de03oHv7wwRtXS+mtIcoMqGIxMDmXWwAEncK4Rug
DhSgiPB3SFh+D5Jw4I9DCZIctJZKnz6VnG7mTYrLgxDnvL665UT4pKuPq1Rwp9Hr0Qc286MmwkpO
Cp+EC74UxEJWJclEyhwp/eE5ObKSuP/jCtzoZcOlrJbp6YA0KaoDL4Eq21MFhkFXo6S7UnP8DaWo
ZMNVwTj+Tcdd/2yd1ayUTqJgbZgi4Wvbk2WjK6tibZt2foyoWU6YXoqX5lnOuJDB6/OTVQGWKNoe
GK2uFI3dfj2t8OpQ/U5ci9pTBsqfcQsumjIy7sq0INNeVO5TiatUzynxzpMcw3zUR7ovjetldvdu
mPWIgENbPszFv7kV9m1IdwTDblbCqxjve1Yv/yDXaMLygp46O2iBBu9B/7a8L7wUuqX8Q9B2FFp/
Mu8TQ3BpbfToXAJ6et431JZ/p1VEV8kB3oOjMxWUWI9hQWmnj45McpEc656Zx84Zx9r129mGqDUf
L95Nvqwh1lPepSkiqykTkKKjY76ZACbbbq7McN3rCLsLswr9tZ+IyIkqhn42yTrt/eoaBKvrt7gD
8U2XNx/Wx44l3TAsLPJqtCIey9ULGc7zrEtdIJAtg0TsKgiqZUprmJCFpZf0PASw2Yh32yItN+pw
vQjGgNMEyZ8djpgIuKKPEMLFKjBd/R96HtwcSGiV9jhAI5YH84ApdiaS2/tSDEYWSBTBupy76Yns
PGTD4E0tGTmkK9BvZjs73aPgh/EmApFpLZbRmAIYX/JeIzEKHcdsV+pmydEKeKQRS/QhI5uAqNo9
xqTxd6I/A0WD6VRW+lgARpOPvO7Iu0er5cygik6dpY8tU8KUlfA8kAx9T4afKYlkr5iM9FBKTYE6
sq/nsFk7OutFWYwZ80dHo+JNF/YFepZj9TgNWdtRdbwAo0FzUNTHpibBHiN5qfeGLIJl21WZmJEy
vYVEeqHZfpGGvA0+vILa0T/zTNl9YCmK3hS4tbpV6VfMTjZQeW+4OMf5tGjos6AO4F2ZArWRc7xb
7EBM3fjlI7VbxSDI0OgU9VsHvNSeTcsPfMaaPVl7Hfuej9vSTR3dcVXlSRLiOjWjW3c0M/O71EKw
vCGEjj/+V/RfKRscfx/u0hbfjdt1Ub8UzovWdC5dNf6b/dVkzFvhuG4vb8kVoFN0OpC4N4IL081u
Hvj9uB1/YbjXiwV82AhP7qIoubS4Tz/kE3r2WizH9GIn5ZuxTU1jvG4r/hTGA4dOrX4R3+b5GYIY
0drID0IWTT2w0RZUygC1HWpB1anosqM7sI87xpZG4tR2icD2g3hrJgF6BgwCKJsS4m3l17zT/IN6
JDULvyNKC+RH48c0EpG4T+QvsKaF8yIJZDkm0q0TiY6MzpB/ESQYA1MGG60a3l4xKysgyGzG4e+Z
tHIXlk/BqUovrXHQnXaUkK8q4EbPE4XfU/4fGYeu5tQpiwgF2N2+YMDCGoqUP4gXh/HGN/Mjh0kD
Lm15LyH6uDJ7XDe3X6y11K2zHpylJNBseR9z5Iic0/ihk+jaDN2ENXTm176FQc7SwXvcVJXUV4We
hFpT7vsVKUMQo3Y5MVyDZcig16r14jnG6p3vl4FSIaCTVK5j8o9chc5uAfmcswGxPFa5qrlJL9Vt
daEKzCUTFopbCSM1U0Y6HH0FsCWy4Q/SWTX0JsaLlns16gZkfy8hcG1f1aL3c9MLOPkl9lq5DglM
+SC9iUyYfD9aFXhlnZ7/mwcOOs6rqhCSGTpJ/Fkq207yB9iDTf3aXgk2/VgjkHGFKeUDFwGlG5s5
/z8PySvZ9AI1eFSJqWrOC7dZWMwLnkkqi08SVy2gJ7Kx+nCRJjr5X4H7hbuTB9Hw0fItgLkLl776
50Bmgm3lEFm+DOPf8Qj++OhaX8W/OvsSw1Du+Doe8lvDuGh3hPnXbPh+02CwjSWlUjupOjDPnMbS
lzi0vEWlB/5eKaNV7QXli6VkYlQ3fsF0au9DupVlEs0jpXAmLqV6qI0WwaitP4QSitiUiwp2vAdO
EHCz/lUsNb2V8u4AQoNvCH3Q7Dv+P7Ma/6/OT2Hku8XC63n6l4KvcuP8uidWxLRBWYwGhnlRz9w/
i2Aqx5IdF+zG5kax4dM554Ih2iId/fGtXjIgELfuwSkOwT7PwQgiNlgYrEfNTq2tCMl29V53zgSf
iy+E3i+LJvCPauIlSqIts+4kuPWGu4E4cdE168Ugjh/xQn2zcNTGCkEPEsqGlREHK6F4+AYXc2xk
62E3qr2LEKHBf2Wgc5vClPuhTJzsA6PYygOAB+EgolAdA26MoTkaaQnPrwbqBklQ8XwTvwQsEGS0
jxzN+4ARuXbQbWMeimjYDj4OdXAGjePA2VGL/dgEOnHDZQlNqWHrTED1vYDvyEtLY0S2mKreG8Hr
FNMbRG+yA9f1cFRvrM8lC05gmkkoxlbcwyREQOQDlTPCfHxgP3ORsur5HGr/0suk9ZGYUskSIlUP
8ZWsCOoctTVlpOhrciiToRKyZ5o7srFRT0NN8yYrgskzL1W3iRWLObDwyIybcObBR968NKdkhO3j
n9F3TaZWRUcJHgBN9fQBlZYTeoEFS0DciCBLcEyGqtuTLNGPBo775mhaqh9hNmpRPGeND+ZFTMQk
zvy1sEe8z7nEMkE5dkGOfhgI8UQ0M3JpS8+Z0vS0OizXxjZNS0qfcpy/iyECShdnCjQXBhi4aE+E
k02NQUYP+J37sE5/wq0S8gET4gCaxQtR0ROQzyaeOhibnALclTfhTWSXg/KcgWVADQ/D42gmbfhP
rlWf52w+TEaHi/z9Ezra8oYB0+Av96+hA6andO99RwfSiEv5xoOHabggsECKtF3XPZDHQ+66qzyb
AFE4X7IvjkV6SrNiOtIaVFw0ZxSlj0dsP07YP8FvE/qIwbwt94bd5lZ2bPTBAxDPZDlvlT76oWQi
Stpzb3oF6eQ2bJ/dDfcvNiHd83M2/WBd8rCcABSn3hZb0D9cqxUEiUSnMMk1KHD5mGPJrLEYaMnT
LMLNgVXfVSDI4U5zxffVbszXR68lL/qq8rL/m23t33pChWf2ulIrXNzg2VHGsZjl0jAkwI3SUcET
1FAnfS+42cp4DWOeQtW0GV0rLZy5diHhvmMZwcCw1l4oL+lp8hKgHSLXf2Z/9BxevCYWVWZd6KVe
1LTKoGH+EkJRydVPonXfW4ktG9PzHadGZEl4IlcUQZ824TcIiFQu4C2zt3Fp/o/vcwpYU0rLhCom
OqqF2iMRxVFidkU+NODldip+onpNcYXpVjgaTA0J2Wkj8yi+aaMv5rKfee2Y/Xj3gLg9SgXsQqv0
M5wzZsJURFKROalYD2ZT0zUiS6KRPyGyLijeUDKtuLwtpm4yck9804VOAwt4GPqN6SFiQKHWOIS3
XYuRwElmdJ47jNM4NrDArvAq0wvsF0FbNxIWeOR7dkphu6u7CL/MHzAD1rHcKa6uBOJPb8MsV0Kn
uRYlVSP/ohgsC7LbHYn9QPSo49xZvJGQKNkphGxusdh1PHYaYFU+KA3g/YdO6HUlZDSDUQhtTjjq
PnNVWLv5DbWShPPUvRfXCS7+jRHbWGofVzVSIdlzfdwnD1RUhCfDqI69/neaMhtF3bKtlzx98S3U
/VLETQRPgBa2V6MI5tvPWuymjXFy9LNqlRu8Zt4O0VSoNFjoEUKNmIvs8lGbDnneokLKfEctlzKq
0K2zUMRF0PtZs8K59fjEhV9XTRcmLqnP9xoMHNg27+aJqQIMrofe8AE0ghWonZcM0STUnXRtf6KA
PkBw9XvUxh5ncYXF84vVEfnToJudBmvZvNwEYhv5SLapPdtQ1kbxeVUwhQlfJ3IlewitmVDX6wa1
nQbYMfMzkKlOI51V2nxW+mcvGHWAPoPmeoovp7KYyhoR0ynfIb0uE/GzsERhj60Vg5mRqgnrKl3X
rPwnF8iuGmo3SoQtfRsE6EUH3zzJRdde829gc6ECh/VLbZs4KA2PuIAsxQgUH3KiUdlx6MO3VcGT
AjyCeA3kyrEwwHgnoTHPMEmdxNxU9G9987wVzWuklYfHWVOsydZj7l94/VS6RNzcBPT7DptqFfXv
9a0V1adT+mpxlM0oslT1uJh3gXcWpw/HNfyc7CFVhHhy/CJbzRNU3rlC/Z7YfWyR2tIcASwyByGg
wjg7OHd80M/9qhfj4YvS3/DurMeQCB+N6r7ceMpLJGpH7pssBaLTwqsjRTo9vok5+OjwFqgWEsjS
NsoJO+Vib2mlu/mh1Zs1K4ufbcigJYkB+z/MwbqIFOXrJgOe6oPx2u4Rg8vpknyYkwvqIsNGMO08
/idHykrvEqGYx1AyeH/qHFfC/QpR0gFEBjsBmta29AeQrBpzweITLRXLYL0o6/0vlIj7zaqQSA/r
DhtnSYsJ4igEbK5Hy67Fq2Qb+Veff7jF89EkdG41PpQj/gLyMmIzW7VeqTVDLHtB+L6H+rd+Dum/
ra6pj0UDy6Y4jBzSEhXUyqIjUEttr7oYQplikxhP/hrJhfjgUHAwudeBSA2SIW/XJaRFpmIVmWJm
K9O8k7rQ+NUZElZ320C40Jcm1NRyOZ1BOztXSgZo0MQaT1rsGOQSykAsmDSrOLLSdIg+OIksiIum
ikzTO0lPrU22GLuRBE4HgjnwGw8zyDd1K5F9+kcvztl948KJrV2AMbegXp8SOYTKGV7OslFdfZ82
G3z9vZUlyxyapYbZ+n6S312BmuJupwowxRO5paccqq8qNV9GgiRTDiZzbg0GaNGaMX4SNY7PrqxS
8ILUO1CaadZFB8HB6gSP//fvoSC97uOnHwNAkJSC4TCuQdfVW40U0zdwmVrW0Vr4zUQiJ0g/0oKT
RwtgWw9qTNilDpch591s07NYPbI0L+hH9wdMVzM7665Qie/VgVBU6+wYEHVqltGwp02Nn0HL9Zqw
kQv8Gd/pCeT6ylmrjJhhVFnQVSDWFOoqOxQLDysPjEpcrNWD+PhxB+SQ+gbmzymNTsf3Pi9pIqHc
z2/4MBl4Yayhfb1oQDoR+droEWrs0+dKZlAUmAYq6ebtJTH3CLrSzs6itrw6OZ6oLdnjp9ov3bLS
8EiTspSKX63CubmIFPuLtjZIhUU2BJDSE7l1OVPtHLmcX9H1/YYkj7VHCKtLj2R2XlYw0hlVsFtc
5ymuO7A4K433IUeW+OtLVUHdcMddYPsDmPm3V4/ESGYaUVa66eBqlePgS/I8F5kwhx7bZb3k1/px
InVdyCymRhEc6HivkPaJkvCQkq2wnuKYDrtkK+3QrhMAyB5/obDP3Y+e387VxZxrHxLWbWPDXq+J
nJQzcmdGoZGKT4KWRNcVV/nsK62XeoDuaoBv5nDxx90XTYFioRgEfrGJml0Hja19U9EjRIxVSH0y
tlOpXd1tYbwuxmJ7Lg5xoABEeacykjpcWzC8vLpldtgK1EAJ4lBkQYgmItMHxCA+aERyuxKHdhbp
BpLD97OwGK4BYoxYOXnv2j+5pcwqgnAjg5reYebpN7NCMHcJ+FmNXu0bixr75YBc3mGt+ECxvWG9
wBHNdjb/cpRklAOJ1gd7JnxBCDU9apSh4ugAC/7oAw9WO2r0P92D6EfmxV4ZAD9Gq/QWjIQF0lA7
0hMW+a5N8YFtR1reFMsKUwEyfmv2SFIpI1K1TwECOta9CVooThUG9ilDCsVcoq6Ug8ApDPRBYuFK
09aRZ7rKvuDdA4NYFYUShHsEnV4ghcYZyb1ZU73kpgeHLeNEIeBPdlPMvr1jbAHFlKOXNjBlhjRP
iBhFTsVDpE0EP4KKWqqejlA1orV7NVZQ0FWhxRvnJK+WxGSQZEWBbp5akKKoabHY+ENr1Bqqvq14
hQ5SKmMWv1nxD3FUVtKOQSm1qhaPzTgm/Y/6xT/xDUD8vAM2XvYRisJG4XFvG/2ZOzA3sl/8GlGI
7jg525nT+uyvZYMbaKrMFZ+h4ETYldtdFB6f6VVKOIDKGZEDVpmIW6aQw1P+ZaL9f2MvR8Xhq+vJ
V3Y3mVmc+a4yJLqmWcPUJcl+GyweXsz+qerGUfd/rXs9J072vH2K//ZErz4KQaZlfAcEio1q6+Bh
Wx92ThJW74UBu1Xhd3iSXeZCNNjujxjODOZsxH3ereul8RtD4sW9k677Zn6ixlc3bOfgV3prJqNa
wQujxI2JuFAXX6/7x9kgJFVaVZHFlk3hA8nZo3GatoGz7xWQoj4/E2KMiSwlIEeI/3WtObLZP0rO
n8RZBQXlCsN8zHtUaGbwJzoIfC1RgqLqvc7AcEjSXG6jgx1YzkMBb4mxBM5GsVgEcAwN+asOh6eY
vF8VyyWphQoHG7Xn2OYDmsbRMNDGDImXh5xMA8FNqIul05bmeM9P7GofMJn9KDR7xGjsBv3w81UJ
6tDkgpJCNzGi0U5SKkBLoJRTX70FwCti7LR+2lSw/UtcR0DtPQKKumH0c3g5KXLekoixlzXNck+P
sPwpD6yER1rLEPdIWlXWyI2nXteU2NsZ50YF59o7zlRCEOx6ry4c524oBtWu4p04t5YnEtK/mPmp
1WPHqLh9+cUpeFPhrT0jUikipcgh3FfR5Y3kXP6H/F6BzlmqLXEgq1ZXkA0HRaGDMWjfRnpybhWT
spg/QzKOSCY9DYSwd5ZY4xFh9g+umnNNfZcc/FfHzYNP/ibf6zg5xde9/OECwD95pm9ogmLMViIf
rfhYnMBfvnjfttvxIV8XZf6lDEO4SnJ5C6KP324486NUadIEB5sBLjnyHY4GFdsa/c2toBSgFEuJ
wOXw1l8LebpwG34uRGsyZGL6PNBujphHxnCokOTrg+f79t5O419V4tnDnlFnkOAdqmHV5Z3O5OgQ
wUS/PrQWafbJ8rLBvLspYVf9hmZHmEIhdA2nQdfYUcNHyJXiiI1SfltMyLo+lIXX6vMn0IP2pysQ
Qi4I/4AAmAHKWNYIhPB+ZHeT1Ftd2OLC0SPl1Z/JQHdZgB8lvh5Y3qxraK+uCggaTR/9kamyNtvJ
h/CDK7a3w3ciFauLwERE651p4MVvfFMTrN5Cq8O0ssjnektJB6wCRveL5tnkwHvfEo8o4lJu0kBy
FUsOxdxycisd1IFzVTofcJKdwZod6PUflEI8HZFX6fs3oKbENMZPy3CW61JVFfwnSMAvtZ5ejkok
pAH9k3LnLO7LLXBchX93JdHCPpgW48h/bwJwDiRumOAglwHA3a9vUH8TYA9n0xJJ0cTjOsrnMxCm
QctUwFxlWqJ+d+1481walUaIP7QCzutmRsosT2OfzDa42NAl+eHnG40PNAV4lMogk268ZDCH5wY9
7nivYdM7k9FlTMHqzXeQBsmPK2DkCIOl9yDsQCSe0PI0K/lkX7/2TdEEec5cMbAYOnwv6rsGWWCQ
fkDT/DIP8waYAzAHTR6+Nqbzs/vXhDj6MasorlfOJFyiKKbYt6WkMQ+yy8XE/TuBzXUeSIoWP/CS
7HpuWms7QvT6ns5mDK/EGwyd0e6Q2TceC5ucB0B0Y3QNg3ErFCRjmpooYV4E7jY+gqEq6j6/fJ0z
h9Pkf8JJjvuGnr1/c+7EUuuplqYd3M/f2eNEMmn+tEcjkOvgcjK0IDcBH9MnIdKiVAKCnQz76zBD
s/jc594GwqF/Hm6tX3HWdCEPSmYUMaJ3OlIMEfhgWbuGzFG30K5cDhuJHuUQ1558QYFzDdxKmkJU
6zyoGH0rNul09LNXlP2uuXH5LiQ4yKiHok2FdoXdXrAR3LXBFXIL8ZNSeYoasYslbd/UYymJowop
/jCy54DVTxw2hLYSNRjAG8alJaUJ27KL4l8OOTrrWGtP51z80X8Zsk7ZDj8nQGBaZHAxGn6xVfde
MrFPMzrwuliDtIbwu4+4mGkIOzxyN1gGALP9FRvcKM0yGSEYrZiI3a7oeuUMzW1RfPVeFJaF0mx+
Zs81H0SQ8s8iQEoMTEPumLxAIUY+I4H+MhLpt0Vqn+PSfscUv2FvYDlbCF5iGqiVwK6Ycz/GC52T
GBjzLtt/nA7RAsa8Az3HkYI9o59rrsn7up2QmJrNe4cHDm0ckog5Y9rBST8iR8aOVtrPpZBim8RU
TUWNoy82X4ku4qPhJtGl+YNXfDjIjHWHvRNkMqnIHAmrK5fiexbgvTSPcelNiuyVt0RV65fn+6DQ
FsgWEZcYxn9Cr8fBOBoJRiB+9kHpHDCmnZ69SHTZharW3nTcfSUbt2ZATX32P1SZpqp2gshzrjli
m2FJeXNVqLiWdPW6ba44KaC0nON9aCi1VNB9Kbgtt13KKGNjx/WNK5RGgMG0qoV3sTW/LcTOuc7w
dRkUbXkwuY7NtY/45xlQlZvi3pBmvFSa3mtNm9WKxFGu5QqXHZkycNF+WhSD6lAnFdkKX/UC5C4d
YSzvHGI38uH2LjOYqmjWT9mVzrNw2viCKcfTtrkMbxjLJDw0BRa5tnADzrGJ2fa8iUaQ1QekNpUt
7IJ/j0syln94vPcuYBYV1/M1WmKqiblCakGL2h/hIQUq3E9HkEf7m5BjGWnWBmOiKlVdS06lTtPc
TUJMqqtPTiaL1e8CICPIU7cKwbCyKpo0MKyxTeozGlFBzTrDpNCH522dBJ3D9axwFuLABVwjuKlQ
EahTFag0PuqdXyJJsBKgtOGae4ZRe9xQ8ruPsej07KAu/QIx9yz6UbZhiuxPKF8DY1HKGqQhLkRJ
q2w+oNaN/GffSeb6kc4qivgrh7hh/2EbCXiMlT0XdTE/8u32rseDr+3fS8Zh8DueeB5notawl+iv
WcEK1w/uN7thzfAnsr5z6IVLB6CBKOuZuCQUpyH6k64cRbRZ4OoyF2sO96YtZ7BQDzMNvB8qUrMh
17LdeiNp8GM0dCeYmJrKJDT1Hpdb5Jrhr1pxv7NJXuLM6UgDbU0XXLwtb5HlvJ8l7bf11PHz3uQe
KXZJtiXlI1+FNLVBqXPlmujyN2+0Aq7BuwPrEzquy4yEgFd0RrN5D2KmSEM3ldNQFf3+flIS6jxs
xXP5BSB9ph1BGYJioQ+WXuzySZLACS6JtH6fddQA9jP607tD9k22GwumU1INivnFMBOxitqZTWAE
8Q8tnYwSpWYo1fZL6mRnTcOa5FPRMfDXB6STfp86TayxLu+yrfLrf3CvJClTlbyrqlHWr0cZoVrq
JNyhHbjhWzHZBm/Yy2qDZhD5lDBrQRKEYUO7iHlXzKYVFBSn6JN2Jr877CTcaRtdrBkmS6ywR3g0
6lG/paEl2Vu/ZyHZ2YnrlljhPzTYoek276NORl8VUf73D6zcCNTevt02dcNboc7tCdWkAXtF096x
4lo9yznuSxFQJPFmcErIED7o/EIqmfZHn4tI8IwxGc3I7wsIxzmFtOMp4Y2K5C5sG8X463CONEq0
lm4a6p+YxeN0mFPFOsxXiaq/rZnkHTwk62hKiO/67dKao6LlukprVQLXMUldR63TL641+/cao+2E
kbHaWbq9mV6EXxmKo0Fj0iLzyq+R70ftgkg0UV0wZAhzA+nk38lmhRYkmFdvft/ckG2JUGhYbbPv
AbrocZ9gAZS3r0vKyrrql7EQC3EUI3imuCv5B0KZaQHSmcqlmYe/zpdrJWyU/DSuXUrZGMCcb3iF
hWlotgUH7gF14Zuaw/ciqXOF3diXZcH/5MBvmt2eoFkgMXUuMRJGYRISM4djWqJPW0ezj33BAhky
Bwik5j4Tsi9ULV8qlgbkptLsHrz/1IZ6PGdHpFLNqkYLRm/IQH6f9pJTJWX6O0U5EjLH46e0mSM/
ZK/fWq9z+W/l2H4RCibO5tN7nrwdIdScMTjhmRBjNlN/8TLe5Kmm1sxJ2kSd73TCqqMZWIeCymQL
CPURL3eaLdWFYJ1MI9gnDxzkoGwc8Cy/lXhP+sph5v+er5NCsTFbw3fsafHOc4j4WzKx9uMNhzSZ
Z7loLOEJd2wJyupN3TEUjWJpqy9XGaotQFHR8+ZPpvHfsVuyFsqP1TBWpLnrpnqa2xbgab3a6FTS
PH63+/DIqW3/CP0NtxxQ4/BwfqO6h7QqVHyBNjSYkF72dX4kWUhbyNJPU8kJE2vZOiv3g1l6cQ7K
zrXmp8TO6OBYmOARiIsWnS6LwNR0BqQp2StR+hSub/MSnSQLms+E/zBExLWROwdJXtWOK5c6UQ+3
lB4Pnxs2r9WRLGDpt/I/apMRWrdKdgDtG2Dle0+03FAddvtrEjBaeZ/2hMAZlEjystMoRPNIOFMv
YlLhwlvojrKc+uE2fTaOayqhYGMig+91XizdwLFA2seYLugsZxldcmX9hboQxNPqY/1hXT401RI/
NH2DiVnz58LIHR0cQ5UG2eXY0V3zN8P+Rce1wxIGCSOdozo8ArybV2ngB4cmapPhq3kgy1VAbNu8
quhYmNyROgm0TXxUM6ZM7+MDQfvIiv3ZZh0e01TWQpSvHlYsAtKGTpSXoHZm1OtAR9aqDvjR0hnx
1bMRcHM+6sCLdVPeQll2ff5ufXCbUH2pQSG5+tIRkgRGmSQYvpeosR0JI1pFEvanXJaxhr3ScTjq
465DbjBh7YBsGvpl/udbLeczO9fhwDamMjrwB2H115ymdQKxtDivc1kG3sqYAG17NTBkkl0/LUSz
U+vP2bacbTpm91eNwyoczBtf4D+jBI/M0VM9vwcedElgytGGyOGTBb3leDo6/pU+f8N8y+kzcm1C
Cy/PHlmHUSKsqvNmULDJ4KeAqMk1iSzf305GKuYMrvp7G5jRBe1jlrMwyhksqDaLznBPflnDyybn
VWvSpgHzbnEdzqMtBHCwcr2PVCLzjZwKmNcFZU7L6mMnCMLGVaej4S8tV46wgCJn1g68oRFS/qD6
GrTozF+TRlJVfzfhCASEsDW7V1+E3ohYY3Rq5zXS1oSXxCDpW+9GHD0gk8mPeRc3a9pEUBkBug8g
ULBdhiOUYHVCg6/qFSe1OaUplE9IPn3ezkHF1Lgn1qMdJBD75wKOX0UO3U5XymUjaoHp8GWhiCCY
A6JNjI/PxdN7mm+YMqoM7HyfWAUaE94YDQ8SSvdXHEQulJY7+1KEUqodRCh4yri2enndcUZC+A/X
P+spu2XcqvywL1k2KDC0E5AOEMbnNpWLZvPQDxwXKe8+29RtvVqhcWTW8Gn7ERZPoLMF+fZnhfdE
mBzAhugQ7na6X7TAhdIE5TJQiw3bA5zRlOT4xrHXFL5Q/CWrkj+oD/ec2w72fLKgShxcU/NpjWgt
KkD3hC9+gvNVOWwswBZ+DOBLzUC17ocFf8/FZiYpnOnviEzCFgc+r1he2yNDznt1f7W0X6z/WD5M
7XWAjd5KIPTRZDVoDIIL/NpuGg8F89G5XoDcEZP3JxGQpmRVjX6m4ksI/u4PQ7W3/3UjvTnhnKhG
dRjN2UfPcB4ohwEzWmN4QJPiZh5NNOGIUXGpMMe6s9bRmlLalCW3dIHUFK63h6lBs7T1SpqA7ydO
9aDvIR5ZRehkiWxq8h0dbvVeFX5rTL8OSaQJYJ328VD0+WxDrTKrPAVMFYxpEw5nnBEj6NTAwbpB
HxQ0M732IYpeOtxG5xkztgMqgKlur9Ha70M2XZUn1O7Jpbqp7q8cfav2u7vmA7coixEvavofFiap
EzLEUbEit1o88+9eusRy4H+Lz4lMP1ErdxT4kzH0GFBN1S9ATw2PSYxnQ9KlwBeaddyt43hNPAen
tnMU89pqCiv0yhFYHEe3r/O7CfOIXPWVsY4YgLtv1pGq32YCMs0+/yUlcjG4ARUQ34yTrn1W3lKD
SeHaXHUcm5odNw1+tHFTpVGfHCowXBn/eB2wogL7fIpOQOErshnJ9oxP1iompGo/SaA8MOWTTzS5
EgS1iAN9fdNdxw3VNaHHPRYUMAhQ3waUqtOq9amHnSR4mtVNvxBZAF3FeMi/J7u8soUKaGvWDd57
FQLdQpLJk+s003AsJw7822GZw52FunQhzt3xAC2NfjzPN34akMVmg2RfGdAdt+p8sEDr722lDKxv
2WuOcRM3ZQv1+DUFuXOTn+7Wkb5cg35E4e5fxODTOmRy9x/1fqTYy3+xZbxlwqVrzT0+63AsVoTu
gVt2lU+XpBAzN1tno2zrhtoHtCKmG1yFzUTY8xM/8Wr71OIbVhq19W0AiTJjDeuTGwQmKC4NYVsY
IXL+iZ09irJtMeN1TxQ9w6ahO5hxHA4fecNjQfghldG+ce+zVJrZ7ZVwCyD5NM9ikEUSTbu79WMw
gixRZ2TtPEzaiVr6eWxjH5qKeQsXiwBmDmHJd8PZ9y0L3d2s7EfyO27MpbtGiqpahR++Y/0ryokj
1nDR2SH8PwwGMp2H4F8LuBhvJfbDF/VJ3+T3zVkGA1SpKNxiQKWUM3XFxWqSxAzTB/FYbgqs9X/2
aDAn97x6RyPAMUvnL7a74dpSHLI0b03+LSpbSvtQxO5AmwGF6PrruO0WmxYZwpWqRyaUATs0zaHn
XniGgXs4qvtgHj3TB77IUkspmrEbLhvP1RGBuFuPAhHSP8eJzhTPncovDgKcp6FYjUsI71Js8ujm
tW5DfYVgJ66r74utyjTjd3p0RjO0vncxQEZxTodh0CfDj3EqO74LzjKgtmUVlQmaI+x+DMKTberl
aTuKVAEBFMc5K57iZOcBfhDkkJn76O9WqJACCqaON17j8gNoGs0yFS5e6jzCCDx2dmhspLFT1PVE
IPYEX5+yjrQnmDLs+Eo+nolbntYpoL83ENoSw7CqxO8uxsNY6CDyPKDdMePwEVDMnS6cgaNKEbD6
H5O6ytFVchln9vzaBddoKFhjsOW+6+gs7jgS3LcKwo0+uc3xW5klutHfBCSej+eNw8HA0ZRye9Qa
i63mCTBTqgl97GrJaBxKczkWt0xOH+XLqPvZQ8U1cRRDpYu/pSiKpGHryjho/XsMtRwP5FTf5IYS
wCV0ZazCzq05BigXeRURUP0jB/NaIEpjIOWYyy/AYXukJ2zau2UyXe0cyly+Auv58HvImMFWcSuk
z4cpycWrL6STBYW3ek48CMzHjhbGUweqtzUCc9gQ/gUVnLAAWqzJ/1Pq9EGBGxNSQAj8Tp9CZqAP
s4Rs4Pxo/QTRJ5+nebFstWJGZaTs1fAsTHZFCUbrIsbSw0IswLY4A5OGe75031sXPUmlresMoqvD
BENSOJA69TGQe+EUSpC0p31/mievg9BzaKYIhHua095c+YRlxjbz4ralklArA17d32XcGlTydZyM
UAWaPdnIp6ElQi/XvTDB0xKvwIOqzKMtwaRjYioogaOqV6miqIyf7vLhcKDKkIjSLp6nU07MLw4/
CsVlcaXI1SKssCisy/pMlfm2kGGatvbXuJ0dlXyiN6FOVEys1YyEw0JN4NR9rBfBLUgoiRFVHxR4
bQrg4X1sCAqErjZ2jZMd8Q/OPyReauMFiathzsw9iXPb0hfj98Jqm6FApgFMSGsrWKWijDfIJlyx
tE90JsjpmQSH1gNTfQVh+9rQ1NKJOYo76EYR0uLruvQlUQbI3F46P7bfE/jKYmAq9GBn26R79UKn
RYbqSLafux4KM1HcX8WLfUualX1TDL0sDDVc7sH87uDwJKmT20kkZCmVGxWewAQQ2RyHoJ02x0jf
Mw7qA7VfDayCvqBPkke25J7n/xTIkyCSicqUiia+xr4xRFoe/UeYnC6Ogc26pxQHx+cV1KXdONBR
LicHJAOcxlD648nOlGvrkFpUk1ozKixIT25VncezDjrvFDaV6YCAZh7Q6Fkyw8zDr8NvV5LwG/vZ
n1lDXcK9wte2Fpq7IqmGObuR9ODdddT18wmdvt3OnDWFvRCDlxBpPjAvY8tksJln/tUEo4RqAO6i
t2zWUTsS0f8djtCGgcMfwFcYxaY7cp4zdeAiTW60ipyNljRdQF0C3Rkv05t7GnRFpuzFDfG9w5zl
IfSVgiqOOz2M5VFZTINicfGG0vFGN5K62sPNiQRzOHjzkeg5LDjnhcbTFzgIAwoeapyoStp3FBX6
/VBPQe5S+Tb0ZjjHpqi849/BAgkzM+X02REQSJB3unvJgzIoSyjs6dB/dgI9qo74r2ArAng67Qee
1KUUydWAcjN/a7iQLyF9Uf/5mbf8fFTDf/mRuthyLuz4vRPECnNiiD3AYBWLppzRfqdhhkwYwEDk
WmI9auo11wQCjwl2htvzxeXR0NWVXnwr2cKaJGnmtBQ24uWUVFCRuu71a9vVFFyhHAsLuTa9maM0
DaG61C0d/LU/1dNuy/4D4PzmjPN9uzlgdW06AtJDUmAbnrP0m5XanjEhlgmVIzIalL6iCqBwT19g
SuhNXNIx6xrrvB4tZJ367MIHJcZZ2KpQdfru+u/Bj81LwFRsVYQNMmsDyfkko+gJqwof+G1CpTUN
AZmy67jphEXqgUFkNCrgazJkhNeYZt3yPOvTQRepkNKPOHcQkZpHA04KTln6k8+t4HBWZ7HCwU6w
ejF8ZpQN/4tn/jq3QGE2fTyd3Ut48snH3UGQZAWBjEDvSc+MgdeGKUEll4Vy4UTpmmH0gblkx7VU
BgtxQhJPE+PHQiJd9P4gKLY22n8XRX/dRTsoaQLfDphdTe+04RnxobRnwyZO9I/g+iPlSrS2Y9c+
ksElB1ZO0NSsUQa22oiB5mqE77ZQf8hGbZkmqjWXLF3X8Ch+5cz4HoCgi0BThDJY6t9lZY2MfmnV
DXYTKMYoxzWkGgVHIaAp9BSy3CELDJfxb9Kx+xk1J4VEO8mR3BX9N0t9uqDoqnTLl6v11pzG1Wib
HA6DuyX/AOqpXBNekPuDq0Fh19KztEjFdpvvX7dffZZNy7BgpNRgOg5q/35pi2YbIR9C9567zcW5
5Xjwm1HLm/h1h0PzpDRruaPzkcFVMbEIdw8SiFfu0l9rxTIrbbKjrOJBNZkmyt+KYba2b7b6ONia
1aR+VQiRwS72Afbq5Vsfdhmgqa2vgiOpzz8cNlsYKe1o8GbIhcETF8GPC9Xd0/PtPr7FM4orDHqz
WEAkgWYnrkzt18NrZcQYaKEAPRTagUp/GuEnxesGOkbw+cmfBoL0zh1f0Er/4MyBc5UIuyEoUY53
BMWjEP5Ds4zbbMWDy6jzj25XA3pGBf1Vl02DAvyn4BYPXLpVya6wEWholsX0lUTsuen1d2ncgZ3k
9+359hA9igIpzgNSsy/Redv2+xirWTxETppJklgUQlfneo9zcArk8UohmLwS5Old7IpGY5GAIRLN
WAjLoNXwTlJ056rWQvPLpxLt3MZQFIqlV427Ne8P3kbvWR5hCphc50rxqbOZUd+9JF1yrE+Gnd8q
XOndx3IcScvRrd1r6TYCJY8pnxSTMhNlQtKgqKI3hir2gs6U80NJ7eXgmZhF+owb7VhMonbZ6Cjk
tzq7QEfNQLIsmV2DIu0K8gvHRcRzWZYOdjbVTlUkao/8tekcfEaQ41TISHBwfoCh7YwIRmr5T9pG
aUTvu2uKSxrTVzrl6kJmGCUYdwuf4JZhbcEtETm+tqIdKeYu7/K7wBfNn7yjmS5mC13A2usSM6Cn
PW/aOAwqg8KWEFQI79LOARmCs+20mCWMVccjM9DszBDIeLUQdUo7aiOQadGnlyACYDq6kWcVUBmI
x3QMKek9FQBgT85BoukRGa6xhKGvJODa2W6Uf/O9JaeySsL5uNEEQP7llXp3ScFcGN7v7wOEJsif
3KEXxtPj6sJt+JO95wZkzJ4R2QcfEzijlJmN4NCgh/TxVhpYUcp0y+qQMmr2eiLgB1kEY+dvbE2i
By/ByEYzNUgr6P3EL0iev1Co1ApyH7EcHxiaPnxE8N6dq+jXvNGP+Ot6BMEOiZxE9boyhvi9d1tJ
ACIh1BmfjICI9dhdGqSisnhxWYkKYccLweyyROYrXtWgq11IrYHH0qlErQw1975BoLdIxJzqcKDw
K4TrqZVzbgIAH2jKnIaKPpjwn1qY9UXbE6jGxDhAFTEZrcWnH2xx8qPg2s++71s8UltGrZiI23yc
GFGzTlIYXsd0wYtz+1/OoxKIY0qq4PlLBghyL5zgfZAig/ReHjrEuJIcF0bI+W4K9S8e1NspBjQn
/Ry0ZAnRhZNApr0KF8hBzK3RiQ6kXMMM39p+4pjp+EMfbz/OwIsTvSVU4RxLPk8hm4Hx4raCLlqp
Vgs1EiMVFWETCs2LKFE5nid6t1yuEpUn3zkPoqhYI8TZ0kFTmosmPcNCvHeK0iweiGQTMvG84z16
ZzXsjlADrUyxIi9F/IswUirzNAam7lzB/eO+FVpGy2ag71HmfNwDJMMrA20A3JBRLMj+R3HFmtCu
AI1UGLSK1Yl6h0wZ/mqIy7549JnmBXkvWglm5O4M+WPCaylVGfFn5W8TLWqdKyhQsew2agZn9Llp
x4cGAxg382GRt88YTNlHRm0fSG5DSb6k45frzadn83DMVb79YkpJ7WsuhEDubY7RCnqnUm1zAvdH
iimI2uBZxijU6rvOBu7GRNt5HJh5AmKD9+7Aa62FIx+ZYLjghuXacQg+0BvFEcuQM2tY/6ooBkBC
1jfhqrhVTWPJYcUfqLvfYBorSWbqks7UoATy/yIvIKZdsUz/OI40guqN1/ttH5TR07he1EqpfO4f
M+ejdxnHZqFySXaPpcprqJpgMjI39ID+lRu7aZKC6fKHX8IhjtlGoy1kGlV5zBFz+cJV6uDsE7h6
JkVpvnTK9puAF9M2E7ikxrrXaNB/3E7KC36O+w1kG1QBTUajFT8AP/FGggUOkFKZzWLhkw9aNSim
dsnhfr7wFDaO4/OBXIfnt6UC9+J3qGroQBZIanLZUA5ILvNjFlGO4GjHTyp+5FwNUKQ19gvwJJEU
risWlJZJWLfAy0zBdbkQ2gJLkG2yHLF/JA8z8OH17v1SnEIeg7wPJk8muZc3lsloawzy5g8oJ4Ia
TBCUW5IS3g9lTsoP90eIGRnQKucfVBUw6v/JJD5rlfbAPzH28mM2qzg2Wv9X//daS/yB7yRgQTEZ
iDvSAzx3jztsW0H1qYOYanRp1jmnMNHlYOyY5TnPeCEzrAj6bnoWneOK+H1KnOHuxA8SUGkLwvg2
9pA5V4WOd8punTLEd/IAG+o5OtI/iVxMA9Z9kdGBqY34yZQ2gJbUBk7xHx5ZVGOJViClKLzoyR1h
pWwZCntDmoutgOpqr9KwIDudjhXYGZCXC2kBpwNYWvAhsCNUR2Jzp9AnBcngS2UByzsdOb7eY6pd
3nGsZkO0UaDJe0K3E/HtyzlMoffKZgCFNArcaOkywwlWJB5ClQLs9LFpVWUE+AzxZnk3M8xmro6+
UoL9Cmz9htdCurtujr+V9VqDcB59H+KlwTsyNzHlubfm7k6uLBbUweIhzObLxNVrKqBzdss1JNDk
5LQp4Stg10lNorqTUJF9PBI1sJXNdsUx5GZ25+ggjDseCaiarIEpFmdoMm8H94tSV6uaFuG9c1Lk
80JNLREWy8hHp20e7HhfB1nwgV0Y5D3o6sXxQ0pj4A2hkyVDeBEiMECAS/cHy5XXh7aG3lxo15oQ
7JccpvxbTOlUm7YV7dYAs0NZxASd6qZErArkRBjvApc3lrO61tbKukTv094XIyyoChY/Dl9Lr/Ka
uH7/hXseiLTakt6+T75C8cuI1i9L3cgWgrGIylOCIf8vmVSVZhmFBIhT/rpNcWvjSu88SXuxsdd8
8ZZElCYq+ihCogZ8wZbpM24P1Y4exUeDdn4yEcQ92gAYPtwsrqbfu6ikswO4InCIkpkVCdopsSm1
FUKBMseTZ52FmgdwNRcTFHx818WZotq09gvlQOyrrsLUKBHdLHS4wryg7P++dn7jIST5QM4/jpLH
WaTw85dfQrozY1MIwbFKxhYfFPR1HVyoV5DijQFsGq4yGfdVWFzSM40cds4/yZcHjSX6Eaqg3Hzk
efEUXX7ovW8BnjHjuRMRbz7CTyE9Ng9sPkXi4xvEw3TD3i5i6FXSEZlyfYZSnyBEIczQtIHZJdjZ
JUudhMFKvgiqZU6A/8Uwd8AFUQ3XJG8MluCZrdihdHlHaG/0zfqd+PneZ1ynMpH/FGI2aXj9sc0v
8NfTcE6z76laf6/J31iAqSKwUBOlgbxu1HwsyEtqDLoSDSwA0n1a8HyMDZTaZ7i7xTU/U6Aec6s8
CFFgFCzgaCvbL/VbGlCaXKfqweHN5hpQJWOCXNwPXtcVxLcQuMQjbXKIZpwhXT5vnvkia9JRQwOx
gAAC5kGu1i+COrpDz6wN28AbBQ6+ckEDWSOT6iz4qTBFt4R8e0PSzzWLC49nG7o7nct+Xvv9H3s7
JqZvJFR1EzT4gd/3a7ykCEpFlvYcxsuzGigvzWIwiST85eXJz1QJ4jaCFCAmdEbNR1TWFUTdxtU0
JDTcmU3cTw6NutJUseQlbdNHhAXw8EFx4OjPIiERdB7R1GHQqvKIV6OJKAYlIdA4uig6dmi6RKK4
g4LSzzaSGbj+L1RlMg2LcMEYpnaPzpIz92V0ki2D+JrXumK8YYYxS3AOfELZCgWZpX/ZGhPILR0S
zwn4B4mnNeM+OAbNFcVI7ep0nwsjHffrl9ucKgNxopy0wbGWSNeE80g2sgPoM/s9NkuebrupeOKt
efykOoHqWwGp1Vcvs562YkB/xQFxsmAZTfH6BPXVHtmq0iRgAhR/RpqjJu+WKSGL9ScY83kip6EW
2a1DKwt8irCR0qXIy1djqZ9VPQOvXJ1PjUyKZHFPZNgjfjp/ePIEV7n7tDKM7fl0bIbqZhIrCWgq
SWnuhLcuscS2ak/BzrsOBwm0V3tJdD8z2qWbkw3Smielnee9KMGGGj75oL3u/Namyt3fUKN62RC1
U7lakeZrJ93AkNpDtfiEQ9XBpw0Bz5hU65RT2QI5oySlh+zzCB95iKfikyw775pN0lXDi+OmjXOU
v2j46dpG0z6kYB0l1iHXsmEIhdjCM64hzVcBTB6II/sVMbj9GWUfPRejUpS/3kXHDIPvIn9POf8O
1e5GDJGh8Y0IMoggbUcQttPHMk50bmgI9BM0xvQwgVIrX9yPdHwifWEk5J5SWtIPozyhvrDxsTBl
Aq9raVl8ZNJVcu8qRAqBf5N569k0jVpRdmwPkhRDQ88BrbtvHbE8y2bLrL4httzK8OBiIl2YvZJD
s+eeuy6mnuuQObejMWRoAxmL+3aBryZPyzjazH3mCJ6yKwsBeqgtGg+8ZVOp7bXxZh/ee2PDnEFh
FAOZTPMon+SxQnTfxy4rSO81KgG0l3WAodsKLXIPg9VbLm8U4GXjAwqjSFlL53I7hS4/lMEIGD5w
34ADc2Pp8olHhPgmZOhlLxos5EoqnnngnGs3pf8i7WdeDUgIlON3EJI3Gc0zBqQ9uCMTDpWhvqlu
lswD115DplLiO/GShN9Qb6r8MAsUBN+63Bnz0ob4iX5OxPD9CcQaVaD2k4ImqRvQNbQPbXB5eX2D
Q71SGAujCptoh/QniBf2qEFvekGyKeVdCRhKltfYx2gHlmR5zHxAAkp96/Ppq4kjpHG4UZpp834A
V9aE4ijdX+ilc5888LJGLc9zJqWPpMk+yRa0v4YVh4NVL06rp0x41lYUc9g65A6SO7PVRn5K2NXt
Amo3nYilEFwnVVs0EwzGc0PFR9dIg7JQiDbDalBAGTkrDOpYBYPbg/JhUwSRx4ashyov52KbEoDV
JpV9N/7fU6dBUZjZA/eDab+8CoEvuYbEK2KStSR+l0et0JICd61JYcHbolAA4SM0fTrYLxQQk2pT
/UVWvHHOA2LSzsnQjNP282zqmzaBNqTQ9/Uvsu5T9Y0jBXfWDXcJyhhJ7yKRUhVYnaDCTCrdshEc
PGmHBqiT02ESiYvY/yP4e9amRIGFMF7DORgQ9WksU4VWIGMLkw947R7X1lTIK+znm7L10d+pvT7e
wQbFADOF966HRgcxBQECH8ckfDPMS8tqykY90U2Q0e/AyAPx+/W+ZEt9GWTvDeNdU5ze1fv8PsTb
D/4b/B3wWFvaHP9YDpiUplWE1q8r7QihArzHxUG376MlUVB91R2R8SRR0JdhrwhU3zlCnfJTkGhF
tRDD9H2RfjAYH9H2STQinMfgTMhhmxehNx+YhmSgQS9ExgUZhxO+1EYUEO+ByMGYUG0v8/TIVtKt
XiW/o5Gr7RanH2JFt5QeQtlP2haPx6tC8WN8LAOn3/Y93tFDCAEgvxN6Zl2AT5qrIN3AAC9Zi7aB
BTQWY9miuLsQ7sPhtemosPYHIesDPhzyTd54rSgYi0yypNdMqTSvDWzZkKr1/GUtxBIiiVk76v1w
80qqrLviroszJhExo0kODOzVX0q4NZsPeECX/kreRSVGAxX6pWcQK2WUXPcdg3yqUeXWOHdplko+
P4WZiDFajaTC52IDITuAGm9zKoqtzl8dDCDqjANPVeBc2GZqqlXA+cqP1EccXpH6m8yhA5VZH3zo
SRiYUSIfmDPQmFawR7J/c++k/C85LSCJYnb3jAVyRyg84HrPBbAAM2nsEDJ7CBogeBLdWFEAxvKe
DnT6PJwYOHbgdur/XnK7LngQrsr08OINlqYqJOhmcNmbqLg5FRLM5rMwm1i6uDvP+zv3C3ck4p45
iEgXPom6EHhRrr2GVZzS+y81gAgQIw8RBTY7FSnxL+LAMpJyN37MzpnzOkiaszf9P2JDlh7IeF3c
2nw+ZvYowQ/43cEfY17DW4/k8ePNIJFXCY6hFq7kOayoIvzuLfQh/5ewt41GuA74d5ylEUnkLBjo
/nI7d28BL2DK3HqLoix1ZwJ6+cM0tCJg6sr/3pp85yPyOYlS7/3KFYbNTgA0KgQbkZAXnxFrDd+Z
0hSvNosxR7S9edNb/ZG88zMReaks8mO3B+jV8/wqB9gyX/oTM9c0NM72sZueshVRb8pkfIiHqEY4
l9GHNZyzA6WIKT0ZCKwjoWJU7EbB5pilx4P2HScN3T/1VvSZTwfawryXtzzgP+6X8fbcLdqBCVG8
jPsDM7dWrOwyl3vu3pMV3lljvUx5zbfjJG0H9/9wGx9DQCRXYkSc4ex9e6x1WRk1oJBukllaThgL
7/1xUZ3KbRxQK8PRi1D6ulYvDJDoYEI3sSQhGFkkFs+7k66o+JEdvuu6lPrItejUtQ/8otQI5gjw
dKGu60daMl6Q8ks02xoHVY/+/ImrCegc1nO2j+NobEWWi3+80HqG4Pm6AaK9qUHTLF/jrToQwUhq
AQUMK4DyxfD91DoAF3zUt4S2ZNOzLsoCkoCQxM1H8tS/sftp24BSR9zfoJyR9vB7vIyUTLlTlhSN
fC+qfLmyhDZe9VUMtIArFX31MzR34f5fFTFN/lRv+k9zOrgnsz5aAGqApOGAmcKvsThXKgvUakP2
0L3jkHJhHMg/gI6JuTUbGdbvPyJh/FA9dYlzOFKg+Sbv+z8ytCpN/dn/APE2CSutrViVFz78LiZj
SAFgrN+o60jD1HeTYAFWKYgj0Xv+l8SH9yMlEOR2YUIkj39un4/N9/CPGXKLqUUXOcFJB7q4LcG7
TkWHuQBALYsXbGZ047tuCFQu1AvrBapfnA/7V6G7Gp3/aIjAEbrbrB+vVF4EwhUb40LkXO52QXUX
jCYPMJL/hI60FLLCOJKwxr62uwZqgIwMs0YQoa40rscGZoDSYCEv0OYbcQt9jEg+d2Q76/N8TeKU
XI7v987wcJLnmEC13XnoNZFyiWVopeNpTcFUfR0TeZnkYYjbLJKR5xqApb2IXROknycIkaz9xGLW
9PNPcohbP1UBaaxlpzgMIu9D8Gm6mjvVnWfog/TpRc7yNykO6yXqlrYADwt5jtPeM/QfRTjHA5Cb
Mrq43vQJdHzB7xzs6pCgt08RUv8ISa6AC2u8EmTCluAbsYZlPzkPl/O8aWOo2ti0ziTaLqlRD1mJ
BVtyi+6gYME924g0mHNy17wcID0ONLBqvJsQhv0Cn3cD4j5FneZbAMgMSjKgf9giDKo21jT/ThZ6
c+Jj+uEwRyByiAHxqpSls9sLHPvgnJrVn5Nx3f4/xGJJ3mBG1VwjYwtPz6GH87sJPFuD5kdjz7l2
LgyKgaNQM37yfapA7ria/R31itqbIWuTYsw6u8hDnG7YE7/XT/+UP+XoIgEFE382qlhzt8oNtgmX
T798lR4NqR6l2U6GwWjPH5LPKn2BZnrqE7gg6wDTEebf+x1+so46WmNUO4sWM35mL9UD+ZnNPdfo
kNmawLBB2C2q+epyUcE4/KIreak2r/ZeyMR5Hy27pD9JCnNboXGjxdnoOeqVQ9rq9qJ8t9kCJPgs
RwfdZ+jtkyqnP40ZWvXSIo7Ofl9ZmTIOvqVC8kz/TYzKaUf+O+N0mUVcYBYsCuiCpqdjt9hnUSz7
mA9W2n+7Au9gQdb8fsUW5JPDjE1SYreCElKc3kDRRcaF6NYvFPWafy3R8p021nCRrbqwO74aICgk
8EBn71d3DfKPlmFW8QvWrhmesZgKY3ifwwp9Z4KOwjJoPxoUPqgtHXdu8t6h1ZCquw6WGXYkl2fT
03sPs9JyKNdKHa+UV/pAvnz+lTlmO4ZRwkgi4iG9hXVdpmUnCqPJoVplMWBaAboTZb9msK1LRIDB
73qeDIR71jd8WimmTni5byf14UqZ4Pb2VuayeAIYkRaX5fhwEo9P7ZJTInT5gJZwiTh5jqq3HRkS
jTuKUd9Xs+VNC4tdKl2LkQcYKePsSrsle5XzIgXDZhnV5aAa3/HyQIdXmR49TIUmv62YAMZzGWNg
wrLz6JNhfkTOZxQuQGeq8QQVm/iMjgWP6iBle8X8/Xj3rP9pYKBAmlfc7Y25nASBwg4nFrvOd1HV
zV6HqdT6Mk7Pv1gSQ/PTgFbF+GxcpdE5ZgXsitMyBtYpQruKzCej6uRz9XNSqKoe8NmqJBoJmYCl
Bj9ya/Pbk1SRd1n+vISpsiZ4XXqXLtT4oGE3O9R6OoU9oFIx0bxfJrnZqORfwiN4Zz6DrRLdH1aw
SEaxTd09yd/MMmz6EtkEihzQWnbIXt/ZBmodYRtSl8S4OaczKL5wGowFPR87qvpDs/f9+1HRR++Y
OWAx7ZQYLEW6wESAsNLiJz2qyIjMMFl/I0dV5FWaEs1XpQobnatPqIzXNWh/SKkqrW3DmDZ+MaqV
uGSiX89ctx5B5umQwFw5hOIvFkMYb4iRPusE1JPKBPwvl1NKXbyBxZUI8nmw8HU5LDJx8ZFJWEuu
V2CdDG+LpZ+2EhIyhDRJ8OeoBM0hTZ1/e8JDIfhGfdlY8e3i0OuzsavcgGSKphDbGlkQyIT2iGKF
DVypKHw6n5iRmsfuOy5FJApJHnpMR1EwDMxOTtCFeGOPjGvVQ3NxE4RJFmZheYtpfBXNvp7sxSFn
TvevIOcmc+g/MVM6VIXVri6obcoNePLj/joLu1Gd3N3W9sKhVq/uhXt/gQZa5sQyt9Yizao0idPv
S3C/y9jY6FEbM30Y24oCcLreiBOZQf4a/9aiC/BmIqgDGIRPFXjKlM658Qcc1w47JFEPM7AYMh/8
mkFZQfLkkSg9ysBYJjd+FZW8pNDpj4k6CX+wzrVgljc951fyyy//bU8eKvQOHETBG6OWbXXZtDoj
yuXRl8jjKabA5K5uEF0lfL3gjJKv7XTvduUGyVyeJASCXBB0gWIcL+v+SgwkRSAUNNLL74SvI7mc
1jwlLVw2FmFo7orMYIclJfIZH52dNu1rID0+dXVsFDQ63RYUbAgz51s2KFHnk2jwfW0XQV4c63vj
HM75xeosMFrOJDAlAgbsaEm8J+7GCCYqbbsVJ1iBhMEqn7lcGJ30Fc8RkfXVj/ALXF+S7QIwHRx6
wxdzfeRzaFNGE2Xqs6LSVGmJ/fyI6i1+2erhntafgpkQcXM4U2DPCusHrNWFf1dFJxRjRbbrtoNf
MDbsjmSTPBCjQI27E6e8FfFC/RIMiEnKRa2N2aTGn+USXOfqi3WOPnACqxp92uyHFC7IMlZK+NfN
FTIQJl3X6ALgj5KsX2+Z+1VWL9UrJ3OaMtIdi8ZkCjHPgacFEDI5H6kiBXWmBnyxTrFDy+T2jkGS
13rzJnSBkDv/EQkOq80b+V4lVz1fNhdrPQRzis7w85qskrcX8rrWfWqHlIm3dJywXVEs+EzsAer9
DdegCKoHIA0GjWs4o6khYlkT+zA0SiVmBqW/lendJ3S9U8Cu2NI1VT6mE7zlLaU8If3umIvaJZAE
HOzTjsiqqvNu5RxVJJphPWdbdgs7c305H8mJhppitj8X6xFUfIzutbiWkSLk7G79CND0R2pO4WcY
o9+g0cquP8r/G5NjAt2bix58R3uvNcaMV4XC/mPU6TBMEiRN1mja4Vhd9Yrn+6yYVjpDrNu3s2+W
iBwLZ8pViDGs2GGfHLrQa23GuCGM0A8xfFo3jYvZMysLKuLHceLbS+gIzFj07lygCG/z56xzyY35
NozqNQk819LAKT61hdggj/UtRQMIw3OXXj3Zp6qevU6S9ZTXw9EbQeFXUnNdMc5su6d5onUqoFaL
mjstN9Qt7R+NRoAPw90RjzJOw36rOshNRjH5kvTYGo85vMDTk2uO6UaNkxtmoe638w5o3Nagq20y
SJwe9Ez2yWR84cn/JB0xv/7/9biTTdvm/O2T4EVhQe4OCpzeh2zpOqxgcZ3XWxZ4JBSYq1GosaJR
XM6p0efqO67e5PBMxlMi9/dYZU5mFrECt3TSIXgchTLYZpcaESB5wPcXGzFKRpQceZhfbZ8xKmSH
z0oo2QSt9kp5JypduPE0QSHG6mhwHa1nxcMQHr6lCGJyJfJHaYk3tlE6Q5cZso1iOU7wIAQbufKj
rxnWir8bqE5MRqqGyvEBfFnmQKNsTSsaiBRliP5smuTyWDaa0MQHjGmR/hcWreCaBikeEDjtpHyc
rzLIn//f6sL3t3VayZl1eJad9le8g6xUhjVKkx0eyyV89/JNETgjkVvgfeK3PC1/zr1ULih5OpPp
Q0HHkpjRGDh6WptyWL7fTlwaOFPUY8LCmeyqWyvjDE0N3B/+XBdeb6Q6UDNvgBfJp4mWQmLiUHaj
z66e4G70biuuhEvxU+QdFB+rvUHS4bLQNGQx8259cCpHxJS6J8XcWp9UJHvOpn+hQT9wz9B4/Po6
uU/6KkpTT1ZYjsRuR4Curd3P/NIRni4Fnr8GQPcN8J2sVdoMu/oWU1TE7Xeq9vKVrgU1y2bAnL0k
8kHx6DozCxfpLpCvyk9TaRcu7tLildwo/G6G7obxDLXTPD8jTBwDj7ej/jozSNcMDPrmE8PTK5LL
IDuJWj7Xgb1BLghbtQpuPakEY/9f6xaiYsQlnDq4z1iuX4OGrOEaulbsn21qjiRiDpiihTBo6BQw
WqvFUgT2DnWMx2QYk3WfAjMYWeZY2jOXx752Fun7ALrNKaUOkz8zHM1Khe9uHh8O0FBhWkzUOss0
a7hMozzmaHqzA9ZfXTFVDpMzyEEXUc8DmhJ70QNEjSZr50ZtaFDW2y015/eZ5kpev/48xQwrENa4
ywwuuAMmaOh0c5Q2rIhtLwF4R0xTzO2JQ2zRIzS43kk3bWi7uTi8Aq7oWjP/JMedZ0cR4QfE5K98
I8DSAXbt+K1Y03m4mfR+Dok0MnCZnOeN4zR0ohyPLWEJtTcFcjCDokT1hfEvnPwt2B/h5zMZi5uv
OO+Pw9Z9L78JAtC+W20yWccXOEXQujQFjRBUQoOqFd+zZFHemoS5Ap3wHeu4yaSfL9MH3TR6Rbsg
8na5rWEiGqnYXPVt+uol7vQoBZn8VLkq5pzV/6ZWzizuFbdBCyKRHXvzEPlHFabOWR+TTQYl7NKy
7lsMpkzmvhBrCZDbQoouRXQSXb+uwAqCcxMZAr4XcmaTc7ParkKRyFkx2xzQ5hHl9e+2AVLPU8t8
Vt2SwheAdfE26KDowEMCyg9Y0cLfmAHjeoT8fEXHGKp6r7H2AyNu28dBg6TE3Xri/ZAGPGnSjJjI
NJMP/TTtF0oSaC6LOMHLLZgPQ/b23F15WYIM9FDsyP5OD39ItEw8Tq/UYPtUrHhUPvhzGSd6T4yo
Os56zeRL4rCK36g+YjAWCzgsywRWB/1/eSPYFrkZgWQh3ddz22llA3amMlL0DEtP3HcacviafZ+X
Oze+oVL/yE+63N9TpQLtcWOjxFlPcHAfdsm9b0SnLHwzO91DhsZQIWG6cKF3j+JioCxdHCDHMScw
1e/8LWNGS2TYISJRTwG8Asve5IiXgrtdqzflUgaaJoJT2LYNfkJtr3oYc3OCTs/I/UkALFhVsske
hhCTi8Huo8C/G9gBcKCMJumafyqJ3KxlTHeRKKSxtgu0EpMYQHpSotA/owkQcieiYJj0+zKojDJk
N6iDcJhoMDGn6C/mzhY1Lc5BGpt29oHOQO+fRdydI+hJlwgIVCKxT/PHYfOvLccxjmUeNhXgLhT4
CdnfvFYzFyqWe6qInxq2SEVWFl46G7+gqZ1K8stlljC2lagXZie9ZAf6yNhO+sQgmHk6e/moP4hS
vSu1/aT7EN2Wjh0oGSXwFgPnlSCE3SUeDbiaXedKTNgu2i1OhXyvPg9PSNaLCQ/hcAJdFaNyu+FL
rO92s/vQqCR+ZvvU9AmfWP3HTV8QT0/jXqJYg6GUM3+Y0Aa8mva/M1oIhm7bnwX8y17aGRJwW48T
LyIIdEE95xHkjlFPvtUPVOYKtPiUFj1MZYPWaUaWiQgn7IXwzXQ1yn8DKGyfsIrhy41aE0hVIAy2
G7Gonduy83MBZEzXfXNznf5PgOg8zWBkQksqm32YwYHy80kcOt4O+2ADnTjPzjp49PKhP+eo/ZuF
vIhbFUrcDnfb6/dfj5uUEHoCux5ETziOdnTbtgpCMa8tr9DfAEhOSFNFfrdlyWnuCSXXhAlb93pM
sxbg57GBgN/Gm2WcLOVazmtcgcJPBoAzAENWwrpGnPMqaIp+kQDwjOMlwyasD7xLHuDnxFleMWV0
r3XZhMKwsdvublRL22MmtksGOaQHRfBxpMPwNX3L8kD4ToCIfdgv5BeRAX7Wa8qEO0KjuTInCPO6
mFlt66e0zJutnh18lNr7pHklHCS9O0czaF3V4m3D9dyM3HRNkdKr9pyCo5bWyG7chzJAKqorR1Af
SSSh7WTmegRYq7Rpk4ApVLIxnno+o5jcos/uKJnR2oY3yFgaL/EPVMEpnG1csqbYUjPmt+XUFtyh
qYeX/arT0AXlx0U8SVNhGFEg0H5ac3CQ9NgdTErIkdQT5BPyhQRh3w+MNUFATeeeV5gbgROdvqcC
alyjUo+uK7l8xKwyY+CVUBrsFfG0EEpYDg3TLo3+BOQJTCSmfXAlCA+WuDgrAIzpFgNu9FWE3QbZ
gSismL4WgNFNogP02c7SMH6AEqb11Zws8fVl/ckTbCbNJmKXxBaxuJ3EszK0P0XQpsT2XModnVZJ
fbHpA5jOmD3qFJ6ZZ5Y/HDXkpvieQ+G4kf5apyEhVZh/7MlfKgnLKzrc54Tl7tQRlhhZg2HXQxtw
m4UDOjOLUXb8CMS7LbyOGmNqsoqKsAs+VDP2z9lu0uzltOtPH26hTYxd5LKzvP+hK67tZDTzDlej
vguNDdvIhgfHaRo4IC2P8FWDntmzDmipGi9HH0lB1FkChBMYTevS0MWo43xQQQFwVtya85NcrVrn
fNyUonQovvrcNDepbxyicuYl8FwV8wPVxk/6jPHkcaxv5n36nLzkSDwoO4pthcXeXytlNToJndOs
2R3+q6ijSD8n2mdvMY31A3nLM+dGtYDz33NyxTFJnoqoONlzkOvcpS6cCmv3C4gpMdsy/Y4rSdIC
cfvNkHWWdicKpsi85eoOm0GqR+Xxj6Lgpf4t7kdd8TS12fwcP1ytRACeez5H+C0KKBTGZecvtYQE
9emoPyePbYR6b9vi26CPj5dKmHWk+y5I2f1AnEZSiI/LqxZPa7nvSqjZqyPwE70vKbeGiQAiObNj
cZkvt9vr7J38ERtF9FRaBTG8zj1wPng5wT4ebTX5O2KXbOKeojADKta3Mw9nDfOKEcNizz/nWXhe
KYN6gSNscSYavLHFQ/gzQuNXWABFVNOl/V/g4PRieVgrnWnjmO1MF34q1FfsrNItzDkNrG+DFmX8
C+b5QTzi3y1e4mGQrm0haVi69VbEYHgFl6lvfyDkMlcr1aUDuwVhr5Oid+f1OOahpTaD18gb3fO6
C54tKNeuNzwJ8EusuDBMhtvQEtQRO8AogpwSsnkAmg/aBDH3xdSoHaJN3SsjqSnWi6G0ufVQUbB6
hFWu6ahU5P/zxxD+jg5d6k+BCyxEVi1EpnbAdS4K6rFw8cjNsBNdf4yFqA7l1GA1zXjMa6Yx0q/W
pHCQuSOdkxicSaDBcN14WFIS7QXm8ZGy5hpGoht/Fm5KzWQ9YLrNXR80y9VXExZo160xl9Ogdc8s
RyqsknA4ZgHFH56kcUQ/Ocy5AZg41hi0GCwUYP9OVnTTgjQKrVyG6MPey5QCBujdTg5rwueWO0nc
ahvAgGJ/51F+Y2kIrtLQLEKFJTG3D9tdRrNrk0b/LJoF3cJIIBxAVR+gv4YnDg9ATFX9TiTJDWpT
EyY3FMmw8glYjZK+oLbWAU6gSA2ySj1oE8lqyF6fboZ4fVzy+WXDYIOsMKeifR19/W8ZPcZOrNkt
5SoywzcvgI29g7MmVJbb+hAWvlxg5OxS9A+5g66ej3ld/Ytqbkbr0KHWfwkS0xDl17WbfOPMbb+S
nYoenngcXco/YGd1lGqHHNjs7sl0dQzxPbBZyD0PUXznxJKCQqxKIFWHVtdvG+PqC2nVAFP9W4SV
L0uB6xYkFvdpxOXBIRsCVNz5yeddFGu84UVKKPIsoM3BXNpVUk9JUMBVhe6YN8Bz5t//CCt+bUoC
nAEDBpd4JgTtx4ILiJEqXuybKHTcpl850iPEemktxCkE1nc4bEpVSGrv8E94XMraY+w59HUsM2Sl
NGB1unbby5HrLgs8qqyYwDJ3OgVdG59Yzyy0MleoOahRC2Y9O48VodqmWomxDoBvXl8fAfDgGG7c
FrmHCTlEZssndIpjq/OWcYorxrxWDK74aAJbkuLkhdlmLtRhtWhcFZA55eHFQAMRsRZP523XmrAg
NYBCdz5saamLWV8Usx1B4QMi3vFi8YsOfXck+IuCoS18YDzO/Fb798SwubjpmWFzfsqyHj7akSV6
hiVlJNApgExsjI2gXPs3vaNiz2iYCzqtb9Ivpb8BXx42qXXc+LnThmeR0H3PGGvsuzMRZmZZgTI9
cgAkEAmvnGDXVmLs6HQhB6kdpfsjUvbeW6H1NH1nflA00NXmo4lUKe2Whw5TOpHTQTAMuoSQu393
+zMak7YKcHxUqMAbSQB229APxGx/mvFLtw2UzQKErZJTSJfP0/2wA13gI2F2mrWN7rIoMtjDXlvJ
Fj8azw/MDo4y+vXjOBr0gEAlVx12ySj/rfYUQwzB5+8k4BgQI+qW0hHX9U/gySrYqO2eYFAltYRl
vng7j0BGbI7UhpP/7jbmAHNGxZmJjI2pK2yJsD7mcniIeW0vt7AnqLGYwveeIuPDVRd9qRQv/Irq
yfPXWFDeDfUgaQ7UzcckFhJRm4Ov+dL7xN/ekX3RSw/4AMdrHOqL9OiHO94HmFJziHXP+dOIZUww
xXQFLYjBJb+NiHeGS5WEZLR/4aicnB2Zgv+7FhmZmhtQnt84ztgwUvIA/fs2C9ZmOR47UtLut0a/
5S9I0HxGVAiAeYfOM9ERpGYjI71lTuK17uejJ/3s8j5F5nBJ3EasspGeGRPjINaQztxt+/5rEu4e
ZeiwqDnkCDaYapxPa9jYR0YCA6AER21f6EizArpHlyOVnQDu2RgaOSxqEN7jlok5YcW9U9Ccd9ts
xV3ZIcJGyKEMG+LnaK4PNSD1sDj4lkvopQig6vEVqgrhhevAyd7H7x3MTgBrTgLp/HJcfODdRNGZ
XkCQHTALSAD/rgQrj2c6OwYJXNf/hyho8gjCQZ3TG/NYhjlfR8L/TlLBfzTsXPGMU4XYiOVefV4B
NGX78tIF+oLntNpLCHglfI4OKhtSnDeObg+1zvM8H+CVXG+XGxtpoRIoxmUcZd7eD3GbHHhMTkE3
yFbSaj8CHIFtl6PLNXhgKiNSilSNfcmqKEttTlGu5wqmD7mQ1yhT2/ifsMyDmw88VdR6XfGmEnRb
+J4DKSV6Vf0SIXMssRXC9P1E3p3sy6sVCtj0mJ4OAZIbHwrljWQUs3lo1zUFpB70QFfI8wx4FbGi
VjrKxmRdMXzJ6y6a9wbMDM3beZg4CP7h79QCFMdQFZ+qBUV4+JP3h7KVOU6mqRo9ebxO9km/Szd1
b978sWeRKfVJ8byuyT36Ad4jDXGYueJsqD1+6iYV23Gstwwv/KwvpK20nARRC6Ew3EDusyx4jSvW
xX8zkFUdBYg1wElzhBTt7MCTKp6wk4oIKh/pJdwx5tjHMAlNgoEY3s+QOsOF7xJKM+Hc4IufGAR6
UAiD2YW0q1Mw9o8l+ZfHtURz44vNVsYwRCU4v+TTzq8smoeP6VEuO+MEqIxwLC7Jc0KFL6py5cqD
lAschkLR7+jM0yjRtK0bIYpwbmSm/XX5yflVxGAgFvU6hIuOScHSVRlEWNv6O/x9tOFjVvTERV2Y
OJm4XOtrQVGysJa7GHsfCITgZFjyWUSyYX188XmMQBKj2QtC9kjMhDL4EG6u6NTsOBBjjhwweHzD
UjOBdsMRbaoJCOZSvJ8alwQuGSSsenB/sNGDkNaZW2zxJrvkf026cJ3epCUbW5wE9ZuEUj+oj7Fv
Y0/e3Czc2vsU5j9BnQzeLqfF9/z5VKM0ZBaFNYxlOclTQZLl6JlJJoRjhyRBnOg9aq/a1iVV7+Jk
zV1F1mLZGU98fyWwa3D7GBUkba0XaX+9y4/QYqOirZejbsvaDwrZm30L9ZdRHwf4jtZ8IdnBxrhI
XCh75MuO8h2Y2aJZvPYGNnCIDJDsPiMngtlD6nfIgnwJJRWML12sWvBP2VYc4aoy4cybfPDBzZyu
4WLp4YSqYr90FpYOfbZ8E4s8RkmuxMWq31QQ+ig9FbChvtVDfI4V4QTpvna/XLqUjyE1VCNb2yoV
LY8ce4/nt8tl1GtNivv317Gyxki2M7k9Mqw6Kq/t/QHQeiRWRbjimq50F2KSMVrEiLS9cinUrSHT
6NuSMYDRuoVp+0g7Q0po9hlRiM1mS/1ECsxT9aMN3NGjnDlU05V9aWW8l5HAcjzyu/ohngMQnSot
HJeCa/WtsUjqfzjwiXKhpYt9I42VGS4QPbqmfpJ+p8p3vIbh8dAF3rYF1GeDKwo8Z3cWbOyzKrAx
ZFpnExSUIPtzJxFV016U1yaJ6WD0lC4uDtB2Tg42V/zluI2+fQvHG09SfPMuQx7AUTd5flgMiaw3
B2WiksGfTK0mdLqHem0G8Gjj5f+romwj8lgmFaWK3gGHp3tDNSbt5LgrlfaiLz9OoRl5ZTjvYYRi
25KQuF0Q7DnDszgfnJMdByLt/XUpv5lqJNl+ptGXB/amtZOLvjizPvCwCrhMbNtqfwMW5tNAixn2
RAfOPDroPdOVUXVcUbrXojCO9a/u8EcIKJWge4jqArZd4RFQGvf6kRphxqMPI3RYHLbZ0O5IWOf6
146cgzJS/5oCbqq6w9eabkH+/7/TCvvCzsdsdnV6kpfvBbfKnj7j2b1W4Od2oD9b9BzrYsf4+YkD
nD0RfVk0RolTzCRxZpZ3ozqwJQue1BKnLKwdWmCyI+a7kByH+ZTWKeIexGPhVSC9ECaSFRl8JezM
sjQgUncUeDsErJztsRooSkva0iRLV2xeehUvgwFBiuk/+i4XBfPKuBTLcosVuzG7RG45Gimye46z
AuiIN/AYW304hLZ3LeWEBnJR1wDhuhQMXo888zfirwcXFWAiB6YZpG0YwHn+UIGBoeaIF4hbMxZk
27L8HyjfrwtsekevHtFOzngDedfV1NQi5ydrRsyem+TSk/57p5qTbShOoWmk38Vw4mxNCS0IFhux
/Sdj4cB7i0iagQA0YLx+Q22UFJ7881rP72g+UGl2McvXRk5G0Bm/3P8wErL7cW5XTsdDlbttqoX7
SYhnD71G2RWERol0gR5Q3zc6UZhsSAMBZCx9FIjRVf/iIEjamhNUM9atoKTvQEEl0KcKB7SJ3MYp
xS6WTHaElwRkaVHvhPCySA0jrZ+eAwUweRtLTgVIWbQqfSqa4XwQ/Ily7y6tQhNeWW1BuP6/HTvk
NoKS2wyMRz8Yimjh5MZNVooYBw8X5hwo1z4c9LoncwrXYeoQE2Q/95Oi8z0KJ/nrbpRgDGp/FvM/
7C2QAkJbpA53fM4Ptf+O8UM5dwxhA8PzHSPF6q8ZjV092wwGmm/9Hjnm5m35+gycKfpRzlpjhZ7b
14bDHiQj+ht2mxs9/sh52ho97HbByE8yYx/vCPZMSqMtAEI2RuEKFmYvkrZ4ME5GCM3wJJi3ItWK
PUTl/xra47NBzx4uVFj3O/UGPYbe7/Q5NW7ujkOXMVdp+et6VYRE0VtakW9/k1570MvR9JFsa2js
/WdUyJd41nQ1bcenMIkg3ZwWqpH2kHGbyBi4UkA3Cq79S5Edv5Wb8aDQejogpargYkjRJifUJBid
v+dG05hgbl0eeNXAFcv7Lfy7LVx4ivNVZUy+SgHaGLnFtS4C+njU/voSadRThhyaxbXlttXESbhC
49vP4gr0nXhak2lAKhkpytaiSWx5zH5ZxXTpGHzc377XZoh0l4jErksbJfEcxyo6ffzxkgb70Yxs
u3bi5AgQJcUm8N8ZLgsdWqscbcYepLY2OebomIW7+Wqn9VAt06mpenr8WpTjAnrC64Afn44HOOP/
3JB4WhfuEukcrRHvM4qd/XV6PVesj/MpLc+1NcfPonImK9wQeY50DFd1pWzLcMZL+J9A0Tfyl8jW
nHlZINQ5kY4HcQGHEcADmGvGTzZoWy26FE/LLNnhj0LJYJhPagD5W4K10AHccTK424XDDKATh7Ei
to8HpE0/HZdQgw2wGZXhnF8OC1SkOh/zdt7sip389ZMe44RXoBDGMR8z0pUBrq80xzxzksEV4WzM
idZSnTv8ELWlLIdT7toCnDgLPsfOydO3HxnRQ15KzyS2KT4cPTgdo2Sw2woIohDCBeZb1urwAD0r
ee7D+IFsjAFMu+/Fnne3mPAAA8QcrOdA5XxfryWJC9UMe15lODHdzFc1ze5yMioasYkxS7upok1m
6AZE9U8MHM/vDuNp9qSM94mNMUgQl0wfqdCm8QCB0r0slHuI5BoUPNCRACbRdmD6b9AXE7nxLj3S
TpQJ+HCEYZq7FYQ98jPBRJwGG+WC7pIC1HkS04suIhiixeS3gKXmLS+sKmEX0dQdpq+yUviS61VL
Ws6sojpthwNPNZ+InBkwm8xRM/DnDjAqLeBWzV3B9JlvCmASTzE5DzcKPW+FFmLq68Q5eDqia6dy
Olyc8+wE0gKPPHt3F/z3Kvs/vTVf+tx87Fyf6/7+tpSXPjFV4j0cNrTOpoXwFUCVVRkLprkDCIzj
rvft3wmCPaIlBCb4X1jDxFhDrO4mCz7V2Sk9Jfoc8qG9RkuAH/ahLv321dFPGfvNfVU5WzPevKNl
yKLHUbR9hEZa+wVfb1kW/988MHDephPNKi0MSqIAY/fEsRTi1JmMpQqhut0cKW6dCotT5eX+biOz
jv2vKxnwYe4plIhH6U1KkVUhRrdB+wWrhGFvdeiCXFKuHtknIxZtx76Xy8dZ8Gf+yGVqlngvq1wr
wGjVUQAVOfEFQvQP7tdlHezeP0IbtZ2Dlgf8t79wzTuEiX63glUF1hdTzyMRFlMMxjrDrsM8/slR
Ex3cfT51xl5JIHu9qlkkNFi1fFKWT9JHTE9GeL9rc7VDTkDEZyUIgM6pLqK2WBPzD01oZG8yp3DI
ffjxP0eg23f2tkx+3UX4TfbcBpTh4YEdmyAyMGUvGjeAKhfVBJyfneSs+CGZzh5z5rvF37E7K0oe
mEo1zB1clbrSVoWaMckOkEmS70eUM4j8MjRE1ePOaMeMGnw0aKtnPII4kw/5vPjh+MPeLT5HPDRO
jPWXdg3eogLWLxzf7246dGoNl5wOYo9AQgHZIPrU7kUMEtzMLDe2dcaiDAlD++jVMarA8/yVk3mq
teOpga9hhen8j1WVCU3bvhzPk6tFbV4tGI6hrptIbcisefi+o0+waBfRRpXI65qS9a5aRZyLrKKL
/bdgEAQLjmjws3QK1rSmnWxQrbjNqmsIh4eX5N7uMAB2xqjynFiL6w2qKER2XLHKB3uOHBw9o2iP
5z7FPry5h+PjVrfaZWxFwqTUAa9f7KFPIjwZbwBHWViNKIuZf+b3iCcA/g0Ypoeb4ht3MjuMAOfJ
vFybtlk9JKZVNc53x2GrZj3/VH0UcBfjSo3ujs3SW1PQwui+2PsTOOcZlF1nW8EoOWU4t0y1mJqP
I2jHc/SKWaSSs+EpkbUisDn7nJHQSCo8ENzqVAvnJZEhjdoDa9UoK71PEjRHzcGdAYS+AE03LEuW
9fEm7axolchZ5BvRsufUiJJpVJ2Rnl16dT0X4g/WMEszaleinKd1f/c/YEXAVlqksQDDhpnFrH2c
kNp+E124xZMWOJhBji1Eb1OOIk+e9axQIDM+hC6FbtaAHs6g/IBYuy5Xi982JCU/JtSJMaZVbZ8Q
l13DNhMG5EVj2rHHZFQVwaN7wT5c5t9i2eXzO/DUqeckp5MNH8uAaNN6lfiNoGn/bilkisQ0uBFG
/S+QHBEqJ6GMiUuOyZ/6FX0Ma/M1NBn+gYn8Tg9Y+PPriB+NXKBXVysGP3doogx4ADJR4uEy7wC4
S1QQwTllTWMFcdgmd0Tcdomz58BFugzqxZWX5ljsHUoPcEd1qtWmUHsG5vCFkWdVGnK7Aacv2dLi
XpOv9TZymmiCucJ65g5tN9ufdgxsr6N5bhhBebou4TXUn3O/XSVGoskizFV6tzMcduNhuM/M8iUX
yp/g7H/XJzAgJcNExvPa1Ff4nK0W2krLTGbTfI4mTxldUt2uYPPdAlvgTd2AuB0nsP0xarO5pXyb
fwY7wuOBD8LcpDZyhmi1XHQLcao6sWC7EEZY7fPFZ7aA6Z9FxWES+YcUBRE88QTuw2+HImOV6K2i
mekkwSClsX4BgS91osljHRfE9Q2JWRRwo508sFh7totGW0zd0p8+mfPYr/uaWmu+dXWbPSNpK8lC
Wz03iAqDrt5B0cBxYiP2G7vN2O4rGdzuLVACOx+XMwf2bSLfNsVtuv2hwSrIXadfw9Eq8TVGbM3F
QLies3NUak9sp47D2ZM8UWGm1znjOn71Bpb07grPV+qXrcmGYITNYaCQ/p24eMa8sza2X39tZDve
62q+vZqLx0JPZHC587+woslgxdhsWTvFqmv+0X6NCX68buh8i8OvjZw93qMx1mrWgQNEmYhatVas
hVFB9nH/m5UbDzxBO9vMBcIOJpEU40gVpBA5nBroNXxFdayRlp5hTrQCY9bXWRnGjjJZbKnKTxRj
i1dDe7yAaQuDFhH/7g13z6UlKkEId6HDxgWvhwiBA+FjT8dACml1tjtHm7wtS5NTMkvXrMcucbJP
5hRtNoJsrMSFFe0DfcE/RT70eWv/1KzugQYC1kUP0DBsJTIoHPTieR2T1FgW8wdF6Su1SocuCRHJ
yxPzhQ00AtgI8WXkdq+TdcB46wyd2nmb5I/Amri1TvRCxakYgElq4GyTzk/7aSDfPaK02stNUxzK
jKEIdSwHwmAG4OKOg6doslvug70t9zbn5sackiRogy7iEioPxnejxn+AbZ0cA4voxwi3A5UdyVvk
UFLfDd2DfpBf7mgvzazw4d9oiHHG/6MxilLWLQlPMZh4akpGIT+KBGs4O/pCv2FWExpyYxbCONm3
NFIyJS1ARuMqEAyzACFd0dQHtfkWybsWnGBn/iiown9XPkONcIlkoaerqTmWPoXT4CP0hEYFM0ql
BUQr1D5aJER1fy91dEC8O1877lzpJ0kKhsxSE6Wm5T2qVm0u0W9ksToG8sl61FIDnuRdheyRExGx
J7/8Is65rm8VOxn6QPL+rIJxwFGgExjfY/8mTi/MU3SH7hEsU+syzTBnrQEJobz3bgI8Jn7mj3Lk
qkoiI/1RMFaLVL+cASrUG7o/ZFO8HijLgMfzcHrVDS0uXqsGu1SyQGCianJP4WhgcV3hrs+PeAYv
e17aa+U+7AmIAFaZCpb+d0K1KPx49pC4Ft6eBvNojtSMBwXDATRf50petZ6QEUaFM/HDDkHRaYl7
bqiYRFW7q3LkpaKvRwuMxOFeZJ5d9xiAYWyYAZ9TCvCLeUiTZfuReM2N58Rs6nc9AcOvxyq91U8G
Ll2waoYTcql+cJvv+p9wcHYGprDO1vyjV8+4XE5DMc8Y3TrEcx62xGIkppp78oJpvE42THUKaJtR
P+6SL0kupb/hE1q+zd+IDsx1EGPRLtLIBzPCEOQakidrq4ry89EVy/75reNMrdVgH0GUbf3Cro7e
ZbOa7U8e5rl+mpcYfjk2IjiZ5qZEBny645x7/1rLv0EiZGh2NcXjsAJ/6yjGQ+kkp1xdn9oBVIZv
Q0O1le5QTJgirfvB9BD3t2ADfjp4viYP1OISeZzhWkU9bpDVyeaDjBa7oERgROG7AARQStya0g6C
NCXbLOwFUb88jam3/kb4yOlLwyOj5X+5el5jkCNyoSdiuwIvweQIuWnBFQnzU5b9uOFgpz4rqkyI
dr3vFCpBN+27Og0vxfHEXE/JV4480UaOlUwaf7S+ln5AjgURzg9GPmefJRxdCc1UPkRhVevGbDDG
zpjphsApjJySTXhF8lofy9BMqkoU+ucdHI9Jq7Vis7VAc/qr+kwhiQ2R//BxSozrCmh7ATGytxbt
Uzvc3sXy+7L3G1OV+hD9E0LUqtSF6qvkWeJvp9NFQLrfWULwgWrpTz0hRfB313bhG8LDKg+A+v5i
5zdEAOzMuIJyzSYkC2qHOO8z7gLY2P6ZB7Bw0Bcsl/P2fY+jBeN1axWlGsW91zCztDDdPHs5vMBn
xOSq8sXCOgvgMmiSBw2HuLJXPNDMipSOxDuXechjENEGeAJpPCtxjii4+4FkZAsS2DfoN9EPyqRK
WIwvi8JpXbbE5yIkaNocc1qLUFkJv+LGv8/zPUdwSHSMdNGLi7mBQ76JaQ3bs5KJTfu5UDEeifU3
tl3FMq0tw5kQUafRl8TZDNSxRIRxsHCKcVZz/VoxKAR421GnVd0nzzZUwn4+nfZ7CdRgE/zAIFHw
IfBUj0C2lbN6FM9hsszO5FMaoJZbpLjCzG6hnulBi3JORJ+yAewuN/RKYTzV0d3YAGXg+CrfiS+r
wi3DyZsTeaZA3c0F7LgagABAITbScXJ3EYRtiCROQEYs2YnlrlJWfd540UpYKpwtM0ILUQSYF5+Y
FYEf6klMiph6qWKKLvCcSjLspJmCytEMO5/+XCkrcXmRclw4wCnFepC9DQzRYM1S6rAK2KAZdzbp
jVkahzyrveMvVsX5ljtM24RqcpkKTrsze2B8oGf4o9fThOdAi2LBDxXLmu+AdQt8iYDJrd4iFjYG
zCvIxvvpJf/gNU+kJnVg15pibeD2seD2Q+NQnQE1ce+Niz9aLH6i8XW9Fo1RqzOmW9zdLaabMmM3
6X+mR9TmlobIuvViLY9wdTkwaOvoSQEsn34ETOZ/JsEn0OTC7eKZ9upj2voDZkZ9nt/3GSJ5RIB1
/aYKv1WYOnpuxqCzoP1G0STy/maDQuq4la/Gh1LcIzaMWk5RFMRPSSp4/Be4BpwV83cvq8NRFq8c
otDApArV9MEwepITNnPHRnJO7pQqW7EOHly5lTAQq487lzrMzh699/pqnu0/88o9BN9xScBsMdEs
67I+tV8mOBg0/pvYEu+ZRy1LQWFkUIJqtU3TmzT0yNHctHJfK5H5QUJ7sL2PMHlyNSA8fESDRfdB
UKjJwiyn5HG/0BIVLgITPENfSgxotXH4mFjKb1Wb0a/x4xxjRO7bcn5/6gmezOEcTCJGSC13tk90
okCZwEv6akZIhGkmDKzzDqIxcE/z6FMO3yogMaL1WnJ13aR5WE+KLljbzhY+NxIpmtrS+/IiezWC
2lgenrfFgbE9BJFvIsOEW/HNJaitEeIiNQlwWVoDgYf+Rqo4Ey9howH07HZrbNG6AEP4rJLIpeHJ
1rmIlYFkqpgjvMY0+JQkFkEEuWz/bGB5Dyp9MZCGzPEpRlIAJc2O/duOaR55SlHznVJjM2K68V6U
X+k2ZFpIKbnahIuub0WLa41/oibbhI6o+wstHQ4E52PzvCWpk+S0imkLsrxQ8RRR0RxqZ/YpI1ha
vZaST58z3sF8cS4vFWVg+bFpYdEMxUBH3m1dKsQM+Ygga7xWX0w0q27wbhAFkPpu9cWyfqNwcldb
MLe4Zi7Jq1KXqUvTLk15viiuamr9zA2P5vqaZAjtKHWaxRclaoTjSTsjn1OjeohDbvvyCVI0bTXA
FL9Yxzj6ZDlv/oupVOVOkJ7VUs5zq0vuwTu1A/Yi9cha9f8D5DfmvUemnjo6AYFHtuon6tBreWMw
K3YMZo/10bub8E3alxO3gFDOFUhH3Ot9i9gsfmDbLfY1XWkHy4AflxjlGWEa/GSLuBnJoPSK31/f
PwuU2LSzS0S8jHskH7oyoCpa+tN43oFizNWZHezUfErI/I2S6670ZqTxWaT9GHzdK8rZTh2o3wIH
vnaT8Eig8H1xMe0usn1M/TpQj7ZyU2puPdQtmOMcd0KJ+dcEONCRFyH1yNAxFmRRR99StC3C+e7K
aJ6+OVHMqS1a4acWcSs6qklEIXLvDNCYeyTagFhCHHKbxOa9K4fK/D9nbF2lSPwDT6okO6whZk2u
xNsMQ+MTYVpLkzB2t0gOJIAf1vFHLOVeXUl17AjTK0FwwItyYai2LoiCgHOg9B5hxy5lNSckM0p7
cb0zz6ijsUzrmebgpq7qc+UiZFGaZajb2p02ylHmuTeVg62sL3gb2nd6cSl7keYcCZlf20wN4EqN
w9UFMd3KLn7YXbTR34QQcGr5NxunudDkwGe/ZNTcx42riwUyI5lDQNR9ofx25yjwZd5JsrKBMsTc
1aCIb1Wvd5Yj2b03s0vpwM0x9a8mryUvp1/BJRKCS54ZeloS1P4URYkFHiYBILrGo/oOZtXyMmxX
+wZXBXePHE8o5pBduzsTHPOWhDbMG3EFHO2GuhXnI889UPZrJDO70sVARwVKn345yJy2RvBS2/91
L2l6CWztk8P4HHZqg0oNdyX1TBoLldla9217DSo1i9QM1xsSzHZhU7pEbcq/NEmumHCkR3+MUsVh
nI3VPd0hA5OTCoAzPT+mtvlswrIM80pnt7tEWg472YT9rnZBhRN0RDpzcJtOQ+zGcsir45Thd3A6
nOLeZMCGIhc2hcqUXa0vAhlCoWWE3qd9QaAl8RSwKp0z75TvFI57/sj2T2bBZ+884jeS8XsQ0n4a
jW+IgYpup731iTkg52Cu24lGMuSIIV1RvIe8rdWgSL1rJ8cmzVNwsk/eJdbQzFtJVkPPlaIPW4qy
H56Lp8VC41SHkIeOatdHPE9p4ZmMYWFS6t4GoueZOqCU8PglXEdf7K45QZ5arQi9HAySQfwIRYlk
Nq42tQq8W7tSNcyZNZLDMnz8eaTXgVP+SVpOdljDGxUWK8lnP4FMANK480YqS+JuvXWFzMBTOZHk
oynIErLc0xdTk86uZG9rhet94JJ/jaGliHVPqhCfTptxHJIyQjd8p4HC03WSCK+DekfTN6/n4mDU
es4C7T6L9boTLMQ7RV0jgFzCg7uXqbu+epnr4xErhufUKUxUYxZ+Nj8RFYgzojkEmQ0oF7ZYzKSU
VTNBXUkP0Hx5sRCUbNuvbdvFISTFv5JvK4dMQqn+PnhGzcazk3k4Fm9jm5QN7NZEFgR0STuwMrKH
ctwGmTVwjdjAW/ADCP7Me5BAxgVR8SarZAb3RNW3xbT+INdAMHmBgv1nsRpTWlSlaNsHRv3ilB8H
zc5l7A2rmvZB68Z3EsGUlHjOXv5N0B1Bn9i9H+BN98GNyOEgudPeMsKMTpXK2VFCu1sk8GrvQdxF
nRICFU5yPpnVjcb3zJUgpGtCMqoduORwUZnZlvI+2AtYGvC9ce+MSiUji8HTm+vSnnaUmOwQ5oPs
Mgb8oPKNubNef4ZJwVp6jFbLEJWfE4go6bzeqMyQtRNdx+Wag2P4NLWEZbBL+fC/+jbDieMLkgyC
DGQqTrqTK6+mcMLPtIzSYVLoGNKq4cw2QJ4dsW8jxAntApooLY+1Di9Vtwb3YsPKpOWyLPwbSsHA
R8iIKmeIu4ac0wJiwgdRkVaPOr7oAqNvBmspuduv12AKqOOLtAZpROz+jxIxCIWWY6IpQjNWlIyW
R/1ccm+k+nfCbttVztVaj82lv20BZTU5LLbgPCEoo+9yHQx8YQNv2XWowmRN43nIB9XpPnY1PL6h
pWHVvJb/kgttFEtY8NEokIa6MP8+ISvQAmYIaclmxNzMo2dtm//AOyoIq3Qo6GJp6cs3keZBYJ8W
XUHpBDEk5WDY8l4uRrbv4iemDwvDC+6CwlkHoUCEVk4w6/j80L0c6zTO5xyf1x2rDtKNi1mT94L5
pTCEvNCWke2LjiZ606D04P7BfCQFBKAZJkpTfGZmeM54SQBiBNY/ZBJbMqPBEWiysjhsTrjkJvdK
aKhp2gKIgLBXHjzbp3H+azXuk2VU4ih0NUOQ71wHpRVImGbMlQbDZyWp5xV2irzFWOjJRj0uGp05
zwsNxJlPop86hWDwvGr1A69z0prP4G6Fz0/6qrrYBuGa4G4fXwCG7WTVNmdKPRAtwZg7FhJkTbmp
aInX2Er3fR3w8e4tSakAbvMfhJGPmwMHST4ocgkrWKDit4Vuzw2p2EcjCG3pYkswu3KDwo6kUdcJ
3N1hbgH2XSvUWrSIsEPr9DlxC1Hnc3M5hsFNWe05ngI05hkaBc4jJF0mpRAzpjY8uJjLILd+5cDp
5Y4kgW9aL8KJ/QKaKK8jssMhB3heITps6X5D8op7+WyX70ogxCiEcEOaSQ+X0dJmG9n62oUVeB2b
1w50MuRajFnkwv5KooE3PEjwIjrzpDdbtozPUMUJTRbtvyTwgo+9IXr69NKI4zWbYALcQmaa5ZbZ
97hVU/8THzAhTO/t/gq8iAKHJygHQ10S/y7TC+2W0AXZSOxKxx0LVYb2SOiAU4xAyX3gxUZ++lWw
ScU5ZJw+zPpBxNxHHJJ1GkmuZg2PT7VQGpmS1CmsKE2zl6UyXsdBBA5IpYjXOXfSa764+OjwDB+x
yO2qmYyeXmTvicxT3bfOT4NAiLhbmOdE+C/HkB2Uj/9yL5HzpiF1t9IA45hZW2eKiUueL5q8b7S4
1B7ZhQr2lonPaX08yUDVIJU0efFCsDig0QWlAoqJUWu8Wen0nasBo+t9ZvvDTfFU3r8KlfBtdKZL
CQ0qLzQcoDLa6ZkD4nY+OrocruABgGLk088AFwykOa8POdR0spA4zK/RCU2nIbtrvy7EA+OAsyVu
KcNd36VbUhDWozzEy41D2b67t9n0o+/27/g7UwApoUM5j4UiurxAhfmZ3eT5yJfbwzjTvnulyQaZ
nYw9zaEqoyz4MTRHg7CIsXsuEAwsM56CkSLTyVCh5Ozr0UM7TFSnlmS/eKMUaR4RfROQXDESmfJc
LCCW95+tApgwO1MoPu5zOKb3wEvxD+4YI9l0duaS9ltXVY8/4LH6YD25p+J6EFO9I9RNfM+kDxDq
3dToh0PUYtN8VGYGbQUELmLZIockBV1jHBN8bbNLpV+izY/57n7hHNvMJ6gCKMEvDlCnwERGLr0G
ygQ30a4rLaWS5/wHNBuYg0wezFcNV2n/hSULxMQw4bsJmzpOwgA6Qe0l6V5m1Crd+rgdWpnISBUU
I7Cwya2RQT+8blyhYBf/B4iQLbuWa9eX19QQUxsvHb2I+bu4r8/OkeplooTtvwuVFf2Gp0zyCfny
lhORcHdxY6RxV5BIj7zijod54GffRs1FV2XTxITMEufqvyEj0KtF3tYtDZqnOsCg1fmIBx5Ro2Mp
08iBCYJcIBplm20LnzIb1DtENmpUxn6fN4wx9eUtDX3o8VlwcG3gIXSm23QX5ZAIToduaKesMdLD
Z3ddx01W6S2lWEKUNpVF+wYNGUzTSE6dHWv4UgtgFSo2LbeF7pO9dtn71C+DWZSAowJy+2V13C1b
SKjIaz263YdlPeDCox9WPxKBy7UZmjHsTke19Z/A6JEkivuKbwox01qppLEhZlD8vvR6Azkw/GdU
8u5B35MQcyBdCKb7bZJgRWC9l9yAXo0UCuXqAdIczEwYLn4wXUakNDmvJrUu4kHehbc+cdw41il9
e+jYlyPbM915dXoYqq1Jr1+hAPgI97MhqpBnax8fGWsRd4pB/3Y3RNYy1F3UPAV4IT+kJfq2sgIi
4o01bncSVnwPNdxRpqJOyRL4DLJkg0ywMDpYeNVIqlhgCyK3CgValu8mNm0MrxatAbA2vpjK1/U8
FXWBXpsdz+HjVvksGaxIU1yijo6/P2qZUi1R9Sc2wH0sbhaosDVPsM/TtqAzj/sbhCp8d2VacymY
sh/+W3FyWHINXB+BFgTdjouQOgOQK8F5wZu5Ry/5WcMltCw64pBtBMQ/impiPBmXsQiqwSzLxRiL
48NTu+h9ZKV8a1HOFvnnyIuUiPbLJMiDctAhYhgclIEmQZ9qDeU1AvYlZwrZP3WA/V+H1XG0teHN
UhUM2cbxNdItx4bdhzBtH5bTFH/2c9CFLwsZnBUtrB8JN51Mfrzd/B1klzwa56eTyynLxNrAFN2L
+fNVrjmHGR5BW/rAGJjhe20vi3/Gsfe6wMBH5JPFhCvdEGPuifJLl3eDimDOHJHLs4T7gfhJ2xEz
PKAvFQoTrih3xn+fOeoAQO9uYGbxnn4XYn6FpWCmHYdzsqYbs19wUNNoK65C8pCWSLNGDtjgaw5y
GAgIG1XCs17uM0fySlzjI2/+713sc32G1Azsa8Xb0vk3viiLpWdvG3dFgwXiX4XpKr4Xi9oBuEC8
EKf5n7b0cZQWSjyNNj2liZVkUz7dgAGSVi1L+BmaIVN2gFUszvt53jSrjypxRbZfTjitDbVLgtuV
ttJfeK65bdyTpOqAQW4RCj7iEf7/89OYXga0ja8FL4cgirhyx8N3Qkoo7IIatdlXvCLrRa7UYDqk
2leeR7ny87qqzCR9kB0oX47zWfUUpndExSlc18d6OvGpfLGN7Ej+SiSfQKsujMs+hYkeIkHxrtY0
uK5OKymZ+BkuCd8O5sVEBEPU6h/dSTovyv3AOmzBa0LTmzEgd5TP6P4ScaY3V4PV5nhxVjiktWNx
/gqYv5Zkl4GgJwL64IiXU5hEC9ifyOM3YvfOhOB+mArhyZZnQR7DhNxcfFzdGEUmFOIFmqS2znee
zy6/HjlF8uGmsdWsfGp9NjmTp2u99rFnJkW3SNxONif+eQsk9DwX7S7oDsc8GiZ9u3fYXGWt4DrY
dxrKJjSyfvdOY2nxpIt6jXY3Jocgo+zQM94NMEG1Bxog9Vq4CdDVUFr2PW1wXBghp5BAYLFnrFY9
9aCjCKbVKhElRUDQrfEpzRq69JtR5xoPzO2XMxdwDRQrgicDQsaLd0YxoT9KUIyLkjpDJflPbqYw
R7pIXQoOGAlgSVdnmVflafo23qDh2wNGzQoUUOSeq0lFy5ioYhygHoxy+rzbD6qo8vNBXBDuHhxC
MV6gGafLoR7Ks422sBwqaC824n0VuBTF8LSmHygZkGXjXse5YOd1CtK8Ojo+lAaKMg0QOQsiHmQJ
Ba4vc7ob86culyc2udx3WWdRd1TMQO3lLlHxIBWApaxAwq207UuTU+JSdHIHE0T6cA24gf0waHuB
80nUqj17UKLIkrLCX9CPIM8xGbsIEixhOyLBFT4TPIgPWSVDO0cBIuyinxXhTP3YkkM2/4R7LcYb
nfgUVpOIwh5ssQpOyPoX/57wNcZ4rw5Ri8+SGkhxMPM57G1mwQ4brvOp/TCeox0+NKB+y8RZi8gA
KS4HcJuT/Sn4Jo5QbEvxfE4LP1qJpPK3ifxoz9gSMUO+sVbe3mE151mC5JiQlqAfHXq5Y8sS3XN5
o/Hu9N6xvLMpJtgkIQodRBXzhPeVTmGRsZ5GVeoWqg7mkLAMfOhd5V40/ftwQcpMd+PZgN+4+DRP
dbRDkmX8udI6CARdtTWN5aelLYS3a/6uoeK07H1LFQ3OXkM7GmFOOPGF4ux6DqsgqrrYY1//WONG
PBq/EvoxE0ACTH3aDfCZbVhH3cpzcMwRY8HvkxL+8E+3o/KmpjjSsoP1zOUCSPMMo+aAD7F00wEW
rYQ3iRjqrx7q/fDAezmDSudDfv3L8FXYK22lXKPg31N1aj+jaxpYwGFzabbs7xq5SrVtUntoYQrf
rt6X5DRzvmAdEhrCZDmqh3UkpWNiN0jArXGjeTCK++cEWTEoKO9ba86Kh3hRgpJF3wOLQRKbhAuI
YrMrJMc+QX9ManebClSAIWMIQB8L071F2fY/8axjuR2vvwbU/vbsYxUd+Rvu1fWV1R23ikThWFZl
Kms/nBmTOWzwVYYPjojCHtCwb94M2mZx362N2ydaWw1pQ2kk79jsABhQsWQgDi4ivEat9k2zNISO
v35R84D64c3A1eQaK8Pz4CXjj+1ZlcyNfbSNkFRsn1v0avkximMb5ilC6a/ngBg3/TtiY5JmAqSF
9x4+9DmhS5UR8uGioyGt28QAwnZkrqXuqO7vfRx5lhZsoV+z+KUsdrlXb1QIIdxxPM6+mZWkwDYB
JZcBQOblFZVhFj7SinJ7RvzzvPpQgVshMFpnCNj62dtAN/BsUiqQXXbcjdnpt2lrHwKNsrMp1MWP
6MWmQ6onW9tWzB8u//VtfQukDg28Zo41+OfAbdBZDEMy0DB657Z4QMSAyIaVTxV7wPF8GeI1wdt5
6O0TkqyJ+YQGUOrYhOP70CPy2YPpB5zxqVyM3W0Tul5IiAkx5jbmooapwjxJjftmrK7TeQqf8Qed
2StcyUtPQhvLDsrJ89VS+ASupuxra6Tntj5WJdXQZT/ePR468mxlNIs/CeyWMAQ0xgJkBQsolNZK
BtCtqcEGzKnnTXnmYPTSTlQZmTrA2gATSQBHnWgsaEfGmuSVMT515ESxUPFEWMITEAfLo+TUle/n
im0xX/MSFAL6X7sObtjunA+hzdjHvHCmsYMW5yiiKiOTYvh8fQwIR4S04UHdgu0dbslP4YyOIcif
BpaTWbb5Y2ZnyoWmBdHKN1eibEs5Qd7jO0w416TErHQbeWRdofDQ27ZxFyQDb1Dgd5tBz9IJ5liU
XP8NuMfy6jbbWgHQ7BT119w1VkfTHZ2SM1e+kZmi0wY0fICIZcsONoo6khHeI72QvB4PJU/0twKO
1gHKHSq7IyQSAsxbFjDRG1hABuuANFXm0sJ2Mlvhn/KXPLTn+PhIa9+LvaL71yl/mnbncc15MQMV
WH9gDzOl5B6XW4xFgKV/4nAAFHEa16Lc1GzQfteg+mZ/IZDEGogCV0MtkodUqt5XUVVa93sJoEO3
8ElYc6TWxVNOts3UUJI5PZa7l6/LDJxYl6capE59YfSlLi6kAZ/iMOncmTaFZqLEnk/0CKtEJpcI
MqHLwqMVsZwW9u7As0xJUB8IbliTWIraKF6j7CKxW/AfoCb2X4ch33j75vWRaEj2pqVozxZUD4d7
0IHKOzcFkPsIYddytyyBNCkAlyp6irJymgrO/jv1BimJjcF+4FPr4h7ioTQaYt336m7Kkn2nO7D9
QE84WvhChmnavEquvoRBAvtbApW7/QYp4SonNZ1vBsa6lz68JxIIXE+ePwcVQR0p0B4vCj/oo/6z
tkaaIMdochimb3Nrm4BVmxE/VpPiIGpoubEW/4kyN9CAHk6cSttboNqyKpyyc4mHshqdtHu5W1WE
oheT9e6Ie8hcYMWPfWc3obMcF5ebVYkmu4USY0fdYpaOcO0XqO41UEdl7QRMjvd4wHLQ1jIQKBVh
eeh0HCG0izDiGZl2tUy05r+pLKphlvFS8dDinvLHWXdlEg12UK2arkV4KhRIRYtaNRDGARijfhux
T95ygmFgS7AACWAY3w7XGKuRlQK13V4I3UXoyRp69553bhVLyoFQ7rH5Ighf+XTANFpM2cMP9Nt9
hDykWQO8nvMY8EL5U3BdOxhXdB2EID1jvbAZA15un+qryzAgYIlb6xU2akGPOGGb5sXvIrpUJgSM
WoIJq4QiDwi9AyjBIVryoeF7O99jU+oRpl0YCA+i3C22lpg5hRlExReJ5OuuAtw63EWNJXXMtrQv
/X7oOAMugh/924tSa0jsvsT2Ah0NJi3mPp+ic6V5iKl9+zJolQv6UwDlmYkqlCH7ohb50GRaCCKO
+rxdQUtsIzwJPBW1nZpXpNhWNYT4AknJZR5XPCI0pfnhh8H9uRNzAXuB7EGYFXdDEhxlqk7iBVv5
YSLL0vsLFXT9igqG1JxLri0oLfIPJguipU2U1us6u+EVtj9sCMonDs8LwED1i7vURXoyHZDjWKfM
IGgdzBvNPJPKgTEU0c6ILidxsiQusadz0uFPooRNoLk/XIAGEQfjDTcodV8YbNyEUykjCJ6RqjhC
Vb2/a1ef+Oaah7VQeAj7btLRJCoKC+AaFRH+LKQFs0tSslGrvmPVbflLBSLMQ0qR3R/9KBwJgwEm
6TTFcP+mXQGLGkXujTJPr+rwSZ1WQXZhLS6upcN/vxfCyha6R3LXMpIfsfiZUpFkVC2YEz7i139C
AkS6LzWCF0dagRlfyy5Bt5zFKxe+H+Nwm0LGKjmNMwy3JZPNqVAQxBr5cQyc4uDS/fbXLlsCIHnU
32agCUJmzZoHo3cU8ciKcAdsQlipDNMAK2irrleMG5gPioKdFQWpg0Zbhjs1Adr9hbTXhTGyZ1gk
4qxuEXNqNrnJrdei+82W9iN2Avhbob2gWY0tnFSVo/gaKPL+/VtQ0U4DrHK4LWFNxP8h3OePHLot
6v2wihLx+jwEoeioTjqnhGrzOwweb1N2K82HrMWzRhPwtLHvKDfqSwuH5eC+hHCqiLkzeo71d+ab
5fEwzH3L8HpYKd+P3hMzCEFb69gamSHm7KcAHSA5jot4+JjMtOGR0ZWCIUtkf9HM82Sbq4pYKaxX
SAgwCIfsCRBl39wbzdhMd+X9OuVV5A3k5Hs84kt+uLBAaaclXJ7AMrlPl61SHhtKPPv+1zpodxRy
aku8oOx83lrUq/IJCYMZMQcXGlVesOgCBfVmhfF7ZVzbXX0DPtEIGLrIVS/3ujWvqbqdMDYI/FmU
ZFjT6/F7Ibz3HPIcfst4008rPPH8IagHRt1EHnxkJ37HLdfFC1yGRMtqYrnM3QL1DQW5nj9S83uW
7To3tCnqMlhhYD5qbVd42J8RnFH6R3dG34WwrPvyEX9mPzGYCg7pSWLo08Kjnr8i4w0UM77joykY
sB2/E05ebxbki7ZH4bX9ei+sXjRaqtGsJ7ifspXmHXVLbFE1qVbz4Ml2K3ba+MhGVOnGfq8OPHOY
FjMB3vCyFoE761dqcMWfY9diaEMVCWrRrHH12Gun3N20NC4zzd1gE8yvBvu/8JME/M/pJHkVBTeL
HAbrOo6Jpc8gnZOSR5mmgyRLOM3tyC/3qFL8EMjJYNjzCYGbokUSX3uuHCqV3v7OfNmC5YobVOor
6H3SeuQ1c6/blcA2IYo86Ul04TnyGC6N6lzzT87ygKswGlpWgwYRaS3bKIk41FmjlDuH96GAENUX
v5KdHRJE3teLi2bgIrE5ljK8tUqD0NQwqYBQ6+tPeCBM8LadPJGl58r1+B/3oFBmX0WwrJKvufzW
ejKYRyk2YeRuiggXLcbTvut40Ib+HXI8riMelrbi88dxWZCc+BuIZsG3tzLTUngJcUzIcqUwfzoB
5f8OvTBmmpezif+b6UpmK+z+Y7OfF7I4KRng86MbGnvgrPoHf3HlKucnFHxOS+3JVpKqwzWK/kEL
sZy5BqCIF54GddHLpvcjMsOE+7k4/z3063fVHt6Uoevnr8hVNAXUYOLxQadJsnC7zrJcYOfebCv7
TAuUibYkw8BdH7IenwnNAr59vHXjm2c8e43cTRbGOeohIe37kMwuQlyr0Q7qPzlldPqVxbqxAgr/
U5NURDjrvodBw1enHKOXbsRHscsyIWbwpX8fev/dxYfL2S1te3DQdtyDKFvpMf9BsYWAP7MENKAp
dumxQaNlmMBGDkUkBjZWPmGcSndtTO6uy0V+dUoIkK12a9Oj4IqSMOKCmk+iM0Y57ofgwlOJ4BVN
JmSv4AOfb06aBWEgcwK5476f0TCO+gCkG/4S78I6JYWul/ja9hDV7i/J/XhKfg7tNbgdq9vZYYm1
84ma8b15SixoZ+XydbwB3qs8kxPuh3eQQzhApHEOYVVllDpfVCSGwaSUuGiIgy64yd/Br6Clv4qI
pCIE3f0BPNQalEtY2u0m2ympY+ZUYcwtesz8Chyf5D/SX/W8Nh2hCsI6V7QFHB6pM8gng9iTpEZe
GQNdl/b/UtTZMQc4bn+LP3aHzQLMibosp+c7demuqBa1OAJOHf29AcEV4FfCoWPcxSWNcbjfEdeW
Y4culTDcerJGB073UhV9rqsYD9MKFPkc8G625FgVjMU0gTo3Am461AkLV419yzHUkRMf5edGEAq5
xm+GZAmzrHN+njjAd1mKxb83zTHTNqxNXPa2n+VIyX50dyRkk0vWAP5xAPL15B1GGjIE1ajSyS/M
a9nzzGvNhzk39AQiOyUkDIWJiect1Qusty6/Z4di9/EjYU5kUDwOZ+MbsDe4E/kt8eMBA0csH7j0
4GCp0v4ukaJRzP36UabJiD+zwDveAOX2DXvnP2m7lPSDPCK3G1vsBFK32yfjT+V1IEt9GKDY0rUU
AiZPgLEc/EpgPDmgWNpvXS7I8ZrOqsD/sod4cUlTwaGza6rZ2KE9U+axcbp+5afv7o0aV6EWGQ8Y
BSbo+N+ABI07Gn7/IIn6oo0RzUJD7PQVfZ3ysQkPEKJawr+Q55Pm/U1pNioDNRyuzXso9XifZy8I
yecMjNz8MWnlgS529yFga9oLnhwBuLL38JnDJuEmQ6uDYxz+npwO/QPNDVT5dcTn14XqR4e/SlVX
GIXl2OE+IUsvbJqne4vldl6wGI5qEusyCVVRsQmjhDgJgr2EjyRPTllXVdZgAin9Uvbm0/bacQ/n
Ya2MQlOx+5bIDI58eouAgagBNL5JDhjM8tLzT+V5RTjgotGhIBjEmEjUXdsTkZ9BK8RbgxxIIyzI
vOMCfa5NkQXIOplWjZDJ+O6S0obGMPcEOdTtt9JK+CSLtNLAsTm847bJkHeNYg8Pb7WfBvtRVdsU
cDRmCDGDoRl9Y9ZQgSIw1V2p8COtc2GAX9pbrvi8OMVf5iRO/2jBWF+kDoL9GW8MEKBu9EEUWEiS
eoPt9SQ9//Gfqi79DYlCzMDOUMrDueQ2ru5pjxJCotLQuwKVt0oD5y3BK35ybuBpGfFEcSwQw6cC
B3pjOLCF7HX+hJlrI10341m3bzponmEyaicEzASO5OIsQokA9MJ4PxqZJkp7a+ydwAnTSd2N7eyo
IZnCI/W94mLlQr8Klq6Ex5CXZL/7e+xBbRm4YVXfhFZCtrIOoIyeAkjjckt7DVyB4eCOHManf5u7
mFKY31bKcjLHqdjiucv+4l9n2Tsowm5LEaOPq9V/B8bbLlKqJs37ajdFoc0HR4bq9PLvSXyavM0x
mV2JgPNoIyVS6S/n251RoCkOVmenBkYAh4JLY9oWzm0pbbTAG5ou9F4jqkbOSz0b4io0iesZU3KF
Gvy8a7SyLCQxhFHBYwaZt4VB5qtKO37ALkT9i+yvG3yepJlzsF66cZHPOSo+lSKaGyeX1JH2PhAj
JygwSVWNxyCANpbVPpWHssgpmFkaXAu17g1zGGVhuOF0W6HDKiCwOBg9661DWLCo5sRbKCyE64VJ
TxZdFthMwLPYMO+I2Cn9R2GZjetyY5/JKxCfuxlE4wn9CwpNsnqozWrE4vwGVGRDznPVH33aOhIL
Wj2fP/bySrrl3AcfYdE3syyh0efcuhJr8bgoy8UvdkThbOELUMj7C/2/IaCXkMpuK+9IbRaZZLac
gag1sosoarA3qNBKM5X9i60GQ6Yje4xs3juVjR/UUBEnZBQNosG3GfWMO2HGgslmTWU3mJlKIg2l
TY/iGpMo+Z6cq6ueQ24JXYYmqcKwFIvHC/JEvuis3vzuC1hxybtdm1oc8LwVDXvt+TgXh9L3MI0V
UgZX/boHFUNFEAXnAJit44PEbEsxrFPkITX6Cpg5aN1HvQVrMEHXSEGFtxja/pMdM2RFj9MrQo7k
L7AcYnmXcizIOwuBLOrUA/34jVz0ZLKBXsvJZvPYXNMVVJEpNGXESQiNfYrnJROQBE4x5HE4X54P
Lf7w5moLTqyYTPw2HY+1US+2OhZ+2pWEd2T0m9RaMXg+PIT1n+JVpYiNV2Yz6QJP8r4jWrET4l3k
xaWmGW5Sk3aaWtjglcCMdpbEN+Di3DuqZo16GTUuSBMFJFkh8juH2xHbOZv24gRA2PDPHlBKlJJZ
wWnxtjjbqewPYxV+UDRhOTS68Q2WHCVSZzAW/QNxshmxMtGpcGGvJiEgS877pgnIq4HraJOj0muY
K6LsvlJ2ZxM/22u0F7I6SvHWF+/H6J+q3FP5aMqrFkKwJ4sYbYSSc021kOMxdLoO96gF2LeCIREe
d8Iw7s7K/PIyi/efnH2QGlx2O405bE09xWTh9SbiCdR+0bfs7zkKB6FaseEdCMyTM2St6tJswzwC
YkHgn+Wt29CZE1h8tkPK1tfEKtOTh5eeNtNyDCxuQTqG+cDNebOZ9WQzULrj8I7EuanzKnuf/p1V
RJya08YqPCGzAKqWEGTvbXgIrBchrfjDhF3vaSy68kWIgTOi35/N0cGwUaOX0wmNdk4GekVSw/Co
NgjC3QJtCwvFQzh8dE1SRpEaj1yM44XgXpHRYO1J3gimsTc4uZPUoORCpLobionX9XCA/ng7muv9
UOSbVtCmo+t67a2B5v/Z170CjOcIxCxSdL3V6g78OqxNpUzEHId869KushEzCFZ18K6snWMpUu9D
NYzTbyMi9YoeLwSMboJ6ZUhnjnBCr24Fli8PNqzMw394B43fQ94F15AC4ZMGK6fgGdvCpVoY2Aeg
HzzgDtx1Dg1oS2LsgshgG2dahx7NyXL6kLsRrVfWg5KA0HQ2mT7NhrJW4zEjR9UdJSIFZqDdlje6
SyMyXkGY2ta8Qrq/sbv0IL2oqK4r8pxeGfaKzox87gmBzZeYywUquAg2Xj3qLfvVgqT5Cml0LqUG
Ai3nQysXjeuqCTfTvH+oTR1nDpLNp6eu53RcvYrt9iaVDNoHzSIkkLWWjd3ylpNHfrOLoAp8o2xm
zRh0m/WkOiZ3i93AE4LEefuVluL9wLXeWAlIT1/GRsvU6j+kFyAE/jx66W0OYx9xPnD5F/ehH5AR
yQUZ2vza8JHJonN4qPlDe8E1K8kCkWaaUWKPMcDrL/vDO+voHlMvI85fyZ2D98GAF2F7EcxLfO2Q
7j/VSEtMJM00jWbxSat+CvFs0Kg0GmQFk5moMZCO7arTNBm5NvhUWDi3XzQRZuSxzQN+9DSHQTBl
wJhqC8onJkxBtI8FMl/xAh6MFmbqMr49ZO1DxckBdsm+Fx8c4G4R+ICqsRGXK/yMmMOCm36LkcY0
d/XSQaUyKmeAAtxzC2j/9fXtnLdIApNYVT3rChUBwPYdZIbAqBbzRpPAJNCrynTrfYU+wNxWrX88
FZVp6KQHpirAz22YE1oD5DUc/xXMIf+hA/LbaVQjDl2QWoJQusx4JSuWSkT69VxgckRGHk1wzhbS
27P8AYEIdYptfWAuwUlRnlXIcO55/Xw+u6jrciGjtNtaztEaGKkqas9833p6Jdlc6SIIUMMqmgHt
XG9yZs3usHg6mGtQ35a9Qt+HvcO6DivPrY372kLOcV3WIlnQHBgZ5DvVmh+hypW7IglkTXwgQiY5
InnztaAnEQmj2Etc5Iqs6yaFhztgBQyRysfi5KDizKODJPVFYSV/kktCznwD8d/g9mYXgFiHM06C
S8DgUpTvsZ0hciZ9iLkM8E36axE33PG/H2kRyV1OdiJ3M8+tKywaQ6fY43Br9Ms4z2bduhZTYRnF
keHPFRevHWtpWoY1BpyDMYIhEv/SAW1j/Dx/6kOCfKVHFJS23lvySmpy/YFwzrN0rrHqjIqTQBwl
pczACu9pieoxcubAxKY3QhEDq5fn7mJ5XPAA1aDC2TIt5lamObjnAt0itFW1neKnkTVu++moOot2
Bezh67kYfaL8VXv3SjKfpeYh3SWSflCuLjO6N56cRwEy0YEc+utPI50xuCNLmL72RkZ8bkgvcyBq
YpzmRHfjBdF2ZzvyjWC6vWteUxZD8o7CCcKDHwxtgIhdepVg+oQqAjZeG4GsznIoH/z241ukccrf
19MfU1oCx8oVklpjItqLAkZtyT53Nms/9sEVe7AHP8ZonDhPRJhpLUSSVvrEFxjGmcmWVCoMJZsW
AWJ02Ftjl4d0As2c9rl16+d7Ymz1ighjqv9o9B6lpcwRYQfwpAS+xcuUYRsEjdv9C0DhKPfwNNB1
2toMNv6akcDa3rerhj/a10HlZE+RCpp2n8uh7QsyVz1GlUUJRW651XCXSGNZPncpFFGR6G1CZyF9
MAWBCpyIT4Ajky6ter6t+7Ap31wX64PPe2yH/zPftNbo0xIu2PWY/DYxu8IZYBP7Xz3yKtZpVJI+
BzMY606EfGj4Pg6SpND5TF0x6igCyl3FK0SZwfLJAz6txgbHYkTsrxnTsJaeeNW35kvLtwCt2hEG
s0utSPMQuf8WcFVdcqLYJLzuwhr0R+/KiGcCTJ2IbiB4tL/9i88uWv2POpR74pD26tC4q2eW7xx+
iYF7Melv8zXr5UzTtRDvE9VQiIAnmNzHmsPOUFBD4M0qOGRska7fB7txGknuT52TAbyIjNc9LwED
GeQPfqeKPlGhg/OwdGPOtUx2SgsDtPCNdjAosmY5EIQZwkkljH/C/98jtz6/OjOCsabYWTY+Ice1
hWDX0NJxxYFwDJr5LA74wFaNGd7yOnqsKps3ekuWUFLXtP3cjN+NMuBcqB/QW3iv+RvypBaKMFJH
jdT3btR/SrviTBKsppn3kkwMWXaWR4g5aREBM9pr6FaGStngOGcfbO1v8qG/X9uWMei3p9uc+W/3
VZiA7y/tpjCxJbMPp2c0yuqBDpi9hrik4nkmTjFfMol1qbSOqj2WazzSkdQ1dBo2BVs5UlCg3vL5
bAQ3KJh1PZ/fQm7ixGinsBpoz7EzM9TiFau0t7PPekdaQEr8B2lfEvj+ei53fzolg9zwmVxIJDIj
JcT2qQSB9TPuukhg/PQaOzFQD7d0i4A6m/RqwGYGYqnthcmU8GJN1FedC1F+X8xAbQnJvkZr8GcE
GefSt5w3t1gPbjPVjhicoqU0o/vju0uM0IRPYGZUXfZr+KO56e3hklnnc9iHABpFokHKu9kKG8tu
9rZqQiHxhg8FsO8cuplQdIkr5wNzmQtsS0ZOb3BxOI3Z4muOC5DzgubvLgqAgLcqLZSqaUYt7Yz3
vreUMBlVC2Ho5tDgVvDSKnZn3Cmd0BTs5W15G2n0N/GC2LAjG0Lm9TjOi8aBUGHpAjqDsSaRVLMH
jCkb58utc5d9ghQpNTs+eQL8H6FFQkQSD2yNvHe7zVI/Il17/4SKfum+Xl/GUOb6UT5XCFabUZh3
rAuo7nKHEdyTHL+IEKuR/u/i/bqAOnsnlQKTCok21Ou2tIyg9L9Ub4cxsPh9NVOn9b6T8SepLuhT
tpP1Hi0yhl8D1F1byn6YhU92hKS3PIi4rtHJau5g5CS/4oIRwZ8eyGiRMDfPETtFKKzDkWOlTb4e
bvhk+citKtX52NVaP2kpVB2zJQCsvqE4BgsvE+vrtg8TbB5ExpoABVPiiAh8xLpFAR4orNN9YQyF
9SDnJ8X4O+CJkxSyPkvQQVSweOK2+OC+vwnIw1yTZGCt+DazRAdoWzwmn0zlEDKlPO/xfKN/gdUO
4SjQFr/Q4k1exhjtH06GIRlNhTJ3/GbPi3E2ZndnVhLzF+K2MM19UM6ST6O8Gbn78jW4GGav3emb
3/oh40b2eFZDkME9exNhmXMPEnkFk+01bAlEjroUs28ewGKJegrhsM8rwzGSeMwMd4ZIUZjnAbfF
1GopXD+XWGgPk+NPx76RUuImFVWjP+aJEpPJJ9B4Oqan7lnOYo9j8QLLPUmSAo/BfgIS/MIeIuNS
oC377egtNK+hp81VKfVpY0hucGOHMZoFV0mj/5IBs6iO2r7ooQbubr+Ujlhn5jB5YGWOQfHtTKlA
uxvRbw7Eyfg3H8WPePswCXamkgKL+16/QQsPJmS2auk9qgLi4vlDhDdI4L5B04VI8E3f45uN+wIu
rdLxAZanayAUkVN5EV0DTLS5Q100XM1dcToPKd/RxuxafcAplyRkqyBmnOqoJlgMUaOgYePYQuzY
mXZK6UvN7wCAL3figNEwdOnbdlFlYIMbSNFrMsOmn6OjHHUWuwt/4J6AWvvrcf7CV1eGCW70257G
SmA4KIdkml7KF6KRjwym1vJkoigo3oHbjhK32KUOBkMKvw67JCfeWhY6ok9TNXKtGJsShSy5lkno
A2elTImBUO5DUL6O+MzmJBNuAKIIMYzosqA3Y39AYkJXhk2VMba2aMdtHZMQNyuIDCSftPPGjco3
mYdDo/zhH2kTUmr16TQCVxLKjRGj88z/kC7cQ1nWzsVTs+FGheVipjn3hXH8rB71dYWBKyswPFnX
HbzsJv/YlsJZMb1E7BM4FYA2hH6F0isv3VMvYWWz3DkFUQdR1J6lf9illif1yShYt2Mx3AcGb6aV
sVdRF/ko3MYUmkmHUK9buQNJie/NZWW7iSKJs2h/dIR6sTPs72eCW8yP782p8VgHCm0VNG3bYOlU
mY/G0FUlqGuUx2B1QgXRq66Y2OPsKD9kHzDFnXCyOOYYqlls6FPWIxymVv42LaXjiFctwY8MwQIO
B8Mu4t8G4Wtad2qLyj7gaJl6g0YX+gyvkNxM3lJ7n6yMfWtIx32vCOOU4hZE+GKQ4gj/kYxp6Xdb
W0BDk43mkOxKBXAxzYtowI20RF5Jg4cEFZ4tKhCBRo3DiXUPXH2ba6bEla3+Lrz9ccPhP7GLoXrq
bT3ue4BSwWSNKT8Cjgo8wLIXeR8sXWgrpLea2umqef41uLF4v50++I6QrAcCjwHMWqiTQ6GsfMO7
BXrqB+IkxIlBAyWDBuc+GJ8/AfDwSBTuTNvucQv1XCf8cIoNWZ/49JUAMZUFuUbX5s1RYIb8JOYp
6DkrHKNMI59OWe3MgR6ubifHsrwg48y+wSjKjB3Eg4dG8gbiNLj+B9GrtIIl1TVQcaOIxMm9xMjR
v0eabZBhk2RmqeoynFObJ6CAC0t7IZtw/B17foz5HtqZsA8EVIXZJrA20y9oqQVbnZlK9bnqfVkD
fz8rWitug6yuD0nZw6iSVoi6Osm2biT1YIkPnyjaFArsd3xVNC4WzSKsprX7/9r4WaX6Z1q8CKiP
kLNtKNgLXEHuJrP/4HFxKXatjQuy8ybHplQuEg0t6r0vpaSx4m2nVujwTZfJBVHM5QruTqah6eqN
4zvTQwfQpEDhh7zMCVhSXVoo6Xyden3VUmY/nohfGFYZ/eNX5fq6hqE+8WjSid3/hn0cdUC5Rhu9
XEIgk66Pra5ufp1scogIwkvYYnCZigKt8RA8DOT+ue1hLLcdgABKpQaRVY5vnwA++dwkY6KAfhjZ
Tl4zAJ/NhLHtbUGHGypO59eMe7oJoTRai++DvqmZhyomUrJbIvyYuC61bVuOBf1/WUW7S4XpKrNQ
NHHzAd8CMYmNtx/ZaEGHT81zYrqSOlGtRNLv707RQoNoRJxfNjNsKIpKqumKuNkmAqo2D4z+g8ue
6CtTzZ6H/7H3k8x8j8UUKDKOW7NWBZIgQomnYg3XeVUmbEPhE/Y+VNEZa6e4Iw8vXg9tXkxQ3OnU
0jut1vzVwLSGOk1C5QlP+R2jJTLIdEo4j3r0HDlHRLHQDovt22sL3QjpGlpfdnBjJsZoLq/Bv103
jwG2wtGUt0BVPr6zHUaNleONuTmyl46U8hyqdo+bZnQLDAG9i55jKLy6lxSKQMIUxaZyJCFrdYHW
YBTHTt2O1yJAYOYlsMvhGv5oTOJ57sAkfzI3mTApIZX/8hIN3T7y8d/0weT0e7AtlCjLT/ZfVf7m
/JNK0AKYSkSKFTYElC28Qx9Rtek01hLsrKrOA0E05dmObEwq+Vbgp8VXHX1yUEM9d8PUOOLzBl1A
HYip0yLid1sRfobRIoXsUPjgFqPNA9+9KRqdVxEP7nkiqwvH8moycEUySSJtD9jtT7UUS5lH+g/T
JZHgoFSpRtrTUO+SFH0xK+w9ksWZR5n8SUNs0YFRNZw/pw/FujqA6oSOFn5VkTOFB7j2nhjm3q/j
ja39+4G4NouYRDa0bfpYU1StFzSn9iKa65NfvDZ6nNEi8qBPl7Aznnsr2rDxvKxovnoooVlhNhow
ARDoxj8gqsZweWxmeAMgof1UFR//UC+Vr4GmQMsamV8EoatAn4WTmZkP2twWmHlCHv2WpI7EB0PP
RiYX6hNfaU9pNdMgx8e74aRIUGNc1IMy1DbcDcvUh9uTeSBAKP9rcCVi83y4s4DvmLuK96KhOFII
Lao9XRsWUtYUiXKF980bHHEKoExDP+YpbGkNm9eXHKu5dxSMivsyQlHVkGky67sdRdKcOZE3b/IY
0qqM4WlgChzRDigzOA0E8J54rXdrU6xS2cAP5tPmVQSRH7n/WPqIYUmA4dYk92/sZtfZ9VRBa9S6
/WNeh460VPwYuRCwwc7ITPqVrqqfWfMKxZtcHSvmNCxPkwSn1s9Yr4cKXY8cUKuZZjmtR+21ybRh
vg+CAuHhtDZbfV4jzGJ/25tn4D3lbSJia8elKIuCuh8HHqvqVyN+s8VJPAJDFqyEjDWfeDOuL1gr
wxgsCG9a2oAhUU3An/MSp3ZODc4lhF6O/4F1NjevhNqOpWqbEGPSpXVoJXLscVLzonDrNgw7LDkQ
NC61MJlGL5Az0K3UNj4RMoS+WoCssCJXE4Z9UWxcfQTeZGCCbY11tLCjs0vmCXkwYK9Zpc6oXop+
VHR8FZYJPrZ4ca+iJVdFR3GYzByF21PUalvS3Syk/1LFUa4eKFxbQSInYu6Yj0NIaIgt+914U5hh
6lvmcDyb64xuThb0vAVJWWGeAqHoR6tsVefrxW3GgeMRdORCi+ZWG9e/Jeq1rUF1uPpdK921d5Yb
goB2Abue+Dl2UypGN/6oFnPOij5OJ/9O/axgxmyxSq7yOdXR2jHIUn+lCktlDaziMaP4xZajb0Tz
/RkGH+vScMUv2RFaEnU6r9zmLNfLlNyhES4cT8XHEQ+cWQORxRQKBm2ahxEWVyubDcR4Mo5xsG1B
bT0yROzS3g31CcomqrqAoY4E36mv/yP2v4aNG5mekjrfels7dikdFDxbNXPQMdb0MJYiHBW7abHE
7UOzE5bqJDt/yQYcxGLc346fw6KxT5mBbGl3ahAUHCabGG1P+B75x98bxOwBPVQwgTcq0aZxZeyT
FcP6mBAcWvV1TEZ/AqyQlXOd+tr9pnoMj50fI1GfBNxacla6WNf0j+R9XRQWBbuTwQgpi5JIj/0Q
hM8E4yS/HIDdGk6D4f6cW9Zu/VN4MLi8z07lnXAiz+uPyoosgvpndzyUdwHyiRGUncPhU8mp8dzQ
qHW5ojAf8GbxbPy1Q3Q8hTqkk6DQdb4U5NF9ODdX/Z+5NDRWwOq4TJzXKLBqUw1X7F4xRU4mi7YI
gNxpgd07d+e14lHvNxQjkRVmAMJO886NnvCDEIoD2MqtanNPuohQT/uGira1dPzJKvL789E2ADMZ
luH6FMad7Uy1pyt4Wo0EwFQVkaxAxykhBwWDTHlreHPnLJSXC8pGTIS+e5XhpEC+Z+RciN8ItpQK
eHQ1z3jbhEynBuMzzhXaWlQ9eWtjT2CQO5mpZOMIGZKq9PMMN6a3x6Oq8wNqxeH19QGScGjrabPW
1YEt4i2Pr6NuRACZ9gnBXnjT5BqWsRmr1n73ujVcCWs/fb1sHLKKRsmnd21Mb2T0xftJRlLuYvcU
sMNWSWBXH2Lkar4KQEYoa5VpxF/tFZx+j6jrbgyV8PXxf/X4uLxTXwtPJ+dAEHvv5p2o/FLWn+fx
NEMNYXvupcT1igxKSdLAwwXgdr5OszAIJ/3AGT9MsPPrpAwJo+sB2Lppnd3S3dOi4LDMbYvcf6io
I3EUR3FMTm754ijD/DooHlSChXv8rmtpNTi+IVOItYYQL3e0ioZQ/flcEwDW1E/Ar9WNl/2ksU4V
SCqxQSPKHtSnKOEN0ZCIdKrTWtQYZpv8Kz3o58OguZ573X7g5c54eD5nJcmqVuP7ptoVT/9Zy/kS
YCyf0Z8xKrrMdpuNsohVf7/JtS/UNiH+xVEOCtVGB7Cf/GMTTa/ejKGTeEFukUHAPXPz387XNmFf
M/ERUYgPCRJ1hyhkAPVipL5pAbn96M1yGVmBgCIZbyv2J99+16z0/NElZ8OV4HOb0e0i42fQl+bG
9ttZGOX43GlIEDG9qEW+ekxYEWwnzh0IxQzDuvS42yfo4ku9ctVH3uP3/S7tWo45519b8Gr7M6NY
S6bZiG8MuWOQ0lVQU9TlxgRt/y8n+lM1C21CCbXlm1t741l05cRcAD64jqGj1tICMTFnwsFAfsqp
AplET+CokKDToKL7Z180g4qKDW6Q85M7m9mucqKtidlDS41lORSsh+cbGVgM+KC9/c1RtB6CCtU+
M8WE2gAOF/E+8gDShDT5BALDK1Nnu1XMExBMW6PW7NpcuuIOxCYFa3h+y2vbFx240SPAJwyVuSum
6khDfEYOhyOapT26GNCY8bGsleaFt6LhHUkNUaSgmOgEaIUAbAxDpnvfbHaR6W2U+RmHY+ht/fY8
PlDjK62wHFpDeoVbGqVLQDtnYmH8MxHFQmGa3IDl46pFP7OTBEJDQT28973c0NDT/mJ904Leq0C4
ykjQxchG6yS6RSntfJHyMCcbCmQdsV8hDbmQBGNEuNdw8Ggoj0gryJlKYMnqtoQILVuOSrvufLQP
8dG19ynPFqrcYk+CJu3/O7o9UokxohHiELNeTX7uyFL8vEzudvueUEFY9XEScJ61M9i5pfrRoRXs
76sHVg14cBp5sQTaNcsE27sinlh1jmSolOZ0jUcUHcOp+EU/9bJWRV+yv8Ztkc/XhoeVEKR4xC7k
pT3fxANXoCfs1WUHPx6NEbDwHMh3aD7Ft8GDLKgIlzmC6RBnMbX05OkKtzm+uVsT2+Ea/0hHdm/v
CE9UYI3cMNsyGU0iQewm/cfm/L4e/wDw8D691n6P1xKYuPidQbJ950IY6X4k43zOJUf4BSYg+C5A
EtjW0OHyJ9AwPXeg1uqxwloVpzTW5Bj10WrwxAzyGBGb/0Qs4aOFSd9gUFELXukIX8G/+egOgYTR
Hr7oh1XSkpU8MAknMJnRrs/2lqwxVfp+svoXDG01oFowSn6zRHiesDGub7Azx1/TWbHXtzSN/nvE
NDP7+rO9V1LH4SD5It25RGWtAuztwr9QJLPKL8AOaeWkax1YypQrbZG7SS6VmC+IqOEXTdWjiAJ7
AbSxjwzJVQ67JoKAZohTqSjNARSfW0/D1FHdLoHAfb+09z6KmeBAnh38/u5FdWG3U7jB5by6vDAB
jY/wBlJLlj6TzdiOy0KJfmoZCll0Fu6P3mvsezHaXTrtT/Jxlo0r4ouqUAbo0vh7Sg9A4SOrLsX/
rNQqu9SldvGIvtbfgRTL2PKv2LGO84KGlCz3cSdy2Okfathac4+JPVAywk8rhbOnGz0LU5XOQPWm
1uQZn48TOdWFNeU3l4ttjWq6KrpBVPkF6CW+Qkv+Cwg7fw5mivFMvGi13h8N2wsK1Rny0JYTbSH7
8xfcHFlm4I5uw+ODz2SMrluvf6xIh9oshBRSaS565pnoFPvUl1FQDcCTlQEWH2bbM4PeXzoQNg9x
cEiaNAt+FdSNFguXjWHs/+8nuw3nXwKjAHU96+LSxROaltNnClFBeJrvU1T974Eg3+5HqLRv+52n
3CZtd0MaNvKp3zmZPFtzW7YOuciIDPs90aoInmYZi5VfEE1WZg/atVaXdvMGgk/GhQphKJi+3HKI
fm5I/n4K1Ck4QFjAr2g+0Zsjfy0QgctfBciwQHoBo2Olg/nP2Emz5Jn5bHrIKsHCHjntCGfhvNU1
ML6CpXyjuctavCGmywI4qhhUpx0U4s8C/HOoW9ewXU2Judw1mUP9QB/ZbqeYc41Fiz2rfDIjVt9c
v0ENfFEjxGJ03ea++WMpoVX3NcYMLKSQoNJr2g88PfdderdvuhRHhrMrHTyJWm4fBZoRBLB9C6+I
cqkZm730hjeRyPJi9x/SxfAB8vUuD2R3L5lX7CUnWb6Gj8f+pzyJY/r0oAYTnJVvp8S1Z2fgxHnF
WTmx6o3VjM0D4vh/hb3l6wgEr4IKY1v0MkM3BqCrp1jUuTvhiwhtpjQHd1yJoyfrU0+yRup3Yk5t
rE4bTGxB8CEEBv7quMu9fpPHgmlH+KFWOY4gdm382ZzEfU02pBiCNql8b0N5oGyl+P9WY6wvHSy8
juJvWxeO+2JqY0J5T0pfa/FJ3xUNdLohqWiXyBesR7HwBzgOlYCCrMr2aIZcP8d5HwlZkov7D+tq
LNPo+k50JGLaD8rH2WMr2USZNupg+z2nZEsBz3CB4/pYq7H1COifCdaoLr83xxfOJuAqx8RjC4xF
uGpCDMeiLg38C0b+OxMS7TmfSuqP079auTxiDeQWXJTtbOSGd7Ln2E4a/716trOtUiUHqHvW/Bd1
/IHUhX1RV3eed3RS75gYt9D5sXqN8PVS3e5cnA6AV2+vMXmZKN4iKhmtKyw3iFeA+l+oORmJAnmf
PMeTpz5SyS4ZgDl260swsLFVjVfdecFR6ElVhNT+gI53b7lyNY/jbwfGKgOiNbS6H0BeMCybUiAt
pcwFjE7xUnAJcijuq5soBwyN7612hsQ58hArFyWEZTx4Rd1xtmU1ZZcaUgpFZG68y8dSMG5zUzFa
k27TcJLFQqpjMntAY0nS3o3OrNqK9HhcagHEvrE+XBYz6Kgs5r3Q4/Al94u8OOhjYE4B/xRG4Idy
TXKZwcDM3SPxk43gTAnCWx32ukjwHDi8b+ehWUtzgp+Vp4YEEpp3C74Qm+umQ23FGcpygSh2qQFs
2FKhumULPQ1bDEm4IvwwhfXIagF9S2HGoJ2ZhjmaYSAPOrABpzxi9Y6EdE+4kgGZxyLENmKrt5Mw
wExJIOd3pH8zhqbVFrAaw/1W+YS+dzUIrfsDEYaKORQXoJM6U03NXExt7Wo85uJ1Elcub2/JIFs/
8wTkBSZdkQ+Wq5O4dj2XmzVmpxxhKZaYaasp561S74ye5HBQMCKCfY+5WDB5o1Uc5/s8A4T4LdHJ
RSQxi/XZ7Ha0XQCdhzqtOocrbjwm7zxK+ZtmVE73vpCn15kBpbu/hC3b0uE/Q6gK+oQYj8+sL+v3
7AruxJN/mGh8iyYH3fMC0/ipg6nCt43VQYjymEp9zk6NxYY6fFBL2aKNVgFV2fH6UYzeRXn0jKM/
zaB8O1VIURhM5MbwalhvwGEZH1r2ofTcp8oLfmkkWmT16cTG1wXkRaLSkw5/W3aU7uZlpaDS4OQH
JvVE7PBJLvwafSc/C1xBFVQ8Q8GfpBngfRWdIs41YEYs8DQf7KLHdD9RA+NDX/QVc0Pn45uIt9df
en0/ldmyGtbrJpBQfTEbSZagR7CKqzwbIqgBx7hrBt659LOzdr2g6qTcqBbCdX0PYxsIyIIXPZYq
/AJ4yHEaIMfJvOEi3fcO2yg6pEHkBoQSMBagjBdUES4ZtZ4aoF5J2rwzNBzHAJwnKg/z6KFkrr7L
u2jsZAv6N4uTm3IcKJbVtTVZDGjFKH9Blf4qtvmxkTRd43XNuFoTgMPo17S7Z0kFR0Nyl+7F5l36
cJo8KKjqXCrIYaPAH9xquorN3ml43jb0f4PHYtPQBvnkH58v/OjXetzC/rgR3EZccg2N165axAj3
IKKTye6q5ygOYXTh5y3oGrEd1NQbdDN8cNEtrZQ88ozjsW08JYjkkVlI3hO2IPK5lKlUdyHv0mDD
JN+mBpTzYfzR5Y24SueRB+WwpHhEp9duw8rwNthdbyvEEPIylwQP60XmimHQ7cnnBkwYB6WK/2eN
HE/dUS/0mfpHHQ/+xnpPWMKF44WckdkV3s+ufxnXmak6jrF8kplHUwTWABFl0ptmHrQphrzGwDYT
wTfIhHUlHzAC5qyKEgUgjVkPeMXEpUa2Kf5tLFvw6Oqgcqv2Sj8JO5SI0C/G7+2OPnDlWXzzLuTk
7k8khDE2NaUMHhChg/YAf7tFWCxLTQr/fMESUwWj/cBlY5iAUJWsr4r6gy4srG0zotWVX+LMSTje
yxUv8Hbn/dNONGdOVapyRnmEJDOUczCO9XUzh3HcYgnu3q819WCrYfOCjc5LwzBi1Wguh0jg2KTT
Cx0YrKr7aQaTdbdZA2mo2s4wHFoPtoWP0B4CV+4RSWmQAO26Vu4TrxDN6oKXZae3xK9AhywfP/EX
lltXihrF7VvJ6wmL9mbcUPrF8JmnzkPp2NxYJRiHtmVe7nM/1P1xmGXfDpjwHqNZ/FXsDWYFH33r
h6bBxLx/ZrgAr8mlHkQVomx+sZctnXcO8AcT8Fy/Bfw/XrWvhVUNY/5SmvEywS7oYBNsLABb9fpN
JhD8N7jWMKEkvP+BBlk6cYKGHezz6gZlNykEedyeYzTERTsMgYJMl7rWqcKB9tdrmkYVeXNClpuP
+VuCqlcfds3qXmV1T56sLOUlkuptrQ6jmyBrptVpS2aaAcrJku/53TI9wbyQ0x5eTAqhgEswULXe
BJmm/P+RwbKnaal0fRar7LM7ixwpPGqeNKx3WRBo6OV0A6VRNvaGGYWgEtATx6c8IoUDx8ZblT1R
TQbi4iw5xKuLUkDwayrS9Mhib8U/CnfQW6L9xDKCNN/MTwMnysi54uCg8LiNqvxuDbBBBuuiKvRU
IbIOaDcuoO5diTTxpWC/o1q1wsr4oCrS78EChUl4Hbf5DYqk2xsC3PeJ9bjJDVykfCmdxtk7UJIV
MKKaPiw8kSEfunx13IMw6OYocqj/+deHh/S89wqq/qGtvw7m2J48iEhG4Pb48uybGvSo8w1w+fRx
Qoe0SUq4+9cw2U4s2o70EvaA7RQfRtuQgKMYY+kokQBJqi1QTaw3g0hB144zrnLfavXnB2hdtrbr
m8hBU+L43hvkBUETsPLg9eKj3hCatPD0/2YtX6l8gXLKc1Djpo1Z2AIHj5GJOv9Hysdll4Kd+EOl
JjjPren2gOlwVEHTdxk2ld6wiFH6F4XOVvB5AuLznfMPpWFLv2d5rgIBwTgNoMGqD+Cq9ljvLyxN
6dYHIyDtf4dq3AJAL4VvYrsPb3WHabEBXFctQP9vOuesHW4LqHr/5LW2zgtmRmpJS+pjDABk/HY8
s/paAvXADwXGGM/GS4IRxyvHHfp3CfcNLtcDGDuO5Nge6bTSSlefwgXzEw2yfvZtTmT+oTxxIvNI
e2TplZDW+caHCMyltnhI0hUculv7dfJw8fTplKA5xqmtAIAqsEQdjPdl3esOGnSmQa2ZzApSTnSF
7/Gx7Re/USZNM268deuQ70ZePRL8JMu5WvpHHA3Pz4TFP/tC1NiT62UwFCyoIpuEu/tA9y3XPxX+
G8EfRuJY4rppbHjwZQWCQh+5baxWXsy5RI7N7e06ExPKY3a/4DIMdxgOdKwCXpXcMUbFYevUE70N
Mm+rWTaUZeBbZ3AECVPU8i6/woyAv0SvR71JDjVucVonRyZX0EMI3CEYtoDY/jJoJQoGwKuX/UFm
TXfaEcapkNw6cfD6ifE9mWhNZeH5Sv+HPM46zymqiJMAaAH1wLs/yFbzYteGVbU9oEWxvHIQlILO
R5jcPlGyVM++nq83ym17i0th18/ANkSJkOWoWuSW4QLXZS+Mo7Th/MoRlE3ZhCXV19ycWi0K7haw
0SJ0y/jJcCn0QYYYgObm9n1htvWRj4V+Ob+YnOAb3nC9/HRf33vLLIfJ64FkLzeHo1EdnV91/E5u
vYEZNanDNoF6uf/FE4sV/bT3juEYw72GRBrUYrtE3x9pYIL1hKb6l78JqhRbwZBNy5SlG9O+TXWS
pEXTgE8tgisSlPnZrW2KgohbYYcNdL/tqvRNGHsvxaQwtQIYnR/zYvZCSiV4PWi0+I0g7tXEf2jw
JKYa3CkqUE4cOEcUYbrJtFxzEXaxszwHGxhQVaeWsvaSAggrTPSXOHXnMZePXgV/CLcKeQ0wThyh
+xcT8+dQipImUkOH00Z8wEati5xnhk/KL+KvB8OTLFLc8yKlfAAEm0vjknmmxDEHkRsNEGTtT9jp
SMp7s1dUPrJOJF2h8RwLLF3tnHQsNLXl1IrFfHH4Wp75ALoyKV/A/oqnHAwBqWkHpWx8AEnYQDcv
4Su64A1RJ2D4wraJjfd1xQh99kbbcqsK8SjpgfKuU3/t0LYbVFZP/4Y9zsE0lEiXVUP9VJIzLgZK
8xmdQMcAg2YelFT/9Rduoxuuj7O81+v4WpVo2CfJP1KBgSv6FkYiFRe6VzOVSYaTluuTA8OLtu/P
pr9jHN+YGc+XqAzF5GihyTxj//Wy4m2CBnhtHJKwewdHdRd0C7mXkdPuheFGW89tQdt2Jc854hE4
4OERtoi7iC1qH7E38aapXYcEx97gJlMKLKf7D0JTPNLfrgtAE31DlTb0wwhM5u5IeeHFplcvZCAP
TUOZ8b9V9whtAmFvkEz7645zFCY31tJTBZniQSku2odbIdOFxMRxQCOAqf/PYAr3K/lxKWZx2VTd
7qdNMrujVVRBpPWbwHRaclgq5ON82ZlG0ZXPNboPu5nBM7j0N8yyHBnsCxN9s6JcjGC32bNoMIy4
Fq7IIu5aD4CZvy5ZrwiawuRyiSIojAocM2U/4eNTciymbZkD2s7YhPAiQ5+1g8WVgi18pDlsBiM3
JAQIjGuQowShN4BtuHEvJI7g1BhKRNMkyw2p1AaTvaQGN4l0Wrg4MXBzFQudbdQamIv4mhv+k8kZ
UbjJK6UPvcsjzE4XhREDNYPlr7czx6qgtOItM4m6Wb+LNICnzezviCG+8YbL/C0OmzZkmryRWiRe
3iLqibXpOoKWKdif0Pnk+pBgqjfpZ7GwfE+B+cG4LYcUEpM+HkCkdjPP3BU/4Sr87oSuHenYNGm1
8qlshy3EGuibxLta0zW+NweGXUffPsHcURrBvvE4qy8UDujUfg1A8UfD2WlYwfM+bsPyD1GyOOnv
L7Q+w96Z7tpZ6RrduU0fJWFIdxI4nb4HE2MpVgEMm6A4JBGRrw0Bo9/I8MyhTkKESyYEcdljELCy
Wq+CZ2CTuhhfDFPS4ZDJhI6hOed7oD4/PRT6ICGutakB//OmcFbST54Mzp63TFiNYTilziNmef0g
fxGDS96yyQzLJNIpBzqYddTQiXd9gqeu1uYbuadk6Oq1YOz70dAleV5dKej90sJUyWBiEXn0pWrQ
0H8hQqj1FgvbVgGpUivbsq+izMXmX9V/ZA+d/Wwz7MWUJt9T92EJPJD/zh7h9PLLUPv61CdCytEN
Y7PNwgoaalzgyyPA7Zp0GlsOwBY2NK64U/rya0NULENUFnJ6EqbqID5YZC6gKO8wxNzCw1OVFwj/
fnp1eECbBBnbrixNR/KPb/I56pqhcPGtsGGXrkRX6Z/tTK9vDezKBzSBKb6IQCALJMIRrVe5v2oe
CW9zfOCURgv2z+7wRWqn6iWDuoM8zrsZXhb31cbKp/nDnIQb4cLE3ULMhz3Ephi9bCsy8hkbGU3k
rFzGBgdog/YSTXURfM8hginUMjXKyVmlYbNM6buAepLL0vSVyjvF8q/DbUlE+CHaUYrH3IHnDvRW
OFFjzDKMAMtKQG8wp+amwSZNxs2KRiGnxiG0pNjqv+o8B8DQLJOlgQq7uqDG54SAYGJlsREWMLcm
ijIIol4DYSuRM0phA+97H4RC0cm4nsMC+9gChpmxs8YU1kbe08Jrj6txJXVgNcayzb+EnNU8GZmY
KVj7GLgRvByzF5gAdhRdIpi8IxY5ZDWoRrNbGj3cmmqnTK42Dr09gh9yKU8qs8d3cKC0u2wsyIOi
u6CNC2jK8HzykZlhbJ2Ql9jc1yD86C0UaZHhj+9fUY/xVnWgh9Tp1OLBijdOvHcFYlTvhGKNfGGO
S/0yx7BuZq9B0gwrXqKVjBNeui2F2UISVcxneCbvhWyiDIiYIQmdi44oJWAXuUYxphzmEi9gEAA7
CpjgJBcbwvpMRsoTv+7jLy5xULRerlJn2XA+3pIMta9xLWuQQRxchOllIDLDRjN6lbLFB1V5e/Uf
Y+baVV0C3Gjke3Ub01kbRLmAPTVoociDq0UCDopyPZg8KzdgugWiYKLOIYpRcsgWExL7t7LP+Sry
0ZkxdAcm7bDnD/Dd+TpWY2eFFF9HWr9TAdORLTbvBvsu2wC5OFun3/ZcAY9mFVHwJrU2iJ/YG3Pb
By5T4njFyiYGe3nb9Be5oyUxXvsc3CHTz//2CJpt70sYwR/3ut7Y5Je/4ihxW48LjWfg93+gCCuE
M789yO0L4TSAOUx7E11P9+o6GFiL2VbNBxACvPoAjjKP6uJtVNcThFCajEein7JBRvKTgVGlMJRo
dbwXor02mTFWNvaDLQODo8R1nGA6ji6M7GuF3IxvYRYY+a5bnvU5q2rezwdCQ7jqfPekhZrE0G7K
r4Ep5PC4jrGTGiaZJLGo+1dTARJBgwQlkp+bh3XtamLqLp+Uy1WTKC6wU+CKbKneJ3c8Wgsh5YAE
4DGnE9QEwi3/VF9aO/sdM33tdh0S86CdvzYSyaBfcEqJ6uIIAGJPvc9QT+c000hYxqmMcPUkluXc
KSU6oyMJznslz+RJYuhNjIOQubY+Y3OZHXXyhAGz21ORMf+k9FIdB9hJHx9w7ijTk6pre1p1zcRX
6B55iahbVCZS8ukRFWhVgv/oZdfhB7xFBLVRK6dOp/piFwU74vKbTH+fMyELyNVc0U2LRXSWvR8g
MtXrH6/KqShfJ58cBrTAlutv5hxN/gGcivACEcRjKXxMbadv/bBMuY9PhddTTMlZaEudsreyW1Mu
dYQURZIJAlFuhKwLNiEOADH2RSD4kXbeChj8lEHhACqgKKJSvy9ECLtPF1zTEQo08WfwnC26wIwx
AQyGpnrFp14YJKZE/ZwyVNKQhLxKev+GaEBzGcjOOz9WXI+3mVLH3tQzseBAnmjFcb/ih1g9U3BM
7+ejpl5Z69zzLi5+w4v24J9gPF/+VkVNCPNah814UyESf4+t2CPYOF1JFbp+4PZHjh5an9LCG+Xs
z1GuPtToR0ZXV5kpmh4oLYL8ll/Qv1yuiFzjKkRwuMFzUquqIN3BP6x2WWSxF3E3EThZDUNZEmu0
BJmx2CzEeEYjl4f+dMRes4Z9ieGS27GVyqZ6yAmaknNB/O3Mj3o64e/lVXRrIPrEWwXv5r4QMoZY
S5dMUdkXFq2HS+Wc3BGqGRUYxt9ys5WBeUgv8AGFNBKTmWS1njGBcfw7FjQVSsQbEJN3FixNXy0L
uVf0y1UcCcNH8/2cSH3unb+vz5f8uDRAXIPNqPpjvLvhEaulY8cdb8xYF0iIKao4/YNg95FsN6uB
0vKO2mPSgaqhwEJi4MF024T8Oy8+g3E+EPw6IYa4EbComYwrkfUxSOiWdgJRrOx2eXJY+Twwtgcz
yIt47h656y9ZgB2sABNMAQP3/pKuzg6W8c8KSn5Djz6blg9V5mTeEzcxB0XwoPk9+ECDIwFp/38O
l+1SGAiNXK1b3Rf2R+jWnv8W/HYkvfEl1CFWG6YlRXGIxt4O9bs3NXbNXa9V2T7+TVxo/0q5gzL6
7Do37P6/iLhR0JhZt7DEYTM4BUp1WKiz7eXRDNrIa7MCPdtpfFKYcCtdez+vVSJUSSzy0Ucci1K8
JGaKVa/UZVbGeeuoXY3mf5Cp8tUnzC/MkSBc/QP0+1S8jP9IGGQ47H0AMhs6YzlOQFFLjopsi6N+
llRIUc/tqa74y0cixSxBOW3/QakSEHN+cqdYVNuO3Z2QHOoNB4NAWW+s9C0UbgS2CUXfRkk9dnPF
SIl2C6/zH/LWqllBWzP7I48ByAsaUW30Kz6cHSFWRTrJLN7ARY1kmYLuzJv96fRtonL9yZ0Y1Am/
trnLCrdLWHwc31+OqUJuWT4Yqg0fngkjE7Uh0IXuIU34wVNiKSPFiCB943ixaknr+OwgQWCaPxrD
kx7Y3dA6SOD4xTewST8zL0zQv8my8Lz30+XOjrvyyNA6PpWfjev4g84k4AhLSnOaUxyzVEpntbfi
6zejmokttFOba6SEheFiMMwO6xNc5NJYnXEk/acaI72Or3BScdYVjNoi+DJgjocFi5G/XyYq9fPL
5a8+Umwnm8kOuwEjZandDi3U6IgHnhRPykP4c1HnljKOOTXinsiJ8gQAMejJMlX+w5Nc/HlMe6Gv
atLYNfROI/s2lJXpPLelfq8NCcTHna9u/YUCVpvZKUS0ilKQMX5HMXujwG/UhgjknL1I4bb0SKpl
zertF7HXGC4kDsCJc7APoUq6xoi29jHThZ8x1aWbWLQL0QExt6UGsbVQHz57E6n6pnpFBvXSIJuc
C7e6KaXBhqZosl3HwSOIT0PHamD72gpK45HesAv4aQchhEWrBB6mTQxh7O40X+mBfE7PoGqea9cP
W0LlMXqa2BsbW5/tl20u/VnK4FI1lJq99wF+2cEgnNn2L0dDsn8SCKet4jcEE2HBI9aNkpwpqSNX
d1MIN92LPZBk0KFdyK2ZrBl6v7QjN3JtDCCq3xwoBQMVKcJRNpcPPokAUoVBr28fili9LItDHZWq
MenoVBITPpvmX9XoMJnKK2md+62qQskKNDaqAgx4rj2erc32BIgweGSkpALVF4QoEhlRQ/ITcaBw
DP1O5vUpFS7mIBMnazKqYqff6MlERS+JZS9mfsTosRmvxz8OsM9R1tHF5qisVchXmrI7ofZbM6er
5uIw2n37H/SopaK+Pcjm8cVC9xqJdNOm06EHXwF7RwX4oO865tJ8Q5ymz0bf0t9zRNNOOeOxSLBv
DeEcEk5cbRd08ZSDarGAyJSYXLnhP0BvZLfD6PDtV13reVWaT5QRWOvoWLHarXtc+q6QGgRS0Bem
4XdwnQ0D4gsAENiZXK5qrPj8ulpti463XK1854EFqD4XMdJ5UtTbIv5M5rKFQlxSJW8hI9ndY1YD
WkIFUzrnMzBgb4I/0Z3/8fX2IDnF+jgSd1l+y8OIBP5wiXBVGYqfFXy3U7OUhUsbxh+rBhjyuuH/
rTPdQY9TUgOS3gjFeKUXQD2aT1EnKGv8i8vLIwXaTVLv5yV4hJPkXIAPON9nVsmjtOMyLUJGE9nE
TViuWjnzG8P+1lzhRt7Kbt4/bn2gINyumdWUclsX7tG7STcoH8kq2tiVMLVE3Srnz6l0g33x1sav
a9tD4xKCuq2D5RpZziDH7J6hPS9PD0vIBypZhLLqufU9jKe68DqcLXPtKOc7YR2luZNICYBt+Jvi
wXlFdZXMKK2mfoDbWq0TR9yF2ch5fja9FTwUqIK9xYTaQJ3tcv5HZzYS3AKEpSYFhNZSjrGtLvlD
kkev+ot920QHtVKsTPXZGjJLucy8aPYryTSm4qMTY+8tKxGdNi2fwVfKUrBalVwwDcyXgBcFCubU
RtEUGx4HPUarHSyrLSXa4qnhh1l7FZ0h5c19xRB91ZCv+h77UR01TpT7K9eiVhhcy28tBjqnC79W
R3t5lkDeLksZsllccMbqtqfJVslrAOnuDHbT6PUfapWu1mFMU8PTRxdrReUs5ltGbbQKlGGLdGGD
VymlihaXlXvjCoTj38YHtd3jHz+145hTF9aOVJi/xIdBuonoH9DB9q/vRTYX5jabu1EUe4KYCbki
SS2cjqtZHmyG1jR4YIZK8TRCeIIcoZaBr05iWsikrK6ajt0L0dqhEALXPc7Jze7VbHoAdAOBgU9R
RM0kamit7plGnE9Z6B+PAjFgkRkbPnyR831zwUgFT52LhBhaehxI/QCnMDtXbmg2oK2wMT7uwiAN
7nz5P1fG6HJaKrdr6boomiXiviFvvP0JMeZGJ+u8HsSFOyeYIPAItLWJSy8Kj53B9JTfFaLr3r5J
Belxu5MCPODDD9JJZYaDieZ9ErxUQ4+7cM2lsWWR/iVxla/cnH8rOKrfWFdyBSfGYelSjXxGWbm7
EeW6lMBLII0UqOpVPadjHILwp5FYWe4JEzHwfVxqDjzdHQHCe9x08qSPv/eYTQsbvgJIe7hC1OfF
TW8rVFpzKymjOd8SpIKSKhZF6hmlVHBt3Z3XugH4KiSJlJf1HvrFFhdb4R/Ll4LgfzVC6xclL8xo
fl1CcFTVsVEkNQ/Klt7gp0E7apdDdTrgYjsNxqSINjM3s6ZqEQ8R+9ZIpeRdLmHIoSAHK9YfiPea
ODPGxEOHbfRa1vHQpFBbmS3qFubph0GpTBIeOPQKY/J+BNHdmJpy+eZHRhcnDXZVbL90atbpHjOL
dFVguXg/bu3fXXGr1lY9joRFyrDTkeDEbPMCYdKbhjrIja5pHSYMZZW4IUXV8xvbGpZScoQ6fPyu
v4/XAjk/wFUCaolcw0MxCZxcG245PqxMDLmIWQnaxAbO90ZghyWP6h+qmHahhO0LepJ7MHB79Uc4
Gzv7JAMeuuhFhqnNlUd+15WYE5WJr7fxlM/GX3cLRG2x68U3tPwuNWsaEfcwAhnV3Iu3JbK3nEn1
2D3xWawI4rFHdz8oPXbxhobgQfsaQXA529eHeBMF4RxoYcJGs3Rf5BROLp41YwmpHDubBA/P6mdm
sBf1202ombDVUe2spxMATUlYOazN+1YhEfTIhHk2ns9UO6Z0T9Z+CcDxKCBxbCwAa7wx+uB+twAV
YvJsLEEvXdoyJeiaSILihbXyRpckSGKrg0ZNdvj//X67EGBHb5UrgwsDloCrn7Q55Tj+6+AJ/QcG
Ngfi5UP4GLwsLtUwmbPn9CXIyMOikxmQPZeZQDrBiclqJPn3A74h7ZBfh2kPEGF+TAg5GSFPGBRo
fLA6akcMGtSIXUM8Mgg/gdCzR65nP1olvC6AAZP8pwpaqisR3hl8G0dhbKcJHu/PKHCpXon5CEKe
unY6m82UxUSuZStzjWWJEAeuSFCjDXCRPdXET7ExoqAlrpZalZjBqbjXoLqlozbulwEErGcfQC2d
24SiMSkKqTDY8sqSH5HnrjSV3w2m9DCNiVI8xa4pj5B2LKB8BjIUqCn6EuTDhaJYrqFsAyoqb+Hy
T0acad2VTGzV89Qf+eMvkZi0V4MurdRBCOW1zyiaD4Lc93S3caReGJJbBs61fwrXKV6/bggGbgSF
EaVp/rO9RWADzgaBI71v8a6IeIdtDP5i4NE2oiNQMKaipZ0Uu9/5DO8ToEzZ4Zgrcn354adeo77J
v26RFwh24IHuBrh5jahFe/yWYRM2UuWTyTBLKvdUfmR5cqO316fuwOeamx4zRwpad/wk6y1OpzYL
D8c3bqP8EjRTa/dfs1iBNEqKkwbpvA5vnfX70LwVhz4CB9Iyfm+/CYxJGncDNWPcwV70qM91mhfp
pcPIgaLL/CczieosnhXSo9SHVljd9h8AxYQzRZ2Q7U00Poc5XYjxh30ZAC48jNxKDFi4P7+rj3Ny
2opT+6OV8jcWkCWtFmMljmoFzEwtuxjZIXVvX1pEvrTeQHGRwILHbWkoOXQ08f1pOiNk5jXm9Gv5
ei+oCMIYtKNFWaz7VvWlgEFasV47bX8kNNEUMou2ckLovfLMLnpNIP4qkkgdBNtpLl8d52wXuibg
wJpB9sgEXfPGB26sipYT0KRIc49chVibez+hdZRpIQAsxUcms8IBxZT4GZY6OiUp1PDqLswigvwW
FTkRN/tWOgylcw0pqtbEMzGhdEGtK7j+hLtGLdXRUslluLwkQGtB6R7sA0FOfoFMzlBKfwJ/w5jy
PGTMbqMAC3LmZsmkMhmZXV+QO5XBPnYbZHxPughTYF1JXzMgYRsK2euOD5ltjfBpgf5YGw9nwKo/
TzlVngyriPYhodRvIt+BYX7fyWBhzISlCLNe8+ZUJb/Bftdix/GRFoIq5nD/RDJfk6Blek/SWIKn
Lze8yGr6g1y9fTm7hQB48ajaUMDcdHKr1g0UAr3xBnUN5htsClLni/LAaJ5tDwZvUvMSCwTcXyMk
xhE5c5jo9Wj0Wqg5vX/SYaMAZRx2m5bTipxakTN5z3rPMvzghAQgoIaWDxtTzEO9Ux4R2ZJO5nPN
3cPZ2+iUj8P6WC5q2uqABJCdlzOS056qWuK10Y4qycDnb1LkTawZX4MgwPqHhRoRdCPP/quVBCmp
omox4rM0T3uPW/loVJwg3kB32tJGP/MBPFHmOH7vMojajcbUWNWtNC3ygCFfugM3U4vI9j3PavFy
MOj7xywmURWsUTDvRCIZaL3qtXpolzRiDgiaFbcm2KjupWt3PUlo5nD1Wh7l6WYaTXpYwJM27NFA
1QiI4aIX80YBBlS/zFGqRcIBCqZLBGX22AGtqQeJm9AqpDgkHWLyDfE+6mhQs+VdKdbgyNyyr3ba
r90313sc3TMyUYPRee76PYrWUIjtSzoo9yua0Gd6ycwA8EXZg8iRM0nTs/GUHMzluS0CgVcwQZkB
pkYaSe/TRKx/CvM9g+mGnHiyyi2/8YUisYpS/S5z/fs1iAOOjrX/JNe8GnH+/FFHvCyHgBjioaMw
ED/9ckyGzx4xYXh4Joww4oydtDRmo0ylwgG+UK43GOW/jYouH53omaByhzX4w50TvnGIgZC2hyD/
6YKgVpK6isEtzPd8iQFqmkHYL8RIot/MSu2bHMNLDN6JoOPz62XhS3+XwHxrnH0quwa8jhAimaG3
EQoovC31UucwwfiURd1Xrp8c6ZBIglww+Awj19b2IkXeYYMTw68pSUTImy1Sb+k6miv7anTxNbqc
sr2I5fKGD0qGIyA4jRNPvMOVi2qaT1oazDeZWrULEyf4jkxiH0lv9l44IFFaZDtbEkxdINUtAJen
Mp8/ms6MW2USEYC58YeiJa7PIX3WQ10AIs0IAan3Qt9QjVkl1tzfrG10/bKxOdkaS0F003cCaJI1
Q0nrSWSVQXyk736GlFEC7BMy1RAfcjFi70WO7XOsh8B1XsH1H2AwAnnD8Ym7eUL5s/5hMQ+AIjb/
i0uzdcAr/Xyp7B57jeWMKkxvhFBbGSzsJZpWXXTPt1zmLpo1QAxYkMGT/zZRwl6KcnFB7LVkcu2a
VOfoM7FBCv/BVqrSlW/7Ne7bpSLvKEXEowwzLNF9yHnjlG0l6SBYRdruf73r208sak4AzUZiwVJE
wKT3B3fZ1yssJnZ23/SfWMQKM9k4QzMZIG1jjLMDo2CQmRzU2UJdDScuq124XZwspQhdYlxB2n6+
rPe+xw3Dd1WezZdPdZ5YpJO3NY19gQe2ybb14nx8TYAJfCl2uJ/l1aMDQDoAyf0H8HRCSIDJSP1O
2coznSYPfTdeD2Pda0sszOpZViyk9ZUJZV7/KxJ+TE0rXXADAtS1aXpFSAaHDdRaBfb8fifx0Wbp
fUEQZXh9wluFcIUgJJwmRUFR13VSDjumcJD9viP3CIVFsKUOYEN1Oc3fVb4ftUKQ5wt1S/PP8DUU
Fy9FKBbmAu65kwR+ILXDuhcgaK2sDUMMrTgdmKE9U4CTHqGL6OcDyBowzD3frD3aeRFwFbJtqtg2
ZYGnikJGbUTGt43bM8B5XAEKsNtECj7dmaoqUg8ETZKRdrOlra1ORU+xRg8Wfg5ycdmFokaR1WPI
/tCNunu6NV5SVIULb8FifPkDFkrDA82Y5sGZ3mCeFT1aLpTg0jKqcOmEP9iqxbOwB6/gFkM7CreJ
WJT89Jj61/DftrWMIwiCzIXD7aQHqwV4ghTcXFuoz4MkhpjJQob/TnFepEQU3lQEnnois7YxO4AL
rjLstF5eQ5piKAF8ZhR8gQdM2hSVLG/j+Fj0+J2x3t4vfdHl9b6/QZxs34N1xGbWGR3VI1o4oznQ
sZI80cHBUH78PlljbPlnn/Zjs99xFYeJjLyohmVyJ0jyXC/ddTmG9teNxVNLf9wEAFPvV0aqUAiL
muxaUxqsVYYDSTiJ1KNJYN+/d+Zv4TDyTYh8ncd2yM52UsEEJZa6UlNP+UtQq87CctJ/Ih92RfvX
2k+rUFcCU1ZWDWt8efmj0fxh94cUf0W2PWIbTd+75IhONjx9NFM2eCbsfVV7ZGkQXY5j8FlTyA3C
ptSis+h1nfRJR+ax6rtJ+5z24mYF4SrYtJrvmvwHhlsgjw5XqgmVW09dSRIRHTkRgtp8dlNHup8e
dcixt/Rx9/AFgeEWQeG9zLtFHQPZR62d15k6lu7yncr5BqsTU6nhgtIlIZDbeVQyipWNNpbnXsT/
flBFd1dFRpnz7DG0iu+J+8b0/mvFnpPRiQI+FGlyQutKi/uUERHioyfB8ZFRemjn90MdQmuqJoBW
vwTmIZp5WOOTllLnIzF2YOJB91YOsP6/pSuaaiXz4hRl8P5Mp+cgLwi+s2Hnzv4rWczh2IhbI0WR
oSA4lfrLaNUFFuFUUREWIRcDuiVGryr3a/imWKpbQe7pMEprxAqym4IjrcE8TvohcZtSzE0QWVqO
L62nGvo2tphtN8Byy1wAdFYIPZ5+xFmm/4oQ7p2H5h2RKQTIczkgMNhpU/87gbQeKDK1kicaaEqK
olPJ9uRrQbqMk0ZKTbcgeRzNNYBxfx8AQ9iZiKaxPHC6U9PnuijpaTRPyOXfCGAbsYVw++TBwXXh
DTvuUWOmXBWorOIp/5QobzjiLhkmGU9zdMnTCmGoTvZde7a09ueobDHQTncf89YTXKYR9p72WIBW
zs1yLWuzMtJZ6pFQY5KrDZyEZTWRtmSdi+vdjV0FJzMWyMrbsWrjSnQP9HqCq+311nZRvAok9iVy
jRpUs3t09SJv9Gyw3Wk5pzcX39HDIoKtX1OfdJJwoOgt88gOqh0oekNcKOjlKUjyhvONMCsmR0St
F3UuslOWy8vnuwCNFKUACkVIA175z0wUJpdmIbG6YU2fiPk5rDlUUopckZiUScyCZwqhlAcKdYLr
xXe9ADrLUZIFPxh21DaYPlA0piV4Rk7qEWV5g433wGAjkhzN6uqDdctA9Q7WbgaTf1P2fHnIdns5
aJ/qKqYZj/LejfygDdeOod9yHU7ggTLtYx/atmGd6q20Ss7Dw0XgP+N3TnVnJLi5q2Sl9ZYo+93o
mNyFs+HIbapYl3x/OCZS6hhxVSrVKUx6824lR8DbISQsJPRQxSuY1SRia6IeywjVfN56UICNnizD
8yUyc47+nuZ4yhvP4uYWcyIcw5eb+USQ7QAbGYmrStuHbDWF0mEebhibloXISvnFt7GDzZN3Ud1l
QPzAGbd89fp2ZZk/+GzVC1HwkLaMmkIBxlNVKpWQwBZcKVGPaKytdeQJUdn0XYOEHzFb4XWKqbcM
3jnkG4+ywIQ7jtavBaTU5SBwoc7MJN/6iZS6jfojNb7e7Qt0c4+HDGQQj9tZgopa1fOxuQQIST4f
YZTrc/CXqfJw7j50nGk/bErFzZZMC5xeN0n9yCGTHZ+QVVIY+vBO5dYuP3MJ0ttL4lVfRrO30Nls
Hg3SxcOytg09t+42DlkLYEe8N1vAq2SAEvflKFjYo72ICU6bUJOGYTfYLHM/FZ5WV0e9AqCuFMsz
ztKkIwd00mfOFT4f7X9bLEUdnk5Tq2OhU1InLI0iwyDLwXxO6VlY8iLfgqkyEFZIKEWdJqrP3rUN
faGL2p0AE/cD3QOpoNORWsG2+iYh1crsapWnhO77Z/cGpsGvJ/hI8UtusPbpasqHz/O7HR2NuTgg
TXXKcc+WTOeDmOVeAL4F+uWv4Ige0L4U3eXBpDeWmDu1boUC/GPC5NATiDVPz8BB440Xvt9p/nHd
KQKf0wIlfRlZyaCoRq07ju1PM3yciJ9IOaCdP/RaUpa98X73QQl5t8eEdLK7NzDsPwq0fhJtLQPm
3wlTeb8ot/mWBf01n2Zouf1mnJ9kNcZEKUBgnCLoOI1fGuCiCD+Y19ooyLE3zNEmJFC/DT0wGQHg
tazROmJe/o25+J+JvGiIzoNC6Qjxoj0MUxtJuObMaS73rKsqd683xakLnaMlPptqkWJ2BisdxpJi
OT2tOFViOMmJHycZaK7rcHqdp16ePJQNPFrj3j4uCCq2Tq/iojBFPQZepKyx8etXHhuu0PfXcd28
RyhaSt5OkCgHvOvZuCe4PH28UJVR/9N6ZbMyHRghjsDycmjDkAqxUGaJJ7wPAfi52tRpH6La9B9U
zDJHUzjB90MTIZqtA5P9RmnwqNeg+TkDM+Lqi51zloLN92qlXdNMGJSIRERCoMBHzcyhkHjXffIu
Ao0cS2pefHhZoH7VWXbajAMJYf7YwXH1UoA2RZYPJnXkxovoE3LCQFZ2gKPRBDsdsJPtKpFZYAeV
TYGEDQfjYT0og9Rh88K8vxFMo7EbYSuEbhqw+fZHropomWhjZDDEjxdAQxBNAdqvl9N0i+KwuuAz
CBclgcffqLaY+0NHNriYvl0SpSoT11mmWjuB6SZkNPtcIvyP6gBNpe7Qpq7rmZji52CZ0dem31ze
BQCym4Nnz3kfY4eMOGTQrRb8yg+lwTAve+9eSfiaQNZ5wDtktne9G1zWiW8bPDQzTu1ytbI2uuVq
VXyt+m6MsAjg+Q0VlEI+dkitgPK1IvLUpofBKvFgS0K/UFM4fo1oolvSpc3NozZZxmlORUKaNhSg
a7ay4H+EPnrusQzZ3KmuPu70hWy9m27XfO2A5VW9IzKjaVz3DLc2odBKmm5ATdsHUT+Zt+4z9m+f
fd06bzt/DGPCkbU8jf0CbEkODkNLDk6bL6NKP3Av8xaz6BzpaJ9gFekjkpplemOgHvlMQTIB21A2
GDV6SZRdvNMRuVbeWPmtD7Xa8EEajpO/WBhN58WyTcEsNEV5zLPzxuMsmnuC4GrxqEGnw4VmHnWg
E7xW1OiQ3SYWcO5RI1dEh7LmZk62VBdE0IiQmrOdRPBKuIkz6oOT34occOaDcHpzEiYfFtxS+Le2
FJfmlgVA0QoWz7rfAzepn+/v0ifqCrcnncKq1Ya5v+BnHYGk7zxFN3igCjp79NR+JVOclxejgljc
27iOXpyRiZobOT415O9muIMPQNKW0qKo4AGwm8vXaWEil8ErUc09IJx+z/pSNgbLGcoieXDw60Va
SPFdLc3OZ7Z/XFIjDrhGEYSIE5UQU8sO9OlHo7MqW9h3j/WjJyqXVgAENPOxWfxnZKtfNJTVnBha
i31HZsFxqiqxprtfTQHczaifWdXHjt/SWHOgmb1Mul4Je9a3fAz8yk8TnLlUTgZJhs1U69s9B2uL
zC70cv+EFFn5zZ/HVg3doWFb0PEjT7eY04BA+526lw33HtXYSXJviqfTZxJru5Ne/a1fgN+ka7nX
405Z2P+HQhkoq2Q+8Cp2ffcrPTYKUapdVCfRIjP0tnvHTh5P/iEFc4Ow4MjGXAw6acqMY0dZzekz
rdTclaVd50EjdeNkcYNar3uhX1Hb9FdGNnDOzIAB2WlajGaoid5onpf4/8aBeO+WH3J+pyVT1sMX
S5AJW+tJGLK0BzLXI7Jk6OyS8lsq4FcVvWuaKorBUevfLlGyuFwitBrINm10yXl2EKQ4BnJ4K/wC
0Rcj2ZRiX6A/xxEItoc1KwPluYSfLQl5BYjEAcmW//8x5QmZeH6n4mpGSX7SAw2QTAdno2JxrTgR
MsbVHmOlDEwwSjWSqPS0gApcA+A9smocD3NIo4jSOAGo5xYpMoMYgDkrhWXbzkLlp8px1oZ43e52
EW5CSnTfczD+xfZzUqtcXA627oPjwOlWmHmDm0yrQ1qSeV217EoyzArw7a4sgSCRdS2I8lSwJXHf
pjBWc4BsAx4KuQpLZJdfcqYyt2H31kO6AeshcRqLuOrgi39wReeH9XKd/zU6mDtHEBzUzjRuuLTx
F1PK/tUY7liW7qz767T45HJ64EOcb1trdw+z2kLMAXmLh+tmVVF0TjhFPsOIh/2ZpS1iOV1TTxeP
AwTXmZV9fwOySvb+/gxsvSK5Gst/uSARYVv5DuaBTQgSMx4fzH71DBbzw4fVt7B0ZJIPAmp3jaaf
p5NZcDx7923FBfMAA9TUnnzuaGKBrTrNWEu4xKxCkuyLwb7tIgg54G/cV7kKuuTbXvRFaq8dG60a
tYCEg0oLET72eF9P2A8PUThLYDgeTJhX93L4YaLLVvbquLmofkOARU/tyDn5ByW3LWE2qxA0GcRa
TJStUxfVDz/PSO5Tn9AcvdjvTuNMtaRgjdMU0PG1N/YY/GKrfVFx7z06OR7j1JQBf/dSog/AwGV/
cnOweeLF4kKJqjmyoqwmTDYw8w2dAcoZazQYGrlTK4P95I3wd/LyaaqUQH5npCwlA803DwDXlVjC
w/El+i1EyqX6OeQzwKcsHNyhDxO4U6OZaW5eMV3xQ4GL6sB8Qj8f3vKByl7O5VoY7QAP7EDusSfT
gjaJIkhf70i6du1+ZSnaMOR4Fuisa5zEXOVJBZ99bWjWKlQebBCmgTsOX49BydyROt3FbjKydZqn
SyPkAISb3uCpbuYbv9D9pxFIIly+3HU5xSQCHfncD1yOCGtIxOjUhSpgVotjlAKSGwpzUojGdC6m
tqPf9dFluLByRzT3ccQBg5HaUxm83C1H+zMLqu8D3aVeh3nHWaSL/aVrwDAquS6WBvLmps8LwiKB
79bRzo9fwy6XmEKSWgx/pPVAOxk/yv6tVXlLjj1R2AQb6p+mRIo5aaVN4Z+v7hWWeY3DO70RRM0P
L9Tg+Y1/+Za5soKAGNZHM8ifuPA0aMs6CEv0oP+B4sv8PuCvqogFYoI6ZFSOrsb1CI4RrsCkN1p6
6St9/qoN82nkpfcCSq7QDZMUpq+YgNKnqieolAVkBFO11azcIBVhHSQoFTTryPKYAuDZUTACyfaN
2EmbXLzF2AUT6ErUodZTZ6wvrcoOsqObriTTA32MZF+GFU3Dvk6hvIKTRUFHWQ1U568bh/ejC6u1
S7miMr5SzwZNTujCEXKwLduGfJVqhUhzXxRfBuzbrI2vvAj6j+Zqm706VLa0eGyfxXR5ddSNlbiz
2Igo0Ujsk7hk5bBIgPA6yKNucENg34tMYNdNwz7SCPCJG80goE5WbpZwKoTgXQRQtt1/3NePx8af
PxGBjGMwi3Psp8g4V9joC/vfBPwt0zkZmOw+4/0rIsos4aaGRv3kPvU9D6llFHhOI2RxDQmwNxqk
qWOuRZlvxrJPSIc9OIMPHv+d9itpR/akGFiFwctN4CrunzxZgdxWAeO8CgpDlc4mDn4fzX7+iRFn
hSRwLNKV/Vt/6PECBVR22f13DuenbSviEGLWeNYL9dJsGTohk8N/LfNbXhQQ6f2glmHTq+kg58eS
JGZcfB/OVUo6wdKQkmXBqbtAyKPKaNHfeuEO9sJYqjEVOz/bKuCm7/k9oUSNMcrVp+EOzY9OBANt
jKcvjmG6FEF2SgKSRKwWs8anpK9gJRNseeJ6r5htA1SHsmhJYSUPpiVRwKOj0qqFjSSd0h12HKNO
eEGnOU8e6mBCQua3hp4608AtVZJHygb24rW9PIwo5XUUp4xUGLUmOsdwmyP+0M7wAcDs/Ji4Fpv6
X2lqgivlTHEqA9Ww6XO45fvukcQlgSQTXqIGcCxXbKf+ehwj83jYdFu2aVYU9GMP/+tjfXZ7Dz6j
Estz6A7Tim0Jf2J9AyFP6PHG+gBpC5UITI8sVsl3iyPGAC8sQM51v2QS/8iYH7V0tAgOLGRA29vc
JiFog3nH5avdU4sUd50TXin0dPhmLv4uINehoTcvbL4bHj9ZgjpBd16OZTSXjKsSzWVNM8Lh8vwy
Y02kBYwV+sVkg/RYWeXbp1+uRCKVc9m6qapyNvsQjjW3X4oga2qYPJMvZrZnEZ8LHSrA+AOfLx/2
1ZCx5fL9aP349SWEMz8ETNBBAHxf3ECOnPG+VITaxne3BdVqr1ghwCIhNk4kiNoAz4qElxwUavT8
i4rghDM2yvzxQSBt/OWn0Ly7HvZEDwXqMbvUEJzH6YwHDBGzevc9l9h+B7fy0UJ4ooLcoKKlEGui
ACe3ehqJuSE7Odhoe/dKhe+BzR1xN02mowRenhe85H1Ua3VNFCXD20QuI12ptmobLIpa0HRrIREn
lRYcM/SZzrlDXXdJqPPqYvghnrYK5K9581sL8H0R7I/UcHwvVWSEKW8IQBy/TT997it+SxLhrAMh
SN+OkS+3UmFPETdyPTv3kOSWMo+0+kRCLpA17mKE2BYrE9WqCm8zsfV03oqe4rFxAEZEmIefasX4
R/yxD0OngDwshMkN+4gRHjc6TUqA/c3hA+8LHFTdgPIelpwLZHjaMJR+XR00bMPGpTi+FPtH2iBR
hNvIdnxcCvfVUauF53X9EXNvsIRYQfw74qYwUaO2dfZvOXItSF1YluN+M6NuYr8YWf/tQU2vQRNW
PuH4oVb7Qu7shtqIhRtH7I2Vab3LQeW+PJFRDDs/NIK/pOZXx+oJ68EK3xniAeybdpeFd4USq/oY
xlPnuWytU9y/uaQqSdM93Uiqx/kbdSOA/YznbSWzAAwSCTymgFsUO3rdltr2jRwW7O/+jCJTdKnk
/0hsRUDTl1/5c4lmCL/W3HnpPBWSg9Xws1019PlMyw/eaCUHNJlFbLPfA1YXd5OallhWwbulICb8
3zSdg4hK3YRqC+SKni8gAn1camFN6IF10k5uXq4kFLQzuVcM/R7C49LLyg9HTeNJWUwx2QM666u9
EUEzau7wK+g5MbcsTPq2JoTJh5M34YeLREokMDdn2+MN6iNjLD0rx7ntfZSF4vHqjCqrSlLpdvKu
da+uF5tRUNpttGHJTXFL4vL0XE2XPd7XpykrVcYBFzHwCFzyTYJR3+R/Lq210WUII5fLwmLI3wx9
Ngf87Je6RX7F2V2/IYnrP8JhpGzPPGyC/NzZEy+Qi9Ug53mT295o2brf7MySBKPny9cjPDUsqAb+
1KNOds5tVE+WdAXn0hTMDIh0YmXfSH9S9GFG06A12+KbUTV6Kcn/pE1Gvwmc06/iGNKdLYOKJdOC
6mN45w+zGLYFpSH6sIPFoJuEQkerITgFg79ZBkRrYG6h+O8R7ejor1f2Edu+qZW4EjCHlCObv6cw
wR6bEMSIdT9F8/Vxor4s/BbpXQ9ic5+DfuLl4zwycNzeH/lGYXYejDPDWTEIW9mQ73XjtOAl00em
nNACQ69nLFmucPO2+DGnbQt142hPmS8xTznN8ZEU5DVJ+akD8mlA9VMetA20fJrJ+fSm+X4uR8Yx
7v/PxLG1gazaTJK/8jOY4YKWaKG7vTdgZvtW4ASyV3M5Sc5d0M8F+Jy2Tb4h1SQRjbmadWec36kg
Mar5fFy1bHIyLSEPAnp8tEx7V/GWF/Lezkye9FyNM7/cNw1uEYHWaqNJ31/D1cx4XA+oTqstzyXd
8MCVgdq0rz+iVU6Bt0yO/9DrsbTOZtnjXZU5oJYm/nPkq1rSnz2EVTsAuH37NF8pEFeAJCgpAClV
wIAP6y4ZcR9hKujZbxFqMlp8MlwWujVkfy3I+7c44/tW7LZMrQdf+NlkoyAr1/kr/vn6wUQTCz5y
JMDl1fDgogmhngkqXwO3m2iJo4nRpI2wOuSuin1/4EShVl7TrU69W76m9Fe4bx7CVOkASsSGhbqi
ACyqAw7pcLJXaMHphYWWS2HRrBHzaTLPidw/uRPDWfDJT+vLyIvpZzrBMdCHxCnYk9ALNWfqRrV5
ttQ7uNgucV1KPkXGqv4L/Ui6vw2El/Etwjd3YJzN+1RR89Ug/AMEfTouyCTXK8w3yOYSuay76aDp
r3wiNyE3emcen1N4WFZvkTGikpXXFIkWpBauHt+TRPmYqo7tKGQfKN/nLsbQhgS0dexcxITB1u3J
Xkg9m+rJP/d1pSQN0KuMqg83fDQ7m4MOl11aAZTHDXAfRyz6rJHm/6EilgMXRYmaIAmJPCVCyigT
avLfjD8iHzpPf4XHl8yiiE3Xr88r3SK20bJ0SqG+RNfNh7SLQA7gRU/fAB8wziYPTZmlbRkQ5fkY
WrR2OXG4P7Ue/yqTCW5/VZHImW1UdFX5Iogyh9zJvM6CfF050hMPyyaqQYXWv69I5Fu7Ev+TZ+x5
g8IhAtKuVTP9+waSex/mHqArCl47+IJkgr9Q3uHIYNadkxCy8QDEbaMYbEKoX1LPmXfGljZatAd5
llHpVcVxje++LC5LCmJROrjVHNE1vI2iadIeotrdJZGkmejZBXZsDRC+FraxG4RajGZ8XP6k38xy
NE2/qYQVqHaqfQQv8tGybe3FLz1OqlnlgxRANofs2Wc4s6o6+ZIUhmoX7ZG+5F6KwBWOczzoHd3z
MZvETztQ3nXayqyzQ2uLwi1SfFk8ra6fAGgGAHsB/EhFZqszTAQh/0RZLpWwNxzzuKDzN5V/mgoV
00BieOS+tRIHdmGchRznHE4mb6/MpA/vKeR1PKw/Npansl5WlEv1KFnlMx27he2J8y6Sy1sGPM/N
ByZ0/3znzVAcSslE9dpySWfjaD5VcTyY0GWzJhelZ/z/nB8we+uw/bITbLRCsHcwF8IH+dfQVjGQ
aIMyjFiWEFOdqMiBNfZoWWCmRpRWCfyAdbYljJ+dz4uHBW/tcsI8kWuR9Vt5Xyd0h8jqY9ioQYgM
4Utn6Iv6UiAPRZYt5BPiKIvqm3HfAVJaPZLYB+2teGl2i8pBNbJ88rJBv8O3IvnrFbw6XQQ2mfCk
044sMgs6LtYGZIDmPiq3xWvUkyTnbev58PPph9iBpBFORjb0Zlagsjy3V25ztobpAI2lBo1rOV/O
X0mfz+OkeWggY0QLTm0q5XLRrdaQasg1W1g6EvnBbSC/KZFpQMuExeHpThrAckOScWq2oyS4H3Dn
jasspUrG/cSkDi9UU30dTqBwUVcHxaP3T9SLzeCEtYNbdQCfraR6NGeyP4VloaRmG4lDknYaBlJR
SLAf8qkVSyX0yhTYchod3tgy91dmSTsQMojbQ/AQrDGrdQIee9J5qZq6+VlSF7LFlweGRjE+y4+g
2F56IBU3rM26PmfcEenMn75qE++E0GcCw+Df0Uph8sPkzVCct/kLG2RnxUH5+YzPWHin4xfXWzjD
4jdWPcEIrRqwrlXF5xsnQ+0IqD2DOn4C+IagPnXGWFm6mpJe2KeuFYeFKQHPWMfcBV02Yi5kaVBy
GU181CNzMLz+L0dV/2WZtz6pB6Xp+6Qy8SCD1n8ieZLQnW10g9hZ3B4KJGxN37q9nvb4qhE7pG8j
ef11sd+/AykitDry4g3UTBh3byAE/vNXZ7/MDnBVVhlO1nwJ9M5q88fP5kp6xRPyoYpl76I7LtpO
cYSuLmZHABDTXVqgg60iIQve5ylxzxq285gfloBYEWhO+XtsL955r+CYupqYrxgp6UIPn02PWLnd
n+RAErzfRzH2hXInh9kRJ+TKJLi/n9npXMAWwuearQ61ill/WpfQvaA91C7KoYGvafHxDZqTv99e
T2I9+/LC5D/tXE2s1uBb0mzBDAi65QY6LlJe/0i+RCNXcvWKVQbvGO/MUBw0VINoEmzoifuLh5RO
KjOsEsjp1WWf05a/gthyLqR8Ebh9lB8rRs2fHqFdJ/o9wTqehzMuT9kRPY6T8zFajtfbs29ByrQo
+qUX4TvCfV5htdadUMXHHefZ4laVGqmVEHApLtdXX5y+s63r87gVhYoybA4wDJaXC94MbdNevgWI
wuCgQq51greyBKg5RwDs8u8eXB0nUWIFc0TcMFzRCpdRRo/G1naGTOg3aWZLzMutwCwM8hRCyUOS
/uozXJuoCmXouA/mIY3mei/EuXjHJBCvlQ7w4+MvieLTPdpA6tel3e5q6yhrMw+ZGtQzk6Q3L8AO
h1gFwmoOXfxsWMjdQKQa8l1kkCK+mxM+R7KplXDfj0gxS6fUnxi01XPIgH8LVK2tHmvhL84XqF+a
mtA6xIWcCV7eBhzG/n5vfiDr34YK5/HSwtIesQg0dh1bM2LQdRnHeF/3Mfoy1hlSDEC1PR6FQFjZ
SXbiq3SWRQiGhXul/VsiNsCzMtgNoL9o4rstrUgBsP691O690C0YJ0WOTZmfI5f/n5POvGEDwO2I
nXBc4tyDWoZX8FZkiezAxtpiACNmdpoa/D7Wn2WdhdcoZ2gXORqor4L0WhNd1AVnEcq9dWtbFdxE
hWVdDDSAO97iEdE+jWXsfM9ehiPeu5mWYM4Bf1dqrPpAzSeC+hC2pj45QRIcPDMD/1n3dvUHyP6l
JBGRzNKtKIgkzVkBzofGZYGzlr1PnD04vlL0UGFNZXWPPzjwkZGd5VPATj4LoI+Lt9pDxff/kqkt
CqorQ+XH5o8VyAars2E6Gv8PjmKBr7IwKMNZwYFTcX31jXhd+t2LcnsuRAOi92TXkuTOcXY2Snnz
xWCoRYkEkV1L6oEYnqP6za6BeeadJ7cuZ0NRcod3tAlX3TDgWrubphV8U74lCAdUo74WOxUVUv82
pUJuN9cqS+3z17k5cBLCrJA3Y8HvHbRYcNoc9N4Qk8+wfYI18p79qoyznbw4QvJDBiDBsThicJQ2
c/GB7Hcvg+8u03wn1JBg6tnoSkMSea8dCdNFgZ6+KpceAAGahiXNRfNIwqtccYMwbGGEoBG+DCAK
KfAKMBMfWRuUHcgVNEg4Ir4ksStiEZQneXqW6oMlEwhvPRVGrR7NeLARQuPH1T6CutctyUqTIoDi
prNcFUjjv1YdgSkyj+A/g9H1xeiy2JucybrxtQS2lww8ENd1c060J5ufHQ25H3TiBrlbs/OARYPQ
6gXI4e8sudEvhyzqBBB6dIy5CmpWjRCrCqbeYj7bUrMY3TPGTMA6tCwYvVjbEQeq852X6psf/m39
9RPYKomJz08A7Nj1U8XQnd8b/TuSbBjALlJbPif9xOIxUFshuNbcbmUYSfnbqc0JyatpoIm7migX
r4xcy/I/fkOsItf1vfFYNdSdT8QBLYGSSQYR2IyF08gJadUi6hUcsyE4XYPDJn9TwFXNa/NunGp8
QhPsPaWz3qDJrijJ1l023VYQa97xUdfYwWKipf+KXB6nfcXEONMARGwhKIyhMJNGVlyFC6ehVakF
NKeafnqvtL640yrYcRC8iDciVAs1DzvFw6NHLByK6FUcSKl+GuA22MEpBHn63KjgZg/oROU7qO0l
gKx0RDapoV/Ni8pql7Y67HpayH3HW+HLOxLxyvl2rR/XdpdEVK5zbmaI2zJwFA/DngUwOt8Yd6Y4
iRqgkPpSz0UHCAJ5uGMcV7F2gmGFzCdduMQTYkIs/u83wu78JH+CI39n/lDvZr6q8C9/ttk7aIB8
1d5S3q6KBGL4XLO72HQapI34I3ycODhzaU0u2mFZd0WJXxNSJs1nOZ0GHK9RT+6eLrU6WO8i5zCE
3J7hOiL6rgydftr2d6nw85yisCe+0u9rQjVJ74tU3sSzIxsgk3gWcZqf5umwq6wzXKiou6OWIrqc
4ip0cZ0ekzYwDCVnkb2hDiBg3591MN2ebYbU0FdL90KnTvp0UfQB613Cmv1tyoWBZV2xD0LptHyl
r9jk0s3Ju2bvuTFYu92Fi+Za8ISOUCNkmpLiNWarNRh4gqN2QiLshD7ptHGFc84KBguRedR8XqeW
15uXYmNDFwv7FBdIO7AEM7xVZL9FHThS6oJABE4AYdM9tIEhLKpkxQG1JYp0s64L9J7fmUAvzbqh
hkvKU+kfttu97bCVU5ci4WP86T4k2H/zFR3sl3qgD2wmn7jaEYcXkESAGhuUBTSZI9J0qwy7ISV1
USMCuxkc2/UZTQ7p9TFBeND8B6BWrrPIDNwMnzP246QlwwqiBrNBKpWkfXqBAsEPAhJn01BYfBnb
XWR2z3ejnJHvLXA4fv4o8rC1kJiuskkY8DYF8R9+jQdBqcUlJ7dYRKlOW9QS8fI6Zpo9TfSHOPQX
CQL4yGNJrDiVc9aFJM3uWBO3sxIg3KxdTcsXKOiJpDr6PLRMDq9RrURTN62IQ+07dCZDYYd+kfwj
DtjJ1b+VMPx/eFdDeg5i7KwttPQTJy5CfBbwfoewAoMq2Dj/mHmW5DoZivtGCJVwsXHMERs2ITLM
tnyJG126+j+VUXb1H3hOT8sYb6eVZ/STVAemLZDx+LvTqr9KA6Ty7UUagDDWHSG097tH0kjTYqVW
jvkW1pIZO7DCx+8ETeIWzIgY+BnjaFl7v1nVyCTs8RPSrv1rebNDm4PtdSPSEtmgwRLi1zDKoI61
8savF2uAEASx2V7f/bLBc6KML/TlpBbDK3/As9hPq6yyo7fGki3mLzA1nAS4AHjTBTA8BZ7U3OlG
RmGyaahrJXWmWbyC9QBWwmN0K2W9JejQ4QKzRQBTYXiPJ27ua79tfkT3ZCP9/5Gd9A6Bl6sLGj+V
hPufZvRjd0EU9WH6VfSd3Bhbq4KwSey1ZvAIOHjwfvs3RC4KYro9TRf4oghW3hhq7FoilVXFQfZF
s4GLZjGK5EG2DpPCGLiv1dFkH4eRPLUJ08AqoNURCWhXPVsH6MHi6MU5iNJgMdHAY5PqUQBddYua
JlZ+5QP5z34yyrS3IWpmW3qyLg7mWzO51nmGUk+1ySOp+1CnzmPnL74dOUB4Pj6VDjds6VYO6J92
0KJn2dITLissn9MnAAEZQDfj+h0/i/o74hdTKsJKNtIMCeFuJg8EiCmmZHnk29zzbUh/Gkwfdv+i
68wU4+FpA+Yyn+1FAhIzY26yFBiVrxgMPE4K0hzyUUh/V7OThTxGIgFVVOYxffpf0fhB13s9nIUz
h/wK5erADhkbB1XmSzYh5oqn5CCfpixCCsD+pvY0fJPZv+MJGPiKVPX2SRsLmZGGFkaCJ2T+1aV1
RTVUIx7UnUBtORrNqph4zFZxuLXtmelIhG739/+mSmJeC1vMFObW3JrnqMRUSesBk1HRqeMLIVeS
IMbaFTdgCQc1EMupG4GB/+F5ahHXyb86R7L/yP/Uif8NWl1nRyOi/n90awuqoZh/1XTNrYEUX/e4
WXd733zPTg4QTT1jhjiewFsYpZC5Q+H5aJEe/nXRyoL+8cR3QLAvPzlTB8Hq9no88TUwrXyPL/Pd
yYgU7+XzMi/NwhzjVaTzdySOMlgG//EsdW7WTInWQBAme4CBYVEqC8STPi0iZZo+2bkTNCaqUEgD
uquGkD6VT+vyFeUvBKDvUkZ2vpouNebDDIxIzhpi22pf0UKSnpO6YjW4yfNtCr7U0Xrp45jyYL8d
UzetO9yUeOxRzJpBKI6FU7uo7Grj9cAihgCeque39gtPFOB/rD3/1fmYneJ8R0JZzm3QttnuRbuC
Q6OQ/va3SR6RAisjGaZxU1n3ri2p3ibvwM81tbTkygrQGyEXSXxrUmj1nrzvUelJ+cpdGAtMoC9T
/KaiWpjtKEW+U2nZpLunDcQNfTlHpYzZXpOC/VOUGScO8SN7RvWV/mNFCwmGsUJ3l8gcLssuTq57
phkmqF35EsOCYI4EKe6QW/MU+zA95uNBSyG2CYp/bAt+JBYq2bBGEMsw2ymqre30GOjrSN4kHrWC
9ldVDLEXOxvE73bYY7Srkl+eTH3U0bDyEMc5Mlqa9ZMXFnzuGfqa8vnV9zo/u21SEd4LpplIC07k
vjwdDRB00R+AXiWh9upsBjFEzTA8q2+2jkd3fdAbZYoJ0tny5WAaDSAsTz65qdmOHnEGeFozLGfn
SLqvKPFFWkxzaTuxM1Rkwj1LPBAhameONCC3ktAj5goPkBZmlmVi8llejE+YX4Ghs0B8UuzU+zhF
JUT5d/L0dyybHOOUu3uS9Igzjr3AfGUWm79aPePZdP4sLnIkRJ8JHo0yfPJRFBP9yx4+CXv61HVT
6X6sp6fGJWTkzSHirz7ZEJXLQW1lk+VqeQNaS6mSbS65gK9LMTkJB2pn9AmSWrK6NMBQMcV1hZXa
oPaF3BOgzq/RxgXVqqiJgvVNNF55ry6u8wAkPXdgNMOGFfp+KswoiIYgJdl8rZeby5dqPGDMQsU2
yTPtmchwzYBFiVMxnzMK5SwyqPQAs7cxbqi2nWhjOo+4ubgKFE3V1J1rhCkpdwCnke8g5f/znqwP
PS4o4NU02SXqoyAGPbXCkhFqvG3j6UXE3qVPjlSbABEO1qR7UoZcqcPPx2R9yRqOYnzVMhNxiYWQ
C99Towek/A2BlQz4uYAFI0CgaZmWMb4c0+6lS2m0nO+cjO9UAb7HFHvcwFejWx0LkzSg854nTfSq
vLoK0YvwFLpe4RR6hJdgrXskX8JcS7NTGzFa0CXFejJGD6o1F8M9jRO+jFwRVk/bmZ5aCEAivPou
I50vyLio0uyxqzpqH013GNMX2MubMc2/o3pxgc5Hlubn7q/VdLd/FXuVXkUU+3UnvrMMY6UKPSdL
vkcN1a2n+q2mKZqSCIx3zpI22US/h+v1TxMQ8WoGBgEyXlRMNToKB9R+QBKdOFrT8OtaVUejDtDC
2Mc1n7yBRKDc2pWYnkXoERF/XdBiAvNwrDGWiD/euJpIvuxFgob1uHb0PGnKFNzYo6rXYWHEVzVe
z9jQYfyOYOaehZ1xcZ6+2ur67AZehaJfXUEm7BhR7bMrVO1iOP3PKC3Ra+W4zOGwq+YBDBVfmI/q
3I/bNBYX+OZ1MJWymoeiEg1v9+qq9SLr9dgwqatIU3Zxgt4RRMtBIv+WVHzBUp7MNti3wtzeMFR7
3qyR7OASxCXnOQoRMISCMvhogx/5Epn8p1Ru2354WK4cMOTQfAafYyEP/URvbgR7a8uusJFgbs0A
xZxM6e+1gVCc7lHwuPgjYNvMzF+T03NsrwmI2MDBwfpjhOo+thrG/ypjaie1EYl0KnG/KcGLV3L7
sWa8lJ8p6kazFkiIWuqLCqfBTOAp/3IivTS7DuB6nnEllgfUZN66as/xAMNVYulcDnnnvlS+gn2S
WPqvJhQYD5yTtBd7H43ZXs7d/m9/rBm7vKa4L1UUGhbthe+BxqpBlfmFYdAeu+UmK+KbT2JJhbmb
648FDSRHL9vQcJ3qGUkX0/yM+VQ6jPJ9mlHM/uirV8D9+Yr7qPXgfi0s2DF5xWY4B5HPstKLNJR9
6BGwF4LTt1S5tlwA7H8nHrSrPWTFZI6A25z8faNh5x2fCelXjvFzGrIbhlHegWI8MvAG0Ood5v+h
dMRt9DY2+WVQsva5tM70ZBd/Lu0HUiOQQnX6LCw4K0WO9xWhkigCiupmmtu61X+DvBjaImf4/jB1
Gs5vh353T+6bT+Rv7SqrXWwwpKpwpgac+HrE3BsRTPzkdWprHggT1bsGpNtteDbCkEQPR1JmEDbO
R8vC/y1hpn7HyBH9c2ilSjj3aEf9ut/T9tC3uxmZvaSP562Xxn0RbBp75FlnEBZU5jZuktj09cEO
qai/ZvjxmWob6OAb13ujaRBaDA9/y/THt5KSe+plT/QaGOGYxVpJLBcBf8q6zqqFyCc+nc+wHzAM
2evr76utr4S3mWtzKOP88XTuJq/2VRILwt7PDWfV2qU+PA42tLShOcoWAwC+nUpv2CvdC4GVHWX+
+/EV2u5wbrD67oMkCai28LRTZb9EO2aIaDxV3O2UYcktxHRnpbPtplSIfX4eWw/xvnLhH59lqdp0
PUllGTkG6XwbIX4nK6i6+tTtdxSfmpPekYgvbg34gvKdC6LE6nvNBOSVO1/iTtrhB/Tg5gKM0DNn
RwipYXkiYTSJ60UyszBBZy5jOJ+z4fFX5OYHdZtVv2oyFW3Fg/7XL/JHfF1LT7a34Xy7xW/nGfP4
j5N+U7aN0G0tJwJCrbM+9/ZgP5SMFGnBzk7fC3tJ7sxR0pkM/o+y8NLaqItBDzEug+aJz9UfsIYZ
9LKUjFvUMxqPV527KLPik1suXN56fATtbmmxPQqVRxnWX+Q53BWYiJCNuAOz9qX6UL6m//BHrYb7
Vsb21YH8e6M0LHpsh0zej6+FewZSJe9ww8evJtuUxwv6BinqyVZqtYBqyeBJZkoEfG4SsBPSNEg6
KevBe6SvCAeyV5D24OAbiNMbE7INQE1Z4kuF7y6LqAoe8qlBgKfQ6A5jT2v4poBSY9d/1VVuVtPr
tO0Crm44rI2m3o3l0oaKUbpr5HcQndMR4uT8hPSb3BOIYr8TCC0/4JtaUBURA/T065R+obog63G+
SkXtEafAjZaVE81R1H97sW0Wk8tdnWG0R9UUi7zsox/ZJdu0r3FaMVJJEIMS+JVZO5rgwcgES44V
9UyiCU0EgJ2CoJZvJ0/V3gKVipij5yRIuu0XFeIqSgMDYrvtnawAQR0RvL1ok4ixCPocyyoFaXoe
ZhtDKAlOaucIqwQcdX74uohkjVMFzcsWXEIMKq/wtt52cCEFyVPhN4pzojIELW0LBxEJ04M4FOUl
/aFBXT5kCaHwXqNtysjlpAH0vvzhMTsBtlWZpE1VzYG0/O72impUX+sKM2aHIE/yhDctmnhEdTAx
SdLM2O4FWfmk3XhVi+5mAYU6Xw68DgbyOJjr23pmcSIVHNRUe6cHPVgJDwt4alNMizMxBGy2RB7n
TnsAHmGvqHTjE9T0hoKTcK/71d0igMvoVLaxKqKxlJ3P3aR3XpncxSxCccF00l/vepYI4tnHg9Ut
jhxlso/lfqC8sgNLL8XVTZ6u2FZxHjNmJ0pMPxDrxaFCtyiIY3cyfA2JOZLWqLJ77/zKc0AZP6Km
vsf1MbeETq3kZxKQnPcOVFocrWLnPpGle91lsMpo6KT+ng399vSF8ke6O+t6Sx+FBtASE8zCwT1e
0Pl0z8+9XpS/B8EHHmVplRkiNkwfQFVqkxsHpTD972/YNULzTillOv/nqp2kLZTAUXtwB4/UmUuX
VmoX7lBxHceNJg9JqVaZfU5hblir6MLJtiTokH1CSamo7TrfMq/wYBrnnJmE3dHN/0ahUr29DPO/
KKAiJsv1GcAH7KaCTjYFfrLl3Kgpq7aVr+uoJh4ARgOo9dJ3BmlpXqcUaZ9r1/vT/gZvwJmZxK4l
oKfqhNNdq735Sw468bYEX3CPzXhy2djX34AaAH/U4HFa34/N3kO0+oTsZ0fLtQyMavYssXPH8xz/
PFUm7U0CwnvMqH+8MEOFZ/2fplEHmf/QCGCzdkxzs7Hh5FXP/xChhSRPjFtHgx2jz4FdvWkN1Bkj
HvnNHSMLTxY4ji+++P5UlxziDaNM7a5GvXV8cEDRSi/bOi4kFBuqXTAjuJEypepvEYqqwh1Ndoj9
vJWKzVpJbbPry9eUq9BsQQQqnF2PtWb3qiuW3Hejse75ud6H6J/uYtJpUzLtmOIG9SZDuGVlTx6B
mvb9vMNNpRyQkuIy1y09bRgugWlGTfNC2+CkeVcZ03d7G4XDdTdaAxc6FSM6pgZvZxhdScygnapu
eNOlAgql937tjF7JnYHis7Fl3gc2H2TIE4PGlj2CH1pDvuWsv2C4dk0f/4zRDZ7mVdeOnOpCH6Cj
KiRJTkw6hfULvnUxzyEGf6E7FxMfcUeMzCN+6R+a/g7wE3aHLtaFQ0CLVVz+uHRZlxqXpolKPD0a
Iw4VskKRmbMn65tYHGZrqAoHKOBENuniLkGh/igGhH57UOhiFT5aGZLpCGLLD4t7n1gJoZJLl9r7
GAKMJE0aiVVbIWTtRv/ZvFW2vbOdoLZF/Cr8scpW1oj3NgPQiL3qf44wLI6tvBmLYDniN7HBiO8y
7v3jVP1u1at8Ucmgz5CTyUjhOvhS6KTxAAf6ga/KE5XTIDjAiDIwKMTnin3wMWL0Kclh5/hdNCgR
sA84guUfnXp0c7hFV0QFRIiuHhEo9pU9eqGQkaf3m4zZbwS7GVqSwe1ctr4sTAdOKngU61xE3OWO
IklsA8EEEuUP3LjjwFF7sQ5CyosFxpGy8caTtKfkoh1/Im3mlEyxftNQpcbxLkOKnw3MfFKCadPF
FNwLUVDn74V6oKONnOPLQeQZTAl+rwSeWvt/VkKuOiiEcV7tI1avpPmbrR8qsxLd+fIrgbzRZJqS
edGYttiBytqxPBsvTNn+/lyx0oU8jScvER7BpZ58aua+XLFUdN5l4RpqIj9DRjt7B17k1NRXP2P7
TLrFxAFFMt6WBunmCmjAuttIh76gQ10RdWmSqrTioB+pq6nW3BYwEmBpFjlbKkT4KuZs3LXWZEeH
sHuz4c+koOL4s9OJTMLhl/AMSK09FVjP6FQ7UAwK8LcqXVRnXKixFawc1AWx8/K6O0OmCwd98e66
SiJ5romA/pHYwTJGIjwCqyscxeSSmfDIk7rOC6Dp9ZhjSHmViXjt4lbMoyg6dhkv6yqURucAcFJI
KdS3fGRhmYaltti1cY80AL2IwJLQSjqoXWx6MQgfrZnZa5xWealorM6E5V8EvnZ3GTSfmxcKahSf
OtB1t+7tHQqltehJiABtkzl9h2gOFz4vtf2/BJDtza2RVr+m9j2ksOwkFBelr88Ft8wyHXfWXtQM
t2HY5H1RhTatx5KnHrr4YYOpEk8vSgDsjoRDoCk08QJ9zWX27thOJwPw3kiRUL9LktaR0xBimLfz
5a6qQDD1lBK+kIY+ukWPAWyHIfFRJafDmW2qJXaHAjAa/ABC77LRaSUY9+uhl3CmAP3uhAeEwtPc
jw8RDvRYTX545UHjDkjdod4Ta6Q1l+SQigAlo72XW1yqWrqM0Jy+4p2zAk7WwOb1/QbaBNr7fLZy
83DJ0H7gZVc1oUn7B4MlhKi1jkcwECnLBOxLRTPPluaOV5E1yMkgNc0jgdAOvF+qx4IAlT0c1UZf
7lSdvmWCmkopit+jZazX8xwvPeHztEfqGxP+yF5RzKCkZTp2r9352p/gDeHLZv4ewTDWS8Rzdhx6
F9ziHK5IQneRvKVfHUBOCVWf7TpUvo7ko1YMPidWmnV4EoHRoP8Aypyp8zlv4sybVh4g3XeXnlBu
q/MqSD+qh3iKYXUin0OrIVgX871C8/RRZucxSIBU0Nb8jITBbzE92WUutwtO3rmUI5GePS8iG3TP
GHas36IKkIotaSECb1vRZOV4ufekhBXKs6dVKPFQZ0vrKT7ESdMSydEbeHoIqcGCtBSlPUvmZeu8
YQX9dMnbFbfDwQTlgAGN1C09RG+jZAtAWGD819J8T/uv0jJ4MdRmJCPh4EhfF9VL4Yha7JIFpBWv
A++HAEb18XtKoXfZ4S3ZJPQMt5v6OTzDhPNUqttDbTiv/SIX6cC1OPbVFTSLWZfMTDqI+fTmIiFQ
GP+D4uaz5BKltEocClnqBc1LXq8fXKnUdz3AwXj1P52CHsz0x7uEFt5pkMU7ST2K2wIZS4OxnJRN
mLJMJU5zomBSuUFc6JdlPxuxuiN5bZC6lXzHGMZNzZJ6yCYPMi9KP8013S9GmBaXOoo783w5DPvL
GuUVL5oX6hIA0bPS9c8qX1apcDemZdHtVU0f+szKlFBm4NtFqh+qwhmXlRiOMYimXTXUXpY4/w49
svWsfdyBMFWrOeBft8wCPLxbzzOhfdjHRoYY7AROJwJSac1/w+slvhPQCyEpMuPLX3nWI0MD4YBO
Al7KGUQ9XhwBgY11b4dFL9w8EfjWc9j7A2LVh/ECJH53o4vQQBbyiQx0X3R9MqTZqjmayg5OSxfq
uMz+LdzHdxxr2c5rMsMQHaKSLU9sK2l0YLll1hHRAdVq+mZ9HC4ve0dxRaYegU02LCVZxk8lDrgE
1j4Qb4HIwVmTHKOPfhH7UC4wPTd3eBHfkReknSHpuysgbYfI56GTQKBNhqJ+Wxjcy4VUFdSThEUq
zbRiSmcnrqL90MDz75jsN+MEzBmetOaN11nPl5RKMu1WsL6suHJYlL5yrM3uy59r9EA4cL5x185O
BgmHcxAzYLXYitoPvBMXh4yJx44TRt9l7tRiRT6QORabKI0y/DXOHC7ASMtQANCn4sMkD0A41rW/
t6K0hMVHegV6YO+TdZOHQRvjDnwLypFfhLW+HrHNgozo3bw38lrQTLGxSt2U7J2WPXsQzqChO+WT
UtCzRoGhW6tSHe61zdnXo7gEMHxFnnbqFaQ5eMF/hQc5W1KvLzoScgvoIubH7kClIRO02EEI9tJ8
fKnhxDieMBITt9CIA2Ti0llAczLmG9UXPhw6m+wgDVD5wlzhy74vtnyF+hBEyOjFHPWrC8Zi7xDA
fcHDp8wxzauUJcMVC4t8jqaCbyUUFcjcIS7uw8S6jF7sM1KudSTXGO7GufsJHE3OMgyX5Uwk6sfO
N8Jft1MRjQhFEqeUz1okRTQzHsV3MG8MeF0uZH6d6KHRxjr05s49J4rhDyAm8PvzgWCmAVP12iqP
ncxKgzz+7+/0HD1uo4fQrApuDgGNblhluEpyRUP1GK4gv5tt0mc0bd8p7uChanyTHrxYNhIJkTZH
Qs83ZobK2Ug6Gn3dyWCGWL9FqVMdKTkDMSG/pB08lk2q0HBC+eUbKol572l+shoulVhDGiVZC1/t
j8eWuikZCg/W1pOkE0kMY5ARamsjPOmAOtupkTdpUJcyU4XG7FWgZutPzjZDwTvP9dswsDuEK+3p
Wf/UF67ieRdWSB0twamESPp9MNaitJqlEifwg2LjACpkDXzQucwChoAYf6UillxzgRWAbL2C0how
mqktMA/sQKhUxFdgEyoVX6yDfeoMzlbIx84xJozvau8C4pnneCF+GzrRwq98hwH0DXwI1XYtLIS1
JXQ34LzDlFyenQEqJAj4Hf+HCLEnHg1XNANj4u9ZhEXsquMg3J2FOzahlt1kvhoUTDEAhL5pde9L
4rJUkNiEf6onFvTYlJ7h+T2/x5ikiClpP7H25pz9w/pVsusi7Al8CtSv+zEkuu3CaZsmm4b5gqTa
yYN9IgKHB9ILvy50URQ0ES4lRxxTzB/ZVMd1wWmxxlwfN979s1OkPRtBjFYP+oTF16gdvrmEgKsC
hKbo3ZEQIFPOwGgggfBn2YUF/5j5uHYKgtxDR7OFuo7fGrliNBf6NZmTk1vrxWpI72e6Y5SHc+vT
HrHl71vk6BGBUeaJQmK19k9s1TcgbXcnYGxAO/Rlu1gHv/i3SUUEDSKeZjNWjH48VmTjlt4XOXXC
G+q1OuWhkLsHxxA2b6ggClP7qldy09XPaNuqgn1Xc3JXBJNbhzx2bkv9/HbltKx5Qr60Dtl314ex
NI9CAv+i6uaTebDzMWfmOouAoCvANABiRuGb4YbMIvHODp/SVE9Ae36BriC5sQ1V8pn4hWbn87FT
w/eOIpJ9HK1ZUa4ouV3Ejr6Ohi824n4WrpSjK+rfcoKFoCr6b1bCurRowMkmkexD8D8eWRXr68um
aINewdPBNqUGMS1XM7egYONxZgBdCBxPOxpFYxD9ta3dK/H+Ns0rMGKfgs0zIE8c017ADvX9NDxe
CbB6wFvqhTjE0zN03MHdUW5SgLzHH8NBhAP1XYa5vrnPCwZu2/WfyZh1BA+sLG/6dhvpcPEKuhTE
aqCJJg0bfvsEazDc4E8urDvLTQyv0F5FGgSLLtQNQVL0QH7M1iBUn4XYz4XfOBt5P5nlBKfLC+Mj
QlhU8t2t9Z4TEKPVUkrj1ARMzcG5lMvK62KwZ0mlDOgfSzqxakLT+Z4yLk9qC3X+v955kDlx7CCc
a7jfKl2t3PcqkbgoFd11xd7jL6S/e+Z26eoam8qhYsTEuNpVxJXCjytNHLKPhClDEGsKz2qsDxTr
vuM2rr3tgbNhF3s++2f+jJxZCJ+FIDX4TzILa//iEDmkIb5b1D7GLi0R4uCEYXpY+0QYUbr1xA8m
78XwvtWoZl+qMArhpSGC44HEXKFwfEK+CG02c5spJ/v6qkSJvnIcHxpoGJNxqtL2wqdHvFjvGfy1
jQuF1Rwd3fW7xMpCPyzQVtEY1lpRWwDUnL74HHmwoL/B+8fm2qtrYxZf8WKNG+9jyjZDBsG97ipL
cpkopsh0z4fXh26qwHCGT3tc9nOF3PAV/6nTvgdBRvlII8pWnDwz8dYA7+tfeYtspmene7LEtWEd
pMJx0Xr0wyz7mg00TrLz73gZqMDqHV254xMHkTNH2gVK0kr8a6GLgKCcOmmg8mphogPpwZ6L2PT0
EoUpUT7M8rqdoRrfKr3Fe2ovBZtFk9GIkZWFHNexPfYWtzy5VCp66YHkSALkmQ+SQQmB8u4u1kIz
jQoNY6YxuPdSTDrqJATIw0XS7o8/3c5kR2osY50UAOAbqWA9q7oNSwT2MEbboY81fiRIGY2ebTGq
Za1+M518D5luPme//+t1ccAaIyDmt6RauGe2MYKWeXdYmRMt+ZSS1joCW2m69UpgZ/14Q31gUlhE
Bn7AS5vt6m5gytMhecitXABcrSc9KGbw5icOXgseUQPiv4A6M6OHJ0lKdXfHviyXgbwzaKrZyKMu
bVHMIRSdxXNqF7+YPDzLjjUprgx9U7RvKz6l+GAp+wZKu6d38hzu73N79PsutZo8sxVKWdgqfTy4
7ru2HyWmxXb2YA/jTqNQqe2znnQ4A5nMx/HNfVYyIY5/6JAd2IFXTRBUk/KoopTHOteDaKPQ5eDF
gCwlYdLgJA3pePLmiM9UZ88lAibBGfooxsl/hJ4Y7+rOZo9GZjif9GpXmK6Q72j5/Fy3RTC0an//
7XhvvQjyzGOihGInvnu6lnCERv41KfcbYLAUiNrHjsEfQTFxn6D67dtJIGY8jyS42Ekro341be28
FGDwbWK/K5ysPzFOrapvnY5b0DMaiESml1ZuMnSb3VV2A6wJUAmNPyI1RaE8eyPt/lg1Al35/gvO
CaewSU4FI4GR1orUTosjS6RVeLaU80BqxISyR1XkvCAtWeitbEjs0183HPlgkDCn8RL7hjzDK0gc
NHjIECGd94mmmPwo+O8Gxfg67F5G4GGAH6/T7acIrCUKnPbasQKDDVUsoG7DipgUaWOxdz1HdgLg
fqs/MIDfHG8OqEWQlCCWZER1U8C+DmTijRzFBIwKj2LqQigrJeQ4ymP5m8+2jQDqlhWxNGAqpyEU
I3Y/srZa5CiI2TaZZ5wdUUX8SHWSn/e25g2geBpmBEohoKJkoDRgNTFw8OFf+npWhmBNy8SEM1O3
pvIyHx8WU8CbCRFt4jndzVzPbb5e8o75bFoTDO7Gsk6hvw11nKzh8qjJ/Bft/Fyrpzb5PCQS8W3z
nDqR9Qk8tdFZv8iGtz8xNCEe+l2VifVID7cDfXuBwOKySfngXpkCtLZKTS13jjBHHQnYRuhejslr
D2y/OAISI++d5TOY46mrA+h++p//8oXJHbEe9ppDQMuTsaAqJ9oY49UN+y2Avm/mkZ6VNlhRaYeh
1N4wF28UoDJCgD2b58XvMz/hwHuSFrs5xGwZUjOhFKwe/A3YYWh3gb0vX9r4p0MF4OP2JYKgLVoa
OI6wY4kqp5zSEAVsDH9gxVinh/4eluMTCuN9dRcmE7nbG8DrrHiMtJwb86uyabDOAf1kckpzbt16
FmKBc+0y10d36/kNwWvG3iQn8KkgLCpJuUpngfSF8Bv+DUAFZNkSS1RDXvEExfdZKgLZTItp3vs/
x2iDYlx9eUDkT+PX9cLwlOOxliBfOZlqn4YrrctM1eVsLCEQbr2rYTWjFyN8Xpdjlv0XNH/PJ15y
7p9CrMLordPLdOThQoXhiHh8+d+rmnMlzAe8le7RbqGppjhytyBE9MOM0LDg92mkCMfOiL9pjp4j
OrhEn4jwsnz+fblzxjqzDm04iJFQY8tjfsiKzKpjUcBZZdRzwpOPNNDBgc+TgrF954+CVABXg1U8
U0kucKkc10qKlAd3EpWlQ2aGoKZ1S6S+jz9U5dmEwOsQGn1vYCOqaT+gxOL4UgumCiObz6h78C7p
uFy5IJhm1bdyk/1Bd4Z2qmFExaah7k1hVEtakeW70KEUzGnQgrVmRr0Vgts1u+jJphc6XMbp03Ku
mZ9Hvo2sEWjbCmkXieB9vawGWLn7bfl+EU95934oMdKjPYGRRMLG0ENcnRVctK0E28lA3ooS8IAn
q4wGh47zPXPW2d0n+b8Tjr3z62e9igkZtyoHvSyjjXr1lAzJIbx4zmc5/n/Q4qOqX3A8qPHGL/eh
8jIMubiSqheWJdVOmQzMdjSSjrOFOfHwjMQdabTr8L/gOKzBAK+Q1CnuTiSSsvFivhfYixJ+6Kld
Re8WfmeMi5SMUsio7ZC5mMJhdIStv5KzclSER4BdfjRU2nLyclfO2T9cZrHg6dnEwz/MpbzKDsC5
JHAFUi0Cz2RIyWgH12hD1xZqR/NpxBRbFeGpu2KX32L9tD2yZws09JbA3co1NaYqdtrsyzSoO9L9
H6QoAT0JMWkaAeLy4FkWbO3hDCF+SK5cNK3VApYK9zXnmSql0XXmKQwy643X8j7pQc8h9YY27Fg9
B9DFfxTYoaNs6K4z41nbNqviQnUbKBdbn4lLaHuTAcjw5/6kYhcVXQP40E34lkFR90P1pRcnw4Qa
sKe88St0Zb7ftYcZjWB8wNiStkAJRZ1cKAkq0cAk8lFkudVxtT2AhYYYTuORld5NtxBjSCguPQQn
C0vWNTb6Z6JWuWrrhpxh2fAp+MEQBimnYLM2lhOKMtGsiORN4Hrjqd+fyh34poaxtlfUd2b+VDv6
k6h11Wh7q3rkk0CAShyl4xbyBV9jYKq2J78R2KlAXpuUClKZ3baVG5EP6p6+srM/Uzh78mpElaEN
tSzv5ZT7G4uGuJKJR8z6yx0FenQdeQYv6G/MMyeasWCKUq5zkQc+psn5zXi5jIll3UkcUMMkN1zI
+ImqAawgr6BRrLzTWVQjIWkovu/iwLBjWF1/o5kj5zh18Y/5VnOUXILq11xRB2nFcMXKoi59owcW
RjEq6mMIX0gOZWtDobP3KMrvpTECHjAlT22+O14jCm6e67nVyvlnOMZVZFXeVM9UFBuMRt84ppNk
70Tl1YSgDKWrjOSMvywMZAMc5kF00VB+fFQ7Wc/cLHTC4/WRZUCXo6xDtVdZFwAmihm8zdolrsbV
9B+0cy0Sq8CVRWnk0ODhZdkcKQpAgf3bHYFy2RJXJ4pIjwxWAo1MqWSVC69MMX1yQ17M4Q8NiH3e
Q6eKQlIXXcNVpLcqRyoTKsPiBYXpdzgZEBat2kv+xL4dRxuL9ZW8Pu9w4EVfMTLuQQKgSI9OTD3a
Lr6ftjc2Kvf3/lcKVWU/IsifIz5BpgTx4D971muVgbq0y1QeVkyhcSmxy9v+HkaxVBxeGgNSssHG
1YILLan8dXL9aPQC2cfMwsGugdyWt0U5jlo4aIS6xzEzq9Mm6MMHFXbu5PXuVxE+yWDkJ1E6wKPO
8NESQNVjkNZvKJFj3PM+hHn78khF/LmvoRKsjoAGpMx2OtcWZbxBVsbivkSALBvYGz/CCixjOeM2
ViQHMaPbnstd9lS8zixuOos0aU54tFXeYP74zI/Pijmwl2oX7o94qxA2uYztjBqIOZetZ9E+vdZv
Sm/eBK6ILQ97W/mWoll2PsSw//6iI38DuVvOp5dvz7TEdTVQhriEpk8z0QVKdrsOPCg6fMqJVjik
WQ6awpU4Nsd8vSDqCeis4406RS6ND2YPxhv7T3dNy+UeHKT/FvVF8WKWw7hM7kcA70kfoZsVcqF8
IUBVdThPB3tlQneTXZ9wxSwqii8p7oue8001Bi5ovcMqcDhBqY2mr+Nu4IbXnwsc4p75HlKegeEh
cB2m8y8nhJly775hRSKdaWhsVvjyL9nfDnPA+1fyYkk2yVzosULCpudd+gHIdqftrRR4r4YG8yNL
hganN9IAArHjJFMYR111Wy721vHuKv06+PKiSH6H+n0DZuF5narL0ikThPKDpqNTSCUP5jVDEexC
+FSzlgHgZvEG2Y5TUJadVcDU1oqgLgq581V1YZkunl0xJfBBPNxOWqFqN7SZgxYZpNbqamV2A/p0
BP1bJiOOrSR5YOuUtO4jYFwSYPcpYM7tmS0c7RhKpCUZy6jCTxADOyUWHKj2535rMzpj9hjkYdC6
0ZKcbxrthdelDqXeDlcf1INtgvE8CGHTVpXU+lF31vqqKP2zgI5uoTU71FXUbesSbdEVDigzGeXw
D8T/BlV96fIhMQQC7+ldyT1X+wREDZ5RESeLSYug001eMVMsq0EvynDXOHqApy7POhcgVSv29taQ
Uocqt/KYWmutljD7YLN2wJQa6tpzgedXRbXMGWnJko5ILLg1plUEhRDh2ohY3cv247Hq59xLZUSb
q+GNuzUMvsAO3nwoy5FtVIbnMN377Y6YwSNdEyCPc8eg9rtnDLDus6tysN0MPUMZH4Q2CiZH7ypA
trSkw9/GbERaEZOYiPxk2gS+aukQyS+eXlBoEeLHePw1tEk6cWPx65rj5JH47a/gOGFrugptCQdy
DIqo3m//tP73vvgIFy9/5YYcRrEnEkMvmRsK8m+G0eJf1nnNjYv+cEVgcrGKw5GXC8qVekqTi2q9
ME8tSonr0AOumHJgFJoIoWUX8gF6zV5dJmD6q4Zg4FrIAvDq8OQ0LI56eoujdtRPjg0sxlaWLt9H
4wEyWonh2zdThER9EBg152Whwr8IHNCALCdF+eRgwPFKkDUCoFgFClU8ON5N3NJ9WD3H+MkGwa0A
BWKshAK/Ws5hfHMi6HwtTtpvVCJI7lnKFthlJlvNpN03LvYV4GZTS8atHMpO+A/tfQ0Ub0oxVZD4
Ddalk79kxnJVOiCvWM4KHxAh5h/AMt1m8UCX4nMNjEvtElU1KvH/bHIBnGInv8pO9mlghk6+npky
wqadzQIjC7vWRqEQnWWd6fBi0bmQOSq12sQjCtYE7CP32lzSvdkvwMgwlw5VnsdclKBQHIoXW3yR
vxr+mB0TuDm08DmhDVjCekLutJXHhSZyuNtC4Z1TdApxMuvhc5DHSoSRb6VjQGhiREWJZhnPcUOR
DiRKukhI/zQzEjZCoxdMHzRBVmgRoV9pvwAToHM/hMfrPFxBUpokaVbsviHth9o3frWrtxvmGsqR
zveVpPaWm1FrQInQh+FAhTCuBH5iGFx2YIBnSREasnLMA05cleF+mOkQKrr9xdkLX0BAAuM5gErI
HVI4mL7kN9KfrrPDDGtYztNT7IqWht3bbn4g4WSnVdhopMTPHSqi5B1aON88pqHBVghWeJHycwzo
HmMM3G8bREwV6XEmQOST6G+a0fOomk8W5wW/AF7raAAdfFFZqVvv2oQeRbj/dn4nSjsCbVXqi9vJ
ymDZX8kP7RN55omWa5Bnw0Sq3VRw9BhSSSEA64Il+ig/D9o9pfB08QD55idtKeWxLlfuqIwq7Lfm
fESMjM6ZptWrA2DlZADPyOfgDcLQPkIzvJctLiBH3E6YvhbcdyxOPeYbwOhKMKebNfxYesYbZuDZ
4pGulPIsLQzJZeiP1RWcYnSW5q/GP6Feg+7iugkDjpDXEap7Z+eVijdWzYM3GdZts4Rmw2g75F9T
pAU8I7XFiTkFcRnZuLyGXIKuYltSVq0T65Rsd3YoopKjB/5zALUUywc5bU7VgqmHaz/V+QRWTODN
Vy9CtpnTF9CozrJ0PfiW86m8FJF6BYFy6XeNymkleH1yj6JQqWFk35p/QR6nyuoCaIz2RK9YENu4
+VZV2n9BiBltjUftAmblfmULSfxWeXu7VuV7zD+5hCkK4cbimXDS4smsk0HT82vPOOywhooUJUIO
KodiCAlTyyWBlg/kLYoo8H6vmcRLrbbl9IKXY2Qq2BkEy3kWFrMoGqPeGi/ZqMUDfT2rg6IKD3g5
kgA22CJU6uTJ0I5RphLXomrOi/wtAxOnTuyRhBJdjGYmLn8Ymd3M+ATkGKoq1qK9ckRUmbekq5SY
e9wO95mfOVvEOGO1eNlQ346aJWDW9Jhl03AE7oe7rGSGQzn3giHzcj2jshcGIgxX+3aS/CqUwof/
FtW5iCYsCuiaXYQvDcr+id/wRDSZYU9kwvby+DWlJ6ViMTO1dAfg0KcTH6sbQoX0CCNs7N2Mz/ZP
VaLNBIfe9VXZ7uEyZFb6gHCkHggt6jGts/sdO0/y77Fose/oZM57Eu26mhibSnNWSfOhlXJo8vcl
/1Po747uAFZP2SXdryXlci8jcYJneinJDXUSrKpF39DRcQILh0MRhs+nRI6LmSl2K2A8n953Xzdl
rRfOyn4s0VVJUeYfRGGx5xGo+wa5j8k9rCM9AVoBldVE/vf8C9AD/aLwKzHZwJT6URb9g43e+IrH
OGvqY4CirWZgDVY3iDtEuAWFNOfL80nqSAYdio5BWo038Ixg9E1TttH0F6pKdehtPhS26O1+Byq6
GEqYjta/U0JIfl6lOGnv6+dqTaypaw5PrI6LRuYxW6YMGnn+AFOvYF5E9Y+fG9INhvN2f8/07bel
lnjdxmGBa67LscBBb8Hjgp/nkdQBCZQMMUxPYNhxym+SiVfAWQD0p+GLvGDbSatIvN8Ti8fdQWBp
MJYBq+eam4zM8LUqxMA8WR8qezYEIXXhuwonANk9/RdLT8o39kUW6EvAVc5OIbW8EgkomMM7LMXi
XvHR37fgQzBqjAlxPkyJa/l473vTTlGWNTwAtyt/f4DU1wbMdIC5yrldGjVrAb83e5m0TPeDqhB3
mbRL9A/ltdrK328sVVra9Uli0UGQcTaTx7DRBZUzWbwZN2hnoSOZ0ZS4/ffqtbydfGhoCrw9Iquc
PuoVdVqPTio2oRz8jVPzlKiX5YVJ/y9xsB34jR75AdMP2EYPDxRCJluTPc60F6Sozm2fVnLr7C7I
sOtr1J+2evkz3kZActmG6smsV3eWTZns4u15U9GpgjPEIOwiO7xxf+5B3t+ClciKB6ybvQ1N/GRm
npWVGwIjQKucko6/fVtUcgjoFvwSKyhVrqxb7B9SYVEBx8Zs2CjLwUIznPrYpZ6oQRFUSCB36hfh
ugWHTsTN314wDax3v38wQH0ZrVPDVzJRe5ipjoJKj0q+Hs/OIuw6xa5WvVI3PoXCHmoPklh2Gm7b
cdDMjcnvvnyVnlj//SekECIWR4DPM5rNr3/jhQZlDAwfGhSBHfZRIfhGC5M6OkN/1ikGku6nuAmx
hfTvYWa+b2i44w30h5g+cfykKifqpHgduTwGORssvS9Z7OD/huj1/W/Vq+/nDflskxYcbfqoS8pJ
2YUm1RJCYIDjuAJyYsj1AUrlZmkUphTfbfFescFXTP903Aub14MsUcESRJ4LhqgdHmjxyVGWzk6+
1j79xvs+FEaB05L/8ZujD45LQqa9hV4knO1ExA9UnrGXQWEGiJ7d20mD6m9hm8Aos8yfocvjXjSk
1Xw3TWqj4Nnj1UZcX+ZT9CShDdiDwBeZ6B04fgE379tm6/FPtu9ri3/ubX0pMnJN0wmgVkwD2TE+
d2Fn3rrLZES0XZtJcOey/lJ3FpjUy5zQJGK2vu8uVGWIm310jFpzCb8G1AEhzAzObPydc+fwpqxh
62nQlbf5IG12+IoRWWH47ZjfYezyXe5QyC5+rKEC4BvDNMZHjx1NJp73do+ccH9jrJN46wrsLzu4
N8FGswwC07ae63lKt3qGXJcYOgGecQsKVM3J/QWjQO4zpoT0Mfbq1KzMt6gM879atDogCyPXNDl3
GF43oeRj2k6Df7JgIWX7EuBGn60wYtdxX77bUFdOL7sqwbBE99QmUN9HXEuyZchvMSKrukHR+O6d
769XbZ0bKgJPH6nFvLQEWXrDMIpG/J9sb5I+wMX/q4BrUjo1iYrdWOomT9nes3z0Ibq1EpBHBmBl
/GOiVrbhaB6amu08EtAdBlK7Vv8DG3NOlG2/irMhI5DXxML1yHHEfs5vw6865X/reXWZzk4h+Eoh
IkgkVLvI0Rx/D8DbztSV9FnvBzQJEFPQXgR7Xlh2CxZZhvpcdOAIQSaiNjGnIy8RZaGdgErBgfnR
xItMIg1Gv8vvBkLvKK32zwk98js8eD4oVHEfB9kmjXoPlY35zrhVmAyyNp7qJkioI8Jn+XOE5CY1
6/gltNqGyoFBg6m7NlciZO71+b7hr5GQlLI3GS8Mn4qgPegOP0A2vrSk6yiIDyzarO3LqDX8VLNS
gs1pSfyNxxqbXSEMKKdQFFdzOyS/o1+igAEHPUW4CoP6jTGUh9+mwkjzqE4epLW5EqFQh8RtJ46X
EVrZoZd+4HBnyvLxMZbkYeSVnNjqGSawSrBV8T2rXlsYwKZbS5orw5taWfVa082OK3jnpBf9BrQW
i9M97HzzUc/8H683Bzx2V6DlAb8OULQ6h5ECKm2WVZEiM2t84RSH4Tv/9m4X3GhTUqei+XTszNZv
x4ZIVhWWgP6a+MJx62srHEAR3KJu1+5K3D85UCYfU3XmcOJ1/f4xfd1GYoJ1KQcCat9VboEDqAsl
945BxOVWsUQZiS0VjVUifqj/42RWdI8Hk8KTr71WoqHNJHmJJ23LvxU2f+J6GeqfHQBSCSqziMVv
J7KR873sf/qWtGdzCT6k0bxTt00bToQIZzoEek0KydbQ0vOPAs/kJG7sJ4eZmfImdZx9unnptmSZ
rFny25ujzwGaKVW3zhImWifJDXJDkdV3qqDYIkFAGOeCZFeudWfVFVIQxpvdCBTfSpmrIzVGqsAX
byu1hnGdhfXwe2dYEtfanhJmlpXezRlUdtMYqYX68ChlvktSGaThVp3QQWenQbqZLLv9W5aSMEPc
kYe+oS3Dc/qgIyDh5TjbE9YUBgbHHxftJKj/ry/ctULQYSOeGXYDByb6jVR990mM7jaillfwby4S
7XNZW7HkoHnC4JhyiWtfWRI265vlj014knaR+v+NjFq1eNFIq0R1sy3sQYiQAx7OLW8ZkZjOcl/x
/w+QSW05Fk+O1n/RMGm51loVTEbpkfYLXVwfJCjicYNVIGiVfgz+SilDF7B80z+CVozcWaeHg+zx
6AZaikcPKff1wsPmSei/SYCo3/wPGPkKwSXklIPGQ/WQBC+SZSPQVB1v5NO32ioDlKXmWFSIUgX0
WAKDVnFLYp12L4eMpZ3bA1WSiBG1y2FTql3p3bq8cRcfXnnjW4Wiu6GaXddqDi1l7W41racbI5Pt
1miHX0PvzsbQuNzSZTeIfzKl3yW8T6gY9dteEh63LsvlF+GPpPsCwuUzfq9MnyRr8Q5trbS53g+T
QgFDkKmzI++3JuxVYp+TA7uh4uifvjUXtOl+mL/xl29KrbekvbzA0/ojrqzIzZOjIl7RNKMSoPYy
3qJkobXJBMsi3bnGwP+X7GWMz6KzX3Gl4EYwjEC3T2O6FETNyLfqYhF41+RNkcV8siM/sJh2n04p
dAEgRyT+CbavTUpO94IFXpDk5ArFamlbfoQ5/cEv5yGqooqc8Lb07whr4dYBWDxlV1hcjwcr8r8F
dCUI+w1+vxwl/LPl64KKlh33L0SUZah11/Ghloje3y6BlaAlEnFjhZUf3BJxxWCnpkSibrIW++hr
+RcYLr3kRlHS6GbctakpYido36x5ZFjpWnnnQOFPgT1NOVO/H7zSf9gsUtR9GRskZ6NOEIz+Z2uj
ORg1Q0WdV6v+axZmuZG28zbZ3ARXM05nl5HWU/frVXK0bSOawvWT1goYvvHYWNA2l5BuGnZq5XP0
Q6ogn6e15lO42nL5uqgINrQxKS+/+YpyxmiiQoVD2RvU5/cS+8wxLYOEQTgg7Z96v+fagveOmAA3
cmNG8zGxNH90+3B6N95GY5MnnqljmoJzSSWJzQLL05o4Vo5OQgjiIPnN4K15TQE2UKwM/2lxaoeF
XYbIAkQ101ucUpGTajgk2cpL2Zky745P8vYONCdH1WHLsz8UsTNKPTG3B4xEbzbzEpdsZ8ZTQWAf
oqo/tBjWOAPqz8cF1GlLKAbKZaUr/OPoeAD8F8/uyqo/r7HqNEDiKaYNDulpA6RR51p6Gq0ygG+1
2ubbZoH707GPxFt6TAI8Hd7dk8j4PM4zQTvhvppupJzt6o+ytyhoza32bfnw0sCYp63/Qj/H915m
qJ+bMzTfPsr2pXnwo8TPkmvX25gAfDQ3GfWARtcMOxmRWE7uqfFrdAG7v8YFNb12lmwp+K/AEuMd
jGBp9egI9lE1WEt6RknSse23nB4j7GkR2wZPtNXVSBtbovKR3oMNtaDeLIr91QD6/01wN+b3+Gp0
Yp/byb5A80LPvRKpVw94d5fB6BKcbgbQcfJQC3JNnI8mcsYamLJAJU2gzyLV3Gpj1fMpxZ07R2JO
Dd81hQBtIV2Q8IwyjP6GuC4J2Ng8hD1CzND12qrOMuYfUypfjG1EiGChnmCI/N0CVCq1LqCuwGkR
DBgQrY4RWXgnNag4J1GDKXQotehss/Wbm2N+yt0mrU0ZTp9GsrDLUo4Wf1/p2IE7ngEuhxSgM7/4
B4/6GfapeZj6IWKQum0LJ9Vpt+UOIadycdzfr4EG2WnRCaALXADCHY7iYS9EhaDy9Y8v/LKU8mQi
yaP63r702dJGif6M2PbnSQJTNtopgZbuP1st9oAQDUkhQ4lnk9HcxaxXege2ZCLW9FFUV1Nmn1fm
nyx+Y6eXkop6klEVMp6tzj2g3+JII9lo17c7c9sDlUCJ1+Pgc2iwAZ8p9Emw3cH3d51EJhCysxtE
7zIY3IcubtjweodxSPqy/YOhtSMW67O/BoFW7CJqULhiI638XaJTMfe9YLFiN28FzGvCuPkRhRpE
o9A9tKrFvRnkqeLYQiQYBghPXuKAdJtzeHscORbcTuKl8tjcNG5Ez99losbUAgHbUm6lAtj1M76c
qEgq/kuZ0ssPCFkNZVJ84UcHwLJtvA22vI1eFpFlVzlx5ittOPJYBlOi9UncJBc/lsSCAWonp7JE
qmGnHAc3cC8JUEM7kkY2oqe9Zv91OAjJavbdyDA2K3FZwST6hunOap6pOmbkPjKPaXAUpvVuis3I
VyyElwXc+BLpWfF28xekRBPctDH9fFa+w3eq/6P242uO2BbXh27An/Khu3TEfr3e0aEv5o0F7muF
EH+jhIs2hcsXdAHIGZrXGpayCSl5I6Li/qCaWZ8JFjjOuk3R8O5HqgTzkNjkxSZgODBNOcEJ29Z1
Y9DKNTXY1wQpjxY3CbipB1/wQiboYcoSmzeTUbkwqIvlnYbIbCbDdgL5bWVhxBUdpxJqTeZOqjB3
e3gwT/acsBRIeKGQ21Y4/ahR1mi9NwhucSodjK1Mb/TAN3e9KDxSesGe8rNdL1WXgNYOAfaMypv6
Ues5gMxlJC+DXFBQk+AJhqVLQhSIchE6izhaZpl0vKSJe6Jub/LkaaCtnYoJ+Coq1z17jCky0V1R
6N8kspKImnlQCZeEWp180yX3tnnVCCUfuQxL3tWbZOlR4DGRLOnHbN5Citffp/pOhzL6w2HBMhlB
x4aObct8HizpYXha3SsDrZIom/FrnViVZEwl7p4BFZutg2CEq+zNeSjQ2H8fbrCJt/CMLkWsN+Ok
GT9sI60he5T1Yo74DotQUWYZJIxA7SXjwI+6dgAcUMCjdnkFJNLRYOjM10n4YsKE45UuCWROkfuo
rA+svsXDp2NEbuZ+NcrOa3AyzfCg0EAZhdtJ4tjYrB6E24rPL3WG1LKINJTDYq37DyJjscq3N8Aw
xxiWylwyRP9TnM//UIXb+bVXssYaksH/5dmNOq07AVyR8U6/+29aL4a2mWQMG0igc/ilGafwI2Z+
wJ7nFwpn+JI4wn5fy++6F1YLDrRdTPmT/mnrjEqm2BppjD7vpcLTMS2eRiORVRGEi12MTcurYaEC
5xKMkWWLLoz7brEUQAUBK5ZlvsIAOK9Lpl7B39bS7ZKPWewk+5aW7iRf0ysQ9J9WEuTGMGSmksqf
GckiODVm5XRhKed7ScflcjfzEk1Bo2oZSyRogR1zneYYkAl3tw65wproqQ64jXVNyfNZlOqiPVhL
GK+6jEMPYrpu+w/KUQGTQ5OF3a/81BNmyrMGtiGJXJG1Zh8u8KdQnm4nOt9dAVjFDfAav9L8s2gn
Ocspne12tbaXm83i6IMHStgIeAUW5vI4PQMx45q41e7phg8AVtzWo7S6xV7/Pst65F3MH4xpWB9T
DPFIv80gg3B0VdF90M4IeJtl0RGxNoqUNyB8RZdy9ZA4WpOYhCNOthE9/rv0cLk/WuYaG1ot8Qke
FGT5zHHJoFx2kbPhXB5MiJrkUoee1MjsHTZTm16IjWPwDuRv1x2w6/ga+ypOX4b0Ug+LjJy2w2eL
Sc/HjMXn1LrAbzWAubE0cHeujRHcBIiKBYIku2Z6RaZUof0HNLaxaHw8hVR5qN+KbT1RgZf47TK2
l1/Dw5GtO4cpFm31cgH7K7nxLyWPLlAhtN67Ff12uxFh8zUwq9o/6alWpPDggfKhPbJeZMnBQLWP
0pxZ6H9xZY357fWHj50KM1Yi82QWjcuTfg32d6lUXQTiBDj4qSr9MComojBv7Zt8zvrSgDSYvLKk
ZuLTF0Ykdk2ILWH+2nvlsAy2oAnXBp2WZWN+PFet3oj7akKF3wQ5C8l6ciKqNaaTgBSgERIsN5h2
75wJfV7a/JVx61RTx0fbQ6Qeb7b61VVX1uieCd/J6r4papW28OzHPPqsJKvLymZqdDdLXbldcwBw
FtqiAMmg4g16eix9r3Iv7MtuRFeNt8i5yeH5c57LD3IuBMPK6s7HkC0kJt/7iLzK3C32eRKcba6p
ACALtxWSJJG+JKEhFgdh81OX8iICceeYfrJ6utyAgiY2PAZnKOn2mPKd61dcoc+LAi+TgETRUDQP
GVmmIBPRgjXqZfikKlsoCBQ0KEzL8kt2OUcBXhhJJymjmqAf+Yck+K3oKv9NgyQllLdCroCGi6Jv
15NUGZj93XqJEuJfdVbTYCzALWp3O23UFsMSgwHN0y9/7PhnwLkfbkS8pQSU9HA4AVjXxfjvJXct
JRGHkp/AvsAr+4mCBsDY2/9t56Nw+Mm5cdekN5F1J1qC1zNALCCbiPAU+DuWt+I961IXVWVpb6uV
RkVyASw/EA9mbK6P7JlcBjtpm7sF/5G/hcOw0R3+RH911zYXF6e4HWvvXt+vDE63tbNL1RivQwTW
OvpGE/O5OTTbysBPr2TdS6TWi1EfBl5R/NqRhwYbBAlRzo69XdT+sFgW3IR5fLEiLUHXIXRY4M63
dZL3JLKPrcyVofTYQf/URxpZ7yluPfvrOBNpEsq/SvfYHK6CdQEsnzkGVPAYDX/p/u2LR/FeteX/
wpzQxjFtszh7fS614kqF4PS5+QS6GFh8yrPzQkY3P9vdfEF1/Ueg8xswxU2EkAvLUyedPkrdbRI+
xZdpTIZBf99BIYiUhDpF3DBqjpjOGU/FIbpYvyT1EQ5W6DACAK7BnpEAef49dyr3amubqUuowxR8
4uCs14fY57OFLCFo+NNqPUSpNA1N03q+jMVo+LzrPaK42RUcMS0GX/BXMz7dWhdU8MFse6uOQ5ZV
EGRrQ90TQtMutoGPw6kTFk9r+9M1XWUJeVUEUu9pMOXbobxfdY3Il3wKFazxCwi9JQzCXjJ5MhEN
1C/J4aoBXArsAinzZRerUKO9XdtCB2aNAoDHrv5fSLUvTmPqUY24QRlmOfLuxsqrxlrM0h8vCirP
a7UV2XsPLY+yvY8BJdrHqSjgGJAEs6A5fBaTcVd7npZdPnOabBYGHBWFCGpYFDNsu+fPR1ypMAIu
v6qiTw5EyXbjTR0xZQQG8GaaD0fS6rm4K2kZJo8pscZI6RgQ43RDFySNUUisiyIRsYGvZAyvmlEg
4ETbqVR4MIWKkfKRdKVVNS9hfyFLgLZBJYrR1gWluXz4Gjf2rXpOZ5LurOXBdAoXLSk5rRM5rvtU
w+kg3GrGwjwLxOb4//x9exiVy+vjyXw7At9/M2cVvaEsNMn4voyxXfVFeJ+JRAj5AocSB6TtDL+p
+oAS6nRKhGbZVpPF6JN56pIw7vpL30RsERLdr5S8AovQjRDGA+4f2tQZt9pMOkrZoHYCy1tSvcH3
hC2mXr9e5tWJ7cB25iYvTzSr/T82zJBf9z2tEt9vlAepnf28otuNnEVu8C1c6QQWMCbSa16NkqVo
/3RUU46sOnqyxBJZqVzMVLjobrqGcRQ4GSReTO/CEAfBr1CiJ3pl0DFgYT/PJDabRBVb6rN8C+1e
IQsNssY+VDmloIgzrKgbda/EfjvT6eY7dRQMygdvsKgWRPsI7Bk6l7e0n/xvJViJGWxBkeGHZkIL
8D4oJNbr1n4Lis6A79TDA1AzafIvcT5Rm+xaFgqAqWMQ0h5RbyyFeYPywQB+B099ZTJBODOTf+3T
tJjdTWht9pO2iuCC/p7Yrf7fHM1XcJ/usu15yAN9uvsh6lwROe0wQ3ZLLkbQAfrkcRu3g0qGpeYA
L6aCGWXPbE26hYENOAT+m5XeawBtkH0YqxwfWx5nymkfSwDKQQU88XNbmjdWgdFRuAccesqHV9z6
I5AA58SONjquyqSOP7aMxH70Lo48/cs1APgcdtAMTVDcsQ6TlU5DnR/gSbmRqTv0MHVoU9nFzng3
G5EH7Fev/cDR01YfYU7IuNmvFTtC0QJhu7NSDxnc3VHLLbhYTssZQhEIREN59zZhSFNTKZdsyVuU
/A+9wMc9AEsUl+5i6evwncdPer+kUi2w/kpnGiyT7UoBl9OsqDB9Vx/DyKJlVY3AdZl0IdDthh6Q
xVafXucO7Hw+I/iGUPvCgfnqY988b4urRSwYC1jdK5QoII6JbR+Hxr82WED3dLaW5br7UglTRlc3
3GvaT6HSXQl9pvdPfOKkbxOqBj0at2ixLPpoCb3US5epLl4R/ZY+aZ3c+Jd3fGCRky20X5N126xh
TqoITR4cc+InSXLCFNaVrCbyUapmFDSy7coYF9150CDDUNVwdECrK6C32cyj5ZN4KBN4jSOLvvrI
UAPygrykOj432d/O56hy4btksPvM29fB1SroYDKOOAF+54V2szM9dCoVxiI3LXem3frkJa0VZUS3
kvngdRkAUYFLorLA2hCOO1h9QrEA5G9+DE2CNHCcovm6pOjvAnakNRHsTvroI+1jhedRgLyN4wHv
BhrL31+Mc89XaQ+TFrpzhJ5z924A3N8xzz0bZ3K1QcuJcCrcK51lp52a8TvSnfkc2//X1ZrOMqc4
p85FWN72QtnZi+CNtkHf194UdjfJT01JAAxO8FilDNoBSzJAxOTfyM1/GyfI7b0Pi1+P/5XNeOtg
STMvnv3SlLrmGeMXch/UPO7aMB32Nu2vGYY0iZ1ZnaQUYCFfsGKaUiMH/Z9kvAq+E5JFyI6Rw3j4
V7BzRTrEH9L0YGj3V6wEZS0y74G9+5kpWtke44BLBFuQnv19xdU1rLkF99DBUkXmAV5JnNtivz7N
EIE713+SetIKSWPKmPPPUouOnYLsGRVVOdN9q3M4szejpDzCmB0FLsnMaYsaL+gv9SIPceEl789w
OiWZqDXYh6MmQQwc0PbupWnrHfaw02PYqMeIDEU5J11sRHTT0YRk7Mo+QbrFpBzmYlpfBWFJKVOf
0ksnQWCu+i/i6UKFMDRZD0fJxwrfokehvlRSK+c54petu5vvKjflfwA4fS9It/oeTAvdVsxgaRk8
WiV+T3umErBvsqRlspBIQBas1FemALvqG8H23HbanrO89GCqpFz4Krao8lCsJvCaXl0gu4yeo04n
mV3EgHVU5tPpP2Awa2GvBtMLCQ90QaUdIDqq9DHKCmIBFQsrBXwQ5bJ5IqiAMkXKquTg00kS6vHV
UUIALQzFxyZ2kzdV0+2jAEkrg0eKHsWBW0yNmN8uBZP6l9I/7+GsM+icEFIqDmQyB+lZ5fPGCNRg
n8meMQSThBwGDLqZV0TmV8EiQcKdhU1iRPy+AyYYD6SBLiZ/3CU/j/uHxKb28TidOrY4Lm1UtEmB
pl8sxsxAFzWC1UIpvtX3wmy7ZORi5wwAMIbyKy9VbdsIFdDOWQPX2ACHH81gojnYQodKaHrhMgoz
lcPTH32excaGCU87qYwjlFEdoTgUGqFxERpp+A4uaSJhD8OmsU3DNTf6TLjr270UvOVeDWY72IUA
yTcM2s/fKSA+XEeLpB+SGjK9GbSNC+zYl4C893nQ04jI/BR+CgsZY6YmvnO1U11IThwBZ22PNKN3
Dm+rniTBe9Rc+hRWx8Dbqjz//suuGY8bLIVJZ1mS5+UKWMsg3/73eVrjBFbWQEcUWXtLzOYd2bcy
RsHvrEgPXeu2NwyHIqnz6MO4lxJnJ0Yt7KFtpC24nJyem0f1Vdo3JmF2eUq0Ut+bytS6cOIXE05S
xj+IvUK/t2T/K2FYQIZ1Je3/r9Lfl6v04zZfaLbTnVSaaEHul9b7ohQHm1De8k74hwDc4V/ZanQZ
rayzsdgLcHdrYrGuqOzi6aRIYwgwja71YMsjhs1p3gkTiR3YdDVfmqala6lAkX8hj17i98Mj1NDW
+yBWPHFoYiBgU2+WJNWbXI6UqeNK9O1jmujKE9YDnV7vGUZ+RJV68wF8RHpDCddonKN5knwBbDwB
FFZX+uTVuyrpgWOPG7vmO9wuj2VlcfAgRQYegRwv5F4L0IQsmA/b2o/xB5o8cifvWWr19oYzkqcP
nep++kBWX3Gcr6Os+S5y9agyAgucMyTUWY7g3FRI/8ZxM+01dNoAaL7AnKTL3YVOvxGN/jEuC/mN
+OblRaRPd9Obi7VTrGdDyp8LaRMhzS+laOcUTtWKLrfltuEkUsC3TAevw04Z/qLVYDEHt/1EuYwy
3nB2oG7uHYt0MFgz+1WDcBG0QVLYBBn7Irrj+Y6fHXY3a2v7hqjRxH3Q7FBBWd3FUSCRxzJogQIq
xsO1yUPOk3KXcVWGS5Eh0C+kDm2pzwLgff1722s24adPAqhWCrRCFXgq/e/PJqoI43EEVzMtlfg9
gcgBEquN0osH4jHsjJARlw8HSkzTagDYmsc3kVZLS/YVb/UGY8ivjIYO/+l9o8gt+kar998XHuoj
eL9ZiuSHgDCWOeFBNdNv3VFUA+4FD+7Zz7mJiEXtydCfyFzs7RbQm8j4auDocIWCfjUFGW1PeBPm
ES9l8n82Vfmlax7v9XD66u8GjExEs0s8O+KIktDUZtpN21TGTZY/895nosOPhXuUHyenWSD3pYj2
eE/CkQbvEXRv3d6zuqNo3NV0AdnA8klalalWb/3IOCRKC0alw5Aea09mGns6lG+1oPqkz7TEjsVt
yHyX6cYV65EqVNaHB0nQIIfUWqsLe3/QRK3BQcGc0z8a5T/HTdJOMS4DdR9HWSlIGfckTXUJFe79
p1E6UJSd94ULzN0xrXFtZoBPi/CfK+2Awq/jHVIIJXe7+AqG1KSKCwJHbPbG3leestVmS0EMdpjp
INPAcuFtX5dy3qEn3GKxjXl7ODyE/SMkeJ6ZveSLoEI7PKqUSmGvmbXdv+97NkIAHVJY3IYjz+7j
j+oakVZFMApcdabaxI2ECXsjVGGpumSNlBmTNKzmE/vnf6V32DwEvm4CEavzhCd5qP+OmWIRWdNU
IDeo+cvCQAWqs/YSgN0XK8KwNtckZZd+PL0f7BuU78lhhMHnk7HHWfpyPlaBmarmygkpXbcRcida
o9d+GNj7M2iSa0plNjWQ8dNuJKVQyRacwHrB3pwbedRof+v7qX6tSoFKuJmMG1LM4Z/+IY3XVnEl
sbMpmQR4ZfoTYQVPhXpHZ+5mi+6p7VyKPY/HhMuOUa4gPPd6aHxIHj/IWstwGoS3pZ29zlDv3EB2
yKFSb1Y88PLRtb1POl6D/fhgaUPRFOOukwu3LqdU8/KDSOO2Fya2nDTjU0sBrxhpWW1eGYo2iZTX
ZvBq5onCEIbAY6YI6BizQOeDJpMIIQdRrcDKHdxsaljVEmdXN476WAQCJcLw6bJIRF9HofKhzHk6
lQXFRoWYaKwriLWBT/Va+wPDkwNfC45CofO+ed0DmAjhlAQuoXIY8NBD9coKbnr1NX4rHptrFvdW
+vD50Rq0ehUkM+0sp/WIJajfwmgvOaoFjqx3oakpRoe20IU3xv0qPRFo5GUKLPaZehrl0vlFKITa
wNljLHpQEvTrElge6ElDQp0BBTPsvUdCcfGFqMDjIBgNvD8/Aq1YptCry9fYGRusVmaiWN6xuW9Y
CkGQy3oSVUcGBENMnpzDKOJba03vG/BtojvkpfZqywh1/zT4Y7mIyT0DeoQn8WoRLMEathiCYiO1
cgypFbkP0pSkAoh60Eu/uQu+I7pP5D6JYXM5PDuoZWIKipO28gqwR8WS8gkVKIvqNVOmgztQUzEG
H7Vveq5J8L7QuTD4qp6WtD1m3eksWXGYP8kh2mUdRbAckTY+o0J7z5uGqsIJcXeERejuHCes8LTY
CYEbxWD6EaHT8tjFiheJqHMKfv4gyp5QL4xTstOIMMKeDBe44osx2GXFu1M5DBVy5PY921ZehgwJ
M7KDGcxdR89niSmZ+TYr4d52hmV7P5iZ7ehtUSDyg4CLpPJhPDYgc//JG4LBYOPbRoQXTVL0FNkq
p3Bj764WpTURxfTfOiPCeBb8RW1VvE36bGSbN+qKEIMgcGMBUKr8nO0O2AdH3El5ui8iJ6CfgVxW
OmI5sbsd2plS04kUGwgp6h0VBKQ1g9sWfIThWDljfddLpcEtlDAoGKOPh6qD03ePDBW9Nn8Vv+LC
ia2m84DfQIpL6PU9t+913uWkMbkaNmo2XEG2kze+j8j4B/is5Q4s2epojLtknKEQBAGGHriVhhye
dl05aceOdQXZiBmIviongrcERRteAlMHwcBbkbIP4RSBj/x609lyn+kaoS9+Vy7DlBJcPY2O97Cd
K1a0n7kQWeNBxiPLMklZnZ6HkLUyeFohCedOO4Pb1kmAEuHxoCmvDARA6H8Jn6lAxDc9z8y9U2Z2
EFCBagP95d5fK6nngKZrw1Ocnh7vX5w8iV3vKZKbXUje7gW8inoo1nS9BeJdvJzF4bzr5h8eINA2
7nrI8z7IufDI+mWamsY7kmQS+h6Nv1y9TNzntTGg8BBvlngCM0w3GUrIRX13j7BUpsKBcWREohb1
TBiQVsOdXPtinzBKPQf/WMrfstJQptQ/sQJNA/FLH1c/wb1L1eUFDbjH4Y1T6FbuimUsst0GctG0
dcgzEJoNTUWDmiIH4uiJ7LOJLrmWr/dGzdN0v5l2fd5g8tMF1vcuqj3BrVZouFwVELML+xU=
`protect end_protected

