

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YWwSN+9l5ahBqN8tuQHA+pe+2Q7Fh9//dR3H5K2w3KRc2pla5S5ifvTi8Ak4V+dzPFwrZE+Uv4ZM
WqK4mWAaDw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WcjiphsvP4YifX33L+r4vrauIXRkGno8B+olsJNjoqAxagaZzNDAFnvGiJsIWLTLoEkntxsgRnIo
WVce53gFCvnJJkmdaYhg6W308/4ThcXkZ2dT7Q+TUTpvKAEe2vDwO0foHspYl4iLWX2KqDyY9jge
moxvN6KH420mg96l6zY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wvng0RPku5m5MHpJv9WwJDWJ8F5PUKDSPU7V99zR5erdP7PcyDhypTKxqOMHkizg+gEusr/QYxdH
b3OK1yRKUZ44xzg4dZxpsvitjqx51I8wGaS5oiuyKX8hGtgTVrbfoHo6u9pcLQZn9XK2J/iSrjf5
dyOg2xTIXw233HzwIrCKg5RT8dfxa+iICMhoGVZIGJ68DJPwrJbT6Swg5gWMje7MS+Ppwgv0Jxqb
7HSKZuEIyqOKVjWI9mOWG9o9+LBatVHO9cQqYlFkeCwc3YeZbVHELaty1PZ3GYbJhCtr7obXWCNH
f42iQcUXnPWhD7j92uOOj9mnGCfQwEtmFpOg0A==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mnRNLVCxq+sgQJhai+B5fZRsJzZ93rdvyaCrmwTY5fIgoqSgRC5N+TQCYgevu6oU/nSzurf6krRP
lHQ0Ztrjgg2Tj4+uhFcaWXWp3gef6Qsz8XcVJ4aB4xMaBhgkUeweDC7vzOKD05WXxyBd0/qZdLtt
lS8j7xW/2WXeJFqpGaMZ30TpyNYKEPbTG0s7zfxCOI79Vadm9yVGLdGkntvGV8guzxeaRo2Qkmsm
e1+jXsDbdOr2euBE7JiOnNqartejTWUhtjRbkQnS4YCtUcNrW9+ObOoPjivEDKhArV2d5T5dFhZd
vZIU/RR6j3BExhd071LKzolsdnCqR62C9tEZ5A==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
E6549NUXinEnqZcngO+xA/zs1xe2Bus1VEuxweH9iD+10PgNtRJtsG9EF7ZdZas4DjOhgJh7DHf8
ndbSlKTeJx/4QdIH6iyjSx9xrJbjCC8TeQlSsBzTcSKNDMh3HuElLUknuM+x5+UC+hkdrw0waGjh
tjj70YkP+K8Te1Nhfp5PHo+OirttOLZY7Bnhq7x3KDxVSyWnLuCBlLcRqRosb6oaQVAF5dnEKVG3
DDqNFX/V0KONWbfs5QSo5gM8f237iV+nwxPmst+L5casdH0vfnMagphcYI2Gs12f9zJ/qipttgTQ
46Pj/rGC5IRv5Z5f3c9wnJBWRVPQ0uHojBicwg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ogp/UkagRFxN6D0Tvatf3PJ+RNRc6aGWLVAuekDtCdp1urxgWDpgdUpLAqv4gVFTloxR/WYTIPAy
tqnoQwfvxF8+1H1sANWUqIMweNpcUZzEYS0M2VRPa5yH9GDRSd+LmMbbrq6RbwvXiR0tPlJ+qF//
xXzjGxQQlbn5MtTPwO8=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WS3NnUM3tGvHLrK1+gyTpPfI4oWwTOYDJPYfQBcc9ol/GaO7Z5AyMRqRkk+WEY00WrbCfviFYMzU
pGl2IHT4VRRzqqLR91kr2OFbN6OGXGirK/a2SoQqoRH7NbdhMzwc2r2DD8mzssXGs2HnjNYorDiE
Vs1axIRZ0Xwgll0Xql9UnW3+H+bZdCSjNWd63t2LxcoNPpatkn50Aa0uZrOTFNGicGTTryERIIjE
tD/W23CkHq3rM2LwJimtfOkZfT6H17TZIlmdf4GzYYEZqzxs/jkYFtiD89KMP+/WhCVPGWSzHT/R
ZumbUYGnUPG9wSLIU2c4b/c9CXNngT5yj0uIjA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
5VRK8tyLX+6PcAmXzZNd6xyYesUvOQ40FYfZYUSslQAnYMn1RI1hna4F3EAw5uoxatUsUmwO31yT
dyr3xOkhvzQZkVBC54XBYpL8ZKYdwofhrRVMSxKKdhfXHoqVeeiCwCjRAwvXEaiZvs+fV4QuO3Ce
AvsSsSaqeMBNXeiRnQrkNAt3KIrLOdWTrmlYrhNd90n8xctdvhqQ8xXbgWfLY8t4bw6QFYH8Mkj0
8OrsBlG5QM5QLhbLdK5sYDVVpOyUK/zh1pXM97qGxrW7lk7DUTcABJAa7zEt3JoOwU91RYu+O8LW
618CIr6l/OLdqfLbibakQa+oW13SzQAd8iOo6JQxTDjeAO6zl42S4kVgqEX5MY6jDzUGxC3UChqs
kuxvBqqcKp+D+LkvCspC5w/FZ230vgwF3ZtP/N6UUc4Wt8edS570IkUCMR706+v1FMka8zA3ReR4
0VWB7ipZzQRPNpfg5Wt3KjlSPwxzlhO3GZecx9964wNvMUWmanTD9J7xmffdZJMaTyjtOQiaUhNn
eDVEcZro+uFDlMlAtR6U8LCF6fSTasfLbbxGGWhMGo7q3UStAoKkhb1AgcmBmOMdpcNj/eyP+F6e
czAdIiCxRD6StrW4LGD+Z++BCbS/fOu5vCpRixmPwZEk+hsGcQToEhaUxkdoKdS/SPlfCdX35Uco
oXbTrt0vpoq9XHKyIKQUfltVcH9N91oeELR3gyrehd/P/+o+voXs0Lx7Vw9R0W3dPqyU1d54tvnR
6XXC9Er6P/KK1hhVLMKBZD3lT/5jv2dFF8ARqvQWhWXGuM5lgmtcvGQ1iuT0fb8PHHpqUlJRsHh/
JRRpfQ3xXryImKi0AcLcV1RkkK3AyjMTBWvNoJUJMc0Le+viECITDOYWolA0vmVzdEzXUCCSdq+7
ae7emm+SAZU1mr31p1LEGqLK/bs4H//i+xlNL1ycp50lqqth9M9UF3EjqnUCquYyFNCI2naJMrcs
4fYSDp4lB/Hm+/EfsrpaUqnMrvezeefao+gWrSsE5XaQZDtmTapDI8eb3tfUgmACiofeIZyU15tV
iHVL5DbRiJWWhHxFOvFsERyx+shsmQ+pMLNN2LOcmU+MnC1TOVSQsJsWvg9wAHDp7uaG1UyoRfH4
FLPJgmsPQqpVRMSrK2mXbFjkWQZzR+6Zj9xncO67ESmi9ePOI/qRJvfcSH/Yx06jS3+JO7rJxYOj
4sKclJVJnZqoQgFXKgpHnS2iL2cnZSoo/QtOXxOybfmC65Ss1r6FjabLCBgW9UN/q/vhhheGhpgc
wEc8go9CkL12pBYKWveV+ebm3/3hu5uG1JqBKyVF4sI3qFjyWr+itmdeCYsJ2JszkyYOBB/8DaVH
npOLxfO0fwsTNtj6AUUcjqjhD48EJ+xhTP9ucXERWOE4ZKvSegz0gDOc1AuAbG01yRfzh57g74tz
YaaFyp53JSmM6BfW7HWmzpeuMXcpEVE9V2ucMUvUVjjfot8Bsu+wx793mmJk+6VB4zShPuSsEu4p
2KRXeiRq9zOy+gDpC2o8w12nEZAG71BY+6Gs1wB9khue1GvkclQwCCUSNkn1ECaF7NWva6LHHQVq
GtMf/v3irTL/44+CKG0ZnH2K96wIIexatmffsTXHqxoh5Mts29Is3lfxYq5nya0HnadSnH3tHjRT
0TLCsV1WDp7zyZLsrh+io0lzEZXLBkxcLdWv6XAyVEQQoMeHxssbAfJOzgmlaRaePE6HP5Dqeo7g
1vH2NLLSDMUg6PVNZd4tP1hnXxPBMrhtUTsLJu4tuCD/5gpPBGKH1fGwh8GNvF08XXG2ejLsQyS6
8i79fYlRNb/0wDPgWKR4GMDBNgr2DMhpvqUj1H4LQv099tIYSLfLdvlPTz59XvlAYpjAU+H91/v7
vciNH7Hcr2TuxjXaFU/Lz03T1mCuj88+dymxKki/B+FVapF55vaK7cvft+Pmx6YdHcHSX0xt+fmH
3bCdfpmrsUxUgPBRsChD8Ptil/prAzAd+YJkwxGs3KdcY8fel/x1DoTvI/p2/NQFejv/pOx7NfwX
JehPJZBPjdBfv/Nm304PpK3/IZv5YwAyfrfyvINcrghnlV6K/ZQahKfmooLeoSO/82fAzI9Ql1dm
fqonkhQI5Fsd+fRoFRbGsevdvYH7mhvj4LeiO/9UdefF11qz9QcEtw2MWaDOx/uowjP0QS3HkIFL
nDeol+DOJBAdoREjMkhZr7MAbi2xANUdg2mvNfCTiv5YpeZ6WDa1nmA92TMMEDaDPtXtMLmuZ86G
rRkXfySQtiNkv38sSu0hhythIK1XhE6XoN9IQZi2yZIxdu2OvmJSSfad2whfLFQt2RBBmIhSvErX
+ZA6u94A4ZJPWPmIiprlssVMb94398CHlSnDkXkYI1q5XERsSlB0jAhX/tE2PjRbwCujIjaU7HvW
yjPbOH/KPUGsfeyaG1VOESDXGjrhKDOB72Eo7gnPI0Rc0GwAdMtqOJ5GFEruo4CwEkzjeoQu7sz5
ux21EcwhKeRR1+y3Qe81ULsVlzT4JPpfolnhMJYitq+OvlJ7CepqE+dOLwx7Lpx71cGZAkZRg0hE
UOObFDar5+/MESqsLWgAcMojZh+OijTUKFkJ9iaOZDyWaqHK9DBFsqo5RZthCXMGoa06q5GvnVuK
P59oeYsuzSPoXUt1KBgX4dz8H1UfTeABpdfCd42wmexyTR3D9Ryab6sJQt0UJdlt1hBmWb4fA6kN
6LWsB73sR2Qi919xd81theRUOg9wWHF7ANGWqaIl6T35La4ujJMzgHOoOKwSuceyC4lCWauH/xoL
NWgoVNkh8vsBObSKwAf/UtRiF1pxxoJSr23qfZiE2Bbejlg4aOVdIwrhnl5zbjct8CmWzvTXQVhf
LkrcJcCazm9BKy8VYim/QYmYI8PkVZSgSGLHV4/ZhzmGEzzsjRevxdjh41XNmmkmezbISNzXb3ST
8qhHSfYwuKoRNvw1+On0v58Do4Oqyp67I7bExM2H3b1gnKUVBJVZ5H7VV+76PVoR4N0RjIftYiI9
cXzF72PWzRBP6se34xl/CgRCq/12aPTr6l1qiP4JOTvUQlMet0XDyu2LQa6j2KL90ZppElGGk2jp
pvBZ3Kf0jXC+0C2fONv52AioDGUGPikmjNLUPSmfPebGPNijV2IP6e5FM/DmmRM3LmZEjNYE7zlE
EEkbErGaKDa/eKeAIu/9sq+DtlZYL8WSr2rIqyac94gBSbnzWy5MDU43lbffWsXa5oaM2MwJlkkL
66Vo5tRTj+UV4idA+S1XiWdh/e7aa3iZwkl/rLtsiHIJAnUQopVBkrp/3DxlAORxJxVJA/UAw7o/
4tBSuj00w6ygWEj5dyL9nrb0AZ10nQlotl+ecp4e3dG70afXWcC3jPFffhC2jTzHD0VGH7y9jNh1
UmYj3oBGkc2zSSWb9aqftQ/sZhmbEVPFT8iN1lAfCxtEdeOMgWBSqSoptXEOx2+qLY3DG2Ywn7mY
rgJcCsB/1bHZlXDDRCq8Q8CFd3N4uZivIwO7sK4E5oMEYsN/AAEAxkJiCz49xay6V60gs9Ct+TJ6
V9oaIj2MTRCPOWjK+VV9ooffRPZcK58zLG6CDxvK8NQifx49AcAEDS7hTLZHbRx3GH1jlwCQphFA
6Gc0gbjU8jCc6fHV9GUafqn38qtVn2QeU3YmC0MiVSKPYf0C8zVmLY8OfO70HXC8xHxWGBrwjgAW
viB9yS2eQkV1nPMTGxpw75zu1w/f8J1gDsie2RWDq2he8kFluKfU0ifw1XwGy8FMf5hHaAWSt/x5
DwQsVHUGpcOMrVZvTHzu3cMVgN9VFkPFib/y8+A2bx2no/3K4cwmkMdDjAixH48LVerDlCpbzvQX
OhD4GDJuI+o11iw6LqjScU4ONnfDvei6mZ64+C7F+buVX15jxKvGr7WpxVCbvoye0V+cNBM+YCY8
vox9xJ9QJ0bEJ1SJuEd6yAypch42vQiui7qQGzb7zVG3TNjsX0t7EHcxaCkeZ4xkrG2xwx9/577R
3fAsTgMqvzjKcZE6zoCazUd71S0UXXCJUrHXGcLTa8rt4LhTnm3pDCSlJLCinxqGqW6LYir/wS3D
l6gZGOhHTsZrMD9pVHJCMcoeaalCVRJ1o10XBMNnpVBhXNBp5DmHJ7aqW6U97fE+Ffb2Tu6A2vla
BVpo2M23SgHfNiKb769dARLjDBo/9PKOMh4ON+jOAg9fc1/Jx70fCR16skBbPho3C3BTC7XOGVaq
8wGwugLBFWqzkIN/f8VN7z5Lxlit0CbOyH6XTQHi9YlH65y4B2uhHmEOx1dnEL0LtO3hAHtaGyV8
z5exL8uSchzMQat8OwOhcI4MPYaBuphjeRcQ0d/5PsnhtzUnNf3dYNEnrZYQ8q0BzqR7iYjG1iJw
ZnwMf5WA/DvKaEQu0jKHz2JZbACIBzp6kWlz8LKKpd2+Ef4D87p4uUV8JkWt1qv10/P0eA+teYJ4
Adu+vIDLE2YbxUkzflrO48yMfixqAjqHOeZwj+l+t2N6vm6I/M9KAycalr1oiVVWq+DvO/QD/RCB
BzgBNY3ngNSfbV7dtC7yQzxlQI8Tqa9ZjXoER9PQJH0Obfzbhc73KwRKrIP2U/lb+qaTf9yOCG1e
mJdPzsRIHLxqYS6BDuS+OEZwaRkFxryoQe4EAp7dObaa7x6Woqa7XDjcV0q7FcZRslcz2eaNfIQ1
HA60W1uzJxtsPZYL/NeCiz6pBp0HGNZgljvfwZZvU5gvsj7aK8SpiulipZTUV+da2j4zf/evvMdj
OFRY1kK/EG87OZofM81Qg5Tw0sRMXiqrIfb4KHsB52qwiqHuOxs5dE/T+wQYX78BpPOfzOPEhV15
wbGEzeQDyv6OyduSE9zL6E03SFp2+ncc2oJGYy3xIIMr5hEL2WM3W/3epLc5Sckf3kJGcTmkJGfV
MdOnaLp6jUtbFhn1quLntHNCIZ6KcRANgn1qaYt41PMDvkRt2xlpApgopuPyFwa7A2XpYkdTnYUn
sZzLjX0uuOgiG3qkot/W/RqW6KRP6zLyFLbyIs9LMaavtbJYagFSoUY6TdVmyAVd/lqcfRBCp2XS
t3zYdG9HhefrOyqmAgXk7l1K1pEww8rjGaq5D/enjopACdyseEqr1ptMC331YNmKZQYpMzGm2/W9
gKGYFuZxoZ7pOYSeRLtdiqhsKoY3BxeJhZaWgsNN0ZdhbieEoZYCoXXHCl+JrFtM6OEtqXLsjdJd
CK09gjO8fWByUDF1dxi/JfJUAg0ZSfWbpjNSxswVS9s9FaDIleMiK4kCWVsqBE3uelQIBFGnC3Nb
cyf3oGUZDS4ULCdxogrd4ttQH/QTlP5YhghoZTnbneQh1+q4FIRRWfGJCNHKrpt8fxfgWgD+xtNK
ZU1+1o5eM+UPTw1Sv40Zgl89wNldechbY3V/JeQr827YUmvSfSkHOpWjd1oFDMVf4+U2vX/Xo222
RpV3HDndbU/maCEIBLzMuXNsOk0g39id6/sFumpOS+wdteZgK5HCBn4eP8CeC32iLenWQCtV5Py1
6QUZY8Flqa3oQBlMv33QLl0RJyXEH0/jLRA0q3XZbKOnTdSqvWvM8RieZJSAT0wTqmMIkSpV+Fzb
/bDXkgRv/ez8vAEa7jc6Fju6vZIsKuP6FJYFc72Q2c8aeVqsi0qDBL67GJyGavzuYwi2SBodAi0E
24E8m3ehZBfhV2YBPmvUN6w1PBbLKCesVsOdwqyptC9KrceQkXC16XbfLAvy3LkEhtEctHIyu/zX
hZli0Js5Ra/NnJHIDa0ezS2F1ykIjsPIJLbZlgTwAuDeqrSSYIPbPIOFPFN4DXreaU6tlqWq33Y6
dh9IqCnSFdXB+TtK0aEU5I13s7Vr3tZJmghNnUkK4kdZLgbUKHfdvvZ7a0fUO6vdvdRnaNnM4j2I
vmIEdop5b6Kf/3CrYR27QKyW/V6yMSo/4JDv8q/pq0MgMtj0nKvDIWdE71QvL1evg8BbCJCWq51B
Tj4JC0sCM/HsGaHJOHt7aOjyonuiQkVucNyfGU9WR4NvKxYAXW1JArrtBMeBWEpSaqPMUYKdJIGH
awq3Sy2TE8jgN/9t5UycmYFj2L78VU3JOBcP+wB4Eqd/mpuoy9AZKqw4djdlR79SQZlZFxKlNlob
GAovKKpWJkXSFtjvt6ZwLuC3Y3/tMv1Of0TcfQb6oOrKaxiOVJFyW+62mEKfiz9EKGhRp01cuedN
oyDpTFu0cQ34ahsgagMEtFUJDWq8+kf8AhQ1qSHJMrYoGsEGVqkmTJyv/YmRX9ZBDHfRqzDoruiN
CCjO0mBaSbHDbcWpIOXvhytUX/BsJdqyQ+3R+y5M49Mj7vfMvm8OgKxyoaMT3psH6QWRa3cXNf2l
MMccQ3sUo7Qsk2ZDxD90g5ywB4o5+LaVNZnCsVdonZ92m/mElnmZJ9Qh2yG4ejq4jRSbEK8NLhXZ
5Bzq0bNG12mIM7M7b7LugQSTqyKLkoZ+lRXCZb11MDKgLlaaYFwWYW0nNIaAbsRZ355XXpUGvZ/H
kCskis897EZPdvxbOOTzF0wxLqR69miAXMwFQmEufa83Y1Oc9iH3Jjx3ckzj3fJjZpRcfRw7Vcei
/P6Qn9PdbburVcx95mrOgelfwQVGgpIK2GEtuwK6zPLX9VZqkKYFd0gVauqz131O13+b5Oba6ygq
KODDZRlmLmKLk4TcUbB7h5GIITm1XQIff6D9755yLrcGhUVio9t7T3sO7SS6tg6hG0fWA55XpWr2
7tWAoZgm4tYr5XaecU7pNQrC/FjCUdpzSmtVYrjikCsPMM0WT0JDOfadvhMjmIsDE9FdgbjrPHs0
4syctQX+pycQ7NlmsIta6Gidmiu+Nu4ej6YfrjHCsdu2iVWab4oEwwraHSIUnGvFyYVSDnQOvhG0
aGkS4EYzVjL/6P4TTBMaYRt2gkUGbAYoJg5eIefgljqvWZmb6DOYD+/7VdjtENJr05IsQ05S7iMy
fCVBwnEcqzX0NIGFuY3/RX7xT6VqA+FJXzJDyf6R2bQujiOMDV9ThIlPqTX9Wy6cbDHI6ZJ7Gznj
9OvCj3dom3vK8RxXx8uCG6Xsx9cIaV7MxSzwhAGaVv/D1ReAW646eXt/Ik+WflzJ8LB/0RGqbXV3
XhPiXuble/wzPXb1k5WkUsNVMDgro59w2QYCqlCty1TJCwyTIaJKLvNm1G9wXGG5um9SFSskQYdA
s/hJ4LBR2zlcTntmhsYuN2VO/lXkgy7DR1tM3nFGD6b9cGnLGQyRCyYJlQU52j1s0baVAOL4HDQP
IQJppvVY+x8RTBmPG8d6jsS9mXW63mp6AJ6c9lOYF2upeD6tLALMtnzRu4CIaSK7X8zk/Y2ipwiI
B/kfLD0cfQ8jfqDakou0V/8wVUG86tyUVXwv4HyDnyYZjB63Bw7abwqA5OBxmedRGSsBy6CyBIRE
D1NBBUfk5fEP7ZITqgtfpnWRbEfM4XQ6vCEOznhdfJ8sZD9MtRBjqQSTUH4288GxQmPAL1FWoSS7
ie3fnbYrH54///gHpP1LNnpi+4+kTNcwM93UHSHr/GhI0iSq3AaKdhgDO3fA8/3ZpIA1BJulhu6Q
ZZ9JmnmkdhsMhbCETLLcXyLjy42tw7Ww84bJ/9n8wWJDlryA+5SVaA4tA+76KkLWpRNm2tCUd/VS
2ohiWzuGDwsVgQCaFdViFpX4IIFqT7iONNn8EdgTzM3v0tpaZLTr+gpGCWIZtMW37lTioe9WnliW
MHm3tm6txPef1BWZLH5nbRb3FPoQmVSb/tRRon1jagQx5wo+BSlKao6JYVwDuoM1eFtz36eCqsLf
xcrgO5Z5Rub3M6kXjElkgWFkNvj2QP4XZknnm49xu52X6Us+3pSCoxl3TwXAyyIXJa7Aow8iz8Ok
xEJOsYD5NYqnHu5sIRd22ltp1KyeyDPeUsHstLVYHgfKN747gRXQ2c0+3XuigR5NbC+T2+9S5oB/
NwQmPngN7BpIFA8Gi8dlGvQeh45aBCOHr7P7UP2oFznTnErUJ0t+Sk3/xY6d7reRMTDpKcICJXP2
4nyadPooI3Utu49gwLqlSAx28tp6zIoH04gfuXBcurfOmm9XMfpnRt5Oy7Br1I8/tZ5xR8Qe2yfA
aBn9IfjKpnfl62Xe88OwirAkIbVgGyskG7boHtRap0F1P1UrR+iOVymhP3TJ6XK8lFrOE/vdVpsD
xJaLZDUsrMa/UPKd3tfFgoi0Q9ceBYPUexveWPXknJK2zwGN81BlVqY84/wj9ib7WigN0IJtWwL4
xlra2JcBoC11/mCPPQVuC+vT6KLxUOzblH0cP/XBxmrweAY4OeB8fGqrhyA6As5Qk4iNH2ED1BK1
5WeQ2PWiuGiJBny2ROJVrpl3dhlWAI/fHv1L3jZlMtCg3mKw8XgYJoX4BnGnhb3WmTu9wmGMAUF8
4l2Z8DlTEigJ2W5Tqr/cT5dx0q1bE+RW2QT4/WowruUYzKTvBl4M39Sv00xPmCOgfthhhuhxjXdE
dSN3L1NMPOXIPI7JIElfrqfFQeRCYzLEiq4wove5p6zZjN4x/zdfG90vUdQ0D8igTx3z/5WcrTR0
5ybr1+If5zGXgcRt2y86AuxoU3xoT3mxvs1mGyzigprDDWR8lLtdc53rirTZfggwZK/M2K2oyMTj
uuyRrWbaiRs4biDtLPpYIBURc9XtljaBNR1kPudCx8HdYaOw8ti9j/4mDZLg0k5Pqq4CEhACpEkb
lEXzd7KttX3AiTqxUWzNAgef0ZfgNOuFkGJHgnoRAaxXYnu9ZutbvCEbMqFCtvcLDJZQRp6jnFwT
DQCr9tFtcBgyoTTEe+sUgfA7274MYS/yr0i+ilSx+wQrVGiz40ALryJafBYnJhSHns5qqJ65eEEy
HToAbUDQauq/CTd/ahFXOilZx59Bta2Y5QExB3FEKKfXa5dv6bVwQf48cZ7AB8LCmju1/wVWeVlI
p7bBYiD/jQ7P1TpbKFwywClFj3gbpuzl5FjOiWTE4XiIESLe3PnamUGqztcDGIyiJG/OY91hBgLB
a9dtwtyV/tIRHZgYauD3s7Mpiy61NI+uym/7G2hmrh5q9qeUOtoZpjk7UyRXKTzSRWMA4O5X346z
BZQOQR/N3p252qjju9xjlep32xErVjlDIKEYmtj0ATPUfLULSoablwIr/ub0LzwuPAJWf1tnHU1E
k438HuuV5OpnZRfkzFLC9U0OtAxY6gbcNGRy3V9XtHIP5rWO+agYrrc0aqxg5+UgcJFq2Otw9EdQ
WqLgjR2xqDEPao/93+HShejnJap/NpcBRq1I3nYitKfEJ9sNy7Ew1Qjzw9DMJxAfyLJf73n8WfeY
lk0iqz0TLjiBmdF+4CiSQuagXQ+a3ENL3HHRZkUozEQM1EAoYohjjsj28lLzgi7cMmJm/mrn+Dh5
Og8NEr0K7JNHfH02LwaVe9k3DAI5kDX2HaWpwYrIxsc99gO/kfR3U4qwXLvLXSNM4HHB1NvxHMmu
mKu0u2FG1JW/cBPXKFp7yV2nr95Ml1AgwcSbh83w2KZvSHmZBRouD6YCcNaXaKOPypHk7mo2jHto
z81RbDHhbZgR5O1antsPmNKi+flDGLp25hwTEeHWXsBp7GisEIoleJv9Bjsexj6N+q/dnTs9mgdc
0OJXkQPD/VqOfXk8Ad/yj7UpB1PozzkelI2ai5iNAdyZoy9y7hBUqboc/vTflErt1swuyyHzllgZ
95iojj5sK8iEHKEole6ble+CAa5UTnikDskQC9CmmFyf/RxNO42A55mKeRPFvYWwpp0GqFeBisPo
boW0Bjy/8jEy4XiXkHk3dzNWCbq5HQgLVKA8QVwM3OyL4QcLhbzRmgiB2ZfRzfJk1Seg1ILWjuqz
ayV+5O45TtfVIwQ6xqpgiRJgc8it55xyOi2fgxKdTAmrntQSDc70tgL/Bdwt+FHjDHebEdna2AHO
1sObvQiCdgADVKF9p9VIQMK3AvLSEGEGgoQlURxjDes0/1eIs7I8uVMlXmAHcdoAPHJ/NfsmAIDw
aWD4Hlw2eOiv6AYjrvurp6SxzsHaKMuHYhwXupEEEuAkz+ZSV7hBFZdBfqocNoxkVSyjDrAT0yts
rtZWB8FNivwZyP9sRD0O7IFUC9PuuxlSvGCXnQocev0V/sDevuYD3OiipfpcAcBOv2oBb1TAuAHF
3WHUc9MCM1s9AM2fGX3seULMV8iM4h1/N8fZyyaMiyVZRaaHS323cCVPMih5Kk+tY81dAg4CWN05
4j4xFcc5lJcLoedjA1VMnm75D4zXRZJneRVEB5llV4iJ66FK8xjilIK4sziIureM2ZwpfRjKDf+q
dufjiORxoiNQEVDsPpsay9rG6RH1SY7CEkC1yuU6tW/IaWCao8/bqh/SUk9gROMqjqecPP62RYnJ
+v2ZLqeaMvfrZ5JDhBohwsSJ9lmFwtRiLkgpJgdxQtVn42xojCjwLWfEinb+RNZe6Sw7YiPVh2AU
XMVAdNSuAwoWGwgq6PAjdCfNFH1WoK/+Cg2z8d1z5SWr4zH71tfGTqQ/mH0idaH8X4BhMFGHRreB
Dck6vSDP56aGGyHnKKJ71SWG5zB/7kFA3QDE2drGAiPwUcOQlxdPpm1thxKE/VPRznzY4Utj096X
zQjXSrhsFaJtXmaL8DK8BOJjFujGhf2YPOByNWlf9gUocmAhcK/Mt8s5Q652+hs1cOR7vxfRquqI
5wRoCrfD/JD6Gsj/9frJvtsUI3ZIyFcKTLVC1ey1r8va2nx+UaNn3cKMT7Mo/8kFq8gfSuHH6lSf
4GwjsBwzbQdop5KkeP+0YR/yA+JEhf30L0viRmdm/+lRx4qjVXK15AK2kfOrAoRrRxviEEioKp9w
S3po8syvd99Tf9ot0GeZbEXOjQNMohamoYLpNSCccfevI3070C0LdenQJQQq1u89fQc3JUbWoaDi
479bNkrivd64sxzc1n4n1aDE2/0ihM1SWvuEZ5HwpUriF1YM21wsY4xbbQNstV6otp//Vv9ln4Q8
wmEoj66W0BKrqZWobsQCJy3M4Dd4FfG09ipPr+4yN9wFQKhJYH64RNOtvMFlHzjx5JeEtIczcrnF
hyPPNFv6AtYjERoEFP+rJljZ7DNdMD1uSu/SdamAx0rCo7gtavopH6vkjo6uZCCahl0lqmuPsK7H
eeDpZmIdDDy8LMYKwcPcSkB6y4fA1p781AOWq/zQZhtuOCKlRezA6D8cfaYo0lFHbR6MjIPMeeAS
KrLbFTp1meLWwwmfc+2fQyvtQYnCCm3IgVtuiSU4P0Qq2XWMm1NG6yJaykvN5ESljPBJ26R1o3PZ
CDjnfEwUf6MpgGRNGThztfAa8Z4gOS8uPSpDGBDrcbbARlpEZF//gw0sm9OjlIqSRKEiKKRF1vd8
xP4jx+rQ52GLjonXtFoNdfbiDt1onoidWT1JXAWbe9H9eyO4CqdQsXDBISK620Wx+BuYKm2PPUmI
936mgdFeW14PyhHKKrO4hMdYh7g3AoJAgE467vQSVZfA+gT8loXT66ofvYmUTUPInYaXnNMSzyVw
iqh2hKePd7CYkgSAR66s1pzN+6MOt767YrRNE8p8PGyjf4XWsd9KVenBpEQVMSwPbe+gth2+Lzvs
NrDVxB8JX4wjZAVPeXl2Lj4GcXRUvfgRwYSnri2LdAgI4UhdFbovzU4dxzb4GhX52LPetDhD+a1j
gCY98+p7/gGr/5nxIDJdMETsczd2ZApp0L2JMp/TZ/jtbgkeIKn3NT2U2qAuOzYwftfpU6D/BOhv
beLaTvV+PQ2mf/XhuCsONa/13rUhDYyzl523NdmY5e18UnIRpGGo7OYzSGYsonjdh5Qkqyzz2ESg
2SEg2tYZxLHkIuG6ktVBsGSWzbkjKJfyasYGDNS9UwJujXN6ZTKpcNGO0fzbfxVtfsy5XtOAP9G5
FzRym8OC7I38PCqrihwrkeMVK9bMSJx4HPrgRVvsELmm62ZAmJgLDvBHU3jLm3BUGMDvgYjRdGOi
zey/hecrLHmkZWS7jxQFJ8OeAeoIY4ysJ89nR4EFZNwhDwYyOOeAvP3i/Mojjw4wkow6yonzc0Ed
5s+HQJSlfM2C21fHWhrzveZ8v+stHxOTjqn3hzVJl/fjQ34Ot66/AJ4gmzZo3GLAT0KiXGvgZIV5
yWvRFR86ywzesCw3NPg0PcRtyWoQ9ccxh/M+WD8MwWOYRhhKmpLopdAEDINoXQYl/AIwzKWroHIx
ryjfEdqx1FyfKw7LpdUrfdwvl1dspFKTc2iNO0jcA1L9z4K2OW9YvOlCGng1OdV0w4JE3QQRCLB2
2bbecuJrUYeldep2o4lc67XDwXjqkGSd/OYDXm8bOuVBr+AWz/0z6Ukf/NasfKLGfzuygjr3C6tw
EZpvYHTWzttl3EqVD9ePP0E0oHXT/99kCz/Et8I6vZLwLKznGyycjEnojK6TJkc9UTS/Jj3ib356
GPDjhGKkaaum/Z8ZhI+JNIU+CyBKta+rZn9/Mc8Rpo3iSeFKScQ7fWpwYpnSczdfl+L7gFBgbC82
S5IFOJ4des1nHFo6DNY053HrLRKbHWxZPHF4W3TAJ/v47brtPPUriJEjA34a7VDU/gIsaf+RCd5D
E1SUrVh85cn+9DpOO2IARVBYdSJdaCMNdtgUOUUJtuS+mCT3EM9VWnlQufjNclmEKLnn/dpGREtL
cgpRi3DKaNW0Lxg7VoMqFnnCipgCMrGv+c1ifWDbYosupTziFHc3JAHyIW0zjRpm206H09k5G+yt
CcR3LnwDR65LK0+rS8MwEKpX1CQCA0wcDt9dV0Gh2/s8y7grRup2XFjyoWI9Mj8ZwNuXD5DFBDAt
hfBeCRSXpHutX7FcLZhhDk+qK+pqNwoFezm8JpQpmngBr3hAVO/Fr4o4fOJ8szter2ihYuAENWvR
4V1q8kDsPHpOlEIKIUd3LDnrikOuKhA14REFKygbBVaPRup5fdgJ410izwf+dFMIWnHVSBu3nPmq
OJbORDmGf3sGn/Jt7epF/20q9kdxXCHI0IolAGIIplcZzghjSvX+SFZkCNqQi3TBpKBSOXZFw5KR
bTh6y7iw8c8br+CeFhjci8iiOfVPTPi+dGp9XARy7pIHl/3S3S3/rcDSkP5Gplig85y+IRVGtcQp
+34Rf6v0pVMtXHj7VC5H6p7M5FUFUmxVZC8HfhN5mDnA8fT5eSX94N2D8vH9MyytNhPOS4fxVzeK
nPuwJ0T4HCYvaEjb1j6F5Hn1/oi+61cbsRJ6rbTkaY7E8UXoEeWSnij77zztY1jOppOlQIknstxJ
qCVNe99/8LqKWGA+19+9/evEmwrCrFzx95UVBqGOhcP+4TV8wzOY79Wy+s4efntfkYt0L5AszOIw
3N4pi5zUwXf2Z6CLaXvq/kuG41+vkdEtFyR+sQzFu6jtoKZs1UpMacvbGpqsS3sBsqyL7Bsqgm8f
GLYakeherSnpstk5IhbtCxjzU1RdlBOw6OaTY9bJFjkKATuxltgvgeVl/d2fa3HhhqVl7ur6NcwA
OVNPIYSrQztNEEtnryHnXQDazdYup6q0Gxqibo8h0sX9q9c4JJ4wHOjFs8pFyrzrC5NCKIlMrtyl
LeYMtZMDPhsQ/HKaAitBboXQBhQNIYY3ZR/88ovtUg4W/HGP1wW1bveM9/fROKVZe17eZAZ+uLQp
QBtB3/Ckuc3HONqoKQYV8D1kpCEZJQkZLPmC2ZiPZiK8p8orUPTOK96+Bv+bJvhZZgU6mo5mfOpp
vpiBcoVKvyPtNRTLmJgdfhvHMD6VKudKuc+dzbhWP82uB9yQUm6EcZVzf+pprElOqCSifRVGQDwj
R9g7F/0G/lNFZhgWaG6TqysxBk8aXzB5VgsmhDHjPwx0slp4DDMqibD8z4etzCPt1GgthZppoG/S
pg+H0K8VfmB1CfXIUnV1d/XAmLvDSYSKZvgBN+TZhPtnSaAwxbXIAhnnOYt9Ag3E1p3i5h9HfjE0
5qgTRemmY/ZubA1SnFLMhN5P+jN5J8YCNVIXZfV100+lHcZipL+K2eve8rX7ChCiJkr1GFmZTGvZ
aiqErG8SUY7Odg2VPG/Rm0iIECpxM9I0OLt1/UeA9SV2K1xiPYLwUuTr2F4MX4/JTTaq/ET1EVNz
ksQ2Oa/ILl8pGTR0qI6KLgZ2r6GF3N3/jKCJdV7abUBP1pP8sDvx51Eogx7l3qilUZohYWNdSNC4
Mi4LzpesCjUFXNtARZk5SFSWAk1PXjQqzA0y6bLSUaxACvtVNTcjqrjmfamrJz3hN7VDtkH5bZXj
1EJi4d6tyf0QX3SKxQx5P2NheErRSnnQMVznxcvoOd/jLMl8nvgYHRGJwo5tBG+YDJQBZ3YhO9uL
nJowda/q16dHV3DboEHl77Kdy9ZGIfl0rOqdlxfgXQo2nTyrOw0HG/YzsQT2Lip9q0+VlprCUbkX
xbqdR3VWvXz6Ro+URSi+2c5743LjaufOVkzobwIWAnoBZZmwTm0IIf0YbFPGhYj5oCyJFIOX2VbS
dvhKC1kPukv0Q/Anidy+0fMRvCjdboqO9UauLzQLTAUqlhVYuYt8/rDEvhSxRsbkjCyDur6TF/j8
MddKU/UOo28g4Qft2FuPlpa2c7OS/87/YJsEYQh0WYPmaeWrDby+ocEv2AG8k2HNHHx10VBsqPxU
iJjdeacEv08JXHaFlWaww/ANFuvvw9IGjgDDa9jqYHU7UZleFwup2jLt1hHH8QI2UhsFmzuzOqot
ApoVCj7YArmBKC/cEJiCFlVlUpq0qnzQHinTtjKqXyZ5YA8c2CUmoGDvhjeoIkOhXDfNj2HfnDkx
n5ZnaxhvoCrWv1uiA8rb/ADsJJkbeXcM8O4fv9ZRbT/nHIPZ/lhfiG90PMqbrTXArlJyfUJRq5nS
zm1aD0s/2A6WAX34wgM3yh91CY2Sa3q8rDjUxVLrddJHGmN3/1EF8TrJV3Pn66UWOYHVXn7Bzv2g
8nIDPRHZkF5fmmteNDihCnx5GnchsYFx09GZKQr+zsQ/Eta9/dKxsXl8W0WOZ2IBZcxGPbsYw/jv
IFJrC4b3a8n8hvhq5WzHLm0xaNuJj8I1Nul6azewcOE2sC2PGhZQrdIn4Ac4/oefe9ieO4bmTMH5
EO2JTvlO3+HlnO4sEMpHuGvWA7n1+87W9miSvW7jpHDimVmUFt3wod2JKKnJFd4uGpHTAhZGOnMR
foSQEwidJ92ALqoGCdYC7dBc9PN5y+9acB2bbHKrF6NJxEw5T5AXBzEjQYGfnENGR5wxBCQ++NM1
kVqR0KADJyDuRXFCbk3zTJmfS2H4ZPrr276kQxIFWL27nySR1SlaHIF3K6B5xoUNtFjkh1NMTE8J
dSnoQd3SDXDue6+mY6Ppw1Neqh06xjRBCK3d0IFjK9Z2X4VlSnkMAt6x+78v0rFQrcGFcS7g1IyO
j+o8jiaRTXzP6U8Y7rnYQi8W0e4KBt48ZXp7NmwavJO0QYxwmGgOeDP7Fd5SBz312QyvcU79BEJB
h01r4YdvnMuMAxcP00cvKwICPUpypF6ZNRuCnSIicYqrt0rgG0P/42ia2UV5ZEwAvvqER32Nx8YK
Mj6LT1c6bqfdw+cDoaqmhcYPFi7pmBjByQnNGglYAMd75244FLjc2I6SOv+VDrteIfoQr8MTC/Yg
hMEk3M3THZe1Gu2BugjmAPE2OmyLCMTxSegOzIRjH1mjmtAWHeTDTiP7low+/xJ68FddjQjLaJSe
Lf9WXLJ5DP5n33inIfY3zodN1IlZq/pIdMh9Xwjdb62cuoh5nmjcJG6x/bsDy4WxsLGhwyUudWIb
LHuYSwqB8mYUYZzIAubSKVzNObgLcaP2vzlit1jQoYMaZQasAd3uN1iSYIrp0Tk6wH8qUB/W8wdJ
gFE5hok7e3RRdeIu2vh1/JKHHostG1x5OEw6WlaTqn7ezmnL0fReUh87qXMvPMv37Fy2WjeVSjlI
AEi+pDFWv6X5wD6udFijw/VFe4eH2w21pbCTOPHvLuZ7miSkjsrHVp+JYIPWZjbi2evrOeNJ7eIH
bwIBBR8XuJ1DThWGVfRMkCThzXdYyPaoqfqYmRCaqxCzrin2mqGoyX39AiJ9bDJsRTvNbRHkAc7p
wnyWdC6HnwKAAp5LNPGmnmoBif3kVIbGbH/IX5ge0AF2fY63yfZ+EH/g+INUr0S7cwnao2+VXmav
TtyDyuC/WH6dD1SKS1i4Tbb6Ht8TzkLXAPUPbmy8WV/9PIWJ/dmMs7yrKaqAp4d05kPSBPYa8bnQ
D+4U677vViD7QYrzMqiQh4KMDN7h3H8QuaRG2kuwrvcq/4+n4xXbohKRlu1MDDS7gZ+I9iwr+/h/
P9cVmaSNdL6Bpwg0slowX2FJ4hstrUtJC/Dwo0PPhoXhubNy0R+zSk4GoOHOqd/0s9b3bZOWfzKl
4m+4EOJbeD1i2A4K1X4LHxO1nY4Q2GY8zTfFDy7O5e89tNEF7o3BTHY1MOrOKKyEkWxDDGUXgGJz
/1qXrtoMJTpfbOxgL4hvpo2m1xglMW5g49NseKVcxR0G8jMR0HiBD61kp0Fa1ra0KnBovav1+UAo
St94iCN6ylfvh+Goxd4A8P0d7zUrjnOkWuDKnJhhVH67Lq90aBOrYHO+DLbNi8k4UeUyqr6c2Lgk
MCnttgUD6n3nRzSAZVDWSHiDie9IZwLqasZ27+NdLrus34zb8dgpER5oafPvA7JQztYuvl4+kPJv
RD2yP4RG2d022ehS4moUYiDoLD79qFGmr9XhXjMmRA7wT6e95CUCMXu6usvswcHN3DPg2CpQXPix
JTDed/6Ge4OVVHlTYAW9JnwQnstX603mesY9T34U77BB+YLZhc+gy5HYYVIQ3de9Y6RlR95Xb9WK
SMdbrdmW7QjG4EHz7W/dLfRdVh1aP5HW5NpV+8BE7IkKGIzFKGywAr/6EkacvWR+NUfiNxyz+Dyl
C91G2iMDZGd/DndPvId5R7D+dH7Zuj43zyzrPBdntLtcaLtKtUB8qq1tZyktgRPxC+4catdUpraD
KWSXguc/2C6Pc82lFfMSBBm4ewy9p3sqB6trVGS/m3s3tMQXDtoTYuO2/2mfexd08JYexyEfwUFn
hIMDLAqP29oNurXChsIWDgkma0ukVQlw/JvtFTNzDO8NWAoAhUXVxRkIXupearFAmCxAyboZ2gQM
fLwkf1G4EWl3aO+Stdd27z+nN+RBU41quxhPPsOOXNZcv02ABGuLOKDepa4ihiEZI0ZhAPhWvDM2
E2hoEFU2wzZmNVJqxK9v7TVA1Fm2NoBkJiDwilQZVxBtFXyhCOe3hzF8KmAsGDyEMIBePdsqefNY
17rWFx3kt+2WUv6iL6w5+11Y2Dh+rMvmc+PAK0chlV+22YUqAfCpgjg1jvlYNZ2//wfK6OI/ctcR
th2wjnwNr8MTkaVrv4/V6jKJsxTlaEuQsgVAR0L+3FnRrfck5j3ryyD6sfgERY6LYqQ5G7Ed8bqY
bB3j2HjVmeRafzpV8h7EWsUefaUGBM9uI4hyADA+1IvZSqvkHoHz1GdRtWJE/JYqSHX19jK4XX1U
Xjg/nmh6WzRolXogH186Rz5zp64UAhx4hjmHwT/PWsgp9dG92Rmk0BXSvFDAcmkXTUu0Q4iKozmK
MHpIAwBup3i+2pTyYDc1cy3R6pN5vanVMyX0jAMpDsrLRmBg8ORSooL7OjQ4+t6ltGQLkw5VdS4u
k12VnAunHBNRCkne9Xr+7Fms+NesyRM3zdjtB4ZgcHhuJQFgs8pJ6UB989eya/0WHrI2JpYKMVGn
iBsS3c5agQILseukhPKOlaWPpMruhp+1Qta8pYgsPy0Cuy3LsxrV4G4JkiOpHwmgNS/Ee5cyKBDK
/ATj1M1+WOU/X/jm6Au4Z/7COWbY8Kc/PQ8TTLycK+zvUKt1F4z8fld0tpY0H1c9ldYsAO70owZ3
fLHqKrumz/S5ungNdpVyYW6RhUX28O71CJ/xTKKfSLzaHUR6GLugqAsuuD4gilZWWDMN/pbHjO4C
vqLNkEVNwoKYUFks1nG9U7sHfP5l2z3W30DHgEI5a2H4kGm3tDTa7XFzX2p2ara2oP41G5d/mngh
iTEZJ2PwNEMec/IXC26pIKDE6AwQSbASejMKZNTqbH+s1wdu6SRwc5Og4C1l2LqviQpFI9k6ZF6w
vyoHaNrgV7C7AYrUxqZ/zRRysok+nT68MbsTmcr9kr0fX/cJjayrAa83i57pDMHF8Mq7a/vy+g2r
JxNEWuYynt1Oc+gIaT17efBXHfHnN7pLHjFP921bVH/iKwLhVZFBXuwZNK4/HTfbZC6v/MigbOjg
Livi5qIpvZ5Yn6MnV2fxgVNYlegyF/aKFjnqVtTOAB4enCJ0PxTf/RMDSJ0AlKNPgJvAioyYhb3O
2dYZj7qsw2iDSl5m9lddRAHjQTo1YPxhPlQhBAB39YaEplFlNy/6QRdfmGcIGTSm+QK7uDE7P8nt
qh9fXRbT/pEIdMNJfiebtxUN68FN1OdJPRRPfMfrpYXs2pgJOC8sMcnhbbUIqBO+74eLQ4OH0rqJ
4UqlMbHXx5jdjLMso6H6c7n4Vuf4/0tP2oRBogHCPj0R4+SVis3/wVSDtjF0zlFbdRLOa6dw60XM
TGgiaeOqOmiWwDkDirmXCtMeUj2GNBMOGA7yTsx5msaYbaQVPwN/yZtG/z2e0ARFM8A2Xg2gQL4w
B9IYXSslR3s4gctnwAAcH2y+P3zRrLKzrpwm4TsggbDgFJWcPEJlpmM1Ry91gkBd5v0JCO7ipEI3
Egr740R5/ih1Q0n9mfqh35vuhRjiOBYyIh9GFfxkmOMsOF2uSOiLUAnvH1e2akgeg6+n3QcWUfqd
I9rXCCN+bnX45M3wvUTvz3aR5vhfjP9nBEJBJZJ6iI0K2qKxc+4u5/jyASZF9TnJNcy0JvOl8VYm
mt/t5B6XmKycdswYLLJq8O/SJ74uZI2hfOZKOSYHqaoq6vCGERmYvVejYho4cimMfaRpn+FDFFEy
F/fX+NBn+EIZd/r1KpIz4uEJdH/rJ1zOPLpSzm/AMW5rKdbcE1QU7llQi+yGKbgQ0eq3z+Y4pEfT
UpjXt/FDXS5fzUVmI+MhFz0dHa6Y5b7K6d9NuSzP5fFwdeyhOG9Z/NOeAdkR0Mvu5cRrF5SnB5j1
4uVhcCYtp4PchJt3VVFiRhb74PLMxIgH2g5SfoWdj+O1012yXIQ7HU18wLpXMVTv/I80ByK3z4SE
BdQ0Zgeh96UHROdxY5gXcuIH0dp6rUHtDw8MqP4J42ZcJyD0vjimNJt+GH2DVwkibQ5bo3oCHqqL
QLlCKaIRKY8twE1rHanLlVb74FH6EK3A04qXmyIc6HUqCKCcSmWCQ2r+6FiEBGctr6OY8OgBrPYh
j8AZ6iqYqefhwHl8SAWbzZlDO43ITloOmlzpkthTqxthrqaP+GJdl9NIIESML8ZMjFTqti1Klbwi
uLgXU2bDkQN9roXiMgjbFx6RxKEvB0X0LE8rGfPjLCaUDcnwRin6Uu5HTpbmCmPSbqb0N+0aBvqg
raa1DJR9wDkVJKIfTS8ScR9Lm9v2yFxqyoAj8zMnRatyR2PkujnieVxEA1y+GzZ3ThpSLurDq1AU
JLUZh74QmywH/fcG4+5fZ/hjU+r96XUMVR/wGDPX363F2cP4bkABOw69xKndF0NYTmQSNIbkUudV
oUwANoQ1SHqAYGB1fD4h6W3Lz7lwdNmladLj4xtT+HYgk5ygVQqDNTUx/u5O18tqQIxMpkjYNbyQ
u+uutMNcXaStM+cnBOpHccGzcL51blibW6TvsaNz5heesk3JPS5lT880q3nnthtUa7A2veDMElhF
fUid2iFYeFspHkm1HjATebPCsga47IDly2Y7+OHHaqJ90w9x6lrlBkMzraxEiimSSeJNj+XRBeAm
qysKmmoM1ccMo775nUYqcJC83sIFMSuf04MTjEaGgvSyEL2m+Oq7j6b+iA1vfLZ/1Cg2FV7gPEqB
0OfdzNfeM+UsDJrG9VuLZdZio8ZM+84blJFLphx/clk/PupZClKuiV8BB0A1vO4zIilEPrlOvs+7
BuRuCOSLbEdUgf4JDR3+H+suz313NQ4EoZN2T/DHQmlseZ1HKchha8ay+jfXFGN7CQTynrSMnqT2
EgeiBerj15D+3csm5ScKLx6uIgp+u/7FSf4sll/Xk26EIs3FJFNVCceIynr+LCpnmAnnxfY1CidI
Nd5b6yLqXDPuZ4zq+YzhWBrromqI+ZpbYjbEPivXEM2ZMoG6ZAM5dDypRo45YulYucBXick6yfCO
xCi5qNdN5X19W+FVUKQUTovB0lYWTbbEhkeyRsDd2OL2Qly9/ZRBsKH9XFXVrBZ10yO5Qrx7yizV
bFmrIuVie1kY8HF+rZPGDsaaUIDOg9LrG0LyYsYx21v9vF7yfXxm1R6SHJlC646t+a5uEyHlVgal
KDxgiZa1X24tM19KO2xkj74SokT8HSTRG+hItVOh4OrwYam3aRK/fsrFL1X2z4SmN+uef+kBqJP/
1w6qayXNnkrX1ijRZRvSGoR73H5w1jshIhzOwMbAG6Bv2fT20c/dWgBMYROrDX+UyOhlIqDU4BMw
c75nOQcSqD5X1pn/4VpeihH1gvoL1X4RoElmJ1WSw1mrwj6oQDr0smmkyTPayQkWVDzIT7tu3lYs
6HlpHH+qKoI0u5Aw2fMFz+4Uq2WR01Yi2nk7u61ttn7MmXzYxAOTlnp+3c1U3+ARbB09BaAOu8AO
XHD4Q9arKMnckwB6vubddjr96EkRZ3aWBqJBDBIgT4cYIuOiHGaIx9Ij//k7chfpAAuBOcBzVhAK
g2h3BubEtOpBwbCmOrlxHc8lRPuzUze6Rjhtnb81OjMpdVz+DClEG38OnIxSoqFH3x2fJkBIQq8T
pySxzciqee1bkRV3TW/pAZnQGlsmeKyhYNNqEzQcM1hAKHokwgB6MxYjR+8cyk9ZgWS9pOmI4dWp
sBTD5colwh9BqRINF8xTHUaomLQ2pBCZ4X53k4acVjzDETbJ+qgtdt+2+V956kmC17gNarpC4PJq
Cjpd53AU8vj9A9nXYxxf2llLev4oPigjX/K8bp+NgqccQ87FYshSIOJeooIOh3itfhnkhjrWJgQy
4UdJh/jh8gMMKdGNBya+YGVSSZaYpn4ZtMx6dyeJzJ33XMMHyF6a7hXDQQwhB35Gwb8WCPmsrf/C
bdUgFstbafIfUfWTQ1gfNjSgRqX3kgEmTITBLcBJ+fnxOTkk2QmOwLRqQE3dL77YsDmADv9uN8Vb
9IjE/PY2fZZbMYPDqxR0+Jp/yGYDBFurTdc5RO5tOz9KNwH1rf8+8CptP8Nolt3T2TOvX09lKY0Z
kZEQxyxFlMYmdpHdfUswnbtDghKBZ7WVVUsYT/hfw+b8z7xsqJHDeDlQAM1yjQxoUQ9lXZ7E6uO2
qGzhtPAZ9pG5Ixct4Lo9ad5b/ila02W61yB9e3q+m3FG1v+X+Ks1zqj9AqhYdPyg7FBDLP6aMxft
3qe/ZkR/WUKm+sXIUxBLoZrY2kJ83pW4oAyr528SD8c8SdBfmxWVzCONwUm/9d/lEQf5lxE9wzUx
YkTHdkSaN/Qb0pYygG0LIF2znrVJk4ogJnv5dLMNGlYMctUgKW4bcbNhbcWqW9t+GPBcL9jRMXh7
KusZ1ODHZ/Hftp7GqeAaqoebONo165MEfFqEkL3y9plhiG3GYSWgZmBsbMRYDYjBKvl70SbBc4fO
yt7fj8iJRtsREOxaPV2Qodqh+6EZLy5p+q8Ko8L94Bt4kqe0AsZuVQaW6SJdCH6Sxmi7DSn3kRbP
9wL86duVclxY2R8AEJNBugktgm3cxllxoIC4Y2wAwWsQmMoeCYJ6HxjC1TkAKRAdLyME8Cpti/Eb
BwvLLUFowsAgti0m4WTaVjlJMi7rJ8nd89s6o9R8FdXR2+SS+yenSfqTpBHpVaj4LKMX4Bph8IVc
dAhADjtK9YnV3y4J0yPjB6eG8DZz4k4FEhyWEL6jnxdrLc/pEhoQQJCsmNxY/BEJyZJ5Ei7Iz7TA
eVZxKGCbNF9Bi8tbiYYCs7A3Rktco/zMUD8+zB0wg0PUjgH4UIL5RkL/dUnH7kYanTQrMUudFyvM
2fbB24ihIusIJKDD/iooUyZycMUdJ+ameYjb3b4Knr+LcI7pQG3/THACE9h4ytwZaNSlen8Je77W
wpginNG8LTBWx4NFhKv3DqQUVYT0/98YP1N0IxzfjBcB74be3/A1Dt7SKBveWPDWHYKszhJiF7ei
x9glJXN0KGLL4Tfkviz0RL1gfIiOrJYz0cr5H5tWcWRLvXtEBrNHI7eGMVWgeau7v9SGiHOPEoEa
eCjHSzwvyU14HuxrceQlGysoZRnVYghkwgsGHLOWyV1dv0btKcKMB41RVAAFoypvHvMufWddmedV
DtEBpIwiEQ1oeLCGOezhbzDIePPMVhQCERXUufEPBEHN02jO2dhocWaqvLIqdBKMsZ2P6f47ybIX
SAFC6z5KMFWY9c0LpGoUg2wgygXbaGTo528oVk7s7sH51ErWkD/WkS8dPi1uUkKS9nDlHky6wOCG
rJ8L15idloKdy+mM40uciol/34xBFqX3PL6xRi1V1sDqZHzQ1kR06dQnggQN4CzpMC8a4nsenP/X
J469x1aMWm4rHVEoVE90TVNaVO7Dudik/STe0iUIUxvIdysxqt40mvJ8Qb8CzKtrI4E/o9v7O0Ee
wZ3nNyf0c3psiSHDD4uCmNQXL+lIG07rwl7l80B3RGVojRv4p98DhDm52d/Lh6xIwqHTEEZZpfiL
NmP+tBbyJRtoc+Q+Q3B6iEV1ZDu1DRmeY00PafZm8bXc2j/YqE1boUzlvAxdJgHTvtXMJjGlM9I7
GdX2QvwgT0rWUUZBobnpzRxELKJn/NqTGSMRoUCJgNxWNjSx7FVkXhrSq504cm/I7LS21nrZPwS+
eCC3QPsrljzzQ0slUoi04kxdGQ7k3zFqawssQTVeQ+LO4wbA385cDOVKiYmqX6nx+aHEdSvMdwH3
L3Np6Hto1uOTedZ4nDYHaySQj2WQj9kvDrEsE+JcyCD7lXuCvpztRjIO7nSKw96sPXS3StCIAgZf
PJbiT3SrIMC3y+ZtMpOeVCf1ynn5NUvYvK+c7FNlfHBHKuvnsnGOa44KTjlgtwg8Ybu+Rxz/8LfH
iPDpilaY7QU54PTtXBdmvbgwL5QX4bymoBpcjA7M2MW10XmPdNuktM5iQod1QEH0aJI640kxmRBY
4t2yc86tjN/6OND8KjJ87syMs2A1g5YDZOu9YNoba+krqYw93EsmEMZsGytvoaHLi4bE5EuTCXVk
n3HdvFUYtnTKB3gxePyS7+9ki1bIao0APEVvTRP2eEdbush4KDU7ep/dVn23g4N5oZQS1ONpRGUG
VCJevtGQeUmRB7uwD9/FUCCVN528VO8fXY16TCq7CHpKEGy25AkVA4atwr8uHGXajwRP2RzxFH/X
xPuMqE0c+kW/CozsWo6bRldzPpLUjDM4rwW2HYEGqxkGofP9Djafdmbn6F8RNHxeOJzCWggt2me1
E0cYuc08KgXVw2wKO3uqK65vm98mP72jZ6XDY/Ef7+wgs8apAK6/vJoKBP5BwkSEggB69emujPHB
C6iDJ74qeIhVMiP9Gvj9AP2DGC3kWIgBrc9BzsFqyhOoIqudsSAui7QypY5ci7uTXGyUzMQ1Z6MR
yp5xik1hOuFzGEh54mDft28YRuphlAnWhOKeaMbzLFz0/6c+WwXAStgGEOrpcdBtKcn2rupew5hS
hibCAH2GEZ8qePSgnbE1Zmf1fOt3ox5N9fRYFntgAPYvo1O/whI2NN1uyq4qdABPQBQ4qoAMlKJP
p8DbHf5Jm9yFP6L3UekoXv3CqON0LGyNKDsYo4HN716kALKGIgab8u90gOisL74UEjrU3xNkaX6Z
SdfitQ6IK5Jqb8UzNfUzHp/ltosHnj9w6WOlEJBgAsD8qVl/TH6rMp/S61T8HMjFy6O7LWXh4EZY
yn8GBz7CGv4sUPxw/GcFkYp8Opv2xWuALXkzU8WyME6cbtThZTDGAi1S/SDgFtFF5L9AiXn1eNPj
PaiOiiWJSXvcwFle3LEnHD/dLEs50G5FYg2g60SzbKW1z64Vcf3q4J9G7eJhPASSo2FRB645v45s
/Y5eXi/8aeaH65iJzZ4XIWy/7iHRFTXU8gnuaFsaoEGcUl09THta3C2cw4ptPWb+M1M7CzFymWx7
uMqv+1DwS/pdrRd62+V6eFtwodk5cko+ZBltM61iDYAzvse4Nhi5A7wxmPDWLSstV31fOrs01DLZ
ioyeFtxGxRGtgn/xzBTrkukQ4bFKrHAbkgM4T1Wuw/WMPkskrpXaSCnNr/teovb02Xczu9QS68qE
+DNnW3DcEUOnJt+JbcTpcCpdDjxXJo/gScO/D6ZdkO70TP+kv7a9UpAcynXkccvDjiTINSugs9LQ
ItRDhpqV4VdvW51/vxXjYK8vflbhx+KKsF2yisfjLx0jFWmXKhooCUM/14hirVgTR19Xpnc/ZxRZ
wX7baai5hUB0XadQa0/fx480Xaw0Vi6nc6459Ip1u48LxIkE/KPBb7/ZD63NTz0aVmddmsFZ4UOn
zTB7gCjVtPSc68wRN4Ep/Slo3B/OwRIuPGw3MIMgO7B24OsHnVlDLsc0yPk+0/+EQYMrmm+abUZI
QOs8dgEDmfCGxK1/WdRA2scyLms2xVC0nbBUNjsvoqrZLyyMs9cVpY5II0USp4o0J872X9oo+PSC
AsKVUsPf5+HIpaz4H+sXLDwX4Phw6cEvBOfCQ2FouGrcgSBT85xMBYwmt6l4dVDyRZoGmuOE1QV3
2xGluXKlRWoXTaA+yhsYg2duxj+BfioRXtu6ON2LfDQv+sY3GLELbCamR9+H+tSq7csNVFDBSn+P
t7ODbWiwkA/uSrKOPcFtOwaalIjthmwZzP2dBNq9i/0dJKkkucnpd+LIUZLzSdvxcyIrOnUX2nHn
zkfc1ozduIeWXFpXOQh6cfugLfUYlm/GXBJ4H51DbdiuNIS1EQiA9O9mmzuoHyjXuTti/QxywUDi
68N1z8tlSisBdkt/mGWt3AVR0tcM3320GPW6vmwljzn+1XGH1SoRoUwOWbfo+M8BaB+H+iPtlAcp
mM87x387vpYFi8a6eN7EffE0sqnv+PDSIzHOr604ErZWigBDe2quMSFwEVN5SYTjxrXCPhu5wQMj
ED8hjh4kzkKA2KnM7cHpTLR8wkSbJCN3ObquZ082/eYX4GrZ8PxmJaqbztjbQbqXK7eTFpIqhUZ7
tH3cvFz8Br0JU43dKPj9jRgUqbSD8Si60X5AFcv2Qhmj/c7Os1O8/JAfOaVy19FEzxEh4Ms7bgBz
pKoFp0MCTSvlHrQp2LjnFdw8pTSP5BIG7fXaMPOS5T6ZeY4M2gNneqihfs3V3/Yxsi9cryqdxF0b
jKOCcc4bf416Kz+RGlVObRdqu2QJZI20EhJddxSY6C0Q5umcaATp/E/N6LyoOKW/33x+W7F0nh6+
bxolaLtqFvDI0qHV9aMbYfTqD4aOAbUHHpecdqn78V24XzCFkFo4YaVncpT1YRnxmPeJ+mcEvhSy
rPQFKgfVjynNDNg8WoQ2fKep5wBUcleIQyNKIbXM1WchPQBycLwf0QjKw9Rp8VpLOr2MjLeKHK+8
rDDPtlF88uatdB1p6axC3k/x77ADYeQIZL4vMGWALLGD/dIV16KG344g0h4sOnJ3aYChB7MCDyJ4
1ILkD18tptli6/N6uI41twuYHGbVQvjOqTTDPHRqrHp6Id8pvFNMuu2WQkWaFD2x9+eqIRUuIfps
NDhnZbqIHMWSKfZichHHW4eguFWR43TwD4K6HZu7vO8PiFJ48ir9QFYLamwumcbBNhG8YXtKcN5N
znRtUIOMONEwWbmawBiutxMF/nTz5g3/ZV9XZqmT+fn4ZcRTM3kUWg9Z1i7tkoquqVw3y4QDbT2u
xexW/wKj+a6BT/WKGxAIIZbo4qfBqv5GpHRJ6p0c5pDigaUgpgE3kcGsvu9/eeiinxJhWcdbeJ2s
CjK9ZeWfVT1go8lr8d17GSJewzyv6z24mqhyBThZSBb7ML0NjgAeU3PGQQUSPQnw7pzzoXyPdpbA
MkJHOwfysCzlMSCQRunJV92SQsOAB2OaMBRlTP1G3xsLGvQK64Ho5HguLdayI6n0C5WVdudFVYg7
tO9g/syTij/r/hTWSReqM0+/YDHLcdSZP+1kK5GwcQkqb2SbbAdlm8+aOe+2L4rLdHQZVTm/zTx/
VhDWxZS5IN+zkvnoz6Zx63kzrOS14bSy0AiBZqzQrs00OjeflTXLeJACncciX1myIHrBEkXbgPV6
6CGnk+ayEae90t0AaAoywLZ8BNgxEjDdixuCXgdB2fEOC+iQPFAX4aFuV36K7DhOU8WMgQZmmSp7
Sxcxtf5jC2Xp96CW9gkwfNi76dCTPrPbVs60VsC1XJL5GVlp8qiO6jNSOxFkJK5S8QcOiiTVBLNd
liyAKsXlDZGOU2ngX3rTG8RuuPSfLN6ZGaYqMLlpkHhE27ck3O1IYpWej2DqJzg0ZJ6SjbxiMKy+
+5Zg954uYtTt4+ruFRfhQhmU6RT9DawGbsjqYwn/tAfW+paOPSZIwtSoGqp+mC7HAp6F4Kgp80fU
5UulT41ZUvlobBoogJjM6YjSTR4YrySQeWOc6KOoHS0v9NXFtkPqvAItKoqNnMmKWveD0nt/lV+y
GF7MbAtWPTF6t6V+eAgvohKnzmH4J4VUVCzEFZgI+djsWqGxh9Zs0p3WmxvLyCXgnO9L0h3ys/5X
TcYSK7Vkl6mGMklFUwPuuz55tI5ALoOb88REU1Ei+ErRr/9dlboIZlnsiYMrvyl1FWwkfEjUa/dU
lyVVrqtvkz4U5BhWc4XVcTaTRRYtlpGJDzdzfd2wxnuGPpzH6KNZcEznRXmOKyht/scCah7W5wHb
tGLH8VNZQ1AwdAp2A/tKZyZIf2AetdvnKeK+fSpDPnml2z6kNDpkPsjyflm4aqyvFXLZDmwbCWoE
a64gMPwSDQx1PGjKafWDKDQ/Co4VfdG1hu0BGdGhJCJVZ62DzqqAh6OA6Cdsvnk1eLFpEDJ7oVBC
ExvY4r6orT1kh4drSU+zuMFhf1/R8ewllNlzuaORdswLmVxsxKOTyxme67lk84c8cFSp+8M1MYJJ
MA+pWhhj0jeOJeuyvFDj4B3Ovj6wXeeVKaxnSt4QSIS6ZjErteTRrcPMJoCuq/m41rSvcfyyHcux
SpTraacPeHRs4q8qePamK95kLHtBeNR6CPcYIA+ERMaJkAWACpzLbWH6FljFOieML4OYCy3IayRM
qnbHT7vsx6kt5hj3HAlPERb/T3j8GlDuFEIf8fhtTCj8vsVU1FR+ixB5LRE9RY8FoQoXpEZ5Vah1
DLF5DoS9+ySGNWua3ex8SgAVUHUYviasXHwDSgTMBRywN8NSqlLs3Ei+OzrJrjauDtrNZyOXt4wB
hLjzf2igw1NDCLzWEIjO9N0FFqcosdWYLm3kyGGX572HEa6o6ZmDom8N+wCpWHBXXUHf0URkmmZ2
vwjQ1lV4RnkpevsPutC/ffagqn7aUmuWKvZ73uxPo9uDBWc2oDArSI7m9VGCo/p0C5cegcMKQ3fJ
nGl+bfeY33c5//qXi2fZPZ/3esRw6XqQmFAWlQRtbNFV1ZLp5MpUFXCAh//OCnIh7tkSO4jmynAt
xMFLQdhN3/85Ir3kBM6FMoLpL88AWZHATAcLJahp2A9xTaJYK3pp3XsEHUFz9NFXBOZoNk/smmjI
s4Rz1hwVZiXKuwNMP5C/5kOMMvCAEwzpV9k0hFh8iIBNLntOzMPXyL5pN5hf+utvJGNpLq2KJPy7
k5v2XHu9fPqEpj/xamCnHiOmFhtN/WAmf1aVcYK/AyY0dpd+PMLTqpKd+ife/dEpnPAZSmO1dhFm
AH4CGb+/c+0qROR3voSnWCNwx+uRCIg05WLRtDLBzJoH5neUucts5q4ojv770qu2ch4V4uJRwzzC
wOuGf4aiOHeFu6V0bWXroLnXUTpmR1df/vkGPzzRMyUdoAqgD80YTjL5IjCj9bXcg7vCjiz0le6+
V0K2KoB7MGqq9gYxqcTwFmGU9NKDiWG8q+U1FlDzYaJ6WuZAJzGrS2bLk0eLCYC2nyYaoSr8mpbY
DDK1yJnFctmX09GIpfCXbYa62d/DlPUBp7GVFBIJT8iq/A0ZSbbDJT0kuL2Lw1OP1s21dK4c3W9Q
LZx06KOqdKwvRrEGxBF3U1CKZ+hic92nyCM5rpBKFtK1ZzUJ5J/MB2RlACAa/QsixlkVpk3iSJsy
5esW2B8WRBCRMqFR8LLedATI+IiSlECPfXDS3SQ7mcccgw+jH/DHptb+HBK7E/N8tSL/z1ABJ5ez
yrIW+VNhPymDhyhquorkevJRiRSX7OHSv7WBJQU4VTdEGnKt6tT+ajjbpTBmfiZs99qfnGldJRSQ
Ylchq5oNN5KDPdnf6XI5G15zjW1oXMD33cFhzW9bTbG3k6SGAIahJmMyMBUvU4ot1DRd7VZyq7bq
HNgWCkyp+/c82hexYJtyM5T3fEAaw08YyQoQqbZtBsww80TRXJun4RGq8Tymbvk+Nn2jLeLqVuWn
OzraHvNtcnmGhmg+JhTkMZWg10CqQRiHwRXqho0cFFI9rYQIapTIl/dIJE9MivCCiz2mruQhx8zK
LyP916uZlN0hnwbioI+b3+fGZTKbqN7Ihwx0EcOZpaNCKGcJY+mSPL4rtSfUVza4R1X03ZntyETW
F/EaGPVUu+K5eqbYyCjofi/QoYwN8lQ7ObwlLTEMtnXviOggL4z+VAgAoHWtqYJYwmeCQMPYvOVS
MZxfoRulPdpXIrThTTEb514/xVLYhAeAkHoMEyfWiUiOTPqEI8WJb7KzW16YjFoyh+AAG3SUggNQ
WCBHfE7OtOI7UC+/rmsxbXOsK4O09SbXeewEXcxaXzp+9JedunDBkXNNWdTtTWuJxL/+H3BC8H6h
4bKxJjR2LAW+L9ec34/peqPRTxneDf4pWHrOaEQElKjDDE6uO8LOqglg6Hd0l7X38SSB6RZns5sU
fN3+UdDAmX+TrsjX0I80eiRtIqhNBH6s1Mt0bEYVcnpaxv5ZZzNBjBcbiXso5LvpOhPkibcwzg2R
s+zWCT8BjhbYLDypiTGaKMTNYZGEwpKHhkJBG79qXOkUx0IQ/iOfiDXk/C55IBikWBftPc0Y23Od
5pfk2Nphe9pvSw17Z/IPwpEnugHU0jRKrhh45XqQJcHTcwJ8ghpcEmUs9SidcaiMKhVd1jVue+UE
AwPtBOWVVGDxN2dLpOHO/kQPJL0UFb2AwPOYc8JkUcrhMTfmhifVUGi3t6bdX8qlmsx5mNdHZJcU
mSYRkQDlxQTP3A+DqdGC8Cy+m6R5a+GUtHiVpQHyGor9W3Ts+gpUMp4S692QOtxFtzFR8Qp87qpa
GzXOy+JA+Sw5f+9ivCl4SOwr6PPXsqyatjp+ZpaP0PgI6+bym2BbN0P74IUHu3VjvbfJIgRUXhSo
zKA0W0+Gp/QvG5Vqu1BBv2Wa2IKkzO/qliwX/JQOFzhDU1JMbbrkCKxILEs2HYvuy39gVlMkQ0IN
IQTx+z4QhlREcWvAjzsa0MrNnmYeVHzpzzLF6oa+IdQZd5VMDjISEGkWfAt3KixlBcFBZNU0PK5N
PF1GUJqWiu2JLYvTsDGqPBaHGQW+JyeGbj/RRiIBhcIgeRFAeF2gBENS+uVbZmA9Uys85zGgw7XM
8NuZJbrpDQKWcok6Eh2LEMNKDmKRJ1EGdxAfT9uedhVd7p7aLQv6mxmRrELVba21DBvhY/AKJYbx
sihvg36/CueFLs0Gj+NWD+ekmluGcpf1WrtjRwX6w1iwlFonkAGk+M+5Q28uCizSKPL+R3p/z7J+
+6NWD2xH9Lk+GsUvnDy+a3inbN3kLsFHjnePEtUOxRolNK3zhKUzUNAXYGRmyooZMsDAxbZHQZH/
xZexJ+FvQc+nmlkYKQlgT+iEjuajFENtedpgy24MVRgOI3nwJpXauh628T9Duce4bz5/vaIqqJSW
Ki1ATYXf+yT9r9o/6EIAABGSNX66/mqxWVWbqImNoEdTdk7IW22T1tRfR3kbjGX8WU+ETzJ54xH7
2p0XS2nYT4ChU03HwctfXHKo8p8+DdTpAvGC7igzyasp3lCrW3WDcQLC2TLo+Ms2beQs+x/uuLUo
nLfHSzkat/vBYl4g9K0679x6rwyr1BdcfRm6N+pHYkunGJTmywK7wToO72JfJkpV1z5/rde/QwTB
hXDrsjqGy6vEJjN0Jq2XKuhgs/NDENRrp41aFCAIwH+nOQdjXkPacGGiNND8odQp6337nMwC9Vu1
Xxb5rLFwfproMiLCWkc3Sk+ae3G3GUvFDz/Y/SMaNRbJoDTiQdHE540jKHNOzIQLDvggTYKYoREK
7esbVRYCpArDDtbU40Eh8f9gb5dt+nqbToQwTZ7hfjesnMUV6bG38vMotZLC8JzBUiRMoJBzpSSe
QQh1MQpWWcCKc/Mh+UznmkrmSZo/9KArO8h2u2QCjNLMU1dMdkbdPdHoMLT2CflkYX4e591UyLYB
gquU4xgY31II5pZJE7OjVULoH4pylMxD/aHvAC48Xdu1QW9F7OXPtlJX6Ec6i6JziSZymWG9ZIqQ
IHGW+GxS2a8NmbEGdA2WTh+FWmo/C85bHlTByt07LdBKuyW6t8P/kjG7TXvNIbcjIbIt6oB2XiQz
LcYXTxHH8YP4uDzKCfqM5gXyrhwRa6pCQ7gg0hd9mN97zjXH/gLdQM/TZCoO76Wj0wgOJNiVNSaU
N18rzJFGqgGr1hFgQ96s2GDvoCeaSvRQQX1StI4smjVFwq2mNJqHI5XbDM666qM+EknQMcYhKwgX
+cluU2aD7rSc4fGhoQ78xcXMLIio63IVlsHalCN4c5JJYhD9M0gUBLd/t+e7uawwDBjHXOUM43Cg
ZAjbptWd4e9zyhIxajKOK5t2bHVZIQRG2F+dVfxXQFkgYH3OIpCOOn7r4/59uJJeaN5V47vgNG+f
bgGVlHFquSA+f6EqFLPA+GFBoZ1d+4vU7kC7pT9/ulc+u6s10N3o7NwKb5u8EicbHD80uez2Q21K
s/72ry/aukkOwAW7N8WpRdATgqsZeFpnAVFRd1gOOZIq9SIURIo7/PAnN7oHqcadB6wyMZr/hP/2
Hgqq21P5N84fuD+/zmK+XKUbPsZcd+jBg8OolOlSOCi0EFa1ZkKbuwngXjqnf2p+WKyJ4vPJN7mh
aTeqmuOCS2HYG+kt7j7/HBBiJy+eJiCq3oPVeUupTmLkGbeIyCsFzV2Dv50XI2AzzROq7+xuPbFU
9Fu+XRYd4MhsrfkKdUDHrM2QWxV2jGW+OyJkd9GsJMEhh72RT8aNWjWZzFMSHG2RUzM2c1IaIuMG
obSm4QMud8U9UFap1cWwYKWGgc8uq9dApna4l0/86vqbxGZt2gqvZPrDxEANh+YtbUDAEt7tbi1U
+gcEU/+WZye5RF0r6hN0wdNp7ikR0uywNyJaUFqUGZc1rlR66o1wLQbE7n910KRXXJTNYY5ImatM
RK9ascG6wGEdRkkQK87qjaPPDg2BBwBn7bKwWgI0lqTSB6cbReJcAOu3hZ/MbFbFJpo2Q8WQuSu9
ainUyvZqXwdx4B4pZfX1yvCh16PBO/xSEwMrEFZdqaaOSBHQ0uz4UjWogNt1RmwMhWEwzYzaUHaz
D0QEt4rAU1qjFnLC+j/vHfbLRmxVwi7Cu96lAliqw275ai5POJGz32LmVZWPg5/xm+iHnJEfkBQx
L6DNQ4bpn/uZz5/r+MCN3D4gTASYeAgLv/jYdNhEA/GEP+47mQC4Bs1hOuIlDQCG2FWGz9q4iPwA
H61INkW2OUGs/AnDDWP03qZ5Mr6Zj1W/W78KEfa3YZqCX1TfLkuLjsCRYUkIA6EpPIQERsGsVPUG
tiKyr+idnqUdGfjvXv72XMUp+MZ3BlEIMsccgoE7Bd+y6rk7WhhisESc29M+nMrk/VKlNO2/isAk
dvCetTBsGYkFfhMyY6bQB32Ou9uAT10RI9OFrVi8j6U3L4RpO08oIQXus2ZuEz6L0lwtjAaU7Imu
E0+GQ9BdZAQ1sopAs2hR6hPlxgeebMTzns96yHtKcvndK34krAKEkq8yLJE+RvU5OUaEFQjagd39
S+bRh07mxLWoCzIew+AfJvjA6eEqfif5qh0wCYImNY80gxp/SxDhDIGWp/C8+Hfj8rAEYk8Wsa/q
lacvqL7qrcrgbF+1QQ/5pY3sZvr91ApCkapswWf3YaO6eduUOFu7M8ovpUqIL5HnI092TWIC67+k
0k2ut0e0mEZMalyRkq7QmqEmButGHCR24d/wIYqqli9UFTmMEtl0rLlxTf3GYJN/efAFmauO3XWd
Yro9I1KKR3lIcy+R+ShMxridUPL/epheOFRZ29Opwvwm7dKG7UyNf0FDVCqeE3BJS3N6b7n7uSv+
C4se+8kbLh+Jq8yZJBoNdcrBWWCeD6G/j/4k59VUIzYMgMt/2ClEnXiQQKBwt6sXXmH+4FEUXowp
98vNeROcYkucTyGRzrqU8G7jy0UHrAcSsGv0xCrPsSmFpu1p/BSX7M0TTTnTtpqJVUJXea13rn89
rxfg7cuGRREwzi/5Cy0O8fM+BCYOt06jNfXBhv9+PxEk3EjED/8Gbfsi+HAdQo2wDVlFIgFTQWmE
sebsaZ82yIlGcIUjiXV55aHDuBySy5lcc2GAxXHqE8sMZlRdF8ANAw+ywYBLUdy3FHIrkisz/VZG
s+YPnnlrh4Yq/pyrmQiiPGKcib2IesiEAdO7mDYm04ITeSCMvYeKmDguf9iZNuZjW/kfmq2NIt+r
RZuWoxUWTjuBJn9fP/FGEL7xykHKtT6kcuZdUyNToe7enqtRWyzEdYfgNP0MIIMILmsj5gw55qkG
9nq3TY2JBqmimwwZMZb2UphUvCK0M4ZtYfVxGwu+yb+dqpxXoe8eURlPXY1YESW985gVREVqsf4k
74N7OoWZxXwr9k2BceQWilBTdCImfwatAJ5csvswQ1cg74bFPtOYsVxezcy0Z694eIAXJEI8+SyQ
iMWgy0LkQUDxHFH5RnY38LDPWbVTDvhRSyWFu8eKr/DwTrlzqV+ZtHsUpeglpS6Sxhj+13d9LgRi
epUSZ82PXYiZFIZdD8Ezz0IDYRP4rs4xEt4qZusETDqAaOvB6bT+/t/xQfnAfMCjIixOHb7bd9k1
SFBORgl9swLZpzvZJbPDHry/iDZUDA8JIs9HFLrOElZxZPGmA6aHhDxVee5nwxUXpc/mYrNxXIFr
6K+e11h06oIb2lizFN/ZZfVA0+JrTbZvIyJjLkESQHwTTfb28treKSM+KoeNHoGuibRmWP5ZV4Hy
sMZ+D/uHRw3Me5l5R69XaO+SJlSMXOXdEvEPW40S4i857LmRszF8rZaoYzoRtaQ+4Ep/CYQc7JjQ
9oA6pHdu338IATD3LV2u2ih+JiX9iQjoPolydIwiiiw/NGmvsfc01wGdoJ5+5/RCJ6Lw+9utFbOS
NWEqxkwNAb/ktYQaHl9uv+zAmALhhKTm+1c1708soMQmclH+RljrHGyfmzcOg6SyAz0N6/Aq1/rS
RqOw5N9vNw+4JEJxV3bDyT04GEZAueU72bqJE8bcR0cvvH2gee1c9ZVjq4NvUb7wyVuCZF18iTAs
Fn1dHHbczcCJLGdjWr+bfYrBDko79M97sNMoZU1vhNeNz0SLxUXUGVNSxCU2syoJVDBEfYQGWuha
GRQf+FgXp/q+wiKjQCD3XmltQ7RVawXuEBF61GFsscE0BlAcDcQL/hAHC4n4JRyFvpNPMZGpd3kM
sO4KuDOdNR/mMEfymkQCZmFMJeleyuK6fUP1/rw9XUXV7vsryTQwtw57TTFSdKLkzC4+4wkENLvB
3yX6scoSH2aOypGFHqQKoA4CwCD7f+xBcb4Ut3ZUSEkSMdeRD4LVTiLJkqNhrC227cf8fCR7LnT3
edgLHeDid7vYc5V6lLeeyFTwDakisOXWXoWiWeiFhSF+WzdljOaLdLNxTruwh4E8jmGMldKOKqdp
GWziLlD8JTEqAV4DK7UA98y+ZCGF9ZuJmy0RoYaTrTEMiraxAb9Wkn2vFwOphZWXvKs3REirjkhE
Y5gBWSQQ9Xh3YSLEtIL/dGu+hvKsSAypaNERdygIkDJR7yZElqT8YVOZr6u8UY5mXVIJLxQJ5f0M
8lA46bCqUGjQiaT7JvD65zaAT+UKafI/YocxFX+t+LAzBoYhxxZr08zzLOk6U+ahGY3CdU6Sj/WH
UidtbRK4910FkkqS9ss8O1VjjIW8pF2pITArzJwrtfc7+L5pLdHyVW0GjIh8FXnyc+6z8W/NBpvM
Rbd/nUVWHn3InKWaHSpVNsHcu1+obpPnmhM1uarpdNbw84sKheCS1lfoLb7/nZpFOnAL9DDYU0Rl
hThVi8gz083FoYMN9w3ybdGgChWLSo9pym0/NE19Hk5236sNCoFd4nmUx99B6Pq4033iR0e9y3vj
dOclTPj5pJzhIcRT1MvGn/WLU88UVXAhTUMcm14hL/Vjbuw91ueyYDncckVUXP31bpG7wHga57qt
CVs6jZgtdRJNAqT4ME1BATfN4AMBJ7aeagGhY6KIXPqUMh5Y9Wyl+ev3c5aigmbio998BJtmftfm
tp8R3Z/duXwCggFO3exAiCmFr/pLDUAsBi2iXUgq7Kzk6BJD9ztmzZ4Fg+2Sx7riQEd0Ucs9hGIr
/onJIE4991s1OfRIXT2ugXs/MKPKn2HmL2KDaVCr5grdgiROOPyC63+BWI+vK8BtB+KPXj8o1Mqb
co8eds+RuWRWbKnVd+xpg2rcfCU9RhiDfaUTU9Le+GeB4MGCCRE7BFUlwAKsgaeQl1ggmwFhJNzc
78Ej/nH//884WH+CFSo6TVTvwapdSHyY7+WVAA2gVTxTddkZbjcKMW4/G2Yl9SveIDkH3Q+SjHUJ
ELRl9dHNYn5XIP4hQnvdTYG7wtocXYVy/JEhMQ4vyZs+5WLTXq+aSYDp1lABc/AuCtETnKCpEnMc
fXz8vsb+E1uINHvACZ1x69e0RI66qJv5hYGQSYUIkqfBPobYJVDrNbr1eugLQvkHyIjo0PCxVz7L
V51LNr9/Ty0QaGhULKuhGyKk6ecoPgJ4kB7lQvwLguNIGEoc/ZQ3jzZcVj+nGQ4BsohTA52o24Bf
CTs5/1snJT2m48K/n/vpHbMoctYaw+dOLzxxp+yTpQql3k3BsIKgDHhIINCo+Lc/4wqzl3n3ExMM
b/XIvqhY8M96RTHuJPPCYrigDeEmWbQn3SZzNxA6GWcOQL8ZyJDtdXqecSHvbAMoAT3fySAFAnEO
wTJvO0mVerbdRhbVEIqUKChlz60XX+hTLBVn1rDT88pyyVqvbtJYhBgViBB584AFAHeyDo2fHU2w
09iGkEgYhDxTTr1jmuC7DyIEa4OumWzz9G56mzRsAwmkioGs3IekjAqLmfFr40Pr4c0/4HkT7UAH
eSNbFbsNtAHZ+TXBTBQeEVgiczw4ciQUWEAKD1ncahYdn0H+4c8pS8x2TKLsQzOu9iDoFv8ydWQY
AnUTkeR+KKBbQ3VEBxyjx0kwt/rjKdGBfOeQ2naDthZPZQZxqnfxB2SZADU7ZEzoUURqJMWZizUU
//fZIDo3FgI1vUQPNMniINVxCGbJ/BOmeLq096KCWhqAQCw4rBIzbJL0pt++bdRWmZix6QbXHevn
O3Rlwy/C9X04A5ggqrhk8SjTMAHqm8LT/FOPTV1y5rcJEYh0AkDqBQkWz4BN4yj0RceTeDhFsjYj
jmjr1MbLmxUjz/XbHZAg1duaCiuPlm4kCrg+CMmprTn1bybRIFmgaSyXHcspfRrnF3S2crEA/S3Z
U+2bN7U1/IDtOtYddcixn+9PqVi4A2hTDpQPCsq49VS/MQV622Zpq7G/+cQJC8N+hE8XlYXFwUoH
Kk7ky+1Dhdbs804V0I0W5wKEGB66EDJibY1Jfc0sj+8RLjLVPntlpu3S6fPDfjnxUXZMdoMkUkCX
C+DsdtWm9TPRcbxSfautImmHaGrqBwPUh+6bqJ0AivjSf55xZ1EpZZrsy8FyDwya5hkNOobALr3c
IyMvz66F+gbp2AJQNxgd4A2qMvyHBEe/z0b/1krdNaaxHBdI51UvtawJOry+CVd6plNK43T+rJIP
T0vOqE9ms+6VV+oYM/nt9CLvcBs8THErV5CK5+wdIJ1WmPTCBlT0p1n4GE57kPaG/6T770x4Rl1D
7vfcv/KFSUWtmV5Tn40ZEbP9Wd+JJZit+1w6FPFSaoE4RH39dxVzaTD8/9KiJGKEfp7HN9qN0EEW
hzYEi3218YbTlLN78tZHHUzCrmvZGTh9St0/NKzlCw+qM99PznPz/4vA9FO46fv1J/8lKdoKBgLJ
puBDtxnhF61vdwHMQD7Yd+VHPnSCV+X8v7TRXgDiTwGd2r2JEhnZwxmqD5NhCasQ9rDmJ60OKHQL
eCm7phscrPjCxeG8a61il0YP+B8HqCqAzVcxl2oWakP3NIW47FE8sLEmGBZuOT7PGN+QFNgpDkIG
v29NI1RZ02FLZBZS0NW6EMfcdzGr2drJUPDa0UzAGSm9au2j4iq9UtsE0GJymQxQmQbnaRF9q5AI
x1wyF+xCiQ2JozIj4ceSHY0GxdkioFMf27jOt7R9KWBdyDd7aP9dSsLAXeW9BShuHcI69ASKC+wg
suLv3Di1J259u3kYSxWLys+0h2eZ3AgggVpUd0fFbSGhzO8Y/IGDP9/SCr7ujw9wJ6+uuq+kR344
IYBvgzu9as+Mhec42UuvmQ3HvwDfECMLmUhwBCARrjeYkRI1vH0sWM1WGeLJYIt7fqjarZknT8Cg
FBjxJHGB2WslBXCUXLVfGPJtJcLSJTLpvg1RmtjHfUbKhHijxZV1bngjbgr1SVPRHLyXLpiFMEBw
ZPIxoBpggN0Buwu5JUG/KVJyWopccGWw8A1mClpqEtj5ewcoNQ7XRjXpfCzc58UrZZB0MQI/kYjV
7KxYgf8it4PMHIKUOq4mCtyyR/39jw8xdJ8xNzm7U55Cvu52nM3Buq2toXNVg9hkyxyjAyYtjD9Q
2Y3nN8FvpckTYuJo4PEVKtikI3p0tvdzhrP+DyLpyh6wA3LYpCU9c6VGbJnGbomEFRzWayHOf5B4
w8gmrlwBZAorKj4D25HqP1XP5OL3sOSwih2ZVRb1ez3+OmFWQV2fJPCXQp13t3OFux8Epgo8l2FR
P24jHzIVLdILOPBwEqc1QSK/URs0hwaZmW1go8Er7+5/Iap+uqfYM/IQFi65wxRzd/PXzzwKl9wq
ls9pRrSokKjJKQmzMyK947ynSo1Gjl8yJTsso5a63YlmpFAJh4s+AEWzoqXv3qOd2Yamp9oqJgNL
4pQmrx0jccWY6WuAz4hZjy0M6UKgqnL2cj/fOdetj6VzVdZ1fbT4zg98Ugd3nQdnzRYf4rhm3Ot7
IrCb6NU0QXHSzD+TH26NaJ2A3T9cJjSmFDN31d+fahTaKZEE9pHsXPF7QNIMYzVVZFTGySUXlNCG
XY/rLbbFraCyXHCN4YdQUabl8GlNd+ElRyPUNtRrso1dxbob+vrmCUKtieFpWJLRIURYJhFBxomi
OyaDLafdxlXL6Zbg7ZR8Jn2zVMPW+Bsfr3/F8JNg/4hIW7AeNoP/xpdZJ1noh0kPzERagIKMxWUh
Vw29j2DfYVueJOfKTtuwoSJjuWGycfyceUiyllh3mOi+I64Y6tdGjz7N4uGdU2yew29eKkWzzAfA
SxEdOULM5tAvp4PWrJAarGos/blt1Vq7YOxxJZ0QwaRrGCINWPuDbUYS55sN/9qVu0HlC3J6gGwo
SimwHQzbQS19VAQiCVBUstCyTKUm6kWYga5QE/cX+lVPAXZeunPsBUSwgoMZyHmCTl8LCv8CcMjo
WePQ3CqYrihRab451ypW4HaStw4CDMoAr0gyhKhnIt7Eb/jgPCtuH4oHUBiDLic/8TLlPJ4V/UYC
TXY+0swLxql8Jq2Bw0+ALurTQR3fCWZXqMua/K0ojmBo68fzNszeBu4iGWRXuNOmbCbFQTROlRR7
BLxOQb/i5Ow+56kxyuFWhKSQ2Tah3nfV+0oZoOVzo1c38uc3ISEAstwwnYDVzu5taHukNLmDx4FL
HIMERzSsKGaqw4RY/kO3hu3GTFLzmOfiSlx7094v+hskcvU6a0AriGSccG1r14EqaDroipYS5biS
B9ue0ysXVaIXlwJkS+7yqq8EfBchMffInqXKhsVzV08wFTSoMgwGaA6mzJ0Bw5JwLVr0HZmNZqyZ
dV/uBbrVV51wPQPr6xVvTMNWfI0rpz+RB1L5tKptZS10/BgUP2XuiUPWjDv3Y7cxf4MxRJi/XChu
POxd6iBzEP7rbgRSHYHixUoBKZyBsRC1QUvDumPszbdKKwJecxCcjiM8+rIKdvfuk8Lvt/X20ccA
GZb79tKN90sn0i5l1aLTYb2indL3yEl4NEyfxX4z6v/HlEl+Gk5TcRN8Vx34QOKRUN0Jc/9+IeT3
6XI+OHJAtdDvEoOY2xW9CVOpeiYSTsNpaexXRndJQAcM8BtMCUlFF9Oc4NrCkrIRpkcU8g/fq5Xc
2G2JnNtOuKesatSbppKQgHVyB77mEziQyJ+PlM7A+56bU6Qlagwju78F43zygH19A9+AorkBRwiW
4qVQMsS7hzT+gukoJ9nz+BTza+mzemHPMeOq8l7PSZ8Pi+SsPvCwPeWtjzOpTcT4gkz1TVz2D8a9
jREC6foEOB2MOnFtghTuqAQjHNWbp4ucwRj2S/+kzh/yVmVsm3W8RdokGLCcvG9PIOhMd6oTJAO6
YmIDDk/dpuxA3F5BwGM/keGQJdng5sTvqnoltcYmXajTHU+mVxKk4qpfIgwvTguKP7uQxHFckdrb
dbl+lH4K1tDHK67ZITuCWg82BMoptMcyZP1yNwpI9G4LA3C0sQqzqgRRZ85dRUtfOPMZPrV6U1tr
Lek+1Y9VtGL2zwGuobVyKQCKXmSnPI+kGnL1+hbusIoOnznqmpwQUBnERMCPZXY89CN11F13ORpT
W2IzTMOax8QE/dV0IkcMuG9OlLla9Y7LlMb2V/7GhUBCcu4iSYVsjakHIJYftCyUGr3iABIl7qEV
HQrzAd4GD7mGXwg97nhCiVqKFmjuoQsUwNEqJ/13dgn4wtMqVg5Xjpkzf1p6gqLR01WtQGSnUl/u
87UX3Ol2VTfK0qOKdo3TXC2SnjTEHecCgA+COFKnt1QmBoui7AiCyCrjd7lCvt9EgO2L9RW8a7NY
b0qBLe+XhxodxL/W6YjcbTXB+Sm/bfkKdxre08Z34K0ipFbqmeHy+uOqR7gpB0WLGQfM5pz6YtgV
32o2AoNnTUOsde3rfxcJf6mfMJdVqRnfOosGc3sdQTvKCXGR6n1ib4G5BZzKm1Zed8ZJuq5Ja01t
okl6lCdBPnGbFPxn+GmgpD1dyBEJZnckQkmi8JP3ePoNWKikJhjwYXNSSxlvjeysN7zwlLSD4X5o
ZGuZ0NLFp6KFbPoaaPEslkAfRpnQZT8cJ2aMRD3B4vPSmtLLnxfViKFlb8st8R+B4OXAxXJfIuDD
Sxb9BsD1g6PttaYD54553Jg/ffA9RDTAQRhMF/f49wNXYbVor19iwAbd1IBJi9uo5IfuvjD3IJi1
jROrOT8pLnKm+3hTstktq3gtdf0gYUS+co6UqzmNLWPXD0rG7giYVPdIOuax4xcjJ9sln7yMpewS
Tf8WO+wojRA20BnM1UDzPMNxKjm3J2pxQVoDfFaa4iljp9LPUFM0AIajFzRDtxwe+M4ZRO6I7akc
S8TqZlskFJW09ETTT0CsHeUjHGXofeQeSV4PNy7y30WIzIzrXBt73Eyy2WtPPJWEu48xIrpMNDfb
4eNVKpZewIrBh0mLI25mt49vlik0Dea6r9Dj97UyIareJo7HYklYmck4o007Eyw06fhGd+XZb1wl
l9TQj/DyzwsNlp1au/NhXvUO5keIpPRmn+tCYzkOMG+k2KVoVN/Yr73eGKYtgu6L/02gAO2FeoOM
h+rtgUpODH+YaKViQkLecO/X5WbKxKrk2oPFVLdF1Ges7kpC1JE8k0XhhWJZzAig9BX3ZAFtLMib
o3RnCwTBQ1jEKGNZMA/r0bhOY6ArkQmewjTQTarXyIErDqEO5hqulbNEr8Gq2UGmuFhXBiInHV26
3IZ3S1GGQ5sytMqxHYxRP8doxS3Dyq+lo3GnfFQa24v/c3hDlQT86jI40FB7G4fEJKK0kDvjMZYg
KvO/31CEZOvhr5bq2yzBgdEHXD5txJZ0kIbtixox2yqLA4/jID3j5E6Mo/uGBuk5fgJ6jcv9iSGG
7suZiGzNqMVkA7OTyNyCSokdfEzea+riXDoFtHvQ5tfzfwOEPnWOil7Ti7Y9/XT8ReH5dIQswjgJ
wHQtsiusvNlWoxnbTrPaJJeAkDmxiiGvYXmmDY+IW08fVEe1tmtOz+c6bqdVSFL46bJCPvyPUOFB
F9uFbUG/wY3PwlbVZMJWRt5H/cjNJBoC9bhZZ7W7JY/snZZ/2s2ZbNh5dGPNyAUmBH0HeQiNESlv
WpiqSwiDTKn+PJ5j1I/f4aaCbTuo7qmgrNkotMl2BqmqE/S3Nkyil0b8fsHzwpjiu8Fj39PNJdds
uQloTCv3VYf0G5qglAkXvHCeG80sPiFTDlF7t6jEiG2ZgH7/xwE45mRv6NUXI9yCycMHhloWHgnA
XuLYFIFG+5cjU3acGvP2G2ipG3IOQKluAcYxBKluVgnL9BqaMOmlXbPAJ5cqwNs14z1L4KQYp7b8
fVHTC4uAakUAXzn3VM9zagLiW1+pM2BvHXeETmea1aG/dDs4kPL3Lbl1hFfQE8v/sRmsVpMRFqCp
TnbGdMKtkVLAPlq7FSG67POK0j5lNLddAiFYw8kAJEw7eJpjMk4+0WvkENmbzUHTMTPgwaHXFU56
gvKoKOno7RN3XlBBBL3meU/Oof85/iMI3213NMOy5q3YOmlkQ7dOSkG2/R4F5PQUOjMho+zj7/e+
5JUWjr+hOAvon8VMhKPq+hESKrG7/7STT/d8yUEdYyKZSFwS78SXZxaoAgg+Bvk85wFqI2fkA4ux
x/RBs8GxKZmGQa1stJlpxR0xjP68sSYvqjOyxnCedsnDG5t1Bwtm92rOcu3iMz8E9sjuiLTIH+vb
Q8qz2Lfbl6eEAfT/o2/kqWLKlNHp0IhFtqGZk4FynfCHC58HMFw6Y0wdMzToCEiyyqn4ZMOENyHv
oN4E2mxdS7J0jL10muQ1Zg+5M6mNojJ2OY7AqsEsshBpYf41aw5Z4wUOGkN5Cf+65lnshvv3Zae3
FHu+JpXnETQKjv0hGZKMHVN3kYj9W54fscoBLH62OjSOOlfmk1sc1qSfGI+yIdI0poMr4QMskbQK
7tl1U6gQHoA3Zr3z4qM44RBiRyE3Wknr+GbBMKnEo2j+f8vE9mRma37HQtTSXW5AM2bkdAA1GcDK
m4mdNSbfvXZTCAL4u/HM1Vj/0xBloNDHPKzfloDv9v2dQddOgpue6gP5pFD+U4NtEc8QMKySopHT
GTX0cd4BPr25oyxpAGdtbfSt+AqG98LwEmVwINDwAUcn3Nj9aovaBVuOQ9cVNiBitdHCwp2PbeXK
3RIi2urr6k3MPU6YbesXFyPimESMNNbW5I6KaPGHqpUemLRz4ky+/X5jrdxDTJC8JPxbRRu8lWFg
vGOgLXT3NdsfyNsBtskberRGUAkT8IePvtU7J/90+Q8yn4zFODyJ0PEE1uliSeeqNd7mlzaB6YO+
IHOc5isNsc3pa5NAqrQp3yHr/g3qeXl2q8AUdu2bKepgOJiSqOrARS3ZhfYS+MR8lGnsBbUA2tFB
s/tmTP8rtKzNRuhQJBNgOT3TRLzdv18QLsqFyI2yVThWzvo9FUviU8r0PT4UeDsvj9jA6lSjzCDv
GWvaZs+6xtN8UvypxZRg4SlzILX2MdsNDFe7vSXZ9fkl9Hc0nuqf/ZUaSb0BXjM4/uI0AuEIJLL4
BWPluGN61TO59r/NVZdmVWZmw4S6icsobgQ8wthxX+REMDL1CGRkCmR1Xep9NEx894ar21FiHd61
OfZoZ54qeSx0UmtaU1hx3Ns8tlaU1piyfvJDmS4GqCbqouURaBU4wrGZ4WRRBB6nPNj5c3pWCq8i
J8rZAI7VKfqR4XQDACwM2EZkmXZQKDJWHy4YcZIEsVdLtXQLWXqfvxocoMDZp0BxG0WsdrcgSJoO
UJwqW8QMcLbki6nHhh7LnXLrBJKvuWf2yaDluDmLQG3Wd/yXk53XuGcCzkjjFDURbF7Jvm4rr7zQ
eSvwQFpadak8cYmIX9WFVPDDGN7Pjliu74Z+H3Cg09os04oG8Kfg5IV4d4xxGvV2R6+rLyJgOHC0
J9GvvARANES8wQ2pL7nM2lzT4eq4U2yAyZJijF9Q5UdO75hw5FnBHp486lYpORjIzsMiMy3wZmwu
zeKGdVJ9u94z+r38lCbhgp2DeKUVZBrODPuUqkhBYVIi437sEgtn5J9h35UfEJzYTWvbKxqwgbiF
Ot+LVMIyueLWB/55fQoi8JK4QUc1yO2aotbsTMTlRfckl0g+qcNbuK6PEUKZ8DyfaoGmQ/liXyxE
FwniavBXbykwkQWeVasXnkKSISTTT3qub/WQ3BWViAJ0R4/elFUcOrlDndunUEdlYoIj9xDHbgPa
aG1e1cTwsxyEMlyAFZFVtLKEIFoGmTrrwNuIzPA7WiH1ZbMGv93mLpSUx/37WeMgUFmD+3kxkGdj
/WrKLBo6cLck2EKVP6UM03Ro44K5OkinzRpl319AV6gYlN+kivmIRhMcjXbBkDuTahDPw811viIx
qOezMEeo8gjizKyySx1ZyrcWM4A2adf5Z2t2uZ+kziLyCr3rQdJjn+jjFyi7E6u03DKg28uD0EYa
WlUArXE7AsCCUCYqH7d7/Xx+daifZprz14Dtnrjj0Y8T+Knh4p89mpnyZuPtGShmflFv+1X6Can9
5fMKlTsy8JoAcgNi0b5SOedz8OhwZRFo4jUEsiJmLC+fp92o/AN3dhSdAzS+jEhvGEeJ/gNv4g4H
sA6Dl1bAR8rOXZKekyMLIaM7uNGWurKmxeVHy96/U+4OyTf9SIXP06qdqvGXRHiVlBN4IfFycWvB
ckq0fxDu9fWklAn1IFOtZURDsfCSGQQZhXKWlg3BJZJVpzUMo2kVD9HbZ8Exm1ZZ96yqe3t4vdLN
MTln20flApAO9s/7wXfCMRiFVrnr5Q0tqkZSlkk0OeFzvm6/4+n19RrRbL3pjElzUApS8vM+d+Ph
4+ShOgeagDEfI4ky6/T2zNoy19EG4jqngHdF+Gd9uhYghbudi53Vug2sDAm3hBExs5G4h7qRJOD1
mOdK+jN5t93iCDpj95AoI5gk/JwWUu7/rT+VIoeZ1sOZITiE+ajXHmdbSE0NvLLnZiWsW9OEWS6n
QCM/knbMq1NKWLmHs3MiWRv5/g8vagaEUztOuVaFRdciwm9RBaQjR+Dz0MKj28k2bCGGEY17eJg8
E3owHt6VdmlmSgcyyU/Wz/mN2I7UCWutSHEmS/QrAvE3juCF3aKwlDNYpIh+G5K7aacjC13MFty8
tsjCgjXE1C0WWvHziHMOtFhF2Tq+1CcE9YTkOabtJ1o+RVng/xQajD0XeJhaNQ7PXzcaPzywMtTB
BG05PuIPNFn2JKFUw6NE8FIDcZl4vgrc6oiVUc6ukLdJF01HFhcEeAptb04miO5/EoAqimeC1f1n
R3d3OaR/FxYEVhBNPATXjn1cCswTYyYVYxHZjUEyaJMql/z64lzNtu9vp1pFWbAG85iAhF0bNesc
TvKMO+rRqoADmxeQCG1dfkePGKhGuU0AnxR5LLBj/rfz6w8r+K0NCAm9He4MnVJtJpAWSmXKzNRE
V9Tz4ln2lxgNJuiiBjxiIQBo/qGhX+vzM8hRwKf1owyeDzAqARoRTpF0bM8JAhB+rJknJqXR9W09
hocyacv3ktq3ck1COCfGv5zxv/wk+EenLQQ4YK0o+V5MsnSEVFjWDha910X4kBVV1lGjMMOo78SM
Lp0FRVvRI8qC5oUEEVqHsqwDQia8Ph3PnE+d/dNqfRLD9qd68795mM3OvRXb7bzn8aYMQybp9Q9A
PWBbvsVs9daxhu9SqY5KJIt3r3EwEllK5bLwy4nuXQFuS6hfkmg94aIoZgeiWfvEVOJtmr7kGrTf
zJhKzjAG6ok31ttbIS+s12S27tv82n0ZvvgpJZ/4n+ZESih/DSt6pllHgIUkQZ6MFVwMeyl2HvIc
XIdr19gdlwiFMQ2LGPZ8ZC/dOfqjWNMInr+lueZvjCU3VFCLOdJBlQFM9vJOGFmIMJscQMOv3mff
jh1QIvrum1WMk6VfeEpdVf3DefrbO2OjvR0tmVK8jLEFCbv7f8eAqq41pgpig2FA9o33t36ziQOc
yt1rq8OiB7xJE/FMjTa7QVpVMRNPNZlSNGxTigDcMhaDKrKhyZSgmHKJI1gytlg2KVRQGI9ZukF2
pAAUKLiAkeWNsj7GOm1I9+B0QPLYx8gWZYAefHi40AS3vy3dw2RbLaOb/zD1r1uSmYv36QK/D92D
rRGYCj6tdn76wFYzI6NbK/rzGAiG/B5GSHXdqpEfGZeKXjo8IEKbrPsjqF1xAB9JbjTrjzPkvj4E
tB7bUIT8OEKwLWr4MLDyOWVzCOlEqnqWEUr4V1NoKzrC3lKKPBpqoDPemWSJghrI2iF3xsV5fuQ4
+hqXKa90YCcT9uXvXbLG901N0fHJxvOJZQJctruzgbrQiIaSjlZZzD0b6zXYu0qUnOastS7gKkGK
VR7tvmxdO3PS8NtJuvdlTg8j+Pf3aWdgHRul7ysV5m4A+sy5jp8PJS07+2Db+xnon/9WuOr+uDuv
zmT6H4rW3QcQpe+kvHFBWnljci5g+z1L2u1T9ca2UcylkBjJSMzZt2tay7Ec7c2Q2ksLlin6OiQH
ZhWEMTJ/r8iB1C5vhZZlahgNkVB8RzfiN7qiPFZICPnEf0/kf5+lsYipf6Ui0uACt9UDWtpAjd9H
J+GdyypydxjD9bC0GACaugPxcFVgNTNJGGYuTCl3a3fAWDnuHDgy0hFCKeMcEr0GOC3t6CMgEIXE
791f0jadYwBagWCnB6zwnwGTsCU5LkSyXkMf+PzAt8+dqBXc/NKM5v7GTKYFhLN1gM1isTGhB5VI
CuqtJI1k+z0CVYw6j3Kry3AkgPjcH5QKsi9o2tTND+QXpWbKcazRXz6uZE45vN7gWKgS7Nk6ffYH
cjkqRC8mrIBFGuswE5Uj/n4OSBue3PXNkUerT9PaL1CE43cUZQ62f3yoWSNfWWCh3ddiEaEAzWpv
x9OCgzYywA3I0gHZO2CCQ99AonPfOUCa9jRpdrLkBS4AXn0blfM4rtowKyvOrvqu3v12IIUwFBwa
BVu1xP8pI6XtKMXe6TcVT54Yw3NfqACsS1OSEEEsCppK07SNrCQp/Dn3CFj15+/hJO55qdTp6+nI
Yip0PTTGrchHVRAmGmoR2cKlnOAhuVTPriVUD1sYGe+/BTg7W3PXIiVXBC9whf4uJ5Ki2AWPfgji
OV71XwQYym+JxbbIVcnxmENFioA5ea3PC8mkxTZ/YGy42D5xRpAMSknUuXKtxnV4y0mElZtR4tLd
tT95UykOSdzjiAybmJcHZyreF2ELrLp33gjJRTPsQyM9hvz8yLtp0lLO5aiWqaykqC1JtJbQzgH/
3InAOWbHSSZivaaFPM/Rv3TKA5ZzFbMnR5uLpX3t7PCILCc5RYdx8ZjQHTKGJvQ/l7KJ7ux2MsqQ
gVpUfr6s2quBFNCwStmtkIVmL4bC2tHkO8z1A1Gd+Gth32pt/afzGWLl3PX+7q7OU7Xa5xYsw/nk
vsKG8oVGaXfWJeHYQk70Ls297kVV9sc6daRU6pSB8O7qPEx+96TSoownWAPD2uy1MC/UmIpJtRCY
gouR/iSMdc6yLGJaEossigQVltnAbMdLG+eqlw/2qa8vdHgOFqZKsP5uA/qsvE7tgFmLQFXeZA+a
SCUF1TiFKoV+pNwcrYxIkwhN7z70vQ3//fuJmEhm4jVPCP+MrZwr1EGqf0NyrbeA2WZyfDm46zaT
JvbV7eMbY8q567x26OeF6TFks5fMp5RIARwH4kiVb6O+GjclfftS+yJ/rTS8D/7Cc03TwZMLCFI/
KFU1nOo7hX1aoTaT4GUqGygQkrvqieU+ewBPV/jD6NoTG2DYLuhIZW2lL67I9Uu5NlzzM09TwiFj
td94T0P0KX4CncIhQJusctl4DBmN9LBr+aQsRwBE5W/wPtALPjZfKll3c+xv7diK73wII/0pB08N
DuvJhcm1WZped7mnJZb9hLivboNe2JjMwnXPO9YqgniwkObBK+Cov00OccTT43+Se9oYilQWW67+
4P+hqeWhzWOtE8tu05MZPd0SpVH+bM7LDF+63bRHMrkHKzUc2th5xXJlD6Hib/YmBrMpXJaxhSmO
ZFjkZH330rO/+C+BgLsdVLTx6zCeAMgIoTLyCAz20isRx69FgqH+kLuN/kAa28/t4Xq/JCnP51Xe
ttVXvVrvJUpI2XX1S1eSKQOS6eeVJwzMoJxLaoQ/pXTClipQqMDBNloSTx2JSrTmVAuAqz7Ki9ng
dIU0Bzb3xP7e0cGSfCO6wD9Z6gz+IEpcOpDE8HxhHdWuKGxxkt93j0529xJezAQY6TisQZZMT0GP
INk18ckDLmQtCKopvwjnAQIg2k10Jyr6Fi9e/Z4tGPqAFV4fnifFL2Oae8tvGw3ITtDlK86b1DYE
3anKWuFsiLCEj/prCf/8RbgkuMFMiXcXS3hDo5q6/j2/2ohY6Al9+b2zUlBWqDE/GI9n6YqFkFXm
cE7arG6kZ0sSsJHdYhJ8C/8Q7pek7vkrbs2hdrVF8qRuV1Xl6irGisEWILwFsOVPY6y7xXyc9U3s
UfCZdMG63E/tEwT4lU7p9vDTgKCz9vjfDG/0XMRux+p/0mTdXDtOJr6fHEHQxNQ+w+XuwXleO4Y6
CXd4TuTfS/OhqF/ZrhDcJkwIi8MJtAC50w614kS5+yayQXpEqn5w5BoIT4j+mYKGitvzc2jvd8hE
rVZvFQfhvVGAVbrVzwMEEJ2o8ZffoFdrYI0RTH02RsVAmJBeKzv+mKbHvmatOTAuzdFoYW1JvIOf
OFvZsL+gBJkMl5j6wp8w2EVmYHm4TmJiD2F8Q5UcYJshf9Q9gF5A7ekjnh4gy7JBwGFlMwAZUJ+T
kkLJsDQFl64gXP8Jq6jPWwZb/bdBd/eAsCcKM6iwr2qjoU2GkWl8GippHIt5vGJs0YsZrxuqQTvN
osHFMSgHAON+ktTB7H88J40jhP1sjipgcf5iLSf5ebHeBzuPBJmyzsGPMHyzVYBGInvEA0ISavKB
N6un8Aij+Wyfy17soJgwSzAahk4fCpBhQKft1JcjN5ojL4b2IRRf817YZnt/jpArWZelpyfMPyOP
o5TosCaj3SGveWG5E81eyeF9q5KzM+u9D5ppH26u+dcnL4CmSaNBYYREZBma1EztzGcmocvZupPv
x1kz2hw4l10m2H4wrM0UPnLP/wilXtcmzLGjSPqRWTLZUeskhwE7cbjwQQUEGSFhQ6oMw7hBwwss
5co+3+RdvkRJMxkdsJIR5pEC1zALnx6GpdztTv5K7YFgNh5+M2rK3kfW+gbpjlEJfD1sj7/+wDVH
MHjs3Ucqnwk8zl7RtHYL1j1PvoBMHphvmLwdwKlKFMH1Gg8Shw/AZbhWx5uPpa6Bf9MaU5F5hHY/
f732WFIIm8CHikPwqWeEzWfxZB5weH5PGU/TnY68fUurt4Z5vhDH8WoE4cwPctAl0a93gVRVoRY2
v6gE5vCTde54ZQB2F3k0AP2gWnudSn/2/c9qWvIUVht/ecoW3l2aRMAggDIveyVNRg0MTX1YIAl8
iosbbARbmLTYW3HuGxunQ+4xlF9qrQ6D9JPEZF3aBRQSj6CEg0nkbmDkC4tYW278xO58P0YcpKu8
oCjmcJ+N3T+T4B8Z20WadkIGEDjGedodG42jnlyOyqgci1tuDrckUludYK+KA8PFblA2Epq5WgYK
pB73QJe3DMISdHbatJXxBqnH/EjCam1lTzPmjX4lGLQq6A38drSEpC1izkE4/K1GOV6Jz0+sCYa0
ZmYV2qf6aBNo5Yl1rR4G34JZeXL8eBThn72UyH9AtMnkKrXIxSvio1PX4pWExm+OabsWAuUG+Q09
woOaC/39KKLATGlPBrUG16Gq0vRf3T18hXlW79OikEPoR0+e+Ht3LY9xnOZkzIarnoyus+ATrYWx
AhtALeSCcOmPbJzaTrXrmR7XwdJfIhVzIwiHU4vba+NmRK/bfxiWsd9tHfYEXxHSFil1ZZ2gHxcH
HjA8Ik6SkSUnCGLfEDuW5wfLhS0AGiLXEuWwK7AXffgmF7L0zl/2FdmRa1QrWgo+FxAeNgt8J7MD
A0xGSqImuvPrZhvZu7bdU1Sfgk0dv+l/Q9DNgEJczXw8WlY6tvk3+gWZHMiLU932Kr6B4u8typ/c
RBTV0lCKMpLmxXHQ2f9hY8Hii4md64mzPDHf9ehCi19g7gNmAdvCTzrXFEV/cjfU1aF/9+Ynm52a
TNPYIG251HyzwiXsMn8diXN5V35OWACbbEaDR+3VtaSW8JkWKP5sy8IuqMD/6N2FOudIxgv837lr
QOP44WfDq9Vn/lo1T9KE5dD1eWLq5JWHG1N8BYNvBos89tE2N5Y5eRBvRwXc5PyxhAWbR5U6z3n1
AWuo4qC2XjsgTRwGVIoyEcCO/9mgaVfo/uARfx90FtIhEvEbRRUmvI4D1hCvuYgIoOh4lHn1H8vO
beko4CkM6rGCQTgKe5orBszxKZh4tjDUJ+KiCXFmfaeaR1bj27frg+tPPnBa7GJ5XZvV11EBTXz7
c5+UFwkv89fEn8NkM6kr4Fy/rVz3PBAkn7z/YIKm6yknVz2i3yEOH0gmotB62RLna5g6mJsmdlkW
oPusEy4xmbPuC7zRxFNhYerpxu3F0FP112FVrgYPE3Klz92k+4L+M8kpf3gv4naZqakBIT3OwD9+
aR1jrDX6bMDbnoMXB+AxoIAo3BOTnCRL7Kthap3x3pm1RtIwEII4s+GOeDpzgH6SDP/lSqzllwZy
MvILGVYjglBreS9Hke/BQqAlI60bD4Jx3KKhmrgcCKh0OKaDrpLC4A3JEpG+Ixpfl6KarG2Vww3y
GM6TWVfJ4efGG9hgo9PhHSzY8yFE0OBU6pOJcoUHqWuvNxn9+eZB+tSed+Pj6tJbrjra/YGfBfyn
QfJ00YMBKdI7o9BY02nwc4AbYPgVfg0liZiLx0+3ndybul2HIOh/iIO4egTMSqksn8rnKRRFB70L
3QK6EvMwM4wN/vfn4TVguGXmgU8rpBYVIjpfqrhEYIwqyeCcul4x7WHav6sxhOw8hO8z0KELUX9u
nBIMiLLe+V8u0hy9znpBdEYYAVJjlLUn0cIraSxqbujGGG8BVovrLhxQuJGzT3i7qHb5gsBjERoO
FqUnNskAWxNFlpM7H+oxRH14jzLPEecWYmiyYcrCAhIjthCfdDa3YBzPO4A9oEpsZhU5tKTxnjBB
wZZKKnD/GEiNDcImF276hU3r6D++jyAH3wlrp1i9I7vf2IgjjWvMza8JLc8Rtx3UFSrdEDw0e1Ep
mSUvOyDFloZzzpHhSxIVr5eUSFOmoLdkR9hnSNTFhdeeWisAbkLN/C0uHFM00ba1d64OTaCUukgB
P2H7UvrwNLWaR9wBW2I8C5kgDSSiCzLOxKMdrUHf9KBaetmqgcPNcONBn8tOmmyAe6CNWFXp3zIL
ItoQrb//40iUUWA+0p+/jhms5ckCHlMcHyq6Mr8UHpvP44zLlAb3IW7FuMCavhB+hMeH6Yl84wOl
Bg197ZWew2OJ0ow7MgCFFdGukhd+qZmN+iDiuaJQ1MDsmONOfGOawvXJwLdKYgBZ7+8cAMmWiiQR
lveNpd9R5Z8Ja5aFcGo2G7CrMKOV89wBaLCQJNtGMMkvGh05tPOADAWzdH0D9MYg5iwmo0MNKAlg
X7oqfLxtlFxI7+s72lXKjYXRVC4c7WPcEff9vbsLqJC7bR3NF3zGvWN9NTlvklXaIbCkttPP3DjJ
Hr4rmV8zlVSopCg1H2AEcRMZMvMsXUQlpXSqixCHJiHXuEW1IqRjlCfmteRcAH/euyE/lFt1n8Nn
MWmYO53UWg0KFozF6stXJKWjUEZvWtj0k3dATiOPKrHie/d9kuSLM4cqkokVNdUR2hRcpOjDoxGN
OwEF42uFZpKZUIBZMXtMLlqonbR/OMCxmzkXCQC18SYn9xj2WYzG9EfzUXc2oBDZp5We2vEPfHxQ
NjEi0nF72k/+dQvPJuNjbgOgx+oeE2DLQicK96yArRIkV1nIyciHBpV9FB6aTPJ4XHkSKhkGjSo+
OtgjNTqgzGVsDRNEVaUqpRLwCsouBEc/MW4SyIlCU9WkKhJUCVh3FnpQWKAEj3LniHpY/PDI40uf
kHIKiWsosqhf5Szm1hntd4f2foeab0UgCmgWoK4Sgr3X/OaBKG+R+ZhlF0y7LP3hyqM7TkdCpwqo
s3HNjDhTTJGLlM9H48V6FigIec3nnjnOppKs5QEkgaBr+GsMZbyjfATxjYEc45uJHkZN4LmEeZw/
Fbg1+9nGdUyrrfYfRgMPBmD8bnWcgAnB6l7mXr8GXDc4AsRDx9G0qggfV4g4xvS5xMCIwbVgRiFJ
B2dr3Qc49pHB+dFzEWTkIWX2Fz3kF/o/YM4dwVy781OdNAC0y947tvek6vcf37HpnMw/BaB/EkWt
wkEg9ZcJxcL5Gd4sQilROFqhGTDL1V53VswSla1tTxE+S9nz51GMzVKJQ4P6yma1RWG4SBiK+wkP
Mi1BmduhN0QxB64NNjDZFjresqvrJGeicI+hlN5ExeeQAZTLgFkHERzjSbmUhqEXndPrXWtUZRDg
6ybfrpAVeut2ZC6PZzyQQpbCiteuPmreo7ul+gHq84QoAu2qaF9baJ6jJOJxzgZcAIUQgqm7EeQT
3KrIQeAea0WHmCoJ/1C8caDHMhaHCs9/8Scd4/2IIMLPXfZC4kMTbWm9WdwqE3L8jzC8rW3hJUKQ
fMkdY7cMLlhKGnnM4qQ3HQJjg+if5ZOjAxgmt4LY4J7HC9isIi/166Sf2q87eZ/FgLgUAqW2P162
LpwUXPBMIg+HwsQkXQrn+J2urnMparsukZ1t7n0HLarL9JNsSPB1R4hQOrX6CQA/WQWxr5ZjTdK/
wIWBJ99NjQkfIh0q2jeft57qD6ICD3rXAB4cJHs8WF+XIYYQgsGhrqnReUIEXfIBEuixNhQrXj0G
h73KzNNZhjKwa6LR5ExpwX3uu/5f8oY9QErehtO1H/BHr/RAAFHJncc8C0fZkrr1hhyJdkJOwBYH
8BT+0bz4Q/fYAyy3rEq8+OBEGox2C2EAq1pZSI1sJMekxpNGAMIPI2vBBGXzJposw4SXmEkKaTHL
wVIvciCs6W4KIY7uUMlxu+PZYV6YsXth2hNC1sFIKaNxQ8/QqTFQJsLRAXh/eUcQOVrjocOoJIfL
AIKiSICim6QS2Bb7AzaaMBX9tga9HhnsCuvSN2nskNlV8KSn1iEHvrrouocLGCj6qaIRG/BkLj18
NqSlmvwj6h9Heay/J+RQai++FuuBfUy3BR5y3lau154gzYCYZ2ES3/uEIhnG+JYcEt4c+OFKCUzh
RnqFhbEx+D8EsArdRxvAaVaQER980BT6Msd67T8vFnl10frYe7ekq1Vb044yegT68P+XhVRJoGVM
4WpflV/gfVv+U8HhK+E/pPKN/8nbTrSTD7hrMTbd3RTCAryswYzU1G0pedZt7KFnxS8kiutMlGhC
NHlheIK/SuBEddKWB0jozzum2ervlJO+LiMSeinyWFugoI6e+Lu72H1iWxh/hBzXSLcgvHawyNxX
/OCecox5/Y+32trcb/BLcMzBWlxeeC+8r0/Y9A3SXn3NZAIxQH87Ws+hC9war5Vdq4lFibuMeTA7
VE8TvjB7HFx3xijok1voNJFckM5BLTe+2crSgNRtw6NTbJfT6QRRychDwUGMdd2Ja7Kmp45HmwH4
hUqgVE+x97JSi/AFzkFnAePa2gAwV2adhT2CWpSc1lOejKQEcus0IDQBw08IuHiGDlJ7oY3Fc/gg
5Qp1kTmJn69UkrLZvffPg6WIYTjK+B1pVVt6deVWt0YTT9ttI8cO6ozuQPSh4hW7caFtnxcJPPaW
rTb6LfHgwFwsX8s2q5ZF0ySNb6fRmu/9cR5uscd8f2XaNPgdYJD0IiWhnQwUtrX2TV37sOr6OgwA
PxWvq3jTvFMKsJ6KB/rdjPurqjqT3RjTp2jAh7NmIMvtMlGVubVPMcrKcNork04NTanG8IhJsFvE
4RzjkmQLiJuDw/Cawsq5naUhBI/Ds9QGHz46yI8ZmAVIKBdw9AE6SYgfOCd9D/XgLkpoc0R7rYCf
txotmYCcMPaILMH3IfAm6WD6iOBSsaWwLq6nu3I9bIc+z4nA/+WPdO6a0rD/123hYOGS4CebpJNY
aGguC0312qj+Vg40+5DgGu6nkZOes4j/TBQqdfeG7yLX/lj/rfQY3n0fc6dMvR9jyZFWjHuz2bVT
xl/CMvXWMGhScEiCvgKJjrzMLOoE/42WFmSUd7WBIhyKlrVKQmT4uuyXuoLgBNuYxrOIrM44RXvS
VxMxf/O9cguMctZnjyDqnGrWc/LhnI2TjZ9gpM1SZhSZwficVDFBgiyyKuiGh8S/pOFWhVVvplDi
kKzNiLJQR+2C2/iGWOpKKhvKZhYJZMtcw4m4ZznRyHODqgGu9r1BvjYkEYGWEOaViQCgUeDqwwyb
wNBD9/wr5r+BZajGKH16AgBK2WfBQ5sDLbjVa050VBP2QbtayohhW3nQ+4BlV8J/YUKn38MMBlhT
XSpAOjnqEcDIJsbEgvBBnfzi2TR4zYjmCH6BUO1uM6qlBnxoixU8lzfh7CXHXBRzvmAmA6OE9RHP
oQxVQoM4ZQuykYRuxcAVp4Bm0fv+ed9ojM/OZ1bzewaOspqe+mpI8NAV5jk/KylhxEWTRh36EFEv
RizK1eHxxZ8QgCTDM4lz2SrWn7w6e4nIv0riJhfFyDToQEcvWCIeSwzte9narb6s3F364Sa5Q2zf
T6m4//3TnbukNaR7bLEzdg2wLuFC6+eYdfK4fq8Ol/FmRX42cklWa/m+9xz8qbqar2Z6j2m2wYtZ
tOBa5G9TYE9Ydk/Lngy2BSzY0QneJ1cqGZau8PCHHyM7xgEBYpgBGrKf4W7SH5+OeDgxGlpElusZ
2YOxS3CPklcTFa4ae6raSihx98KoKNcIzaU8aT2n0c7se7hQGUPXuoP/kCyl9dEuTMGUUBQYH7yP
fHG0Eyg+L2t7iZTRvRvDctHUs3ZOaeMw4P/WP+94H5+0PeFlxsl81m4Adh6nhcAcOW2WLYhChbEf
88jfj59nq5XrRajnn+SAkfLoxKmB/BaZ+fAAtyzVLlaBUwez0U+vsZAhy3PuTGQJJtPYnQlyCkVo
UHWwUU9tv98ogJzNs/7o52JBFc4HrXJB+KHb6sU8F3nnR1kYVZOvuEWQcxvZu8Vm9XUfiUydyMmh
tB+vhwxJCMWVPxnuf7e5XUafy7LlQMe1HglXrq/asbh1CaFgRxK+hPcTZKpTkCG0uAeRGs4YwcfC
iPUMlQnMq2CJfuX8RXqpJNFGPTbP71XIqKfSLk7S638bjUAXVdFhjphKswV0F0tye1r67iKMxDeo
a+qA5BNEpCmzecCMynzA3Xy6lwhOIoeRUwsWWrN0iZ7AUeyfh9AvM9xm9cqZ7gKM8i2mWHJTO3CP
hQlyyH/i2DiAO0+0LMZ8YpGSpWjqdWZF4gJBXlKfxz39GftxWx6p7dmhj5Ay3NjFIdpGIEs8eqhJ
rOxe/ty0zC1XLiHvQ/W0Md7tfKG2mH0ZG+Pr3ZsyDwLXeQfLmbfSY75XHkHOevHfh2FCLe8GAdMD
0a99vytK8pVl54U79RWuybmh220eddqsPX9Sir9fMEkf7J75smnSmxapJ14kdFc7i4EezyPpLy+7
oGl3ZdD5tLlGO5y7IJzNrZDMBW3xqAKQLnt+asQlBDlLJBmsjO618Fu+SAG6CLgAuJEBjrNzcWrs
H272tC5WKR65i1o8iTTW6VQLT1nYt6X21lJFTgPIBSYJtQUHfyQOqfCtPkl3v7FM6LjRiDugLolL
5zt9bQGlT5DvA3uJ9sF9bZ46IfWXYS6/5JZqk6LZGEXg6pV9i5HeoJGsbiUc2jHNfuves8K5FMZt
Y4cdKeP7EwRvPbqQMMA1+ocj9kejjr2KRM9uIKROr6/zjIk64HiyCbhhcfIWhMmo9HReYeynqhYo
sABDeqtuLbxBvHTPL04qtwQtgrxxYAH9vRLps7iczvmPgOgfug968P1yXu3sYeouR8sj1t819CAn
8GESigV6fajgye+R7dV+bSNMbxdfzmpmTaA6ED3LANhVpzlBNMTodajCmUpJOIpjAW/+Kg/YY/jh
c6g+RefFwnhZnWIuc+6s/mmWM1Inlttxjj1KUbJuclkeYOGGsDAR+6prbuVsQgkBaNcnrdP3Fvtl
RbngA5NtxP16ANBnxzhU2tL2oh7G9/g9XBGx26qWtyr+qmukVUAaS7pLKlw7kIYdtnIVAa7LP2qJ
hAZCYuUJZP8s3ew+AZVM+O2BCB63cGDcaLw1dQT9lscWWd46ToJCdZEy8YmihLrJJ5PSsjSPijHe
oBqooJGHta3PPGSVzrJMuaPkNLYp/tJWHnOZBjGuUD+jOsrgsuZAsX6xFr74IHXwsJT8DLhIv9xP
p/p2NQo4WMnMuk4/HA+/dJo5jpyg5fOK/e58gfIZfpiLi5Wmu8RQP9Ucavckx/OOCUbZHsVnk4yc
bIouA0VmKJUmUcmh8SwqgUIm7/knIc3fgittcPrtMfYHpbv++ipBJECphAkDRNmOAbvkTAI1dvc+
s2szb1tcPrz/COHQAJUpst/0L1iqq3IdSPVe4DuQjd4nhnkno3GgWrGdVQ1iONVtgYlyTKlqjkFQ
X8FOmmHGHBM+2u6NgmJRB0z70xRSWm1jTIQrIiA4y2dOKUtY+u5ey5Cx4uXpW6kf83lnftcRCNOA
2AGs53tmt+AUyoUJYMm6z/BBtimE+DxK3j9T84JvuSAOdnBA4PJFR6qyww1CeirYKFh4Sydxq8Xe
y7cEVkFjQ8aU7wqU5Padn+JmXABm6uNW6u6rj4BwpjANDvUhghT14YB8UGRK8lx1sLZzhaUZ8wbB
vjx1DeNqyhNsxQ0D2QZoXC/MTlKCvckC6yYarXHPyf5Sj3hsPRXpgQPiAUq2a+tscN9iWGMGtNu+
x9pXDGlScHhsm3x8iKL76HUngBisv2FpHdp68dScSfMLEmBw2H8/yiQ7EZLWxAFJXl/+fQXgWeY3
dMqrWDHc7KK71q3Onv5F3smw55IH5u3hTgx5VRlFPtHkgDBykuwHztJXR42bG5xkUC21gsfKVDD0
WBrsqx0HJYyINK/iRV5F+aKzaKpNScnZaP/MmKH9r7NF8h6E3ksmOTosQiFX4s2+PFaU8vrELGfH
dGXB2J90XqH/n/x1TzeXlH4iPdhK0SIVAmxIjxQlw9QJI4HcM6/kZ6HGMLYrGJmNUw9XTzk17ReG
/PsKHmrVYg1wU96qBIqU3sEf7yEB4LpdYUVncxBmwn74eMs61bY5I9rk46faSUZWwOhX5q+Sze+Y
yx0kgVI7y3TAEybJxl0FNVo3xGKPFdK+vMQyjPxnY9xxPvT0UPnMf9dX7+mToWC0heB8h9fH0a+x
EDgD6O/RPeOeOl7oSe5ci1yPIk+EDnbBNi585RMxeD8nzIwULrQgZngNQ7Ko/WnLl95lEvwJQfuX
g0nWxJ41gLxfda6VUonNpJefqPSlJA71CPJtSealk65RtQABSNcQOUJv1VBt230j2jm/ThsRHwD1
STALzxY/LrMwFavMqDWWrmoyyXxmy+OzC7bW0IcsHkkZDZytFbsm4n9OLdTTbsE7s8S9kLkwck42
SNUsPGZMmlmj9Als5DVaArpm7HGXLR47tO+9/oQiFlt9vRFfr/ZCIolXIZlQbV5FdnGI/A4FpNsO
+gOvAev5yfWw9IHl+5jGonxZPw5L71nkz9cl8YMON6huGz0toy4W5BoEgxdfXXy4cH1GVILVz0BB
GLbj3QLjaBunpikX0E0rFUWFWBgE5P8spC0fcQvzpmuR2nuydiQi2bprJQ4GF2ex8lAyco23xT23
H0ATW4bEUWKy3g1T3LROzqprIMTMRU6gJ2Cgl2ZBzV0MLpcmGaYxT+ONBfa7E2VX21XOb94R1SsF
c+d6uufqeGF1r9O2gxnG78OxPSR3teLwNwzoy80TlbgXNgYFk1QfMUv5XdW/a4yMnNXCCmruiF3p
Gx4wafws12QlJ7fpTq21kaHpEzoYOMuAJRi8N80ZLYG1Qjc3FB6VCgwPaa2alORqugazisF9wLM4
BxPEM/yWA4vTRHCKvjCy71jgL9CqjzSEBthBEBGaTjYitxISFRgwmSFxl1My4i5Yh8SwOQIvx8UR
UT+1e1wd3rPa5RNBHF89D/NCyqlN4xsGX8anl5CmlTpcnneUg8ThnHWcS6GID1nCRRFtzI3wHJJm
N6pUlNevYP2nkyVl4FYllgSmwqMHdP7VVY8OSJp04Fhy/EUzrCabgv56l0HtJ+YH7pdE27b38KeP
Nvm1ssNtGxsLQyaFoKRMXJKPMNtoWSoEo9lIFTJ0W51FMjuQyaYWmdQO1Fwn4ReJmqqMHuo4U2nW
imN2mbfYBJ58YDyr5oe9tfXgqUE7SyycwjysJ5GJOmsougGH96fnlXcaOXEjcYc6yepBe5byXFFJ
43lUI9SDDCV4NDLIIX56em+7lkUkbMBtP7m8PmIW2zS69f45sF6NkX9GsYCFBywhDFAhKhkOnqKa
U7/MIaAT+xtF00Ya5I+ao2Qa50I2+kfca1/Jvsfjia8RHtS/C/8JDTI7rFrMznwceJia+Hxe/KY3
ibim6LwESSILFZl+rKTSxhjBG1zSJ4IeTc9IpnnR3VRTHAqq3cpjs9gNmO2ZiZdZP05zCn5yEGEw
EOzwEDrL5gYbC4HluiQf0syvdrAKg0PvOMpz2u0NZiNYhINVgVQqmn1Acw7BT9bXzVaQyge2N6MK
6Z9uUerrw1s9LHkyI9t20jq9lbCvcok5V01WdZZ8wph/l1mCmAHy8uF47m4wddl5m/++V5u2CLlw
ikJBJhiUsdMMq17ouwZjEfBab/l5DEJCHDlRxxOtOJTn4UMSFIpmyRLBS7HeN87wp9TY6yQaIHuo
bmfy0uj+5If+S2X7zznqpTUHWis8lHghxCQXyUXA9OJueGjDj7rhDhlJLMpgtdPHTfF50pQfE8w0
F4vqPAFZaab3jkhY1fFabecZqMYkvMA/Y6Mv8ZGTq0/wbHcRdikpj3tg8dLZo3evMlOur6pTG5TD
m2ETEsET0BxPeJqmByUqeUCWh7PKMYskWnBCPHHSivPYe2Xg+Gx9bmTmXZLZgq70wmegpW0UexZa
3EnDjENLUKnDzbqdzaLBhqqf58pRLFkZlY2TY67yonddd7WLoOTa8fSaZgSZsRW1bT+P5gW4tN2p
PYcGVA09rB0RgctZG73WWPO/pM0AvXO+H81AaTeOBDRt9FQR/8QkDjLbT2T3AeNUoF+kWvC+eQbc
tbov80XU+Gntbl0b6SP4aGUsMB9QVIMKQmLa+TZVXVenO4fWCOSsp/o68Ngye2uAithMDM+p0Ccw
hTftdbdOzo76vdrNA5084pYe7y7l7ccoNjlPT5MusUPondlmC7U09BrjJX4RBLtLn7ztsSxgyGR7
xfp0O0C26U4sW7ylhOC9IXZkyMb2R6nlKijBMFN98thrFP75MIVAXD8Fw1DUHweiKqJAozufcADg
E6IcZ5AIAWCEZ+hYh9siAILXby5nXKxqPdnIVdTHYoar8gMoboGf+xpZDjj29KYmhZUKAAMvFra4
dwfNtqgEgtgTh6FtfY8DCDdnpB/+xK+7aeXPw3lgkkhsIf7yj0ZitxMiih5m0FyGsOPnyUCuzzKu
bX+dJR6lx36iFMVuNpMltTU4bWPSbl8K88iMEr2Ypw+yJc3lhEEzr74EAUEMP4Wfd2IZzsVvWAj6
1p7+AY66lEaME6VFYapycQyGrBFP+AczvaPmmTM4fOLF31HF/JwY1MWhfqcc6+tmwCnPe7AJr4lf
dbrNC73NzYcytqXCR33xLXE1Rv6HQCgrGQhQRJY1KeQeLMXtgCpOXT2xoaKAst0MJGQImaaxI0NK
KSiWSHqh7VRkbAMMnskT7JhZpAd7tprGxQtJKKZ1ylng6hdC84jCLS4Ffie0bmurYROpU79343rb
sAptcrVf/8knAwh0Pyjq5BrygOxO13Sy/WzcPdoLXCWRwoSiWwM66QEBEP7EW7p33jcRCEI8n/iM
I9n22s08gXrbeG1myeKIWa7IkuHeKyQ7ZjuzffCMnZdzMcRvTCfRM4SNjSu9o9x8vhiN9ZxJVA6q
RWEAM/IaTv5U1/97DL7S3mK3pIGX1JvthcGYWXOCoknoTt6mVJzCxhsURD44WrNgKXINyVzwz/z5
6R9Ft3QFEOTRBpaXmt3WZ9VHKIgcqyGM0UN+fsYWzdmVBg8swXo+k/pvChojvUFbDmjHUjOnqtlp
Od5QZwcDN/Sw8o4lt4b3jrOcJE4773shiTI6f7HU/YfBmogTIALoR/alzw2ssq15a9vfUY73eSMt
IWtSgUYUN/JI61ZxoVpJr5Suddq37l49DR4QC8wte2jZxnDGkkEqFAnVqFeUNZPkJwBV3ky05e1V
82TmQ1XNyV3nyuvnXGVPLMvhsZqGg59lAdRUzjygGW0rDg4J2zoNUni9BKy38DrSRSd0jGmWbhgO
/PmHxznYxPtUQmLfXKZH2jm3Rq7bI3gdgcoG9qgse1PGhNKGsIxwFMsQFKZyo1waaEOQmcaFYvjE
M6ZHW4jP7OgB6MKHXfv61b06m9fAUy9bW+KFWe2oyoCKK4YLaSVFeaxc4pXC0J6o2HPAFrPLGJsF
yttU0auq25Vf6y/+aw5xJ6ZxI0vOvgpl49BJMUTBuj2I8XJAiK74urC5MHu1H+KA0nJk9PPyVHhd
6j/+h+ec2OWKC2AcFIk56pviixN6vtObGR1ui0SxGnBcd2dWDHKoMv3ikrqh7GyhzYIIlBnMTzKs
Vd9Vf11x9lG8symvGvdesx9pm/73cNsVeUFHtVB7jTX0zKKudTP+MjdHePaFA6l8mfYL0QEg1jCV
qDbegBB2h6EDGszu41AaB/2vC/o5S/enLKYL4zdHUVCKFroIxSAb6G0V9+eMA8cexGZkUXgcnrlA
S24i00kTTanpE7+W1jhLchv196JSsDxFTTw5sgz1kc42oaEtcNmyBUZpKHaINy8SQinWd+CcJk4X
cj520kkdkYlv6EXNwbvTbfwD7BazCFINey+r52XM0hhwLlEItNPvCuVJxqWtqjyivrp6XlcYITit
86Rvkj/br1lbd5J6c9qRb/SZlzds9XTKrClMRHplEqXGGg4zTD1UXjNRxmA6MNt/v4B5hycQjJO7
LWnDFTO2CGEf8w/AxHf3zB+mgblo/pUZkUWBfiDyk3S6Lk/dmo6GpUgQqkEePBzRPjxO22bixEPN
I7gq9AxJ14PZSumMEcKCpVQpRyHZvDro/R2WWD0vPHgPrePZMkNORKwwm0b6/i83UGCC0rkhYCMV
P+GisBSstn0pNbfYekndrPydU0PoQnTpe2myqekUFoxJLOaxCGGdruSIeAD1Eg0x3J+l4+B/I2VG
1gHFVtPc23Io0aLPK8vrtd1BhswN29Jnz1TAlZ0tRqxFEygvXhcRGfEf1TGIAIcO5hlDgMjbbqz7
LZiRKw5RLPdG7YKsg+SSFLk+3GYCGDfD5kmEWqiMkKKywGCxuVMl3ZmNQxTzDcdbLATRdZECgTC0
SDhq1dT4dUlY0lJeQYFc4QBfzceyhNlQ0TdWA719zRxmiQo5lO35r61rskfO81yWmcL916rRclc9
+rA0ST9rULGf0KFwm538ZVQd/G3tL13elNeBW6XdoJec5cgvMtnCb6GQRkuDlKAsj/UEhsvUwWVW
XHtHr0L1BsfdceCOOE58SYaryr2xE9J7Rdvwxvpj8trtXX+M6FjvOc6RJBL21RhlS3gP8g8Lh1FC
BQsYnYmepdqxRj7+6wcNtkU7k8h0fKFTQb72ngmdlwlvJ4DZNvR3nV9yCBBj15q2OnbZmOMx0ETh
ecDOOtS9ELE1j4Zr+H20FY5DJcly03Yx6tc/OpyGiIGpWvtXb5fcILKP293e4x9zyVR5abW/4h7m
4RLSW4HAjjIqYMM17Z9sXU1R2dcwmRPUoB/PBK8/vT+s+UaPtKEyR+Sta7mxRoqTO0FZb/nhJuMF
xGXyN9TeI2HA7H6i8796I4N5DzZ895lU1k+AV7JT06hnr9Gn2LtCDqwBwviWewULkultqyMMNqJ5
npAldRCS5uvLsX84z7S3fdVR6bGndOvpAD7OCwhamsVDau1A9XnhWjbRNvFEo/RmJiDZH9VTyWLH
ag5ZyV14RPdXQkSgmsFkgeXUG0ahVwgHughZSVKJOhkT52XkW++9XAHfC4KcevyVDgvkoCAix/oZ
+50cimqE2l4eo7MoopUg8F9kS95Ed5uOG7sE03JgOM45YhRMe/mM4tRP0QONzRfHW4MzGS7nDLIC
js4W1PpF7T0dUMVnWnnxok/AMqtuBuor5jxsgyEddxvkA+ODwdgACByF1NPZENEpdSCpJgJVFG4v
uAtwEsy6LMPa0MHbBfpWAeAgrM/hIznd4gfN4wPf33er9mEn9TMwfWLmiZkT7Ow+i33I00LZcqPS
2/6YYz8dr1wGSmAQmjZ3dPXse7D38DR8nWGjEzkMA0hzhlnMXc/fDvR8KN+SUurlERmLrUTgRDEc
262JKuloaZgpmabYLTTDbHqXObK48fdv/jEJcQNF0tgXzPIyEXPCBNOoUfhyTdc6B2JZxVwwS7ig
x2qEvOkILbJnioGsPKCe8uO9NMu+9fpJEIrOOWzKDPgGHCkWGKTQAupeSxZsbDw6K5wbcdTgjJIk
TfG8BnQinxQ5ne1a6YsMoUq1jvD61IQ+95BelWlC0crb4NAWDeNTMjGNlTk7OJp6b9+N0AZDnYIx
W/Q/YTt0XDaLjFSIq/aGSANHSS2qnIeg8SwusVSkG6MjBQyEdOfpHvI5WmT2O01AsJElmfux+NDd
UQfSrMzDd2SgZq29QANZ9a02OBbgQuWzq4qcksp15tjazWDVGXSaHCXFgTbqWszK14r+NpMPUsFX
pWLpbiInn7c+YBcl1APc3wd1/NWsLZHRSr3GR7PKV+AN8zRg1eDwYomkl+M7wuj0swHTLzTPt4XY
46vrU7Uwqnhzprj1WlkSfc5hWv0ftVStdgC1i/nlcGsaCPbrzahaOrd4iNu6IdMEX2Hbt8fjvDER
hS9gIbYLAtBm9yJinHP/sQIxreVfH/EXC89shCAtiOGuzoBYFuxG1EJmjtyCoHzjoAOKE2QZPW1i
pXMZz3Z33QwG0Lkvp3rXupvD7J7SS89yXuO+SwOlO0QpVb4bChuLle3GNP1xeqJ3ZTInGBtWt++q
0q2YK+z0EdVil0rri3XT4zj6jdni1ubfswKvy3PIMUDFnYUtCY3BGyLv+SZt1dD3cCx6/0/rnkq/
3WoTsLYDWVc0SqDyHJEjFr31QWiMmQ4p8PMjb6G2RacseNKlc7y3f/UBMRTxeHC/oPsmy/7cU/wK
c7UVOUOWoKIG9dKKB0j/4CA6Jvi5DG5wXDMljDdBo7vKg/jr8mRjplWt65FSUyX01ZKjUzpy7v5S
hlKPWztpciD7rwnU5IiNfKyTFtSMRESgZlvIj5k+/Y2wBhvKzw/a1zmMCuzs9H+r/1evFegUYoBv
1LBUQuyrSYPlH1NfJK0rAY/HTVs73k574zm9Db4XmMizBd9uG+fm8KU/VDMEypkDi6RkqXNN4Kfn
qwZ0+5cYmCq7VUtQ/7MamQtxgqE3bfZ1wmaQmGy65g3//vYmBrWc0UMPt9aeKAAfHWNTWg5yA8zq
Pw/kIrOns7cWRPXoO5Ta6IqO9UGmHuazGl7pn0x2lRV1P2BHvZ4X0XxrHnpS/ln2il40ixOtuzOz
QxK3D/FNhBejb9c4bccl1RFzUpn2/ODtYqxU5yFsxeRls0zTj4D08+0P/k3H7QsbLAYZ7Y3gIqgX
CkazpD4SAsLukxkBa4EdASeMENbyiRD/WfUcL8JR81QU6v+oTCejhiP4aqXo9SquiKc3fzXn5/R3
AJ0FXXWCyvafgpRSF7ccRj2b+G4PMFHjsXUPhjPgTEU3eJG0zOHpKi0fpvJ5EpgR8UyZUDMj2G8I
hw61g26ZAeDSMXnFtbfytVr42NJT7WLvFHI9diwTsyTf5hsByznTsErMYBiUv0w/6jVnNJpwrBfp
Ez9669kfvw0TV4REsd9Jgw+8L+mIm8PyjzFPvg0xA7kK9rCoZrjXgKlhdcU3TqWE3Ln/c3YchvcP
HeblQhgzPqTvU2EjYc9dXVK1/Eh8lUv0qRCGkoc0BmzbpM8N4SDmcU3913iRK5bPtWwTrWG8W0uk
nmej0h14vfbdFZDJD2YXslr0CVhzf/o85KRDdHRqpqbPYNpr+8OFU169mU2n7kqqxqRVTpD+3ewa
zxrJ2RuX5lLrJV9rsjLRdi7jVBvMojlWkNobZ07Xml0KxVebevDUbib1kzfkrrg1i1FCu0yG4ODE
VXDve5sGvhFx6PEntpQkM5K5MlKYiQxXtME7L3Nn96t/RbpeCs5VCkYGBcZs/ZIatxCblRSQw+jm
pCJ+80P+E8Oab1rzjnFAXVRJQ+9zQ9yEm5d54InY9L609KLyDEVO36dsxqCBcK4z3Fv3CYbhqJJd
n/3R8cPi/KlXksUyqk00aOIZ5pR6pCCVjkzdWN/7dfWXbA1G30EskrwsgiqLG9lex+RlgV14W7/i
azPYOkEsdKPZ+7754uKEdXVzUw6yZtuC29ACUb3jHf1j2f2C43utASdqqA+sHrrFrNx/QalZb1zN
H7iGuuYq7fVIJCPvqfoGkA37RNBDtmfaFvoLd2lJjuBUVjJKxP5K5YogLGt3+PR9EWrurriNHgCo
EKez++6J6iuQXflDsobeNRshlaNLMB9ZRKBPWgmcOcRoZMu4OFnrIAMkC3OG5AiHItmZTwpaHY/m
g/OJ4zbOSxt+qu7G1mPqbjA+VCUmDNvgtgJmqdjCcafZH8XqBLVC4sopxKoa4g0ngmSzSBZMLo0v
06LwXmyWD9y7T0Ntj5svZOKuKzHWqH8GfXQW+mmzfcGI1oNbP7d5C9YIsGWzNnHnxwxpSx5nWW/m
ubGQ1waPJe0u/afrkSq/0n1LwaVNuZhU1HxaYmV2rkDklJRg31xdD1qQff0QRCrbima3QD4AfPPC
YLeQ2HRVVjUNGTsr6kLiatYWUGCEBjOrDAKrZeRAaiGnY1e5D4j2Oh+hdx3cnwGi/txbYrSeJUvt
nCePru4wANDY/xJi3DTFDDjvVwGp9AGbuHwfj2ixgWT8rVNQf+t6mqIQgY1Yn9QUtkZAYy4/bYQo
K3fH5NEDZCnVJy+ldZ/u4p4pLNEypc32VOrgQj5hpdJ4IYt6Rv0gKAuwZ0YXRSgecEXcAXAltTEA
rPzbulqsl5fm6YCzRaSECwXQY3tt2BWBrO7jLHUVW6OKtB+ITK/I1QL7KNCUTiwoin9OBrdgb2rM
fbBx9Ka+oGvJ7c6eA5HZHFLTgc3oMZqgkCTuoHmWZwhb5jJ4nS8aZ0oHHAK2iBzXx3w+xbw0HsWs
nQdiE0BR50OdS4TCohvz8/8f+5gdZaueeQ55OJumFkXs7r81mqYIFTrAM5LXrElXmLuBbW4RPTiW
RqrLd+fRjoODLaN3jnl7SdMm4cMXN4O0F5L1ix1zZFZ5T456b92c711X/Yr29ogovofDNGNjhhx+
eQeqWq9HQ3sS72Aq0szlXk2iM+hCM/NCnF7OcD1rk3/NaKiyySG+lqZE8B++37pvgXNnriiJlAwE
QYung3VnCS5Ppo1cmMOVP/Nv5z/JJLvDQccDyObmUmF94soJdLhCqondaXHz9Ssr5ZkHdKeGlAAF
UL2HUeRBEDsoDVm2PvCclctG9IGl4NtDfEMeK0Pj6m9pym6FXy02qjS+p0kabSFUsDxB0+Usrh18
sK7av7vqmQt+6ufZSLIQfZJEb/q2/PmTIO1b9YpdbhRKddtIgM+rL8HemsGrTpEj++QZ5WMv3/ix
FE1Ij4yF1SdJt2E0SrXrOkCdNFjLcLA8Py9ODD5L0tu1HcevcvnJ/3uBX/Ws6A/XYxUnuVJwVS8P
gj/N/HHtZVFom6j29OykxKf2oOZ/eqlhTskw22xpXVlKjErx75Jv39qsFfGPN/iAU+XBUBsZA8pz
FSW4A+w0MINsQKsKz/xz6Iu6zZNbYD29/CXpaPUUm8eMzrQw98iiR+ftc9oCxs9Nb10AoyVZyvmu
L0uwj0DM5oSiL7RjSIN4TnVt7RohCp4E9+wOQ2sM9weUQM0ue4toUE988K6NBmr3FD2QdEGTzCNF
wHBka71FqPkISY2+eLyWaswLiHklGswx89mdtw80BuxSuDeR0Hor7deMMTu4F9K774DW4EdNBL/U
pn9btVfCd3Hjs6za/LYBbM66Ohmi8E54PRs/creeSPtF2LuVj72H4zDH3Jr/zoSd2v5uWAyvU9IL
hRbGVwlQVgv4HdokMThScLmApFw27c8dFC9RM81c7dBfavKayTJ2PCnEHwLr3Yff7n8fyxlOOu2B
14tVj4Pc61d9iMEO4Swz49KOPhhhwjcxgX+tfcQZvoOYWoZKnrhuHRUCvu3rQNQQEoL2+h/Dji1k
niyYTiTnzIrCuO6YUElVztrwG9BsslA2D7LhUE9Gua6hwNYDqOfiHxVC7PxuTzIosDnyPlBHzd4P
OXexJQPgmKGDEG+HWDwuSoIVa1ok/B4Ob7b8otetcJ9V8+4jAUTCXfmcUIUv/AQ8XpwTyayL5eYJ
6uSPOr5W6tn7i39M70PIlYAs8uD9eHmSJXYfUlcR5jmiAddbFTYKkkj9wMRJErKaQPSHzvSrSt3C
Hmu4M8PWLw73kxehumB9ARcBwizipKeVopYMPYJff3bD9ToTeXwL6Mx8xPTeHVjFILP3DzR3uE04
VDIKnA4VNmKt3DqEgjGtVHXQIqpOPi6JJC6Ek9ijqYyXGDiwE8l/B7GJkvMYLyNCOceCCxM2ZQ8m
rUUdCfkpYy7FavGgPu6OBYG+UXZSVZagSDszlJkQ4gOVS2CVamvfA4wDIfKxJQC92AdrGQV3RNIM
wKyJJrCBA/M1BU9sDa+KB7LF8KiZuJcuCOzepSfldldi92JAGKPw/NVUbSGEFQFz+/Yd3Tcj8yUb
aOhJ/ro0boXqOrF18MS8VdZt3M6ch6M2gI/fhezAI58qA2fAwTHwShf9r8DWF3JnbeY1kT6FXU4G
sdZxWVmvBPo2Ks3qHtk2PsQu8N3Ov5r9eJJbLE9kw4CsePMQb5l32zgV0QFve+f4+a1O/NNVpyg7
NfTxDbAaBeBiPWkXpEkAwkhBQCSqZcgZk8bLZfaA/45JuWwMHTb+N6Lz2jDmqg3vVRo+v+An+3J8
uVIc+76E++p+UcRdv3+YEx28GjggADwZVG1LZAZkt2y5eLzCS1+/q+mg2aCxIr921Sgy+fiF5hxB
4UjRTrJVv7sSerNNiC3AjFfr6/siLzLmdJglWQe2bKk1Vcf3hZGNeHdGXnJhCicTD4sWeboXgkCq
wO28ym+QKeRm1snZFujQmpzfSEtwjT13LRVPYmjfc0YJ7oErRgx+OSFZV/LB+92wiWO4Cr+yexTP
lVhloCY222/7qgNl6pf+uHlUU2RBeqyOJ9BNGHwqoe3KcphZCaj8hsl8artVMJSNANpDz7ic3+JY
/STphpnhgY4MIzFXi/nRDANFAYxM58QkrWFZf4+7nc1W4KDEWb49FexonAUNZwQHgmMDhPzftDH5
idxbeByX3wRbzV7Ty3dh7AXqmrF5tQ5o+b2oPqj0siRZj3B+XQtV5eKC2z6inttakqjYGlt2+DmV
HLYWBGxaUmMTtK2FDjQE0i/DwDt+gNC1DQ2FAqirmxprioQARATq9pnB7Wikl6+DWdJDQ8a5PtqT
vAOIcTQ3xKXXtIga/sIrtMn0M1itiMOFq9lbd8S7QecI//C87XUwzRUwsvB0frsx8+C2oEHsQW/e
+BF+XLx7pKATU2LGN9RkV6GCLeBWVlQi5X5GR+CkvbZx412TUigJj92vTuoaKtrbRI1tC73ouGjr
SOC9UxT5Z0PnGpx9Cxjwz00+I1wl6KlktLJe+uPLc2pYZik+kywscXWXZ5tMOjM2aold3SlhF+p8
R8sVHg+kIFfPMUyb8aaoLc3IILj/7+7qIQMgmcgF6vXjUY+iDXu3t0KxE9hReP2L4ILCgu/AIIgc
VEnXVUtksMV2meSOsfXV2ImLRyC3vo9pqwi7xcMekYXSQUnPhSBRe5YpUsLUk7XL6dpVAxRs/IkP
fUwwXy6LabnFAxSxAhPPsX8eqfNIzDXdh+IgIc/cG+/zBLYOgX4tcFjwF7P78IDEruX8Qxoy5Dqv
XS5UOQF0+PgwZ/tjDmOOwHX3baJ1q3c7DXiwUNQHmoivJPSHPVKWnUIHoIXZNVN9YOl5DfBd+g6H
TtZX6ThtsukKrqjhGYv7PfqpugAp44SB+gInwZfBYwaGJ+rKIiteXPmi/xh+eak8ULqaqjkMXkuq
TLd8JLzyrvHs49lNesnPLwI+rvfDs+QiZaxHjGDwtHEO5YcOsavFd/wG9AY++yHk98x6AbCR4deU
obUdhG/6i7HUWPAavwcyBUqwjgef4MJFbePi0T3dJSeRhFRY5uwio5+lYcQC2ytVWJL6+xC3kA+W
vKumk2qDJwmo+hGXaGpQ4BWStFcvktqqP4A30jKPiEs5/64jvV5x7Cl98QXypfNkt7RkqjzQn/QF
857b5n1JBBuzSjc/SRXS8rwSKBsPJ6gsPgjaDZ6/gIYchOVjqm9ul96M2lg0V1Duz4VElbXsLeSh
fTI5gUY9+rx5qM2vvsVYB9C8ZN6gilnLC5nlw0jKzWIJLi7RJL6WtNKlQzvNej/eXRl8cscmBRej
gVJOuddu2Id0lPnA1D1sd70NfZs1azJlnyYU6Rke4b51UQa3za12hlivQVFL5sBxFnXVar9ZWIao
up5kuw35sDmRrL6cGWnOixhIcAw+KU1HEL1GL8XPH9HgkZdlBD4xxGG+pFwYb1QIFiHgBNqzAZX7
h9jZ4894KNoC08LU7ziLFrSzzkVeHZMmvnrXyAP2h3TEvjjdxk6FLo1XoPRALJOX4mlwr78ShOPB
c/XWKJrSGFjyGT65t/iGd7mth8204dGcqHUBUcJB4UqTHMOrRLR3u8ysTWcUDbgqOllyobm96Gc3
kd7AsEKrlLsNq8lKhXamu/40x6bRuIeAHBiArN0dm6HgeZLsCoViuE++bbMhrBt9lwn7W/SKt9k4
ynsJy6TbpClUY5EsneWDI8rbYMrWZlJhnbxQIk6qAU5WKr3/ZUoSzo+26Tyx9Q1rAnR3WOOcP27d
lCZAsoMObiqvPvW4vOQb1SMJgWZiFENR6xqmKwKQt0oTJExrU5ik7FuQh569tF+r8YwimRGqzVNE
m7vJDvKOEBJ68plwHvyeq2lrwBL2PIaEoCyjsgwKxykp0e0P9vmnpF6V/5AE4+Xz17LNaIRprSKD
Dqxvvb6jgvJdjohceyTpaW7dcDwBJ2nBPBI4+X9zBB5rd1PBdVpZ+cvQFgetXSlbfIiYyJMsYGTL
r/zl9Rn1NJSbfQRoZaWa1gMeozYkyYZdvW4jRrAXXi731WdQ9z/e6VhY1q54sAJ7mfTDzBBKeNsa
DFoKlryJLB9TD2kKkDiP48jf9Bg/Qd3IzGNjktgY2g4enQAPy9Fd6cO1pkjOVQ/2E1N19+3p7d7e
U0YYGOrGpCCL5B3/gGh2ZXaIfuWPIOQo5ZQgVMP5wsXLX/ITxwtMIJZhqw/99Y3WCqQUleuCrwKq
/6O2XiXH1iDO1gyWqXo2ONygg8Wc4rLLh84016/dwvLPeILcAvcPXewx77VuBnXW6cwAEmXE5AKJ
UDz8okxR9zfGWTy4ma5SdRKUHbnVEH+CFiVp04e241lC62Lz63/Ew9JZGO4LWA/7Zt3D1ECULOXJ
xJzrENm3P22MtdMy8+/m+jpE2zU/A2fxKwQaViAYLgRSuaqY/huruxGZUarX+FJ+M8CeQMBcfvBF
gfmCPf9NI/Oiuj3qqUxBKvAEJjvquCkUwBENpREJxjE61hTmetA/vN1cENbAmxOhmcwStsstWZek
vPyaMwpCZJyXFB/2R7DpoSPwdXqtibR+R41p+k6OLTMi0scg9vux3c5YwGX56I490rYB216ql00B
9ut3KxUsmDx2CREBUw+QVHPME0mdOvsVUBH6YBHb3ZqgPl8rLStP2y10Clz7GfewYAQAA/MQE2H1
ULl3ypSkqPU7PT0nPfCarW82Ud5iz+zjMPRLDy5oAK4xeDM4hhTpZqPCd7Vrcsgg96+iIccTFSJX
nLbNQJZLU4878cDvhLfUl/Q7w+YZKF5RqJWdDqJB6JVRrwFBdKmWdGlmjxGWMc4KQ2nox/9UTnZN
ZEDYvtj7CKwQQQt6GzcV31Bz1ZLmG4EaKn157VL40R1BE7lH3+XQY/bAFsFAEdPXYRYAsjXWjnnO
57GYrf9GWLrC2nDi1+cq1CkTQS75PNzFayTkiAgYFdYDU0FZj+yQEVvRjYcGVl3m4OnoWSn+QNtP
R/PLPS2IWZHwU7hIVeUGOgGtslXsZubDtEMILrJAE+MgJnqUz3KEYgDapt/JuCrKnEgtY1YIFmzO
bS0KUH03xop3EOrpbA483oWP5sjjMWLkUvwgSCW2hRDvk+d9+/4HRpHl4vqRmgwhNRdKc0JvjAWX
gzSr2/UC1y1UeN6lnrsKcuPzaA6p9AEzuCYKVl9GX23+63/OMK4PdB/YsIb26xax2xP2zigzNTCw
iXNQHzaYyo42w5q4IBYJK/isFGJ5EdCxMLQPtzloqWfE8+K8pukkIQsNswG8oqNpqJ8wGVfQQ8ss
ni1xNkxstoj8Dh9euguEw0juKSKacLgXUCHSYHjk5ro9uS47F48pMO0YM3w3v4qffKlT+zf1W+Ha
lhVfNsJwgehT9p6zF+oWZx5J+s2tCLlebIA757iJ3iPptC+JStdNC1bCedEpGsxTYNu167+sYdYq
ao5nNxB744uDLCAlWzGoF2w5TSChgvtQNM3rQRBjgiVXdj51EWGHHVUymi0Rk99d8SkTxx/KPNfM
RMmaqPEKIMVg2ZgXUe/HWIfqYC/v0oqGPh+85WxEYIgc58V6jiObdyb2Vmff+9boR94/YD6P28kQ
GyHfd6H314Y0he1lVAV9+IKH3alzwPLaPofnmCovxHTQtTZeaQ+Cu2ZJCVusMcq7z7Q+zrRxm3z6
eiUEcsR6BRmsm3LCNwtnREsaMvKQxFQ/aWsEZLwf4yf5NG0Epqb4qvJ9XU23Y6ERKqGjcqBRn3FU
t1mFcdo6uzbaFC792InGI3kudReTTDe6HodmAysV3UdW/T3RXlJOmU3Cq7oe2bvlNHL+NUbDt22i
p1dlMvJ7bvGgFVHDNLG1+67sQ+i922iGnAxvvT0afZ+hTvB9imF6ViYdNcuiTMsmx/mVAUYxUnpe
7iWM5x6iUz8Dkv7rw+JKTxG9zMC4oaet/NNJqPJBThUJE7TcWZYhSSfL4spOphTctxp0/40jWGA0
ZHB2L0ee1ijoSIWsDMFQ0aBoQp9zmJvo3pmZ/Q0eeTj8e1F2CVFvDmtM5oukCkRdEg5jwR3hSWQw
PxRy40ySnwfKvf7AEXFH1zIGnVg2+owQTdUO6SKvQvh2J35uS4dRD5bHrdMAmzawEHwDp2Ng19Uw
azjJpXnYSNyVethkJd6KQlIzIES1a6856IIoEwOBk+WWNGIVfLstSg42kB96TH521A256cDQzQQS
NVQ1r+i2z+7OZt+Kp78+ZOJr5NLvEYP+Wz/RKI7YskY1NLnSFTD6ZRlwCvMhrvNYEpMUcKrzsD6k
Z6RxywkegU58g4zM9jPFRoyH5zNsx1pvggIJDa2ahQknw1DZhiVcjWmMYLDugoVWF/U7QI62uO6F
fPFHjEgSNvvTfLXGBD5ue1B6WwyIUS844KR2PPDrOwY3ebBLfU+piXrMzaMizQQh0GLOcfJ/f8GI
lPTysAwMoSEDlY2fBpUgMVle1H7y+FChJxM9gPn+TeUscfj6p4khcPCo8cB2wE3iGP+C79nbRDeM
bnSJ95AYTXcLA6zmsRTTTLDjpcInh/Wz9rZc059jRt+vtMVj2r8t97QY6zto0ijve7yOSohEgacP
eCts0dwehjr2+Z6422kVPETRaCp8EFDlz3Xk/HpRtRbBVl6dqlUpvxN1k13AAW5JgNtKeE3mqlCE
MZ/eRqYf8Cff0jo0KZeYnKrcclsolOODQHx1v/vsrvlZlROIugmAd8vuWObGzuEwDYHNOuIVTKDI
/m20AvqLIbg93fw1urL+6yaOWtnJnhB1H0ghphii50/KWfxeqHd9FNIL8dyvtQAktMrriNx/UtYF
pE7JzbtbupWk9JlwN+cwwjGPIRUp+re2fU3IYvfUlmQS0RYGBTrMCpOdcX0drz6i6P6BLHKzYCpU
phQKXTD6PeJ2tNvMY4AZXRkDKVClNESDmpp2gJaTMrYaXBU3LilTkNu88RlgGsfA+a89w9gK8mG0
x1la+MQw6gVXdvstm+GPG+9oaJjIL8wO2CxFVaMHWGcm4dV1biCmViUJY8S0sxGFPKIp+qX8GfLK
dH3zBGrRWPu8gXHxFuktC3qx5bvGkTlOlThjlDbEy+cVWJ3gegOXbUWExc/7BeH7W/AphZtVTe7Q
PCAU5/2awg8ntBumpu9QJcUtE9C+dpWSIWU1P78X8GDFugR/5gAD0flJE06YCU9VfAhea/zx92Nh
1XBTOj3iDKAAbJERMJz/Tg4ISvDfU4XBNScheqnOUFNmDWgyPN7U7yUz0I8FGeVoFBMkWQfo4x82
U289lN/yKkyk89hKrWsOIWFkwWQZd/UCtSDQrPYbWkVGWXjG8fS4YZkBPmgsxZsixdcETAld77Uk
HK+3RfNQ+wVkS0ny5jKXQog9VhMwqnk6mGeB0sftxfe9wnvqdV2yYoMsL7QkwjYtEkx61wGHNSNI
CXGPHje9Ne6PvVeQJys5CRDhtrEXlBwm/PBgvJb36+QOtujtpUnkTaHiT6tlljv1ZeG/G4+0jf2w
I8vBi5znKcAqplg2F32lPew4upNw0DojqdRD1H3ALkMdvJTe4NGpR9dn/ZIP/sNcWBGM5nLDAGeP
t8Sc7uLpXg6wlWxiw0H9k5u9tPtne1UhkJWdtA/alTuqZlO+QVtJv+7yj9CLOPPyT/3+EHeLXVG7
9qmBzarv9psxKf8cM/L4ogPdjnbsOTVBOUyLx+lEKOEWvAnsakvGIIggizvfn6i4xPzrRY/AED+8
jkdUJKe/V392up3fh7UDHW8WHlQcrDX5Cois/rDk7UT7piCSaNObU3TD78jv84Q8TMkdHXWRlT7q
XU4Ow1pRWpzUBDpK/hPiAr0uHG9V/tW16O3zcgBgjWOGiCEtj0XU/6y1n069LWV3lex0A6oFENxr
XBBf4KRDfrAxJP4M/4DP2o0TZleO3iZpN2CQgo60fQrSm2QQAsHLgyPknvz5ixUEfoOm0Ati+Jb3
gu4bP3zArx4mRSULKsrN+MErVUi9qSy2iV8rl4/FWa4XRKHQ1qP5Hdo05JtNS4MzBLePJ2SO9jVR
iemeQuIVPeqdpGcfVVMo9dRCgXpcCQz9TamibvZuHus0yuMn9wNG2degfsF58yFe1pLW6oDvkLqo
aErMe645YWNTTtPKg7jMNR6F8+4LwhcaSunY0YSCmdfeDLS+nX3eV+O1X7zt3Hy6jdTUup8Zptxk
LMYm7nlOTgwOM2sQM06XTVX7tJ5tGnIPCnv4PHGLlxfGwEF9BzJc6Wtp8gYA3nLXTFU/IbgYyWtw
ws44jBTgv3jGWrc2HhfLMugPN02mfL/FvQS1TGswN4T4FbQ7k4HOBuZ6MqQEXz/2i8TmtHUv7aAB
nmNDpTKiuSlhU6I6ENLXtHkuCnFWvSDh5qmnQ7meYhtMnRoHjKbMHIQqMo82wiGtlDmRiYawbmri
78RB8oz3hglEwLvgN8c+Znn5UqIpCukAApeuBZwac7adYf2gn3wHE+d/vyYGKkzZh11E9P3JJz9P
TzwC+pQ6399PG3sArCtbK3Vyf2gXI5KAt/e6XsGpu9yEc2P+FuisosOcyRs2bhCR16LJVkqNnbU0
UIvpoPmsso54A/4HR2XVGKcnJHmHiBPpYduo715DjE84ybK8znlx7214efn1ntiTNtK+KKqRXKSk
SovTFhKESMqq3MWbE/3kTrmKdqxD4vsj1WqMBKkWIDEFh8weIwg/0qRsHvC3osnWrV+VGTRzZv3i
n8lEW94ltc2HmhV/D/6Ed5Scy5o019DxOrHoe1iMTgAWsO3NoS4pMunfOPsfpEF+AQkfKqyMsakA
d7/K0CVvYXfN4D13l9dsKJSS9qQNdHtw3Igeuiv3n84B+w87eYLwqWRlPuF9B2GGb0eHOg8FvSxM
5z6XMPqKvwy9DL2UhbcKzM8zz93XUjz2+0vOPi637HaGet8TPUmpDLsmVqeSCiXTVzk5xHodNuRK
X762ItyxB71FX2aSUAioVcIwvw0RTnq8wopMQM0gFH5LLC9H9GULRqekLu+C0pJF8+4N3stOKyxt
bI9YFdQBAPaI8s/u4Eq3xrN3kDH6OPXrwzO5XgDZEsy8gi0qaSSgNcYqT0FnTrAxdyXHX/xLpJom
EiVw3rV1E/TRZtXzdQswNci+3IucD+pF03G6hbNcVq52m3sh35cqcWz/rIsoJrK6E4cqlii00t/L
l2NLtN+uNevZyC2rC8rcK5RvAueKtRTvb5xJ0gxHRsQ9C6JZghU8QQpWVQwaGeH9glTAhswfFAoJ
hBunG4R57HVwmcd0+3nuw9e16LacBivxC9clTlAoGrRVDUa/S8TY8ARFRPvAxb2ky04S/wTIKqlK
UDeOaipTY+0Hvseljvg43qEaqp9STcdZqH7eQ9l3ZtQb6wP0oHepksPmTRTuX6EdkQWMjI+HfxMN
xtfyetVL9r8Y+eyk6L6owJSTHMcBAL06tTVy2azgCtdYFDDATIfLDiurNtrfS3zGokL5WHTI+4sW
8ckAyr7QDyA+IRcM5BEs27O1Ff4grKB3Mu2EG1KhA5txuKd6M5pk0k8AUupPa3vvWZr9ZeXMbUYJ
TYgm+eyD7m+LEgtTBHNYA5kbJenw9abhPd1cqLPHwM2fk89pK+z07VArxyS+9sPTbrvOWnch3qlk
ETwy8Q7QgED3SfSVOD3f2qy2DwJhmNvEqjU49AzvliUev1h7v0OaXr/B4x+2rAaHNNthNmT34eFc
BTfxL0QTYbcnw6FhhX5IwK/cKOVHhVc2Kxw7yjslKMDiS3qZamC4NUQI1nRVvJFxSVYQlFCjRDGc
W/K8TWeJFsg5dn35w54xzGZtm4RX5BC8IrOEAcItlqzUI7OltWf7l5lcSFM5Uu3E0ZflrDA7NZ7l
7eO49D1SKdn1cdCT5GAW3Qjm2zQFG9EVgN3u9oTT6s6Op9QvnAHsS0UPs1fZR/g1jNKScbig/f/D
65N06lhXJGIfibjDvh8Wt2XcsQgrxD8ohhNLPQzyZKl/UCr1xkb/u/1dbNrQkFPl8CZKfi0FoNEl
X02i2BGhuPq3wi0Z54p7ggt3i46A5Vwks7T7lTBn+MPV+Mu6C/hZj9IMoDCxaGE17Jhy9wANscml
0bOnuyeL9MtMoyNTCd0qArIFZsFRvahtSbs/3fwABXNINXFq4nJVmzOZa/pGyFIKt0xX6IFDMcaF
zV501F5U5eWfEElIfgLK4yecvpD5Cp/suZW2WVG+dm7KLpWmXxxiqBfbPGqDJWLZrmCAg2MtnA6n
M7FZ1V+1zfmNiHg1aqXJZ8gNlbJoxHuYIFgkvq8+Ew0iRgn9O+ZtRuVLGWVEQeWhYAsP2e/9QdY2
Dmi/N6Pf44LKrxgImasff1ZCaj4EoWXNuoHpM0jkE+UByNrcUyaPtm05PZI+wPCWXTxJsH0y8gKk
gSxcnISFwjXn9Sli65bH6b20wMQanoO2W8ht8hdRta5SIOS5NVW9wCEXVGP9+3NnQw1T7jlGoFh/
vACBf6EDt1jfqI+vegy4SqcZ9Pd3QYt9cjel3nXINBWdblfGg6gRctD98i0DfbMIfFJrINiL8hWl
TG9RtUrjFoPwXM8y47wjozC3yTBqqPTcQJVmkaQBBb2GlLtZz154odXEgNUQbUL9ykEWRBKEhWvO
eolR2RMyQHlTpSJxEXB6NXfeaoFjNfbD451y7OPxqht1a9F/66RT31E4arwjrijJVfC7o0SrASf3
rQA93fNFl9ukNJmK/ADX4Mh3VZDBw3Ei14Yn9uHXSNYFR5u8JQYNf0xfFumRZePOysgy6fs4G4St
cAJnC+g2qCRL5EJjKZX/KemVH6fdjdjolbZVr7L7X6mlEp/tRrOwmtHosZ0Ocs2klBCrt9t0KnJZ
hdkzj1nFTxgfFF4a5xr8H3XSOapcFgQdqCZ4OsAQMXklRgr80puh6bN7D04QwHtuka9QFQV70x1t
2kkXPT0BaaGT9/bgkHi4p5jVXFTEwoBqTfELG+5b1m1sXXeuzY0WqRCPFDOScm/WXX7LbQ6ohMU+
7x5YFrQqLufoPr1CfU/70kSB02tmU6QHt5+uYrHVbi2HWPjyxtkBRag4CmgsWf9jmrAcSeKDuCoG
R6xmRdcnkf8SuyVhr/iKRHIBdPHKwAMGnwA8wDDXkZJ8y/n+qqm/GQT8MWy0ZxmxphipV/Sk2lhL
zpTE0yEhGeqjZf8hHOwfb5s02MEjuOCLR8tyC+9m6SNAhLMHBMTyPEKL0M7eKN2Unt5hm0DQGmX9
9QK+Vp9h2y6a2tGWEoKM7jX+nfwXHTZycMquNC39gPI7FYk/K9VPMOSsoYDloQaJMC6VB4iHqA+F
ZlfeGwh8epcBhHFR5hDM1DcQ+aYCT4QrNHKGgjGq19Tpq7ndJxxDe3lI6dPIoigh6eOvrV041D+2
MkO2xZ/NGEfOW3JV9goeICFKpFg8hMlzCVwqHuLujjDrMa703ofrYAR8vB4vgexkeZx2S/zyWJxh
mdyQgZ0xYZB5z8q4CvpUJEAz0KqReXMqelP0FYhYstOEo8aCuTkjxb1RnFbrV6yKVix7E2nJbiyI
m1hXWAZLLIL1OELK5Rcmh8/Q6xh2CMuCg4Zeq8//LJLovb/WW2H30F/hlWq9Q7hdKzG+o6edYwFi
40UUQadbMsU78S5DkO8SGUXTFK5TtzZJCOXx6jKF/JiW3T4BpNRnZezjdURj3k8vyVRJy5PyTObI
GQpTjqJHiLy61RP3QVVERHJ/1Ss7ZYWJClapJwJrvLsV9UZ7jDGY1nYgbfJ2OhySW9j0shPMBXFD
zOX7crgv7cecvli+Jk9n7Mpn/p/GOfsXIlBzSMmC31W8AZk+8UXu3pj2XfOXGjda8uY/YNn6ZNcX
k7C7UtxZ1P9rfR/ZgOBxGjDSXxLhaMvtLmZNMG/MwD+tgEMMF9nCYstDTbjwI7GKcStbZaiqblyC
6yezKJsNFpHhnoKQzaLiJs/2Q/Kl+dTghk5hZiqb5PXajjrPE7UZJOZhq2IbT/XbGUPE2BcGq50f
om0zIt6ZYZjZto+r6FpGmEf7Eev/CqQpTiBcJtsdhOxQeVKFIIffmaFQzc5M5BKlorI7Du+lpXmN
pJGYvfuL5a32k04rcvxFpfGqWLyc7rC3HR+SqIuWCl+9y+FO68RrZRLq+GwTi1Kyadh2paUJvW3a
+VKjMRHA425I/ojxDAeB/j18H9EQwsFb84pJHWhZFHrCQLVokuAoMnmnUYR1o+xQs54fBPAwENlG
gwWLmSkGVaJMRVdlfbI386XKq7HzR2A8XrnOaSjsaAnyW4pyCbmJb224KgqH8ZxL/j5fXsvUVwQm
ydrhSwE9zfrhCdvJIHvvxV1goYFx4+z+BIySYTVhZnYmW81zvljSFweWBwPR31t3v5KQ2JzTIPh7
tbykNCFytbv4DeuLYlJd+6ixbHyjBVQddJlvzzW+oGB5amjGglTgdCz1dr9I6jJyqFidKJCO1rqe
YI/OWWPBJg3UEqckimY5YcvRpKSa9KvFw2I0xNcvkY7LBcVXUsdjGXkcoYjQWBySsK7PdPER/nST
m4YcOOZ/NRNlfwuqBGzZETMZs0docICepe1DTiMVII79FIrmJceAhYF1cgpbxdBr8gTFZYp44Qyl
EURf6dY/qQKWedvqBAClkLqA33RimIq4O7lzLcUECvPKxSt/1mkQ3KOycv+lPWl+VeAqHLwKqo7y
9gA60XqIQ8hwdsoQBC5gTYIu/SJMvjDfU8bYGp76+2HETeOXqp9jt45XJJvsW2Y3DJlGVkEjE6as
3w2pq3IUYlijHB/qQJKALY9zwdBkaUt3pexycui7+FK9Lxov2HaWcA75e3xC7beYPN4/34/dzL/u
iu1ae9NLH2GSDG38AondZ/7YeR5SXqcvFMuUH2heu0dPV7Eauv34ynNu/KvFr8nsmFZbU4ORI1v3
c4V0enmFxucpnAf1t676Cm0d7EQSqE6KZqR7XUybfXXEV6Zcfj72zeVsov4yaDK07C876qjJ8l+r
jKAw0lkCqnegi5FkWsnfAaPi34/DVh6hdxEbcq+PLwv/Rvrk+N7accwKAzuZBvyHpbPomMtw1Hx2
rhdFjKBKu033XYv1+eVC18jJNv94jWJWxzUZkSerLxJO60+ZowEG0UdXVWCBKhwmk9UV2+dZB3WM
nediLmCn4OFPFKHPAEWQtHsUFgy7Gr8eu91RA8pAZrj0hX8anbgl/r7YbAfCb+wAdm2qTIvxoDH0
wLaV8LyiNOdw5uGHqIDs7/uh9Ptze549D8oyVLZgpsP4AlysgYsmNMwmDD9+VUwZUB45aDrNC7dT
4Ax4hZ7MRYhTiS7oJeu4ocBfwQ/kJgKrI2Vkw4Jd7oIcogN14EnPjOyP5518NsuvbtHaOFQJpQIz
qTszLObUHuntDQGda99Q/fHY/e1jUd1W+agxfzw8inm+vsUOBvP99M6So4TJpL4pYNnMYDz3wRdv
8TCscMyVVrDnRHXy6utzzL7cMuz9usUzQ+R8+9AKeE1q4pnx1giFiYJsQfWwpSveRLk+qgMq6bkL
fUYAjjlYXuVlyyjXDMkRZGEhDk/w3yZgcA0ybwRdyA8gC4swqHdJcDI7NQfguPGWpqJEe5bgoS6X
TQbF9wge/SeOH9FZlEcxuBHIWQfeT6eV4vtGV3tm4+4hfS48zUqM2KzUTZ3InxQSb8qag4u4+KZy
Z5mkyFRZD7MRmg4sFUaxIAJws/ShXpt5r0/vNHMzcAmQQeh/sXFIkMqMUDYtCFvGHIazZ88t4A3U
Odf8FZ5FO986Ilq/2s0LLv5sLb8j4BA1TX+U6hsGjQI+XRcPGuPMUdN4umWcKc4lAjU6lc8xP6Px
15I78IsPGfTiZC7ez/y9pz0zwSNF2ayNZgdVcUhTKKJEdg/OpMvgtOBrBCxK8hI3A0JsvJqXmFRH
N29U4e+lEtO1+lTlZ5YicEAM+9tjZDdOHUVQo5s0H+ogldTuGbYxT/vixWFASg1eF3A/coQNbSk8
mLOSiuzJdhMvgRbtIRLe6WV9OM1u1i3tHJPIgJxyHIlp5Xlb2fQhfsBl0DYPf5coD3jXLCQLAVRi
4As5eXDZ1PtjunXTs9zwTcepEKT8qkRwsKKX7bsCT28HhYDAukJhs0GDNPLAdpC419R/J9JB27LD
0LJLHmXo3YDcbJe0O/uqjKBJTJtdYmEzzYElmT7pj85P4AFDUrmZGnZ8Exqy4ufXyaizTUHc+Xd+
2Dv3acqlfdC9XEiBOwSAx0LqcwWfQ5rjqtAdx4q932c2zutNz1p+yIetK5imb/CrJKF4j720Lmht
x8i0i+c8o6jLyFjJro3ZAB9mvFYZQj1hl+jQgJM1NJSqNrL0JpdtS3ech6WE/R1ws+SZFQxh4JLN
FKNZBYsMKLidb+gQD8jxEzNFoFphbZP0GkEhNJLXEeOxRT0MG3AG3g1fl7c8/Hu8LalnOPBaHnzo
JKT9GYDeoZBmj/0OMJ4BIAdXcwLgyMA1xNlq/IguSbZWzTBKCecpEB8E2mWMpmM712BHnt7ttmDa
zTGoath0HMREDhTmhdfbFdhlzqYIkcKe0ARui48nb6GGzXF50Vw1fahwxwVN5AbDyn/+gGdxp1OY
e18JPBIse+GzlN7nYXQutnS6EszAQhFbuywBBfx+BmMapDBE4exZC+jtMADwvjAQ/tcFTpMrkytt
6sf9J9R8ZyohUNoZq5sh3oUNP0AD9d6sB4PGGYsqMIAeHJdkaYruQ2KRuN0Ug55O5FOpAll2YpIw
cFhmpu2PNXzEZhUqj6PF4xYKiEkgksR98KjY1k306gkkXryA/+lZzgBdUswFuJWxZ5N5Cro803dW
Vgca4kG9Sn1uYrVmyqV/3oATDexcjF53i9c/Fq8ClbpQ8Sp3bydwK9BgFHLV7jebrTEFLHCb7Yek
BvOl/lrQL2cQjE7Fef8j8f6dBSf22DP/OVwTUFyOxwEiPcn0VPW7mXTuGd4ZFS4/ga3jNsbKRUWQ
OCD5bL2SLeDFzTfUnhajeavy2ITIKrXXVRKRWvpSXgqme7SpXHTLYEnhdYlA56qoeteVjQrP94RS
2WqYccHT/pt/nBGcwQDWJCivNQC89YorayX/h1MYCnCjKpQXBp9G7dr1AhIQ3o6eh1kRayN7pk91
jUqGN0WH/vu3BYsV9LEGsXJMnd5uoQWZsCaFtS3nsSWZbUh3tx+0wbZ3jhKvAxqT8qfEbo8/vB7d
xPZceDrB5BZ1eopqLDicbwnaliyUiNHINXbQa7yt7BJz2RVUIVWf/h3u+Ea6Kpa1yRvGwEOdtBiw
UytyWzn2GbceCxH/1iGEk9c9ufulOMJCGhFdjxTgwCCl027JP8n6blNs8z6TeVfT2uvGtUYJ3kvf
1pv/55Cg90oSAE3Tfu7+Oks/W2cQqXvAs4xc36kJOaDU4kmOoRjPUDHo0qdM0PF2tdFQ5Q8fGqU7
ldSRrYBOWaZyaiGi+qrRXu3K0Jz1CtFvoWsdWs+nX7n7fyZgPF5bijNPeVclg6mpZg3UupTI9m/i
HGmCTj1ibTZOEOEWgZrPaRqyjN0K/GHLVyf5gL2zjNrzU4uOc4885VMsuVLs5KE8+BZ20qNa61NH
SsCNhTB3w5VZNYiBywWifDpLKNT5ukYWA+HE2rdbryHBIQBNtsP2vCx+rpAp4rY8RBweU0gbobwX
9BDgcaTHkzd8eCJNEKR/m9PM4CdslWyuB/uf1KbfdMkX0CpmvanUgUJZdovm4p2SjSaM71ED6Lmb
PitdhaT2Sd4x86PRIh76JYM56Rdgu/QHEWaje/bN3kGD48R1L4zuW42rEMMcpqz+7LBmVgc/zSNR
8jCMI35BYdH2fhFZhYnQ86OdmCcLP1dZXq/wGRWTiDSpmRqbJ2w5PZDWaW6hJs+x2F07heEsHZYA
CWMHLawunZSPqtBDMKNHGd0QHpcVO/usu9qW3+yuNWL5BJ5BBv/QXMU14yf6i/Fcdt+LB+CZCuwG
K+jb7CzlGvP+QWftVeUU70AJKFfy8y8QGgOh4ql7MmV8JGW7Hn72MK/Znp9vXFsWb22qfhGNOu8b
nbQRHl57P8SMJuP248S9bS5av4kTcnTWiBSway7xlGiiYPVNEExaT/YIJkgb1beE7ETBBPoaDC1C
EkHC9RhsvFHBX1FEZhUvjfxFqN6L65nwl60Ulby8UDfApxlRehBYrvZvi+yVUd3Sn/EHtCbza48D
SpTyIOSX6/AKnOPPU8DgdpBrMbT+lU/SbYzuPVnmh9m3cM51i3VeJiwR799LY5s8M2q5H8Kiy0Hv
ydu/vzFMptvYo1ktrzKLTy9dhiaq9zW+5LO8TkQrSAKRMMVQ/jXxS5ufKGgRO4/7iDh2PPqs3KYF
WjVpIOZZXel/E4Eu8qBivSWjYWdvLkWQyOd2vQTJGCGKvVPJnTGphyPiYVb4+Q+vy+pYRfwRx9zd
IeVSihgMUfg2oIgIiTs3OsyjfiF2tiDMbiXM+C8QHi/oHcoC9lFjolF4TpMXC5BxFk0Le4YMJdH4
xmFFK5ARlQM9gpdKzqpS4k6YwMnrr6Ao7KzPMO/bB1eJs0Hs8svc2H95JQCH49zg2tEPl//IEPGy
yXiqv+ePMQq5iCTQMgOMhKIrczH3ubVM9ytHSA0mN74rCrLrFSKtCvxZ+uzRwpgX5C9NtRrhohVx
rpvn59Dg04icPAAkk51LnMbVbLGd70ZTMFfzSE4Y1j57n6kBMf29jQ9s4pS8uAyyrDKAxffj0ooJ
9C6ms+yzwBDjaLURvC+KSXGPHOw8yTHd4MBapEpAT2UyOSFNdkf96y+fwgbhIwwc7/wwNB4upEfm
H6N0JycthbFVQQHP/TyN1fLl1uJtSLW9uNfedNn1DvxOhDLYtqNKQdR4VSjIe40AaSqfpgNuD44f
xRrSX88/cA2PGXAztd4QHJRZ8d7iH1TUA5ARB/qVZwHZZYUHH68n8OEdtsbgDVNj9Gd8OFmei5An
UMiEOiDVexNpuK2xes6E0/gi+phJWK8BY9F0nGWuMEhGmpqCt0Y8m2sC49YObWEV0sFnLUdogoQx
n7s3FdTBTBnTL8A3DvAFGJG3Ji8Iga89imZPvFpgcTYXCfY+C1igMoe8Vt8O+dXAKcar0PeOcaYF
5dWuFZnz3Yiie8s/ThD10p/TdUpgP1N8X6mgn2dYPjoU+jTBk/bp17MM4Xgt56r+XMH/PksJ+rRI
C2VY7ozfRS9txo1QhyKSi75E+thf34W5QblKyZhwx5vKtyN8WUo1cZNnO59EWKNEWlkB+sbl4CCu
xED1PEnFUYjobOQY6i26RdqIRsAryKUY61Hk6OPNOEiPCKMPEmiy3PHNu0F9beq8QfFdnrXok8Nc
XnnMoBo/fHNcpKCcWdWAxdZY/qiGZfLgoQE3y+BvrkWQPEpw4REJxtao72LInNEG8JavTZrk8q3W
lzReMCBv8LvJxrjsXOY7ztAX8p1JMoGCUqnazOyTf/Qb1L5lAZiklxpBs2A6fvDNm0kE3yhfcYmv
+vqwgzL/sw5ThGA3reoUT5qzGyYTexX3ha9aYak897+h2Yu1nRCTWa2uiv3xUWNG5QUpSaCSeExd
tOr6ebhJJQbY3yf9uN6+rvlcXWm2jwHQc0GvqSKYd70Ar/UknIKzb9xL4npkk7pvYVdJ/PX+0un8
Hqvb/oBlDovxD0LFjuxaIhYCySls4ydHa6TcqvKC+bZYrvp41Q7ZFhb+qyN2TH5oqXhiFpQlP8Z+
ChfVDIdZ4NyMfmePehrYquph87R4Gx9rB95c6TKNjOnIt3wIwnwsXZtjcVMoCd/6/b4I21xx5WYt
hpnTmEYwU55ANrh2ItbBtZAt1rfAHty+BdP8aDT4dnGyDzOyzYcnHh1ehuDFnLhcTht0Egbv8h2F
SOBGnaMu08GBgHYN5S+PGkAzzX6DH9olCAwogEsRDR6i0gyFC7JQnC1NBMjIcCv1bUiwpCNRdJU3
AdqJ506C5NLK24JAykEWbVB3fgAR09JTkaao46PQGR/x646XjDXZgwVaAhsOCYDtv0O/H5ojfTYo
mYwQzQ2RqrlSZjDIomIIiiyXKv36XozTNkptMq59SutKYmirq0XqSvBUUJnVX3P3LXBRCJNL39MQ
pGoCUkOZLONmALSF8ZxyNEcVUw63jFgQ7WjwNOfr2693xQx01JWoihl6UQggFDhn/r8FjSMPNkJ+
scAM723aPWyQG7QqoSOwcsVvaKN5faItLHSmYDeU9TJPKJVrk8P9SYPb59MyxJFhmxgGlaDhdd0s
CsB1oOOccXBqAhHWDP2GzSg5ISOJFYH7DM1Wmlp/6sTqTWzwPjmwhFhQ8QP6/V8h/acWL7LCRzPV
NE98enWIN5ytzOtGV06Xpwuqp+oBg/W1AOYRcvw1Jd5hIPl+uARnI48qKfCE5IkceoeP3YVbf+Zg
O2SGPfmPG9U9XuXiiwAAXGGRhSk0eCBqFUD3/eMoKJgcU/VFQQUxsXMN2VcQLynJJkK0dquoPcg+
2JdY/3oW78pmtTtVAIBuYDds+My6mHL64l5HLnVBgN7arx0FO65fWOifldcA1MIgBaeH5ys5QiUn
twNoL9UJ61fcgHA52EBFrjKaEiz2TOehZCXPCEfuevF0+UyoldJCfbVSh668V0KerEpoy88RRV7G
NM/Gdj0++ZT0LkEVR7zmgtG/E8hbKMnJYDrpz73c/fDMVA2OwPQy7rrt03SK0i18WyjFYEHGMCEW
1plHbIex7g6bBB6DI+5cS78q7/i2czZJ5AIqcCpU9bf1Po2BBPNMxTP7LohJ22kQ0RHWPxIN4zJm
/BzJOfCr2EMAfylRUbUHOL/35XrMedFFRrXuhRI/ZbXNBEufqjYFXhaRCQUc3WRJ1qH5we2Fzik4
HiuOuLwDh7/xiMPvxGm52iiJE7uWTH9ClzjBQAHHyMAnyM0FYQTa063Pke4XsFMK2RAbcDZvnRAD
+bccgRCjM3A0C25nW6KSqw0PYI3ZW3yEYeR3+Ix5oixHpSEC57WkkHRoLsTy3UAvySXThfvHHU8D
Wos+PBLs/RZufhSjhQmB1uRg5NP0jhGb86X/TrMXJBb9R3OC/QMO2UOCK2YQRWFMyVkgSQPno9hD
0AJH6/wFzFQo8+zRM5p9NTQQzOLulOUvRiI8ILLGnQESKYR+qOsI6LNNCIsYIpIgpH6QNyh2fANZ
1svk6uiJ/XM1gPFlKwa2AQvFWHTxzaeBxHy6pD04UrXMD3qFVSTeFkDDb2ZJdPPwjz/quDV+QowW
QM26qmIouq7m5mB7aczKLqBnNV93NYMSSSNRUcoPYtsqT8pmGqD6VhSfPZGNMTCKBZvOji8OJIB5
2DM7IQ7xOen/bHQu+evDCJ9Jnuf9U+r33NksjdCELH9e9pkKhoT562xtCHhHttoDsQwCH3hf58tl
RKE+hfwuYmB8qHUqcy32xvfRwX2Ztr9ir5WI4UDLTDv8IzT/VAMkE+dvsVEU8zQb786yqRmOuq2F
2u5hzub3lNSa30z1shS6Fhm0Dkh2whU9m//7134Lkh0PlqXkJ4kTut9eqUg2C4VVwqoS0rk12Dka
+DwJuoVMdyDh2SumNUsidOo+B1exKGnaPDE5RBEO9VbCQGNH5y2c5Fx2BjB4Pfduo/ODfmcEXJBB
60GiLh5ZKOG1vvEJlFtAbU/kJB1HRnPb3yppSjXZAu8ili1ofAm3+YFeQrNntI7w1b8nzbZmMIgh
JLUuQY44BW+zSrNy7tluXlPlBIbDGakRxNlnGgrUpFVA945nX8iza/CVKTMLAqrXbhEgiyX8L3rQ
QLedyyFlsuydFEyifKHddhcz3Z8GJCZiPkyRzHoPybaU0SbWe/7cxG/Uve7WVYnY+hZKhg0+El74
O3RsvHuCNTBftTor+OWIq00vfSngYait3Z/HTDBRHiCX4inikb7N9rKU03N7qbE3/R+QTU39Qoe4
WMElWf9nPzFkf10TnQkPst5io/+JBrWcZxDTacFanrR/bo+/20TX4ZrlDdKsbDmqfOS+wlJjKLN9
7CQQ8OQpvLOVDzCyF0fapQeADLi5lJt98q5mMMEbQjZW7tI1O+SpnSZrn+F7SQNeZDhP6Wky0ALu
slgPj3kmECDaXBAJ6fjr+SMRFBRD2gN/B3FYDlKHapip5MRWyjkf2edO7oXqBB0COSu93ds4SjQK
fh86jSvqzvj6fbORWEubWQmEoKkv5/cgjH6h23MuKTdhfC2dbEPTdC3PltE2GwwWnzXpJFn5y+45
rvTMemYHT61qu9GYQUVdoKKzswCC4rRfBZ1TtWhNTOcQrLEKI5pfqlLrMdUE9chj4cBsAJlNXmT2
Yjk6ajAfGKxwuU2SqQXQIOUk7mLZ5yP/haYj0KJjF5IFfUumTgFe6SyPfFE3VoKZv6fAS07q849K
JvwhPXjajq7R4+gK0thpmef+bskivkXLoOkMVhnc6EU0kwcgS11sJrnJ2YIVeraZuI8tqj5tRD/q
pzgr3Yzogr5K8mkFVeyTV2A3FsgiIx7nbHBeRbXB8EZ7+Oolmio+Lx0xVDUADqBh3++EaY7347KR
z17q1bbi3V0CvX2ls95+M3A2spWmuelM8yvPZ9FH8d7EM2t4tzdhHpq9oAcNNI28aG8D4m6wvj8t
B54TqT0+1KjebuRkVIJ/ug+BaUcKP/cbdLoKEU9SR4sqVEiTrGDt7Hv5MRP+E3sODBHE5dOXOzeU
4w/P5xHCJ9Qvbr8A56ow2xBLYEpInHB5fEXYIqZROtQGIXGbsgMy5V+/48PpfDbdG6rE7rvlcUe6
RZ81GyukoOWMRjCDQh9ZgGfmadnidJSy1z/PaFPsZiwMS3lenkLgqdwmSobw9WzPovraQKR0iZYM
ob4iTm0CNUBL/HD66S9CV45+0mW1Ax4+syyYLk0b5Vr3ZM4L6hBY7z3LIEJspaQ+wfvyo/2rPYsI
cME7yuOyWwPysde5k3b9F2/7jhMMMfSxy7ySTYrsPA04ucjitopWFRn85h8lGXEhtZa1vzW8IRn0
CGCOifUX2JIkFS94ISz/X4lk4ww/s1TlWQPD+C4NTR5HILbD0olCL8xRn7rBwJ8VT4vrHhEqwRRv
Z5XO1l4uTSwsuNAwtv9sfk0s7YXiLU2nUxzGCPeK1DY1h4iZqgyg1ntxcly6w0G1JVfPbFHphtt+
jEJ85RQ1E+RwRmBMKLnSFOD8BQFgMREpRalj60XChEGjfGlWeCLysUNf8VGa/E0NJ/+lXjpP/Z+x
Xc1coU0oeEgwqRbIunQll69vhVkZgELS09/ZSBU4z0oA3V8qyQtJjdvgUXs86ug/xoI1gmmnoF8i
kvmARLKRc/kyEL4GheNtkcmMPDAmlfhAhFYKGPhm4db90eVLlEiwcIhY2CPU85fAbVsrlJifVvyE
1nU/nCYPNXZVJMDsnSg8gHpDzjuxP3P7ZniwT5Bpw08Dn7Zqt83n5BfRQeTv/xmmMKOUqtMXcdrp
e5V9Ocge+XEpwBtG9NX8Tg6yMzqHk/i4yVCGcrHgMPjsYAyXVkNjWOoEll7f4yQRfB8i/CEzH0LF
NWv1hIS4C2tZwZvy/mmeD6Yr2hQVDYxiLpl0et4txf+0PbkJX+pkvoRw7QfKd3Tm71CyWdmF/SzN
NBvd8MzzuMTYbs9B+zoliOU9j1LMNkgFc5h/tRMWl6W9L+s4kcrCwYexNcGA8hoONYgNvGv1b/py
PEp3hsgGa+HL6ZWviB9B2EnclivUljJ3VVyHz+Q3SVNcso5HVNSrfpmG7WvXIrNv5H5eZBaxMy4I
mzQ7QgQwDZTL75y1VuSERjaTHFy3I7hrEW7uYeBL8dygrpH45IBLin6dWTvWDKLRh5kNtSuWGTGg
KaypC38fQBC+MjVj+xE6W+qpZHA+uyu14nJ6ADIHTkvf7b8xaFX+0rdfrZbdi2URK78QYmdjaxBY
2WIPqmXrRIkudNnF3HJIySh+bpTO+etFDP1TIm65kJ9WcXrIjHKTc4mCcd5dzgoxVa+8iQekAcY7
IgyUacW+4uAXyIU+jGFi1+LNtcDA4a1bfCEpmnKnFUfixv3NazlBAVVp/wpCqUe4ucOxgJvq2FH1
aiZK0BDAg+o74olJU6BLcPxwSu80L7rS3ITQyaEdfBmT6aPInDf7lW55w/6fR4pc1tAIs26monW5
ticg/cRjEDP+FjtIYvaK5iY5k4kDoL/BacKD2CmyMXCC0GWiC+BOL1arpcwgZYRkOglxVskBuJF8
12mSVG5PlGhMCh0DnfwxjTZg/VwFzwQVYzZeEAYpxZX2pPlJASaHRElDxxYonO4Ub7GYwMAtdKnP
2Vd7nqijE5VviX2myGyPMvCJxRUrqmSSoHD5Agxnthlzbo3rIMBDPKMg15XjqiY7owa0kt62luAM
BAcKo3dU90H8CXOqmGSeef0aDridUU35gkHWogYeyKnf18xDHv8byeAXGJF0tLaTPMxzRzuqmjw3
sUvaH8GEYAgBRMLU5x9Lvx+9Bacf+TUMVd4zO2btyw+zqL2atqpincubRF9rI7bLLY+I2lfcrLqm
5iMmQuq/nqcFXWGjqoyngGqb+rXwtkJfAz93bTBriUqjVgSF1go3BhD0awYc/9Iam2ln1NupgcE0
BFzuqigAfIZa2buKyOZYnNBYXS1AVd7Grs0wz50tuqjQmVhQm4kByRTE2Ja76nRqEVm2g7rH4048
8b5H7CNAivWPXDhN/+YtaqTpQCeUrZ3y4sJ2ewUjRYfT4mxrCfXylaE+3C6u6qpBNJwZtyrIX3v2
Ko2Did0N79YgjZkCadDmyAK4vtJUd0ePslPB3CxzBdQyB9HK5hKUNVc7r5vf4VsPbfM6oDKFvvGb
G9S3tSftBjVR12wCZnlg//asWTxTmOVFEfMBz0pmCKxr3X1txXVZRVfm+5CQ35uKknm8AEnOjgRk
1nBst0E2dXg+9+P1XFvLaIwvmSUN3LGRqjYpRhM8K0CqflrV76pqOqlPYZmToVDgJ/4DNwf/JhlA
PTyNjGJIDUWx9QkvkPhEh5fvFfV2L46FLAK2eP4VeNPqfrqj3t/wqSt5bpTvBxcguUHrZ4KCFrq7
XQLMZrp91FwzxY54bb1ffNsebF31qRUoU1FAD95mxAdpuOhQeje3so4yWH1mh1ToqEupdIDZgpCt
5eyIHrO4TKw6mdt70/e/C6HROTgZ0qvxiy3+nkb+d+7fFuY7nWtU7IZ1n0xjg8uapTAfJZUZWS+8
0Y9lt2bU9zu0tGtySh6b/nvdwfwDezZWjUz91wSJlpeJ4dKkCZXfrNEsxRgvZVOzlAC5pIoQ/B0k
ctCtNFK1QtE/rn9vwqEmlL98O8dOCaombDPvw/1d+LQ3hJa7DsI5NH2uijdTgLWPvkamlS2B3skn
+m4JmA3XwwMtWmG5Jiet4JLaPqPp0KRf90KvKAJTGdKV4cpsmD0hsLzZxG9maoddIfwTFi+l4tHn
9JwDUXSIGxbZMramJJ9NF7dZMOQfwRiOgnE5m5YEb3ktqn7TwLYYZcGrdVhBpIsokIwNNATVUUMe
QahRouFqOm68rwHrbjkiQ6zrHMVwYkHEWwYLAEJtL/lMVJDmqWnOzT738WKuk4jVmmjyeFGwNBr4
V386s5MJ5n0Li8WBOpNy6c01GKW4paNEvsJdNbf+zneHbN88mDKVmUtNbjkZwyWqEf7ELO+ieU1+
NavallRpTvHZBFfgU3e2c5kEFw2MBNmx7HvLRXWyg8N0OkAYBHAoDIcis1mUA77hiBhcebVRj7Zu
sXZjLnbOfjd+A/IoqBh3bESGRsVSrQyaOiVSrnvUZiWLkM0IbNpTATJIg/Ixp6qkrirJl907MCHL
DZnmXuXtgpFpiaPOOekHFeWeAwTCMJh5j9qbB/xKS3ICLd48xLCCtcaVljvyaaiGrjH9eADVEKUL
SfGIPQh0T0jyGs6f1MniiAov7brpNVXVtqErfBkcsY53uCAx/bp1C12Oa65NYW+RDzZdbds+6BqR
3gwykVZj49DltdB8KXaGY2j4wfi26eWXkaKJmJ6V8JpbiX7BPZbb3wNe/fxRSou3Q0lXIm9OeR0x
HUP2BC7JrtpjfwAMhtCnWXdgB5IvvsuGj9i02fdeTRosRT9W+bCoF3x8Z0xFnVM/9piV0xWpghKm
pT00/XgjjYzqa/NtVRTeFergGiRyY3uwOgRoBktssK+NMJYcjhpLx7/jLuGBPoFBGvcPn5iS5an/
ER38B2/CtFZjQWheS7/BOtLW71Al+e94BRPwsMzQjsrHdJNYa9HuC0f2/rBDoSSpmD9Jkvsq2z7w
oim9Tt4QB2wzAvHvlF58uz41X+V/n7fYy6JQDExUiy+sWoAEGhH03loWTQAlMn4A8L/u3sJaFVJp
8a3CIFBi7jNjmV2F7jzQkHqPYU3HpCvk9M1eS5zVXg35V2Sj3BoD3Eluo/0Z0nZU69Bcjpw8kc6n
QqTpBT3nozUpGw6r2ZmJejiJs5juFD4Cdz0VJbcnh6m/PZBELeRHqzReQN9TYqA7XrnAEIk/+ly4
sQr2MqDbkc7Gn8wacI/P1HLicpzo+UACyMMspg/TYY0K9ykvz0i/9cJXX766r8Y+tj+BYn8ltbDm
9LnI1v+8eQXBV9hZ+Mx7ZzoDsCVVGKlmyme94LUOH8HNL4GNFtTA/a3TBzdfUBhaYbQLJKehbssI
618jfuh5YaTp9bJcDGQbiKVk+doDNEupQnQrsWYdz5VyC+p1jyqSItOOZE1x4EYnuisuLuBG/ewr
KkFROrQJkyUfdUIz3vHQvyXEpNd8s3sinTYerFtmRFSveK5TjkZU1Ff6X14w/Hj9/KNEAnwt3jXM
2nzFFQmUm8lbNRZkKbhBAXsqTFHbSXRx0BrcB4u6PI12vTRQtNpSEnitzrmvNEca42LM5S0WeC+U
kap2zhXyCy+WsyKlRPIP8UD+W8aqo1cYdr6tLAI/m4cCfnx2XhHlKQD+7gpPFHmP97sCzJWI9KvJ
8u1uMYkd8VDs0nf0V4x6w1XZYaNDXQxUNhMQLrPuc3QBPpocKaFKzSFhrbkJWFtOKM5IMGQe0TH8
bktd5/wizlHj1Fb4oOJ15N3lI3BS1DfRQmsF7z0u9qrZIEZI8A2Uf3iP8VufN20lMlmnKgjXZ0Ab
FJiG/WIZRZdEs/LlV1+b9DVTHqt3wr3i4FgzptYwmGr9trXpnIa57t3L1Jo2B7KeeTFdGWACqmD/
c19H0khDZ6DN1iUAclbjOFJ6p1zcAMx0RZje2M7WDTPx+PTlt1JnZGFuwUJhDjVJ6RJKmIZbj5II
Zus3mPfP5/+MPR0wRTlGce+3614r9uwmKZy7t9jhCWrRMDWWUgtS5oRMWI+BKRNC3n8HCkafs0xz
sAQEcYDMO/CN9vA5qk+N2SGiqAbz4xqP919VO/avj7y0hdO676M5LKUiyvC+GkUsRV6HxtR0nsZj
XytyAHjzF+M3CRHyXBUpIJlatNoAtLH/o2jmXWNJVrvqaGVFU1YaL5yPDEWBDOvmyGT9lt1slYbm
gQqr0sZWeXAjVBFrzOxEEVgAJ38V05LmDPpLtNUEELJBx6nPEI/R3st6LbtfFdo8A7bnrMkDVI+8
SAlv3E27tAu2dumwTmpOWXjvLCEnoJ7YP4wM62j4OuaAy6YpTl5ds/QSst5KaSY+FAvav/NLLHvh
WPwdfpMraO8bUxMTcPQ8imaL0iGtf0c7TkFD0JZhSVCB/I9c16dSoLrQpW2LQEbOFgygX7xilWmv
raa3nKXxAQaEHacVLSPL8ld1Etdexzm8DXZ2RyZXzXwMV+mndyg9z0cdqMuNyc7soKAQ70mnHwfs
oromvz/Rk4//Yyg01U6bqAJzt8CG9nG18ADvIFX6WQRCoW13sN5yjH3fM7ouhOcCAaDj5vxUw1fd
vkduMRBiNJKTfkRVeYI+twMUgjSiHmaQd628d3U5efxRwb3w2v/Z/BOeA8zpJMkkIvPn/hskjMbr
Mf0z4odQVOCJ4ZprDLZCWMzcOCw/YZWO0Vm+ZWd50h6kUle6sKHlawdkCGEWam05VcQmMsfIt8lw
lMoH3ZxpJnkBOnYN9s30r0iBKXQsS9VugwVWIt3ixqqffqa7af9TaZItSMq8XMSjvrkcUu0QuqID
AJU0NOdzd2+T3VjZaXAaAc0Bkm1ThUeWQ8jJ/4ZnmQzzg3QeqfALh6oWlL4x98unCqI16CyL/SEP
qQjWHNI2LSLptPtEbAllK1v6aoI+d+i1yEXZwWMBk0rPf6TrUkUWDRr0A59FYaMfGpcJOU48lt05
nBHIhl2lQk5l1a+ZUJ4AlCeVCJBVqNFQ5nBB4BHbvfVL9rfBx4SFlVN1qYjH8wDhkzBxvuP2Pn2S
nG4LDYZI/lxiPnWXRHP9G2qjQ4JTBgUu4MUNy8wLSc1bKFTIqPJZqXRKNen6A8SwpWEeJOljJoMY
zihBLc8lBSvAgE8QDoaWn0p1KxGhc+9CS2SEYK1EepYoeavyuB39AU2hKGUA9FlHTyCG1cgnIhFC
/Soq6o2GI3rdfXqCbJtjRz8tpyllBsHlJd8+AEIhP7ptmrWhTxJ7F8//S5ecwb6sj5iCLeYJ9mxC
5amP6RIwQ16MKxUe3W8uR+I33lxWGUXBrRqGQ3ZkStIhkdVGQgm6FzhYFWA8mnwCalDduNS9RL5K
hcqeS/8sAWDpvIzmbZ1FQbFFVyky92DnASU20/tp+Sf88/73R/ndJBsH/uEMEOFIOg1i3a8z/b3B
W4VzW8+Rl7qSFYIc/gy8DV/tlcCxP3ZCCIjbm9Xy32Xze5fN/beljrTcQlE5p7IOCwmvME3uN7sz
8Am3zGmA+z+kmwOZaOQkl3Ln7epgq4sqzvVvEbCbh51a06W2eObh2oc3aeakkBQwMGzUoVqPpESC
QQ3ma9ECompGcHGSF9Y0D2k2l19ZQ61nXE4diUm74DH5RflGTCIBVbp2HDRcWFytzQOT0s9ww3Fa
Mj9BDV97J3l1y1fLONg4V5heTdPvtkAnt02zK9Or0CZF+aCcNoTMIswaF/ZAwnfkWiU9P9CfI4lt
HrMlS8GSyLzakBEF1GY/ZcS1GZJ6fpO5z4HMYclhS1uW3JCZVJtOnXBPmzBwbfmhrXJ/c4235I7q
IjnFnzNMLHiUK3geAY1n7QmlLAK1IbSFdPohtH7ii1vGdTm77c7aDobZ6tRmE0iHjGojvWDEmUvI
v1jPOHXuvV8WzWp/I5VLYZxo48eW7jQL1plILbJ4K5Rr5Nmyr6lCicVQ/P9O809/amI+lg8slpoQ
95WFQnCa7CD+oAp3hUg+KRJWnZzqWW22ROx/EqsDVYHJiHVPpJuqJZHjgpbhv3Cd5m+PXNuitdmR
/y93VaG+Po16h5I2TFQHVAf0XDnwZsFG4kMQDv4wHm8J34G5ktNpPAfD09bBCOgWnQS1QuC0NtUE
7ovz8kiGQeWoVTqDag8JfEF1X+MkfoIsa9UIlZq+kt4M/CHMdaBWTuj0RPqhPHkNhBN1D79yJmBy
hiOchGuCI2KcEZlLMRHytE2BIx6aZ6SoYNynpX8moRmqKj//a7+i4gsfGXFDd1+inIwLlGXT7itO
miSswIg/od+4NEbk6hoM5tmu25pslkQe45jrB/k8IEstSPAlANH4MWa3aT6xePew+HDRdiIU23Mg
ptOJX2Q414KZblzCzcS01+gDkBP1Ect4/k0qQXG5N6Bu4R8ppdpKWJKCNsSXy4pXwyGPNqut/akp
/4lwzEinMLtJAiZXQoZAyHdCD9PwtYW6cMw7mEcMovyCKUssry9bFKLnQ9t7jEXfaer/u14xVT/7
lpvezUOVVa44wUrsd24/nwz6lusPpwAV8z06toD2WCrVWtTjcI7iqA8MiNAjWxiPq+eq4I2rJrdV
9FRWZ9lGW5gvm1Shxzu4GwY/wEHzWTjTdxaOIGGKmTTPbn64B7HFEHnhf79DilL9T1u+Lwj/fp3N
n7MGEDUTvSzNyDpM2rorEOVDbnmqr1wIwLObmO8Uh4cbjuRgu7Xsffzxy3ZqjMOctdsf7wnTDrnI
iGizGApSgC8VYUo65MCPe1DnOQHrpV71WfsxjAV9opq/adl3Z86zb7Ou+EtvSa7a43jXBwrTUGJs
sZNsmUmVFgmZcSOOtTKcIspHvyH38qWMkNyqvYx2XK9Dk9ZQaASkJx5+ZvyWiDDiDmrMrDC9D0kv
JRUUOd9/E23W4u3qtNfFG6lFzTtW8QRR9OBwSKy2Ya5LTOll8vmnL3RvZEx8I2NtIC3dWFLIQG97
OQleq3Oc3dEMTnCWcdMJKBti9LpOmcH0WMRnPuBVETQw6Kyk/VDiZduv0GF/EBD4if9eObA87IHn
6WGIoCM6G4ltCDyPNNhcX3QcAe/A0D3i+WoSV0b2VoVSOZBnsfUnHI00XTKx8PEPIOhHa7TLWsXC
O+qjSmQZ+xQMXPHMPOj1G4Aq7SYXWmqUU3/QE3Ocx/J483I935jQ8+9bnQxJo9fz3m8fNbr6Cwvs
o9+7gRvp1WmtuKF30AV+wqOaSK/RySIMseSel4fHxjcLjOTOEehdPVvG57rGytHqM0sOoZFVI/sb
dzCY6dVV7tT1ZHBhHhTvwXU5DQL5C22KOc2dS9eiKzeS0gYOySMAR5b5052nb6FdP6jQ7bnOqcWg
vJ3T35c3uWhOAhUNBaDWrvFWAbUpcjKZBXcpxoTX3d81L00zetjPm8Dcu5kiKHwZBRL466DpdEO4
CnrK2/3SjP2isOqLpyjY2p6RBDbBuPGUsWWT53HmixpaScor/KuIbpZpBIkIBFzJea7V74IeVmDZ
TzRELnNCGxb6rQhFcMQfp/oAHZHvGaGirSiH+sEA0tyLbLF8/fpSn/TqxOT7/x26IGmFtLfPioG3
Iwc3k1LPepRjGw+q+IS+jseCKuMpYQbT0bET+mK9h2E66CYmqHsyRuXScufX6FGI7Txz77+ssZaT
HPE4RQXA817hcaQ881RwEPm6UvsCd9wqM/wWp/NUGd0RlF09lPhmrxVhnVV8Gc61meondo/uZI5T
0I87ioIGd37fmHBfMkyaqhjlPDiFWjlUpSQbFLdhY0xftPxweIQy69t18JQh0qIea5q0rDX3qGTu
bUGqs8IpsnOYfO2dQPcLKogOAkRZUhjKhQHFh3XIj8i8exNW/dxdSpgnjV0si25kFlAir3brCr9E
0M0V3TYnn4Xb6s+D73Ef/qQILF3VnjmWtrmy4fRnZfGpBTKvya70mazmile7DoAUOIo/JiNxL1fk
92b3maMm2rGOF1um54JXfWUucmAY+jfhtLNbEgO9/EJiv3xx312mJ6nT1du/yv4iPUeDAY02/IgF
JfLeHu5qbX4gBQ09pbkkRF95Y68qXNsE+/CPUeKusqAkWLPXEcqFWSu/eFo8C//cDAqjkO6CWx0+
H+H0vBk3jKRiFgXbc600hiq+qGfYtO1P0owyQC5AkLAVECaofAeINp1cKPO98GgByYJYs2Z8qNtW
tWNqK47O77sWQ0M0h6Cs/tLuNP1+LenNaJe/0zwmQm/CO1sLjFRH5zOBnVVN1Xeb8DM5a/lD30jt
HVOC4bBL/rfcjh6R2wRw4qyj89jC2xBuBwzmAxaLxGVYcDUxU84q4CrUts+9cifnDck/pBvx1Kcp
NxtTkSOY5WCj9hfp8JeT6xBkLp0BASdOD/qm68FAWIfzg5L/mEysOTNEdkFRIDOuXzXKWOHbrqAJ
1NyR9jLoXEWtn9Gh614ESpkmv29kQGYApIDtObWwWOf5CamZHJYfOSSnfU5zzC7C9kYX3KUIzpAw
8HnSGOeJNrKO3xYJIptqy66c7+lSfvExL/X2vRWqmy7C2JpEWdjEgWnFQrSW6DqWeu8z2ON4cTL8
BhUtRULIIWSyXCdP+uGXwWILeNQ1EcqiXe7xoFLr1sEBEAEuStKMtQEuNbeuZoSdgWIVz4qVcqB9
bdaQx9yddHzJClzbW6vgNB3duRa3VuVVOWU1174oA7SqV8HF5pw1X88S3mbvJSVNCTJnF7eMgHsT
wyPmQgAOrkM7Vw0VEVOIrzuyYn3GcveCXMEzlvpSskMcmkdzet2RmQvMjh3q78m+m29bET/Jcn02
tZBizNgogC1k6Li6+TgGv/RA6nsM7SAWoCTcyj/Vkm2zfvHstCh+weCHL4wQvA8mXvnmNGm+XSeT
n4K0dOyS7lRy/AQLwrgVHu7fAepSo+YMokb1OO7iZKmp283OgNKpT8KiRkPvnsp9V4Pr15aYu6ZW
qZz7DbPYhMrnnDsA+f9zmkT+hoG01bJqCpDmDICyOfKMSZBdc5FKbsrK6e7oNkQ4BjVDIoPerPZy
18yqiUKl75swVP4l6SfsFam+w0QtIS/Qg3xP8hph0zmBDVTjHpYka6yBvobOouUkYgsK8nyY39g0
HrXZRG6BE8HeFMePRBfTGwfvY/0ulwSD6MRFts9+xJBXwYvO88vVk/eGNVkWA7VCWLZWuiP6dOyb
9wI/mEoow/YCqMR9JTjYZ9W3H7P0rTAaEjRY6ra4slQgw9husdTy7RwosLBwW90zS4fX0V+yD0rG
fN2HqyaDDckCUiJNof+BCYL4m6cRtwgYDtXAAN0ZfOIh2qjWU3H/lnq1W6Ktbo5ltuGZ1Q4RiAVp
1bwU/BpBQ2/bFT9jlNmBYNW/b2REzk1Qt0TqtmQijms2Z/Nq7gzd9/arUiY6XrooOdv5fZ5OGyUC
UJLn1Qc7TpubV3NWB6zkfiLEIz7FcDjUwtvg5bWy7GWKHIXhNDWum/dvyBFczINyj9tg0F3UF0ey
pEO/MYCudnabwAqgBl2U2maSWf2vzs8BTIBRwGHp+VFgcPJoaepupuKh5aX37CFozhmPkT40KJ65
VqWZuMaRVf2xTsmR1nIPJoWyaKHPxtGvNnH/2RjGJvXUB9cg9YQ0FT0vkmeSPonRfLmA2jwqAzcG
7OMLcbmzq/LoDTTsJjt0NEUCiZ3ZVcIEnpdVf8oykr7Pnnhd4Cd6umBj1FALKbDDHhTsLpnukhvA
8SnQNVeO2Wk2xK+yfTBPn8a4bbme7ou1V9eauntHwrZy5+a+LBU4XqCr5ylXw/KYhFIuaYngGJj8
ToAr9niZM8cSwGP1YEp89OsaBRtukO66uwqzYZkHhoqnv33bX3SmH856zZXj2DNwimCtIQNuMaTe
DTaGiHr94Ke93Kf9miwqZCqrE6xHHl/sbGeOyCQda4XogrmaCuUeA3Yps1Lg6Pz932XFflodclyv
UNrBWhDelG7eLqqW/KxSvu6x3R2/yaYccG/dY4RWrCluist9WRY5qHAz3HZbbpj/U/gxtWPIi0ef
GlQNoVAi4ZVVJGp5wtdyQIy5UzZ4rIMtAV4E0/ejWW7dHlSVQ6Mj+HesI3AK6R83FHz/vGZjvEZ2
Q1EE5m+CVL0856IJuPOkQ2fFKpzqr1k1w43vFOACdhOafCE4/ove+YfDW7nO1TmeU1/63WP3pWqW
KXq4CIKXir53zu02C50o1ErWWnfBE5P9ZMg0vJJTbO/hJwbD7+VnqgVTZ3/SNgS/83CFPmoVyOM1
1doYYxYtfOSpoxzgtxVIKHoqn8Zo+HfGu2T3vEgURSTcbcDw1KnwoRGbhsdawFyRMU8NlwCzIct+
yornss/Y66Eny0XyuphBFwXQXBPWtzxSEOOjiXZkd/WVHdjDtqlYn8VEQUWgqEVWmR3kNtJ5bWUJ
1iydA1MNfCNi5lU+DHbTgMtkVZbGPTLhXLUJjF7zuI1pqFQHdf3kZwPjfogrhI+xHV6a9Dyuo9O1
RZd6I+1Q8n+3KyVKffMBDHz7jhKpaO8nZwaThYTfNAdFoaRMH7rbau1DoWxVgMQOtKaUrrEBntlS
6v5846U9TUO41FTaP+oR6/gIIQeNWKyFLeUcHvyfeL2FBAeXyncg4UKh5DLB0oFnFy+G1B3UhPOU
JR3a7rlJPxPWIoXRzQWJLQVTgtIqE9GRGQXNosO9VE+sUQz7ZGlcqDv+Q6SvmKs1eVsWBrTJuCtB
l8vsROAyaa4kK7s7w5uTk7esbGULXmua35piAs0adSdYQSshuCcBCPL5KlIILW/SEv4zgjk2De+o
e5Wua0xYA/OQsRhfemCmmqpD7g/sJnuUgfbwk9EE7Ncf/ZDlLf0zQ1LSyxeIFu4TSKALyWQzm+pl
QWgjQ1cQVv1pGh6y/TfOPCvmdnA1JI4J1sTaar1+kDClwn4hSjHw+iz2h2gtUVD9svK+GJpbRfit
lDQ8TN3GIWRRYq9brsm8q/POpW979j8W2Lw28kstk3tvbQvvmoZO/QOPS3Ggv5jcimXXiETpbGSt
2e28z1oLhCO4SQWia+wWBQc/kioHkunCSBSk2KJdP7RWzIAfNzzJOqWEjCRHEP5NsnLvP6N9ZDrQ
3Nyn1mt4k7Y0CiLtx9s5eCtHTzgVlmu1WkMRGkk8vhy74KSaz9Nx1IqgPlTxP+X1DwM6mZMKKmRR
Rs2V60i51hTorHWt7a6Ff04wp8KGJF3nyR6Hr+OGFdMpYLyVLGboLxKMHWnSrwEv3koxlC5QVUzr
xl6v+HFSiEzxyj2AnC1HmY+LjPL5wCVkl2mgGqI8TU7bGIgQSk9DFkFFI4xOuR7/9zyJyXp3AFlT
z/isLGFyixelQeQf/xXGn5dg2gAToSgNgU+G7QAZ8U+8JJf8JeDDODUTYq4/MhQfYbrmFlZARqYz
j8H7wyFZ/tsz+scJwar/i7N4cafi+9OjZkmwiXzxwZPT5QJI8lvZkFb0j39pHuMFDdXkYps0rqOH
PyunnA/WjiBrZkg8qfaH7xCY4m6BMsSBb55IY/zAM6VuNOqpWPTypHRY9IUGMRemEEPhoE+jqEzr
d0TzIyAI8EQuvwr7QTf3dNbq79/bP5Ko37uZYDcadHoHYyAeFXVtn5y0/tfbcr6y/A1Xese4BC06
0fdGQ3uMMONcRqur5tYW3OPfHUa8Tsb/NvA+UgBCNbNEfQukjmFfqu9iMFklVvt/4u092B9NDX08
aMF/6cDKHRVb79ktlGmk616cwP5iOb12fY1oXEtrQaNpSiTVukg1HFtNXdoav19VyfHVhAOOmsK6
dfvHvcrlwlTCjHTOx2jgj7wscWVdRznlBuMLoIaTTngyW4WUmiFpeWaX1o2mko207ypBIbDOpdIU
PlVEKDcPYKG8b3L4ULsHsa/LLs3KX7mGDHZAxLuhOba3aZbj5y2VdH53NSljD1WXfeHrEO3RKAJI
+JwUiEISQxDo2ad5IENSzV/jGWDteyY3UQwao0uit9OON8YHa9i0x7AGFSqya9VBF2q7ajegUAKK
JeYnnY5oy2hUm/w/mYjDFzgl3QMNd+JdkCLgqUVh+fLTJ5Ce2/VCPwkCmRWGwcXAnS7PsAzQtGnZ
WUBrz1PlwTnGaulrQeDY7uKEm8jngMvBjYIcXZPo9EPlKzZCJ6CV5OnBjqLG85p0r+9TsHGAcRyO
3M0UgJABuExfG9tbwPsbrKbKiVl2vdTqXoW8UeIm8XhXtf6laRADxEpW14ABlu7mYrPTFr8twXWy
NvbJPUuGZqHIAnZh2WmovdfhE6bi03V1aBgazWlqwkKrwaeklJWSVSytoIuyYZVVe0/gsM1rZkDY
Yp1u9PmchEtpB7Nq4mnI4PXhCFr9M4794PAWmaKELeavmqNTmLP+cgaG/EYGpHFyQpfqF4tcNnIZ
5bRZYmbSHMHtIR1DbW5lL8SSwWAqDRWLS5oMW54Li+jksF4aYWbzfHmXTwSIwLb6HdzHPZNnfZ5a
8aqGxs6we44lEWaCCVyXCOGgAJkqDyk6qMDfVVKrwt4PTcNp9JuB5W/LBuajgYwGTt7qK+CaanYL
kU2HAPYwQjwgRvo/DxsyZLX6/XX8R6v+CVW/q8bde+7CuwXOYE1vv30kBMsgCqskWjJNAT/p7dzT
WtAzRLCrZIunDmgChPK0ZnANvLLCJtMB9EFrtUQFUFKldBFNjKs1lEaPyX5uS/JAxpSvzdDrSmbF
dU7Kemrlkf48MVcQjORJo5YCM8aZmWmu1Ya52CiM3k5cVZhlTey68/rp/dMMksOXMzHFD1WycZow
Z7z6hB3lr91/1sBYB3O7RquNrvkyLv9dy/w8po9rCDKA+XiVoDEuCgXqSaaEFu/ZF+/UBuS7zxSb
P5HN3MvXTyiaaK9ZzdDwtCn8qZxjI3a7w+IYLgo0IS+Or90opfQizsW3sKVbaInQ3HsjpA66mAY1
Dys/ES49RSZvCHHyzI+QF0M3W066qEXkBp3Llm41Qv4Lk2k4/udZVQyI3glEbxYkGMlJnN4gV2ul
+U8kJQcB8vlu0ui6BFtgjB50At932X8CIwOCBImAM20dzUd0UZUDV6VrP1P1/TTU/7sZ/pRgvbCT
GC48aZIFCbrXE9KxzoM9LsIWkkfMehoktexnTfTK49/K5H0YwYVkIUnl0Z0Cv4xfj62SddI6FQln
IeQvMHBYMImb3AdXKuhUiJI6XolCjRmcpbO94r9QWkhltzUDmyJg5Jz8W9Sx1oPbvP03LuqGdFXP
gOBWN6urQImDGkZxWOCwYUIRa1LmnJzI0Zwl0sqlbj0Mq9v5IeXbYwfM4GRXvzgTEsUKrQeWIad7
PVSqbGv3hqYyY1DmPB3HHVfmqLmQAS5T4L6Nah3QIxayQu+3VbFLP5mZBmji7O+qT60P6X89Hs53
CogHyosExyeyVeHBCnm/aR/2uwdnFHnsBV4+oJ+Z/4Dv4sL3RRpK7AEjurkX7X06fCnXrQ9/TEm0
HAUzTp0Yax1Soh/jkd+LT2AhwKmg1yVJycHQzCcliby5wtBi+QPD7LL7GF0O8O5w+F8a0EIkmSNB
H4P7mDJpjrq6wNXSlPWF/fO9GS37CHJAFG2t1yz4Ufj90OtBayKlEJWJuubazTOHbc/HEBCjRN2J
BQxwNf/OGwHbjwDbztZ5mKYFW2nJxga66dVp4zsWyA+abN0r+Ap+F1VrV71jBXP1nzQMahrgMOjq
PxUSZRoOYopR+q26+vySFtKXPtR2EFFKJI79XJOdQb3AJ9jCl7tM0xJMXMmhn7aOo7Nraf6BS9RX
XciM+8ZxdeWSRw==
`protect end_protected

