

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QHA3Ex+CmcwhHYj/Cu3wGvj9D2Oh5X/PuqFEaH2NXNQZh8T+UDvbmRy04SPk/2ZNtGxTEFpvVC+A
OCZnLDmVBA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EpCFyIVFCjVsV8JAoVIvFxgMicPOE+gA797pZe0ptQ+JWzBRfe+ko7I0AJCcVXyK67/23E/Rmn28
26K0nfbqlZMWRo08GQzdo2Pvg+0zdb5xynhVYesyBJF810yAmWPUXibisA0Uz4hy5us4urGRvXui
1VlpuDGRFz8HEMlbkMQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
H91qDFpDLhLKyu2zO0jS/sr50G0AneZOioO9iB+qoJcFLnwgo0vpwwtqzJX6wbDVN15cu+R/IWxt
dEt2vBf8d1vLuMo7BshJZtbUM8fTrhTZcFoSdUQSe1qC2oLTy/DpceJuEMWuDApMg7w81zUOWyVZ
l0ZQx93l6uEMApiR26abzikEl3AMNYgld7204pP+LGkuQpEm5BNdhJ2R1igYEH2SLr9PoNXl6Ybr
Jw60dHycu/SF1aZZvyjj/k0RqWzkWo9OF2bMBdwweatK0hL4Za0tR1dkbQIVANMFXr81aRAsb+LC
ySA4CauSi00Vi5Uc9EthY+ZLgX5Ay9HkzjDp/A==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UQgJtyN6NYDXy0tjNwGtkb8soUmLxZJVzWlNkhMS/C4JfTEXUPg+A6vy121UgFOz3JMSNyezviZf
Mfex2hTID+DH3Y/f+mS9lvkRe2ugr1UrbCWMuo61hHhoeO3FlSVy5OojiRVr0pFZAlcHpyRyAMDC
2ubNAtCqnKhJ4O0W2nXkasQr4eFt+GOK6JSg9BIu0PcXYnr8Z96U14IqU8qoaCFnjmOffa4iFoKt
fCItpLPWXVs7vpK32UsZ6CdWATv1DRVa7rvpoKAYhB3pTdLEGiZwBFovoFut6DljSNKFNe31ZoBh
ZvEnbvlCLpTfwwRuxQIxsF7NsbghGxInSwNF7w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GLlPz8clXjBHUAybAGhYboHKfTw7ps5cfHItKbfGW0Maog/3BI94ghpter+alXbAkH+8KTGFy2Ck
42pN270kZeA0uP8+FP5FX9Hdxx1rjSJSYnLaETC59zrF0zNRHR2eUpWdzjk3Q0IyjEcI0hzDMWpB
BTUA2W+6VKIt7CwOChCNccifqqqM2/lE7U6SRri20DGmnKYCeA4SLYKMVgbYiwIQ1WpXXJqIDpo1
bsC7dc9a1YP5bjwk8u1LIhPncODSxREUNUwGR1Xb9he8Nu6GvsazhQaKR+ckU3zv9ioeFohkv8YC
6S+WxXXst2ppErBUJHaQ9VRsWjop1VaIGfPf6Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NOuQSwyLor/NCRAPbb+hLF/fWkzD7blUj5CmRCbO6PxyE6eUcw2hCJ3syd0WNFx3AwuOr2lG8SgF
2djEMbP+862p4gxkXmmNOf7tGqVDHgC/fgmOIsxfkZ95hvRAcEvi1RVx++fS0h6KGuC39yN9BrTt
nmZ8JjVs3v/ky9THrn4=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BP26diD8XpcagtcJpVVq+RbpugiTQYYy381rJIl+lewz0g2oe3rZrSn4SemKHDAtULgIN2oNIFYj
pWqaeK5KLTW0n4xvkxIsB7rciQ726nTjcRddBUmvF25tkhA3Y3UhvL2S3bElyqF4lCnStpJABIFq
XT3R+Lyq40nBC3EXTPszZosjTkHBl3uO8EFhwXxLaoSimXXGgappLzUn6dp03J+zr78NjVyMcx18
lwiud2D8+5QyO+QXigVTSDyD/Zd1vaDmZ5CVwxsypJWCKZ2A3qx4HCL5RoXw/1eLwI03EXKqEgVE
P4uFzHRwLGNImIZpDLhj8SnU8I0lOUFiGGuDRg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 132672)
`protect data_block
5iNVtA5/9aeubTWaY5BFEvS91wnCopFj//rR/nzbiwBkcP8CbYR+zmqaXLh/3LgRxMGwE8gyHk25
YLb4jMbas+6BwaP6LIxBAOaEsaLc5ka8B1bwTA9ZlxnatYHqab8/d5zVU1e7dbpSCupAgauRyL6+
6dn9t195j/60XIf7btBwuJ6ovYUOviYGn63wV0PY5BMCNHuw+y3yJq1JzKvoIKjtwJ1KCZrraS0j
nDcRN1Z9PNw7IKpiBlkNV5uiWBtOYodMKCwYV4mCiarRf+Fkr6SjL8OO68s6TIYVR+L3AxUSrk9R
3v1147B8VCqKM/1omBmaYGy16a7I18Eh890vxePfnv4QvYqeGJtiwurtWnW4aPwZ3etlySJJ/LQv
rKMw0VdUdFLpaxoapM0J0ypYPw0pMJ3MmQrBcyfJ4FSLTZO5kFZd1abU15VeVKDFusRyA+VRxFHU
C9ryQv3qz0Mx+rWH03BCJbLNlhtYs0rOnYdwTK0KNb/zg4A62wZoV2IPGz/Yp+3OOoN4Y2p6TzId
TRVCbUBvD8nBW5ukNSwJZHSSxkba5oPEkdgaYDk7Jh4Qp25E8P0QumXRg+VwxI/cI7qAwFishMBU
jpyrGRsSJxoOD/EgTBpi8IE/qLjHVZ6MhLzaX9R/tOEGPyd6UfWTlZ6Lv4br5GacOgfiPBvMAkwB
8TPqA58Rhtly25zTROmuBt+EmdChT6+Jb2zGO25YXqnEX20TwbrRspN+k5IPalDs/e2RWkaoi5jJ
VnVDDfBK8Iwe0KVIh9Rd1B3zZazl+wC2E70OR2Q4xNMDteR5YMddt/8A8EPaZOfa2FzV5fMuqEb+
Qnqs5mo8JqtrUG2luJq7mUa/8O2dyTrYlw3cscHaKu8vHXJXqu8nLQ5qzj9rMRUQdIbLPhQ6Qgvm
f9Za2vyqhN1k3bgSTkwMDt0C/Lijqk+ipR7b7vwb1xhKlEXBRvl0O5H7Izwv/uFCBiTTMP4RlL2j
RNZThdVGQBoGwwPmuD4rkqm9j2iGnND1a6LnHZ7N+A2tPEmKUBtHoRbPUy/bK25hwy1CmOsC/ZmV
qAd3xKvOzykRxtYZZVwGkMiNFdf9ennS9cuyn8YuFJf8ecuMH9O8WBL/N/ck9UJB4/r1s3LXOS9d
fM7KZHiL9GNoX0+EPHMAEGozjpekhXF27T/OOTpgsa0JS18hRV5zvUFEyHdnZIqaSpbVB8OiQJeg
a2ZZ8Fm1q94KKsQ5cHzTQnZvkEL8vIprlPjewRZnNai8PGt4N/PGObnJ8ZknL7syT2BAS7xuDuBZ
Uyd0FXLfHFR4uOFi0J9cQuRciyK7c2MbzWD5KyFHcS3dUzJZgg0BSOnSZLdoyttbecuZetrfqwHH
JpAw+86fdJVG6IuEOX5WuRoGuljQ3iIjQ37PKJTIIQbHjvRSFf7qVr5JN1jazW5DgLMs12axtWYG
s/+X+aEuRkgfkR6uXLGG8vHOdfIEnJHaypCJ4Z8rcLEWFf8E0Q9EZ2xXnHIYr/fiJWOmcAUSuVg5
6CYCBi5eZRcaM7DEciYkvoTu2b/XfTqPDSDML62l+nyBeEDu+U0zzKR59VHQcPq/ChouAsERyM0n
XhTaiczaTj4ala4bsW7CSbFsHNDcI/aKtWsTJHQuE4KwbXm6GfOx46V8QqtEaw9artU4aF42Qhgi
nhDxUpaZIPKVEk30G/U/ExRPShqlbIadQJMLAHlJQJ9xEJSt42Egz9Q2g/G1Pmd8/ynwRwgbcN8U
rOHKtvrrXhaN1aYd7T2iOrClLdmJQiExYXKmLNDhSzg2RW4gnHJGqpYFp8nc9AwUu9C0UxbiKWq7
Mj7sAAbJJK2ajVvjN4Q6fOetFyL+HdarcHetzFtwwV4UztNMXukjpob4hxdybVOvQpy6m01Do0ya
RqQsGwZfcHATLGEQuIqaLUz+P5FA6h9lBwm76ug9abwhYCrgs1gHkx2vMGpp5TBgFu/k0s/trZY9
S4e2Fe4KE7Ouv77YRR88iIKiyQeov888vJo+vTBoExJ6iJwF4VQZGb04mvKxYI223E62GNqIlpzg
3yyUHrpzosS15iUzmDi1fcQ/braKKnZWDBqxKOSD2bF6OOfh7NkkxAR40WegEpdj9ELQqC8A3ibu
/7hhWGkj09RV/CoOwrPoNjKxmjo+wkacM0NTBp+Nn82KJNdXBRa14MzM/so2E+Rd5juIjPVrmNtW
lyOHm5ZcI4ZvLriA8Ttedjy54B+XxPhwq/D/J5MC3JLQ/sCwWOqg3RG10GBdTAHv9csvWgEBp73e
T/C9+twyQOU4SkdByI1oL00MDoePuz7xHHnLR1jyekiReyMmU6i6u/84m6FhYztnw5NCMocvh0MJ
gdNffy9Iaf6KKuT5I04/QUVW875iBHYCjSffrgnnLy/w3g78YqDecZxY64Hk8Tv4QEfVpuEdC8v8
r2byv8gtUG0qZSKv1uAnPVSPV3m4nYtfRAD/R7aFObOQB/FzVJh5NkXO5FsfjNz5g/QC0HasOVfI
76cTegrWwckMbsoGbX5sPXpMndXDZWFvFrD6DDEvnKmwgAUaJRdgEBusaFYS7gbJ85AosvjA162Q
tjEBpOUn12OCTpiBOpatZzUWzKxibQTeAn7WSvBS6kPpNpS1+SnscDZoZU/uv60lTG48+ugxNyiy
IcnXThYcvQVXirL/GOVZMSjZKJRLcoD0rSKQRU6QMLy6U6jlXCfBbLM4nsBR2jbW+hu4jwIz1Lxm
aNo+I5u/1HXXM81cqRHbNtWZ7JJm+v+y0av3rpHkxTDVPG/BbWq845ezKbm2+Dt404JWt4xbu4Dt
XrPmy+gEGMQ3kpfR+xWHy65XNdpG4mdecE12vFEaa4RBKgcARyhBoxJvI2/NlN9tSTPzMwhZEbGQ
xwDQQPEM6g6inmdIzJ99uSTAJOtlB6Qf0l+XutGpLTiGZTlmDzCw+KgUTBA3Qxghwcqu0JlATG1G
WCM2CONIEtQXpA75qpRt2BydN/kWmlLY2aT3eRJBLIwDYfWr5qrGRs6ZtP2IOBXJvE9SN/KyIWBq
RXinJ3eWIAifvTodX1eDMXHioBZdcNkuRgQYwsDN7Ayq2YjiNPdTwXIvd1MklmmWkk6XNCnluyRv
iN6uzYYzbGzFEeHyMjItUHnkkHgEMdJOB39yUn3U9zMItpWihYRNiCbmP48uxKInZmXD2cYf9oi2
8t8vRPUKRHfaVv27Zz2TzVvNxh1+6l6xDE0qrbI26w2Shv9wqN43W0E5YPypErxApTHZtxhFr77f
0c/5Gfey/DmT5b66T8SgiZ1r1r7DidlYfZWDyhEUlxb3j+Qf2HwArA4ZOGDARueD+XowLIJ4wLoo
gfHBdIJzJ/KawKZ7nzx8O9nKaRT+DT03SEOqsFcr9iDXQYStZKoAJ1EQLeP1iLXjMk3YuOpADJD4
NxXUXiv7QRzAb6ujtQwGm+GWrsiTr+NlaKjlgNKtwW/L/JYJatsie+XNVy4fsaNmdrYXbP/zcZh2
1wZrqgVR2NGLj+GMrOZb2eVtIZSyMrnzUKTAyrfhcIQQAFawQzh6FgCG2t6V0Dv6AisEJccZwI25
uJnoULJDepL2y+VCp+P1XyZiHUzt8K1jh6/MSR6JmCJwyZZgpdc2QELp+bof0GYjRXxWZJqlNgVM
64zkVRxFaWRtwUiciuVwS0okHKk1/b7vou38iIunA8XmYCyVR5b5qtDkzIrb2T1gUTCFDSdo+xxV
DNC1Gpk+BnpnKgi61TKatpNANz3MG6LkVwVYY8L6d+Ex2RqXPiRvCeBBmxODMKfocWmPEBDIrglR
c6G0foY9QqC+X6K9Ig+vEnRbHyZPMaiZYZRGXBpWBKYkNStcsSeYIC+u01Vue3crHnXEiP24WLKs
fHiIUBw5RScVQQ6ptJcspD6t+aP1DxpkylEnEsr+aBFNgsoIfWJE1g2D7zO5UQCMIjkYkwx5chgf
yLkBldI/mmyM2Kdw2iDmt11Z0fc1aC0tW51X/sfa+QPwmIrERb6ZEJo5LZXve/Iy1E2yOmkJPnYn
gy/27GPo/ylgloaB4s8bA0+oJWROK2rb7N1KGOhJE3HCS0qiydQMQDV6X11wW0Uqqpjwo1Y1kBBj
T/xIZjAb4dF0nsrOMWtWUehUsE2v9fYW+d2nRjP3pqbmgy5u8CgHYlSv9/+LnyBuOKtP4zmg6cb9
blP8cmYTzaBNBHX/fbDh1xhOg7UN1pLg+EyS4zDN3sq2N6HHhBCABNsABIho/+JLIMkzE5dXNu/9
p/R74VgNBsD/PYLfI2gAULTAaEoMDewpmfMB064TD+lV32WEiwMowcyeK5tljV3HJ2xz8dlBHlIg
0BS1u0DO8R+rBM8HOn1A/stqlodnlbWUWQQ0CoNseNTHjUOLb14JKcV71ry7g0d1C+CBfe8pfD9Z
Ylh88Z/lpKJ7luuRZ1OYlqc+GnOq0MqcLF5SDPDOL1OJFyU80E3r245b80zz3rDNQ9Jg/lQ1xc2k
PsLshetujFWiuaWQkdLqLFoanilteb1kQLb3WAJItCahLaIkQr1tGOIzV9VQzHA7tAvzw56mgTFG
6cSRlLPdFSSnC/B6FK9IvgR/XILT/bLqkYvZJ3uOYl2L3TfGGxRm8YgZarYOdFyUDvkPTV2DbqGM
MP6+H+RCLe4CM78mA8STDR9ZQM0R9zsceSjggdRt6+wrHqBfYEQtJbygqe+84mERBmMNgsupqfyF
yxqIOud1PUWcPsUXUSo7lfoIBvmBVLVZDZqmD0EcDdz9kv9t6DoKoAFt1HI6QQLF6AiNGIhQc3g7
//9/xcFjQMNPyssS/kMsoASWtIiehdUoJpu298SeNp5s/NlVVLlTAUMSJ72DeFIvv7ky6X28ip6h
1iNHEAqu4XThN1f+9hCtnE/mUDQSdxqZn9VLzYP9SDvxkR8R10k4uWPniz0DbYEtil5LbkrNXsJu
48uV4Bviwv5Cb6UYGuq9ATiiMHSavzsjMSn1tmz+7/Qmwc0/AP1FwUtewHyjXJALBzesZb8Z/Xxf
17x5gltEgCRlgcak6AHpZlywPxWFdesMT7rsX5yLwlpH+CrHsKyDPYzop+4UwMPcZFlt3XKAIVFJ
8xuDwIeFhfyNH2JwTZuLZd8Y5NDwlgyB7Aykq41dArTwU/KaC4Rmrt13y1vHbYeww5X1zk7zmdk3
3Hw2eqOOLZjRdiwYDhuVBZPHDt2qoijDmOD7LS/Q1rEweW739RuyFiDdKm1wsiuQBeXcF90qmJA2
TBYb2gTfwCGuLyRn0zpHiEG8hx5r85mjWzEfrK7v/pKIVoH8BOeh8IsvpGWBrySEj5TcPNy01ntF
az/liQnxGKQtCYSkaPuf5VuUUnkU1mpvVqbM8vWAIFSzcy0MmJTcbjXf2hxYm/OHSQhfv0Vq72eh
z3Uzvhx4OK81RKSglBvXPTk2qqIlulO3fbE6bK0VCXodBV8MvF3Bj9P/twT/YkOjqas5MZGbd3hK
Wvyi4N5nKioC01x+hXxDmHgZQS2NkwMovKf7h6mDNaqOWjAn/g+e+gBaNWGXXRmS3Hsb6n7VxSCP
1QxKdicUxdCh6QX9EnPRwhN9aNEYTF18nKQpiw+Z0zQbXVZAOr92yhZvNSBrfWJn/prgKzLZ9jrA
hVwNbeizcVkiuAasJu99GTqPsiuLmPpzgxW9+YoWNSdkk8FPQzlVc/pPjyQMZz5kNut4UvuWdpNF
w2gUh76z5u827J3rpY++hgeUj1kdCCTWe3pG00+SBM6Gri1tzPRmPYV0cSBP+oLSpQcIFD8fF+Yx
2neThtoffleS6Yl+XjZ+Mks88PJvtICE46VlPYjoxd9c/tFEmK0gMa3CMzivOv6B67wOKV81sCaM
M4ZZ/TFJb5BECh7xJKexC/2V9h5tal4fXAbnOtEtuYFvXU7GOYYU8YXNCZZnUnp4SsGYslAlc9pU
UhbIYcb8et9bA/og4KVwZilyM1QJGSpCgOu3yGlaZH6C4/LZZW/OsSidOOUId/ToyjDjL4dHmSiI
XMBZwBl8vuphvac53JXnctXNx7VnnyK0bg9vyWsU7hdZk4sqjp+thKiS0694SuNCtDnxlQY4x5iE
4xNIowEcpmX2yKWRIWEMXVV/nTNrs/ezdji/cKncdxUN+ewClvXHplMjuGexLzfxwcrC4fqWlZPp
c/b618dSqLiGNVuxRtGoLg54l9Or87LJoCWFoFyyjzO8b0gwtRMonVnR4mBYqxn9+yoVKKjfM0jR
Bk8+GCbb8bnBXC0NxJKS0FSXSiAT8VPHZAAf2pxv+C0XZOi5zBD6uPNr0JDAIufCFLsX/30S5cz2
BSbJYCbL2SZrRqyO6ivpKXDEu8HA3Va7q/gXwuhefICOl9is6JbUZuuG17Y6g9M031JkixSqLhR+
J/PXMR5s91wkXoe33/KwfkjyCWR38oSTYZVEX/CqfSZlgdIwGRdI2E/ZAmlDMXBnvLpeQh5xOW1r
XtiojR2RzWXWpIxvBHBQCzfP2ojafjhWmP8ewVeSIQeNr2LWsXM8qqy6lsWSdogiAe7sp/Es78Z/
ksX3u6EsTK8P7v7xhyS2fB7GWshaY3JRmD//Aast+VDMIj5RTrzsTLbGpOAcGCYuY4xnn3rGgNiz
eWkUxWeV/SDREEo7SKwwKN2o3NqHNLPY2BfofKfW3Gg/WHNR7mRRtsofkvAr+lnw0E1oZAkHbLdx
ioALJG/1IqsFSEhNCYx8w3xxheZjBznnf2IfooQ4YmovA1wmqRNucfwusq60eFhW0K3Sql0MxdZ0
lIFs/dd4w5lebFbfeqRjXN/6T2iNga5NpALygI8xcRMOaY4mx0xym2HPCgeeV5oiOwmZOmUGSddx
OtbeFZR5i0Gg7dHS6x8DXHvoUh/ga02uCFJL3Xm2GJ4mEJaey1tPLKpVz3KrOVGYArzCVFlScdeP
7gaSbmzPqOY3+eif/jYDz0DSV4H1o6Iuy3UG7OGyMNTtWahHIx09wicworuag9bHeYcjXk/G63rF
5YIigRRYb0Mroxiw5aqXSsFMa64x379QotFhxfXZlJwUATZ7FR24jjVKc4BxQgh2OpRlzk+Lw4RO
hWpkDu0CvAgf6aO7/91cuQ8qoc8guunU/mCrSGrc/1fzOt9H79pw7ebwUJTnuD7GkRzs13yjUBgK
wJ9TZ14TL5buzvvquSVykgdJ3m4UXnY9XPjEOUcy4Ys2GsYeMB5wU6i3aUy9X13YrBGD0L3Tb1Q5
Sq5Zp3G0vFwfBvOzJTrjCRRQ4R/dgTy37oeU+S5c41wXLTSSLxX6pFf6nF/745jHlUWofKomupIs
CckOA4xXRoSaRTKSr9S1u4zVQCyLMcfyArE8VX1FY7XiQEIWVerLis7IrQV0GWhYcopHTPdMDtfm
YrSKJMoFq7NDOkuxvQ3l2w4huaFo9kPI0CZ1DnbzsDBpjyYv8FEonq+x7Ru6w1IxtEJ7/9Li1VXW
UQy5oto6R2exeLi+KT5AYCQoeUiAi+gqpb+Y4/wy/ub0mWcneRWsdFxd7/4oU9ZZETLxzkcEYeur
Ob8lvI/0d6UHj7cjlZ5YoN0ShEY7RqYDwFWpD6rKQRVSjxFLTIEx/41pNNTaq/AB9HAZC2oRrKaY
E7blTt4HtELKd5QZ0uzx+oMIWqJ/NtfVsbpqwjJJ1P4gLiCZtVncI+4oJhr76vTFBU+IAqjOX4dq
RLWI6OPI5mQ4HM3zriRZ4I62O23MWrFME5JCJCqasEMdl7zTaF082/xLWwMc/AirYjF/HgYhmScb
sLTTSJWWEGWD3jDp0PVl560GN6WQ1UP4VPR4W7TD5PtOLs8exOPzpMsWTPy3S+BV8zpVTNK605kL
kxXz9Uo9w3tOsCz0Ivyfl5A2nMuj1l1+8yh+wxJXEEkzZMDuyWoFGHNIPyXpjWgWDcdvhUxfuepA
YikpOwhI6n2xbrNLYEMKztDv9ZVVCzDs9twFEckw/bI0nAvR9hCw5TkWYHSsDQ9uKBMvIUcxcROg
QY8QvJ3NHDExdcVjEp2EMd6dwZMPLe8Y1XeJ5yl8dC/WtbNUZCxuO3LUxr1Jl4OMhBzL+nMcMvWl
Y6oC+NcBin8/ciIdADz7NCxqqCVQRE41OCf4CEg5DQvl28Jc2kch3ypSlbzxmEH6xihVE2q7XpP8
kmHFxdn437LNszjqDyylvB16W6LFcayXw3sdwBq3nqQLXwttuelDkWWt7IwhIqtzZ0OOxKDkqYzQ
M+Fjazzb9fmxtEgpM9Nqkx/aGr/EHyktu9xLOBG2U0dRSvG4dCjzrf4rfwxoM6QFKwmiqqUovzKl
dsC5ovvY41cq04wJDtO5wRmrgQn9LBTCN4HAZhV+4iYmCQzreUQoHnVBtu6TILVp/wkfIC5vussY
Kb/qWwr3ydYXQ2mE8Ff8aZvtUHQSdIkCXA+ekq4paOFhQd3eg1sTrJ4WPzUH2YpLWTWm+9C3/qVC
ybTucVtQk3S8eav2GupBk3X1mkmAVuhAmCIohjO2wVugxaB1qe1kMcJnTGPa68ovgZ5QklP3DQWt
ydFP8cPxKJx3VRYUh7U0gwuSj3vk5FO2C4uoKMI2QtrKmJomvYlC4XvgG3xwiNLLT7Nn1ipXimVK
qgSpbxcsSJSzSg/V+tP6tHKctbqAL3EnS02qmBXXqT9dQQAW59kiaojP3/hOnxmEiwVceIzcMAZD
fS74059z0lXZb++XbD0a9QVqwTWI8o/klnW6eb6Uw+IjHvXfSOHFPiRCY5/1jozdmU0OINGi87uA
uxqTmdH4MX+CJJGhB+Z0z9q407PUlhCK7GOY548IedTes8fCr7XM/Np12VxGHEErbrGsbaLEShmW
+ry5JqyMF5O3EvaGMqLIyzofzLcvMBUM6YhhbjGofmudod73cqB/Wu4koVfelfapR7Oi++PWVz49
KpI9TMvHWtQ72GuFoH3A8Zq7IoaNkCrOqF325WxuWWIx5vWSrBzfaIUaNlcAc80/5TzJsxVYww+7
/tC6QLr+YgMC5U6gPOIOvs+WV1n7kW6iGUQ1NTyooMhJYqzIQG5L98yteIYl83Np9B+020ShcfD8
E5gpeYGjYEL3WM3Zhkf7iGgVrYo2RM7Aq0m1Ihp0HRw96PIvMTztZE8vKiIu/t12nZ9ni452LnRr
xQdOwLX4CxJA0649FAZ+RcK8T7Ae6nrJLrUF1w9R5t5ulIYy/MsaNCaVucP6H5jn0RXVNtMnzJCN
Ojq8qcR3Huqd17t0NjZFM6gGsloHrXmWdTGYIEN/+B+vSS1hfun+pmEZpo157mR9HfUgrPZVl3Sl
Rja02rbs9NCrXLgRz/3bLLgYfWANN68yRs3Q9j1645FN83iSVa0Ccb82AEI04Zzd1N/lx/7B2UNE
zAYlLWT9Y4lZrcclPDy4j8cFwcRmxuqtlt9/jvnRLiroTyGGqTpbrhQIu1H+TTt8v7JnZP383cYQ
vm0mFWR3UI6zlWktoCQAhosOLP+LxZkRE5FddHmoIp0tCqB2/Am8kXHndx2ugl9FQX8m68y9DbDt
OAc3BWVxO6Qs/uXlKFMjuzWEvx1VtgF+A/ZukgM3u4HS9WBU5KP9SKffMzcUJCgh7tEfiPg9/ZzO
qYOiq01Yrq3dPYjI23ct7NR+W+ZvkpitVHZuk0Iv+T4Ft1gnH5Tfp/hvyPsOvtdZ1Hz47k58XhZ6
xM5eH1Nsk/fKZK2xstfX8vsKnqiw5pwPx8uC7tMW5UI4bjA6JM7o77FWHaKXl7hCGUX7AtPUwKM7
yRRf6wQ0Y8OLy9rBD726OHz9xr/cT6nm7rQvLPadsikIy9yFZURGRWxcpedoPepAoxiw2PnWU0el
LhPGEOKBQ5NaMVDZctSUn82pyhykkEYFR1Fg52c/UOhJeG9w5IOTmA2DXCm0iSPlBHoMpwOETINX
o7USKKzGfXcX7+x+fP+WkEt80VgeKOUjocr6EhPUgT+nz2xbFlQJmQUT9nDmhDqRm0ToRUBGodK/
sUz2rvzbfnWlc1+0o0GIKQzFIiAI+xsKymJZB1lBi1j4vlwQM8QBJdtTHjb259UTBz2CMC5PQ9zd
z4cdxXD0YSp+LJ1vsdAn7ZVnBz9p42wAKhSspe4blpon/S/CLvIClQpjfPjmosDV/yndaCW1Kv9k
+ohfwKD0TwFMMtretNY0IBiPaNEanwwOK0mAs8GPEIL9ZGg2ZXJRSeZu1Ma76na++1J1hLIVzE9B
OuwYAq9Bn/tRWaMfR9CVX00qznvv4EbJitDxsHZRl9RPlHH2/qzU3+PFgK2+3O1xJe2/E4jNQ/WW
m1YrK/hEEnLucTm51felVJydXZUT2rtmGCNoDh7WC0lIaiS0prM68CKTuyYYb+DdPuWPU0DAvJbq
mz17JXKVm3MTEV/jJErCSdMaH5CbxZpJ9bmaklUUlGswgLj5BXFKN4tAxHY+1asY1sZ945kuYet7
44EIpBkeVC1n/wPnmzvBINC/iTy84xHCjGK08Ag6OZH9KXMo6j/hhs+AvGN5zLtfCrGkmNM7MKLY
yLJ22YpD5Mvcgx5iKUmPj+jz1IYOkB0u1ipRpIdwWF9AusqlL3WE2+FkaLwy8idlvSM3H2opyTCb
xANwlualjUTrbPUwyt/2sefgTeukiI/FzoUi8a5KrcXXEjSu40FW4u0+ZGKNQjWGSJ0YYF6Pw3rG
QLET/dwi/onAuOtlVrwE6wDQY0N7DVeXZcNnQ6K4E+PyZ/6cu5m58mMDfa9nq24Dy8DUNBcwhIVd
o5Q+yGYnLAZE2a0N5KC5xAoM1IrSOCchLFH/mA3qukpowhMF7n167AAVJByoKWbmNrhgsPwooWXp
RyEQjkkzeSBm4+ctno7rup4LAUtifk1+VgRUDatbO5oVLf0wdkYiB9sLjMlKmwcNLUe0fiHShDGY
peFcxLZR8vWuBki0Mwsm/iUttmEiE3XqaPMFBJHV4nMZt/+jjqUfh2dkF39C6brIe4lU9Wx52Oyf
Ejm/4syc06APtAVNufYFFk0zp3mrmoAJow1/UKf1O9eCvZ13O+Nnr50w2hJPCL1YtEDaR68zfTeP
/g3YU608avSBYKHuCRlDKQi+Vj2XKQ6V3KqQFb1MeD3FzYhcvXP1A6SIWXJZZ9bA7lK1b/JyU0M0
zjqQUlachlXB0l2AIgVP+8x2kUJouLLlWZmkmuGNDjJ0ZEyhaPnPnF+KMW/5Aec7Z7a1NEMeUAbq
1ET585XDKg6HSYkS5eRPlzpKSPGBNW7o5G53X88M7fBY2MU/U4TNPPUdI6Qg89MuOyHw0PaVyEBr
XHSDs0hgZLxWSWj0S+nqc00d+00LHv8djz/d140H1xikFHwpsPEFpM3mY63swfO+5KtDIla3wfkl
IzIE/igN/K7jEyhcmRlGg1p2Mht0eZDKKB+tJCcGQQNVpOQ2zZusCdmPvaaE3RN88AmK/txcbRQy
TVS21XieQ9R37Pzok9FGQYbQZJYeiwYySoCoWFBAssmZ3FKodI3gDxEakKnZ7EpJsw0EqAQ/yHHD
soo7MHOhRnd0qhofK+AUs2Q7wt8xgEmVl0ujXMNAbEacIaYd/wrH2ad0rBGgqFupNIKDEFXLqH38
KpUmSO8Y8A2pKtaTlRwo7HM9HxIVQIYAmgFLPC7YwV/hBJQwn3RxAOPMMULb3D5bSr4/WqfutumH
b7tIXmOrknd4/CpjVYNh5UJJ7Y2qryhDtWBJn+9TAOFQgylkhJqbkehl0UG6pw5esC9QCEbT0gdI
3dxjHyQPE4WH/asKfw5sboKML8bAX3aq8FlZYK8kmOBUMS4YV7UzTkKUGrIpU5+o+Ob7JfQ7dqX/
+bBNnDzFXNBsPOzRQyru0uJSzipMEAWyuacoNQfcdQGJ6aJJWHu+sWG0ZVRiUOwR1lxCgxKBmCqW
XFEImiaD0IlAuTfZhbYBbuIdi+W7T+Uhht+oTodZFntkqyLS4DnAPpd2O2FJj22qooFgmDYqH2Mv
/IoOs01JrBqsVUR4V0JSztRSI2A9NO/cLCjTjh+Izwmf8Ph6FHjqRr8ivXGenoOV3tgNtb7o5Wa5
FyZVLhxIWrHmuoyHOOQyGNYN/Nf7RnGJtdjKemKwvHziT1y3F0Zj/kvW7xSGYR/gdBC272NDDown
Cd+L1B5DD1PJ6FDiT/tosY0tmGVNfHzZH4wg7bdvRWRTvwn34TcjsyaVrLVdMzCP2SWpPBfprqcc
VodafjZ6wv4LC7Nzh2/73Chz4dpbwk1f3STsyQqYpws7yK2yUG/m1551zpMJXuRxEHXcjtA9cV3M
oPLzbx+4qNWxn/rMLthyCanktwL/ZXybYSAYE/TmmFxB8hK93e/DEL2wR40O+vz0EPLWjqEeaWvs
Dze+HSW4RCPKHFjw67hww76MlfT7qhchiO5AZcnY7GXbq1yXpOAnzk5XchKitG4w17fQqln/Ov99
UkkiHMW4HWNMRiTfJp0oWahPmBrGFzS3jpgHzuOLIlCZP5EChbCWs4DIHUQgyDW6OsJSsJZMU0Dh
RQH8tTDmGn6KpqCAv4/R0vXibBc4V7NIrwzHGMNpkU/90Nqa8rhMrEtRvvKoJVngf6YTpC8DZ57S
E+1Jcrn/c+qlyua9QlVZCkY3JPevvC+9GIrb3D0dSWMAVxKLzEuKWkfN6EYMDMqgPPccqaxm9BqC
YOcTd4YB+p4jyS3Ewqwxe3UDCsbAbC2AkcGDWxkE46EcOfJquCQHPcvT7E2jXxgb+F7G9XDkAkd6
436h1fn/9mZPZajGfetXSVOqFd/biul7FEXMv8GOZq77Mlp819jv/YOUvFP7IwGAx28Yy8l8ydtw
+FjoF0SQzxdv/dW777v4FrLTHw9wytz6Li8xQJYcBXjvcg2m1GDKsX2mt2+XKMorRP+6m3WW+lI8
EWfHuQ9ZAY3aBB1qUgK0DSY+p23NzJTEXydMK7U2vaQuvQNslV5/SmJEhEsYgoRPQ0GVoAs5iU1Q
RZ4xz0ibBZfo9xDtMZBMU6ekbbyf3dfuJSbmQtcvLpFgFsImpRDca7B8lp6+8JMwaAL/sFu+Kfz4
2awnBeHcNDcXCnhciC0Iv4riqYSmzznNT1nFNHDR8ke4epTvNE1OCGvVL2A3h7dQDUj959toYSPB
bTbNTi/SYrZmMSiQnHZgH3tA8RwpwbnWLg2jjPwMqixXPbFapZqy9wariGNCS+XlbwWmaAHwsCSp
AXqLYzWK6e3+EUO4msfelbKPTV4ONl81mzBx6W9ChZ2vll5PxBj7P6pJMOcuPkHgkga+VjSfXNM7
UK9m7Jd8jHQAQXiYLnyWlZG/wrthCkLXeWIutZ0QsZcG96zfZuv3jRf3zQq2q2BM1N2wiafPPHVF
Q5yUmsxip7IOdqxAgRqjWmRvIzW7JUQoP+LRHkdHKkCC5cuaq/MK5IHJPBgcqDD84Z22v8Ec3lU1
1vbq8uF70pVghQH3QkDdVFYXJGhTkZ2dRpSGDt2LlWr61SC0TgqbK92jkFlPgraJfUQDx1YDkUrd
VkYP91d5EOdjANJsem5sU4ldrEQLygL1wrptjUIs/ypxh+No5FKt//IlZwJIHr7tCP3+cNB4AXjU
q2Hx04JK1D2di4Qw0PsVrVRDRMBnWi91Yn0cHNURnRnU3fbchT7FECIEa2YozGSMwd6hT5nuBoxt
h8VAbQMI3YrirAJWKnk+x3f8AQEA1QvuU1GkaK05+G23xryo52Zs/d7q7P2CdlMPEiZGabvqpot5
JQtty3qsyZ/rSO9ODbuSOSp3SVFHRYPaghI00JJyFO+hkZbpV8qwnREqa5GYrjTv0Au8+ebn84HY
1obn3IHaw4VDWHsJjKXw3vk0RTLHczzyzh4teP2214I8uBzJAAxMJRqTpP0RzpDayZee+YOGja6b
5yfG6c9gdyp3boMN+5oTzuoG0GyJRk/Iq7ygxYilI0CZDrHaw1gJ+YJJrIVUfHqmTPeTBsKFdUS4
uTXaUjJZK4/RY/yINetaOqq9TG7DnTb4Mjfb2VImUGnwCO74qwQsbPHr/WsWSycG+3VFJUMoZ4De
OAzeiFsXMM7E3GrmUESW7d5VYcysGMTHBbbBkb3VFwydvEoLXKfWYF/71JOsyDNsGBAppfsWsIla
jo6U8/yky+bmGYLiuxteCKHhwCvESnYP/5kt/MR7PDyMuXN38prn0dsVrZpOAOSm3D61ZPjCD69J
yCwAMvANhlNtKq7CHXM2iFj3bdAz0lTUpIi4bPQmGOgK67k7BROFNFQqAZ1rFu4n6E3Y4M6jC9Vg
r6vE539golsv4DygwHlnwV9lIOvK66j8tL9909FpiyX/UIljz+71hbF9UztRCBHGw0qxaWeMGgYD
3TA9y2GQPoGsaooAMXtlo1QVjV/ka7nt2gBUTA8MyY6+B8atd+8wRQhgI5w7RtZL1KzdM+uSRkDP
hLPvA6cT2FA9qTtY7fOQIx5v819VfDdMxVx0LMsAX/JVHQZi4gtfN7Yay1bRpXpf/CO9RyYncHrR
HAuJ/uDjSsgGpHkAvN1xj4cg+gsUhy/t7Q77wuw5vZCInFfgbVnevRZ6kwQYeUpAF8UBxFub6Uvk
qPBDcHUVczrtPryqvpsAGRilWNXQZoPEfZ34c57n4dtDpxtjWoRP61W1J+J4mKJGiZk7a1lX8QgO
emRH68O4SD/r1AacuLAx+vGbXA/izUUKST3+1bxw8frGZNXQNgZV5tFosACpR5VvUq8SgQn54YOY
XQtLB4O9Q/P7Zz2JvKY0AmnzDOyAxo2nfJ5xCDSl3gpLhxWusSGGq0UwAo7EbVH+FnxCEp8uvpyb
MmgQCyrlXJco1mcIGXUVdjHF3EdksnFpS8ELu25eq7/iSZx5A9HPKoWvPbBaneGxf+QACBN970Tk
b+yqjW63c/k70ywssmuBbIwGv3Q5UKtm2lzrP2ii7tJsWhkPhY1yyH87TPrYgZsL7EVVPo64D0Lw
2oB3aOoobJv6lMC4N8vwwPUYXk3tRmmayRXFA6Hgbgu5vKOJDT0ZD9oyuDcX27unZ6SfDJOaoYzx
+7GRf2JHFj25sFg1nu0nNUNnAIwgzMgTGVtBDsECbsTHJv51mymL7PPF+vVKxskpj2FnBhqb3CXT
2Wsj8TfyXiXnwr1vFlP2Ji8IZgUIMsRDO19GHCOuTIxGVTmFmzSwWGTXQV7sdaQIqMNgEHwrAsBP
9uMeJn2wj+/rzDCHfBaUxG6mWZGV6PDOnfrymvfExGY7fDn64tcBzfXWnBxWor6i+hjI3WY6zxni
n63yd8T+3lms07D+x5XIHmbsa6qjpZHDMHA17tYO+uFK/P42DIBI1vi9yPBBsUgFZuXhgXTbbYOa
TdPMsUuMwmsuPrFDaRDY7HmXftJa+EjS4Q/aWILyrwunjBFiVZrky1t+d1o8sTFRvKbmkV2u42hk
5LDGkNIpFlGdiUa6dqzH2i7p8rogR37IFnP/5U5Mp21u0/Jq5gPjBskkzRFZiTt8eoZNMqpf/OJF
ce1MINGlAgLG/TDw+UD34Y4QLcBQD70me8uZwcDaEzPdKbc1ILslPgo3Hb30X6GUzPdl1LOwKu/N
2VaZ/HwkP5+oD+uagCEaXa/amuKkRt9sFOMjGm/EagnLjdnt+7e5eqNMUwVBmbr6I9tz5rKlyQzZ
V0h3zz1xkEhoedcNZBDmWeqEaZRZn1eJ+H6xpKg4HRfb6CszvdCnxIk+2/Ap7OGHh3RzOGY4n55t
CsGMV1vnExulBPblJ2Wl6ELTlmRVG3YcVdtggPH31+FpjlEZ99bGjdCmeS4cfVK8OpEJUxEdw6hr
dzGcdQo6PAFbNi5xLHHEKn0LNcEMYg9zi5z2Z07DfFh9vfv72FBEpU/djB3UgA7K2t+jgUdwvBnj
lHW6PQXIqX6HlFEoEOXeH5KQ8PTY6h+8dnAPeGnhQaTaA6G9QIkcUdmPtf7cXUSCzvFFfowCSbgq
99R0/VOI2TFJ9vZ8IfYVjKJVeRgJtV7awHVqp5W9X6Gl2T+kARFVzOJihUlyhpY4Ghv2uKHDKIEE
chpOnoFwdzixgoWSpOuhz9TaFAg5DuImmecrM2W905GoWVnpFTKPAgECNupDwQc4emvf3R3eVnM/
jPGRXGl3dtxoc12NaHQBPjl6HYyGRcw80Rhw+BVuFxQ9vzY8JyYfxxLC9KjPOL5tOO2LGicoYHOt
5bHRtqugQfdMUTlpJx8l6MauxZj94lVma7yJucpoL1LQVyfgdyfArdK03qSePGn0BnJEaBKMx1D1
tDLdIP1HquSCRsv1P22oV5v4dUpXTUBti9gfVLIKtPPw69urtmjML5NH9bf+WDMjpMQFhF+77Rxa
Zo7cAFNXCs7iGOXwF6A3oefD3uKIWcf8YqNGE7bt1DDjxBXQEcsVuJ68TqbCFSvO+E9Ss9dSsJKR
83l/q65g4BRvMeQQCTgl9ComA6c8IOKzMtomKO8UdgI2v5eNoonTedc01Usrjl9E7pYdnIrSCyKY
MvxGRLb8FoaZufPbW+1icWHsG1EgeAXrFc0rQUXnM0CpjnDLginrScp5AiBbrxrebbRfMi6UQiTd
ylpETNGLFcp56iTTDtXfElFYoooVO/EUBNJvoyV3xb0SP5emloekcz9If87NB+IK1GAL0b593/Kz
MKAM1qhbTJgaI4tQTQHyReyPZinDF5Ffy3l4L/EoQLZqpPjtn+1s6pvwW3OzygvLlg0Yf/6Krdwy
GW69BNhmVltBPqhL1Xd8/m4s5Ehc/I7gD9lzLGLU3IILIBwvtnXoJprb1oibRcVU2FYhA5Rzltpo
eaBt6pjUdRXiLSk8LtiU5XEqlGwGdDKq3swffdTpMY7hRTEOWKBhSSfgRX03PBnhYZqOC64FF8us
dW5UXnJXZ4j2IGeJ+ZmzYLNncrJ86UqVFGm0DbuifT8q4jtV43zxvreSC7XLM9OoaTwV7AVJBw/u
3ThfeQB9NaJO1tLf0VPdhGMmPumbHQsUOp3EdN2iJL2+m7KqKvXifU3kTPa1r9miAZbGg4zozFZq
lpiASj3mIyi4KZYoHRww+/nCNaWknaZYsI6cZEG0KF6gRXyFcGeZChwLI9bG7+M4hslASfalg/v7
KMIYAJ478l/CIEqJJx6fMoPC1X+LoMJRnOQnY7R4/yqPSVnZS3XqqKmu8wadrpZLFFbPPHpJY8z6
6W1daiB46odHZKpL2lRMSLtWwoq2jwFRcvIuPe9tfXjXPs1Cy8MRuirRgCTSOpjh3lXU6w3kD7WM
cJxmNKuGpZABBKN1kgS3d9Qfpq3Rtl/617HIpMeG5VaD7vfK/0Tp5QTLmrl0OxiV6SY9fpXSgUyw
N3a65+JcFZQWwxBZFptBdLpEgKRKDrIqe69jKKd0YKnjbVrr+Be7a/0UrIce64YOAIx3JW64XrLz
lxkic4l6B4sAh6nlyLUhVexUCjODtYI6+ALhDQOI3f3b6IJyuJ64pVsYbi9T3feNzJ1UHBFDuKX3
FgLeNicPZl8G7ApnkY9Mt6WA+7+Vj40p8nVMPnSvcb8jsi6OuNB6ejcbt1VcWbuug3FAS4NAuC63
9TOAvhqBIsiZB4Mj+2eeHDqqkGmT/GRH4cata1mHUiBfPvECA7k8q0Y370zGkdGRFYuzZbsuo1iU
lvnFG6r+vf0nLNBWajsUhyGcGU0fef21G/ldQURHbyC+Sb1ktoukIRvOtBKX4YEon7N2iI6Wpg+8
4kRnaWno0FecP13MCd96VHyB/YxbfkoJe/fKuqyPy+I6/inkFsza4YsueJ5RZ5AnyNhFxHkZ3S01
/5JQuGR5gbKIKeWfhCSYfpiipnaR942uNh/CJeIWuUjnQ+Z+dLEJSE8FZQBDoEm7I8P24lDnfJpR
0kJrs0nTPrUMC7a2eJnwWwJtddOtSINNPF5lZhXQt+gdq11HNqEsMblMNSnUPRAHTN+UHvmH1EIf
jJu4JhFZ0H8bTXF6Yb03NqpSCodenV1rY4AaOwxQUyp4wEZT9Cx6obsbVA9lmfqCNmjLoS5aauce
20IpMiFun7iYM1geaIoYsVNGeYbScD6MKyClLTWW69++SmQMtEHPQS9puhZtbtTkaEYs1heXjEed
tneP9Gs1jWe3ipIxSb6/fl9uubPNUrLPlcqVi42x2vhb0m2OnMk8kLUvSzSANdJDhWyrnRGG39lc
UsUUwPybVIr8XfI9ECEnN6GRbe+kVPkliPWeceCOIrO+puXw3g3KbUEPailXqkvbEcwYvaVUUmMg
hsovsi4UbnRV25eBs49irEz7yX19i8cCDDpQIXtjVb/IietN74E0e9GrJZ6EAuXi51HMIJJqVdbd
dO2YQ53xdXKXK/xEhK1Uu+8fPD0C8UlU4Zwkbyx8HHldLlPKwIWJZl2s18peslH4MFn5QEKWCcFh
Ol3OU36JCEAMtICW2GKeNZw79lbKPXNvPUv5xPg+Vy5pZx56U3sTLbEUT2JsmnCcNd1KcXVqF5RM
9ygb7dd/u9vXXlagD6kJAYgCLo720o0KHW9AL0/wqqMM5XxrOtujvFBQ1k4gZJsy5/3PM3FRmq+y
v1h8UXGnttSaAsE75vORdIzt9yrMW7NaQcaZ0zEL7lQQdQlHPLbCBCt3O7X+JG/JfvB3JkdEtdCp
EPV/OCS8tUbIAu3mphohcKmT9UEQoNpwn/u1FzrxwrtqgYrY7XUL1al/wtQysiqKSy43KVF1EEky
JW2yLIiEDgomqZYtaEMlXdEo3+2r9H86wKpjVa3nWCQvnXMLhp/J6KnzzR0HXnhLfN2v1luSSfxV
/Tzq9KCoUSOUbjnqR8SsoJkcOmMDj/eJ5BDgJeqrO4972hco+02j1/2qdJ05TAaqcITCSb7IIqNn
LvtODYS0TscBPt08zvBbHbMH25hhKD6w6ShHi/vfFs79dcoZsiHP8lOrHNZHSb0Kr4QDrK2LWU9k
B/eTa+s8LyjM8qptCQ/rNASFwZGp3UAtGanAe7gxEF5DegAhDFTXBN/DTs6RRTWiKR7gJx23A4li
mGlCHgEZMmTL4f2hLyJkftcgXDnDuj59Q5eHLStMpK59pCN+g8LaGQ5CMuRGrX15zYyKHfciJYcp
8hQDOQCF1Mthwxr3ylRNgdKU1I1u46xc5iM0XiX0ANw4+/5slwo/Q1chYxZQb/r2M0E1R1y2T4s/
lXlvJW4U0Eb0fY1j0OHkbpLIqwU58dXwf52W3T55pV+gCR2tfHJe5Pkjkc8joqUirY4xYo2ctIYc
wyFhNne6Xhfg7/jazoxOW625+xhEuiNGLqHqTrKhAc7cZWawoLZQbDVu70OoEEde78HWMmkl5LY3
kis/A0TCGsHW4/diix1PDrq2wjmOKjPfOlqsqAHxtK9sX8F6sIPdR19hMAdgpKoI6pUz9ErU1HM0
nEBskZ2IoUKGOcuwKTLsteECT0eKTGwZmqspL4JT3qjEM8j8T+PIBWsSA2bYvQBqQSDabWWZqtwZ
pH03iOdOQAdpP5u4Z4easFeEjqTBZTOGRIpZbkURJYWTz9bi05k6UC4BjREM22kIKe4SqArY4NDU
gihSgl4+XkD4FttzlOno0EGwF08NWmAKQMBqC2bOYbNgTp5yJcCpmUnQQqJJS/T1qegpwcmYG21L
j9EJQqgSjlpWJ1LPj/ZhJK+drBdARAbAKY+3Q4/gL3ZulwlIHI0YQ6L4xSkBZZzPlWis37LRfNtp
2VT16l8QUFMDRN31jPEQjgo/15doz+MIY2rwqhK2aKjOW9wt2zwbbQq6V4lRb3sWwX49osmDKOzD
5ytq82K/lmEfcOVdv7Oko9e9caH/q6D+0DR98CXL6eUVFOagR55CYDcF80qhB1mW1t9BZt+MQflS
vZA2rdTZwWxJiLhIi5+DlNn8AIHoGfrXGPe2m7QmFb5PaBk/R2MCUmcmwLVjkuzO3FEYk/PO4Hbb
EaCgMWSKxYp7TNaXs4GR0umfs3tvMFoE93dSC1RDn7XAVkMWawuk2I3wORJzw2mHB4/LIr6njYsg
972pxxluCn1Bq8RuWMu6qshAiZXxd7B32ezlox0TS6lY4yOFPVUy/kQpNIJgln7pMvz8FbrQnQha
H71KW+Ub04TJo402aVTcam99bZ3jHD1hZip88GNeHrCKNug/aaJn0a9Qan9pM5wLAlngDW4Tasd+
cXHXqTk3fHxhWraAmciJLVvGaDPugNhGpuUuq4OCDMGCDlzVWn7nqIwy6K0re3oMBpzpT0pYqP3P
NUQiThiwm2oIck4YZZ6zdcgx44N7JPywP2R07abv5D0jVBYXb6wdNeYFQQnt6CLj9B3rFc+/d/pY
WGIN7t4KzLZDCN4oNgu5Mfq/I85SJczy5x2fLz/d475j3NzuGEADCNI5eD5GnANBg4H6iRkB8AqX
ea32phSJs3aaIuxgaHtpBAyBsEniLr3jZfpmJiaYKUTV5la0afYbQGnocxG7Uwy7W2x5ZehiFJCe
rqg8R5Hn+0v9KDlEJKrQARXJ6eamPqVdYCPOPHFTti1tttV2AmVHF+sooKzVskK7LUFzXy6uPBqZ
djYfwuwL46pogLov69oc5GrnHCHk6XFKSVAJFfS7ANTkygY5GkS/S9slRVOvoTVxJDUrxlf1LZsM
b57pUzZ9Gy3WOi8rhWBgI2vSdXA+s0iCZFPM5Qr2DzzlnJRSiipX/k4G53dEiomeY5khw38yiM0V
wn7J1G4MUK/rjRakzJikYo2mjKDBaGQdiz04KvhJ0Fz3C0gpTpdMTqBtCR5wPKVbnglSV4q5z5MM
UsL22j4KKae6K5hvAGHF3XFrxGI2FFeYWUSy1voiFA/R8fgNbc9zNNgfKrBaHRj+9+qTKZ/gZInw
2EnMCeiO47jnffnC3K4jdIyjlodX762HH5qCDNHaXaJz2cH5xnR97l6l0FTHOfZ63sTTt7So5kXt
BKbWcK49/uQeeupIcQMirlCYoQxzGqf+hXqsv29qwxrgXR5SDS7tPuCJqTzB4urcdjbDP0r5Axre
OF80GVzOfRs7mTzFOa8jnnP5A0fEqFpRrA2vEzjgUwVQdWQrMQLSVLZyTSieRrt40+G0icb4V8KI
g10sGoAQ0RyGYfZzmWfhtFN0yu+4TFJAoCaZJm3Pb6+LS1gv+yzX55LIpFXbyQA6mbEJ7fKPU4ZU
mqq+YrAT9c8NalWdBOeHgd/wKCrlswnlQJh1RX93CSdvqikPhvHMdkYPZTQ0/yFIdMSFvflW+iQk
kswaxdzhCxU8dZHs3ChwXg7+yYrJfqqDfNcpH8+udrbvXFNBc7n3+qZktSIyeDw2gLvRBGr06GwW
ICeUk7hCZyyAvQwH53ewJtN7cNTkry7Yj0EOgFBwg2MNec9I7MlTBN78gtnbv4wdLL+81bIyQrqF
6ZaE9qzLyS+0bgs9LLoIJKAgmNBHIdfZInie/I8ReprUgI/9QQ5sNp+559R7/OF7hSeETRptadJC
3AMjmxLc3S+fmHJg4t9FwBmAUCo9kLLwZ0HOy3TWQdKjpZj+xVAAWP6063CpOTlbW5Fi0GN5zXsT
/QqZCoWAt2YSgm83o7vh5pkz+iAd1KrKamw3eK0pEW21Y7HBUuoB8GGU1SUo4Gbj+8boVteaUbG4
uyRlHeQmFuFefLnfwxKJj0aOg/Rmc8twt9ma4EE72zanhBoawEBgluEcEEyd0SP1EPL52RPTguRI
AYaWr4P0lHkyi0wvf8pRnb2/P+0NxzBJ0RaGY9vRwu9JZ+wUHTixcqqzsa3Xk0ccUZNMUfW14IZz
O/cXXmEu9UwpdjyH9h1wW0Kp5QiC09wk0TtdShH9i8/bvm8UxquqIvCfmn3PlyHctazlcVAljagN
VDPE8dX65pwX3WuHY6PUlam7cdoiZrf4TClfvUzO+o/Awyh5kMy8Ijmmi5nJbxdwqug4vxjI9YcJ
dR6J+e3fRaN4J1HS9nlF21QMFRF0yv3MFzCFREevaGIvykDPtXL8YS/LrZunxCl9drntaYZpP58S
nA8HjWrss2v+LsHuq+ZXVmGfo4j/CheoqCK/wOyA8pgaXCZ5mOsheurCbk/iVCmzUEkv5uvnDqW0
hcgF/lBQtOapzopxREoXg9/XG3NPzrIkhxKIXbll44/U5B7lsJFW1rtVOSvS3pWLge7opXtXVu5x
JA4X39/RWkHKy+lheFJ/bAj6r7HVrouyB2Z+rRghdQ2GelT7FovSKV9LSqh0jLXva5YmtRUrhgoz
OYo+JNdAkfzCnodKkLynawLY6QTbnAEQA1ogvUlNkBwpM8PO7oWF02INkzJ+stQ3Afu5l+JL9+gM
YnwNHq6ehej5LqXccjp7181iciZlrB8GkfUCupNV2lcFQhUNciWIzThKSYQ4tPaX1vDQuwKP34w7
oXoR/BYN/jbrBQHvGkjjXNtOe/Rpr7fdVzbXotJiUgmqRJPpWhWRZ+TMpAnPxcO+TH0LvHL6NwDm
x311aLsWQd5hkEQ9xgRhvoTQtGJF8e3jtlsZSc/NOkB2ZBQYdd4pe2DIIgX/zn2RooRotJ8oDYBH
h5Wnp5zQM6bkCI9l5whCkilqoTBSxkkaxCisb46rgTfqXWl2dBn3CFRErX6l+zDx8Kl7o7ak3jKz
lWJPqK6+BrAHKUq/mb6L/NxDulZi6iSSk4XaImIoZrBEUIZ/j6xhjKNtad2UIddjkooNVaDs2h8i
p+lCvsMebrJkSl3BCCBzjbgJJ7jFcKT+KHIAJFDHTrBeeWsL9HGqvif219R4PY5LqHZIliwLRJBz
roKeOPAyeVwjFPZxU/6iYzI2W3eGTqocNTtTuqn8GHHGx1JdJCb5aJtD0N3ykdbtwOHb8Sgqk85p
j1aMncHT8MfSlKh5n8Q3pEWK65aNiSBDGoq+mNr75klR9O2l3zPzDCgJEkX85PA+MZA9Q97NQuGQ
t3iemz6oUyawTYcCtb0th9FtognuuphHMjbVyrBIvgKdW47LKwrIAFqkwj9NsvHMMR0C9KooWeUo
TGuKunQ5IMSLbjUE+GkN3QSk+tXcMaoXzen8jrIbySLKwfl9bgfHAhJm+zywIJZk9ZeMsJRNgxY+
9rJ7u/fW529uKSCZjKgfz/5ukLkLPHCTfHZWmMZNNuC3V50/nGUTUJzU0Ui9vdUxLWyOm9bpgUb7
zreN39C8YcPrRUaYrkAgnvqy29bC7Ieqp0WkKafLkwm9ztu7xynz2cR09hbG20jNbP2qXGJLaC6C
KBBeIKS1T9eXJkwmYP7RQv5LK8Ly30upKT8cujIH2spaxsASpIPR9gvu5A67LRUJBp7Ld1QE9PTt
J5r1Bs2PgBvqjJP+uVr+WJ/RKCI1v7qA2WKfoBBmw9Wx+AIcutRKTq64zap9Y/2aJ5pM7qlLd69b
+cTStlmkV7Tqop8q5Ja0CWgBUyRS+Wp0ig7U05xq9E7eBYpOP+AQYgfewbvm2PgNOoi+c5siAkY5
nAK5hFrTAu+TtB9PCN6+DoJrQ1vFeddqeEQvAcPV53+1yQKNYJpIH4b+sPpzFNF2nhd5WfAq//kz
DBaXwM8n8yEOU0xNugEDvgcYX3kIZrbhW1hyA4ws7RgCEo+MirJjoXgWF8h9kK00gzcjdbTgQSr8
Lov1pBWhlafCBN/I/35sf0qknGUtBsh+b3tHnTgKfqWY8cSaB+vu+A8fx1ZYjSM/D8U3nMjeJhjs
kAl1mwa67Sd8acHsE8Dd/CrnrkV/G3Aqz5GsR16d39Wohov2j6ZSGaYzQKECG2yEVKyeNJHl8MMU
PPROj6VUPS6hiDa4WLdVtrSaQ9WZaJel0aD5OhSzVprnnLROC79zi1hut4oDar7YFhmYAeItigTF
113zI5OHWbOf1JNhm8DFyBHNEXyMEUiw/xr5OD3WWfdbQHC583GD6rZ4xOq36L2122NP69fAkzUG
uHdAdIUmZ5/Ehh+aQ2EFLtZVvmPyPh2J1IhboNI8rh3CCCkV9nYP8HG25hNPho4FAFO2uFBpWzYa
/aGtnS630gfcMYbrsQAXa99Dx6djb8IbYPr0t5boyPQPBG2MsQz1z6cjJy0nRQGD9g+1xXvHvEJJ
WTIt7/vgkYUPNO7MVXLkiXwIXmRbdstd6O8M5pIp0I/OaBEBaFipgMTwqDu5yY/kwhlkVkeVfDqd
SNVRnYlNvFw0xeNBjleA9BZ8+7x0ZpaNKhHJSd7ERhr7C4tDK97YHn6D4BkNJ+Y5QN0vN7mLwK2G
0HQGJvfETasIURn/3FRNSz5ezwt9dygxme44E0rso68+63XvzmhJVbQUOqFjtrUhpqsvKqz4legS
BCoJE+huhNSBcAGghTcmoyCYAOPV+83sWv1vTR4VnWEwnTX7ifpsZhRkB11d12lox+XVlBMHrfeO
ST/r6c3N8aTUUy96xFSkNVYMvfiGBMQsbx32ivbujsnBcsc9mMRSzxY3NLMdkerzJQ4gA5xVFPru
HeKCSoksA4hEIlN+V5p4IFgxQecATkQgqRivtHd2Dm80ipbSED7lUDvgFlZd1ar4YouqhIs6JNC0
Hd1v/1+6EHTX1QBUTrC9t9lie2VfL1NG0lJwEKH0oDFZ1+jJMho5ZYc/ckvjp4Joh8Q5KDTQuT8m
aoBeO1AoHfy1qLtIsEKiVuU1Y9IwqWa3v/oaknhfSM4+fKkPeFYrDT41DQ0nIVKGnWorXAsHitox
bvLb+13QfQTJ6A2nyfkBj2fGmxwwSeBd5yX6TcpPLI/wVwnlP+sPyBChsYtWsgcXfm0t+RZPFWG1
6lDB3Sp5bW2MS7NaX/19PqUhdDZ7j8ia5TJiXz/2X3TlEZd8FdZUrxoUI7+LfpTYGblSNoHJtnZt
hreEVSnSZFMqqe/grJRRK+RhRzDjmAXqXbylBHEcC6oTV8GuHtoKf3aZzbC1p/RbdUhXBEbji4+f
4SQ/zFEr2TYVFhB2IcxXDeAF/xvi7CmojNJ4Wy2kmAsnMYZFWJikDO6Q+dOoHzCN3kBxO+UMhjCh
+3TOfklRCJu8d5mbw4vT4E3g5WBYgegGK1gRi1uJX/Zzp596FOIbCVCeIs3il5QU0v1wzIJOgXgn
I6bGKZMV/WVp2SGAF1JdimFozaeBKeYrOaltK32kSYF7RfeAE5wXgam4jAhDHNpOzMc2V4oQkFGz
iCpl6IucL6/F/RudwSekkw/4Xj3xd409/9bmF231fWmOfC93Dv8Nsk4wbJ2aADjvlLipnchwCOne
ygyscmSODh/Ib4JogGCUKAly7H2i4aYY8VyYgdGGHmP4TU4jLFIKVSx7GQQ4f4WStvoJSxxi3S9b
gzNzhQtR8L05qjNYyOlTKKK1V7d9FhwhGKK+6tsX0ypDLcisSXVqmoNUkbdGi3enPqNSRrf7EMnL
rH8jkgVkjIZBE3GyEjU42lxtCO5VgKqzDUZ18wbO9FVn+QqPD0FWgPzjhSirOy/I8p/LceYYgRuD
QAcZu2B76G4QspR6FB4BtRFilpoQXbNwBa+wq5JDlR0n8AkYCf0iMXAfZ8fPbXmZ4Q0dtdmw4N2u
X9PkYy8LOsXL+KJIrpYLnn4oPjvLlJes78G6ehBlBLofClx4GxBDyUK2bhTrJI8wPm6FE6rNbRDP
l7wtBsDBHkjVuysnXzJE1clLTyRalk3/zkvEQZmb91y71qrdRPSvOum0el/GIVMBrirvICHrz/wl
WaA07iwrXf/1llmVpsun57aAc6Fdpwio1dlIYOOBS34fDZ5FR9O6zJJDKzl8QJPDVxjq4o35Flgu
xqDmsx47iAdj+e9J/SM6w3NkG9hXUdcMFDwR8OlKMAj7Fh8IHIuGRN5aBwNFwYv2BtGJKmRXZkpt
7gjTgxFJaLgURx4UIxW/gdBJ5Up77ofy7GwrxKWXMPwACsal61aKPfdWclsURNHeYnyJrhNTLfTj
tiJQCV0aAu3Ocjdf16Kh2IZPzwSywTNOUPGkU0ppylk6BNJjOtJ3/9tiHJlMD0WdCznOPXRCc17T
Zl7C2sPmQ0sk5g5j3kMRAMfrsYLtId4WwYOvU8WOATjNSs+roFQ3AyU6/NsVd0YOGJA04YS8QIrP
QdWVsvl47Ndd6NyjzZKPIY5QMwxnii9gcgmK1ulBgaBIkU6K1cyBXM5eUADe61wp8oC7SRDrb8v6
XH6BrefZtHJB6uF/1heqKL5nwMK/qHpxAuOIJ1ez63Ww/nXG1pk4Iu29NvRhcNfUMgtDlMyXKi5w
CFCZKHERskGxAMzcXufETCBWjaVBRvzUbc1U8u/rkWKCKp2U+vlsawdliJqb7r+Rhy7X3wtEby6G
XI9MfRaSLAGeOxz6xOF339i0/F4fMPQdyPZpXmXo70gvx0xmYUalAjgaNgLN+4BSUEegs3I6HCGH
f5csLZGmmpgVxmgKiOTTkIxUrXDkD9/jvL664Tx8NqFf8oTWZS6jKz24/BJXe22p8HNwZo+vsvt4
6SUQFuR04Sqfy2lZK3OPGtgik6RqmFYweex+RaYJ32V/ruEOCKOelpIl2n/R+vHPrkNYaoNpibyd
1hHTkq/ngvCIltR90XAasPfBwk10+1BuKRkNfCr1qbAd4XX1PnG6I6t3gScrUDGpb1kUa3F3LX4V
h/+mp8qatTKfqK63oEXb3JPiNzX45O+Lkr7tW4Msao2lCFawQ0tb5C6H0+CMaxDlBuGHUspkfYOH
oWdZri5ysSK8nMS2tZsg43+sKmZ3RHcaKeRq633bC4nBghVOnpOlpJZgXoEeJX87XFXzRyLyHUKE
Ve6sT0Q4ODByjDYM/KkeAK2vVD91P2RnZSUbhRiNXoGPz81BGXKNX47YWPxnxrdDBI+I94RqiQFV
ZO1PBcyi6hd8BpcX3QUr72Ojox9O8kKdBC8ru3hnoUAqrXHf9v4u46AbYCJqCPM6ffws8Ijw80ZC
/xmVvK5Wr86N/XBP47e6M/TInsOigPBTEWsaVMnjrNx1/eeDmfmYhHr1Jqnm2jsaS9ojvV0p85dI
4puG/f+ZtghGGDKqsdcAP9s2538XGi5TvP13I/YBP+Nbb792roDyR/SP50IxdFCVd78WEbaks6+/
j7+zFCe+W9vLjQ0NiEqFSJeotpMbIl/duRSU2R04004JB6x6ymtW3v35bauKFv+bs49RXG40Kcqf
yW8Y7ri5M/9wpujkBGSNwCASkxe6unTSJJHTjUBYBnvItHoq3JehMHtxFzcXVCoMSwuMmNVEOzMb
6FyMk6IYdUEUMRaACLqj373RB/ntjoaAPP1875PeqineMekmAEy64w0um5i7uhvTsZ8D7KysNl5m
2tjHDUfk2p9XyFY4Z5N9tKPgK4K8irQun36fMA/h6Jlu5UcjL4+XJI++/5osNY9Xg+97ZOrKM/2m
8iGxwo30L0LPPhUuKiOOiFQKVLGBlgzHA6Q+PFu/BcZ6E5nCwjTx0Eo8yAYcSKtLYLeIqlfDtvN3
tR9k+rxYgiRvAepUiRuR5BLJdCs8vzyATWyulH+XfDJDTdeaEOcQH3qUk3bWJmyFrP6L9uvZ+wjm
Xz35650I8B3R7tMwCM6p70H3iaktl+hcDE0kXvqkKtVFzSYog2gGpA6zrXd0QnCzfMZif6lPWaGB
4pHKqJKhtDTSO/tQXc28nD8Yi8p5uTWEbvZsdSQBQrw9n4HVJeO1cdUbf5xZhHnuVZ4CShbifPIC
RYjaqiicXSMVhEaSgNe/eSTqDF7eXw+7YC//KM36KpSY32e2CpWYtc0poNog2I3WF25+shJ9bIyb
q/sVXdqQQy1irSjttQRo48tFSrCQAn5sEvWv0jA0MOhTqeP1m2Yq8eaDliD/DGkYPYN4Xx7ITEWM
ZtEVB77d4jyBffh3VnXYLK1NhKu5r/Vu+Dbz0A4NuLaJ0o783C0pdDQc6f3N7h3LX88ihjm7na+B
cp87c+GYDdk6NvJJ1CVCPQKidd9Ep8UkMZ4ANooKmxyUiFZ/YnPAZSVF1tThh8L0l3KHaQWzjW4F
RjffbFPof/w+5an3a7wfztHCnr6623uQ318YLk7ZQJpIPHN8iayXOpVykTL6aw3G6M7CcYOBNAit
QZ5zDW3nmNsOz/AWE9BAhNynC6dRdImj7PUxqLmsB6g+WyrpSsl2yA2TKi6RAsnVPwJxeRqlpN6M
k/E6kmj5BYgL8PuirP+9ieKGmXVoT3L/MNcJOpFw/fwVLmnT/CmePmeoAPPwBZZjbAUWrW3CIz7i
B0DBxhqeEecx4ZJVAs8YzXzygkduLStQ9mXXkG4+nGWeYuUjmW4BGlcrcbs83gOl1ravuNGmAcLj
j9PhqrbjVQ/haFPONxRr8PILMBG5JHmQvWQbLg+rRDuEjdJzpifApQMPXm1v88fqMHVS+YK2B6R1
QaHBDQP2TuTpLlFLgMVwpYO1+8AUtinxRrxQ/Pg2DDQBHwrKMD+DW2BaqjQ3mTrI69mBcGs4QaWy
hpgypiI4xo+TUsbOPBsrKjZDA4DtQTfOBei8BpepcbO2jmFO/ZwE5cbpwto8bUDfp4V0GGXHWbER
x9ygUxS+cRKBWPi0IeKvONAFeBBEJKyA0Vg8iYrf+P+Zm3jK7L7p4cOxEI3+9knTlb1mFMh7IUyB
GDVqx79wmSgj83e13a/R2/lQplhsqQD8/+WZAx8PySBn9SQ2nC60fshW5aUTxBF2xCdkKCAEqbKA
8X+84Olooyp8SjwCBiX+k89zegj2fM/OIxA4Rdu4GBSQEGv9yapJl2+pTCfiJM5AqIwSLQc01ese
k/0BCNWc6GQssTUq3fv3hWHT7mQg4OGlbalWMRLmHxRT5qa82mI9mBzBGE4EU7OyRnoYA35PQdth
vKeWsq9d5LdIgrvREJJpKACtE6kQwKVS20hoCmVXdf9pK3EixFFzjCdXI19g4/GDi1advAmV7XDt
bSkxpHZyu+QM8ZjJBolWwplb1SSdi/Yf9uAzQWa0SNWumgdHJjN3dsaeIXKrgsvvOxnkiXJI96Tp
Si8//6Bs3bHkxbtqmIx1FTz53UnVBagdyvoT9/eKVngsoCN0zDkTuaKqkRmKBl/3RH7Noi16V5j4
ZhhvgvLryf5qTE8AGxyZYt9eJIF9l/xIncZ2TkUzXnvBNgisd3zjAuIOeWjtIST90mGpnWRJucqY
qVQ1Iqv1G9IwYNI8A4HjOq5fs7lIoYHfurvnXgCwqCrntGKFZQyVwq1AdTq25b43VD+/uyX7Kezb
E3mOWzVG01AOfPGV6b8Kb68RmG4bLaVkKcw6hYzWn6PYjdPALyzoYagyKz9Dvjifehucl7kPnQ6m
kibdVbZuTIDZ8zG76oiHHh3nKVLF5FUD562a9BbbUOhwFYDgaP6IPVcygMtXEQOwuy7IhEJsGJ8J
zQ4m8sigTSDBJk4q0GcOkSlWBYPU8/agcgCCvfTPEoFJ9GJfrRBozn5F0ymw+KmwQUDHbXwAIlZO
MfqQLrDZRc6xNPLiSPAkL75hFrUh9lfVDZ9ZjcLIi4L7O+DfnMOl9WoSUybugQQDmoQ5Rx+Ow0M0
y8nXTYUYLSSKkDK7VFhNlsrPatkaiGQo8mUH6VDXbtXAkH0X2wA480pWP53/SCqrehUWSnX7kQ4X
KZQsxY8TbeNacHrimrmSpBN0tgLSBvjBo/x6jWunPJqUx+OmwEybvuxJFjoD99B/Fq+HdNQlBpZi
HjSL3sD2cG14sRIr3FBHqhLVrkWgtAlvw+16uvVDKlnWnr/8gXlS/vCVjuomjIkJ3NG/ugXefr14
9mTtDvvB7rP7fFdRf96M9tqczVql+rbCdK/IYhFBjeBWLsvniJhpkp9CH6q/tKhgwNcss5mb9dsP
GXRmzplpyj7oyUVG6NN+OtbUU+3m+x80puTIMCeZ++/KazJftl0Z7sB/meobJEOOMf++6Z+VIzxc
L2OnYrHI9VrSG74QhU5T3VYEjoCu9+JnVh+BZyJh5CCdxMUa8NaoTyDdND3ha1Qxp0lV4YI6HtlR
/ULBmX0Q6B1hgoj+D5aCCnZM2No1iBxTIkTp4UoixPIC3A79fbDXZAvoRICPJLdbnIEhpbZoVis4
ej8cjUmSqGh6x5B7zS8sMiqPW7+HTL6WG/fHUaA4R8HgB5yj613SCukW4rZqI5mcdGgr+ACyNooY
DDIIGjtI4aZ4Usv3SRUpgtdmCqmwLYtqj6CCMHC9eq4dFoEjLnegKJD0djcM5cOY73Nkp0g3jRPm
+Ze42320FFXZBgNSAY47Fn8ag2Mp1fDPyVc9AKIG83pMjCjSNMzUs1PJlfVvd07zAcwkYgb/hy5i
oOHr1gkVxef0RLcUAcFXNKhKIfXX3ZRmFwx8PbnzOoA9zUEfAVlLa2OBmd1pdzgrBGk9pz3i4PHC
tEvloAICciANSfEvxJR87cNfrLIk2l+kraCjt8+PHIzsgKOAYn5lSPMXUVw5mcPOBx+unHaPg/Fw
Qevts0nwCm+aylWP96ooO0qz5HYn5LljTlRMXuXhvMXsJXfOdFY2ruwCJim+8fgSEi93dxQDOwOh
5HWLFy1F6Qn5czLEnAL0uxoe5FvG49rq29Y/iM6tmD4FD0ng9Y89/lkwzdd3QPQtqSxUB+AcHkMs
OO/w4B0sgfKVpPQrmXdjkn9GHVwsiWe5MzKveG2EHektRxEBv1wiQrGW2b3no6y5DlYfPKAlRZyr
97yE9ZAJUGvcMpIK5tS0YgWMWFAEkPvoYXOc4VFWvhjz89SqQdbqL+BcjlvCRdl7h2Gp4ggAfju7
f+yx7BwndVCzcJlZx0FtohKpi1ff5pfyjKEe8cmTRmNHmZjSVoHJUON0D7LBESB8aHsgqzRdSZu4
DRln6ocmiM4Jt5TVBXerYTFHky3i9jYHIYOuQA96RWCNbsNcEZhJ22ed27n2wEHj/jtdWJ29klGv
mwYyMsglqNJUswSfln+3VMkyXp6qm6eg0Imp3ZSk1Uf1aqOdlsLM+XyyAOQjp6GIe/x/vqqNjywH
8Qm+BBn7dkfjntTaqV3LLe9wYPPmaGBMtyLHn6/DqPjPFP/0tMkoKVIZQ4AhzduQn5CxCEayVCRX
QfRFwTnUINeowKyLZyPkwMyoUj9Jvs1Hs50YxqOMYoZD1hQpp19v5a1ffqDW8eo1cOyuTvQkFech
Zwr5i+eYZVQ7w+5BxsDFjJdxb/ASPRySc4HTiOD3GhM4+8F5qTQkZrv55g/RfRG4y/k7vW3oGWyr
R5VYwr+t8HOWGEVPp7fk/m8GyB9NqIhu8N2QeIOZ7ddRdhq1C/luX24RjqsbpIAAmQncD9YTMQ0B
EbO2IIqMo2rBcld9KS9R9G/LXj0taQyXg3xyaBhwqpQhy3KJgyJA7CMICu6olpuQgrFZG8cYYoCy
mkH1FoZfcJeoFHWx1wC9uKlWBu56dPUZIvsNyU3i8OmdZhOo7VPDOhlwvx0SMOVnplD5rCw++8KK
/GLa368y4sqMi8lb4idddQzA/QBN7wmWpzeoGI3lzyHniKga0eY3Gi7JYuwtl+/gEcne+DOy966r
UsxCVCCN9TOYGVJCs1J9OINKRqtpd3jYU/tI/nmO17QZFyiW6/8obEeu3YQ5H8yUeIAoslDDBZQa
YXJvFCknJ5XEtlvfOwKEPwh/5prE2LPyNmawqMm9WBc0RydXcYYF1iBr4g11ykfAWDMprQwPbQjb
i+r3Cz4ntm7JJhiw+k9DOPw8D1LTOY4jiBK3VFTIAXknj+AiTafntY43Xr9wKVELGRyQ+vot8+cy
jtXRfPKkqMYaRTll4AUYV1jsD8HimEGcC1zk6ThBR44nRroTCieDlP+4APrz2qEYJZvW/rIpVYjH
+9rlPwz0hsZQMMKNJgO9VCUfLiUFdKCfxsitaqDsvbMeDbJNMfDtgZ9ssLU7ZgDM79OPA6IrhciJ
8IvsItOKlLqsSrk24CPg3XLikOqBTidjifn3YhzNepCyW10XUDJcuF0N2Xml2PvHXmK3t5VvB0rw
ouWFNjoQBgq4+dTcNcMGeScfZ6L/FW6ikxKxVb3+kA/MxqFg93LK/FfO2y/XUDvQS82g6jWAQ1nn
Faz4pFM025uPHAAHX7HRIBFHl7xfEavEe7tHtMKN39mK1/tmgzqnEBDNcnG5e3s0dUPnhI2ZHD7w
p8djgvqF907UlWkMdaVcYxesrJtDdGvlKWW5OE+h87PzRDj16fAPBFrWpScJJk/Sg6VSrwWnCD0M
EOPWMaI4goCi5rlKqaH+W/4TI2WODyZwUUPfuwnFK/Ohx2oQ52NYqo5JMMgPRICFZwR8p+Tscdw9
KsiB5NP8dYDtzuE9I++C8G3IRH1rzh8qAeJBHUExQ6cAcw2uFoodYvYHcpoQFzSepacfBu/MTCB4
Dc5aK8CiglK87m4utB6wtERc0yl4WnXDmxiu2Rw2nvE3trXo508FbQ9J9/hWhTwcC+H+PuB9LTbz
xX298AKPf/UuIIG0302YmWK77USXL7c4EZtffAIxdLe+xAdIdmrvbdNTxAcBtyemFSZ0DKl/CLO0
74LfmxpArNBkApMJUgjwIQqdmARoUvSWCdvC9uSuvw7xVoFwDu3GuPE7EUj+QUkNReYzErEZrWO6
T0lA3yucA1cO9K4GtgD6pGQR7Qs8o+XLzdP4mgJNINxlMoSvyEhmSDYS00lPcGUKNI8bjEgaRiGu
kuXNYJxoK5IWyRsblIgWp3K/MUsMJrCh9RLRexCtH3xN76lZRoO0DYA+fp4cPUJiflbzb8zP7x+p
qsPEHJuhco507dtSWW+mO1mCY/aKLEDRS4nbP1Lu04tLGF9v4P9T/gUp2jvCFqveDCRkjKUUcguT
9ok6yF8fcQyxB/OVjVLGIKBVmYLi3z70chyMRxGSiOq/rYmlSVUlB/SsdFIz98KP3C3W3U6y8q7C
tFc0bFnN/AiUSlQwyzRZQAkT0heiiZuUXYyWO673iZqkNdBxDrS+0JwPmXNLSS2TSIWXq0ate/0l
ZelksBfD728DxCQzX9bWVaHR+9ZTvInBMfZsT8AUiZ68IBy/L+fp25GNSJPEUnpM3KgX9fgMK5G+
zUAFPw3FX43Np13cbTSi7W17jX7pvpDFruoWf7ecXaekNoT0NH7REC1tdEZ1CXdwLEAIRJ/MzZok
lB5Zpovlv3ZnNMCJbe6uCFgAcG0UTqdgM3Mt55OkSqg28eK4UZLEXfroYzKYLOgl6A95xsBMCNmj
609NsY5Bm2ZW3tIooCU8rSxIWyX0yJuZH8zSupbisH+h8Uqw/8hdYbzH94ZP5DSCxtfx1X8G06sO
ftVb2gTIjytsg9Wo71Sa5u+39KgA6q5kaKDJeu+04Q4WIXgJXdi2xJ9JetB7KTut3hY3cIZdFNuq
H67+lCVYkaz6woXqxrmKOosOOdU7f7ZK9HExd9LciVPRtOP7LOkRbdxf8HPbLx7T01IqTlKDiKxE
J+FOjAQY9Em/OwFk5SZvaSq2NYyoh2PcCFRpON+FRZs24qbQlxsTooU0TPdlKoJmRdz/c8B2xfeW
U3iyng4L+gI5vPV/LpFP3pebjLQ0wcE5VrUpQFalUDjQWZsoGecz4qKqF6uxAFkWEemZFOualrQC
u7TiLugspl6Q/NCLdx95QxkCEpIGs14NWcGwUGCWirMMUWr746no0O2eqRYK7aq6f6MWiMgOqxgu
Sgv8MU0KjpYRI6uVRa+yHuwNPofxGJM5wr+nfnlbaEDI+6b/OopztfpnlQkmnRN8OePqBcCtXeHS
mKq9RcYqSwDXtW56RgiyoGyEmSn1YWhtMlcys9y5AumIN2/XwWORqKk3tdXA8NpjoAb1ur5VesfS
vpEICgz8Huma2cK33Baf0slxhD31s/OUAJHsY4/pqza2s5Wm9mEYaji3aGOGuiInYZuwag7VgHBR
Oycs5afwVAG9nGkinrDCb4gtdgzuGlEMds+pegPRVoUMlFomexQFmdC8ihuOFEQ4sPQuqKGyHLDQ
XSkMxwZW149SgvL9mff3aVm/i7VTrb3YNzONq9ZvJF2HTvdj3F/wBCnNf464dsrLvU/ST8xGQQj0
zInVNhT4vbxA/7MDatDoQL8YNNjC/hu9MKP0FE8eG6wYwXhrkSLfY4SBAQIfYb3jKrZtsVP1tfPq
lINONK4H5ngZkpN/2WwschspDuHJyknbK0fusOPUPcmNSREgKVNFYmDk4Z4X3vRSK21aZEt97385
aftNwADdvPLWhrf00eaVhhwzsf+WUCpW6xDEAzFKP+ATEDUdSu/6nQUe9BBAIueSnVNF79VT8PGX
f8ktkz60MVeeKFxO6Ar7FaTIhQnhepttItKtiTKSiE4ZP1vWczGkp661DFE91oA5BSUOMuBKFgaL
hi5+ryMCO9Nfu5ao2nBBdKm3TdmH+vJSecrPNmL8DC4gG1wc464Q2KfP7pOaU0SThSldA+7ikOt4
kMaPmHLc9x2EXmVHK0JbSrmxTOJJaZ61elaxJK+xQY6zuqXlmUA1YRURdirxEJDsyS4jpDn7reoq
HUtvImkH+pjLeN6qsPUyCbGoKx3pr90rIufKFMEn4RlrW/3eiEHuY64Q1N/8zM9m4HKTxYrnPc34
nPRT12T30nCRqBKf37Dmnn1aNW8Vi3fh1K8veWQ1xVMzVMb94Y1mtjhaghSqmIJR+Sb6edRCnb/E
VPjvZU66zAUd6DW2/hw4D+aQYya+Hi9dA/y5NwvN9pW3G2bJRpDBrCDhuaLBmfXaRmmWstBLEFwz
0qd8xTP7bk9UtWwgMSAtr/Q7mixE8Ofk8StEYcbmg9/fDF/Q8XwAy9FyF1wO0TA/R+n7cUKNWFAb
X/pId19D/NbJFSLMV6Zw8glxBBoZZJbnTKuxBuvE9BkAv1+qUxM4aR+Ow30FlBmOhIGn5TyRMeRO
9vSoOS2twfRG/hge87EmUKjwPMyxm8q693Sh/eZc+voTAbihRabWQ0tCTmAE5f6ZJ2oZKf0+kaZX
UFtkwENYgwSOTnuaFOouLB7NJpNGFTZOpT26Id3F7rplAUQVaVQWwd1HIULdlu1b1o/6jEjAAtHc
o4hk/BCOu41KxNZ4fQVTqEV02LyqB1j4rpEBZ/QlaVmkz4iaGxsg/U2Gc45CoeimB/sYkympuoVR
Pz9OKkETF3ItlcflaWF3AqlIaOqKQSLPArM3iNQSoEKXnhb4A4L7zpEdGmDPqhkyHJVuQ5djqDKG
3fPbc0dP/zv9IQslhVM26L8Fs5aB3C2FV4pyf8TDplhffn1xED2p/erm8PyGL6/unJUXw3RXNBNu
RUbkXIK1BhrRcoyW01F8DZwx/Iy3ZSt3Khzx8QAHbF+rHMkssV/nRiEPLqGnyNUtZahMQYWvcDQC
BLapNuYBvzuTbHqgQRPv2Mq5CobzemiPme18izDmfqMec6j5hJha5oOQ2arTVx27TaEcIhTV/EAQ
iDe//zGF1H8rVm0btujCfw3u7sZz++L5mTB+WBbKnvlSN/GpvKpe7QAqxeFSx7M6GmHIC++ZZMe9
JwtmvF5vTsLyGpwMzT2o/6NOzRS4JRZvHmWJFSWEHq/05ok+e6J19JdQrEBqF7ds1Th3fkltjOFf
ELgGXuPg+9gjII9pMbQbZZ8I8gHIiyNydGxUD/FVBmFLq95KGWrpAOJGv73CCm/BPqcnygU8b1bS
tGAb42XoSDIPCdaGygY09J7ldnP2Si7uEdAcXnyCpE375m7O6sfxqZq5NOO8UOADJ6KRPWJ2RvIG
6RkL/plhBOf9DrXbhkrk1accFzQrFNIVP8sVJi+Es6xUImbG8il9jGzVLz7T3iRApKb2GzSYu4F2
YETVVFaRaz7aaHTwJ2AoSXmLDGjqN9iNkpk0xPE9gCcFTZSfaACnXnfWY706V4JFD/mu68MPLyG2
EzOWXsT4juO1yvioFpH+PLJRIRINnMt3mIY62dNW7Tlp4pbjTTIx0OFOaL316L/gRCaLLzzYQa1Z
0Gdg0QUsOJvTAeVD/F0gApsu5Z4/khiFFGu1A1/7msjhpu9iVI3nE7qBWpO8B848zmNNRevk/7Cy
0Fd1v+QSZ0+muDyRvb248aRhez03m9et3egunzv4YL564A6izsJSrskV4SWEJsxgMI2Aa5iLJiaU
97AWg1gvGojCcS2VKu0IWwfcpOcEb1AJyjUKbLNlLiXmQP5a1HfoEYsd8aj1x39jNnOk1yZc++ab
dSQrm7jiLHQ51VABKOVqcDy+TC/OusC4AEbCToxUotUO3xnXgwy877igr96znIixS60SlVG0hBRo
YdJfcRyASpvrH3IvRUcV7flZqEqbcIWYIAS7HThSuAHJDjRgDfTKWzeC+/r9TnwPxe8n2o8TXiuH
V+kvnAUcD/pjbMbKcnLZVPTznL9FHgAZJ7HC1tqnA0KGEHuqdjRECHHonusm/iwTbOJebK9RowvO
99duAOFdlUeVNmhjt4Q5SvTgk6MqE0DQlurthh6RSWzc35+kUnhXia+lptHvqqS+RTLtbczicu4/
OLEpnaqV1D3tLmy5fRESxOZPckFM3IuuOxyiJ5EbmEkg5Og6eLkF4PHY5m0aw7RuuvdnLSP8Q7c2
9MJVLegcYiFGhAVfP94VMrr9sN+EaPh/xC330aqgdDxxy2AxWonBT0eJ/OkHRnb1RT/vZ6cFPXpX
jMsHBb68UeiT+p2RslktIcHgfeRaJMsWfVszxUfc7bKIaCd9qUrWOX1YbI/3rm8wu9ts3SbH5R3Y
bkCyKRMlnmy6iwhGGYiL5AmR6kelPcIxgL67Gm5THos68a940fHaAhAQ7Po8POL+BkoQJ5VMisR7
DoxExxbn1uu1KjP23cZp6lmvPyOzxXDboHc4Gv3b6A9B3fzHu3dUl8EHGT9Eu4M61wahB5YU7rCd
oi8VXXJU5x+DkqEit6SycBrV3cUGfDGey/L56q4dogiZF2wccgLhIKQ9q6NY4OVlJPbIvSTcHLBy
InhGGklVnCU/mIRCQLLNEwhrPF0AMTP7jiV4YymLDRsjKpDLe56VQSFCyaV0Lu/TwBxXbL6Efk/x
4BhGt+6HfU7tJ9M9ABL+YwStYaltT8S8onAVeIEI8RK7MjsyR3aH/KwvqE9wURN62lTXTfHxh3B2
8roJYUxH4jTulTxzkEjDIfgxxfOKohTUKr+OFrG+tVouboTPrPabbJLzWljaqbjJFMfiB1ALrV06
XH9nepDqt0kJTzeYQPpNhSIfV4D3Z7YNZTBFhE/Qtb5yAyrmn8CX4iSFXzwRzDX3uodNJftykA5S
TDkO0ZAx7recw/YEVBA4PeBFGNpvRlgsJqC/MTzVVc5vaWmOaCOWgr90mZHB5K9pDKjByLaNfxSp
vzMRwAdGpiU+/ZuprlG6Ncvn0GqDTZTF/JSyQEns0OQ7a94cusCMifcWS3Wuq54acfZMY6eFiAGF
A3psIXZk01KwEIpiyShnQJ2bteom4Ym9/nQlj9ibJPuNIKVKh8BMriKK2YU5kGyT96cnvLmX67mZ
Vioijk8kBMWTvkAOMwy3Qsdkn2IyMj0iyIQOwgiAIvlAx8E5sU5/sHeLOLw4+42eMQypNgBzwDeF
c891STYZb2soQlpbAIJcvlKuanArIt+v/WzDo7tjeI6yhyqBSckH8WXLg/7Td2Fgo7wew72JegGh
823yF5dBlZP8qsKNGR5nwSwDRdzZjOY7uKNMcEZcQMaL9Z0O/uNR7qT2wLLVqbAvXCF4gl8ubLjc
NKglflkBqVlUvbCZv+/yh8AhLjL39IBUDO7z8zb5KpnOqCFq5pU5v3Cxx/XlfsX4OYFbOK7pfpaI
/wUuj0+0VTqS9Hv2x0b2CnzoUAxTb4LB60u42gERbzhtFYrJlUVUIjF6q5+s/9CRyd2iPnGIjlw4
E0yVv5GYedqAwfHfYGLd01qLVfSN5vCjej3RJVOqcWzgU0I/DhMfjVf27LA0FkCspiwGlFXlOOho
av3J4BbU0EyOmbdkjGZ3axLYNnODgFkjqKIGpLCRuFemhQPqVnAhaL5uai78JiAdcFlvCCCpFoIv
pQslUfpqeFPVbPdCObjfB478IX6x5FEMgsAOzlfjoZJcErRGNqZDnSYSppRQTOyUNEvb0c7LRttT
balL1qGXRuSQGs63jxdMFd29tju1HZVjwTMKbKVgPkQW12s13YfxGHE+lmF55ZwSKe6r3BcgD8yi
xXQ0Z5I4yf+FRo8a5Mfkmv8KtW+rVPoWFeZchEEMTHz0lm42Y8jVDBreFD/Z1av4hIU4v5oViIYa
LvP9dENLIYf6dqmhH/wxOwV8vXhBbjBRpCEOzCKCGCT25xzx+nk7mV/v3KLAjmRFf0+UK96HUdXz
OPBtSTjAIgDnAwZnK5FTTMaYHNo1qXrZWIOa0eSbMxkufjd5fHhDXMP/45xZ5fRN7E84pg1TheWM
NzB9aNDCzZ8RrJ58PynD/Wp52ertidxoOIe3DNsbdRksfkOU55jPntDZ7PXNEglaigcU63qtxxAM
1/bAK4VKUMYv/FpBUftv//RmzVc+dadFGY2Csw/YXHnJ/pzzP3vF2hJD4MaTRBonZ8KtFk5xE1KK
voHwcX6BTrDdmh5UtJUGmRQ3WYfqAu3C/TdDRESu5ATTX8iWRbGOAxVclNwFfhAqDoiOWhnj6JHg
QflATtx634PfajNIOd3jRUnKplqimuO+UfHrjRHATGy2HCAz4amP9cZw4AaEyKjp1HIZU7vqNP5m
bvJM1XtyaDnsz/5Z9r6V8SOYzCHkfAqhnDspyDCXOg1CEm/p6xKtQnWl2N/bF3bmFN0PdpH14g34
/jnZqUwk0o/Op0aL33Xy4y9s8sNGa9b6+3IZ9DnJ3Zqg0e2+uiLP9WclLlvAciNWqv+VQ38l0HTE
itwQGMT9L27pYFZ93AKmndsh0JA7bWpKfEsnvkpvYfikqNVqomKTLUthErl+6bDz1DZZnZ7o/NzT
RLCDp7t9GoDkj4pfsTY9Lfc1iJanaAFDWL3e+dFc7Zm5QPbsluROIAL8erTVW9wnrfnKEzAiAD6U
0+FPKox4E35bkTWZRMhFWEYQip0PnI1a7tPMb1gj5u5do8N6RT7rM99J3RXB6d/S5Vf78NQSwl3d
464eCQpTf3Mr/tflKIJFKFTb/poc26e52DNN7MS6zfGdp9R/LARx9+b1JJ0dwMKTZYDxDyjBS8DS
M44qXGdbR3vCvDIdhYMt6ZbQHm1WARrJAqEiRWuzLMesPMXptd7mTDK1XmfG9bsG61akeWR8cK8m
sxoHgbjjD0UBT2UBcjAM1ouVV98TyaMP60zk+MoQF44DRqwkUsAZQ7TAZoVEDmIKVh0cG35ZSnhd
u+ezBSfhF8c17Z5d3ZjFoNGc4Oey0ivXqd9FYHaUMoSl2SXEyXK7glwvV8mU5cu0IpFYrilJH0f0
FIJoTezCJmfhjI1aSwsKvjLoOKTb5TyX6/upELQa9/B6fu/hDOOyq3LIfS0Pguc96kRFkIUgXngT
oJkcPB6dKFlmO6ytioeLRab1JARvc0fG2Or+mIxZEW4G197RRSJWDTMwYTXkwVUko01v+UCimUox
Pw2sdYD9sMSTIzAK+0w9qckJndbWU8HTMQ5xxdux2NajyxDo6CFzEEskdyChxK/TSD5fHZuCxvJ7
53LnQJ3Ano2rVAc6BfhvJenaahuW204KM/KgjWxML+Po+f21mWociWygf5OQwehfexGz25uhqOOA
luz/5awmXQ+5CtgSAQfvd6CvTtLR+OSihNaIn3SgkEAP5/mQyBqSJrKAMdyyrq0lciqyPOf1EJjD
kc8bhVNPXH94MAgx6kqcZvidoO4lbWYk3ixLqYwaFVt8eM4ChSBa04TfBDrzx/NzGLK5pJ6qEB8+
bUYp1gOGNWjCUqoex4YD6XeOp7Zu9HpE4e1I19q2tWyA05W12zq2vjV0VbKkTKuwo1rRQ7rTKnTL
eO06JoCgtPE5FMDHzHlQhAdjvVCpHu5i+/dOvfAPkbJn3ywI5BxoVN44QfAC56zEdZ5wWQWffuY8
PYqf7hOrM6CuFXQaB9645lBME8tfuo6bKG7rlOeysp7hceDdAcZWGk6wpUVyQmAhY46PCn2JP65S
Um2DWihCIbYB1DQdR3Rk8ZU8DUIaXUPPxDIDy8sLTwVNk2FbwSn4jp3wPlxSZQtQGqWDpdSnESFh
b2Bwe0UvIFLpscv01zwiclWkQ6bEAe+hSpOVzDb861SY38diPp/MSQQUls1mmgDtK/uBhi6sZzrU
X+CqNcKsKd2uGIkm/+8RvRA4Ee5z+AG4QcckSUo34LX+Y3wweUzkL9D2sLiGaquaqxkPkcumXD+Z
uAe+1TM5+U2mj1I1zQLAjJ5NOeZafePrSLiqZ6QUtGdSHLLqubPheF/RnlYzP0PtMVsmI11Obo8r
qRY1duzwvLXIGFggusesbYbdrPX1bwA7c3Km9JWkOfqhUlAP/ypLK9/qHzgfDozk5gSDKJMyApXq
/B+ztTkc9UsVd7i/raRVvRAPZNByQ+YjNoHlvXhtjIBQmkLcWjdLK2Goz3slQTnGng3zXYUWQjTL
iV/SI6GL/aNy5zRAELexxuVH7tIeLlzJi+Kfhg1RpAIiQG2gYE6GCPMQLlz8hVMnijhG1Cz267zO
Tw+b6VHTfWsFC1n7KFHoN2sIr0tKC96iWjCtmwaiDxh0AhBre8b5NRQB5sgNwlrLEneD6nFTbJxk
WHTDB7BZund6QXTiQPbKn4Fk/HpMqpU1WevwPThyYDYePqDV6qIDYvjuDNWG3SM6+CBXNeFqp/Ja
3Opb9OT9pGabjMXPyvNP6uXxiXdCDnx/rlEcl3PnQOSwpjgFABqc0Jdu9G2uUeh3U4IXmxKxmjxy
k09v/yzJpGGP38LybnvDQUQVerxyYpAEzSxA0aQqtSdA/NyBm29rjBhnhvZFpsB5eKqtUqT26Tto
vzNaRvoPN9HHQOnDbmEuZ3FJ0zOyymzagDanaNux1+bxVvS2hBKEYks6SUcc30zXnQyylc+56xZG
NARX/0RSxNVjZk6yR0qYnIdR5obDrWersyUx6VzjUKWQyiwOWHtOpKmBA+vxvhaUjvUFdf/NIF6v
co3MSuiwXPZv4hWAUOkf44GIYRtT+4fUYvE3HT2WfK7or3neA61OCBL4/0S9Jgc9Y808IJcba/zb
7+g1jmEH0hNzNTVPhNL/Ts36RYCNo1d3khSbDyTWBUuUKSxbAihCaaDwDLdoTtjitSMIDklCQWcz
5Cq86M7SYbvul+WsIxkiBtQjmo2UkW5ZW0RMG+5PZwhLJHjVbXRSIEdO6rYlOlU8hHSIGaBOkBxd
sJaYA3LrPMur59XMPA0/GraZRJbvH/NCU8YVQjmRQe5kCQUQPZnD/P7PMy5LoYIP6e9JTvvC3gHS
TZh5t+tYBp8IGLqchymx/0P/FOrgMCF+XJun7B9rnB3CjS/TTgs8JEr2QRkHBb3szvt1iL90Mc3f
OSjRaZVNJxPwZHX5e0U8g3AnxVdKp7IwPClWMZo4+YUZSmk9BHMwPei1t4fcq43RfoK05uGJzTc6
cyRp6P4PjNRsApRRp/u8ahsrxwm0u0cRZmfi63CBFUeD5lhYapf5HIs74cyYRlaOAKNe5KLX7Z2Z
XbLPmSHfcGU8jxj5ydQUzbJhl8tvbL6Nbh32ocdiW3zMEW4rDsxK/MpgUVXiIKVh8hfDDUN+nQ03
nGFFHROuJzyrzUH9jhYtec+Au3MVrydY7rSZBitKZwOj+xUe1Zt0GhdT5DWPvl44+xSaVJqBt/wa
z5TEC6gydT6Q6P9qhA5dY2k2Q1yfwIb9btevq4sLw/6rj6tXWZEnolqBwDa2tgmvJETMrLJVl/cn
E7ENpd+QQkhE+4TlWRKxG59KhEv41ZY2MKv5+B7raCtVZIX2YcfFA4nFoJu4w7QG7djq8HY6BVPp
QIU6EmnAg+90naaW0hORlN9j7hL81BWtfGCFpZlqWDErgrxMhTcFyAE49co2d8zbHFWGYOkWK5y+
UieMwm9zs051r5/DScbMqSFzcuux7o2oZIZYlfttjgZ98C901juITsW5pZOxZ4ntAeUYM46SUav8
VwteTXdRZMj+sOx0iy+JbxUF2kzfz6YvylGae3Rbx8s1U18VmwCfHPxLnU4fUmVnq9bIf8PDJcsK
RVJ0LPl2CSf+TL+azjp2JlyMFfmB14s4CaRELBFF+2mxyPu+bZtnG5eI1lmeszoUDK61l2Qxlp0I
mVoPJP7zzgGWbhEryuhyyYS5R2F8lH7WbwZtV1U/r1rNCU1ByCsa9GCieAE1U3cRofjjJP3Nn58I
8ih8JeU/XoE2vxAKFlO8i+dTlKOwNG+ANHJfBVYFLT+i/172WM15YDbWTCMXUgR5gBGa1iwcbDIL
kpEhHILTUCGPaewid5so1ywPUByQSvKP+xp3tCrldl1S2ju3Cg+eDYs00UBtF4kAyjxJFX4fFpx9
KEpn+sv05FeDw/ZIlcR/Fi50CXolJ7BZNXaymqeMy4833qphcoslzRNE/feZLThm4StDS8lsb4Mh
1MO+FrdQXaEvrinB/55Vo8zjTK5FGtSXa3V5+elHISjMjCsXDrQwOsWtmX4192Kjmts/QaKowsSu
DHZljZEpRIOJMjm+h2ez1QyawT4Sq5dKmDNKSmgEhn28iFqZSDjTF3b05hW+cRT4a364/siFxD1D
N78IqIEP16NmiSIdQvjJ8aARpK7ZfyO01cl+VtPhhX9NN1TMyfG/q1YuySxdsTI7wbDfs/RCkLsv
FRV+oaI1WdHkpEGSqZOu4BVm7qCJ2KjsCKjv8auEJpVJBO+B8v9UWdo7w2XRCxIokUgGf8ZjOgoj
4e+p2WQBJ2BDRacYnXRVwcVuNtMOWBmCqlsdZzvvEHVqwN8/hKl1lskCH4Qbg9fpULM8HV7uiHbT
lCt12AHTDptVMIS/rcOMaSz4jPiUhoMrZc7X0V/J3GGosu/X3vyiMvn0wPDLIylkpmkSq90nclJm
c7RFUEPeWdFeVBlT0Tt2T4UUjF7fQE0AO7rrqCpKLRujzBPj3CN9OiPKzNcf6vfZyDYkS5SP1UvA
EmyNM9nJsnM9+XwnQAuEdzCzz+5CRKWhXx4hpuKbhIM+G/rBxfIjdUett42MXYbfSk831QoNFc1r
c1/PEsfchLG0EeWskxV54OvwYdnMN/6bqyctR5Oid6YnpGgbPUYvMjbQLMF0bBk9c7gQaM3dDD+f
nOHiHtZnId9FWiAWZaqta/9PmL1cASxXM6cUI3aGpY4Fn2FvyN+oS+1uzVlWPo5/VDn5cFj6LWZc
78wApObcpAG1HroeVut426vHZ9JmkkZ4GRA9CgS255tWKy/CKuyflRov/DpO7f8OfwNcktulsA2C
uBGok9BwVl/FpHIufyfUfAtnkR/SY2xY0AFIBEHP0h0qLEOvL4Sq9it8Ls98GOHHFjM+UqL5sJhi
VCRH8iNEFYs8ePJMDr5b9p4AQ/Uzp8LdZcaCtfEVChIKBYXWHWm8Bgkbn+3t7WMfLlF2hDqVz26D
naM2jpixF8enhtF2zaaqXiSY6Zk4/3OuBv3BPLs0ccOivNZmUK8bqQMZutyUvEXRTGxeHBwrmtvB
4hA2ludC7fIwuOd7i5qBKxYulxVRYpkgqi1fHpOmyyuaugYh+wbQamRh+0/8h01D1wCe3mdHrCmS
uba1dHQntBzwkgKMTByTI++CSB/NKpcuU2m77O0sTY86L1gUF7X2OAsXL4UhJBn9UnjLHgbfW+5/
ZJ2cH7S+uRXTkcU7o69XVE2IWEMcK+rw9vx8gSz7KqMnsu1MOj7bCIpF2zgU5TvCcki0xK7/0hqI
rf4T2EWX9c4KcOKNWvaToSHgZSizBnvpmwJJBejNiz7ckTD8uDFqdqYvIWLvDS8VTSZyU5IgQ+h9
ZKuXoXb9Gw6g0/gx78N4x0mjrCrTQ6M9Vt4+lmXofkg4BlpvkuLI6ZnqPuLimreqGhhYGFJQrTOT
y15AU+ulgeqkri8hHD94sR8F0ReNZKaUiN6CejIm+QM0+kFrC48DcIdTOsRejRmS7GgK/hyIrofu
q0nlw3HCflCkKHQnyUuWrF7K76UcU2zdYqQOItSL6aKk9nEmVU0/O5q/rg77DMTIdqmbqQ56p/yC
thRPVkaPiCLRQPsdHwF0NIilMpyh+9+Pdamzy4xDUpPX09MMlfcjvikK5kCcz1hMJMv460tQIXiu
YgoJImd7k3Ir0i01PBY+Pq5aOrRtFiU04EaE+Wz8kpiiULPZJF8j4pRreKk0kgzniBMD1GF8XrRI
F5VyK1ozjLuwTL8TJ+F0UG02aXYgiJIfTXQMwprBlgtEOKsoDMv1UNsod6wq8nBY3NFBJo2iWDc3
VV8Yzw7D2qkooNt/MPoRzjJR8zizCbSWK2iDh5+kaIJDQ57Aj2wbdbbWXmeK8JrV5Tr1Zx1cCbVN
p8jFRozFywJdc0p1QXq+A41osxMG/0LlXLHXBwYpRGRLnAY+xA7iEEakW268Ya8tdZ/lSDj7PX1k
33/XsVrdv/E2PYEnrhFt9N44rnoSbmGs4bLtJuCMtOdtsY65tSXIwpzypLdEoopLpNlNURPeA9lq
GQWXWD8AFkGmzzUqsn1ahAC17/3vXc7dM5M8jBn4TlPeY284uAqmcGfsnjB6TXDYBhxhrnmFk5uJ
wzDdplZcW8DkqZzk9fp7TbmC2zuP39tMcehTUIqrFcNeNTIRAo2j+R5Lrrn7yTfNiYltrTqcJULd
JhJPnHnOelI63vxgX75zyZ2Be9U1xHT7e9qa/szvYhlR1sCYgAQrDC2tdTmmYPG75mkXYdFvJQaf
IMC1JLOYakqC3nzaloGR59dRZnCf4H+zIDen2+HF0CrEf7hTflbKY38YJnj8WprQri67J1Xh0pYH
LQXMPs3qrtM8ANjR15FYHv53AEdrVK2ipPes+Nzuv1OfAoSXU0TeyJBeLjF5ZF59N7PE/MM7uZau
4JtgXI5U44BCQ6zzRPxeeallyDSvHIh0dqQ3YjievXwTK8l6jyRQOlr8FNc1QSwe3ovROcpsMGuS
W4FvtnRB8RfnwiZh0ZzaF/UsQqkR9qkGIT2NZ2QobUe+4k059ncTtoWgVr87bAZk0MwvIDANNE76
fW5snDVbgVCa1upDt8QYy727ShIYuvE/IJDRROefIk9MEN3vsD6KeNlpLNgQXWSFbKQrkfolABl3
IuvFChVGCuAYltrB8rkWPg4t1/e33w5XtTlAW1huLALQshpZ/Nw+CsMW/hWwiEQuQs29OxwnivQN
pQqDmq/yJ+CbSE71RKxbWjLHx9RzDjgTTa5YNhfU2okqwjl1NxOFO6uvG45Rtk88J/BqQAylimAg
P/4ReDYeXfa0StWHZCBEqQDRSqmGGJd5eyxiXB3zkSJnpjJeTa+hAaCPqcRbVv7M9CVovEIY/oAQ
1us2xHNbfHNNKZ7+OYiWM8oaERHwh27q0Dli7fP3VDoWQQ14GkLgBZbXpXGgaPzh6rAhhg5eK+Np
oms0zUOwLyMd+k+6JOOf6voEWkT7IGbbLqzCICuwop3HQaNFwyUL4vqQ9FjPeg8i1G2wepe5B0Ho
LcwajmCV2vXp8dDUtEcpM1+vNfnOpWDCNeyaCT3joyTtoQNsXJvGrF2R7WWIoCJ/W98cYCJWG9nZ
iIgdec+CUw8KC5DL3cAmMtxtRWerJXT1rmMQR5pOUj1ooGyM6+iyeNBLGT7JP83FXWb4pYEA1G5M
27KIRDanI5BpcIf1TRDNmN6opqsXZsHLLZUt+Q0pCNfQYCPbBDa9L1KTcGlZsE1yeI64s0jiA1ko
PPflbBcA+nURQNQDTPSKveD/JIvhMP1AbUAHef0MpkTvG+okwvL9w6b732FYm5bOl2vD2F6CG8b+
HpE5onNPfu9Dj63zcB0cv4emeI3XxyfatWBojo5JDdJDHoN99/ZyNxZatVOJdIg9rQWrw36OO3Lr
LEJQFXmQ71yxTFnNEJtmruhM0lJ9/5Ydzgn4X/JACEYzLde693piN8/4bKo2QLvk+gi64hb2630B
9iABE6SnQtu0lScFlKDox041F1TZTR0WdS/XFDMq/Jjuo7hL/gfUGvzl798K4Bi50aRcTVBd0+xY
zty+bMyu38KeTX5Umc9tQ1Vfdi+NzbX+bcJ2MfxcWcSI6M8xok9P/mAt3vSuCujzBzJkKi+E9Qnu
HzqqpwqGvfvnqPWqzf35xUd5CgwIEyhfanAv2wkaq4KnVL7najEQinXxoj+WdZx5zZBqZ3qn15l3
xwQcuPPY5VDCXHqxIUBNVxpTR9ZO8O4V6tEhn+PyA1MfiAMc+JzloWJise3YET8ZN2UhmZFv+9oH
EAq/UxYb3DxBawHab0kh0ZYqcvgQKGHymnWi/g1965c0oL1jzOhrmYJLKI9I7RgVvENPowdpHHo9
3+HoVwOPB5CO19Dq0b+pozxYhrt7y+ZIuETz5qh7KJrNnOmqh6F/sMpwQTCzKCqFTq5wJZmTBEs6
0v+Y8EO4Mg4feVDSUDPCjh9Is98sOJXDFx6pJmCxtKghwn2MKmPB5Te/V6fPn0El3VrjEDWfTE+j
3jcub7HTadxzVCGa1eKzRcJrYrvjj1p921yim9sC09o6g5Ri70Bwt3OoCb6yQyfCu5qK33Tqg/XZ
zgxjV61SZDOq3s7vavQ4fSKdG1NXrHwRZhNAYSNPiy1p7G9/ni5bo38kHibJ7iF29t1a2DLorWg5
aWb61PUQjnhbsCD+14mibw7omdsftdi9NXSKuAaw9ygCkbY6iQZRwJWBEi2NkzJtOxBksCO3AuHr
cosg0d8sctMrXWNtb0piCMqGAXG8psYXZ0+M7SrJ3ONwXF527bJsEqXQ/NA+yaCiTNFsWo5pi+vq
CpZPYkEUadTmUWvGdISDukXyodMaPEihaJF+L0I3nohSKUF9juvdpta0wthO/CREx1pvHGQcFdOF
oKJt/xoMrd6XHfrdWpKT+VKnGICyYgh/teijlK8THN73hiJG5hixRi0M0HgTeBqFT3eNMsBYrvK8
J3uDJa63qT9IJLBodQRY/zIcSagwaov70WRI79OYUvVm1yNo2mfT0+l1OYFujpdIjuYVf/9GVZAo
2um4t7DatrB8ylzKT1IK8CJNq4jsyE1hxDXpykrvwf4WkMqvztaVs6UF4qXA1yTVV0LmesoA35hb
VrSvn7xqd0jmLU2eyRJ3sj3SiBkm+lRB6aSKu+/94hTZTiozGi9306O+wQ7BZMg+kI5JiDRd5RCQ
cQ9ClLCGRfLc8ydD25/8Cji6/fjbcy2jqTa6RVK06HMWzJBRtLaQ02Ranwa3MJeUMV/1OR+4aP9P
ek6+ZU7O5f9aeaBwR41EqLbd0/9g8htqOvZjcoyJH8AgF4Qef9m06pArXtouITDs7ppYfU50Ashl
A7efS/HknjVqWEFE3k3uo2l8n8q9u7nRetCMTx+bKO+p8aFaWu1HotmdkBGG8P9eB0uNoqC73a6l
kqiv1O81t4VX2FEQ6iElwR2fspg0loqDiN7E67BclBSzD0K0bntyOVephAi5tegvPr0sReaaJr+X
0QhY4tKI7lHF7MG+LzhCN2nME5eoFseegTwrRX6sARPienwohKE9nB0mWZrh3kN8geVK0nQJCLpT
s4pl9rt0vjvNTrgiju5hO+edqAYqBT8vqqCAiVMmI8b04iR0X7ETAfLT9ghnAAg4Se16VPk0Nilp
VvJNQPUiX2wbu8aCcm8/773kD5S6KqQzBzAol3wZXexGBtM0EJHa/FSXGFg6FvkvtHRGf9XzatQN
chLoTgiURNV9dxOmzoQH0sAt0iHficzTJjm24hXBYCzjqfJQgFpn6qsqnygFmUtJX0FNO6fEaVHy
uBUh6kDdVDDV5H7bw+AWSy3jlz5KkIST54lYFapneSzNyU7+WuUKvhfIirDyC4n84+FUNZjgGdRg
7Fs+thiK7H102TqW7wlpYPZXuKuxHxy6H2AOFFS7KOZLgakqIXErnNUZUG2XCQbzc2u+MiVCY2E9
PMV3HelpRfBiL4m4Yjr8s3X5c1f7X4vr/FGaPGM/Eepc9chrdvLkqBUzq8Zv3scVTUagzzkPLCy4
e+GYVw4KFt1PA7zBf6dJxBVpzAkukRL2tCES+8SHM9Yq/TJnwbO6HAgzm05eHbJHXZSsm9qEQI6o
FQegR36cnr0Oaq79PSmxFyS/siAPW96ssVgd90Hu6boMTSlNbF88+HurJYPd5ZF0AcaAV7cjI2TZ
vBLoxV74Wkrs8VYjDVhb/G9/dJVYnae20NV5QCbXSPSxiz4TCMqS/agZi6PSQrcpXOCiP5W90hdO
pz7S1PWiAnGb/JPxXxuyLadgNUYSep4RiSm4jf66rb9e082OuEq/gUJpzbu0u0F4kAfDaheM9OCo
uxQ98XBVUX9zxpZ+yIXxYODJJiNHCotB12T0Py5ylFAZSZG6z8Kpcb5nAr4wikPfopVVNZEVZGqe
VyVgbgbBDAFQAnBGklwtMLUznN1ZIyqIEXzYRgTGPSGBxCJimpH4AdWQ5inwcLjh4SBvzj+xVTqF
kFuyY3Gw7HhdcJUstPF0SfGLL/OWwrDKyTMY9hPUSDL1Uh9fpk7AhUq9x0zTxaG/8sqB4FsOsSmF
bEHA00KDQwqVYwarlT74poHdoe38hTDdgEMdxAxu6vWjRsVSrhCBj9p61za8CSJukoFQD2D8f1wJ
SEq3ZUKx4mdJPNmoXopWgJxKDxNjl71iGPCMzuqypSz1BaCKj/TlJhtlLNbNWqH63g3VHpOOg8IL
C+nRa3KB77fam1zhbdeYiBSRx7WoOxZKoWet5jws4SZ5zx3VVMDFTtkkXczufoDJ7xP4g5RB7fPn
1PPm+Rf0XuPdRtHlEy0NHas7fBSpdNZaPVcIjwMb25NiRG81pXEvmdzM0UysrqUHUto6kqOzPDgq
6MiB59tTfYdzbd0mlj8Sr0+mpsgOWBSGp0xBg4q7Qo6FwZV+G5R/M9JEbrWhFSG3yLC8uUPj8Ao7
6bt2Ca/S/Oi+Jbe/wrLJhmSHswDl9zND0ePpUbaPBN9JIAwfe3fvtNEUHuvAAV8DMuM7hXbgA2Cd
7g1uqOpS/utEKALqWpshSAKilbuEnJRSCylBl49e6IkiAV8d/kGOURwVayAkg+Sp+hUqQuMbWkVo
Z6XtjAOxzR5lTO9xunX1qAyYHWN/5Dh0WaA1d1VGUS1DA2Jx61kOIssClbKF/b8lS0JXkgRsyrBK
ImXkZk2bOTEgUHBfGrjeI74dBMU+5lqLjWHri+Sx+i0tpLIIvYWZjixw6RYINWy/Tv38TAqyNmTn
BHEGNKbpxTv9VkUGk4fca1w/8WX4hacboNHsLSuvp6DOWpQmuKmZ8iQxhQ09zD6Fg+l9DoPiUVI+
abqBcW8hv90Ho/gbc00hRi6vE7eJrNUQQjAlpDd7gkcPlTGSDV4aNbdLBZ9t/TJ+x5BT8zDBVVzO
EkawXnq1nBKcEFZiMeMO8atGuBx21QtPmdLDBAJ0ysqyn2VR5c/nzhrL77LLpXQUshibVkw9/dVA
s6cJWucCybCQOzizMzzTD3jouKB7izH/8KTaH26ch1wOx/mYEBqkzfsRkbGKgNbkPFZKTQe1G8pf
eafjjFAiPhRQ/piqGu1hA+oXvEA5xpk0BJFsEAM7Yyk31U5JhdTN79zA0U21Q8XWzt10Ex/AdIId
L+qZ2etszNs4ExHO7klVek9kJIF0ky6GkM2ttiPRGDuwEeH7K2oI6yWXcXlMUpY6kXpR9+dq6ymC
LmHzMwZDqtj2JK8sIrfcebojaMnr9bjrrC9QvCLvPyEZOy5MGIIMn4s+azFOgc/uMp6D/f6J8gIW
nXIxgH3YDZXAnsQqVb6yMvTZ8tXfzSFqglCrBAhGm+ru58qO4uezYBeM0GZa/17vPwUWdnOBnyud
c2E6aFvxIk+rO3vC53Yv3e5Qot2DUduPtQlSw9H+iht0Ytqh2JdKMjwUU/43aw3aRmcm/Eim89Z+
azL4jMzXfoDJzdQyiGUy7Kpq7VEpQrfMi8q1Gmf7CMhpsoFiSdQf0lBKE+ldzKGkPDV8irEF4Sq3
Q45Ul4elc5j+s9vwn5lzZvvPRBDao7hFxgZkKmaPx5e4Atpn6/z54A5Xw+I37jexq3d01i0Tb+2R
3USGD/Bk3lLt1VolXdo6m7dAB4C5Tt5AHk9rj9nKxrBwXsQ8+7fAWq5yco74EBRXlC+w8z/xWriR
TGuOmbCvKtgkKsoslwXaAJiqq3x2GiI1qqajO9VpJB3nWUYPMfwGOtDS5zsbaB5L7wJupafA4Q6S
JkCeFHjvbCQRcGwKNY/iYfv4Wy9WNzLebYOgsdiCOl99UKWS7ydYcv7EUhxMt7fbljmftjFidGhp
zECNs0v1eVGFGh1Qz6xt3/pVKvSyPICgGdGIcE229DLKlFapGir55brhWP7SZn/BEKT8qvdKF2FR
BWwudTcf6ziQuTgc71eJjpywqY/+geChprFg7xads9/jXA4PLVBlUMcTZLtZxNL6mx3blA2nvIkQ
X805vW+2oZJOCG+vygrtNfMetmQpplYIWHmoWT9d4kDi96l6l6fhFvvGiAXaDfv2p6rIVnjWZJMv
eOOpXgKGGKcR23pSZyc4cOKGVCxBcSffTTtoY9Rrp9AVvwuMy/zpI5t5BnaeNKflLtNtLwI+ai4J
FKCadFr9U9vC80FbJA245VyfhBX7HwlpPS0mHRjwmf4SkhL6I3ZTrdQ1vtUR6g3dVF3zWZY1zbGQ
NB6X8szDab25Hmc128Q2XysGSyGGNK3nZNK2q2uEvitQY2MzFF9qOAylliRAlI8Q0iXXvWFciz1G
6ZFzCwD0VPcioH97fJIPXIp7boPnnEZBLYNfoklt9VqFWT5OA0mFCMmbam9PTRZH9RFcLoquzh+b
7z6LTf0H4uct6JlkT+N5Odnz36PBDkwBirzOlkgG3qbGsVRFsXF8EX06KXiZS1JFUWsEyuBFjvfX
bX7JH8vvyWB0JN4D7ResOClt5YJYg5lFPyLWldZi6tTJd/QETmAvm1UJc4z4Nq54gh/WxLWQNgOO
x5YVhtpFBgCSiV1Dl4xsb3X8Huj1539YCdJrFKKXwvQYCHWANebZhstoAtf6tnEYPL4zeQ8m0o91
pBntgeEjhsMd3DbcKfc8vtDziUUSb7rx4f9yQoiPN8UbYMMLXjpymgBlSB0z/4Zt6dpp+H3kR3BT
yjqmIHjDTaMVb1mVfaWAjDIkXdo15T+YEBrl4qVXo2Bpd8elusty5+oRQIxX+FsVEXDVuk6oQQzI
njXpQOiFgiVdfqPdiPv53qn4aetdaGuf95XF46qQsZdWrBknLIxhTrtDtImhpE3sdb74ZQkXcUL9
Rit1IliguNEYPIXPodPDi5D/AaggTlMs9TXWCi1ZtiV37O9vN1EiyX+V8QGgAk7yyNrVN069me39
kGp0TXYTsLoiRUonrrh8NCpnFwMHFeGYIZNN1Pdypu5bnO448BhWp7QbRQR4fw4yib9McUDNCc27
cqFeUOPTFvRwfHPvFCjAL5wLSrlScFcHJ6PrgsIC6+rPF9dcN6chZ9B0l3BOFgJRENL/fHo1xJQR
sT6tEsFuRzPWf4XioMeH7xA1k8E3m6tId2TRPRrDrWPo8dV5BpdHNBp6XzAFg0PebNDb0NaQI1hM
vvLdFuKiJUmq4SuCzC1SouljCroPrScBCfUtFXCc4KRuPbq1aSaBjgnw4BtjnWRhNBPzuPsa1ub6
ACgcMeVqs4owFB3etPtXB1YHKCOK9UaK/XyFNGddchhb+VY3CfB+j+oydDsOY/WIAgBV3VtC5kkS
uMkCI84IyGxdkpuDfUa3/AnfkYRTsKB6OYcL67mIa5kYNRwsOXWWaH0txG2A4B2C4Q04e6G4MZbq
sSZqR4VEmuGyMP1ZmaYI89wdELt20Uv5ZAINXWS5MM4LRR1OuiNu4u6QaM3oGF7OPFXOnLFWU2MP
FY152pXhXnWmROafo0H4YibpQvoiGO2+n48M9xjxRtsLuO6CwhTkmeWHX8ZnGnttfVogB8tqGhFJ
JdM4ZL6qq7LWmFyZpMydlQr7W2rt30vxO0R20DkcLieOSzo/lzhWau88wSDcgTozkyeiqJViUClo
IEPN7kUp3UuIpIjkTk/SFfrJyq7P5+1p8BNp7nqt+J08quL0HndyOstFhY/0F/xVsRBCpI9+L6OC
s+Fn3K9eIEAH84cNkuszWG2u0Lw0iK5OhIKY2bK8+hVT5CB25JePYx/f2Bsgf7afGXaPRAaeGJAT
uEA8I/a8tSyupXlvba3mO3la9W8i2nfWyZSkDHkvK3mw5i55SY6o/sjBT9c0RJyTpqktD4YcVRuB
WW9CLqz5g69SuVcntfY1ZP+UUayPH4PjpvaoeYO9cSVX3Oo5PuuuIjNBElaYqW18ZiyBK5toDZji
tJZTs6jIzjgvzjiQ6c4POWxDb3CkHK22bd6SywIb5rFRaYDBGHiTKOHPo0lePUsDj3SI5ezgVGwd
BlZ/y24WjPNBtgYvhsnWv4r6vfneK9gDm651CSSL3DWMouApW64YkQ42+6mu9pGikCxwumrwLGAb
6SsYhOfWuS7RZxAcnFo9a+YaRVdRk6XcJLTUrwZUKrj9w+4JALkwjsHATtHCHFFFhV8HNESC5XB9
6z6cqlO7QAf0TkGLHQSCpSzJD/HWfhgqvqnbPb8n+4HAo9iVJjDqdBKpctPrCMPrqBQaNjtvRFI+
wowWF/fgnrH7OkgmQMn0BdA1bOgXFhKKxjoLX2RSy6FOF9q7ABFSSMqDcpaXlTyRnA3lxXvV3Q1l
Ft2ouN2XZGwNDVsdgeEs5gE5sJQ8NiFN91q/KBinyVXHniQQNFslnEVgZNJLWG4oLSGzkYlT1G0i
2Rs0K9yS5FC1oaT364qVJHMHTr42DnjJh4AGZxj6XELe41Lkg56kqM6qKqnmXtbLOXiUh6alKstU
DMCORv6wWH3AwJRO2EE+TUXZ+BkL1CbqQOUqNtBdivZGsEbTMCBdO0lcPvAdhj+qZwcLIKCgZ6jH
Yg3VMmU9SHjqtMb6qrQxZJE5hk/R4+gjOM/4+gFzr+XApcgo7N1f0it0Evg56GtfNl4PnGnos1Eg
oR/QzJCnYAgZaEiuoE6md0eN/QRHKFNZ/rIU0s5Qf+oBwaCxC420HLHICD+M++daTeXhm4uyz9pU
HJACnUKiCf6/Tqi7OsQYz+K3Q227shJ2baYSSnDp9dTzWCN+9DYIRl9aVuImW3w90wk+Yd8mr2O1
hdk6/54nOg5ihppxsFkKZkQOMIbNHtdVYqtTHWqPO8/kkxRwk7jk6NIkxyPaLa7j+WH/3PpMd47g
6NdqPJWsGt8ukAq1/ht2WZoFxr6Pii/mhGUpCa7HeWARowQfsxx/wNuBjUp8DF5d0hUnov5lG760
HUODU8JiKAn4CcqlNkxrS0QbQNiu0qID6YDQ/0YQXXK19Ed3HL6WK0GD98rGVBfWt9pxDF8SFLhD
NVvGs+das1eY1JTAU+oKo2p4G+mQW9otDPMOtst7DpwrgcuRoRVs+lK8+IiFaW4xkhLsRhUly/vN
J/cdi4/2x5WQZeL0Jm8PyGy6odlC69EcWBxkBVeJUEP96aShUcPBsTs2rI4Y2F2iS2QRz+ZGsvIZ
+3iI75Ba8qxf3tRizHj/kJeglPAGY/uUC+f3DWsbhZ2MMKV8mPxD1O1881FIR5h8ThbcBvLILLxA
C/V38ViIIS+H46WVTGHwBiUcu2zfHlt1pLOyjsLJCtsts1JcSDPoCiHRy31FyCPEIGQ2sHgri9cW
7L0Y8KGKJ5i6TOEp+xObzth/Tl47bE+Lw1M6sMFagCc0YQA6MDlBPRs/yLjklMqXw0hh2y0sD4zy
e+L1EtZgZ19D46ucvBd61eSxENtPmXl4h1Ctjtg8jVD5V0QE2zvRrv5jPp++VoISbMNDA83GiQiP
hX5/R72y/7wuEOr16y2MG9O/779ZGWtk3ZQt1kQSh4B8IyF2XhUoOuXJ4irF7A6gs7YzGSOccpQG
Gg8KaPpMELUZPtN8xuZXHvGqUk9BdUGvfQ3i7mxOaQuFjCyA2GwGTFQZ7qZ000VdB2IFBTaJqrJP
J5c7i5kYWPJVSaBT4s0PlS4VjZuehmfPAlSrlR5Q+6AbV3yoR3EHIGQ0TEFU4KeVaUS3gsro9/Db
oY0KS5R/gCquaS3nN04qEABbZD1w1ET9uqzXfiKVwkC20oG6B6KcnzygRxw/k5YT9RszCbb2Q68i
pvB54KOWRo3AZ75tmVDAoX/OQyIm230wWxNKl/ZiNJ5HJb8hPN+q8yp012gkvHTrFuw7z8xsC4s/
V+w/yMaoVLtYxyFfHRV87BMBfCRwZYVhxQTTrTRWyoVk4uSbsCLA2duZun5LgtZq9OLHZoJwmktq
0guzKyTsMyyusq30it1/fQj/SQcweSTjLxN0nHjqX/ElZjfdlKkKw+dYpHJ2C/mOzMdeZ6yRLJqO
/wDoFlIsxXc2ypHUNskLJ/CsTpu98SmAey6e9swQh6OCK4WdqzgLQM07yon0a4dNi8YzK/kG9R3c
i3UIwGAdlKIh+yPTsOB+A6i7JEQ7u2qYzWP4uN+5rAwr9tGSiSJ7zazlxOW+7M4IQH/keKSe6rsc
hUxaWCOO0sNiOA5av3BKMcYZ+dTX+adpDXgmqiA8dcKqlZLaDA7UC1uQNz6FRCBPOaPwC6f8NlBV
EcwuD90N8Ajit/FkOPaZGvNTqpFs68ZXCYMqzvTdLVGbNrDFvCv3JkHlt1DSo/45ruW1Hgi7a91a
0rFFKtj/jkYkmPYyxIfzPzUyjCDtPdQ9VaUl+zJXpr1RkBUnCFKxZq3lZF2L4CDT00xYbWOsvvPp
6IsHStaTsoQtv2olDLmIGqYh56I5Aeg2pzKEfwmEce/r+7CpguOPD+ctcTtnrVadW00Stn+a+5pJ
D8YqTRpb0FcVjOudpLeXKJB/LK4WqIn+YHXjCR19atGll75Rk9hRKh48jJKFCDbTZf5SlmtwwI1A
QiqfnbwKaL8o+Ct1LnlDeT+wemJpcBmv57QMgfHsop9Lpz7Rj/sxEmuiYbaPfKmZTiNMfOAxWxBJ
+DNiC5KI/2DBRAP3v0IkNWKLP2+P+ayWslxPpGIjzsipQAOTlRfrqyYlMZLQkvhrxwkIHl+vn7ZN
uDSsLD2ALXAII1pSJn6Ia0EgE5KEOFcrA3crJx+u4nCs/r02srPyZrPB3MDoH6KQVxeA+CnYhBWz
JUY3I3kOfhJVwLGXFvf/bN8VJznoo1LeriG8ET2BP4pJPf2E8dsQ69muLbXJFQ+1qAQMsBBYjsUP
pnZ+Si/Ui4SuM9NJ4m5XeVki2BpHnNoHOoX1rpRfaZyp2t3DEWiTB2q7fYZ7lo6sNcVL2oKzD7e+
Dm7BUIkgHWX+fTQVDD2KrbDP8M0v4rLKiYyrRjl2XzByPUtIvKPQ3G0i5f7eikrGbPfStySpppzZ
qA9eoxrnFZaZ7wLbIKKtZIrbaqS4yhDO3snoxgAOJJj8sSOJW/nuM7wlWacjg1f5q+qj19xTJvbj
Tu4ZvYVJn+QLTyfbFYJ3g11+irhQQ18GXPSHSU94hqAFisL4ASpm+4U6BtDMs5CJW+l8LQFz6tmT
3w7DpSG5WtDRVecdigEj/nFK41FUuvirV0IsQcRoRT9AOmvHJdrQQK7yugCiL4nwG8iaynZC2/zz
CBlIyeLWTbW3CDNx6HI9UNsumbkx+HDtUv+95CScKczx3urgiutiBoUh1iIiAQUW2q9SGVQBix+F
CYH5rqvWN+OB91/I5PNmIid/8JsrlK+aQ9Mcr3JHg8zy3UZez63CfD6t3YoJNv5qCg/BxhB67n3L
O8LSZ09nkLRdsy+RqzQKtB5uGwLm560GHZRX7D4M/7559YMZswtRiUAOPFcbueyL98tJqIBhGOfw
LU5wtPn1VVGAA97syVLiFlVnwBp8JSPWjl1t9iObhRK+k2/sY5MtD5ek4VBKD9CHdGLxpCDRnW5y
YQdMI5sDsy6ZdajDNzxqlgFythOuum22EMLvNMfSBjn8Cx/ZRH9babbWakSKTXMXre+qVm5om9B2
38LtICusQVfivlO/QCuCgHCIGjUfkxcyY3Vl//GR86dCzhC8NMCYXE5aQTMwheCSFphU2RMBqjf+
91PXuppzKUc8f98DInCDFmNtrqCSKunvHINmeiWj/arEv0LV7pMvx66f9CE7M5N0r3iP9Ue+qGLE
lM7WtyF9frVJthtvBvj8nBv/Act/yyvNfoEObgqYEiKRhuTPhAURbnSPXsuCYa32MhFKoJ+rwIHO
gaVw8scsKo9wyC/68zyM/Uh7bc2kFQEytXIcx9obmYyeVJfkumA53edmy16vdyhb4e8okPyv6OCH
3VUZHNKz8YskNpAYI/i2VNiOFKnJk+ABJcDNDFHhrW6LnbaTUq6uMDn0Bqpi8NAtrSWfXItObbEb
Fcy8FHIDzX2dLusaEf2lWEaWsn8+FtW5mGtVg1ocPpTzVyY2oIMljry8+oui7EkXZBPpxVJSSReA
6qQjA7gIt0HH0ceE5YlQL26aI37hZEjBpSTGU6BHDkCjMU+0nNJGeEEWOS4ggbU56wF0ihfzC8aW
HzeFe3pImhJAHLmujIgLV59JqUvC/p3LgG8Sp87WVU+6BOtnfbSyWo+mH2k5fkafknyqBw1sET5j
tVx9HEJT/tBKSumAcPR3m0K4sYXUbjOykXy8UGn4fP4kvLDDw/fik1vB4fPcsZMPat/tBM6GV/4R
asuZsUg5utbERCZW9/M7ClcHRWmpRAs601hoBTE5XR56AdjUxdlXeDxqE/nZioAi9x+xI0xDNxHa
qVpI4NJ1TU0JcTASOW8qfak0qwnwiiNNIH13M0Akb3aPrL8vfG2V6Z6sXLX8gT0Usw3qlNnryUTX
9QxIHWUkEaAxHF2ArF3LSpM35FlDaQlIUJ8aZaByQzBT7P71HIq5QEAiOizq1z1iEHmqWhwNDwwl
xbv5QoyBMC/dxrRiPTCKFv09QVMlgqiON2i97MZaerBa1UNhmmfYdd7KeLiF9Dwvew7XPdLFbvPf
xWyq3g4Ha8EoPYGVrsyVdcDl5UDy3fJdchQ9eft8FMBo+XWmY4FxnJdpnR1RwFXX7gT3P605Bgpd
RJ/MfZgV/5ApqFieqthFDyk6416iNzUKeFMC+wkVYs5U6bY3kBOlkj22VbDYn5bZDzEV2WfdNBk5
F18s4NQLjOt8jW2zgJxiEPVQVynEqy/jljKPGd99dCshoL/8OS1IgeEwnU4WQXe1ufBe3VIsd3WG
FjlzR5sFhVWX58dnfSDMLcx78T78GeQsC205X1LDbltBuuB3di+gj/om2WHaQs0X5rfKR+B6AV1F
woO4QXcZ9+2gXCUzGj26SzJ0tVO5urYrFMtxwZc12ievY8vQFxJWVQEnok5xIwx+bnnMXITa7TZs
Ude2CVb8dhjkTR0GJiKPXbGz2lUIlo9T6qcZPGHVoQjv6UvlYok8La/g4cryaJEbEmAlRaXEQ13s
PgalOzwxx/8ylD2aS+DzksBOf1hBizNVM8i7U8acRWXqW4rHhebIGkmwLa5rFcqFdv3QPUZ6v29k
GBjQVQoLOtiuBGDPo13xaEKo/H+CdMzBqzIKinflSjlkcJdbhgPTXelkQgY8yQ/aU2h0bkz2gAe+
sQuF952OOJese61Y962C2/66kTwDHwpVVX+ED7FM9Y7LBrrNY3Y7134+O/IOskU5fz4fFcDIhG5y
7wu+qwhgt6da7kBtQ9ULrvweDB9t6mHzEn6phSq3M70SFI1vrndYFMbS0+BJdKyhb6Kmb6s5/9DA
ATMwSSrBe1BGnoXnkKfbMXLSO/12F3U0CAiGTgFXYm7WkwwSaJ/00ZZCL2oB/O8+jd/SOXlZt7I2
JJnt/eOGPcFXODJck/JD2Vs6MftNkJL4VxDrxjWmEKEusIQ0/2AUViPls2y4k02xaMHQdu3Lciu5
AFbMhwruyF28iJfzwkZdBaa9g7B4HI3GAUiqmruejTSHT7x8lVDirQ0HOmyR/3gjaYNZ7eVd6SW8
G4WP47nUcxYqMOTQGqUkUYXit9JEcnz9aMbBshfoWilwCSNXcvY59N53jQCljmrTJzCH/BPYGGCs
hhNlu7SHAlF+YR8SuM7JMLTZSixu8KdFlVXIVO4cRLHWmjuT77YwvdgxFT/fxTGnQzXuFCqG/k74
4vC9DNAN3eBP+acZa+3gjJR2u2+gizN5MOKz/hsUxv7F6CHhZ+QiOqY8/ia7LJ4avRX5wVzeRpqv
qT2ie84Ne1DJBk2l8RjezgYqxP7/WZcD1hhEtWXtqR2BaksneV1uzYRD4PaG71F/F7BUZhmVvwGg
BFNfyiXlJQFV2kU9Bj4Rr5dhYPsD3etM1Z2ecScTDFr2enuVdUYNADisF7eGP6aCrNZSkYoIAS7G
1c1f72lnFdkMIxljOnOYaVBwscQZG2Z6TjDPEfw7YJMurSvgui+uOROgcRkFKYoqpzJC2F0YcH3m
CAp4Yx/WiyDaP8aowvOvcTkbpZ5iA1wYEYcDfq34pjELDAKargBX5SyRYc0XLUE2Sab+u1wXGfJJ
0Wq+cS7gT2+nLuu+nq1mFrRSK3VtFP2NWEXvXzTQbjK+uxqeXKI52LS38HNfoOjA69gIxdEZyewa
6nM3doa+yDP0SPe+AKHgLEaey42XGEx+PiwSO7wRR5GURKH938PEvOVVxQtPJGPP+Z2LPMAr2biQ
4e0lycwphad+1MTOykWdb6QoLUUtPIXHxO5kPR24LAKFDFKWIUmu1AKMx3NOPTdQjzfn6tokOyYg
UpK+E/dUVgTF4QmNeRBpV8a3IqILYt5pd2eIgcUhnYqaFr6oK9G9bxqEVWwrMcI7CUX++BmWTu6P
Mg7RUJVfLLOhZiD0ke9LamBZvNvh9GB4nvmRdlAr0JyTveaWhgNz+o/WilAqVF68Z1mrNLctokaM
dgvfkJe98QvfwUMnH8WK+ujOyc6Gs5o+n+SOT1WQJoy5uuTynNqWjNc/AVucNw7Ic79uUvxFSLY7
6epI2achJiKTP5pxYaakEggRxGyE/YweJEQ9nqUUgkIqWOTY3H6GZ83uTuKJFn1/BX0ipeNSVpOb
+l7fVhMQMIFOrXOlkUfS2bIHG02VR5E72Rhc3hRGTf7Cv8XrIYGd0srQRU34gm7cgBe6NQr7U/7K
Zjl/hdSnZLNcW37HGVCzw7xP67b2BywfXIC/XeuvasgyDAoOQr7Y0JQufe7I2EHWodYKozytLm4Z
Mrd75x0ufYtoEflDqy4s6Z3zi2IyHtLougks35fDn3hzjRS/PZDB+QO90F8fzQZ2l0a8ueNnn9Ib
lVnzbL2vcA9k6A4iUL8DAE1tQ4/wY3G/Ud2dpZphzrYb6xqpBlRfQh/fuKiGg4PioMbu1UMg8FGH
NNTAYvM0hd3D+6lhCPi1huO8Evm4XHoDAX1uCsjNjkoIb1w5JQWs5+BUuorr5GaxylJU4sZMW8IK
U/IMqZtBZVYddNRBGlWJdieg+K8ogfigVdClkLKzdrebGvMgyK1PNOTNpLwY9q+wsWp8jkMMgqQg
cJAkhJZMu/i6IFh8AyI44SXkU8Nfpk6dZghGA1ny2WR7epnIK0TZSLOCL31pmbBhnxFOatnt8C4k
8spa71PSMJuuD3jFqldeXC5+wrWBKKq6sMl9lLwlgTTDnXrrG2aQtgKsFZZ8dRJNdTT+RhVaKUcp
rFWVaoAj3jRoyeVxTN3tsEtZcWgd9cavxDjU0mumnol3ZkD6P1uG2VUukkb7VfeT70heC4KsA43Y
PClnMaUJH7UAnP+olgjE3Xu4l/OfHwE1kCqwt3NmrNKgVNlKrZoFeZxD3ZwA+J7Ju2Ah/rz1n/1g
vH3OpcAILz6KAq0m758zpjWGeTgE9CRv2/lBq2Hip0VvIk5Fp9srBJ/O/jQKtFnWwWE2MObLH7CH
PDSNyMeCL10N3jqTuUg9OJsVf2nEsMnEbKUI1XlEE5UaZc7jcIKHc3RBhYcdF1l3h7FWMpuIE7qi
IzCDVliaPkS+9Jg99sgAIJpdWZ/pJhzORV8vnCqFp14me3zyDk4F0wd3bUORc1zBCQ8xwabWqW9O
HMRyTceGFOfyJz801eYo9Zu0BqGgrGQZjONxOXKrxKa0CJgje0VUOK5AucGqfWPNArcW/KgKDklz
/2dv3S1MFfKp+UZFckvWkfbL7huZoEQMCJJ1EzJgnQ4bq8Gm98jLEvNCM9pcBYZYfi7/l+4hyJ8u
73Dkowh0d21hQdjIl9JxYiTAzKZA0qlvAH6AE85+pPGMBUG1/VU0UX146vNEDMJpmr87yei+vCea
XceLTXmTSR+ZO3qqHuvCHnCOYJ4ALnLkwOPFNzLIV7NkqjbR5Y7djMQuHpiZzXmCK4m5FQXJqTkp
qoAiDF8UvPqJHPQnSDDydQ0G/jAoChAoHDwA3jdTgepyxhwC2ozNqJCNl02vF2rP2TOPvRL5Fj35
89LrA4STt/agZ0Z5DIREcF8a2ku7mye9BFDhGDiWq6RfDAZNzs2+du+EZb0+FgYPZjw+4WzVigI5
ddLqhayOClmvO14gg8JlRkNSY4F74BQM/jZG8L7NQpOSuvgTEhPvQ3+kVsJdGNGGxcD1zh8FZHDb
+LmTbvWj9Pu7e7jOJxGUPF/hoYsdPi1Ihca0SyjnGSLfAJad2oU35f4S5269ovH7NSSqBCE0asoI
B4tiwk/MJ1SBSJuSbyz4/OAzKvYW6GveZiAhkCoI/lCuIjH2+CTS/wQp1697ViAN99G4GriJddzv
LbmCLrw+WGU1K6BJU5oIFWxOsG2qLBD/tKjchZR+Umz2rYk5M1rdrod5TNeUEw01PDapdchN93VX
M5pc4lSdOXgavDF0/3A24PTUkirKg4bMQ0u2Yvl4nRzX6xv0IEo5Psw56YB432hfiatMYz6WMUhx
8qDVgetE0/MLMJjpQofM39yaeHxkev4oUJdsRvmeCT0tEZKMq3hxmhRNV9wrV3BT2eVTklkLYAK3
VlHahSW7qkZJFx05LeFSY8GWftUgaLPMhm2qR8iK6JJdyHK0zYnLuB/RnxWPFKTj/Df0npW/ayPx
bsZfmNKTo4yU00tWGeQmVMEz6kyqb0/OexW2D7ENuIKSQEMnaC70BSherZLj4CKBD2vWrOwvLyUb
z9C9ZokC1cf/JM8ZsctUMJp5fTZzgcTkMhHd7FdNfJx9mzzsCXhG3OActTlmZkmaVdFiQ6aH0hjF
uQXCEVzkGSxSQ1NzF2sZ4D4RXyNc2z6i6CefrxWHl7uKxIIayW98PeT6PFhbUrSS2DyvIA1OdqjC
8czYUUJqhf7vi4ZX4bdc4iYRLzuv/DaBxqEF/3D4WQMRAT/sNTNtTBr2vHpBccCKau1wpHcDRXwL
hvJCkVqzPqUvqZb8eDx2TWMPsAsbidjKC9TURV1+wDg0hCll6597+021IYRUKJYXqjr5VcshMHtj
ENgkFlU19VWcT3XvDO/9dMteTrxTojCyofZXE+EIobg2zd+SDnLdP8nuNOZRvbQIljHgPlNogS/q
z2VWY3C+3NIAWcZDGG5Ot5xCl9jIxf+JDBayhRKNtvhbF0rbPxSq05DAWLx3Jd9yBBSwPxLV3Su5
zVIfI8BcCc6/cvPBOSk7Kr481TZgtYZxMMg6LPRqybRYM83NEx1OJRYZ2nIjSx+Mcf8DmT4+55Cp
UUR4iIYvQqTZLXjR5dMjxKUan9Ju9Ya5UgyKiyFaIk9hYq0DpZ8J/BUWWq0IBH1AjEBX3fZk7NBk
l/4OoRjiWDeP+AHlkPfuLflr3yLqL8qIAM10XoifGwnP+EYOuafKu4J809woTnWdvruAC9OAifLy
O3kBI7GkwQ5FLlF206f8MoVVspvwZB6TeCU7QLfbB91rXXmE5hgOcIFZeXKrvjgWsfaKyuBd5fwb
4WwmbBVxslDokRZBt6YipacFA4XvY/0d+Bi/+CHtotZI0s77D51tGEt+uWV8m22uI7UA3mgncfZ+
DoWAYU/7YMR9HW2saxFv0lGi0M64dhATPVRF/rY+U8yylxLrfmQ5BLnRJLfWM1CfFAbRVqMGPcHU
DAo3jDHExWhvo2MEmOpDPh+7XLVeLKux8WqcTiPaOpK5seOAmxVLnCeF0woP3J8inO1QPXwN6gWt
FnUQUVrgOY0fguzpbmJjn25n97G9Zj11rvjglXHgmjuVkrt666EHxUsabnB5fPjRaD/QLLY7Zayb
21VuAsk4ERmplaR49xVWvIV0BVB4Dk4yml3ZlM6NIvTOUxV5mM+tQS6/JJGPMO8Ze0PfIzVcOSHl
yt132u1GvRjRKdiVWIXiHlNmCsybqPuRwc0XZYjqTsUg+wtN6GUPUFZWICwAocZnsCBUVvevH/m0
5YV7zMe59BMXpRRKYuTWAyvKf73rMYHLtAa4mrrsA7k5XGAWo+UHWHV2uO2n9dvH3ejsUx2H7bed
R2YpImJWz7aVpfjg8nShA/VX4mTke7dwyp4dM7i0pDXkMuaD90+qADeRQPpRjm+dICdp4bT6lFvL
N8KpV9QPJZRXz9huQgaAdJ0AbjR9BgBcCv8KuKpKgWomIizzHybGVtNdogvcnSxuOTq5oRPwK4Mc
82ITKTrDX4y7iZT45F0sTVCqrBb8QrEqQrK+jV/0ePo/pYtjzCVPn7emtIwy2ycdIlI+jFMo/RYy
NAtoIjqaABx6aLJHFG+Pjj2Dpf8sDn81awkIpIIKV716kaTzvc5akOPEsAdSXdtunohYELy2ugm0
Qszu6VU6kw9HYNbVg46oTm2HJSPV4XmWBf6DuIOu0Lyeajj4/KevGr4cqWpRfRTL7xqYB3fb9oJN
z3UqzMIvRuQjiYSOWSwWrUQ6f3CDiJd+/6MKoso2hLy1ftFWOD9sH3G5EyWzSVoeJksVLK8apHSc
h6c11AvQL5SShMqiK1n41S/k21hc1rphY2m3MoqW3jElSDodT1qpfY/8vOn62uBYMswm19trD4K9
tcjVV5Izu6fXlW1KtI0MemgjwKSsMG10tYbLWJ3ZPU46DHjuybzcoNAuvcCbANOdWehqSyXhnG/f
KcOzhgFIhyCz73DqzkdNtk7m9+DtYc7wTdksNvlurxBKdX7L/0xZ/8HaQb0E7FVC78zH84f3S5LU
SyT/QAXdgaLrueSzVFTUKI77lnAZBMuubIOFVe0U7iR2aGK6ipm4V52+gACNcbPWxqVTUz8awEy6
/fkkFcUTt12dLwPUzKVfpixafT1pT320JnhgROGbBdXOxhTvxEpE2/1euxBolbMQ/Lov9VwQldQp
vjxwtisu+q/i6ZkrXFNmjMZLsrK95OL6zTkdZMpdbKY2IGPa5sHhbIkJad83pgB9JSVJCKhIxfNm
6V8SpSm0acgHMPbYRtNTXhMQCZv3ma0sGwveLNbN1offo++NEcbRNiHcxwZg6Jpjq05fA9W1Brrl
G3MrPSO99lGnD1U9ZfpTHdtUo5NLy+hz2kK3zmu6OZfCYQBVVPYI/8gUas/FT8IE/OwciInRFErA
kFJemJ4NKdjMjKA6b8JCAQo0++XqUizNCW4PL2kZ1PiO/zGnDwOYLBp8Fz3H2HZ4BsGxpZ8+mSPo
IcUZHuOukXesOsg0r8bSpEsQ/L2renPG+3rasOmACiyRPH4tDi18joZ6yg7YX3u0yWzr8dKKg3Yx
BoD/EWCjvxPR3xlQ+JuTUsrftd6b2wRLH+1kKkQW1rKH0XsdVfi6WPSQktIcsMB/h7skG/x47F9a
FnjDM0eGp2auEgWTQSJfp4c4A36HdXT1IUSsUB8Pm1rsAscYPkTT6wuaDjEcgO7xXMlGgwWt8Pab
VVGK2TeA0rt+9vu0n+dhRYK5gf2uH/pHGMaKx9U4pTGaWdk21xmnLJCzm3s3dsLDH+uHPKP4auKE
5l8Vsgx6FX51B52frYyTH+In3WvIUBXg4mVbmPR62C1acYpucI8+ncJMIW2hJoUWMonyWDPff4Aq
8vMWfjOba3dGten1vvI4NmQWxG/1ruI3rdyjLffmjan2WLWRJCeWMZ2QiLAVNwMupmBXtDPss68C
TfGtHK2/S7A4a6Q1OfkjqLRG8UeGBbnx3JA/HzSRnaiiyL5pfz7nfiiT8rQcNLNA8wqrFld4o8cM
yMVHsJUmtenKCNcUOs1MoZoTqJpFVzf6/d8+t7VxmK3vrfrAi/4no0zf67z1I9GfSiizRDBSWNkh
zYC/CaffXg2Pnh1wQfYMU7IbyT5hy5yHZzUbHDAdwjFNCLh8bZzv1k0N2C+RndTaFRlW0uURVmDf
pqK8HsZLJ87InYjcDejp5Bv/imdmzqOBg4Ox4lBJxu8+2pHfR19/3FA6lvbYrE5FYzb3c1D1xBs/
+OcQIZrlthxOG2AQYYvOnIfzsY5b30btkC0gbWis0+i++f0Fn4iBrVWdkYClHOLj3a9tRPQoV5H/
pJ3AozcZbG9FkyynIG+/hnC/Kd6f7y0PAZv2wbOoJQPz4o6aANiuV4F92j5TQB3RUzHYIl+DQVR0
sSQhq3ofCCaeL+09plAdecr9D2USdmdzJTzFMdHxLol46Jqmop3avHeHFeYPo4Ey51IScbz3kdPF
XTwOKpx/B3AfUDxdkua9M5hqDK8+dffvB1+bGyA5xs+ZVT2DkyrzFdnd4ijuyGdpYK4v54/uUet3
E5lGg25LfcfTQW34tceiL5Ms1Vf5WZ1CLAFenXFB5Mr/QU7VGB2j2EJL6tugszTp5LEZaAUEi0i2
3k5s+vjkacUvziXx4ubRfAvW+Nv0MXdo6ESrvUBf5W5MXTbzn+JhOXfYso9cEsInV1JVGYyKNCaW
9Oh6GSB12oGjtIFTctqYAh1aH3GOMWUjBwt3xjjV/oimHrDIU/3z/w00jIBwriC/bfjF7FGa78e6
OkxTiUWbzk7n3H0BMDWdemUkTtvs0hEklVd4ru79B0MS70pMTXEzreA+vOGNzBlQX5xaLE9HW8wM
1nbr99E7BuW46HiXqJZgmWU2uynKvrMPPyRANtF3zQBI1kEd/wc8SKS8s4R9R5lSNtVkhExJOZMj
JAfFlRgZuzAVqE8/ROAXNRCuVCCsU8oO4nWyqjKnqYWRf+ZXH4G4hwrwbAydYRGFIi8al0Na43dn
Lnm+kxuRPDUleFMw1t9/8dqrvhwnyINMBzgHiPD/99WYP1ZN3x6gP9XvioxFaugGL5kuwHLh/atI
t28ZoNLiYOHKIeoVgc6/+/wuUUgHHSPOZ+V0DWdw8JoU/T8+9RyqIZ4hdLwXJ0tZ38lydb+DdvEX
FjoGvRmB3rIXxThoqCeMCu6IgWVa/OgX3t0MW4lsRZlGeZ5MbyzQzbn3Rv8Z2KhvJflIia373T5Y
3CVqZEtfyc4iLUeIo1kHbTXbYP+OWU879+ELzwWRVqWKLHnqaWM63HxBDuXCaDmjZHCK1TKKoH7w
QQz8h7+WpVnjoVEOrXzJWBArGKlcSgUm4xZUy3IpBxcNiTBFLflJmiGwgtTLQRcyOu21zAUUaEnq
dqWMCq8fbgx5KeMW2NvY1IRwfpNMRqBo8KFBfxFggLiNEuAxbn/9ls0jH49/dV3xbue4vmBhq6r6
MEk7wFtz8Ql0pxYVrNLXdq6IXk4xoJQ/ULNtQEdYDgLRLaZCyBBkdkYeaN06kfRpRTI0r8rPmjf5
zeMwsGa/b35wP3PxoBYwodU0U0yGJhYPl+T0BU06NIzR6H0xZXfpxT7Xg7iS3MZzCgJFe7WFagub
0qqdq7u4Q//ohxjvGjyqSpKBXSYfFGPA/QLME4w4bquMLxmFAJ1pYtV5ZwKuZHSlDUKavOM1fOdU
0u0eqMq+xrf+mexX4HsieZVzV8Gc+q6TTVrSXebNYP92/HMe99DrRCS1bBTXV8Rurlef0YR07NPJ
8qphVfaR7ib3W5E1rozeKRA6ykp/L4IWung1oNnOCtUeU6VBNqhzrIOCIGrNM3rcKvzLOVNtjMEy
JW1XBVQjAtjbTsfzuotFZ9LQBmomTERQOTaOJTSkKtcFYI2StDUw505gZmPTDbZZjNDccGWX1+0p
fCKzs9aysgIc8Ag7kx57hTh1bz0ja1yqiKfuyrarjj4kgUUBdmjqBbx1U3vFepWt9phNv/D6tg8Y
JWy0arhxoSpINjKSBPbvHiUzry2YVaa3XN3hkO7+f9zsgpXxmJ8Te9a2kFhcGiXUtBMo6iHBCQYS
rDuyL3j7vNLWm/2Avjz9wOLDuge3h2tpoEegm4FXaN2GmYcu0qPTTddX7470ye6wooMoPC5ZZntW
q6AwwOIF9cSimLF5CfO8yM00eutIv8E8T18r0746nMF84/6jRznpIlgP+OVkR3ANrxMommhLLz7r
VOYA6+DLS5t7pp8P+Roim6mWD/TTlnK95jmZy/Eb2uHWdK0Jlg3pYa3Lh71M8CRrl/JP06SctmXD
s57J1rFyi69ekUFENARNyZz/xnZl2wG4zxGknw/MxOQG7h913XzgWcXPm5PXnD3l9+K+r0Ci4v3w
dway58Aox7pbujCiLClG3SuXOMzZ51nMnj37LjacE/nxUmAiCbyZLxuUVNXpoYIIkAH4U//S+hzL
xF5hqSWR5RHhUwQkr4MHIPfppvgyNjvGPmiRDmkSfAjA8L86CorH35BsJpLQua48F0Fx4VQqT2sU
2T7iaZy1817Q5Gm9KVQxLXVsi1rFtIsswnzmrTGybo/C5aEjgOfidTRfh0zKLar2ajyGKxidntTV
Tm1cgSGBnEsRXwauiCXEF5OVU/lhknZrhU8j6UtJL5N+wUcairxac/InF8tl6y69Tl9Tz9+DwqRR
4rCIRLYM/Swc0aycc1MuBQuPCVhrRFOhxRsnqLr2uc8n+GrUxa2wW4AU8dWkkr2kWllgRMwo9l8p
VC+tyd3lyFoYQ7THds44DNjAFRoEgrsKpG3TuzgYLcHmBlXTznOrTw/PqdEak/eUAvqsm97M5+3u
RoIz+sA3fnhOpoRimctzQ0DosUn7DDrnFL8El0A5Ar/hJSN2bVk6XPI7XyZHbTP8vkh86cdZavSG
+ueBHIaLx2yscANEFA5qKx2F1RcOlY0abKKxAAKzDHxI5nMZEnFG7QsTRIp1sEihSk+9di5EZCp0
x6qUOJUDKJllxlEX2RRILQx0UdnPtl/vOz3l2b9UhEBlTUB6TER8uniWK8vKCWEi7mbcO3xCEzhI
xVAtvLwhX05FVhswuQlbPHCC3T6L+4SvhJ97ilNimFmfRuzISAngU94MMMvcbx3OokzPxAfdQWbq
hqw0OmZSbUu+YeaV+lADCG7+FewR/+7hUps9BwQVVZ1m19GCZgiDVyIcrSvmu/AENk40X3vFH5ew
KHPwjDpULNBPeQ6QUXAJOPe14qEug3jbqt1ogmfupZBq6jHtbd1/b8A/mR5URUtSeavqmNyJEJeS
fPUrCvPsh3v0n9IhxEz/xdmAoEXw8icgXwY/5o279glsvLDVXKbBS8WBG0nquWY5Y1sNLtUA49iy
nhLeBQlwXqYbB7i0TpMe1EHpF4lodUMpgT5owYIisFbui51QuMetXoNooZtTebDwKlziRBUGz5zF
SKg73emjsg8Q/xxaMkkm2B6ETb9c4T36yGFFi6T6m4E7yGwxQPMuQIU4E291Gbe7xlEAGaD8LTpH
/FkRhqs52LbtHq0JHU1xFLjkQBKtvscazXAK/zGWkCoVa0uFO9fZXtOgaifVicYvjTFW2aKcMzjD
bweckY/mt47ezRQp3dq1hQrRKFTTJi+79ST7fssHahIs4xAHWs4zC2QOy56tiSpEdFzFrt7y9LP1
gQ9359N4UWMBQY3OzwTIEOplBI4jbvw0hONQvlWk8QoMVnfm7I1TGf8bj4PjL25ohEGXZ8buFb5e
p6NkvhKIkEXy8mxAW+ajW8iaDyPBHReIwUKUunHQwo3qoWFMJQ+b1IitXAzy+K/BZ1tbaT/iFDyL
7LRkNb9nGjajPNY6goy7EMUJtTpVYnHnra4rTYa9UtPigDS4DaX2VBqxzwwfBEGbp5NL2+IkEy7a
7QR87yrviIQiSdcr9hU2jK7gXPPwj4snKAf+Shca30LL0e0s9zduUi8Y7ZYLDwtlh/Y/1zJqY294
2+uu2wX5na0r3ua/XIClaNOscn0yd67uTcYOPU44mcr4F2krAzEdFOKEbsShb0tcvorQdM9cG5I1
6SR4MghJL6mam4Bjhkpppx2ss6HxxFWPtLY1sVjiwGf+ahIhpswOJpQ1xzKDmBBbdn1b7aowFbtM
k4xTuQ4+fftOds/fY+FvCqlrIt/VHc9o9/bWdQ/YSOS7h/ec/5R/vTpFH+Yu/cSkzlKcjfdW+oQm
oaH7tRt8Yf4pnRKXrfB9neWf5pWnLrH9lIHJ8Z5cEqlSf+1l7rjY/aB02Q6xxRFS0TuXxOJEjpYH
jpRpE8SA7aAqbARDMhbMXBAV7nKlosL4KgThpraC0jCt9m5YxY8OZfQmLAI5xn9kjOR7IrfwF78Y
jvXpAsV3cfvk+Ucklq8f7shFJK31tCesUx2pEMBNlpLnmDyH8tuo0yUCj05gmYJAov1n+DfMZAGC
IgWdj67uqsll3s5wjMrrtnutuKaxRGrT6mYe7PYPxm6SwiJnkjfdwgnG8IIY8peFiBsHa7DAIINy
ZHtIv6yaS0N1Suxto/AAgq6rgUTKALi4ETONJ1Kq1/YLqUhnmq6QotqzlT6w5RP5XaAHDnrAhPhu
p0WUu1HYbA7BBTypdPN2Vu5dh4+XToCzca9GWFU8sBL2hqI1cetn2pWY593NNJIanm9ldfUgnoKA
KPoLX8/XR/P7XXHpJnqhUakwhsIcCy0g8ZfkZtRHJKJjOMneNAe3ztNlbjAovh2S3PN7iNwN3lse
NCZLFQHe64BWd9Xyc3koeQl8Pl6scLlx+5KTOO78WOq909QQkCiTvChtKwdf6/G1qIeoYVh+0tYS
IOWDVsIokxuW5WcyVWdvUSuzS7VMotCY/+ALyMNu4zh4bbUt00tT0F/1GTvfLcUVaBQ27lzuB90d
ghJrIvy6SdNZyZJ95Qrqo0a9R371bJGxB4bJECHrK+Alft3mPch6ZGo2LUAZJpyyp3VmN+n471X5
GlOCHny6uj+zvI3W5QQyjnAW/2nDS06Fx3eVtLIqmPbPnhjqRKKWrn0Sfk9hj0RGURK56g8Af1X9
ZgVFtE0tu08T7bnDRXRzu4j/1VL8bjoNuxDP/AVSneFY5e7SwSPDwszjJLwKacQeEdfkcET7bojQ
0H/IHMPAQZJiFL2D459Fo6x6h12vEEnSQ3ANZaJj7GznupaKqFg6+5jPWg4QSG7EEUc4FLKIRwEY
BBy5KdetHEf1Njo6EUfJJFh8hKgLEvN8CJflDW+mw65jGLaHUXwAiR+XydFUUE0/JWfsejuP+ze5
9rpGfcxd82tPuVo7QYnzV3rAu3BF6y8Pso7numABTiTC5N6mvjPvGKHevn2ZjfxLvDpsA0KKLRXh
0NAqmkx+ljFAGMyH+oSTTb4dhaMYO/v32LQoiI4lethalkOfqsCskxczUUTrge11J+3odJZfzk4o
x7v4ciVQGF1XDwXYEjkEXJI8FxMH1zffClHN/uQJy219epvzsFcXuZzrNDQMffADbonGKLGjOXYi
KcMddDGu6Y7NRvqqZ57670MbVppwCh/7wJhG9y9/4jbTFmi7NJBqlwpH53bWivZxETiNEforyu95
yq2mcM8COUlkY+YYDDm0tE/f3oWszxD/VDmiqoct5Okjkl1vXW9HQx7LsZmCoDunCBIpjK3wx2Q7
tzg2iH63oRYvjYgzuNSOXpOsgMWr1rDumRm6Ft4RxV+qKjOe6Eg9f+VxDjzuC64C12mdrNuBf/ni
peT/UebvxM74uT79JmRIbq6LMo60PVNg1zTn+qska7ll+GkTc0CMPzFE/V9pZVUpf8K/07zqvaVJ
cuIQ/M8eIz0M0WE+XoExKH9sPxT7BpyoIpfnPWinn0AQ1ELhZVnp4ID9/65Dt9hejUX/Q8oeY944
c6zqFVKi1O+vS1ivappa9wKdILA3tUewhtX5X9uMfGiSxKEYBRx0Kxy8W60bp6TNX4GpWmCqP7O2
eLgv3ZVvGNYdNdUEJXICDCEgXDuXq9Pkhb4YMq8xWY94fQhUMewiAqVKplVO8ZRUjv2pc6B6JmRK
lYZfrrDW8Jf8gdpPYCnKxAiTinknhLndFJi/OSemhbyhZUZf3LBkSJKt9CJ1sqkda0IrmF6DmeIx
hb0wGVe6AUhInNNWuiUDTYks5Dt2fltK3eeXIitfzLUh6T3P6UISBME3xrOl/Nk37rEKLSnMlvz9
nBeG+jUWSecXrjjA1w0WQk59EeO3cx/aCI7vXZX5TILdF01sAyL+tcQlblttK5F30TBTnKuSQ8Af
zEux11hn2HO3uSynZrSQCfpgLFdsVTtW24cxlMbJ/5K+IRBXy3HEv54eZkcDNTGVX3ILmmlHNRTR
mDnMSridhb6MEv4Nbc8gfw+Y0DKv4K/JOayeeG5rtWv/jX0Ipu/j/TNS9TTAVBqEK2DPpyowIqYx
hTbg1DM/QOAIs+oaGiNsfSQ2MJMX01ejOhVdt4zDuHD+95fMNO/VPOEY0JH8oAhuYgGRAHHTxIkH
0ELYJZA5deTVcBkYqn6I+YJyVL4RcUqVAR15kkpYERyauSGkZs9hcKajMu+oc6vRH1OInjjrFYlZ
I0gyjj04zd5ybwz0xIjs4w3jCDdQPnVo7+zLUj1tSGVDb3dHKHL98UzYbDOWjX7mzHAKQKLIoW1O
/8qTDLlgdBk6avH53rmOdIwTNBJ0YcrLUMnnd2qtXgELwwpYGZqN9kYe5Ep1CgqHFgce4sowak8N
S+wLkDvGTq0wJonriMmG3Ydf0vIEQVXCcyxvtU+vLTwppZtR4Cmq36cObHiQdMn54FkFSssqFKN6
jo0VL1lnZsYfdhN/jAcGuiQ9r1J0KeE6zhsjwHIX2pCnKaRYbvrO0k35ECRIDwL+LNxBgBzW/upf
iWBWMwaiYyS6vEamiELkCxRC+mTq7hUZacxM78I8Js/9/wNlsbvjs8qjZNBXKGxhcrJEwfZ0NyhS
QvNg2NYGk5hzvsRxrVMHWda4KZsTtM5EoJr3M7x3JYVc+HvzL5aVEJo1no8b/lbqIkmbk7hWAPC2
E9+CPkEK0RwPB8mfGVL6doOsvPw625t7oY+l+rBgY5gYM2+ZYNtEcP4X1sWz0sOjJfYAkwJAhVwI
SqTBMx3/k2o55Oh4qqA5NkFhRL0mlQGtn9bBZxoDKIcTEHHPDKUPrrrXsk9tgGDGtS7ClLDH0vKN
iTztCbGkn5z2f2dPpdGnbZQsISJd9P5hJR+nN/V4K2lHF81EMr2+s+VOqiCGzjEeQsPkdxDTT/KU
76lb2kapz5F88vtB9tLoL9pcn22X3bmgcRRDB0M1H0pw8b5Q487RFWfhQtOba4UOQXlezXbac268
8377w04HMIJMvKkxSkDMOipQ5ytgeRbwcP3Iu35fXfMtlWL73COmL/f2sucJAG6AggH6OZ0RVVQ3
/EU/J/1SAoie9cgySQz0ykD7fH9A4UqdSLrSe7oRvYPEJGFpvtGGIzcRMzHgWP57/95snbpLXpuF
UHSribzoXd8uLxRTQvWnM/Bre4tmekmkTMLL/3wbXXzsDxn1AFnmR4vMjAuW2PyZG3LTrXH8jUve
uHpAjuoM6qW+11HfTAigA29PpSV9v/5iV61GAn33qAyfA24c4SDUHhda4GO4bcSryr9VuQY4L6FC
VrAvLeCdm0ZBeJZB/55JzzZ4cCWi0H/L3Dyedxq9nvg5DFf5IcwpvaBmtulVO+fvBKJnkehyfqHh
fj2zcFoWPtW1hjTvPKYxQSqt1FcwmTf0pHLjUH2cqN4cbwnDKcpIurSkZPAH/P2MDSJj2dW1y6N/
qxQA+ydqo+sNUcb9GnYWDeCRxQ5UNAdj2qQwJLshMWJLxyoaraJjEBBPXBqAViZU/5vNk92m3pLI
Mo5l0lKkSPJ3Ac2WnfUGxym9QhkaWD26fAugJfEC/jhhVCSIfAer0zSX+flGDPns+lJX6pft3VVn
6uk0ClwAYYweGU261G3bylqigjV036/gCFm85fuDtRUxOqyXpCIUl6Y+8/C9jjchnTm10qvyWCcu
AMmv/tFF6rwNYMWDxfcnXSfLF6897Gpm39J6tZfefx8NpaemgDiZdByrg1RjZCXvKvQnJrZgVj7D
sE01CF2Jej6kfVyBNxF2M53H4HBeBIGK7mvcUAA2zJwdmZHi1wr5QTMzdZ4S9A1zcb9sj0AcqW3r
qmgbpqTeNXNUFDxj3DC9fD3JptrTfiSPF3r+YkmxM4vl4SuSEa3cgl2714639NnWGM0ga/IAezKR
CIuF5uRGrg8tdaSmoF9E7W2R9ONNzWccz4aTEeOXmssHOwiJkE5zn7cgwUCWgzaVYkOrPBDuYlOa
dv3AZmFnmr7Amxf2Iyv64BE9cl5pbIfjG7+P1kGiZWUHyCr+Na1JaHDh6b86TuOxIMvWYIiRUFz+
sIciQO/QHnm8Zv72qPsHxGEIXsb/lrym3CmwMxISjCyHqpwVDS72uADUGuLwowhy811dCVg3o5As
zM/Z/8WVyplLy9BlmuuV+sywTbOMGtjdjfF7XQl5PCDQvcD1U9Uy2GNKywX2MnMpXmX/XmUay3S5
9AfitdwmCfKHkVScOf4cm9y0mw8Uoc/RM9pUkl8wYWFQsvt4GzG34+TRTfzKjGC4LBzqtJ0cjBre
XK6gCvo5JzZs6U+Ri5n0taTuftKqy4T84DfXgw4OOueaj37mT+vBxHfeHjx96s5IuJjBqmF2TI5B
+hE3+tXMfMOy0EYrZhCqnK5J61iC/I9xiB2/qcJam0kK9OWJn2qSnLSy+h/IVdOOOw6q8ruYzoec
SeAab8086VxLWjhxMn6lt9CatLn+ACvAqUYa2JB3/zLxLUGQFdSwD4Ri0HN0P7Gm8Y0Myn/GcxhV
YsBJqx8MgDhbu1nJoTFE7SUWoTTKKPv3Se8lnBCBY61iY4w6NGV6GbXThkA69+EQHH89eTxMCXBF
N0lalfB5C1nqW3UBDqWwzCplN/jTacLC13MKz7u6A2CkqR6BE3PdC09aLNWucCRdKqoC6EAULKMK
mJ4EO1il7ZsvhriIhQx4WLtQSYTJD6wYlBU97gkhcR3XDkX0d0joLLZFKCHFRcmSPk9PSgwvguEA
cByuecYKHoNCBTrQzNN6zAA/6705tvrhRDTYhJV0x/KCO6uTpn4frg8cVfCzTpDWD7g6UKImujDs
61fiu+JWM0TminPdazc2oEfGsBAb3KIxwenhqFm54veGo+z4N7aBwugiraBmNjCZhqEEeitgglbY
2rAZa7K9/oxsm+yz3eHarKOF2IzAPpH4WltFyal0ogtNc/yUFM/1AmHvXzQMMmi178XBe2f1R/2R
9x0d3Z0X5VBy1y0sBSUDwsoPKO95rrs26TTKkkyETttEZ5EIMAy8LqdmhsuO+wBCc6CtQJ9/FL3S
6pSDKraehWsWKgtf+DNaUrSGv5CFzQatEoMiSEMn/Rb5hXDQS+5ni5Uj5e2X3LdCn97yhViXiB5r
g0NZ1DEK1NNEs8QLhbwZm1AqMELexH9TyOJv05GMwSOR4pYVmcqp4QtvIGnUD7b1aN5EhpEd++WF
+/Nc+FyLj3FgAGgvq4yZmppfsEj2QrYxD3oRsSiB9JPmxfBU3zdi3DZu7Za0Wx+vVS9oQ4wYMpkV
OiCNtne2vIkBHvjuywXbz5TmMW06oJflrg2E6ncI21zwoDbNxukJrj5KHRtjbf3UUcVBtos7XxV+
xFdD12KqDYMz6q6Nnckqv+SAHegy9ljwY3WlKm1kkVVku35ijhvUKf+19Xq/coavs1jY/OqunqNj
4qI0Xc38LMZQfEybeEIH4e6PoTzeGMtUJ9p3cwngK2tWedtSsgFx8m0F+QkyA3lUyOqGTZBH0tIY
weCqKPpTl6cxlglG8KsKQWYCyHnmHnupHM7TApYkqVvGJ8tmp35CVE+ArkqmZuJOOF7wcAZOpF9q
UnklhJvnunl7IR0Ti3rLMhi3tpYG+umHIEKhHxfpIfHDzTqB4MUSK9RGy/FP1jFQT1x2lDN4W6KM
IHzOZFpzlw7rEKBg/WFfzeQl9R54eD/IDRXeDQwZKXzI13bdRJ9HbtKF/5/0PDKPi1xNuVc2MUMR
GsoqqM3alrbFiCc/zjCbo5Bq5ZlHuEH4K7PDwBJmpNumgAF2qU/x428/yhw/O62lEUJULC5i5gw8
vIhCd4VmMjkhLZ01INtftIvTH86GwD+huwCADeX2gN3AkvwDYG/jvzVRIA+21ksNPh+cw39cBshR
Vu0zsdK2mq4+P2OO+fw48w1lnIpIraP1ZGDeZ2B6yP1nVSqFHSos5q+kEa+37regFvrjBV4xXwDA
oTIZiGanGs7JCPGE+z+yhtdrTFTqtmy1WNtEDAEXktspbvr/my0npQRCcRclsFJrO6MYr/kw1LsQ
BUAc/m5ljzf5Xz7l4iqniKj8SZS64fURAnypOa+gwxTMmHJ54iVL68wOK7+QiQlNGQuKdVD55nrt
/VNAfXIY2imU3tne/vUA4fo7R7dlFswqBBaA/1vNAyWYGHJ/eLeFYYTUxfg1KwLKo8oDXJbxx9wQ
ujEZbTVuVksW4WanZ5hhnGKPuh1ltgWNceQXfEGnWRB/KfuHfGjIwc8gNW+v7Te+MuN1zAWajwqI
jlpiSRFcLcIZ1/HgG+HvRKqraHHPhURuVQ86V1f4D+J0hep3saGsKiWCWlkxBLFRsHds7vtPJ6kt
SXk/gswIxRIqrqLF/pUV1bMEf8aWb263btlWuGoA1zl5cOUGoZUEP3t4BsYAiDggmwu3cZ3y3eeL
zZzLe9ByMeOwAfwZcpojGpm+1K+GyC3kM85m1jFhfVV3lxOrWPTrQIwyGb48uHvHMwhpj1JxSmuy
6Spxf1INNReK3IxTI/eKGJNamSzt+29vOAGgadEV3Zr/BSfmuiz/OQIbs1qp1vPeYyujw1eWoEgV
wW1oAaX9chLXzEdDgMgSDFgLfVDPdiU+3it53fM7DR/2U2kjFbn6VvGnfBf5tNS3FjiSSEH0jpKz
534Cu/T1bB7Bjwij5ZJEzBxNwfZJWJfSq8mPRASGquVFTjLIldsH30yF6cGHQFiXLIyQIYROr2M+
Xn05xNcM7deT1JOhrHAjvE7e9i7pr13XNM5FAB1juteS/HmJbGVuPorCqbFR3qmhv/XYQjLsUIDz
LJvU5qPN98Yxu9g34IX1ad9pBeUTk6cTwWEccK/wqk8MzD6CFqBmuZ8TrFyog7mtHxtHzXofbOF2
k+FmeRBakU/9A4E6UR5snu31bK0rfzeHu/gcNXTNJFi31n8ZJ72XBF9ps+uqqgWGbMfYlMhH0hio
qx7n+u6bCa0y1dGXKd3soBJAf8ZJaQgLrt6+py8nOXSinc2DfS6FELChQXsffHIjjEkwqLPeqijF
hhlSZgTsOxH85zEAe6xBCZkjzGA1lYRhW8T+HoPTKT0uOppErw2sYhnDigmpDph0bkCCXdvl4Iu0
zEthAHmA5EG4yHYJs4fqMpekvJZHP9EgqWfs6s1s5wzP6C6HIZf3SEpGPPBD5l7Jodc75DZuBZ05
uRAbkAh1dpgDctRiOVVcPjBCetEefIH+sAoOfc9/+4mSqolA8TjNDIxwmU1pFf8fSnHuv37Xz5kr
THzNAntYKii43EduErT7MLCckymdQmlbL/q5argOv6f3hfsihz25pchEs+8/yCcB5Dvi3pn9qvcm
K30nVFwupunAz4Q8otEkwgUyOjIyP2eufo8B+um0K7qnZHWTIPemvNyvan9/EA8f6HmtyvEPFTOC
KBWRW/mNbVd5o2KAMBzGswHTztFwLH4jgyXkCuQrBcxcHASVN1EvqRxpbSbjddjgOG7Zi7p62eS9
q3Ur5FkhHdGXr5hCnN9x6MEmlNjDGOYGDXPVDurxSKST2zl8zijf6i8JaKDmQF7GEdiMN/WNB554
TcMgzgCqfi2Llr9qG7agUssR29jy9ktWOgeMH+DHmbxjBgFZjyfnVVmbro6i1/ziBIbF3mUhM9/Q
LqJOZSKswUX1BlYO2LJLX0HKrzh9IyJZaePc6uQwPid+qp38D1XEfUT9Sl5pXnlYJ8rwJuuAc+nr
U+QU5tHWYIcvmz8q2XB0jqfeb1L+WMm7LJes0FWTXexOImpnjDkzsu6snudLCY6YQMaplcfzGFEQ
sbXybui/Efmv8sekvsZDYQ5HRiYgeSwmASSO/jDCbncXXqxkOs2GmUoaG2X0pjgsoRw4/TkcsRyd
WkYhyKCfeub6RNsQM+QaJhLAzcHlrc4ftafjjB9VLNFsqQYwVJ0HM6i2ou8ZqRwahqnHkY4+zpUj
EJmsGIR/Jy7DznET0HqCq2O7gNzKBakOZfnWZQc5UMmshajyGvB3/e0XvroORPtYbIsXnY1rXVuX
BenptjRG9MFYv87oZybKaVSMeKzA4nxtGlNO5FkLGfhtwOyctKcMh1NnFxokKywKYgoTL7/hbwVG
M41nSC6pze+ySIhVfIeRbiocqyS0sUbYpFWZXZvPt55IOGna7Jr4Ov8zSu/QtI8mq7bhn+EZXAtA
hg8Kpux0hStnu5lM3t+FKHqbxE2oupZwHJsrz5bBE8MBKj6Uz7VfIHfAZY22vWCdW9GiRzMUBpzT
6jceEXS8Xsd7pOUeOEbZ2A0hLkNvuxZ+lEfLnDtveeDFPXqNIcdeWuPqjQ5usb5RwNHxBT6lOIJC
1ISsd98hXQ5ezvkarUIlO9Ou1twUoPGWQWkK7vXHyAuhhm1MwPFplUCkN7MxQfMkyhUrqWPkqolY
BtqKqIaTWIxeqoFXwM+9WUfhiSBjTgb53JcuGX7x7LRfafHWJ+N9PXbyE31tqiMjgfgUkO+73n4G
eTHhWo4TVreANqGez2k6h+mMf2TUKj2gj/OetFZPCtlN2gVd9PBYuPuiFq3E6uxoYrtSRHvAsz2X
KqHWd3cOPIFO3HFy1L4EW09j7IzcdA02yY/7opU4UYoXXxb+0SP3QNJQndwLgqkJ0g2GPL3TqK/4
p7nLu8/9o/9a9skhP3ot+fSQG+ka6fGaS4kzszO3J8pdIw0stQUohEb+ognx0Ql1esPnIDIZ/7mz
iopNjaxI0d5khdAf5gydUOuOmx6hrEra88o4wExoAymgA12bsu7glP3hjbyr3UWW3o/KVuW4IbAC
jvHFoZcJg+O7DYoO0G9K8bekCnAGLNPPtxGVyi7jAJ2R3KqGXkhDYG32vlq0sEtp6p06PbAXVm13
C8ryif4MgWIHR6jbiE6k28QhL84PIFeKZaqIi+lu8e+3gYcap/G28FEVdQBllKvGMmC3ppdZEWbD
42PYz8TSW2ycexObT+upitzdrrx8gZdomx8tKMI5dnMDpqo5PhZ/WxtcA8jvbNOFcH1WeUUjZdqR
6jkSFDH2dPJIM87PndN72LcxnSTqciEEaUqrFZKnANE8NVlalhLt8BqE/mBOyHpAMDdwDpK5dqKD
p0xY38X5SCab2eD6a/jLGW/Q78mmZ9Ud4I7inlG0OLqCqfEYgLVdz99I/lBJkCYKhN9JF/4lA2zA
J8LDmj+bBIjXT6nlck+O7hECQ+Im28OMAU/VuXY1nE5chq6E/bIBaHxcKMVLa4ih0XMYkymWKCkp
KH3W8jaNVcS3yf+UKJCpYJ8r7WL4Ab+AUDPc2bF3Z5RF7Xw77qCpxR0eE67gYJLJmgXRyL9xhnuA
zctkaLopWGCnc8hGc+b8Lr9R2kK0dOjpx3YRnqjtSfAWUEVWudmTj1WnQTiCaCE0Og5vyp4JgvC7
4rGBqJLGIUp2rAU+ua3HCki8IOX42lnX9aXT3MJOS18812xPLGcjdXwBBTCpn8AJg0WRFMy3U5nN
hofmqscopk2sL8Uk8jdpsRBDIAhwf6vK9eY0+s5bAfJvcK7Gk+HwHT0MftUqImfrAXXG1NZ37T4h
K4OkfwMycNW0H31fEePjRSnUft3DdcdT2bCMUshSxL0ajSyURSQLeGaWvmmZMsmsH+fWsZOpBZ7V
Ot4JfO+e6Er608ScZSfrPGM/fz8MUuz0J2PpNgcSkLv+McdsYjfFq7109830lxncj3yt1PAaXm9h
sOcDp92BVhcVWWkoQpOmHCxiGpnEp2ygRXJCjsaLSbUItWvxlXzagKGwrjQ2ZUt5sjjxg8BPXjYT
OBSAI0DaEndbEl9jT68KWeTNnPm/rdGCt5x/8nY9PfqrBn/4gG7LRh+Cpz5ldEta58euCfSsxH7c
NazP0tlKPOdrAEMNe5cISGm9IJXqvW65fYvd3K0kN7tKR0m+SX7cOugcPFasNz+i/Hgh7WSho1dj
v9A4WKCIYh1BLv4KWsxKO4UPfqaMZxdZc0Vvn5ZbM5av2HBKOWSTj0S3HTpMmnfi4UGHztdkliVN
IQ0mjEcanQd/yhl4W+E7XY1Xxx9Wr9cJUOY1CKkFQzcwbQh65KNSybo3fIwOcdpL2bMb8LtIzsiG
JU0d/EIzEENCmv5SV2R2GN9dJUecsOAwLKmlwBM76GvAwFMRsxKpChHzXBOrF/qUcExAmddoaCtT
YS2CqSdQQCSBjm4BmHWaIX42fm+BTgvOrZdU+qE15QE6Bht9U3KjHZkOrJhg1XKsVLRYRQ9K5FhA
NZXmCC6d2B5OtbDh7l8y19bX9pZbnCPoXKBDmH0UMMANJueV38jtKj++kn9E0COXUjanXX5r52NK
GISxYG0uyD60n8gXARBzYlF+BLKkTC0Abv9Xwe2oSDAhQrctrm/ebT3T+TbaUjkLqg5mkdHs3hi7
PreRr7HO4JaKGSf+K4z8W4ucEEVPJg/MLBeybUJwYEMInGod0wbOMqq9FERWBDWknPBDodl5LlCu
QcBw4VC2ZdxCuyRjR9WGz95SXZyKWX0kyEk/zuGGgHU4TN3hjoSPmjMRTu7AK2Oh8uOoCiQCztXl
HJU2evm3xHQdRqDRqfDY7HkM9/RrS4APG+mQNeBIY+nz3SA47L4Tys7wC9Ua7MNlT0EZgyDPmnGF
DihLAtTvAnpxe7wY1Y3b7DBGqZsD+G2zb6cZMSq7yePy8B+3BaiCnsrWEDQoM3eVr0D9ymSXERsk
9WR9akqZzEBpiUeATfeKbwJ3uUuzqxlqlwgv/lQl2FanPyJsFzXS9OqL/YMv+/QWO+ooZHs83dRQ
2pkhYokPxNLknZnBJ7aRKzfQfy/UzUTuXoUNYxtSBI+3X3wh9nWP5l5yc9KW83qfF621l7ltkd6K
UoYXnbskjitH25u4O+V0fo/IfxPBQ5XCrFugYkz6fYbRncwHjgX7a8S6Ed/iIOOC4cTcYUOCMcJC
4CiHelDlLgSWuQyFdZYGVBtqTJMjl6VBTifycm+0v1ME00BUlQpI1N/Zq/lpQUQijIpRHN3JG/dg
kCDs8DDpxzTBHGADrFledD5RDsOp7mAzssTZD1O8n0pXr4NMyJSbkw8hVKZ7DMn5muc5V39rQCoJ
1+OqCBt71VErg6U3kU+ghR2K3IsiulRXgiiOCaKxE4oYMKWq+UHSd8dwAc1uLib89JjLcMSK3A6p
2mxXd82OFKVNO/OWkpsVmR2jmwmB7WdvS0QpUY5/Es+rws5F1gH36DFvgdeCQwkgFxmq34kpu/5v
Wh0pjVXyfOfFa7n80a78H7WGddDjhsQ88ZtuLjt0Ur3q8JBe0bLKFDl6mKm08PBFsjNoZBJokcN7
YxrRBHG0wStcEYr0h+W4sUHRu/7uQGK+izQHdD0ffT0sLi6JnRtGmZd9JX4GWA7AztXii7L8X5Ge
BXi1MuzP2/Y6TQyl2S46Krf9FqEy98XYnHEc3nZQvuTioXvC+0j4gFscrLtUUTwnrzSHJAgUqQJZ
6memv9PEyZBpLNDiPagu8fU4smuERkzF469jyCZYESNgTw9nSuGNze9NNh+MIDr0c9o42ti0V1R7
BSpN9y6TdUX0biDdxNc4qL6H/q06ye+tq7zCPWHo1s9o8vBzi30kjfiadGcLxfS9CS78KSOyaxwW
ydSljM7ywp0ADBM/7Cr2UX7sniZ4HIF6iugiKa0DyY/16DyFtEuZveQ+GoINlBlpa4dgD/f+wHML
i5qaW23dmbkiYlhtY4xeQP7WQtdFisHmSto4NHt8baiFblu3CFH8tSzTInetA4FgvUfLpLS3RoMN
HIy2U2zWsyhiHjDKwDoDopNriIDsenGXyHBhX3eUpOa0UcnxNSqC88ql3EyvW8iEjleRCYbchavj
uuanVOHraVwRoRPrVrhXw+pHBFkxVp2pgrhxxShJLySPDIf2ux8wiqpK36IXpffIpxGOCksJIQPN
PTXQwhO5WuwIZFaSmujFJfrOUq+TNUr+wsr+qmZew5mznlHVGTtTr3elIfwZkl3vJSPSt2Zz5gWG
SG6Zdo5UxM5PncHA9ClDnhPBLiF7D+fxIhzPdfWEGHd9jvKUyVUYO0O52ZygSHLZV1qgEdmppV8M
AqEBQQSDqyaZRJ0C1XAeeUPFSDj3dlUZYbn/Q63tYx8+mUGbHipgaSAcAAUJy/34B3lpOby7TUn6
n27TlliC+lT3TI/fQvpZYbKwL1d6u6lR11iWlnY1ahzdLti6Xv/s2BCNjI7DlrOm/XhZ73UzoBfm
F1ueh0SA2ppu/vRHxRhb/MmhmLnfIJCe6CGTR+eT6TBur/JMyFffqPnrujdldw/UdlUU3jUus4N4
0Y/acxLubyd3WFZKB2bjjnexKUM6wypHgJOy/jQLrWjdkkB0YV2CHngshVIBv+jRMTQJxTO4u0UO
lUsFOcf8B8p7+DVBW3QJ4Kc2jMUNi7Vnfiusy8HAhOFtntqtiGcW1tWqUbZQCMrUgCZq5mLyOsgo
csfKj1/N3m+C/79u9dhUB0RsGRLH22E8M/8FMPi2gwM9OwcYHSS/v8YmrDsjW8fvFadqPC0VEg8v
FmucUR3eaL6eJ+uuOqkGyQoybpnd9l4JFfe9M6hXUw/BQdMFNXMf6v1Xo37+ni7OnpV8TDJYoFkI
0i1NmZ8nWBDcTt9aygOCEGVYq1NNewMZD9a86q1ocUEQVhB5xB02uvpjP89zWP1BuXY1L2khPVUr
EWWzuobqMuMEoErVILcm3Z2rElhOZNEGt20/2gIND2of5CNLHzbMJLQTtq6xXg4WZfoZMdSvRIoD
eBGwc/jSWzZyRZSUOi7/v296QQvTGY5eKfwJ9VHXWVKMdxDoSsAsdI+KwJ8gl+PQRJwmeEY7mCQF
a+LVYKO2CW5CRTar64dJ8VXVOHH4K5qzHEheUzLNI+8jqIaDbusMMMaPaEg6bdRy81jQ84L4xCTQ
EewhJW/ZVdJ7wNyil/AffUAXYTIzIUgCWGIevEHI2CltmVtRhxBElQu8VZn/ZhirvP5eGiR/d/0m
oKZd5vYYsPUdA8gkNqGVljgEXjFTD4F8G42aTuwLQ2i5yztJ+assJ5azPfzPcFKy6G+6RFyRlPUM
bAw0z5bW5Xp8Plu9PQPgOCSrn6GkiHqUIkQUWUsc5a4nqdEuKrNgRLIhEPycSfgZQqW06d5Npx1d
GMdY4vKTSyzcN4fjrJSCGZS5B4FzVuAuZTaiRFKs88bbTbeBOhYg+30/Uo9kOScPP15CUpyO7Vrr
J21ulVEc1RtWnGvFqSkjD1QewFfAKM/IbA/SZpmYv8mFx0ut2+mvAg1Np7PKSZLt5OTELKgzSPGL
didtkL3FXqyJasaZhwdBWX2b4lG1IQyyH80u62A/M1f9qIfqAcF5ue/y4LR0/F/WuVzqlMmWY04d
vBJgAT7obAOQ7hFaI6F8hEmF6o5bagOWInZSoM+gCNSfAyPnXqxTRX8ZKDrGagRMHagfhteg1mdU
M5LJplHY5Mne95pE8ckXEi/4G8liaY7GKrA+bDor32poLVZRB7b/iM0ucqxbF09V3qeB4DGKZxPv
MFoKLjhoVmJtiFTMRUzqoDlK4/g3PD9SAOhaueg+ja1UlPht2Z56Qal8XslmzYUoGZEZq79OgcN4
7Aw5NdARVLl1UDCA9W7daqDDkoBvLPBWgt15EgecUIfv/7OxJLZu7aakOau3O78Mxbie02jyTO5m
Xao707mT7hnkhopYaEXUlUZxSHrViAOljF5l0zYc355tbgUXegPTU2TB+BqpOeg4MAHrKO3kZLym
dWz993lB2kg4O5P/l78t/AG6U4Z9xrqt15AcO9x/CHXi/1mFTRy39q2azXAUJrzUTll0772wy/hS
ehZtr2+TcMoYVyy8EUJJljwecgL9ffWYTCL24f7wQJO0IyaQ/9rf+Ac2zDoug3J1kHHYpagJcrzi
BhRxG/ZQSNsnbvS+u94ln/DoCUwZYfMr9RWt0vS4C+jDcYmWa9o3IcQJaKnbUoqwOyJ25guBfurj
xyQQ+vqcwd/XaIB/SFuHX8dmsGxNPoxOYIM6zSfAqaoS4XVf4d50liAa4MVx4tPByNCj+m1SsSrj
7ynL2xeHUtZwesQBEZGPrwNeyypAqClcGADFA52JDz7Baw8JxJpZIR9QQqmqMc42HppwnYhxaORP
0TRh9eM6aDx3aE3YCAt2hqok9jLTneQcwvVwUgycoCzRe83FWpMJ9M+QIXIA65nLsz8tjnvLKZPG
17j26C6i4+G0Nm9EYyf4sdUJySVX1UZpkxxpXWiNBwhi7azLC2vkK8AAcy6PGtuIp945er7Vk60E
xbRExqoid9D+wUwRXnudHDjOE7R+euRZjTuEejlP0DUZqtzEfeAo08tiF8JU1+huklMh92a/A5c7
PnRgfORJNJron808XRt0SeO3ST+CYNeGMxrEFfM1Rq8ohI6JiQOzcEoznstM/Xo9t13jbP26FQSv
HJqhJcgkN1EeQaPrJSxNkVQYXg047JzN66YCHyThy78GRt9aOOSq/v9N2Jr6OCvM5d91Xzs+U20w
5/KVEfa0nZFgr6vek9D6b1ywCPwH3n6+vzMC8I7IxuG7MprCxjqjTxenR6wQA35uSPJc5Ad6pY/H
yayZ0KLOUPxv709lzvffrQalsYlwb2buO5ympLPAkW042YOLlnnWAAj9Y6AJquMqaIlALXtpoEDt
1rsfr36GGVMPqJa+7AWiwVgzRZmrpKynXvyMAM2BS8x4JtMR//9RdiaXXubsEu7NHhRVxFCUoZa/
KN3NHW9NmQASclQRy+sorv9AX2qp7cwAD9Wwk++hUs5WuVKE5JzBhiLghKJgXSCBYiOkoimO6Zp6
5+DX+lBfY9is6d/E7Ofiw2ZashvQoUJLsjsBe5u0OTL9FJq2C4gYKnZWTT/UUaUj9D2NxPVEhro4
jFOSxhEvbcm4/7+sRdqfHzCa6+QenhFEkSjWDZFdTACpMXviCYU+olwohCYsqhZfg5jWZzYEhUUx
Q56kt2MlHDDEc9WZdtnRb1uHPVMmvzusJKhR097jiUfCiwMX6NP4iIbBmcheXBztFsSI8OSotJHP
73XYl1TEpnW8uJjCHviaxI7ToMySmSWD9KvOJ7EMHGS1BujJp4kFlEkXCJnJovntpkmfapwsG+H1
sNrj3ryKijnFbs3BME+VXzL0LENy+u2I0LGWr5/CFR32BEQNr/aFvgG+1C6cHeGR+P4flmu1N4P+
PH7rZ1Qyl9p1wcGRRAq/tNusHTQzkA4kKE3g+K9H825kykl3ffXSDzFEcepydJ2rgIFALspKxcPF
tWNq9rJuK9ETeurN0zE3crJEXNNLLf5qRph32XCjTzgdezbtgecQvC/q0GaKsheqdAIdRSSaSE1b
ctIw2AGcdqelwyS15l2sbyRq3npMVYFrbd3DclAm/qMqFKTJfD1cFH50x1kfB9Qj3HrF6FBN0ko5
bRhVb7JB4fg0PjAtPXdKmT6s4o/qv43NmlunOT03uOjTDK3ebWZxW4yQHV2oABWJdJpK4+SGNwlz
cQrjrkCgiMjCOH8i9Tsu38O0hjaJq8uk5ntjjbx+4rBWhaxctJItjAa6NsqKzAebM5CIwwIF3YPj
C1HFvblxTdwqm8Fttr88OUfXHa3K/yDu9fmRWCkcUBIpa++UiwhNm74Pa0uYGAsOyWVHhfvOjEEV
w9KvuSZYYefNBQ5X2QS3KrwkLoMtGeO9BIq7UkuLT+RTai1yeB53kqZlPMdcFtI856uArmUxm9RP
YSoMXiDgBLG5TWugWtga6LICrdBeXhO4cDEK4xnw7CNSwNvTuF+XNQGckDUu1gGzrPWw/tXubCwy
hly0sAgf6eMJtn8Nk5nAcTQLKeHtsAe/wJfWV7R1ytI0v9oOK4bzz+1S4p88yehqiHHVRKXMedhR
/9amH3eu50edObosqyNbqE7htZfoVbjm1t+rRnDvl9T1fluaMKejm9cX37v2W1nErCilIOfoQAvG
X582J4bzEVwLeBbVx2fLHXaEK3Lqns3vTC2WwaWT3RW+RzObi5DZg4UIk7BO/d1/WF8WKQGPrpkr
HvHGbXMmOhlOOhGKvhMYsvGHotALIpqsw8p0jQ5Ax5td5TxRQSNP8fF3nZzpHrtKl5zQKTVXJls1
1SMPArw2tC7CBOcUAQjx7dWaL8QGjk9bV3kQ6MJcX0uO+HdPml2iEKViZXPsxDM/7wshEPn/DEbO
dX81Iiaa3iMpJtKyKn3/76DAN8NGSB2n9QX3BiJ+9IPhzYQDR7911fFcnlFuhDJTNRooFeetG7u9
VeDUVobX0EDn2bTs8mHqarZeK6BGapn8tB5YoNfbSaSd5t1fy3ELb+JCArKXzdDJEWQl1sq5XXY6
CTy3V1TEKCLHFc79UqmDCBvSch7CnQ5MLKgpaei/kpoKE2kGY8rbftPfz/R4fnZfPTGa8tv/K+PO
OQllh1V8IGtZ0EsU1QZvKHs99ShQ9Z/aIjm0paU36UXuUpR1sSJuQkm5A+y9W4HLe8btlcjzlV28
G6rKG8GyN34OqpP03rAy169a+MiEyRCBF8ISh7VDxm0W8Bt2JgB3p/v76uWUAwdKaWWbxnhdR6QI
rHlFT86SmkUvE0ztnIs421g6+fiHKV8GMs3IQU4NbTa+hytpfIIG8cHvWWRLNBDn3mMFsNtyyUVR
/8EqqmiBQLpas4dxQGQdoMnUFQ6kBKXxuI2SwbdUCoB2UQeNTlL+/2gRuBHiKWTbZwI/czKhCjeK
FXhk+r3rqRLdnT/H9tlKjXH5+NsjrpHZBSDZgPQCNRzuzSqLztM/4Knz0yKWhS5mUoUgYaqbnJE+
vx5Qn4akOejP4qv/CYpGw1Qo+V9Jm9bDL4OUO8IDLKAodZfr4a7wJ5JrkCQ6yODJg9+LHEHV9jMt
1hXPE31GMqOqhS/lhUyebZPgxKqTpELUcTIEYKIniZTDFcxabqOu/bTLQuOgwEXAkBOAEA8nRYbI
h5lqQ4UIYxTWHH/dCOQUvrn1Vyb5gcysRtfAkJnnW9H2eZ48GCe5xFbaDHFhA1/u80jhdvxLAJvV
ZG5xlCd2NCMUA36i5tdV79HS2W7nsFnRDjUqxHS2XEHPeqEQtG/awPfsdnF2fKGMUpyGTqWl2RSU
178+/1LzLUCLpSTsTS57tIP18UCDYmX+9FMkEMIDhuwESLNJDybzLQDWyyzZcUZeDaVhvudoqdIG
CaKEESXr3zgiyXKQqeiu73r5saD3o2/r4Q8NWrV8FuwakVMdJF9heAGkVGdceLakM6zT723Iu8qR
685HaDodl1PWn/YtKJq/HFqTlwRmGYaipdcJ36Qk98wFWboVaoCVyZ9ev2aKf5+wVqWeWI4HiuWt
vHpN7ytMX57dpmlxKmIZKZBN1llJCH9kfwHNbWEBihoXShG0+mlfd1UDmt2ylyQPzzR4glZrSpzE
XlU7IJnp434IFZABl7v2MwYLtExBE8Z584P0VdJkXCj3QTfFNB++XMeHltt69abgsLBBGtchtpzA
wwS1IbGGUpicKqpFDGOIV70QjLcsW6NK7aE/ytuqPhauKAJRlfHouLkDoN4SHhDkcxsohM0qxpmI
WRz5NR8rjzmmpg3oKPKyxx1YKbMhFMCZC4gfo37E0iN99CatnMb13ipJ83X8lTH+/tcpZ5D6CODh
DSnPHIwPaDMCd3Gn9RDKsKetfyyedN6vBlg031YkcxitkqUsWYPBgUHAgiqM6RkRZF2ktptHB2HB
PQAkiJoFLFuJMuvrnKcgLrqR1LQ3Q0ym8jnWt8R/WXxyo/U7R6k9nla7tEVoIh4Sf6p7FppleBuD
BCcdFhdYKkli0eaWsBSgpHPsDgCIJVmiH6BjeHxcfndE82Imh/tn1fQYYCl7IvSaFYnKICgX23Zp
/NGykdsHlb5o1HeF7DDQxh/t9cXHqbyHgX2GUsTfOvLVj4PLDi0/HMPa2TsG7ZLcwGquT0rK9PtA
4C5MMvZ8ChiKRLBvwhOeXraJI7NYLzHZby9yTF0xX2B/0Ty8/5SwROv5wt7SJ5bhnAVJw1zt5tNL
+Ck4bZeZyVIIdyiw+T5IfZwGpFo/Vf1pF0lymEcUu4zUuGrxl6DoRa8PcL3/5CwdntEjtY5pwYEC
KR4Ll2NN+YLwgVfwPWJ/4GtAX+SNkoGYB9F6fy/sgyG6TtgydQtqMzKOnMR/jNblTz8UVv5Mg63y
E6wy5r651IANIGLZ+7TQydvdcoRHvnjkQ3Je0kbxIHlooZrd0c2ILgoNhYvoEE/qWPcH7CAfaBUI
XOulY6LVAHhXoe0acTVL7tk5yvyDnAHE5HlkCaOn+JloEW0XsMNFbnI19N+1j+4COifMMboiN+2q
iv5DKtac/7Mjm3vFI2IGhBeKp3rlZ6D6pAd+SuTRXOGw9V1WFgWUQSqzG9M96BB4mss2L0ozkh9J
G0/v3zne3r1SzIxTfBFoHpUghRcwj0BVp7EXDcB2pPLwAXExbA2sGZIHBn64hvV3OwBqOvaFwDG1
c951PKtqqHO5Knos63MGOMJGcT0Xx6PiDlKd430W5D8JkqQQB77EFz6HlmgIMl6yNfaQhu6kUcZ2
hBha+sy8KhW7ytO0aQRY3mVgr6wB+DH/F46s9dJoFbI1ELeQkf4twga4vX9grGG6xOgE6Ml1qL3S
4nJXQw+qQ/yAa3rBZsu3dwBQQxByoemDnhtvd5Orxpk2o92E6BfKvylkjXpg8JRFqANZ14TRendt
XgRyz0pCwTJ1+dDYPlpRrUTcG034o3nShXSLNXSuK6kr6Uw31mxxaYyFJVEmZEfhxvJHvhwVeBAL
ixx496LqrXLFbgq+UOR3heYl4hgftOmTbLgSO1GBftJ0fzoe2UZJnqT+O/o9EAKVKtQ+wFZYc4jz
otdL6sOv4A4EG1pYpTLbg07TzVvEP9YEr0F+OZ853gZKSQ/SllYy/8WGLiWfFXmhAXszTfgUTLED
zVXTUTLp7aBMWB00QPIDadju2NJx14jwMVwyK6buVne4I+sH86mAmaSY0fDi8M5Wc5kamX37ofAN
DBDxCi8YYBo6D2Yjgq7ZudNCZjJ5I1zu5gY6lAvT+lwlp2CNd40KlrLBvDTqCYxKCS3OA4VDWixp
nA0CbqKmuQ/RChZREqxLpXJZruYfOovAxodXSv5TtUFlGsviUTyI7qT7A9zc03BkcAgDmLJGt3he
LfkDtcihVFI2OyJJJ/UlpMUDnF3g5y2btuDJc24zMFSmtsMbwiNwrg5GSnIbhfM62R98dMCfjMkv
V+qhqiISSpthrZYRG3COwuaNNqMYjFMUw6BmlfCgsAGHGJsxjMEYusFshcYbW6VVaZK/pBw+SDtx
DUFvom8umwVNOrclSlMprf+FyMUnWQYtsqziMekSupT49JVpx2UQGEnD4u6Pwflsn9wHv5XdypXz
/l2M+GU1Zx57zGVNfDmvWij9Qm9lLM72ochp/MR2BAN0D/MgszTY2Clby7SxU9YJHLYN4Tw4Havp
+DJRbxHDeiJFrUXsXSbFalGherjUPhvL7XznQvKJJ+FvrC+UCZ0ZtzeCI9DxEuP1oYotg39tRlZp
oDPY5Z1kVafGVBu+Z+IIp+QUoPkWqfD3sQ7UGMEY2fNDoqbsjUf6ZfwNxPiJi752Z1eMOsxHc2fO
rxo9KVd6+yfRXsY44itrQUafL7v55CYG6G4BpsUkRLb6OgGPE0ufB+Gl8We+xRp97RgFvp3dmNVy
t8UkY14o57Br2jjMp9+kEZGyK1AVuHLiBjg1JDFlx2CXv+IYslJxAZihTyFZIKkNG95BYGaHxl59
14tGjWKYN23kSjQh7f596puKjjo8afWSdDka74njNT8Pm7Mq6NggYwpYrNgx0Zw/jRqiEUyuYo1N
WKmrrFQ+xojdQlmwbkg711lG3gLbGnx6/kRKaaAeLrK3W2vUoxEFpIn13nkd3HLAfbvX0cvOue4N
eotuOkkFB/Dk3//iolEDy7FIP/Kw5GSl2p9ph9yN1Fo5LOPUSuv2vWzfc8akFYl8BmtIBpgjvhe1
9UNQtnRFWWp8Mbgj8HAegsqiDKvJnuQBTogoaClZZA+tu9XxGsqdQvmdelTBKVxUoZnplbkfWov+
XFnn4Vubiv/n7cVjQ2/74xpsD1gybKPU/lXhzX3NvAFZqNu9XT9fANiMCiq3yx9f2hKjudjUyNSH
WFKu2LUZsKi6/VMEefYpTM4/8u0NHll9B0lHDhgRwoV+Y/Y5rvrUrOYc8IIBaFVvcMyrr4K9pM+b
NhXolvnt4kuigR2LFyA6xGuFjVkI612oQk0eRvQflJGqOAsvSyCfTFKy58C9DLdMWY5gTEqDQA5q
tzLCinVe9x3k503I6uTPcJ91wBx/Ax337xajox5R6rAB9vMT520+q11Wq3rD1oe0UPkUpqXppNN+
uJH7dv+YsmpLLPXoeb1rls5p+qtOCC4IU9GfBRhTxStRkZYS52BrUbrbZYy/0fNFi6WU5J9Muml3
LawUfybaQQBw050903SGGZk/h2IugkzNv5kMcKW39ECdJabQsbMf+99z7wKWjAID0Qfhdb4XrBb2
mBlK3HfKvH1fGRaLyYtnvFH8VQgD5A7puoPn1l2E7OWu6sRHpGnk0gDgNtBxvEizFWQArOQA418M
113rUl/eQVn+O7ZiX0HkyU2gg87/G6URLi1Hkjr9ydKcNMyqLB1GyR9sPeYXC8fzHndqHok+GqZ6
4UdQiEZDK7ZEHuND0WAi4fvhp5G7XymK1uVRRwV8Rco7TVG6j5ozDlbB92UW+FCOWJvDWyUTmaas
ccUKBlOzoTzEaMNOqm1BIIBYDGYCvuOxuyNxY/PqoGoKSLwviiOtr7hYcIkZJjZUl+E+j2ueb+V+
FRYJ4URq6181bZ9oq4mP3MQFj9/Nc01TcEjfl9+fB2ALmsX57FnfHL9ZjjOqja9Kx90yvkXgox3f
KnFp+FdhIH6EOsGvCFmlKxfzhHDzGMkuj+y26RDmwU9Eh7fajCmRsKWQKjt1oIBgXJliwgYNstaH
PBQBPuqLLDSp9R5ImqyEQYgtaz/rBkYjPHzpKNPEuIF3rjUvIN3H1LkBKQGdfpjK8A92qv5dFZK4
hGy/HMsM2s/k3moA+qcmpo8uKciUWhbixMQPbkBBXmS8/OHkkWQYcw81MJ+mv3KhcZn+GfRIuQ8y
XtRq576AhGS4Ise9QzyFV2OcDQSFU31Tw5tusnmUzGzvfmHv1IPEZK4zphM7g9eUDIATuH/Iz5OA
YrniETaY+LgFbYdKvv989X6npN5T9sXIVWRMaH9cZAzx2CHkP5PrGOlo9nOLGjIUTsMrpITKmQ4c
kAac+7pxSSOsOHfzhfajAA2AmN9gEBMIQkVzjHuPLerzwwJ87pIBXMk/QLLWnEpbF47DfrHjPv9I
QexLzMABNgSc16B6IvMgxF7PDdGgh5Er3Vc7nFuwoJ8S5dD/7+mEW/2wSv5VeJsSokzujH3Aryjm
F28ukz2O51vqz3f3JPoknZEoe3WF3H38VF1mXBALE/cA4dMkMHx5QSg2Lej2c0g/j+w/Grcb6IFa
a+PXb43WTTBsyjuzJMT2TQa1ck1KzaZv4CoWKfBHpclr05cP62e6gcIgmTtZgmA6wSsqvF03kljd
ZgbxcnDJb+WlNVM991zD/qT3G+ip9cdoxLmiubCXYtuGgMjKLFH3/7SZ6iV56Fp8KsuhS2YQ6X1B
+0lEOcYZ2oIKkHDniPx6NKiE+duc7PEd7OW9kEB6DqAl34IE3JPFTm8yt5NPs/TE/WVyt9CbzheW
kHYSSp+edbDGRMbOtL/8dNZroLbYW+o/UEmS4aGfZzyIpSiHlzJgBiMAtGJWMkTtUQZvTZbh5IjZ
jhrhpxs49dPYiMS6yR7r6oKNyJLRj4zVfNJm1huKB4iZ3u5RDGlMS49wJYxotKHFJsEMYPvUEHTS
ql+LtgW76NE/u4XHygPk9dPukIw5pchyD6tC0rFTELymdUo8uyNl47bRF4Xm1dq5s8QkDN2a/lLt
ahgjzkU587xFdXnBgPuMhCDn5i8BJhcxf986+/Suzy5OvrpoByoHGPamEr0kC/Or8n0/KGXBvHzs
O5QN1L09/tHr5ToZ88ioNW/H7Hk99eHgJQ92e1tjnddCHt+DMa+ZeOAMR8tfBjMwenLRQILvk87z
GK4sjUV8pldoko3TP8kSDJjb0iginoF89NEuGrNghqY94ifHq4P9cZSCVkpL7eduoi/2E8XDGmx9
EEGUfdQXnTa+1QmIlheMJ9rCrBgx7hnuiihTfPKhZ6p2lDHOcCEal3McCEyRuhSxzzBD4AZj2aXE
HKNbaBzr1ty0vdkFZSOC0MepwxUC1quUZB+RJTfRKbGpXknp4KqAHOYKOa1prRN3XQTJz4hqc5SZ
HESzBEKZaNiT9ZvTrytFjRP+FZwFKE3ttCGpzWgfqy6N0wUsxkoM5bcpf4jdfQwVtRYpDJWiVCjT
tXYw1erWRyf02rr725QuI7UG0OEQ9lT/1qU/U/NAHDMSE0AMmTwCjdKciVDPc7WUvvj54BdWToc/
qWGji3zbdCbnuz0kq5XBU/tkIBBx+2q5AfzHNNLfizQYKa+ICv5Mto6Fa90TnKD6cvE0ZOheggjN
W1z3AUIwwgso1nDjrETiRQWXDLpw0GyZ1coxwp0YLETB1rXQIL5cyopshFCw9EKRsnbCVZYA8/eS
zRuCjARaakvaRHdP4GPhF5EardzVRgM5lGygX3NDIHCttA4foW0Y8kQZQYynlKoKQ04n/E+zYQqW
znmMCroquTr298A03tUwATqrgdqDaDslROSex5dsfJuy0GZtbGJ5XJ+XOrWtFQilhBnaJn0abjah
3p3wHyENr6xS8K6GGCoVpZ3mgfaGA4JBZKw1O5eyk596veir+Dt5U28//1PwqWjsS+anEcspBOr0
oQZj/GRhuqDIxg9wlG42q+PHwSq/kp5xexdqUJkLJnWro+/TY1gkSBhzN9+VumWBtcZrXIoOaOTW
dVPuHiX12om/irymCnU9oNfc7HSGCo3iRQqgR44GhMO30PoJ4kcea0cNj5YwiFpVbkOH8H/wQ1aA
oPR9gCb8lWxWocvU+TbwxBfIHtzPuy46Xn2OOimx+ayG7ImFPloGwPtyss8IkCaS06EXuzFgXj+B
VgeOWVR8c+Asmdp+NdnFpZpAXJF3MS9e6TEo8hymiE5mOLhxBM4OkIBgv0qvgkw2uLkiLmCkua3P
LAlgZqjxWMlK8NFgfmKZW6uhiUkfvi7m38/IHKFCBHV5q7AvTJq1rnxEqdlnazCs5czLsgUaTyXc
X6FVQmfQhb9hJAqD6rtBrGV/8dEBoXI2fvzeHvHjRVwmebHG85Wl/mpnt4B1H4w8Un9zSXp8u5J8
O0mOAfYJ1SNT5j8sJ9phsnkIZ81MHcCptpGztdowmRcyiT4ZHOJkc7ZTHHg+qE6nkwXnpEhC3xS7
9CGkntvz9hDH8VVu3YtJyEyTIbrU+ezuiop4vwqk6TY6Im/JSTfNnxrLRsvmwvivF+ScZutFUTGF
NB0f1FeGzqJ5fMfKqEgYSeRhUDRW+L8qTidHg+NUajux4enx3/+EisW/qAY9NMnzh4vakV3Ln6Th
mbRH7ESpv6k7jGtB0aogvOP91XHSzBC8RRdwYBBq5AkKV6N6VhjYE2sbRwgaUfUEUWs/uY2W6ruz
GuRvGvR5sNKUlU4YrFougnS6F0z7QpaPSD6ZR266yfK5RtQj5zlEwvWPsnA0SSH/MUFDRygB4kzx
XX9s7RqCVad49iLXKugD9IqEJJbRjeT7Nyz/bG9vgdCHLmzYKY3HSIidB6/hc+LptnYbFC62F4Kz
qzIxbRtpujHR4Pu7811wipveMUOXiEDqMwg33J9McRwSxvha7J+VgN4pgJ2veqGzFdJ7Eeih6/sI
41FlFYNZ0tSJV8fB/SVqSICkiPth4ha364Y+OyS4MC0Ak8AldTz1FS3dPKFHQ7WVolP8XVXynSrA
sw3oCC7qvJVd0zKGPk2mKiEVZQj247NVubpJQkO9T/o3xMdUgD9IrOfFuhZmgjylE9flWoEIFCKc
eY/Cdhd/cTKbEecCjHOD7zcC26k/zO3RgdGKJEO4QTdBRcgZPMAsENzlZuAY5MEZxqN9h2udGQbR
+BawvKOSHHLS8bfcQ9CxxoYWDmyOFJ76IDCU2D5DFFjraS8RaNoYpdYPGmdAYdfRzJ+tCGzD9102
ICSecqGkOE4Q75Ip1gzDSY0FvCawKCyYOz8EhKYmiaVHpoxmTLgWmcKOlUcdgGW2O7HteFmSxM4p
GKhrBpTCPfLtIn+b6J+TIHDPEG1Z+Gr67/Fd2dE1dAOjQ1e4WUjjngJrwUpNZUGQXRFVgHYZ1h/L
y4pZ3GYhNlvmCeFr/Ud4gJjpta+QJ23rm0qCV9Gk06jdaSdxbo2+eKYZ+ex2RO1Repa3vbD4yRyL
uwyK3D3yzLUvDQRUHn8Suja5NfQWSG0CbftV8ozdcs0xMdKliPZzc+UTSf+CX4/6pZa7opPzUkY7
WaJwjNUWNu8xO1Fso3mrBjegg1CNqdq5ap+uJ9R28YdbEC7jRNMtgKFPwh+kiFBxQqE/HmRiT7QE
m4tN1WMC6iW5QJliGNzKHG1lq+69uFpos5Zz1Fmsceo2HjzvJPsryAveyMTdr6InPqGU7PQIh87x
nkICvqb10wc3+pRjTMnApN1bkp6vub0tMGMQLcuhbtrcSBY8LSypqqCFiPBJ6t6WgqJ+mnrVumtR
NER9VLaFSzMMC/w9ssullfMVhPrIuhBUqOvdBK3vAiryFakQQb+iZHtxlnAkImkNaC3WxbkGsM6B
kKmLVGvK00F21vjfMSiLZ71DK89WF1RkSH7aiMSe6ftisBlqH5BgtSXgAQyZBItjXg75vMgd4evm
DbVCAxhWiddr0SQr0O1Q+1zSmF/EXFbm68TG/TKbxXA1IA5+7iR0TtEAASlTeHiumezUVod2I6Me
6t7h+PoDRqnov7sDqjb6o/yh6MWR0UI802S7M7hBpvHuSR/A4FRJBN+vUGhRx6pNNxqveM5G0dLY
StF19aKp4XL7THkFnb6Zt5efp+KfWok5e6yhQxKL30s1tspOXJnOhDl7KijrZZ7kpbtb3EUHv7ff
7KfkjFyQ/r+n+6mfiRwTHfdwR6AzwrFwTuYu9swhuvZkhwo6/NXfH6bN+Ohf2gNCvcB9jdRpsdtD
nLV8Ab3aDGkNBytpOCEYAkjCcq/5IW2TCApcgDTpkHMwIYkVPT3bRB7FA6MmRNxDCPK1rlPHAAny
6fzjkU/4xrCijRssUONJ5jgzhxp88BlmoA26rxZdO+nCy1TFMGC8Qmy1wRZenNTFqE2hLZNK5fZA
IpkvTlUg++8ADi8PAO9Sw8dZ7p4v3KLbXZ6+Divf7w0Y0FP4XJHhm61sAknlG9tOVITj2p6tdq6s
DlH580hDjSEOupk81n3kcDio6izxoGeYlkyZ7jdpmCvE6/GZg7tw2ErDJlnG3NCe9lz0GgSL49xG
72yLng6Ss6iDi3xRugeRYlmG2nut5SM1HG8i/y3RuOauQix+ugI6DmbRcM9/vaWubG0JNPtVjrfF
gbqA0n91Jm9S0TWF7/kWWDzUVg1c7FsgzMUIV30P66LAetRuaUV9y76C79I2CLbsCqCrD+CYASUn
IGsHfFPbBgeoUYrp4MFBlWMkvJ/28kGkoVgn+aKGyO2bXXUvhvQlmFmIqZ0vpITke3rTMV4Xv++B
bOA6nmqOJ32VS6w8FIAgX5DlV9AyaHREhlvzPpR1JYxSP37uVtBDjPGyP5IIjxNeEcKtipCeTTB8
WLmIJa8PAwtaUdwtTk3ABalBqyvT2ynuP6by/31IUs2iCjYmhWEWFiaZwfbhGpFxFl0R5DMulrh/
nU6PKcdOX6kC7wx6GYxbQjBN1QJFI+PzNst5HBwUdV7JuKF5VaeFs7t7Oye2zbRY5zK86RsJTrmx
ZaItBoh8ir9UAxlAHmhc/7rnXrwxWOLpu8BUSS6oSGLYwCDoELPYrSK9mRtebKf2W2a8e+MQPbeS
zf2YqyzbrvUv7lNpjUdjIwwb51uNVtXyqBbpcKjHsEtlXDsQNw3YpFGL1ZXeegVAerZ0Xq4xG7Ot
RGS7XElYGKxQAibAn0CY7L+qAAbdiX3XktkJjOSTAF/U0nXA39V29EnVcorOwxONpNmrrzPGLzGE
2jqRNQHPZNErMjao7TpA5kPqaGNr2/n+eqmQ4l9p2wtaRP0I+ofKX4Sam2Fux7ZWwh8YQ4n0jFke
iwztsyl+AEFGNu9mdqMOT+FPNDAsfhKDwwIIG4a9q11fz0hMRQU8yaScZqKy0OYBOuUW8xwc9hhI
+k+T0R5BAswxYIHWIwl8oIsqOxYdr+wECZNsw5+CiAS8QTa1dOHd9NRVRuXyvGT0sLoOUgucQipa
Nt1PeCGjLZB+fCiudFStl3zFkY4XHklIEBChUL1mbe7Ei/GZDWE63GBdwy9mIdnoQftvPPn7TDJ5
fJOkEV5Vn9LT8kBo85YPf6mZcEmCzXVyPhAzZMlCg2FXYAgKHI9vtf+IunzSfk121sTaQFqIgFY0
k/Absm3SqXencHVt2leM9N/bILHSG6qmcNuMz3LdGRKC5abcFyRgHMjnmngeSNlxJK0UNhhxB1zG
3y8sC/t4rhx4Ei3oqnGx5vpZEsvJgmQV9ZcmQmP6u7tAJxtdMtjo9ZyzWDuYMiaB0yhw0l5mwGQk
HjGKsy7hjDZg9Dvm2iVpiuqYBc2AphZy9IoDn09pI6rBtGL5KrfdM2lZ5RGSOkrj9/5kWrfTHERt
2/KnazCSDsnnEUKsxYIhRmyItuSTAac9svEvRk6/25BbFl0M0kWWPEBJFV76xLQoy6R02CK2MwV3
01k7580s3+zlzzF7DnVxvPbOLXiHFAXwT6dQu3cJHE1LPPLImNWqmQ9PPrKwunXUl8vtcTAuzntX
kEqmcGhdqtNSVFRwCh3zJVj90X1G7pkDMqv+QAcl1gSH5KoL+YC6msNIJlJJBVi6/4+NrObs7LU0
UntwrzQQjp0BLKgi/+7xKwKQWoNPRZXRrKdAWulIP81GuiOiV2Sw7TobV0ICr8YTRPYZKtn5/ODf
iIihuDAg2glMtQRKX8DwUa+l4iQmEAEZY3bbRtuo28Mr0lT2zIow2p2YTDOuTyX1y+C9V5b+oVZF
O92GEEAscj13R4153LTg3YjhoJBlUCBZBbaZNmwpULb5j+ht21EJpqbf39k7dm9bYUR7BZbKREd/
q1SurY7sWyaY8LVoEFJ3k2D4EyIPxd7wQ2uGxfBjYFJJNvmF+HPBoN8hnNB/3ePf/WamVrkeKhm5
9mmg5GpmgQ+tvfjMqoHsuZdyVeN4Z+QVRY6w1U8ItTGsyYuED9+u5kZIhOegBRxnJlHe4qgvs4d5
w8w+NvqD8UVlQWJyaOpsFeeYyWZD4+U9s7mYi8Uz7Nb6tpFabGCRL9dHydKUTAey66AAVzthdfpL
s/JVoSdWO2PnMrnj6R5Sh4XlghsNh1swdF49UPq4+I90WgfUhFDFbr9hHXtKEtKXr8tbAHuFZbSo
bfuJAwMD5uXTxC94Bxdc1FV9jNm9Z8RrL1HZvmV/xpVNwljQZ11zaQsrx7zNoaNM5spts3fmkuJL
eZHqqLnb+sYhXhlAHu7ddjAK2gv/sxtZvDtrOw/PWIiPA9CiwwLwGAtYXzRVdRjQOiq62vI7r1lT
96cRTivS84NWwbweircMHn8q3cQdf2QT/yLBrpKP1Qvrz89mpDvpTxgoM+w26mcrba2T7T0bgIqO
KmXyz5E/fDTYxH71S3H7oWPdHXIBS2uQB6Q6erd3sM3ZaSopqZB0JctFHEFGH8jAXVOkPJ0gZwLC
0p0RYGgoaXjXP6liAnGEqHErVC4SBa5KeW9sqgB96H8vghf3be79a4zmOpwx1DcntkEKSbLQXLEt
05wLvh1z7eFjSZarCgMALKSY/3Hrom0wMrFvYwBHEttMfy/k2woLNeX13RnDVt+GmbMSCxqIfO4J
+6RhZqI77XXLaTopeK3FEH0vI0/OEUXrpdTgZGWjT1sKYkmczutN6aP6jPj7kSJjjJ4PFcQcNmAu
dPa9Pw1RiG6m3vmnDieh49hiPMosSjW6cHY+RxoWmuoIa5zYtZEgEyRDGcYZHmGO7vgvhqSJtv6w
VxsZnAlADrDoZZPKoWUaA8xhIr3R5YaE2EQNiFBZhyKEFpLQVEO2mlggYst2Zprnay/C8g8OlyRw
K+cuQ1M48uHUb2doFZWGjGeiy2NScoq7ub2SRLgtGJTf1dV5whl4fVfafrXHtuuVATQDRwgew1hK
u/MetWzDShcwbO+Lq3opn7fFppnplLEHKeidzogWkomQlvLBMYzkzl2MK9c1XFrwQXS1RdQ4RQBQ
crsWsqTB7eN7RbPCzGl8zy+OGcLc/Edq5k638B39I3cHdXPKL44OFa4/h9Py++USKDhJG3l4SM5V
9KSYJ0wuXL/1DHfRCJJStJGovNdIa2eVxUPSUATVPW5T2j9Aib12UVzgsvzOZZeOG7zJeLVSW2E/
3MOPAOyhzh5CykR/BUx9xW4p6p/yLiIyrp/nz8+U9R5eyCDVm6dzDTkicsOeWbhn5W9YRo0Q3Bqv
2H3h9P5MlJnhUZZCO347jUKfwuvAsbfYBFpmSIOzEBYb0uou0iSNK6N+5kv6mAnTYaOso0ES9Hbh
MJXtM/Ds0SOr6405gajbjw8VbJhi+3p8fPtJLYZZJvEp5B2mdN8rJre3u68tnYjiajG36+hqZVVi
5NGJ4ljsylXWsEHzPM4qOKWXMjZNopqIwR60U5S5rrQ7YhcF8j0yD2QS9f8iWHIz+sNd7ZiOtW0a
NZyEYSJVwEYi+YMH7/+hDkJA8c25lkId0tNdciRvuBS9j2/nBYcHoclrW8DEAn2WvazH6KjFl7Vt
R/9qgtiI+sJHtboYkFthxoqZZ9QeTuO3/hE6EmyF+Z/mlwNZHGoQ8S/rXJmr3pLhijKMeiTo1TDe
1P6t427A52w2M2Rd7eAkxnRl16smngmbZrNj6S0zE87Hf66qEZSJbit3c8vBjUG/SGBYr1mWpVyg
Sxs/tp6tzBDawiSBLuXagp3oz6Iup69nkbuUMeOBnc+8bf5FpLFSNlvX20aaZPDnblCZpXxc/9gv
iYAR8E7odL49Q/LMZLxvS0SFPh272zwYI+ndHkfG0XQsAUUYm7XtLI0z8rClegfjGD3swS71XeDg
yk748Xhr6JBMiXQiuPvmH7GBP7IJvjXAWxmqv7S+TgRF2TBW5ZPqz3j5aVyXdzr6GtenrQGQs6ez
pTZzPsuMFgQLKDlhen8OLpc7XGPv3Ap8Dg0yruXC2COKBlJ1CsvoF9IZyOhtG5IIG784EbKmJ/Uk
cQ8R9oiTGw1HTw4A0q4bYytZFuJBXAf7IW5mJ7EYzrVXbWg6ZV1oamXdr6XdFAprdOfePi3sFWS5
j6gpUGB2YANMDCJgTO37wDD7RDMXuS3TYs31zSGFItH4Zli9rIYQU4UfaDA9wMbOz0fDLDwtA41B
kUHUMaXv2JpSbIZu+d2ARfVoqzo+ZXgWwahiT3vvK35PbmrYtxhni4LQsQD7dDr1LPSjEc5JPHny
eEzHHV44XGTQ/gxGUykhvEqJDvOtbUrMmK3oE082FHSkGJd8Yg366MMoix023v8iGQgLREd9mzUH
xikWNxwiOtWh1/RtvZpe4+MjL2rsxJPlmqjQme+pvK1Mqu4Pm/MQ5EhvRWwIuzLsic84vn3lbx2k
5GMaVLcj7799UeE/ExLh77GZ0emTTmAyXTfK0RtBAUwpnoibTUjivIC7ACGfVqMyb+sHC2cOowwr
BpB7tLmbxK3sSi9kSz2uIOjM9pxtl3bvwc6XFza4Q/0uUtWkhmwnfIJfNgy5+zONWpryxif1k2/Z
fo0SXzcUTV2O/6nJs0kXSlKFg0p3WlBhGPCO5cbkWbQwoJFqzS4/4SWm6M7n+RnEuUP9E3u+gvNV
BASYKkBfnHc8HtTNGJTZKMmlU28lFRI1oESTczIUsG2Kjf7u0woaBhgPNfk735bqqrOouy3dveuB
5bxE25wblGR9t/2CN1sRxQzfagQcZQhm8imsjBWWkfeF1o+8P5hF5dFETBO1rXt9CZpIy26G2pkt
3KYLbIrzlGMhpbWqyXznl+PjUzf+IKBB2JmC5R75Jb0rHWA+cttUOrA8JhRiz0a6y42UQoYtravF
d0XXK81aNoqT2t8JeWAxLidkp/ADHxqY8cOFqIDj9Bj2wYE959NB6fzuOF+rg/9ha44Z3rk4tYof
QTIshJaT0RifLzmcdOaPjSi3YEu5GA0Druyd1uOLprIulsf00MPIEsETtgM7uE7N7ah/Tp5qrpZC
CGcwxET6cCEdkN7uW4E1UB03P1kXpWRTuMLU2wHT55McfhRC0OmXyqd/2b+gyzxT7KUVHSp4eViB
Y3hwE8NS7D+ojbY1W9GsNdEB/dVV4LhW5CMJAsViCZYjoaqAPqEofZB9Lh9KYbjXQOFmPZaqzKyB
t0mRYRDCEfwpTC+OkFD7fgUACODz9MNAUImGBgBrBEvy3hNDeJo2tKt1XGeIYuQNwI3kd2EdzzYD
+B37k/HCATLNk4MzgYnQy7h5dcAfIwKHsQzG4/uLfY2JLBofslPFun9idJ+yGxzic5+rSyx7zZNn
k9R0MahyYVBX5EMD5cA5W3N54POqpKWXgYPADV1UDwVapLgt/2CJNURHx9oNNqjdAasTlMscKrPv
AJOLJejyilQ2CUnQ31sLn13CKFh8BEGkXQcRvLd4+fmWlqPFH6a3YFh227EhFEDDFFml9+EFAQN3
ILAZVLXxzT85INmjykiZiF6cjSjdU70UOo902VmOrxL9nyGmebU9+yBXmavEYADTFZrTCA2EhsX3
WVFC9aLH3JhhZj7eduHD1SVhaZyhRfMXsG354SOvOCjE0vSv0r0lwT576wkNTLOoXUmQqsIJw82y
wt5zjeKGAvyStf46Oo9gZc+vFqkF+QH3eKKSoGCSMry5MM6c5lsC4AtMJplyhsjIi2ITRVn069wb
85n3sLNCAM3F+ye7AwvD7D8f28uuu4E33Zs+USH0J1BFh+gpkITuy3iPxOA/sej3T6gPbkt/xfD+
k4ctDhoH4ppvRonBeLjHvB8ZIgspGBYX+Ux1PynDaXX8UXj/+L2haTBHa42wynET2yw4B6F8OMkj
veBjK5AcxxNQrJGICQJIB8BPNbR4UPGgEkGST3DkQ5aUhucV1D47T/pdJ2SrTwF4XFywRLo+yvMm
ZXWn7n/PyfAR+vHRZPuK+dKHWoNWZ3vI3z8cws4IBVmngeND9d6jHxkJTiS5Y0HKXi+/W9eYa6sn
YTSZZFclZ+FQsQ1LiSE42F8m0HrsLJTUKZwAo4R2gCFwO5XUs42FL9WhZDLOp2z9LWbotS/UPX3D
NKisxBppAa1RGcAnnDm0oRqnqm81gaoWHbvoPg4CRQPbpykeVtHNBCMllThvM3YsL8gbWtTe38ZP
yZsvpUTL4kSeMTAYRWB0tD2PUksZIS1qT9CaW1xDs9C+YwXAPYMdGlpkkH5E9/1YKvN8W9zamvRj
HBbRnCxhHzs8ULjv1qyczGOjpIewaFfdrLJTQ97I33RMNiO+ETDlLeSF0ZHByoPiseirvQbzBqOU
aBuB1Ixr+J+J6EwGaLHBqN/q7Uc5mAmO8c2poFWT4HcivoYmHYGiZMnockptFhIOlURpWjLB4puZ
DGuEZC89Z4qKotMxP61it0WqIcqXqimBsjp2qzy/VwfV3OTRowVjn/9l2q21qAgj5hTaNF13fukK
4qm1rfOtKIKCwxLdOBZTUWKZfxv6LHMB+0RB0YE1M5GhupcISk8jGTW/tCri+pdUm6iltKGd5Di2
Qkkry6EroIRWEit+Ye4wfnNVduRUV8xGCK7DVpogjHlUNomw3i1FiEp/krQoX/6nEqB00UFukPmr
JDx2RbliWuXieVVh6ZEbRRksrzyDDJQuMhR6xVk+3JmWNlM0TX7yoTz+i9jyy51Vx/jEuSs4sDPA
Ky8/zeEz+M3+p2vsPy0Fr7e0WsngN6LOXkkZOX9Hn2zQHjQErxoQZOxXmoSGgo/oc136QXrdklnl
YkP5WFYEI8LaHNNiQh3mKjGsNn2z9MfKcGD98nWPufGDfCAxzg44G7vj4vw1/9RJAWpZqXQNKNJ7
9S4XM3FyxYaCMlKeAslw+2qLAWCT/YgunPMJRMG0Sx7XNs1EAK605ULxmu3qIvMhRSBR8hmXrY8F
fM6avrzMH76SolHAIHOOQvLG5YqP2aga9eQsfrtrlOKN7qppyq3wANAkm29fOP1JCNiT1UrP8Gu1
B1aKsmGn/oEZqoa09cjXYAN25s9OCHDvbfQMMbnC55itiV2Tf+nnECqjRI/cTGzbPmOR6PAMCUux
fkXiCdA2Lgh8nqKJvcYDvKBm3dqJ3I4t8QM4XD74pwp5lLtB+SeP7ZVJIMXjR44cuWvaeqSaCM2g
up51fa9Kir4tY+GTXiiaabCbz4pYBA/4KOMhcO9pwU7SungjbSdD0ztqD0ORS6JbXdB58IrpS6QN
nAqDU+MNH1qDaSVKWgG1aGvzJCjQXHnZvw4EziKhby/qVLtCOz2HKbI7QNAfETSy00JmxSaKfr/L
k2VxZFyMLGd9NpPnMIgL4MXhe86Y1X/jZ2Q8HvYRwxvTLVttFnK8u0lbv1xyKGnQYrrzrArpBZhC
5Skzww3EMECRf/Obq6NUfld0Qbc8iNGqxAXvdu5uDuwJ4En/PyxA/aL5gU2WerOIRFlpSSkngWzv
stlHpPB+EovIHu4EFQedDWInCywy1EswZrADPC5/augoSACiNrj2EXR0EwdnUF9cqH4dADeA1mDY
9wyzq6i7KBBpervc+pZY3iwAd+OgM36poVUUrfo48ramhUTI4zNlB9c7INMszFvGFRx/qSvwbcYS
lGz5SYQYj99kr5xAfi77DpIjhUnA8OlAZSygl3d+8PKwpFnCuhTnT1LdlreW9rpG9bICV0MS2ndx
VKsi700R67Vilin5ySTZ0aRFH9UMgy/g76I620VDJcaq8FgqJFhDitEUouOSrN+05qh8QlrVUqgy
jc61IgOCwvI5k6mcVtWH8OA5LbN7KDpxA2koQ3KUgkgpXtKFBbuHTKKeXE08xPQtBHrBstEKVsWO
6Rai67uHmsJYqNRtUndDvGyeNc9b/c1NWGkh17f/ZKopbXBgyAnsSEWzg/HrkFlqsNHPyhVFPdCQ
tmTPmaFFZbSpgnCqbay9Ak/U5CCEIGBK7Yi0trHeXOT5nW9FmAhIIPUAO6P1OsO1Xrz0tz7jewv7
FsmntiMd8WUPhgslV6TQ7QRBQMNg0RTIltx6Ewlion3EoZVzCP0NfIsKPWWHDijkLf6dTaWp9fky
oAKW0sXEcuFyibu9Uq85ooEIlDSRxA4Z9ryGuIzrbq5K2+YAGNwstb8XbBdo7UjZKBbZ8pLUpwA/
/jEAY4m7rbYCkIj+7+0IId8H7nre5xB7lIAAXNyDlkmChpNpitNzq+AgpaT7G0P3BdggSBFiiGnT
PfAFEAVsPXGN7wdK5UqE7y0KYjKKmD8SmvuZbxoRm5EuS2FvHkFM1/fMjyvvPsl8aSufFDU5x7AG
TwXxMQxCPhmJOAQkY4IS1hF+M4KEyVS48CKQCNINQZbxdCLA4+V5OrgHKEPqjVwFMUYMcXZWGnMF
Otbl2eKVSCPRO9UvymUIeSodhbbgCZWzyR/QjbPEQJmLYq6eRH7ENZqauKJC7fg1gyQ3/BsllIAU
q1GIbx9rnyDevqi7XlWHYmdmA3sQzustCQbJdcwb+RWzs22DfCgdzrVLcpCKuz6XqBVntxnAiqz4
+ExGqPUWrqAGfpElndNFOckXvjaFnhd1hpqK5eir8lEUHHSfbt0G82lyxUykuofblU9zbGWJGRXN
dKXf7WdZ364OEZaa/JW5w8ZXMVnM/6FAknuPDWqWGru9vAvEh5LFzBvu4gxVlx4x5jVuskjYwo/C
vR7pWfexct1H7PK1WXMXryNEI8LoI8uvQh5QxR38wkBY3cMW2L/eFKxWVprj8mS0Wlgv+u3P3z+1
Lnz6RHrSvEmRoLCYuHUFIGpIjVttCdzC9G3T6BQvyA88QWIQL68KldLmbZtbbH3MJLQk3hJqCHMJ
3dAe/1et3ITHLsxamNi3zBAXwufUiLabvPVXIQaRrAeSMOBFBO0WfKOVpT7m305Ce/4mqF5cGfsl
fn5vkDA79G0LnRJRigxyJVXEoBe8LKqKgZHF4T0lDUmwnGNNrPVyhSnJm2yAHMIRnHQ2XxPNojvt
2Q8H9vXoZn2jHpydpmRVCUdY/sgoVs1buZ9ArNCkAh6IBUr82hlfxn4UsyxDBI4SXGG69WorQlfJ
t/RHWaZ1Jxr9QHOEIqa6awUwyf2Z/XqAOo5IGu14Xz+RkuVD6EKf0HBm2kK2LSmwJH/DD23xGFTb
0vuG4i9I4tCSYrH90Gn51Cv9sVGMcljHaX5Z4mhbcM8i+B7bp6ex5ufZcQipUJJXGlmD/fDdwh5V
MiOJbyOEujocInkZ/uZfCt9n0FsmLDGW+YiAbc/AZygJ3Q6bbOc0eyrhLSUNO/lOwxMzMGFxL2WU
+e8DQQjbOS7iI98UNuxDSMSk63NAuQvvzdxG9iYVLY2t0lw7eG1ONjV0yzI4YPbIMx2HYoLBKn90
MzUbj4KzwpnxBz/+g5efO72iHxtj4vm+mFHtQZevVIFUgALw8Ma//58v8Zn7Oyi9Cv3dav4/utqR
qCiY6uLttHEg7HZoUmEZ6PJjIF0LlF7tis0K3Al9Gz3joZs6bkkax3R1VCKundZas3gV8x1l601M
PY14MGvHMPzdgjWO8MTNhGPKAhaJP3pw3PdkUAbZKHyIRkzewTiihBy8Bi02vybLrPveAIxQXx10
7MDLd/9UXMBTAHYFAFXfzrX8KJMTmEp6Qxr7oHxs9oIcLfq0NM+TMCF0BS6dJVwL0YmoqurAJfWW
wHFojG9jbX4s9nTc7qN3agdvi48iEOmA4pSo+fGivfrc09u+JgdSuurCuYlWHeySEOYucYsXYxNs
EVY1eN4I+KNMbnH5yjSe+HrzSByr/5lgSr0073f4dPePcX8XzV0If5ky1r6szmUBbEs+AiQjr2wx
yTuSvmMf8/DQEAdZaFqHwtZZZbTf0L/hFOhcd5iZB0wsq8nQn/GPQpQQtURVLHSTzdPPqISOpvFy
PfsFQ0pObwZXLQAL0EMBkXhQO6uWTdY9P4U0n/LVwpSwf99bML7yigmxmkYOjjcJVrWjv0CwRJbm
TFRhbNCY/W623QZrn5RX8RS0qpmvyK8tiOyjqO2baNtAR0nHtmkDzvY/4a7jv08TNOFY2zIFp0Bu
KZgKGZ0NGX0N/5b/8qxLePtKZ9zptakBAZo744Y+7WngSTWQE3RqAlyToztPW58wP0XdRyfLpz8x
jrkHM3MKjjjzF8FzCJE/Oxo468eCu9E0RQgjPYWAs5fDUYP3r9wl5hWOs8OL2HFupBmWyOz7Ua69
DEAFB8v1acXZNUvwlmPmR61ktrcO0GAaMvuSOnrqt/wKXm/8moSL8y7k7pywysdoJP0fC9PYgN3O
jvB0NAZmlNjA9lg4aui7KE7cLaI0rJS/gKnu25AJdFsVWv11IErCU73s+dRzu/KHTZbotfH6CHWL
Ob2SLAcBWbYGxMj38gpReHWSGZl+mMKcJmjEJZ2hYvebP2N1ixh2R0+WavUy79NyHOLc88I3D/xO
fPfBdt2JXQ6MCbbOtJdQK1mGzJtIIMEyO5qErQFqOKtOLJCxHKBnLAymvup2rXE/YJaDhuDk9pKC
2c+kyhAgUw8sjT9ubmAQogL0GYQYsRRf5rVFSVNFLQkXfGNLIBXDUg3afgO5TZL/LFkq7RVrm3D/
wu6pQC0WpsdJVyOcGwZk7e+kIfBgfabkCHyhonLz0GteO7Uni3KmIsO35E3nGzDCEzigyU2p7FsX
1JdTFcTAdvXWvRxMo9v6U9/LbabnX9jknp9UJZLTY2P9TVEN7OcLU5b9oew1T1E3x0u6Jfn7+DIZ
yf1beP1W14Y2EK804vxZwS6zV8JcI9xJnpKdQnsl0BLJJA1sQJK/JHTG9bJjKvanc5Vy4wcQkxp8
Ez1RpsdZoQ80thQQ23KD1w6VhmTXrOE9fyA9ncbCC8CXatIPgIHCPij5WoAceAQddFdQwUdL6lVE
dqRxLj08iKwdfDvvRxrUaoQGhUejcCZOg7YPTican4wb8MhogMEUfN/18EEiwtntclFEzW/Cy+Dn
LAO8pUtwj0Vyl2mrZI7siP+3V1mPdXT6rSOrPa0LLq4m4NHBGjUpjjJcfIkOse8aUfonIuH0ng9b
EFJYHR+aXRb6BeeKL6hP8aN2/PsR+9vuxvrggH4HFzMwUijubx/IkmBKMbNWWSCu0rMOmUTt5Frx
MKEai6pEtVFlGyuSrlAYfASfdNTPbgYvbj6LDLLJGPsoPjk37bopIRK1DUQmsE59jaW150IpqOq5
4eO6PcxP69x+FH5ZxfjptZn2ZUQNrEMuHgRG8C+ww4l/R6S+YZRHTSR8R2sSx2OzypjfXNG2qX5a
9oag4zUgJ33OOmBaUElsY+gChsZHWargBPMmzCn14DPh0GvHuX9VJalmOuoFAuZVXZYS/ek1YSDP
y6AH5VVEB36AfqhiDiYoeIFJlWilUvTkmCHbILGsBFv5/JHhOtMzudtLHVEI0GLA8fgsTifIvScz
tfYZunHjHOWl71ND+gDDfjsVMN9Wmo8KA8dGYZ38vuFL/pxR+cM+OD4DrwVmIdd41mZb2fd9TItN
qIKuHJJ0K35AzNgs+PDTI0W6U52Mk/1E3ginR4St7qyjpMHG+LWMgZVEU/aHvbiXmHwP+d9KxuF9
A1d6Xn6HvRiWvXN1PEdetzmN3jxp89B4ESn+aXxDvsjLRYeKM9kgEtO3k5RKq6IJKjuej60IZzwa
DZvH1sAK+sVC1tKstFHevWYvSXWdX90ovPQsMw3Dnj2aofVv07OEh0k2TbifNtj/yn2RzdfMMI2Z
HCdfhQsYnld2GDtgdbDZQtzBYSMI/RWnYnn9q62IoAN91jKa4rGozJPy/UFdFYdyInrzn6SmOyJU
dxJuo8JJxHbiUETM1WVs1tX1BNdJ8vkhjBx4Ab54ERdGwYJbojSpso7LpxIR+C9xbFFjs9fEZ5f7
fIrQepTL7va7/pYrUQC3JBwKmp+Y97ch96f6tzS9y9M7I2qRU8Ekk3HftVKjgBen++UwoSx8Twnx
TRJ3c1D6GBITgoSLxjl2NV91ELRy4Xz+1CBWsWgvt6mNvwzeYcyeZ7w20/1+CDqwpmrjDYI+uZfy
uOzhqkj9ujdp0IucUH94m0Q0OVkta7xwqC9nNbddbI/Td0OLO+2gXvgC6QKqKrSDiJzvcKK2G18i
f01EkUjQhci6nwt2bAjKMu1V1PISxbJB4IxtX9+Bu+YLUJ0GCouCVZ8kc0qDiLvGJK1DR2Lccmx4
6ytngMIasuWsaszZaYFwLaCWKt0+3rFVstL+SyrGhQ9gk1juSv+P+aREfer2OBEnfzP7uKLOCpJM
HvpTsJiKJmtKA2MZDudZj3J/Ktybuwu1I3AMSNrB6vYfs6MHW89bDNPdSD4pn6NvB81+6q3yUNy6
OiEee4hCj4x8hiaDyNZUZEH8EZTw2Sm39xiSf7Zh/FlI4cGGJWiEeA68JgGAe7S00rsws9dqTGzr
P6xn0KVjiRjmV2/BbxakYk2elDxXJIonGObRYQqxkuThZ+aPYNO8e7NjfrbnYl/QBF7qSq3/OB2q
vRNhDsb9WoPqEhWv3pOCumMGudj/tPQZfK53zkVVwv9jdgwSP0i9eRWZmgKsXH2V10ODNeCSQL4S
yDdpnC1N6bW4xvUCdHxi5oOp+lJPYud66AfTx2QqBSORqkdOuBQYd8cRkwd/UQ5+SMkodzPe77ry
Bn0B/w9CQhsM7dEq2Tusv2bJ6hA2q30jZVLJYuQ/msFktKPp5XVfdrPS51NxtjwtNi4A/s77SLR+
VbAKjBJWmeVOTRxKzxDjQIgReiHTHRXCf4OVriiVRv85PvpOu2kF022mOPXCl65TdYh18DbEL1zG
aqjiu0ma3V1LjPLfzMfrG2ma+DVawY8WEyU9zx5qz10HflADPthyLoENnuPFSdJ7fD+mUUBs5lSm
6o1MnE8nPfUWzygBGuc3ENT0r6RxYhol8KfHMRhOJsRMEzoksX0eYz3hiCs7+Uyt7IFmtcoLQdr4
oSu0j/b6SKbEQ+CUDbJqpJrHRQWMblnaFaF1K25BCH6hi8JrRey0AaMwBMLahdO1SyK6IHikUOWW
VL/Dov3zmOeJdaipawdoD5Vm/sRVBXeAmzTAFvW48lm+ED9o8eRYhesLB6n80Zj+F4TwJVt4app7
s5riBx8oRJh1UNtQAQ+CeLKjwLgKAV/MRrkZzRwu6Y3t53nNjPRalrHpjoeV2gm18i+imvBrcZjq
JIMUrvH7gGgy0XKJ70RMgVT5fq368XteNHkqPeKPH0t5zefirFpW6jz+agQYjlqvLeE1WLhJK8r1
Eq7z+4/PA0GjSdJ63EkAZw+u4WRlkYk3R+5pUy2qVlzmbeJ05D8YWVeqzBZhCyqIhOLBwIzm9XEE
IATxOu7De2EVZnL+CY+XOFDQaa+ZPRVpwtF+2lXrbrb/7GW2+cYCS6SvBDkv3DQqt965BygoRoB0
Df41oy6XDOhHGfWn2mluY8dYuljnDzIDTRW+wMFEpXnC4Yunl4HQwOv6KCH2cliDFc5hcQ0Ib6QC
2fBziO6QT0/Kkt6JvUXPzELZ3sHNlYuSGSquZfuOUlYXdRDk765JdwCmXNIHymKvhIi1WKvjCCVn
kGv37Lbkv17exWzzbC+m0pcwFdq1/9uCEqdhkNWDbZ/vH65XfAYHwROds8yzYeH/EUs4JxM5DB30
BhfwC7tJj2gTklm4DhXJ8an+uXjstNSh5ebzy8HmxfIPl8THwqdVpni/jaBxs/iJy69m64vL0MUw
BG/jk7B/fhkhhTytGX61c/DcyiR2+E5EwBXonGI5eZtEREo0fmeV0oguA2IJQF8c7Qi5GJ7qwGcs
Z13bwNM3iRv8A8jqsboeUdKLpXqQhKsuPySFvhWn6oNUENSUQascKh2I5KnawIOr/YUyO69W4T1f
IkLYwy+S7nknYMEUbWZqeCz/X0JTgRipDes6zQ1vbjkDDAl/bU7grP9VmqWFEzcsleRyiI3U3zbW
Zk+vBOtIxqcLuL9HyeUdmjn+1lmGSHHUOnmePDsd2k7l3gH5W+xcedjYm6h4AQVItwdHDP7RqK3j
uGfdzv4dSJIhXR+wAHVEPbGMVZJwSIHEm6Ids4aUs+dTCETvJv1eS8Hv62Y1A1Qpo82ILxlUZdO3
rCH6QR39G4Y/ohgoy7ht5+92t1QPvGHd85xVdyKUgXf9jpohdfVzqIccz1eadUi3+A7Co9mVqYdY
Km55HXdK+cV/sbNY7i1qaHnoS8QJyM7WAfcyw9u0mej2f9KCEuIDKRgKk/CjqvQPSKPktwSfKoYq
q7iZJLlAKDAR5jv5MgwkfiOS5xX+PWz46eD4WE4x/wtv8TptDAYFjsQ9cab9u6RYBhDvKFEepl+g
6HR9sXGtCsTc5Lkj98sVzeyZFf77ll7dRPlekAKTbb0bv042+WHnUciJ0pw33p+Fk7+fftan+l16
4lVUdRHeaseGvw3oMqoVFUPg+HYCFvcf5e+HNcal8bz6iRMtx4gUzeuiLvlBR3hxRMdZos2k3WTB
39CYmczAx4+Mx2nkj9B4LkGTrhWX0teopiTY/30kTiFdZQNuKoYbOzHGoRFT/wQT+K9dD7zmfCPn
Vpm1Lste/mze+/iGfDQ/rCzYWc7I52VXjHW/kVFGUCuSn1F6LIfKJfTy1gC/TjwssvKEn66npZDZ
8chRkXarTmBKK64bGeSo+WepIfoFcuDgthJJbg9KdFOJA2N3Ea+IYcFswIwEN0Ixx1fVmGsfu127
FGOL1crjiHXHlEkeiWqIDSY4dwk+LjvbjQkqQqSb1AZ5sIJgtcZgpZX0umP6qhmOoLo2ZZejV9BG
M2mwNOPOxwTb8vnt3cLLK79K6oO/WhKGYlAQxmMTYH7SvOaJZICbHooWfnJqX7bs8cbLAmp3wJbZ
NL187sjb53JwWQFZnGl1tPUPGlB2lGd7kkgK8PGUvK6qY2rHXbPXMYLmyOv05ebtttuOK+3rgySj
NLrH+xpzvfB5UsnFFgPT3zhqEcP1NR9S8n2sqNJfxPLzjlkVPjgb2jEU7+aCF0rC/u8+vr6FFXdD
An8cod+KqIKKGFKVc6KoFGfS44z8aLiS1WqReDIP6+5n7B8GLChKps7VGXZN7SQ3ARWE4n93TQKV
Nmh8ZmRNTsrrw40Z80RaM29fajxm692AOKLQFLUgGae92h8lZTkTwOiYrU2LpaEQDLWAupGi+bUq
bmOiZ+I5BAi6+8LWwKkBpXYVi7VVGbnBsowIVGhUyqPge8JvLFaryH91PS4n2zVM0JhIrS+5EDuA
fUhN7gatwibBfmWMSe39YUq7v/HqkCsYtQ7v/jCjJl6/kNcpUSAPSYoPvIgpky55whnUSfnNhD9Z
i4R63Tembf7LkS+ZcUvDDwk96bftXX7jyd4Q8mOBbzCm5vrXxpD7WiFyh5l4bytOtm6ljD4Evaou
AAFfPIUZ8M3bKvPY8APLR4LSfFx4sfzKkK9tPtJFTD0qfWZNTHYzW91Hg6q9IyVXLbuES2qMEDr7
QUiBlVzLahDbPdbZSdzOG6AZREs4nlLm2qzVaML3jgPVZdespnJhirAWuuCR/4a85SpsKWUYez5b
BrQF5RCS4O0GUJC5/7LI5ECq3YfTOdoKJNPwOneY2xhyjquTZG9Ip8Lu5RYosxRUPClDRmApqMJK
1owAs6vIWZNeu0OR2XQ9PyOn3O3KZwjqNvHaSRO3FbVp2LRT5K6wBr6TtXli4bBOgTpMR3fjiqfU
Clb7KoWKy7xD58MjaX2CXFxiXCkIb7SPYDtXvppUSLmqdWDbzRfsIuCUhsu4lu23mSR7ZNE+1XCK
lCR8HTEtzzs/xWwH5Jm0oY9+voR8cBmQkigc/a+0o1knnfSYc8M8Jrmy910OQc11LSLW7EnpzwYn
mlpY4tXg3UT7oA2hmTyci6rWL0M2QccjxQLb0UQFh0CvBy+5T7s84t2f2L+vqm75NM3md+cpC9PI
cCfIsBb+hRbqCwMuRy9o4e4hX8TLM5wH8xUujlCofStkDZgo0qzWJug0QpZa8aWYQ/3xk6Uzd7O5
LpWRbDhKqu7eC+3AyIVj7mUgrsRD7JehsOnuq7QQJMlCWnkroVfDBc+zcF46Ik8FqG8SbIG1P4f3
jj0M94oQ0B61jZWc4byhVIieE61dBfMwLFkcpfL/Ct+NIcR46cxsUTdw2FfvIR47HKGsT2ojcH7h
s+cYeIK/zZJLeGKMdxcKNkNi7fdgDSR1CZLB+987X8PpY5GXc7pSHGSdK1N/5seTcFKUePTvSdqS
fETXFOmiUCWY01+xFXlulcGiEI7wXNECOa0Ec7mTQ5/ie/Gq99OwaKuDsMLv+7s8+QwEBqWSLoUS
0WFYO5Nb/QYx+h3BeWeRRwT8NADjeRTvjRpkzkZUnNFkm6OrY9YPL+N1YOF0wTS05iIYRWsZmDOY
6dtbdGIlfptkqJ4M6IjSUSRFk3WF08xSsDcdbTDk4UycVyj/7AVu15y+N9d4gaEaEprirAh+O9M8
pf9+VfCeOM88LB4lZYH5QrECWBhYCBAgOMxKScyvzPGPkpxl/8YvpSSdrvysFCXsJdRfP5/cYLIZ
uo8VXMKd55qs1Mxh46xWsCuxsPRxeJgCjlPXpyvcXtlWYhqiDKIMXOFWzb0SUU65rXKzH7MRHHlH
SuCW05dPKP7gIOhAvUsFJTd9uStokFuq2HX0qNffKjXNzFSwhs4+8wZGOGyYkfJyvdMJcrLO3HNr
BOiYq290r/c5OGkkMsCI4PUlINIfq5CTbmf5zvRrUCavvKXh0ztOmPQ1hWWOYrq2OjiWq4L/KP2I
Fbv1qPqjNen0tuTDDiZAms9/Kx/gdkp418gV+o+7q7Gx3BteueeEdpJqmjNKaiqqEYTjwbUOmuyq
LEW4RBUuD2gf/bVoynhiNKtb8EZ3k5tp9C3FsY9CNJoFxh2ZRyZ9bx3DMU43dpHxk1tx3f4iczJa
wYX5nQpONcb+3NhU4tWO26ZEchvDnOawprO9TcYYGfPAdi6L7IwnQuloTiMS8TcCir3bYs0qRX53
0HpgnF5MPLMKZgt4kZzl9ErNTHPtDeqBgLOBtteWNJzzdeuJTcF29RkIs8vfn0+uL3Cwjd4g3bmT
pd0wjr8Eko48BgQKPBbMkr+jLp5z9rITp0g1E9d3MOvRFsg2KkYjD3k6y/4piGyEGNflma5RZ4UV
HVNZMN6KWeAMi4fxjDgCC2WOPJScjXzQWbvSVuzTFj7ZR9OGbvluJzMKQsPxsKtM4NeKZ/IymJpk
4F/7rJ+F/bgyLbR46KX4E1FzeCi0LLNJBiZ8KqRx9AswYbwXpr20SotUcjka8f89LE07GJgxBwxh
DzQEeMi/Q7bpcU81lkRPr5ggKtiNWlCsGuEklD2z3/Rt5i+TTGpxU28bjbrek/b4iOMJPpHP12Nx
nKm1/6dsMtHl4zGzP2qzSpo5YnPuBk2DvlXrbI19pQoA4Mhtsqs9Q1Oofk6YOszwHqQrm3cnOzKM
S/Ytu68Aw8b2swnD/fahmWJ5rknLBJOcp4soBxo+BjqSs4pMmjK4gzvyEx4sDAmw6UqUzWF9aoaJ
JPAW7h5SWsomzAk5PtYsu/Mrhdlr3okfl2hGEaTI2+TLxNKPxwMYeaX3IhJAGTiyg9rR5ttfWx4f
JCfSw8qzRmljU3jIWjyY+bDeiDP6Kh2mCxHGJi8/kzTMlWTPa1Dom8cMVyIg8LGTGmHj+xOS/Nk8
gI9t4p9zfTcA+vBxXjZnBbLakdWroejxALEJmUkvN5Necksb4SUvd0mmm9AeLHNdaiAuI8sYcB2W
lyQdbZ+fTHgOuZ2TPyKbQq8if0ZyzmVVYXGV674paNtZABz3J/jSuiaUjM+ZyXDN+IpHKcvvfgQR
Qs7JfkXz+hSj3e0OOvcOq75uoW7RoouR5ZgudrJ+T5vbTE38UWwn+Qt0p78LoUrYKRlrrqyT3y62
KnK/BdVhct7AWDoErpkdvYPOJyXHbM4D5RZdob2oT2ef9/03XQt7sL3yCHy1xz1a+O+jbKZpy2J5
Ak0/pixiCRBwQ3nrhFZGngDPIce64TOZEQ7roC0NqXfjUPTuRdSTH6dczX07bjJXBqZ2uWPglzr4
jLy6MXV7e+tYZmCy7a+z6bDvazhgFVDMahIqTJ3DmUTQF8c6hkSCud1HuBC9uBZvew02CNKH0m6H
XTvKG8CGQYiPQYzRTCtlpU30xYDO6c9LKiUIBUhc8xTvQ3DE1Ah9jlhru2Dk5SEFJgWZ8lqcYmRn
W3bTfIc8SQ0+VIt9mo1RgQYdaKSPmQy9gFRQ1Yz7qM5HCqH1Ee6u1RBOZFSCPTglbL4e8QjHJbKl
1Glvf0PqCMBRrvNrR1YikXu2okCFySQJrYLNis8b/AcgdHQCj+ZkbLIEKOrgGEE39XmX9knrxofu
vLsFOoHRe4U8KBpqoNzKRpdWm75pTIong4IGLRjMeteCYqKA7kbgW4dZemskElAySnE6Skp4vtsw
4nWHKD9kpAyhTL6mfKM4uS9ZiBBXK4tJfTG+3FS9VYAOgAlTR8NGGiBWfTEDNfOssw85v2+6rOBC
PfOdux2O6iS2y91NUT542Aqq/XZIH2P2BhpxQlN4gK+2TdyPIgjJZCCNqn9/9ZHhMXYJwQ/NgwJv
2hqsAf3wj1uql6WAkU+GHZ13YkSR9RCWKdfNCYrHrbnwpEw8MQmps9kx4idOW51EgPpm7osVfmPl
Kf5kD6qIsY7ABa2eOku3XbEiDEJeZ7w4daa6Uc+nEAsgrLJzgbrhWHku2Iy7ZEqd9eZRtYFZfu4M
+/lrKZ7NTRj9m8kQal2T35JwCqlHsAufK5Y6eQ0/82y6XSvjgxCPBX64yd8Hljssp1Em4IY0m/Nc
JuqcnSPWNDXjnIVTDm1CeWW0oHm1B0CGWHA/wOz4kyXW+H45g+XRCFC1yPd7M5vrxJyy+wFIZcEE
R4RfXKruqKcC563ljquu+clHdIObg/pGU9sxbY0mqq2gsLM1lGQYKM2Tigd3t9M4L9UomQ6+dXmU
vuZRiqg08HPsZuPxE0iFTUaE4yrq1qBGj/yuu7rPtjy6cgmxos1UJ4uRD1GN9iYCCl1UabjAkQLH
q/4rCTcyO/pCutgxlnaKnhUpH2PKCbY/aeVLKuA4iBZNEsk2XbeArnQMLY3kXfLWEcjWeQDPKoY4
VI3+mVhLv7RUEuVsm1s6tFaZ+TXJs2g5VeOUUH3xxB+629YMgH+hPQcFXiVdX/QrjBuMLx9sX0Q5
1XU6kKV62Z22hnRjALbyYIBKA+a8SPsfeVDh8yz2ws86ENJzEZ373YzeBeyUmu1l6vXAUUuz8MhY
kl0DDPET+P/iQF03cqIaRXjWV7CrNKC+GignelPYtqq+Ad63aWPE6cmaUZexVGNQBNmKlp6FvY7B
cxO9jbpjm+VObf/H3llDpxmf42zUpxUlmDM9lzbo2cNLTwxZCtvdDvzjHpio+TNvyPRzT/EGUlEi
z7a8eAtxg0Vjz7vQ4BZDgxBUlhT/Og9aHGG9sVcDtu2j0K210dzYe/EUUqvPDvhbs2BJC1pWPc03
nzWRo8pSrzNCiNp16Onukv4oyKDLyTYBq9xkuHFoPkeApWd+1b5Oc+TJSjo3msu0Ot040rwq4+Tj
CbrcCDKA7f6YeVky/aOAis3ooDeiipv0Qebt8zCocLhIQGgb3/JLp4lYz3LN7tjOlnmoBVn5rl+6
pvoKSwRCxhNwmuzKL1uPpIFa41jWKC3W7H2bfyLiu/AMvha9Hp0ZilRZajgYsH8JwvM7a3guutTt
9cXdTKAwgCHgPmivyYUiCdPz4lb899irOv6MpNIHkz4DFmbS1e7dq8U4ZIPBp2lK3+Rs7RsDZ5p8
oxdYdV8Zm4JMVdaxgnYe33NQh1XvNzjOVVGPys+zMjPU4bwwg3G2U9Xk6iNwNHJSAMJwfNDiX72y
CwoXbBgh27FChtMS7WHl/YYjHpKNgVk6Sxd2L1UhV33fovDjdQn9zKC+h9lODyjfm+ittqEa4mRk
eviyhvswtL2Qnz4KcV1SK9cCF/pzBDKZT4nG0s4MxYFJfemkj3aKCJVHepvwBsrkT3KfuW0bG+H6
BJXkd6zgPvL4QqUaLCq9iYvW2s9OSU/Nqj5T24dnkcf6EaeKZbyeyGEk7We3oD5QlNjg+PkoW7E5
jwL/UL/Gr9p2U7TctnMzCWNssekRQjOQvhKmrtiQl7igwE51S4+hnXSgDnSIIMx3sV3NY1z/Xg7a
3AKfzVrGWI9WQaXjg5aa3viMrLBdLIx4tGpzADajLgbupqpsU6UuCGZl7KHaHj1jyY1JV9S94dsL
3jsXc5jjte7YbL2A/qdkDzp08su0hc77aNycHQglMjah3jSd3RBco5FcdVtHxFIyxNaqOftOY1Sc
evYJs7+EgHEDX5DPmrR7jzvaW7oNatl+g3q/Dm6VMnfTlVkF6pZR6SDmndaGCbTzXiMhDII7JQhu
JJq5ddU+qEgP9RzHUHMBf4nQElVuL3UaBG+FmCZxvhV36S3yhujPH9I9L+a6cHmdjkvgCk6Xj30C
66M66d9XLqf33HtvieULgaoJRYMldlBYiF1a8aMzdU7MiXWvf4t1GR/dfP1HoahaG2xbEHpCTNAs
PgLf/cPIDiCcRpDVlefeSzmP9eHN/hLIBPLsVl+I73wbSK2u6Wm2Jhen/V8EIA1y7cDfliODa9Td
jANjPbwdzTKYWroJbOLuUvsiOoFkp253ZHKuVHz0Rf04g4bGsTbrKmoAD6RgfpZUcHF6a1ppXM51
ayMBxvNSTxyHfYseXLl5mm0Xr2F/Tf3sAFfWmFwQmfjJcrZzzXz83RxwLite42J+Uhkb4sAuXDoj
TZzSRs+cbGb4MSC24zrJGAVbYgsmqmSpNm4Ypsh/wobGSC4Bzp273rfqiEA7H2n45ITipp1HkRhs
xOHBxiIV9yLhonA8Chxn4bkCz/m/6snIG2GpMIjC6ErE+5svVE8bbj7e2am+o0Tfxmlv1ZcVgR/G
D4xnJbMVEovfff0C9WcxN7TPmNh3g0+Ouyd8QqXZnY6MMflgYDgylwXgLFGeFt4/pqUS1ZBlec6u
mV7CWbF5Gqvc6ZkEOp3DlrEV0ikwruCyqNQEjp+8ElGDzWLe1p6KcYP8xJBvL8aEAqr35gCqq7eT
jJq+qSzI+p/o2ZyQUG7BCpXR3G2G1ZI2ufkpFN2DSd2uedl0cSpkPlXJv7mCmnvso3fsE1xXNg1R
+l2uVo/BR60G1CoPCQswgFC8qeAdU9+WyyKSbSfuj3dNUrkQehErqiO+4TWCusd7MqfakXVnBFb1
4zg+IEBvdtE9e03aYM10ZTdzzIhso/LJAQvW3eToIMST5KYwwi2zVqJlPxC++Gb53kkpC6rynXVI
62yGzFBjbvs+mVzHeIWYzTQOJl6wj1goM8CxDEwlAcPDsdYRbBgAlEVUY1P/qb24lXh+5uLZPXmj
iFANVR5+jEwfBUVYtm1o/zoYyE8oWwOGXVt0nL3QDQEUcANWtsoYwJ4hUO95S9EcJW0izPzkx898
aqN7N/n7epppRuRKwUg/xJuHkW9jGez7KUYbAWF4kvpJkPziOp/c7Frq/MncK7XzDOZyLibwOvv4
3JttLPzxbsIH3CdmS/D5E8nzlSYLkoYa5Lo/ivNl5gDGC5IXKLl1bg9VyA2iBGzZFTYTWSFMh9jN
i61Ie3fNdv9dKaU6PeiaanckMKOcMuP6uWymKrL6WVcmyT1rTJYRBc9jMEfg0iN/XKa6ApYBiseq
uFaWH4Bf8Ue3cFNUjGFZaSKsLsB3zygwSXitwm3j+kTkjriVqkS6TcRouGUL8flv8bYJP3TuTAbM
4qj9eY2/YhYNIC1jdhnDYDdOnKmIqNtwpR+L85nEojRpj9Wi+0uO0HynwboEjSnt645rErfFsVOE
o+vd3pUyb2L/CtUK6WK0zc/edlRXADpLz6VN6Oi6EmX2TEo6Qy88tW45avNxLAzHlxv10oX2topS
iHuIvYQZKxUoOJqSzxTKw2Mt/a818el1XvdawyA+hUQcwfYiTpbXPPhkDcMLyMUlZXEao3XhKt2t
bVo6y34ASm84Yu71aKzeC+J/xuDOwoJqYhoe6ID0M55LLgdyXP1VzcjA4u+D+JTTt9ffECPs0aV/
P1zPszzVrozhjTnPfkdjuz/Uct0jZLqHKDqGvisF4mW4lJabLj9dWpb4WGvJ13VwvnRfG98ArmUm
3RkCe02ZjUCoLFRaQ6p+QtEbA+ugG+R5XVPYpuLKKK3AOO1wWU+wTJC4ze/fKQY78YQu1pm9Dnsr
SCFEbOsTcM9PabxOxiQ0/e/cpvV+PZpyyRMcRIGjeqRDmCnxlrdNxvWWFwfAyKxbkhzyBziHWKUf
pxhmFVcEkVcrZGT7VHEMSLRWv68Sb3Jv/HrMFCnyoC1Xh6AUiyl2dZMId/UwZHEYSnd2izzn6goU
gcFymRzquGBB0VIY6PRnmSlcawwl2+aZ+jU1wKIm3TxKTqVP0AFOnRKqBT4BOWnyJI7EXwFWDk+o
1mgTXz54QxwghJcKTt8qA7AnzChDmUX+PAD0MOzOimLK5k2ffC5uacyXicSOdZzePgpYYFOl3tJ4
A8mqBb1stA0yEpz3jbISkXw/p4vKt9V8KCUFf3YeTu4vormAI0VdtociGCcJ6wgqyZ7QP2q86DQj
QBeydPRZSi+EScOQXMDK0DyJZRsysJtAkJ45rM2lDXHmUZ8Rd1Y1gMWgFU/eH91zmLpwruvN9aPA
eHbphjRD1Jz0KLu40zOR++ZBGeoZtvjwXpnJx4FhCOmp5D58LsOApMZD/nD7fqdAkBGtZoDymeLQ
qQ0PX1G9BltRX6dBqAWaSMKUuExpgtOvl2iBomWEp9gsH0xNJ+x9OxnMuSlp8pV0DbUwaY6Vrwe2
wMF/wa+wrqf1pKu9sO7R6D+MjA9DLaFgxr6pTzzOSEs7S6TmBIB0FIq7kMSFhJtbiSTj9iCb05hS
i7n11qmNJ+z6gaLxpkOdLxKSqBVp/+aQf8uwiRMdthK6ct0Bdfal/b5fjE9331oshAm5mApR9P9q
XgHp/ILIxGwy6BGkwvPBr5DRqyo/74YedAN9xKRVkvTDc8pVEKSoL3AfODVRxYjYZAHNQBse1pQF
W5E2zarBcXBHLtOGiIEaPGrtunWHf/uTB8Zvhj53/JOLkKSj4rjYSIRXrSz5PF6K3jvurAcVhCMK
+BqNGG/AOHWOAOcoiAAtlb8775XhHvdtuVmOyEMnjKfnYkFEspbKh6FdC8yUpZHuOI3tVTsT5UIw
MjHXaW7ik9yHwtu9grulBAH114pEULkfHcGzYBik/KfbK0pufKM0LpvS7Mh2AOJL69xggD17Z3m7
fZd5Od7CzrlqkQ8N1E1X86nzRVvkfRtpgkKzSdMzE0AMcaQaSEuiwM+EtTKiPxs0OiLRoMDOKZOj
+cmOMg3Pe05oIt5Lfy5Mzz8fvLugqmExEB89hVurZedNxVgtFbQBKz2X3DldjucYRWbZsFEGA5JI
c74hpXdy7+xrxalqLNUbexSwknJH8ZPli7gH/CUrdp8ENM/0iZJLQqUGOGT1rfXENnFo06jL7kOy
e3w71NxN7ybhev8aPnBXjjM9R1XLixiCIbmXBmNEK9SJav4cvoUUlZivlq/K26k1SvPk9tRdmvj7
YKF7JM0lV30nIxmWJm89ngbajkDW8/1vmpE8ggfmdqoDKqDt2R4I5eUiu5mjJodKqEq7B2o0PnUa
X23azSLFSIUku/kcVIBdNvzysYbu3F0EsBs4Yab2I4T8piFABtC3gUeQMISsLo3K/dlV6RlGHCHY
NOEk5DYtLJA4oHttAHx5dnOW98aIJYKzT8D2gMSUFG5dkgZ9CHm3jw9E/4SfEE5xom+htJsOEPNB
2O8HGD31nVtRYmYHo4AJnIubXbrlLM28zfs3LhUvkm/+YioTkHTvVIX/dEgPS3ApXMavp/Mdf8TY
NRAX76d+WWgKHTW7ROiUIRAPqp2/uNrH09zEgUtQLXQFHASsK5Tnf25QCqRn/+hH/cGH1LXiEv5G
RWDD4VHpINIrryK/Vsw5ljFSVtc9jF8BG31L5YwRnGQIA1a3u14ks5E2XPy05dcgNHqWT7w457YX
lXl7qKdJ60Y67xeZtCAknfxVDJzbo2QiUlnd2I2HLZ//q0zoG8wq6OUAUurIZS2BMYC70yA5T4L8
gFNpbBvMadukP/2otrkVB0wzl1NAcpc/ecLz3MNLCppZRuG6s3fGB+gaIfQvGI5NF95o86YzTlm9
mL308pH+3Enz9Jsm6KKuG3WL1APn4rUDcyqBfkG4ajf4hADVTYlZ9h5NnabDi2evp/tZm21oo4oC
za9bm/xw58VnBoAi9vQLnLWVG+mUvwFtUbPbP69jDrttCiMm0NeEa3iKoPD7cTckbYNVkSQ0iKPN
IIMSFMUKK3sS6cwZeETrrc8wyMPJ9FQH4IXZs0h5925+eqnbCIPB56ZSg216CGK6uGFsNnqFqO67
IERLrBv3Sg5C+Jf7TbnXWzZcGmzDEEBuADYmPHkqeNeAbt6I9DhVbbRjMwD6SPR9VfjK2cy67f7p
2mvNhFXXmE9SRXguY9x+chVTF0e1ZWYV+kqv6hfaA+G6hi8Afzea8UuFUqePrcNrTM07oOx/ml3v
/D/FtPfaFaiiB8gMBOH6xXc5005GQFMrFhj2J4vPb3ipad7KbJVeFntXHNO/FRrQgccHyJSMx0TW
5MC26ZJ966gqU3SwZySXZ9HL7c8o9NX2Tx+lcpW50rVebnuL6HQYZAy4EvXqNACVOCIqexd4kLXd
3BB36W9jz+pKjz97pt1c2A3iW41MPOTbUcvxflyDEA5tmhrsngPlxbeX6mBObabSSl2CAuFjK4dF
TDLxjetnHh4wvOVW8D/lG+akiag1JQclX3B5WEYsW0f8Xx9Yaz+PaGOiPyvmieSepPAuFuWb3fWT
YKHtBtJaJuCU6NozE1n/3k0/D5hPZn0046VW8+n8A7Lp1tTggd9ZHmssOa6x/+3c+RDDMSO5h4k3
tXwiKwIWXOvFMgefjgBuM9/KKJ2hOo1CYezGwYZS6T2IiMh3LhGdBEzgcVAoda4JiuhmqsmwunAj
rvsBS0SWKBj2aJW13e603efEo4UhKVsAK5ApL6uR+Nj2DGsRqyrHcR5fUh5J8uyaaomFtxDvvP+j
ar0K82YpNkLTGf+FQ4aUJz7zhpwoewzqwctWgFx+JwfR05K4bUMK23bI3kKI6L54+Y3N2K5KJsJj
64OAwBdGIWgfG1tqIm8Wi4IgPeoTkKjtqtMa5BPcDXvySQvDP0QAix+pz40cONAxnC79ZlDzmRcC
2csLFdg4McHCfTihbuzoI7MG88iapuSNDMaB/RHqWNafdfg7gFQ6xHMD/RwVA4t8pyzO824vg8HO
JnSESWifEBABbBeZ8n1CzrekEoasdR8fjdCMuHWPScQaxy/DQ77B75z/Khmg9kChj+jjSva3NghU
s0MN7/OQUqItzgY4XizXHnAE0iJ19CE4+c4/0RgKYzYKl4rPgHqaJb46z0kw9F0oePGcJgyYgbHu
UuZlakHzw1IeucJwFL38FJqjYmVCtxcP4Y4X6giTTNGcMZgx9I2j6ujwbNQlngoccX8UTw/d6tiI
QSqjNFpEVjizJN84dnALZx4oozOun4WDL0U9I8kmPxZK3q1NnoWotKduK9eNY3LLUPd3CCNGczrk
xMLKftDGWV6lFxXYUFbgyaPaMcXLpdZIK2ApInqr25ivwxwSYJSm11+/NMip+TLXhIqagOTAbk9q
+1nQjqUFJZwY7ZP7p/eTFYRJhEX9hLkAmxIpRNZdC4TBhfKIEvQPDXNRE8/tRQchpukIn0Lik8th
M90e2VZjTNIb7I7Z79IBgCo6gMI2n//5UgSlqnKr4hACFSnmbpvkQGEN9hsfCptOS2zk2S94/ybS
yxKbzmtHJv1dAvKC/1FwDv5BxydxkIPLpAjFGOnxW9GMEZo81h/JAbYqoHKya8uAqKFS2g/VBgJC
0s4F8UU+Fvkm32uSgSb2GZPiYfb72ffZcH4nvI0afkSIu1cjjXgYuo0CFBy6X14Nal2X3S/8xra6
Btls5aB5VqsSdlO0JIN0ouMTU4jOLe0S6lXhd+GtZFXZOTOnc3QdMaUjPbJTJPA7Thlc0FPmfBWb
s39lvDoHzFTYeqahSYliBTl2ZYYzeI4RzIIviwD8aMdIK4ZFVksfgeuL9QQl9rKKYGReAJAX5h1t
ZPJsb7Bev9md+v9bQDYLXUh2/HQwmorwtg0mInTQznuRpDCIbkXVypWgkH3uzb6MV1CCT2QSTwOu
apjp1ux1ciWyNBvA64rDgtD9RtkddAZDksrNIjmpbCrG5j54n8ttv77s0bFTcDvLWjdWDGXCWpWR
egqcqPScs+sAwZGsAVlK5GF81buC18qpfPMovbHv2hYOgSuNbVEH+hgxUbOSXs964nHJV3pKydw5
3998WVqLy1yz7gFYuRuAUmF0wAVnP5oxBYLYiZzZAaAGsnXNLcgOgX7oQAbxvGV3h26naqyvvDtJ
BLkZGmfu3xpatN2eUOfim3X3bVcCGcgY+bL1m8LjY3q3XfQ7KxcaTmFIgLyUK0ypWnAppVja3BBv
c+28MY4kaRFFJ2Hp56chdBgEpV4LJ9TqIQhqo/23IezSktaE6b5TGoeMU4sUVV+MtBx0XT96m0jr
QzGfAuNYU0iOwUyVLUx+z2g+2DY7vusulOY8KshFHGgBd9woM1bbpMkHCReiEYTVNumHTaf7C3xh
N6ZgVm987qeh0eFYu3tJcyePlkf1KnwWRCQIXacb3kc9fC2Tym9WsvszaAh02AheXy+hxwrNL0Tq
qzsIxnoR92zqvP2EMnchyZcLQ+h876xYMYKrRkgH5zlg9MzS4zYgricFEVgJ0XivjPg1FLBonC3L
9+xc8pwRiDS0vdiY0tdx6GtsO8GVPkuexAS2kjD/OgjFBlUaobvlEh+aXVt/6WbPSKpb7xV4c8VM
QstjYLKTpBkV9JiobSfWKLx5KNX9Z/f2LBVXy628DotZv9TDCT5V073CSDD669Jfm2hc7kkr9/pN
hxVXT1XW+SCWHvWVs5ykHEp0YH+EKnf/Hw3DdtJ0YvfZ+T02AJBc82NQ1jV2XHGTwQLs4buL5YjH
mOOS2XMLkKfujEExIs2C2H4LD7iBfRhu9WWvivcpmXoxV2oUeYqosntmc69QdKD1lAYV7coMn229
hxJFeGEaoaoRDZaDbcK8ZqURXZmrdp7LXfA8Xnw8XAqigSGBtpXwKWXWjCLXdEs+6fZvC9M3ZguI
gx+1tP0Q4wONn123bAdG1D1gFagFjYJHjZbHMKw+qelAZFRNWkz1OOFQD0lOA2BIyx9Ij2Zhslqd
F8YsQ/hd3TbLp+dgMPQERqdRAUSpEq1bHYHRx+TcelkUL/Uv2IPMq1c3HwXG30uh5R260p8GFOQT
xuHtanuhJb6RErgxTaMLU1RialThA9z9HzuqZZexm56mRZXspDe3u80Dfpy27zXvEfRe1si0CFMk
KxK46dqt8KTFMOdhZw3ugzoFe7AAIKitgPgpCI0WGaF5aNbBH5G3jCnQ0cuMgN/rzqov19VrXvtN
OIdpv5Ku9wmYI22guHGVRLyfQIGCve7+FKM1qq0fiK1CsPlAp8Zl6S7dxCnBjZn3veTy7kkNnQYb
t2GHvVEHJrjk2uLL6hfJCeZnqUeCORlerR/qnM5UVgejIjsMLiPYHWWZt3BqLcmn2/pr4WAwX5cl
MxX3PhonAh6Mq2aqyZLYuA+x5lh2JG2YTu2NE7VAmeY2KgRsaoIKtxlUSHJYlLABnbYcaXOKE72d
Fm7zWwUF1jYzT+UnHfTyuhyZxrPN980g7affBpVahfPSuW56dqcO1YbpHPRqjNgwKGS1TvMLl3G2
iTWrq3FS1W+CGNptwlhDLsuYKOmjAZjbM1LQ9xBbXLEHCmBSN9JfSnof1n4xGK6CHIOKjanUVHGJ
O4OuWCevI9l+rT/rikrH27A0dsYG0Krb+tS9dtGvsE8MgO3FimmKPKXkalE2o0S9XTKb2LM9fdcC
IuBKGNcuhK8jcO/BZy5RjYH8/m/NNxUWt/MslNJeQg/amITLjGEl/Vi4DIi8kNw6x9WVuQzmTEUD
LfXg+Y5x3bNGvSg+AOoA8YQVNCGWzVvzJEeDzo3MY8I4sXbllDZW2qQtVkCmk+/JqejBFT6gA4zS
b8pd2jJOK8Weo8A47MhGyjEuA5whKubYIxoMGynJdA0WAwnENMkuVitbi2szITLH0U+KgA1l0clM
OQcxQdofZLRxSxxv3dw2bCxzpDFzX1ZqUeT3MKAPJV8u+zjzddpcb7eOyz3tuCCuQHX8TLsEUiIT
nHfvwqsuAi5L9o2B7rU/OcYxHVfWSgZZGquNN/HTdOesJl51SMJOHA2HdzLiZuASDm7NXlHE4F5o
h0MFBZHNvUO2TrjbFK7H1Yu9SBFtGL3Y4cuoMgJjIWaNicJ58cw8u5rfKp7oOB/XC1GKglaWtoh2
t3rmxYOM8lHYa52fPrg+dnJZwT/w1lZjvV+W9bwOdN7hFDksv/vfh4dB2xVGNnab910w9+DnAe6v
oEOx9SaCMZQsui4BRuhCExeuBXPXHziVMMher1piN5S0sSmnXzIdpL1gEo+QjqwHmFmKsxgJMNSl
eK66Kb0ur31Cx0HBBe7HfXZNbNsSlE3Mfbh0I0Ll++2AjYU0I+OMvfmyxpLMryhqRmd3pJtxBITi
zNe7CCgxzg/6/PyZcv9mMplQ3g9h+hX4GktNksw3XO8mAt2ZbQuQwqJ9/zY9+FRAYr7cc1D2TnvO
Xp35ucgAtAXDoeNqLJXqMH55iASqBSevErukq8pBEb1CpLppgkRImGnECctNMjV0k8x5tKQxxpAp
3c975O3jUqEylRcIhGZf22r1Q0B3r0MOWbNJEx/7ZBujzeM0xaExetdT5DU9pENwFqI3IXXhEGmS
Hn7Ot0skmjEYoRIiYJ89lJKjolYa4IPTCSHQbR1pO5m2zj/wHzAV/fg/XrXV6jjUN+tyQdsoqIf/
SAdsDnOm/eJHfQevhtJhSAjww3CwnUXQDqdttbNPQdIiFIAMxQoQOsDn7QVDkwPLa/FCO0Xx5KHr
tT4eJ0j51RZISYpxc2zcScn0UFvljVDvkBs/f8S31v/qMFoUJqfFXMROHy7OkZz/Ay7CuLm+pwxN
wkM8iR1BJsYLN+PjbdrSNX/G/x+cDUuT1rWOWg8PxCGebBLG8kJeHaECmZ+PhVqgh7q42GOMBpdp
0YxkwU3j14XiiQcC/DM4+kJ2NgHLZTnUApf1TIo9GpQQU07eMU2Gmqu5GKYlx0VEmIn5skKpjBmB
cc4MDPusvpbz4WQ9qzkOl3paFPMEnx1c9Tj/ZgGIQxMrXZNbgo4/z6ZMm2G8ThahhVWELzwybafp
RKwedY2DAp3hr9IHTRBu4U0enauPVo8D00mFRKXccTFHSm1CMu8tItka0ggRgy/nL7ccOyvMONwO
Et9sSIQeUWkLA8Pq6PJhb7YgVPc5fIpbKDFl9FvVm+pCvEFodNoqsPckyd/g1gw6j3HR4bj3oA7G
ocxH6htAJ4J2hGIdymiDqFfGcxq6Dhz/CpCZeMD5ZkerqAsxkBIcJJSMafd9OlX2XESHwEfDKG0i
kmzJ5q2jgAOXaLoSq+5G4/kZAUUOP9exVzXs+nUslXWhUVcezn0HBhI9gn2pDBcjyoOuv6waTA9O
6r8eTTY0txqNtM/+3Etw9Ja3K3hgcPGl9GxXjIMyXE+bF2QBXOfGICDvlxSvlQdzQYvuf5czGj2J
rcbgQFxa9DU7IBRKRofpdoCtSnTSfnlWXzQvR8d5DU5V2LBlTl5549HL+q+C+Sf2sx1bZOBwgKxI
XOSnDdXXf157fgL9XLGGFieXVtJf9+UXkFL7hmS4/ku+lfuKuI/+NCF5UpjlacGuRUpeoP+dKVuK
ZBJORNA+LffBnE8x/zqt4+ke2sdH7X0yDUUq9MH4jVVNISOMLJYfDA35EUk4ZBpin8UWHHz1C9cp
urAtdWEzeNQGrqomGEmBR2yuSHHqpSC94JAo2TGhGxrYS+/j2LAsObcRJpkPotd4/w+nI/PHieK4
DmQcnZuMBaZlaT8Qrnx5rSthc3zYDNMItkyIbrFDT9Jy9c9SGgfmQYvOW+UIscGNo+vX8MoNJf9E
Wz9Xs85pdNOOnjawEuVI5rHNxBhoFuRA5u9ARC9XgHfW5OGEFDvWqef8PbJMf9LOPlrNnHiJ/yBb
sDa2tNOaxKv6o5nbQcfdbaaMfaysjf4XKW5OM2OKb+fXwEydAsYukbu8HRF5Xo1Q5BpmhbcZuzOO
2lwvWouBalNXprtsD4IupDbfwaS2R6klITKfhWeDR01eAIG68Ow2P6gGQg5sAicjKdy5rOtI2+Iq
RAW47c+sSFsIualQp+I7isWa3to7knH7JN1gX5vAgUFQK+O8o3QTKnaPjLa69rrr1jYhBvQuHCHg
b4hpObpq3b5C1FzXvoM0bilMAFmYNvCDnRy/6+CjZOy0WL2ivu0pClN6/k5zM4LQ8BJ5V1tOcxkY
Uf19LmcZUTVjNOz+LV3m2h9bSztGUqTYlUlytWKRk0FbK8wlHMRbA8lP2/uZGSS/Aij0qVScV9kT
vU/aBYUhdgLa2cvavnkEGteyzXEw6NWeno+tUe9dIW3DdUoSzZKsPChzVF66LDPSv0fMOYsEVtMU
AKwmCsCnvcT0Etgwb5h0Ogvl0O5LHqm/Zz9dq3lHrv+hO41XUPxtvrDB5E2knlt+Hr1zLHKOhUBU
QiTsvCs8TKoCdxxhm3ukj0pZ5e3sk00XuuO2vKnfOQvQNQ6Ql1yYE0uieZwCAjK0yL3MMcut5+o6
iWQIXejuED1h15KqNqnxHcPqxDizUYrYYLPSdpyyT7yssGYj5WyKKb5vepzbZl1FvNn88aPJC3wM
Up2VqgLl/kUHO3kvomnhBQYYKFRtPmcuz1DhJqr8wDIJLtpaaIMqz/p0RCOrtUvv18gC7K3yRvi/
XHro811d7ydjRNu0iSVUXPdDIDeDxvN8efirTZcg9Si4nKFBe/Hn3nxCwFKK3fdzhdNJB5A8wa4y
zvAItgmVYi+VVhNKxFCz8MHZZMXaqLli3oOJ5PvYGmWoYwFdpMGYfQ3GyA9v33+MXGWtdH/jcnck
YsKhDA4lFPXGy11v07uz8VbWpy4K6NU9Se57YIsPK6vhbNwyXH9DQHocD1tEe16aGzKHzTqbOr9z
6swD+G1tovQWhmiFgQqdD8D05bxLkFm9o5apeTFffwcwTn1Hpxd6aFl7Vg37ttoYiOO0/9phXKua
87Kv2A55m2SL/onTyj+dwrRvzVENQxrkw7N9VifpEEQRjWSZf69zYQH7y1JdStxSK6BWQ9YDc+6k
NFElO8Hgo12ZlhssLLcF1daSSDX2YT2yLUQ3jMtqcR9QrmNs7CmEQssLrYEpBfmoji5FWjs/EdDw
IVanVvJypxnDbZ91uLJldRbt+OJ/+NMrQ3gTwB7QVs+fIOOqSIj+KfktNqQ37YngYVBuPH8qQFX8
aiJ2fkt5edc2ttowsTF9a9r14KyljW7eVf8OmyMIr2VvzvC+VjsPGAQdxJWW4ANbG5n5/vCenYkV
JGUBa2zVsluwCZwJV1ARLzXlobzThwTS0P1J41j2Ov53URCjlXY6Czk1kCw/42//hztbPngVMauf
5rPI7Y+sSUPblu9Hwm801p8hb/ox7rdnu3cvEUz/ClgOcpZziSnpKqSu4tVOltF8iheCT6be+PzF
nEkUjLeDxDp+q/ZT2U6ZsuIdgBdowwmJrWUALGgzn408p0jNMk7lBMIs0picV4nYABOFqz9ri9Bi
B+kpEv+kiA45szkK1uyAxTy1AoWa/0+/t4YGpbyKrbwKAw56kd6ltoG+rMafEpb18nrxemKflYZW
QkwiwyVZjlC5K8u7u256iGsdlVy599mCy+r23ZVGiBQvE+43YW9+XgR4sfeoZwdFaM/6+LyxzD3v
Hu4p/dYEgSFkgFS+v/KOME87YKFzTe/iCq0NTyG0RIqpZogUb2MvqtjgljyjnooumRSLJiQ5aftM
02ZgsQ0u6B0H+J/amvGO4HlMbVocCx7yl4w214Lek8wcsP2C8+9oZu+62BSGfFSFYMfycaojuUCH
P9BI/oG9ZR2gM+kX5DxY0JVvEL1nh4b8QPhMVukbXC+gRDgCQLoHvyJF+7a07YnT3dsimAazXCKp
pL+hG9LLWZTIR6zwRTNlZ/IUBdeTpzTinC97rVpB4DKermQ0NClXDeJ5C4SbGs8ODzlEaTXxf3dE
PU7V3f3NfhGVZGpqNclTQUqxLLCEeA/7LJXPvDpIDwNfPQN/OQCrorbZZRvxVxaREBV/i7uwH/UO
qLEK6Gwf9joE7VKo09OlWxUBRicczXY4gB3yl6/+5srKe8Sbyv/oF5ycjTq1jEuLUNqUDGJowHYW
SD9rtTNTLW8+fJJTX/vm/7GHnXdUvdCfsvQ08aE4Fs19QeOsVjHXdGtK4BUOHFwadJFayE891uIC
AkBsKv2jiEwj7FUndzVkqyK2UR/e7WFhh6T8JFh5Gf69EJtCTW/GXzxN0WZiLzNO7O0NGQkX7i+2
hl7QeRa08LhGpejLtQfvawHl/f9SpPPFeNw5szjZwY42xgs1cCdsMjyEQtDDoKv0b1jU6wgtI2x9
wU7RXuJR0GgJK9ikUdulnKud/rrN3Jgh7qtYqoVibVWha32AUw10jPxx3vjzbVgu9+jp2Ud4ZU/h
GiNf28W6mzkAmS6ssYvo9WQLLkxJ6MVwRu4XVl5TptT8/gwWV7AhXduAG8etK7QWHcicS5hq7ZXr
Jbg9csJRtPbxtMrNVqrg8tx+PYKhdTLZU5JBBzjyrFtLyzSOIL/kiz9k5WiWSBsH7ZPTEZGXcWoc
RbQcUey+reLjK/9UrTNNaJX+zGi+jG46Ju24klmFU4fYmRgtEEiGE8CGIMwE8H2LAb1ZcReRAeb/
e9ETk7GVeSOi4FimSZCyb2iipt4yU3ftKs2xLV8B6+Ziwbr7g6+m/O0kqICksfdH+gU1G/UeEbSl
de6Qa65pRX5OLg5bfV8T9n6mzvcA/lZxp65sUzK2Bkdl6yOtbGsHj6MnL5+QDSTKkAp4rueLOJo3
mP2vgnBxW0eLC6iYiCieWcTNWitPT66aGftXQpTKEqR2iHrEpScZzU1zThpR1Lt0TgRhAXyzD9bP
sDAqYDMYHpgZXKAWaxgtEMZvaPiPRTx4Nei8NDNrIzjICN/eI6QYSqtHW9zJZQlY8OIx3r7xvIsy
z3giE9g8D0p0Zdzya1BcNKZbBf9JxsR7GhgCLvWwKg/keSk8K6Z8yYsUUrKgy0wm6hB+8UL+HHTQ
yr2LZM/2PYZw42lGFArF8xdLGSiZBGXrvgerA5GiFltkrEqBgZ+a54lj/7jTiKr+WT51sG6/VY+3
lzr979R514xtFNtk2osPDStIAgDQhh+Uw5KRCEbZ+0IbuWeTWY+1npXJRKgNE1UC4+mDTIVYPvYM
N7C9MJ9yfWh/jjYoR3hD4hkJib2Xy8xabxVRZz7DXwFLjatoqllmCRH+og6XpT+B7A5eqE75IYVR
hz/Nw3VOKMiQpEOexVqIwzZLcL4hLODxUyausELYlweLp3OMkCXOvGFPDEHELmxElga57FqNOANi
WFheICpxqiitZotFx53k03qPmzELuwT1RMrkdthuzf9H3qeL3O1d/8wDeZ0BO4Ht4RzWguYJ+ofI
akibruZdbHm7DVWL0kzavZhF0zfq8ZvwICEa83T/EnCOv9bOragK30V0S+fHnzZ5U2nXg/EURyhO
Rsgu/KZcd1wZLYQkJvlCxt2m7nwPjfmMJdHbA3knbUPs70ohQ1cYeCINYn55GSniuaksq7A3xH/a
+bM5ZgRnKldlIrodnRnvE+zawVT45syO7CezSwFmPHUUio/dgMs1WgolyMNW8c/zb9hH9eGb4hFD
BdgcF67Fx0GStGwbt7F5tb1DHeIaJMbGpjhjPMmbVMgRNxNNs1EnnrCPiWhFr/esW6vV+WZpnRg+
5W+LQVeAVbpIg8/KXyQ+C1ceqdQff0Gu1m7xXFz9/XFPuUaMdv62SvEbUwHEyCWbPjwHts/gU7jf
P07k0hNKOIZgL8LKFD6cPNldCP/brPUsSU1XV8R/PEu8NwFH9yBUBuH+Q3y6t1zUeYrgwXxLA91V
Z13q4T6zXArbe3HgKH0ElTwSlwn9fMwo+0x2XBiVqBB98OX7dTtox6Nv3UP2pmfQQUqaYyNEaO9U
xOTvf+jcBGIvwQ4t0yPn5K4mcWZEyUWat9O5QM7ZPIgCorpbERIylXut490qje0p6LtZaKcJ8/Hk
0n0baLKt3J5bPPugHdLYRyG/uXiyo7THozSa649PGPWY24qmws2Cy+Ez8VPVBHxSnYyLALmIeYqf
j9HfOID+SM1AlYzFeFMc8p1+P9XZSJG5S2Ox/Lokmo47Nv1mI5HDWnZyNRwypdmXLOfjoU3SUSF8
Az8NC1vaaWuXWKhNSYmWBEFi6I+c5TcH9g+hVfpXId4QaVCsSmLiTw5QUMbQ92GBU40tqa5ZQU4j
sN25UybfoclVtX67J++SwMikP9pkAPNXv4kLIbfKQTeYsbUdSSO7SbDVZplEI1fRjHtCtj0NValG
QjPOZNU3bzmEaX+rap8uh2EvCm+xX6XS0QtSXKD2KAeM4uipBkvr1R1y0vFARi1/dhz8esG/pZPH
m4F3REGjc9dmOCfmUjbXgc0rJfIueMSD/NYdYOdw2N/d3gpvmrodMLSX3uR4zvZcUx+IMEWv3qSr
awfsE0uaUfqowE5ZC49pd0aN+olGFA4ne8VtF/pQRJhUyJk5g51uIwCwlvrMubzRy4pnuG55COti
IX4mXFYvOmy2Lx5jrXXA1+CKUgq1+QcQuYHSf+QiwX6xZEAlTdA+9CDZKrlMP71S+bqukXTMDZTS
8zXaAZZXpibsjcaKRQJaWJ2sEjZqdFNh2eDVt5+B7Z0I9mkrddwSUPXj1ysJcSrNgp13N8bQswGM
6fU3I4cSdgWkYce1u0+oSi7lLyhufoOY8mxm7oj+o5q458+8bK9FqGAGj0Jb0sNJD+bOKJoPsxVX
yn7RDR0SyTG2FLJrFPWCw721A3NkASTyLLiiaORh/mvkkZzF/Y1Un22uvwi4YJ+BE3CWXKEzBpQ8
yhynktr42uyJF5bFj6L7BrrnvXZZwlh1iRzqAEq6psOQal0fEBdZZxpioKcmYwu6D+QYIxoODFHT
lneEp3KZqeTvrQoIWf1bSeE4caQQ1bZx4x38iSnJJ6L8+/BbTmaBp0birz/gXoZCgWDT75XUsiqF
mM+iPcEeEZZJ6ri6pZslDPEE827TCz3hPNh9olr1b36ISdRj5aOg09JzxDbRkNFdrZ0waLK77lMZ
5+pwpApZpUSHJlrNZ8oIO54Af07NW9WThtdQHv7SIYCdyLLlQkh2SnElfueNanOhwLG7pFbCE/L1
wz9k79YQxI5pGeuji7Vk6DWbMlxM/PTe4To9m9yUInBZps2QdtNqROw33VCcOw42+H4+G1V8rYhu
aibHuUFm3Afrb/Hx+5dUJgvHDB6/IxelRLMerYf+IfI6dy9o7hXTvnXDoCNeTr4xFk4XYweV6sQt
vzZbIGfmKrXhUkh2tEHKosEHbZ9inHsGeGrkzOvMrtFdEd1DxxhymcwMHN/w3cPTPjBjeRV5Ypmi
SdvRoHt/5GK0pwZQYgksLORI5UhqIAjugZilr6EvSJ87gM62yceqObs3Sg6gtiway0dLXRE1evvh
23nYR12EoDDtF5EG1YCzs4nXafMzcYInGD+KXxFYn57zsaC6WuFaaxvknNbGL0fKhFYMTQdMunph
VU6ECJebVw7zUxIPoQrULQgNKWz4C56/09I3C5XF5JTMnvEq6CHoMOd0IDEtZbf48AqEwNUz5xVU
7oIYIj32FM7RAFIPxOJKdtkJYegEEYFoboERWhtf82akfUjH7vuwpceVu6noS6hz5pahH8w/BLRG
zRpcm6Sab3Q5BIKKzjriUByiaITDMSdZCjUxTH6usTrdQcPw8iUGzX3h0mhtuTAS8KAvngFdZbuw
L2jt36W3m0lhygK1H4fZnMhJlEJBo1r3K5PTYK+UhAg/LoLRiONzaN9kdcCbpsw8WxR0Z5nO/mJ8
AZiLCkahDzhvr2xJ/cH+dkFTvUdtoRC+tPzFaaZEC4KCkmzC9zHtdtRzWtZkJBLIyCQUskraLnIP
guODSJ9giZQm3n5qmx7auKAX+I1f+5fzCajCN4/cWXVwXsvIMKpIpWgQyApgPZSqCQM41QrlhvYi
MHdzBKS7iYmP2kpi0a6f5PR142R1BA2LuQPS7ZDruzA0KzqE0kckun4uaUaE5N/yHBXCRO+b0zI8
LykvK0B2nlaanCkqVbogYRR/l6sdSBB4R576r3N56T7CDcr2dpqfgKR0JjZ0pAkjr17p1HV+8UvM
CtTB1P/LtXiHJ1F2vOAktGuB0BT7OXTAiG8ys3HyqoLmC8lTDxz6qE7QvN0++07KYqCi93j9S5Ft
D+HgWhJHvN/6YvAvCmu105Czz8LubWa5Yx0sTFK8uXpyRH9/i2U82W2f/O0wO1/bfBUvispe1rPT
0no89MnOad4fmqWwuaobMnkJ+4e9EBi7SKhCnZYcHn95KOXpYayxcAk6hMAZrllPN9+mCPwA3m6T
cMQkFUDASCgbSWDNfyDhECkzvhN/87PTtuaN4bvBxCiD6u/8P6gGaFQsGSPJQUqQlho/tX899frR
B8YEiX3fgk1SrUr366/f6tFL9QxBz8y8TlRsDBl+rAM9JRUvwlPl5u1VGDVN423QylQ9zGsApHPd
LG/t9XpotJwglOgZF1iqE27NHNPYkudI6BRiUUXJmE5h595dnnKQshLA9M/V05sTyjGzbAhy4uQn
YP7VehwP2UjBGOcY4pK+drq9cMiC/krtOSnUUNvvI1Lzk+IF8qmbZOJ/iqhkH6yVicNVli35MyUk
v7IxLMan5xd/YNXLwZI5H1pShnNwUxvbZKN257/jTtCO4vhwYzPmRIO+Zo+RrOe7RDWs3anmcH8r
h1sr9tgmFr//zgfkuYmqPSGcYJbKhhubpIRWMjxQYjQEkZqxEuUYoiAT5XEQy6TanvgpObAUgmLV
bO1foEXtqd0Mhv8ihuDogLcyI2q27lcWKyXSZMHBaqr23DjtCYMadfs+UgW3gOnJDxL2aq8bY7CW
34MLIrsiSnj9RVJPAz3oRR2/PPIeIryPI17nAqmFv88TJcQuaiYC1krNNDVKknS/y8KMJrO9KEDR
aAK7kOip/SToJ0yxJrKWnfaCunOoyzn+43Nbmv2cikuTY+Mti+Pv5z9My1MZb/CmNbfwlJHWSZq6
uya1ovQ9YhJi3emkpEaG28kF2nq52q5nsminhy6Api5SFCXCiywUvFe+sLGMaCogkmyoNNNxGaey
AscgtTHGklie6KIBZOZoJFB4GTN/E4CH4y0q+XzBH957TKXwomGx0IsKVqUWyCOj64zpSDotjodu
6/Ed1WzWMjF3FcK3FtcsPul8f407f1brdnw3/Wm71uOKirhL/tzgU/ujgv4QrVCdeLv07DmevYsy
GF0txrPwGBfwUUjGsWRYOXdioZOsSAUEM5jO3d1lajlgQokq9aEWmXe7cZzyWVM5RuyARFoLhYKC
0Um776L2O+Eb3WLExIZoIFbyXazwIbZXTAe2Su0FgI/LwXnWtPjEDQ2gboFvTn+SXH1N+NxkWBd0
mGNGjhmz5V3a0ieaVsKIMdrvFPDYFg2x2X0MHZw8xapR0yToKq0YWd92Q1kHTpvd8h00rg79Yk7u
2agtym/RQHaHjNXmOLCmf6EuEgHqwvQPRsyKNMfQ39bqstD3rX0fp4uDUzJnohyrL0RChAodRiHD
1DSTMJPIeTUFperNKLynpMco/kNZyjxy5Nm499rP78cSFbV+dvCImGHLfOQLbJv3sjdrcnSMLdMt
Lfnl7ON31QHQUY6tH4Qvv4XravSrY50O7q8OlhtNyiehqVM46aFJVTSAoIh82q3DqGed7gCnEObL
irK67slwxFl9rfaEgy47uUubjPu57yYyOhc0pzTWC5P/UaWPDDAf1zMSLKhOJWWtH7ncRq6Feu2k
sOUH04bVVwbpzBnkwZEFd1wCQCeD/XB3ZoehIp4HdYWsJLgaZeEtoyMxKZAv7kloC/d+jbE3nkqS
adovNZUch75Ocx+Q7t+dCS4Ef1IGeQ3EueQUF016v+yZtvvpMCf9qNYz2kzphquOS4s08IpGGs+x
QCIzAO0KKeLi7IDJHuX22H9/3pj7tW5a4zZw8gRZSupb1HLOYMuxaRYXDraI28A7ZMZelKsFUx0+
q4lNI9BnjsUaBrWIG7bBsidnkXIzTOEP2O29G0J5v+aweASQlsf0GjwxNVKVgUhH2Szz9CPGUkCZ
QiIjsVM7QGuhQ8pV0CFXt49d0uz/Y91uoekTzF8Y9PEBMK+DgbBs1nn++L8PhvvZP0fwnCgg8GND
TiWlcP/lNtBPMNRospl4JZDH5VWeJP6ktbY5W9RNXAMQCEMiOm+HSH/RzIdFXoVBVHHKDnRncLuo
vFMAfQuLPl4FELSI+wm9a9FWcpdZ8qe8R+/MfvlQC+VcapVbSKvHFkQkmBRFYuuyK49ietanTSkh
jotNDaogzNW4bEZUh4FN6GEAk1iN0p8E8+JFqPyedMQhGeQxHq1yef7riy5mQ5rVCJHJwej4oZGm
iop5JACQ0AJ3LWh41IHPQOdli82hy44Q7D8TWxzVRQ/dzBmNtL9amu14Ts/i7Gy0MqKmz/xVRE3L
gl2mrr8qgxquAIolGeFbgyCMzWrwpw0+bjWsGqA1PKIIo/lW05QQCvj+DKvgWc3y64K/f7uvZhYk
7an6PN7f6ncAQZ8HYqnfb7rMaJXQWtUs370a4QVMFvexIPoLmYP6apZaRiCytdjoGIf6aZ3mIW4H
LWHrYROOh7gfQs5c7RNNdJfS2elbiiMniktOtYsHWIZxs9GNlIxPqELgoiLVjVhBmzOnDVTKuYX3
YHDxXrZ9YHDhB1hrrKoMo9KgD3q8HQkWknIvmcIJCHO2RuFA+EtP+IriE4K2wOLYmBdGI1C9XXfF
LvFW8ic1OO1CoUMtRVT4fD0iAMlduCUE1bTXDQyYKSLpJjznQ778XU7WC2RLryaovdgf5br7t5cg
d+E/j53sAxnFaA31VasN6ghqV7NxfaRIP5kDlsfdnmqBTGKAh5OGRVP+dPm4AMkkY7vhU6ZHJESG
ZG+yJ/xzBB9V2XIdK01XS5Lh20ZANlP1Lyy4iNQL2UG7G7tW2aB76k4CGORTF4yL5+6CPHy83GEO
KD6DSdQimKYJOVMKzza/IkLuKpR3MD/D4oaPMiud1YjkSHsKWt5/aC6iHDFU4AIklXOeraCSrLFU
Y5mkLPuoMJN38Aw14j7pd2ObM3r2P2hNOFTeGAxn56ozFc7sRoYFa5/efC8ot7TaNl1KbOKK8hQb
53P80t2fNrNSpi/053Egh2kAdaSULQq4XPQZ97ryVIisU3fUmEOC5pKBgkCRu8Wnlh4PEHJUIYAC
a88YNRGbBN/p33AzBRG1qu0oYPiwsVFfThvLDZZmUVYOZ2W+QGZ7PxR+5wyE0Thw7e9brnjoNfu1
GK0j67iwOgQsn30XxT+91/Cr+bjLGukw4qrMnG3HdeJEHz3HcUEZuVgXOhJYWUmAp0xle/3ZJnr1
RmzrvXMScylcD3TJQApg+zrj6/WghKMKebQqe3q0uH8S7if2niIDYysz1HIyXyp4Fe7TTHGWPytQ
JplWcucFc+zwlCBOgyV8555r4i2SK1X2QaKovLS309e80CrZfbziCvPs6Fplh9MwfOkl1l3VSe9U
MWxbGBsxo+R7T5THbcMcygAES5zNEoYKqx6ZBXclulHSbeJNxJq6HgETuIPXqAk0vpVl30xYXgz/
QRr9MlYhB2T+aYwPDjoporFi0aPgE8ymUG9QWLoVnxqDPSUuvEebdQzzIjjIEUhY9G8KQpFGx5bD
KmYBxv1CU+3U1hdqPf2OXALgAaW+ZRxROeA6BG+ARHfREWipXp+ItXp+4cLTGVT3ojJ3dTSOFnfu
xh1kIE2JIGAqDK18+i2LjLqIhvjB6IOVGbo4BaVAqlRVgFzPVLy/KetsgCh+7g9RxfFzLJgxpy9J
gtvEh0VtwpgK6oI5kmjv/MOuQ7o+fjY5DEx/NgHvfzydp38QGB1/6Uz5BSAMneEcDvLlkrkvsZiX
8LVsfq80N1M/egcB8AgBlHHIZanYECLlaqmSe1Tk96GMJLzaMAnqpPGXKgekQUt2vHkm2iJkJpZw
TmCuqIOj8OuBSn0MiMZLMgcK3PtgvIL8zbTM4XrI5KZBHyirnoalxXUpCQjpGJdpVplRm6Wyje2l
fYLH8J58eKOJLD5hvzBpsDFHJ5XuM9dMuju45ydM+Je2/2CRAuIw6EWdCMhYUEpSQVPJ4ZeJcQhQ
jhIcBXOTUBtBRHVootg1m33Tst32QNvFnwn8P4Tc01tD0qYrrk+kLda/r0O+cwUhtfaSce/pVqz4
WHZrzFn4hQm5EC/uFON/ceMEZ8uYq5db7uSmOGfuRsRbaNfiXBjePWdbH9XLAVLDsRVr6jlKoK4m
FQYQcXcIK9zHcbkEm4XEDCmz0qmjc4ZtGcvOOI55knXybhSEaoMsv91qkAZW91jbYU/LFuC2mdEE
i96+CYJnNKs/ep4UVqca9nnuMiBPtAECLNwLVwV2VvMGHUObjnF800IbJ6bOw2QPv9o7C4K50Wkb
SBkV8I2DM9nGK5BM7XpofHjOS2s1pqzmErNJpNJXL5KYoSeX0jvUm4mzWQYQ5oepKw/3F36F8Ss7
RG8uBhdBKalxs+gH48xFquzdnUIenvwtZ6jmhP9K+zzOjCxJBJffFYe+uI2AgZimEVE+9YvNpz1V
UQXjz75l2BEGvVgLb6MSzruCbHW4taYATRO77f2OjObfWooetn4vgzKfVu0uUxjTqp5mPE9Digct
6n4E3EGMS9POywwjWUsVekb634nwb5lVrmuUkfNNs3AjFUsX9h960ObpX3Qj5n31SyLAD2Ch9Ahf
0e/CYlOCCbKEM7GoLQF1yTFcMtoYqf/GlO9wmny7n6ulFsjV16K6JAr9jlSJbHW/oHEcwjbsm3+O
uZ079npOT7LK4o4gb7iED9185IV2ihi+W2pi6OhEiQA6TQel/Ca8oksTWtbiWpQ+00ojE75TjEHp
VwfeCDEIgtw3wI9JjnaJKsmp0OCrr+zQhmR1ZVJ7WTufL/UhejgeXqgJSWM3IK4ZvkDmu9/BXaIA
yqgLN+HAZi6qM5hWyU6Zadan60lhv30GU7kCikGUntQsCM6ZYlKQbuujX9+LLAiTBWTheeYQFeG3
TZ+eMM51aLY+tlj/gZx2nbW2OAnPcNqpoZc5F0L20EpUEoZgew5ynbOeK7XjlJdILBx7f/I5ylxg
InbARbDhNWvfE6VJwOC2m1YcAkYDucm3lrvxIxBUiFUDLQXvEhGwKv1SwWQ9foBQGErrEgGTdBG2
OLNaXhKTbH+sJ9bZFzhcTrkm3Wp9h1SD+pNJ/r6FS70cPYDXpJA8aTvSrs9I+AupoaXFYJPpuF70
HZBqUb9iC5WiyZBYKID+NAsZWRBWOcJd9ADjElSdGpS0wNHT8LB9b1G1aLQW88utuuZc3hlUOngw
bSVSAmeJ4XZVP/c9PI2wWA0qmMJPxn6DkfEf6a7ADx97X6BdEypWWseWpFNHC2yenRbZMrDlRBVt
ZpL9ttE5zkushq1OnHKHWBV+3R0+uurDrCoeZFOiCzcxeF7NzqkffP4lUS9y9dLrXogkOTakTn2T
p5YgRt/ww91DvbG2IDEgv1g9nzpOnTrd8zDBKqJRc39DYedRQ0Ewk6H8cSiOXASsXFcXQ2ynN205
Slc1H5+KRjFi4SLqpjbCUfSYbfbJm7SQufV0MMHH+L/GZK4B6iJ9nSA36GKZPBYQ5XENCd9ELAO7
B5yRyGYA2Yd7jo+E4wlW7ubDOdaCOE6vS5zxgV9ar34v8PJIWUEHLVeMsFAAcvNP9+5KxaIwic99
cJC2U4zyxoMUuIO6CUxDl5gBSJGgClqzUDl3YxIwm7+UONQdahGgmzqJvh4tGu7NU2KwNheI0rxQ
Hn4e1yAog/6wqp2qT7lLjrRpmZZ8gzBQwpDkVcrcnNHrMfBraaTKxNwZd7saNpyBljviRJMdCeUK
fYxt+XSPPysqZktw5PJigxOSi8+mN0e1SjiRjwxf+xyLtXMwwf0h6RZQkmSGO54WQEMTOybr8H66
pKyQV5wRpTtt1Y6Vd8pXaGGMDuxHeZyusTc2Fy7BBlPncTS6O9ZTQM4AMtE8ZxPHIDNuRh+v2G99
dFmfqcUi3vJSCM+g5yK4tIXhkyON5otxbXp63B73FgCNTR5E/v7ZhoNkpw9XN0bumuL4GhEu/mNG
7D+vhdPDnfHuq7q1mtOa398Q0mC3z8x4hoM+jMGMcUAdQJqUgrb8k0wXTmkkZY37+mo8Pb2qYNcb
kReK9G4/Laj2Jx3KLr7ZJJpHn8xSP1m3IvbSogpS29biYyLqZPg/fUB8tDyEzNdeQhS/joDCwYZh
stobY+zuS2K3GDdXKUP2+lo1ieeQBlG5au5RCkCNMRUEgpxZrcAukti5VNxGdLNBMHAWPaHIPSqk
HMvp4w1O3CSOc6N0SFACfZlMKSyTXVAzGqLVOm3OYPA4ly516QWWkq2fqGX4NfmhaYQ3f5xRevDM
Hio3gOdZy2rt7TJllO+aSmQ7yFnsvQiX4/9aEqKeoDbjsTvJc7SGVam2jqh5wxijiVWwfVhpdMwR
eudFHs/mLN1cuBf/rQF6y8jOOe2B5nUEP8XNPr8v+W2aqXBP+wkTjMQ9LBX4OxBCVYdllJOo7aWQ
xW/WeFE60q6o688CgfEymhoo2FMXATjfU/TPYr4BKtWXXbfCSyq0i582ek4sK+0SuP/bXX6vzn03
/rabzf03nuVaaJngKaXlF2TnoRKeQ5PPUTAXMUtEjrOGNVfQIipRGwfJhQWsGNWZYV+r68Ip033v
Jg0OZYipdWYE3xSJ/a+p/+biDy5JPCOL0TPSfCOcTduOj3+AGP1i7Yhc2+6nEqM6coUl6I1lhrTK
9F7DtkQM6r5DhHvHgphNm57EOJEo2TXZE+8aINcCwAERlh3z0YKBgtL3H8MnIYS4DthAaI8FSYfK
Epr7yprO/LvbpSjxnUHTkHiVbupSEEFNatq4nGBDT/bzhGGKL+UkOU7aY2Uf9iY/7beJ9Zrs+F9Z
XG3J7aYMArX39eNLQ8mbgEkT8N7A/O4HBybGtUH8es1fD4Oq5hY+k7gYZKM6IAmTSYphfV3QLjfR
Ps63ow04oWXgztX+eOGKD376fI8T6qX23cVY7IXwes8+bNnuz9iGEo5/iN3rgTJxo5obg51DE71W
IHstH+d09bqJjcyjP1P+kHUFP4HL+Udkp3REbRFnc62n60oWfsaJI9hHOw92GIwLmUkLrXjbEExE
Fh7gvRdx+8Ok+K7PBk54Lai9wbc5KMhv1UmbLJ1ZpD9kQd3lGuOWhKczpm+e9lX9B9FIoGyHxEZu
18o05wpb/XCMKohDAHDVAIfDDVzOo1gGauuGsKl6UiI2CT6zyNqGCwa8wyDt5dwCT1V6Mdh0skRH
G44Xf5bMqCFHNcHv+H06+xk82/KzwtRTrhTL8nDXtpbnJLB1gLLiHln7vF7fddV1z5FLFMSLS0qU
ZasTJAXoT6d+r3pICWtskmPPLJv8u6c7qaH3f2lTebw3WhGORcniybdPw/uYdPztZq7AtnovlINT
b4TTjia3AL97AFlQ/+PxIAqKGXt9a4JQ4a0w9yo87pmUAs0O8MzGxMjbEuWqmAFjIJFmNh/a0KN6
tKSxYK0iFIkW/nrg/sDYOzKOu+lWP6SGLNl08N3EyqmwoA/cpFDlXBCvHH34Zz4bD6BFchqTD9us
cGKpornzORqQaX/ktfE5CLqWG4lWeIrotBfvsswKr5a3+uL0PRQiYfTzr4pG3UtNlw/hzAhylfDh
9PYJEjb66LazTO/sB43Wc2vWL/gUATt/o9g3wCJOko7CxBwPqa1F0ocLzc8upM0rimaWrKz0cXlI
yU28hdHdnT3N8i5ysB+qgDyKhMvmdOOWAwQMhlU/c9qZeWoL/UmoBFSfxKMygy5xjeT/zGYg4nOF
Z3ebIvo4GKVZHLrbBMfWxuTB1y6R/WwIX7zPP3H4NdyOjibpz+FNnJTCOAMzUiz4kppcS8s++VgK
q3DnMdxzkP5XkafXnXlYCqp/U8TdfcWYDQoAuWy8B4fQ2+BBx1QGDiz5Z6MRQDMN8Nk2jqUe24q6
I9leuJhkwFbLmioITnysUIT2TeEzHOLnbVGOwJEkVNUIQJx0LtcATZVJoyIGLVfjCc2X7wILdqPh
UdLWHN6Krc1BKZkI8QbrE2r4/EWjQXkWy+bnZDQ7oTmq9Rle36A2J+D47y2q6oARjyc/A8xVlFCS
DE146DuXUDr6/EQg1eM+k5TRFSO5alQWvCdQKaDla/Zk6ZBCVAOypqliBUmki8Bm2V4lQ/wx9q5A
xrCDo//wbvtkjQnuL91egMXZs/Na0ZmYY6bUaCGLiq45ym0cg5oeyhD25Wk9mzjphnrI1UkCbHX9
gtl2/cXl+MWFY+0jcyZqdl3V0WaJeuaag2HmkMk+y36vebSiVtrrzkMJYd/+0h4FI+91I/4HRp3y
8pTAEcxFAw+ebIBzNGAZVL570lKMtOMQnRTYGFFWb2eu9CEeJg+DXhasY06uE8yrMbn8uAxuVPHs
J1rn2aGL/07GKWTQ+mUZRlxMN4HuSzKynCBBBa0o0FeCo1BJdamq3J55D/S1nkOQ/52Mat13Jwam
qrXP//V6OdIbO9woT49Vm4KQ2bdwBOBB1UyN7Lhz4PA9o4RD3qkum9zsUdtxX9lMSp3lWqKwIFxb
hItzUiqYNfWe+0iXlrgxeBv1ahXhhYl66XiOuYHc/Ttm/Gy0wBZ5iGwbjYVzFHolfaJcvTVBo/VA
UWot3RetsE1Siu2hYVmlJCsg2nZxkCD/nyA5L8KOJar67GsJRYIRryppHWM0YLXloOcr2yUgNpFV
uYBlLjrVoYzSMrnHvv2Y7o1fGO6TtmFPeTbdfkQzZ9sx8DHKakrkBHH9AgTN3tIX9/Ueqw6GZqDV
prNd5uT05PSJ9qCt8rxPsWny05eo4rv4nhUQwrCBtL4LAx57YjqwLNFmHkD/Zg3sXCppJmMObpvA
C5GJGVq+QAl5YWMkP86gU2fmP/4oYwtEzwAydzJra4pVoVSa7CBy5F4ZCD+ZBkKQzL/FSO5b4mkA
6Edl0/9rdADKkDOEmazAUJYABRDLtBXxpQv+je9vIdmU0LuhPBrLHoxlVqzWJ9N6EM/+m+4lVZJ2
BQZBEev94+8VrCdqD5Y79d5nsJ0skD1a8+X3AnWLv7VBbAicqvdKyxAKqRKRrGgWD6plC9C4ENQG
hoIPJVPhofOZQLnP1vhal63Z/tSjNiYd5N+FwzsdwlMMWu4yDzM/dz3JNGqEXZkt1hBb4XtE6Kh8
1ViQuu3IEv50kX0sg2J1+WIeDdPIqQ7lqDOyzETEk3Jl+WWdyh2T4U6TdBA/Yrd5rpd9fVBNrdlt
zrlcGVZXMoKylzJRp6PP1T9I+KIq7mtA1WxxBBxLovodI1Qlf2yG47AaHbYieNHY2/VwpMfR8oWJ
KUG/gI0oYng7P8cio+f+0DyeFTYMQZMJkAR2zsFw6ZoCng9g8Tz90fZM7TtO8I/N0LFVVcl9yrKH
1HzocoIYYqWqjAWWNNyDUD+E60ClsRhp0fhF9tyU6lLuY3H5oU1BjDXadfJk2uaFBoBIbhsTOnV8
MbikCG1x7WGKzKWJ+HWPiVYLqBVPLKA4+3QI7Za8TUaqpbV9YtLslq+XyiUlcchD37cexIy2CZu3
fF0eelF7QsGnn5XuQ/YRhilxEyip2rqRhgdiTJx1XJ9UU1SF3gvyQX/AVukiaC7621Q2LCR8xLxp
aRGZ4UlgkuQmCH7rgh4v03Q6sFdxlaM5GoEvlLCH0vS8RGi9n917Gi3h11iNO5H7pxyiCOX18y9S
92NVMjcW1yHWU4MfrvnBIrlNvlBzJMexPOAMtUD8ChVyNswiCw9lm+kH/swpkrsMp9S2hVrHibSV
QGL+RNjg/HVF+oE95SwrVvSuUL/6BBsWDmSQZL4UI7dOMq/4SIC7KMZDBbbnZ60NDC7Y7+qDGl/q
L25mFV8e0nlAh0XrhdPocU20nKqVYI7os0S+hC6FK5r4hGBRM3AJwMSNfVZ1G52g19E0EV04QwI9
SI/6S17kdG8HDgFJ1OHyb3u3yTL+sK0b/GPLY4dCf7VKLDcH6herzpoX3oupJxowBLCprUKBrLJO
oJOP5mKYkWr3HiMqc8UI0vXDE7O9Xoe/9GviS1GLAszcdXwkFMQI+sy4ezzoTxbRt//JG5v5hQ+e
uDqI4CNohJ/vJzfkjcNS9/gdt3f97J/hCciUpXjYjuhYN8gPVzNwsI0ZsP+aEC8U1ByMeC5Tx16K
qqb38WRLOoEXKOHxm8i+H2qP4breov4UBbdP7osCr4zCRgfLcO7whn31K+ifN0W6LqQuO7Rd5u3F
EemnFhbpMfS3wQzYRCuIwHMsxnEwCAYgpLq3QCKyglEuK74qWaGO5iGcHAdDCE513usMf/nmOKeH
7nDrUn0Dw2B+/IJ+qkeJNvSR9Cfi+m2o919CT6vBKgeVF02BdwYr6SbpXTW1QZjNYYImpQaMYaph
Ofktgql6F0XHEaSw4Aq2OFPpajrOLuDetWmpFYjNznFVosLBsUVtKmg/BkGoXwxxs8nifgLkYYl1
JsdnJ7psx2/4POLxF/TWdCrt5hvBC99QCtdXpmU73O/zuS4cMMcQy7NS1AjwdRsH3sHFOrVehYxu
Fi/rjD7liw5zTzZyyOOyCAaNaOqALJJFcTwSxiPjHVF35b3dEwpp2anibANQjwbqFWappNtcdv2Y
aA62nlyDxFS6SaaeH3318FeXYkRBIvbb/SKPPd4+IUwHjDCSw7Apum6XLg76wS15WRIxYRyn9/9k
ndlcxejZLuK6Pa26d2KVjD2A8p4pwYmBc16AGNmyU7Bohj2xZqqeJRxQsGIw37hp0+EuQKvEbW8Y
KYSg6vpfjsGN3k7bX+hukSKAa1nmnpb6xnjNwCfY8IfhFBMRL753HsKL8xFLWKX0wuBH0UNIBqi6
18xETq2w3Ss8a0yO1j6JOeIQCZB4byIFo3js5rozKnzeOaBtSUiahbiOFY2n+fJo7W0eu4dXPC+W
iysXOUHO1FODNH4wXAV6PXW8cIz6zYsAQwetEPfeJ2iSvoqt6FzBLXw4xYPnozjGvkBZ3ss2KNz6
hSXlEhbd9ER+e71xbMa1DOn8NhCBtVRuVoX7/0f7JzWwEFgwYKEaLVtv/isYCg4bHRFqRzZsEQvL
3M+6deKN7iaqS1uwbBrssOTuLKtlDN1QP++OW3xsni1+ix1YSos8pfsd8o8uNvVyRWJfB5nWMZyZ
yC/AQsu8aYtYASEYeR/WohxBy0rKIfHSf/prAVFVPi7lMYIN3Ldpg6lgFQTkf+Cdd9EDDnUt+7Yd
NMQnxWM1YepnkVPMOZGVX+WMEgJ5x+P2u2rtp/bc5cJQ5P+QTauecNfJtINP+29kwyqJ4JLED4GI
WypxqydvTyKJJ0FWAriD/qC+UosQF8EtdOvSJJmAe5VLs5OIKTNUlYxuwrmwa1+Wc9CtO65ZtIzP
4W1Nle9mxcrTDUboxKqusJiHB/JDduHGqQNTeUqCwm2UnkF3xmjV7zeDWo6moYTaaH2N0BHIbwWZ
cC0FJWXaQTJ2w9BTOGcpF+GJ3UcWngNP67g0MK6JyvPtXxO6q3Ly1jQa+rWeaAOsd2G3QcfhXZtt
GIva05pHUJr//cLMxZWAlPmkZsf0AJ/Lbcn3TJZzLk5uTFzC2iA/0HQpjXP279LYlsFUnx4yPnnu
Ifc6cWYDXrJVHwSN9VtxRmMrDacnzR1E1NL+T0ZsDZ9ezZviiPrmVJlcuqNwxjNXyfQB2jeyoyoH
a3+g3ICSLd+hzLXLH1VxH9Wgp1b7w9Gpk2spX/abysQgMRJG8YqEMUnAzklUwjLmheE3t8PHsWie
E/v0iEcgLLXFgKav+hw8vtyNhxAh7f/JKi+6eAb2kSEYDkEQoe1l12Heu/ICMCGh1796HND7Mt4L
MGtN6+4iZnAbOJmB7e/aEA5UXfHbAtRIjgmB4yPEuLXNzp2eL51FYOWPHEUeMGt9dY2bYT7+7emF
ToXP79u8YaoiHTorEpzj8oOZPJjWtoAxo90M3+Jj6L3E/UlCN1fJ2yTHeZ6RzoJVXzh/pnEhcYOI
BI2dcSFfisbC6eWcecYpLWcqj2eSggQHrEhIB0CY1dUORBM+k4kuA0FD8eptsoLsnt+VDj0GL6Ex
qWiJLZFR+jm26F0ZDVW01wqwlP4n0mDx45Sdm5SCm8JDrmC8yGWkxtm2Vq8m/8fVRDLMQdxE3UBv
YCPdYlQo+cAu+bdpzY/hTa6gB3MS03dJu5evB411iIKbILjTTtUlXrOWoTcXU01sjv5FeAE6496+
VCDARaZsyC4/leO087lglxDBzkiZsFBXlEI+7jgl+WV+hdFxxTT8vcLwK8OTdcZpIihAkp7IbkBX
M8geew2QMvbOyAGNNfozSlrIRiN2Sz1imIprSw7e8y9yxRJNkSBYHXlzGVuOq/cK6v6loqG79iCM
n+zruyE/wnW+lCk5wyFMLGygKSK80Adz+sEf+lCc8kaGJ6HZ8zbm7m+T6sgiTIsIH9B5B+1Eihai
jK/zFfx3eewGRb+Z8EEczuplemV5RbzueO/7+H5LWMObHsRGrh1P7ibeBfgq0YHBO4hhDO1DMC8A
J3Xai5AbNXxnvhnHhgPtCcweD3GEayYeRFJQWTktxJ0dzJcxpExOrftvQIeiECufydrMyELEv0nz
RT02+tw60omVnGN2xwydYLyjKFPPdsmaICBuxw4JPcRG9Z3Lze/U5nOIO7yfaPJy7d6Ca5TyyS04
LUlTZnzjN+ALt6NbUeUxeGwzvJTpbtFYk0WUN26iXmQ2O4Nd/xHZ5vzaYClMzczJg0p1BV9THh5q
TuQlsR+KgMYOkdWX3hUdgRFaBY3Ke8FjxisSpw42SaWwY24qdlnHvd9YUMiOppFy/SUmNwJz9MMW
Nc36LigbJewBmYSOPntLXX3GweKMq3MDxCJHCzqvTf5p4nMTlFG3xrd+WwojWgr6ned1zFnso5oT
EDiClJOAYfMdgzLiujXvS0luGd1PIAPqb/7h3qtoJcfD6GEv5y+h+B4EiFWPJmWHSmRC9Aj3XLbq
VowChvyQ/OtIjuim+y4xWfe6jc+agl5bCFDbA+LaoL8VVf3bsxsIz+UlBIZH6rFySmvNicMQu82Q
xSgSyh5bQlp1UHqO1eSuloIj1RjvmrzquBA+Ga51+FXK+O2ybzQnn65PLq9tXeQmzV7BNaLXSFI7
lk9RU/okj7PGD6ai6/Fwmpnxb2O5ma6frwB09vNmfWi29pBSCKIDuNO/XqfQQMSwETffI71ZybtY
9cngbg1TcbsBqWezU8c3VYotDT/LPFiYctr6ZnYflpH3IAP7vQwsf7o38q5dwMqXhFd5l8KonC7d
al99EwC6tO4YGB2TSmkF06gike63Kwh/z+Xb9nEOxml7lN8Y7roxqwlakr929gxWmthjwgylecUK
m0unlo+AMfHdPSX+f7cA4SmO6kO0r2gah68ltD8GQDixsyGxOzZCOuZ/rh2S06IIyVx8tEenR+Xh
4iWO6Dq+cC9pwXMcRkn8K9uDVi87bQg+4v4vmkxVbQnnMqvzUDTa0K7fZYmeOlzPH1EwJiR1Jdal
4uVFtF2uE1zDwhp1+bolgO2LU8iiT79n5EAUJeGs/hH4MRw7/TzsRuv2dmFeu+VPIJQc+vtuUNMg
0UClpjsFT0Lvf2c0Sfin2vOeF2zyU2rDBD9UfNblH9kUzb/rYeKHYJMe6S3W2rpSrZp4b65TgSp+
4fvzE2WAQCN0VSWEMUDccm2aWA3RJwqeUnE7x09OrN12iUFHEQDkijYIKnHRtMHd36URrWRVby9j
izyhWQEUmlzeK1RUBX7wKaNvWiTCLe5nCoofLyUqD5i+za3WrTcWKa0j2VP07RUVJiN9Syvvi5pR
ne6szvQx6KArVVRmxj9pmYH1+q5e8wrAycRDDQjREBqDXc5lrVf+3uYkbVVbLEPqMFqKGQD9cJHI
bxXA08eCTDB80yOiCKAvTYtvPIMHu3Yr64tRro2ul4o0j0yb9x84nBcwRrX+C40KOHzaFE5wqV3Q
ozDUW88iWXsVJhpPqEAsE8Q+gEJTo6+u1AGyGqvkYtnPhN+H493Xqt0+JZKFxSnPNin7XOJglfd6
mPdKEf2lU/QSv7jBe2fCXdCPNYEoDqLvc2r7NjaQBoexB4PYJp0pB2my3faHJZLBo7AqZgOyvf9e
RHOukBVipekOdZVBTFeFQk/3O3eCT8v1ETHD7aFZT5pgrj5VYvDXylY/20s1s3Oq+Am3RJTekbGw
Dzuik6UdSoouIqDQRn6T/1YfXBL3U616eVRQmJvcsvmPMaF7qaWxld0vS0fxsZZzHhL38rjRNK0P
YWUpY58qqP18dKjTM618E8QNVOYp8ZHNvZJNLAnmtfvA0/6gBdseNa7r/yXqqeIuW95jPic8A6fM
V1UForCxiMeIlAX7kimICgebFIzyX7JfqcCwDj57ORwS2/nIKtkUiOTkT+p7S+NHeSQ4vN4qk/k7
UBQ+BF95Qou5qOx7Etzmhd34a9gj+yr9PqKswwbSqhenL1tS2orkJ8j+Mj6GWWrcEAh3kfnidDOx
aWERuWZdxPXYbHee5SN2K51cmyKnozuNfarWJuRIuLJheafrZMGfWdUstdreyKa7RjauwYl7RZSU
Gd7mwLoDwleLj6mpz2DRxw7nt8Ne7kK/QtTBHlbfNYG1rQgKbMajN6QH5MMe11sXrB634CsrmuST
vFYXeOxkH0zQ/g1aB4//8LTKvSAMs1Adr3bMn9Itu3pDeq01UtO8/PCWvAEfOEy+yeBbcOBzZg/p
gfrmaNQSX+E8rV4Q0qMWEZJJRzKDi/EZ/2NkHwIqHU6oeEalRzMY9tOA1ynDhc6f2UyWY9l/pDeD
cMLR6RikYXUy9zjkljdDGVAH/TlRLm7c4xLBKT1FZXohaDqxProFxINlcYkBfzkFA20pYbKP3DmX
GLUr+19WQl7y6hyun54vvIOvz4OlXoR5zWqmXadJydjM/FJWQrJrPVwc+b2LPDvBC2CotrfS6peJ
YdkwXFMtyjMEo+ocjTEk+eyTnClaPy03HZpwRYqMGk4NWlmmWhj5MbF9pX0XL0A1JWwmWIrRK/sF
OMjYrtPHhjE0VRzznJ3WGpmOsz79Y1/zUZGIQ0Wh9WVSebmUHilE9AayfPr6N4XR9/d4tKKH5UI4
UejloHwBYWvt/Rsustv2SayEWWBp4lFH2TVEGajWGC+tFYMLfslXn0R4hNukXbsn44zmuJGxM2JN
Uf15HdZsBW1tysU6PGg+IaF4buIqAPnzrTeAI0tLoIGdXI8/UMz+oQPV/4wo+JdMYvEVo1kZrHO0
tYAGvds9YNnfSyxu6jGXKotLJoATuwP3c0BnVOKq2FW5RNz1Z7qto0QerGE1KaU9icEiICT+FDo6
6w65qB8XJ3zEkX8b4SaWqC5AeBcdu4s68G+s4eole0eB5KMQj2YjvOAX5FF6DMbE1XwOrir8EMDK
cjGZgX5OkxFult2ck56+jOOqKds45PuVg4CSOJVrdKBbOVWIt9bSL1jauIEUaoIa4lx9fAR0inpc
dztuZe+ODjk76EKn2CGmeUX7+M4Y9kuWnvKYtBEQMLLfBYjUPu+WBQ3eLr8sh0sUfL3SUBK1kSjm
NsgB4gAmHRr8mTLbTGmLmE47unvaxtNdMMJ9Y7OONf3g7eg0e0e1Llge4BpWO83yMs0Rgtt5MxvT
kJVOHDtkGfZwstZXNy1j8r/AjCj2Z4SQ43J1p2rOkbhP62ASThUaE0EPkJy0LksA+huOcIMyduMQ
1pPhxKJS031m8tqQyNX/qFWW++5gckDhLROtowGJKVbQL7r/W36kieZo8/0Zg77sqAUY+iYOGunT
6tUAhblhCXYH4rKMOhqoX17tjPkLx47wDvVB5kRX2ScoFutRbQqkweWtrWS/TWpBD9FFbARpFDRd
bNUD2rOFZ5D0h3peQDhBoiDStso4yUTbC+VVdBW5iarZk/iD4bOyfY0ptTlgdAA0rDuOjsA3dwzL
06MYbdJ6VMQCr6ODpliZNOb5OAUb3kHnF+E2kmcTKGm1F+/mTxnOm0wKA0eYaYCdfgzDGp9iMGOa
4FVI3IH7h16ZoRVxP+AHz490U8+pVU8D1NNxmeHu0wSpkOhYKae+w/0TD5vmlcZs/QxqZAoGRgpz
Y8A4S8m8fzgD6SycwGdgyRBaLu0fiqu9CEYE63ORURTt8/+GN7KXHFrWLFiTu5bbeoNu8xPjDLww
ED6qHBCQkLbwYRZxUMlPGyvXm6Bbs8Tp/UQi+rHnywTGc9DPwNW0t8ai8jisDJa/InkN0juvE6Yr
kBvr/gqwmpP9p14P9vQgPpgjapdD6DL3tnnU7M54k83cw9dEU72vs4/3/Nk2s5Wq/l4yvmkHNGCd
5udPv9UJVG5DqdfqvLxZsmyDWGjBY3+nqjYwInahchrEIfgu8WN07+bHqTobAYNpj1JhrGWimOlb
gQ2IysmAjVfPxEqNZ9dFgIOFjTI9nAdOalYdrjk9htBYmeiJbGvB8rCBJ+cPhgoky8PxF67RMhEy
qgj2Nz3IMJMLKac0vHzt/PPc21BdQBb0jROH6tD+9PipbYeRStcvpV2KYW4apEqUMYTKmuq0pKgo
EAhgXK8KAryJew38UFFJBtpVeLfqmb0c+wFi54mZ0oGAo9/FarFB7qc2v8r8j6DPRHcciZBZF3vo
r+B/MGceZ08H7qYpTP0qnbCKcwQHYpDtRh274kTCQRMjnuD9U/cp7fk9gguSFARaL0uc/O5iYrXy
vkAivaFgIBAN9K+Q825zupKp0IuPCBalQfQtPfrWyUDdB3ruA3lujHAF2nYNavIEp1cJIAstJ4o0
NNWvX9c0VJvq//3/O9A+7o9VNZOBp/M5cWm+3miQvk3ufblC6yG6epD6DAr41a88XxXiUz+CTY3f
xPUSPe2vQAjfe8S+vpZmpjR79xzJALxkW+NUeeHr0LvG+O5iddGlMmvEOqhgOgmSs0xfy79f6laQ
rGU3V8z1J3WQxFXHLwaZAV3qf2Y8pC4Tt8YQeBXJmQNaQJL4/tX7ESSFIpqNnHkfme4P7tCabqTB
hh4ra+BHGxlvdTzfpL+6P2OAY15W47V/IKZ+NPZTlh7FuGVuB+ynqb+NAqovhndHJDvbWSAn1+gk
NsVplBspENQwqONOcOIA+MmI4aU3eiDgK412j6myHE8c0V4hGI4cz0lV3OQ0/RtacqmuatrJCBLS
lHXaJBeJ5wq72pVhalcpV0iTgaFztHYdxJczAIk2g6Png8sr/2FA4OWOrIqfbeJ3YV1rehJUaSW1
lge5up0Z5VdH/DDEBXf21SMB/cQSUupuQsLVSnXo4i5jfTskIARunL5YT3vxsHT7qXHPS2SIppAz
c1YciwbtgRjMlEggdGZywqrSi5WOj3onWJUyVpF1EcLRnfXCG4DVBhsUoe4qRFW2INJxK9Idc35+
0qcOyXFBN+Ri3BMmsAeBRkRixspvStNwV5w0i/BsmqQpNu0GW04Y7w92KuGM7aKli21ZOfi7XApF
7x/Bs3AdhaOGruKtVBK65LPf3j7r7hpbQuEmcqyXB6bWNhYWoRMrasE4LhGqYYuo+Jlb7FYXC47g
Btp28m2TXK9aKyCKFtjO51XlsWlZOfQnwpL3OptWkxSkfC/OBD/izTPL53lnkIGzD3riNYoSc+r9
V2MHDXxDQz717JAYEU47/whyFICc0wAG5qVOwJcduDNU4Y+UI9EwqBvLBxofMT0gUPIAD0YKlwz6
6lT4coGtV/k8rjGAz0vWfDtMI6oGD11fTX7vtxGri6yqLPkmKJ/mDLB/E8YN1kqsybS3yzyQofXW
NJrapqUdxfiOelQSlrPrhNG5xikAlSNlpMV3aoqhW1/ZdbGHsFpEmH55Qo25NI+zkuy7ztndcHCW
IaXyvI7KM+fIz0z1vRMuxUwVJyxSXCOBQV8eSBqSbZjYtL3IG5/KfSara19ZyGexobTkHg0EENeN
msuSFnzlJA9WCmJkXptyMxRJjRWBa7YpmKqVdpfZySRYbN2bRmIKu77o5FHdPfKBLOGt8G2QxSlZ
S2AIJ2pSWpVoQPn5rn8s6tR6GIWB1FepruvxDHFPrYCGWxN2R0rbIHeZLOX17AgZFuMNLRjGKACw
uWXAfI4EhDC17uxn4Bp+MfaxHw0A5t1+ecSGreUbEPA3M1C2Eh69VQq46tJvqNr9THTHl5UAYH3c
bkmOops3LdySzi7+ygQ1+9HoQRb3+bJg8P26FWFv7FwjBJvEdf+tZGd0mmUVu7SJ3ze9Pw33jP5L
1ibSCnOnHxDgHHE2vgPEZSdFBKTubKnBB4Fgie/1BM0ZOEFgeHtNd/kAOUJuN4HuWkXCFo66ApPf
3l2UY0W8i1aTmgFjusl/evAwcFzlojuCZKqq5kyy7lolblxrPbGY1Ypb5By6rmyVq41oihqYYQOr
OZ1hel6BZ3pxVX9V0bIPrdkHNHPhtL4IFxd7ajBNS8hp7B5AKVzRTBRkfo00GPzi8ck6H0jkOXgb
1Xto+RzHiyEmoqS7QTzIp7sUPA1p+ru7tUI+qm+U1S+TKiYr/w5/xd4MgESk+3JlFJHtyzb/TbF6
uuUYMGEJFvA5wAcuhdvgUxqhOeZJgmBgBGMXBmDN5kOplzch4wAXcLbEHWXNsBAR+yJl8mNgbfD6
UgXtsYgYEAx0cf+PWl8VMiDcAZZi2rcV9/ra4mMXm05oYfaBrSA48Aq9jcvlc04Qdha9ziBf2YgX
QS7GMuKkpzrxPKIZfrXAcDeWKtqhAUrl6bTsxnhjKLEmbeGqGGqrg7P+4kVdVwDI4HwJutHH9VXk
hwPBft0AQ5cFmaJWiUuX+bwdAtlnm5qjd2Ie+q8OTti6NGFOHo8eB3CmNCJlJB2S7F1vn6MnCgv0
4uukwQaHSg8H49BjcuFnR7Ma8iS1UQoJ3uScEQ9P98smLrNPooaNmtPqFBiE9kk9kIBDvzDi92vf
jim9zd/T3G3MaXyt/QHRrOakiQcqUi4IoXqyW/y2bPavuxJAVxU4QuoQl/tWjYlv/mSkcmbAeIQe
QhNdBWcJu1cD1GyXPblSmLo2ndEBQwpEkfofpDjr+SrlR3YCV6HQvzYVQu+7yMgjpw+gTSHCEnW9
2yPnOplBzgLadCIxAqpd3WFLm+e7yvaCGkiaIctBSfw3w9d0800Se+zqqN+xR2h3lzMnDPUjYgc2
0AvXWTcLs23QFx4gLqb3CHeDlaXlC9UF1K38MM2X9vZ4v0+AaJdotq+RviEANZQQOhmNfp6u+YzH
M9xwp+XdiR+pxBno8OyXJ8psY5mT+wiCZX8FLGVAC0p4MgA0kpoO4JBz+qvShgE+GoAPWNMtI4v3
YTUp4+q6oVEsDONw+ArljJIY1zawm1Rc9Xe7LcenZyOoemrNWwRZKR1XBJWVdCrcKiMthMxe7voV
5FFayK/ig1xTTNe2Wp5YNJBTLk05x4oFdgKT6nKnHJoDZ9hzwHdxcxtvH9La+vtTZnwa4VioMC06
tLY1fOpSziIBKiFe97s230iS07WHo8JjEx9PFYkDFChbkFjdKpZyEzWYBO5bgvcKPbUdRlQL02dp
IyNi0FXIyeWcma8MEawK9NzyGiJQow6hMwoMYWmXqkOWJMAlYGg5VWVRV3bzq6mAL1/l8P8Ycqdj
SnaLt1+Wxhz3QVO0OJhDqXqvCLnulJ9zXA3+Fv2EKh2UdbGhlZJUbN/zhRp4MRU1mFmPzqQfpyEg
YxQEERAW65GhhT4OmbyrWRKtrdLtNKWt5NevR2Ks/Z0pT75x3iODM6mZhkjf9GJnWr5FYEVNORR4
rproyGYqSzAG9QK2e437HPKgfStUIU2tDxR5xB9gVqW8rPhoWnEAztIi9t5X3IEBGzIuqCVVbZZq
QnMeDKTEgv2CN3PoZWNhqZOBFTCxkCFYMw489Dib/fNMwS/7TA/dnHGbVg4BjUy81a85pC24smak
pVjMjuaS4DxE32JJXYO03rCPrJIYxotdJVfQrzAMkcpuPTccOiT4Us8dwmZ44/FS0/Yr1TU4W0Ne
eAnqUqHwy0qn3zwsiE16S4SdAvAB1EEoFHXu2SnAhdurtf0l9ZPW4vc6mJWBmSQ+vn3hl9J3h2Ga
N4GLT9j3NBae/lkYhX16TYxQ+lF1u9Y7EZ0Hy0ifxR3qXJDNUidgU3HkNltvAof3R7qldXRMsXm+
CxRGtI0db4wTKMwsRGYiFi4zgVzZogE0urEORCamnuLtfAzQoGs1t/SjKzYg0m3+jzZauJt+24jH
UR3AQy5gqjlOrtZoNaeFppHPRfeTFQ2qW8I3EWni2f7W9lTi5ecjuhs0EjUUSiyX6SM61UK299vd
5BrBr38Ge27N++uw122i0qcf1p2ooW4ziOgTEKIJP+VclhoPwxPOdPuHDZnI5VroDn+CxjSQrQJn
Mim0cuPNoNNajCPSjH+5gx4dTL4eT0dETQgtm8ONcoSVijv2mr+w97fePjPKp4XREIWH+6/Veudd
F/145M7ObLnSdS53IDAGS4jl4gXbzhkM4tDK8DVb5aRzYs/x4puvuw+nU1YIZY3bQ9+mhswozotZ
JghXqCOoEais7ju7p6utyl7rOotIkMkrxl5SdOozqJyHPFQfx2O2cqXkCa25HWI3xXjOLbiN+DRI
YAF65bVBPHDBE3QqcetV5rb8EBhy4Jtmhs+wqESc00HRwEqMtfA+nr/p9pB0A5X+J7zA4X+j6Hl4
zmSwK2tvYxuhYDIRJsmobcKuAdgr3h5ZtaQUzlsU8E7ZdYFQJNF1xGmCPOYJ0NvBZkY0Q9KFrIKb
Eig6jz/tjk74gh0vZR6+8V+xWxM3J7w/AvURzOHjUiSNEfrRH/3hDAE9GUA1PnzmpcKcnJsgCZ2l
JnFk+4cplXVxfYJNX+WqLQ4YueCQQx5b62csTd1fTMo0giMaUXl4h6lchNKoH0N5fq6/5TNJesju
ddLE74yT88yTvOp7QBH2CLD1JLhrlWmDzGihaKrZe2Twa/X+jR4jicbZyBeLfg9oY46fudSJ/5+/
Cscun7bqX0J56eDH8v12Xo47cJQnaP2v8XO+jmcFpaSSaCItxNjzGJwyr8ANy1jpvyz1rngI3CF2
7bhvzqkJ/0opJq30kNDD3KGN41vbxgoQLxaxJ1lLAN8Tin1A+XkQZN6ELatFcRaqPVELZ9WmlCPZ
4l+L5fTazUh5oEkLJmL/HfveSW4NaURA99xpU/9efTfjmphPE3RlWwPu3unbZtezEdXzkf0+nhfr
0sqXKUlLyWmwnV+ONkurd7PnTUxnbjqbs7EoRa8IxQgrZCZy0sP1GZq0htZZBZjNXaPkTllU7ETA
3oOSHKHC1vJa6Vg+B5JDS+s2eoJYD7ncQKIuQM5iAsyput0A84/s/CZba3/vFi2XiDXfi70wroYb
8r6NALSSvm8mO0RS0oWIlLzQwQILOIn/3uqb8Oc1dDBZoMCNd3cwEZUC8DpdbIPelD8CU1eNk4wk
IRo2n6JlWX314JJ/+sXZL9ZDsMmmV9qt6iZaWS6e9jg6kVB9Q/WHpgBvrYvFPZR5VGYfP+7FFmxo
Gkx+Y2MO2W6EwI7oG7W2xGtNnh4GrIOhe4mtb5VXyvjLtRIcB/r5PMoGPGYM4DyqX7PFlJdzvSQr
2EE6NpqUL9d8vmhD1W+iaPNDgC6IQQHVN0zKqDHgbYPLDuHBASuRNpO3T4/kxTlVXzDtu8Jn865N
1lTzyqE2vxADPoDFdiEDdHLw6ozOL5eAbB+UL51t4Ls/pPLvdPJ5PaXtbd7FmjrS7FsiLH9Eaqkd
opJq4PHYXv5q3Z7j6U9q9TxF+QkFDO4dgRzJL4HmijZOWi8r2Ff0yIyFEYBDUSY13Eh2EgqF9NQE
Alyl5M9Fi15tDT5DixEhdInfLFZLVFJOb3wmPWpMPYgkjKnGbozaBH23tKD4kpHv5Y/jqcyiQmVl
RqlWFdskfFi4HQMTk11ITLLj0XjdCgLQyAmXMGnazGUQrMGQwvEY4cZ9ZhjgCwk/q2FnAhBWz7p1
NUduDSxE01C651Ntbr3doiRFtYsnkWAj1HSbEqg3XdpHpab5t5u9vQ0bLobRLm6YDkmDnXqeAsoc
siYBAmsM4YeZpG5Bvv6zCvuL04JGNJYaY52b0wE+1n4ZuvsLyZ+f5HoA8o74yfFggaadnKrL6Ee5
quV9y8h4eIfR8qpLjbN9OHtKtXEcwrTbHIXC49KvASd6LoI5g7qSrHWnYgo3lHLm+QL6UeyBrtAl
iYzmb4QaE0Gh/NU4TVA4NEQQmuKVNTM+9AaKvEUXzr8CVHx5gli++DFGhcKgcckyCHIzzzlHu0J5
0N8NeS9XMBHCTBViS0xlItGHS/XVzRxLRWuNE2CuZL7S/T7G7kA27tDijcaIiownh+w0+sqOv616
G7eGUgVljHH2oRUPAyivVpt8zyRoIsW6Q0NzTd4O98ViBARYPYmp12Gg6qPqu9/PmbSZlnohlQi5
ILJpM6c/JOzIYg/TjEV4AjHe7WF51kCQgSUVj7ZWGm+v7u4W5arXUJxuoh6SFzDD4qI1YT6XluCg
EpbBB+WeHTMoer3nmfuShHJexa4qR/DpcPS8wLf0mndYhN9XZCzS7ixkOrv0X93aBCc3OHD7sZM9
sltOpXEa0RzA+7UoIEUPH96pLEUro/JODrDFK918akVIT71/9EyJWY2yImRZYFMUk3j3xycbxtMn
IchvxBBnvQoK6ROpJzNBSELLKAV05u1k/AMd9l0iBvf6t+bkzdmNeBFIxtB60Jjnb/CeMXKBCBDc
cbwdGNc9xfBN3/GAbv87TymzVGQhi5j+F3qmm8STUs/IaIeMlO7qHvQpbCCfEz0kCwAo9yDOsFvt
yDfF4GxQk76bBtgkU/KOeYXCHpN++k18AUD5KyZSPHqGk/JEukiSBLDkw7dlaSeIL2JqvPhWg5zB
bq3Z+gZ97xmeL6w6eBKw4LibylFli0PFXIVPvo+UdYv6Ee16JcoMUwV6TT5Dg+OAHy4zjEJClojw
5mOANUJzoRam9520yHes+paE94F0yGhyhakQQCr0WjZjpg70v+FKDRW9UrTTeSbMfbyS/MKCOsuH
Xc2ZOW+Pjs4YlBvxn0LfS6QRniQ50MZ43rK7vzR2O6bplO8WYL8l30ZLZ8etubm2OS7aaJ0cYGem
PNQDfE1akmB8X9qZUwphinWrQ6fbR/Ibm6BtXuZkkKzi7kppkXqG3E2qh/ANjVTWLMPWrtQ9DtJx
rgGzVLtkdSzVrTxz9UggEbAAxzHZFyvv34pgoeUpybPCgH5w8n/nf/r6ZzwXP2Nu/vKencdOwRtb
t3P3dZrEMKTnuiLMl36z/Mx/SkuruH3pWq6izqc8ELCY+4h0DVuqkz1bEw53/UJ8bZGZIKh0AASA
qqZV8CfN0vCpMH6jbqquOja5pmDCZ6ki/unmibQl9BGEH3JRI4pdOowTOZSWhFa2E+nn8/WPgoYl
PxI1JWHvap/QPfKAed7aDOmp4MQLhj1sAwAHoQeYBSQEHnNdoNwdEy8jxtbQuPSM5Njofa2+fDA9
HN+/bRzLezXi511EYsKzsIG/QVg9sc2GfeZ20+TpOz487m2wRf9Adlc64tQrBt1zxJG0khtLmYqh
kEWSb0ow70Ne6I5n/yGtisiTyfC5BJGl4fcrpY1bc5StFq6NwvI7i53uzG0rrf0z7gDDYGBXAZBj
ikZCMjcnyZjTUnZs0MCOmwRyCiPp9fBzo25nDfcAG8m3YN/eFiYx/L7iqfPPK7uO+it3kZMOpUhn
dD5G85il8t/ubhIzdayxkOL9dpLZetagg/wP1lD77/vYbIGycKKetKcYNlNKHCMFiT/vmshIE0pJ
KRynhFhbXaWLgS8OIrPGerdqoehxGR4v6ZPnayYNpH9c9l/E7mVvAdSRA/TI5Gs5UYNtUclZt1+F
/h5dLDlLE4P2S5D55+8AQp1NAcr6uuTA8ZAQS/CyaXe/lLcpccxFjzLEQTHkaGV8y8EkeA6215PQ
vHUQvkIf/FO/P2idzHN7YvzSHZ5OdVD7Mdpe5kYOhw7F/vltVwPUjExr3Wy4k9dQ72rmkdFz3ti0
GSXPFtcOMNxuosscrbUdTHVD7x2QuTRqM/24+8oA/b2/W93ierhAOVjMzL10wXcrA79FE8cz4rBk
VOCGHCrBW770Mn+DbsEyWvIIKRPPsUaM7YtTGalqAGMKfTqalgGq21XBgLS3WmVgHabXKffdkdxS
CXN49xeCupZmkv+WbUlg8yk+sXIivb61OyQI0eTU7WHzHFPzzw8wAqm7n9gKs8/M1ZNFNdK3dmGv
mJ1F88yRclqNpDy8xxNoa1tf6T8fKV52681T4vP7N3paf9KQN3cAWpqWMra71FAcTUM67uZXRPzV
d9r6q1jvRZmtRbTXQtoOQvsAsjy2dgL6Nhuvmkd5wE55YuuXvHG9+uQqTrWQurr86EgyDPCUXd92
5WUmWKdk6+7f8MFMJEPXaAh0gNCoXGNYYaYng9IQjvaNb98WIFQ9mKLqxg1AjLSmr5axMObr+J02
0srjvn5mroUP5V5vljxrJ0Bku7kLfOlO9LfMQxjmm3q5GI1nAQiNgjNY92/Oh8qckb4CG+IOnZS+
zGjVBeZ1btQY9lkw10CFIMM+Pq4JJtVCzB//AzWmEU+Eyi+7UUxRxbCWtYQENfpcVAUjCDKkqXtZ
KeKRn91kbSu9clgJu1NaMPk4wK+I9TMa2mhkuspH6fQip0TJwKGe45MJkvEkUJeRJeGksgt5PhyH
Z2UZI/6k3BguMRqJXjyEVj7zI232Rhhv8l0wAxBKuXE1iKfzUFWUd1D085SFTjtjBC9OMlRo7VPu
Ub+91llKbpkAOk9W5sgkcoLBPsy8Vmz2eW+60W5eLzlGWlT2i9idpUb1gqUiPpbbY6mLwuvt/jgL
hIPg+tyRfGpxcdryAq5EHiHaJ4WvcIbhnQ7xrTJM8PnZtB/DW7fYbtn59Xkqb7KftIzRX+ZDmyGO
/Cg/81+lO0BdxJkISxZdneC2dV5lvaM3g7diB8bSFfg4qLrl6EUOhKNtWnEYbhJ6YU0qKTIKbJcw
EL47vSMJZPrOTS5U5EKPUNsAiQ/8JgIp+RY9X0fadAGs++LcZh3SRQ7CgDHYiBoQ0CHubzAJJHsC
csxc7UigG7NyneHSp/R8EwpgSi1+Pydl5LEgFLB2PN53YErF9WyF5B1oZluFrHwLBmJJsrZnGT7K
r4XBJoggzrALDNBJgtGbtz15G1ZBDJ5dyaFVguCOT3cKGNxgEPLY+uXpxV965m/37wX8E5kzkyZg
gB0asrZkC7CS8L1y3TcrYeQGRTVE7yN5HNeTQnxf1va2ON6csGvb/tbjNlBYTirYDcSY9T38QsLN
YsPhM53O1uYWvtf71I//U4UEJ7sv4uEukVO3NXHhAPVbmass7QoTjzl5SSiT6IgZ/x0OYk7K7o2+
XHGJRuyhCGm1b1+cHGNdUceakMG4OsxGblcYhyGhG54ELrr0HUjDir8vdUCuukrVYknz8xMUAXkZ
2dKzDl+PPBicUB5VSiD+ChMZplU8Kt+vO79g3GrrZ5InCMZzF8WJH2weLXAG0YGhjjHj4YFo7mJ1
j4JpLjYSJgC63V+ZkcUCADgNaA/q0y7Xnoa8RqSd8Y9PdDiIfnACXEQ59YKJTl2g110ILeqmLUzB
sYF/MP571duHj/V8ESIFIqBBwoLnhFa6lsNMFx8dZoQoNI2XGQYBUlHQIssAHLqydztH/kG8BsCQ
KGC3TNNHifkqo5NTUavofxQllAJNv/W661jgpVLIPUatxowQen4+6KzRDs6RBhRpiSpmaZLbFOS9
N/l7/OSzIMfF6wBYPkl1j7VGWO7m64qMJKpkUzmOhlf7mFyE2nEXuUw8JuY/RIrtKplwMxbXaXhY
40VSBZSymV01ZqhFlwUQT+9QbShp1QK9R1SxCsEBaQqaH1wNqe8UOCOtDf0z2azeuL8n0nav8AYb
UVIbR9TAVZJ69g0ulvjHqpuTleROZJWzc89hS6FyexriF9aamuY4NvmchErnMgzsKktHPEorJ+xR
CEesYp7I2dpFqRz4vKXOepou+I2Hwj8nsgfWX6wackk8nJ+kCtYRz//eXyyb/U12nJAU2aSoF7Z8
CIdscdjYHNwgkrbxB86HusxY/8cXZ7BUyYs3z/6CFR6FheW128CT62J8QI5ww79J5X1qJCLVuuKH
x/ki0VNHtaDh1AChGZRxeBFfbRW9SkJiZeJaaszBBZ6hirfA6JYNwlsvjR33hsdQtTKn7cW4fWVR
Ve5A+hjR+iV/Rt/AuGTILvybobiRQOaHBT2rmW0bSHpE6qMzg0pwJbeLqRKmhPIHxBnUmMwygD6M
GQDTIQEHYwt2U2SpXlLxEgpgg5zXInkeG0HCAUPCEuCmOrKqsziG8BDc97cwSZ5ZXTUyd5NYVeXG
GBDeWz7X2+aYGI6hxhQI83j31CrxZQdkWd6Ulz2RsS/mouVLKbSxE9Tk+HcgXChHEag+WoYr8Nju
DAWZmVmXQmYmTtm9a3hz1yQgIR0UT54Sw2nVyAtI60AMRL9gvahtHZuvFKU68HVgHEwhFdov+u8A
Rg+re4v0XcHAVUwrqbcxVXm210dJP6jw4BEz5alE3Aiw5MBCHNpN+PvVMtqou8iwK24n4EFYDjBC
CdCPCgOvN+NNepsYMvzkWO94eF7rgopqxsvRfy0IQiuSOB6Ck3wa45YYa7LXl1ul0inNQ4tInvui
xVXcZ9eAnTk6j/2ewRJwwkm1q5CG9OIKLwYE5ygUVlIIph/qRvEpcSdRQ1GbXXuitXkkM/fk9Ia6
3DyO4OKR4o1crvoW6XqW9DuDDfN5i2MOKUdoAPW94OKUQW1nrWovcMTJSn7DZfZw/s1oFDLLU3p5
bQiC1aLwCEPIBmCcDkiT9XAcepr6yKQh0nVkfGzKzxC0dmx6uhRYCPKLAA67IAlkdlu+5dqdoD73
O+JiDgJ9AdNrZKg2bqMmyk+a2YIJ6qJGW3Ml8lA09laJi2x/whHdQUawX+KDBi3M2Se43s92Qtf8
PDEX0mFPF1RCnBLYMYKaJnfZN1N8uDZ/8bsY+SC5nm4x5OAN66IN90xci6YoxvaUCvkfGO+4XoYf
DjQKvg9dlUYv7aZg4PCmiFx43veKSg+ZNt0Ztpp/hIAqH1joCzLyWWXzoQvvFq/wprJM9Wddqmb0
+ZrjxMd8W3HrxD2rwIdvpPk2lem+OBKESoU6KaxZ9J80wyz9yU+LB3mrNYRouirMzHC6n6rNUgNd
ZBwMPZnYS8TcdWAPgpnohsb29VA/U0+ITQwYPoJykdHhs6vmFLyBg2+yyPN79wbPlMcLDCyP/A3d
Bjzx3/zE7fEbFYfUhdOqPKAxZTYQBPEc0e0Vl1C14HuBbvLxqyLSPSs1OsKLfZNC2uP6p1p+cmD1
/G/2D8fmyCF76jQqmNl72vJvNocTSz/vyMtEntxzcLkZG4w2CmXCl5uSKZ6eR8FUQt1pO064QbX6
92UrIwrKfoTkSjaiPIwTNJd74m/uiWRiFPSMiqJmBvfkMhYMfNJI+s4aUsCYupPy1GNIKyYasy2x
pF4oUze5I73Rc1luUpdlDiAErERRIYgd8NWDiYXfvBEbf15p0WHvT9Itgbhm3zvIMtdMtxMA44le
Gj7P8tJE1Ks8bQSbZB4o77glO5CyhOmVGlRyIfjFaPpGBWIwmMqfA/VeJzpfaE/QNn9bb7oDAarB
sbd9hNMcjfnNP2hLvSfXd2E52jA1M4s1mtIJGdprNxkUQd1IBhzwY5LkMqQMZLZy6Ao+syBpmpt+
wZaIw/7Et8czp+uhiF7v0NZXz5skubawxD9uWcfAiAd1r3j6N/elokgjcwYloHZaa18Xvt9OGQyd
o5BYc5zKqrbn+TKHoRfCysODPzy2vRpDEsx6muY3pIwNB92HPr+OJ+H5N0TchvlWBvcIS5m8liMu
wD2mG1Y/GItcNJaUc+qjVPo3FhMfk9bnlXG0NsaTy7SYelj+yAvSf7ygV7a35OTCTq6hVpH2xkFu
Lf4dq4fDKyCwWuFRyasLa+Bp3Vx1JWL9RbSh0OvAoolZ4M25lLf8fnQqDGy2aRIw5P9PUBvUp0mx
nrKEQl0lCVa0NU+ciKQwr1ATXQOQM+M2ghDh5f1z61iHvVMsF0t+EfeDNXavW3TfkgWF/aAExh7n
hAkArWhyhY3G1MwoBgg8UIQ9Xvdqm0U0KVPZRIRpvnekUd2h8byoh0jbSDMH3yhgo1IkqwwLupRY
vZwZMpxbePdkrmdBVbBmPPLyl3+JK2+ShFlDkvMygQ23ypmDUJQPaV97QDxkFURJEthb14+NEjz3
QFFLYFyrLH4h2aMr6PNFFWH811Ur4wDvcyXTtDS22o3X5ubowdUHhbhKbtSP7jAys5eRnPxVx+ww
aS2IGWAqghCKHWCDGOdM6vAPSrcFLmzLrwFrBIz6Vj2Uyzqke3Y+Owp/fK301na+SmAMEXbxaPlD
GUX40yXf7Ydk/Q/2SfP/YKswPDZAt3KQ87yHq3ioIuaPfAhM52ZpRgn6SOttbyASWGCuGkKPBtP6
g2i1p5B7bw6a8D2K6dkx57cLtGDyPRYIS8gKJBtaoGs0OQSk8cDhl+mjF/FD3wIHXREp3AGLCEyt
9hI8XYyLDrs0nWflB51i72lhSY5jxhh57JZm90vkAf23mRx0DgJ4JZmg5690S0HoZQrRcBmYTFwK
dbo0MIFZ2r7NLqKZ06eyJrkpm7XXrMTDPEVKxK9IwOZtivFFbi+jugD9Gy3MlHlZsok2x/KJ+Mm/
d/pC0iMjumM8DeRaHEGU3toZan3TeSm1Jru7SB/DO1DabWJWOE0XO7jPTJPO82rTHOo4tdbwfuf6
gIRfhOz6DGifQDJLODZY6Dl3dHGWiLbapS4A5np9Y+PNZSovk1qh35X8rYnuHdhQC0g7E34iQ9e1
AVa3v4xXHPMPhEb8FrOCDlAaOlxcAwnsDBl6+ntmTv1cr3CX/N67zi6xhPURy9yLNT4ZjIXzh8pG
MB2D9zR0iuwHrZBNwQTtZvDNJbR3rnUDsHgKik//ylUg5O/cabJas/SA0zqmmmf//zXOoLjdto/m
aL+vmUN+BK46pyUT4vYlk+PGOlGeP376iCNi+81z+SSmFDTPZDvv3Qur89cFaFcyBsDeHdFOOY30
C5aB9z5Yd/WatuxXajVQzowFDhYdPjS39HNVavMBq/+w2vE3USjfCEHPCgqppwWIykpYhlvMq/sD
n39poo7BWzvbFDBfDBuUl/rGmnDaiQFZx/XT5j+A7pIILiFsf1WCHTs1ynIS/s+XqUhVe7x+G40c
RIIcfcHbDXya4ultP2n/0NjdwNCBU4p2qbA4SmmTnpjVqXVKwfch3Sudl+5FUxmJYwqCDGNQCur6
jMKco9a0aTaGA4C24gAPJRi5wp/KqzYX32q0EyTKl46ojB3aY8gmZqIZvVfuwlIJdTzcMfZx9PSS
W8Zmnwe5QwGMW5fGHXfAMR4GFXD/jx3fLLzZfWSOLEmFiEUGJmrNF3VSXAFNv8JahlwFfHStTB1x
wGhWh+HAqej3Kt+9fv8jI8CgIt0ROa6MhgznpPEH2RoM5C863fRCVSC7/vu0bEw42gBERLQyRXNa
CY+9vueMhk52pvkcF4kK9zUs0Z1bq/qbV1So49wj/J59WVH2wBPWvrNW9ia4KNI/vJCIxNTr0XaK
xLcndZvL0lTS/JspbbNVAp2nNPFVfLKCA6u3DXHguVH0gLmdDRLaQBQZUGVNyJvpOF0pNfmXpsfm
07ONjmvEceBG2mqAbLTjS4YdNGWUtb7YP6DYShDkl3LusM5hkK8CLfHePlKrAwsB/g6YL/xD4dbZ
bWpcmfOx+TNZ1o4op33cshEXujvhwNhkfjU+MZa2UsSA6to/IQuWSkRJCi4JkD4cKDogw9BgeJZj
Xao9bdvexNeRAI15CKpiuW2373Hl5Q0XjEiyvgtYn6bhtpj5F+5vlwaNhUGzLnbuAwkCKDHSBJJM
ef13zc8LEQ16+Pe9Xi5VSRUsyn26vFFXJpa6avw97mP7ZxYMURv2TK8Xc6gPVfCzCapd60UIS7XA
OWBghze60BZntlvGZi3hHlYdk3JNrExjeZMKJlStNfepq7B8jPYQfzkDKkASxht8And61YlJmjF0
2p1p5yF3ZKWq8ELRp/iTp2aPWvLNSJ0BM5AfKBA/wOBGwuU9LajuDU6NSE3pJleMfCKBE+KqBCz/
CeBejuRwEeyRpT5eJN97gVbQedNM4+F83eN6jOuGweMLaHH/dFn8Cz3twLtG9poF9MRwzWLtbOOH
Dw3MfKAGWa3bGLUowr13Ougfg13AV+bN/EeqbqR8vmZpYxzJ1vVv3oFMfiDbN/JuK8cIStJ2uZJK
B3VpsjTgz06BYJpvArdCH1Hvq8tuUWSh7mhEo+vrLCIUmMecwXjUF6NDMXjLzthZIX8fTdvbfubR
RvGBY69X6RYMaZnfQx54YXe6rWmqQbEZXwmiQ+XPn+s/XXkT4PC3POh7ADPgAYObKYt30kIl+Qw/
b6mPBAdCehdbupnGlygzlic8cSkZH82uDsd2I9YrKahkOpAYBKTrdzkXJlquu/cdbKiKjZpyLVrJ
9v6Nu4p0W3P7/jyliGmt9uguF4nwoSuwIdFoWd3IIorne5N8KiuMUAEysue6qRs+lSjsBDNWdPQN
Tt3jMDV1joG7SX0Ix/TtN7emBmcCz3xUWHhTJDmGWAK1GWceXMhTimEyiTVT99+MRPQ1twYA/eFn
OYODuj3BGrBDWZqRaS5SRx/35Df//wWGyM+di8/N/ExqwCnYuWPKL6cP5+ilD2U449um1dhaD4xt
HwZXfm2Nuzp4+7QuJv1Ts+IIO14ZK03yIZr6yNjl93Q8UNPAaJiP97bM9PhXAzHeYikT71/oxu6c
xTEhwpiFpW6HxYesm6NEfHzJnzQ+wGQa955BjAw8KEXe0MIBFE48+i1F0od1wNDLnb2/K7zh6xj+
lDgC7nEwN+NVcWWKbzK4L+DhLzOBNpn97WuPxaM9hBzrU/IudRSrpcitI0BD0HWvudfDhChDgEwX
OuqPK4OCVTfIbpKan30nN20jfokAVOUVvNvuLhLmttFhptZOC+nw8NOvWhN4bWfb4aZhXabVed4j
qjmITMZ/tdUA12oAtcSNHCfZslk4oNX6N1LRsMDFK2EvoKGyOA2A+Ipqik3qxUDV8icOkKwIGu5t
dIjpoTbnWYwne8pBN22WdVni8aYnopDj3hbUnd5LXgykYMudmfK2PG6Xyd5DmsAYa7hhClM1+l3E
Gr8MJ+m1yJQOTE9SKhvWKNvIrjaNtuUj+NMQH1Wcf2oTDhY8PjTfAUQnnRAz1Fx/nyjPfEGlodTs
qYom6FxJShWl1DzednOs99pb6/z/DHKfZM/2ImkqAjxjk1iQbvNsHSp8+BKltEoddYxnUlzlhDlb
WNIXb+NuKkWgPZK0+8RY8yA5VdjbR5V37ZXnXeXnaqfs1OPKFO+eWafPbDcEtq5UxmWPN6n0iRuY
DCBl5eDqI3BU5SMl3iulU1ghMSHrPgABMBKrx48mGth3uYPGuaQ3lb6T5K58d2tLFARkI1YCxfI4
EopiCPP5YH2l8knhLPXs2hXDUFMlW7nEUCg6ypxLSUbRgzilLYb7GVn3Zed9o8CyHA60Ih4EKzU3
ruClC8DkAPbzMvIUsPecrb3fwAoiExbau2XqRKDCyvafufWFmHGyXQaCmwZ7JQrIARtlqJrl4FdO
VcAW/KcGncsz/EBQ1vDHTvn6wafklYMT2B1cwnopLxEAKS9214SMSlJ5JNnon36jVO6as0vnLRwP
n+raFGLANNGr2ZaDw5v+gYS6ZEbQsw/HQjXxQfru91vLk8TjbNoZ/YZS2umt/pHTFtcMzbfJGWkc
FZbmsUQNRT1zmgoSRvpjC8Ic4+JrMbDHfVyYKzZfldd9se/PoxBYXIAQo0v6c86ZJGemq9rPYpcC
5wvvaHvRC6bKZQW1XiSAvsba0It/tzwgMIysqgr4Rg/pnv6WIbfVVPQiD/hOeEDoH00FUDBqMblt
fkkyxFo2uSbkWuQSDDSSyKI2WVTwo39ktWX/3Q8YdRhMubqpd/ACa5JQvLt2DZKa5r8AInekduze
b8WUTZkoWy7MIUYG0pUXYHPXAgaCy1AVJkSGU/LlTdOtS+AI6dRwweVjr/NMhwB4j9oj+d0/3bJB
ZcIhhRk71FQxj1Q8eipW96G27uOqVYnx1dNpX4YVv6Tz+l7xAd7WkPPL+/9oriqg8QIcjrxCf0fT
WOoWtU/mClFP9DdrWGD4JTKJmd3EMTFZHd/wrwBudhUH5ylCjX4kKKXtDWVd3ITVnXD8rM0PIVNW
T5marFh7YfxUrBuAkdlrt7II72IpFEoz3SLTVWlGiPIUADQdvs+zklUNvM9stkbj9Ca7VzIxHhaj
ERCT2KiONil8z9txIcyEEgrUveEBl0sm+ZHx2G1wjtQPfEkuUGBLeO4PTrVeuXD8sComIskzDm9L
/nJ1lRihmfKlfDNR7mUgI+Sx3GAGSNr3bs+gCwH4p87kMjyjYbRdbgP2P+ndzjA9LDpT1/++O7H1
/jEcr3vKiuFthaDCPSBZXtmWnUEyph0b8wjlKD0ycV0wjDI7KcXYXpeFINIeyQq22gceicz3RI8A
fUyMgxreC2Km9RH9wb7CGPbyB2YcRGW6xHXKgTQtEfgfQ8ESWmopBCnC5QWedcJq/EpnJ7OapQlv
gKOYe94FJv2PiA2sliBaVwIFziQ86Ksk1RjXEy6E1MUhp2Ff8dXEqRK8Qx2w28umA+g+vap3ab8i
bCbRmshfrvJDeOO4ywS0C9sIVMV7v1pp5WwdMl99rPJZ3P2Veb2FZvoUjynePLokT0D1ApZwnm4D
TCMTq3w77dDO5xGJmxxXZaZQu9kHvOQ7r77pRNA0TZllVLQvwNN7iGQyXXPSzaujNJ/1cq+k5Ryn
JCVWCwF+fxaJJ40OpAISgUjYKTc5mRg8Afpfi+tW9EMpTl1c9yWxHpuZA16ZWzNWWAsaQgBzD5Qa
v0PFY+BBhE2Xc+Emp/LuAbY9OQzJY6iWNWeBoArhhOZu/cC9dOnf+TrbbNtyBzmP06wCFAqtJMRE
YhQToLadgGY+/7EygwKcIUsGHxnmeTdw8Nuq1vbbeWRMSYA3h70Cs55AWUrKAnXGp/1Txru2BizV
67ksum2SPDKTsMBv43KzGQxKLqV/dFfyvV3w157J2YI8uFG3gWv203qKFFLyD7KW50bDdw50t+8g
ZO524eCyQQZNuukgu4PYMfBIiYjql3A+4S6HdRpv5pkkHOzhtXu4FsRd0w0L+AxFIS6bbONiW72g
2Aaj7YbhA1JmZJvBRn+LgVS5PfH4Lm23d2I85/Y4lAQOREpFcHJX433c5d+MkuCCdUy+lwKcpjeo
EZOpS6Lfa9N5vR+J6EuHYKnzwomT4ZWNl7IMxzky1dIJv+f6Te4zfI126PzNnphAsLQKvnp7lCTT
dBoE+0CHB4PdT+ZNgF1sANfwhLoP5EZZTt/xJomhsbJFsv/BV2hNKWzEX5Zodyg+yW4HXBinOhgi
p9VQyxIMMHP3YBLYD8ydEeIKesRc0zr0L0ebjTHRyCqq2qSjTIGDYBHoMDW4dvANUQqmt95T7EjW
3CYjZJCIJrktG5g79I5Vg8Q6XEXjgNKQV8ItKnaHo1QVmrSb/Du8c3MAh0JeVdSK36YPN6ej+Apx
VC1MNHbkWRX2v4a6r2warGuUIoSHiWYniGNx0eE0BK8xMLI7z0x8IS68QJz11GFNI+g/dhNt6VFz
hchAyyfTvrWi+HPNjQiDtMHF5G2RMaT9URBPYU1jAIPhPMhtFXeIodH/cjuGhPfqzrRPXz+GngfR
uF1/BKatU5k4A+ArNiQmwrRUOO0mlb+KdiiH9B4ULyNObIsq6zUkJWlHpr9pjvlTZViJBa1Fzfp3
JhjYfPDzylzawNtv2S1ILrMEpEWq0EFczwMNkO9jtByajdVGfZpTtvga5ztUerqR3PtLll4ePwo7
r4WfDszS/yLoglJhI2sTB+AlEVCeVAp2VX15nTyynlhBNXHE9A4m6IPSu0ni0o9JAbabjfu+6kLK
PQL/8j3H1HISSiMe40oyPcC2TqRney3/gHNpG3PISWARJq4Qkpf7UeovNegKtX6dbY1RqddfSy/d
pr/NY0ACCeDvzTr7U72LL/nMO19Qo7qDjypnf/m8rke/rfKiCmvrbNMPxOzqvQjwKE7B0TqXt8oI
LwJy4siyelrI2ZC9DcAAqMvcrkrqFN9+VFs5pjA9jLZyfAqlwQAhyGdnQdzRXLxfX4mPnp18/lWm
85Nw18kU/sWSeF5S/uYJsuFa+7m29ObjfM8EkFaTdGlWJOueDeZCQuYgzBPdphoBrJZqtKL/vjU8
LCuqEq6mLMphqnGoys/6WJR1yG/16taucJ4i3ZgwU7JKofu1/3E2/sobrB+aYyEXIPZMKobcUHBX
xtleszqSQg6eBfTaaRgW+dWPasnQ/JjY/NK1RkQHwEsoZVFrikIxqGCaPmTg25rNjxzQpLYCp1c2
Rtzz8Sg/1xTEVVB8DNHyyDWY+pCVdSDVbjHMNzbVl1TA6x3iE+E/ZaZmmU9t4iF3LWRHt9H/zReQ
h943OaUwnX0uFfPyXWZC/eDmwAchk5u+VS0grqTvctABLewHncWoaVNyfHmPEJk4DWkr/V2E8UIa
f7A27C7q6WUgMkhHit22f5+XwnqFdovp6zWiTXqozgc9/Bsh9TpJzMvjO2m5Cp4dOUS9fl/x18mV
sRtJkAH6L2Z9BqHkmK3V01FzoycjFavuqaWFksYRicdfu8iVUYhV7NWAypfFMjdQ25KhPizB4xPx
3uAEgNVB2rVgx0P4Mi4zxU3AIImwDz9QE3ZzH0kchvwMcrobf3IAB3HqSn2tYMbivYG1nYeD0F8D
ot8slLqf9/tR0UGAk2pW/y+zKAxy1ueRS+jxiM/Z0NahaLvu21ttpHXC3lTIcKBuOod4dj13fTle
2QywCmU79LR+Y3860t8WuK7kp3MhJIwcRCPHX+3TzU8nHNj/XIpqCbuFExuKDR9a/XHR/T2TsbNG
NtOvBBg6ppjR9ODsBT5Y8rQ5s+M+1K1g/R4bJoDOXGEjz4y5hgUkfcJeYF336cjS7rWEpOWdmIuL
kYGVSHfJY2tbLdPb3N9ipWjKGWcXiarDBRBMzifRBQ1R5GoSabP5bA9sZbsjQOJvthH/0SfyGhsa
XsaAcP8xZZ1gjmYkAC9LGKLxKVyWF0F2wjbaM1NO+bSS1qQxFK6sIgP4Re0Qdk7FL7g3XtTtsezJ
WFyTMMMG2Lnzt1UDHVBNrPWo3uETBRLHUikiyDCdaE8tHANRe1ppw5R+HOEJkw5Oxk1b1JEQzm/N
1LLiJWtDUlvGRJwgSylwHxXTlS/TmcQA1JcFusjvktC+guslj3hzX4LyqkScyHd0gWE1tK19Pqet
F9p9WgiFpU0Lia62b+rAxqETyFyxBngvhyD/7J4ZsPGk/IywdRxw8jD/b03Ix/jdUXTvTyUjz+fY
M4rI3rCEjlIyCRz82AwBksXv1KDZU8z8lZ7/gXW6bWqoMkxmlzyVdtqV5Ch/khaqiOHcR7EHYAaC
RQvi16KRhKJR+kT9qzmyBp3rz8xy3JqZ/jQ0fKKM7V+slixnUjzWbsS5GT4zboLabzsZt+YtYeE1
k+bnvmtG/EYCnFfLXRNnsnNQhh7zVCkyhhODmG7NAg4hR9yRcbAFbO+5knxy9edddE0Sb62ItnGU
90qjMdQT8BUrOSkk3lFWpAQTJqB5kcBf5y2au20XRDqJ0b7a4U3k0Ac1QmN8CixEEHBnr2XzbJUT
tiOUenx55KLScdbfrjKuFBPJg8U59FvNVyITstdoLKUIY33ZhaBEbBlyFFUIDPfnZHb7c0VLfARu
LdYU6OzyMzTPrgMpoVU63CasKyrCKFO9vUwGAL2oeXMqeuW/3YmOFsg3Ev+WnPEwoQnXUieZg7SV
waXJ17qjb768GNw/kZe3dn0CQ2UH3xCnUWUBd+u2B5gjk0gtOCEXng3BoUG8wkiW+LJF8ZTLVVLU
SVrQ4ilTxf4CH/QcCyjgx1bM9GsFg9L8Wp7EcUjfmkb9ojxoaxUef48v+lt5awVozFP39/sQBiay
drZroskCpQGUI6mVSmSp7SS7gOZMf/l1scu/hmHaIjKyqa3ckffeoOtu5HRUqCUoObQKlhjCg51Z
CFtfuvKJfKXcvbp4TAQlYRvC/ND817hxXpNlz37sA4rmZRG8ftcdTaZ7AP+crO0+OiqIF6BESXCf
xGTUEDmBPc4e/uzjjwfPfwtSQqB36uyHJVkxMzdSJ3SBp0eyHapCQUiWnS3dvxBGqjv9Sp4NvTNY
D1nAy21AfCYuX+9Hm0xv2ieNmBjd216aWdKIXApy8ZqfqXeFm0m3YmWrIP3k9rNV4F2+GAs2A6Yg
rGcldqvCtFRXfJkDyN6uLyJ8nL7jUqnreEH5gHsCbLmsnTDghhEPda5g7FHTCd+tr59VwjhWzXc4
CgnjxDR+MaadK2gecK+jqmqR2K7NAOSVl1k2y5QNZTk6PCC63m0doYOX211TSxkLvFb0QuEjuxdW
faKJ8oANuTOGhs6ccUHq3NHCxtS7olitYQGuQEca0125/vkgN9U6gtkWeb0wXpLsgFccl/uZmzzR
M0iMuFFzWYedyr9nnpQrUjiBO/dt9Vmk4EJJA+yu29Ef6QlRo1Q1uVaP43d3e67pDFKuYb34t33W
GF12yBYgK9jey3JH+0zPbI2lEYD3qTliGP3E43Cy6j7n24VzIg1HVqudCQUc2diwjoLuC8PBQFVY
dXH+yMp9e9YrSMhD1RZDLrMSsNcHma6YPRGeP8WQi0+8ej1cJI8KbblFlN36FufufGyz2ymv+Qwc
Azg6yFhf9V4/QD3OsXGOfeNL2n9XBa/l7TgMhrV75PtQoQJu/MZNPThfifcf8lDoDb25YCGUKijI
ktlCvRdYMwC+kVs6tPlqKc7Fz8IuuCBTiiq0f8VLoNelgslXE09OHyNvzkHT6Z9MJRUaWY473/2r
sh55KisyH6OUY2rQ77UyUUsyQ4IEPI7c+zoYQCk5dqeXtTdnv1s34/Z4Er9B4xzrH/5MF5XuF8no
Is+1yyStiVcchhWaSUTIEYSO3YAUZJKOb5eRSwMUM6sOUij04nU4xdZW5WJnaYwVtDOT/pOtDhk3
Uof3D+KUR/qLyKg0b1JzWGHWnL4RXrhsmSm/9NSGsNya06XHFzR/nr8+DnSitbvQWt87BZQ12nsQ
xgLKzDe4te71c4UP+4Qv6FuG55mp8yTVgTSRIEMpfSFZlX47XEgxfSwBgZVIQIAQn4bmPtQ37xJs
5nFQkxOaWaLXD7RJCKTuEBFjU9sKMBl7bJKDAV6Djh/OznUqVc8aX5YbN9Han05GOpgmZxZ8Wf1m
slAmBuPbBpZ1RwkrX4+znDP2ULyuGd5fZhs7RctOgb7fgpj+qAOhnq4xR8IBAMU2HMVezP2dCrk+
hnI8XhsZhd6jKTRK/8o+Nr5K+LItCY66x1AVqsOE8+gP6VdYGbgq+11kREylTxjxbg4EBpuDDAwf
LnjWJTeInns/qf3nOhznxkYRx2I36OXvo9NrsdWYKOxUPM7RZ0957UZv2KWwQX3pT47ogbS7G/0d
fJt7ju69ewGafscfrj/kQoYFw0MvnTh5Lp/oLZ5tN0xiT+59f3iZiaCIxPSFTcbP4ztXpQ1roNl8
1NEck+OXnuNDaQ0hYhIcQC3L49R1fQn3rai1rmUw9s1RtkAzpusDxKFEs5C4uTu/2seIWzfr/65e
WU0+Br+aPJAqJ8egg1dMbxUjGLUlsxpmyTd+t4SkkBb/QxJdh9g90fgtIoae7vnLzJey7K3QgihS
MWf13oFS9mbc9ZKr34a7UmJGSwBEsGSMcx/HwP33ZrUzzAv+ypw+s+BGuW8dX5v7jZqg1LCd1s+l
aNueLI+0/DGQo77/zKyzLdxQB+HLkyG0T1vaIFuLOi76T2AKSGffwS8sLkFC1HReNUP1ngdanRfN
ffVzNFZhhpso9eryuOZvmg5ecVnGgsylPA5emOMrCFHvh9gitdYPpGPMmLvKZLWnZrgq1nbhQNLt
cxZYFpSEcIwTK7PzTs35brHk3ecEifqfvS8VlxI2jG27hn2TV3tY5rGF7JKfBn1g5hGopn2SYVa1
ERUp6RPvjOr7oAwEn567xd7zPttigIqvhLqiHHg0dkJwj8ybpXi5eiEbyEbKQpYgmR45LNRLBAiS
nDTVGErZFC3NN736oFivUPj/Zp8uSU8lz3kgO74cIlgCsyYKH0KrC9mHNV7AssNzGE9rD/MNKYjz
uWMVH0z3y0lUXaVro6yIb6UuuXZIRPP/SdPabdfHXsZ8mrz17VInMg4yfQNeq65PQ94uCbQv1iiQ
HWzfdtB/yQSvszecpQne12Dl/n0UIpye+AIHfszxDe7PWwURS9yGpxe/yRo2MU4eQxhzFr2E+lJq
XCm3m5A9finbqIVYRUbiKBTUWte5S3vli1IKejXJu6Mi+mrdxGNVC9IG97c+BnFVpDUO+MnlO9pi
os5hmPQ3UjFOdWAtkueedGBfmDK88zgi650zehaD0/h1e/tIGkboTWqENe9ocWbf5R1edReihtaU
czTgaA6tIYE8WVzsxOUSoHZFVECFs0sTJWarwG6474icBzwafScS2CqVMmcIzwG0jcUIglVwmc/6
qFetGxrRVelbETGIvsqQcJwkYSDEjrqFUcByPIKhg6hiBR7DIPqUFnxq52m7f8dhU5QeMojWWS8x
wvV3hfO0/H4W6sVmaYebVfVdJ4E9mo7jhQpCZn96z+oyCM7y7b15yIknnkGDBj6pW/B2wk6X3VB8
evz0wdpqAscdhCb6fD9AMcOjPk32vqHw+xOQY+7Mn75Z5H/tgCBPTNTtHw2KpH92dvnulgKheJg3
waeXcZ4yGiAlIdZQFGKLcEWSR3tg6RWfrpZ2xO4zexZc1yY5zqLU9nyLI7py4BLl8QyAjkR7gvvP
T5bNgRjhd5qJ3CH3WZYM9QnecSxlpLcbOymuLxrEO9HygkwYPHRya6if/O2OMxDyUiQ+To8KlEJL
OHjMoV712uxVvHRm3kN2Ivzj8DRSp7Xn87fP3dF+o1PXWoBCF3+2+Vlw011MtMllT5tbUK1LoeLl
GXCgZN8QTVGTw62jE61aGuJKWIRT1N8byWUIllaBBL7L7370QrgMXjUg7A2k63uVp1a/5Y1rrydg
TJF67uNEajBGo/tcqCCs1ClL3/AM+g1m9kgpxEY3JkoAKLSh1hwFFeFjVjivHSYtmRNJxCIM2JIe
KUBDJm5cZ78o8z642Bi3xrknNPAMsZh+cYNbBNkHI4QfHHujnY6Bxqs2kAcz8eNrNKbruwYjYx+U
jPiroOwZFFV6rWVSe7DQ2A6uyclBq5XMxdX90IZX440g+5lD5UxGY4TP79YByVv1suk+m4IRF13C
minZD77ioR1CODgegwNH8RXtGSjYzGBj1CxMCDoYmxEnjHQ7vpt/Tqbi8s+JjjJh3+DBxREOUxZ1
TdO+fntBjcpX5xhe5cL80bHOkE69nqbqlDVdCIhR4bH6Yp2y/V1V6tERx9TtMCvEj8njVVXEuhdg
tg3iycwGKiB4ZZssjHZe8GfWQ/cc/MtzLyIJTdpOqP2ewz6GYeHx+4lcEvUauU1m7Vz5h7WjwKez
3BxPa5kx+9tDHlQtLddCrDKKAeMRGyvOQLsbf+g8wIP+7UDc7LmzfMswIR7uffqxcIWjc1E91t9U
hoL1oPEi5jYY7UzlbX0RJ1vi/tZRx7otIdmq1nLvxBWKR07YMYQDA/JG8Y3ZxiTXnlIuANhC6RjU
koj3YQ9ObHSHZjUn6RhCZ0mxyLC1e0ZqleVm73KmmDzYSGax29gl7QZ8p2y8rp+m3bb6lwW2ClPj
4ASCXQNz13bgwVac7obrIAv69Q6YzUoOf6pLwaq5VKud5Gg8MQmo983Dmv58R0M7CMPruCnR3nkT
09ITQ6BWrlkqGxR96aQnCQ3Fc1/LuB2CwTjt1QXzivESVSjj4tD+bptmXHPsoT62d5YjZ6YzKki4
QyJJfv+GjQDKqeSbWagjGatPuCmEhQfsbhixdAb7+6J61muEpejp2vBJBsch3K+xruLoxBJ9w17s
dH3oHYFNccdF5GzaxuxzKEHGV60ZRk8ER6/ZpebGp95U3c8aGOfV5X9EGS5v1yfPbm/bDH1zVhjC
JzEG23mNb6jRLgU14bnRmElucGZ7YoZ3EQ99WI7UrAt8tWoIiyd/5MVcKrogm6bgvswMdZu+b0kU
gVQKXI4TLTYcK6SkLMwO1nrNHB7lhr6i4NZPzhjQNdip9S3oJxv7jMP/9DEp1tlMK0UV9eRqwFUA
gsNbtbq8gfODNqdTMo+yGrE0jQ4rcC7qRJA09cKBNUklJkHebn3V+Pqch49hw2Apbe/im1MGEHbq
ytrklwooZChMXMuVdkLrA9owQLFi7M+1Ll/Z1OulFGNoq6Ccarw9C4G4odRbWpksw4yvkoMAVS/S
6AiVjnrT/aT2AXdJZt0+Dr6C33mT41hFuJ7MZeEY0Bqi+Ofa4kXFUZU8hIOseW9ONp9C+SsGS/BO
E/Fn3IH9kS+V1mXwfnS1L2VkRI+rR0zL6zBc4JEYvciPakgI4EK3VtybkBWLiJquiVNyXsHptT2A
zg2Oyl0HwuQO4Ei6elrGtwZ1Qs64e4I4jJO6LS774epCk5xkdvZJJQCLwjwq16EQpTwPM2djbuZg
gp7WjkMu+7e0uf2CP1NmeUxc93JCvyELAvC0L4ovpa9pj08GUi8kpDD+0B+TgGCTpNmyLO/fU/WO
2pUGI89eBJcJ86OoXC2tLtusNZN9cVp2dpwdsDJdsSLQ3ADmP1ybr6IuJ0lDpEHlxjWRgsgoHnKd
c92u+el0iQ3/kSANzULSC/9vqOwKI0erDq0tSY368V2h2Nk5lKeP1a37BJqk/7kf6kGitoXf0FjK
pHyc9NBNMb5Vn4j306hQYj/3NRdcll2Hv63ppQGT2zQzZKCHyV7sZf4RKjbETu5VCM+/fSyMa7DB
x3W4AsndqiBc8tTQu6seKiNW8H/HsXo4Zg3fkq2hPZ7KZtDTtmxKCR+eXkB33PywimlOlJqfYQht
ZFxUViqlExlqKBuz/y3+MfJWvycerkmgK55D+HfyTaoY57Lc26dLlT+P9Dn85aRe03rWiul8f42C
fuvVMWaSbaNst4WbGf7L+xZsANT2DQyIJTQpKUMyHXTw8PDCFPWbJLjRnrtj7gHNSyyyWg5/PFnD
YOe3sL6XRKIfPeUhJcs9uKwdQWzhYyEhY69bPPZ6Rf4Z9xBKv9RdatiWFupFcglseGkWiXddlWFm
F+LsLNu+cDQi0lFWaZAMSqEOEvp4qwCtBCWfdaVydd3Mbg/pZVSWHa6lfOi2ydQci5+PHYjNTdUN
Vyh+2iU1GOW9/O7ztov9YGMUosb1agG150QjSwjEK7JRZApFXtdhh7VXR6pgxsomx04NguFvaSGO
6ZCU/tSFaa9KxcruUoScR9TiT26ksxZeE5HqTuaDXn1LqnuNaSgAaJZC8hJgejSAuWZvVXUwW4/V
WGm2e1PVjUzAYM9bCTPSM5Wygy5bXZTvR05E/e6AjOWTTwUZdoC/Uub1wdkBi+xJ/djEdL8EDSke
oAUBMh+5tMRL6Q5N6FI4RObUC4xZ2GuNStKwf7+fH2gDAa6CFV7joIWAWsvak2lOigvGBPyWj/5N
cg293I+oxOSghcu+kjbDhDXTI5+g9+P2DqRoP9nfDOa7r4H5HlNkTZPiHaypflgD6omqxLIcwZlL
/xFTMcPlqX94QLBDBi1+xB4yIRtA9VZ2KlQo04PY67qXHSYQVxk+vLtkZnEC8UeVGs8s18GgFVsL
bKT1vjAxF5PEwXk2pCc6ZsTPYb2gY6FHE2ZoI2FbLoJr8vPyhUbAQeWQp7GSZmYVTGbUTlnwzY+A
aDqHt0JZvNDPHNpMc+637WPttuvz8XSAeff5L/BKxCvgUsI4F9jO2ttZDTBJ/BvlkuwAB64OAlAv
biszlWkbankNqPEnFju1C5xdOwO5C3EtgTKITudU0fAXUJjXGUZwo3mZ6aCeFSb9adAYAwZ4xlwQ
cHz0a6Aa+cC5GUx8VVUz23mwvvo//DiaOI7l/7B5cpcM5q2XEv3z9AZkTyNv+HQynNN6JqGLKWJU
lsaTEcvn6xC1PndVgjiIVPPTzie2g1yqXAUiJmdfhaWRZHjV5V7oHvDaNDE3WP4sEjfLdZACCfUR
W7Q6MM4CFmtidHyNFfX2VR0S8MkNGcP2DVso8g5AtaIw8cKsLSRh6ZsDF45dRJm/lKoZjdQSbOCZ
xt/iDjgOsJsF0aWyelQb7UBu6/hm8aDRg6KqA3que0RWIi4XSO1tSaOeVgvO3zVl6kX+zZ6IVMJE
LfNuDBIEzzIjYvcpQBs7qa2PUz/bo05xQIm7LKmIfV7Nyj7nsV/mpgTq7J0lgOt0tmJ0euCbwh3x
xKxUvyLkFzDBBcjQ6X5GXA+D4l1NoXwkeUetk2pYCjEa3uHeFyUe/92UdmIy5vejYxrABLkzthoe
4UM5Xpaxd/umTABci5I1/xMmeLtfMu2XFGLmADWZAi7Z+b8QJMK+7XK0SYdrAi29YSzKAyErkaCb
7HSn+KXVhITbSlNO+33BsnxHC31Vtb2ODHPJKZYTlraroHG7UYQOkD3+OXCQPLkeZPkuTy5sY/ve
WFltI+T5dERq5YtYUKpbPTvjdUyHpEsd+IJ0KHEiKwvGgEQF6osaUnb7e2hT36WSDX53pH4Oj9aV
FEW0HNsj0e38cpnlI8248mxEJY9wAvd5v8RXCfB8LnhH14gyfNeRyRgg2DZIbxyVZSiLolNI15Ra
MBny17lLbniXk3hjpXK96pit3USytcGe0UOEah/fMAWYU8uMqHoXlO5MKLJyGBeoMIDcSK6pYKlh
QS78pxdzfQqcaGKAi/GdNYN1PuJVS9De5BXzwJVISWG8vVgNZaXAsH2klGQRSMi/RSvVsxNRXF7t
V38x4r5Xs9Zrfvehc5OhjYFjffCxdZHx4MpQXmGLeOqi8bDnsfgqyit7HvTtDGnhepeYmx4Zibr/
fhUcF7QrpbcxvDdtqGcBR3nZKBzwLMGyhaU01mN8uV2WedIdSH2j4ptTtjWsRY7TTaI8oI6KHYHr
yp9heZcupoPT4+VKrLKL3HxhWSd9cUIyZqsRVvlg8tKXJSERahtn7nisZAe8i+kuLHjmno+aVGGK
SoQWwBWO/N86tDvkV9EdVp+eC6T0NzH0uPdxwQb2L5zY6n8FseUJOc4mSkxNLZGPxUtk/XzQaBP6
Xbn5epc3/QWmc9I1+ogC1yQiiqEmDkHF4I67T1h1LNtA4fM+yxHw/+ltxd0CZjomDDKQL6lb4ZZw
x9oPOGjXWtemk/qaGZQUEhtwN8IcDOvs4xR2oeTR4z+XLgJPDSsgJ487PlCTOmhjg8DSOp5tG1+k
/Qzmqc/YJlopHpEl+i4gkWldCdiYB9tMeTuGvcn0QIZusEGgddlbQwwITHtOArYk3ebE+FhKE2tD
QGBU/UTr+L1LYtAmGsRUbrNPfv5N8AUzoRbVKnIcNhryuUIq40fzWT3XaCVxKoxMfpsCT4MTh9tl
BFtim5lv4hx2akOX8wEPe7P90uW5Fx4KW75yub53zhU5q1Wj4ijzgGWiWOHmSh1lY2b/9CPc3vrp
JLjWCFmr0p0qb9Aqhy2kP7WNnbsNVCYpP5R/S8RQrHIxBPAOJsVJLOR8OW+amGAnXL8F4wD/eC/t
3j+fEd5ra/R/bLsMPhVdDa37pBU72ZRD4gm1cSDU8fRm98Ij3hWX3Svi8DYC5sf33Q82QXv4/Ggm
ojf80CmVGh6YbfAA0byMqhrPKYTbKRGJHzMeyigtV8Yv35FJ5IV3ydvU0SJpADofKDqhkw2IlPXq
TwkUiAhxs55CJjxGBsEyUOjDGsOwMWM3hB4Wsa6sxMa/Qc3+zrEnwsc5W0pq4kDvfK2jq/GY5IOo
GfuQM9AwF+PZGdtjT39AC1Ac7rxVxLjPK5kLElj4SnIY3baKIU4eZefuSIosLGZ9/s1vPUiwiHKr
ZQX0P3NVswsXzXlklgN0RQakIV1bsGIz5JSv6YRPTZ4gKZPgYg4KLngTCrZQUjh4P14sgRgTD9n9
dtDgI1zF9iPaa8msB0icMq64Zs4/eVWw9jyfdLVETmJZm8ALMmVeai4ZwkIRiF4+SqWQsLgWk4OT
XUi5uCnLx8GEmr7Z5ShbMqBjVgTazRBUhuyHueJ+l1+FYyKKuokIAfwsZNmgcB8QB+i42/oMxKMp
7hVQRS8vs5j/OHV4zL3e5ras/CdHElz5ZqG8Xg9AVK3JXDlFzQ9bNbWa5cT+Gd0SjyTFuKQyj//N
OcjzKJdcmXKS1SWx2C5RFERMGgUH4sg+rlgx1BxRm6jPP/ZDW37YR6HQkqHu/fDIs9mTNeKaeK8i
4aBmSj8cY37MnaL55Wvp6/VAqlqcyFLiMO2J7H2ZUnthoz8s2dEYNqLirByCsZtfGJMudDU2Ivpz
gz36uY8Wp14uP4kqNHuqgebppoNtsvAxMCKA9+MB67Slud+0Gxf0vvm+eOEcEux06YCiXUL2KMwf
6cYAeFdsm8rmg0v8ESbBE6RWsPP5riebT27l7NvMWVCfbgslYNqpKsf7Q9RzDpsWZrT6+wCT2QDC
/ZRZy/C/qwY8bLRAEGYco9tDwp5hoIh2L8L91U6lWRNlqS53WfSUExDqxKQ1cAg8yL75IMdMhzfW
3U7y2kgv9/FCk5rczUtMzbYXwVWdE5CCMAoTFj5EJAsTIMsWfcX4PnO1ewiKAUOC0I0P1K9wu5Vn
CdKRV9omDroVR8PLVugBraoZweSaiGV4fmKfnXhPw7zXE7RspWjQdcvOGub3d9DMB/dW2BKS/aWh
21q79uwUrEBKmnlvVmsvGWECjDqxTPHtmH5l+tquHQCDAYTA7MH6manGbMM7jUk9zATGAFExNCG+
46Q1sQXiZFyVulQtYhb+f+BBnrpehV2booLEnuyj2XSaLCHoNtZ6CWh5B+XF41zOm1PAPlVC+Ybs
rSLM+zV89BmW+Fpgq+YUnixia9hdlJzInpvbnd97FItP4vzsbcGOumBzisHbe4peuUvqOmNsQGzS
jiAahT9zsmEbKt6RP5VymDj9ljfgPTACTmbMvvxBuCOJ0U4seq7bZ85fmprkmrAqkKT4snCLjnRb
jiIovXTnjBIJnXuEgOG6oTHY4WRY/P0JwBUKOtCMRlUyDBTw6mj/7byv6iklxdDygrAuvvkGkFit
hSdFqoAktjH9PFdFmfgzTs8f08pT5mCrJUsXQ55+eswVNWAVSiKACGCjiT0jrbuiIdFu/6F3dKwN
K/cEl3nETu8TLXxn7XsSt358xQhhstPMEFiRYO9B8OidL309sZbZohiW3/8oBEor8Qgs14ZoMLHx
+jwnvRqK/OWsaod8Ok5nlkmHviRTEBZAz5LpZe0dJXIBosATGBDIxVF4deL9RDjlkfMWN8X0zGkD
0BmvBKSHbpDwKqil9/5zzYA7BCiNNHD7zAaH1Ce7+YlM1nufmdodwZgmVGpYr0+D6dfNKEhsiR0b
zQaa0wM+E3McF7Im+hKwgnai5+1+3bluiuKbDkRT5zQQ9OoiW+a8lFYv9uadJAnzPdsOcx9dVCin
3zC8Y8AvoPUBbhEaJa7R3bNgd/OwNdHZUdehLfhUrmUfzZNjcUKWxgj+5eONfrWEOZasXKE8GE+j
kxTqak4LH62QdCLUICTdivGuygw9uLsPH/8aCc7X/Erg4crt/izy9pnzEs4CwVMlISf0ESOguZlP
ylxQQzWqtGkZ2q3ukCFAfHAV48cOFZy7kbjGoCqPb1Lxlq7MnABLGV3lsFF4NaKdaZpbaV7ELHjg
cVzltAxrFVBUHRDf26GJ+YZbPzohYWe9eNecEXph1YnL3sT8C1Uc0YR06aFfyMqp0C1DCEDdG4gd
XzPHu7mGg+lS1xW/W7bCPo+7OhHIInarXx1S/eu+dK71xF+wHs8Z143MNIPeBKhnhuwJieqYVJif
EWrfQ8gat68qlMeAfxJxa5Kw6+jYFHifkw/WlBmIJU2RNiEHu/gg0U/0jy0xq+wkNfq3NiBvUOKV
swbLpfppmIptMSAmZT3jKC4xs+87Y1Ob1I9GmZIZpGQFDXBEfJ6QHCOvMLjUgsdONvSAngvtIr7W
IHLHtbUcaz4mM5irw/TKOqPZBY8prfEe6mdSliNCwiXzUqxvRQW+974FHG0h1x+/4zpPe3IhecC4
D1v0snaiYeKzPmy1hd9DXj5ZChM0ImSf1LA61eyPmIYvkMXmx7PEEM1YglCrDGvuwxTRBg7sQAdO
sZD3oAIcSsU1i8QLKgezAQk/cD0pDH5VM3I/VlODvTUWBnbdKT8gtpo5hsNjfb/rfLuULXsn9S1m
nT8Rf83rxIpHHGs8tz7Y+nAuz2CouTRBpVkVVpSiwEahgNpmDmwH1wNhqIgrKDHXRNLiI0lmdnS5
sxR9AuagJP03WOLGaHxNA9TJ4w9jyGMtUA+vYkzUMK2xI67bOvwpn/MZHZQkQ57WazG3YF3SOPS7
PneO+9LrHtE1GiMRq7J6oXxGYID50Wxs/PFEms5lib3lYxxbwrDT7tQ7aU/LIzoFyv2SrYAiksnI
KjGcHDBiXa2MEXPM3X7wg9CXNoG+WTax5AOhHyj6MYAQQmcrbZUP/v49eQOvdPAEUSvpvB9Si7Ay
M44i01etDdyaKkgYrSeKmM2W83AT21CcBvmQIH2TjdL8arbUXKtVA81/0203vOoIzX8UKSJysbuK
wjjBEIeCNFwLTV/o2/FifB6e4/XeJsd6M/4WfxAGLp7sOggR5hZjz/l3nqZ4bgZYeKJIIER6+hdZ
4QjGGIpO/CheRKqNB4GgiJ4kcUclCYmMfk6cyNt+66inSiwTwnS5zTs09sB+UN/hyJGi+aMvfTUQ
2pSGqXALRmu9TGmSubMjQrZo1wk9o07MKHiyJBJ19Pq9dfxj6pyRqRs/u2MmB/D1oUFtXtBRd66g
lGbpbjI086dfHcQRpIUK9qH01jhFB3cU8Ut4VOmrXc/nxLqeIfSKNI1s4M7o1GC5fdXO6gUiBqgp
Q5npKRW+sYeBnhjh8a/5mMYZBPebs+HUB7xoPnALbpPg
`protect end_protected

