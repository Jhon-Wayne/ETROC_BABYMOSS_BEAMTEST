

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gD7l84kB+WAh1ATog3H36h0/cMgn9QL5jGe9p9PjvP7N+FJAVvGVlrxcgBw6dZaWDNZqNANQuRFv
ZSE8fsSCFg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YQUcxim/tlzHeVlJ7otHN7u41KO3Yg5DFb1yF4GCsbXGLtUvWNlkFjY+UPIlgYImR4Zo4dTHJQ+j
3BaUNSUOqAVzT9CfyUelv2YD2ZTfAtzIe1Mboyb3+StKnuzxnZmIhVPiZlowdW5lQ1r7BjDPOsge
ztxOfUTbvYcTUE1ABIE=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eu4MFD/NMz3pssr62VCh1XDd9mthYydX9VaOq3lWUwHi5/7e5dl2SAWHtYwTnBgGPY+jCcMycJhy
WSlkhQxVj5BsMm2aAItwXFvH2mSbjlPggtI0/+DNGQ4x8LQSFLTDYnnQbBrHlJymsS+/asMkXACD
SJ2tF8LF5tMhAlMPZZ0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rNAzbNlIFUMjdhvgzZ2FokzvR4AuFtV+1AHGDKa9QgeBsZ1e0Fom48uKbJ9iakvqUoUcKKAvRzeY
OBkbx9P7Imx0gvIgzFsgiVw23cBYWOhbhSqVb7mef9aKx8yeF8T48n7gKldUkwBHIPeqaayRI9/Q
HCZO+k2+HCjRZE6L/Gzd+IOdEVUFOg3NtWFPk2JFkfZkxs8X7Vg/xxtvH7uvp+/EbVyiMbnwDT/p
NSqOyA+rJwBJYD3xRIPTFDI83XJLCF+1i4E8hyu7Y0F9MtjKugqEHwAG+JK3jde00nzNNaeLVUQ1
OfFMZJpkk0Cg66d2cvJY/G11oPkmvTq/JZ4+5g==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
apuTRT8aJu0TR7Ciy6ONiGK4AT7TUEiokS4gFf1g+kDg6PdKk9VRun4HKszIadRtahjPQo0of9uS
yvu3GS4EQo+Y+T116wnAIXnZSa8EQaEsDkziOI+rCvXv8IgaPYN8Cq0aRlASFL7IHOWNI49V0c0A
FIG/+5U7ZyNQFCVwuE4gCgK/pA6apm5kY4FGJft/EdZ5YAbR/nCTzK4P53+XsKHrtGfw+/MthFWz
tI0OtloKqc7laKZWKOVFqWq8Qmq7UL6utFODtxEQqzczH+q+Gw4rkUyOosIY+cbB67hX+GlmXXEF
jMwvUcen9t6c+wiH6rmBDcUIiuUHHz6q+jCwJQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dfDj35aI8y6zqcW/IHFxmCDw2mpyex25qQAUnsL+tIRxivv/85PqpCOrf3b7NWnwUKMrsxtw+JBY
mtlPsVxQKR1gn6VkaHwbEgwxXXxFe71Z+1nWQhfF8Nt55jGvq1joWKMrurSV7Mo+HkvHMSszXj3v
8ElD0S6sN91oml0nObejOhxzHf0ybK+sGag+CFA7aBr4k4rYglf7AzOYrPl3nNoCkyrFDQFa46/w
SXJm/os7zUHbsDI5GGUH3BU+NktHZV6GK3iyhtHTwrMgDtpGk6vKHMKULM1Gjv9g1/jp9Ao4cUhr
bCVOXM1v2e8A3564rmh3if78zTzCKamPRAB5Ig==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 962560)
`protect data_block
AabbJR4gDsagM2rIXw5Cn3fsEgtfvAFWDEsk3bt/ic5XPdOt4RpC1+4HvvAXNrquG8eNK4+0eHVp
B/tmPSroCfRZo8zCJuIKa+gaQU0GACfGnhARIPmk7XT93NH9OM0VMWbCa4w0xk9MUFa3WBpKybd7
UPVW1h5Ns5F/mfFqYy4057xW9Cb4Uf6ku48OekDc+oHZHc2XbThfX43cp3/rfn+cLChAh+aozOJs
lUZXQZ+ejsImVBVpbk96Rld/fsAVlBU69KFp6ZiI4j0VstbKXq3/w56CxMf7AjjGCyxhGuhIatmL
kHS+H1PpQX7UkwPME+c/asu7ngeYhPOdlK3qHkTrI6EB9mXPy9uhMhtafmHG3wsrL0NR5WT+yidZ
zuZlZaCKFgB6hPAPfzw1JWGTT7AzPj9qTnTHQXX7NMnbyZJHK51dtQcIMZ22gLdeZHPrZyPFrG+T
LpRPUE0kdSpiDxejK6AjSmLcsXSglVb010w5yPNVF0Nf5IujEQc2y3aAvdsC3GZhnRPbKZ7aM+Nx
voU+uQdkhVOp2sGG+dYMcylChHvtetdpRXuzUoFZi0tdCKxcO7i1XPrlpPbeob+OV3g9uGJFLVbO
8J5CpN2I7PeIy72ibduNRjndTynlpO1Y7Z/cN4KtEWGrA/MK7WIVTKjKe47ABavrp4/EdxOvgz4u
wH45erXXu0aHjN2Sdf0FsftfXgHhNRRZT2NozU1Px+a8INusAal2CLojQkAxZseWhAssYjtBKUaU
+rM8hO7u5EVrLFpwFRbk8thyZz27ptBtDLy6r8n0wifbsjNwYC5tIjZ0h3k3RkVj6R5sxGR+VCzG
OyWw7WdMEstqGAs6z82Y/x80uHHMsyRab5D69YJJgG3PpEwRWlAFYQ1ViTVzA5MR9+CG5KojVrVh
RZaGDQi9UFHfL5jOUX/+bIXXE13NJOZFtTvCu6Qszw5roKtlrJwHNigsnZ+//RD++jmkgk8eq9F6
Euya2bhRNvblYC5jPC0NaztxwkU7EoG4SpNCM2GuqFbabjaWTNhtbP7cv/wKdE6LyFpIF34INdKE
eFoDVU9bpXBP0lgxeoOmcNZxNzF3RZRx8xDA2y6oKcwb4wL6aFHvamo+nr4Xl2p3EsyhDmH3IzDH
62F7BoosdRn0x5HOS+Ca8E04q/ETDpOI97oa4JNPMzHiYQcmbKhi4vTmcw30PRAEW6AqEAe/bJH7
oZN4ZmfEHt0BG7iHDuEhmyIqLH/4V7xmfjG/uS64gDXBpYf/Ik8cR8yqHH8UFVDwYHnf0vBWThN8
vWw+OZ2r8+5pQFPtGK5UduXoKmms3N3I1jPNAx1weTt/8dnmEyuMELrdbwYnuc/9z5MB+HnlbfuN
mnfoS5IlOnvlpwN1iYo25RLyAncmnrInxQjbvQA5Vpr/B9YV6PpgIXfZ9WN9mEjJk4heZ/H9YSZH
75OxUJ/F0iJGxhXjvEFAcM5XbzcBH4n7CC9LdmRXo/s0DOoW+UNWo8gsAVfzPonhhTLc3un8pjXV
BkPole9j2k/nqdXyvMfE8hxpkNjm522pRCggwBenzPzvO3gFu5EUGYCzBd90LeHkLOro1KoASCSR
ZC/5srUzWDxKRm3yatZG5u8QML5up7WaKGS46uPyQaAVIDVa6nrLMt7LCs255YE8H5POJXHzqxLX
rfa+qErTnBvNeUySuK2k3vqPEEFV24LOwotcmRIgfiXH4Cot9vAsdO/0k9477YX4amgzEkyQE7kN
1tszdVAYz++5d4tuu8WnRklKGiQHzHezNmB9LrU/13j88F35aKq83noJt4ms1eYe7I/Jui77yBCz
gxqs4N5/C1n/KxTts2BV5WM9lz+FoXwcXg0DI8Jo0XgHAgZJwQMiOEho7/GGIwr/GHiqGqdzC2k8
6PHWUGPpJG6Zoz8yM/HOg8t+eJGhAHXpxRW1XHsxhWwgVDqbgigG7ERtHYfite9M0c1HZMC+7lDc
4p2V+V5ynWrky3tSr47HwfUj0UqcPbqApFr5SsWt5JkHy3FFmOgrDq5CBQRVi6+fU22A23uala4A
EVAAfidqb78DYlRgF/HJXVYf6fKXBjd0933DOUlN2Goy5ab5XdHfYsTFKeT+t9Ur/utEOqr4x/Tp
rjfw7vUfOEUeIzajF7GD3w7IWQTAhZI/SZ3mB0r7SBIuPVj1xJEepcvVtQMkwNkTQXIvdhFF8lNr
aklSn9OPaRQ4heT/CG3WVT8jz3cUnATZPsAN7NoM6bqviqsmSExQtJNwdrbc9mnlZmjsgX1TyNKd
ty+g1RRpSBCM8bhjbvXt/W3/tLmBe1XXQGJELEvJPRM3omZAA+IoTtEY12c24d+hxDh0a7UmyH6f
F4qErZrKZziWOyloKFSmqwXkK3vWxzrhaYItbf+q8rH+P0pZDxdSsyt1ah4WSPp2PIcKHbN7gsrg
W5Y5Elh0gTu2YsOtbDZ1MooLRmoe4woPbGIAQjIHC+jAl2aFBBzPD0IU/s3FhAg6I+0sGZoCqcsz
fw0hlohh9ceCelLDPgY3zrU9vQy5vqUnyS6X5I0uoDA/r38489wxXozIbfwbnum/uU+iNpLuHv+k
AKH6MZklFgE4kKO9bYQEI+ouvbo1xRz2XvzBUu++pqhtUHBRs+yT9wXVke9NW3XAONgckyEFrgei
S8E1gTaEBA1QT7cEKsZFwyNhj5NblEY1DbuV9OlOJuhozCbDpwkioC5wL9fs2a4+4gJRVV7h1DB2
ouTaNkQiMfj5q+GyZKPm1v1g5+Wm6qJ4UEoPLIIc19PPtSspCImSbuhCH63wR+y9ByLFIiIjJcGO
wwT92pkg7f4RJqU+uejcanHpUUUniyE74A5Jz1cFbC1ItjgDvjobfCkvUXVSWydwVFJTYd/Vw9OO
Qd9ToOaP0xjVs0HwKaciTMA6DTNX30yFvnPODM9orC5UkpLqtdrpxoAudVTysGu0gmrVRTwVPr+E
tzdFH5a3EjdwgKFv/c/nRk0NOH8nNYYooieHbMwGnixYyWQYSG90QxxkgMtObMZsXO3rG9w9D5me
iTlq1k9TXHOlMZFBVqg2AAebAib7hAqkxRFNw3CFsGm43otsJ3NPz4+pk5fmiODfuxKZ1ygE+B7Q
oTC9P+28QDAgWptRIk39F0Otj0x1Gqwe7FCaKTqvK+3tR6s7iXkPDm5ofMlFhQoIuwVdpP4tBxuc
O7z05paPEoMYtBl+fuAl884I1CWlyAucdlufrctQ/wPjzHGWqxoU65xbCq1dXNVMSpekB1CJAJUb
Pz5B9U1MbS4h79pmJtGLhe3sAXt9jC/CMiERnMPfgjw5Q1pUofSgZz43CnLPlDdfz+UAW9hBEQko
fEQ/UnF6wyKsiRQP1TJL22ywFMTdnVWVb1rXq8SQuGKkYVQSUAHE4mqLEMS5p/YuFVA278XF54nz
lh2MCoy0RoiGe7E5pmQkmlrzFSiVET/jn8vQes7G+SRsvlCQsPWtwf//T95n7n4P+JyobJhbX0E6
A4XIk93PWPql+zsr92+e+lyQdBOlbXK5VTdwElyaHLaBKu3an9LJLmbJxFn2G44p4D6fyFIT8acP
gQPnibcHlHNO3jIG+hGWgnZJiCKl9/UeYfetYX9r2bv3btl4Tqrqqa/i5goDcqd7+mtSWvLs7aSh
H4gmTUQjFfY2fM/1wqrh0urxZ3lZBoDUHEegI4SEgig3+AnOJ3Q5zQ0YJ7Wu28PaMfuzUh6Z7lFd
8LPg8mUenJJxBNcEzAvD/8790LMk/f4MkfAKGVETMuuvwoqy/lV18eGdH6ql3zxCc8wdbAzonp6X
tiEnSKBNAa25YwfG+BwbahWNCiO5+BkA68QM+PwwUTn3CFxGa4fubwUr8N8liwC4X+ErKyjLIR2L
xz8gQxEw8jL/G2jVRrGBqLARBTnnJZUuYLPsdOrDx08rrs72ZnfbnQUsYspMdjYGj5zEmPEUufyU
gaFmWOd23WYU9/IqTTcbdM41qxLWvSQddSs7GrXiAqBf6MeCCo++/4W3C+3AERZzL3S0xMSgbKr0
3bGWm4tU3v/VYhczDYg2IB2Yz3Y8ea18svLR++LgWGAlbUpR1vWaF+zM8dv/42+tXpwUD2vxaz1P
0j9aoCpAE4lI6ozswd4e+5aqIlomiWD/BQdtVxpwjn0e9ixc329B2Fx141XGfbiz9m9QDJe+IUH4
goxG4uVLUmKgSNyYcknE0fTrJIrek74agZ0qnbLfbmRxGLMHXhATZUhI7r+J+vuwpqDQWMCEnTt1
NBHtDVso411f+LK00Z8H5W+WiCbuoOPnXsIv8jMQWGaXNZpTHvzgBjrGHZecno6yrggQxO5nTr6+
gxVrhF6q6XNmdeeZjL9bWbzbFGErCP0QbE4m4MFX2JK10jtuJgMQAUdNCJSLR4PMvSs5iOCZME8q
kWvYxWY7DNMg8odD22SiePRL09lz/BS2dGIqOmGEbuuo0WflEaXDFFaYSnn85YljYlxixflxh1oy
ywmw9PT8Ac6F70G6d/Kg5bDmTysrL9VKl/HK4yEPQVqIKQh/+HaYu3Zt7s+l2DgrIEhxgrkHzIz5
i21D1xE1cvxqQpLg36Ptu8dWx6SKayIIUz+9ZnL3jWpbjCse6x0YU2/9wTwud0nPwRDYi8ieXaZU
8/Gk/LGHlLuwUJzx24wzBUHFHTejSR0A60TZVscf7DGu6PbH8f3GOPl8/NZ5X1Q+/87fTcImlz/w
SbbwvcETj7MXZ6mtU6rH04hDzUUhmyxFfScqu89ZuQtg7S7tp533xI4d/r6yzzuxJ3vAWERy1hCZ
Tyio3yHc1VlNszBMGlo2d2n6Cxa3luoxCz1p9H0m4jfJUUss0FgsUnXAyfcU65JZBuaLdRcKs7NC
lZHsDF4yLd5NzytAshPSzT3y+JY0AvzTSN/qPuMCVl2GoVU+UfNyIBCIpf6hHdCPB9BhiVkZe/Sa
Ork0cs54q95Y6RmMLbx9DZr91UnbufeYTx7l3D/xG+LgtnBkmfcRIUEgk83fNED0b1eLRRfu7ctD
OXB9Yxy+da7ZfRg17Imw3pRPPsLjZQXwYsR2dJEd7fklAVCVNt/h6+GkShegEky4N4WAmp1kWguZ
spBYEPk1qEyOR9BRY55MJv+s4NG+B0jQxUJRHAJTX86DVdOkGpPZz6z0LbSFz8lDht8fs8zdyPW9
QlNOdy40iTWi+vWR5h6/nWWrxOGDIMXiW/b700caQeE8JDPcvneU9wBZD1+HbWZlBV1bz20M/pNX
aqmQMFQlD0rU0lqFCMYIto6tgVtEErEKcpLQl0w0Z47GrF+w8sCGqz7IcpiT4VE1xjHvZlKtmPB/
tQuGEVlgPnMmrKbZ9B2Q3reNKzDRSmH8sMfGIwmhFrlhRtdt1XmFObUm53saFMCQfeL6rDxGcRpd
hDEf4flFyabKRWno4HLJU6mSd6AdUuMUgmX8C2nxeDjLhyVSNJ//8l7ICBarHKx9xYi4BW/0TZiT
DHPmUD22uc+qOZDK+byCzLw7SoBTCGaD+AASc6NzDub6PNQL3SmIZOAFqX2RWhGKcndCbq6HX2Qv
I4zfnuZ4cqbkaG9w5a2H++1Pxw7iVeOr4dEqBnWRNw1fGeOaqHAyeDKP6wbOi//T8h9hfMYRMikQ
GsEz8ojP+3p6JxuvD1muW+PVmN12lLzZboClBlk6bst44Lw9uAmutLfNKDDGtFS82u321UfUZm5c
eAH3Ty3fVGSQwHYzp/cc4XyPYzmkcb0H458LBDkqIuq0Y5IZwfpFAfLisgfALi0U6R3Bl7TZNf/N
vURqyYOgElU7YAQLbCwUMQR2hc27JJF6++eqe7Xcxs0FFnkGOI4/Q8vpIFHJ5RaJMLXHIxl+zbfl
QzNagTyYu8pqRcPxdRLVxO/HqhRSzKCOUlBK/3mVffyCab36/Qr7jRYUcE32IVTw9zh7P6CbdWPZ
yrv3Mc8CSJppg5/3VWL4FVo9mjLBoGkcaQsgVRSpMMlZx/0JRy/n36EwakPL3pIZszC8ZMqMPnMS
mI5FNYxPeRHrdFRs3kitXdDnHEE7Vxbt6zhOQiy2OtV4PatV29nCtWzlby+QDBB1Wcck302lnG+i
r5ZBQPtGnUBzTSn+0zkN9D09SdvA+wZK4hb1WeWjz1wkLx9QZbyacYh5n8/FeoxO0CwmsHYLPNtv
vwWy4qOcR6QC5QtdFaY7Evr3aFy0g4frAhA5hb9KN19byR2fjYqv646HKro7HsvFSY0a+QMza7L1
bl4pfFerp39QUsiSzMdvpxaGS8U+flCiRV34N9eUZX3ilTPlQ/Nre7Qfk2zE08jzg+sm5XAVwsBi
eTP+K5VRajVyMomY7iTjYqZP4DIYpQQIbuhAJP7aTQvktSeMyiT5tp04UhdVsGJiG05Uymjkv7Qk
Vr6vHnfhUAHz77w4PYi+yoEvP7ALQDPz6iQowKDiU+AwuJPXymKwXRgfNRiiMMQ27GEJ2R8IRHhu
h80rcF8Hg/Gh4aYDdzY0Fu7NNvCMt2xAuQA19TAq7zpYEtYKhP+tlaaT4IYz8R4c8Xa38WJFhbhD
A0u62sJ8Wz3wBsn035pvHk9rDAnoc2Et/k88oGmzusePgJeiazVvCP83IwcjEznQ2S4aVd6zOWcZ
6JMuycnbU6PaQf1vVhxORVYMtV7J9LX6csxft69lyvS90KudC3sgSsceukUDjKcE/0Js3Z8aaqfI
QAOCUdBwsRtCOQd3dOjAzcEoxAGqvtxLf01ETLc8BkZXmEBbLqjhQ/3+1FN8yh1vLMCaqz2kDcL2
GaUui9yrclx8NPvqQShw6e4956qgPdP2X300yRTeu2ay9l0zkN2IJ1+E8RE0vwUJtcK00cKV3T6b
Vf/OF3yMzElFnJPMseKGryVzYak3D3HBjpQ7Q/viY6gJTCkepBonvrKtjasEAC2caoDNTMLv+S2Q
7QEHp8DMMBO8QDzQft8ctZkEA66bWQj5nzBahUadZAivGaF78iKoAbf/JsiYy5oiP/t5xOxozVkd
7mc4ZKWw+UeLJc0EuwEzveBDBfHbD0IzeAYfZOEwb2/Ub8txrU9/x1bYy8VsK0x3w4z+dcC4Sh9L
TaJPiXQgbfHffVEfk37vNsC8m0ThbbkOTDmw0G2pIQHyb7SGgVGbHN5CTZmAkSJjFF04MXvYQO0p
qOvhtIUtJIRax8Sn4XbcCIomIQ9bkrO0Od0y4cOE6+MgMo8zMAf9/nwT0gNNOfc0yftaN0wntVlz
8/WzZSR/FjcV71uqsXVqP8jME5FQeAhNn4n1D+SFubGJmdal9f9FnRgAq5xR5/OQqpMgVtFNUFLS
pDhjqHn19W0TthOT4TTxDgRc3aq4k1eH7uktERCWSUUl+adivCHxZck/+MS1/v/U/wdteH3tcH1V
e9cY+kFiTMXZY7y+dc+2SHkQlAOUE+5ChTwxbsJjj69jkpUh2PsMG+hybNdraNGTYvIbrfvrta1y
X5ITo4WzU3d9Cb7ktE76SRzPJ54vW5+vkaGBaoZVZypYlmAihg0U9qlJ6j2EvFhKkvKhrjwOMG2E
367XTGMK/r/zEch/B12R4BdYRLNsWi81Pet+IeZ/ld73qgrdDXAnzKbWrbPdWPFEifFT6BfOSoRI
grb7MWTvp0W+Yq1VWoFOD5plNb/QxubekHisDIKGD3sOIW2+WgKqvaZIWajk4rrkHWUXE7+jazxz
1Nqwca+G2uDahfDrsj+GPY1URSQSKU/5IdxaP+cr35+omxfHJFK7j7LqHyR/Dlr4Oo8ZVtQFd6UF
EFmjHePvOlYwAb+gxlsyLBx5egQyYwtCgsHJ0bmYrVwe0X67lbiEvCEqyMfrqKu1v8no79DtLcMC
apRpq1Opw3cZudIT546w4YOJIWi+dZlA3PER8lkDjfZLmLDtUiUXP0liwjHkaWDgVcCeTAD9PRLz
P98KBfHWyYMoLW9bFPW6nlG3e+X3n/F45Kt3GzqrjBp4S5+rG7T3y8PJs7OCeovqqHcP6XzgMHxN
0MswHYNzvsXKUTy5kBfqIOIwJ63Ohd7dzs9OvdKi5kek01wcr1h0OjvoF/dWjEkIm73sAJD/tfDw
QWHd05g4GT7v+7Rgsy9XW0ACKFeL2DuqURgiBw+Ky2kgIC5nEV2oiitdZJYLbGO3Q+dxuQU6dKeM
h4BBBAvpqQl+ykgUaI0qXzGRNHAB6d+ljBIef7BK8p1O9/i56bsio9lpbCPWnGVsHXMo/Pn/4Gge
6dBcQZqPm7VQbQF0zeS2Gxh2RFnzV2S3EFnvNe20WHtjIK3LAamryk94kPWu/CStb6mT5ubPDbCJ
04wAlORgOdHWKblnsH6UAUAN+49ZOezGSgxrI//91Zqc0QWIXm/MmLt3kIqJ4c8il1cc+0T+XppN
sNJqjn3o85ZSLzLvmDeUSCb5oe1dFYRrIz8DiZJBtDey5PWqjDanPImorqAhdwbGJc1hsXQ+IRCy
vPbeeS5FCuhZ6c355ufLhJu1XbrhF+nL7NDzJY8e/Bi7uib5u/DOXnaSISxySAShUrU5kNTvg8Y+
t9ADOPNf6QGAmJmdcHCD+E0IPf6CLNxY4YkGtgGX7aFw5itS63sJYjh/NASYuJBzYN3o2tXr275/
ghxUcJvAtELB27OoRLKaOByvdKn4zMu13qFSe//WG0wv/GS0MZ1APZ0sLazjBzP99EtgKHuiF8ci
pZxedkDnrmPjEFbDB9hV8dEWHOGiqmw9fLmQ2fT5Bp9S77drkLXfhsA0cpo6WtQfoF8N6mpFWRtS
T1SHoJgJEgF/kCzLpyb1x7UiYpiZsFgTWTb6WaU04PfM+AT1ltbzVFhhq8anbazbHE0EfS21VWBU
TEnfN2q/QiBLihCWWVC1qgK3/mjTf8bhCetxLS5sjXQda1IP4P1elXDCIHvnx/EX3dt/2fn7dGWg
LakEMHT763KpsHZWKHGDPiXK0ftetrfr2T5LhrTH2akpbRtdL4R/QUytcJ52/Bjo6gbNiz9Kn9Em
8jEVscibHSIlZOqOYOobCw9TKKVD3oO6a1BfmVdm7ljuFQ0DceOGDF+RQqbM8njrkIAAzQRQEDK4
IJvsiF4UiySKn8DBpQ/ZgTvLVpg7bs108pHjLXUAo9zj0dAm/z5NjyvLK1qHerAFy0kAJdaJp/Vl
uAjcyKS/2QXBFwFMF4C+XD+vuHBA8mkY4YJADH5Oc4moSqzl07C+W6MydsHr1VHHhSa9wM3MVWVQ
VydFGLlMwY89PbWvIwiof+jROqz/eHkFfBcX1B7RuV0oH8BxJ2cdKshC6QoYHMhZW5G5Y3ehKzTi
h4EIdxdRfpWpO+9qNUVwuANOjWBhBTApHQGpInOTkPUSOB2Jmweb84RZ0ZJU/CLat27Jm7SvUXvI
2GOCMBBvtNn4ZMVPYrNZOfVBZTwLOF6yZxtk2m2ZwzMgk4ieXM9BRoVKkF4wwfp4UsLM7rx3/C9p
fxiVKXE/DSpJ9T01PuhmhFEvj7IxWPKDkRvmv2jlwJl6c6K0J7x5U9bORcad+pmpZkrPep3xxC6C
fmPUjRCrWDN1X6db3d+V16s1pTNH93PeTjfGPt88E3cT3DkvqQMyBTWpMnZ3/x9U+cqbG+xpU9b/
v/4w8ALqPSM7C9qmB2ZDIIGOJcpsC1AjE2HD6bvXHhZsOTxaMBPez83+WQ+l5JaCFZfn8wzD/L+8
3xjlnNEnIqNd0tIjbBFp+pIVMBPdI4vp92QsTHBHzJI/OpDEysyS7yh4PaoKskczOul7e+1tLDXR
k5yCqDP09wxULays5LXLSKYuxEGSe6/M8nN8Z6mvXxas7zkRITk7m7+/ynIfzE+MY7Q6T7we3rOI
Euex6qSqWLzU9v+9nNSAlVXVfNHccRqATTC/tz3x4wXs/RetB9U97uIHrm9lVgP8Ssp+CZS6ivuG
yg/K6k7D3wu3SDd6csnr5mVy5uCRQau64R2jflys1THDEQMddXrq8FmjH3RLvgrCJC/YFF3TvNz9
FBU+rQ54t6xL/TmsrGZdv9CBvgV/OGTtKaqAZxNTk13lFNT/7FkEAl43nP4l5kGLpDOwajEqvujw
dHQdQRYWXObzd5BPrpxHbglEalQ0was17GgQdMI+4B8tMsCOZC3uaNpcsusccULHw31b6C3hwlkB
sMVTOUoOumE/ZCNykrM+cGOtq3atCHdU2gAyPHAMFPzUt4SVQjPCT76Y7g4atj6k8jjBA6+1ez4z
5l0aDfHEkgpau1F86Hm5zYKP5F3mG7sJK09Z9vT65FO19XB8+dtpAHuxrMNGWCaulHsPwdNRxIAT
EmH/ooP7PswRq9bLdGCMV6kUUetusC3TQj0Kh4QafbatC+NYv+I20xkUF/+bho/ZuwworAaJsu6K
NpiUP3JmbrZMcAzy2nXWSObFzyjlW3jw8HYdJ/k4XtceSMDmtkYrTjhJBye/IwZFBAJM+PovLWOX
Bzvr9HkRpYgXugm3aeAikm7qWzCG6JhSIMjNhpC/f3yGcPIgcfKI282+s9z0v8+Oj49DAJ4KDmph
3KY9YrTaJ2nhgbkXtsl4ppGCIh2bkWclfeIhaiBsmJQAyWL1YjJnzTk4BuoozVauiObJsRpyfMzP
/oWe2wHJFn73wTyW8lA1qs0DTgcEh7Cb7UaEimZFyeRVwV54eY248UWCZ2hoR3DPSFL/liRHPDfc
63vLHH2PUzgCypygFArzTbksWtdW3W+UIzn5NrQhx2DxsXwa1nirB7M1hasBueEm5wiSddPhH4ud
YM1S/6qJ2N/M1TFaLn8aP4i3ZsMDBmwSE+jnfIL0Wl5Ae/qgtK1DE1ntz966D/2Mfhx8gmNRsJWU
HOkT7s1T9mgupAOYa/7V4eRmLjLFcGWP6Y2iSiXnp3ZkZavjU1P9ECYKiYt6q1Z+RV6+w9iU0xFi
wZXjiPQQC42OkzUyLWL5lPPxt/T3CLqdLs9H1T4a8vIzTzWqnVD57RwWCqUzPVJPhbZrePAcbKCV
2jf7OvxVxgaPpw7urgwhQuZkrHCQ8B0JyEl5e+omPbN1PnzhdJh2WXmVnqUJ+/GYwXMs8bo+WCtn
Re1mjrg3beCY5Si8l8lksO6OUqVuuhvhhU6FmLfUwKQdtYU/zsi+KBc9dTNi6W5alv5GhnHLBB3j
ymh1BrqxO1XoZ5t7xQw+ntbbOrwFeZemRMayo5gKxRroZYQo+dnxQyAQfr2ctXbbpW8ujPHtBAuj
CABM5uzhBwhOUpft73wkFPkBWDDgQpfzvXWiErrSc7WE94EfmanuuHT93+MXkmBVFnyu0R93uBjv
lL6SWHMdCqzZgWtlf80ufGIHiL92M8g1xd7B48GRuoionOKyPG1Pa2uGvsrsw+r5krgZJWARy3Cw
DIh/+8BCrpPQQYc8wCwMW41YG4m3FOO89+bo1FIssiBysBGaAVXKJAlIoLnmN7BSTbZYjDfVSeas
rkKmjgu67fuyleekxeUhL4f2VTf0fuOxIKvy3uqm0tFzPRBwax03gRVYnMPTgVk+XMlwNfopN5oc
yj6ZQEjAvUWLQAnV2Qvu8L14DWg0PsoXF/In6bUwe+UGiAClzoyAWHCWPHKKbHOEV2aO7G7ngzEk
YJxWMuv6Xk3x7da8Heu6nUoVSDJ0qYpSwlRE5NDUYJFnSEu8QMA95ba/wzTifxgt+HeaeL4zAddq
P0ML7oGqSWeb0G9e2uUxcN9WAdCM/27WSAlMAdumI6xpWERxR9SmMSfAG01Qv4on+B0GsMNwhKiy
oy32rc0F6IXcQA1YQt2bfHUnUNmmyntHtV7sbu+Mi+d66wVzki10s8jFzzhY4HK0r7DtT7I7xOic
ydSLp6T47XXFEXvDqFTMBoehXhCEh2f6qavzD2hGjHY40bsbZmHIU/5FXzs4sJGMk1CbWQ+vUaa4
7yNGbCDSu1yIuNJ37pk7QlLSfgRUiVc5sd+HZmB1ViFL29+jTqqep1YlGNimXi+vRv0BAR6RFtCI
VTB7kOSgVlMOflHyy1wsIhZVUf/ev2q0lUPvtTinwR2pdbs410P5N4n+wq72yK4bQGvb2sdaVZUg
jJXQYb/HE2AC3ye1U3TK1MBWalA83C1m+79sQenI55H6cpEV4iQhit0viO/k+OCREsFSbKMM4hVo
UU3BMjISycphiW6rJK+hysAVr0evNPfAnxFOCTGXx0Qxf5ZgUiWvYVTnGoBn+YH0hF0W8bZMJDYf
Vv+v6gNgAmHihacI5Sn50xpAurEE4Rk2K0lHibs3J4YAPiLbkJqTpDGJGgHNMfiKU4ii1XmEBlg6
AnL850880CZnsaytvOX6VJKHwJwHbjB9REeCZwvyqvTjMCj0axOOeC43TsjFhSg16y/wLAR8Kt5z
+qCkE/w1pRtbe4/DOAzK3MNH7BSOfINx9u/VKAujGspsDjF4BxPY3fmsHJcQcPoAyCj9Vy3K+eCL
Bi1AmhjVs11pG1L/iA7h2qikb/CimLNJBPBVk6fAFWaa2YE5nI2D4n07lbXcXwymlj1IF7zyjDXS
10WyluCdBDtKRHdy86YTRTI+mCtmytMaSiygR5aoGrO1T3APJfvRA8Mk7QnN+8lUoCspW/UrHd1M
HAX/Wt/Idfjr5efjZfvNg64OAFBqjVla7YR+HyQp2F/61wjn0c6AjQaeBs2LoGTFLwkTi4w4xihU
TLAsOJSphhhePrRSk9QIkGT2bc2cT4GzShnG2FWJ4ybhJizc6RCv68HD6GsFSZPDAM9wLLuzrsig
4ttUjduyixxNCq+uJep/wZLkhzt1tMR2VUfVuOITvByJmJxHS8lXEIq2Se7lY8LDIkCb2+6xopub
V/APM+rcxJQF8avKDHoeIXz2yu0EJfy2Uqk+dshLoNxM/hz9JEZCg1kIhvh92b54B2/rAHQgVESy
egmqsRi0QdKsQOZV1JIG0eBwGSUBxxJ+FVe4zVu2E14ShpUhbsrKVJ4ol/QaFFBo8iBDId+ZqgeK
3tjotMJz+kj6dyyBoMAfyr72ZOpOz5BW3mQzN4LJ8q9kiDu+fWSEnMpO5nW6cgga1uPThgmyRBOX
G7b9f76nhMuxzHhTKkQdQtsxkPiSb7praCQuHEt5CMSllrhcrl/PfN0CP0SLtaCl1bwxL9gEMwCQ
I2UeHICMKy3Q5lEIU70BmswkDnrimO1GpzdgpslfrRqvNzajSyuAUTyZw1WVGQeJlwvi5JkTLX5X
/xS+LjdtOpwsHL7MZSC/7Tb8pnkXlUoXS8FqrYHJiy5gXbr/yHR4eflfu9exETbYfUUoFsvUop+s
eGwXgVQQ5fH1stMB2UzqYi3bPoYFRtTm7n3/OUGcClePiXpI0w1HNyi75oXMvA3Qght4lTyWUV90
su0UiSocKlNGXjBfoQu3Ey9T1W+d6hPk3hdUE81Otzt3AwYYHeSoSBTjQhHRc6ggZMV4Icst2J/x
c6ElZcbYITjKYYuRWzlaItgap807aoh7ocyf16OhU3UqCnBtILf9gsYpdn+jo6pRFTESk2zBWYU4
C3JChrR3s2tbFkGjemEhfMj7PVoYq8W78xygB87/hbipaPeZJ2FDu6nAR9d+k5qMLd7MhO4Eq36j
eJyOV++vU+DL6WrzafoJAqe3+E/eEYFRbZ3eawK9mishi3NZ2uvFPVYcVkz7bvcEhRq6f77rKyHu
b3CF0Q6J2GQx3U/IsB1z0a5vVx2ZopGbcdUVVdzOZOC5grTnoh+2U/g/lANj3SpMtezmpYdvGdlO
vZWRAsaOJ4b9Du1mApIvZXnqTqeZB7x7P6M1fQrt9T/erWGJhLMTyJFsod52UCH54cMx9T5OIX+M
DBQYZQkgAM5ILsU8lvL9GJzlCZkXwtUXvwdGG0+YA276TvRPYZdooPEUsqba2X3+QcvlWRQ/GW6K
E+tCgxTribZOOhVSNnDc/FKdrzDMYIeC+CpaqtwafRcROQuEaPkmWKI5rvwC73Vkm7G7Gdxq0io8
F4A7dRU79sH9CXRVV2ot6y73bPErqd+dzlg/kD7Y0G/sUtx60mA4QWLU8HumsXclSUdo9XVM+Mpo
F8qzWJRHPRvH8YALCfnFW7TIVI+4TI0SBSuWmrvQfw4EetFzpJR0h9lx57+6EniDcMH3zF56kiZC
xdAVBauEHCBXIIOWhpv6YKs9fjmOnr1ki+R4Hog9p5Zdmdi7/E98IcEhwKLYlWP2PDuvuCcvdWmJ
mbGPLEQAm4Upo/AHa4/hC1B8iJ/ry0Zc7gxUaVjWOZTDJO+Mp0jc7Ay4b9BqoTvbZlO/tmDV1Mkq
lVhYq7czc6dzZPuxevoYVZtt9XhEUt2S5Atu4mtP9ukQyWfjyHfiRdD28RTrvw01or5XloNAIxc4
hzObrrO1YYBfGRv6T54c//kEnv2jRhP4ghbB9pEPTSaYRjUppGKLbMr/fIx5DGIpFMyo7YGDebri
q9voTbrGlmELhBcVxtkvjtF5AsjTV2en3lAacEk7rDw9VQ+uq2yqXD1UM7KqigSnes++ufY+vg9b
hylx0lyRTtXEuQjhVcS+yxE/aG/MmhPyH+5YiNgxWMfSV+5G53FpGvTk8rZqkoWznXLbzpLEZy8S
yhlXHC0QtxmXjP20/ZlD/wmRBYdFecLynK2Qkfxn3Csl/5k8JQIChBgfKF3vxOQC0wL0k7XkdS7b
RjJ6o1gcRZK4W+1JLKdH4Bsy+LlBdxmUi5/htEEE2sQEwkJYHMxU2DlwFigkEPi4DNGhwAAruPCu
EQfh/FKng3D034iHBVgDqwhHIuyFzSPTKQybcsR+vy7wulw/3v44Q5PDWWJ5hc010/rf212fMKkB
jTbMy3iQct1aYvRbPTQaWlUBNIcol+v2Ug44UW4T5U8FxS/T2Q7x4S5c3oypjNLKKcCbn15KVhwX
nprck8C+6m8V6o0S85Jd8Rjfbw7Uh5kaC3HL2qUqZH8ZXUhIHvkvP1dc9OjfZHoSFvv2Iex0bpmd
dk6y4q3ec44VxHquBze138dgk8E+W6SmmxRRmiNMWKVpmyl+L832k8eCmmxFrwYelbLqDWsGn8e4
YwXh6C7pKQQPP3xkFsMNm4jmeaOK9VdNpxEoapNuOw0JMP0IC+uCy8Z8B2n9D4kfG9isJPpQHY7Q
tcwa7KyLrLnsTQTo6Y1j5DPcQHLnQEpTi/QNuR7gAGIF6wCnX3L6HX6zy8NUY3KM7mwGum5CXvVS
WUUVKmXcqnIVi5wv2Oe+L96aLJ9wCF4bqHvgYaXloDYhKzZIsGNlRmis+ZjzUAwca+lDA3S9SEH0
6NRSG7FzvbZNUYzLXpnXHp+m2D8FRD5C/HivDoADAf22kqPUUUr7y+6A+G8iMEKoGqQv2jtnV/Om
+zosmWfUuJRXBpNiaa4X8dTPXSTXHeoIGivp2BBT/yNxfzBxJVRs5KrJofWi4lD9jQyJaHJF9BqM
b6iz2GE0vi/k/hSrKqk508e21rOaVG8ERsJghNZ+pJWMKPTx9InwIZpexYFYWUObQsKDylaMjxfl
CSjUlRFqzfikDqcaDx+hhAPbMjIF2tiudsi3hACIl/H8vqASrBe2kg1OVcpAC+l8SSDSOleIO/ND
0Tz8gLmWfn/mgbXwEGVbEWHY2/duwxLdcWAvHp0wgEfWGVdjaS6cfhO3J7gptMF6KQOIw2JrjJcH
RGvCTDBhnVqzFzHMikORD9pGdm+TJ0auVfwBppIpQDlUt4BOUeh5pNtXQUeBERVLdDEOSeXwtg8Y
PAk3Os5TwcsbGZDEjNBVNGu/jSKGEG+LUBCQWB+8hwR4icApnEJDPPviGgmOMBdmEL+4wSpfSvxw
6TKRvoGVLEY0r3VSHUvh8a7Vn4y8JnXAgeBSSAUWTKz+WZEiobFd7IwsbDClLnvYn8Bj+mPJvf0e
N7pK70fcTFWAz98z9D836gjOrS4LlFvN/0BcBF5hPkMvyiFJb6m3Z7oFRLeyWlpeflJ6Cw5w8K4T
h69j0yL3SXh9qRg6Y8GK1LWno/FH1PJRyeEKOXDpwE0AThlHrImISTZEQ0OAn70Uxq/Qpoe8rWRv
XXJwewnRw3kMaLxUmtzhFNwVkzaWxeuxofreTRup8DMe4af30d2CYBNGEHpg7XJljmoxlfN6ZFwy
ZXYKwC4E3RZyKlUnOcxQo2Suprba8WxXPmXrWkzT6U5PtGm6XfoWDolbN2ZNR2OUdTpLxFvY2Xfw
DfdIZcaedszs6SeucxrvkUSYkBdRMWQFn/2o3J961XUIIQK8X26ZlFWOdiSBRAwlsfZaYuAjx80P
xhnfhlkHca1GitP2eCHkMCTHWduFsGov6iNpd7dDcFnePS384PbWazKvRtpM4DZ90TdRiel3ZFCU
fmiknCHNMa7MwhOdTkcYcHn7fFZMwbk0Mb8QBRpdqoQFEfSgArEvpRNhdEPTmXwvfjkCB0Fts/kZ
jxZJylvBtVQ3SRCb629m30dZ4PWPSZXHd6zUaR8Vk8ZlP0j+QnX+gngO5IkCPwmeJI8s1VK8A1CP
iAGPcGqvnvlazCdApA+1eryG3t3Aw19LeR+fEpDViBgqcBj17e/RyqHehXewgSk5gLQWJPQJblY+
6i10SF16RKzkY2mw0o+cPZeiC+DP8oeyz5c78DiFb3cKWacPBnG9O/+iBSmuLx4iLTzJomE6fIzg
/bWTFFeG+Zgntjo68yZUIpqux+AHSlvPxQ50FCOS0ityYrUkUf63V5oLhdpsNZfjxzangL0kLi0h
t28qW3b9eGHumV9Lsh7io/L+I3/YsqrsLZ8GwsLDS8rspVpOVAo58aTLLUn9T9Gh+OZglDG7rgpa
Nt3YN35kuaQ+OYL5oew6p1Gsclra+tFPfM+Yyh0LddGlYxVW28Ee1BibA6DqGBuQ/GsqiPIH7aeI
MLdxwzp3hnHwXQqVVwU8MowoY2N2qXbYbuQ3mB8HvmBklCalb7HcEjXFQNAiVR7dj42W79X5E9D+
bsLcX03o94H08goiuviMbPYadHiqbkS28V/B3fXA8JmKg8huSSeL6zJLqa5Q7RTL5o7pXfipIKjU
lCLDnbrQ4Sm2vjae8ZtLOZ0PBHXkH04Wnh5myTI44Y5xVEICrmoF8a6E9MRnZ5grvDN7iXqhD7fi
2P8/72SNVpONjg3pgFYudRPPGbCEyiphOhamd1BvuCwphjgiXOPq/Ryq01b0YluQae+BH/LEGGdr
RtckcCFyPM61JmdUw8gXduicPworB65KhVgAc+hN6+HnHt1iT8m9pmD0aUu+gz0IfRzVmYvAeCmB
35ORf21mEPWFeieBYYM8jjhh0BOLa+6dU1K+eCDUXvNyCVp1KD857hI0NNT3D7rvnvIYUET6DuQC
zTmXkCWB92HyF+5km7hvJ6tXwM7sr9zGXOMEKPwyJXFNnr0TvykRcSXhVA1fnQP3fOZ+gZRh/Eo2
0ea/vJbQ85Lwx56yXEsI5WRGEkOSTFqVrm4YJ15JjIPjuYIqCDbnGrFG8EKoBj2TI8/QjqckdmX3
xwD7rfEcxSO1ZA9Rpd6hYpY+ggYqJZccV32aDMXQx2J8k91H++rhAWxqVJMRLOk2ho6xTadYioH/
Nk38azBAghuIj38UD2H74phoqr2JpCOZMHwUMZmw/DzV/RoepRReyIv9BBHYTXXRrMuB43v5sS5D
FTrNtS2N6kgKrtGWMof96DR9W0Q8mXQakVszpFjLtWXjK0C2ejTzFRKAmi+GW+lMymGrQIQM9HmR
l9Y+Ts7+b8sQ0EuE1kY9sl+Ua/FnB++u1Xf0CFQB9ApDVMwNQ+8QYLkTxMMeI9X+g8vxkyzVOgdD
m2eQU7lpAkX0T+vtxbtPEzAUap0/IenRC9t2ZfyUQSEcmlDnFMdpak8j9UkR0l5zdyzsrt501/1q
3xRaMmIf0ru1L8CDErV9vQEbxjYZ7UgTtlw9tFRB/29GNNVNbdgDn8LtfKnz+M664SuGUxDwld/e
nH0kbzLLVHTbuBE1+lAK+eI5zNcfY7RPXKOqqWUQV2fR16RDTdegne1sr6DvWWefGRvOtfigtcsp
TtURylt1VbogoIXRQKkaE9plvQln8yh3JsnoDucaVRi9Fx/JElOSJcSrRd9voOVDO47I72g6YcRR
7MpS84bDWu7rbqYjrdIx138KY1xHyKgEMiS77GPVDMpuM9bZpNcDAlSk8fndXGDNXqGXRhuygXc4
UHq5F42rnH+jBUulJ3UDFM2oiPSKsj3VYQkhovvIMBmA2P1UMI0KholKvj86C1BTUrqEOShwaI25
kkbOQyN6563+9KhCXsZE6fsstJgz4zO1TRcz44Gy5YSlCHWtUg08zLpNGp4HK5hYTwD3UJJLL+yI
0lh0aZdkQwhK9SzdK3kyF+XDnKQ11lIDKcj1fvHSh3HkSNRijWl2wB8M2gisEZm9FRWCYPL/K2GF
sGAQzNZxfkFX2jkqh7u81sPt1+trn6d9a29wLq9PRsM03hSPKURuVSgg9/yZiZy5oarQr58EGYW/
18aPoE3oVE8+CxzaCYtEODpMuL6eW2oepnHtkv5zgi6BCP3C1fnDR/bcZvzZkuSsYroXrFJGKKiI
CHTW5arF30upzeeCC6N08YZBbkh6DjfKIthI6TI5BTsFMObpbJw3eozMzrwwBOygqOBHKc9kLRqh
MjKf/8Owz0E0tazz6tQ9z7dDAu9FVoWaMbQFCOEYNtex3NW9wkHlUKtFrUfYP3a60LP1Zx4ZJrxW
xQum92mznsqiNVGYShUjIAIewgqG1RK5pDYDcaD0baH9lxi0Xk+GWh0GzD1OjIBwC0ttkueUdcDl
jrWmrZ4H93qS79qI92n3UycHkioPPfUM7soNtBaIBfV8/yAlNLgbw7C02As8epmOEEigTDrLN/1L
Oo/H0C7t4eOd9+lr7xrc3xdEWVK8vEwANZ9yQK1DwiGcCTu+H6m8MvOfgO2oGFoeyzvzqHzHAsIO
hEPfljL86NCZylOAPDNjkqHZnKl9LCIyRG8V8ugF1ytKh489nH+LICYn4BIw++46bnoa39SUjEyJ
ehCWk86qOrM8n7O2SXMAQJBWBi2qdNDgJHb3hBUME5wG9cVlWp4cGcbdW/wdJkPLtT9U4DRNjp4o
pyz71ZNoD8i0XnL/ZzCjHh1eodh3n2OaBXKBAk1bJMPuoE08NncAShz9Aa7cK1hRxyo3ay12R2PK
yg43lpq1FLUqWVtXsw5ZhNF7ILRTLmwDOlaHzGerLiEdha3oZf8pJo7imvgeRiMmOvIFl2HNLyVX
s2K2xlcwk04a31UTDPvrnb05+OrkROV7RYbDo/5BVEo4SHvWJilKxiof1UAA7Vda7vjzNbHYIpd0
++Dz+7mhxsQ9vXIOboE/RJpJbbpWizoFNz5b4az7MbXn3i7oPp8GBwOzhzvaL0njmFYUxcUmFlwq
q9Azl1o4KDYmU3lS53HWByiX1bxrJJMkkvG0g49a+2ZYrB5ORDrQcw4G9EpsG5ub0paH1hePufAg
OSsD/fwLg2lTefkDel6GuMepRq3AYaHh4YJbHQ9vsfpiwyjPKv2/yPQWTjfsrrkwxQfouOUCf+8V
N5FXOp6HXDmeSOywzqKeTv5wYwgu0/2hSnXXP2xcsI3ziuQ4+JJ9Bd905PtppT0VbPic6mcgYv/8
efssPvvoQwhdUYTprKiRKYJ/+cyCDLadGGt4ugWIhB1jMRa6FIcZTD5mmzTyW6wcxZLLDvHioJE1
KXhepgTmsYNFqnjOfPzanYcpgeDQO0gvTSiJUqMeRYkIyZQbhQaGNAwzNt4QdHZNOF5VqYyxHuIw
A8kIrPbS6w1gvDGnV7Nt/zcZCA8F4NHMM4k0koosUwg7+ffE1Cz/8grlS5lw2kcr2S5oQO43Uu3J
yLV7fk1un39r88fH7E+TzmO9yYcFbTUN4OuEewBmGzDESVygGcRYO6Oh0tBUDpKkQ/0T6wc0n4bM
yt81RlXku2vYynjwak/EzgT/b7OFrkGtxgefmPiJh3U8Lihl+umILis32y1HgzM9oHSqFGxeS0RD
8uqdU6o5OdXFfoOM8CZs2aziskk5KUeoDhqRtkpyfMD5sy8FN0fcT75sDXgEMt9/v6rX4PE32i+4
ebQ2jCea4T1sdN7qab3LI8ImX1wt2zSfF1XvAarQxdOWAQkTFXxadychsn7wvP3O1nYaduHqjDrf
O1QIBfGLCmXYzn+dKEbRT9EvpkUJRv7nSC9i9HwZ7QFbAgJnPvTItAT41oTOTjlYT65L1jaJiaZF
qGz68nkYqy4AZP2zChjPdtCMIpaunqHWOoTP+5u8jagOothOo0VRyCHS1TFyj/rArXVF150bmoVS
DhWB7VwtSQRXWc4PJm2BOM2iAHLKHJAA4oNZZ44UcP7YiObFDbxBAkhiz1L743uaoocf7tjuse9c
O4H/O68NW0odIzhKYKgDIpniTUDX81Sl7UuU83x0RlFTVg9vkChYphUoavezZT4g9ub2xZchSco2
JYxStWtz8/8oiO6H+PBxLctkNpiS2wq5wg13WouVmtrhfxpWa2p8JS1TRx9ydOStuHhKobAZaplp
F5TKgalbC8TeifQECFd54nWZtSFbBbOygBXnh/rfx0cM5/399QT+u0F83ABy/yuMB46hCfGwR6Sa
aGyrXQagUJTKgUlbzEub0X/2eXOVQaT7vSCTZWExNGlPupnoNtkp+LFP9Lac4pLgtcANwMGfg/Ym
8UGDZQVDvZVG9g39saehy0RLyeWIQl/7K5fGUpu6gKOv8f2u1Uyu4N/USOcO8qbVDwCvfrxYPVJF
zgmSI7T9zUandbbu6jzQRwr/b1EkJHwmNMFHFnwLMd7+4dFWm70/47MjGeN/VapYfJL/u/lTM41x
WcAg5ksjDE7zfnAWTQPcPxCR8LeA7Lu8333PVwD/2Nm+kkiy4sJ3wwPY+HDg5Aj4h92zzPfbq4Dz
mmsk7JPHaS598XPWvIsz++k5z8QRf0hBD6eMKdoctSZ5k7wQeHGJXVMz/c76UO2A8j+mbEGJVbNY
qPS5Df9nmGEvO/7a5SafnIvxjVorsamKtULUmL1DB1dQGqPvuSX3Ejpq5WLqZudZTR7cmRhd0Lyr
X66BfZLGiSdCKsyyl7XdblRW6zCWbJoSD5voENYh8lKgq6Btq9elFLeoRJsCml4xxMWYtYyheQPT
I5aOrg+Tl6ClNx+YbnGtoH/dVsA4RaDk7CM0pvNvQBT84UsJELyu0GS3UGFAwx/BtyMnk8sb4AhR
EpBWa6l9QNWtpp5zLrux0P9m5dydtYA++Kb7n71FhdeB5VlLOmNokwQv6RZ4QXFkH0n9SdCmjWCk
9iXP2kx3FVoYWQYHaEkcjgiq27yBLwxH7BeSXvuaQtfzTQs2YKR7Ch097Y2qJsCPn9GietflIbkd
aVQU18iEGhWzdryg2CspPe9lxq/c1Z60p4/pQsvyY8kd2xXlHnFyK/e0SWVOYiqIoU4T3HN613uC
jH+WEFB6mw4HW+QiufJENHmc+lhxMjSo8DRomHK8dIQdck3TN6rniwEamzenoNqQqiO36h4XiIRS
kpzMTXxWD2uOYlo8himua+k4jX7hq38HIiSJPNrC0MjHXtE71OSV+5kMiuzhqWUwU1qFTlhIMjq4
UzxOwMNbhSrev6et1A6/cNSbQftnC/QO+R1ssrez7ZtRTyc/0mB2CpXfg8Muo8D1yoicB2twnBpk
FNi/YwGuDVY2kLhDbGSXIJJDhny5dxlMAFeIqI19MGe/mePiEGiqIZWH2DjPoS/d5VrSSUPRJlhq
JNbPrAADohpiRkNfSXZJUS6luJzO55xJvPmFNoykszl3c+zFqyfPcUFIGKbCCKXUmFF8Demd4S64
7LWVYmFocyxSwmYHzh++dT2kF0IoSoRpg9TYdeAfj2H6HD31b2HtvsZpw3x5jLrhWhTSlKmD1VA5
eAMsFdKa7fVuzBUfUCNADxoCZMDZM6UPlpa9ang+L+ostJxVI2OUQE3Y4YAoYlnb+ZhJw1JYqSAZ
yOiqy96R0b+oNl0B86ccl9AZi4/GvkYGQAjQ0yjLwOLsjXjCg5lE1j+PCkF0wVg22TmQpJgqGe1f
1bhHdExrOxHyJ8xqF5/LwlFpBLh5ZrvFw+b7efy6TjFiHKKnxQMRf6LeA/24Ni/iiE4PDARoSM49
v6rS2RqN7U8q3tjLze9HDAru0iDP7OjcrLKAZ8Ym1srBzYytH5NOVbGfncJ/LvNNotL8pm58U/Rd
r6JsHDSUfwhLmFuRgZxZrdXPOvmIxeJ/wYEyNT+SiIYdrS/u2AUNh8BDY0UP0gIc4/JOyCTgiDi+
G7vr4Q9vX2teN3WEq4CnFBvOa7nyeHRRUj+KP1HF0Pt1nFlFxon9Um9UosXPFoizIqWjIXTR/Ssl
OjjXdigqUX+02h7y1c2EK65tbsmL2h3Q+GOiDz9G9wic+CsHU9i1WYuMhA51di7OGIXo1Muf+B0r
hrbU/9CGbTcVxIpYuRO/VvNQWjer2ZOC15mkybxY+XWZbgHXDqs1IdJONa3h0dbetO+lxTtGYEqi
uVffoahV9vIqlm4rp1hSQYdPngVDzbjWZW6Ix7kpttadcyIZ248RtXP0RA+vHbDY78zAZi8KScOt
Jc3DHKIAFSXsX4e82tvgzhGCE7/sR7MIra2bi+7ufV/0hWhGGXipaAI6SO7QOeXpsailgcReOjZI
BD41vOBrap4740YmDw4FkJGMn12Gu+ZASYmtN7+yJxjmQ4N5chzST8cAV/ew3iDGsIO7sCKWD4rV
mubqqJYR5VttkxuNnqdJPfAJKXV143ECe79Bvc1g/f/NiRQmdkaGetvN5o7X8opM0dTSfS9yW0cZ
BQ9DP4d8Yrp4Eevaf9TISJ0t+CjLh2h8a6RKcOAP0/NtIMA0SvcmVIh2QM8fV6natOWX/cjsdAh4
nP3z1sxTWvli7Xkyuqj2woYFlQFdhf1MM52ErSo2OPQVk3H7pZ5OhBHB4ZgEhzYt1OFY810PXAw4
noeLR2g3wX67Bj57OZnrBIw8mwT1gm/b0//m6EFtrUqDUNyvYWmdBtCuoZ0LNcuRH4wdc1cNFBpL
TnsC8+QJmuaUYyzDCEUOKEQysv2d/wTqEJ3vec6QKU3Rfm5jaGoHDLGPCunt3Ks7uC4opfQtGLvZ
WlqZamVmo1fKixTS1yLvNVEZeOOzt4zmwABp5MMzrteID0zDhpaNepRCHULK+uDDDYjgWqeP4tkK
in/geFXtn3Dz8A7zDlUav/VkP44/oGig7mKJ5mrcLrdI63MeyVpNVV1IBpk96ueqt5lSaY9tgNf6
dn1+nn58jA7OcbyCZkcoB8iAynUsLMrTkZSujL691rh57rn7cEZFt/glrZcLuUstNN+H9RmhLyqd
+i1euC0+zn+ZMPxzNagBjqpgHmwGk4Qcr49CbVXXCX+Xmw6PZrLcIznLYbgWWDUbHsdLTqg6HNcE
RmfbxzVdm/jDENEmUNfBgCorBmWmNI+IDsTI5KPR466fZzrhCwi5lp8O9vpSu/SD5gGMjoSvSglG
+6EHShXLheLb9xqg5qk6GSYt+JwML9u5dXZDo6DkDNAEe9bSZGYhmD/Tb/NkxsLZpSc7qu4v3Tfb
GGMhCgJmHxp2mBkclG5+lX4QN8N4nW5MCm56WBjNjF2dtSR3YlQVuVxtKorzp4BjtpJ74T08mLWi
Xx9iKwJoM42Pucks3o7dTKfNlODs3ZdQDskRT917jJymeFJgTEdvetHNB6cIp8gDXXGhRYPntA68
k4S0cF75DvWRHxi5fTK6ki1MRpVTPPuh6qAz3SLacJiH2gX3NNLGvbNLDKjBpDZq1zTABj13P0R+
tAKpM9Esm76EB/cH1KmVnfGlRBeqE1RF3a6vLLkM3na9WVNiUcNT34KqSHOSs71mDCMysMk3Bp1g
jRGXlRgpYDQrprXs138ZQ5rtTPMQlTA4KK/SPjzeeD/oR0waxOgAgI4uHvDobSJL1XqCT3rcB5L3
7CTrYlc5P95Abm2955vUDXWH5Gc2kLz2tADRs3W4uKFE9VtwK5g62NOhredbR0Te19S0B54nuV1T
GCU7S79keogrRygN4WvFcUZp7L5AOef39+meK7vYMc4gH1BM77hjPQz//nywBYTYLM7uFSKxuetq
iP+YH8xrGi30hxpdLMmAM4SEyGywjFI8iMgR5ppAZywNqLN83dxY67UgLe9fZ4sIfu8y3i4Dx9oP
miZ7KSBO8W6aezrESTmkkG1T6bR2RXzFE+dijJebTzKU1Fkt3FOTwIddBX8u4iSbJMGHFy4fz2ML
+2ru3CwytG4l89MXw3W1jPixLACfudQaKJeO2//2CRfxN8ijaWstULocyMZirEJltg7GhcH8LY0g
0M3NXUSUMva8eLN09FD8qSvCwBgEVu9nhpd6y3jhiAFVx3a32QQ7jvf2Uj9pXnPIGtRwuNSbr30E
S1clFEECHmZy9IFBt6d3ESIzwD4SLQhomK7QIrijfKrhq5aEAm07TI2XkNEphSJlBetRbryFBRwh
jddIoosO5Lnl2MMTVhzNB7qrKX0iP//oZEqrBR3+4Z2U91sW1NJylNKfGaAe+xTJl8yx/3ua4l+m
sHkAtzF+z/EYPHjl7+Lucx0prTJl4AyC4NqVHb/VwYfl/RZg7te7PoJUrtSgwl4Y4kigKDClmIRi
xpCc/3nCpP3ij09CS3NIlc4RCs5Biz35sLEDH4YIpOgfY6cvqcIQ8Gaa0OFv/VmHFx9fKhXco+Ce
Ob+YKBANcEUZwjP0xck4CSibPypN3cwIdR1wehFR3ilIJj49T+pd4vTSl8WhWasioWQ9hr/wnl75
qzur2EjMrYNDXIMi5LzFBIAsT7hloAIHPJ6l9fsk3zhUH12xgoelgawCkgN02j2PYX1KmAi1hA8g
VJ6rMOlwSPYc1KtnBUUnVmHBO7oUkvX08hXjmMWksPC4svjqU9Netn9iFLoDho6eIblIQf4fWNxK
8lJQVLzvwC7JrNE8gKQvx8PD2luimJTMktZ9K3bFCB8Pp4OQXQFVBSKhbzijymmMq84qJSdYQhXr
K+Bpq2fCAalfwo/B9w3HTs93TrEa3qoNzQI6X71kGA3Rf+qts42daOesVZF2hak10gLGNFRL6SI6
dJYylY4pb4dEAlbAjU2+0kBmFhfswIW1XceVlFuGt80UE2Yn01XDFAjaFw9LzLaK2IP8Cf5j/har
qQbz3Xu3dR6laARr/sPuTlqEbws6uqPw5nO2BhqcfrJPhQrmQUBXqnyqzgzqkF/4MvSCthPv5vrB
rLtmQjPq4oWQEyJSpRaBAqdX7ZbBx0uWm1x6I00slzK13DffgWzt/8fkonN1ydw+5CLffAIl0mnt
TSg0JLARB64sNXtXMbZzdkK6dRPZeT+9xOovdfsQixfr7XHygvCz1i0DCaYM3J3TAXfA0h4lyM3Z
n54sytM543nxdOyW0WBP/GVR0ku3u1hkjzmAJhzzml0yb8VRgPibe7OScG4aNeBxPJaJgqPTjwKd
hZakoV7jpRC9coMaRhUO768eqieAlJlT+tYIDd/2knG49tG7avAS9KD2wrQow4Z+yCsPx7dEAtU6
Dg1UP9sUTAtehXnNtuNVowVXLpnhtW7fUV6amxjf2h+Nlk2TfWGx4BP2oG2FNuNefBzfzs9bipQb
3gprpaSBoiP4f9VIV05EvLvzJc2KAL2auAwCdmd0LVKJJPyI4qP9pIXn9tdFN+a8hnT0Z3gsOaYE
K8hmYKZ5FYU/75bACwADLMo0+KOthayJ9R4H36RYSuauXF75ifRk/bcsrIErLSLvKZdnK3j2ck6t
aeb0QOjZQHMThXJLMA2rhXNJhrEs5yC4e695L3wfMdI19hh9IKgcdo2AJVGydrphTnT/UiKJyJoJ
VCr1A0WLabUMDgLJgj+Ip6W7YiL0Ds4+jbDRdd6rvvCAmc5j/2zJ0fyf17uzfQUR5ZcO2D1Nrdji
9MYay2rNmwZOCZwy6Zk6yQx5JgwA1iormScx1rNZ/pRncsVNhIwe1wTXUt5Q0dSrpvFqdDcnhNkz
wiUUcHJstfHoq/zTlSgGGE5uxbP2lyVMbBwsNc5d/luvNOBBGhAsOS7DUbd+OKJiYSNy42nLVvZ/
L7/EdcIRZi/RmL/r2aB/dHoH0nY0bhdwXLZZOE5YmRm4mLFSUs3HndXHaaAQWmHVDk4Z49Kwo+YL
26sCFY1dil4F3I11fTvmNvohpJTQWBFawV4ox1HPMG2j3dRIxPfc7g3VVtkOcwZC38uHYMUAQpKE
rOjZjn1pEWMNsMKIE3CAzpuDQbZ3P773F8KFPuv8jeTj28y8GjqFJ+90dds0Jh93o84thSjdOEAs
5lDHFYTQmZ9qVTHWuK8l2mAIHaCOQWbhY5HFUdXRvH4zNjBSyRhcTGgzQSVlNmLYHQ6Kdjg614F8
WTtlWXHKUDCqnLzbXU1MI/N41H4uaRiLW3g7eMxZJKV8TumHrbs5pbF8vn2OUUdbh3pku9iadx8r
uEljgBl2lCAu3nWdkwpapYUs3zkJ6LgrQmksiSE2nGvVz2DYdOee4qIXjsKHwKuLXRv2LbQMkEUn
wEpoZBAlyIrHJnLL1vNYqabfRwVHFfKJ0S/RdDwD8cIEppfG5UDj8e2sDAk91pmdbA/ATSdVV+xV
MLCACuW99c2nMARhz7PUnYx4Ml6KrXFKKpJ2ZAIwwQ9cK1qIdXcync1POJekitF6KSZX+ZmF5Z3B
rAbSnccnTrxnmFJs4rjL3hYdFVBRpPQUmAU17fvsEV0OYKMO0bOHcpoLQlnSmUJY6C19mit3I8Mv
q5XLj46iPp3PqD6v38w1+an3dIjprX2HRQlvmvfhPQW+L66VblHZL6yAZuXFAhRKYU9hWY0JAzXP
QQ0olIqhV3aiJi6MzAbpUIpGPdwYSMREROlM0kZAX9hUsVCILNMBhNZ09jCYBaoYgfrcPsdiGk8R
LjBvnU5QT2jD/U12b6KgT6fEICD6G+zND0JQX8/8PYUU4vlL4IYNcoiUx2E6aBhbewBMVXLops5y
gIdqxe3oqhDEmdTlkAFlBD2xK93ztbc6W10SHCJCjW4cZDk99EnKCobqZWowfW47qfrzH8VH75c7
8R9EIFLlBARqE7MSfQqlSoiE/Cy1KrErdEV5fvjPQMo921o0ufT8THuhDwRvd1zPGhh/lZiV7vX8
gK75xbXFItKAPTUToWBnsm4U3/+ujZmfY1+5ahmhfrV2qiuI8yUfh2r1PPTZb1SgFeLKh0H0oZVl
yaTAPx/IJ1lSnZXj9TyCW+YNgTvi80ti7ksfAPa5AOcz3NNbtFH1kjFe5Q3Cvmrg/dYh5R2VeDuI
IR3yoqhA97eR5VKdahROq08z97E7ujXZP/EZEaUoiJr03YmFW1EVt202y7TubmFSLsx5MFUA3ZRi
qOi7y7lC26MwP91U6Xc7GPAULdoHwe8YxjPeAoz5Y2o1lSnCDodDhNoDI6j6ARrdGF63MlAjs3Nd
y0qr7if1wq6wg7DBSUG3cqs//UdLo3JoiENS9f5gdPP52SdfWJZF2Q7U95Tz2SWJRHYgNPVNGp+E
6v5jJ+qwNaO8WEEY1+/MftsjFMZpCTFotR4nfCKPsCFUzOYaVY5Iu0OfP98z24SiLHGdy1U+/ywU
d8GaBd9wBogzqPu+ivu6QbHKLO/7s3948ikqxffqoeeBWqnQY818VNKnkYTIrhsYITsKdI79CNVa
TIiIqu9sS6Yg32pXYHQhGi+0ehOBAegzDjUEkQk3Ysu2aejpZAwaHIjz1h+4MGUKHFxCHbEeTBj7
JGniprRS1y0g0gWj+mwJC0wbjf+ppbYRgaWRpphZcI6vN11ml3tNCN0AV7VD042gn3K9epZ1FbFQ
z8mK1YdDhGqgvulrvJKTlQhx/S5orfXjWNHEyBc/g0qVghTge19MxrXCFJFBgm2yU6F/ke/VJt/u
w/eJmqQjZSSebXlv/L7KhXkxFIOe79wbFkPfRmyhPCeBgbyrSlLY0pUMnWavqS2TE6KsWxUONJlZ
SNUCyDY61+RQK1nKxfFwHOrXDukZ4WzWBAHVPXovaifMiJ/JSv9CMcI1goYqY2uMn/QNd0hz0s9C
PCxxcBS1MEkgpjpiFmBRhbEtY4E8vycac7MtZRXrAGpo5uBWhMZ7UhiUgLXrExunaSIus4qStPie
SVzLHZfP4uLZq1S9A6jNdZJSumYAENyORW+UClaIham0BokXWNHXga2S7Hhyhzon31ICeBIvOGBp
w0yOtG/PpZInPBkju6a57H4DFSnM4wmeIN20t7BWDCcg+V4NC//Kvw0r7kQrsYXvEaEky4roxzD0
6KHz33k++OpVdxBVazO4ipaqOYe4/nRp+1qTlEyzDOT32S1y+5sOUXWef3dodBRxenTqVhi4be1U
FmcXr0Q8zWBOZ4fOupNpOmbAncSlKVe+ObtPQHyzQwYGnHNsVNGCqdhx987D1hF/J5/3PUfLhgsW
wTeSZ3m9dZbeNO3j9wpYJO+Bs6rz76T0X82HF3XyBxvlkbnMZ851XlF3EoULpyeduJssTGLkgjj0
HOjA85upuUCdDZ3Rx6e8sdamjhelSYyPo5hPtCE/b7rGgi9gZQUzZyM4K2eqEFUwjybql1fK3Ycc
b6WmIoyie4O/Y4cnajEAAyUdE2dlsjPzFdSepuJQGwZjkoGz8QXlt+p9sJqIEVBpwO5hUJSmutI8
p/KCO7kd+nT7KNf0R2PO+ltW5SK3ADo/B29nZhhJTpe04sAtvBUAGCoK6ihyL8qd8vZVj4iXl+RO
WyUApJJtKml3C+iQWiyTakadkVqslllyo+kf6yINqY0ie6gvSo7bttEXbzmc0gKTMhmFuEB9hFHB
uf1gtLcrkaNo1ai7TFmKiefh0YpV619n/0LJ7y+uu7OwC0lwDi+1WwKjKvswlnLOvgknvhmUa4fd
oNCHdJdI6JpsWlo6SIPpcf0svzxRnJ6SHZhHYwS6xj1AZkr+Wqz8vzBkV3icOL0wQ1OHzWVbrBjR
9bkHILJ0dHgz1tb9rAgcYYvFJUJ8XXaOQQYXhn6mvL5L9Ys7WdszlNbiILfDh4ycXn59wqLyELwd
IymFH+Pa//cnmnRFBv+tUAsCsbrvjDlCQ6rqjmYn4QIYgnOf1gGHVUuhXCmyz5amie+/nXCF6oIT
/TJgoWHIGcGG9Kt7IESkGxnSaEq7lUKfmAFNgUHrj9KY6FhqaquEzsqIhmx3wbd2kBJmnSucaNfc
T16HqsBOP+ymx7jRarMSQRmu9OID0zbURlF8gWO4vKPIBp1z7ahC7etx0FSpqdTbLM56suxJyFwR
erFutXA99Z0m/3udXxoTSyVrl3wKsr2s2pVGLrS5ymxw1OxosOMVn4JWSJmsR62FqMgw/zNDsNp6
WYgWYYEKvom6Tbeth6UKhD4n1ola2HEgtbswLUbUpJ/Aii20PZAkdygHorZliKOroJqXBKGRkm8t
9846D1zX2B53qTffgxYkvCcR76uYXhnWmKHM81PJDLnrDwhr+iKp3LZacJOGndOK0m4SevE2THqo
Y4YtVjlOJ45GjV9q5HYpNDSWWmPJznODqb87sELjzmY//zhUvXeW1SsifH9l8Pd4TfKyURjSenQx
/tTZjvrSv1hG0llVdmopaiVVDFnUMa6Ghi4pGjPq4ymdZ7E+vP1aqn4jrTQ/PsrRKDCCforWoZar
O0Q4KmCJBoblkgiIQVlc2QDKqUWnZq7sdRY8uaBjqXvoLm22Az+sWYnxame9003xB0kOpRmMEvmI
qsPgvh/slTouCHOEdZpRnPJp3m/iSy4RDdNCKv8Xg/+TzgkVRD3z+p+9cpqdySfMr0Kp6kscApzx
xeqzMbe1h1C8Y+C8s3KioouXOdqZXzvAahiVlLtMg0T51TbDh1lXqnR0cX6YiUWua4fBI1Q57Lzn
E7wj72zMBU3GzoI5jVCxG/uMT1NnrWwAs7cSXUMPF8VFJdvTn3x76Y82B8ntw9Bd54YUnLAcU6Pg
stBkNseYEHM0xHRV6wuSBqlA9VZCTm5ZG8p7zFMEvIL4sDCt8HispI+4t1LTB8kPVMlNH7mojbAC
n4l+2I4TSGq3OsZBn0lqJZnuBeoqssmqn7ubDklCmcZiUCUUz7nrZ5hmaf72UBT2EI1yWBF+IGJ8
HsZuySqMkAc9OIajCZLQNX7AI1z73Zzpiazelz+fSzhFqz6RCF4sHFzwpOfUIWbhGiSPeCynIBjH
vohHgtDLKsj0yRzdGjRDKVqiUTnlBFwPTm+i7zi3Gmrm9AN819MJxqfp7BTIuywMj2LbhEHKDaMU
v9gW8lZSARVg7s8Lsl1Bak0hzrvZOAE7dtRYS+3CughFjb5W0nb+uA9/Wnihp7/eYHfsfxBGDpqY
8LxRZALs9GpaRYzTjU5HEG/iL6muNIhN7daZwxuZaRfOsM1vpJh9q6JyfF/inugxwHTccBIn1N+y
PKIBhsyugF3tDJ4k69Yq0leR3gPepZU//nF3GYhFBOAvInvFvEcSTphLWU90n56mUbG0yIk8XWz6
1oqAHDCFfg1kBLTLhiszOVz/4ZToX4OwCtyJ7fqhPNz397KcylHRGpMrXTJZbe6Yx9oYJw1DMb+P
hfomzmuM84GzUtjDg02X1/R/UhMKwt4T1/z1JsSwZzNAtyTgB9K9PPwOxoTeFE1S/WQT8lRL7CZe
0SHwrx6ovHyKRCejePHFsoS0UMDoGgA2FYZmra3pm0Zp2dJp8wWzauDz2nfR8gz685sJNj/0ZgiD
VQM1WV5LH6NcoQTQrPPyP/KoA0OjL8HntnjeyN0bI5XsbTeZE55byTftVojwmR/KVptxY4/BOXfj
5ZoWxsj05IqDh7RVmKa9lH0YCRXwZwxk62BBE7uIdWRjgP0QKscztJq41GLN1lkpFuN2tmV4CzJf
tk3zEYGugdCsf1oaZsGKmtAEzaJ93fuUfcv7vpXHPc2GIwnmNLO5P5+ft0xS0IRDQbm6Mr0q322a
yZBkifRWoIHsp8v2a7knVawNLHg/w2KZ/cFl9LtpHjw92hhKm2FZvsh4DMdu4/rcA3txfv+OjgA5
zXXx3dj2MPuWagOCNYuX372jv9/CXX7oZhHA/hZGseXfjf26WQC8Pkz99AMso91kwxU4bYfjnJUZ
DrEbmjOweQngm2QrO5axFYjpMSQ5oxuudRO+RMsQth4L2SoGi3aQSGXUBOp9g898wzAbHrecpW5F
J1yjzit/P9tDpZcgNdT9WL43Mw3bAYEvewXHphoiYWbLYlL5iM2zth+WKKDZUdRjxf0RYqL07/hN
LI21W/yplNyIz7fZNYJ8eGAHDYviNQgNRARXSpZEFkLr5d/3Tu4oL7VrzTJHtYNrDKkVcKQn6TuU
70ktvKbF3sS3yIcmhNQvgNfivKLq5flSKyVrIfEPl7uuuVEbWF/qXp+P/cnfIXCBO7nr/T7rw7sw
VgIJn05kAdV1exS9Sf4PTwSaTKdoLIH8g7uG/+bt+57EGFk6YtQi/d7WoU7+1r9bsMbp7t5aptgJ
1V94U5MuGGysF/BUTzBaMg2ukeZKHqz5TZkJkE2cDklX2/70GAOgJszwauNuUMj+nFQ8FJA6hY9S
t/y6JCp8xZosWwQ9zlsgI5ut61bnG3B497ecPsMuHmlDuV5fcuCA0SO7fjBkj+3zp7vRhu//b1E4
oExIg48QCTEbIeyYeU764Goh9TO9D9Wpkece+Q3l2Fn6atSZtlHzziWWt9eSj+FejDql8fyovA1L
v1fyPD7JAf/Tw0om1ba6Ec952lIilLSXJN7XyMWZSZivXQBIsl39Bn70VBlTuH3MCPfctSSlswjd
MHIRrz2XmW5s4cNWjgpujKegW0lytyab2yVhQBgVyuo8tPv+wZAaVEXmD49AMYU5EDb46cf6Ybo4
zyFEdGopeLC3dFmZuUwbGbZOW69zXog9HsmT5UBxGjYfwfaQUj0JYcv2xsj29eMMA/8dgArhiEtV
oCH1wDrpUWXs7NA3d0HjILMahhxXp3W6yYrThGEr9PAtGyyXFEsYeGLsk2vxDpaJUwHlU3WEfCGu
3w44W8X3eeycIn1SidZxV9OCwFS13JNSbINMokN+yjHbS1r6MiPfgf5GqE9OQ7IABlThLQSLsWH/
Nfd9qCK4cga4dOYH0NbVohf69TG5l3IDsOrty4pkXJ7maGn/qE2NOxhWeKivsvoIW5ByJeip2b+h
dMZ/6Q+xETkI2w0BpTdVTS4KuNj5imYO28HZE4NmUun3FEumWrMTnuu1T0tP+pn6q9figDyt90wa
Vp/0rq4CdaA2AnpL4IhduHZ5cp3BPDeLu3fWb4rSAJdWSO2I19LkxHdRgYf4Fe9fu/HzcWHlgmp9
a7xODaZCTiWmFoqbkiEYzWTbv2gLml9JwBYJXF4TkGIPCJBh9+YHLX4nMo3RQNgsTMI8mFqJ2Tem
G0bYZSdHMccR93ZmsOAW5AdigdVmfrxc2aqffMpszZMH2wT68QP6bx7zLbyt+Yr7S3enXMqRIWpK
8TpizUpdHaqsNQusP7cDoBM5Zx7R88EbEUHfB9JHxu1HHBGvjwpyNFX8FEl6VM1BUfrK0hxY0g+R
7gXsw4JrTcgEyU4m44xmt55+5Z/9DrdO1IAJ3fnK2HlfqaxcRqpqe/QT7lejJQ8rh6UZLfpKZC6Z
h8tN8QIYuR7oxizUmITvqR1LID56/yS5SzU33jEKePL4sghtIq9w14Tw2zM10uEttWQmrsbgwa+F
QaJs8cXRcW4gwNXqnZ/7oSkkyQfT2It9sZMibfRgumCRTQCVzmAknztpwXhsnd7M8eucSkNDkXKw
eutXqkjg9EL9rEI5/5Tzu5S7eD/gOKoA6plYUfGIbbOenCjlli48ItXnvLUPmk23h8DYzjco7NjS
lMz6HRARSxdLwWs/jRQhZNiFqcyTeCoP3poce6VwrGeKBu0w4uKQKP4tPHGsH8v6M526834fBnZ5
GvJvu5AzZXtxr5CTuqSxB+GPGXM6OG4yZyjNL4ENdb24GoM7I+FcEue6LX0/MQwkVgeWQgWQ0I+i
HUVNEW/8ODJNUjfpM4z1rldr3CuWz59NVms8K+DKmqbjGvGACuhukqFe3ZGrEue18raEdR6OnS1z
oJsijeKrkVc35Y/RUSJWfGX/168O1SUGdS0QCXP3ObOaM/+Vn2ztVTWZSU+7ATRW2SubC4hmOHCm
X+pgWxblcjfo4e2bKILwaXd5tpBF4/lsOSj9tcSpOzemmJ3pJWCAyB4LuNMHBiswHOW1gjtYFX0d
0Fo2FSPWDY3OLALX7vQAfzis7WtMSweV4k9tPKho5MNrVfEwiO+3D4Nc6dUkW+LHW5NKiwQG4fby
wJvYWxMU1V/nz9vTyG+G5gAhiAFuXnMtcyMVv8kprOWN1+Mq8XtV9DNW/PoNu836sTfA0tAIvl/h
MWYH9oNZqZJsSadFg/V+7dnZlflWUCFntCsaNmRfi7mLwWIp7U/FrOTW3jKgvP5S3lHviE5p7WAu
vtR8Mm9PP12DfV3yVL2XIYUw+FqNLcDnzLXC1UkUJv9GYEqSAShWvimWb+Z2AaRpS2HWqBrjXnie
YFkc8tADCee5upNAhFpy9pe+jDPdpHPAGvb6qw712xQwFt0Bb+ygxuYcmb3Si4yNlrtT1VnRNeVS
EDo/AoQKnaDG+Qq2ECTeggV9v+hUL5Ykj0xSn0bcDZK8y/vDJlEX9AqnodWI/60PSpSfcRwJSc3L
aO1w2+w25r7rz5NXBca/0tUcsqhsIbJyNM3T6eeU9tUS/YAbxGaaiULAjU0kGzBAVFQYDcI2VmlG
hXa14GEwzFFEQHaOMZYUZbaiz/CpEtPVooYSCxzUfqiPKbADTLz7QhMnQU/41fF4i8z2kjJ1HSFe
kaPLOHk3ZTvP8Kc7la6xNYmAXIMOSn9MPNYrVhpMaydG5B/fgVx75DCjgnzOdviMcIeFubKgNYHE
wQvC3a2BwzZKoHQMv13Z5xCTbK3rHJUNiL5VHRmIuOcZJ6huERLlAQNmtAcDLWr5MM5VzQk4lGft
7RTeR8D6GxCRH4/gYbYohOhh/OYgiV2ivXeuQunclkBGKuvhTp1oScpb4jcZHjATyJErlGpGAMbu
XXk7sxUmLZNwaC8fdimU8y5MdJwtzucEeptzq/qIvup1Re7/2L6XmolPz6G1CN+lFBH3if8K4CAp
OtEwpPufcoM2CQNmVJ9IVelav09AeMuEpRtmriVJ6vg4QjVljHp5Gz+3DiBYpYnkQ2Jkxr1vCVIU
nexgWVtvCTNYg8tGcRhnlNLjWyBofeqooKEzdmLyGHsCZlTodURpmjp42rMb2V+k42gVoCtpVz1S
x4KPUxKYDwiGGvqAFw+q1u0gfTXrOE5zyfk6Ve3AKJqeGut4q4ShlOq2F2Uh6rsH4no0JeN/AEnN
ahzzXhsGy2QPbQj2vvrP+d9Jx9tSLQF7fVw4+vXRdarzv3zkZFKv6LNpTEs3fl2Mrxg4aV5JcuqY
OzpwAJ41iT92VjQV3d5ISIiio6VG+3tpQAvPIVb6q6rpR/7fmYqakgl8+x4tNH832q3HPegYvogR
xRxOJEbkG4vj9MTKFLXPPXvpqFuyq0ShGWDopZhRjN5NfnyXoBpVAHLubHb9u+a+hRexX6YtmwaQ
WdLazyYk0VR19ndjbrUN5X+wzGxOzuYfHtw16kUKP4uuwV4rqj7fxwmV6YIL+GDbKhpTU3H6fEwU
jnpshXeRIGA4Wc+jUx/XZ89jvGwv53TqciidINHdUzMp6msF7Fge5rdUyhu5dDToI7WjsDkdy/b6
wzeSIYW/c+iQ0QTh2SQXzCD4AuVGFjqznTv/H5oy3xAo3R70M9xCjmUQdyWHjOJbAlvVUzj4jlhV
wv+VvEbi88EQOISP2lyoYUeOMsL7fHoKjUS8rMhtst1R3vb9vnisu+EqzUZ39WtQpynBYONpfMwO
BQDdPciKJ//mYKFHJQ8KOmFN6JnNrQFZUM0JciG1ApIMrOD7mI1BDuWhjoc7hCQNOeB0VdpOQr13
QWok9nBcE7EWqzDYxnzOZT75+NFB4Cuz+UQQolPOEuK1Yni82PL80NB86CFJjZuSlZlZusYMH18h
SG4qteE77CY1Hv34USykkZBweDOms7DHx6bALJIjI+zpUPrSYT669eu6jKCoCUF9pp9qL2XHABCZ
WjAF6UudYZ/gp1BvgVjBj9X5/875oI3YwR3m1gnfHsFhpi+1Z1qUacdQTS6YmI01yvMa/hve+CqC
wCHfr7tFp5bRL0sZAIvEfiKU+fTE47yEdEnelbueXjzebpelndWKSGVWQNl+O5Y0/u/8fFABjIsb
TRmu+8WUhSJiiEdrEme5HspHL/hr2jaVrORNeK6TKi3rD0gls0kmLxwcjahYPmD96WIM0Ucg+6vi
nfIA6yrtGAw4Y8uWdHoFNNWd9Ehgkcny67KdbEYiqJaJiwvRLmUwShp4qFslrZukcxmMWw7iypIF
jYwWwGKUQlfPMhAgH7QeuWOP+2sqyGaFn0WuY0bdEnCWnllVcQkjN+UVUZ73HdYgS+dwwM48u4Aq
/5ZEt9fAH1F0CPrCtGFnw+E/o2E+H2mB+zg3oLzNs3ktgII8z1RjmsSTZrOCTK2bBqVDR2IN8OeL
Idn6+EslCPxHPiyefej8Tbpe3lQri+3pUDozOSsJI/NmO+KwnvfXydlzy+MMU1K0PJksOFtA1Phu
r+qIRxtnMXB+t3VRFxY0VAq+fNTvbRl+QuQoU/EUKSlEDaapnt+pcC0jGjPee882H+eHkg6PEznb
M9VEGLdzHn4FAgGLJkWLYEO/tLJ/W0aFcTjoBagHUe1KP/O9l0ftyxSiUqvJrRHIBs9mJk25bqzO
9sCJL0dgOMTid37XaIaA39i1Q30HcWRyqeETMJ1Rcxwb3c8Z5IyCat8ti3v7hvwXUrp5YiC/epHJ
y1/UeTYDkER03N/TwAxx+gv1mdz3/TTX15fDAwW8yaAGXR1M/llipaJvc6W31jH7TZSM6MfF9E+K
RZNwyDKMUBwvyUr277Yopc31jatoAQU/DB8++QlUA4VvOUsQhY8dHC5K59deZ+aaOCCVd/R5HF4X
oVOCWS1wU8RiL970bZUNtaIqcNQtOnvIT/8sJ8Cy/JNQ4Imrmg1TQXjnqXmMcL6glRjLve+p9XAm
dc4i5y5T2I+5msyk2N37pVJltCaaLJV496ZkhQ47wlFxx7NOrfZyREDc4YlXxrMW2kvASdCQSrh/
1hKX7MP1ZEHstO2DIw8xW3OAvbE2ALbj4a8LFtPAep5bcOYS9Xzs2SdbJY0MetEL43pE2prhdtJD
cdyWEED2MfSel7pFOpUR26iKwlENIRUiwD5quZ44PMTRcohndH9eA0nsHchN+VRigbMEsBqrgWhG
LBBtzR9Ge9x8ljIOZ0hhegCWiL2aSUS8uJSJMk8AROX6+bwDERJS2WrCxK5i2nK6TX8Q9NqiJpUY
hTAfQ2B14veZqLq0wnWQM9Mg+bjSVsgxSSOLKj1y4GBH6GzldJceaET0q4bGWT4Q3cLrdf+bljxZ
aN0c8gaCUqTxRcRVN5b2TVIn6E9rbAbDkzyNfOU93ogXvwo5tHBJKgR8RxmnZyzJ6hdFFBLdh1w6
xnveEmU5sDqzPvmZFcmptw5quyrC6fRqPwVrNruvuGkCMM7D/ufDBaVkYXK6qqIcjm42pRXFPs+m
78qswN60nLWNkxVMo2/KkPT3NJ3HSJRrSUarM63r5zkOX9Hp8Xs6N9cjmaWs0uE+6ZRLOdHWp5Z7
XahPqjV4BU6NZafOdsulW1U2+lgSpB190Oh1JxIA4/k/yMdCoTMkz9O82oopRQ1KG+dnygcxjEG4
8zTz1kBN5qO2NquHWpNwkZVxsdDPnpdKprt7EfQa+tqaX9b94f8zS4PsUhVIcbXr0956r+Iwbv3k
wQTNf+ExplO4BrKPnmy5I2+uTkbNk0/pmOTUiVPRHs0zn21OpYplHGPdTNOSSf7xGa5tlTYUw8a5
+ehLekEvGwdjARFN3JCuF5D0R8Ypwl/f6nCokr3o4rt2a7rsIqVsDDm4wxKX2HJBAiwFASXXj/+0
4yf1oOL0/xnh9AdyGZQ9CE27i9VUMXoFeQZAOsNS1KuUKA3HGAL42yeo5wFo3G9lfk/WDrgO4GyK
stZGYcJS108fWDjmMYC3TjsfepK5VjsWxo1tSAbv+O0IHY7MCFFShTecV2p2gh/eWP+0zbBBjVRM
apBupkKAA+BOEVklsijTtm2bhxU90ALxkHbltFucNfYc6WLwNRwkoKZsFBWnFeMhXMS2WZtx53xc
xXy7fBSpPdl99jYq6cEjrRrHnpMlSsNI5/qjWacKSLBjrtpz8rdAUSmAEF55EgBfXJGOq+Nj0qh+
3CV8nlM68t0fPqA509G95VWmMYaDFb4e4JKprAeHu14LZ51iVGbVjkG2zDcm18uxlCcT1R1qRgVR
BqNUmqiTAAlLWl7liJEeIsMAr3HYjxrqdlLGhgqUqpINtokZ5rKl+n2b9XKS5ZMlHM1+kcQE95lY
cxVKMaDhks7z7BsD//lLjlWAnn2fdeFklYFGXKTdeKuNuglq/9Qyy2bbm+DBxXwEU8nJnH2iTEgx
LT5np2YOEkegmKr49YKQzdbGm4YnfkcbC4A4MUGi8CfOOfjv+9rcCLpNgFgoks71eO2OTtsmbf04
k4X2zf8TSfteuZSNuJckxl9sVKaFRx+Ns/biSoiBhGhWkf0dGArS5S0PWbzChAw749vfqVkqmx3J
3Xq/VcMw5Xa64tHABASHNkuHpDM9otKVXiTF+6z3kxCtQHr2/BvHp/miNDwg015codL8TDbz7IaB
njBsgQdwou1/gBCXIJbxzah7Nz65hiPjaRdLrjDqKOFQE1ebu9ceH3qBffQ/q+/6dTY7OgLMCEFW
rI+CgG7500kbFObwmFGpL78TNMHfLyk5mjK105Tn06ktPZTZMTO0WR/Z/f9vK/koxUoxKNgo+5Nr
IGneB9mVSLMjFXQNqierqBdVnyfPzkpkHoqKzQV8jTH0p5kyzvwLNffP6bFxgFozcBI0Hbc4yBf2
/3LQtuli2g0UeeEcgE6u1xsuHm3dMfyqtNKqACPfu3tnkyZpgqhuIRDDEwaaGBYoGW/epDkQs69H
yWPxVbkpW4M6xAv4KLn8qE5fq4oXg87SJl+atfGNbqObpwp6/NjQlDrUdZf0dl4e55MQNNu5mWKC
CT4AXlFdJIiOJIRCJp7d2THgXP4WID/QNcZli7MWjI9sw+PazPZYqdbknzggZ9NgZxc/hc5XR1P2
9qRF1mgNh+oYyoYZyHigMTHLERPKUMtFMu4ufemDlisOJ9tQoqT/QKA/RDfV2eBxDnnZKsRJcFt3
VAi7O36d/DxLW/JzvRB3k64ucu++6RRn/pCAqmpxuLeE6FRtkECOFsIFQvn6pvOBB7qvJDZ3LIgJ
exWsh4cLdU0I8z+pl6oJk+J0hLqU9l6TGiOb3wQ1w45D9bPSlbjjUS+eVI2qwl11hNTgXedIWkj1
k56hQf7Z8h4c/VxQ+B8O364wZX5O64AqiBSm2tvxtK1LTPQDk5wSSvgClIvu1I6VEyc5n7sefDuz
hQObSLoLr6vgMS3OAueQMbGj9yefV38Fu7sRDdZWZjGWYN/P1sotUD2+tLHjCxrHCg7Rawq6aKR5
B2Dju8WAe/ZedphIG8e+e0sFWqftdnzhqjudZwb8gVKyeci3sr+A1q2wPidAeEtBfVBnuql3oFfs
hiIH2sLdktPp/wmjwnfTmfbqxlc+DrJnWM9bldcfvxYidArYU2XSPPt8SakICeUobZm1DvzQnN52
Zw3LXLfDy8Mb1O0OqyTyxUZPyvnNz1+yfRnV2Wjp4dlJGfZCI8FZoTZE5lHAsfXmN0E1dp6zUmn/
saXNgBRnmBYLAjZfXNp0+95zBawEuXGG4G1dlomcjr/A21SHUk++mGEopZ6QGsBaf/h8wSPuWhqb
FabnkjBid3byJJxVW1IIUlmitXWfmAmv1loS76dlIDbZRTatYH+KpbYJX1O5f+Evabqrz8CfO4SZ
O+jfSIQhBBeNXTlmRHFBANm9rThBnS4XiJlZiEM61kTZGvtEpx3/mcvzT/yClpI3VKntNgU8YpEA
P8Uc2Rnrp3js6tIT0dgmSdtDJx0ZlDIRaI4NcyZT/GkEQfiIAMjbR0banFx/3w5IjNj3mYme2tVt
N//qxRePvrEVM/xeyhe+BKGkPv/44twJYQxaxzD/6O4oiqJ39whUAdsK9i+kH79qT7qUQ5MX7g6I
tmH0B1Z8mnpxB0PsD6zlKVB85hOpHLz0jWaxBUBQqFG15te1OE3qYeeSCltVTRllxActo6avm6g7
3NzvqpJSBFTY8QzG0oWhudtXcwFPCW5S0hVFMIcD2BxzhJqnCsd7SkVP5Ik7/BqTkauQLPibZyhx
+xhvFvOs/smjL3Hefbk9WODRlbjByc7PunG3s5aiQmhB9Q3SjZDyIWFLoAhfulleth/FNffyeM0e
dwP0myIC4Et/9+oNMocYDwmRzp5lXe2am4u1eGEgpP1z596YSeyRsTKjBg8VYv+fUBpHf5fjYDd8
tbfKqEvsuQVAWErJChIoI4eATb2R8ThRW9WR9vbLwsV4h7onvxsko8LFu+RRqFW+XFUBfVnARg9o
ev0hs7BoPweqI6mk5yOuKw/1IUJapt366tu/8tlr61HLZLsCW4yiHd1uufQ3sPADuD2UzYvdGNrk
lYeS8s05ETh/Rk2yq+JCIL7vh+xTVtInh/xZNLYscPhDAur95xNNAZehtZciM5nyGIdwOjrOkyuy
d3F9sRgv3i8T71l9d+ytoJnWMjFWmBcxCkVjiB9nYkY40+GHeoTnQAre9OuDPsR1w95UE7GVhKaa
XhOe2WhhFORGTVBhv5x5axcr5rkMcCcHAtWGvmGg35qbi6Afh2cxWnqqUbGp53VfIHMSlUxlGod4
g9dlProikCHTZvwlEKLgu2mpYBMkQLFtcrNVTPt5PwFpwqSHkPZoYRVWuqzPlCzCWoYS7h540QX3
ne17Oue1mrdKyKLa1hdXCPbO5vuep9ifudiGTHL3Q1EDRJ4QxoKah+nMUDaCi4GqlFnpoRapIxRm
/NLZTKgIR1ZFPEx9tn/SYxLU0iwRCF9bfhrjKdzdSCPpjIwflg8F1CCtwPNqy7bcugOArddcJF3g
EQZmlicLJe2VC9f+q8MtDVmcDTcM7yNO1z3xrXMsEqCVlQAXbfoU/vK7B5c5XCPffY5/8Do2Qdad
z68SyF5XOb8Ez7gQL3YfDjlBcElSuV5QdqFpFxB38KLUtrtXj39PX7J1OXyHdgLVKMLOPG0fvvVD
DhQe7lN12hINCoUBUZnlh8MY5UxA3HIivyZLZAxkfqLC9HAKJlmzDQLfa8nAXoyteUR8o/oSxOhV
cLqcWnMW3fKC5LFi28a3ofWzEXOIqnQa6ByOqsHR6ptSYITDaotVfDta3EJQ/LOgTfnT5ra28jhC
KdRuC3smz7XKQKS4yEY84nxAdzIEZ9nQjhzKmRx16C70ZjKfWaeMvp9JLfIoPxmT3ZkPAnK1iveD
dpyw9NTnhlmuGULYls2Pj/j7DT6z0y2/1+Ej7tSMn2x/3Nc4DfdN2hyJTSYr1cwcT3z4jRt4Hn+Y
8vUps2VKKZRsjh2FBPX1pMkzq60Y7NxeYC8mnAOizCy2g+/4iUF2ck+yPWBal21nMt9gy9pc4Ug4
I7e9FIiFo6rm4Dz6gn5KHIdusAr0tzqSRKzf5YmYn96mqM2gm7GX3BRB9j+Jz3HFi+a3/jb6hUTy
0bSZbTH+b2hbx4jD9NEN+Jzk9BFlET0WK5OK6uXHQIJJsfnqr/zjl1sxQg36MNv/AW4l6ZAMFRJi
42IQKEgCX5P0ClNMTsUo72Gjpkp5V6V9M05ptBe+THbrOabGIkhpbincAuoGU3BkvdotDIMZ5924
C3+35L9K7cUv35tFvBmIYTTVyXiteKNBa+IjOJQ1MpVc528uHRxyazK1ZZUYXLntcK119CE8Ad7/
QhdF8OzY3zGLtZ3DWTfx8Hg9sKC66ZEDm60OPDFgvG1cPQvTMGwCNxeNsV8fSK3fIfeobBXshxCI
CyvyW3x2QnN6HlJaVtPHLXo3DnNfwEu0RsaeK6k561OB5OEa5zkDd4kbmm3ZWbMBCdwwuD608ixq
DSRMlbtSkhQAWBPl63lBlIJGI8Kf4bay1jpMxgO8QX4xja4cM7IVOrh+5pIFWEBplNvwa5nU6adQ
MPcne1q7i/9SJswjMwZAUYyk38X5tfEVVwwgNxYKjE4jYfB0soZmJKV5b5AAyTr769E+0MTfmlPz
fyUAbM/iiItQwHvn21yI88TcN582NfXMgdB9Zru0zG3/5VMTdDPA3s7L0Y0h6/SGaUQGSrSelvzg
4MqYZsZmCOtlgsBrW+3mp+215FXJgMeut0xbwD9MifUj26wXsNdNg9Ur4kTuTuBh7CkVJ8KTwb1r
MYdQp+1OppRKbRE1bl557jeTrPyvZwoOgsql2G8T2ZUwb8ifk5ieRxon+vANZJLS14O6XbZE1uSV
9AvGMW2wtVdNNAde42oDgd36SlBHMqysxud52qSyjUgHay9j/kLgZy8j2JE4s5WAwQk8yVIza8GW
YVyBCS2QL87fV7So9L9aMvZz38V8ytDfJMrWFgzUnM+niMu3WDZy2ubXuRaQh62IzgPIltFOCuoi
SkaPtWkL9YKefYrlKNH0PdIgRqcV4oRie9A298n2elLeRjoqx2bU9cNEMPE6/X4CMMHHebgpPMNP
5o6ENLSOBpSS6msWolw6+LwyQ9V3NLpqmvhxO5ZOktgxmhRLoLXHWuMusKsZ3EjgYaWF0r/XtQ07
OcMBHzlHrqa97Vzt8WcmuNu/GHykg5UfRRX1ylZ/DLiDC5x66ckja27sGvJN/gkzXzMM81AL3Y5F
4jtqLj0ZklAdhgTH4ZFs6riSYLqH1deLNH166O/erKMMdX+mYNDC1NU1d8w7qVkDmPByEl5ADFeb
hZgXgVTsJG5sLdLgsg4UNK+LMqUIEI3Iw9++9ktxZHejLwwn2t0FNNbGbrQZxF7mNN3P2k++coz+
DCZtDWV6y4GkMUMrXHL9EiiymDvTIVhiNXw6/OGT7jsMMtIyIQuILKt9EXzTMGSKpWxFeKRyxBvf
tYrVcD7kxy8yULyTx7PHurWp87bNIy1y0KCdoeDGi166mUlgoTpTnyIziPdfMujtZzHWLcva06CE
ZrInJrWG5Ir2nQ9koflhmQg4il99MRoDOv0+w/1V9+twEb3wxtkupNEmw+FrqWeCoUFI4Zrdl1s2
hf8YaRzmf48v4aGZwiUWsLJO3fSmy1LiglWQoWgA1lkdUSBrCk4yC0EvWfR4JPLlod8EuKsduJ9E
k4LHD0SkdBVtaLOs4XSC9vp9BAWMw8vG1yNHv2oSZvfsxR4O3cPpKToazQod1/i0EsLeCvkOMOl8
uS5WwfMP+AdNyS46c7yW3a9HESXwC/RGd4PuEo85orrBtK9jTgV4qglcCk3kgkCzGfl2Hqmpj/aH
riTCJxU/mndgTgbn/r7r0W7Dl+Jlu/F9oPymGLi9pmlFNZMAk79Je1730eruM7QFnWT9+zLWh4J/
Mth7km3Dqpv7g6dDrb8Swu6VA/2u3IZSJND+vbexA9EGQ7D4O94S42JbkeQCjJ1jmfD0kR7cGHBC
QMwBjmGZG6aHFzYgsRuBnjrMozFSymkxxgaGplgUxBpki85+QOiLyy7TZAVv4Oc+QXqlhfG6IkNm
UgoWEKw3FeDvETdtzHWVsHfurdfcVPB4/MCzQuDU+3jM+GGtfObuMkNqXUyhzohGDJKCi9DUhIv0
2lKjVUgDhtBLhH4HKspOq5D0Q9t0ssrhfru1YqJxvDUlgaBW1MWzHtTqCo6S5oaF7dRWRY/INaz+
vpk5tlBZawoMDIgpCFeGBuctE6SpMj0lOS5nBU3LiTrUpBNz36gNCsp6QibuksBaa4Fkl2dsBqyv
ML8nb/kUqjJvCl8JPluDIcEAm70bQOL6Kw8HF4okV6uCAXeRiFpovEPEOjydW7N4YFfrYPgEoVjS
tssIZzD8uyeHArBrjyoYq2gMXY9Pk+XPvyR0pz8uk2L/EKrBJteMaxUK/mlXix5UDb3qr3jSergi
DbQVdfPFSrY0cdcfbimDeZYHtrJOSnRzekv5PfwJ43bRt0xmgDtL5JUPmsGdlR4WmuTWWaxBFOXl
OltUGvjpWQcilURSrApqC9nQmSa6uCL/0f38W8wYE1HxISqRzosfTJDi4YLlOHLrOWmVgEpt57lh
l41SbY8r44V/ZaCJ2amVICOXIiMtWhgqZay/yufqc9uciLyrqjcmwrizipcKRkTrBrYjXIu070UO
r8OQjpXHjJrxwvfR4K6dUxzbw3Lv0NMnydgCeTtHIJ3wiN8xC2iR4U8Gb85lUX1j7X+jxQnvP/0t
QZp6RW7Y4CLXzBJWR05jX6hN8k/AQTglL7lEuPT3gFAhbgkfi7Ly6EFSg2yTGaIv/xmFpYd3ughc
i8uZbMiAHE6WTGy2qZoy9vVMLHXCgUaJgGGc6XwdF+aEAp0UE4Xif+2tQsI/W9eGZNUSwkisq0/I
sVxOE2VoI/s01ab4Vn3X+WJuYBV+W7BA009MirVBnOURxgN9wCatO+uWCidgbS/uba7ji/nn9C+D
FmuzyxdPMxJQzcbHdScZpRfzJ4yQOx4AAytkF8foeWN/imype1oA46NUXHLm00nf5cjUnZbq4f6r
udumbZ1s0F9hzy9L3JBfDv7k3bNEmfii15VKhhXRsOP8kHgmdCiPDu24XGJTw8HmSpbZdqLAqRfI
ektsd31IlHds41+Km9k0qSDwUCQhR01YtyR4m5EmtHKKyQF/ESp5jGNwSf/XtcqZZMuFsr3/7bph
l+eNBSO2SU4e3Yg2TJvXVqO897HG+owpPMps575tdnCCVBHB0GXtl0GYbEcXtounHHxd+jecKCiP
dlcAWUS4Un4ZEfkcsG8rL7yLVTufyqTLj9tW7yyUxc2j1NEQfK4vZDex6ynzEgLWjepoxrODwDXI
c5BzPSaMox2o3j4UNOBz6Fljv+n29q2hqJhHsaf4MO65jYgU1R1sDvOWzI9gHrMUe/TLGknA1yC3
lldqKzdRLRz5EHaOO97Vg5NHugB8Ov78FmfjG7nVaB2TLmSEOOm8wWzvv514f92unpf8ysCK/7hp
AJso4HOPAp6UbhpywWJnhAS5VZe9GyKeYcWDwpsSqjjPYVF6Z9ta7Qy0Yw2IOffvmPZAD90mQwQo
DF/ATKEE+twNsULEwU0YJ4dfRWx2z6di4uQXuzLr06N2FaVNhSd9/r7SOry2AFTZIROxl6m7TZvY
HiDSR9mpi9P16tVkfCzHvQDt7CT6W1UsSUzJZxDCyhcl7w3AVR1dKiBDuxU5zIdFL9UPURm1QjAx
Mm7EZVxVoDnmh4tPS7EaWfqbu8ocQe01Dr1X/y/r6hVH/6q/ShzMqvTBl+P0f+kXYaVoPPCH6Nzw
BrkKoops7UOJ5rtBrMidojXO922LEHcFkZgGAYoHoh4GxPMwZJD8FoMBIZS1+tPosJit4wjFMG8Y
7+PC8TMBaQMogOyFAmIfxHOFkWdOCJd5AqQ7Bi1DCutjdvMRq0MPRj1DaYCIR+v+T1JR21V7X2v2
WwWKELYNcGveYh++3pyy2xSdPRN+j0mqkz+hq9jsv+ZumFR7nvFSV7Wy9CDcJ5CB7cQ8VLbMuk/C
BPA0qbPD3rj6f55I/IXpnAzsYngqgSUoKBIqeeDbVIKfKZlNGcV/ZK2DkacNW4A3j6P+wPHbQCE3
PF/AfFCkuv3aebRWywzQjHiaU0/jwubBhqxrbPh1S/0a25viOLqlGRWSVSNVEPzITyehnOub0zAp
cRRbvBGhg5AoZc/s7IRqMzlgXGcLkdWvC1F3Jsx77kqXbdfu/n8FRMf1IFmGYhYx7WR6kedcbtPq
X5q/AXQmOt5rT8da0k2a9WGbl35GW5LerzchOmJFKaBpnobh2TdFcSqb3rUuGuLEMKUA0ueHlMrs
EGpuYoyjry5amSI3rTUD88mASs202w7afxvrqOGYZVw471T6MmxKVhZYPhyotzW74BDtbwFxop+8
7dHyA3JVkhea5zCtM8ytcwY5iYTrURDVW1rH6tmKr+4nWfCl6AYjuxDj+exR9v2lvQt349efUxYJ
Yk8/QWhmhkasj0xwp0k10puQ+1r2ZjYcjFoxdmuDFz/rXl5HTvh05BzL2s4PxK45VAPqTmZvaQ59
qEOmk1bVIpm3cYyVvJdbvN11Y5KYI5dwx4TcOy04m+qzOIed0wGti7Du7+4oSfARhA18WSQKMKr0
duFpb33negn0+Cnn4uzQA2ihqjE2gZXk1fiZLawhgKOR+28Cftj5VakwKi0hBbyNq4NXkojvf/4Y
6704ADdqu5sMcWZbboZCAVJXGRg52JAGQthbGAwelvzh2AEdN6nsNj+fS3cCLIzlwrLY5gTmnfIG
x06EG0cvbFALKAgEyFaOlPT69yOYfnPF7oNU2pVv9iKbYsRBBrtBG0SHlaqg4OAKQucWpSAYWnd2
3VhTxuCfPaTOGIKGILLM+MGVuXSFoBxMpt9ZCRamh3KWJDK+qWr8hMwgNd3+FR7cnygYF542w59y
LWLUxU/NyhSnDMYAJ02XzKFOPUvkCHJoFixjbF68yVD+3xdg2SM2STm5uux8S/NZw9+ELsBT8jnz
vo3dBVIggz8oNnz94EgF+EF97T9c1AtJO9JNS1Gb4/boZ92KEvLDWMAcz40pNJ8H2YZPV3IXhgwP
hbgHUsJz7SSPUo0kNcm/R4jNdUpViwkHAc/sZwhCnNudj6O6CGq/n9t7wDskW8jB9ZuD77gcglB/
dsxMM+dP+0keHakFyOeZPM458ncdGYodJ5vnEBGxY/H5b4XfMIvdfp9x4cUSnB3fcA3KPRdq5+dL
NBIAZj68EmP0R1fgXNGztw+7Uygr1CtSO+nDxQGrXfvDRHsMTv+sRJs5MHQvGaoPO1OtlQeLeftf
mboODDp/i9U18Dnvrq9N8hz5FUFd/MEff+DnPJj/dcwYWsltD0qCwSYfTDifsZ+XrUbs99fJO6rw
2Ke7qql8s8We7RDZ7L08sVLJGgkuERMsrMU6S//Irr/48jn+N4xLfF2YFizxdqLodjzAJer+AYWo
o0SInJdpEPRdcUYSHvaoD7rccEK5MeEk2PXj898U6TLd7eibO5aAhbYIAlNkP0C8s+FI5EVr8Rod
PXZRWrXozq1O/B5BfVOGrV8jkgcRa6kH3VwDLemTLQgXaJTddS/1bJeQ5KLSN5FQBkxUBo7L0mwK
NOd1thxeOUXCRjBtrMa1HCa8Ca5nxk78NwtDg+TOC7v9heWrIRDnIrUV6SXlYAmPCgRA/c9rNVfs
lG96I+YFrkhd1urthDlDgtd3xujxJALPVR0KOtRbRAKDUYHz0joZ6q1w7Lqe3Y8LOsTtxoglkN3G
ESHmCOeIG9jk5cTXSLTWZEH32sz9XBK1dhs+lbDeby2bS9PZ/fno5r4PI28pwmNYw3zuK3ZfdCbj
dXtqHnxf4cBoe1VGBa3lmiFZvRb+r0voTYVkHsfUnkteQG5Q0EINx+Oe5ZpEH2Lvif80FKyOmrHB
tcrByIznJchWlyZU/P7ubF9Nu/ggM8BT1dHSOLVNgqXU+ZutDDyGZONMMOfIrXQRoS/AVersx4z0
nSVdXe1oN3KeJmDXaw5hZrwjBxETayhmuc2lENA/8jjmTx2Yz1YK8j0k7C8fe6himYHHenAqnuqc
EeTbgU5ddq0ZTRNrGl/IHJfb4zhOyN+fHCyuKSVMji44DXVulEDzSjehX/3MBTzuAD+pxdIJdvXH
q0ZotDAJddSHpzhr69Ph+u4CPAroPnPr51dC0VdoZ/TdNg3r/EwYDuBMBeTBzyFenNLj9woZ+lSd
+FLA32EKqKxXvnnK7v+C283dIebJXZ+ibDr/Ur0dlvS8C/91rMsKgJUYC0waHbeDln8VshXsyDIs
V0EBQQ+JzgjPrPqlKIcRPxXtRAtpl2GaGYSdnTK+5XvRUtPoe9CQ8Kp0kCp5oXDkbGfiw3EzCEXg
/ePfDPt7cVNi0lH3xNRLcSTWSeXIrrm9YsTtajCoyeYAytSGrI5v5zw0T0JJOVovGHaLXLsxPdHH
AE27BE/yK3qJNeFQSWj2Y2PuvaV838BeAVRlqrtgM4q2v0OJ8XAZ6FILKURUAxGzUPK4WI6NZ31N
BD+m0iTY4bUvLTz8HGGuyIlI84q1UkFA7f/s7E1F0AsH2ro2BIKxwl7dZD8ZiJGsiDUAuLEDplsx
ug2S34ub0v7cxPdypNnqZhd9vvjBgoxVczANfm6gLUaPmrs4pGbz3ZWpsTwx5pH69F1Unb3HgFqy
aDJ2wNOqU9fwa1OfrKtUKyjwzI3hBAKTIHFrJ8xTaLB7lKEGZADI28QZTpJ1HkklHuTZa5YzTCnQ
YH7Wx7JGcmPM3WJ+T2XtZo0mp0m/0HjNmw2FQKjgsiqfno5Me84TX1GRmc/8VIYujXWnDd3jOiSd
cIvv3USQymramjR+WxddWTy4Q3HczKthnWyKRoUdHzDQJfFAtkYCmKG8O5pPUKOEcNcf08EWhMhx
BbWIupm/b62CKMqXuu88bFSiiEw01lagByJvg23rJV6vYcmDZ0dWq/MjNJHKyT4N93LMcQk22MyX
BLF8mzh2BKmfSh6zQwUcXdeAk0JE/N7sgxBqF6YfTBxaUvO9pNzdlh9q3qXA5jRaoHFN2l1Fneyk
QJWtmjEp22bxgFKKPON427Gj1QwlrVTAXy8Bacgk68HVR56hI0sO2Hgjmcoza02sHHB+2NoMFeue
a+H395pAbexumhH+cfRL2WI4OPJ9JFGqSdTtkxOpQlKeiey2ikNYnq+sdatdiExZwSjZ+sCZSg33
x782/nL8mGDfe4zN92dr178nKEAx3rfaVBOryUOOdYN6GGsvernpF3KZXO0MXgQOl77tmSXnLso4
EoIOwdEWngDvOzWBbuSLn5LYeALuFb3U1jCUuBekesYXM8zOFL/ynkUOl5BWQ7RoLD1NarXQ7hLU
ncQHarKI1Mrz/3VErS2Gj0OTHGQlLsNzCmWDT9ue8Q5cXcl0KUdKLVzU78z5FQcTNHdeOXXwAxis
XTPToy+y9EFgixrA8LOZdqhV/YY1amQFaBqJEaBTdzxkSBNBCQ+PQAb0MRtuJstGU9RVRBKPh6s3
KN6fohpDKm6lOK1Ohfrteh5t/pwh2IxDtZEVotIuaydTkdT0G5mu0vu72jvw82GShYT4NnmlqREM
B4OM9EKD7TcoH0b10f4PTs6tpKH9n6eQRUOWnC1Rkq1vOORcDanNFYV/qQxSJluiu/HzJ8aqSKpY
HXPoChtAYDVM9ctWQScWsDb1qS5xr6TYO6THSNlk7ouZWRABpRACydbYj4J3Czqk2BgRsIjPdeLc
gXIWVgox0UICQtz37ZWKVn3KrwTH2ZIQhHo22+RfntxeuG+tUAjkdv32Kh0bFw7/m86iJ5ArZZYB
p2BQeCsZKJuaXYcyEHflwKkqExu3da1amF8vKOngIEYf8gSxeLprZIO2i0oN/r7BabfYC0ZUg/ul
lQULjoon0/TwBd6aloyA5EJMP0xaemRkWlPxHh07N35xxpWySQRwVJOQf9Zbf4H1tNbO2VUe5j3s
Tj2Yi0J3PHbn9lDBSqhID3RYonASNbSwiHBI/OaobJzELF8Yg/Fhsi5cWHCfOZ6r9UdfS9VloaW8
3rozMuQHOb7ZffpOoqwiEjG5/iFOsAoPK+SHhVzA9/o4oEZRurRe7sVS/sks6w4CoZrxBh90UQ/8
9g1UJM75lbwzmlmZ/YezFY3LtedFUhQm2WHo6CDCsOTwm2lEiTbWBDm9zWy4oLYfuVVdqbBUDfpu
d1GG7VKOMb7M/OpL6lQXoOTzVQ21eR7g0R+DGk9AgC3sItKN3YLA755kho1Y8W074yMF6HH+ujDG
09BLHZU4eXrtnvknzjJBFIInM+dSi2l/gHIMWfPyXmBsN8berzmENMDoK0hiVcmyM6wo+s5mWQE+
GX7L1Gv2iYQnzt636n3OAEhum0IUCNOE1yo4x92MHGRa0aipwdxB0uJVEQ4+4gBMetFV58jXtsvx
Hl6CXgo1Q6DmQNwSCa1WfsUcViojG07qO1cO9k6L1wbbOcYqa3ReIAbkRLs2hprDhMZubK+rh/y3
I6UJ+DJ7aTZs9DgRIG7gJOoO9gYHwLpHhy30FxfQhrLS3DNhD4n+uTac9kxedK0gK92IRlAhiysH
GRAf4bhwAcNO0D9o67EVbmOZlDzQz3jUMmWl42W2U3eg7LAB59DeZAA4mO4Hrn8LbL6CjbMJhkQN
+TmisjryVRRWkJEsZEQohPKpJZ9W6iRpAeP7CFP/soJ3RSN/a0K4zQhKKN8KFH68tgoN3dBEU+0n
kntGye2bO9SvM0ffE0q9ryXFT7tiRLKyJBIndRnvbXTCuHeaHPeD0kXz3whD8m0y79K+oRUM4VLQ
d/Xlhcv/G/lMtxepM9z8nvQ+cpxpLUK7tpWyjoPPnpNp0fLPtdUnI7CW9z0RolGYRWnHfkJ8Scex
xyx3Wc3toS0q5hJ0L3V6XIK/dgCXPvssG42kdW8Xj/NZqdx1RHQJVaQarKZVM3dJ9K9vnNSZPEGa
4E4BLdKTelGv8fKPakjCzDAIWP4r54hP4wxfDlnx9EUZK0AcFTLLECgmwNSRwQKa2RA06Y6CB8N3
RPDEf628iNrxMahlR4Zbg1A4RFbZb0K3R2VHCGB9w05EoPB0SPIREpRVuzOexwqW0wa2r34zYna9
RVzmml5FDPkYhSEX4t85qDVeMj6fOvB5jogDwcdlXSsBFWMrHDzOOsPL0o8K70Ko1ivftnp0e9ng
lWM/xGwl5naBEeC26jNPPucwUEIF96g9M7a5D3wLbr1Cle+XwxHN81Ett+D++3xgaxYcbbiGjxCc
zEFExA/s7NLNheRBDJg16kqRSkjJ5RDrqV+v/AQMQPaL6qE1ibsoh7zlfg/2Cya+Z1zJpg8Du8yB
GO/DTIibzk8caIyxwlGPtRIa+Jltbi3GXf0ZxMNRPEzVA+5/n9Rj/I9Z4x9HlO3sFOeMf6gAWZkm
B375sqDiRbuybR4mKy4KNFFNt4pRxEa1bh/mc2onlRJ/loQwoIofR71FcekCiTRqmDnMT7nbwplA
Tbafb7oknKgdB2CVyKnljBFZsQJDjDNWqqZFoDoKIUOEEfbPq9BjyWrrsfhKwW21QslpsSc2sR2u
z8AZo2IXblZSifWfP9l+WczepO17C8eJd1UaV1od3skDItt/Vz3YuE96pZqrFAVO65YGBMUmkEIV
xCUSWfpBcLHl3xYDFUJFXFEPxJ+1TiMRTFE/NXQanQmJEKf+f3rp/Zou9LEtXoHSH560/+QKeHZt
1RZyhtbX1tA7atLmlYaE90BDZ3RbLBqYQ6veDGd65hpAzIzNqRkbYToM4tNhHUuQ0qoOnfe5fgcE
hcKDtfcQA41Uhx8sRtgXFd5VJQAqMsoa531jNpz7r5jr5HJaQdM8MgXQ1KZpDDhbQ0I2PgrX8twQ
XYN8tOfRo54sdJAmHpM1Z3nvxlj3x2k2J9jpMxrA4oW1kS7W7OKLEswFmZTLiOOpPCZOhPjzVosO
u8Htc5PWmnpLoTKJUZqsiLvcPrp7iQGdJHzN0zzLKEbcR+5UKcal/7U5PPqySFQUOU1TWCvvo4Wa
5BBc395CSHL68tlqYq3svon0O1sMa6U2BGVh3nDBAHN60JJtchi03vHLCV9gdkylSU1w7nUiaAt0
nWnIrWZvZzBH2cnoNwL0wV1fKfg62C2BiFyHm0DfRAgALbC9jncoXHeffjFOWoQwY4qwAEpoMfXq
VMvbq202NOgl4H7ytQ0t2eGr1RCQfEhoDbdGLS/BpvcwbIq0F2CSgXGuC69xuL+Pfr/LjJxgrMxt
6Hs2qGVM9ZhZ+lZ782lGzZFcHuJc9UyHzTagSOHYBRCkYw98uF7GXJEAaogWwa30VLld0/WezwV6
bxe7GrqCKDk5OOmD7A/Q221Elr+U90eLivOishXhCQIHXlWU/P1yjCEBoSyYntuwBER1CB7WpGlQ
iI2pEgcYkPG2ff27ulVyZ552KvH2q6NAsl74mD/9hQOJy7cUQYJ9h5Z9Vy2aI7pF33d6+NyuMVm4
VE7rpSa+6lbcwAN6JcGbNu6KTe6Sah1U4pw7YV9YJy1ryvLuKJfAD5Hxg+JLYl3LRdTQOdN71UIa
cIJaASigPTQoEKn2pQonS52IqeKmQh2nxhTV7HchTkhy4BLBI33pqayuvkoYxrcibbCwAkL/dBs0
DIFByDhNX8CfS9VHR7IUQe1nIWpLMzrTn1Wg3kEZ0xMl5g2Rz8uWWB6QS4lZddYaKNK/dlmaFcU2
3CB4zsZuN+qTrgkz/QJV0XrFEdccmREU0QSwoKKqaH3AKDewLP+DBWQ4lhayk5f8gqqlAah4fL0I
wf8YN4qdSUJ95fq7OvOdcx8UriMVEW3cH+Zc9Qi9+S1B2B3huLdvwt/ffLDDk92zVIKmY9Ts9jVw
3Q6zMQEiwt+4OtP1oaBSmDvc8lmQDX42MSoA8NiyPCgnPF567vUZEuHMMkFDnz7Us6+v43nLeKku
VCJLdjhdyXZlGwZqbSJpytu1IFge3Y4h5CZysAFt3Nf5IiHzj3EIz/WmJDu5FEb70/BsqlzG5Nz+
V29dNjmuO4FCltghYZJtrGdwwEYLOAEMI2UjNqcHg+SvHwzWXYV33fJ4nNedf1aCdJvHm7r2w7bp
Gf4rjzQqgCVhBudjbnd7MF1Px/mo9iXvi4SWSmFEEd8vpneRHyOvGjjF10zE103KixFzPYlyO8Rw
IMTk8mX2Shi751SeSt/DrZBKPrdqjW+Ru5fUWu5TrxLMGHOQG66cWRzyJJZzq6Gv3DFzi4wnH09t
asnGfz9l2klwSbfSQVTXq1niyJTnWXIBo0A39NXW4LZr8zl45TOu7DW4OwYu9z2vO0Kgf/LUYahc
uh2zg1FZcCEUMyCliXZDbrJ/SyTIMVWCfDLXvxNx2jdvJ2p8v+RpSezZo5U417+tioWiTodE+ICL
LxI1JobjsrdktjwzStbjDYgWyB434xuTRBpCqErLQm4Ze8oiExvf4EDGNW+X+e091kENVEWufWgD
XACRytzj7C3TKOE7FKOw2eijWWvlMcA+GxPNmHqxhTktUPs0r594GZCTYI89nWRpd12Uila7PGrG
eVAmqi+ek+TRvl+Jn/gZNwPpfNGUfOF9Df1EN/Sbw6hGvrfmWoKYEonOt7kXavqdgQjkHGDVdNSx
hL/siSsMPQ4zeFYRwgHtQm7KTwRJCOZTkXMEUoN4mhWiACVPipq0lzUA0MLSMuq62LGcZXS3BH8t
Xvr7smlg2ZRacSpe8XO4YbYNWRksAekHnPYFqjFuhH1cMUncrGKD8RS3M8TXqOTHZQ0MrcCjRpG4
9XlY2fqMtUgxJlaaOBFyAG7RQNMAiFdxD38SlEu/ir9ydG1A5RrwFtE8DhlQSLC3wvODEj4pO/z2
IrtPIcsaKZuwI5YZbpnXI8yqkUXf0N7LqRFGzbxvo060rPxcMbuFmqzQXefl8VIYeFISbF6OFoGS
60Vjw7Xd3wqoupWlhakLeWbCIMxEVW9KdWeJz6nJvRU0WrHCDqzLGLwee2MbW+Gzj3uSYJKDGKno
WcB08/LmLvxLbyzIwv6ryX+utujkVMJszNE4tJ5YLvz1TmdDgOXTQS6vHpMJ42zMC4RTGcyseIZp
yDIzsM88V/zl3ge3FLfUcf+5DluBs1pbjm1yEXwDkmanucy/V0ymq52RI2oP+7X8oxo6LII0zy+c
s/ZK6O5Wx3gUqUfoWK623nd1BgsLEqXCz/16pqQ+Yl1JHonaRHIOErY7ty3qd/XOSaea66eft0y0
2WvMih9lVYuw3rYWpaAHz9/j4/NOtUALcvqSRBcZmSIxHZTfSGt0L589yHW7gTU2U1YjrTNFlO1j
+vtoTD4zVCXFB8s3y2eRWgqzVr3In6iqpXfesDBUOuk6K7s/qPWOw3z+X83yOBcYaQ0oUHa2EMbR
NtlK5vla9Kok8bhSPjEhiKXw01XiIZkJUTus++a6bYjPg5b/d2rrjbwkpFXtUeGcS+PLhys68IL7
8ZpVE0Pd/0jXOj7oww5pFgPSpZGE7QSeCJBRd8nIKqwPR54Ksi1LaZ82+GHduQLqiTuNdrmbNqsA
GrtpsCPIx19YH9oOThgJd1sEP36fGexF/WUUvBLat4896zDiz5+8LUctNKSK2MtuMOpoAYoQZ4vY
MF8lDhNvvo9thL5hCNHiWA5myOoq70zhSqf6m+cB33f0f8VVBSWzjJ4Fkoo6ej+xSu6+grNpv6sq
L0+LKKpCPn7B+KIEo985CpHguvcorZzgb0WwCblSpjJ0MfxXHOYxL9TmXnZ0UfwkIqHROT343pqj
W7PnSPdrI8e/OROq2+srcwXkvTglw2r3tq31aI0JdROrIGdu1+xQTpC3tBgFQJy02uRrYkIZ4hMa
0YCL3dwyYgYufib6NDrm3Mo8V/rZMr1xN0yHtiljSCm2L3grbVAG2vS9c0ec4Qb+dGnAXu16+QM2
7WVFJ6dcrrdb66hzKSsz5C/cEwHhzwcCNkbMwc+PUX0OhIx19sAOd+/jgBqHLOXDKwF3bXcXGJF1
J+EaLshB+sYnPB22wmRzEo9jbnTeZDj7w+qRtSeaTIqIpmsxQVd2u9vv7de+vzV5jUlfR9DAGmES
WFVQuZNTsskCR9mm2koXHrq2B3fA16nNAtXLDpXLsBJlgNqUbs7rzmy3D2gxnUXAUNsQgDVjjS2J
Fm9cGxqLD1Uet8Pfkj/HLu05OHxiuwp78nXWUsGS26ylMDX8JEgMXOJrN4NJbWlk3Bx/RGRAY6cM
Y3TTBqw6zQ+ceTG5qnufg78erFeDeDcM5iZZ6xwnOprOf2GzjOaRZr8+hodbZb2bIs0tIGzri6o/
2YwTN0mKj6cY6nsm9sk4hMyK8Ss3fcQasX2pclHBXAmu00VSYgDFlZxqhBvB/G1QQPH3FUWrlrkW
eX5f5CiXrHvYd0xs9LtFoJzNCF9hF6OvqObgjotnU0NNMBi89sXAtgVF+5rzNiVFENfm/VLhfDoG
NNvmNZ0FzhSIW6V60f69HWLHQxKLtxVMZR2OvU3eYhmNSNVpxdYp5rnqZt3JJHKB58UEs3uNaASj
oBsU/HUqcGOKAgSh6uxPX1sDBRdsis9EHkaL9QskvW7D0LWMx+YJWA4tlD6C3qo0V8/FofKoj8bF
bvDhRS0QeQ3WKdxR7I6ST60dZqsBQFcR9zuMxAUl2HljPI9CLnlIyzd1pOv1u2REMvhl2SEB4Rn1
fFiMm5K3TQ7EXrDdIj5/RPsPTE2KK1FXZxz7V8xZs80qhihhxFrwn3zxnUlyBIVW4lBNYx8jXChg
a2QBKmVeL3I10gXotPp+SE7xQ1GBqP+e9ber/bAYBuAOeVR9M2/83Yu5vPSjde7gFV5M/6KOUTjR
Q83ZQABklQkHirZKIJoas5S07PiRg0h5AAt1a76RSMH+H4SePAlaKxazlX7qhT3x++uOZcub5q5q
kU1GyoLAUj0gklKuO6vYyArK4SVJbriCvPZlPCQgXe/xQJyz2YLOSW2CA9b2wzNOxr1Q3fKUKp2l
1DE3ybHnVufc5avP5wn1/TpKPUkdCgYsxy2A6QjT7Hr1dYHR/dU7HaMKL6sLM41XL1/WOwY6dMyF
oDidAZcgUtV2U5OImiFcFnMDKm/X4fq9oDzkWl6BnqYmp1u8jjdALtpqLF5g+FkDx/9Ur1gyBV7p
dFTgl9wka6zG73jftdjAKlWbPaN7HxQH7u79xUHOJFKBRl7gVR3ZdCWmKfPblSkBkeW+xogIVtKq
xOgoDg2ZsN/YcVhmJTw21oEABdsoivvIOfPcOxsyu0xHQAm4jvFJ8NlLWUzGuTasb/CUpvCGxNMz
J0KhhIESr/cqpzYa4rLIpm7RQwmo+73oGKaLBpbo0HtzWUqUiV1ikndAGFb5/JFcaQfutwhluEo2
T85eZGEZtPRI7Ei53VguUNsiAUzrKugk6F/BC7UIQm/eEKibZidt8IkNHPAHShaK+xbLJc1D2byd
VSxXnLaI+DqOwQUHlpEWllEbrQCSLqG0dTpLMcFsYBIeHrInmT1OGchgLD9X560rHXrYHscge6Cw
U7ToS/vlBh2epFYWZ+3oZWkRbVXBlYsnhupIWuQXDXy2bAAy2jFHfj6Hedu9m5uNvkBIjXM13rE/
uqpHNuaiS/alllgCk87pr7Dbwak81KOV3MneQV+OixhVvruQ5vClDZdIKRUW+gaUKxVOxCP7kFVP
wWAlsLIvdQmqlU76cKvepyv3kPYp3N3x3qKgumAUeXlcG6OrIsaz3Q60H/gwt8cjoSFY7GjAflW/
DUo7saDr0G/wMKZKTLcsOpJNXq1Gou0ySjoRvfEhiA96UjYhWYEwGJHl4NffJDzO23yDaGY2wiTq
lLCsD+Egk0GPy10DxjUUy8cYASp1aD75r5Fp2Gw/i6+5WDgVB/qYDbE5YtDCkJwsRhjnLpbokEPd
omkvBD35jLjC9dGM1rsQNho5XtaUrKe4bbXg9Hvu8uzAaNB3mj1n0lA0ZfCFIttp6PdlZhYOcIiF
b4xR2eO2x2JVZEKjhXMYtOJoiB3F5HZG/x4e2aJfDEfUhlgOcxt11WKvqQUCwNmeCZUBjeoCA+Rn
pBwcpsUoOsrNrnhlGHFCfQQDWtiBHgx3CzvA2Kl/Qk8E8Z9rU8xr0HYYzLgI6ByGsEgiFiHvC8A+
A3d0uOafgi9FNQ5EMT/SFlNp44gOOA43NgkAWrHEKgthk3ZaMpVRv/DjBEqfthTcYfJhjHb6/Kmz
Ib6TNCRr9FqxGLEhbRT5gKfgtaYG31xmNHWTG3dAkEoXmAtnhvuomph5vyFeaOLthDMvk1J4xEh4
jhdHTGM+UDvVuvC50wcohihyM1WVZAdrcTebfVB5YsXsPf21F/B7ZpOXnj4WOphIx7+2jDbvgeip
fRrigfVCTW1HbrOl/xKHcpxbujpswH2wMCYDGSGEaGEbJ0IIq2rC2GTZKFFw+GIEUBCymGtZqpDe
ylHV7SY21gMoFLGz1R6XtVnYPw3JGAc1SwOJA73ajgOxbJ1GoIgBJ8np11wT4Ub++yLjWj0Q34Ok
HHsQojLkWsfZD0NQ+mCl1YtBymAPd0ZmI+ZDCMFI7js5MO34+e0CoYw5TnPgrsyWHGZZKKM2+4U9
nR/XE8IddS2LzM/+UAoGGWOz4bbi17WxltR1Fo6i+vbNRJ1roQQGQshryKdHsbQBjUrlZXjaGGSr
ap79ri1TVzS4zNo9lEsrO8grCe61FeZsgil887RhAKtcs7eZoIGc8EnuaJm8chnVGq4QY9p1oIZP
r1QxzYkjSrDblsYWVAylrLGMEqvjCRnh2ErqFVOjtkJpmaT5fUzDrqZal8iHgWAyQbIDp0j6roia
6RaKIwjSUgQ56AkkhGvlSTULv7ZPSE0eBHFMigW57QST2bbt6JQZA+0uzW3lq5GcHaAqOjeZ6f+o
P1eGPPhQfudyzNcW/6ESCSbhSnsTGpNPWHAlMyJNxqUOFREEwF49AujkNXzaDmU448WKXnkaZZSZ
MTSWCADkZQ+gzMXN9m7pCZQPDupicbAWorPWfOzgGOUr8/oW9ZTm0ztj19rhe0lhx4/CYpJNGZ2U
HERlpyDRh/GgT6POQf2/w1g04CLN3T7ku09IZSKrs84hDQvb3QtiiN+1w5AtCsex78WHfjtkV0iX
N6/D1c581QAK++kg9DlmNgX4SFQ5Ex0/Sj3llEdz19nCy/pA00hIgffEqyhOa5qqMaFzbgxvQIUi
BZpanVXcX/65Yb48BpN2SCUYQurvGlCvzXOgvCS1Fj5M/ce/CbmLrhuw4KprZpTlROG0ZAgyw5BL
SYsf7gVCw5huqkOMfIVbZMVSgB9Q/ZS6QR/Zk3iZy2WqTvGu4R/RGAzZFixbpvL0MPgv6aCUxyuY
0RFyTc7fUytvBenFgnhm1QKSMOLHOqAR9IsPOcn8GCPj7pz0LfPwiVmby4RnwztdRAW8vJE2qc86
K3lJZOfrM9PWPO3SGMYMDUZxXuKZ7YjzhHHlwIImo4m/VZilgbV1fdZn6YU+gpluS3MmBNCfP1Qr
Am2qrbiugClG8YNrejl6XnudTuswf95R2DSUUrR6vesVsft/axCl/t6FfWtPgLY8VlSTbQsFgna+
oLjdZrThnWnJHKPIdrWFSoGe1bQsj4TdgBjyVa7nGTuIE7rlHSm3sQ96xUJHxRYfQ1366TMxnJEr
v+W8acHjiQB/uI0MdRZnNmO16Jp+flNDHgr+RGuoWZEjYvCF3fx7K8WGru6WtjNa+Hvut7vLocq/
RfImboivOnFbvistAt3JN+Zg/fOvtx2bbwXk0k1TH9VCEypcrWciAkRstKYnWGkV02aB5KF2GdDv
dwaLpO7YxJ/R6tb5ggaXUXBN9WDfSsZjPpBaKphweeCsMDEMed1wBdLCqRPnPWcT1ZY/2sjLDnt4
cvuFUK2mJ3TQLUj/pJrdLkbqZDIoiWbCfndyo561ax8dOIx80cPsJGQ/Z/nQsjMZO2aF+LPm1bZu
AbQZD5zE3c8mGQGfUqbZBxihPKX/ZUQzkXjX8cjPAD3iHjbmuHIhkpE5n7QfzhN5I3sDD50Oz1qi
ud6bmJVRx9g9E/udewOKqq8wHSG39Ts6u4AD8XbvnbmZ7eQauOQf/Ansl7URu2fbriecTND5Rpwq
O4tnSPDJ9JrP11ezvh0if7WVGNYqVaCkcGO9ktNpNvTKLYXbr1539Rjr5qqjdFfmqui2RvPmN5sl
ErGJNy7yXhpnyw7ZwTR6VbwL84rEySt2uNJf1J3iN6K4kCApBFz+ZB5EyimmI/BKdACOzBT6bWMa
4xixFOKLNJWZDzJ2p1vlvQpv3GLYluZXNavkHz3NuplmxAbEq7+PrxfdHPoKEoPhPBamagLRQdCH
Gyyle8XUXct68WgCF7M+hcFfpKLRgL5uqA61vbqq4USQ/xirZ3XEOsyBV3UHIRFhxk91xhuPDFtE
iLOKaRmix69l/HV1PUZFPaIhkV/TFBv6Bq+ax6Uwk6YLVwe/Lq5ujt+ciy7hBBBMGcPBMqFSPkGw
H4W4T0b4QJqfW2uykou9AyN8m0T2EY88Cemx++vHN2Q7DOBcmjCRLwtNbyAkFq3EVF7nCom/99Pc
2o3pJ7MxOKukVyX44Ej8TgxY+K8pgG2K8UHJHp34hMJLGwv/wUmU1EWlTbQF6uG9E7606lWdRYHz
yLHXzC/T3pdi2GxdbIae/7oEMvMG+ztvHFi2do64LXlbJ8E+U7sH3Dyeiq4Udz7dF7O6rmF+XmeC
YRKpnhAmqgl4VEtdQsrxAynIEc697VQpwIhgzf1KiFo/UUBEm2rovA8sKZbVUsJ+JBPHuDN+QR0G
XYmpcWdRFmIz0YoUD+jH7v1DTQDpU9IDXxFvuz0FEJUr3Ng2vScVFxdwoQdYY7Z6tjzwD11dceRp
66uSbot+3Te6B2MniLIhQTfuZ39sTmxqvm3SZiBK9KHK7sv+4zgmI+m/tqCqfanrqqiT0Jn498vq
4Fiq54CRJIyewKMGgOoVXSuHHW0LwnSg/joi+dLahHr61ew4ajZQFybw+WW+UH9+JZFP/vov+f3z
rZQXNnrz/HXebO8Wh7qJYe0HV4RCRmUosDVYMKQD1yk633JRIssuSWr2+eMepk+mC+jdxWp3KE0T
hVV3rGZAA/CcmzG4HHceVMuB+ZzEbVysUsckABm19fo3NvkNrqgfAmqiGTVHYGuQseTNnoQrXqp5
0PtAACClNoidkV/WE6m+B3mo/JiLhsO4uCkmaZzkRU0fkvi01UxX2B6a+waVUiAU8WewnXBG0NPd
7PYS47/eJFfaq6UoVkfjgoTzNFamvcPDTfSC9XFaiVs+UZnPR7uHkrb055U+t5bXiK3d7PeyRWKB
LZ7wZWfgRQpuvnRah0Odp9Fl5EFZkq7Jfa20aTSI5HuLTyqG+E+HSnRglt0KgNsP1vot84eRSc4X
m2hNiGhVUZVn2uFLee9YWxfRXZKSWVlAQPAx1LFRmdegRFokH1TIA+zTj4ZIwX6pUFhE3+VBWG4Z
knXN3d9+hWhWrLdVzlbMnLo9Pu8Ui4tpNCQGoyvjTV0L5PYYHRa6OP/LaCH3U5jBNKNOf6b88oec
n2YMzb57KGV5L+6ByBdqRT4m/VN65os4zBi1oOeTzUsE4+wDTSAEgoFE++sankwucwAZqVh3RYmB
Cfmv2MzlFKp2h7Y4rA2FQM65georut/frdtkQ4C00CS7LhYjs3VHUEVP6ySdJSbB3YOEVxx9aai7
0vr+mnQne1o50CDJmB7DLt2UKHAV9DkTjzw1Bpkl8Uw22K0ITPIv/lP3c536AsJ7upK98Iv6c4U/
z3XCwPq5WVjMudNuPeiZLH/GVfnVRtp4B8lBI2QfunB6qVd+r6SmZYTlic9t3xMAEDvfxTwObQ4Q
axnANA3erDvKWl4ZyCd/5jqCfmhQ6bjrkgH9UmMsNx5BxKr2SxFLXB2067mmh6Mr9CIJuGMuT1/I
956P+exjo9RT430BqzR0t9MbTRRLJNuP+OQx19kh23pBZZTOIENPK455RGXxPFLkJrxK3g/SZVda
bcomhrLz+0K8vzvywmNnUzc1/9Cr09nFh7+TagV1oMUy1+PmrkhJbJFV6vp51I346ZWZgtKWJ7wZ
xH90fwbwOpz8+jLEVHMhs03mVefs7w/aD1498kikzqiVUpYHmwKU9QkCG4Iq1KkXINA0L2I3YJ4F
rXFRlH+nbPfnvRYg34/iMvv7S2dW7VhFtqScshaOAXH4MKNtaTap9e9qMkf0dvCj9BdkjzrGE2Ko
ldzIpiJXHGxnYFriflewpQ/pnPfLE5G0iFamMTcP/q14tJmTqgTjlHC8CMYj5vxsVAhTjsVPQBBn
Jr+crJlSZKo8ufMT9n0UfxWWeXAvOyZj4lnH9C7K9cbV+ngmQ6Yew9Cee1fcdzTvQ5QwGsK0OKYk
td5AS6xEkUFGSitjphQD5FLTDYMz/r0AK5Mw/eMq5QLu3UJ3uWva52C+xk9QgtY7YkJeUwkjqbkF
nJW/ZuzuzJJJ575gbxiE1xu9Ct32PAtFawilBE+e98gaeWCbEp0+EdMtXambL8u/P7nv0YKVySga
DY6FoZ3Lx6PZaUNcYShjOp0znpp584qGw2I9Y4/SZeblVEfXYQrC2Vb+dnht/gcL3pFojvUft5NF
is4jNYIPVtpKs2aSpg/TISrtc+Pa+vIb25sHqPZ5SbKMI6lsES0yez1qzjraLjws0ozEaHOW56oE
DpU2/EuH8r5zEnC2HHQkarou/+dvMYLkHzvb0R+RMWtcB8BtzKtHk7h3XMPvKXT4mvjsqlS6YfIn
IRAtnATuiHmlY9TAgHFx5Im1XBPec0eNwt2Fb1cKS4B1lspaO4iqbL8UBJgmipcBNwKu8gzKCINO
esfh2HcCa/CuYyoJ0u67t7GN0RLOQf6ey8REjt8+/+vH0QIh8ALmQgoxAemmwAkahnqVQa5dTsvM
rRUjEXR+C2vq+4S7JEzznEfzX0tfWL3o4Zbzom9+dAAUPbLj6uqKt+n9BsBmLjeqdoOLt7m3z31K
GDIf7orI/BuSrnyQxyeDsDGkNhEIa0w1jiTdrPkShvh4evEvVVZGJzzv9xWNKXiZSNG4AZS3J1hY
iK21cjeEJNWfWwsT7qbxraG8VSMF4F9Q7/TcVG/hqpl3gdjG6sINKBdq1yxFv4qCWKruITWKdhtY
nS0yt7XcKQnOCvsAWv/IM0yJ/24JlAV5bpejL+g+443Pc/jooY/vRUKwQez7yF4Gi+puLKRUjWnI
lP3lSy6qTdx2KqBnaAiTPEp4jojQqit82KmHGRPhGfyvUH+6LP6oPPTCKrCco9AJgLikHBW0cPHM
GD0I1w3hSL7p0+jOmGk/aF4tQ1LVh+wzOkhxUj6FUjyiXOkf1SNkMjVjw+dHMZV6ZKkvpgIoVc0M
wj+lVTwxZ6hnWYLzI5St3BFkxWG6Ycrq1dz9KvEzxZ7KbaTHUG7Se2W5zU8x8mh4eBQBFw54UxSo
5p5aEvcN8xandw/OUbJlta1IQfnvb5npYIA32fFjwWAb5kLLQRdJJ4zOFkmhnozts1jgjKl8ZB4l
VMR2HtOro3pJt1EsgsD02UhPtkkzF/PWuiwPFSBy4Q3SNrw/5wfu9EPs6VaIganEOjKnHS9s7ke2
hw32BCirp5gkWGHL1+wxT+TMW4NZ1bZ8m0lEJStNpW/wwauMlKsc9kf8N3fo0PpS1s5wmHksdI+V
ndhJ889qeM3TKDXX1MOIBa3q3yuAm0e+Ug0TtHyMrlKwHlhHVtz9NgrfCeWHFBT1gIPT+diK0guW
FKneaoa8c8nH5qt0AbA/tEY8yFbuHmlCq6QxVqMr6D9BhwS+N/I8ll269tSN4xk172H77z1m/LBv
eBqBTBg0avmtDVUVNBPv6+Zg68ell3xUa+X980IJKjVN6DkJSDfMAfZJYLxjrxDWgRRG/cAsar8f
4PDvnvZXFoulxg25ALZTLHOrtExa7yOFPKAQIJ8YfCrLWKYUsbXub5CNw5NSwdrPLTNl4me29Ocf
pgO3LI6Qpzgh9YZ76K7HfCiCPW7nKPOjmA6b2UD80twOzgqkt5FQrNW+75gL8OX7jAiHbC/3CY5a
mvHXYEgM4Jklckgfw9Phvsv0xXq6g6FYdT8wlla34hD7CB4r0kivTo7ACbYUQZo/W7LA/ddCAU+w
treI+CjRKRxjGmD/KJHfXynbCuPZHniwN8QicikQTSP9z2Z9KWWeIVy+p3KB2s9NJ1v9S1FZyLIV
N9x28mX0Vwn23Cclv4Je3p/deSWbpb9sPb0tZ95z7xnb2GSyrDLZCtDayiYfS/BGtPCAxYGx0ybD
uV3OIUe3YKGeaoBLAfDIyytD+dMjClyIV8mr9fGf1ffnguz63cCFtbJE/bMKA4D6XpJgzKsp+mnf
b7KgBLONAGUmyaqkE2e/P+7oUfQNufMLCHpH1ze7xDGbWq9uYZdaL1cD6HCuD+EjPE94dCIO7OiV
OfrC8AdZSWnHP1/ypGy28kH7k7GCZ6OFuwUsRS2x1u6R4rTBP7aanOhNwAqg9oXXM4QMz1GJfQna
KCRFWws2J1UxPX8w5Z9Qp5Y4jP4fKxBTcDyxOnHONone//6ytRmdXadC5ry5cKdAP2LCSwtWWVOM
akHkGEQ4DuBTa3zW8d5rbM3ZcNJZAXYPjIB/vWI/UPS7AWRo9j9wLDSdVcdOwihNqdEnBBZ225jU
bxHTV8i3Wa3aRJxIRdZjtSpkIjJEcZ9nP2ybZ6ysboZPZFEL6j5x1Kppoi2CmRdoJ5xxByOk/r+6
DygCaF1TwMZXEPXItQyOU6BUcfAk5h3RQlOJbg7/bKeld6uTVVBNB1ILCktvhKlKyKP8o7xdY5PS
USftuHW5bfmDoi4IGo9vCV9ZkQgazbJRD/k0pcnNdk/vNgMUTNfFEwsfZ/0IDFoioRJPt0NS201T
KG2ae4bPtHcKXhUFAbHK9y4fHUtlkK/B5pAcXaObT92XK9MxkOV8kmVqtgYyCZGpGL70riO/Mv0U
8KmT4W8SGeonaJs2WMS6lU2NJeKPOkdtfm4DcloR+4rIArimHJ9Bue0BP26ka1QkBH3xJjg9pDcv
5lzD3WBRkIm+dSMNYdg8o83nzqF7OX8VAmdoQ3VV+nAlkf0li7jd8Uo88Q+scecoaAFu43wcv5ud
tPB1XFmxSfdMrmfr39It2Ia293lOxzxU8xqCkbIABvPwPtz0GgVTlJLfonoZGc0rewejBPwWN/O1
9i+8+JO/Yw+/rCuiICa9F30wfK3ZiOfLWQ9wn/zqfTQfgSvoE2B9t9Sxu2yXjfC2r1oYYezyZClE
4shZEy/82ynTFJo1AvweY0bpKlFHY7Dg/KWzGnOKoLwVQCiR7Rs9HlvETdqEmKxxgUajr1p952T9
ZzgBLvkPH7VZ6VlFHe54HeiOerTrzNc7U/6v7y8TVeht4xKGbYsIItJ1mwA0p1i7A80NyrzqJ6Mp
UqkFChcqEAXkKf1uvHFVlSGGGmVa2Kv3Iget6xZFMm3brMyzEf9wX2BntqFGwu8TjLltfj/J8vEH
xLrI+t/ejgPVwG0iTZa/icCwflWtyNajPo+9TyiIUnjp/vUHbKyeJzfiTpYh/d8CxqyI60sodGZy
rKrgsRSsTqcR/RqjGeacMvBjQ2qWRb5LK2JJy2a5opGPwZ3pjJmeXbja3gOkQka8eQVwkwBSD1X3
zJjUzV83BQm8eOi2C3UWH+8xDZo+x/kJVXF3tj2iFLXCMXu6j1O/pthJj5xjkjb8DsC5IZItFUnS
XjhiTiZ3gd+Nq44X3tBmavH8beUhjMkgtc+qhsbrDNwO8rynrfW7JKg94vY6p0OR24MTgQDxz2BE
lc08QfXn52E3f8E3pp0wGUwajiX07pMP0f86ied1rF1k5uayMm+4Kk4dC7NK9Dn3WubDMHCOknc2
3DdVi+hZDDoZcLBD9z3Qlve5ZCx7TepO77YW/NKr/Z30jCMgPDQood9LMt4iZDAjDz7LgUHCc0aI
qLuYpj+mb9eFnWHX0ZeI0fndGaBNRO+hOeTSiFByVrkjOeN/uPzYMfMXocwoF0NwnuAC91zNgMjc
KXE55UUUoWtZlbxnYnHIkq8ouYZTnG+JGQFTrMLNFzKVKO6bACQ7N0WXJDmMxdmDK0rKuDltj1m3
dnlnEPdKZEyDzPBPuVfJFqGU33jor2+2ZP+3ptq39BB53Ti2ILUnj3xycMvHI0q3XgNr4J6UPVRA
ibtoB/P99DKlQP6822DyzX4puqZcCehgtygKq2m1evqnVyQCmi+DnyotZSr4UB0Z8gafMXoy1Rrj
5lAlHgwnAc+abznbyJwHO+TBoua7IqVLv+PeJb8fdpuhoaN0xdap+badWrKiORjAEsqcoxZJpusy
44v/7FgN2V6HvJGXCff/TGWGLTPoryHyq32lkQvncrhHXGerqV5tSgGgLG/Qled7mv09kk/vMR/I
JcKHym1XIhi2ijaQLLficPrEchKHSLdF627cYVWw2XWLAQQbPurdigUUNV33A3e1FEvnAWJD2qP5
bUBDPjgnmj78vqEvzNkLCnnnlIDQnWqR52CwT4LCGHZOB3YHHd3nP1y4lZlx8Jfg4a3B/L7Ei62Y
F22YfmDS8VCv4D3fmAzFyvWHxAbPM/TLcb2Qxtkei33dZJjeq9FEXukoU0draUIrV8sjJRyRKEos
/iiBnTjg9rgd1iba7hvsNthTls/g/sgzAAe0630bK+vxauXCdw078dfmG3gZtSyXUN1xeIRJCBbc
1MD0PCy+tUhlMxBFpjInenXilz9viB43l6bRlbTICd1GAdEVSLkFY7+1vq/At7oBP5453GcizEBk
w+3S14tS4h/YHeqVGJl/YvVIVHhNp5ZCkwOcdL+7tEr5mfJiLDz08u65t5H3ACls34GcgB6Fi2rb
GZZ2kON1PpGjVxonAMNcPBGHJzWPAr0quuM2c5n7Bqkgt32ztP1eq6F6dpSTFfn8XaxVVuPT3G7U
tpW7IVLIpUb8YJcx/KAOx9X1+WigstZtwtjBbvR02bGC7GaeaYF2TEPglzTbbuIUpdbzfR84GsDe
USfASZE6m92Il6GFGW3jGBzdua7bDb9JEL9P+k2GCg6MA0XodiLkHZfXT1cOA4hcDY69pRWe9lg2
VgtJQ/BAt0HPeaHdiaXOI/Z8TohLoWXG9QptYDyrV8EstfzLMhS1HTNSYuA0r9ZEwAjN2Rk/eVQK
sYp4AURipti7K5eJOX7NMK0Wel8ng8GKU4jLgQ6pEMR8PgVFr7vY5jxotRYhsF8s3+NkTEGkN9LS
OLfbWAutv2hhMyZTRteTs6UccaESam9QP0ilI2G+20wdJD9Wqh3CvRU3n215qd9/9D4U/G5A/5bs
padBovr2zi9Sy/WK6X7PghK9klLf7u+Edrnt3HaK6+9oIjfPmKFkysWSPW3RDaONrcSN+eL3Wi6k
krmgQ/0WtMYoWnodsIBFIvg4m9hsk1DVw9vEitKpKxb42+dVbwOJvtoYaJero+yRF5TVLkPBXfGz
ZonomTqzNc5tjyitN73fHptQsRasctQLKQn+kXFHGKH39FJCvfSh6Cb94FWYaCwSJyp4SyrHshEb
+huXB1h4IMSi0+pchv4zfJqtIbOc2SyYLSzFBbI65gdchvNDtK8gGs4nSkPj/ckCc27WkUzSZOMu
WTJcLqx49SU2nDB3o92lT26SOC1KubcyNFrPxKcmqYcMWk0nMoLQnTEgtaAAg0h+ntw5optvUULS
wyKJGSw+SwNQKLOGNWNETeFd6jdGowOECnUrvaDnINgZLD2RztroXL9QbNrnRV2Jz6jW7+7lZZaR
ZJky00qNuQzkvmwVr6d3aF1pt/Y/SPREvP4emNHzdc+SnuMMW+8sXTxALkNbls8k9xraUPMx/Hs/
mLgXJTrDk3tfnw2lznBYY4xBRbZOm8913JHelxxFA897tpjh/YoiSYsBzLP3erciWchUZWoKqULh
OWrkYPzUKZ75ARAWHW/THzkTSK4v3kXTcyPix0rPEXjh0vjwOywl0NhrlBIx+X0Z/qF//RSU+Vvm
Awx/VjQv/w3XcHP4fUm681msGdAot0D++yVC6gHS/OBCJO6V1K9vUNjKgA4WnmWU5UU9kkpbvawh
7g+cbFg1GFLHOM5z9o06SWbxm843lIcQnm4rLue/gTWxYfCdJ7ri7CcjGJ3NULdRWqmJWqWreJei
QLlpJEIUmZOCzKlp1QhmvP9qDXHEvYe6Cl4Lp2QibLw7wpRjTbKrczIRWlLl8f5Tn+pTBQbs27JH
t9UhYI/7nYWa9SoHaD3z2S9PlDb6dj999mKrjbHC9fkVjbuUfFR4VavodkZmF1xZcGIC2rxgaQnH
JJOcBFEsTmNLXijaKR6GfU6e/7l2hoFiHTFEMrQrksoCCv2RTIrw7Wf+LIwhVGdAZMtXvdCW9XWO
lEJPLzAgwFYe3XYCZYK+qFeOhaQcxJFryi14dzU2ev0fJwMLN88T5oTlVVSDUF/Os1gybbVT30fa
Lr5vNlAMS0OYyw1lX/qHZpIx/h1UJq4w806+0yGgXg8aMWJ42ijE9dSVhFtRUwEBGj6Fs5QMB2v5
yNdpqVKsBXRrvxdCtgOtCYj6fOnr4UoaKO/Oh5EE8IKEsX2AsybOsRvzzf80K8BIiTmmKYKfT9hK
Z/vm8KZlJRs6kv1D7eOEunfdYMDNwndYcjUNx/87u03um5H2mnh/x5UDi/TqN3E85bwA4EQGtnxH
eZv2Np1mBZ5qEkt94r1CKbgQsa5cpFeXhr3yxnQFY+32VDuVFSEduG40Wt/WOTGiNqw6x+DbJLsl
6pww9md8cRY+9SPKfTe9A2UBd7iDm9gbyTFa3dGAIC/Eo1dtkTN6l4NouH6y92+ktY/xjS+Lzlp7
Jkjkvh4w5D1yX33bALSBxwbSFI39JGmimYWS5pLW0V9tZV3k/o9UierG7Vc9LockZ2RIzmzqAlgH
8a+LkgilUjXOojoq8IERpCOJRuyGYkvPY4xiz+vWqcbZog7KUOYClcVhSSXLH009iBkmjIkStJnx
zLIPwofvyUIvFUnUFnPEtHlwlbmsRXGWJK3hwiLrQlBgAHjGrrdQhMWawGwrGLDjgy1rGCBQnBpC
F4+Eb2UpFIc/OXpVBTsDhyd0vOg38xavGYx1jRZRev5tcJ3qhLvXc/86k59hWZG4DvxIrOmO4mZe
fu1/nXBE1Xvp1T6MqueAKC05ZpUVGyGFjooZocvHYmYUrtp3UlGmPJzJ9yUU1gc95hy31WiQ8roW
DSczoaUkF/b5BRxjVohX4FEg00JJB9XkgpHyExO06g7ojgOfPENhRhqMlu7z2S0ZnCQW4BO2x90W
9JWrHVcsCvBmUXrIhtUKHSXd4GkOo+i5Mo/VEqPorK56oo9/xBp1A4xeHK9qskuQHoCZc2F5JEHb
B5HYuvfpu5lr2sup/p6uKGepgG8uHp6234nuoo988iQdH5KZcyYcP56PRVFucqHkT6AlWL/C5OH3
6CG5dxC0oX/Jx6OV7u8q4eO1DwbxWePC3Ix3kKM6FJUqyLHR+k12ksu6hK8pX6YFbMSUv74Ly9ur
uUhQ8G5zJNTSpTaIXhaISXw6b+mfLQ8JqkbbbwsVaE6RtBwcobDxoEDZZ1VMFIP1FrxgysZqYGxp
rQ/4knNUNMhEWNkwnwaHE5xB4RDy7T/d5XCDjkAH+KvoFgLya+YMlfP7txn1GSqf0AU4nDj3MIwQ
TyCmkcL0gbpDqhTR/4igtoJiVYagp9lDkEzrNWhgXb7s8LvKY2carhRhVqeFhAtQPAf5rt25KcFk
FdxxOz4j802Aq/349AlD/Wwsd2DVT0Er5HYSmdH+LQmKF9GUDLdkSNo+FESa7eFD/20ktXV+50p+
MJ1mIReGiq5dvRMkbF5Be2E0VJ9KKdKqVVMMZavDeaOSKsQLchIV6DxCL7IVm4fjPaxujICWQpMV
LeySYv1AkQbI+Vwkb4WGfinZ00mhUMtzaXqec9p7QCnK9V3FzjCTilqKIigpEDbrBHRXW8DzS87R
YO2vVrRJsf/b5qccvjHgKoISpy/AETPGB1NBurXkk7OmjCsL/f9BV5uio017rR6rh5e2ofZYPUIV
0JSNBAtw18ANmd2NAz6pJHRoz4fiCsW9IlbDBgCJ4ETi2NQtVfrLgDX30czifMaRk9l2MQSC7LPe
brbERWMmWGgF6c0yJTX3Ig7priyKGpwFKqHSzXEHT/KNAPpPDyRp6Nbr1EUMi3BPwnM7vjAjKbiP
6S2/Q8sCKE19XRWt2OLRjIzpPal7i76v8KAtJbZjLKnPMPpbOFVib0GxChQW52zzpi2gbGpBxFxl
pMxipK07MX3FDXbqN2KuueRw43RIO7YGGq95HxB67CjJBbcF5t6t77Yf0Hp4PQ+i3dg+lk8OWQ2m
4IFs8RHc4B8pX4CMBVfNMxZfudfoQ3UpJdGT9yD/mShi4AVKU5WvDH+VpKnyMAQ5tCj2bMnXaN+U
xykN0A85jY8G9aUCAMoX5UCdKTUD2DuKFV0veMjF0ihybM4UXUn/umzlHN86kchDWNY3nGksmvpN
Ej4GemUd6FO+N2z6DU04jexEe6sdqMyAv39gcEZFZzNiBO+iTEDfHJ69KTNXiOOOhECahFIJHD0v
4gjZEXB9yM+6c5JG+FG3TU1MBUiYySgjNToOzfmP3mZzcsVaitg41zmiBJlce1r/gSRepbkOhngN
sURbRYANtOK1DM9OEjpfu7+wJlfaZlORLTRdBEawiscoGTA8e603Tg0VOF3n6LYL9ALDTWfWCufy
thQ3+X5HH5uagurbFastqiPVueT3xRdfLkN2qABciokjOMOpuJe3BiHzkk/q2BnkQAYMQrKTkiRK
RUW8A2n5tRS+ZhIzTtjed2zlldy4aQvTGI0elfzsj5GK23ER0vm4Yn/Z2kAfs642kmf/KmZq6vs9
mBKawS2XDOP6X2FMJnWjTkl+F+CTxGCG/2C4nYdBDtcgovWufCRMAQzVO/f7/uOD+ZREdTfUxdbK
scoChH+4LJi9s4JT9XajvNvGOvTHPbw6ROIG05PEBC9muCArtuOqxV5NxyceGEg8HQsRRFWrmkta
USyIZvA/mqhZ166vi0VoDr104ur43DFrAaEOCrCtDgOfrW1tSX1JBQu/ADtLjRSdGX64cfQ+n+Ek
+t9zAeb3KWUcVorT4FCpJKni7ka276dUx0u7P4q9ytHE9xCS8amqtYDbxu0WW+etNivbmqCYint2
wUZQc5eoydR+DHsG/lqKABcDH2lhOFghDMPhcIJrgq4wZTxrPdSEuneK4PJuhE3wLuJXHBrLwSim
rtCt7AIZnYt+QE0ISrOq5IGbNSkQK3laOVsakAyv6fiJbRaS5NJJfQXwhUl1MTzUrqx+5hMZTrwY
Jgm8sDHfEnDu9v/3myLxSyVv053GZKexN+p51QYUmT2qX9/BMV3SlmL1cSRkqKqvw7W1aF7IQd8K
Ukg4NM43ieexHsq3rYtoDBKX93W2UrkkTCy36hX+QKS+0QIdUECquXiK+ddqSlSFgTpOID2MKsAn
p7dUnulp6L9bQbMr1ChODEXU5NU5RgpfLVg8D80aUstbZ65eoXYWyRI1PlmOe35pzW/GKAbgU6mz
N/G9BB3P3DbiCjAI+V1GUjMq6xI/SGmToA8fHbDmDHsxCgkRaGPrU9xAWRw2/Xymog87+ABykf8N
Cktup9J/H3zdYxWFFQU6RBJlwYpoGzI9kg7NASqTgLv384D6n1/RVFyfEqc/j//OEoBSnhuzAAUE
hR3OmxGSf59Rs39CJvOoTnEpfR7lJp3dojlI9USNoUfPKP4xlRuLkcCbKFC57cj7LzpdwABUKAe1
1dgoPwT8nDwyw1cmqA90PCm0Dmfwqd+NeL94p9LxzYR9nzg1nTLA2M609VwLQMwgjORwLQh7S7Pp
Mw2OBRung74nQ1D+ilyIQSeJkzoJJ1eajXSPUHSc9wxfe+iaJFP9agkdWYEiMBgS6AqkkaBtBwON
VcGO4HeE7rj7aNfCej8W4I9+l/sYsKee1TRng+XATgJF/Wbqz/kFpkrNg+pt3KV8Vj/qfG+gC5VS
541zABg0DpOBkcV1Hi6NEDbcN0isTx3HcqIICY61Gkehhozhbwn/fqL/ozQUdTbTaHOoXY40Lf0D
cYJ2qegHogLqdQhiteqhF+WdpcmCS3Gambu7AKL5CtkFnmZrAZl3olKy4nm38P6ZPG+USsFhj/SY
cCfO2Au2KFjbzXlrzfc1AEhoWEbBlVPcvxITbuuJQJBajNQP3ZviYKqsS73VvKZrXmUVvkZMSqNG
QFYND3lvhlnyhm9FaSesztLUqnDwaiKd5PERKwf8VaH6+5VmkiqoNVF7CmufNVjpLZFbdhXoLO8D
gViFJPkDxhYWxKWftgA8cjkVvms90Tycn92IjssmXXWxfkzyodfg/R4Qn4Ceq7lwFJRRy+ShC2ML
QkTFsygIG6q1tIYioWIEoAqpvzmiGOX35EXNMd+nbk3TNcfXgaykzn7vpJX55SRTLhjTL0maMb+s
tEZ/xPSHiLJvVyNHKDofLKRw1T4zHQE0A9OxcBLWJU2mZN3LMxpd2IhYH7x30eAdWTrKdcy2Gh1m
N1HwmOpFBNY0jW2InDaCpepe31xbFrznNrCtdr+ZgNV7RbIIvhE2WmJLI4VYtYrcqWM5pEZ1gX5C
YRU6ewb76ddMOUaZwRLtlnUfno8dBLV8Y3rAHQWLxY211XCNCCy8HwiMQztN7CZLb6P/CX+ES54y
4rkGSiKl2P53gXGLCuuvIqxhm4rGXdRaJFfq7PPHNFXtT34XeAsdBBLB9kUuucqdABcGZj6sdX8l
AW++Pg/mGDYKE3Az1uQzqKAqMV/dHZdXHRvuiYfWUAdIswsWaXhtUJWVgTv8lFn3BHZqRub1uL6U
qcUcy42FEdjYwdGbJYpnAUZ2IL5mM+hR15pXYUeC6VcrRR5102MqzKxNtk7s8MN/NJ9wfDhkUz2z
3RunX60wUg3yeZL/+TMN58UL2MIGvczQwXGO5oTexSnk9t9Ss/rNkCv/L2ZczV9wz+QEggYM5aWf
1PrZfHguxXTsrhD5XSfHQpLp9bdY1jRBsTf94V6RdaWQwvIJrrsg90bjKbAHOtjwrvHCd5I6+noA
yCsuuKQm0zTIoz9nzSGPoKVx9Px7fmIzZoqGrAK1IrmAYP1ea5lP4Rqi88tyJd4R6y55ZzdZlK6Y
245psmTY0MJs87EhplJQzqdQtTsHzeGORzWZycqTdfKY1weDoKdWrqKImFJ+1eE2X9zTdetkYAd3
wy98RsVIJyiFRVrRKlN1WGGMHOtIZKlix3ehxFyvf+IUuJqaC/NhU0GBwhQDcAZTkQhRv+kzNH1s
M6yvplYIjzgFNjwpLErSFfFMUtzgB5YX6Rhu7o2ZaAdM+Kxo5Clu3c/rO0+yXcD9uFNCMxMqMAx+
KmuQlCSWqMAGnUbdf0KXGR8Z7nS31uZGgv5PWd4FnEC4xfQxmSP3UMDPGlNfF8/VGIICjbyYZVGn
d/4re3NSElZq1JmjxtcWmH2ivL+U+MPYXHimhuc1QySvaFqh9IwKfcCtGcxvSFb6z4RzdBwuZnou
4OrlMOsaiDEUZKP5i4ci9LK5JgK7mbdPMGd/qSH+MDnJI3ucg3J/BRQLcraoXou5U1dDp3Hasr6X
CS00ApYpACXgUKH5bRS2kR0TaEAYNeAfBUC9aID7QzYf7A4IJyaqojk7kLjziuhCCC2bS9MdPO+0
UUK3L04hJO7AEadlN0T/wOi41jkqoFgNbNvCvBIyK14JdeU3vssyT3J5l8AFzkFqyIcYRY3+Z+Uk
BjGEs8BsP52x00m1CeMHANzw9/Bqx9aMXh/lNuA8Vd2HZj4gxQPnasr33Pf/iIiJGm5O28zDhVVh
NfH398n8W0MzO99AC7kh+hcQ+LD4eFG674odpO5OWUyco73Yh3nUsTQVUW7MPZATGMKhecBLaWJv
tHu6lRWbevLR2oPBZRsQy8TcJoep1l9Dxt6RjwYWnrQbQebqBXchzm6360ZFpZWjwo8NkQLN9Wi7
G6/qEqiGRQjKPOgp2UUErsUTbfF1haeqQYAQt12xSapK7mUFHdbnNlABPYv1MxJ09OhISrXbT2Sh
eW8V+OsFCwDa68KHWL+Nzxjl+zMxuORLxk3w3amVvk088gHM9Y6UwMk0tPyvmlrmFj0aaoHGOYIE
QDDT1f0ERbAn3afZGrk+C1V8fVxzvvOVgZjtaDZe4/dl8jyrFdztHG525a7TsGUktDidIvK4DSJb
v9P+ya3JCdFhhLMba1/lErD6yArdK7qoztMX0IgK5mZtxW7WGLVLXo1Xsixf2lgotmjhrFFhrWkm
C4zPrjsQBL4YFO7aR1PYI3JuydPxarEtj8A8Y1XIap4fA2tBLv1SPlK62ZSeYXuntE1ONm/wLjmZ
RGtgGVvaqPMN1TUKpVPLY3v0anc3EQ9LfCe8bRJNvfa/wHRNtvT4m6yQQ5BgEs+Xoin/wVGSJMR0
73gakVSXAfqb8R6jNqLrdPAw/3zMJUFzFWE16vaKuKOGVd4TpCmB0OCcy+FMMQV5x5I510N3uJZm
cRDRIF3ZsWZjTdiDmqbaTRvm3AFPpx52WxJSeHGwbe8B1ppH4SOJQG73m2cheCMfseumHVOa1+ns
O3vtfJR+/TpsWp0lcGm46l1PHnnruVxaPHtz8teOwJUALf1LWwT9B9IOWxIRpdzMC6IhG1h4FcUs
JNC6ZdZNKFg+gyQ/1f09hrUyDxlwJ9ZnVM5HZBQMFxG9p8Yjyu/7YgGl+7USHj2pHPWX18r9MrLY
9RLL1TWW1VQre4L5HSNgi6jXSbMEWdCIXauDbDG2yrN9nACIL7ClNH4egi9lS/yl+HxagopRutF2
NEbjUJ5WpdWsak1nVrSl0eXinhgnJISuqkOOMCY4zW6qVch/VEwN1BfjE5Jefg6k+V62dHpXkbEC
fYTmEsvnjgMfviff/M4tcRydLs3vXUkPCegxwP6QG7IOQGe9A1qKXyrrd8AX4mN/rtASnwRLX537
KBlCph8MQMHtSHa2Mq2Ka2LEDc1hfuUE6AcY+isixAc35t6ym2FvEWsXR1t6erVT1pWZENFLwc7j
BbWp7CXGf5P2EP2tdIga9ldc1W57FUg4GLrdKwLiTNIriWKqFxBWiFtGa2nyfqHzeyVsGn2roU4e
ZvBV1LHzgRiuCLAIWsZtsvftYk0a62vYBOh1uVIFfORkpS4MUuYG9ZoJh56K0L1CW9KE7iTf5UST
NLyzLE7aMbhorNbPc+jA/xgnqO5/GslDlg6ZOccouY4ZFBxqlLUo63VisXMHDmGk1t0JCyIYdZ+A
hFaJ2iTAut6GAbDNTT51HHTUIfsdWAePi8WUATKgeI5mn6gzYsVLq/bIt7jzXBX0o2IeIRup3LVq
EZc6SHQ6xUVRCWbPTkN7aaUa2fxsnsQ/U/rLSwYiuh53pZBua6AoTld4vkh9LY6YqfdSPGFv3V3N
B1rrybZDGUqngTJfst2RPX4hMOXJo6cEFHd8GAqdmh+MxI50cOiAyYAIomqVen8QUKJlmShChudi
aS2OyHG+8AmIX0LZv3/c5ECp9UfeWhzA1hZ60Jb+TBp6ljNnDRSfaWX7U/z8Cx8M/oUhSiRO2okb
jdnzqD53ex6TLiMrVRiepQYho/Sv4osUl1oVVMaArDzC8N1uPG15kSBY3vohI3CwvgoT0aiRupit
evE49sw5DEx/Xfwa+TCf9I5GO3vjMKVdnmeYOD3XL+tlv7TittOaY13NkJGMlxbZ06eF9osiwVwK
5rKrGInAVFhcFAqQEiRNCoazXyxWTiN6MiBkwmiv87mXx8u6BnaybCyQXI/TCGhD0G3TNBoed9Yk
Gx/eMgJ4tYNOc1Ymxz4fO8ZDp1rPP8FTIIZZZv2oGCebUrXqmsADer9CbFskA/1lyaz8W6wWCZgg
0RSPx+rZRwVVWLr0j3tMfPo5c42guxcl+tBBiOkPwCJYlg1SB++66L8zlCTzCU5STOnV6IendTH0
d68Nq1OLnu6ydbowTlQcIK725+a+Huo7CTyfnRMq3+1j6CaA6AXAyWrqzIObZqPmQv40GW4Vj7i8
byJYF1lTmqC+xiYfLuS7SUhmIQFQfUX6ot7lHNGOoe6jQok9lYhwQgtXzymabKmXtp3l3I9kyeM6
S0FxByxfAolCzYpHo+X4KOwzV616uAN4xEQU139cu1vRcGKo93chXYJHxkxBLMt/lUQ6QE90zN/Z
WVuwM1Zgzzt44naFunZ3uLOPGb/7TgWjX/7WLHhTwO7OrnhE2fl6z8iyK0Q3nfojUON10N2E1LIo
jgnnxMncBf/OsPZFv6ij19m65Qwl664o7hCFPVn4LiQ8L02O0LVwGvOd+1+PxNVZC+Rand/eo5KI
25ycr84bq6xrESO7zKosDWFPjZJQYF3uzLoPlIOtQSy4uhnW49kzlrqXPWlyTwknsmW0Jl1/fDYE
88PEWslRJX96bz3qyEk2vL1Dw0uFFC98lUQ3WqMZmwLoypdIDSX3+yXfv4zj27L/OVLqJvdaargQ
m2Qo5mr1ExnTqBEF3KaQXFHt9i/PR2Pia83vHa+Z2kXKVZX9Tftaufw0dxz+xOHM5DjDdpR53b32
Pp8gYZyzSoNNseobLnbSj8Z+jf+iZpAS/KaEH0ZnAdr9qGwisoPXhMmzCqFpzT/FitoPzMcYH5uj
NVAXmb+U7eLoFxv0DvGMgVUBqDNaaIjVHnUDnqjoCkDBFPRelGXTTOS2gv/3YQRtO+aZOO5CQwW5
f6h1MtrBaHuwtY2A0nJto4+ZEaxhnpawy7EZH/nbuOCR4+b5oZlNY/+9JJuiFKNryIeuEifgKiXz
05KnQY6FWqvBy+9TePMQeqohJ+JMh7nqIODzertce7kkALOB81T6mjJSJMjjJkzmhjX7JHCM6cEY
AhbJ4+3MQ2DEod8nOdEhjcVpFUD6p5Fly5KyVIJBdfnK5HRPjfNGoTDhUv87NmTTabrGRvKgIGRN
c8byW/xbHA24eL45/dm5IidwGCXrjGBFEPYeXp1wUagRdIbe4c0GZ2VOPfgk4L2/UYD297FAZ/mR
OSs10Fxco6pxGEqNX1A96rcXJvN7Od4Ga+cIc6rCN+3KEw39ztnDg6dWeIUGEiwAWqZ5sEPda5Zb
8OOjk3CFLgVASL1P7t2CV+N4AvuXs8Uub80KD3mTsHWzVlQm7LBogHRyEXWbD7yPUbDxtoyth3uG
qYg4DnWY0uFpy9QmJkcq5A7lWxGyES3EvxGDNyPmzBeEPX0BHq4m+k+mXgHPOHKS1DA6v59Nfsh0
9gEOknVykVi2qz2LGRsh+RbKYFJv43RhHnYi6H0bTxFsRO5utCBlmCV4baYyPai/LgO0dtvQGN+L
lF9svc7gySMZ1lPo/sMByD2SLaYmRlgrX2LrkzofUockiRolS4jqFEoeo1pwHZd5zLgmjVI3bo5J
1f7RHK/3Ci/WN1y7tMIQnOdAenqEr/sPsWPJlqaq1drrBxkxU8L54/FkFWm7ZnEj/IUtohk2qMaw
idMomQLWIgdrI5Z9bHjZ2juhgW6AxbhmwTctPFdNwd4HyzGgqGef0uMu82XPdLNEbxVtZ0R660t3
MelUc55ikFeQf2/veNmddM7tyS+bhx/kvMLBarmkqh77ECtF0FEF7HLVssMpesIcccF2DW1rqmOY
NgcsG5Cf03lF0vaSf7rqeyTiWeqNVj7E7/0s/K8kGDrgfbQWyaEz8TibNpodcTt7GkWSIUGKU9Rx
Vg/Yz4KBUWgCCSaThoTHhaxG1dqCzobnG5r4iTmcBSwoq3vjarA88JUlOQS6+gfxo0X6sz+YlJEG
ty7++FIUXUYKT7BtabNU17ArPZbFyLmZ+KfORCTHEgcPL/jYHumtslafppRQCF1wmf4+W40lcV6D
HkHSPUp5O927UgfesXPbj0/1z3hj8FzVm/Gfr5ruX7oBWWPdzIM5LWXPEx1hywEJDw3dS7x40j6K
f4Nm4jNTSYzDWOM5sfEo/SWbfo/0C+9gbpWAvkbKf4usYPS3v0PFHiUuk9hKA43yc8pXHs+mQvQy
DY03HAsM/TSjN2Pu8BSQDcYQ1YpJKCyIULZujU02aLgu5zs9Dxhoa48gRXgHYU9sL72ZveSOkYzY
78Ah85/n3cAUSXdu6hKEcDhdoran2AMfDmEek0graAxdsFn/4a0rMk7ESXEvfp2IPuVqDYWDi0rX
Z9xpRuR6cqh2tm4aeo9Xbdca2I8bWcg3W5nTZ/MAF8y2/7e4qk+r3q8/2HoOAtPwcU9dRUPJcDCB
g98fjIbLls7TM7YaQJIr2OtZTmKFqjoQQgUT1RPHfGFrIOlSLhcy3W1yN9I1dX7+PWOnIZIqtz3S
h4jZGu4nrSY0mmh09UWAkdTXSpGjIgB7v0LHYp7ufhdYCH1V2kFEBnA4XeSInBPCWoq2w95vsHHn
1XaaJqmkS735BJo6owpZYynUNT7b2d8aA79KP+xM5baGIJQBvVPcitHbDxS1IB7WeoKtWA13QMBU
Kt4+cwrk2c1M1rZnN6rjoDch8Sqzz5C+hhN5lkaMXydeB2aDe3JSNF8oZWJUA5L+81ApY09liOP7
tbF4ujdHXdAWQ11rQZTBviKoCvABi0WwkvyYhTXxfA/KITWBEe+p796Hq7xiJddLEhoWnNYvg9v/
QnJDJCJKaY+I+DOYSpJZ0PR/CNiR+w3wocfqgKktBL4gUiXeDhFW5Cy+QamNoaE9ewDJrVmEib2J
AiNB81HizFSbJgLWs9g7ld2r1k6fdWAAae9mopO0hno4xjVs41gU0gA/oxPTsPMUpSlG+HfMha64
RtVoJkdIp1xyS0KLv/1AHOfbyn8rOs43Fpmrv7dC89KUkpi5B3lkgqOI2GF9wPV3nmiBqSW0QHPt
IClFAd8Z5Oi32A7KqKQ6b39f/0fTRAl4pLQE2DCdlbmnRTmImfH5GHGKgbx7KvilVAZGi3gXc24o
h5uO95UAhNKVrbyKmrVSWAcs83SH9lFJ+lRfCQwujcq1DFhsCMyORhWUSnzGBZoDshZOWe/fDEZl
pNZcYiMPRleHZGh13jOXyjI3epwfk0FxVa7MmouD8A6arRwwYw3Ae8UhSNqSJgG2NoaMT91FvPt8
SftwuTgST1dVaPDMqHQIjXmYVniQWGwdSZ7kmvYfHINU66YPKRgYsWpGWuLGtAgr1aWtsXYbp09z
KF/k7v8AEy8Z4gqMUNEoGPau+MrjhCpipy2XZ72bZBORwtBVPlEiog3Xk1hjMCsxZ2o4cAcQX/UL
I2BhaFAYYPRKb5//on6uVMeDUb/M3nZwynMIuItJTvDfm3rrcNwprkqArnz5pawv1nVqGH3wy3GC
8KCUtibEt4hPfK7n69OMFNJUKUEU4cLfs54SBEZcsvp7jp4/FOStVUiSsfP2mdVgIqnu1zsPZ1FT
cH+JA+jeUw+xBkzmbATCg+2k8+FFNZ56gVIAIUo1X5QBvXGhLG4N6rBRc92fvLtHpTMJANbbB5qV
58rIO41ubZ1wvR62cqzWi99llEPLx1hXnY8dlWWk/6atK+KZ8ySmJo6dU2xqEWZbAYTBXlITdmw4
3cmlSYZ2YHSGl9kngF1xvSK4o0+Wy1gtefuv49c8xIHSjk44z0EkFuVimluOZ2np5nMjOZA4fOpj
IngrMhS46abNx+TEF0l+QfS+d27agSBhnIzuB/jzj27+jHmk/comqoHooqCLMP6Nzs3sQ4L1BDHH
2G4H3T90cXu3/TchG40+UVJ7aH2QL8HCvHuZRbnjpb16RGiDplMLizo5juasQYSF9MZylDaym6nD
7TisFiYVs2j9eyTxHnhBe56W08eKnTg17MimnsNOjPuQCGI2EdMON8y9/zFqpTG5NTnlB3fbOMnv
Iv5gCgGS+NdBZ+kDgSEhEbRNFz9MZwPtBRwGNlPXJ3Srb9ANxF0MJAFu5MAESR78ym/AtcVIydKU
KXMPzDFRMGZ0ZYkbqzuhY417TUNtF8y41hGkqD+t0vMHc01HZN0G4qID8gJfp9YQRBuQW9brHks0
m/H/AxuJuW9ZncCXkSvWJZo8wgtjbRbpJsSNm21H5dqbr7nj/gnep+hiTCz5BTd9aCkWPYspKHD9
nBH+EGhTv5I4qLu8/+EmPi7zRvMI9LIp2lZnbgX906NiO4CgjZR+XQX0077epYZZTgukiYoo5Drh
dZx3pGX2DJhrAhn9T1PKOkLQg7/IrgeE1akb8qu4JcqZOwr1hKg3CyeiboRuH0F6HoDX7ZPQrgHn
mL0zCrGeGuGy92PwD2iTftA5+h4qJtTX+MGc89gLKaIFAx1++qLtM0LKqWv1Om6sQIUr92gSM9Om
1yQWmubY3JUpP+KE8X1BVAPFoAlUuR8DdNwyAURHqwhGJjXKdNA03GHSaVTfZnJ/SQdOCpqeIaZk
JuBxAl9WGnUTCliCEjY8M42JBQqsd+kcom73PHTYcKvKGxvSDR9/MfqelDNkXqF4jjSAODWATNP2
97E8p9829erso+TVcSh5/IsnTKFpag3Vu55bw94jXm6D2fDrVxIVITDXMti6h7Sogy+9wbSJZ/MA
bYH2XmYhmBlC0yMLTiEL329Zu+Kmy+z7b2LET76lb/F3l8Ur2j2bWydCszVGpEW4qdJFYPbffG+n
3eFgrDiQYGIbigybqpb0qGIc9Fz/bTiKLsF56UwHWjDYyozKbQUMa4HBlBjSODZnpD287HtNjJiG
U0T1+osF955nWrEumTWsiiz9n8AJHsXXFOVtJRDAFzIMi9Us+WzFenn4is9mFe0Gt+XN3gtmBhss
cZVsOfI9d4Hyb8r9Vy41CcSrP/6z397q/cUbSGaDOtZQV1IyagGnYUdXWeTG63suel34eOJ02LoM
2hcsY9AaY7zV+TgsxtVRZwyMZejdDiHPYrloBA/yx6VKiLok74GBwPkduhAOPIvyyvw/6D4yuRx2
4RcjdN0iTQZ8jTCVUDC7ycni7hvhLFHOJBwFJMVZArcyxPrIDyxJnanUq0P5n+IwsnD4myiT2N6Q
dFboLVyBJ1LSpGwn3BLhxAyY3IlJT9UH/7crqEOGVobtHvOM5W3TvcM+6CPhVp2FfjinUkBJHQg9
L/b5lwyOqxkO8kaPmu9DzfKpI787m9CB7+Ia7gO4jvQFSMDU+jIAZ7GfiH6/I5cmOYg+JYq6qT6n
52IrU4NiLEdBVM/DGjELbaFRDBZL7ejMVuLx+o+Nv8BXnAlM6AhbGp1wuOFB1SnbhrcAmDS5DgOX
1lzwxdAEUvKGkR5GNVZxHlRfm0E8OzTcC6ffZShnEjICHcpxgyqLeW9gDIYP5xBQuwjVcVKhQGPK
USsyeoUr0eH/TVDmsvy+J0ze3wLQlQNcucKcWReR2aHhnKjGUhg2ZheyT4Jm5XKxD12V3IYxUQdF
JhNzYvCrKld9usM9g3yXcVBVDjLNU387qrTQ4Gq6mhzMhY2uZ7nsx/Ee0V1fd3FUjrxnwDaRNToO
aEOKDIIt24fDypbQ1GxDYkBsdyhhXfkvElv0UrAj+9d25MH+Ji2e8enpWpdy+T93DZ5bN7zTRJ/T
syUSMb/ohI7CJK/hApHU+c6z+tShO7qsCEdEi0UiMDSR9oIKKZddq/yozYuT4h9qRTJAYweCQjq+
cJ+aHSex4S/d2CNMZzwIencOtMQW3H3uBBr8TyJx9/lF9+y2+Zv4ct4KzBjUothL55jlH2p5zmXK
EyhL6ejyx4c73Z6f//ZODow7nlIBNYhPBDWm9h+2vdowQ7SwknplEwTtVc5J6xVxSKq/+MV9qjBl
Mnkgsl0XhMjpaOqTV9+yA1RrCEh32nx56Xz6/44h3W+FyZWVctbmLJbqCL61hxffR3TLCD+FIgfx
nzQMGXOtL4CS8/zf88IasgsGwfmNzTytHPX5Un0s9aQDHommKk2OT+oTqnJLmXpP8WNqkISTFGq1
sr0Ag0AXEqf+AMPkpXoB/ymDWLBcReCes2jA4EbNixMdcEnG8YRCFgmRGoherzkNolNh3/1rRx6n
ZUVoiNVIlKO1ZUGd2KgFGKl0EDhz/jUdZ6SQG7Kj6I3n+QTU4pLGhjH6EEES4mP/Ny6Tji9RaOqu
6f8SrTwsFOoxnGJokNiABw33B9yh9XCxRxd+OYIoqu/kJ/0v/K+YKpJjrtEAbqsIqBn3O/JEW5FO
gtiJwf1yEye5lCBGR+yQ5X2ZGqBTpxboHavY/z/6to1s5CYoiX9XZCoueAOPpDwnI6JDtPoDNKJ2
rtnF0nXmt5gi9l9vv5FjEAatm6HA9q5chQn84VscXN9Lkp9lpk5vfBmkJw/AW+NomNWQUB1U3NM8
SIxH+eW6bgAPYkUQT/x2vN5wgw523LPlrNEAEbVp6v2FX1V8aFo+u89bS8KAGywKLyzMWIa5N605
Mvm3OG+8d4WZW+eMk26aAAGKUHEWsnK+otgvI7FVoPFcvu0JaMJuIA4xjTlXyNuA97n8gcdThHlb
yhOnSKREUJzN3PK0xlpOEAO1flvXJVDo0RH1AjOubRT7V2cH9eiV+mhBS4WY5AEhtPOXfZTxPXZ8
tYkHVnG1QdoAUjLdrnQtCteonokO931+mvJRa6Ui8XYqe9M08b7KAhC7P677SeYcvyO/06NhTB0A
tZbK6zUOgAz8IOYRJ/q5WZDgb/EZGhvOugSzbgd9q5TQxsAXC/ZPdBbkucfaiCEqfJ2UVzOMhDkN
wNeN+eVUlXRZyOJuytA1za9JwoQChghXUqv3NnLn2P1W7sKcbMJlSKWQiB+wJmRbD4z9KctuEcdr
+rh1JUwZcICEsWFk4ChOfIyoUII20vparPs5A3R/QPhi03oEHkSLWkgL+v8QakFrom7kxbKMcW8n
sFzctA8L89b3Ahk50pi6lbEHk5OfkdwXc1gzmy6AU8Nd8YIrHsM4gkXl3daJpOePC9qaepzOpFmm
T6zOcjpqD4/C1ghFFnEXk4RxaAsqi1MeTKuKNrWk8Xi7m/8658ZzNTW6987UuZZBed9QxhJQr4PL
TpHwy6rkRJr0WflXPW8oWEdWlXsGt3rfSBPSUI084Fhuvxeen/lSIGxmxYIfeK6zXODRjOhqDMDV
+l1ULixuCPGeGo6P6OPjsqKkGiCNxKNKkTWd7/nY3BcfGu8BA3hQUGmOUhdh0Uh2xBXEzO+DjB9o
GJuRfNVcHPJPnnuREMpajIJZ5B4sYd/y6J2eqDAd9ReJMUK6XoKQB3+FbFG/2aCFN5gWi5Rm5ZdN
gPlP3Wbae817d0CCTROqUYEep2AUIdLDSxmrjOBCCUdXEMbA25PYHc+FMdXc2QeovrmlDkuEZ9eT
6LzbfPzZeP34sHWP325Hge4sjdu6FvrPmQmslGMW2aFH1UCoHpLU6Gdq7WTU4sG7EvKEe7TaIRqO
kBPxw/Ssb9hHImRE/cNa2IgkKjVukdgQuztkTXOsdQrrJeg+wQFfa/6C5f+aOvrv5JY7Ns5Tv06p
0lCLkURf78qbc74gHCYvhPzTNYSTfh8ypOmxFSRyu9/WWQuRzTVX8qUPUPU/dhmPoh0UWHCBNuY2
5kGS4Evhb/Rs6f5IjexTUKj14asqwMKBe9GI/CCF1ME2g38UV6boQWWdazgiBUfMKuAdG9xdGUDp
jFSkFYjZ3GUN7jr99H43yhe6JFEMprXU9qq+tqbW01SiU0TM7PkCGeK99JE+hc3/JqLlOr0lmYsn
zPuifwGdB2a9b+InRUwJnmDHXnwOyBLkp4oUQt6gYx1XKxYB332vluPXe3gBGC+ujjbyzlSxWAFX
qrLHS1QUkL2CyTHWru+Kyi7od7tcjdk8fCy714cq97UvXpN1d6z4DNMs7yhwgx/ZX0Isi3OJu4HX
sgrL346lhUrlVAbLVU3gPw1btTvYHMK7wyU/OXgmpLg3yikmnJA+/Jl6B0enjnQ3jTmkzgNswHP/
WgRidpgo9+vQNHwXBKAv9EXuOFq0r/+H9tia/0YPwrTZ+HwCeDmUT03d/RRR1iR9mJKwu2Rzky/G
TTIy8jYb5PNg2fkx/ulQj29m+RDj52fQa7ELFKdl+IU36kJD7aitk1kO4YDN2E3l1Mjv/Kf36xLP
Ul2yw/4yUdq39L7pomimgjPsW+ZJoK81crTXq2JYQFjye/mwVIZLFQuITKXi92z5JJrWqQbKfR7x
qWbe5dBgS2uLI1+Q2Jl+tRWsO07NRYjqQvRmU3UBK7zI+YPhT/uTZ42lK/tcck+TcV5A9eP54wQy
f4UaqoNLrdT3u7mY2/00V6CAKYxlZgU2VJOA4sCP5eTkszbN+KDTlq+2teQIExEnIdd0XDDWcelR
4H2M7/OyB7d9bQQe5tpsjvlpXEJZRGlh/cPloK5CciakVKR6NWrZFUSDMceJG/e53EytYYjVtAao
3aSj7xEOyPkiv2Q3E1OUYEoyC2l/ICrAiwicPwf8zIQXpzgIF3ZNYlD4YGI1mexumugVuDjH4luU
OM1pcgW51nYbZHdZTr8skE9L49NF6qPdDYoThv7nlJRF1uKuXUytkKc/cgYzRX3Nco7jeJmzRI4n
V92G4Y7OHI9lwxCzdGYomVbV7ZHGM6JguXN/IODRh6v93JTj1CXC/uD/4Mg8w1K2KLz4DZ3nAysz
xV1ZlZDgTvhN0mY/51bbWFVXqpOwvdP1GcJiPQrMTAjPbHt1dvQSS6/ROf1mIZTM0RSHRr+jDv+T
CDCMbpyr7JCp3NwD0IC6sWHGosZvDcaU+mMFsW9J/455XFaEJknssFyAsFmbdVpH5xkbDZ+cBbSZ
my3QkLCFLTUsxKsIYjoEotFC0JngPWzWhRTOwNOkHzQZmybZ9iH+w1jtOwQn79C+KFpt01QCTpSj
YhrCyjCFj9MdxgFy4PysYjSSG3PKcRFwipX3JGdoYC9OCzYTy0icTfcqnZSViF1Wl8A/pqB7Qgyb
UmzNeg3A+RXgOl6U3ccZlpObuslj910EOqOPMbWtJkhoVL2aXfXYD9Zs/A/uM3uV0PuFMAMxgdZQ
7jvrCF9D3gdWeVU0iKj/+imq0savaOIwjrRSjJQmtmpJJQ/vOIun2thD6QvY23/eyAChjTAZ/nJd
KbhxA2rC1ATgl7TSy101QeRWevMGDIKztZe46wm7OpvoN0RMvA/QNwMwNWjh45Cnu0X1etDJRykt
6T4S5bB8ftc29qCLuxpV8e44PLTa495maVbaxABqQY/7/tF9QecQ60YnmJaOiYYO4cQDyMfcVXQX
i/8f8HlYhX8ZSbEWUNlht+FRPYlj2t1BagBHu+gcqORili8XPyclk6jJBZ3znkzU+dTBcwoDNef6
XXhuxeiXMREA7vOWjdm2EiUfZaz1Yyi71HaD39RSy7e9kzCnFs2suNhdiN9GCzfU6bZA/3XhuKrf
Rwq+juBV8xzdgMhWoTRTWub4cqVyP6SvaQHGdZFdgMiXoj6BLyDr0woASZCzCwYSWd3OgTrls/1i
XBL+WY9vQ9aMkDxTnu9rDjSLwnMk3WiNjPLQJHKbfrkZvfm1X3J6kyDbGaiEdm/wFyl5TnO5e1y0
AJM7oR5u+JZuRSTo8c6a2zu1mSOPQtDlFOWusNPZKkMedIV2mHWWHZnudlvJ1W2ToS7Bxis0oplH
vil/eIEdM7jaygoVKJ1HJQnm/MmIrFZ5KNqunMp8JtOvSExC4VQ7Wrh47EKq0FNLP2Ww43IS0Yfp
b55pJvaVXGoaLBzytVZICouv+IeY5/aizksKlwDQpG0Q8KEgECUKOWqKKsSiuQELScjSmY53vAhs
OLnfm+dsbMV+1L65tPjcVXv9ZCrPNmmw4Uwnu0jJ8L54JLGXD+YHwjXLLay5GWvN5UKzEX1s2VPg
qwr4g4gA2LjiqiTSikZjDkowB07cRYJbqhMTUlnRD/LpMCFUvM2Qvk70Lwc1YsrZ+zizbbn5QAa9
03FCSLzTviTjzfdT0TXMBgPntxQL4SrridwbG4s0tCXel7bxvnpz5qwxgCDaujY8M+kcwg1YBg8Q
LUcV00PqKMJXSXlJR2nPpICu/ZCb95ToCgu4xqe0SW6f9bcTDeLluyovUw8VcKTEotY7/gabrPJ2
tQyMeL9Hk40wCqqJSV6Cxkdrp7BePKsW1GtJxYuZgiN+lg7oyMyVhAMIaU+QDDuwMQMjGgZCKS33
X0eYnpVQwPT8XioangbhM0M45AX7U1TMP7qB0+EQzJSbSOxXo7cJWMCZyVE5r0vIhsPjZc6V8gIj
uC0YlFj1xVEJ8P8pSrL1r3haZYCErxBp3lUM7z7IxPQTHMZCY+vnhGXV5oJF8Ru3KV7f2KfZwpj5
gtKKKs47GpyneqSaGov8nXfNg51wxPnxMFimiTS92h9hG7r7Qip9Zcs403YczNw7QS9U+j6g/MBJ
SvKTAKEWuUsFjv452Es60IchpTCXWVYMN7SaMqju2uxiA1bPM5vVXf2VyI40Jr3EPVAGB5jLaE3l
Qt5hg1Djf0rR2+5GcsbJ3JGrYSKC+QLlIVsrqKDTUkVt+UqKdFdu7eHXc645Sb1FNHtpmgnildIG
mJPT+b+K7YIVJZz4US9faJpXXN7nRz8OLMj8YTecxP2Du+BxHuys8P5kjG5aUyMeGqfdpaKRjuov
/LhrMbvsCePASctfbG98HOX5ijcIUXVD1/mdGd+meGJceiPjkyBcz5xSMf9sczN9lnq+NAQl2QxT
qM8MtzdL59SUpqt5MeZnOdyAE++orkvNGtecTvo8Lo8OOt/+M8RS4USAI5NYEFr3eNUIUeeiDIGO
qpOAYIcsJIXBkDG6l83vhjfCLYhew+1+Aipkmr4HPXdyFW363BnNzototZXlIjnN1NnmkLjNpWWY
WOqYiX5NskUf8w1cCq5mIWMZaBfqXa2lZjJik5v3Vca7KaX+JXAa9jbZMP7bo1U8XAQHuKAP1b9p
PZl7qqfjPZlX5/d+nHGZg7mZHMQEp0z/gWoHpxzz3p3WsGypVMaNv3Q6sfyUqot7aKIrApcwT4fR
E4FcfTeiSQO221khQjbuleHaiinDZQzJZZex5L8kaAkIOuCP9mZ6M9RrjHjEqljfmB4fZt5KoxkX
QUHJW6v+IYiqy5FQ0WguhiF7z2qdhHPuevEWLpURPUl2srBmDOr/f3+L+CGjmfrT5PE5ivHJNZlE
egbnMK2ohFSLtpRHrsaeytDoXRV3BQxBI3qNCLquyXa7Pe65gn4Hgtxo+njUK6oq4Xio5YoDWQTc
KSvlxBkSubrN3YSBZjAu7d2qflgdUipJgnb0zJ3117CjxjBdN6rCu/fNKjvNk3rqwwlsJKVr8zcw
25EyaNvOcQ2CZaGSyGa7YV7R9LeRg6+rWmvkL6+zvSVOOxUpLdIWii/1fEQdG7UPW91KbRTLhJ+K
RaxtZsbNRM0FU6xKTP+REEN2AHh/yCkX1iiLs4JWE7FsA16PcQjYvQuplvCOkpMwDMiSIOpznAYl
GJ+GxBrNReotxudzj2plK+t05pCb0EDnltwK9APnUMN7Pew6XC/ZmG67OJyUMFf06wbtxP6jSf/P
yks92mplGQXgHc/TSSWoAdqy+B3CEPODAgvmbOa5/peYTNl36AljDvMKzPjUoyMrPnUR35lPWdf8
cCewt9nDTwSGftAfj7FSUhW7BbQgoD92KGuNppBxQFsWbd7xQlePj/umCBLD/h4h771F5pfDQRXM
B7qI1p6J1dox00To/70K7mG9/wEWMtjkS2piI8LqZ/eKgQPxfgxFmr1SrK6LNnj0SXHNex8TQ7wF
/PyBwWL8ejf3SbDfCa9DiZEUklNltl/uP7jiwy2J/x8nlpSfrGr5cYdJfNsoN2GiHMc04N3tc2jm
t9eHFeqXSO4g5u7DgASrr8nScSz2TMDzBOdZ1JcO53JhGV6LfNuPQylf+dWEMbZV6st1DRRCU6/N
BDur2F/KehetvLuAeiVDS0YZNU7Mj1cTVykbfzu16q4SuDXtvdg/9gARn9U68NP54cswY2mH+oiM
cV9lgkWQPUn1YB3sm4moSZDFWl45pd8mFPa11fpy+zCvV/CTflSCpte0cqc5um6r9zCGQ4VWHHdy
UQtZgX6s90wLEqGDVgajyvxVDOICm3b+VxHwHdPBRtSp+eBo95NywTSuFHU7yif3dQXSSzkWWPFl
jDDwICIwGJKI60elRao/r9I6yA47ww7PJMcMUvPS/n6cfr63CBn7g2BIijG5i4GlM+qpaHsor+8x
94VzLbH8AD7Zk+SwI5d3NTPHBEas6sEgnoZ8LzjT8/dJG+YQ203jJ6CsQL5Cer7SKIMQHG7ClQOY
HBGYOeTzBwndK7XYXanqLxsG8jD75PdW74Uj6JxT3zY0KTfjDHceFIBsG1kl29jCg4bfGyLEwaZZ
cMr+nB3c18X6iwHQXLLIJ07ZD7TFOo9ae6+UYlBpfM6Ubj6LcaXANjYXlzddl3+CAw3yqmh8ZVjS
WyxXhj1AKF8SKLWFVNaX7xd6QRIz7VARkr2wdU7+9LOrvcgf2eHHtaydMOUswJVMBza7pplftTZC
AmC/VeuJ0Jlpi0A5+gHm7L7XLQgRsrO3idJCYibnh5IAsGgGvntVjFfOcnZoBbXcX6BMnDMoNTK+
LnlP3Drc4B467+rQMH0D2ez2o0dbGjXfd6wVB8uE221wDUQU8bf5wHdZ5VY/tiwAh1wVwRKqHEAU
d/WI1/e4JzPi9XVw/TJGU+93WYmt71v3yAA5Kj/iEDzbx1Tnm1Gw6YYKvDpYuZj4UmTgYDtWHxiX
zM3YXWgRm9/SpnaZUMFw+WLEI3i/dT6bSSGvdBRiFvPt/7hojci5jIuvAaA+0aiBvy5x8p7KKjdS
lEkF/l7WhW1qaPw3C8A/Y52fKQiotqCjs+jAW2z0ry2BpsJdGr8RlpsSZAwdxNmzHzfF61tl9yMK
vWL0WLTJVHDLCTCbs97WCqIEwsuZhblgdJIce/rzLy9IvuY+x0mCedaQjEA9r0izNOb1MQ5aNkJ1
vQivMr9vhfGOig5zzL8olezUrHvEl89Qbr2D6jVsdIJ67ilGB6Iipmmg73uUEkpRptxaKDeK4KM2
OKy50tze6Blkx7ZbGiGs7AkApWyFcLn1Ps43OBvUQNbChCz/qUEmH11P+id52VYMYmeOvlGvdIc/
Tqf+9aif0h5U84CpvbD2o8KQCnI3izJKvx9A9w+7zs134MaD1hvDeHDAJTid8vctN7OrX68UhjJL
L0c/rRHWyv89XFANLzqWZ4CDX2UHVggw6WfoNkUaqAjsKelo+amGNFZi8gHEfnB3zZcrnS97FK0c
v8K8s+x1dfChr3T0Xo/p/q5gE4Oh53B5RXAo+T61jBTeburngNXzO4oAE1wwueX3WRLE0zuK9nhW
hHL4qRgcjNb0IaapjiNzyer9WJrMU7m81131yhjs9gVgjkjgNZvOA5sAVvjQdAFvk57+6s6pj9cI
ghN/XSBGSNxxTiVPm6pj+Twlwqrzo1G1svAiEQjZfxPpYXZ9sxX/sh67vhqJ7/c7rQhjD0rLevTs
robjz5zwMPK2n7RrUzeOK1XfbDKBOhr3+tkdgSD0d/bLTf82/myFVOSJCz9qIKZIMg3kHtp7idKa
CXzAvnlYWnK4asSHV6nglqlCUQsrleC8xH4e4GpKrp/v/RqJffX9NZirb7itk5nJk2td83TKebuT
AVpGHuv8Mq0MOO3QZo8Z/wsra4A1XY38peG1XPUt8a+kUZa266lMYaorpjUsXCQaCQ9e9QpP6lMS
uZ04nhGb6NhXNexqhVuk5NQoyS+OdYuPYdN8hBOG8EPdnmYTOyJiTKmobMZYDEWRE2JGN/d14tCw
no1CyVkDfLeDpYj6uJcuebBAJxY7zi6WoXtUcZKw9XFosCZRoBkiAZh0H3NmEmvPbSfEr/Kjkgqc
uNNtGvCwNJnYsa2rFftaro5UEqx5LE+rixvoX3e5rUWdkx61XCG1mWAroDl43bcdENzFtD/Y4ZZu
xdJutkpgtTh0TsquN/Pqk9nvO4GYNDgijjBO6SQJ27Z8PEnOzNlfvkS4q+qy+b0e/hglI1e5RQC7
HibBP0Qsr2tyi2cRKRvPQu/epiZUkUW7jaGBnvULHDKeTfejsdQF7S+PnHphYe6dxO/85ASIN+FB
MHt3S8jPOpHsMHbZnmKV4RJim2Q1E3tQjXLCF4K28d7g3PyV81uqhkIpnWkaJb+vRoFZDdWgIOt/
q7XhSPRwNkgWbzHhcmGx9aWGsiOLmdysqynTfub/q2EeWDQvIap7wj4fC29uPXvuv1lIuhw4bh5t
aHuVPY8hkUE0iGLVENBx/8znxETDISzXJGLZxlDG/ZuMtQ0DdSprLS//m9+sMhu35VKKqx5Q1/bt
wdyjy4bc1+wM40StCby4Vi55GvVjQzi0SyDAM0e3SLHi3o2XTjwHO8QnrAZd+7VpzxmR7Kg1HOmO
zfgSTBXCx2HVLYwznTFZOmkzTBuHXXet84mytFHACljwRZPlMkRTYbwZ5z0wNzE6MUX7SU5JBCwn
tIN2HfqMXFTgPiYIkDd9NGUVixYxLjChNokTiU4VQrgxOqtUUi16HsJ5QRTczhUC6Z4HOpIAd4T+
hei66UYTF4ieAve897UN4dxMUdGRSq3jVPv1mJxO/2+9YpaBfTYvy4Oz5NNyQKQRK9HbsiKHHEvY
ezFhHhLxtedK4ghxataQfLjRP1IY49xoPgzzOo5561B1zSokNiUeJ2TWan0aAJIzCymzxM3F2V+g
0LB1FnIBijIikm2AZaFqv7DOGI4GPSeHOPM42zexKJjP/srilEp2SDaRp1GN3TIV2qIxKyqx2rfq
yUdVrJ4vKyrDycXvLdZX+ZSkvpJQMldUmvplu1QqnO/mtrOcpvbtE8MZyATOOyEAoaAQdEFWZfqy
hMi6tK4uQoSjrDHkD7eOasWgkqvoziLJI/Rndx0aqxZGD2eOF9rLmUIVWfKts4jN2akm7w7etB1L
BYvXUp0f0CMo5uQNRrWqmYZUy56oMQfnQXmh6jAOwLAYAwfQ57oiR5TvnjUE+KZxfBNekX5koJSn
EchiagD/hm1fdiRQJsnqM9lXfvPYW0hRAuDqqgKWn/FdTa66mgXdxydqHRGlqeKN+rMWMX7v8+7G
WmbhNyOCorwNQgczQefRMbgXlynF2xLpAH+TqEWLE3waZ2DkrnuKWrGYHjQ4k/dGNfhIbKNKFHN0
AULlBmOS78JH4UM6UAfS6mj6g1V0KKgSPp6K+r1v5ue5WFy8s8QoYfPDtD9vMmXIc5N6mbGFeMfe
fRL4Rd9s1UTCSIVbCbhp+w8wAR3JU16yWR9KFC43DybUyXdtykHWWv6VFux42zk9DK28Z3a7ER+b
+XPpW70PJJRK91+PGhYXyuBl53T/fiwmE9plH9zhBKVJmpk7yXs9RAHD+QVu7OddhK46nEuTLF3z
kYsmHv1q+n3U3vgjp+HWeGwbUmkx9QapOIefTKTyNDzLHxRiSgLnJyruk38Jyaw0LYiUjyqZ9/UX
0Psfkmn+G3oNX/l/fH5W9L/uHp0LeGAXLHV6g0aYjdGAU+jBDSgyD9Lhh7sUVj/rzdrTmXWG/cso
fVWwR0SHiP7DqhfTZ5UbUM2Rg1PsszSHk8RRUjQtXeer4QkFDYrO8KyIjv/wwVbzvwv7J9XlkrkB
nSIwkF3JYtoxXK0RbbdUcmLVaVP189vOoB3PI8oC8pPdFaSNrmQYRpaDiZfvbg0NVScPsXvAsBKq
Spd3eX4MxU/YFUCFU1BP7Xiyf+deCBKpr4DfvX0d1ALBRQn1LxUWicJNN9plRzOkaQDDWnPxooFS
2pTCnwGZd3qeroRgDhcLbGw9wS0fEv3rfW10cHH/LZ73XpmBrRmKUFmeiIVWuonyhGWvtFv0Kudi
fk8T86n61Nih30d6ehmzcx2JJiaNf2a1wCl/I9Qxv+naJ8JzcVwtOfUhDWr+4mmhFRwvlRzYZUK4
+HqmAj0mUtsTRcgwia8fy8OXEfokHbbfF46Ir8DzO+rlGiJnkYM+9uOk6ggFO9QWICgB+NiwtaJN
+xEd4wkUPbEPZzcz8XB7tWeFAwwe6QxWq7l8tte56rmYssYT+1VLq/UD/ZfYKlGDA9d4fCWKNIzD
JgwUR/QhfIUTGWpDjo2b0T9lV0UlmdpIk3xDbEf5iYrX8ScNx/4c4uAUmIBp77VZ3QzFqsjb3Xzk
8A/fDwCNS4mtEqBYWcJcJ7gsyycEWdEOmKa/S2M8ohV+tElUSSwuUfK2+0iDhvf8rsqq9ZysMK/H
P0EVAn5Ly1qcH3nbcKnX7KlYvOPZioTggxJk5KRh0rlNX0dTLy+G5giiFUnCFZ74y7jtHE1EHh79
qIsOq+4K3jbQtmv77K5JEtQJhp0mA6BeVYDLNjsboBoJAQp7aO5VgoTn/0d8Vx31mBE5GdSYzOrp
b9EVpM1rkhnlQRGL9sJAuNrALqZbwvZ7UwURmuA1Gr8/cLiXc8Aj5deUq9cwgSRG+pLupNuv0Gpb
W5J0Yl3KWEZZPILog2YyFtIk6ZfRsOE4uAaE1Ea9WDbMfXve7U4dLeNHYlG0toqrv3cBy6+zvrCZ
bvuUavCYGepsJr6psrj8vYEEoatly3hEEZTS8xnWQRPDTBzPOsHiFg/s57YN76SReQTRKmPLn21F
Yf+qDSd7v8vSyefTXxO62HSa9/IJmZZ2EXeXa6T/fWteDqKVEimnS/TY3kDWbWTYkpyX031gYR7c
WKSzHAwHX6Tc4E1AMUtGNJ9K2XhhlXg9hcPWnrn/xlYyrbuVu/r7iOSsylb4sYbq/8cB33KuSVit
Ed6o2wxXXvdvuxVP3HJjzAoAyHCX5NYemC/xnqGda9SgJjtAil7279VgAmJNSS0BiC1szYMi3oOp
hcTqSbn9g0xQiuupO2PuifIu1Bw6Vl9nWtsCBLFdk16pW5OP9OxvJ5rbw1W4+0TALCo2UYA0WBRT
K9mwRT9dqOx11ZuKLH2pBjDYo6OJPIS4q4QV79Xo1OHEZEeqcXnuottkzpPsmT104s8XZiLKl7SO
sH71slWi6Qch9WooyxfCxD2D/iF9Op9PPjvFRa9izkHKe8S2NqpUC8iG9/IlJiy8QSfWOxI3+DNZ
hMaXpJFO0nceTrFPh9LMzHTVCsb22Tll9HBNhyj3C0IYHHu8RzvJGYwSKA8N809yc7DJqNLO1VTi
oZGA+uQ96DrH1Z+Gijh383tjJTKG2gdnrRZ4EV/bWRgQpKDZwP8LLtAr4dV2D0eqZulq/JKfiz4Z
ru7JXkaKkuEUjdDLFIHCi20bL5HHCxsaQWpTAIrxvV3qcduPR2USFyLvJPJhX4bJwJEBG6IsGZ/5
ZbnegE/n2X4JdwP5+GdLK35fJrgtELy1TATZqyDUg+JU+WQNNOjg5h7qneZT5DZkVOo59uJodiEf
soWd6D1CUV1svTUSPIgPqCElW6vNGmYff2QHi9F6sdUB4x/hqr0NY+Hddnb8FynAVDW8S8odgIQg
ueeMD/XihtODjnyNugEso2e1VgkE827WO94SLpock8Pg6JqHkekzUezYzXqwOrLIWjOyIUFqEjyg
hWfOt4VyJNY1u94FsSz/CHgNnkDh5FJ5hvJyILP+x8Ym9k8As4OS83Ba8ohGVbcb8tbbqZ/cqb/x
UstvCSq10GJ86fr1zSlyypMYp0J+j+2Qw+kA5JdzIfEX9cbh5BY7YrbCWYCgD5222+n8vijZheEe
1+59RkVqiNrcg6TzBg+ahJj0yArBdfpCYv0jXCQw5CulXxwJzNwR1pGdbFYdfWmZdZ0C7Y+YQucj
ol92zypkvkN4yzIIYHOPntmHdXzvl/SoppyAETbzMmxX5tRWHabCxe2krUd/CjNA7jbV+dJPILmI
UOzmGQuCOC/MnJS4XgWGZU0AKu4OAdnKAeeo3F0256bTOODLwMKKsFJoOS/mqQ4MsrrgTT4VrFBo
C+Jds9a+7U3m7mksmmYVoI/no3perCzCZLQPF+gZoRZnFLgjUH8Ne3uMOuBqwKTjcFgpT8LER5qB
TlXbJsGBwsyh2ipwr19/TYpD5KK6jg+ZF34K56LuX01M3ZdOcIXB+0qKpG9mSG63wGnCLAhshLKN
lIkR3y4RQzGWMSA/vKDUjN7dGg4EFRlq/b2eIptR/UBC6QLChJpgzxb9DoYng9GJQXOC2/MlYozJ
yNchDvdwOhFemYQhb+M+//t2eUCyTzaj2tyDSfvjQayxXPbmYGdAPPI9SjZp8YClaBj74iGEez3K
TPMOJqyltsOZEbijpSY5zQU9eqXKw9XbDfs0EQ9FEe8NY0dCmCIrBuhuZYj5eU+S6nH74NiamlBf
oprfR3VResm6sTCrA+2kKEI7WFVzRh8E3PmwaqNhAx3YAeCIdYJTBJPYVXbMA0s6QSGGtxHF0DrX
FB51d9ukFfzaxLyXyeLAfiHUuPwN+sV2YSwC2qHB/pSLJG//qN5T36hQnYsS+R8YJrTkqEO7RzS3
VjH9GnarnoFDwUe6U3xecjm9B+IjzRfnL9qaPOW2iZlfqKecwLew5SZ4fW0KUVPyrjE90AFuXvOj
X1O5wFc8CnqmFKnzera+5xPjqhOS81HLKl5lKy1qf8cHrZ6g0HMc7Mai2C6k0klICsvfPbBHGJc2
sdzbVtTw2MxFHM7JL682OfUawNbf5JrjKMovorQCO+94aOLbW79XAAd2YDn2N6DatZJT384fzm/e
W3/cGDq9NpuxplI108TCDHl+RRYzkgjciClq/3uJfHwlKqfcdZuyuI+WyKgW8FYUsWLWRQp/NGWp
p2dYPc+t23GdH4z/jOgzyDHYtl2U9oJADvHpXJ4wTLa3F6spmN0AU9AYR148yFgr8GjIVH0HgByC
pKPflZOD483zRSrdiEaEw/DNlikFLCAQHmM8aKGpSpZ24HofctONOX+wxpa+2Jw/oqwNX43fzuOW
p56uxICFLyCCupwKG3gw1Y87BLu5K3XN2L9a0mfZNF+2xxHWvuEuCw2MzBZAKPw+AnMxCksxSVeO
31/e7GsTEo/3mzKvIO+rdipt5t4LsO47rgWdEhLQmbGp1nVicX90HPSdZ7toeySdX3zF/2YzhIVg
eWu6EaJPonwJEtdAsug9P7aCJcfdh9zRPBgirAE0gfIK15SehaJ5eVaskyYuuGdNMT+ZPWsN5ggH
zS4Wwk32JkUd9FYrUNdUui5GSSUV/EqEX/yc6WOtWsf/0gf9VQegOZDiP+clRdPO2HUdlxY3IY+W
nkMbJCfsOtxD3EzCfeJYp2ej3i0BQPrYssHfvN727rdmkuMbw+x5HS30ZWtfUnn+Fodc77S3cTyg
L1jdjWQqGeVCKbl7Z0l5Pcxi3S7oqPkjH/q+Uzk8XPTYfsfkhW2/qBlksrWQxNhiNiAN7RL+ITMJ
P0HyzHT6yhAmoXNdhRuBOmSjlYS2dW8i8QSULI15/FfxA9NuBi1ZFtmxomYHVJkdWQKwg6QI05wl
S5QmbU3+JxSSv1MZMlb5X6fPSgkfjV1JIClf0Xuba1chT6t5JQvswi3NMUUNiUsxTd94Ca2ts0U3
pt9i0gf3X212m7vwTXJHo6txjIzPUF+3Nj3VtnqgpqEiJnAji5DkYBwiu2z8G9jN3Tx3sKIymLY1
8xiLnrinfhCw4c3gbeG1sX0ChQgSV61FiO3torYf4fmGRFGmJFoFS+7Uw11A9DTfadZ7hCcgw4Xu
S7eBXECANoCPJ4hSSLHSgQCMU3zOf3sHjpPZkDXIeDkaU3xzbDMntCBWvx8BXNo8sC06L7uJzq9k
O1s2wSev2LY6sdAIlO9kF68BplqddE67rsoJsYSE3e0SFeF855eu0KIw6NKiwIEStQkCt5DrBkGP
HYQkMQkvJons+/UrSYYTBzFTKHvcsQ1CQ3XlNkw0ZZwdkgiEQkrx0MeSJfr9A14DEBG93lDIaEps
3DtEzInIN8+/Yrg3IiW61xzsnWxaBrHiA0m+Ke0p7LCw1DUyLAc+ydohYb849nnxEBklufmrXuUr
Y3aEXkoePCxCL1g4tnn/LJKBKLxxwMtj1JF5dpAkRXKMKnCY96NiLXBPkXtKkLigq6aPK542tVq2
kmJTYvUBrswZMDNItb0WCUvVBYax2qwmVpSYBLJtUWe0ShFOSxjtFTDCRHUPEOoZwT7IpLh2pAVm
zdyxvHbXgkyvBicRuCIppDPpG8IrwYd8Kncy2M8f3pZfjvjQWom1kTJAgi83ikJerNkiqQxQENAx
Aa5mesLv92IDG6426c24sHU09WJ7Am87AomI7ujF4R8ycwr9K5Z1fR6usPgHAbJ+dhUQRZZrkZrs
p3N4DUlkSlP6afObEC58Eg/YATdC2pzTKTNNl+h7QawpDLnv0FjLCFNckXxSMYPUCkqFSHr+MonX
HRDPQRhQyKJSk+7Zsv16pKG5Npav66GQB8dFMnJqo1vfWsaiIdDiAHUaKGeFtyZJMWalnFtOsBk8
DkRmIFzVylROLpqzrgDqI0DVJyUp4ZOQ3wUZ0yS/f6/KxdQJYDVrgcGzicdIFxFEoQwkq6WN2WeY
X0uYUO9akUD+m1W5n+RZuX1IJMDA9vFY2njkTHENNc3g9/g/buWKM3L0jkXM5vQo9Y6azBH+EqA9
a9GAszBo9F+GNNMAnaMB2mG7bQ3DhUl0SxlQnse5Lyb2ZWDsXmf/p8GOwCp57e5VbeNUwybRx2Sd
nCKxlBMI57zUFRJvUChRhcE+OZ/1rJD6ghWhQLIIS3BNyEbi4RKqiWy1t5z5Nc+jkBXgzPb82doB
p3zm+KOv7BeUwWihD0XV2X5+bNsisx/O3ZmWr16y2WA0j4jsgq2TSPLEeMSWYdScUuHpc6vFFTKU
ehMRtZ4Fby1i5n4flkaEdO3t6ynbkTViJCTf9P1cxM8xOSx7s2LprQ+Y76oIeARojp5G7wYLb/xL
T3Eez+u9/IWMr5fzCxTYlp6QULeS/1Z0qU2BlnV7PvH7/xR19r40wTrLmH5g5XA/K+bqFBVtDwJ1
94EKU5+NW9VdQXBbbrCPrwlYNMJCs8DInzBK4TVS7dj5bpp3fdgM6weNzHIjaj4FiJCmUDrUIhfG
ky/+45jPuW1Rx8xRXRCadzSIVZR/8+iI46v5T9htE2I3PVMSK6E6jjZWGsbrlqN4zatQh6K5z6vM
D74oyiccePjyqz6BIov8VA9xLdG0I/2ozKy2jJPOGx63PUL/Jf94sd96280+mBPQjH1he9wV0m/p
FUMiqZ488fWMX4D8fNRYzkjY4MJMaU98yCOiNWPOIF90eMl8G/mjK+FUKaMSOW7sB4qxBNBLTlH+
oXnJ2CF4wbD+L3HSOduoQ5rX55QttK/z7dT1kQMkIVZohwPG/gdHLbvSHdfme7CctYjOr9KWc06X
4yTJ6DpKKMDu2KK6CvMUquok9RrWX/punp1s3ea03EtLq82Lr7q0fsAiq4FimAm9nyAoCTTnHfTB
RRGbV6QIRU3Pp3y+bbuOy1k6P/HTQN7DJKaD4+K2XgY4yZJJ9Uv9EqL2OYQdla5Sy0ibRyFEAWEV
9wKmUF1VDdWhgQ8cL3dOjNvlQc2XG9J27C/fFhXzJV7jknNp91k83FiCQ2/VhrTLNo7SUPMpIxnb
DL3kYYubmh2yE4TaC+I9cPVmswHamWE2Ofg/SMgDHJJkZGZ6GgmwjWneCz+aAn2ZxnIiIz8XtjWS
/4p/Fa1T+L9z3t1p4zofIWh/zRJXrBvX7YypzcROCt2W5X3ghHPJgNcRBEBubALa1XnbGsAlaN4n
b5lSq2fBqWz88PD2wrJfC1l5R5Me10bXID6YAK9FmsKHZluxYPMNKMtBRdbTf//34u50tZHQw+ZB
EYeZ0j73RbEij2jcg9S4h8vi2nXVSbKSBXeimS42d9Vi3u2NhcAlRu23Nqh+YNI0OPvI7s59SndD
yBeIObuX3ZmfgQA7q5LnFpV5uW7/mmQ7hSw6ko3JhhEBhFbmIl4wIE/5o/elwpfhAwnRnVoGs3a5
1U5Gc92RShske4vLK1ZeOXCMgbeSW1mPppr/VD/G9v0lLr9C7eCJ0ZNL+ohMCVPlISMDf+YC/V+u
a9goHKy9xRZzx5FJlAC3s+yxSn330c6yOxF2BsDH7Btyl9RwoqU+2nmn79hcSdUFSuDfobAk0mfn
edJ5iMvTBqAIfKRnz+6b5jcTk7n9wI9aL+alSLGvEAEKPqvPzsmscYSBofdyC8xPjiQv/VBmrWOI
uSjEqw6VvRLmN9hR3VEO0K7ps7WdsI/tdmokDJA18VCOkZG4cWAZk0xWPuAtpnsrQ1D4XgpLgkTp
XZ1y4E+cAu2j2/RUXWyQKYJ82gGo3FV8HrVh1LjhNErlli1cOrEgQlUd6WzCgLU8Zye5kMR2NHE/
OvMJmWAAay83YjfCt8DL+l7af3HozgW87VwvdApdYVmoONT8pNQIrxy4xKAX4+/6W2rmE8/fxS4w
LzaWXk/YcyGA/w1rSbIbqDFR2c6+eQIPQd4Rok0lCS7FKnLDKT/aEig47wN4eLc+D6UOHr0qgELt
hFPJh5u8or66zjUsXBZQ7yZCwuw2EBtuntT7B9g75ZRxOFYO2Jq7OX4XqXT+1jxKqTSjHsDpvWMX
PcY5p0186YiMRTT5z1zLSiVclJerpbuKloZhPpAqh2c+jKpjP07QMar/IXhbCJJrSWll13GdSJ+T
qHkgoPVh73IXnPLM41J0tVdEks2yYJoK0k1XRBARQUoctRHk/AYaY1kYEmgARb+zbbITo2ALRrx5
MrA2+lODlntEWMw67ltHn926EliN3kMzNiHP331JM2PcTh8QVVGNFrP7LTY9snor73AbHRX7elRE
mU4tdchsf8gxcC+D8w/aGvMKnfEvlL1LMzlOGMX48xKHzo7tIZBM+SaYkZm+5FvQmWtEv1J/Pvbn
IumBDhDGK8xOna29MMNTdP7LT0XdGaysrAMus/wKW8rKYVjrwAAKVn/zk2YmEmAFblUbz4oHkv64
VLwScljeUJQrRy+nUPvoPAi0XEwdc8Y7xagKyXnqoZegNTVzUT/1wMk1Yw4BHS7m2Jjt+wmWSf3C
aBUfC4Nsrh5qvuxduM+tw44hyIMo0Xx9f45ubeOxiKXRexNVORqhperU17RjsdwOhn0QRHnfJ6jf
50Bw1+IEOIMy3h+1QkLx1Fdff/T2eYqvBR227chsFsIiuPM2M0pYDXJ3E65pXLtDjJzRjeur2/Hf
MhYnMZM59JNsUszB3L/ZUl+J6ZOPMUJe8psUP2v7GuxS0q6oBMj683HU8jQDLdcqyiBPr95uAWLW
feoLjgo+9+89mEzvc9ZFGhNTIaqwBlhl3UeZoA9newD2Vu3yhixsxB65DpIgKAv5yWi7sxpySggw
S+TYNaFHamm/mUD+V8n2Rn3SgKva4ea3IvRjnXf/4hrdZ/QHfr+8pxwjy/ghmj5bbt5RWr0mwSOw
6Z6IcudWUUm3aQXkRvbis6rUxLxxNlHdgWDnvca2Div1GHI4UYn1Nd6zJ7wUNpdPYiPXBaDuwtcV
3X4gI57/yJnV/VbDyR9GUBLJ6HoBm4HJ83vn4hcewZzI8xjrBEudBzkfkUGRghFRBxxYsRSiZUqT
yN8cR6FQT1mynI1GTCh2geCe9uoxRk5cim5KsNo6XL9ENxtpmq711t1xLrgIVMTFT18h40N6rv3P
0mOoyxH82ugrdOOL4kgXD8r3LXWqwt14vtccHES4GIpRYJ9yz8JJuyvykqVCCOTDwHZxvbJ9zCvT
+q6hsFlfrPCEMuxQsD48ypYtwsWQX2Rk4IeH1Vv2ublqc4xQ3TFli8iXyo62yufdoApnd23L+AXX
17Bz5px+J1kUl4rsoT78VH9cc9yVT7JfqEsx5/EsKqhmfNksaLAshiwH2K7d6znAtCV50qn67Agq
l9/z9aBQv8kodRp2+n6mXAyGuklwPlpx8iRl68+hq31SbNxRdWCHB1YRpMipgb2QciPBs1TsrfY0
+h15KCuP4iW5kU/qJBNE9mBYhsrsq5XeOG7RLSKKa4NkmKsQadM11ckSD8TgewvWX5YeSFtQPvnL
hj4hEyKTQQUP4kWfYD1VlZDyFMZnER/Ne++f0w/vYERL2HBIZ2TtRUWgEcoNdlqTgtNBmuFSq8hK
4xlSULLu9/rbenSeko8e998yZFM1xoVuLkbAaiVZOdL2NzVqez+ao37dPqHiagRjETq6JoGovZc+
uXjNG1T9aREbxe70a+kquOZH/ojLewvfRaq2urfdCAEswetMPVFdwOb87TgImvL3lA9R/Kn33v33
xA+M6nMacieVcRnRkwqKF/8nGR3LSck4TLaE1wtcQyqEYyzH8St3rFuxTayHMHFqM70jJZkzFK0y
p1NB1jSxs+ateIDLPnDc4EraQ4qOlFAjrluS+VPY5HMK3kgocuYReYh+P+h0y+Omh9rBRGRD+zqT
UCyc3GWK5PheymAdH2kXCJiwsNpo6aXw3CLW1eP+Vb9AxVUjAxqPwMh8zXr4w9w/9zen71ehvDJt
YCfcH8rMhS8mmeopEcT+jEU9bvNDTkR8DI0T5rpo5CqifMl+tLOfP3uqbjH+rPqWJLxQbKQ707n3
jC5QQFxERwwePhVAA21085NfihS5E3yVTZSakkaU4G2bKIuUFemGRkd6lOeRSurQti8Ne2lE4mC5
vnwXAgMz9zEKi/LV/d+gzOB651c9UCdprFdScXI+pR1TFmjDkFftmte8E70UVfv4f2X64xcTXOWr
iz2+Qzf6rw8BM+cUj2TsTIcdmJQ2XApMqbZ1phypbFl57u/kS5mfMRbxBG0erhR9bTdNL92QAm5q
zimS0AsGuGzkkVo5/y+tahj98Vtc97/mFGRNOZYyzKg/v0dL59sPc2NVzgKzD2P7peONUuY/kKmh
nrypXnvMbgZ+RgX8f60CMNOym7Yj+zyp0O6v4dnyI+QrQscH6JQ4a5frpmvMm2Gbnr7Tp8Q1U6a5
9yEnNBrvK25lbjVFppNjqGdwNHm5g3goOms1NCnMAlAVb87CQnWMCNN7c4+2G0tu6jNC5IL09fqO
1gjfjmbuiv8wvyd88XaCZYQ68DwBqYN1GRiBkh0BWrMY1v2n4zOhd9wahMV8Zg/neVnhjLzlr+qs
WvOt/+nCYSAREzPf4ZJ6IT6cDhrKGnVMwQGEva365vgI6uxSHhh6Tz7SgGNOFwYHdAJwKKkRtNPK
zz7mT9KEetfdZQXa2pGZTMleA+sbt3dU4Me0yehTBM9935ByMzisHUftuEAAHqDzpcDwv1HH06F0
i9wDB2/iOm2zhyWd6aS31FwqyJpOIOyK9W8pYEnxAsUmukIFWtrTlf5hGqaZa77ikJ72BOgM1a9D
E7f1j5klIatoezP1rxS9+pzup/Y5HXgl3lJzvdoBmUGQQn4oHPFWt8S1T3lLojK/RdsNaygD57aI
5NXnD4rsjaCdC2AIDU4VFe5nlAE4V3kCtTcouyjLGEKsj9enJ6/JpvfwarSzNVJzlYVxuok7YGKD
8kVrFcRoQLH42nBtkO3JTpW1ZQ5SN8pct2ctqcJw1EYwfzb24HKlT7wrzY+o0ZA+4/+k0gLnhEwf
ew1JehnDYjIL9v8CQ75BIbyjju/29/PC+A4Re0rPzZ8JLTof2rjd7+6WCGdoAv0rE/l7PaqR2Ept
5OCfPStmSRszdXaj3H4oim0iNDfkvXkIAV12/4upDNiQxeeUaJAEp4dwLZudOFJfEKULwRCjJWyA
OrdKXBOHIMkslUjOWi17nRl9vBw/RVx9xLV5lAoQEpJdsLSFi9RAzm1K5y4CnLCBneAxq68T0LAH
mHCLWI+AhmQ71nTNzQd8m//o2WQEmjK3CcKYc93v5/Ae9DYtxrOzzFiPjhg6Hm+Xgw9L7mE4HRx4
bfFKxzviwn9tONDcbEsY04aGjHrPpp/J64NUB3zD+V3MEgmY6/ajN9GNGRKRmSBkUQKaonGHfAuB
GAMCKdRuwyNh3DGXCKPD4q4zWCNSx4T9eLheFxQ5Y2ZS5e53pqzunVL+vuq1RWb3P63zO2bXtyfh
pGTOFqum6dIoArRe4lG4Hxih2dKUBLoA/SbVMHWuyyReX8J+M0eDBxHbZ3KOBUcYVbGbazYY6Xnx
25tX0e/6hfRk/Md/u4cfdnVKxTC/pOkBll46lyGnpLBWm06rYW/WMmpBQGW8qMfC1x+PrDdi56kH
ODFG2/jsBnqzcuu1Mxam3YUN5xqeiwwPf9qnWimzQ0BqDmpLf3LTiJCs5Dm6kFpXPaoG4EOAOzvx
fgeG9xw3VWSy2kYiX6/i/mKD/DKc6f/80miKdjxlZZE7vdQoq986q0uFS7h65wklop/I1tlxTapI
bG6/QNuVbtX/f27q1mlcfXBSOos0I0+WzVwsC56yY1uJrBSwKospdkFdno8CF67fT6Lcws2fhhRQ
VgS85EpoRiaQAIetFOLQsXMAANNOL/9JCNpCHCkmNUi1yLtunC2+zYCYNqyFYf4ReebEpfBqbwqF
jFVDCaGlzBMADo5R1Cd16oGU1zgnhf99xy6vWoxX+I3Wcrcd0UJFla61QwLUkVTMWCQ9X0zPfakI
7AOzKVJHjqjSgc3bvdOIqPAv6YryezXLNRnvUJEHnWYXHW4hkOxlH0CqVsAcZjrgUCanKmj/xjO6
Eo5e+cOSEbvE3FdQ/tv42d5+hX+qEhJQ4L7BMt0SG1M+RMz2mCncN+jXJkdcpq/ZIxkiwgQCLvU8
Qmw7DZiVGtLu2l6K5t94kcp3hqioowvvmwTFwuAF8Gywe3snYu93IPdj5n7hiPLGmFnEwvwUy4KC
ZqSkxyxBJi+gACQYLPQgVrsXt5/vhqx1JRDJD0LhpThsMSnBf+Ye0EToZmvBVDb+EZdMGQWEFdMl
dYWhpdNfT8Nt1nZoYSxIwDGdXKSSxGENm2X3Yti435pot311TRLcM+BQscwMtWajryisp314ovnv
cLljgsXPP/XgaThcryZEvO3O/bY3X3z2b22wQZpCD1ep1bXl0jPAIOI9kGyhRnYpyRNwaztHXZnk
eA71HxgSGSghOOsToZ9Whp3Ar1/GdhocPCMLdHPmJ0wmc9z38+yAQNXjEReHKKtlTRr1962Dqr7b
aQyvug8OR1I6FPsXM6egGl78mwh3w+dwtGtmrSuCg8ZkSPto4P2dn3JuXQLbiyNrzPdeV+J8Jgmy
Db6aDbgN2o+L1gOyVGAd7CmB48eeC5s8czjQv0Cv9vV/HsP7sYeqzm7nebblPitGrAg/ZLOu4HN+
V9v33CmHvzR4Nzm/SzPZRzHtFsVk6RR0DyvyxkTUbWoto2tIAwBlRkepRID5FHOwsIzfOO7BnPAV
oYYMMXQlXk+faQY5XbJbr8JnOGK22rzx6mQr9r6PGCGryO9vmb3DdHE0HDxE4WHvreyrcJ8xaOL7
9dmtT4qSlvyJrLPr3bxyFcGxgF1rrCV1rKf3d+W3W9zY02HqfpmWHetYHI8WACVux4nco4BBM+/+
G8L7bSViNISxXpzKoO8kp+owKO3uvgtE/qvrPF4VJt9X9jTwZc40fWv8BJRDIcbljiMjx0myCzu/
AiFABVuyI/xMZZ/jlw6yDPwhb5ZpBOOU0kV8d3fdUk1hg6ftGJr0Ozmr/9io4f3UOtnQyVYPOE8O
BOQI9aWp1GYP6CGWdhoxyFMqr+igg2Hq4MCloGJXBfrz+keiQCidonRiOd5sTtM8stzhjd7m2X/R
Ql5yEd66OPP6oNIVVOXqvIbePyCc9cLMbFvPvfRTB7gpjJa+ZkhsAuMj6uU4mjnf6fJHmW1PD+9L
ZFidK0ftrwz3aT+VjpAskD7vYYLn5AdpM+j55ewMNYjYVZt434QehyBGdGRnTgovthW6YXoXxm7N
5Y+RuO/uBFOUP7FAxBYzQW1SfLl+WKkwMCWy1AB3iceR9Arte7gmicBhrVZI7LB9HWxoxG6Fndkw
1vXrGS+8nNGu22XAe62cv0TVsVtBcArwhynr5sXAvMFMBzFbrQ8F+R5LzlIqcHw4j1fkPWpxlw5/
LHRNjNsNGc+VyTye6DuxTR6lCCWg1SFdM/Nr/LzciK7heFvs65crWMp0u4x05uMFvX9bye3TFASZ
eJ0FVU0qXfOEi8CNU7e4hu0EwALBUOmkh4JAGFmp+HzA84z2CeaT6YSkN7KfE2CAs4u3S7Gz69s3
LqHpcSCSfWeDQUtlY+q6H6JGYXg+VkuxG6EIwLlw9GMLYdMA6O/J2Rb5wyYtBYsUVuyiyq6CwmQE
f2OcOQXa/9W+I8kt/MMyWsBoK1d67pp0QlEaLL6HoAeMV58IQMzRPz8nKsIzzG9kuRifs8KuuiU6
HhijMnGJsfG6Jji+W0+Cp9wh5tHNhPKzDizQ9pGt4PVHcib5A6ZI0+Bu4Ftd4/pvGCDF2ZfxcFwC
4ZtiSEFDIvF04szEUKP1J8jF7R1NnfRaarVbgtCHbtCM30SqnZjOpH9m/4Ha06euv3O/ZZUsTyDv
sDtCjS4CnJUmRrCwEOUe0x/aDPhUmxptRIifnRjGpbZLpzwGwZSOX9SplqdBj1tUXtYX8FbzWPgn
XZVnpx1MeiPCDGn0NXNND4CQBt5hOsp282VHpRZDtSB/V/rrKbPvNA8KACZvM8UT6Kf910s5qZz/
GJmbSlULgrO+cHW0H9qK/v0/h6Ea+BXCXXM/p2+2+7a2ntbBXm4NQN8S+I/PVUQigCRGdkPgdjSf
qGbZLNAOQSDDeXc5e1twK7Ahw3vqqktkTCWkFJuTUvrlPfbyadXtVcpHEYHZzjiPehTnETDQ03fw
DNrDavt63U8Moy5a/jVqmxpnjk/oQoFUqWGGg6yVbxOrsdxER9hKyL2A+lXkuJ9XhwNJkbo/4t90
N2vrbk2gCQVdZvfovA3ogjYl43A71Lws7oe0O4gqYtnGaz5CeDpFLFus7LTracZrmSpIIyEqFEPp
06tGgJx5hGjMOHQcTSAQUxbDmXTPuUKbUmE2L26GLcH/noVg5eNPs7IIQSQYnmkMusxqUp1Xql7V
hhGyeAoOn/nPhyjvA7kFUMLVJ+nCQ8LRv9rDvbveGIeUq2CX4b05nPPoldDPgcd0pJRdMKn2p3wk
oMAD1VwthbjCzX9zffSAKYkdkSMgFjK0YPd5h0wuMy4kFME0VnvIKcTJmrhBw0O9dlIZJoQD+Mhd
CLihqmj5bpPmltGrBcUgQm/eKeenEwgIqMPv9dqIaedgqstl7N7YXoqW3zRZa+0sg0iTFEGd48Wl
FyliH5s4D2WqcFIp43ZhkEdNWAugeBGHAjdsjuLNiLYvADmduqu0H6NBmuI8pm0EdeTsFXL9fjzJ
HeKxg9WC5ELbe53jADGWrwDxgk4Ug9uobigVsUduwVnfvdS2eebVKBI4MQiyKg5cVu4PzFHapqWb
66b0jTp+640hw4CU2ksieymSetdurwdf7p47bNl9Uvai9cU96LfJxDorHKbItYCMUwm57mXX3fAe
n7Iq/dWd7Cj4Ovm3CALDvKWMpsW/VyHY+0nIGsc3O78Kk+pInDBr6K40GS+3yuA6AyUzdfYOOlgM
tf8aM72vYx1O59vwmjzBLOMyfysC+PWyXe8/X8/dCenfxvsKs43x6Iq953pjsqHxkyoPUTKZu/9k
htanuvdy5VjM+T8Or9TXgx2IH+A2K/B911QeyGQkMZkT88p/HOojcAfZgf0WSy5d5VNbEdcqUYKR
EfuCgmBYSRLg6qhNLZt5uj0lb6HXjGPClLuzhWo9yPhh5lcHpcqnsRmRgTIF6/v9HFMIBMwuwazT
7N1LlkOyGeCHQB5f5vIMEJmYVJlrXkzDJvpue0rHUoqjWI35yY+EVIUqx7dVpqmDPmfDROPrRfZ+
l+K8C4cgrQ4SfOZNx+dEMVOAk7kIxWlBzH+UBS8BGQC5lHhK0CC63v1Yap6u3YHApseC+gIPd8ev
iFiVgX/EpQaTOYf5IQeANlRXEwZp7GIJNZAa89H8HNTM8TktiQ/GqRl+hGqZ0CoDA1jjJvrrCwqo
HH9heHRpqVgP+CDcgUw3vPG7b8i1eqGGLw/PXjxsCmnd+dg/rWPxV253Ak+AjX8Zf20TQmG3625Q
BlP8QqJ8HYTi8xiFhOq/XDIthO6lSICnk85KSX4/ktKMvdQ0PtCb3X6xbhQfg/d6pdkOF6bEbhFA
urKE9JvNXTbma6qDGeO4oltOucneBKb7GhwTGJRIc7QkiQF+SZebiX3NzPQvjP2Q0ZSiYfIUDnIA
7FbRRsYwErsGxLe/LAwYvHji0Bc9kjaCQ+Jr+26vmyzQ6oMgySP4v/33k9o8eRSO/QBT8HbC+akC
4Qz69DpOWypZCurfLM0rEmjjV9jMks4v12rc2/NpvNS7My9vhvp4CmysvH7TKF49fhHOaoGTwQSp
WK8eV21jst6QpRU4FlXDko1ppreAsPRZqAbcLLvx6Gtd9ceYgfuDvm64yHJb83IUv1U+Rpt8wkMS
z/HpK81z/W4B9C8IyKXX9645AFx5kDj8Sb2Y45Vo2CLiZE4GH7o/+rZLPGbpOMSCvwQf+LI/klca
NbgzUbqJwhyTqS27OvE6TKW+KlvyU3kKh6JELYNjsGLWSZqj31/iYhySic0Q0CiVv0mG1Rq3FLgZ
qKEeoPTWuKkS/0FzaA6Z5/s6LLXSPQm7cLhlscvjmh/CJOkyCmrnmLrQrfBccpzhHGdkUeruIxxU
ve/O4o/A20PRB2TU2kS6TYBORSmFpRhJA51rau5o4u6aEBtFpGto2a8MA0IvsNeKHEFX8vaewFSb
j2dVZTsdswgtWv+TJTrfKfj4qfvO7H98z1Ni43QVjkvzCeQVUxVh6XN80aa0hW3djeNmx2xvl9xr
UU0p30H9CcZ/AR4GcBTG/3NE8CYZ1DP2VaN1kRtLUftl+ur0FnPo3KD6rs/DhhmxyRGK3Ix4UnGt
n12JmXDw1jGGQ+eq9lgp7UZaAGu3LOROCcNLaChbQ6OqnBbEa5AkL0Uc+ciLiZkXimTkVGyUBDMM
NuXdDWfJafFwCpVQ7w2gvWHkhtTFNv5NTk60JmFt41Sir96h7aHLTzZcPM9LlmHNoOboG8xOP+/m
H7kaJbU7QzAliCkpWyI0NVz3DWF/FGHnfnzl9Z90t+TwLA88OcHG3keqAETxax4TLwnxmsmzLpxd
ALD4LdMR5mt346ZDc+7Wh68HyOZh99OlcCSLcWKuuUiRRsIFfymg+QLUi/oq+jERtcz+Ij8GB8H3
vliwzjLGyYWwfV/PtSZg2YE+ecZ7B6nSPIhwMjSBAzyEDfO+79Nw5TEtbtkE61w8tK1BEu+Ypole
mK/C7fBeg7sMYBgT8j73wHzii7yrqfPrlcM2XEckHSei6TRkaJaR8JfR6JpQUSK4D30idNy+pmoX
MJWsdpwndS9o4A5PhL4MVOVhy8YbSd5qi3DhBOGcaX86NIi2ULdlQQypP0mfwf1Aaz0Qr8ZN0xeC
Wa+v2L/g7QCZvBZCTmp6JvP0Zl9xxDwXEHWzMuRD3UWZrkl+Yze0AASkvL/8lPRq41AJKEzT4il2
dvZaOEK4vLRpkINSTg7ZiwGJGEDBh7OugnjNQX1Zgi4X6G09KEIoEKFYP56kg2BWcme6Tjl9Dxaq
/l1NlAEq1ZbDsVCMfyZWi3mDix0hPKjf+OHpVgCA39oDW2bYNx44oq3smxwHGQyTz5/ntbx5cXCK
PhIRhVDdtmwJ64QdZqOwuzkmNt4XjscUIiYmaxGD1bjodeE5sIiJNy0RVYDPHTrtpkLlhqWsyjvE
oSzk5Gh7nO3+RO0108Zcfez02Em9ZFAFHTiRG2NQ42th2dZ8bjqgbhCsfGOJHpmnMHPRB/LCFoJK
mFbPt9Rg9J6KwqOGSTEWP6g8n8L7KGTG+7UexLlubS2eqA9ejhbiAXaZDuuRC06qzXuvyD1zpvJ5
kR19qEl5aBn+O67vjTay7s3Aa1kkU2JJDX5orxshjSmz4TwCY/wf3yA0Jw0GEWVYb3gfklW1c1J7
Gs5OyAukg/oTGrdDkW1HFtX1KCkQbB2LjJZaUy8AWs6MmAPLNOjo7R/lOyJPxzENFPvoKmf+jocP
mA4XSMVWdQXOwLe0kF+WJ0/PsOPRE8bgRAJatvU+3R0v6EmjQrhT1s62LXshQOKFmrOlj3V52D8V
O3AzBAs1OlgkqeQJ5dM9W3BicZdWQi9vJdb3pHuJ9yucV5JEJHQ/J+3Mw9ibks78h1LT8MXwXqVv
vzFXDNSwatMMOMDerb1Cv1hjkMllyJqkzcMHWIQGG5qJRgS8iei1BExJFGf7Kuhe8by+/+tC5+P8
fnO6a98NuX3ub5pqqs3LawN6CoMuRCXl+k+ZenKeHiWmQ4BWJI7uxWzxHKt7wa4WzhaJhcaompb+
MbaODrbjvrfXztsL0LaYGMBBYMTX8y6g1MHKwUh6FWFgZkhaVqQs/r6Gcqhb3TTvJ45k3XWxk0ZD
L8P0H4dnFNKTJZ9113U8CjJ/LlA0ehG22JJuwh1OMC/6AdEkOgoWA6Z9Iv6nE2Lm7CPT51cFoHB+
TOdCKh0+b8UI4fxvrcINL5+UToZLbWmvV2cqyTN2xmugjwU0VDjGOqW37kmYRe7KKBMEC8YSWQkU
Hv4IaSEZegknShe5k4GJrR2CJa8QJHmuHOiZ4lxddvYgtQvEd0nFNqT+LMHxcoUCqxCUeM2YyJHB
9kJp3W84R9N2WkOQnZNJ2vPlFc7nFSR7Tk9Ymq9GxMMnRpGT0KdbElIltWUxfBEGevVgl/aioU7R
CMiZZ9z9Jt9oU2VxV1gG4Yu0OTStC6L+O1++GJCV3yOQehST+m2CI5cd4h1drdvtm53hQMz3aHG8
8d6I4zv0mPropTCSH4lc64qIu20BB8JgotAmFqP78ocSaDmhFNZWRdPI273ndzjDz6SwH7WEWpZi
nw2Nh0GN+krLlZ/i4LaWn95FS+zzq5IjK6b53kWfomqvyI23v1h5WTiTlbXyPKZFaZjMjIpwdVDj
RVpvhLj9i5286IthfkdDKQ5vFVhF1TW5dLKfiGOyf5tRLMWi8uCLG8eOhj0GcwBOfWz6OsPfVX0m
JNvfxbtGbXq08BUsk9Cx7DpDDRqCWD5XJi52vWsGWlsfswszrY9h+AgwqDeYqhMMnptDObabjXn7
KTPhbAB2gBGvRrWdv+vZBJTJ/A18JOVWvkAPq1sZ8q1zxWYj8zUAbeWPZESWKRZCm4jtfxYCHacL
6yvq3X8ngb5yBAOK0nJK0KCjE72DQ5gQzmKkPOhRR2+uZXFl/YjYmMTE+plyswV/FznOqpNxuEaB
aK8zcp7fEGgKHJlI/CT/mX7dC6Aelk3vLSov4ZsN3jR21bdXjKYoOr6xO3sl/H9Dmnae4ZVgk+rx
1yO+YvUC5lwFJWvApwID3LZo2+WH1XXpggYim9v3HmjCQEcUgos2H7cgszRjm8cPFwWSx0Bq4gEk
/v2M2RbP51+OCDA8PoyXWig0JtQ9KfLNJKdEhjvSf6ha+HA+ByhpsZrtSLWkX+VDrTuJH+KdaRMS
f6g8bCoxIauq/pxvwMSVdEOisf9Q4trZGyPep3yjPyThqLOHX5qiIkK8HsAgVoHAcv/VPSc/19up
oG+0O0zu7IjsnmbpLBXkBMMEskpHq2NqE/GRCxxqRHq2CDQDodpvF6tQOfR7LVIdkVTKbwaUUTP6
5xmeuzB2Ne8WAwx+WsrFfO8KeXclcXSDZqkO97DVRQOjRU2vPn71AkD3UtyOtAHsIym61yYkF1D/
UPmUTzrGVaHj/S1I1yPor99fnS/cd7CmHk4DEen0+WP88hqVJSRXdzump7k5i7lpD/1aT7SV/grf
/RNLskkDwqKK5bc5PDej7vUTlx+zmF9OiTnDsO7g1vK57sNZnbQe0XkDbit93HhtmT/nVlTb4kYV
qtcTy7kHEmojdChyHxqwo2OZvzdPpkwfjTuFfg34Wt1BgxG0+tQ5O5KWT7c1LJ8j5AJ1834/cdoN
WqgxyYR4IUBDFYsKGZME+cqwCAyzOpq7No08dq5TkVYhWdcZ0Marmt86zoxnJfFTa3mG/hJ407zm
biWCmWhhtmJFO2L7mj+8nA8Cho7d3D5Zyj2PZdiP5YMiEeQy5s1a8/9s5VEz9m7hkmGkdj2W/fzH
4R9XNyh60xAbAKMIzVZwRJgPPLGu613pZULPVd5OMuaxsBTgPiiPUt52sbiYuGa5MzBiDbQM++I0
LsQmGXM3q4LoMiOmNOG5AwQDjd1KUUD8U/y6R3I8+AuCjAc38oKM1mxmGxQRmFSHwwqzhW9YPxTp
65DnCigBjBql94L2ByLRRdVl1AhhG02DgLCEQK7ZTZ8sqGj8Q0+9GdS91rnmpJUHoI2JOb18wQGN
AAaozzbJWzgC1iSD3NjQk6iIzhqhsBbKNCHU4PowY72W4iNFtm88CF2tdpLL+WeiWi5Iwi9+rXQE
L73J7Lfbhr9NUXYwCwTIrYj8hLO9a2rsVjdeM3SYwDpZjEnBQzS6hqsrJtj9Yp/LbySk910r5uK7
NpwHEF3bA2wInEAYp9TFNO6abIMq/IsN8PEj+OnhMjRogIknJMMexf/uAKdxrwVyAkmcaIlXfBVs
Fe6GJLAvHnS+Z1D7DxA+iUD5hrZsTLOJ6EmN1xLS7y85ZQglta/aW2Yzi9fUdvxBvGvK4Z12e1va
f546DnEmsBZVRTEFXZV+a5fxkniIjK/gGKKur3gGsZpRBLXBy4IRqRP3NK4GT9RyxJcmLm/x1vIg
b2mo1piBzPO93eRoGrimfdOXvcnztbGwTKlrgBstGTmYMa5rY63fArwAYn7qLvltoyo8+sbQron1
I2/NoStovzq0hanFpLLBodIKoPi3RWHL0bLbSaQd8YQSRH0NMP7hmzqe/7x+N1cBhbsUhlUxpCNh
VBxpCAAwAmX4OWjMEFso8XOpnjkdmrgE2HWYSGOujSk5F+HxNiyu7dyg8TxK3NMe37WwK4V5lo9s
blDuFUsYxuyCTfd5etVTIFqAvdBCEbvx+py9XHAfhP2tEPO+w80IMEE/3rDTWx5Sr5ldTIWHeVqv
rGpT3oNcWtva4UPpWqmKpxoWmy1fNR21ijIR7nwTeuhRC5FutqKK3fF3Ri22R3a6lgSAls8BF32S
3UBUMOLqYMXJ3Ks/LYUOCoJ71sWO4jh4e6F1Pf61/4dGYxL1JLcYW+G0Xlo4Ii2bHuRhPjlFGUs7
AYH0OIy1dkQ9gXrcYU6ATtDmHpGsZR4cMxDrUfgYW7O06/aT1fVuIHEdsH/+nwmYksy5FSBLwwqS
1UwkhBwfGvolszSqpnAI6peOe0EtImcDJr187U6jiz3MbzJBU4kU/0P8iL4hFvG6znjo1SdD8vCd
qGESCFA1tjsFyr3DnW6fPkXJSQUxklfTFq8I1NVRJpUyU9JHejqLvri5/+4HOqk2VFwSTphTpeXc
LssH9+fiPJASKBe/klFRt7mWvmQ0hGSletYVDYNKznI82EFBfNVs0duorrzUvdEciH0XtziBMOhI
K9TjyuPxQwQ8Rprz87bDKSmgz+lFjPtd4wP1UOZ6B66CQJE5j4Gv0WkvstsUPfGDVlylR5JT+6t5
4hG8JSuVNX6baj4TYmmQA24ocmHBy28sf3I2UnhTNgFRsJUyHBpXzXrE5WNiYS8jxmmvrTz9jZ8b
Ju1DoKs3YyfOj9UUDwAk5arQXCKtAq82vYRyT3MyEVD0ljOyMy3TffEihU7f/ZFlrFaLC0K7SNSG
QHuY1KivGUsXL8aO1xCYTn7WhctCUbMZAU2p9m/qjkg5hXZIvr0dsSPSORMOgjKstF/SOShzW0vZ
aaRxERzvQa5rLompiiM90oE0uKXxzDZLcdV0KBG5E70r3RIRzoAVxmXi9FnxTIkickKzHMmVusE2
pc7L4a4CybAFEhMmCHpWz53ZkPqF26189SNLzq0HVTPptvgZvDOHCbNhGXISfujqj1iTEhXPsE9A
2ZGzPxJ/jsDBxJCa78NwqJIYnHtBTPHmICzUNxym3c3C4KC32ieNf4QffvVPpYTDxqXpo0Micj/Z
/FcedT99yKWl/eokF8uFH4e0NSxmDeSG8a/Gpr57xhvT4XH8lXmAYVYAGJxqKk3gWPi+G6VorYvf
wf6TZ3HjPflQ0bDhLnxpSU1tkOvr/grCA/xAzZC+4tA+wWz/eee5HQhS6lnU/E9LG/dV88fBKK45
91XYoPsCFt6ELH+S3/R2lNRam1xDc4QJPf/FJTkmBpoeZvrn3++6igspCfDM/m39uyCiI3TCuqfy
M/s33LVjK8rHQK6t2fdV47gbjqvkYiSxmBjyboUQl4e9zhTMP3zMTWPc8jcs3KHHf4hzE7FkjpUj
CrfbdBCmZKQVPeM5hfKLDabrylRJt5XSmOKKvyqb6NBJ/sf2nx0rV1VeelHI5fbqP1Ip6ssE3uUU
6JKyJ+BXeGMlE7hcNWVvJcE6PWIxJH41WXaMutGyRDkXFo6denhMzrHSZUuYQReNobAU5vwLCjie
O5cUqjw8RWDvj6WW/ZzBQwkjnLgPMBpFNrXmn7m211XRu1MsOJ5gvdFoy5e1N5RdhZkgNVQvgEca
AfebUO0lTkOwpvN+GQD20jeM43DR9+rbmi09O9ozMBLjKMLoobau5EDkUTi8h9Jam+pSIG6qnRcF
8kt/vlmDkZz8F6OH13KBW5/PFmG6mniME8LtNRVG2vA8QLwV7Hl2QXkYxQTJ6SxbabadJZ8gnp5B
HI4GtWgPvKIOa/X0ycLR+sj+zzYnx132I+FY6Wgtj6CK5DBOLFIXf2SxgpUPry/2Cu7V5c6eEUOW
mG+hpZZVZzblXZZSm2la2pjlzQgg855bZv1sMKOqwZitZIlpeMqid4pjVRwBxmmCYwCP1jSzc4jC
AkgWArC41G5mIytEZuh1hQir809UYZ/iGp5RuWxxW7VEjf0gT0ekCzBnwINkMf+VUt/jy8W009fF
naSLPMbYktaJbJefyC6FyyUG4MOMRK0WvsGv8j1nTedT6ykKiptXpGCBWoBmkINAIiZXRG9hUoa6
ytshK8jUoUxaEf+OvDyrmxMlZKi8SOylO9mwvMLKVBRfCQ4Y6DEH4YJxsc6oJvWoW0M369PtsIBQ
U1PxGvm5Y/nudohjXa9wxojyNGPLimsRy/7k+rDeNpmfUOMVsYtHn68TSPuZmDrrNyHepBI4+Oai
4mkIWS2I0aCfpCj4L+zyYBmKl93K0D5tKfg8UvOkdPFmHExPtgnr1xcWORXQdaJKBn3i5zyqhS6i
3dUsSxqrVDwT5Zd2CemwnxDsh5ffZwhIOYPvqV8+N2Y6sgDg2M6WSpEbzlDY+kYCjVwa4KJnzls+
Fdym5y3dUMkH/WFbzfXKMixn432LgMVJ29LMgJFokJ7jXTs6MmDw4TRtReAJclNyeo5n13calP8g
uggoBmnbJaQejS6EFfc40UWo5rjVfZqTfxghk16dTI8jBcb6g7WamDXrLKZyk5iJpGA5pEvTmty7
21m+hJtz6/oQlasKK014Rvrlmqi6mHEq306jbXd20aDMWWxH6NHBAAbKVopSsJza5Ul5amyyqEOX
BkgcerSv5XlEya8EGntivGqqhMfLQIMEjlVwPvG8kdZuo9SVWIuSvMR9rFG9UGTV8bFG4LAV4yBk
ZGfF2ZXUHYiN8tFNGzAgbWuPbxnyP3akHM0nBSGkVh1GmfLMY0U/RW3RGUNdMWSq3iKcf/vCB0HW
Ogqety7enJpu0VfRFBrgvVFK4CNTf7ec00a5FIxsQRpxCgDpXgBDg/iWIpbV9AEVBBHtsgqJmERQ
XoYP/moOKlLXgoL6iV1NRchRgpTG0x3B4TT1W+Vl2DyrLdiNutvKryYRbzqVnGbfZtMtyfoU351l
Z0JeIsW/zbYW9tLTENkig9WlICsc/BI40pa4mFTXWbqKzsPceNTu+V+Bxau4dKY7Tqb4v9Q044IH
EA+jdeQdkExiG+H3JIFSLUUhkCA/SpSPbp+250SQd5dRSYzOEZkCl+v7vGCMUlYy4OKBbmxdX/fY
aP7m9DrMA7aqSlCY8Tncf7mRPWTiNNhRsVWd8EGBaZmRcqBLRGjB3Yj6A+0N38pmbDMR8a51NzBY
jPWW5ufyZvkl29ccLdm+xOl0cnNSoC9Itb3N3YYMP7kHDI3FyfbzJczhxyynH43HxVjF/n6PMPn8
Pit6+X00+00KYMkL0fPMq2JV8ACeQ2W0SP2YsGls7t7PtpN8pY77OQNkCdFrToXzaePbn1InfAcG
wWmTkinq9T8rBqgDNWaxGBfDZnFe8VaaMXMXIxLTgxHL6qwUA1P363yHs8TzMRZ6G8va2zLg2rqs
S0xAxGXCGrYzCZkudTvO6g7pvo+sdHmcy2QSMAtegDrWiD/72tJrQTQwdiQyte6clj3iQUpSJKsD
Zn8uDFztlLW2Yc9N51Fz6q8HPaPij/YJvcP934e/8vQPIHNFr7RvySLZxgljfOLJvT34kr0q3Fee
OuQ3NTsYnTseqnrCnRVWgTUhw9ZDJ/JCt4hpqiHJoxgDhMcwQkdSVB0Br2k/ohf+VcoMnIQdmaDV
iC93/VKugwptVnlZ/KfVwEYI9FMtsVDBZCz+9CVR3zwvM4vmyT2JMaB360ai9BKP3TYtV8U05xwC
+6sd3RgoZS+TPfjIZa/Pbl7BmAqN5vVjMEybTtDENk+X3Rmzqe+sCHNy713hwUpn4hdhMbH4m875
PYh3ZZCK47xXd/JCihFC6+TY9RzpLv9jdl6zE3aFfxZaS3G41cJ6RYlvoDn2XJEmEwT82XKgYp0i
CmdvuSJ4zBQs1INmuTaM5Pf6EdK/6rGCLa+Y6pGATe1U5H2U+i3turvibEcsFD/guCegZYBL4NTu
GeUotengMABhYTuAovvmmD+PMSSVeSkyU6tpPPrTqCury7OfKWhmSfP7YHAvl2nPAWmd9F3OQsha
YlpBdvhCIx4NgrArfjPJYr0HsKlgZZOBxuuw14CXnrrtzbQyUrmBaLNPTAl/BBuDyJkWwsVvmNQo
sy0fKNTy+6xRtqCtbBZoUBZuBhnjdwa9FFAst4mXkNdVpWpmlcAUlLm4yTHX5opgisa9qOLi9pN6
ZuEK/pqmk9devXNlEE0Uv/plUmO8+JxgX5BhUvvCRfVqZebbMSFHO1h4/SBmCb/YCma34I0mvvfy
ApWV8+DeYdmh2bCssYz+zEyaUj3kJpv0W91qkywLlziuKiA8AuAeylAc0yClAaOgg0ifIr31rzOG
gHQ/n8Ayb5L5BLiuWH50+HHXw7+dZE7psQONUir8bfX2Un8FUUUxNnoUCM9NaJP4VJrBVxMJ2Wc/
wv+aP18FHMhU5ptoyYPDrVjSPVV4Zf82hCQ6ZeaONJkAdAe6nmlxQIDwbfpQdAb9zEBkjVtdgclZ
F5QyIRdb1rJnnANOSJr/L1AW1zZjDv8sLMfqk7GaU9s0cNpmUi1oQWUfHw9apaIPfqOaZzjqJtD+
XB2LOt/ueV/rLLdWy8fWFUQCofuWvFHoeKGpC86zi9pQVsUsXNu3h5laYfVsubLjjRPCZxwq3zJn
cfEs8d9uxf9sBWE6gwd8f7USxcP6x4u2tTWVPLDPdqsL/HlOMcN40qVGoP0jiXBi4AdJHgI8eZR5
snoXnj6WVxW/CZ9XaK5lIPFa64d4BayBFbdTJcXpAh1aLg+4ch0M1tl3WKRE4Gl4a+STqIhftrpl
aTnuYtWdrtkr47V08tUPRbNI1HWQRqLU/dhGPpqa5fcUKf2oItk3BQF3Ur7+t+bNlYtR1azgAbPW
8QLx7pGIlZaBv4cmt6nW3q3qFFhkmrZsQQJKHbMoQ9nfbCXEAmvG7K/JRCvxJ6NVfMPbrkJVLFVS
aRR2rcRoyenZi9Jkm6r4r0Gw36bUuyW333dJ1N+4X8F7Vrwmpx8srK4cdVKBqKTf5ew2nkomAIVY
nzS6gOVX38I49str0VR8ENUbKuDzz2iAv4CX9rDG2RL5xS6z+ZdzZawg1oWdb9+Vr64HQzeeIr1i
KSyfWxpjbXQCUgkQCBd9I11q6KgZQ4b1YV4NaEqZX6bNmXQ4Z1Pvu/hNIGkLXXUDGmn9rkhf0Jc7
hMQlpB95N5f7ZZ4pgSxP5q3UrOC/iVTXkTVQpXfGQKpTcMh9P1p1Q5y/IklM4/Gtw1ofKMPQRMrD
RY/hXm+nxBfXTv2B9mUOXtWIJzSx1HFir1/+d7q+JciU4SHLiZtDm/TBNoMrSlOy74Bdn/t8fsUK
Rar4zattaJCyzA13sBXcmC3/x4SccWDbMcckxKZiOEja4jDyckVBUYlIK8EaTuwtuANyBIw47O44
PeY/zKi1rwyejDFX3TGi/zrZpoeAmlI95RkPbSGxgj5CRR/UC/8y0UaGvoutDU0TxMv0R8RMUXB4
M6zstvcs+WucFksYprbASpUZkTavqlkFmh68DSZOfl2haaJcuEf+O8AqZ9HfJ+swuXJgjijwYH1y
ELPtn15HJXTYKBDQo5vFPs4LcDZ/K2Y8UVX29oQ1nx7xJtMXboMJx25VzWaB1DZFxOdxxJTsJJyB
O+4CAItH3jX13jskpjL1XNhg4bPEZomFKYSX8AIb1UpJpvwier/rCeRUKziRE0DJYu3tcTE5k1BD
+gcEYA5NSY3M2JoHU2Xkp3T62HJTI1d6X9CXmjz4Bz8fvGTM7ZxxLaAFyTVz7OXxZ6AAnckiigcf
HLIYc8UDp0GBBafBdsH/DxfqEEK/ccd8dBxmPSmdX421GrrX04YXqpQN8+Gfm4QerTgIkVaYp5KD
tybhn3Vt9UL983mILhdfezXndzPgMDm2j18HgD3DyymS4IytoUz8ON3RDbvcakEzDKl+foYuBqi8
ymjSxHApt4u+9uenwm+DTt0wkYyKUVOqyg9HPjybjOGrY4OGrvO/YyOgYiCoAc021jID3rsw08VX
oOGAvLmrPbkcCGTC2t3IPRm61jwC+N99p2Pm3LSKimhoXbzwQXSjvDcXJaI57XU4kadp6aWikes1
4MFs2ggbPX53qPVCrBCBuUyd6YTT/Q0S/pvDFL2mK9yCrq2pWHZOGciKj3vK9KJYwS86tabooCm6
mHfkKIugfWbT33hRh82weE8NCITuLIATvQ3RW+iiSrCvRyJVfoVsMVrUF7QOHXAiLcvgK9SO2XAL
QRYCa/RE2FbOeQ/BY8GEMwy114AVmMWLcR5FBOsvQ5s3+7aXbzNZy7J479+Eyl+AB8BxtMIdc/eN
ILmdLlzGZbROb42gSdX4AyJIO7pE7nyO+LCEabKV4aDUQYZM6Xddc6bEjGFJZCJKhbxXk4DLqKqf
mVMDqHlfwjprJu7yz6Q0vyVvXWai+/gTAHphT7BfNGxC37fzY1ng+ZRNG4KekNT4YpwFUkhlG8QJ
5rhMKo+ugBGKVKvyIAzJtLM48eEZF3A1zbBHCnviNbXdJmzNdTo1P3beek8gs6IhnsGo2PLhzlDY
yXmQo9iU3vU66fj8JItisoDB8gWxXRF95zKvS7dXPoL4FA9C49cMaD0A4bCgkJBCcfeVNKzmbMtp
gPV8TTGCM+oz/ieaazRCaiRP7K15P9Mjz1WSnLHEG3TtCGS0gErNP7gv8fezIPbHXGWdrm2FSbNH
RF6GjlHPwgXOMznL95uKn3hgFge07FGXmS11Ao3WRAG+kexEvUxPi6nggQmtu7WR1PbpF3lTxitq
X3xd44cBicjA6a0Q7ViGsfyY+O4NCz8Wb7vcfMtk3NhSprEJv0YK5hCe3SODLirmjnCdN4Eq/+Ic
VH7ktP9j0SxuJKLo2eNzK4L0K6nnN+i+g/I13G+xvI4cvJhT9owUCpDBdO9Ky6eY3vcZJB0tgdLh
e63//F281ZpKdPvEpcOKxlKW+ZFC8k8XT1fXFvdXALkt125wQpYFzO0a/DCBYaUsft2BgwcrAUMz
68oFN+3+w/dVoHDMEYxB2QlotsTNWLgaeNg4XzDW0SDgc+BzqV/8TNrymoQYvHpM3R2hHheZIH2v
R3G0uGNVI3TF7F1+jm9soLgc9CBpTzHoOUzdJud11N7EGv+ff2JjWYc60dzX2byLAWRy7yrWlV5n
A68Vzv99GNg7IZjkpRbwtAcAQwra8VA+sgsPntQQU9KUeZeIluWUz9RofDq9XEpeRp9tHWytcVc9
OnkoxBvah4lSamVZ+DydBHv0XPWapj268va/VJaw2vxTBn8dXUgxPM1XwN4jSmLuFVvyQ8qQRUwd
1pRpTg2djknkzyJJ/WJ2B9gqVyrye7s/2nwY6PXdMuFtzekta7Mz7rle0BMwGuk2TTQEzvwgS9eo
CJPaNhTBC3kK3OjVDxzvXugkuE1ghSdzAKMfiEEfrzO5m2Y4CM9YRotSkv0Isu2U9LY3ZKOEMT7o
sjhsaEoJZRdXzarJZDysYP1eFsbygbP9FD6tsxAeTfhzH+hHPrNwLkwUKludwJbTEFLSoT2eMbPs
9pFmh1wtMH0YIWA0IY7+WF94errc3HM0VXLm8C4960h3Sic7iwhveN1IvnwFTjPrhDjnImu+24Gj
rVnyY/ubac5YomBYLwczvW42AF763o7W0JkNVjnyYRecSXrMAGud+T3gxKFPGv4TYCJ52FLZKgDq
zSRddiIMSGMwfoNdR1wOLNnoz4yHV326jcW1s/XND+7Xgi0BFACQvEkGAcRfhKp8udR6d7Vg+HZQ
1pxw+8dJo+QxfwNahHgeMNoztHmbQsQmgSNek2IH37sWE0zu5TTVI6O/x8XUvdQYGHlvpZZuWUMn
oj0SknCwqfSLMz/gl0Mz6JaH79IQtK6QZ4/HEkg560rOBhGf9vcQCuWT1dBuwXwEhabPh/pJBcdr
cgcHO2tTlap0vgyt9kkbI1uU4Hx0bPVr0iajlgpfJy4BW1O7OpXRuA2hZvuHD8DzfNhN1QPjmF4k
qUqt86oUTxjOryK7yh+NCnbwoYMHsfV7yQzh+RPW+jPrjfIXFn2yeUGnWk59PtnoHrJ+M3/zx6ax
7FLqGUQ7Dan/SrlxNLhcjYDx0uiag4c3u1UGb8CooD+6FBODhMUXf0zzWLyVRuR+5e2+T5stJaA7
i5x5bCNAQcKlNuBWNcJtipf/Of0CT2q3pkpW09Rh1ODAgjqooItKE74GzakxXfiRDUTV+OudWcZW
sOrlrug34R9kda/PLhENB+fj1hocxQkj77dDad7NVbAGhpVClfPfGkjOx4wZDyLye9fRdRELsApZ
FsgY9HMl+OLWVUi+Kwkzmf+MbvFsw4XDfnHQmjtMTuvNyNvDyoz4B4b+Zf6+H1NP2PfQi4/mifjC
onCeCzI+QL0OgAf9SawuQ3+BkeBDtgnbMUPSx04mbq/6Wohm6aqVy4HVA7oUnO+zoUXW8i9o3DtO
tNR+DluQ13zYLJrJMXgmm5ntEQd9IOr211Xq1Fc+ocgdumEQCD5uCwAJ7TC2GWqsjXX3rEG6Efxk
SOH8jOGNO9YL7Qfft+3COIZUPv0h9LZjIBMimpwrpkwXpOl2Nw+0JplNE2Nnh5HLD4r6+v727+QW
9uSie7T8EeSf0V1EUMb2RSpzj16Zk8sMbyaaa+mjlPPTpSDAqVNxfVvpJenX5i2cDMDTq33wwYUw
gDGynQlNHglm6ZTkKVQENWoGG9AdIoSg27JeFmte5wRKSLLd6sMW8Czlx1vho7vMGLoU57wwaLcE
osL8zmkRaMwW3/NnUlK40XZogg4o69DhH5RGEi1cHkAzFggP1oMGhBE5uVdaRUqnwbVVhx44Jjih
u7W406he9AyNi5PnY7f2Its+yqRwIZhq/BPZxz+/AoZo+BmGVZKJyzikRJ/7n4OH3ZKSnkgF54li
QDEM4hriyHlKaFUrhtHD0uJcSoVezwudFZN7mRnxdZ1LZuRk7ErLTT7dDEtsE37QPS2vSEMzpYdY
BIglC9PFOwhpWQIInzXi8KzAKwom7NWKFqK4/m7QbPMqez9YEHU0LFMALgcvRzOKrsS5PEq9A0c4
nkkLWNAoWaS3glazbsL3TH3CjhymVPuupAmH82VOEhFOHtZJv4Tueumk7RIqek9l0R/hSAwR6GgQ
R4RI0if9TVna2RsEJXe7xkEW70trtFmFK+wdUV0T8hgQkos2glSz3JYNlHvaiKh6xysyiXk1/TnZ
jefiKV6YrRHJTawvLuAt9FrXt+azIBcLZfJsLr+ZcmoR1NWKbpW4UVaBcLOgah9UKVAfhlASx4iX
ILXgqmGN4jKSHCoqz8NE2dbfBk+luEp/YiZCLyrBganoOTlGbbAhU8++GTufQmtrfgW/7QcWegMZ
sjKrz4MZOt4i4HtJQxMIZAXgN+/Scvp0FUDu9yXMBLd1Y1FzYHsTj+g40Qeag93UShWgpRLxj7OT
1QJU/KwGzSzbIMHtPHHt8xYzaS2VeeT4RukNc5UDbthIXezD1GwSCuOU6kcKVtgMP74hE+9weSYt
xcLFjRGaA3KnQPIY9WxkrI+VXwt8iEHomtVnYXIZ6Tf95lV6ApQrVkk5Nc+NzdFrwGUaTmPomxet
1e7IqVJvYQT0sy8sSTSe1vp7mpiz2Gxg+vTuf/cyTbA4y8KvT2rFTlTSWWEUQgHPCJ9vL+a+mxik
OndXNz8rhw8Mti1R7d7MFDgzqmcSkP+WBIwvrAr6YRoSYqQl0X8h0N2tkIeu6QY2JW4rfbaOzbzT
oxMFIPUNjj7Ks0urbUq3ltdh2CoXrrkjqqVy5Ht/X/cmjUKgUG+HiSMJBKDBGfLuGeBiFkbm3Ufn
KKTplSG2wliTLxlP6KjIQFQ6zUXs012jsDnAc5t20v0HUrSY7vort9g4vfH6F9oQTh6NSBcPTQ2W
RuA2c4XI6BF6+3pqUi7/BwhtMjJ8hgr6Wf6ip40Wt/hc8a5eVfPHjO28HBYgrJ+dkEHBxLeSVjUf
nk7BwlTdARE5UZsHzaBiZBQAjcnH/bIGv4PeJtcZrFjeIRiacc+wKHzCMRPBii0fsgLWhHbfTa8G
8RvCylbiECj0jiLCMHcujmU7AUneOPPmNg2ia3siVTXhwmUErxO5CA+QQdQE237djNOXAnMJfIOf
8eV9XFxXX5A2nFracnXJtSPNiHx6ONNfkhgRT9DhjP8250dJch38W2mEr3u3m4vJJaEb98bOK3t7
Lz1tqJJaHAZeW96NH9800rqgT1p5hVE+l9jT5egU7HTPO1FGWdDIw6TqvqITMtszi+MHbbL27v4Z
WkBfpYTsqZSwYKTYY16Ao8FIdVAqmQlGlwSw2vFAjLa/nHfpB/Fk6UxZRMbPCVcSi2nr2QCLT58T
1tsJCDcZNsFeOn+CJaBXnjkylMSLPlkp70Gyz1HFoUT12LjflQx2vKPelJ3/yfyr/DrQDja3O8Cl
s/R7N3rH8FhbPrf+x7r6jmhnLv5cwWBd7q6kkmScNqWro9l/F9gKTCFAWam27xJ+TzH2bcX4xA+d
HiawPddxjtrbYXjWOXmEUYdSdlr5C1l9c2E/WJ7wfaoWCUqGLtgQ1p6cmAisxXhXZ+q+VcjDqSw3
dF+j05yI/fiXjfYQMhpjfw9xTEoJdZq46DPzAw2WJq6hYmyxIpFQ9advR8FPyRit/oVSf+bRkF9t
86iwG78H2bmbRhHdOFUConfo80LI6cCXw03nY2mALLO8ilLSfAGrA2ZIyOmDwEEN1hrpRFfrEE2Z
IvuTRGBZjvue0Yjtq3pOxZYWMSgyI8X2rPKWz0hsgXOBlYX5pAv45blAHVP5AcjbX/HNXIsGeGIt
V94ebdfn30GrfjiSXhqDLmrC2eq0be8y7J9RL66vJicXKfh/FwK88kBhZYInUYiyr9yBfaa1uk6E
4bm3mj4YHJ0Ot1WAgVi2u/lwb0RC5JIKtQpBioiguafRfvbPJ7ZObujV3w0x7KeeM3K+o04bNOqZ
zEcIdeVgsp0Hh9uz5wPCnMoXqJIi7orDsKm70sVr4ILNVKgDS/QkxeHVhutXvmP62HKl7v3vu4wc
P6PG/6FtnDtMG9ak+C+ppfxRNqiG7NVY2vhwwRKuThW7rphEKBD7nyPLclQaS990Ql2uKCNQgqFr
463uRUQA8PI/dSIFwkgOVvjp+Vl4KFa25fPMTeSq7KFAZ68TrX+oQC5Mc+KlCueGo/6QWlW2qwaq
GB/b97OZMHdYDUdf+WQ0GWhINkr0XaR2+6LTUt76KEXTqa1c2qbgzOckcndfxTG2ww/bN9I5MgEp
ckAsRVXDFgjHP4B/03TbbSNDx9kngEen8Nf57iIiY0fBw+cmoie147IuhsWotE9MPcgM0GwFTKYV
oBr4GS3GkFs8OqtQdxO/M9HVTM6cTHLRGMHgiqnxKphfh6LpKE1bBSYMWPUAyBLEMiwg01+yj3tB
ZueK3Wy0B+cAEJL3zV4Z+lS1+bqIaOSCJQ7HcEPrtw/ucVaDocUcW9Hzoj9gsUGPLK3/g2sIS22f
NJHm7TmpE0+h6KD97n8aiq7XZhooRw7TcTzOXOMBHZ65X/7g4jGC0SBM5UOf2CTTmGlpoCZ8nd0I
IHqb24FitvMi+EYHfSAIqxnzjS4kP56voKn2tVVrE6Jmjl5Sus5WybSzL6+FHLPYaa8vea+Zq+cJ
7mmXbte3exmOdFaayKHNUQa3VQD+f7Rl3QPTAWPnhUCWckBJeWTZiRevQ6fQkGl1IBsWFoqeBvO8
/38eTGKh6IXPqt5S7/QRamI3uN44LjKBQcVR932pDuQpyrtbN5yW1pfloWrznNYvtKV+kQU5jbgd
fDVy/DjnPtZ4VQra/pnp/NRA0QbYc2agP3gWQTTmCLyU7/l9wgOFWjPHWCj0qWTPbj1W7SGGJTSU
V0r0zKxR+g67xupLwvvg4B9TIBf45MYI3SbF9AYkrFA9mDCiaf7Re5MhxMVlVTTIEnQ0yciCp9O7
gDHzoO+0IM8AtYAc1cASAZbdfJtReLs8J87R+nYGi/4pgj2UoAzHsZR2JHYBYhE23B9jlGPd4S44
orWJFYK2kQCERiINIINHwLKGAQXGlua6bHhoYB43DGhwNcaWfijDtkhnLEh9PHRbf7mfvl0tbRRX
AXCO85vjdsVD/fyH1lxNzR7wsD+XbZ0QekTG+050KJebCnTg22DY6YCsn1P2dFblMK4JAFuQMwuT
tWd9OHLsNZ0suWPw6MZVF53QNWKebK8CIvXyWIN2USvbfV1UxT0SzVAXAl1m4Iw2QQPw+4qZQ335
OGjhw7f6zP1YC3CfUajVvQtbSoUfbi84b36o7jbzzu6cdEgHf/TqDNHmxJuLy5z3OBoGWBp0r4nt
rgmKkKrPmrSwebr0EqaZjoYRvKmrV2wTb87H0ueUKPpMu1cXohVjg1qRFbOAzGl5kH5On2UOPq9u
PrtJziqai1z7SmiOP60vJqsWrQwlE1CTu63Nf6dUEcxGKYPbhDw1H2IOoodxoktVUKKFlWab5z8B
TE7EOG08Sst4sT9MjTmD8K79lSDrSDQ+YyNlTZ/uYHWZCBesc7e2tceoPPiA5sgv9C7goKW+Z5h1
g7PZZqnbtCwEv15ak9bWjeKYjZdOQDZ+UPoN61KE0jkubTSckjsHSIux4zgRISxoCTndb2Nfs1sz
LyR3PEKu4WQOSXMdbWIqiwjqv170b4gWff6OnD7+LrlCADGZAdgyRKP8t3U3CcW0qRfSEyjyz8cF
LCintGrlSL6yk6GCQfFtLOW2wGdEiwJdPL3pAv/CvTWyaHK7XNvwkH+xRpoiC4ZWQ5at50SwMRZN
fjop8n8ieTraV65Tisk5Spj6nyR8LPpdC1CQqILg1LU0fHwwXANZpCk1HdN383n4fD0LKu1AjbIM
IwuTerKqAcj+Qr5LXX95PgwQq2q+EegtJ/kOH3CgmLRXsfAiVeaqfs6AeH6KaO70sWh3EFJFdFmj
XDlg4dsD5aFR7hsSF5FVpUfG837msqZ4O11QbQRVs3jhEQZTdGU2EDyE+bot4O+F98TN1orqN69D
MLtr1BtEeRPpQgYcjSZ0/FbRgfTyRb0a9gmhbaMWPDApf4SEMyQqCLnlWid0q7ckDycqT6LQxkB+
GSSUbl2+UnEegrngRmODVuMeLKTAfe8FfYqzLr6wqNTnLhkmFVdFaQfFHAP1Q4OG38n5yg2IZfHN
1a2XEwLSDbEKpYYLtHJH+i4vdKaIFcCX2D3UqGa08xpuV9FlS69jUg1eC/VDAwIUiSfeC1zoiGHH
vWjFazFpBfzgYAJwPUXsYJlzbtp14QHuhon8sM6vKUt990iq4eTb03ZMT2ZSEazXkV1xqBvaYhXY
SdwuvYWvw5J1g8rdvvTrK91F40KA1A9PMCOvX6YxINIYpuoZuRc8cTUwSnjBZlUMrg6j9R8n3LzW
3QmuOIOzScU0lcdlmsMapxeqZT+SaLHW7Q4/BvfeaI+MB9ajPq8E8mEvOWJwCwCB0QInlJsvD1G+
uyXgIYi+Fnuphcja5UR5vd04E78R/dzqvUcfdW02VEjOD7yGlsdkVdn+JnhX4ldVSwvo0+iGbkGt
+dKy6kdWiP3WizIvAGtRZBVKACCiztZpEjE1bqR05Twy3HldtcNBLXsPBhM8BURv+LnfW2sRWff/
RDE2dzh2pHYmcXnvWP5Mt+2zgEaXkaigJG5mQvN9+eql45Qs+2fNrUHf7VhBdKChPPs5UwGSfqwI
X5H/Sh2CVWbN1EyyI3mb/9BVAKkASMQZeDBmzS12C2KFsvuTgzQKAVbm93K1ReoYjW8eA+MCiU1l
Czuw54QgmXJnOjMpGxFviAyKySvpVsl5OvOHpZ9/jv/KE8GD58ACGjLzPF3bXDlW/ltc1PNP9wkq
5skvijNMJYhDkCYZxit7G8meF51Ef7Wto6FaPShWiiXKAo8mjdISIaGaCU16lSQpGAWc5CfGtLBC
0dx+9gtFPWCdWlVC13Lzpm82Z8N6FA39UGpn/R0sugEKplifnfE13sT9gLZaCf21LhBTLv7uU4cO
//W4BVGtX49W9SSf9CLR7toySTrkbgP2waBHUC+4UtfizrgcOAZ6Ate0IR9t2Rl+7q3ZhXrU6eIO
xDT+rTG99Uwx7TMakWdRhDc9lr+JaiF8gQpjn56tczXi8mPM/mlrqDMz8IuWLGVS4zCzrZ/PyrVE
pkz6dXBekjGut8+MWJ1mAEAuwV4JeoF1/6atPd213cGgr2qnX7k53v5/DEP7Z/6dUFT3shmRWPaA
CFgWkNuia+Ja2WfcOrBqU6YwAkHKQQ7k3gyfQbT/WdcPc4s8MrD9bxwHvuqXkiI/cMHUMKciESDu
uCrFD5NS9TXXwnb0UAZXL0cSkZh6HbjEQVh5fPES/j9g17kHCQYC8TSrU+d0h6uc+K0hJtafaoIU
kpiOJ2buiUgYODc1yPyvPrM3/AGN+w+eUdbaNFNZHokn9N6TU0vZ7ziwjZa3jeCtwifzUAtJ/Qt4
OaUFT60s/BMV9vyqVWrrL0fr1WeuiKozN6laGR852wPC8tz/dSFOp9wNNn0AiJZ7+/DjSnchpxF3
UvO5YdSIQLIvJOg67iubLxnkSd1h3DDe0fph68mfBLIP+3PJdc1pBMUBH9vfpCq1rChhTZL2Mw/6
3CnG6rwPCVpdiYSX5fG7y8uJVthv2nLLauvAFaBFeVFSyzYy7isuRCc9RanpEmm5G+bsn/mSRzOL
wByrl7XCHt/JYxQC+QI5UwMhhSUYcqSzE/h7Drl9Rl05IfMZWUIp8HYngVY/H28424wNH53Rtbtq
YC/DlHmyhDPbU0JfRxwynbn4jdBhpBxmEf1R1meWnJ2bHc6uMoMDsbdKbze4HIGav6twaU+freTy
cPH0wVdk+8Mz5P0lDcwOkCB3GKsamrse54/gv4gHL2EShRoS2PhxuF/XARVT8ZDouZF7Js62fgo+
ujwwvivUl2FKKgeBbo5TR+0wqoOrZJgj75fShN392UdM21jTHWWKCKxziBscratMvshVMRuDqShX
awsltNQq/TR0UVTxpyfxDJI1ennTfYcVjJ+eaOXiwLLp6QwtZsQAFOXd3WcTuuW4sK/7doO7zmzS
cT2xg3Cx0PE3mN0Ia9MSVvySDsvWy3n2zEIclHhzgTylwL5eIncyVDwSdpmogA3XmSf9Gi9jHd+H
EWkicu00Pe7tPhOH89se0sISQzOUlPgEDXLu9ZXAwcPtWN9DNKRNV//kF/pKebZdwH3r8rFf5y/S
zIu3mUHcqRzSjazhd9fyTl5112uCFbv0v3LY0nvP3F2xICH709k/ojldcwjyQbbB7P7Z9DRM3kVB
n+t7CzO9SEnsHQlHoux0J29MWKzSuEEFvh4xMdlMTo8qVntvxpfKCAL+wNW3KSf1jJZ+Xs4ntWUa
WJOiQnyO9rllnXN7j/je5CtibRnH7w6CDFuN3ORTdGaU7aQN8wt6rqUwydUH3YdE3eaeLk274inB
I2fJsdAWlGUkzZRwbyDJ9Sv4SMk86QYCIKKmWoUw4KZSMtJIJQQLqew5EQr/JFwy2IqWxWUFYjpM
5nd+kPMQVXjmsd5l0R1v5ZBdK2JXR1DeY+bgwYp4ecCs0doIOjZI/ik4EgZaNdDfLWTd6LZAYUb4
gLKOcRddDhPMka7tcEpeO8/wpSXaD9XaksRwHTHzOkJRHkQT0tdYuUK7b1LcDtZoKmgFFvMr3kZa
edCEc2db8jjEemoElyLHt09SEVXPunaabbv6pG5mksZ8zrNbfFUacPpbRw8ixUGmhdpK+tD5AF4x
YgzOse1RazSStcNj+19UQnc/D4IE5wYUm0LvafqJRceyfUX7yVvgEa4CtGpz+k/GGugMdobjI/zk
MwAjj6Ym1a8ej3A/qkuMbVP47PHG/hCDHgQfQHvPz5oIw3Huq7BhydDtyt+2OYfK8P248hKYzOai
MWOyQu2PPYP3bbkvNXqdzODm4VoSsfE9NFi3juSbnU85Oze5EzO0HhcevwkhIDGaDsWAstLlhdoX
akHPpNdY4640xoH4L/aOiC2sTU3NQk4FQsnqzEuNhlMKmPTPMBhkqQOyDPEZ8cfDLEkkYMe4ZYKH
bInBeyc0W6FK85GEdDXx/oVYdsxSef2ljTJW7doS2Wt0Z1sb6KrNI4L5uaBuh6ykaTi34oWj6880
syt4jltR9tstSxGJ5Yu46m0Ah5SUdQNKcyo3oQq18F9vytSHFz+Iq2iixEeA04MvJ2ZRS/LKjcbD
mxaAgoZC3uLuxTudgYyJAn7i/sA8fSLTqzwNpyhp5O2LZgbTZyBBsTnGY/KGaDeJG6WSxdpCDdt0
R6y37EwhDkP9+nSLqxL0yDE+0fzwfJIDkrQv8kJnbD8DYXpR6hVS/s0jsXeP36hptdHtoR19+Jdm
dBa9g0hidmhUidER3hL/iAgJt1IeWe8LGDWeWTVBre+6dMhim8hfwAwBw9QA8RAcKGAgmp+2p67/
bS0IctrIyoQ43bRD1yVIobHB2N0b7D8dhCXlsEhplCmZHVnD0VaZBcnxZ0X+uZjqtoOXVjlDPeqb
83CnDe6rZOVTnfVydLIVX9sZYk0GUNPYbj+uAeT4euZlNxOrOpFGadt9SCV1pTtHNsMJlRyO3OMl
qhIpHCitFBFFh76nyUAiLuzsnvnz2T9Twa1uqY2Lpc4VUIzsT1KCaox2MIqgK6QQ0VNVDL6uUZRY
lTLpiSGb1NgCUsBnDtAWNK0wcB1TOyZ/m7Ror1kjfngKP9GIF02GJNRWoPHZJB+8GzyhVYz5L+WK
mYt9oyqh2Qf0jx70ovqVqx01CSRmoHZl7dg386TRZ5s9LHW/qYKwufhdNoSYOAsMIpVojTe1ciWX
7HZDfj0aYphO2DtVs/UgRsBjiB5NowBf9V3jis4kBPOV+IS0EbHieXgeH3NqGNXn51829ORWYeLV
2uG9RYtZmunOF74IpTHxNFdw23va4MtZV8h1371MuLRZWN3b+JbDBH+Srb/aQHfmIjQxOfx4G2iP
pZu3wZXPbE05bXna5RQ/N3SnUIERYsScZohRP5yQ/uz8jgSMlyljWUDpH/0AS3FmlHuwpXlB+SZ+
pBz02buHapno4kp2oBCACKJ3CaJLv91pxrzPSIVVw6k5lP9IuWD0QX7tRAG9Tr7LUUJczZihG/lf
hwF0F8B/+rTy1FDDZdBawXqMAkOgGTM3SEJY96gcwQeg0ECbUORg0Q4IlQR/39R8DuSPpseVy8Y7
3vQHs3wPfhKeh/tg9YW7VL1Pkgy23bDTeOezplp57WihrwSG9mTWHegxWL6uyNgO4zNopGYKhddY
uQjt7lqaOoyM1KbmgEF9dBDy0aiyzeGkNWCKEALf4pFE5obHdonmN6l4WrtAuNlHnFGM7jTh2w0T
xF+jIoCniq0d28nNBggIbn7OUJj8LLx8EaHCQ+cFPhIediwTwSmFAquqKvmSpd5HvltIfLLRqV3+
qIPanhRJNK/iuRBbaVsPg6uWn8rJrj1tsf42neiYZS63AZnjH3QPcWBIaT9zrnrW4Pk4pqIHoWda
SM4k1DcGh9+Lvjn+Q9OvfoVvW4ic47XTcpAQACgoz+vDu/wijablLueqTchaAAJp03Qd8stnwFDX
gIdWEjjoB1yUUaZpEZsqhVcdPl2FhSF5eeH3oRGUfZK6k2BUXXy1JAitY7quF4IXtP1w3micJxD6
QsKzM1jum7sYjBQw1hqe3TYZALxYyXBYKUHGsd14fcbWL0puXuDOFJs67tJEXWGwETpCvoB1fvLn
hiPc+RQfdx2oTOI6xiEjuxNF38udFsMUPPWZlpY1KeW2Ntl+/91ijZeU58GuyxXUDh6FmS2nWCAd
bDB6JcxFEw8yiWpjStSto+UqoPgBdo6xut8/MlxhAuxs1cQF4DrXJk+I/hmipa/l6cKGxywVkhab
HtAlemf0mdaXZQKIUK1r0vjtS8a+yLqUlR5dqxjs087ljRRvkpv9lK3T1DO6z4XJbdGXNWMdRh54
CSym188kF+nu1mJLS01+qZXCX6V4FKn/ATBcwo6ziHQbWYTSCgu2sv9jYLOG2pv83gAPlB+lynmO
bec72w4szn2xBeU20V4EtTTyTiPfBLxuBZhiosSSZHj1g0q79yzCYkiHjxOP8c/+AKsmj7UBoXqq
67UPOHbk3PHygDaKYXjHLQE2JSRyxII47unKGvCfMAbGmXsN9k7rHY8VPyDieHcpr/sZ4CVDMaGz
0zf+Aalb5nSeVM6a/UTjYp7SnESrAcWRIyUqqc3FUjuy6xp2F62wfWZXz7uPAPNBVZ8D7zI8nxJF
ImDxfGqefbbZ4Jufnf0VbBnbYCZGujaKatOeub3sxMbOHJBu8chba22LGAgF70ghPQ0q8Kq0DOMC
L48Ns9noD0vZiaqkmnchlUKm114iT3/wCTYQ/U8iBs0YWx1MKXvUpo3Rw4c1Btj6TX+jeUt53VWd
9wYTruk3CNd8qrZOumg3j/9RaBLDa5Cv8cK7nOpABaBpoT1oMOGBxuRlXJo4wxMnnviSpZaDGJWn
mS2Yh4iKxXF2vFoZHPXIyMaSjpwceWJLlpnYNii8yPSeC6QRUCOHvbjaamEADjlWD2HWA0TSZkhK
qDaQCdf5E4xUte4/ErP7xxwGtlka/4C0be/CavzxhZswgTTVm0F+F6Fzb30X7AlrrT8pGQfiETnc
99uV0UpFOEg08nyUfcud2h8Jcq5/gKexefTvDz9gZ8zTVQ5+QlBKr9/dy22F/Ph6mPOcv65U+r6m
gELTtX3xiBlmVpoEzWvg2J1Eb5+6HXNrsOW5O4TnQVJ7zZsh4OXdWPqtwtWGTjoeaxDj2YAsxIUs
o/COHBoal0Lk8bOaqcynZKegpvOhn8UURlkKsaKPFKLwWhKCSTP+RlzEldyqY3NAaLPFU3cmhPDa
yvCAoNvgdLdq4cEsWpSCZsRNVKmnwdD83AZhZzmFcxyjqbEpn4HslYUb6DRmOse00y8TWS0tDgFr
MBxq/bHKVvLyuoFXv2KBPXiuvt4TXnKnav0Ysz0SDHzuc3mo7fXj3NUW3SQcL+hLDkd307CK6EO+
lzzyJxatb64pSXZOdP3X29qd6Y+MeJppe8U5nil2milevI5fY0dqu70lWr3BH3Df6QNjshT8aZyR
lHJRCJ7810BdPYB2L72jz0DY8L0MIch3NHCWyBee7Zm0jIVeBs9GVWGS4+So1sR1hQK3cb9SvASJ
yCM8dwUmFkgKCOk8rxDQBlXtLOa+pRla72QvLCWDGDNgRS9WF1HSTFIssUOEk0ardUwtgU36NUOG
SFaVosRgXX3+0QAhuVyALHaBwvk10LlBNf9blGBs95yp7TTK5ii8qRqsdN+kMj1c2j8RLKrDxp8e
qQJ4BAyGyrq4j+chy08ycUeo9f/VITtpMGo13Z8rXnmVE9KLaKqsbu7dze0mtpJ1Kr5QmbMVEy4o
EsUkHRaASaQdRRSqgua+0N4VrUksJG7Gu9b6RBuKf+vNGGk5DpFHcT9TXUhh1Jw+zdehY6t5Jhc8
dE8dh8PSfK0j4bg1a4xO5OnI7bB7xU2x9DTbuGCqzrxpd0XonZMSS7DQNjU1wYn6Epwuw5M9nOAm
E11zeaDg4/AEie4KeXGDc99WShMogaw2M7wo0Rg6GQicyqtHNs/BJrOrQQ6r4FKxTIDdJ5V3ow9t
glc8PCOBYjYub37zLcgDqPZogYSvkJHFa6wkgJas6HjIx/j1g80I/VmNh7zMZSQB5XqujHA1mVYx
V1PyCl5CiV85bUf27Rf7eb/BAhAutO5f70Ov31/vOdAmUMGNZI7gU6sESmKSmmWiWIRodZPO4iPS
TCoIGqpONvrQzCiBroNklYl0VrTrqsOFospq4Omv2fUktfJQNKpCHrl12oPQzFs0B5ZecBpa6ckZ
wlfJIIhzZhVrfe/HOU2GWXt/mAokvP7h+U69cxSjRz7hLW4wGimBgzuWct8N5i5UsKP+2tDj3CDt
tWFSap4zydI2PNbIlAZtLztoESSh8koNH3ZleYciXuOiLq/oPvgxmDaZQwUrSUgxxOr/QmJnl4jl
dD0Nx2uT0EKurVkkQLK0KFUGfNdSFlYvwrKI0vyfKphtGeULJYOoE8QPF81NotY0X8xToPgRY3Uh
wnkXzJ6HNtu5L9cJLm2a5WPzoCdJ+N5+4Qh+OIZ4uK62zfSvTVsCJHjoYe0RfFDt+rhcStaqueT8
yNx0MTOFMfe0lvLXjzjTzb/mDlKmQjWAQ7ddja/nhUu/CPcqGmILHU+osKvVjK1wE1qzp7gjHlpX
nYfDyhr2Q2861FXokoK4bbOpjMADFzto0cTBc1ToQwjVHJNDHW3GW+mSYRJqulECALkdBItfNpiZ
IzqUFfpqVbb2wgzXjdpyctikTiOF1dhLs7+gK7xGnaaltICya4BxPvFEtrWOT1v/wS6b4l3R/v8f
Z7xR6c4NUP7TK1IR49SfaGm2zjYPFSvKow2GIYn8ZoFot+HrsfAigXda8CMQzJERyzWoVNDghi6I
PIEVcWlz40CDOpJ7nt1BhENQamWvA00KYw5XQ0KFa2w2UHDpzSheFsORxv1/ktN7YJkIC/cXrvAm
WKhkXlLl4B0A5v3180J11kpDf8THk1ZNHgxQb1Y0w758MecvFNnkQKX94cqmBEW8TT6j1/z+Yaqc
mo48jjRfH12apXDPM6wsa48Xva5Gxp8SMMHIamVWJHN5jjMEkY3hVijqx56YscUhDs+r6GMGA001
11stPzkQuwVIiP3aHdLfgQSNVkP09Sip4MYy1VX9mUm/xB8RTpi/iujZuJdflzcWO7SR2Tr2toNl
T+WzDSPILhe6z53e/EhiqVuUb0R3oM3aj9crPvR01hTaW5wuwhu7IeoUFNlogxPsBEGUQEJK2SDJ
OUATysi/uTaZJHXZ17WCjZbaNqfM/v9K/gy6MlFisE4CtlmDFj3DoDgi2ps3OrrhFyAUM4HFfdNy
1UkQMs8yBXToxLLEo2YyFR9VQrfHhIP2p+v4XgtCczSb40n8SqSGjVIEes6pBPxbdJo3qYeu9z+j
pB8wiMdQ5irZ+rY8MkYruVNS3yAI1eBrr8EZY8eA9+mSKh6EVYwZJbInOAeXXFo1N7lyYpXc3d8m
tO7ImZHZeFeadzturRU+rX0WdoZQALNrWcxouF9DMW2GKTAFSg9WfLlCmp4v2J2H0BkyhnzNEi5S
HrZ2bhEJorvkCDxqR2enLw0gTDiouJx7Ty2cgGFDIf7mF1dIwt7EMO8SFW4yBCUOA//0vPzJuCLy
JJsvEe6al/6gvBJ3rcTSEaxawUiaAIItQ70ByUH4Zg9UK1skpOABTGskK8jbVt+1ruPits5YNOEb
+DYYnai91Q7LYp9IWCagjESPyWJckiTiyRx4hTHZIej0MILR3wvV0yzipGC09O2xzV+PU9bxV7YI
r7SpMteV/8az7sINHqcTBEeLFpIyMGWkVST1VvmhX6Jkj6KFxxH8AuHOKzH5pz5cICUwHGjBrgRQ
YbdiA4oDcJcek9ZSZbBhY18JO0YkQw2dN+mTb+j1NsdfwlUknlwJNlEkwo8h2pFqxT0Y+ge8D6Jg
kP877Kex4s/2cAnJZnuHknmMEnBb0Cfs6dWkF1Vn+6keTWZyiv3tjQEADblT7VlkPe3bATz4BG8g
Gt9b85VyGQZOvcOiTE1n7jT4EsNZDFTOnr5FmXGQ64xry4+PpWdbO5rcANmyjbtmfD8O5tWPilDv
wmoiQAUF0zAWKDXgFtxQb3Eap74ATUQnbSu0F1K08VJXibVN/n3xN1N1fVdz6d4W5CIWTNZn2wuy
sa9wRd9sKhraTM5oDRleghZlRk5tyvGegiaAl5qnwQbAHAFFsllsPaq4OeU50PEaudOnA/G8xfZU
Y1Kwkx6iZEEExAUkadzTIIf562yay3C90/AGz8WnNubwT7gxDy3LDUtkQQsa43fXaVKy2rR1Vl58
zp0n3S/9oqKRSm8NgSL1xlgLrbNnft7pc+LaJ9toW2dgUNdzHWhqeziLG9LsZnTt48CSB4xisb0D
wIAjEqkMIWC5CDTF6fdEkEiRi5MbVRsn+zln3SU5pyspS1ku/KhYoDr4ZMtWAbHTw+0tTBXNdJmY
b0A8GQrtk0lsI2Rw85WsL/xipX1/O3wxmIlk5lIJfS6EYeS1vSoXCe941YIU73RKBX0hZ+J/c6oA
/csYUUtuPH9cJf2CC2hSPn/vgeL8hVxkvj1G6lqyqa+HQOvZjCKRDLEIc53F1BVBTsoDV/BrFhZH
udYTv+720HIceuF7UvkyJJsB6DN9mco07xo3mP6wdMI8czHscTvUmyO4xPMMGNn9LIFx3HLBtXlw
LITdq0CWy7SMcLQGvHiFT7mQJhQBZSX82RLUsev27eHK8q8+Am/vywhxx6PtT0S/eOOTP7IfQXAl
XGtlubPluRyFdppuBPGAVcAgKKELky/HQN92wJ8L6RhuummyD+yMYGLtTz5ZqTuIkJvMhElGjEuL
E/gCdq8LONnHKWDEZtmMkd3Y8BlMUpiPqk24UPEbHp3XCxg2cDoBM+KLAmD6NRGp+A986BQPiqKI
6rV8LncMW0nLmtxHMyuc3o+tjhOfT6US0m/5rtTZD3iwg7SOz+215gX9WWhJXZdra0nac8xRN1+0
yAz1iuFd2VuGPK3JtBcoqZdRXYdKMvoamkAopmhTZ3dahneJ6r75OhkzJvOjrGZwltbsZDmWHZEb
TDMiOXs0oZdCDLqh+6uQ2v9ySurvsrjWggKhCSbWBnoXGajo6UdlSxF8v+MVorlEtTBBduzuVOWU
vb9cgAtRAsMQTb24fTM8fcqrIaS/BUEkVkbIwrjWG6FUMAnPy67AbD+WWQzSsoZHDDzYgSrwRnak
tYXmqUy+WpRQn+qTGTZ+sCoRJPzf//UTUu7ZgjDYlh+NgxPD1dKkZ7AglPjhschBcOFUFtTudxl4
sHd+/I1cVFE/9gLyx1SPgR4bHpSZHIzpyEd77YGDeO+BGSKxswhIwZgzNrHpR+HUejieMLcmj1TP
jthe4SDtmvN1w7Xbp4RRmcuqpa2lL9654I+8x3IFN9ajWjPvIdPEHgYp6+0umiFHS3nLhGrMyan5
3K9F50ktFSXd+zMk+APvWb+uVde3d6ZR41WcKvpVY+QhoWpG8yOt6aN2jbLqCb5n57DKyq2f/4FX
lKx3MFQVDxAKBWKa/1exkxVJmO6Q/UNsNWO9Ihf9Pv1U3NXA+x9S3bKfRI/c/QsAhwE+G+XapIwE
krVeKqWa4v/fLfyv+Z1mRuXcJzEroqWMQxtmrF0TC01K95Hxb3Gw1ldrs9Sd6Z4uRmOi0qcVRccN
DKAf9cFqxxtE0q5xJQ/A9yEEOnpMlwOat7cBPH/VQhTtjAWKqoE4TsFx5SIaFXIqTwPYUcG50cX7
m2eA9ru27efIyAsVZyqWtmfO+PFaDd2FWnIZBve57Ss2vPlREGFPqu0izJsTH6ry1b8PDvqvJYCJ
79ssf6aqqGRRP5bQH/CnRwrTslUG9U3Dkrn20YYwN1gLOaQzIEwkwLX7dlGowJ10wVqbAr/1Bqn0
9vRx4cfmZwI1lRwTNfBU8eFME3qk1W3jC89J5De2TimnCuScFVHUbElrjNEn9B3Ux3t4A/u3wfQx
L1mOGCBryefHjkqUx4wl1KRvtIOZoSwgrJuybYb8w9YuzppEJ818wOy6/mFcbA7zOd0c/oAiP5Se
FdGMCE9MgsAKrQujy6/i8eFGLfVutTkuWH5EK8tm/QfJq8lnAYO1zAxp1Azt4Z6DFyP5ZstSGE7y
W36A+Rd+eXOwH84vmWrw52QffljanxScQ0j4e5nnkuJAXEIH85y/XPoFmxNjxM9X0KpqR9hLNZle
KFRt0bhXltM8g2TtskW4qFN6xLBGibCT3bfIAptZVRfM5bFypOCaMOB42DvarXuCYrwVyeLkowQx
OifM1CeDh9rs3AMtFWLw7ZgzsN8Jt6KSGrsEVvuXMhdQTUj4aB1sULHOzlbDMvzOyHlXwlOuLXEp
2FOaNY7HxJApsq1sR3ntKwhOmHqOMW/F9o8Ck3LPAeJjMCJYMuPSLb689Zi/UXraXBQKJBsDyVyn
gq3bAPAxyEDiI37vMuB5yPwoynSRb62bnmknyiQ6jydjAcr8Zi/RWY+J0rcD+fSSl0zsOEg+GUbD
WbbhNygxO4Z9G0P7xHonSrZPD4GCFiJoY1M+p6UjlPWMMk6vEdfXz+37yNssx3e0X5ksgvPoDHGV
xl3ck9t1zQrz7O1tvgj9Fpu/hAyJl/+eyXEGrZ4mrmnytS76Ra2YgXB6iyx+I6VaksHp4lnHpoX6
K8n7B+QF9+QmV9CGzJWNQVAIFn24V2wRyeDp0osIv8fIFBQanAFMSgVL3c5VvL+6bHqvK1VCgOyV
V56VIz5XLjFfUwiJ7G7f9GtSEsoKyLs3w+LrBuQOafAkXhPB8aGth60cS+DUx3B0wmGGB1vmQY7n
GTF1vPxN6hAn6HOqn1UIkFCRxgiuVbPcGV6LtAAzRCM/XRHglahBIdd1/g2ukBUqEggsmvlewunM
4/32JFX8iJ2R87KW6L5+LgQdnrtPdhHka7DodwbdHxHiJcy5cMHrnLchRkmO/8lwB2WukIQxlZ/1
4TxwZSm8qiGAka3nwJqX5r3oSgMiw3F/gCRZwIbc+qkCzDrc1QuMnu9mkKdGfoYlPSA/4E4iAeQr
vu3VjIcL0JIGJQX4bArhN7a2Da5Saf0ojgGwkBFk9PlQJr4Rw0aARmqKhV3Lfmm587NFscuRgVrm
Z7BjrIrYes/OIKofm3KxOfBuTLRRIJZeIssw2vF16+YhUTcjYRFA2n2BtlOnYo4B5LemaMGJLLzC
MPq3UxyK9sa/u/mNbSIaT6YtHF9skFhYAsFRHaWEMlgJmo031w3FpDtwGDi3FZeAVPPI4qoUPw7c
NoU1NQtpNI8aXwqvBixnLs1TOauON1S3oIIHpW5YEEUdek8DSBlLs3sy5PUoKD/WFD0JZupNZY5f
pNuLUq12LV76K2dctwpW+N8DyZzFGavsy0iGqqLjkrhC7R4fI+YP4VHwplYj7vGBrtRWuq2R+d/E
fXNQaaeMY0v6UL/WFQn89/CRdNWg4cXd5D5mbCLTILfgy35QLaoXzJLn4zXqPHfXEVgvOzZ/Igs3
tI6ph2o8+Leo1a0DA7DJ4K9xAw75anjA8NCFj8Q2WyzsRYhuj8ra3EN/lykeG4LJR3V7gmuBCzXr
6KlD8m/A9wGxvFqhQVHiVJgbphnPWqSpdzYRN2bDdzEK3jU2fqsabvdHmHoWUvdiT86wNvCbbWBh
lvEB9SWAc4+k2BUDlCVoV8qjEMazqSokT6m0Ct84TxP2Glq6G+xd5vXcxCdV1QoclCD4LUr4dTw6
1h0lGFO8ky2vKkyetlHbGFoqmQNsm9dbNRI8vdFRL0WJVOh/E1N0NxqIBLFCTWWUbrJ75sPdAPV5
ewp28MyFg+Qppb2J90ik/oxA1Mk6/sIP7wzhaGzKI7elUK0To+O7Gym+u2LGyA1+TrnfcGQ++fNR
Dcl/DX0g3h+NbpXiyW8BvEM+Grc/3r7VDRb1BBwJ3rbfIJyOaxJvRDtH3dprtH+KYmwWdAg8Tci8
OUJPBvqlQJ4O81PcvAiDfy2172msuDLKS1cuv37FhaFgO8YpIEvB2ZAqawbvPfI/WrFe9zLF5ekj
QMq7OGILhYRDXUurJ6u6tsZPKuurGmFns9mxLZPD4rowOXqy9qC1qkvjSRxRFk1sSEf4GX4rwKd1
VTN0Bg3aWPFr5dE0TrtRpAcDAdQ3RLM9e/EOh7v4DELGrzAVBW0qIbwuSSZQQix+8ez8rK/cRzSB
4y6IlVJ7zpRIRRpNUEyvfi9Rdrnz0MseVUsF0K/d4YejkoIYjJGpKUuUL7oGY8l+RNl8WdkZE0gn
iyR73wKBivKJLFpdtUVVzaxoxVygMV+Qa/IwEhU3ps7qMNcg3IbrDPhdFJzwxtkL7oPQrmp92iNZ
xaUhuRDyfq9errDjPG4lLlA0sGMpCuQABXkzV3QGrQiFCHtKSlvbJCxqSrd2RpGjkhmW8J8m+8CF
Spxd10raoFYR82sxxEJZUSS/3V+SxBL9xBQ9oWEqS7Zjak2KRDEiwzIByX6RRx9q8O/pye/02zLP
YnPY+45uMWObnWXgcSJOU2jcq812hLi9pRKu5PnslOyj6ytXzn34znrI1mhAV3cILX6DtgUAkUx+
C/SH/3W1ZU/nUyb2zbJKBeX2lkyxC6BEtrrb1GH5SnBKWUqfhqblMTFUu1u5mpElpJkzhds9xM/X
w6QDeBlviYpBNTu2OTxYaoWgxp8jVOzPAHpgI0dlTNYucIPHQJh3zi7NfHTqKlQGGSEjZhyJ56Tq
NzMtDHEfHo0DTkPojggD9vUv7qqFAXTiZPr7BS8AiSCN8dP/dbVZkzmvr1c91oz+ubhodlgfwo/Z
zGyhemBMaU97LYKjkijjwcdLjdpRLGkmVLGZLB34HGGs0kjAVSrNLLEe6RUAF2Ay7rw7CbPLeyCB
l3ThqPUd6iJAuypav5ADBGFA7NDP1c6RkJTwCnLdpTIpgZmkw78q81SOs1mK8zAjk1HOUUm8IsYj
+R0KPcftUNJCI9EtExRuh4mJOqRSabSUMxv613mcW7VlW45Yw0X18FweHQYJnG7BkHoe9ClOuuHP
RGq9ZaF9HoLQqgpwxmKgm8HaI3MwVXuye/84vWLRz2gTP9sF+QmycqFyyLR8MN+GPORqMEmjLnmo
R/RIi8fVZ4xE0GL3VdtpKm7LY5in/EKLdo4VV+rK3lpv2s5jLyogaAB1Py9/NSF8AdQCkYSveM05
78JZs3O2NXxGpyIeuOYXMcX14/eILzcYEk0AoqVL2DP0Y/HyJjeEGHNMwKlRCXHaW7h63YTXKck/
/UpOU+w2WE0i/+mVVygKfYT8aW7DOxnljCoZMm6qKMc0BuQCt0WzZIkftKv6ewu6P+v6gle1zFkj
WLmaO43a56pJNybXprpUM9Evr+gx9EFtegU+7fsVnawzND/qQElIQKsvq2XVYxgfMnD9ka7Bgg3L
4VwDgi6ThmViUFFzsl1YwUZelQdi9+7kYpZn9E6/iurz/wwQQ2+2haphsRdIa+Kuh1GkWU7B574c
2aNxLmuOg4bh0y1+hSXdVk8S2vHcOHvnvRwFnh+pwDiMtrEUrnf21iRFttFiunBO+xtEf73jaYyl
NK/D7sy8YZ6yK41KoB//gSmvejNvp4Wi/juI1ZQsYo4Fp26oUb1ELLw7DD3O7ABYd66PL7g+VZEH
bzlPcJL3/tuFuwEPBa11ovTh6BwzOdTk5b6VRkA+y1j3crLdcP3JCs4UrPwykaxDm7UQTKy0yyoZ
4Dx9S4L/UdKGMXtBTEU17Xws0lxBP82FuVAheJK3UYXKt0PnPam3a1lYomvhbGd6JeQdZh+RIL2b
vxkxE+zvHfauOKe41/HXfJNGU6MjDPBG6rrOyMaOs3ZXxvH7SCmdnn9L88yRU7NnrYd17oDfsaJV
HDr1GNMO0oI/2BiYip+DvlGp/mdXyZPMmPE/XiilTEHVTF7638NKOgMCGzb49bsZp8f7bMsjzD89
wd+BBD3VnIFnGI2NFP6nn6FFdE2Cr+tu1qY3+isE5F9J5BtZQfav8k9nYULDIOepJclSNTbT8N4B
O4Ts00AkNz45hZaBRurt+NjVWQLHBnMF8orQ8xQ4TYNUPEfLcYmt3hLPFwZbsuOQRZh5HANaFrmE
ENnl0CR+/+oF3bAjiTgKeZeUj0+8UKEsLldJ5NcdcbDRpA57eKfc3/DC8r2hOFAbwouIxoU5ltFG
T4ehcMYit0RadlnSVBgpR9BsauJu58PA+j84ASRbnO+nCPhg4uUyzyuLh2erMCXrP76jhuLc4j6x
D98Vuc7DoNN7qjNueBF+HPm3DXAHvAqHkzng9OxcpgzcRgKrZD6aaYjvH1nE3mCX+mElfwgLML1v
o2DzA4Op5rAOQ6qDLLZaGu1u1BZJGdagjR5MpNBWUe0IF5Ar6lIKRQsfqmyBHZwCkA3DWdjwF03h
g0c8OSMUC1FwrOtjOYsPv8LLF4nEtXG3VXBIMWoPWUZFTupL2dUafwKr1jlDM+KmYvZq9c0Bl9p+
CCOWWSZwHOGH1Y+0yBFuDlSL8fQPEeia8QPOd6JHkDxkwKDQlk7RN6aPADEDpV2KMIy5NJQH90yh
gUTtIQqGAUYHUKDAKIs4bmV84IRy93aNoP3Ut7iu5U+AgmhHoMZiXV8DqTe3C4tOwuLDVGFDnddJ
wyleRtKuq4zCudUbv6tA4jlsPdhrrQZAilTEafTD6x2KA31BeMoXT6R0VDtANnNUdbuh0UOddLfz
af+D9fiA14Ul58WEK4/ZLjlOpa64qSiYL4joOVHEvbsFjTxoDpvyDP7LPu3ytu7he1j7TSzqB6h4
lcNlkHHgsW3wscJ68S0OY5jt5YNaTZ7OdDmlMi36NlZHBgUxG5+TmoA68+U/P26hhsqokqd8nDwl
Bo/n6kNypwQt6yfHoSrxsNNAg5Mcs7T0zKVRYpq9XnfJniTqPWi6uH0ksREwumro+AvIPk6wYAEp
fjvDqiUQQ9yAxLXpQLfQbTBS/lRG9D5ZqNzYHqEw8VFh4+N5kZHSDWcCr51qIvYE1h4Puqd0T2Je
q0gRbuyf75hgDd1pPdsDbusnua6M5lyymwluv+CGPJZfuw/vUgRZDf+w/M/ilH4fpzXfZqUPitV0
9KaHj2tvqaCD7c9BozK0Kvl7f5wyLOu/3zXJGvWe9tzQteJ4Z0Gmh5+7T1adsirl5YOlNVySiw8k
W5Rlk3JhJxJRpu2doGbrxxgBDCax+1N4+/z+0zFoJWeLEkATRzxp68rMTH6qU8FcKi00J8hPh0tT
C0hkSA/DaxWg0sJAJaQN9xbGAhCjVhbsB67mRpGH4GFfwI7NibiQ6RBEJ8XkDFa1crW7fRNEdoek
AtXY/jo7RkajoMDoK7761FmYKAjbJftZMoG/cli+nRqSPHumy4n3swUcpdI699/jGHi94ntaFwna
gLJViqQEr/mOL4xI7d1hDNBXHveM+Y/mZ3assZo/IkhoacHobtPZ/I2BBXSD3EsMtxRCudpLALZC
Ap7VtLTPa/l6aE2trlIjPSDt3gQ4LPUFoCNXyejHM0b8+EjYwLHAvuFanwS+uf2eerLx61uOp3pB
ioz5PcgvMuoXH4anlEzuKZcT9XtGfe3q9NM1u9efSN3ONnAbfL7TET1iWU+3QAuAs4HLwvoEwyas
T5wF6lpRNtsiUHzoTlBgbtWaHVNv8t/BodRqBM5+C8dSKecBv4L9PZaBNkq8k8VH85sJL/2fxuUb
98QSGpvJ5X9l8p5shbNWeuEs4s2jcjCzb9k/Ae+7u4EFh8l0yiYzlMj/A+jEClOWCgCizrV/Zkkm
EpsRIvWLS+Xe8tJoZugfBFVSjM68gkvDbxjQ3LzH6vtbnJzk0NsxsR3HIUDlvtmUZhOf7qXKW1Ad
J3lxl2eBwA4ofCHOyH+PmFNKGDD8qGbvhKVYv4zUeNrO53lY26dtD2RkEa+W7hhU4+px7rZv5Av1
1oY0UpEBFxuP5iYtKs70P+MEHif5fZVAQBlGHIg1OQ2WCKVFdtmWDDOmYD1SrIvbwsM2ZAgu8OvO
e8JX/aJHjjhJAifrQjtYNMJo/MtMXH7cvvp6OZfU2NTSzc/GMVOWPxE6y+2V0BsN6Ywbh+8QuL5W
0jR1DLinPe8Om/SH+eX8o98ymnY2KgE2PoAtCepFkJNWYU/W5WrNNU8K+j11mgvqGZO4FRpUckmR
k69FoD5Yx8Erz4Lv85ZMSm7LEKfLkn110C0yPTzVsZKIwkkOl49ciB9C+lFxuQ8zZGh+p60mXgBB
WT3dw3YK4cCGiLUqVuPTzghtz80PUEx8Km6WCWVzghrhyApAJQKuhUpQwa+oZ7r+2lic96zVhusj
2EkS40uQL6zuDv7hwh8+6icDv8hoR0vcFXFAela7v7aREBzTrbqxJL1/mdepnTnGK1g7lu9OS/EU
OPvN9fI9pNktnnFNNsdmLGOlPxNJjVg8acQMCYK0F0IXIige8DqUuGQ86I86aU9SFEpuqJvh2/KI
BCMoH5YRbu3TW7D/jockP84JYoxGm4WkOnGB91y4mSHL6Z+7ZYsMzcoBers47uHeH0UKXpR5uIzR
y+Mzj2LcsQCaYf6w+RoJ7wYrr2OSoj5us4BCIpcbOzx16AGmJ9zOWy02lSzbQcbCTK0upf2eVmHB
mhkvbnP6xc6Z0T7qCorKKl2N0jFwVxndoC9ANQFi+x4OjDcAZz4Famx0NJJEJEnWHfwE+c9eVwPM
zGgs6uh69oL/5pDEYw5XV6Tb0eZbvBQKwzrRxFWyPMhW7e9nACMB12WFBBsS2Af7OhAh+GdnJaP3
eWF8nl0orJ10U1Vgd9NB/OfspjHmJ5LtvZN2h21JXImwiM29NQaGz6zb1D0ZXqXpxJbljn/c+Ynm
HcL8Ykoy+hwlwl80/GDUxvcBJ65uUiB5JK2tUO06G3dcCxdwYZ60rijwj2WoFi7X+KwjnQvugRjq
Tw6rqmeJCccUeoEOo9JtVx1ZydsILc7CNOkcjdotGBz5VszP0ueptZgb9mhv3mneqU3eQVp2NjPx
IHDXk/S70gCciqBkdI37RWYHBWzZ+RuUpxr/O6Y0Ngm4I6pXMYoonB+RW+h8je7BBznFcfBGmb+d
ITn9k350fGnG7qqsa2rzzDTdVkgR6vzpQphOYCXGrGjOgfL3Re3bPQ4tySJISrHT5m9kQzaBkiqt
9hGdvXj2pex+2DWPugHFHx/C8aKram8kam5ohNC0If4f4ZpFNyZTmNoSMJzp0xRZRbFijyKgzL5P
1cdtlR876TD889uIiA/U2qxE2EZsQnw0lJZvrYK2CyRO419mVMLI8oukpIuBRAlMmrsZoCt8enai
NXaOkUv5PQy7K+J3iyYGZ3JxYC1/Fx/j5qHssYlhyj4mYnU8QBSJW83E34icCRMFptUqzCwxfMfu
yKadq9PeY0LYNmdSXhOLZfH2BXwTaZ/4P3OPsHt/pfTZ/bGOgt+uZ4HTMaGACbieJEBfZouo1t6I
5K+VdIX5JDgCfwhe+bQ2l76XLTimeQ/BJfAJ2Oe2ZFiWMgxCx4XZP3gib4r0GzPS7UF6n+m18735
en6cpA4BzU/7AWrQrkNcPiHO84t5vRso3xzwyiVPL5hfTwHeC6QaG9lb9+DKbh8EWK4Hy1KO+RBL
t3CeOuwcHUBD0byAJpAhdRVFvnMr7C//J4njBa5/z8Msr68xOrVPPEEHqNKHzAfGzO5TNF3c4o5J
qIbDKsbzl+JsYh3k3KrImO8Zq88oNYn0vjh8xQ0YSIvNa+9l7n1Fr6atuJIAceF7r0CjnGMbUmwj
zzJl4rEv+fuLQNC3l7j1rw5f5fvcWp7XOzdzWT7gteB9rmt0O9k/ASsZ/Bns6trhSW10vu0PxeFM
CS3THWWR+MO9weL5kzdA0i354uYzgx48sOlY1pXZFbLOuHM/7WTvx0exiD3S/Of8ndY3WCQ412mK
nieWmI3tjXpLvSo2SpjurhPD4Tg5w/3WkrzWg+NIdT0R63pk7KPBnG1uCkX244Cf4n1XvGN+NcLP
RgPZd+LRQlk3maJjxK+At6u0WMC3gf5NtRIYe3yYExki0FGWt9yr/ejtVwTd5Xo13PtB6UGHcUUd
bTxRaSfLNEkWRmGR6xdjW6cShFd8M9jdDlltKbWyfAc1OtEth2tLWU46Ycd50qFSLhoEcho3toia
kHpFbToIJ1RaG7cCIdb0y0m/Ayq2PH+nT+eQmkwTpGFnPjWjEXKjv+uABlg0MVWaTHijjUUKVotQ
njMamZvYNL4+92po2LNXEOZwkXmq4K/KsSXASKPSVlfE+5GhxWQr/SJ0MCEPMnYiJmbuP6PG3uhf
KELrwzNNQMpICX0a21OxfWXR9wUEbJjsmBVZnkHGtZledyN0G9je9iE5uRIu78x827E8UHygAHXW
3ioI4d4IoLVMt5vwIQXy0bgIFDXBHxjRvaAIJArOzIJyYNY5CPjA2XTz7cW8nwsYowqn3M4FYYyZ
KNhEaDmThbC7Zy/xA7PQgBmoLoYVlUgICLGmYdH5YFXVTd8v37cQyBuvZFig7WQnhWY6bGtwZDVs
YN3wczERi21ZjeXL5blbhm5T+k9utF1wsVPDohHaMQbOUbQQ/D7w5pQVsSNDQNZCNSx6/ulzCO49
B7qFmIN896r5PYrX5REQhfTGvWMizd/R8Ly2BFaKPsVf49n4YE+U6zZwFG5Q+DN2aSWU14g5sCsL
3BCyoJ7OuC8SnVPaownAMwotjoTUKbmdUERxFGkX0kuEe87WfOr5SktQxjLjlSE0spiNHlSHEoZE
TetysYIZ5K31Mc2WDSXb+5VmK2plTrM0ZQUb6Eel20IYIluskSf6yxZgdNnoQTqsDQ2znWkrpzp6
Nz5o/Nmd7W4eqf3hXmEoZ+yAoAaJ2Um/SVPUQ2Qzc9LmNNsWZeY8+31X2yA1FGX0WIhLRKTCQ6au
pcIGtlpw7GxGYMEQSecf/bfbiBz+xoqgh7IPzn4+PMQzeusKQvUup98Tc1P7UQRJFnx3lTUDL4v7
DCsenjRK2Y1zj68QG1DSaGPoF1djAneDjQ2WBteGH1ol5QYpA4QLzSKpZBBrtFX2XFzxrWxzKeJM
WHTJn7r0OMiSeMJB2Lj9mjjIDARTY8QI0XlM9BFwi0r3ajP5K1xTnohSuqjfH9VesbFzCdX0q7mJ
nExcsHMpGCF0d5W9OcGlDMnuEblzbx6ZLkFgiSJmXytEQnSK91ma28/5Tc1y4Y85N8PL3UdnK7H/
QGeM69tWYeIP5SL1Jfpz5wCUQp4XKphYWBn4z9NhMFJqJcknpzP4RB6xgcUCbCAojprlDjWQ3dQ/
1l8n9tXZWP3OQo8o5KPQdBdgHOuX7JrKipWfmG3Nz59/7Un4RPoRS+u/FTbuHMuGuC2pePb9sPbD
spY/96YsfBXWmkpD2XOc9iX64Rq4XRC5KTO5adIVFSiN2u8ZPFsE/YMs05AW8VtqXVVHlAOx2Bdq
oSWLP9AzQE1JLV4Agx5FOtMf5+/+fvsricEXDysA1qOseGteqkKewVlJnSSY44mAQ2Qt9TyxP8aL
8blVXwsXgbmjMsS3G2IMfxYnQH/pvyhgUAYIZx2OkqwXIHiL4pfNWKGYJnZZBZA9gIx52qvLBFik
qWaqUjtyf9+PmpK6kIIGzwGfpbDr+SFIlBnMTo6uuLlgasQ/Ef5gB/JDmcTQHAq8g0hNM54x+E8a
/48qGV5Djc5dOd1e6GnVhuKOBr3q59l8WfPne0Vpe2pb4nLb2KkmuFcVyCxZiZxiPEY5ethFsVVw
sv9ytyVUIhvfcMLcA5DehJRaDsk3cQs+nbSQ7vNhUDeyThGuMQ94IfrVLHtm2ka7zUIq/hv61A/S
1ytZrU+SDI2+lTvlqgfNPGHbgR6xnu/2ig0wzo8Z0+XI3c6Qs6MMAC2mjwehDU8JWOb928upHWST
9gNsTNiQKTA0d3yDX35/4vzLehkwJBYWYhP8aQzJAZkp0UC69+fHfoCk78QY7tXwMBxQMQ25Zzif
0AxCQZEYZlYToNt74oHfGM11itIjykz94SShOW9IZgW21NUAaw0DaJVJceqYkR9QlROKHL9S73Ag
g5DmAE3c8cwEa7gdj5K8ciaJ3HmXo0eD3XxCFFKJ070hkt7po62AAXEcuFiRpXzx/LWo0eZs5lQx
VFtlJuwpVxzTDCvywAZdqW7shBRtQLKUl7miQLdF9hTBEErCZMR4jHt7qKADCYx0rCVSDNbhSjZf
mSYCf8RzBFynFBvu8wloqvyyep3No5kB1aw58WpLpEplw9PwWhyD3TTWqnrmNg2YWEthHsb0y4sI
ZYhZQsD8WeIamVG6JKCy216qCBcd1kgsjlNMYql/pY8V2oT/rGHdsizWpmAdfJnTm5M/8eosyywC
Z7HK7hF/gqzzrITyOtJgs7b9jmYU0lS12lKhcgaMoAP74OyA7bZ/ms3VZaHernVKDhXFiwQ7q5wm
4OMyFXTHJcwEp48DTh1NOdwzEnSmK0OkGyb4rbM+hflx1P6c9D/XO9iYacBXYmyBtM2yfHimCvn6
9s1xoZi3DVZcd2ed45nwXpK4Q5uPGdo6rNxPsh/t+y2lXUq77v9ibtEKwDKcfGexZCdG5DPzgJ5Y
43v8ELYS0UnIe8BeDEObPcYW5Fv7DbC4EG/QOarPYqvvVnFahXGBdNSmC/NEcfO4Y/WSDUT933ay
K0N9h2mumTYTuq4ZezKArV91woMv+82GEubYmFkLSvbGrI9WdWVnaS9N3jU4stR1/6i2tBu1zKfY
Ph5gIeBHNTvB0y31tHgIgKRezmYSIBWtKEvAr1L5qSEP/7vtH0NlkAFvdi3bRtKCdjMh56a6Y7PU
ZcImL+N0vQJGYxuXvoiDGfKB8Xe5MrBDzNDagn1/N5O2Os1u3SvcGpykZN8NvTOzbn0QHt9ytnR8
plXsVwkfGil4MNOe4bfaR8qkZaRzvFS1zouqIcr/cL9+spzzi3lQhE09/wGZ+tpTbsK+TXW+t2S8
JPSPYA1o94zkIRCyRzqAMVa5uIMQtwOxDuDzAk1DIG0bKNTyZjNRuh2JRcaOPPydqeQbmTEZUV5Z
Pdle89B2gm3LFr1p6abclx64JH81II49zW86bcW2RR0FGI/vSvpFoo1SU0ZcWiccZQ8M/si2fR2c
nLeTPlJFiS1uKXEoTNaTYPLSmAuEwOrZ7HYEgcDE/hVpu+JdWzf/gW5M5jCIe3Wfc+yY7l+TJMWG
6FduKGKVZjkznprgbsTkMbySeKIcgltq9bymqTB8wZHyZnJsqbf6yXP9yLfIs/kOJ7A5C3GZVWtq
owd+iSMx5dTQ3YKpmzfV9EaAQRDK3DmL2IqezrKe1aie39dXUeF1GAtgs/cIiHeOAcO1dnGuHyPL
bblpBR35txCz+9dqjTiYxgu+yvOSLBf/J+GiCaQkkRduFyRD/mroQnepHo4pLe48NIxfaE5axFqi
B1+JdO6ynG3L1Y2GWugv7m62p2uRgqYpLlpeP0Ea412miBmJaJpIHo2aXokI/DhgqaMoH41YLLeR
baTyo5q4Aoj5JjJeeQjXTXIo/CO3BoBrxtPrtiM+a/ZhPp2G+ph0hqS7q5cLKpCgLy8vKRF/keuD
Zu3GpuFSF3n4YxuC5kNdGxMQoBlAM9aLJhf22PdpvQ2UGM1f2z1NGAfYFqzYIsB1DzzS1ZZ9zuWx
+YLQOuS07pIgGm57qrxjGDoNUmoL8725ERQuI7sIkw2bgkVEh9DWrmVR2aA1r8Rr/kvQoYx6CCbo
HGrjAGUlOJBsR8etoyeazqiFrLMGSq8I4XuFteULNhJfNzmTFQ01E0kDCnlTtTA4z/+cAaAKD8FW
JfmYvBI4eLYWszb9cv2+r6SjS85UZwK9h23C0g8+k/t1Z4sOi3SKnhpU3jhMbMH39U5gi2qHKx2Y
KcTanXdXsNxQp0nAB4vWBx2Nwh08ADXoAF1Vmq2x1oWAItXAlKkS2dLWrQawxRVoc08h8zU0RolI
psx1e16pRi5Dp2L6UxiUz4sSFgcTCxj9Yol8xSckR18scEZB6eBDsYKuA9owRQcedYEpCYvMQqfA
zOCv2Q51ZHuY77JdNey2pT5Lnfd8/2ci5HlFciSAJHP4DB8iQMY5K/ow8ombOCDromiipLPn4WlP
INpARmSexhcvueHxyzHKYmUP6KWoHG7TWbX/X//hGmUwd9L7DfLbN85wLPs3/g1ICCSRSEKQtnoJ
IA7lnzXUobWNoTwECSxwNt6OhLzVHP/KF+UrnyUh63AMHohgObG+xvw+FXPryAI94/mi/aECbvIc
AxHM5KAs09jZH2y85lL2ClIRsDULFQAZCwIeBNWNG3yNipp35JxgEzJMNeaKEJJvYxmKzBm3B9i1
cEvsx32+tahp+nbycGzepC7P6yQMcj2t9omVUDvrCdYCYWdA0MwfaMX4izGUno1NsTxoN0gzJZ41
/apTjHcK2k4uGfZU5wbkN1Dn2SH5cPW1LE3lKonM9kZeWLVcVDQox1ZviwxKatxvcRQv7W6rAgyR
CheFN8jllGWoIZ0SPJsI5/WKzZxzbyCK3NW1PdFxZIwDvLck7uoKAkxJU9VrCl021YbjIZKIw1np
xc2hz5FpsKuTSrrA3888vVGASDHd4CuV+Y2vDxJOx2BlBFYirQEGviIsRXAZ8m+kxznu2Pn+iG9J
+cDH1f0QCiMfYlUBFTivMkupbzCYsitRvfH3uMtNIQDcQeaJm55mEtngXtTYygguB+12emNn1Jva
ypthkVWJOzmJ3gJvuKfh/7z1aHqlHmdB3HXn4AZkGCjIB3rVTdlQY7mdSGifv+QwGiwi5m3Eq3NY
tNA4Fp6degDNsYI/g1BHhuFbHIEEJ7Ftii5HcxsbvLrZ4qTA2EI1BfsuOlnRy7Abc77spBkOXl9h
0ys6BxHIFn7v3m2aqocUhPzQZXWpnsm1iTjAE3rol+ixK2hs9GbcU4+SZ2B+7fxaaso4BCrgneaU
7+0AlzRPzG2mmxbIYP28L0DD8lMaBVUPVoGbdKhnFLK1QEWrAV7IyC/DEuJuhqA7fg38guOhgRak
xYD4nWBu20WEDALJrxasvOL/xtpJ8dxLWlZ3sSMOisGU5+2gn4FBqtOy96y7O0WCgdv98E/8+isn
eRDw5nrRHn75Y3/P+lF04nXRy0dyrg649/r7lg8NeqpzieuBMzzMoOiLzhSxjVuwxE7UUUErKNjJ
02p393ivafGOYFTqk8GBb8/4Bzfcrzlba7J7IufLUYapPEUeEjj2mwB5JXGDrqeVcI1Yen6gmQxq
bJVwkZG8txhKDm2zpkdAmkz/8SI1fKMxF7eH8Y2QcHf/9SHNgljf1tF0zY5AdObb+Hh4TU6Bd2b6
dK9yA+XPi2vz/V39bWcLfn2MWh3HgT50HJ6Qx0i1iSMpgbQeFT5Aucrx+QR98Y9Fs4EWurTO3NyT
z+htZPTzQZ92Qp4xUFZyyvcDMoKAhHX7ocUV2BY12PWYC2TeJLRpPAAkL2hXq6aAsIVH9ktGbjAS
oZZph/s5o7n1O1eC32TzFC1kXPGBsrnaDW2ofJ0vt/aiQ4X6hO0EbGsAqKvadGFOuf7DBWdiNzCi
IO4WCFtdnSjWhD/mZbfPmuz7Tm9K/cnTGnkslWHxzvMAsUviIKCPd/RJysJvAn4LKnoeUCIGz6Z9
dMWOcLbObVHwfM2A7yKqP5Bi2Rc2qOERytwr8O8Xvpwz+GWR1m8tWbUbitt/SwayAz9oILhhcAmd
HsEznYDqwhhJUSazeKhpeCOSsr7/Rk2nLw9Qg1QXbRbsHSUyP1tPD8MVz9XSgaNLZTl/eYNJgqqQ
RL0AYmYmnNsM+7zN3HApENiGZOsw92ivG9S7RTUSJwSbMrCCRhqrFLvAZNb9DK5x6cGGe1WZRv0c
ES+7arzhWPps4jHP6ceTCezqWv3we0w7BO3IUKzCHFx1poJWFjx17kQIw2C/PZzhlzvA1golnIlN
3kwvib1O+e5pLmMMNv9kEXqB4hZwIkP7aswqJr+vi48BV9IyLvKJShxzE0XVGRqVvDKzhePWb7wa
upGOe88UMWfZu12hyPIquZJcIursxux/ml5AJYFonbrkb5Y3eDxWu5Va0PkI53dgxFsrcB1Fxsml
TaVxn+qfyrzDqGy3qPwvKs4CpL6+9jYE8M1XTj3xwylunnZ6RedI8J/uoQsTiY+8UMDFQFpUBbVq
0yQ+eLl3y3mCsqB6dP1EDm2D0xA7KlO7Kb+n/J3/Lv+WFgx5JoFaiTIgKllafrEglaTSF2mSD7FM
uXfwVOwNgzVtdsHAw1GcN85IqcQJjMbBGF2MT6BCZ2w6MBr+pLdTsNvLzVbY5hMiclZQvYadXaMo
k44KK2nhx1VqXfsPDceTybJyAtJyLu1Zrl4YFpz+jEG8b0oD3tpkeNGwwHGqnWlMVOTPzFYpd+Iq
WFjzMTdu6yiOaFKZlux6j/QZdgV3p5+VXc0KYf+CtcKJNTWj5AIOX3MBiHZtmkpd7/hszfLFemu+
tB0+kmddReL0o5byNylGUQLQixGXE6y5a1KiKBD74eihaIecwdYCT2/ytVMRenR/shDBRQk0KJ1f
dcND7j2jdedG5keAhHGJUaCAhKDy8PmfiIWyFfw77/duzNh5OPw3G7i8AePjjYcV/GgJYS1LjYcK
SUcicgqTvRKDsDMIDboEMNYTMyLV+rxQWlEafLvOkhiKBSTmfPTbtT6mYHbxp8NAC9GEgqlmj4FT
6l9EETTB7AUwEwevnflhqVuijKj5sJs2D+iDqUzPTMgdSIHL6yufhLRjHTpRq/EAL3impyv6ssHD
Gx0B6/jyvGUy9MyFIC1EWn8iEQ3GyUXFb2Bdc1OPX1XByWgic0scQxUxGRBKsrithSmebxmRyCxE
ce6WIa05ENGCsAM+RdiziZnnj0BjzlNws82GLDlQt78t8rHi09nyR9Gz8ZAkksn2GqzJMMXGL5Hj
X4LieLQ/VGLL2zSHcQYtALYbihgX/E+jf9SzRN2FlLMAipo3F+Q7zrL0ebdb6b67k+TmgLZE303u
Pd1JBoFArjlsqk2VgPtjTDa6IIQnzhszR+VjDJX7LxKF0Kv5rlUCIxWISenPPJj/p9d4uFKLZevd
Yi/znVcc3DiXiRQoOYIcGdzGRc6aPruWjA29B+PuzaCDIfG5BouFzY3XJCd9cdPA5ucjgslNDsOi
x7LDYgwI4xm1mopZkwrPAvuzGmI2darr6fxx8Oul1HPPjKSIMjLioKefYBGStip+cT9UT2uHJzOi
Vrb5qHBMe51n0ay559HJxawm+0ra1tB4Q1WvI9GWS8ipA64RtTL9S2b93ZIKtcG7hMr193cWJvpr
b9wTq5uUYdUZ1uh7EdTM/zLOzzmz/hjh3iE6JED8jbP0MggYubgGDtfuf3/gGQ/GBfLQXc0dIBxQ
JIJ47vKE95NBo8rSu9/VAHFYUNYNKDefa4nB/G/3EOYSuwATwQush22Lk2aVr88TOSh/ukAFuER8
MjccNEGXpb4HAJCNUtLXpp/Nkx9ImMBVMYmaHXuk6GukizGXf5IkT8VHYT1RkMAdjV1SDRTp7Cou
pkFJdR/r1jDKwkzvkUUgXAPAQXcMQ7RhCSsLUofVHlNDd9P6GFcNdJ14A1D5Vq2gGGL1lt7wvKpn
yl0gBUXHnQGnR9M8p8FhgqK42GpfuMbCikQaL/HOxWdxSfWXCAlx6BuVRmRURFXqQnHzQ2Da1Yk+
gq1/I7LTwAKNWXCb59VOgYHF3vW2vgz7yHxZFfei1NFlP30B5+py7rsRBdNKZp6FHWVbpXJ1Gg3G
Dff8ByDXzDixy+KJhc5xtP+xil9AYlOqSUzoZTOwiNG9yGz0piz3w5DhSGEzy69ImfMaM8p+maLP
dHXu/e6C86aALJbMJ+FHy/svIdXbTpT45BwArpHdfUek5ofYbRB424VxiyHg1WuR8TLhl15TtdvH
87vwWjce0ZjxVXzd2rUx1Lwc99m7X+VuuVEQbLjx4x4+ldqYQ4MO0KxnJQRupmzVAoivJ5YC3vff
gxpZY05blRqxbLhgMKSeLRlLiGCJe83kDpz7CNnb5NEsAVMxDFaCB/G2EMDJBukH/QVi3SXPOwXK
FAjAe2QdNGxJY77dZ00UwKBAmi/DXt6p2q0l/hd3w0YCvHMgKBVkDCQr6s5yNrZfkZRO3cRPbu6r
m8DL2F6FCcB7LcMFgPQasztgCzwmi0AwJpOTcWKCjGB+4PzCwuQsAhtRGkKmmBaQvsShF6B5CGIH
7j2awvqQJASDiCDwiBjsNG4dVeBQRaI6Zsv9IRT9qeQeoCxkz+1womSPGzlJJ677j3LyhNFUpVAg
5BTmCs0VioBTnGsonVhNZXbXv8OGrQG76Iwt3VUkO7SxjyEM9OarlIKRCqv+HbV93wV8Ky2ZDpQk
zUUkKyzXxk+ueiaS+Q3+4QyWVeCrQVjOsx3bkxfuIQOMkdjGbjOPTsbyeClKI1pd44m3JIQT3i74
HMGmrn0qScoQNhVpgRgigyfi3C/rbLRXx6wxV8pO+6JjEsr7W2Z76KPOSfo3VcDRh3otRo5mTfPj
3kweJ7aP0JFQTDvngDOPLDBtp5lugF+LIXO5WNYXAl88VsDVOfpdF51kuAl3qRya7fedU85JV00+
stvAbeg8dMq9DmnfmPXD2iUGkftd6T39iIcLq7W72C01ecmQDJxLwLbzSRVSwFcKI6wJ0NYEJ1Ew
dK0EkZaIpg0eT6biiIl+2dqGvgwUmvFAm+CsK5sbWzd0fLSTiOADdqyuOzvIcBlYucjMAIPAVHcZ
Qy/w11R9itlCffR/ardtcIg8yWbiLPMnTF5M7ngU4Q9ApAQUPnUMluSO/hoHCuc2iSrI8HRzH/qh
JPkYeZfiNRNN+p/eNXPb5tAYvlfYuXQqZOPweft+bv5tmrAcEdKu5WBVWt0wdJrXI7edz+1JiOz1
oXyIWoWX0DuHA61shbafEBSdee8FmiOVRywq4Y54V1NBsO5g8evBtCDwa2l9w7lkCtxyIEbCYOI0
2RymKJGbyO+L1L91zQQAM/BxFXraqezg2wpydB5T8EE0/vvOGy47VYI3sAhjsZp92DTn+iFIHn5/
/xVeRDZjJPW9cfTjjM73BMxHJZIvhnaHAHSTMQHCGwh4sFRjjvzwvB9n7yFikts7KcS1uyU+qjYl
VO8zN4d17ryauQuPbX9ZBWbA0kX8fMwL9A7W3FWkyPPJ0fSeXas9F++ZtA/lIqNUsSLXsO64RcXH
SdF0YtoL6fS6mvIPFN3fvp0wV0HQjEFGaJs3glHGwtpRmbDc23//s73sJxezT56akbrYLimZBcE5
8/5C5IbEpY7u5SsyIeH4btJ//A92cxeANReWh8XfrXdJ1eglNYTJBlDi7hW7tLKGeWh3hwgnJNis
v6tWq/OvEesMiWUDh5GZqdxbqfbbRI1JvpSKX3TvItJa8kUFd6gbwZwtdqm0xysWH4S3KiPQuvyC
EfAhBUlcTjo8swcmv5dvySflScTrKPKmu6Uvg6hRoGI1X5Kb1rx6QfaL5zttnQHo2cdcamu8pmHs
gFGfNjwUpI2hzl603cA/wAdgoF2RbYsFCvT2ZKXAygeIB1UPJECuJ1rWfsI1Rp7GyogZfLD8bShf
06MIzZ3g2WTGlgwhWYkih/GKvQWgg07TKHkUEJu8VJwW/GJ3t9mOXq7kSZcZYiq3zZ/pEIA234qw
EtfI47fybO4DSaHpMCvunYXPt4QmvdaovZvggEN+PufYCZ1wt0EXVk4OFa4vzAJ7k6BKVGAvCLxG
fmNp1WiHMTzyjHSBgyqxFRvhEXBgvrUPzu9/CsBoWCIKGgO2E2rCRUrLJvjSNgOhAKlPU3ytDXy0
nTBP7plUjE1pDU+hXECztdsHXZc9Vc3kI5pyQuIDwhgGHDDJ++Bd8pMkNdCb6vkVjr+s+NiE71dW
vy3NKjCip3QNeaIk935uq7lDLe9bNclhbBZcpLWIWL8JX+kQ1MGXBKRO4DtZ2bppPkgr7okLbppi
h7CejzwJ3rGjEhVU+MgPH28a+Zi81RJHRzduJ0BbtRG3hsfHnXheWYX9Ru0gz0PKlcZxHuivOz9N
VdO44SD1jjZdjPYCIsQTfVCRH/AWL9NRIKHV0QcM0XVdMsTBMwGcB2aJQ3nolENr5uNQyGZdCmoI
FUtSUdiXrEcv3ipbnzGXVl1I0MVYETD5dgt7YY6sRhMHXjSm8/CPmmCCU0N2ZAuV1Ayl5G/oFhlr
0YsJA8/+g5mh6h8e9dh4qQwj57vJJU+JEHE6NUhvWHtCyRpSK92mcrkwm4vrrq/EqiMDJwTMyn//
VysOjABNFi5XErrgu0O18AqNUCk7rJZE9gWlGlPSQr6A1shnAAJ2L8FyzQKgluH7xQge8hs+eB+U
Nxgg2nveHSgSYf8YirVZmUMcb358F0ltML9mmWLcM2shZ1jwpUQFkB+W6E9AApEsJi4O+w3s57X0
oplNrLlNwvXCMCEH70hHvDnsy74L3ncEd8g9m27ZmFVpkBdLNlnhXmaF7sDZXZr5uYbJlmbDKxdD
tMY0+LMKMtaio1PRxVmH0bmGqeLGbpVuqlz0Dse9BlbtEVcEgUllzAI2907E5OEZZOQnc0im883z
AZqHVNM/k9loQFE5pykNRjC2RiDSOjiqWjJSzWe4UNcpYl1dqIGjF0HEtClkOuMdMqE+l1sRNXwX
+9YxeH4BIqjGmPdrG4NRtzPIqBJ7XHf3WjrqJ/fD9uy5+2J07Wy11GW79CVTC0/CoIM+wjHF39S4
+aqnUqzfLfR3/TjjjNU35yovsQyeBR8YUkMZ64CnpxyqLlVkEFhwYfmIFl+/DrDxmzeYGOYW9dKL
vM4Z9kqN54HnPsHJmNJoA18RMCYKtZifPH1Ylp495CAobWhQmePdEe+R+08ylahBOUu1JYHcuMLY
y1hhbBe0jg9/ID/840B2zsrCeTkkFuH1vPaNoWW+/2EhqvNcrXUtj131K99io1XGhTGH8bKgDU+s
hKuCMCXk7H39elzfioE43Qn6FDIz8rWbeQuQPM01J9iZVn9iQH1/SyeNIb5tFWeFUynStwVoDGeB
oLoe7MQhhMWgku1g7Vk4KOPTbu6iKVuLsJpi37kH8op3JKoPa3eVIVj1NLOwiVakfWzDX0qdpFzu
0vtXFVXVMVuoieOnWNTZ5R58bxtEB/+oFIa/ebuFEpwVkBGgRhmYespXql3keWrqwuBDnHXBBCcM
mWZum7KBNlKSowqjw45SHbb4HK0FogePIKAyx4LF34CrKRUPeKA+cBiwdirJfVjzR8/cpogaHypx
7vqGW/E2sBOEbbNRXG8Hoqdeo7XBuagoBw0wS5rC7by4Rr1QHvEGCV6xrYVV8vhFBldJam83sa5U
ide43Op3cVFUD98eb3dPVXPZhmmRhwjMjle66qBkIcrc1ALrt8Ua/ilx6uqYotW4/Ydx2mTpvBSH
S5cQfKLiTSy9IBUOUbWH8q4x+YYZjzbasviZUxp4o/axvH0GBguXOCxiSyZK1Lk5q6Q0ODFXuV4Y
rWQobgAql+Sfbj6+00ACn+C306bmVvrUp2VrUBkjcPiuqqgn/agpPZM45C1hyG0pX/Bzw9amKly/
flks7tPwm+nH+4a7rQYdTO3c8QWwUt2LtR7ntCnT6ZQv3HizbpkxuQ0TslQgOzHqTZjwbzapiM2b
zYytZiY0K/bIy+JuZRrHXqARclBqqGgDheIIJnENswfRrA6AulnSFcmj9Hl1fg8VBgBg+JlkjKg7
lNdrf7WpTuMPdn1bBwvQWA/3sGvVejiOFJ3x08o7CCh14dtHeyYZVaeVaQGPhz1oA4lkDuWDL1lP
hibDLtSfQ4dQEPvnChVGDT2OPVEZhI/jtunkLpOoM5LRIDeRxR1hOkMaTJItKeQqnOvA1V6ksaTM
4CaI+tihaqzOCruv+TaF1fPV+vYIUbVD4J7CVRkfDV6reMJXTY0tswiTvkfx4/Y6W1vW7KKH9OPw
dHZwDPHmWy/bInZQzzNBzf5nTVZbltt8CR1l8X2fU/H3PdTcGFKxAnsy2Ek+wV26EaZFukKqY+59
LiOy5LE368jzNpzwfStbv2Mu8V+Icd9OGTSYALV+u8mz7WuLgaU1wWs55wNanbqZdLGUIjpTPNaS
da41iothqaA9fHIFeyADq915lqxg+rGPQucuknGP8Sg6tqOeahnQXIBBkLPPirq/QYLCZFqWSjf/
w5onmlE394kdOif4bgrLX4LFlpzOmYKasc1ohqlZjZ0uY1BTn2OMozh4g6tqozwAZtEGB6FKw1wQ
QmLp8ktQkhNNlYw9Dy3d6Wk5wpvq+xQXqPVZubocY3esT/A1YW1sqZp9mz4oEpha6UtaRtpZYlG3
Gl1tKT9u/Guqztw6VakDUZ/7/J22I1ZNTZuO8bdOI3i5o6+O3vFTonJuMYylTVO7POt0xbya5VNT
CIoJI4EnS5QZqVG3zHdvihh8CdWC+WX+pudOCI0m8Prx6BE3spEtH1lAh7quakHIfAs4M3TREqvQ
HcGODeQQQ03fcJ4XQaYguauwGbl/RtNsoumcIyFEsEvajYRi6nwWbZeNVwZbwGOaqA8o9NAIpkQG
IEp/WLA5IiZ5vM3U7UuOKsswXgyGnBJqo1eaE2RlW4ur+rHpxxJkko/RWzS0kxY1kFkJeYTkB45/
RNvPT8YRD6TH+Oup7U7VcWabTcrbom1XxVJLV4rjwU7rDfp+NWN9mcOiKWUzYw13i1jPCCjuTCXF
Uob/dZq0kYBVwIpPn3+7C4KXZZKC1KeSHTCWfyxbG/7T1JvHarvwMkb43cSsUdZDpxZcaR19kAwk
7TmSfpA4vytUC3NfJL/QtcZ+sMCI917GDgIuxy4nyNwfaO4g7a3bBFJLkT3Eab/kpxREo19YGCTD
Xq1Lpyj+tj/BCeS9WdaqUmM7QJewkPrFkNnET9QVo9T80avEQQ4fQohfZ6eTDI/mHfCttahy0i49
TOuc+f/g75P42OqNMuKCHhjAgEFwbS75c2+jbJ67i91j2DsPaso/x/Kj17ERNcIHoXCuhkPs4WEP
CIG8HybZITw7GSBdsfEQDkHShNoSBtxpKlLAFYZA+tU+v/1YNpICT7v1/4T9guPFjjEeGzMihYUP
vWMbUsCBPiAzy0BmCDKfgmury8a+KzKt5Dy7QG9mX1FoaNsxOAonBHjl6qSE+YfVyy5OVkKkqLXI
vxMyPOG3PAL2j2WkGSi8dVtCbZJ9RqlT2VLOJLe+fdUhE/uJkc2godEUpBNgTQG91Aslua5IkfHC
686dw7BHLSQ49i/kQ2j9dhXv4mLw66rD+rwB8WykKZZ9NiWcIRx1lAgGTi8FM3RaxUPXamNwFq3l
sxUVObuay40yb9aEo1zpYodTOzdgnkKGrKvVm5io7tlHAzynyPyiBH7Cd4uNBOGzSsNii4wAyWpE
h5DOasZtMvMo8TrUGZ83wlzIRXm8jDSN3WrpKtthrwzydsHM/gsYh6VegODsWsbSs1bYpwPXU5tj
jCmeMJpt7E2ToWufe1hS3TFjVvBMakt2LVu9jHoohlZf0gRmJVgrdcfpYZdtUo9N5oeWG08+yD1U
QhMku7u4PVlY6+YyBZT/Fp8QGe510j+cqt+qJXV1NYIwGlHEMgj1dhIheM1JGsk4RE1lbXL4IFa4
zHA9ZMPzWk63RZtOEb2xgl3aYuRButS2sW3zSZxH9LjTtlydenC/tXJRb+LZ2U+zvgsOttIEtZ6D
KU7LVc6sGBAtie+saX81XkkzZiEvNemY8UZqVWxeAizJmS46j2vw5IQa0HZqo+UgiwRJ3R9wjVoJ
/rWH3vvwLDS/fLwNNFz3CjdwfINnmhc7jY+YX1yLfXOsdLbNAnmzVM9prkMwdhi7roCidP7HfhYq
J+GhYmXMeDEzsF0hIa2jbaVuIFVq7Fp0YogQB79kkPYJ8uQNBjaFayONS5/hqJU3SYy1Etn1/zhv
JpjxcxctvIRFO2CU/OUduW6ETVKyBkF3+AFGFDCkxtAQAkQGSAqJeXnejw/Swpmw3mbiJXd8llPS
5deRA3282BUKjdkB4NNhP83X7yh8ejU1izpK1/y9rwOW0y2XKBae+5+HB2wNR8KtWp3GKomBRoaG
XOegQE0/0EXXU8THQXeq8sTrBMCyFp/HOXSsIo6DSCHdmAPoXHboYxq+MPie1kUKzFfUWsu+aezS
YU8vLi82qQObfG97sWKN2ej7hP6Fhc8YCeVEOgLyjw0nc9jhboK/QRce/K81lkLjYSeh/SiZE9ej
M2SGBae0WxN1T15O+5ohnSC9sOrBw4Dmxx3e/AqiMwdos6C88xW7DSbfUK73q1148A/eCN2fWAeI
nVkGxegEVJnkvtZJLzCk6anqjDckTrtAo3NjnBsWEp9CEhhEJgq2NpduJ2Kog3GlAAlScvRmjAhE
mg77vhVu5GFt2hv8mOxaBHO2rTYrZ+ZwIeaur9HmfLioLFA4SWfpyHJsmJciX9Iq1N0iT5KDVHmL
wonWNNS9kUj3K+//CSD1Z4zqs8DQziOd8RzerjSDwtNgGDiaeqi61mXsXzbpEqRI1ogZhFWt19OS
scZ/ETfr9EzlUfI+qDekUsqYqs4jI2v2zoIDMygOpQzvgnFqqii+VdO5wKtgbqtHTcbRTRG4va+d
ye4pLMkzt/0bO5OF+xF+VWkxMxp1gxYxBYdRbvcDD0IbTQVF3Wp46pkBYKGy7+sU6Q9YyRVYVCFs
3IMv+VHY3vXcKz+L80c1YWCF4+7H6APux1nAz6T9trbOQIjZFQg/d04M4BeGPtTMeMnKw2H2tUQX
IHeulSU/QyZxh/myCW/i0tCl2bja/KI9kehsJriUCbSQKJ/PVIxX6+dB79Q+BL/eaZCJVIYyEZSc
OcRdo+rMfaB/eXYxDSQO2am4JVUmDsiP438jkw0bf40SV01Wnf6fe2XjboQq0bPXNUA1+PdOT1lr
kilVrRcLi7OylOoX85td9KsmkkTPSV/fb0EG3ccZ3+shNGTRE7TfJ/VWnHimS5xKrmD22K95wX/u
pBv+4oMTrxhWGCWjmoMQ3k2nmg+eeJQrSF8x72esuOT8ttBpnIjgsd5Ar43tW9YWH7fARnf8emgx
R3J3GvRIZw5/Rlp8NBFNzov9loO10ZPoNH6/zNYiHlL+lqQ2jlkN6neudowNoBD7y6TMXDsw353f
wwPf5v8J7teSvMOevc6NeSV6OJeTPFqyXRISG4PeQ/DeOAUbj/DUxTC6uv6rma+OOFpswwF15Wfz
Fh7aD39+kBmO+2BcaKKP8jiTUHbymL7q69Q2ALO76aqMVk90CljX18z6pEOnT5BOxiuuWinBmJm4
iE40s8gB1i9hOV44hZ+c98sKJoC4lL0E6wDSV3/MQTogR2KnM0xSf4z1BSy7PMq7uZJNdMjoXQh/
eC9auWCtP5SdjV4up+NoopvU5XbOTCemtTU1UFd+17psznJuiJf0l6p4lBofmiusq9FdEyoY1/c1
s0iLzdxJze9TK8eWXp1wlxs35Cuf/sAj9KxXqpvRyQxr+FhdpvMy8NddFclsYdNTL7JWeGJE3MYK
1YRgVZV87xU60Z4xtUqtsvT+9qnqRBAN7bB/yys9YxoOA4Yy+GL2DUp90yRiVqPKNesuGtdeDsHt
+cM5f0UmNsHSldEiIYlAcKkn6vuZJ6GySS2lhdK9UnbY608xHOe+vl7kj0MtRguEhTmu5XW9NHgo
sdrceih7mp0t+TtTQgOmoQ58a0ACKe7E63G7WZYrDwNwLcu/H/xnNyn5AKeRWw/o+m2YZpPVci7u
ctoVmcqFpG3hYK2bAT6rrEk/v3oEhlV6VPC4vVw+4nVZLSBZ8eXuCNk41sza/zvmGjQJ1UYTPDv/
7c6klv9ydiws80XTqwkS/7wO4sI8VYZz5ieRitzPV6onvSBtMtHMsEy4ZBNdVOo+puEdeQPaPEEO
WbjuhJQWgBuCy+IXGOyJC/nmpPmiNiQxj5xUEMgursELPTlZ1mMR+XljPEzVH0U+ziZ9lSRl7j7m
NU+HNi/TRfP91Y894MsyPNwShl8HR2Uqv3NMpDW4w8laqc227TiSvQW1qvXJ7XxrUj+g3FYvTCko
966jgfi77JRiivbaXjHGX77aePIMHRXcKLUFKZrhoMPKsfbgcCLJBHdglm+fqGqeqRYKq+xucZal
7A6qXhTOco++r5rbGjqp7AFr13RAs0MX2wysTtrQGW+kjPj3pAjOt1vi0gw0GMGDT02OZpSlHLMX
t7rKXgc96C1SSdTJ/SjnUYmTtVcOV9pQnfmWv6R2BK4ZgGAfbqLut8rKrf6era/8+Q8/5/KWSuMB
yQGgUIzCQ9mRrra53j/OZJqGiytPuFann6TNDhGLRozixn5kV9OuctJtGm2SP43Ez8nxuEO4jVtP
laLicANOzfe7G/+IayzBdifCTVvlFD3kGxuXTaoj4cet1+Yd3D2flNugzH9hybMPE+YMIZrp47Ap
GQyIpmbhd2SkAsVtpNdm/eYlflQYU8Vbe68t7kPrhTChcaLpRfA+zDldR8k7nsYVBxMgUQJPiIHN
DpoIekoHkxFQ0PUqQBNEIlyCODE9Bhsy2NLuNzxiDuvt7RXAVZoMXnHCkacd265qcEJWNrQ2yl78
0vTAylSsOg4U2nI4gHVA2sprpv/jSn8dBcgi7dtbagvrScAAKtvacAiUdcGc8sbd5V1YjEGKwGM3
wjrMwtMp1yDxooFZeGL4SLHzSda7LtJgRtfH1eXLIBJDmWGZtR04bKqzTyAp7U8WwVJvhoQUCq49
dTh1lRlxp2oDFB19Voeg3VlStAB39S23V3vaxZae/Bf30mWG75s0gYxMAiiBBSGVn0nhMGjbLUCL
FL/YkrEo8Rbr5wPNQHAG1aByW0Jnzoi4YrObWBxVyICCk5XUJIBRFI0ug/ODWBsEOj8x2jQsSa7e
UqYdslhdgClFGHqlzyD4kqP/2/QbVAi63YJ8C+kgC0Nl4kCd3C6IO1kT6doTo6SUc/8PHWZQkeo5
yZ4xlZcK8ubAJ3ddEg6Cg+w8MmuHN0DeYLXukCTwgVB/z7Cm4RYgZ5SL3/Dp4Qcc52NaDTEs9r7h
/wUcBMi9TyzkPaOAaf+U72NyPVrGEjmmDyBhB1nujlTG9e2RujcTX6Dpr3Yxg6xvAGKZrRn2R0Ky
mKqHPKN6PlEfYSzgXzqD1jopzd6qLXAck/hCNX7IsnZQ3k11qFdWbRL4P//F/ofPbi45ZBiV5XN9
RRCU6sg/leUejphukq+lQscCYzxm1vyLK18EAAgI0TjVh25tVwggKvuOMdjAHYaUwVy9rvWWfguN
HfdK74XGAmGWbakYPtDB7zBVpwa/Au8rAzkVdGFH8mgdUJmgoKBfVv8ISZmi1pffgfg7aquZXAct
fNNsPZT6xQevXQzPxYpHDyYSRltszbKPY0T9dZ98nJF/bz/g3GGGSMDR5u8a4BdAyGurasd7Vf02
AZ6KMPzeMsDtnmpslHpHNZ9Wxe7X6QKbUedTNwAKPr2x99d0TIrFACgSTSkyAdeT7Ja5cPzmFO6a
j7GIvTaEDtRc0GUPKBip6Xacg+J8+gL/WIfAgl7vy1Zz/EQ/ngsVDgRqcjM7iWuLTmFYC4Xen5L+
9u8n/40kO8hbRAD39OsrN2JV63SUARi0kQz03W/VSUXd7Mt7zsrlEQnM4tiEnNOgvpvp6TXnhC4T
UP4FwRxF9plfuPqxz894T4868ZK4+A0UgYQFsHswpT61EHrz60pAAGN3Rsy2rEYKOZ0Mo7wDkuwj
ZGkPNySenQemE48BHQ41DpGPXW4utDK/4vpWJBd45VCTyXx0iVdpkFKczcdyUtwqREVzhytSrSPq
CL7Or7tEHPW1pp4rNoTihhVDsLyE5fakqVr2kTQjxgl30B/j89krb4nkqxmAF7WBlrgVL2eP739o
3fmnz6xYE+zrRlRynS1Djlge5Ft6FhrOUFjZRld/LneLL9VfHi/BnGXm55qWFKXsU9tyG5tqemep
6RipORNnBDGnbFX0eJzhXw2xWgQOE8Y2JP0S46EK0ML6wAb3L/W+P1syjj+oR433wDExyMiZ3oMD
SvOgNn/t0zsBcGCDZrTKLovXNllDHLxs30vA1cOxH62DcZC1qEsXcDSRzfjR34SsWQMM2GPdzIIf
nCKGgLzGvnuULRNDRDbYkZUgYLrTho9Y/UPC6jciAu31fl7GpzqpiH5aX9ie0DTpAG3hEIctUUos
YVoRRVEfTavndVDjnOOM95uoeFQC4dvnidDVhTMlIaydpccEQvTBA53q/rotcfG9yhomX3On3MHi
evuJ9lLfut25FDd831n7G7p+LZFniZi3idENrDRQQ2VbQzIeYKp09Z0bFlCd+/sliX0uhCcQiGMF
36H7A7WuKVaXLV1/h04NBEmh2P7p7dzKyVxxmcOZ8nXyHn7aqeSnmiJbqK4LAoG6SIDJySR2tars
bGvC8Dlf7d0nEzJ6Z+PHFyPlZ2s7Cay1wX73g7t0m8M4FkufRZhE/Gj0W43iAvbJIt7HCGC9o3fe
CEp+qS4aQYkJwmw0+IJDmrFIEEdvlPoyHaaouyeDMiTd4m9qgIuWITV8RdssKaa4pp/uUCBv20kZ
9DH7t90Bxf+NHmC1x0rEjzTLighZ9DagY3JjdlGgCj2WaHuhcW6F0SYHDP2ctZP4cYNFclZS6YcA
ORTMlruAulY6Be1M0ojoR0m2PD3AMJGWJMS3PftEFw7r5ElEzAXF3gTqOaPcjsWOS+24/8wJHFpU
IyvCDrXvi1xtNoEdswxqE4DZ1r9KvppUSOqthk++UHayG0IMwEX9T4m1DDX28Rdvy3aWWD23WNxo
mgMTc9po6O04ZyMVrrVP66zq2E7FJ1SyD2mUZttbUJXMK9vdZMMK+Pe5hNQaz7DzLMsUS/b1CWNB
m0/MoaSCDWx5WW6x4u4Hatl3XMLQC6kNrMpOxutlieFPFyFf75SXzz+nMhPUTwtAR/M9igNlVnWy
2HsefMoB/CYSsi1d2PaMaPlUYDmSEeqmPbesSdBk1oG6HyRe9PnlWTA5MfheZOrj8V6oF4MPKmM9
Tlzv3Cq6doHmgrl67WU7OecqQyIBDeU3jrKuCkILy2vbR9DHPUyrJd8M/U9ajlxNyVRXkLdNIL4a
ZR6xZ3TsmFnWf8CrJHgZYBmEeVobeDZo0KPZBkqmIuNd9081jVvW3m2LkUrA1x8JCKaMQzsqIhxy
uJeE2TcqeUWgGBgc7Z4RMgLk3OOHwVzt0WPMAcrKgZEGoMs2YJOmLIMTib6pSN5Z1oOWmHjPc9AO
XZN0YE5pOe8bzQl0FYABnWY2l8nfJYM3ta/zAbDX0lhf0c0b1O0a9AxtXCQLo//xs/Ik5peizTMd
+1iCG7KhukPUKZqPB5zm73/obIgAfpARy2C1rGqGthqCdrgtfpY7WiKsKW46msoqeP28bes2BXwE
hob2P12rYcnoCF0MsCw35OJX4MAvuumsrFWdfh8mncFtLTe3Vcvfa1oinsHK+AvSIF4dt4Bpnamg
sjJdOh4JvnoVdJhyIDcbA/HIe/xVNxAeBKO5qIf7wv0s/GPSpCAgMIc5g/g9fkPavpygF6augqLN
sOb7tglfuoYoAZM226J/rBlAPTMY337wHhqu/M9uC8e6HKXAE6pc39MiAr7AQ/2pgy4rMQRbLL65
VKKxOHPXxa4mDIyTUM0W+WbTNjCtospzGmZGc2LPEE/NiBM5J5Y55uvB+sTl+l3RFAITEbedM9Ub
YUv0zxzHi1A3Cocy4jQcyKXzSe4v03BYmi227h8loIweDNbQyuUvgiRGrZnfnyx2aGf1T9q7EVWr
KkvC2NQ4pXdCEeSZwmTgQv74hoS20xihEDSgKQcKtL4NxrKiO10AmmFGjOKXOfLdVLFaQj8ms1I1
K5eKLKBxjHouoS+PXFs/wFkDi1WS26QaoJxriEJeTLP01QP98sapJJjYwXF3JUi6240ZSH6AtZN8
NPHTXyAEs/NZXNhJg72yNr68D2AHchcAU54lD7gsVseJNfjB+S3xq/khz/EPzL6iuWoNWC0Uub2f
c/WV5wQtPGLvT51lksyHZNzh4kEczOlghvQNUy0TzQBj43pVuKZfnsUJPvtpScDICTJARkF1x3fZ
+oEtxRX/29hQn7mJAFYl/C+PeDSOlALXJ/l1cOvo1iqe5R6bfCi8HJQVkVziSG1JrX2ZFLkHSsJz
yGgtFA2O9jVIcOKvPnqkpIq5y2SZ7hT8tcWiik4gRWTBRlcM+WXRuUBRuMIuTAGqNLX/VOl2ROsK
0MtTZIG76qPY8e6jBTWwQPWEXK3/mBLpDGMWOBKfEDVvfvgE2/9Uy7BJx4au2HfhQOfA1ZsPrYx6
RHgVWYgTWufDfew7u+dYKJvUOsYU5uNAot3SMPnpRIZEzB6lN+qUj7W/lNs0MPzCaufU1WRPzUm+
dPVQdrLkFOrHABFcHUzClDqb/fJXjCSkxitjNGAiPD3pwM0SJwPGV3KGgkDzlC5LDs1aC8YiIIXi
DxnQALco3TkMK4HcK6YruK3de5kj4bIzLYn9EVHoERg3zU8PaicJle92K1X8sUcSOmmfHdXTixkM
3lNBZvbiYremd4DUtT/uXrUnJRjGOMbzjH2ZPrhmKmUQop03Mmf5u0A28SrA5nk4lMZlcX7bWQ/V
HcnViSSApoqhcm3S5svmRWrlwgEu0u4U7JOWz8inUEMc9nTvmayAG4pxFWi/blwU6lLPZT3hSoGx
wnBiWJFfhY3lzZnbxSB7X8/kfKkwmdxksu+tZTnbUvoeWM2jDWMnhHYV95+nowgSVj2om+Bx25dP
iAdoZNsKpC7zAHEyk6L2sitB8OlKFTuCA/rJIgHjs/3gN0Y5fBV67+k9Tt1aU7LJmmt8KbH8pWh1
LIjaRcdmCsI15JL0m/+9PPhM65mNmlUZOWyETqPxQj9+/VzIp+9M6RVL4J54KjhG9ep43rQpWlV/
1gvREraLE78OwLpF1XN9cE0QCqYoj9SumgQMYMrbQUwdtbjGPAr1IWyXhnLM48fCIAAghpkezdBq
jvxOB3nF3tROkRmi2tdmFZ419RzfX2R+AjTUh9PDiHqY5Oy1Sxg4gJxsnJuLFXV1x5kNFjxh/X+d
ZWgrENc5sW7vd/LRGErLqiPuR9X7Uf9473uMmasiVCbTgcyXiWN4Bpki86tDZxy0eHR+AbZO5nF3
p8ZH433yHsdd5Bur9g/Cwb3NxC7zZ9i/vJwPPWYMGAToZsTPrRjkZ9MLV5s86j3f9RWUK066rGoT
NWJcDV//l2YdF936d/dXvOXEAbotnjRiQDs5zVS48ypNWHjyu6Ab1zY4Woyv9ecJnFH61H10YIQj
vg8ucRx8ocCPzsEKu/e+YaUerdyi/8XgMay74KautZadQkXQJ10dAshpmBs5b4+jzha8DqtSQOQi
2sxzD26LeZ0vrrNPlJtk5sExg02JJdQHUME41uz7O5hnfkZqGzykAxFnKzqdxGyUSlOQgsCGVZhG
0wUz6TZcAUpgH5BYD7Q+rA0Z5m4596MSawChHUDUuC39MxbzJHDJe08nG36i5D7WbPrL13PBTMBo
RN4/iuLqBFKCpCaqjR/v7yLNz/KcSPORbqx/VJrQRxOKUTjI5dfUp4uSYtdp4rA6kxjCs7tkl4Ba
uOf08VFa1V2rNHIuKOQvGgleElzC1mrv3F2XQR6gtgVw74cwh+zW/L1C2rrj4gywJXS4+TdYOJsN
ByL4DARXtNNm5axRCpa49KV1QAp58W9Lw2KtSZzsRXF3tEGIr97oSuvyh3JrX6bPcHJv0WadlDza
soNR3zjAhUks7IZsEMPddfzMSeNhogGneVMFh4eqbVeJudZJXdhDFOADK574OrEf6WXnGtofvM1u
3ZE7Mb67F5gT3wWMF04+J+MSZ1U8OjWOfzhdLIWhDyUpfC8GdW49Kd9b8iE0vt3qbADRSJr7yXdf
LKN+H8+97XtFgUMKL9Wi+wIPFZy0q06Qw5FXVwBmFr3Twb4eHYeDCjRGvgM3p1AznlI4NEI7d3KW
ANDfo8oQA+evE/zk7TU+E8xQJU6abeS2Q/j6nPW5jOVypnhyCwaEGVu532G8nwaGxfHJNY/zI+ep
Ymjbi8AxpuCoNGzJ65VIpSJFChZOTCZve0S4CEnR/poI3vneGKHamfDyJVRTryAdJ0IbMN5ygD2G
Wh36JVMiWE9KNShPWcFdWnnZFDumc1IyIxbhe7jdylAz7L+g4rRrlBdupBbuBzK5SWZllwwInglw
Voa5H4NMolo2E0vzzUsJzud4lfJKwXkKyT4zA1qNP4UepzYxpxgh7lb+x0zkHKBfKdmwumMBTTw1
35h7XD6DfqDw8XoXnvhoZljhfLHan9kNBKSze2WMHCxAMkV0cq1AmCci/AYn8xdeWxUwbMKlV+Wc
dlXaAhTnuH6Dlsi9YsXdwbvEX8KEm2+7N9TUPaV68tHx4HY6N5/FS7D6ZPODvphUAaHXysmhOMXg
IAMQ25r47JdaJHPirueMQa0umBsxU78BL6VaA3zL78uFi/QAMt4/8AyFCBPGgsD8qC4Sk0dYW2CB
Qntk0CYGSGz4K63TZB0Gd9BJNtdl6DvAvyKL8zy9pkCTw94jXe0lxPRDZzbokqR3ezDlM8E2pZVN
fVbsbGWtz38/LAC0q0LS+HB4U6ITnBTZbX87Y8jJszQuwU2/65aZGfqhcWrNYt5ehMoMqozG4kCf
uUtr3s2SvbI7ApBFr0qaaDd7uC5kG5whvyaGYleEvqraegvBC7FX4+24tKzIClpOMW+n4pCNqr91
Ai5mAcN8sQ/sYGk334Z6pECfDb45uOPnziBu34vhKfVDr3/2giAXrik7r4fQw6X5oBwZ0KwTThJg
fcfq7q/jW/fggTnOKn2g6CdpHzw5x2kX/nd3NhM8CAsnwhe27qkNedRWQG79TeKmCD0VK25Fn3wZ
bZr4Gev/tRl7aEMi+PuZDgjLXhuOCxXgMT08Z7rPCfonHmqk1Ys3P/tx42JejaY0Q1+UO9CThDYJ
ti9UDxAsHdke/fQsq99BipxTwP/ARZG4OXmsxGXn2aC+IzX8Ci8zjL6gkRJSUyTRBcEc1EAW+W2Q
ha0wMiQyz52zAwCNOZkWzuk6bQPd5MNIHf1KrJw3vj2mRTbRv4cBN4vIe8EDRO/VijNKIV6oNZRg
O7PzC3SsL/lZXyaNPgm9t9TFdIto7MWPhHoUrXfP/accxmJo3OCWuWSZY+Xx14VBStTicID8fSfH
4YRTbBVeBiuZyqO1JVY8hpVJfs19QPR3NkIQIiUWUHkbHHAwpKtIWP1TBGPZuPCtCL10H7ZwnBBS
zoXYR4VvJn78ytcuSI7eM/Mq5EeOYl2rSEaziS08GxwElEGCl3bb7s/pZuBGihnrPxEfj8VywbLX
AJrigITPz0p50gu1MRPYQ/c7AcGlPE3frNtnrdnRnorve8p9IN7P361eVPoEv7RCechEO8y9R9Yu
+9kZNa6ugcvDIIEXPxmGTDsi3fHcI46+5qTJ6qUlBI3wu2/IDtvqoglCNj0rTzmd92ATqo6Pbv+5
odzBP91+aeqw39AoW4Lx1La/siQUK/aXMm6D2xblm/Vw+Y7aoSt6N00o3OSEHk0tE8EZLM3FeOBk
6uUzubl5rhGadCGKNrnSb0jwjPru21WF5+aACjFEx9jkNRXyhKO9FVSgu002AvtCvnsJggjr1RqK
U4rTqqEsgCt++5cYxIsP6YSKlJWuOvIrlCRCHipRoAX3kaRAPyFBIEpGAfLWBglP/UWcJwrjohh+
oRrqqEL/89N/3BO0XU3fIiRW7pE4U+elmgcGzyALZeAocnsuDah91L/Dt/Z4u+QSzGZCo1laf1yz
m1JG+wDCrtekp40CKGJC3UHARgridFQXIxS/UpnDLjkqKbU0TB8e/UZYXl42hhJiSI7G/TEGfDNv
1w7Dk0PFiSov6cj9GnNzphDgJKg5k/0GWzJHEbH4rqA9yVdCLd3HtDD1R2QSZSHYTEfI38kpOQSc
LEveSaThPH3FW6rL6oqabodyEMlYXrkMc8iMEOCFcI160ZMdsfCjEQqbXy5cfOo1JPqUeXpvaXyf
BtDS0IVoD9d7XMkouS8jEtYlxYVVd9UifIdFwws26gO9rZhwsCanuUCXJ2+18zDetZgy6S2dgQH+
7tGJ6zb/kt/nsNNN9cP4dG98xuCSEUtdlktOZCNzVWOpDUJPfC2U1ncdJ+UmjrhdARO6ym5LDAFX
4l7HqxQniy7GFPj/B23OkN3GUAPRQzKR00aUOn09SGS0ISV7wMvGb/AQmNVNcRU9ueFdrgj3KN6g
glKOnYhuaZQU+4m04X0ZG973wxBdMRBNIM4KKuTTpUmuuCFwk5vzBJls30BZj+RKoI/JT1Dg9qLA
L0OGszoZ1buWErr9LpJwiosM5v9akhCqEBrM1OQVR0Z/bSqIYLIt09dum1uB9KnPhhoAoYsL02nk
j8vTEUDxfl4UG3IY0zV1ciL8QDmpLTnMfFxCIABFLJYGI61OTEhiPuM9SgXWA7b9o0c262NaK9bO
bvHSjdVxlnCR5thDXunhcK9BwG139YWluF9gE+S5qL423Ws3Rs9GzIx3t1lUxHdewzTb9a5Xb/fy
wvGwzkEVYC7hA+UIRrqU28ubl8mKEctvcstyM5ve0IvC5mPcfsXcHMjXk0z78Cctkz1sw2mewQeG
yZLajuWgABdLEBOvB9AWzrewizxLsZivsf0ahxQNIwfOdx7VPHQiLMZ1BGrn/KSsiklPvAQEOzJI
qZqU+y//VCiAZG/pLOR6/FY6Ink65ngE21ZLQyY1Mi1n1RaLexhMC7NOwf+FO06bYEwq3xUbNROn
JAmdyvqlOYWR8iYTnhqV0xgwWmqiz8T9yO95iDu40RV8dnaINzcjx4447VcnOwhLEojMFkZigICP
DR9FcFKc4zfWUQJUCR7WS5b8PQlqpTI+ScCXouct5XLGdH60vHV8l/Sj+x+hC5iAoGW5jY9zEB8D
6emFqXWjqz7X56qPwsmoZ5afPj8KY4zB97VTM9uGqtHtOV0QjT4QJ/uypkc76NWUgEtTP47y7PUr
NUABP7dj6vaykYkMOs8ZvyIfZ/4t6IljVUtITV+8dLYymf8Gu7tErA/hxvD3UVVU0s3MEJQZS6RZ
SEHib23VIt3jWBEuHfCLcdoQnEoYtnImpmH2uc8QwP1pnOokkHJCzPh0R+jNRyxuW2sAdpijWDji
ulzKMwqSuJgWWWKSXbI7UtlIDZpTkOX9XYexgV6vl+gbaxnYdw3gKPPFkHglP6iiuRVcyw/D0HZu
bLMOH7BR2PCOWY0F20VNvhpDZTmwxD7wAyb9OxoVROUjOdrPyFgX+xVHhphznduOC5UtpljGlpGQ
rW+5q5FjmWbM7Bmh23clcRQIbX8NNm9tz9zJmLpK1mzhO3XDRek+jITVyK07vT2LC7whEF7tMBRr
O/uTrgSykll0P2TvSG1z/9X+/oavFK20b/Ut9WSSvzuYBaBVEIQRttre6LQaiJR1PtCCvcmi8z/S
XiCtYby+SKvm9hUT8xYZ3XsXsGuJxmSvjOf6YFIOebZuzM8PifGwCgNa5egIx4vd6wzUW+I+op/X
8cgInzq07u6VH7+bhlbMwK363c/EKwYzHvmMypx7XIJO9D6J/Wshho1nU4iEj8y88Zz6DtFB36KI
VLg2GRfQxBZZpDiYsDe/kLFRDOJ/ezcl+MwUQ3+wn73FOuRAzPekJ60qFOewGBacUj8wdvgvr/PK
pZkocfQH3GwgJ4ZHucXieSy+3kHqVZzJAneJJi+OUU7xu0FyZwD3DI5RwtBdK9bHyUPxazexleYj
+GqZlA087tLdFIpnGT5S8c72DNqdY308qsBXliarjq9SYCEeXNuC5nj7bD5GefnjeJe+mmtAdlt9
OmHgZYhJ13suyO5U7Xw3O+KteH8o61JWD2NJtwtSoKiZonpzTxrTBsjkVC9KuHldjsZ8UFsh5K//
ThyLIasMqagjRhMhI6Pr0QyOAnkP5l52NZFfVpe/k88ptRdv5NXiRoVwIBQCokVhFf24VsS8MkE/
F58hhxN3SmKv+EaBw7CNnoWfJTOVATMFzc4InCbRSHLZupqHUx+p1uWSr86BPNgIVFGhX42WqXGX
hNm1qpfVTght4PsZH5Rxit2Na7hkoqbe/xgFQPn3KRPCDXJgJxSQa23P8dl3MIxBvYqDlipYE/e+
Y5vMk1N4/TctD1JGY+QFIKpB43aHU4/RxP4OVb//v0qYRxkzjo69hzLWaAP4CKLMdLBGLvNpa+Yq
7MHWkyxY53VIat9QHOX3PgtcOpcx8M+nDc5/8eNlTz+Q7Z0/MdnF7l8pIIghvShjAD0hg78ZTamb
lqblgqv2uhE2QBq0xi26doRi48KwgyGezxF3i5MxVIR1hj7Vl6HZSU2Iemuf1CdkzvJ4bhCaqRt8
cQrp6kH8/yk3gNEr1RqCI8Vs5/ZMaFNQtAAw4SelI0nVc7sAyIseIr389y7mN2F+nC4Vh41TJ/gy
wnnXaWjhi+S5dF5QRekgaHtzVoGEpOKGUCYfLQx50cfjjijDmEIsaxX/xebiiPAud55kkSC5uaFX
xHbcHHLybKtYxb2f9uhPGyctnlp11UGur9kcfcwC7A6BDWz5ssUa/V2kfNSB5fP4tuKU4de53FWB
meKxGls9e0pShEdDig30ydCUIOIaoAoU++tgzXkwSjNJsilBN9Q0/W0GSELAqs6RhoTpZpWyJFqY
aRUGG/jEqUqK9xladfy4J6pch3hqDcUxbyXdm9thiBxkbKAZK4heYT6RSwlbPjgJHgy//SUCIP9p
MWV2/ceRvNqx/VUMKxHGARbI5zOD1pSibXI2khNWk6y2FYq+ub+mUiAZXSCo6BLkCMXNz+vB7y1l
6/rbcVwVIFcWnAajZgbO2QlI0UV/ikZ/C8T31538mlVLIn/l95ohL2dP7cgc9EczG44rEBUwXL/K
Gewd09NKWmbO8Tlre3ZivVvPGKZBACqo0Nz4F6/6V+e18HbA91oJbNeqFaTBfi89i9fhEfzQWoge
0ZMWkk/hkzYsDMVFuaWddbrtzy8STCBH8zBTS0gP0/16V4guywhhA++e/KW7qaY1zOu8D20HzLo7
oEcT1wq8J7TagGi2LLxHzLl8U/bxl5tSDjpTse0vS2KHSaq8wzlnxbI93uo604fI9xo7BwVAZAJx
epYdoYriPJFVxPwATJbBknYeyP2JLWKTLfPJal5nHzE/XY+/q4grW6SrUHatJDVBwfFVzs9mu+m6
x5Ebaw1K2HPatfttU2Jq5cycwmJi1pk9oSCakrp0w5KyVY3NlnhvTvcuY1aUM0yVo/qyLkKR+jYn
d27qERGzZDs+0hwKljoOkaa4qP4D+iU6bAtuZrB2coMhLJO/LBEioojV2sWlTPBak+XFHnS0iCYQ
Kpj48mDZZSSUrffIVsoBrmodFZZBVjyMKggFOT19yS/Te9C3eiWzpLMfupmyxNhYe2LTtCIQQynN
ITMdW3RSZpiYa9R92tEN/SXyLGBiKuhdA6uC9mYPTEqvZoSYeprksH3tvavDWq8Lo3V8grb6bVkI
weRW0+odlGcVnOYMyi9thNVfGmNXANOeBfcoq62uEkmZ7FJK/QfnWyS21F1gkGhPyL6E7GGwSOHf
E0kneb7Rx8k3bTsMBURKUfg7IGvG7+aqFQC8+hwNp8PX16mq9huSA4XnTXOMAToWtrwp7IZfnrTu
pDZHeTN3dROmchecDPoufw5ugihS3F82EuOQcOBVgz8yKVJ/WUzCDBHyQB1a1kvW4S0KBqMbeVZT
IM6or8UZ8+PLIsAAqXGDVpLt+gF2JsMNlYhEiaeJAYN8qjoGiuGvN4+2q3ZGKOpj2glz6LRMAEPF
gmUsVxs761/9PvEF7d2RLBAXLcZJsHdyHHFsIQRIqPZ/s93+i7l6n+LLdAlbD+XWQNVA39ZuMHSb
mgf68MiduJe1D9lSTl4F0KD2xMt+VP3WaajoTxVTgHYWX71gY8lQ2oT8Y0E0r/VaLRoIEwVLJLoP
0/nIEswMNHtpCHW+ubbYl0ytHElKW7aePLo7xUHq0JVzDj8rNTI1HVbFGD4SL77BS5CagrtCg1H+
q9ExlV39I2y7NYcJBQZceArqT11R0esLlzqTW4+jzPxxjf/DwdwWdhsPTDKliD2JWLx8+MwZnaLQ
TAa/96xzeuefohfVSOugIZ/zx/qTKSxNOyeGO7c7XS/5EPXtxFILXTYPDYRRIBzVhL9MjLu1VTLI
VGx5Ok+bayck7iRxKAZw73Y1MfHIozWmbC9cSW6wKIGF8Vc/VMnUHEDd/wXOVZ3M1UigQg4Lj2b8
9WY563xN3hFM5fwQODNlJmoHbPYyY5isEiShDRDts1RCDh22vnH1311FEvv4xG6SUuGvHw1uboGT
23o6rjCrf19XU9uuZvFqmB/hV/QvZ4Vgjz6pi/qlsGU51kA/L0H9DFYHUrRZ3ehfPQQI6SBA7GTf
rkq90ZpRFC6qAOTuOndH2ON6VV6j9iFbm01Uj+Pv+RYtznRM2f7Wo060CwGk6teLvVj/TQXkJhyR
LXIsIr6owKl5FUqIi5TAf2XOCCKZIT3EZGhlcwEDkT65u3MpBdjlzAhSVAivJJIxMBK2K5ccSusJ
SsHNe/tijQZAF3l7KsLZR8olSlXVPCG4qjHitcgFjcS02lSKCkKX5gWMoOW0kQjiiU00Hvs5x8Wu
aFMN4eHagBDltHanw5c1ADJh/ReOPdZN0FTedBdyypZtf7VQYcflLiBtfj9vuyOEfz2fxFK7fSnZ
lP/73MpDY25FYtro76LxN7ofEKKU1whfX9iic2JCBYiCXcZAC8nZ1H7q9XC4dsZ+PHLn0nJWgV70
4Kag8DJU2iUvXz7pEiIGH/3xWYCtOSTMiPGgjFrXi/YqN9MX3tZj57oYJwxM6wUPQCubxQoJAJtZ
e6zS/4heqI+M8E7+d0kiddgecNTbbRv8OUrmb/xt3/z3VFmGDI6NU6OErBgxyYb5uIJRQQNfRHH0
NolFqnhd2ujMQbMG3lAEoaopgj3wgaXgfkle1Pwz2Z5rvQL1jDD7wgblnaaF1gRpoW1o3rfYeh/f
iIFRTU0I4FLV8BYTkMbBBLkPlGQUFIO0w/UzT/cYqe0T+TL419G1s0JJVWnhfzwFVfoGH398h12f
gDjlthOz6rpRD1NZf3AQV5Vh21FqWqf1vyTS4SqiD5uyisfIaZjzBmiZjTVP9VDUruWwtC0e6tLr
jhVL12CVtrxzJX9bnRHijPMu6GN2OTdpDyHC+6Wg6TPyBr8x6V2L/lj3Rk+qt13do7/1PwsWvyAC
GRF8VMHULySkqBmc+nL7Wg2evGlt/AAMEV6nmFHA7LFdQ7xgu9ZXkh5DFwiVU/EwC2JqZRodH9Cl
r3sVrYJocq+IAAMDdpv6tVr5g7/jfu9E2mP0zbk89zeptOEU8BfrHQzq5nSgG3FxTEVw5R44vY+9
7djZBizOnahkVQFBx4lQBZqlDPKp/5+9D3B2/mqD7uDZSxxFkRJRctkefx/KwjPDgn4ZrG06aLwH
jMjPIV2XbGzjlSakdjj45v5Jj1Srjp9RUpeVbmfLqmfLnWTNVWYAZkBi9cSEx/s4KVHBunYk77NE
zKs/S5+pIROFHaiW/wCh7BSnPg4iMamaNf7TH1nhVzj/a0d+DQcF9ahoWSmXOmYYtXEYh4uCrtBW
a5GL9HdUdoaSDG4HLZv6e7fVqd5kot4AWcKCzwgc9u9VqHx1Z79gmmcJ3ryHhNFUKwpXA/Ge6TVE
T8+JepU/a/7eZNj0SNUsQz8S3qFNZe14z85muHOerDGsIVSfwY0zLq6xh/r4W2K7UT4qRR2P/TrO
iiGlQTT9TnMpYOMb2nZQdBDSGHjJDGdaaRreVfkHeSj9ds4XTxoYJ5/ZDlpypaBxgupZ4E7uRMdr
2QbrfgNfLCzXQmZkfuitg/fPR6EIZn2lg2wox7ELJbHcjsQrEg/LQGymlL7T1GoKWONAok3MnZnn
Pr9VRAp2wTqwF1/WS8RHuaiSyPz4iHptoRqksbiufMDyLsqvd3cmCV5sFpyUkpOGX2T2GWQ0+a+D
rw3X91+q3hGYvC+jKAgmPqnBg0xtZIOFEtxbrvjiSO5lppKR4w2Oj7ocWjbMn82nSOYam0ZC6vJ9
BcDkpmnbu3wY/eHVEBEfUXHVFNp5iGZIqE5fnuyBTsc4Qtoip+1vGI8CdakmYVpZjhTOnSgrQRjh
kiVO/6Q42c1kQJQ1+OAHCn0ECYg3po5nR+qjDKMb1uk0OHgTv5Ds4LEu9Md6bQ3eKUg9PE01k1jM
X5MCII5hVXssyTxMZAfB2XL351ZsZydkxaUsjyuBy3eJZSVou/wcgb2+FKEjs2vKZc4RQh+3709a
afu6hVt/t5K22gqngqMcOXV85K6+gmXWrmNdwYy8G751J3CZ1Jl7Wq0sq0s5phiJoqwgEi1bRkDW
ryaHllqSRojAptry4hMPTxPs2wl6PIZA13YJCGUYc4hUDPWvTsq4dfaUCxX4ZNAbU7nZy6nA95IM
sLgvb3xvahp6DmgPxJDWfGB6t9U1ZhvJP16kCnLSIAc4Z4keiV928UbzxIlGSpkgFOxLf7jGE8+W
+9gSVwyNCFyhuwPpa7WJTbN3yRAWilSo3wW5q8Nh91gaGBJ54/xngjTpayrmL+FOupfIN+RIxJAM
hvubKgAqu7PdvTZHzne5KXzNnemU8u4WRBHSGPv0vOvdxf1rE76dyyajkyOtJ4kR+4pQwAUmRrmp
DP8/sp6p7Qbn4Zx1dWxxnDGT2+g3xHYGicgzRFu6UvyWHXgYHUzvtQ0v3UX9ysNqpw1FXXQjZqJI
vMsibvyAiyplK3GaBXvi3+FA90m4tNg7UZEOtUbbGo5vjr6BmrxSy0EDTrL44Z0PRjMBykFtoDW4
CAo+CLlqNKP/VnHCfFYrtCdkR+75MDV+0tZ5Nq6ppj/kZnCbNkEPPa9O84OzzyntwddUN8m6jLl6
1fNVafwXpqI4qXRuQzSdePS7Yh/MawN51nTRlvD6Fny8to1ocJ+ji6MM1gvjud7Xx5nQz43o/OSd
O7lICzXNU8tKDXr2yjWjpOS9N12L0lgJi77j2EHBl7Jf6gfkNcRIIhuoSUcLyV/KnXp+OK9AqAit
9Ri9Hb7Kd7LXSrnfsXf/BAfLzoL4Oqf7uJE8SbQXzL9LmPNhRgtRSI7yCt+teWY/y+Ai+wLK0u1L
oGMegf0unv9OWj2y8HRJ42QrVia8Dc1l3B1PcKDIxwSEFPxNG1iZuNkAeK+J4YG5BMrwMo0OnyGY
z06OINMod7pyejlYYTKujKCzSjcopikclhXAiiuac4VSXGfMNXs5AZVEYlUJp092/gZigCUik29f
h7xFjfX5KYIKnukJF2PaL9B29+R4vh5Hs4K6Lnb8z9P99omvd08jZDEqbVc5DGTVkwn/pECal0wJ
+vWiAzk8XrgbRK11xcpbxQ4K24RYrDoagReMXOj+lEJoYPoEq96tRD3fF2BOTUxwISnXJ4Q5fv1S
YH5C+Ub/RlytLeCFhex1P+69IPBn83KKs4i7xgmUrZ7SviKej8GFrb4InTZ/uibXYNUIMN03z6Hd
ZReF8T0MnwEg+J41JIHTLVKYY65UN4W1o6LufqbSfvVA4E5jiR+U40DFfJinSn2K5b96TEw1Hljr
5++E6PZibHGLMonYPp4LPuceFSxLl99vAv4SNITGRnHcV1uIz+OnZNLyV5H+7pikJuO4fEQisCUS
Og/nUDUwauB+W/yi7bkG1Sx1akc0AMCAY4UU87poXGu8ulk2OsmAnZ0rxwe2C4GF31J7Z3JhEGD8
8BKGokmVEXFeiay+53aVFxpnLFM+G3/q8Z1DrM2l3bACYJGIjfZJFF7yxtBHRDVRLlMdfpxWlB39
1EXWDoCtlHUFlt36YW3DNbTJtJqcRFDlCJv9rESComHx2spbDOeKS+GAhYQ5LikbAG0MAt7hL7Gj
wlUlyFbbAlBLJJ+iysKjvcToNAyPLc2Bt8p/4b7FiGfH4yjZDyCCIqFvOn4cZ03gKRjVlfA+rFpd
4TKvFwOtrexHPeQ0yaWDnLJuqIjAtEHFts4ewUC6KTUVaU7lqWV//GOhcEuasVlqJKDH72ozdqyE
LxBk4xwvGz5hZzCSF8y/1wrREp72QMcPFTzZC+N9Rqy1fxGWLvxpNyUbRbWv/asuVIyjYFRcW4tp
Q1vPso79Qdb57W/r9U1HpmCZKEHsJJxYuA1h5891hCrVNWivUlOgHIkzbXCMgeZ1S9YHeC7RMoJ5
Nc/AlT12Uk47ZPuCnZyFHGVFjBPKUlWMAKQUlIdasC4Q7J/g070E/3hWDEefA86CgImxVNmTcw4y
lfNro1Lf9MdeQGYWwnsPApyK0EIDL3fQM9jFCOmeactY6jTbzfFC+xJb8sRrjm9JlGgpNA5jVkqy
y2H8JAa6hGwBLckRHFTHAmYQEvpJKZmGLPPKvD4C7DUwpxF/vNSbhQESeAdlSlhwxfVcPujYGtr7
IJ1nINEV2pzC5xrMReg0Z3ScEzRy6JCjUrh66iyhpHDh3Mr3kzVS+72Y26nvf32jEMyXXqPrsboh
8tMPITaDokDzG1JmHs1gV1n9W6B/B95UJq5hfyPWC/0995h/X75PwRzeMTAM0mOEXJMATV0qHMvi
hLZplvoRKZ4spcn5/bp9v9kDuy80v1mOL92gvJMlkFLYAnh/E4Ue/zxobCLN1YISQszgh1VyzDlm
VACLHOFDRP1ILvpLidn19X6bDPDqbrQkThgN/up5Cpzb1zrHiXlY4Y4Kju/8bzyfEJQ7MPapDTR0
BQBbxlz459Rp6x4NnJH2gkEAJkisOGVHaKvqARqZC+QKajsdpqdtl18U7TrXx39QedfMabDYip2R
e/1kQGruY8L3ePxB+JpEbkxCx+bM2dPSImJ26rzoL1muPSmDoLEbE1EwR05a4DcH7t2R2EEnz+qI
5TLUFqIiWNTUAlPkzKt02I4OJ8m0XoF3kk3pW97dw5FHA5whM0yqPOPaAXLguZLmswlIcaua7msP
jpx0AicRNTTPm32UXrVQJPdswvSHNlNXKJSOUfco2JxHOjQiMjk2WBaecXahazr6BsJl8cve23NC
5QYk6WAdcvD1miFfi2JrFWlUm3xTtZwMea0Rt7yIt6RMlbDuvbGncVFJgSGSPs8E0ByZ73Tz4Rhe
uY3CU5NVVfodn7BU1zDQhLvLjeJbsU2pow1U1bqBRKUGtA3LzhbAJL/SkpaE2IgUk21mBU4tqj++
576S4yH2acFn63oJHfNKJXnuN/4jSBGp0GoQ5DyzSmdBuFCLBvZ9G1pscThnQ71yMPRBErl0nEvS
nOgPco2oHeUyYMPOPX4vSrPxip/PPGAKlutOy6nD+FPkagmzbDx+bZ3bMtlqHiCOXpfGOGp0pMR/
P9LPB1r8SywoAKA5TJngTG6eqSiG29XGPyx5EZRwc0vFJysEZXEKkobHQKHIcin6JkJ3cueGebog
AlZXiweP2RNgmMkcLC6uP5lH416yyWwDpn66EcpNZEHFUvYF3O44crG1/hq87oPsXoQdZjWYCpuf
X2o2XS0TMv1T1lrKwAo6r8td8aRuhUTejh4mPTmRKKLqJhNO232vqAuCVM668v7KdK+OchZOtk4C
Yck12U12UDkikNQo5nl/gCJpVr2cfQLLRxUVYzhUjqGLVky0srBBMcCV6fDiXGgepmnkasDkHuRc
Kyy5zBMiYBnijlZKEwkfLiPvj95xNTHmGA2uP19a7wBxcZEXRKPcURMwOcxXmrp51ec3S51NCMd6
4BPhX2tw4bGaMpu3+R6lIjMZyvKGeoLO9j0gjA66SZ7ENwGp0i9drf7+ZbTVDr4nvJRnxlmnKQbV
efIdwBZbJ0R/USA/VYzn4f/hUYTyfyChl9H4JOINmsnZKQt1Hw2mTVzbv0cGLFnPh5t6kQsio+kM
efYMxey5IAaIIAOVkqNYxXyJNldxgAzDQRfcNK6OS70Q5XU32ThAtzLOxy0RrUAV5APOdqGVc5pg
tRGyUI1C0SMfaPCRHqq3yHsJQsW7bl/J0rZV6o6KeEIyWYS7z8yvzQTBFwYKdgzy2fdMzTkWfC08
PyENdM63lkiIomOvbOKjEB/Viv3YgpFBjwav9/QBA+mtvKUOa5jxfproGOJfECQB1e4vHdgb3dNm
bqVZl3BWFqiz8Zs+a3e7+ZvIYzJaZzcfFeFvNephPdImufpUSBadtbFVpI+MEACp0zvPEe9sLSsZ
Rrnh/vke4CZJhQzdLUVmNNMSCClbpp/7Zprmm+0Anf0BoPXtzDctL/x9HZfvdqKuqWLu1J7Gjj1a
okE+2jcerdvy5X/t3UkKcbIkUzWlpOIdd8CigYh2jjn5fqeZCbSk+fpg7DfOR6XY07mN1YHgrF2x
+z0jQ4sazuL11/erk7KrEEo1dveGUQdvEymNc+7ZfMNo68RRH+3AF+mtH81p6E1V6TwOLATGZBab
OFnoLHJrA2OBZsLVw1Z24ie/0uGSw3xgC2dPXRgNYnhSrU2RbBwqcDSsThNktNB5KBabcf11bVoE
rmyyJnVkqljZw7ul0gXvZKKW1hZNYHR00Mht7eqbNQQv60OWXWaAMXEtKWQrsgDyvDjQIkCh+sk+
UxMZ/JQVBM/8QuQLOaqUmenYn5iWEa/7ucNxHKYKSh/A2N8hhqrB9t1MbfiKxrv3cpNMCHz9bRXn
FgWOV2MpywUgrYV6IWyL1x+2upAatLFeSI0gfj9GXu+5fTvAa72vj96m5fEgzXtsH4aaWMNpAB14
nWnU3hj8O89jYsTmAWwvrDqjnko9808H7yVIrZj+IjGnOqtLaJtKswdC7/+boxqRrfowT+aMFx54
yMmDjkkateBpACMJHQZP2zJggZWJCDl4At0N5Dlenqfd6EB1zkyHOtVcl/O9wxb8oQ32yGL6ur+r
3YawfY5m3YqKhbVlP6ladDYk1YfVHdgHzQ671Qy/Lfg56EeTOkO4IaNvAeFR5TxbHwBLouw2QG+S
yw0dPyuTFIya+tNNqZuUlprHyJBbPcGwdpPmbEs1Ec+WRB2yU5NlpXnwfdwJeqDpjUrYE3XYdRog
sN95pYYHUxmSjvNwfOmf7eljC7ODmHy6ZV49B/QWYr8f2+EalaUAyu5xae6goQ4YR7qAzCHLSz8z
WxK4gQPEU6XmlAerW3BbjMM1fy3C57sTwv5CEmmtE0eVDtwPLyWKw69Ji4TfgOztzdVi0Eg2v+IN
r0ngFY7cyeNtWlED9nu3o0TJsk/lzrUm861Hg4p7TIndp5PtVEt1PEXrcIqN3j6ZqXR1RC7/35Sn
Q41bBzMAHIrwvha+hzdEjsS8wi7gKz8c9UsRmO+vuHxxLU3j9bm5Znx393sRAKlJK9AbjPTP8ssu
n4+Df0O/23SNtemG6R+BoUCT3ZoFgbl8XD1NGB9GUlEev4tpMQ0xY5V7Xj7UtfLh2MGxa9pU0u8r
RX7Sh8TYc62ZtwPa/Czo37bndb1/aGLgtaCxDcA2Vsgs6Mc1lTEKPq3VmfksvKsZsihU46/EdxeX
bf6g//sacp0HImGAEqWKEQyDBNVo513+a9Buzxbdv+k90F8grso/uP4p3IDH4R7V6VP0ifeYw3Cq
DTMZr+5OBodGIY92inDUeC3MHlBfwvO4pY6wtMJsPy86D+ZVT17TP7Y0U7x5kikUY9IWHboIGgkH
KWC+gTh+6LwoKVLQrKzFYVDGCreaHOCBSB7lT512oNQnwnqmdZGJthykuQSX8RlHZMHT9yDX6VHT
e6WfV7G1Mefs7/PnBsQUAiVatLmlB/y172Hb/ilMYFUIaKwE+xXy9oFUlY62BTWrtDvOyn2FrRIG
PzGXv1UVfkRmBiEnvo7lERVCVUUSJ0IKu1+XbW6bw4l8E8MCkAi6vMGUYjeoRiBPUh709L4HaM/A
CvRQ8WXnyECK8JqOIpuG4dbx6uv0TUaxSskhMKqVCR9CUKkrG/BG3qqXc1gSin64szhJFSM0PmmX
wg2Ev+O2eiDRJ25u2RxJIgMPuD4UBwdIe0jdqbIUD9u+l6P4PSqDFkbCr9Ca/zpAooXbEx4B8nhN
raX8t+SduEXY0g1AZUriwoH77gw0Bo0+4aRy9u2wBwLVXSjWB3ew3YWbiT/JDWcMD/fk4O5cnTwk
O8bsb+vMk1J7hU6T3QC+40YhJZhRYG2Ee6iE2SHmFPpafE8pn6sMKbwT42JcXtuMZvDFdwRFm7UW
jfXCZRNQVELeoV8IhVzLp+5DAJw1SFXEVsvH00rMrq3Huw3UnQr9t6c5f7bIPZ2fPM3PazbbmIAG
8getvheJ4kuyXNPwu2iR1KU9iYVd28zJKwPig4SXRU/GreLtswkOlKDIb1Dr9hI51N+euIYQDGdt
M8Xxo5S/nWaC/lt0AXdgof2p0xXvj3jtKFja14U0aZ6sW60m3u6+efPedAuX6ezB9Xp/CsRckjSq
hNCKDBnxX4wlPCv5JlAHyJ4Dd4ipK7LULcfC6dTFy1bL8PTWEtPnOW59NC5yNaaay56LEG1EhdmW
6Ng8RgwKFu0jqYc6kYtTkofv2gI+seKE/JPWk8YuPgCWivhTHUdMZJ8x6Jpp2Dmen4zkgYu8+wGS
npsiK2APwGrjnJcbUXmigcDo1DnmG3KbtQ2D0jCLIBpfmWuKHI/HElnj7XkP5Vi7nLVU3r2qN3jp
HkQ5Mr/cit2k0xjLsMQFxtEOXILayYqnhLPJWWT3KMV6xLjofLcC3uaN2CQvshwff870PocBKC8F
n77THrf1nP1dIGuclnqJ3uqk+PVxW8Lt+l/FZl4X8sMgnk0dDHejtqtdeEGC9WA3RFl9H/2XP7Aq
lXtE3xOiufo2Ug+g6NDojQ1V1DL8PEgF4vrBoMpuWpzskFHNJj456IY9Z6ydJ4ZBcujPvbfW4jp/
rtquzhJT7Gw1Gprhb+XVhszUUcgrAl3ukgRBmjCL/Fv5KAH95DnlTIHWm2tmaej4j9iJU4KHcZKR
sefZqUZQ2FyuLH4UZYhVUTsRCkO/QaSYE7XtWdJZ/84q9tn3RBEZiyyPgksgezwxKGs0CeGY5Slx
nt4ryWN/uA/X7NxBcmXebY71oC/i6t7mZrOvbkWIK3+qoQjykkxeleg5TX+xDVdqFJ1BFW/tOnag
E/cQ7f/vNFq73EsJVPrlXjOCuZl2W9FwCwN2ompWY+hkuJSg23RnSVN6UxxKMzDBwqTwxemmXE/D
1oRNGT9mOa8hJkck8PtwIol+8IZisq+kZQtZ+jMfCoDWyOwROmx1kRwEYL9j66deETmk/ybfEYBz
ZjPH485RSiUmYYqdvkbFXMLSFJUPgsoIvST6YqozxLXVoRZXz4W1G4hzDhqH3pb5svbhsxO2G4VT
wPrtwWYawfrzXBY45hD9B9HzD+zvR4nbc/PTRTNKAaLf+UkkU7NmT9O+QNFUzly5a6zkngyDYF28
NJJRrH3DjpFW2gIH+JrMySjCPwJNXyh+C06503HjJJLKglX4FwK5WQ3QM2N7OxRh2Mr84GAGZYUq
aMzSkQbTnmpVjPRXdQai1AP581L4N6Ug4TsBulswotuv9K6G4vlCTiXCv/uQ8Xi48ZB266CQ7S5q
1wNGjNZ4b6+IjJG5eh1sbPp42IyE7hWGXTQbYi9m3UF5UMzHUPfNJsP3BnhIs7SfnOjr4ShMwTvg
wsiK0V+VSb4FtGfQaC/i+UEwWFeaCipY2fHUgN8PjNs/OcRWumFZxRY7gi3MOQaNYmU7sgbtPXLf
domdM74wJf5V0AZhAh+HK2QiZq77HyQTgCq/ro1j96f0bi+9NY0uxHK9IiHo9EGarILB4RKxv5PP
yCaW8+sDsA87ao+Z/vIJT62xAyiUkhak/tMj7QODFlJQzUxdAtCaPnlRZ39FCLEIwtuvE5uvzahp
dlY4cfdRX+uU9uNoAlsA0MqrH/9+z1fB/Lr8/nKglS/ZEiIYQ2V2R00quVHbS7DtfVbxbaCeXnhX
l8lz7Awg1t3rl029iyoKSvz7yGjH6Eo55/oB94xeOhCvvyGpdz75tNN4lhqn9h7cJ0/jvq6N3dtG
oE2pIV3V531sbWvXaeRxB69lKU+8YzCjr77VqRKRrLgU41NxNaZzhhHx66Q/UnyFXOOl2w0HiTwA
ABcIP40TCB177uKQsZMoW+K/VrmMSqHEPRxKUuICuqQAM9RfRhZUBJOomleJjtwkvbV16EYxPC1J
HAZnQ14KfbMW1NPnXJKO64sUC5q6BpLNJD/71Yfh553SELe63G6SEcduz79dUAdrfgrGe4vcZIuE
5VOWNgl1X+608QEaYnPA0ad1yJtU8o1ATzzL9T7NSBmLQZkawW+A4cIdM1bAknKu9oNQ9Zks+TLy
aQtlxEPgnnt7kQnKMPgtPozgc4PmVcg3HlaxdX90IPC8SWstApdkLVt+CXphg7a8VL/UiEmiZEo9
hhZ9YqcUtPM9jfRR/b6ZVS+CCZlM94aSsBjYzYG7ieOlfNhbeCn9VohbZHJO+x44cYm2czT87ye1
BSvHEZZC9rhCO09MAyV6B7XbQbLgDTeQqCBqHRS8DzyUNs1E0Qi5FRLn5mgLsDaqG/V+hvWwSBjg
hYewjDBgN7YgjpbHDTtqwltHB1AFhdvN9ZUFo6XAmW/0kw01O+ZuKx8fR/wxpqMAUAccCYiMKnTw
3UdLVDFyZR+hZEJaymJVNridQJ+4svKRJjYeflYAV7O9/LG2/+py4QEhKFkHMXcs8hkttNzxozJ5
noYiQJA8JCCoPwJtzJsvf4CIheXzwGpGLSC9jUDit8ObJ8FZYgjrQrxBc0PNCQu1SmuSVpqwtN9Q
KhU5qWny5NfN7yrQwoYzWO0U9YxNCmMrx/ckvzujCCyB90kUvQWJmP77NyLHEYghWUEFNW8Dh5I+
oDUYi3BbNiFYFfhfNcCLagC2b5IkA1RCrR4QjYTJ6S6oMRsT0JSVFt3msLZcZVp0PRekrpq73Q1s
WWX0po7NEsMw2YNWdRpx622VgHad1WoUY12yoc7NkThrNvUWsrs64MHOpYJxs/LCV8aY8dq+Nuz1
LcQPbVRLhDpdpiLNMD3XgCcNYDpIlKUKgVpJAtgxUz/0NdodWo6VOiiJ2LDxOD0ewelZovzf64/1
py/+xQU0yTN0ub9OgxNaNNvS5iKar7sK3CU6vAMvFtbA6rgheDZQ315eFggURHVflWE0u46BoOaJ
zcsGE9OfW241Y2gU9UGe9G0Cd4B/6+0MtwzKFAjzjRE67kGNsgFSON0c2xpvlA8+tS/5BEf7AHLZ
KyqBrlx0OdsCgdnc5t6wt5Gs9cByWI5Xgb4FPUxne7VFGw2xN9DwpqRuu19GEuAo9EErbaB2/jK4
yDkDT1BBK8eRM79Lr00ug7fHdn6CQ4SKD9KEY8yIDhDcY2H4KEdyF5FWfW7oy7wLLm+kzRMqpYFU
6LmXnm5epnNqYz8SWRUKh4LYDevBOaj/UBTPtGwgI8ZxWsDU5WdkMsA9qw3zDKOd8LJeO9kRasXV
WGFqNc+1TnC+C1Xs8OokjLFZ5TLQ+2PkUYYnsGQNBpjw/a1f1IXDrJBiVeGIUNAi/hpmNMyOBook
1PEk8fF8ev7PIWXyGk5IUwYXVTWbI/Y1mfWu7EGbkP8gaBzsADjcgq3qz2vQewchGeqTW7zIrYHv
3vjDgMTc4adYsM57DHxlvIq/Bzvq/LZfZj5S9/5nOcQE2lpNev5PNgchpw2f7T0INoEzg44pmhrx
MgjWlAAKMVxvFv6V8VLP7SpUIl5VZglAoNkLAsVNe7jJ9zlfWxFalc+StJoqOdl+6oiLIp2onIiu
fJSXjSSUF9tP7L8YYJbUi9zKyPcZVAMTMgqoyiqyTvMN2qtyYOXnfzd9KJKsFuB9DTvWmAO2b534
PbtlzlikvJtpigK6CqqO/GnbuMtLB5i2gnLpGG2kW5Ntx9+FK3ngITJ0SatP0olA2V9ZCz9LKexy
o+3zRlr0hREfDwzykOlfWjpNTluQXuw74bsN8Uf6mrHHpl7IJCGwGs3ueXfuqVlIQaQgBF3Tvv3T
mgVAeCJivkoUfEdJ6IurfWnzaAElson+PzfR6rV6DsF6MhGRsHLCJNNG7QyRJDSFbIUJ7EjTL84m
IdKPIwhD0rkEBahYpYtDjtygZT/t4q5ula1/8lFsxwjBaYFVdjT2Wn5UvyQ49xp83zYmzsdtm4Bs
4RE4uOLR/W94XzERObuJUCqOXD3iNcjUCshyNXKWMycsyr6uJrav0Lb1AdijH0hgLCUsPSyYNf1D
CwQYgOCO4ZVlkm3loH1no3+jwiczAGl/3KSfOUmD5rdazi0uYa/4PRkXoygfp6Bw3oilCj9nLUPQ
QZuPxAc4m6j2RSpp2XdCACdnKQA5u7KdEUlJqLvWHfWxG1FHeVJY+oTqlWTY5ATqm+FEGUlglrW8
8Bl9pLTICYzVNLv2wL+5uWRkEdxpMAH+IVJJSVsjHjQsMsbNiBE5jy2kZPTppVBGwREOQrjTw/7E
4pKAzpY8iXxixI27KKMkHNd/4WuAkUJ0+MJyOnvuFI5rPgbXMVoFeJ0Tovacdd68CBYcGibH1rKf
D2b3bfnKAKPpWRBalGZ5OLM8OP9j9/uCJTkibGvDAMJtCy+cRI7GLw017Qka+ivQyykOWfPkrhel
QhfJDqfZ5bIv2VK2LRbrgWgiK9poicYmtdoOcr4Y1oEGUHFUcoUC/46DUvQYMCTSKlYSnWWtk547
WPBOnaE7Vg1SfZfhjf2VRS5OenUXDmMVyj2l7FqDt0F93KYjuaTFORR3fmbG5ccPlJdTdD2YjTUp
8EJutWKKJKkh1eOdDsFpBbP1enpuQsl/Vb5F6gMkIRklBRbtMbLmWqAhCgFBPA3vmz3IQEtVTOnZ
YTZIibq56FZoab+fRC1BW69C+Lmqz6YhTouiNSrRVCQQ1JJUUFfdZBtwF88uk++mBQp+dUouCtgl
3OtP3T77z3GGggLv3lhTKb+hT8fESuPDlRF+Rd3c9/8O9267XLEzzA4wTJmJcn6KvMx5NOtTGnL+
eIeWOH3chgdVlPQXeI1sjqX9t8/2QEGkS7w8bq1PU35m10wcPanEJaZ9C0JUkgp8UPyiI4H3DPmM
5iVkzAIqWYhHNYta/nzWI/X87cS6CIEIz3s/nSIwtGmBg0pYJsmbCraxFX4dtoiMSHhr0a+juYRL
Z37kqGjDgGEFTlkqqtbTcR51ebaGMru6ssIK6lUQPHHdlRa4074LDdkZSnjkxM82LZt9t8ulebRq
BB0gcozUPd1Km7mKfgN7D3EjeXgIU9d0aUia9xZNiMeXFGdcwcYjhdWM8RnkFAhF34AgqztsoLaI
E3lCtcLviec4EY5CkdOKDhk+N73LpW84hq+8ZT+msqHHlAiY5sNqaL0PLrD+t9iAuNq27qaYCZE5
X4shLUTJ9ocxSSQ3KMcVjicJ+RrSWmIzG5taAJP8cueowhP/VXa7UlHBMl6v//vw1Ks7nM97MKTA
bPvITYpaiNkZXAC+pjvv6YKPQD40wUp3WA/2dniC+UQ6ssVqSQwVgyW5BqCamdbjzdAi95JVQMJr
avXwEBGNC7M+XRdAhrmJ/jpr6flobrddbeDCotAc+OY/SHugOfxgDUhxLXMaB3OXmkpOUSWco0MD
2tJXKEhinWYvebuGZbrn5JexYdStbVtwEom3g2WF2I3E8Ob7GSwxzevNL2cCrXXWGea0PbYGOAJ2
IT7TkkpVHnJ2TCwiOkfe+3nuOzbAhw8MFZ7X1JW3TUemBtYValg4mQLvOOMqk4k+GiQG0/IrAKr3
A5UdSuIJ6QGbs+J+hQUc19F1w9E/UYxNZ1Tc6VambzM9Stf9+iE5KThlbIummMskz1bjykVlOYUq
n/sAblgCEPEgkugq61BtICSKFO2QpyVgYo4pf31VR60qQySecudiYSUpREt18SBQdWdfQ2k9idB1
yWmxYZsJk3TqL2u2352VZ+rqEubyTpL5SHS/5gtCOycM/W1eQPQXuNmwS9M3Rz/HB1bYCwMfN/uw
dnFQqfyUgm7hiEV5leH9d9uvU2X7jlk9gJbHNZMQoY5QHlzUU6/Qk56yKWyPhu6dg65l3DMFeYXL
LjeKGSsjTKn3ODtE+AEczFF7gVWXWVmIHFPnRjHyGu62ktzIJ3qebVh5rl0yJdw/yTJbQ/zIFv31
8rsQpm8b1Y9/Yu6muCPYCbZhbEFtaQmmHGg+az2POWS47wM2hewLp+zb4GcgN5Ni9Y3lJL4DGjgE
rHIYzTaw7Ip/9Fq8QFYdPRP/UZMHvZ7CDGhv9hDfhwRPfTU/0r2zIQN6HhfA6fU7hWJND3S4sDl4
dYHhX5Cjenh3SglhlaAUyd3h8IFxkgQo9AkDpjxTKxo2fCjtZ/gJSbbGgZzRbUZgq+5aND1H6Nn5
OxmhQM9YSzSqcnJkJdqjtOfm8FzQ6VaDsIu0ZSvVuh4BXAZh4IszPwIomUmlS4hGtMCTMVg01K9s
sVkIu7z4pTdwm4wc7ka853wTUvcL7Z93J1dSIxGdtR5uuiFGMFY4SxyBaYynkdOhOnPIYmNTP5at
/ym4O27HbIS5quvrLUcmS5/2yq4H4+E6I6Z3xDHj022gWR0GYKKXoFeFYcPaUOzra3EKnoA5m8pH
5quZu3cxy0tsqbdaN/gxcFOcwtWbLaVcBulRiLvxspSWNx+7vJa1xAFe5X/yUPXyUSXExd3zpr/M
U2vYDg9t8L28IHRwV3kddHKhutAZQ6Sr7QBIJaPEqxEbxHZI0wLNPqihU3eNZPeekhj80TSpbHcf
7Q3kqjjTyOmk5UyKWIqCbSXtvTQ1VvXY23OIRgrt4S6maYoOFvlaBkNcTYorX4RKjb/oSYvq0ZBQ
XcVxWcKXTEKtfffVtBVi4rmdlkfsuJFoDL1Ew9qxtB0oAY2CQ0QsNXnfr6xb2WpYgJt0UjcHfNTo
LzZMyCu+Dw+NsURYwTPDpJzi0Gfbb6kZ/JTOgsPzFeengy7vH4bleqTu5zn9J9/xpFA5EZAErHKk
qQ4kk4ran+ckLH/M6a0AlbpU77IyaY9yez0uVFjrc0FB92qiN7B3+rbNqGWcvrIdKZNNgwJoc1Po
XgMzslR+L/dIP9qmiO57KcZwwE63w2Pi0knP2j+OeIupGm6MPG2D33Zx24iHX8Hm9uja9VnxL0ES
eL4ghQqIlYElSGXcu9FAblY6ZTNqBoSXuEoRBUv5ZLfuZPyQO53jCPA6qVYx1ohRTtwgdbQgNfqh
HGHFwoZkjsZCSYdQ7VfLzMt1rMGp9I7vAd+aduv+95jmpytaPGSTp8at+BMsJy3Rtu+sfVQhPN7D
UEH0mKrXO8dHjQh4Xcvg58AmAjnwN5eazvtHkC70OW5lcjBUjzNvO/Ywo/UdMljcubpQePIEgXhJ
cDD/t3Zwn1DTApXMqgzFm8DrCtg7UDe43NJYyxt9r13f1rIULiRgfq8yBy6Ox7jTFwfDfXh4LpQR
9Nr+HEpYiXVq9HZUtBP3sftIRszByvy6rcmP90Sl3nbj9Nlr8dvW0HsPpigFSufi7rKvKEOHud3A
m5BOIQoYb3yg9P+p1mbxy3rnL50ebln7fs0ApLTQ0hhF3pq79opjYxG2KnMQw0xCc2AB/4k3lhFb
Fb+ZaqIfykWcLUB7pHLkHcuVEmEl3mJaHSv0DeCCvMmisLm0jPD08K4cRAqpPYYBe9jtmWkMkJtq
9aRd4ZA5th03uoEyhsOHFKU/2XzRuzhV+Ns6qPZ5LyUHD+/TFvYbtTcUwQWegurk+g8EUaVu4EgS
WOTr+gza0BYjt2k5BG143N3mSUjDAu8v1CKLTFkl+HuXWwsF2QXUyWBrQNsr6CmAYJ0uBZYrSurn
DVfNTRdp3k8XABpJeXHKcA8259GCt5BIh0bwx9lEhOXulR5aAlx/Pt+xuEZGajaFaGGNTnau9svS
MUmfA3NOaaMY/IYs1S2X0LcLBZgSlIkizY+hIZPGEqaWnmKxIDbzLZMgZh07K+QHVmYlwGAEzbp5
NJDD1MPll0BT2ip1H2RdEdfqrO/sKTkv4gAY2eHAWrtQQ72yMvj0p1/1esTGhu6MueXKPvGT9EtZ
5X2bphkyox9I5ctxNaNbCoPnWTQFcS30X+R0D4LhSwvNB2Zpypu9w4+f1YW0Jb9RYzdAIPvpcHjq
32Sb1nz9VY4fMJ/z82goDoPtyN6y3UAbmN1QmYoK+82y5D+/FkWpOo23LRMAA+mroEbMO30DGRSS
LI0NBt+lZMkEMGcHKLZpHwURzALmjpaIfHVAAXTvcYrckxp3ySAoH6Q+SAisUgG5ipVi4GJFl1Ck
HyrZmvfUZYaGQ9a7UJx8sM2fWBMf9pdcIgEJHBeffv+udtiD9cStxB/WIfrpW8d/Yv6k3lixIFVM
3XerkZHum6APJ35wJ1Sf7Dc3cyxCnFBvCgyWjZRv7jkykwgoaBKAfMIO6xwwFEDOX6/MjWfKXt6V
jOfZ/DoBS+88lQiWI5fZvjx3fwX4uj6mXUHMXn9CItBoFhIuipXo5J3J2od+3R4MKiKsYHKTW+b8
WvBa7g04abLJCsq7y99vecs31mJVKT0eHrgLk51886ywtHCfPdGJu2fMXeLyp49as+NdpAQ6KTqU
Y5rFlYNZKIjSGplcemkZadEHQ1HbBi/q+lmHhmHBuHd7Wuoyijx4rBlohoefc5dfq6jBXJEnTTjz
Pm7QlfoGzAXQsPv4NObDxcB84WYkQF0IPNdhSDa5Z1gYWlVtko76tuNMkoRftrVIZlf607zRwrHU
OLaNCNbKQ2ma36bkQI4g7qfA3OdBGoCDKMb2mvS3U/AWbnqJqiVMpdrqQFN12aX+SPHAwlKoZIAo
E+L2/Nljrv7UR5wtGJsEtVl9+UR1JzK5UIXTK4xuyDBeR9IlVQN0SIsHLiNznVtesSYjwpaSSin9
E18nTjihZQaHMRQiBt/Cyckt+Zsm5xgT+jYrZGSAd5kYOhmjYBIIFbqR5T7L3h88mckOCKqRtc5d
qdm0AlLxmmvIUddew0ffNoR82tFqVQnPYvnbpm+rxlSUpyO/+ML5ovIjcpugMcTTPnTtX7I+VX24
kMlWzT4gKO55BoWSAufX3a2C0GsMnCoTzbmVgDD5VU1g2i6pmu+FXU+sSUlJccv5GT5Njfcf5UQO
xLcw60SiUXy20b20oWUsFcmZ04EE3jir3AP6YNWvCtAKrVFc1TXqCOlzAtocaq1sWj1/9+x96nIz
zsgztG/xByE9AqVmlySjOL2hOsJFWLn7suOrlLSjo7urogGZLky1h2wO5wmrVggq1yNg+xQNw50v
UWSYOceXKAGSjSe3LmWdWisgLv3UjyQkiWt1IPcln0GPF5gP15VXT37o2Hvf/Qda2GrdTWXH+XqO
Zk4njrh/L1jYvK+7FNHAdAyFbn96Bkwbxg9u1Y6J0swOfmeMaoDvmwIIW3RZ4wdEEfaGggy2n9T4
Bi7S369WSrw4MQ4rNnbKS1Cos5QuaUx58UXn2zpXQhrYwoCFyMRHxaqZR3DIVeOorg9WOCxr/jfs
QVVlXNI0bWzVtns8WKwaxjVPANfQopiCO7j+HggcOdJC/YolUtRf8ZRgxlFqYnQchCihOe2oNODW
HvrIBC1NIv9YxoR6BY8KXeKoLvG8AbTu7di63r4XRHNHsG7hWpcWuG/EI3HFumeDeRpMzR/BSe7M
7znx26FgN6+HtOUollZV+5HPsAbRS3AjZBzB03jT8ghAlSHBUXTq/cLVa5tEmHVXzCbQjCwliLMT
EJgd8G5hO9Sbe6EE2n2JwNlyiYrWnW9e5Iy5h4OSgNTZzZuI23+bOc324zZwYubXx52wpTvbzlEf
Lb38+6sMn5IkPr3/CgHi8dKp4Xye2PgjMeC0YDJoB1FdrSp7JQ6sDXsEAmn1NiKh6/nDtAD93ruU
dSS4dTQ2NRnFQngKTcyrBalmxN1geIs5ZwzpbSlyzNgagW2ih2mnCND6cAx6bHUeJpUlQz2duQ9r
/nly6NBZlDwj5gRAAJY1tFxFNcwzhNgZMGpClPwzILNvg/cMmpdbMJ1JYzojGgwwwc9cMZQnVQfE
wDpso/1DTH5rz1H+ev9h5/0VXDodEFa33RO6u3/ucnlRtjOZZGG8zpbfSepSQmUCGQlncKEUf5Ti
2cVgkyktBsSmlKqsiPDBurD18TJUxd41v2XbNMU9qKJ8UhbDHg5VdSe8biecs4zvj0Z4+K1hPN2C
HwBAGDvYaByOk1/7XsVNnXfaeGqrVdXlsBSO2dWzn/VPf7nBY0sbPy2K0+PmCEKKWQlYUNitNi2I
qqG2iYB8JCmjxJuHH3xZ2/VYR+Qm39ZpRk0SO+uhq3SaW/FIHFUFycF7P6XYFHrl5KPxR/3M4+8D
RiieBmcVU7sMftZR0TNGh1zw+1PJIYBtWWtzsrNItCAKlDkAJBwlRjtH3TzFHJi86ksnf+iHlPzK
89tMzfSO9VudeI3tOxiLZcam3Zkjt5mwTXSP8ZNjwwb4e59Cz9bSWmO87whzPakBvlwSB91YGPwu
MdTP8AT8jnsKK3q7gnUoll+2iklcYxjhkTXZNBDp/VL+gQCHssa+DexN2pp78Dj9Ts8CrU1VcmvF
q9YMqnF9Z0nP6F3hzJIKQ7oyw8VBzp3MM9HGaKIvxdiSwkRmDyjgkh6IZQcq3MkryEXYzJioMgnc
URKi8WzQDdksbZLgLVDoM1X+wPUupzFoNe0/jVFT6vJfQQ5Z5yOWwQ+dnuCM3OgaISjxve3KOCic
8DSem2OQt6VHmC/09QXbx8UHnyx8qE+7e37D0TmUyNqM4sBT30I0tEPNkTEnoGOOPBWUh/K7DsjD
Kp2LlAk9DrMhfANHLPvdXa+CIM7j0JHnyPFDq18PU4l+nVldUTX/dQNx6tCVAU3Hgnq1LRzEUU5L
W8DQy/jMzmbWhSxNK7ZAul9dOCqFxpyCxSWGWg9+SR7SCfI0y1DumWFhkjECkVPQs762FEUAGGgA
R8HC2Pj9tmyeINaFtq4vk5psZZl3mmW10p4JU/sKAZvQZDM71ViaJjdi942AUuXMI6PmUP1P0UKD
L2sewBJrNSJwme/TaVdutsJ1mqkmFfjH6qMBdIHjwWNfL6iTXwTgTcQPNnm6erkaZl8UlEcgAz3y
a9NIxaEWqK7TRzNiVkJpqSfWg/JiYu9H729zlvIEjqKdkZu3m/mwmwp/HmkPLzPa8BTpQjdb9Ame
tcuBOlZnFH8lq05qSpn3g3gvy8JnxyHO5egmzWq4bIDodZJ3mk86OFYdMk12ooknplpJvkPLm5fj
lmrZ0gQb5sRfLGrIcjKc2CPRdQRPiZdxDWSQ0/PiFvBdamB4uRX88HSnIz/93QpaVqVzmKA4DH1K
XTbdF87yUxEn3xzfDrhvboqtXbBLVyLfeiaxJzX0rlnKoedAGqLqNxELJQgSFQosj+heYASd3AAC
Vi98Q+5roti1McFIVyUKlIcpG+tt+i75zjFFj/pAzd8Io85gANh34JwZWCZc+2SEMrySEmbps1hd
BPJ1GLw8yZ9kEW3m81YHmbmZW73fdE/9+3xBy/9eUgtRpi+C/djeMtqASj07L9cDcgNPt8WIqJpq
QHNMR4NQ5HGItnH0aY2f8cC93DrWz4sSjoz1SP5H13LTjmV5BZgRGH0bp3kh24g2oU35tVnl24bS
19df+cffNZTHvBNqHuD0xcnLnS/kf5bscnH9kvpdy7g8QXG+Ex1qlvHBH2hnM7RnFRhyAVoE1iQf
AeY2g6kk+yf1+y+Tm1X+5DomOQZXGOWWTRxJB7aEsw1abDypt6qxytRIrwZ13pwE4yzHpez48CJ/
P4rj3v19EhOZlE0NrCk99UTILT0C32AXGyjhXs3CX4XeA0akA2e8CogBKb6XqfmQDZiAuqRHxPNw
Ga3tmaVCxEd+v5tbEXu8zvSpVCbjoeOM1mGyQ7GQqarUDKFkxUwiAghqcfDnfJZmgTmHmQFvQbGG
4JBD12haYwr9lYbZoyx8Y7POpJpIZEHYexQ1WEIWTH/v1hCDIv4xTFGvNwXFvws0vAWU6D5JbSVj
0cS7iABVofDK2WxTAfoC+Udf5SX6O0e4oDDDQQaBfazUbfyLghFjJTkKxjh4/uzrMC27hhmOs+Xx
xO4yfocScVMMnXBbHdQ/jRgKUWNF2CsKWDmNVKMPq4EdRe64ikNHlOjm8FbXdBJU2RVkj5NsPyuX
lBXta1/n13YkkM1e5jJgrGStv64rV765iOL8UdSwpqdYUcGRP7tD8ZAG+5qAQmKTUCeVKaLhDYIk
I7//nIScdBiUjfD3uKSL5r9CPqeWqWIVdLv5EQjfqewem8zOZLgNxZW9IkbwQDe5+Jxuc1ibr9Zp
UQmpHIG0lAwqWX8lo8/NZzgmwN2CELhLsxSLQ7E6GulKRiSGz55WxJyBrZwjdjrOWsh9FQte8qMP
/byUM5r7nQxANNYJ346WZ4EX4ExXVtC4gziyIFTV/nO+/biFz5dDrHbsqFCpTGXSqXk/lZsloaeD
kabogtkF0zgXZCCwCQublTCMA0YMd0VESdcl3yBGBSofboBMp98jNm1sdcwME0VxpgYOXe2NzK4+
poky7hLBFfJ3nlr+HHtimjTAHo9FKI+wGZlmPDY/n/Pzx3iZUrYTPR9fSjhwfCkmSMMBlqmP8dv5
lLX0QM1LJ1BPD4UIPunITQoRiyen6JPwIGIHlYQ3W2phbJdJjiuwRr469zO5oDBkYD+KuuCadI+q
Z2yFoydzQ+W23pJytpcDtuC/k7woFfC64dwz0SCZKn8It3sVxscwohEGOMu61jP9X5LYGdV19HlX
ZtD2CJHoul3C9bC/OPzeLEbanuzyaOhxj/87zEzAARlhDDzVqlPHO5dr+vhxAc1JMSZu7gAEbgON
QjHMmCCWRXkKlQOcU1EWSXi0TG/hfbtzlmV5zxqFt8GOny47c0pOXsZSzhAUB6yxyD3FtOQi6E6a
x4398hinRrOfiBsuMoROGQqlfofcZZ2brDO+aPcbsx3XxGwTKOsjkjCa2tBiwS0kw8YrbK4ipYV0
ROWLPSpVqi8hQMwcDcVeYc4yNfphZvDFJnWeik0wStdSWY39W43DNgiQIqjbbdAw0Tmf9wr6sSWi
2PVpLNnILuTFX7P76+g1SfoqiPmYu2qLx9kUQm4KSFOin4XCThSbgUTePFDVyq2Yg01iMPgQBDp5
uHm/wodDKsAEFielsUAXn5eQcoPCcNjby1nBb3KSzhWwPIV43ICbBzhEHkpbp3le/bsSyOcDhOfn
AKlg+Rnv2xTl7FNlf9yPwWWLEHmfIiXd59gE9fAAZCEwqGhdL4F5ZXaSzKy3E+dNIXLAsjySLGT9
wjfbo279Loiae4FJ55++RVzjPHcLegAB+QLLAk3PB5yS8UK/tGCLkUAMQMC0rYoI+ZzdxI1nxETr
cU3HDO1HFs1+kutDElyfiKT5TsnJV1l90y3Gsghk/8qSVZvXKYQt7C58pr5lYMtc3ZJzmxZF7MCh
T+b1izBx2M85yNuCRsvlmP4aUXDugrRh/q84DIDZU6kymUUYH1u1T64Ht6mHwx+dsyUbFhrjpubA
I40FwH5gtQ7hTkev4TEitOv5CDFaoKp6p/q4pYfJWDfYDhlQVO3AmpErmdOl4YFP55qY+m+ta1A8
gHmbnw1h7JeIkHet9fPoNyFNpQIZvoCfYt69/+WpztC1kaivzimLFWICrEA+mbDi1qT+DXyD27dH
1pL0M9BhDAENQ33EGpSk1OmarD76reJYEHXPqAS16kPfP93Pfh0LzxFRhDSHyqd7ZU6KGXfs34jT
jMa/YFu/vJy+J1MpP6F8ROaNqdsCnTJAZm9Zu3sAMRRhU8kwnQyhjcBKl6GerYKq79l3/rsu3sjc
W7zXMhNC+Asa9eGK0asB7OmgCSEKUL/MurIEI756/g+CmzrHHNyjE0R10ptzU+5m69ox7nV9RIaa
iEqaChQTV5kkwtTkkNQkjzxg09IIA1AIuRq7haVrafxGbt9rgFnmr9+8lVi4Scp6++peZAmHmUM7
AwJaFkAR/xiq5u08nrQYAw/0/ChtQJHW9++u5H/oQFrd4fz9rrT6kItUjgyqs4ocU5RMvOLFzD3G
ruuOki83+PcNS0mM7qeQ1/K62GTsZnQkDZONap2PfpAg/fTztpDX+mNhB5bS4ox2/Rprihui9Scj
a1FoB1a4CKiZHBM5QI2HjNNzHPN31WFpR+EzzMWntjgaAOBKJvYPhf4d3twYTzwi0zfPcsjAlt2n
lubFCMZNiC2pq3e6NkJvsGxhYG2JC9Sh4P3diviwSyn1cCqXF/fJmuEMwfSRN3r7EcduINvyoUZ+
nceo6GoTnUJ+sfVZFPtTILMFNOuptw07lSKRTYL9BfK+hTZN7RSzE/64FavPM1zaBooBhrUJbQqE
kZBm+cc1FFeTGknt3cKWYYLlQNW/hIK/t8zSMTW/YSzWqqEXr60/BfKfw4K4IQDZgGeCapM7XhJD
B8mBpTJ3Ara53Su3vzti3yH+cIE85i9+geXHZfL9/VGBpe6aYJD+3UyXH6MqJBWsMGLXZUNDpibL
UUye5BCdwcXoav6mGgum2KfSLyu4hpHgJ2PySBkV3f+/8B2qPHM46Q2n2u+VEhvc5xJ4nnlBXcY+
N1D7UWT43hpcM4kfMbbMrgZjdWSYMcRWI3VBmdQVgvvefYbiNynbPRUPnVRMaOuZ9hUfHsRb3pDy
I3ZDXVmAfV9+r3eqhVIxr5O1wbQPhEJ5qp27h+Xwnfaq5iDEX8E4LVeiVWyNBght6Or3ktz1QRfz
cj7OjjrqE/gR5Li3V7c6s5veS+pl/NECGatQyxvAZYHdFznswOKgYYkRNWw+3NSMycm2zjT0nxNd
Pv2lmCv1giKBXcy5EkTTf2+JjmNxTzs5lvPGFo9kifUKB/0ueHO3b+TRz/QtqE13vOScUHuh79Bh
kKt+3K3dPjm/3RIwaf+hTrJ09nYru8+TlcWmMp5IadGESCpwpi/m3HmtLOR7oeqYmjDLxNzwGsXV
BkpzNA+uluak4c16sBc1EzxkOw+K9DZRBpsmCvuNomWcDPuMcVT057aMcrtpbmsuVHya3WAeX5Ux
fsSL0w6Igdc5XtdcgZLdE0aVj/NHnBfB0SR/Jm1lM9w6umc24kxev5RavsRZkUcrVEUmePvSstuB
e4Qk7NiTeXvI1qZrfc5+LTaKTRkam4AHb72G3B7inArRhJO72ZP+RwTyQqtzaj75HVXsNox8asAh
/BcHE8vdxGK5xoYbalqoNH5wiWVJzXcGf4HcT6dV8hpBwCO9giZLyL3rt/17bVFXXzi36lPSt9sS
qFcT+jMP7ZDMhXLliNdujTy7mwbtJfNpcSriW6eg3WygeUdqrHtsI/zxTzKsbajCSyiRmFa3cLOo
lp57rLqX1qEJgQeJ8BlIJwGs6YJifKA8FVgsZblfYWPEyS82aeS+RO5OxqIhc/Blxu7yET+28Nmg
uEc4EjxI1yBkYpQvhDCMS4TAW8r+DqXCOee7MOkOdESHpva+SY/Sz/g8o38rjcFUuClv6tzlnua0
WxEt3c7s1S4PNU9UuV2gvVt5FpuR0LJP7aYT8p+P5W1o4xlNe6bYaP7b/i7+qWEVrAwhV+mYuyZq
ULHc6nrgW6ARPhc1OwYMWm2mdvXuw/HKRgyqAOm7dUkWpWiQFrkYL9b2XPchOJTPJNMFK/OiYEXz
fjClL8EnYZg8HfaZfyNXYkArz3FcDQv/abOyuw53PLKfnrhcdCfbYHwhm4f3ydcXHFaYpkTjKVzC
wxNqU+J924CtyGE1VRd/RDzE3J6uBLzZ5rMvmf7aOQyVccyMrTu9t7XrLqKbEeCgVZI2aJmOGjfp
TtvkfNYQkX6G4KMIj5Mm49WvEZEDr/5Qhdt8CPkjLdwBsQFQPqzZ6Q1CXnIxoxtGw2MJVgya+H3/
EwiguYzKW/7BV8Ky0FJpxHLZT1qr5BCkGXpMeQw2q1dP89l7fF+dwka3dz3/NH/l7DEj2AiHfBss
/43RlhIMpdYiiqfeuOVFlPPBo81K/7fDwuWHAVFoEhchbrP7phtLTk3zGtgsbQNOnZ5KqrEaR5pu
eluy/PM3bszDOqmGqy/kLt5HE1aaXv3wGJk+6Pteyn/p9nZAc6UmT4PhVpYmLH9D3DxSVaHlkRAv
6hIIfVPjnnnmqMS6rKpBbxYTfHCIrIb1yK57+JT3Hl8kRHG4bRja6hqKjjYjEErfCLBh9H+naO8B
WOEr4xPXvq/9NcInm6M5+nFAHi/gQPjDabXPVAyZuf0JWRvnzP3CVok3WKpFUkXSWFD+Xhe3Ds3K
z2xCAIz2K8a5S9RMzuYl72LtvLDLEwoSxUV0SeqRPU6KPW543S/zifDzumDwrhRzOc26XTJjF/U+
vgyDY63eUFL+N/wzR5WNrj5s04T+fJde1Cq7eOfRTEmcWrsnK/UgwpdA0K6dKgTFGJYAdCoWyKuw
CGpE1teSq9BfSqySuhzqWnMjmoGJbdDE/3ce11P/w8lGbm5rWTcBLcd8ZAX+wsOngvivhyAF2LKu
8sPpKsVwckwvfFBsI4bc8N1Pmz0QLAo9rkgqSRzkkA9LlSiNKPoBdPWv4NGtQ+YAgIA1gXUd4Li8
hzEo6wXQ3YGUcPX4zzaXnwMK7Xj2QFeePghX4GjhedRPzo21utXGl5NvbACm9NMxlw8rl2OSrGtO
j7gzSmaMWPWzBAmW+lPmQOgtGqL1oczEc1qrIat0s6ggXIkca+uegk8P7Eipy6lmBXxYBjDN62zB
oAtKr9cm6isNBoV3K2GA2Zh8XoOMrkrIw8OTnNLKyxXAA4FzcO7ySrqo29DoNztWgTYtUb5Igi4c
fDEXQrn3H872oS8uuP1pDO9/hjifs14BguhiypZH8YIJA4+6z+BErSS1wXyQc6hzODisti50MQEQ
JSYVJrVk68BqJ4KY6pQhetd6d2ZSCmwbmU5e/TSGPBC0K3kFkEzq1zZt5mQDKs7g/XoxatiVa5yV
+3/0+u/EtMfJBGfo4fVL77zmIi/4V+DODqbPWr1tJY5lGBKF3r/5m8o0rAWrdZmSvzRgk4HCRW1P
f1gVElBYxK9gLFzSVJu6wKSZElo4osvsbxZlC3FSoOz+Us7+osJklVTn71EmsmvJ9RTl1GTnEgxd
GUIZYW9VHx30JYtulVPSaTtfwPAnEGNZZGYbanzaBCvzpK0hFriML55dX9urKTJlpeHmfftFOFCQ
5qmIjdFhjSaO8BjQM5YYeXRubu+v0wB1Udd9Be1HBNJr6+MLk8/+IKIOqeXIls0ACuBMEcwNxN8S
uzQgFbcTCFISsoizDMvaPhsEnHF54vodTJYOaun8E8Hw6X939370fLS4KWMndl1xi59p3jWPHL2e
LcFex49WbQ4bi0ct7874ZU0jPWkcfLhOckHyAi2rmYCG0Ram5cNb2Jnu7UWB0TluX8TL80dDpkSq
/U6jAO4b+ZFZTfX/sWCtAlg+n9Z86qDss9a8d0laD6o4ocR8BcK2+rrbsOo11TGiD1GnXXnPEi4P
9M2EqBtiJ1Kkmxvoj4VJRo4GBdg7VoPv8z7u875s9kPlgwY/iFcz2R6X9gvkZeyUdggjTe1ib/P2
ACE0pFvQroe2XwbTKmF2JZ0UTmPjazB2Kxu/5Lt41MHW81ba+4dUYp8Lq03hhN8mwWBgJHTjxML6
7VzSgkO/JjLMkovZQ0BBI6bAXMIMqNud2zP167UxeCyM13Hsb7ZaO8DvVNC2ocTpBxZBgZq2EjxS
nrQwDRERVaed/J/LTmyW+sRZX+AxUQ7phFmc3fp1ma1tXcZrca6gTZNpQifXOoNIF2pj31YSKNJ1
YibTs8Bx1dbBLSFrHIMnt6RuOAKSHdkP7VJIg8uM+Fig1lDBZBeyxFuappvEdw8vnycLJhC4Uo/z
uz+GbhjFASyl+G9ucEswmh39Pk+itfyoYqK72ey/9lOtMkG303tCUnPIVYwdwGl1XhioGCriDxp9
IjDmJRKwH1LpbwOkC32jJWI9Bnk/KVGHTk/JGyaSfd+oQrqJARfzqEpCCfV+W7yXI/lvq5yNYWC+
zi5/zLVpUB5gfgqTDk8dHEwdZ0NWU1qPebd1QNmCiEXw6BEiSjLLz3nnvcfU9ifQhjrtqU7xtvEC
sm7UrJ1AYg2IlSLXz0TlVQDTQ+YvsHrnEiwuigheYjttVcZKTAKtf8p05SKOMFfUAzQfB6NS2vJW
/cG+jlH0YiEbmTI8kJbaW0CrCRBJvCEwo1uifdCK1pMLTX/pAQO1lQI1fug2/2sme+oj6XyAVyqL
kI1dIQx1mSd6t/AvzFX0UtH8kruWjKT06ns/cj6J/8X1oNdIGN3GFBOJX9vVfIURtNW2RCREywF5
/6JvH4mEQyxcdr9E9Jo8IvHB6XoDLrXkgOraWTQVop5zhaWyrTjpopovK8Tz8aUgoh99BpZ29kvP
yGcs+mubKLOuGXRkr9X7ZsX64T6+EIneE2f14Bb4J1tC23ATNQh/ywZnSXoOg1hbw+ooa6fG5jyy
ACJZtBTSeeRc05DBHFsumpqGnd+s6g6aXrOb5+Olrw80sBuiwM21pV+Y9YQTMK/Tg8aLNviHDEdX
IUa9LXVt/1QEj8D3Th/br6D/IyAKYsdWSlSduq5GZGJWcCX2f2LbFiCOn7NfQbzPs3pQ618otTmg
pU+8N/UtTGiQD5EEFxaBpAqwAP1xb5hJ+VjDGm0MeJHC5Db32hVq7o5GL2XbjeLgR2OEAKZInm9R
FOPeMEbL0n4+rOd/AigsK34JBtDXwMn4r+z3JnGAUkuV+/L2BdFJtIaTeq+gZZ7NTLY0G8LLHO79
esCR7jX0v+faYY9X0HCJbWH0+RqSr9kU3T3xF8xR9S7p9rwI053zuMnvQn27/PzHjeE5k1HdB4YC
Mcdr80RMdnA7cYPl4v+8KXyoWFiJl5Hc6MI8AlzyDIIN57KwWMennKWOdblOIOOfUbbyej2ombJE
nls30e/cAcmLt/dLcaWoyHlGmSdVF6OnEVUmfIummA6ycebhKjr7+QRvbf0SYrdw9sIi+NSgU9+R
u3sDUQf+kPysttBavcvugaNMSQ+x1RoJMAhBBqsV27QTT0RTzfALj7uV+J/6rwmDUqSllQmg/cjv
Piyl8Wu4i5l0jk11ZCI1V5gl1RGEHDl37vGfS1voZkk/ZALeLSkHXjSBYwfkiMl6s7vzP0XRHZfM
ynQIYNw7Ig+ncwblcT5nmrQXkexlWmF1QcbbVndRr+qdjac/DuYSYA8JHqln3e6YtKIxQOmD5MN5
1et3wF6Q6N37nWX5a9Dd6Nbcm1PNvbKfq+6LO2fwD4q0XA4t3lbaSNH/m7Di0NpKIb/D6BvjEMcg
sLNDP0RlWTnbZgefHRD4JvPRUHtgFde0N86ou4FrfUY5l79mBRR4CV1WtreKoHH13PDq3uSRZaFR
M2H6zOZUQSnyOr9gnY3ByLfFdfcOGw0uM911zBNjuyBP3i1SmIs1mcdBwrREj0Z0Xiw+hyNeTeNO
aH4S95yqtWQ/OxQxPJemKlJ88X+Ia0gbZ1YNM3o51yghEKCid64c5kDFAgA5pMXJNGDXnY+P7+oa
hnHRVYa6xpH2Bsi63BG6HC/OA390ZcV+/d0OYsumjFFDGyJ3TOa92j2nOfjINb0Ap/jaecQS3VnV
GLGlTE9QcWKEM1DyzNXPK+mVWZS0XPxZkp4pQy45re+damEEkfR9G2D2C2vb8Y3rObiEHeIe1dLK
uLbq4ER424hy6aht/AwRacw0deZlajdv7CnxJHRLrHdYj3oyhamnM4mSZi9/ToLcdih6yMfbzv17
L5DwItUnQojAMBqhiFkBhyzhltYqxC+k7tCuiMNGK/FnD07iDhINBGXVdAL5Kq233Y7P3MND2Kbo
RkYf1MgQKx0soNoQA2F+8g89tika2pMHQkH4de1A1AfhkaBKfvHx0G4fLMKwmZJOm4WfpZU9BZq4
+0ZpKmILSxeUMrwUfmlD/nnjw+uPLWPQB/mDY5oBc7gQlZqCTcERFrLcOFgQx6FFsrrTuXelsV58
KWnbe7gyktuvC41rCwrX/qXp/BdoT/piMMhXLVNoiAhr5C9T43L8EutURhTQ1brWEjSrOWkTDiAU
5nOonKf9jGVC+IznHbTtc1ctH9hplvTVnpfM8yog8X8skXZ0VjKfCvH/Cd0Dn8RrBxjsc9gAaoY8
shWE+iaSf089g0QwX1WZ4yK0IVBU6uKD6J3mIdUPpAou+rc6mWTTKH2BbtxWYk2kEKD4Y9Mqc77s
2b40nm9UFyGlO+ltvlQ8IavKoIdos2QUHRs+5rpaUvOOsE8CqXh+Fo9YsnYahLaq6nQOn77cm93Q
lCKLVg7Uxaf+RCS1w3K2ZxP+LhOSWjVqU31QvJV28m6h8wcgotVTQBznv4jnWciBfbRoB+YXeK9G
8zHP7JoYHZuqwRWS2Pg/dWCc3KiEe7KqI/Y4uhqS2Qo4yXScsec1toVzto418tPh/9b4O/cuU2gB
t5VJrosTeoVLZWfxivfgYGFqMYT5HzSjOpGe05+EkOSQi5OVcvcWq3+3S1uc7md++gh3IfB03pFT
OBiJYO8Ra8NnSP2/i5z7+drqQDDkiacBhkca4kLTnZ0F8VaqTz+5fpFpKkCYc9t9zAnsWmHew9fL
1EpFTUgugJ9QcoplMBFQ9fLEFa3BOXwE+4huaNE+AKLqWBdvxKuBCyLvVx9GLnRhCgVFQSPWkeGq
EyDQFKPQlIYxztkIZI0sQYSfK9B5XnTjb6KoVM6Ub2gGHCLa+7XPt0urpLIhGGSP/jFVfPLQsV6E
k5jUfxSQi4KPpEp/Mx/znkU4xEZZWSwNKnPcasz8DEGQWdZS5HBsXPDovyYunDsaO2QccU0/oxNO
Yzsn7RAjeZ0XQ3LSsk5LpWJfPGt46tkMmonAn8M/t175qOARx85zbT/KO5pks3hOyCHkxlIv6rz7
Xvr3+90Ma+dInWth6uJGX0dfJBg+HeER0Eu0x0YrY8SV0YDll3xNQqvK+lZpzD7n5AkRH99X5gd4
AxOpVietjgsVuqyMjg+bLWz0ODY4nhXF7TPo+2GNf5StHAj5dH66piLSZ+AckeyYKoiE2pCmRnlR
njlsoKIabp5P+cx91gG3+S5o6xrtb/Zt5xiFPnhx4iRG+ZQmWKy/yyULQ/di+fOuLRUPyvM8QjKH
/rntdfN4nLXWYJxk2zRk9zBLSwfvcY8I8oTIxXNLoUDq+u7ZZXgyoXoRF45Xvvpr3y3XvNyRSDBU
pT6XXI3KYvJzCW0w151fsPkGtoa7KAMaAIqGRgfjYpWRT73/Tp31IA33m6cQQx2H6lIQlOp76f6p
qwme/YeFdEXiwDO4fsMfVkycS/Dfl1nKhI1lZeUL5irENu6Qu77aezEPbysFaV7kOeqZcyrmq/Gr
mG/PJY7x87XSwU6PFOEMXVotJ/NswARmsa857b/fHnKqKgISrrBQBczfg8WVJ7wWXeF/dimhIAqs
oj8xpvqdZnHfOBE+ErTCOWWbNHG8stDav45eooyxxwF5U6aftTmJ6yZU+9nyochbWzS8D+BWScFq
io/J33pYIMhdVRA1fpeRzRxg/RczqJO1EamnrlPc9DbJeYMH7WVb8SYm9/9nA6a4d+6IBBbrPgQC
UAd5WiRv/+6yG+c9EstfQfOtJQ8GmCCD6mS6LaOG+mWv/bk957wXGJC8nTqYPNaUHvxo4PSqK+Z0
PsBzyUdMwhWo0xe82BfbVxC7GkCCWTL/7Wo4g/JPmQ2LTjgqAmLeHG+NiQHw5XkT0pfMhWkqDFWT
RIR0pAxMIY716Ejks9Kec1lX395p/75T9HkoFGMOQCQOV3Bk0HW2DjAvLtSULI/OmyguOhFxN6GH
IF20b9saRJGNVsjSJJJ7HNZ5Wkn3XEheyX4rrvHoqLqf6Rd8mGw04p3pcIEfx/13Qj6NrbR8RPcr
8O37Jl6/O90v8KbjrsCn6MVyMrzqZ/vylwh0erF66gIM2GoKFgFxC/sFpopZqmQPbatOJvE4rl8h
fRxMp9yVhVztwd+Gwy3UE6Jv2taB2orBxY9tlQz7fqlXYq1+9/xEul7g4UYB+bIzZbt46rH1JJ/a
OrxkgjBNR87Yt4PZmaLprPJEZ+MRaAGCE9eSTtpItNgyuI2mWJUwk0atWwvpAZCqhdBQLtYP0qfs
j1r5J+n1nv9hxd9ZulgykV/tJU5xBDphY5xnsdeSmvdkkZoirFn7ekY6Qfn24iT/fS7uG/wrVufm
YvPqSPaap3fFWU6X2/l8bj9K068Cmnova0L22E4Q0wHDAu1gvqbNBT8g3prTxEINA0Zh/W5Yfp7D
cUDwXzJelnx0cmR3Oo4sWM2nnnZCs57MR1Ci/V51CMkALJHiIAkkXUYkAsWJ8NtBrDZh355ZpwYd
HYupNsjYm5lUT23XXPLzEdFkKLDydD8eCiGEp8yD64hbxsPhTN27Dn98LwGChftb3ugVtW5UHlLd
Hwt+WcgCJqSNvhHPXbPZuaFRvQgqlALV91s4gZBiWgmhmAKCKiMr0f33k1J4GxRIrxm5B3ENFjhs
KpHGUhWQWNsh7npmUyQwGvOqu58wcpdbUXybmLIcMnSDsFG8xQVoFlrPPaB5NO7thMcKq59scZwq
4wazMfdcCf9ZMfASnnhRU7PWqBZky52ZTBG4pTiQqc/saKE2gV1wKAmg2XzlFFModJkbof+iYyL2
7yORghS9sWS4yt/QEZ0EmIfJ1qlBkIz2GxnX4EL2gAlmKjs1OPDJkLTvywNy3yy4o9ttPExwYg7V
RHQl8bgvEb0AlDp3JEyFfgPnTEH8v1A/b9Y+me4gJbmjs1+tp+qdn1vx1P9HllIH5huiPP3env9H
CLSNJ+OTv5/0nAPxTAHE5EvwhdX5gwmu7Dm+cElDEFJp2/qVRB8FCAaCWxK+4dJFJH1NumigLr+g
z3Z8fpO2hfDC962WhjMtEvU8SmMypFlyHj2FAJxML42nSpPNtv8JLq3XiuR53woO3mWC0RxtILDL
hmcs19+S1XHB5bPpxh1TOl7rN7zaqDNIUVYSr3gUMIDzmcbOjyi0YpTkrA1ziVR/USqW1Ke8xBPa
ANYk4LTK2JVkBw9qpJsx8HPiOWgXq8zX9eNRff9UHWyEXMglO9yEQAQOfhCiRl94o+JZ/K4bYuRs
s1kqLpWkIfCIFxLP2wEjTrByBoCpR/BAQZyXRuhuJ1E2q9yainLi0wJsC+BhBz3UIOAtu7Z50HJN
rwaymtfPCbS7j0tD4zApRsyJHFV/+fwI/TaG04vKAhNEjbCuxafRpkFfR95OGgk4HvVeGN0kQbow
pjqEl6mAWohiQqlJNPs5lgMcILeZT53nIoCe7AQHc2SdjY4wFbKZFf81eCeVjf9K07J78BcTY+im
JiL5MAv8MJJJZf75wqoyQv4xorPSEwe6+vFZav5WeXvTxD2JAF1uKoPSBNDad2x6JrNZMX+RzTXV
p7sGzwaiyRR3c/OJT55vz6yFYLsAuwpg13o5WeOHTySlxDc/FNZ+XE3t31pUkFW7Q0Op+EaQXh1S
eLUEdNrtQdhSfpuAJ6j6cPb+1H5oWgaiDmnl8Dh4Jvtoz+E2IwY8WnXP9hrEfqlBukG+jUy2GXMl
zVeOIWXm4T4UNbu5XyjH1Bv8CQBK7FxnfNhEir8lQ0sAOI1h3TOQakwpaXnOQHgDgIgHRNz2nVnM
Rqa6/J4Vm3eG1vIo8jq/+mIp2678NrqP1Axe7De312rZj33oMobF1QqqOf1GJualfVVZHUoOA9Xk
tR1rHx0fjmGfROR8zPz81RGLvLNgZBA7dz8dIqK2RLTRBS2dADmj5Yzhh4ctI/STXy1dH2iscqhJ
QobXzZDY5ISWaSPZcDUz6VD1/mv9MX5JU3k/qDOplGW08yfBwV2ITODiBAcuwnWF4JMW261rguzH
aWLakjjQdZAVpC+wt6D0gTvMGgGCIlmswwAssErc6j2C2SSrUDRNiZHcs8T1jqoRkfZD/H/UB+rR
6fZMGwx4Xjzqm0ZXVMnXbmQ10H8wQhOhoRTHeMaieLhXrIM2nbPlrkDgnHmymUYUABJUfoaIsKhi
59mDcTRSlcmz32gf21rgjPSHF/l8U8e3T0yVf5o04tuAX9TXA6Bc+tgaWYGzByKvvuj9tqlAlkZc
EVydIv1PbNuz0CqDQV3qeS2eVVdOu2+9klEXkn9GJ2FiR5gXVdqtsQIrxlZ/7+T4QNLuvJd23bDX
J2CKEZmuj3fILDGN+rDGFUEiuOFc9ls1ZrqziK+NNGHaSxOtSomslvylrR3M7qG2oJtkk9OXLuJv
7040aeVWJAb6vENHjOp/8XecdULok+ta/f46YWMDDSyYd0/IhCO/aYwQl023IBhRjp3lMhkIfiSN
+DTXQQJqfILFJa652gWaqpYgLE+gsT5ZIrDgnR/E0s/PXhavo5cotug+IUpWHng6DFSqgpoyDA3e
mcl/l6+y/Nvkcaic2CO+Pl2g5C9f9MiIdbN6aivKKMd0qSBnosD3+t6dY2WjRDN/Ya2EKMBVGFjO
xi/2ft8OwIpQ2CUv44aPZj7PZMTkZqTVoEU1CpclJLUdPu2RFrGjTQM2Hdq3x+zkSqfjF+O4cOxS
Sx/jyLs8qmFOkxTNTigCBjL4VdmG+gfap/5aAqUNnRpQeAJ+xkjIwPY6sfiJvY9hhgBTm27/VEbK
mH6zoejsI1VFmbMOQM2F/cwIXVWN8p1LU39Wg5eHfvKmbXk7K/2u9qaupeot6khNBbzcr1rwhPRI
6t2bIZct3T0TFnKK+3jdCmb/G5nX2OWTNHdrhmt4xHJ+NUsifyICxs+IUhcsZd9JvksQec0ZYBtW
M1U4JpQoLCpjlwAH/g0wmErlv6WOsLvNDRG0idt5bahd8rM6+BV1H6mL1z2eFGzWCv9wcpxW0zzM
koS05FG+Rxk+4TkZkCpTQXKr0Iy4p0EUjwFrWdbfaQoU85u/MB7gftGtmoCCczklmJWGk/06JScy
FEix1s5RsA5E3vDrtYXqA9vvV57h03Aihd0k+nslTYaL3aA0Y6+CnXoIl0KbhLmhIL12zVz3Zc8x
S90G7yOXM5HHuOe+HVvB4rLhX1EBVULnDN9nX7eCKA7d329KhWztfRwCt50vddCcw+pCz9ctcs0m
2ZBwTVSCu1CeobcR+WpD4TvPeCr+A9O4ZVyRTAohGqiGnuKOj4O1vPLSFmVQaoGZDPDQ1HYjgYYJ
8xZ0qQ4hlIdkD+4Ij0leNwCMF53TKLbJeN+E3PJoC3vpjsfe01sdeLHosCzTViYM419HTbrL+lO/
cZI2OXyG5SYgbyX2awOlpO2yvqgxRO5yYwcCM9PjxS0X/vT92ogUMOhEzVIuG6U9vKORSCxT8khn
AqEoW/HgUFWDP865sVMdYxkN6xcOi10Ut8Q1gGhWoVz4DHBv0ybwU7zOwXuxLmcssmNN1HwlZ0Lk
pHXedmJ5FiCmyYOILKNyxcdtnReod8HFZtHTzrxrsztDULw3OvbebETQuAVGc5J+UdT46cw6t5gZ
D4htRcUuL7d3fexpUg0dw2yr4OhZLoI9BdGuGpHqDaQbUuFE21vBQgGqC0of6rzSAxsec4d2k5CO
/vXQ5Xyumd7uSls0om/vHHnCgjw3JzP4J2nj2FeH1LZiUsWoJgvKSpC5tjqgfwwJs3/mQv25uHYm
ZLQSHOnFGcH72b3d/txBf8o6YqFL/Odhr9EwFKQzF88RYqf1H0kWH9uQPCFrpZr689N0sgnUwKE0
nNmAmKIc+17PUKzSgf8e5zq72Is4/64pcxWmrFkh6i95Ou/S5moUG/w/Q3tRrCZx1ZQdTR1k2ars
8wwBh9p6/6t6pknClXWefai4zbHaFCtbPVdhCWkmWF3xKQ3YfP6J9ZXWyjuXzuPfQ5TLxaTG9g2X
373WOm5mX2DU+4ddNeP9rNOLgaVNERJnCJ/CzwtHA3YoM0E1nbtHGZGrZOiRALE0fNygQZk56Njy
ejqlmrxaUc8jqKhDGXHEVWqSVvXPeJlym6awZIQfT255f1n2fwDu35+weNUoueoporayMLl3u2RC
34Cjw/vjBAhJcN0Kz0Y1KCLKpZL4G0C4IOwcF97sgIhxWzrZN3lBzFlmSnOK1CBwhkozVfGe916i
HWUFE+X8l2N+Gdshg8+YG/aKK/pSGCAvyP9X7HLKKGNwDbvYR/csXS3zdncwIDLUrfvDJfrDU1Qa
n7SJ3zk3QvZFZb3Bpv/o3cd+OMcvQVMtNj3+UEBJiSaRr05gEe7kFIB9ZtD2DjKjPqax/Vme+rCC
4l0v50TF7Ww+b35XTMTpxtDIx5FzRX4TGg4Q37i5xtJbjq1iLC9UVokyXDyD4yauNEEnyUbPxxj+
vUQpoX+31dCsK66Z6d5L9MgazdJi09VylWzDTC8xcVj8rhy+cAsAuoZNYmmxDJgXe+niKndYnS0y
lYCXVera41ujs5gFes2+PXlD6+U9orESUWQp6HTUXfkHRyME7+fKs+fRd8jvLOQZ15kVwIf34Zsa
w26ybxdct67pn/vD0H81WNBKU68DJmO4Q0SvuMIu3HXl27Lsz4i2HlSap7z65lrXs47nM0tZvW2k
IuXy3CYzjbPQQq9HeheuXfbWXc12gBIDPJNB1O1HBZJBFnE3AKI3k6pAZSDJVGJscsPuWUqKfQWW
VbrXYfo9qMEGBv/OAl0g0KUzRWLHewnZAIJ79Ql+CfsrkIiOYEQimpHTlJpxviW312b3V4vTz4E9
nh3Ek8dvWR4gTiUVR7OBULbdj55NmTrAq4LUFVnbCPNgNlBv2apJrwEBzMXM2VHF8/OqhS7M8dO9
G7JTrNLJ5vLb2c0nym8T/LftorVvQOahUUY/jRg8LyUOqOAThLvGvQWehIMH6ahrhlzqDQ4W+NUF
S46MGUIQEx6wS3oV2J3to2SCt/lYdSW3hQREFlRqid5DGSgPmkcOrkufB9o6kY/Qvxs18gP02ech
i5duvNL0Rkm3Q+80/ZwirZsOMoRrLjqCHU93iWqz1Rbfk1wZUo8EH2CxWMm2s77LooysKFjsxvqn
KP4jbWvsN4mt3ON33PtXHSBEUbf2sbU2RarpDbnNrDUN85qx2IPrvwctdIRK2OxRE5jZ4dkGlCT3
7wAYRpwqYcPCCKzYMRVLnQBGkm32MKwfdWzhSnwF0gQGmhThhbPYsPowEGp2wx2AaFP86rdqwndr
zuhYweFn9hUUAyPbtbcaw0qVjjnBBELgwRaJFpIkZG1qVpSIvzaxMB43VKtyf8xgyLlvtwdqw9/0
sMx0oO5bBMDDYcNHUHKf9a3YGOScmExtfXRokkO9wJrk5N102JhHJ8Fce0y/XaPvzlQEsJezy1A6
0tdrayDPxGI+kR6FAOS0nGbvxIQadgRaaZSeFKxlNFJvfYLpgRjgIpg3aRZJhdZ8W9+Bbuj/Ujrf
wxWJOoWMTqlb0lncaUW4GGjep8RWaDBplt9SwcBW2lksMQ+ctklPjyH/HH4LDVxNxAy2eUAPd/tA
B2vMuv5yuuYIKkgiP73oG7yD90G5PubxSZSfmDbO3vXPtjzWldv+scs8GXqstnpZ625J9JDwSwp8
8E+VZX0eBXFPOEMrRqcteV4/s5IlZr21SLFrIS9WijPl/ikGLOHaW8TVXhJcmmiOaJmPrla94DKy
zO0swDP7Nn8RuGM+7wSD+AKpyWW7ZlbDnVNigBmsiu8qVa8mZHPjEpiQzihgjHnb0BnF1Om8OGCi
cGwQqYD85lyICvIsCQLfKa4tW1CZk5ldJ83UBvt4IPZYQDQJiLzzArpuIBMl2YSnbzHXe0NMA+V7
AMOP+1b3rBLRsTMDoEzZ7K2AZk2w+DvnCpfg3EE+fal1p8VIngCOzWOFqFOvZrf5J6DH79OsU4pu
6BY4naJDYwRdq2RO+8S0jvqxPaI2E+1JAsMZJHaFqVz29rJfllkfSjdPfOgRo8DjG5J/4/FvFg7x
s0eTDfRJYK4HLQup9ytQPzX6lz45+BaIr/LgYxYux5ixJenv6WHRB+89BEPtpxnJtIlXglSCLO0z
luXBjNlClz0oIb6H0SAoGuddQchxeK9SAJCVTqW0A3/G6Fe2YvXKWzn8ixu+JFDA3j18wILruMFj
M9yMEuKWX0wVT25OwFZPyYV2JL/ongbxgENO4zl5bxUri6UylmbT8DSIr8XfUmIi0kbZeJEyVBjf
4Gmy3kVIk4bdqpXr7QTzeyvG7rVSzrCyRyD9bkvtJ/hQlCtp90AkMcyJxeaBRh7cStskPU6YhBec
jpTZg+l5pqtfmAZJxrXx+34Q2mmLJpjNveRtCIHcS3/W1Etp66hagJXAeSOwaYd2xSRQhqlYqamS
TLjIQyn4/zXf3nCh0AnPQI4g8SPh05GgjF2GrfqcShmjRrvFZFcLo1I1vN3WEOOhsUgy1Qr9BoGH
yPj4zUzlz+PqS6r2LCs+UICBVyyB/Z7W4OB46gQFYUJTK2Ex8Evi1byo288/YY5vPUpi1w9Htaf+
9O3NYjR00tIf1SgidZQ4Bbyh/7otp0hFb/YMPpciqhpZWC0vL5QGL2u+gzLWtg0XAPnQMlrDHr01
PuO+3MFXu6amZmWYhwgqn5i1e6ZMyfBXQI7Ualfe5PdyJ/E+h8MHoKDmNq3JWAsU0tf+TgzNX4o2
YzfamXmm920adJIroiSA+4R6On2nw1SD763R/U5WjEtr1Y1e8TEUDrFsEX/v7NmkFTBtmwyAFXBd
1z5yKobZ3WKWBJ99XJ7JDStjuvkvbfOp4zjSpZoP/fgaD+TvvlaAYDrdt9n50Hpkz82drbKTCZGh
ZJjg/uDW7NI5ccm/0TIQedVukBXU6Av9Nh61/WpcwJ2s+tBTsWycadXw3f66ByO8J4HeNJIREk3f
TeoN+C9p/7q501j2NGT2Hs04HHkYbiqtRaCrSd6bIMd+qyeoGYKeGgswPtSCa87Ry7dyA3B6kKu+
FwZriyW0XKdzVfpkAUvhcM5B0CqIYL/2h32WBtoaP7v4O9wTWHJBNeL+FuPt5G3oPbjLUbT7AveT
1y7fJYg9H/XKAcIYUADRXFjpT1Ce4Kj+iCLPiQi4kZbAuTDbIDPPVUx1jrVZ+Uun996oNdBF3fwE
fmcypLCXsoV12CbEjM/Phbxunfoo79nkKB6mBT0kHeISZQCpW0mh8CnhVHJFGpwe3OLO1Bn4VvXf
IcIafIrRj9pkv2kqOAOD+jJxrcW9uYQZdxiU19s24oYbv2mTn1tLm0bOz/k6pZ1WrsahUur5sulQ
TqjpLYeMZSi+P2yxXlZbD/38dYbUUUla0luB2ix16Bs0WEbXMcFchewH1AG+MzZsm8c52TLjEVNe
XPYO8xUZ6P/OVUMcEZIKl8nYNT7vyVvHPTqN1RVW5Z7z4z7W6fWxblmNOxYeIygxsnvvvITztaay
nBtGejHQtU44vgVm0Y3swl7kF4ar9ox2u9X/d8MkwI5vhljg5cxfZ7QChyqSguCM7Q58llVjM3FO
4pcdua2dmB35hHmAEYmGRn1vmp86Io2+V2a3q/rMB5/0QbbvcEDdonsY3huYUNI6T1dM0oPB0Mbr
poBACNu8XdkkUi59RgmGMvfkhiLKJDFyxBHwyCA9w9LxBoEkCK6jg5X6MZ1Jh77+lSS9HeGOtjq3
mduIPSTmcp8fsouHyjWGgLZ4fQnaiV7o8s/l7L+nNtPlU6rU6P5vkUmO+Si2Ao73au2eS9x9h1rE
Lr2te4tZo3FfJhcgpJwLunDBpMk4jmFzHeKd7oF9Ln1X0naSv+Ak5CpPAc9+decSQ2h/BEdYqqfy
OCXGiS8+261WodPy9NmAcRuMq1U5Kwx8sfkF7HAwV15c15WzUskV6a6lnLXNa5aiUXhH5WmXczEo
rsll/rLClWsOAAPf7t5f87xfjV67apstWCQF8vrTOjI7G82HxU2H1eiyEodFg1O8Y2Ju6asTx5p4
5HCWPWGAQMQRVX1781vRPfJrg+TMHqSNqoMQPaSoaYM3Q1YTzgtjGGV6+pKYwTEzoVnp3MOcmZmi
YgebU7KRdH+1Kri1gqqWqgijFazt4hpJuUCWZeB4RqZW4zKn0/MFDIhUTTF1LD/aZvV+YRIdg5iU
3XfFVkGZdpoMR8WWZ8DIX3WAVpt/xuoY9JSdsjO8V4cmllJMf4xgWnKSkk2zpZKCxIhhYp4HAlUR
Bev3kNXBOt2w790NAVVTRDOdIopXRWOweB1MWUQZq5kLksCnbkECmjVoXjczr9JhzqZrXE/A35b9
+jUkk4ani1PTIRgXsJdMlLWSX4xXo2EkefFqJsqveWLB9Y+a5qL2NUwQwCqGW2ixvRZcwxNxVYpt
gJfmV8rLPMhQvXbqqCdptfsoabkNagLnSQKw3VmUouFNK5KLaapHR3u9mfPBYyCHpxp1liiepgBR
jpBXQrf+TudyjQfxQZZAEqxoPjCgzjTGumBhmXYgtcyqKizkh/RFDUyI/rhxxWVVWiFBomPwtNvN
9kPsOFf0snsLc1IdMVAqfuth4t4h15Bpr/dAPdDx08oJejb60dHZPeKUyQ81RENhkMRphZhZmcbq
it6Ax7TjuRJkg/lwhFEF80x3p8xk6ZmA1fvrt89NWqxAxbMFZ0Zo+XYRYEEwsTy9BoGDVftHF1Yh
sMQOl1sG7uEjFKaUZuNAu9A9hH+/NU87ft0oROQvPpEdjijDMOXy187I/q7P2EtE+77XmokKPg+1
3MJvKect3BTmG9/3pSzYBrDmJc6Y092mm4uWGsoFOWqMXwqNJZOytKkTTASMv1ilG7tGmWS9EMcO
Q2Rw8eOo+nrk4/PKLI70WW2nvOsWWxf8fx+AYQV/pDHNgEc9tmxUXoKJN9ylqE9a/osbZhbduBz+
Zms6Sf4F9hQIT+raQVzcHzsl0KZC6IdJ923UQTT0hnf4q3oRpWuxVSPHK+hpRLlVEN3P46e9tNNy
lE7THUWVwuykVtFiY9X3ZmoRsQUCGkCyGe65kcPYRONO1yhJ9ud+loaUDOP1KrVCFIFqptLiAsT3
pmIEz/mV1fbu1b7IvfQRdSD1Wzg/kKrgh7zB9VeveNBmr1vXJpVpC4oVLHV9vwhLebC3FMlQMT+o
7NGS5NOtxSSxAjvw9OvfK+zi7g5VXSKrs4e+RLV4CZVMdSkE4uzGqEUlrxsdsHYkVoIhbOj+EEAe
bu2vOByGa/Tz8ZccCwY1mtlewLbEtPRH91sd35u/LU5SeCIE1s+Y/CXtM4/u2YdPwhmxokuVurcO
LNjbJg47iAj5qKrt1qAXQbDAvf3g0FPNpKKTuheamJCmk8la1c0SMQfkuiEdpphzeICkNnIFIP3o
HcGT0EaOscVLJQyfL1YDogr39ZPjtn5ZeMZ7D1HcY+3UUY1u5paUV2aK/CsGl5+0Iya/Lqbnskeb
dr2ln0UDMbBfpP+7Q4Tgvtq97lrr2ZH8Z28JjXU++g8TOyIG5tYa1yO8FYNRhBkkdGlUUV8vX08w
aw4gxqA+DxkZozKVTWOEfBPrHQY6SlkhG3geKhkiIs5jv813mEQmgnd+2aXs3fwtT1D3trIbGdPp
xZ0b0l9DKdtzq9Tr2xA+dhZ8p1YogmBoaFCzpH1HcxxJJst8jgxm3p6QbNi8iuSE+5H3sYmZ7DdW
mi8wBHS+WnwudpvT1RVWleGjVpAvZrBRtG8bcmyJ+KQ60ngbtS/q4RsLwW0Cr1YZh7aab6MZ9Ckn
ykjCFEcyhoP6xWWubBUBXTqt0zQ/LQojRknS1lSTXB9nPWxAHGIeL2SsbR5SC8P9aOX1LLrr5i6f
LvLU3QZEOR7hu0MSuFgy8smo+DCTxIylTMmpu8YWUt/gKTlkOsV5l6b0+R69lALm68cqmYDPIxcA
RgMd1P19W4iT9PHWocIGrajoS1X6c7h+Qnj+1SBWz0Q1TUNOuB8i0lV6vc2PXA4lpLtbsKIjnJIi
Og0ADO970/o+ldk22WUiJnRxv00VXzltBVJhnQzpCG7KkGK970L8W5y8HPSPOCIwjqxDwKyeQzXx
OIYrTt6jWGQkHNRvCsCvkQlbKGSc+oSK+P5h0oT6NPOCqR3u3WGOYArJHi3LZphok7Yb4QK0dS35
5XMXJnoenJM/00huLM264khv3GUrKsOhydFv/fWIEJS6g/DgwggzA/5x0WEaERcwfVFIWP/NAn1U
xpYEcxMz/uSQA17+7ik2xWBTj4Ibhd6kRuI3xgAA8bBL+P2snhv3bl91EqqfuRWPbV64M/nh/xNa
oVeRU5lghFJRTGIS0hk69hTrwRd/6q3hexqeUS5V0dhPkruIFH+6cLj3IpX/nfz5zSzC7oVdJnsN
I8YseSfT0H1GwcbcaAbycfSx7xRZ/sVQQTtOypHOy9NV4M9ad7wC4RM0ywVjnbW8XQEJyJfzbNTG
BKiXb0PeRDOLVIFC/9qQcALvFsO6V28n5kCy8PLs86utkXjfN+vorOr6tctqnNt4is68QbgFgjos
uXW+6hnTGHdRYK6bXMzaKWABn2Kc5hCcQxrqwfBcE3KuVsCrqSTFUPq4Vk4q0fEEj5Lf5qhCC1yx
OjBMF/lEYr1X7SCqRtIoi3aDVU30P9v9nBtbvyxxNQun5jZZnOYme9TpvSWJiDetJ2hLO0zZ3rkW
s1yMdNmYhi3Pr37X3kNb0TQ/89KLqZ3AQg31dbPW6/6aBgLCsfCkZ9BVyVgCmxcWoj2w3lgV3BtV
KtGH3uQ7aD24S9ZexRNV0WfevpWW9uifem/oJp+OxqwrLc+nDDHO+xBap8B9Gr/hUjWJDaBZ8Bnp
pmOfbAwila6WeGcwZg517+K4tvRkWyMbm6yteC/eh/w1nM5k90Mp8qat8H9zAVNelOfdNyv+bmuQ
NpK0VvNk91sNTPnQOVWeD57parwmyS6IdSIWswYPvebQZAhA79AJgUCcDcMfKtIRXuQSPJhEMRIz
FZWWQxTRzFC1TYn8qzfwCmL/JTC/GUWjoQqjU5tzOczGVWcnTV0Y6HMnO5MbbTJeGe9M2OtG+fGf
aIbfJ3foOZIM4c1+9Solbm48tl2lzXjIMSd9Andnh5/gUk/E2UrHfKwBB7AuSeX6oUHEr33PiVGf
hOSgnjrDkRld6yIf1koJkNSCQHDTgNrCv8Tq3bed9pwvyz3qlF3GaOhJpKJfAmzbTb2VpElaCUeO
PgNo0AVLsvy8Ifn2gDbAd58BH8MqyUoc+FwbJHdo+b6L2wvNK3/SX4pHe0LixRwIEHqxNQBjRtuI
6EhePCE5ocvHs1sFL7w5XuoZnMOLhJdu+3KR6kdAGuUx6Edd1yDUdpmGcyhYv4/s3b4eXkIB1Sq2
XUQAp+q0HIVisVeNnBSNs4zysqVXYkbDdLV3iRZEIqSpy93nZkjjxNzWCe61i2Sf5ZRTzNlDFbJI
RBsVb0eb3q7j0JGNree3jMGPZx+JfXuOuU8gsVyiglBfOnPXEdCtTHpO8SzmfkdVs3hqluRipfzw
MK0KguIjlTtAJI25YnswOspx2Rr4FIXmeutt12cj+VN8dmseepPVIV/VcrriLyYVj7sBDnKbyjLs
M6WUu0wf3AxpAwlDMx/dlhKH+pdrEz8w2AIvROUp6g3sxVWAPoB4kUztxN0MVos4CX5dckq5dGBc
w+PY8Z4fN1u3irtx+gwP0rRv7nmYJi5Xe3SekHoEJsUJxhmXhb44zieCTI4hSILyCCXh+UIL6PeI
5MJ7myY7jTqwgVBfXpm6jRCE4fxomSw1Df5K5aAUroO9cnvMwGTtBCjcGIfqV3eoMe8UFsZnNqsn
1LjcW0ujVwb/USVu6+aIIHz8WMY1tHtCqb4KN3cnrEX+xguIJ4MnFDOQvzIvbOWoUD57PiUtl498
2p0BGwX9DSx+wf4i50XpMCEhND5pNJkx2cKjdo1jfNmGGDx/axnhD2Pcb5hO7LPmMhtPAmIw2/8c
1sbcTFbzvzw4As5wR5OZZ/bKwf0kwYlPkLvu6GfFTrJxpbfq8eNCJn5FStvfHrvI0nyxuBO7D8nG
asJ6C/ZGAmSs6YV01UmiayTXymiJSupf3ZcTSr2J9K0mrAyW90zXlxKbwgqkGpdTQlxxMYb2xMuS
qPmMkdLeftXMxwbYIjtcKK/5AKbM8ZTjYLQrk3QKMZG8j+1JJgCr52a3m8mdwgBqw9BrKeiugYqv
0x6hBh/JlDMTERGuzKj2vGmHfFu2BXPOmp037jgz7HqUC/7JUPAim4LtpCQKK9EaU+kuluREI91G
aoIcVEtgpz19Nzn2HtxqbpKcsEI1MwKyXAh9xvU5tWyROoeKbXZMStIa54c0o5PWWqIkdFBKy5RX
59LU9hqt82CodbERSJvj5TbaDF7U9EhYCiCWvlzQj/psRv5ty+r9SyMOISpGpXbCe5/VA6/LN34t
TtpL5R92i63HV5axjJNK7pRN1d5K6oescJbPkF9y+4t+lM/UCmX/WXV/XXcGIx8MIzYRLFCS9DdJ
alOfyN+V18LZl7vHNCsGsRO7acbmP4/7zv6NbcqW+7yWrhZi2jzH9h4tOXFZxRl1E+fgbgir7OdS
fUg9oHoisoSU8SgH0MzAd6e053jsJKYhXdUfvk9/3w8uBNPjjhB4NK3evsoQW3XlBuDSpp2bA9zA
7dRjD3srZeVwGInbCYDXQZ//llPxGMcqueGrH91XC3XATx1lqjd2CvIDmOsfqhzGiFQKpQg80dCQ
tle/Oa27lNYxOd/7NZxaQ7EuJU1fpR9eD+PiNg1dc6nkp4BFM79rYuWINL+IAbhkFTL3of0ghCPS
JE9qd6joiNcInAA6/hKqMUFbvhveJN8TA3yRIvnj5HWWSf4m1hx187sgAqXWFY+kJWhgt+LTH7gP
+rgYBr042WhAduq+6X37nfsWrbo+GNM8EiGzKtq1gJORywbFs4BqjNjH31IQpTsOuoqO8UdP2eri
jCvabwPEskxmu6y4cDjB8xi9IRZ01xykS+5rE3MvBNNvdBb3nnXva4ASBTft1bgy8EMPlwNMy8Cj
bf8jWWZONIp6kANu7p2hfM+JQbXBO7YQEf/3s+rqlF6BBFL+Mn9d4xiGgToBf7P811/NC9G+RZsM
3JsMztC4BTFwy3RrW1qPw3ft+OsFGIci6zxYTsqKIXGLljH9l69vU0q8nhcc8P0Nsf/plQvGsRG1
/gXEO/gNja8AP5ckuJoOKmyUjsKlrxAT7I9VlAmJdfazf0jgnLvZYXt8k41WH+l1Z9P8MiKQsudp
5QuI8iKKwAkexU6ru9FUJaZO4kDG7ms3TEPcuNhFvibfhq73TAiTLW8P3OE7pUrTLXzsWNcpoTUV
QD67LuVNR4bqwv9p1QEI5Wy+NS37XhTPCDDV6GLAIas4OuSZtM1k/MO53ZIgVhCJewvnU8aCEDo4
Gx/ms0JhjsiuruvrhVzSbrfuqtiG/IdI5acsfnwZ9VfAMZ+30ngUl42nT9AqzYi1EUJ5AKUWlZWk
OvFLb+M+JY2eoE3eZz5jloahXZPy6qW97IiH5LvzDfGhIJzzg8t2qdPNYxSc+vT58KJZkZ67Z8VJ
j8omaWkDc5/9kNfdQeQM5pq6Zn/X4wfKWjiwyOrwwHB/vr4GJyOZTKC03mGWjgQ8ravYk2xNr4V4
u7iDUXFdEGfnSSaB/D31VC4CV86QA5xsaa7ncDm8Kgvlv/mUyNb+ZrBsD147g/nyOLrOkPQ9BiFT
PqJVKBdp02pjg3ZuglG+eir5ITXwxVQg+r6rxp96DsHsYv92LQgSM+wEzktsxY6vUi4L6mwgIEKm
ZaLS+NaXG26Cbb9Uk2Y8oMnI7UhZBUiIMkiSa0k6iQhJRXmCYtONgI146YqgCE4DPS02yVoahNVN
PAOIqRSRuU+tZrR/p8yq7Gk6PwF+J2e+6XKREvawZG6lG9zA2NIubcXwdxyu/65lfTf54TtcdET5
ojVR5UI6RlJBVJXfS5VBAXuixeFfEyVQLOLwHRkTSZ8bST60TzECeWIYTAk1a4nsJUgZnXIOUNGz
UYeYRgn6bSC55qg6ovROLBZ99+pnbVHB8NAilKmfA3khDo5IeU8BIXZpSCiWvLgaB5IIYFqfBl/A
lewJwRZ5H7mFFuuDcqXVU9iMvmZRhWS28hVtVttK7GDJ54yc9mgKL+ZN5K9E7t+6Lz+CvDdTwK8S
Z5bSz//OChsTgig/fs0tkzrp0GnVVHCTlfXiDi4IHD4TSn/yyH2B56uZG6QqMqfKEtNV0Z8GI7My
lvQTHTyYK2ZFSeeEym0oFKSCOFofHlmY2fRYC2nodCH0/IXK2/RAbjncFqAB3dNDu87xbBSiXkD0
4pb2rY89dC2yWBZYt9SL+3vNwX3Sq1yS9N8SYsyo8CJcOQQRpC78x1FMWh6yAJ+Jz7B3GkI5O/vr
5va1fph+V1KMxiJdz9arqwzuftBCU1H+As0n4hWoeM0A9hFC+7fVA/rt+o2JbpNEUF0KOD6Kjitb
r0zMZfAOeiVc4Nl0wp71INEMHSPC/J1tyehD1vEFCtwyrQ3aPw6qyg1t81j3XMIYYDsHbjG7Nrdw
niluiwNfLn9VDzuq3aBqsRf2bX/3sZBuD3HdyQRQbd9a1s3F0MFJpCyyLkdSfMlm/JEeySpsBaku
EUAIeg10DgdD+7k3pFn9b2JHeYpk13elwMN/h1za4GKinhWZbaMxGCO5yUSRyzlvoYcFXWxHM0ob
3Y3XMh0nZLaRJZN8jaF1QqBUjVLohGAa06RbHFUPhNvB8A+IhIQGZO0Y57LiU96zhCWapTMhDJYM
5NVWg5DmlppAZ1MSqBBo6DZQPyKV0hHCYx6r9X+2eJATGacRx45qF6tp/kJnedoILzwX/OF+z8AL
elYAbUIE/G5ibyXZG3sPRRSM/OBd8wELOEN4/jgo8gfQ9CvTntpDZgB5h6uNIFlQabxRaJzN400b
45E8gkT9xUtPCC9bLayB9kbVot19eo3DqaBpIzMsGJLpY0mQCV10hG/Mu+cjQXgIbsjqbMsnHqxc
jQ7gadj/DJ0d3RYBBOxNAiPRjvIpvninL7JJqQwFvUtmlPV0etmKRHG2k7EA0JvKdyWisaJTGkFb
P/8Mf1I5COJuIAk9/i56IlzFYauYJ+yXCgiKxTrtDZYwWJp7X6ym3NN3VkMGy6Jn/tH+L3OZZoMt
DH1A2tLMsNuFZdA7p0YPXkJFPVXoEUuhDxtqYpq0GjMPNAz6sb3Y0oRl8EtoH/nxcl5RS8nrEq5K
Jg1sjE0R7/DAbX7Qu8HBb1oVcnKc8NSCjK+lkr3c2mhOgbC+8Vcb3xuhUMsGpdhAkOR+dVUBGRyS
gAFQLiPcDX0kkJidVfVyP7sKtMCvUNYo51Mk2zImwnXCtuEQ3Jvoh7QtyotHg/k++sBq083qe/sF
B4Ny2rGZ4kJKp5yNcOJN78LPiFP2DAre9zg0yOlSy4+zenEO13abI3hhQfaDQWNJXKp89TtCaAgy
xYPPnkUEXM/SQ7tz81rzgqVmHr0kGHYH1xENqpA28VTmtlDcrhFmGbja/zgaNs8yzEQV9L4IukgW
aEUsKI9HvBxKEznj9ullh0PvqNKSftpLsk3b02D7YJkxEzTic8ICvGaerXVnI327/8SGEutEXDsF
zoCaU7XtA8csq/uQsvctHxxy/d43OWcvFa5I/VK9rZs3Q5F0XSo9gGREZ4pnyA6E0L1796Ah/V/9
5eZ+TYpa+U92uunnudnMHZXMv9s+aenT8lAsyMJG7Jp0rjKkYoZ0NjFuZ7lGrxS9NR1sd5jh8w1r
7EAz7NjTtLoDNZ++H0s9xpi3OcNfRGC2ADiNXuYmPRglre1mVR2p3KzRdxsrnqGrUbCtgBMUVldh
aJkNNybX3WSgRaB+PD84rjesY00tVPuYXLZTXMBf4Wc4ZjV5nYHuNLU2XJsBdY1NWi2IyOQ6Tzlg
W6jUvxJx0r6rdCO/of89he09wwQxT6xgJEKVLLY1EECt96TUm0DJKbHjwZvbHm2pj+gTQkQnxdma
sDQZ3aXjIY5Gmb5xXxDkZhmNQ7niDTaFR5tM4jl7xCbX7Edn4ljVTHCSbDqAbYPo22BO11C9YlBZ
yLwBL3It3/FBkXVpG3Vi1YZAaJylvNw3Hsfb1MksGaTNgDL99YVskDujs0I2fgG8fi1znSfmsSgl
ghZHnH3mdVEaOmVaGEJ+qugpU/nA3TaPERMDuKDbILd89KqtfIP7j8vRn/R6eXRwSDmDIgsyIAq7
j8+Bf3G278viKTXNYylpoFifSeaN1Xv9UKRWEzCmg1rpjdFta0QtJ375ECoqXtjWo0f+QsiAVUPd
UekB2wTM8CMzh/vQhHvTgrFU5pEQ4if967XEQ2r04x+x8t1fmBkNCDBOv5tMpr48IgLz4aLjwqHA
hO7UTu2sMKBawxyn/Iv/MhNJrFIpXDSEAh1mdBZODikXd+0KTdvhKipWN23kXMlqduzGq6sWTAEW
nrzmfAtYyfov5orw7YMq5ENkYtPsEUWC7DL9Zdjdyb5tHMleA4dauR14wgjx3up6VL2W/PEsOzzw
64Lq1Vjn5FbaXSEHSqfa3jJcbPp3oX6tYIXTFGhle6uTVXxQwbScn5hwcOCxQs2E+0wdaX5rDDZc
SFAjPZb476VVHFPSIU7oCVijpugBbxVlWnGcEbSfNf+iJaYPFdKVo1/sQcxkwsauXhoQ9e+W7SFc
vaMBWZJ3LQ2XS3Dnk2ygZMufY89jmM9h6e39+yvqqpg0416s0RZaIiM6ceb7ilwcCjpYEmWYkgJb
avy+tYFmbz04u7WtEWDC9geowo/wxlDOWQdq5hst3OZrhRRnrsubKtIfWNbnfrwpsZlCadIQFoyu
gouRW65rWdCXy8qoDU/j/pxp9zqDxpu24+vt6f7AF/7wQn6yqjmTSVvb/bWz4S6ptIUp0ZqNyvEk
ruhtgJS2e/41yWnxkbnZDhcBNOZOr5g8AauNDwve+ZUXMFuZas3qr+mHI3n01VVCXKNKSoLs55mU
tiDQUQyQ4dm7sHWZlKkgv6wBZltv+wSGU9xFovGrIqxkt2WVLFI24mowu9hJAKCXaZ6iNoMS/+in
uofUCwMQaHJ7ARVZzPODOFlJlGT9UPDK6j8S+rpWr5velTLEvt/jIknbAfDUr67Ny2OULulWX4i0
QCU4m6HDddXQ/fa/LmHRhxiHWoCzCZhhkCuCKW1fy4v5MSNWz8MQbd+dDwHi+EsEXeupHQfnhiar
PQjF1iFKPRz07sHNjkgRpH6fXX0+HnPVIzlUlk/E+bBT3hvTt7ozJdY6AyOz8vhrj5pYm8fcDZ93
UH+idz9tZQLqLEoZR6J6/gBrCN9fazYSIrCw+NE/SnDD6UiM50+ozdd5Ci8h6glShF0Wn9GOo1uP
wIQupTRM/5mmo7H6SE8HVRSe4+bQH5tDBY410yxs4kCnWVii0btjsHMVwR0lOULCoTiuADXlaOdQ
XyMThb62fSsooSoBeYIN7aebK6mKLCs3qyCQUKoJ9OhAFVW9JQvD745dZBtGUYD5lvYkkvYhErcW
tWeoT6vtUFjeYxn1mnf+I2mTdKJRsja9aouj/jcfRSs4kpxJpKrEDnSeGfIQxrDjxPVCqAAKnf2b
YHN4LDMGMwI6ivgOxmihiJEOQSK4LNhgev/RVRWNVfU17o5KuCQZ4JVWtP4Cxw2bcdPIRV+B+dCg
9gzt7JO9HN076L5wUR36mPUquKe901MCbHSwgqrlQ4DhiII/r0sCkVgxO2I9w9vZb6cj80SK2zhJ
SRt8gk0DM9eGWixXerF2PPyDXA2h6vSZy6fnBda5ZMBKPklr5tuaOW8pwXPGtzyuYeeYvJRXDAXw
AfYsqrZyjX9p/E/wX5bG4hPGRGSL0gA09UsEFmUrFPHUpOx+gkRzgeMrIgbAbN65h5vMda45TmDh
oxJtf5UrSyKpzCa4Wi48WcPTZBNvRVulnMWLdwihvnsVBFjcAdEK69+AGSxGAu2mmfZkBGCd9wzb
UCzr3sZlljcCtSJGNwkX03vOmyT+qTDHxL06KpsexsfaJrMLpATaNEe9eZOolvcQ76hnBQ89kPqV
RH+WpCPe2kKhYCANkKdudasQ2VLCqgSWxM57ICAnFVLqSp2zl0O1upBzippRfR2XU619Zd76YeFv
H6fOswetSxTl3XHL3txBodlP4eXPFe7oIl96WxIv7fCZ4BR4b0XvV1gJ0/XkvXuiB89vH1ekCmUK
/ZuQzW/0myvFjdtkbgpyoyXedLkHhb9jMHdVvQBI0p5QiraCnNUiMcf/9xKa0mCi289vwcUJj7pZ
mHnei2XCwFdrbm/48WpiFf7OzhWTmgJLh6YYcBCDPoR7gZgU8xXuR3nnbRk2/dGM5wA0y8kwTTTY
b/F+23TsQrXd5lufcSPr7/w3qx77G9E7vBavmSp8MreRr5uCTbA6i8bQ/Dc+ozGvacorSeEDmXPH
wPpVUhXZSH1TqvzHDo1kmYnURddoi5JjHmJRNlvAENszji9mr1Z+7c5OzEM2OUVSBx/HL+xf8LH7
GxrSehT0SgBIxXUR+sMDqrODmQHY+igEm+pa/yffacpkwx5yraftMOWHr8noIthKf7gCV2j1fh45
ZBSTPvCREaY4D9UzerRuspfxS/9wKFu7g/xVKSVjDytydaNCPUdIYdPhQ9il6w7INE75q7LSA1Ti
BkPTPpEdYWHIhku0QsNQe1zaog/d1NkOgtUbQ9wD7PBrpnk7r9PR3VywVoOdCoYUukUsDrAs2D34
R+wyBrMh0hEDwcOXyYhU5EdrslauGl/grq78CBrhg3NxnDDwe/YD8T9IRRmA/gBFcAw7kljMvaid
LoqmFvkMOwSBHtEGtbN1n43qE7qrbM+yll3kmP1EfbBvNK6gcWvzeXibBDpzsoDPSsb8vCE0rAfZ
tJjVWVcdj9Eqm/wb89Mf/hiticgml2lF6WuMHdVFm9K1whDGzOkCOioE33PEMvL4LedaCPMEUl+R
lUjtIZNwwvLoUbXyt1xhlqcuDpjvVmrqPMgwSXVEMRICEdmumMIGdDwJS+Mb4DC/XuPcLJhHIikJ
AjOfOqj37c5d+x9dP5/LVbV0x1EiuxHc9Rpxei5JCkIUhTzUOhTpficKLGSUT8cgh0dGJbIVV178
3j5evAeEvo9E2xCEXs+eb5fOQgpuKmTbXMJ8efcHEMmW+99/PtHDtBp+xatrCJ7xl2+4Ljm9jfAW
p5zOqR1DF4fJdmbBo9gAyw+WlHoj0y3WNhb3DhAJdxN2X6Zr0fgIvbqhi19WxQRhhxJVLeXPjmir
K5l4PxdfPMUOls8wF99/BRCBUp9ScKro979YIgXXzxVY7MpZWloMDDqp+m4ArusIyDJAmX9TLWrt
CcQwq4796hY+zRKo65+HPSG18DXcTE3mVMS/bep47LHP21HDcFjaaa9atVQlb1ZG5f/sAo1IxKQa
yeJjnDiBl+TbntuRQR5LftrOMMbYeFoJ9tv0qdKXWk20+HeiUI+KaaDaotMGZ87fV3Vjt9HXQjek
19p8pwtWLB5oPaLpHTBfXq+ezE1pTZb6i+LZzbbcYELS9tHjPkLSRl0j0skZ6dMp6MTB+lypXt6f
Jowq3cfHbBfZ4FncUPVCTO6/To/BZI+xHdoXYI72Gex3a+kwIG4TjaWlr7vc/vbTW93rQSDNkOVY
f67FVgiaejLKwCM3U8ob779uIoeTnClnQ7/3FqxP9cs3I2LITShZACLyKONW6wtD0zGY+mHFl6pm
dsk35pSfEvYSVvBh+RNA3qrFO9uoT3rbuL4baT3szJjlJS2hE7gHpdOp1Kq64vTWkAYxyeaPIqOn
sGkra3iwkKCEp9yeBxtHNfAs7WFgUU7SidM7IzFgWq+PuqKiXbvndOy1SUEeq/ad/S7hkHlfY35s
lYByZURG9gVIv8YkzZWmz2Jxh3+l4I841XUNd3/GCI5qXmqEU0UaJZI+13LI5kyQJjwj1jl5x6f4
Wln9o094q/7uOMX41ypJfcSY2dYk7R8NbA1PSme8HOxAgiPDIs2Cp4/Kg129aHcHX/A2EpXA7jMa
ldGDpD3KxBuv+1dUGpuw4wxfa2LOpsenaMzX2K6rqMIQmevbB2A/uuKaKBPPvjoXCyhEUNLfPMoB
4g2YsqEC/L1qCo50idnkOwvLJIeGmSEHvCsw/pGYsLckkpAhqZrAdlviS+OQdOL893x9/P/Q/Nbn
WZFTBK/PY+EXY+4wRF8RkjvG2UGTBAhwYCIiD3aW0838A1Bn5dDKeGHBteyl9W1eF8I0UqPM1d2h
/au7oPLvD/UWkdOWN2vzSkzwcKXx+Okppiq3qC6PNKD6aU8SfA6hgwitPOmL86HjJZFicPwE6s1u
Xq0tPju2v4/fEZVCGVSML/t+ud8dbz2g/azPi4VPm5CgJGFD2OIFz1NHsOdvn5aa6Dyy51ATv/0c
y46nKM3gClOPhwxk2Zmhiz1R63Yh6W4921Ll8Mz+gnCzP8sYUZFNMu2dAJgvdTVP4yedezj6yTXd
YmNfCzUEz4QvssqllkV7wxt045QoXo8UBIn9/arpV5uN2mXMkkb9JrVC7+4F1nLTbhhtyjM4r6i0
9H1IgIto7eQ4oIFCT7Ao4qPOgz6TiiGW0GwMQcwBqqrdO9+pSln62ZT3DBC7zTVJ7Meoc59PCmjX
KQazl45NrL1tagjV1SGp6wcuBmfjy3qY9XPNh7aMqQnWUrYdF833yCR0I+R/VnYEu+h1akj7AKck
7fyDxikRv4GNHQU0UtxoyJIBlpScWvD79+82SBT+XDm85m7N3R6M1z9k6Hnc4AaBH5Xk+6nqqY4b
nsmPDGT2/G2vkM//8qVGUTKlcm/+oSlmteu7T46m14AUNLZMjZaM2WT4ElYN/la2omISJYpU9oAl
bHVhR4dEQm4mhmzrPmkmBwh28XIsvwkwwoj0rwr3hTT6j3i0mbApEGtOHW1DhaWWOFpmVMudyQZj
a2Yo5tW69h2pmanYQn2rTW+tjNW7L0Z3EdxyMmjXf6zoUsPP7f0pHLLFf6J16uLJNXQvBFBELLUS
3RI+fWAKgkR4+bznS9njvjnf5ZfrTWPg5V1XljEZmVgHsZlY3cWKAXltkJqmor/mLDf2KEszP+UU
RX8MvDLJo9Et9v2D+qpMWt95lC9pwCd4KFqWmUOjC0gHAce+ZF29RjXRJilckGv2BudlLqUU9P9A
rF/Ca7a7bTdLCmu02PSKTPsVX5cEaEnGD2a21/d4JjCbFS1fF8cp89ADfv6h3k3YSj7MrqHEBHb2
9E4rP5LrWwDbHvz2Ewd7FFGHA+fHdtj1YVRndMAUklTG5QkbD7FvuyF9MDGKWSGkjBWdqdyeBlAk
1dtCX4UEAiiDYRM/REUAhciTdrmd0+iY2HZ6xEw5wsjshxKVceWZNnY/fzAkcfAcA9GFh7dfw03d
RziIGP54z+xM/pCZkt/O1nLygO0nt44jnArr3rKdhzSK8dyBeX1Sn+62GV4Itq0TiKcqBf1//Q26
aeFLZ/jd57PHus/SSE7RhwkpMII4vL0H+HWETKdx7zfxYew0JUvVVSQN+1Men0wo2FA1Y3L2w7GQ
4Z+95Za21sG+ufDJ6tdbICfStjM9ITFsomutF2+r+WiuIWoNXlhh9mx+PYickwmC1JfMPr+Wlce0
4PMPYAb/rq2NmBYsYZ5KqME0bMsOCrxD0OSCcs3wc9bdH38UiT35WMS+CnniAVE9oBVny/it9iZg
om0fRIs7iTqTLb5ySr6qx32Y2PUcNIau2fcxGSsVYcES9m6NGfRH+/bCg1iZFqmTJ/dm9RJo3aru
FBGtfHKWbdNDH/xuiRwfoigm0/SPSjHtcg80c66laZI3CWS9hxBdI+1EJ1xrImaGRl0I9ptu7SVF
UO0N0YBXKJd2nkXk52AfPp6LXsVtMgrZA2RSc2Ma9MZ3rItdLAdMPDiYrjbk1Kd+tNsip+YZoqLQ
SD2yj4i9dj8oULs8fP49Wv3qBGoSg/C+iw0aQbHJMGXDqFGfhLWsySnrV1vpf11nm4EH0HrrwVuS
sBrJgk15wgJpsF60Y42QIRZhdRLZrLC+RgiEbQ/4nJXoJz6qUNpxCPNWfeXn8ZIznFb2I88ABEZC
CudJ7/fusO3po5drE91TZgnVucEKaKpBdC17bIw4z2ojcC8W3T3t2kAGCj4uXN8QPaTMCiVdqNsU
yQQkMD/YkpvmXpWn50r9P22G89rO2mBhtdOQcBlpHmAfdE4SKauqLQG5amzzIzEVHmCcYyBCSq5p
6G9NN3wXIK+SbTNwrGlP19rm0SemqOUsJrw78xl7ZBZNcsxEOht72DD7FrDmTQcnPZtMqlTYU2mz
vZk0f5MqZ2avXs0AH85YqJpVMp+d+M5mD6O4bmyHnTNfmpsehYDNwOe1hl7DOvHUx/7LMJ/v5O2r
j6pf2t8so0SIHDEClaTl093vZVSHQN3uL0g4bTayLx/pBZZ7fT3YastV9EzC2tLOdJ7irive98oa
/i8gk8LUleAX4RVSRohUCajXaCG8519Yp18+1jPBwiVe8JqsFK87N8ZIuXPqbNI4RQbAO732Xl6o
G+qEj2OngpTN36dTPUuUQ5bitSOL7LIphmwfDdgAlxAHTVTBBRjnin0bCyfhBcmXp8XGzmScdO0M
mIOt5drY/cCA0RJF5dLEGMXsnstRNL+Y5CadWYBZtGq0W2gxtL44yRPMBprECZhc7ONVZOsqJxLy
nMRJ0viL7CfWHudTqyAY/lwFYB9RhDsby7ZPk+lzn8awfybONMr2NzCne+BZkEDCqb1vzF8JIiEI
vodv/w1Xjcsgz04ZP14OPvzD1i10xxZcaF/ak2A4XYUYU1wB92mEPV6+S3O9kl7P79UpsYCNTS2W
AAh5Z/Oa4/+iKs6ZbWQ8wSyw13zzhDbTDTR6L7/KcW5zDrElMGWJzc6l/rcmi6Ojlz5HUn+mQ5Cd
TT0I2SOZTlvI/h7DJFh6eRexJNvNwcwYTgFSSPnKnmm84WcCrZQpxvB6/A9y9LJs31+Nf8AqrX9c
/2ViFCuYfC/n23NeaTfKZPFj5Wcj6bY8xiLxTZUMdcWyStTvn/PWgnBQlVXAFthK2K+dXixNWyob
u8kAbTPCY4ajRylTStecgXeYtJTL7mL0scnSE6H97/8JLpB3BIgjxf13z8W2sKUobnpC2rDMMXLQ
zckw6qClRRngyGiP1xJHGGRWQyoDi7sNlFNvGivNagZArLUYtQm3B1fgzffRKrxkSStueRry8qpq
nNiI7uTZrSgM7s4vSPveomODJNC3XrKKFO67MeabZL8+GQNXwh54CAu6s3SS8bu5pjBwFZqsRU5b
lJuz4UOq6lkeVSxXqLOPIwGdnDHWguhDMG4eChppGe2rkeU1GkeqN5qzoZ8t01izXMh7vBBGHzah
Z+59vwIvVamwFMzVEokRYMWKLWvDmwPfgedBJ3OS5ZCZMfMAbIyD9IOqw7yNsv544uicd2sQXMt2
Dn/4lFKgtFWgwJ+iZyRa3WTQYf27046ojz/twQ6n3aGxj7jbBSKzYgIAoE2ofkjilQDWGw+wvD2a
/gvClArpnA8LjPCOTryx2rBQJYpHx5getkxIFrpUKtkgNjw40qrVNvn/OgP5KAsJpZUQ+RZHMEcr
sjVW4u8UTGTjWKPifi9/45AfU0GItcfDASZ41zboTDl9lc6Am/tR9QEzbKMEJoCdGSmzcOHook+p
8Uyqh0XezVW+r5H+m1bdecJozoD042RT8vy2HrcnekfzUTIueR1TOF+UtGQ4IKnED7AetMhy7k46
mnNh47J9RgM9Yxzz8KrcHXcJOsMdF/heefTgEcoNGV5Z8LyKqc8GJLGcOJa9l2iWmoIkyqmwxsUA
oGBLmbLFG2VQLN6kkXoyaW1yM6Mzqu9ifZAW9KJM3H7W9fdKzcbUV73a624IRXmWk3jicucA0j1V
hvxcJRhaerXHxKziBQ8hzSVJk6N/jJhh4vBkAlyrj9uYXt6FdrkiOMj8OGYo84mIp3osE7hlxLaT
LxRH8oiAorYRxQm/txYxTwuEX72KfuyoNwV+++lkRSyq8wJHCfctqP9aURtp53eepwba6HmnpsQG
JBdMIaSpYuGCamIfhVrUtkOIDLlj0uLbFDTkAnSDZIoE2Bj7TGGUy4uVaG03WEfiy8tDSlySoeyc
oTGa+tN9a49kFlrl2CrFxJGX/eyHK9E2z80QJAIs7S4iAbtuLNjOqey5VFY0NTuToJc91hL3Yqih
sOmoS8Kzgav4DXr9ImzmW0TNP5CY1GPzOzGjRXU/UaXX0Cug0dHKqx9rknvtfspbY3Hrd1JNtsxg
eR/VWe1g22oQ68OFlfRVNz5GSIRONhe2Asrz463cULAqqfzaWhTX0JCb44FMPPGYpbwYn898RRzj
RDCxLH8K1AiSDxzeujHx3JB70DMOzvip8gb0OtX15VSBoMjJh5+VXlKRUIAJSXOx15ZSgrGGQjhM
A9rqYFCOwf+qvxTHk3pIzsxWpSaFqBj0mBCHz8IzN/5ov2LutHdgaXuZCagnDeYx7xzFVqL7eRhC
J1l2EjcyzBG5txpMYPsMiocZ83+pzGbYl1PvcfMIakIziwLUTqY85YrWqyAaTx2/MfRXHVcahGlo
U441m4p8KEaa56HQzqow5gu24tCU50Q//zyHb7rWx5a3LSAsqKySjpgf25bqmZOLfBDrPPAVrIEN
KhCVD6AeM4jd0gt8G95T9kJ8lme4lvksynZB0OQcfQ78NT8KG3qX3DLtJGL72tCaNxiV/CZKq+9s
KKqM/0IWF+sjPa7txkiLP3cHrtqPkPeZup8nif8sUnuddC4QHC5e+z+j51BweEXAoB5wG7jSSJTX
hi3X3A41vM9oAfRgonrxtmZs6GY31+JEpHRZ8U7A0WE8ptorHYaeh3zhgxDtuBmLUium132b26Wr
Go/9TRU7mQvLDx5N4ov3PHVVr7rdjozkwztnuOTTjGm9y83kTZVRUoXGp3WQ61r4zTzWvJQeM8Dv
SLzyAhFQS7anIlWFMfxIW0fQxbjWvFX3s868b7BjFpcd+sSKP//KhX0CR7HMPCxvNG4p5/8QPQW3
07YAaCVWHp5/tOvjBY/bKg2/LS3MrlPkk25HpkuMPDKkX54Kl5oExXXQ7gG25oPdQLPEEXqU3bQk
LqDgNiHczahCmwqtjn+vMC74zTCSd3OZKM9kg8D8otjCbLVXIicQAwmAyI6XaiCPSjTc1HzlY/2t
apS2SMox5/1uOyVfA2bqzmWm2UO5UXnQcHv0naC9zFxZ7OcKVx9io89hO537LFpSuNjl+7KpyXqS
SwGrpnRgpGdx85wjJbabAi1ntLSfbXA5tWPp6CPKe8gKKFNYTF3uKOqv3bJWvfKTXzx0uDwUO5qk
zfMLpDYaGvGjUM6jX6RQYCqZJ9e4AOE9zxWGyXw03M1jtNn3VCfRiwrigaWpaGWRQdLwpd9vuCRH
NbnBXRHgGo1Q3/GpaLMbWefhFmM/Yp54/OC4xvpl6DGCxMa+yukEWrhQxspTjTO8RUswb6nEwCtX
DR0ZNj+J0hOdOJETFelD94XZ8kUTKveML2DFas5A0y5x+cEDGRKgUpyQwLHQkreYwl8zjl75v7vf
HK2GFwi//iHimaGHMKHqQzm7hiseXl/BtMPOIjCsJ4SeI9OdH5T4LeaBIpmH8YCevJiSoRSuX7Qt
kPiHa+3P1+UdDgvZijCZtEnbufXKhg0xJjGbq6aIfEini3s81C6JgrnXdEYNiGmGNO3b0YF6p/z7
JfLPURHIGrvqNF9tF/hILhASD2hBgVEfmd8SthoVXVhKO2jGn3bbpDUipayaNUjBwkn9FWxeUgwU
K9lPrigYaqhBGlktrqWJfPgdYG7iOD4l6gKV8o0zSGBOB3sEc2WxPJYs7ij/w8QzaZ4TJYHSiahk
hE6oQAzWDKbOHtHtK6aaJl70TEDShF7JdOki689o0bVwG8+s1d9PMJz3u+aIzD8yA8+0n4d6+H7m
bvHAnilEtQnvwi/A29GFk4cvk9C4zl1UaF66ig9p1z15bf+hXydywbZ88cazulgyj1IgLnPERzXm
0J2DkHvXqbOKXHxJBGpXvfhZ/CKUpq9P7J/zZ37R3hVHdbKeJIVuUu7RKB3xB7IHK3hJaDJrEbkJ
VgBQxaclnrnSxKZjzmLrdQfQxzZgSrdcx4c+iuDpzjRcRpb5K4D4x8j3OUGRkmbJ8bvIcSuaWRp1
WHXdkDPwxpGSE9QMRPUHvPIqs1sT2iySED3bNE4UR1AlexWRnf/NIW0Jc9lCx1Pmura8rEctmJtB
jD7kUnoeIpKKzxiM8N1sDI5NYVEA1PmD79g5iI9QM4YX9Q9YjBTcIO6G839F/A62P/Z44GGxrSjI
RBOgCU9xq480wdmSiCcrZUP34LNbdAMYUxCBEQF3DGihdKp9i/+hup24lwWlnT8aCOVxYfXWyPJH
ONUKWbjiElskQpg66mQk9A3kgaNCIC5GGMTLVT3PsjicIznwqcXHjCblWKSbKn3Hmgn9P1xnpdHP
JEw6s3LW85XXUNYHrq4iKNXNfbfWiSr/aQGIXkJ7E+gpVts3f2edwrRpar3zUYO19qfyKOrmVDpT
x/NI9yTlZ95xkhVOtBuW2KLVgos3Uh0TgKa1fdM9QzOWsOgBCHI/YNkilEVoDitdDWy6HJpgqhaX
wSDH3e0+uqKPhP+JxRlfmoTszxtsfhBWu4XMq2agRJ1I3Pf0VvuemhKCWDTyPL6ykNvTX/1dx1UH
epMRhJw88GvPyDhcLnkGToPZVvQQmQGZQ2oaIW3pi0UxPGuKtBMUVO10UkbIJ1IR+f1tLGogOh3H
zLNr1BlrRju5ehWYt9z6AZDBtTxreWW6eNnaO72DI/47jtRd1y2zxMO7g5rxmEvPlkJc4GfrWTWB
neYb7WtKrWf2Lya/hflHvMQA/6LfHGFeN/fJGNKBngy2/djM7y/mLirqsNsFxUqfcYKB5qzlytAV
wxAA743v45VQ9bHrhyP4Ygs7EYkCwWHlG7lgzM1lYqeEVBKCqPTmAQq/9VEmlmXLG7BzHn8LOIm+
rKXxda7LXJCjHP5LNxKY490pZQu49RVOdP+rcTYa2FT6BkQd2vlClL0m/2dHp/RswJQPJo1NLsOo
u628tiuTiCwhXuvSyhnxDexcWpA20R/+WVJ4lna1KBY9YgufNscbYhHkan7bP7MrdOd/0Rxgtsz0
DpOWCCVKKg5y8J+d5bRokoT/IuQT3zeicOpbkjqgLZ+98YeU1J0Wu9UtGSb7/H3A2ZpbZxh4uMka
cfdu6RDWKQpvPMHLAkd9gpLzve91gtdJ/n7WeRo0Zl4beNLS5fgPNyhnXQHqC2dYIcvqNnjyLxC/
wzT+haJ5y2wKurBVonxkRd19KbMaHvuSS0gyoTuw7aiQ9kX+Za2Cc9yNtiUDftouejDetn2Yd6qb
yUqPrcgK5FhiD/mjzmRN2HaaYrT5lBTXKfpym4Q/0It4czZiwJ3kr5KdvbXBYfUmEkG/shkGMCBQ
ew4MiH8gSv3Vs/2AKMqHzOGd3a9kPpfeN2wspKHzCbA5buc58uCJ9UNhy4IEOzm8uImSrIepYyK5
SvIe1SbaH8FjEHwZwRvOaTrwCY6QIRe2nJxi4ott11O0MQHx7oLFOS8wZHGlIDhaYd3Svr0mZbCS
O3SorBOAlEIH4uFjT2MPphD1r6JC9z9eSh0aopBOscRtDr3+3tpu3anr4NzoIGxpPj7iZ3/ldDFR
A4TfqFDlQ6U2MYLJVeCnR17WBjDjuXEokauigx6bO/L4YbwW0n6RsOj/tyld7mFqb+m0bZ4rymLk
Yvjwx0V3K2Ti9Y5vGpliFwcQFboY9TRRM+tu0hb4Kim19QcpKhxhUdy51gQ8YXhXWzHBsDVJIPPS
ZFaQUra3W8fNjbuyyRBkd1sz24/tDLzywCsUzO4ho9SO9kItieFrHpx/V5BEGwQhqcjXvF6U5MHB
bZnOD1944o6dEssf18RuggsE9RKfaVWjV+fiKQakji7cO8l/+k7FlLY6XgPllybL3BAlIw0jSTUu
b2Tfkpyj4cqTkJuoTPYSIpBc9XJ5EgGmAFMS/cg1bJQQ/p+xzcPUMEXT06kdsHKrMn25lJDmC7Hn
wnPl73B9zryPavkeFTtOfOcQiul3Uz1GL/jPN2wWX1f0Eau9/Xarw/RAGn3hnRQLjhGuOGFbZ3m0
AWxVHx7f/mS2vUG8ydU78gjienTLSQ+i5ueN4zNpkKUhm3qN+sb6lqBtCByqg/exsYuFYULpy8Ok
aoXxafH8dekSMT1MDInR4qReS5I74T/SFYrVEXOQDmdKDkJxZjWma/ZqTT/PmL4J+rhR7w1zlBv+
Ou7u6d3V0er3w4xUWgL+sFjrIh57/M+zIcfozc/eHZ+XTR+jkZSFdjiJwUEaTSNEnS7y7InBk8se
CEgwwoKwjVqC3Ywl//VLJZgSvBPOpLLGrfNXLxNRkxwAL2+OSzVdYOXSZN/L1UJyuIml4lrk/+vl
zM6qT40XTLjmAnNLuZtnE9CKnI87/2tVxdqBH/PqmpmCEcTI9+XsqOY+I5kB8hbkg56VLKRKcQ3R
2E/5kZOBbA3oUbXUVbdAkjUxDa+2xnSL05Pxg8j8EJ4f9Fasp/krZV2paMHDUggfoY4Jj2pItTjR
Lu/qSCRpYvnKAoXZKiDKvcQkLfvRHymL9ktz/m+/TrcXUfb7AxL8I3LBZynTXgOWTy2ES6mHWF3E
6zP5XBqZCp9yvgdNF/xDS5UfeO7r0XKyxkhONLd3MqwQUnV1mrWtfMh46spoz2CtQ9oLelOmOoaS
g4wDZIclgSmSbub1xNVlm0xsfyn/jryI5fyCHR6iOG7ptYnuN+SIB0hXODljBlK8NiOjZ29q/O0A
wwFgOGlttLjm+WDjHA8LnEop4pmxyCt3WH/sOiK7V4d5YS11C7DJjj9wi4FxvzhOzZGZi5r6ND1s
RanBQBsZHmxqXQ68bFfqGWxWtll8vV1MS1tdD+7TLfoDbBR9ualdvkSNTf/K/xjP1T1SMWJCY5rH
B/ARzJ/IWRZLL1SSylAZWNNFjiTCCfxeiNhezBdQsfoXqlVMYN5UKal2FrOS7DP0QhC6bCyNXQ4g
JRL3MItIqAZd0ZAMFwOP+0JxUCkIPjlS8yjvK8mje5totbI1T1fEj1SHnXloGUPi1B+1c6EM7KWF
s+UTXxVyy4CUSyA9vOeyBbaplFkWOwu79nf78KTWXonpiS35WD+JN4gmIapIgnVv0ArSdFWsiwvu
Tk2VBcDLoRJPIWE9OGKTx0qA4dEjcZtXyEbc/RV9ZTos11kvsta9rjs+Rv4mfNkas63YpUIplfPU
b5VRaLeblvlbtJGnEifL8+PZhIMW5l/Zp02PlrT2CEP4rgdeLhjNjB+klJkLM3G45C7cs6rkIbgJ
/G6R2G1rdHZTuGfphQ/Cw3U9azm1YUmozq0ku6lfcXxd7XnZ7qzQx1kkwhSzc1aX2ORQThBmyqNJ
9L5uYqWR15c1a8UlY1i4fq9F70Tb6Z2i2ubjQLK2/aP4oToStddCRKi+38h3hDGe4govR3e6OGLA
7t5eNcNU/i+jCsIj3/cjhoS9P6g+Keh/UW2qx2Hmov+u6z1IKNWQ0LCJ0IobslJJq/KJ5Vw6sJAg
iwFoxQ98efOToYmX41ht4Oz5Wur0n6U73mC+iBpQ8ELacDwKwpcAVv2MUSTfw3jmMUK2geQLjEK6
gQ1hbRvvG1LRjM/YxQ/bWzr68ayu2XGZABK+HzzRqfejmBh2rcNA8B7dru1+Gs8zO8OPXcSniOxc
yk9BdGA1I43i9Hn3tjb3sad8B9GcHC7oVDMlP8sNXVMaEmvp68tOSQob9qwKAOa5C6EnA81sTPu2
aZNjamaJbgbZpPJUPoesC0od6lTUqzLrB3BXXfb/qvqd9wuM+DyiAARHZzaH9oPGp0L6GIhE48db
Na2D9Mw6pSREf5KiizPgxY7fCObz/lQ232v+FqwIgbo/AJrEEXiecfBua0vjkB2FxofC+2Q89Z+e
ogB475lWpz61aakT5aBf7tjreNBZph1ZNLS6S8uCZ8y+iEn8IGnfbvnIQFcKxg+gwDLrFstmTnIG
JAQ/x1VZBL3Ks0YxZV7k6n7Jh1ekUAfmVw2kchbnLais7SIO6oGkp7FC+pPYxppScmmBzN+iPlxL
gFGhyGFSNy6WDGto6NaTT6Z1g0kAt9510GVkZlBB7yal+JyYcHH54GT0O73KDwxyqbPjc3uh1GTY
yR5ILySiaN9ATdl4o+4oHlX1zVfTElp1qontmu1MziBT+2p+O5UneaIauF6CiystkMoayH9faznu
+YTYW4j22TPEouAED9FRe5SAZYBQbfxtf6cIEfou86pvzZpRdM5VhDSyUb1SI8uYaaHleYInpho4
eODmGaVyRSsdTU81YGWTHqBIPmPm9Aj/55038ShyUgdciQyIQ8H85pMb8GVYgoOWFfwl9BOQ8rev
yXnTSNC/RK4SkFMHBzB5uZDKbqYnTYIGx7jqDpeDvECAl18cuNVLEfcHX595aSd95sokyMcyfs+F
PtPeuZ34uRcNJFCB5rWYIHhQMIyOwZrHd+8vlcSqRBXOwB4Y48wReKxOWZtn3cvp3cEURUJUvMGW
V/01GPKYYVdgS3Xe3S7Zxdtj7c4mrgo3WlO1uTzl4iTfuKZ4o5Qc1U6EP6/u0RXoWjjmJJxAzSwo
2uDkPfJgc3qfh+Q7Gn+mqq5diobH3JehlzhBS3T9KAjx1eQRrjB85KdS9IaCI72tMb1X5hHSxCxu
6y2sT3WceT5HHxIeWY2Gy4F7RY8KxVmscAuRyB0Tsu7KGUAW/gkj0bFS0O4t2wwbbY8duVDD3CsN
4cSrpGOK8lAY2jGtQ6ZBodTRymerMove+sRVIL/UOI4qyPks3OAKfH1akI8l6bhn3xIbmEeeIcot
V1IekY/vDz7O8LPz6w+8rTqEb6ds7oreIozlByUmk55SeffoGfcRNRI6vTpX1wt9TpT0mkW6HM/a
V8jv5jdq53Fz8IybpG4Ss3LCKT4Cc031kRl9+SJkXmFyp4MulNCtnwo0l5k9E1Pyk34izyYOIaqx
JvrLjnrRwbmtPnn8g0gRRS/NI0W02JwNqUs3JyuffDIyGFw3S2EgS22zDpUgyHyO+6lYcvjG+/8o
LGIm6kB5iNVsn6LCIAXBXk6bnq4VJpst1dNELzzimEtxupfUxgLqy5QiGiO23ouJNZF2zINdZtg9
c4eZ3QDAISJBuQdnqXGs/xvwXbjmliqAUPpdmm8Z7aMnurfISGAdNRPp4SS9qjo+gJuGQPyXsVXw
NBtreejCun9iNtnvrzqPWb96wzA+2kRGa9Y9PKvJWIEcH6Sg7wLnFPxZfZNjYnRUfIdUSR3oJjNa
HBB/Tl+SOV6aWVzgc8RQUvfz+dG+tWxALhIu8ze1ZprDpeZF0bAyHAsOlxEX/3qFD/A6dsf/8llV
t/y6RBWdzO23HZzCtVwH3v/EpFUeBQACjkjIj+old9wdDrsMevOqN8+ggI34cd13hMGw/prvaWih
p+j4YNoMCkh0TIRXeQoY7JfUd55Sg679QMhvm6jNVX1NKhhvxew4SqH34HYCizirB6tIxfKcYQ0e
8ckuDxA7KVj8ekt+1ZvZY5pKH0aSdYeRnRDTRsOHGh3h/URl64Him71dRdLyUUPgmGb49cRRvazt
bx2NVYILGp8ErdqFSr0giij3wkiGZ9MP9uU9VUDdQ3kel/fTl64ZxZ9PZQCJBZ7ZbzhTcYq9TIfn
XFISWeVfaTANdfNL5oBOr6yIC94jwYbNo2DLP6E5oskCCSbsFOb0TqKTnFJtJ+wC6x6dvXB8Q+79
kVlMbqHEeJoLzNTQtCOFa1ucDie/2FnTNL2HHKFub0HTjBF3fr4tNGsO6k4indzdPmhe3tZN1XP3
q5PWL4lHdP5YhHbZMRDRdYQmozc+AJnyIKIIfeYUraXlDzsNEMWTyvKvtjO+yssHXh+2CA2IQJk0
MVC3ruGhv6kRaJoTqzkaS2GgfBjFS5E/OlT/1xnfsXov8yJAPd74CeHDOAXxHZcPOcApjqYSplSK
bG7GwqWX1+UmaXjGOgk0HVdGeuXqGDhdmF36e6PJtrsBWdKq8BfLk0NhJg5P5mGXD2yipbo2nZAK
OSkUfgY7F2mFdxxfqafGSWl8e2Gp3u3e9snQyLCy6cbHZZPhdO5zgdET/88WF0t9oqXCNvYrhOlz
6RC4yeEnDhuDceeUJpIXMkhjI3MVI/capeUKGSwRmjSEl/ZlJGDsFRd32WZ/LAlDKO15wWRCs6LA
PAkq7OHRix1NYoy7bjDJniC9f9t0h10iOFJ+nPz92iBsfU6x/bBfPTiYaiACxS/eBots/GJjxEA1
MrKIdebwGHbByL4kmM2y4HJYMrRKdwEeEzic+sXtqD6lzIYDM0KBpfo987kcZ7UxbRAYwpQqPb14
mC46T5drj97yDNtiJcpHZggwTjnb1QzUboTlD0dX3A+B1ufUon44A/W1OqIlozoIW6DRgWXF3wwZ
81ioK/AbNyQK1FmwxIKGpcjNHm51EfP0n6euIqZ9CDdGcSOw2HaQh5INx7T7AzcoBKCs9QL0U3kH
t2Mz3EgZf+Q6e27l65dg1A2/P4e/vHPHT8rhykgJw9IYqS/G5ZZJp990xTWiqY0eh3tY4/FCh1M4
Kwo79HRbjNVp3FRrHTyy0xCO9CIpBxanXqCfGbGWDYoAu/xVm02pTEG7y2Xs2dcPDPDf9/pf6QFV
lXm44m7G7SXyqWX3TNQ/chRYgkkyB+r7UXxpRfVNZDZTUfS0DfgZ6WNOqMzI93/+lY77xLCLTXE+
urujqdR4gT5hEMDUKA6m9rTjZSYjN06rV+F3qxZ1Y6h036e3QI5LNoPWRIiQCMQbE36a2S8uP7BD
wdR2oji4VmEdR4E5plVhKcZWRIZC3Y02iWDfByn4JLZDC9NDBnAgR6cxaWgY6FV8R1028s3AbgIe
y/MWDDTYPu8TYMAfQADOnb7VO088X/EBzF7WUmUXHrM2JiiXS0GCLDwm1dcQxpnTkE9p7LEYIVRE
QFaiq/VbGT+3u/AVX2+X51Sh21YNMDg9quDc7TP6c9FIpfJ14R8HfLBtj4tbQQyPRRXf2TvlFXdZ
vRjWh/I9w0gdE/9unf5Kmp5mlXuyA/Q7kpf/LzyC3++A/nxE55stgnwtKuXvAqusKjn4d07EJT7N
NlbBpbS3DKuj30uk6FUe/cOjqI5NNQjRkf31hTIEJRCJFymcAKTuO9yyOFb5sQo7S1mLpW1IIFGe
yA6c1o94gTI8us65rOpSzufuLKfpi+aKIGTcikEUXLSaOvIDyQqrJoiRyV9nm38U8qQ+2duAvRoA
1AviLKn9DNG1TId6LqY7X2d2RwVPgh/xeOfWlEoHIvFBYxL6gEkb4Ukwgxob3YwDfEpeBUw2pKbL
rHD1fED/Ha7C+HBOJjFqbd9Kbb6cdyxVWkk0R5mDohaG6QZPoTKHS2f6OTRcdp+Tviix/WBrx6xP
smzKqSdXacvJhKlfjBpq3Gea2HQeb6dZtA5gz5KfNKWqytcRiPzrIEV98UZ8GZCIrWUG/ISOr/iI
4oOLwf0hvAT+8/mPmvwGmqxKUFcQjwSceNM+L5G6a7R+SmGakNybuTRU+/AUW8mOjahrXIbHc6Zg
QrFq+0I2ENmQk+wBBsbOtUb2trhHoxtf9pWoHtSz+zgaV8kE/DiaWFBWS0Ypn2NAkyv2HFZ5eZAp
q/apR/pqKyKjJQ9PoR2Q0vlFYJErupVfUOUoZ+othlsELuT3ZxBXvLm079bkxQqWZW8fCZy0MOkZ
WwgEhzrmNChXK2IfCngHEMk2VikqgRg9ErXd/p8zMKyrJ5zQ8FS6D2VAF76rogP+3WP80qoDDV7l
XaQoDXhBFWXNa4XQ80/6b1tM+dB0+nI0/xZR/MosWnHxyC/HXPdEnCISy4F7aeG2R0ZPkckQAROx
kLbY1S+PhaWlVNntgmXzTSsw3CxchaGOwodQTtyplG4Lf+fN/nBclSs6T9nZx4MkNTjwliKt6Srj
HPuSo23gWpoPkXVkvWbdiSgr4MQvbu9txl3c+7lMvTCMjrx2pgkOVW/2PW2rqJNZgeU1Ddd/9vXq
PESvmG5pYUilxWutNNLwYrniQdwv4JoGk6XLCf6M5K3LTvVUGHyA06rrdrScNPXNstyfjfk9iv1w
yRFLWUtOdc92iE+6Wig824NOrR/NMvvf/5bP06kjq7bvgyqpxAmHP09EgWmRO9I92WZJj9DfuVqr
GeDnQBztiCkWYcKSDhOWvyFOv7TT0Z1x3CHgIYMflfnKEuSMajDe/yrvZAWX72eWnt2r9+EjglYc
474xa4MrFPmNMYFUBgRrhkzLlZ9pTiKYjTTSZ4PoyG8EuB1KX4lNaAeb0crranXdkJjucTRcGggg
zrn7Gh7vYT/z99C0Yk4MNYlxrlc3hg9JGH87+2TxYPTjzZw88v4i5mrxKFMLSN6DLecSOlR6f96B
HOtMtJ5j9LZW1oLDZDNLadqEgtWdepTziQ1H6orShjOkwSmUf/p03fDk75nRZGClbYLIcHAro+Jk
lH0joCAytmiJO6b75By6M0apGJHyq0KoGXGoJOtu3e6Ih3nmjSqbi7TP5KKgWT0QIjexWyCnQpaC
/jty4m/dk7w2To44K68HTAfOKEhAm53bZRY4J/oJnN7jEylR1iU2GXSddN9WtQsG0VbhRjRkihnX
ddu8i+GDC9DLlKCXuOKz+X8Ae1BT3eBTnb/rnxhUa4aug7JLqdJoGJz9YXRJHzX4zfPYNCALf6vM
FTVUuGCQImHQ4l6HE7k5OCiEmCTQfq/pmIc78tIR5sLPbOmTY/UVhVM39lDOjRE97dwRS8ZFcgkG
73zS1lafkNaNJcUdJSZHzU74VbQsK+n9OqsWOsYQrbhRKM7Cm7//buBByaMQvB5c4rl4taOHU+Fd
+LaPcBd0AxCCJNEZvW3yK+tQaUPNP+ipRBEao9UUAXMk8vMVdlcCU58tYwRG8mFaD7Es0ipE/L5U
qhNV9eSpWBfpKoyXHdzNDbBs/zvJ6gRpiG0Mzjac4ih9jw8M6UMDcS5N8T5B5GdmDqvw/ON9CGJm
GAv1N5fjjoim/CdgzfnttcVOWalTirlzQNAigW7G2C7DdEzrI1g8J2GLTpRanE4HPgDgt4X0V0us
EBKJ9AjCHLBkKcMehislgP32qGw7NigWqaev/xs9PX4nunu/rDAkUg9nUXqjSHBqW4wVH/rvGLJv
xuSzNKv4JN2Lr11U6DLCZyOmupY3bDshwxL6iMR2NG3GxG2jEi3qoyE4XTZgKQhhsuV/fzlOe3Tr
WIuNTlLxcs9pDVB6uwLrhaQunYnwfCT9+VNkWi/f3+eDUHLo/CdiFFwYHHt52MXO/Ehr7my6b0L+
8cf/OTyZ1EtUq8hLlMDRCvJQi5MqnPOg70DV5cEv7Dn2kg6kkZODZ9S5zGqBxH5Lc9Rs9Qak0kJl
SUXdncxE268QMM7vyeFtVl3CYtXeLPQHrilSkBuv0b+194JoL9NK3y4o1hqfqNX7e6zjWqPoD7e/
M2qg235ZFc1ynwTR1VCvYMWonjRAfMQgAK/2ZxoaQWcCHTX+EoWOxkbh4WBBPkL48BA/WA7wpd4P
H3PF+alekz4YxOzVylOppg2lfgCxkMKRk8ta2Tb/nU/oyl2+2iewBAeJcxtk63SOSaCGIToPWTf4
zB8ISt8jeswOEw5w6mUuxp+CLyRuCDVML47x3BdQnwkFDXC+TbljxZiR/ZnJmXHq0apol/i0LcvD
tLk+aBJ4SklSLCi9Y+iDhvKIbLWm5jj8+LtmOAuHyNTxy7tRmhgNwCmz2qCo1AJRiQhzuCzQTdMY
/T9Qfjo5PgAKmtF4o5EQYKp6z+zq71YE6GVgf8O7ktYwa/Jc+ecndzVc56OvkqBURWEfNv+tiVda
QXOi7wkw3L3rHwisSfMDpDTDPZO1IB3GXIPemJ01jJVpC6MhfokAXRpXVLFqnXEgcbKn9ULEqgmE
oPxCykpJmaflmtY7R/1qgCNjsVexELRdCq3Vbkd/kVUU6MJecJlC/ljcUe4//8VDI4t37ISjCNbd
scu4icKJqCB+Y5X8k9od0um2IX17XU1WTHaQSRp+sZg2RQ5EfFwdkm2UECPbJVWKAJmy0UzqTYCK
LLso6Jq4IkLZoddy4nz95QbE4eL7TmGqIAC9N2aLZ/as/Fj9U91/KRDfyAd+ubJnEuOeQNU+fU73
rRNC0D+gJmmPBpG2s3z5c4xOC2I/YFBtO+S2Yc431Lna94hRrIdt75IGEPkAr+yw8XmwC3hLpxuJ
V9v1XANslF7Jme6KwCpj8Y+bEsWb5Gew2Nim6oH00IbdkghAdx88KqCnnLB4F7nsU82ZAOe6QA4Z
avKap9oIje5O/IXci8w0dgCKc37I5Dn7NPh9HpxOzXpzW/R8e/1zFOgMRmyi9Uln9XdfdYyx9rTZ
L5wJc9SLuX+5N2j8Y/l6cVOhy74WsJo8JhojPbLz/+678t5qwnZeqJ6ndwAX2g3D+RHBCyqD9vCd
YjGEoM+4IegAyt0HJ70IaKKiTJ8bLEGgTiJ9gdKmXO7o1qZkdHtb+zQ6NFx70Ts1lcXtCubAIA6e
rODEvQEkpHA/SQE9M6EgvQAkkFI6MoF/P5l4m+CxhYdfdHr2oxFbY3kMrJ2F6c5L0NErLEiaUh3l
D356M99OWQteolBYSsH3oVM4wW3/yR9WOZTGpKjLdlD/1byX+GYbzd4VL21pKDk8WeB971+dq2/3
4wJs67VryGoaync2V0QnDPaflksPaXC6yc0Gcr/2jp5EZvQtAdDtAP8DcX9nM9NIknBlZNaGsGjY
a3BTGP38TKTak7wDfZxxg4/2hy11hL11YCQ6yKpIIWyCDhHzrKrxC4+mdYkNnH4FxDeYAkJ4G0d2
QPWRFt7smLvHtYcJeg7UCUGLK84VeEbklEsYl36gUiBg8YaCKLyLWE/cQ5wVmLVrTKA4MpsqzFZi
PAYaIkDkH6B75T7YzCMUQoEfN/hwjh3xvdfEnzY1f+tbIo7yisWMcxCtuAiUzanoICdpgU2/J+Yl
VROs3s+kgDbqmXjS3GQH2E9pu3TnH9hM5a14jMJUROoLehRTyeNcNjEDWge8lRFyhKrdlQLIU14h
ItJKRFr1z9fprsNLQqGL25nN3Y7wHsIOi+Aa31j7JSTbxla+wY51q9hvxR0JxERog1EnD7d7bT/H
xFMaQW4+nzkMIe1z2x1JrzILlKd4QW2zLLMKhjgP/lpHg+GZotaCg2Z1L+ez8Kil2LTwIkkp6I6v
TtQyGUkaHPwh0buHZslh0fwuipxdgvvtJB4GYPbnQEOr50eRKEoofTGeDfPQJD8JGgIdRByP1rNw
/IkH7h3jlsuedC8jeN6OywbV1g8O81XizAmdBR6q7QlHUgTl9LQgVj9ckdA5HN756AIdK7LI58rT
cfLQa1UuffTUZdes77OwBQK4zwLjm4JwWLazhrNYgSbX7l2takiImP9lF5yNrJqTyqXg+bxezR/Z
NC0nsswbLJMit4BfUyRZDx3qKYZIH9lhrdPNLk2YqgDQFD4BtR5JTvpvYWbqtied2d98WPzA/Fch
69d7KzY+YLIe3Cvs3iN77rA298vNCAbQ8rTctsSQTVLW3IX+VqGkLkneugx1jzjk/txtqFx6hVOk
O+ek3enStURQ8FrWo/kt2OcFOxZngT45dTHDoNZAh9AWmFIsyYjDJ8KaCZJElCWWTQfzyHKAzS/k
tGewu2XZazOy0pVf+E3bfpOUQGGgwUarflBfpmAtPjLDhSsiIv5G59spjqwau5cGhtuQOlwHz+/H
E83tHvriY8JIciNK76okEmx15gI+DggIyWF4dfSoMjPxQF0YPp3IcAE93OJR9u1P+YPbs51kNlnE
vhs72qzQUSmJejUWwNu6eSdD8mYyL72Ie7g/p6Fc7iXTjWlQHrsUkvttjvfI0yD1F75UqGEXpNFR
jkG1FrFsb/8chzC5tyJNpwPDM6SuzT1izvo6kAmmKHa/kOprifefUDzu4qRLIEjO2dbwZicmO9ZA
XEj06fQKXucJ9FoOZyl6XnWdJz3dkKZOrM/btX0gyRFmImr8RbrVRJA7VJZRFiMA39rTaMf+aYm9
bGapyMHtxY2IxV2lsmmeZFMbQ/bEmzYy13+z0woTJcD6E0/yuqOXJapuLVQUJRpD0A9BzLmcx6Oy
IG+7TvT9d6jlIwuXxhfRkkOcOqLlBo0FYKzdcgwqmgCuiYSkYSuVeSSzVnJA1+p487q4gmu+Pp5W
vX6wRJlR6sXH/jebBtTn2HIxru1v2kwrVdzwk6FUfhTB5MUrKpZA4T5lfftJDS2ZubRctSXe/3oN
YNk5yZcFJ+m7DgXNyL8ZCEehhMCB97oLIUfw0QLj/hDf1prSIO76ayi1qFMkxnIEBsm2YQgf92tj
V0t8GdOiGK/1FQ9fsDmD0X7QK5TqrRIf2qsBVDgjhBAasM/0ngUl5CpAboAtZ6f+nl1KXtDfJycf
n63Lt8bNHtlAaxeUyw9mpsaolkcd8lQ++1sYK0ewXlW4bsckgOm7AP+GwUqh8n5wBMzXNrx/rwjU
QDBB+wjOL+egmnhNMjwMp65LMhRVYgvvffVTc3DuzxwgZXFw0A4DWpK7LPHrzr3YhHzvfS1ZpX/U
XAG/aldHuMPdB5bspivNQP8AGABJs9EPcYLpapxufoVwn3rTNohcsb8NXeuPKwOkfw+V5jTlDd2Y
dxGJdR7nCG6mJ5tkzyLH7K+Iv5E8Qwbt7u1McUSoPBA9ndQX1eV0hmfkwocKWdTKgbEQhkFXGA11
D2omYlRLsql+w0Cel/eGH6PZb8rNH7SCDM4+/M8U2euLoE2QgzTe6jDn+0EUVyX8dHKlRRb4KQkh
0SWavumy21a5fGlIu3I7Th8scap7ks1EqDdB71DBuN69qDuyiQZW8pvI6lhpTtGBVeIMYQpNNyAq
2ED/bZ7LoC7egGYDc0qUcIkIVabD78QmzO/o8cT6UJImT7NxGBkZojywEgWIMYiyVAzbrzGvkohL
nvzppUQt8gL6Fu8RSy53nOsF1/WVQF9/p4/Uy09/VJT2f2/CkHnDDjSUPDDw7nzIYS6kpVCkBksP
V8qJzYnKSRWuGcXaA/ZUn4t9sVzYur5rpDOLXcVlygo5c1mPrYoMrY1VTG9mJ4n/FIXccbby1w4B
vkm9yDc5zG03hlMZx501q5iQqdso8O8ND/4wlo5940WidCc+5ZDKeZ8+cJcpeORkQO8rvyNlcR0V
uXCH2saDw9Mc1Ydfm3YjCZQbmDrlBhhcZC9NTEhuJdGXk+uThNqGVlFrwibhG3WT/ILweL6T4OJC
XXm3IDfmj9Q7v/ba5oEUXcqM4/6LZvKjD2lU+OBYUuh4mLkGD8l3pW4EDlcI+EovvPkDuUaQrF9d
dWHaP/cSLigOVOQEBTNlARZtn6IFS4Z1+dNpyohWpchFsSy2fba1EfrLNBFLa7XsHRwQBEgPRhgL
O0h/s8fxEc5JzHVNKWdv05zC2Xt+jxHi9u5fyOfNnHG0I9imKjlVBdTjucqa14Ncr+ukzaA3OjL3
yTw8nM1sjSffqi9VodvL8iGcjdbE3gKmVond1rZ12kJiNN9KBVLEgloIgG/uA9M/0uwu4Jj7MehR
+aWUsKi9/PWCPw8lqh7CjbWqsjGN8bN8XuBgyl0zXzjj8+2I2p856KRssnGMzO98hrQf4VUIBKVT
fZG4lXTKagUVuikgP9tGe8k2lXsTz1gLSWYAVO145KIUixwWh02E0HUA55NCfU3LX3KB/6pyKcyY
3HDZILFMfIWpllP9MDRqVQIW7zacznpH//wRXlRF79qlueGeSoPYfUWw0tV5m+PQ4DWlFG3kxCGc
AGHEZdA+b7byIt8EWBxUqb3oKekboWNuNIpbcRMThixKdkj7j+U5PtkcOaIhoTLSXKEariq8VrBl
4N8Gf0Xpw/DjiFpBbNLEbQQHr+ipIiTRHGjGFoMXg/HSBzCOwe4MypI24vmcGwmS+pzmJ3P/LNs1
oRtNzbhFD/1oOQhQwv1B2csbC1AYxmEpFRxjUx+lFZQRuz58VggQhEvTkwIQXpZqBfRQAp+UhfdF
EQ2Jv6bGw/rujsoi0H79tavkvkTtebd7X9NI6SfaDhAnYTkgNk+jAXSt5aF5Tu7pWtw8rS3rIVJp
iU1UdkNSz2RxD6EVJgcFbTBJ2IMsUj0oseIavq2n57NkWqzilAu1eTOeOMWP9nZ7BAOmmEzYWuk6
xJrSntQ2p+u7K/Zgjx/8/MCfT2DyWzJ6jvgim7gSGyN/cggg7DA9ZNDTXp/ZWmCWmZ3PjQdXaImr
OKnVDLZq7VK2+Hd3S67ALC2UNXrDeiSyhoizpUL1ytnr8pBgz/8UXH2FYXhggnrPtmfxLbGfmFFf
MTxqAl+ddhpEs6mk8jPbrmo6lTbwlFK7wHRfmAKRqmPRyKPBgtvhonurktHlNKOvI44V8Q+yCXIk
XusUEXcmEm31XwPoeW75hHSG3Xfy0o7mnaerodfVd3vsOcX6r/mMb6h5Ra5r0urPTNbIc4LubREw
q1lMmqAIA4QememFq4HnJuJhUdAlCvntD/7wt0/XidCKmUVIp+J2Be09BgWr2tmu8ZenTZ7AU+gZ
P+8jfJSnbwp4TnujOTj7sckuduQxAS44gyfhpIde5GXmAQxap9X/KKxZ7Fhb6WRJhSBHgE3T0nDm
bnq1MF8zpStmSPpzMi/A84w3EvRkFnDHlDvbTDRDP0Md9DVdZ5AN37C8z5HgCKJsfQn5vj4uKta2
pX+OkxJejyfjVRDCs90+dnyWcU/5KRHpwYExyBpNRFPQfEVk+ua3dP9xBEKz7wyn/TXx4dOzwIPV
zGsNaJoowCSsTc2OL/8ejIekQhuzbMtKSLXxibaZ6tB5z8pVQ18Jfw84jFmHpFb6ciduBiPOUk4M
odsid5vF5OW877ZYFHoI7liBqEFvPxjR4Lrqt41vAp4oH2gv/o04raD6E4n2FDIOKzX51xmIOo/1
GKhXj/rfAvyHoz2A0XPU7uPmjqeLhj0Y4TohBuHBi9Gq6XV7HJMms9iBGKkhNOOK9TLpG0wKuB7M
xk6pvos79F4fzMhdFPnx0zeijJ1qcsBVbv4UoaBjig5TgMz7r6lsu4qg6qJbeyAsLZnyRynfiYCx
qujmK8J52veNId2B9j0WmtjnF1M3sqtjWw67tGco7JYA+2KZix9mRKTvKR2YIEd5lMyf+g+jUyPi
NV1lnTHbcYfjF4QvDbuCu0NsDfCr0UMTxNGKpQY98vGc5v+uzE445LLHannanlCwVR1Nggj0Ltxk
QcAWcyBcS3oXpJKerNhcLUI9m9Sl/9mqR89nu6DVSIfzPDa4KdGflyvmkbGdItIjHSKlT1aTa2X8
/66jca1fu6OO47GF4+5DgPb37GFQHgouZySytvmoP7D2Dq60pvEJdPX/yPoVMhwALcyz3gFeYMW9
fQC8SjoTc0F2gTqk4Bb4Ii0ShoIGrxyVF8PJLlS9sS/0/1J+XNBTbo29kP6TosjThLpwgNGfwiW8
riAQCPoGGw/DmHarUdatISaOPQbGrQ41GGtBmawOOj37le2KSqArduvpAN/qZEyd1ILRxuTpi3Qt
t838nDlkP79RRWRcQ409FSK0yG5zj3ZolqxEvArJLs4JenYbTET+XqW2GZn3IakuyxfgUhZs3bGU
IVHWxPA38UI+XcyvewGrUy2Wzoy8Q+QZtlrWh6J2wUFHQIsGgWprVO0RMv1AFQ1LENweBaX6UTGH
I0OGoWhFP8AJiU/tNBxnvOAKrP924ueur/mFO2cPa8psbSMXFvi2uP1H61vLC3Q7bFIq/Z5FZT2H
UybdEJAhSfxCeCriltMax6Ke+Elr/T9ZKxUwVI6Rx/xNgrBd2cMz7kELQ+Nkk7pG6u6ORRv4R3sE
XgIV78d2ECMN5fukBI/8Pa273xgVipQpqzRyKOYVi0j2BhlPlQ21hG2XcXrtnfBLmKYUCsePCis4
fhT6qjJXBrQpXaU7hruOZIf1XfyCf4WOFHetAuf0pbGuMuZdHbTCIWrzc4oNBFZ/zYOmtTAlipuw
tZr4T3gJ2CaEtrG+SWh/2jXplwYDk4D+b80AuCxo42Gdtavv7ejSAFGKjeq9j78z/q6dKTMGSquc
hLXPw76mOqToVBgtU6JEFM35tILqd9l6jYKJ0x2RcSmrZLFDJQOvweXlEmN4AJIY8iAicsI5hfTc
N+DKJDxp3K2peAJPXMVn/3JNQN96LckIjsa9Y4hTFvEBOW7wpkRWebai49GjKWlF2YCYjLPOepXv
1R4yYeIBnohgNKGBqSNqT+eM8/LNXT8uHnUcUHVRYrPPNJywEjJzYaUJpeR6X6iwIu9Qa4rW0xh4
omc2LKW9b64n4OgFdwETMgU+++iviyDTly6AFDq1BtQP97DTPfWLFIEss/6zbtHcP+0JFZyg7Exj
1PsbF7TBxpnvxWyKtYFSFJ+6piCSRWwTm5swZwLDQjfNS5ITB4jq2SO16S08Ymsrlj6QYLo4Wowp
p2OY1EfloP4N07AL1Iyk2MLdYvxrCt5NlIIg1Rv/e975pCUCbEWuCFR4sw16VQRfX7/xWQ/7FWw0
zNBKdZ+10EZk+ty2uNI9B3IAwBH0zSvFqLyS5YvDQF3pQdJQwGZZyUsbyTynSWhmnYbHzARnestc
Z1ck868hETu1+hyGN2U3xaeSu8qdb9g5VU7Z8xkV3mfSkr11IRg+D4K1nmBec2d+0ipEY7Tr2QJl
QYei2reHL6v5zfvncAumiBFK51UEYXz50Duu5XRJS/c1f0nCxzdDiSoa8gL/uDDeBr5qo0+7TgbP
OkeEqkFHfBop7jGr2hCFoGZzBYPgrE7m3K6eVQT3plwMmofQn4Lq8YBrXbW7fRMl4IrlDKyB0Loz
FZoSnt1h4JcEtLXLK9Ll+JGXv7GGqkIal6gxkA+Sv6UsJ5nBegI0WJuJC3rkEYIF1iyhTRwMu7d2
2oU7v0jwAESri7grhfxiqTdoQR1q4GEuTNu+4OJKDGQN4iE82yKLZIxblqdfhKZciWr1IUyih23b
LoWDQb/XNq9drYD5bEJ3IfFKJx4ObCp9/u0CMCpeTTTcNusmPR+1FVjanxcq9hbfU6CHviKFL7pw
558qrmyQS007Bin4nLEAFJKdNzpvDmBoi57MnwTKPfOpqJRtJiwljxC2AWwuYbyNuqvt1MKDn60K
2wkMU11F+5qxMGFdiZqmdl95Jjfznj0ivsac9TeCDBKunz/sAj5MEvivUFzXgj7MGlOYy7WKEoMY
ckOoemcAehc55MDUPrRY2ywznCBzOBqTrBUtzVXltF51GN2mtNUau9bW+gathrgiAZUyXjHMFAUr
A5uvOHtE1gaGsHr1GoBR+LbVjgGpgKfaIZAjjqEvbKOXZRATKHuyVY0YgZ9wrTaGyGXRrO+OVIH0
PX/vNVwzwE7TCeEMFX5KaEhNQ6y4bgufxNLrGH3B/s8+HkZ73lLKEyhHLoLZS+S2X1bS2X7pCZiA
qN+/UX8+bZpoaq4R8Cm+RP66tZcoEKaTr89Kvlpor+cR6xBm8eomoMSfQqe2XWZRZLMvpX1b6PXp
HG0ROonCHPtnYU2lE5G2nufcEiAsDg7fI9d+3MZuKreCK7b1YgxdSIIa+b2m45kDLHWa8o+Tpgbo
1VO8LvwQluo7mZHHWR8k+357nHwROAtzvp4pfREbQGOq7gGr9zko7h4MHEjtY30R+43JJSmeHXO8
Iqj/RarBtTByiLoyvnw8uGFouUBjHOdksGsAawwR4BvgAa9Jr9rdKdRGKYOScMsP1wYLqTieezoo
06WRyKXOqMI4AXzqcpzUEZ2j60uhHbS9ZhVjIQiV+db0DUp6fg/WLHwaEAwXb5TR9xg1Kd13fcZP
JdmwVv6wsQjzI4yWFBAXzm9NUL6m1FaJ6iZMhuFkBqn85RXmHvpr5gySbEDXa+yZ2yV4cIXu9Lpr
tKPirGeqXxdZnOf+Ubut0wzMnt4j0e9uMg4rJoGvBcRC98P3LxftTCsZo5Hpbj6tN2Zq+9k5tW+W
Lx56XUF3vThZdtLAwsPbQwucr7UY98dMpAsVyoWcoFsIKzQwvxVe1P2inxFIOGDYK+eeXWuj5Z8M
FzMLPwiEhzhFIwwrAoQqG8v1v9LDpRzq/RND9POtbu60tKITxPu2827eG+ai4ZK2w2DN54mNj+C/
XzyzrHtQW3qMoXMiPqZ5+diCFrbIRCzJ5b80qE9x0u343W3MpbdCmuE8ebQPUveIGYvHNG59OvrI
Tkgu6INLMZCaGEaHkwgF2WUIHLeujz7n1hBofAEA/YRjYfWSAcz4g4Pk+1QGx2zMwZ5G26Vm3LW8
Ns9S26l67ZAnQY1xN5UHpB8UnXzisUkGuLC3J/zbe2P4Kzzs5sQfADrGE6/te5GLIoDJbR1R89H5
uLTMySGJ5GpSIUEBKi0CZIfvka6g5owX9Qbm9xz3c762WaEDRBmLSlgk9+2KzSaMN09nEJ1A+V6C
O/VlNIZ/ItOLoJkn5fekwhwySaiE+4FSJHkuBPOA7fkGxcuFXXHqmeE1UEWDPqsxQiMtG00VjSK0
DkkkIPrt9/GQdhImoCzyDAixH1xT3MkItIPYWzpbOKbftVTNojnSTQRpinRAmQC36C+k2tw3ZM5s
u/B6DKyEYmsd1fpYWL8ueHFiV8HW9gMwd0Ey+rM0hoda4aeEnXIkbUeVxsq3x2b2ZZADNYmPZhcP
yrZPYehEnggvCfNMHIInNefg6COcuOOgSdjHr3z59Lp4HU2+/9PyN77N5vkR1qMRU1TA/ojSEIF4
GCgoeVvo+23yHJmqOH4WYwbWuZctHsIfnNbRnLlNGduAej3I3lgfLzMdbhyN4OAkDhTshc13UtLy
4d53kNRinlugTcK+4uN6DUw9Z81y2bWmliUMjYRxxzBCCTPEy0Rph+nAyB609XlKBmhOq1+6mIgP
Gs2QxMoqs9TeWg8s8Q7OkWwg1tHrY8GIJMQdX98J83TTl4F3ZXeISSTEc7GsM4APFR8kYeYwR1YZ
V1rqalOyvaFdu0Ar1nuvy7n0tAjLWdD5oLafGafnFZjJ5yZKvK6Z30F0239EHE+DMDNO+klFybCN
pr6sUCu1z6l88mbXrMIFAZuYGjPSadd2vyrh/BDpoJcl9ljP+3zYVs/vkiMFZZllZ6TDqEN8Oxbd
w/oDOzNDLlvZvIxJHMmG/I1r9DDiFAwg3pq0G72Cn74pFDKtCKEknT1J3oT1Z8pTsrKjCX+f93RH
4w4KO4pX1iMEcS4fkF7njWkh1iehGykpnvhaE4o7WlbiHtDFTUKAtRwJT4suDel8VPpDPI9ooVnl
76ohAPJDmNUR7uANVYNahOGWfEmawIhGm4Fomul6wHlZAbjaHn/GO5jEp+rVT3rBtVgHhYwoy5tP
1ross+RZO1ZoYbv4PULGr6e7TTl0R8Ts2Pqzk0tmuJDrWkto+EDNSngOJE7i/Nu7brnNL2unACme
Px2QB5qwdvrADfNgx4PMLvgzZIGwgeTssBptive/8zuD+xKOWK9jQ4AiPS1UG/Q1TMgrnxAYow/k
e4BlzVjrdEIbjfvJF6LvZGP8rWeKcGj4Bpdbe48Si1KHSN/6G4jVNyiWaB8B6xlnOcWolgzuWz4h
mSx5kRyCs37P1f7oovJnyMfhlGlIPHNcV68IB+fVQwtxA9wbc89C+y+TAO97itje9kBeWP7I7Pu0
86ocTvFEPUXHQrz0n+ozKS7e0atUVoUm3aF4UHc6ctLCjFbbmZ1uD/HviOvlxtl0+QDJ8XWuAfiE
wWDTXWgmefv4up2g2RkBwC3z/O3PJyYlRUhVkTcbxXMUCVKEXTCxfJ2UzEwR4TcLlc3j+Wz/i+QJ
FS1GekKsLyrdDiKN+B3gNKh0dWEG8aGX/ZSsar+cVm28KlFDbHk4hUa6y2E+ePn5JF1XvO5F1Wjr
WsJVwJ7UpngH/UD7e9kbpimsgBDmPgXaajPJiXbmG9Ri7t7pNWuxylOqcxHCqJOeI8spp+gq8gtR
QF67+yclVEdmesxSULTY0nAe8F2r0zByLok9Y/vhwR3uLsUQVMvNxKmpcLuFS7hgFP/kS/o3SFtR
3okMFEdQzLUQmALRL4M1+TRpgddl/XnNOitxIgCmZpT2d1JFu/54qaUsWaVtfSzwJoOwgh8I/aW/
vVadVg7w+JedEndMGRPdgNeKO9aftolQ+coQ2YrPEVTM/KMwRB/wY4cqy0Vg0vVp9lPIlBem2Lvv
pirPSrUIkcDpHURMmZeNrnMOXfEUet6gV1kQF26250vucbkCDbTvZUPrI9Nyq5773UPbIIj5/gdy
X76p+FJPt5/Zr6X+mlyywchcsWI8GrExilD8eR373gXbOJxQbEuUSBe12ramryL7V35LZJuTbyGC
6hpswywpIgahLW/ZZqgsW228+2QnJ1zw+FBZXd5kfWVA+ovR9pBfzOIgtKvUpHZNzux8A1ZH6uij
3+P78osgSYr2deO55HhabsMMREFqKNBKiq5nFNpW11o7q+1eghmDAExQIj/SXfb16zS93hr9aSyQ
QkA2D52kVksNJmEHlFG7vyuckBIjxuG4J97AFXZ6K8J/QP03FdUlGPVC06axC3QHTBJMhI0+5Vkq
JopvGJhNzdyZIkw9qPRvA0JI2e7Ac/9KuNhFg3Wlu6pRX6VfUVe6aQPEcjxYgWqsAHZBp+MoPia1
t7gsXF0o6cYa2wP+QU82vk756q5y5J/KnigXWq6yG5Fqc9ucBrNkLBG6xTrD4grMterWPd2J+JvT
rbsG/oWoTSuuNpNoB8NRE8pd7raVxRjC/e36XLoXavc15mxtJvw5kmQocMfm+FkHVf5SyyDw5eEe
TWopsVWct8bFhvK9URhIRiC08CCwQy6OVWiqr5utV+/GUrBJpWbOjjR+XKm8eX1TeSkNnXcl9s0W
IwbAM3jQwrmps2pIYqDHH3bdnuHX84FpczYV7+2nb3Q4fuPm7P4h42PwCmDVcLMJYJug5BaKO4RH
/TeE9fta6Mr7xC5zuowqipJCBFpfQWjGXWh7ziVzsour+vI2VnEQZ0QqkI6sVCXA2f+6zbS1I7Mt
irlqJnHCoB8Eyxa9nsRlsLDZoOPu/js6JGO5m7CCmXXDVM9hTV0PdzUr0uiqQMvpUEFDwfoxwGeq
j5kTnTfpMO+CXYu3UAhTHFY/CkEBtNC/VbL+sxcSoj2JIAAa9kwgLPzX9lTjKZxJFe9O5GCuzP5m
O+Hs1TwHjux2d2XdRVLf25j/haSk61NCnmgfyUCYdmamNpVFYuxgGnPJk1c14ha+N0Xx7SFqNJtm
bNlp7Dw2QWtgbYWkWCLs50E8t+00j8my/5htsQrNTDUL+S2VJvV3mbbD96IaEwWx0TQ0ihGexUD3
OHwzsZbg4XPkfPvgxU1S1qKb7xJsuJ3RqT7ySADbMFh93HA0DxEfNScEuXGv09cktweQCIVWVllw
1WkIjdSCsTHPo9aCW05PjMRg9IFWngUlEvDGsO2Cp6h0T9dA6GklxVeiryGbZHv66UF+IP5O4AZH
8NNK5ZpzadRClUHjAzv9bYuWSOXUUjjZEam+PL5dZQcoKPG1ECMcqlIGWHreJHuidH52Rf3wuO88
JUhfQWUxLmpzYhgfkhHgcyC6U/AEwWQGkI9FDwyOG62HNvlxcWtRIpu1+RXUPtmyFRl8I6ggAgAl
nL4rs3cLPtdofSEDqHWnqOe4Z+HGMcCfsOs7VHAPHxURDcg+UW81uPG/Vk91LVvaWhXKXzMsWfKK
0aB1dajaSZYiMfjz2hQ/o3poEn4/Ghi4+BZRr+S4PKKc7qaxHs8tq2mLhaZ7PO1ciUJl3BrrLqZ7
iZc0gf6v7ozh+RiLnE3z/9aNJp2WIMP6MppBnssh1SoOQ2Rd86G9LQfQb7KbOIOOggqqH+GFdQAg
CKS6nquU/n1dK1YQkBioEtsTaRcY5Ux41Ooun9sPdhrC7FigHuhCrNFqfBi603E9R9usNCEzUBXq
RLPlvipyDxObsQKJqiHyMo9mjLPomF6P7cFgRi6y9nohaESrghc9Y8ULYk0xi3g/ZXGjbbQKHhHB
bKFyw5hgwjteOe8Qfcnrm+Lpo4Jm44+veTgJXZcgIyL+Lufi1ccLyviSsk0AK8odTS3pP3KApI6F
9ntDjAZm7uTHOUwuC5lTJRDlfB/sA65orhlUb43M7aUDUgcek8EngPHSnq1zpX9bjb+Km3adhcTc
fU9MU9jIVz2fZYSu36fgoVOqUJfshUbIq93pA1GCzmW1rSmz5qz8v6Z72VT7VU7TZJJovrCJD1rV
YgjOkgN0DeqK1vvOOOCDgXz/lrYsbuFJwunnvrHUYAMI9nkIbIBe+CPajFU+ucUTFOVYsIYMSrAL
Y+am4I+889q5KWcXtmR8OcbAlzGEWIY7vffqrIjyRqKO/tp9sZsl+L2TaCQFN+/yD9RVhwrMNj/D
6gMDwhfOAmOFZqHaGK/1ureaarf3uonhYPNG+/iGsnrT9fxR7Oy7ITVwNy5tCfwFW5PRBeOeSwrO
V/f2bP0UunIRrZD4t1OOlDZUuiGRYj+Ps1dzXxTIyygkgQm/clkLq8Pfzpp6DRxh25v9yi/K0Ez3
qhqvRjCEYHRtKP+BPv2oX9Xh6PVOTA2tuemhKclgw/pHfTzD5RtVIF833oEI5+dz+ZaD8tvW5vvo
TIaIVnxCSrY+aAg6oz6i0KP7ghEHjIVNMBfYA5TDBD3saXX8LH8WeQb10342yGf+gMY2oQghUCUT
u+Tvl/TBs46qNSA8faN03zPxbXqUrx64AZJHIh7dVtPkdg7qm8cL/1r+ddg2YqmIv06eMFc/0uCo
cfnMMqXLJKeRquhogO3yJOYHval09Li7iS5XinK8aS5eC1U0+MU6j9Xr68zsEL08tcNIrLyLEPAV
JNZRuYWCAYQ9BYreVDcGul18YDpRn5k+POF1KZYu8y/lTcAu6YQfi4Bmzo/S7TT8QGCFxLDSXPvx
3WrMQ2rOAgBdcbabF8jyY9djnkQ1I8lczX5kvmpoqgpQPtFJb0Z1D4NB48cPl2NvPmCj49+HRFIE
HLyRKERqo91dq40tqCpbmkyyyM9mgmpeahz78tJt/RV31f9ENvu8xTDJsXHx0NMnHUP9rtTLptQp
RX2N/w3vnC+B7C1Fr4xCjF//iM3InXg0cMoZO08im/ccGExf3wB1IYr6LAUWYvDwCZ3DXIbyB0RC
lus+D3fSsoCOa2iTkJgNFPuAf0WK6sWePODnanIk+c6MvDAW9PgXTpko7mfcI831hVYRPozDlVP0
6rPbEMcGPk3/L7ixoWzGwb+D398+puW+VPa03DpK1UbDwscuAx4tncJFMeoSAwuFeyhDimcMKoIA
0do63dUtFGy0VFVSO9rmNRAl6ccCzDfxYfnkXLzI/nuM9HP9WOC7KWclguFl42daBPH77p+/iAMC
uyUcdWe6qyz3Cbgd0BoF1u0UBg2qz5IMcj6R4R5JWAucncwSnjyxPBDw6QmHk1sqytXXYlj3qCwB
10LjSXUO4PYv0kVJdz+Hhl+32Wf1AQm5LUClphG6k/sBee/9qE9iQIZFkyay2LdrdPZQxgIHBc3D
JXoHNRQBe5Yd1OsVGAEIRmfs8JBx2t0jjdFlPElAx5t5veQ08zLoCQTUBFfvR7mXP10oby38vRmp
CYJzR5SKXCgfKcvqYlZcLoDbF7JVw/FqiF5NTxFZMVELwJM7gPAjlDB4YEtsLQ/2teczdO4vOXuw
E4hQwMkXe3forNd4loSMB0cBQYXsNKwf3kxtGfSXJqjeIoxxpnXHI1engTqw6mbf66x1gweVSaYD
CI7hgOP0yjZSMg+eh6JjQVZirX0HEyShgBUdWqR0cVGQTu15MbKP+Oxad9m617T7c+9+Cxg6BDG0
ca6G6O8Fl5w2VLJSJgkeDEAnAINTOhbVxME4QA9pexR+A6FR/MH1PoPMKAnhXyCK1V6z1EM0OhVt
uewyi7lt6ZWZzm4rHpnalAUHIICGwtGZYA8EVyBM+XOKl0GGeD/ZDjM/J+ruovQHoy36da7p4lhP
ul12X/D6dZBpx4giTURIwLfmTdflNwi2xp+dy58uTZgbru5K7nd4UC4pNEF7xndA1AA47TDmMFZX
y9DzHCqlB/Ar6S2O4KXLqLi5FJN5tTzGA4LegUCRtCMSJ4VKgCaE/3+XB1igSaAfY4KSTrvvYs1U
gaAKTaVTvslfkcVZHn2Vrya2GmljuhU7InRgV6XMLG3PykzTJy2YVcpccCDjQvLnFnfhj5fKKCLY
WgJlHvGhuM3Nj4h8g+bFapmnRyDlGUA6qRynDrCxvECIBpeLEpec/6n9Epc9JqG1tI+CTYBjSll+
VDC2ogyAGrMaLFkPlVnB1CvkgcIQYYPbjS6N8pRRUIRYLdOLYVQC/MMXErBcp10GwXU4CTWD+Zh1
IbzUgB7z+m/sL2HYtrrIil1KH93AhUXbj0bEXOMfjFPDBOkNrv8cQoMzCLJOUzM1yNeLVFxLNxKo
GeXjryNCv+6aSQEjPsiYqxtgPqkJ+CPilhDhNJ4nbrNQin+lCl4F/Q5yCAsNMh1x9MVkOZllpNdo
slnIZckTAYoG8LEgvtyrBawFUJt6bD/xeO7x39KAruGqywAPZP9iIE2OauP0FBIvCHQkHMYgDVI4
gieIdRZLFqc+4/pR41rScny6mevXJ4GZgBspJX4pxtq3tdKd+4ymiDXhUejJyj2Dfdw54m3TquEF
vH2zysLSA4gFe30lO8X5xatIB4H8jE/enRir+dz+oldywyEc2rTj1F+K5jbI9mKNI3C5pywBlgE5
qrdwf9KAI499DIqaqRpvM7rANoKRGC0iVJYGmWSXY7IU+doZaR4lRmkC2AFqpQrIPIayM4dFRDJD
vf3SI1UnTbfrIt1npKK8Of89+MdklUYxoAt+UOeFVrQCf9dvAqeBZNBesczQTGmO+wivLjYZ9oRk
RTPcHBJQR1nRzPzsKo2lXgrWDRfJjybPofJiYU7LwIa4HyA9K7g2TM85IEP6T5tk5VJ8POCLEEgU
vfVfxXo1JL2uIV2tTKkrTIAN6z1UhsqEz7kcI7hoUsbulN3Jq+dmHVVS50RT8ZcxvhQeJRyWSGu5
0bDGKrku3LS0UfRq5Jdvzrt2NptjXB72W4WaGnIY3Jzw1YTfJxMtOtxZkyQwttdQL8NQQ2UxAUDH
RXvvu7DO4gAeJeUYH4V6aXrSP8Hi8lv80LGGfRRbSIY0TO5pwlkFynlyuo+Tf+WiLGRExWulGAvJ
nvCOS2SGPJHbr46YiEbSb+CFJ5GoB5m3FLxZgEh+BStbtN/S3vtPwfHxzs4jC0MzGfmcXvWbNUWU
rLypmWINAF5FZKZpp40d+eQzQ/oUhY2f30H5OXvPeATZFOYeqeCVptPN4XWfsND9m7Vr4zAsVn15
XbSP9tcLMe7OrH1RwTuUlNvFN8dxVA9VxjY8pJ0021K6h3g3zXEd3jmO2+cCWQaZR8bI6Ya+Boyb
7VInc6LXJspk34fUE2Dx6kTUhpFeRLaR4eXkrU5oR7hSffunSn43SJSEHtk1WBc9B9FgEYwQ7LwA
CeVwG/M8czBVdDYqn05HWMQ1qFWMS91oahlq7jSJOGvPzjwNowSES1xTOMJ8Jw6/ab7YmZoXD9Zr
7l5SVu6K7W2OaOMb23Vut939PQ3XxA1gBeGrCGhkBxVFm/u1SiUwPioHiXbLPekQcy61+hP9eyN2
1qC/ctv/RZpLZxdUzKm4OuJYBJuo1kbLpITO+2Sjm1lzVKuyDEiatfSnMjpJVxDF3U4kufFySTUM
8/vph0H3CPucg+ZTig3NeBpq/c6ANacBcGNlHI7f+7YogF/vLLURdJorlBek09f5xVNtDZRiqmk0
58t1ufN0xegTKo2TuoqByR/ksio/FC/dCEOfAg/pyv6B9UGm/CO7KGO+84EYNCIHuC6C08LIxpto
dhu8QTbeaSSVByHNfqNfOEd7DfoDLY0tKMgt5s/gsOK8gp+fCYhMj6ncZ0dsci4jITxSY3uwmWxA
SzWi8LylwVQJG0YJS2TZW7mjyFQ6tgw2xO1vTjQH8LeL+yhUjEBxrIgInMoG2wjwOCGSgpw53Yvm
TJo5wtM6cbD0s8KFRsQe6bCgiExF13FrhZo32rN/tJ3JVn0rJvq12ZBLV0LV+6PvoLnVQmndyQMg
64NsjV3QFd5gRwrROj2VLPCdptScLobeO/HASSBT8ybgW2JVwlKk/DSA6xQdERMVsZBipGsP+GF1
vIfgy+2cqfrYdyOb8U/fWVPsk1c1RCYkOhORjkHVYCmXKDrQHvh0wpdwlYV4KVn2hWV5iRTAibAh
/eCJlW1d3P+La5QoCA5A2EQ/SLlUA/5xXFp5cTWQIvxOGoQ2+Ra2sEzVBOoRRTgckdGprDE4R66O
c0Le2/qSjWCkd1LlB6iEGExXTgnHJLeoldRiflVrjtEc4cn9kZ+xdIFOrKUzzX2B5zFFmsuuqiOw
ovkU5B8Yw+2hK8ekkZQ05UENvN5av3DM/XFbySudgDAzwd3lrB+NN8Jk56LzrbdI1WZdwBu6vW9l
UD9HyU4fuV9E7M2fTcBjCHaRBym3SLKbf/4JIFgMHvx4QW875ioUkGbpvAmPjZmC69n7VPsxgVIb
etCg1sBk1jh7hYC0/5sX5dJQetYyMD+s51JhbYYlknnoBDg4eyN9OkxYHeekOoa5lZu0IfrKya3d
6uYLwCWpCXYvogN1eGCRqdKvQMki1j8e+eZeXN1/Z4CgoKyDygAWMCKWcRlbBpGPTup0DKPjhSrL
ykTuByLJD1ACgfkCqY0x5QgwDiIA7fJDT0zrpMZ0qUPQnuclDcqQz8kx/nIEROBhtcF18JlC3GTf
A+Mrlnk0QGfWNJ1JN9IiwzY3mvBg8ntgJ/r+cKWRzJ4A4Q7MsMpKQif5lOXibSz6EuvTt6OF1Cnk
dPnYBLuuNVrUwVeQgv/fjdTlUFd0g6YaREru2bI9YUpHWTn/YnuxPLBBvG9yGdb3j1u0tUyT08fG
s4h4nHb8gYp7gHgntKqYL9Rg1BWQ4Xhjpu+Idh+vPG0D6KjMNLZLanlBV+hD6NVc/LA2e9ECMfr0
6X7o8VgSJ7fWhJaRQA4TIYRWERioRTwk4tizqz7NnNs7Kuxoc3VmySuT1XuRUhC7mx2/SCFYA3cS
6MxQHm0cpzSZLuMT6/SfDRwxD+w11isyQdfj42GalZya39Vh46lizCUkJvtPiu+2ZF7SpcthglkC
XVfYY4RH/caydrOsVkqF4fV/2heoufMcjozjO1Axuhdld7zwwbDFb3qy4mN/sy4FRZyiA4M0bigZ
MkkAoh9TZ71xEHkVda8efN4Xx3Jykdgao08Hfbn+x7NnErWwdprdvYa7zeS8+S2ff5UX23rSvslZ
X2TeomQ027MgTLrNGNECnUN3zxr7FwEZ2kugm8Fs1od4fKt5dKZU/Z2Yv31H4cK0XNP5zZy9vUmr
SzxdR/9OUfM4BEW2/xtlDwU+Q8qDjim46IUm7yKQu0c8bdu8N/NPYpn5GoJLkqbuUGeP6aJ1bkxW
dWAC3ppEPRapG0qiqHMOiufD0SIhJNZ+/5hwuQeiVYjfRZMkqWt9uO2dKFKv+0xm0mvdtnu36hSA
iESiJNe4suyRcl/swFIw2NZUTLwaj5GDcBLJA0kH6jQQQWiNJ+MQUiGK8EL1VQu/MsKhT6s5/ARb
Eyf4t/+91r45zjIlEBN2nBdHrf9QPwYTsKWWxCSP2I2EL7HtJ6UAcNhgpfYw1fz24TEAXkxaYJyT
GBhYBhEEmPXbcPnjMPE9UBtowhKxOUIHrKefcWocNXHeTRHTSyOrxIWjIjLRkThG2H6lHTiqNf6E
h4Tdadu+LCs409GH+N6pLBCMAviCz8Q+C9x1mKmckfw7OKbSk1qA8BWzzSnDy4Pg3Yti1o0+0Soo
+MGwyAkgPkZFlg+z6dRB/SOuHeIh5tKbO63MMkK0678QnUOQycFZdqNoRo+dQX3oxroWq1VRO9EV
NmVZSsR3mphsvNAkIOATYiwtYQGdIb7QhJgt7b+0l/p/a+TdysHuXmMD+D9kDMn0dpX83vV/jsEh
7H7HyLfDcq8766jgl97/gJMh66Yzf0/1FHMA0cNQlO9oPk/GmanEoKO21H92RrKSXxTAXI4g3E9y
hXBVUuwaiyrNG3pI1BhmgGoMC2Jmqw4wlQSBGhvzwSbxuucxEdbC8nHf1YxQiYDA2KcPubQx9tzP
69qSLln3ShRY8YvpPxFwFKVrk4kxobz0X1h34M78qcZfYbZv/rUW9bANoBDwYRnY9ONovcAQDMA+
5jfa2GFrJ1wStNFQ+zdskaLnWMGz4bnI0tB1UAaGWLsuCKh4i+vOq4Ml29/KkK4lcsBf7BDnRq/Z
2OM9J6ycQRgO2/QKTn1S9U2bE15Q787FaZNsV4OPGGApN9g7HwX0y84sy378pYHtUWgnwxuv5HIB
Lf+gP2bLrxyH8v61bvqJnVxrbe0g5lT8I1/UG3eAXTKJz8sc2h5L+6jpc2oLpOpDu7s6pi4CocPU
O13aGHCwFbJ99NOwjUEClQYCCwG5RK5/DbPTb8O2WJ/wyWrOgMDPBAILYZCwItgw6fhfpAwh9bEb
38OVZfe4/HSLrFKFHXOvLgB8O5DwbnHWRNyD7ydG8F658kcuzKRqUgLUti3ZBMod7OSvEs52RgWm
qqwhfK5kKLurEYoR8BFF8f2mZ5Fb2RNQLj31tcHDdq1daASHcUUtxNwBr+0qGHBvIOeezeDa5Im8
xDEX0OGXpZhmRp13L0ZxFtveHF/emDKVAlqfXES7xTt1tqTmTEmEdGnPxwlDj29MSP/W4aLIA1ks
XeDQIPrufrtHmpS8r6UwonAPHz8LNcpSmp8U/ZOVQmXmx2zkX9qDJHdgUyCNNFns970e/hhFuBWP
jgkMQnBqykPILwm3W3vGTVzxQmWO1pZyMek/DmWj7YyKVVvPrgFeLXghZ8TX+gkY7+A5KPmbjoqB
aYB3SgitVtVXIMi4Jz1pjM71b306iB5VOwpBidKYgdOIgrNN3BtUr6dEOOmUVsA2TdqhjxHZ+Fmf
ahaP9iGmL6Xi74wed+tN/Wbcv8p+th+anTcyODz87ybQ/hv3FIy6L64UDpHy4yI5h/Bhk8d8rZNV
SGG3cY5+ySyUUDZdl2/Ba+2JpyZfO0ZggV3KpTuvxGgc5NpbtYwBV1XSJcZrpWLcCDYpI1X3rOkh
fYXk6yykwTmnT5r4HqG3LCVR2bzTGdx78Ah+ee5PaeRu9dkgVlKrGmlGdZhnTSy3Ys3IdfuFIwC2
Yegh3G74Ne1xLUfbx8ozoQlgCq0b1G/CnBmfOBP3DF2cfrrsdVt2NqaoUXprloOqyZwpwEdaXnSg
a29d9ebsTwbBFNcMuNZo/2YFJ8qUDGCusvYpZDqGHXrVImyc9zqCAhSq5CNtmMl5jNJLECJ1/XNZ
bvtQZEQ3PMl0JejEqIVPh511BTPHvdmzezKqlGd22VOP3TLXNjVOfPL5n6VZ/cGjcPtMaZWCJJTS
9t6ebq4EbZEKa70wE/Npf3QjPS+VirXaSpsQ49nF8rXzPOjOH8ztlBUyFuFf2bz9io5gzali6sJU
dsAvV3ccLKe/1Kc3X3SNqEqZIVKyWs0J68K8ybeEvGGZMfxzMWhBz6Iv00dNDNNB+nZkmnDDWCBE
G9n7wfKqbWvU++Z1lRwfFB7SOh0LvqJGyAjnTGeOS6o5MGI5mVZLdCjREr/Thq1qdJo/yZTU6Pwy
Ru64BClQI9XMbyoIkGyu9FoqTg4QjnV/L6FJ26VItYqmDqlXL/QAXW8Y31N0mGSoH+mRb81GeVWP
xFkLxOamyHE5TqxX9WhYWqYvEbUk4fZaGXTrJGWvcWb0JbGrPxicl4KmOVc2M0es/7/oYLiU3a+8
v7qayyAfvISc776174NdiZZngoBM2AlUczgT2CW4BPqb1+WO1dwQoMaDvTtp+4K3HiRqmwp+SXAn
kZe5XltQoeJ4SSGZByMnGza3V/9yDEnRVLslpD6aK8ARee+JEalJZDTiiR3/A5iL+lOz614ZnkGK
hX2b9d6sqZDee1MzvbPILMsjo4YqiAD6zMmkwV7FH0eln5hm2GyI2rGcCdQG8c96IS/0q9hL668W
cjF8Tn9ab2WMHILqj+iK7tCMAy+AKIj4v25uvn+B/4xG84yAMSa7xhzNUjCuTKtWiNXvNEni0tDq
9N2OuloZRghOpXgBnNborDGbS/uYBTt66BeSt9RQWmJ7PuNbbWsB/RQphbPa+rgFsB/Kac643klM
aHtxrwDN06aud1dka9PJbLnLyhHJNSS5sA7ak4x9tS9kns0oK+EO7II4BJZEwdi+uHjHqOyy8c+a
WgyJWEOK5U20KkkKPS1mi8alw+4KapGSsgyGucxmltLyVlg9zeOtxzuVITvo0svrKMSHgIZGL8nS
HRHvBidS3jXOkM6UoLx/JLRuzLkxyZ85QCgBfP+O6CSe3eEvHq7ZiueGxaxYBNdsgGqYKCcRYcgF
bQopk4Jp88pnqCSwuROmcI/kNHd2vBxLBnOa5dXGwmr5VVy1HeFHY4ijpW5x7vRfV1jA5Ffunuoj
eb+7kPyZXITf2ImmwFCrJa8mS3Gp/paR5Uy9Ti2caaesiRcKPIfKsz18Bn6KvLmXBEL9iH4+C8du
eAkx6Rp7cf5Rwcpl8w6wdHsUO/uCRrjMBInOQgJlGiwAtz+etB+YnS3W5Q9wRMV1ASL3EoWzUobq
wOfrCVxHCtqxGULROnV4NWbweDr3yLcIn4DSVAJh3ZrccibdVVZdm+zRWnWn5OqaA3c/Hk+Nsj09
wgp2UgqOCZZQRF6sCRIvMIM7Rp1vWE3f+0qBwY4xHJxfvgLXyf/1GiNO9+o84QO2esKyKQguqfhc
d4bXsj/Aq5XDTbF4rXP924D5xfAlPMfqOloDNPH6E7v1t8h9MtL3TYOqDs0vl6/nxiFxoFOhbiOS
l9em/1rtp+C8v9f1FEd0e42sJLkPvy8aSV0RXNKFF0vyDOxnjE+XbMbqwHOznalFjkQatL+5DtUA
rP7Rqqs3DZN3JQ1AyHzJNPtqGYphuuilMp5GaOC+pPoaDkkIsyi2N3Br9NOYO5JxHYx8tuUBCZ7E
QU3RVci9J0snGXxaBINhCSZl4OmO9rQTjfjBTjAPRZf8JmC/dyrLnkYD/Tj+cm8QL4aqpI13EIOi
uHHPQws4ezxIHmQOKnThTsmzWfIECp3dXk1+nexvPKT5Oez9m8/dad42YaRu41nfEIJZSbgslRvd
zCe+Rh9fbjYOwmsLkpABVYES5ZRRMzSDMkyPFwn2PF9OeGC4RHFNoRjJVQ1WFGHMvNJIplyf0PGu
VO2OvA0P4LeKzoPTO33JtpWbz8543kH5JbM1ojH1XUDeNFHTpcrJHFQg0janLBDeBbr8A4/EbZKa
fqxzQKoAR398gr75t2GozG/rbMA/Iwv9wiOPQ4ZJp0e9Wd6j7AVcFKzEY2hrdzMVExZBAMIuuDhT
ZGydTcjLy2xEPmR2PAMnFx4lFuTVvCuUVenCeDMjPYtQ3uLDJn85WBh3tA/n/b2eUcrbk4mFA3oA
1QtqkCOE7ogxBMKYWsWXmtMW/hmsHhZC7mrQfkYnlPxDcZuG2Dcqs+XXOwRUKMq+UxalvJpuLi4M
jkfKLBt0XlfZcjIIrLkAbtaErbg8jwkWktpLZ3HQ/QWqp9QVUNzNdZkT7VBSOBy+yjgTRoAeilH3
x9YPDdbYbwpHnsVjAsUuz5xQscxXAW+ahGBmDp9LHNpJP2/tE38KVPFOxZlqfgZk+6XIc4iBh6cX
aNYe6us6kYjS1aa4X2R2fKNxUURUqW4ucDOMZSH5y/luoLlvOMnLB3CqYd75pguOMxHUTt0qSp4g
SCkU//NdjPwb6KYsOhL5+CMqH3bmPU5ln0J2DUi1txO2rSxHFD9wXGbugfEQd1NG/zOSl1/Wterf
cL8JJ/hBPocRBQVLn7LBaLfXs0sNaeCfW8wEOwj8jm+kOkk37EvAdXH8//45RT4yvgapzWLow0La
mowusvA3urf/L6BU90fzrHoQs++0jnnvLCfg//cJee/rUKdPlj1+8ObhyR0TIVyuJ8S0/isSlgPw
tuh+mAwUlohoGl5cP+qR/XO6ragCjzZSbffTCyHJj3Ne2acYw+nXuaIrqCFgPzt8nAunOryULbSa
lYbFj6n+3o0R2hbBt/Kee0ZW9iyfbhQx6K3BHrjX4GUaFMnmvVbQnrns4hV5rPcjOhJurLHL4FcV
RPalGB3VK3FtiPNFcxT7rL6MzwO6Fdw9xhq3d3VHUaSUSbFtct4Dc3TEs+3LLtmxrZdSQi5dJLJ4
y6vzNmsBzriTwr5uhPrS3xWEBBON4uG5y212/7ihmR6+XHL6du9OR+SKOwXy4tD+0ihFtQ5rQ0bg
5OSyA9Egb7V0Q8cpsAbJUhluKpNEKvpu0FWU+iCvgQwVrcUtp82q3U5rZ+9dnzpG1Gr1n6MLu/Rv
OgHtUAQ5oJhrEhW+5uR/TbQqRoJYAE3j1R+CJZ7sRh3lfw/UiE0V3b6Z7l11anv4mj7Mvqq+3v2l
/1tMBNnRvThfyI7FGZI5F442714+gj2uKaxSZJCI4m2H0GNotUwXdp0AKjSGqG6MLqoI1MwQQ841
UEcLKNLco+G3GjwVYuYOn9I89FU1MjfWxP0J1zcqd5BZQQDuCP+eXPyB1PQkJA4SWRccrXPewQSR
n4NzM/UQyKjCAGESFvSxW6wgqusW3NKo3hV/cY18qnxd39nuzp4R12Z2baiwgchNJWZofd84xMJ3
1AK4HPoL6yy3yrO/K5ZeV1gzhiTsXK6vtZXWPGS52yK+rFR/G9cRut8fQ9vt8Pe0pHGuv/Tuq+B5
N6U/6MPjJvb4abdc2ZTGEuN+BqEVgCvQQbUZYGkRRxqbJe9UGlalEyzrReKsK1R5i0rbKSUobGw9
/889U2osdf/1RLTqTD4gDsNm6pGOQ8/pKoiua3LA1PF5wj9ERHYEWfdcy9V/AlUPr8hRKSf0y75U
GohesIN4yr9nq5OcRQz9nKmJXdc0in0Ary+Wn/J9O/fc/WqylmFrTZvehNHDCO5TinBsq4pMygAu
k7kSGBbK6ONPlya7H2tN2lUGPR4T9IHMigda1EctOtwQ1HjGizURqxgmqRYjiOjtkfRVapXBS303
7i2pVcaehp5/FCueuYilNFyWVbw/k05x+aPCMc5IALiPwna6yVHI2iyN/j7tecYzfzrCh8UVpb6c
JPVW4c+B/AQP+n+S+4WTiamBz3VgoQfyq6KNJeExGIPvH0Mc6yLhksojZuu9CJ5VFkaXdzFby226
xPZWW9eEb6sDzSd3iZn78MJo1gDFqAmI1Y59kqVOXW/qvF0Ll207zXmiGf4tWprn8pRmhqkvDxSx
Cw+sfdTCqe5L1XyL5bhpfWUt6pptyTm3zpOfZapRZNanBYB/wiXB62C+KqPz06DoBqvyDoPJCsut
Z66krHWmeb36T/LW/+GMVlCFLvcNAsQd2wQ8uOBDeXOc1IGH5lIqHd7gDwNKfDSaEJKqYHT1E5/x
JJmfd1uwReKaRcWSbflQyvWn3P+sejOVCaJ51AAjyE3NhbwdKxxR26uWTdwGLcLLC9frjMoDkLIx
PzcXpAR+0r0DxiwS47xtJ1RegEAW8w1yqHEMpIodijI1qPxVBhwzGcNrlbTQb/Zj2oDZ1n7ng5Cg
GjB1rUIwQ3aAHQezPSC6WjPDGWf3E0Ez9X2UCK5h/YWgWvA3QwuWyGCx2X46XKeO2BVNj7sCgmXw
K9UAF/vseYw5Poo/LDCg4f8ujEg3HljqSXBJ/FQA0ZFhGD/dlSPPY6fC0SsvaP8L/Vo6aRdTpk0/
s+G8zquOPztCbvT4a9xWpk0kwMG7KhwaKYJuSviW/n0L0TywUMZdf2M2/zl/E7OZp2UIvI9NopMD
C/eWhg3Hj6GhyddBj1Z8c7cdf/8pUm321x+Sl1NSORNMvidRDkjsw0InCSShg7sxbnFawQpvjj01
mpNmCA+U+LAHiUPF8gb8+daLIjz/pCLWmbv9Rb5mUc+tFNPnZx5IY2WViqH52/kfdWwtHKBeajFo
srIeUyBKXPbr7KZxf3Vf2lzgHfZljFODZVl7bcY9x32D2jpnv3i3FuPxUfW0bO2P2FUhRPLz1jCl
9cRd8gTfV0hOsynngLBMzkLhhMaFn1zw48clwRN04fWVQg6R78gYX3aUAvd4fG2nTQwf5hhtbMHK
2FR3r8msx8JphhnijQGJ5xJQqhHsaY930Z0cOfMPUEobIE1jDaA6ShhljtCa43mCqaUvZ2s4vKow
t0It0WhXitBCSQNkYRcTrR6cIvLceLV8gicfwScejDXJ+kgUOx+aJTdQ3ovHDikwxRIgKGh5A6+j
S15R39Xb3lYGNOaToyNc8SOsnhG7KF01tr1RVIdUqarJNt4ryxdyxMOrxETt/xyTHt5MDnddX9Ik
T/pit7eONwg4eCYMTwrQYhq3CH7UhohoL96P+jeQYaBtZ5y7xdlwJy8EuKv5z8kqtluCqjJXaHc/
CMXhPQVXlNV9TgLkuObJWDWz6O5KK6Vu0O09tzgUWN6jS3p+YqwOLdu6J8Vn31Y0/0yWghxAGSQF
0lF/TKedX9oDYOFaHbhsSXeKjiOqNO49loLUe0w+L2wp+6QIek+qffTBOxlbEXtpKaa7R9Ssqo0U
dHXBHdl0AS6ghlB0Qb/aLkny4qz08NfjAumD8A2WUGq//f3E8adU9ehilrK6n+lpVhvFvW8YUeIx
JZKy2oVnnB00WsB0WrvuCuCfPdkhpNzcOXJ7ckg6zcedENkUNJqtFI8004TkpKhlW7Epg/lEmUko
6IkFAXqWaxhMkeGTpGDFlfR5V7xDcSwA/U5btNSYmnB/S5hP/PjQ7NUpxdRlQ8e8pn5uMzIhlaCm
nEzyQrqzbOrsX/40F4NJ0J57OmE3vVvTEUSGHfMtzrvjmE8VtP9hR707csK5w1elUdxpM4NcKFXK
1i1PxuoTwUabOf78Ix4I9YnYTlcgFMF/WhPFwdcDyiSaz45KK2pUkzrcYFP9KD7ADBzROuCKa/pE
YrYD6Sa1WiuN+nC7GhJSZD2+cqLljIcANCtUnBo1OruZXj3LEfM4nY6JgRD3dG9jWqUcNMGZde0w
wFd2kOmDm/8S6R/O4rBnGZ9QFXOz7Itb+s72axeudbSUsJZQPLRupDHeCgoGwfdXwROQ2vPK8T9I
PEIE53bFal1Z8164jAPzeSQ06K3Lhrf7tl0HSV3dcEfUZogZmjY4AozUZNVvSq+zLTHOVaNyrfdY
dHy98AG7lPF3cHxszbpLURvVdAnqH949silh8EIH11k8rSVWY107XhQ05e7CLpI9Vt5sEB9Jux3Y
6QXxEBOzQRDB4V9ETeIL7J/c2E0PwTI3cHsgrmFdFq1v/+NPMG556CFfCIn7aVutiJXjquN46H6Q
Xuq7hEKT90UU0HpQs5aknUaxIQBlrl8A5meETMWs3ljwjbhE1DD6zP38CK4+s4oamshHcm+vjuOj
LqjomN1XKVc5G0HD80Tz3u63uxOtqTfYeyAEv/iExsifYaGfcKy+XWivPfe4hQAYqndqd6Sa7bDH
2R5QGmJSZQIIBX1GqOBejkbpbFLM03yu58WHFDNzZcKXnv7kPrGtCZSOygilgcj1XmSji91TlRcM
FCtx7bP8tLf8z0iGarMpBas5QeHN3ctf6ZPL1cx3SIx9Of12DxR9V1uWZEy7DwE9qIV66W+Gv2ZR
QG2zW9w5BGwVzgyFEuvqtCoKA0jg18Xxj0TBCTB0K0h6SpWDInXhdyPK3Mg+ikd7rni6z004iOjT
JSEuc4YFi15e4ZmdUGbsbcuic32R3wQCpnm4EqFVugc4/q3IBBcfc0LxL5uNBOi7yEAb2j3UHEsg
jvd6Nyw1225jlFX3syvtzwrEdZWGbGkSYzgfLVLQjNAYauVQ1HM9orRSqTrwhHMMMl58RuebgZuM
PNCxyt38dWKqiczWFNiFiO6Udh4cuW/SALdqvmkEBMVKsH3VotIjrGoIjCkoqpafq7hXl64n2/GK
5JsSRlvdCHhWRi+Hp0Q3xIlDpT0eUtCZfudwU8++FI37xBusw4CWHyKRfeNfO+a+DdtFdDTAYik7
30dFFAo6hMd5TODX7sj4kJFQ6MMAy8zuLJHuZpPuXV8p/J7JhfEytHJLIYz0Yxcfnk1cj22j+exE
KhekLdFI1HzQl59XbO9Z+FOUY5UyU03Y39URTkGkvRPIwiWjPPJlrPEdsuBR4EPNq0m2W73mblC9
efv2Z8nA0X6KAaeYk+7c4wh/fLhM4YQwEX5CDHO5Gw4/B4tSAeB1CtlADo4/fj8kw072C1pYneGO
RUccXz4JO1izUx/+HWQu8OqGfFWy8BoHvoyH5C9yI+J/L5hUArkkNfyJHHbSxxY9c7qzvGErffps
51LZ5pX3/m1Uh8c9QJQ8E55v+6IgqQBsK7xigF2EmXeuu7MXaV89IFdYrlHckweJ+fF5aZHAM7mF
yu2jhtIzv0besUdRxCndoRqXwNrlOlT6U2Dbww1HlPiRIxITGM9NFi3+RU5vgNamE0csA996j08c
oBD+2jrnPniEA2SFk5Zqz4lN8Gxf/ojoEUC5cxw3Fg6ZFSWcRaHuNn2Nsksl8SXtAQZwazuff36J
XBdsTbVLFlm3EsW8obmY0pCqe3O6QAYWflNr/1NuoZqQIVNEXJdbiaT3H+PbYEQmCRkoTO7TqtrL
/dDzEXS0MbdjFG83vD2z7Gx6gNxK2zX7Vzs36hYgYsZF2jroIdrO2qBt71sB/8vNznWwoGMnPqi3
9TIVMG5KCNRtxVdPSRPudGEim0nND14Xfi/u+X2DOYbNywLbQJgrvAgAYlsN2Hl/DMPl7uWRCSMq
REwByidDcTrHzTQL4B7lm3wMFaShPCEq68EYa+0i9kDTLwYmQP0kZxYnAes6aT1uVCJeEew6Vq5P
rtbvUa1Fo9okXhMPb9NETu9D5DMyfgQereQ2FJbZ1p5gguVNMNZivebG7tCfXU2TV8XS79u5M1Bi
JHNMokeKmtPQR2XSBePttFAZNBwE0FuK8A3oGXVwj4hEsoIYrgLRk79Jhn35nDrdiKgoBMWV9qCn
m6ZHZKpCx57F9F9FVSOE3ZQwWgNVM9d4lRhPNOa2kb33ZJdP4DiBu4+7nmoFWFFnLT7Q8bPzqXTm
OpqK+5SWTaNu6AbWE6rqMIJYzk3y3D17KqU3IPyppXRY5dBHGEnj7YN53nZh6L6mh8YZeseSaRad
YNHTMEWOXC+qe31lM/BT1/riw/3cLIPu92NVoUZ//WiuBpS9pRVUj0CBQn+hNH5EAE3wILxA3WVx
GedcPxg8wQwp1elkuonBHF7zANbCtjpyJHvweqiPzG+Xc1aEGivEvYAvBnTSo4+koejnKWHmkzh4
e7cwwDtnL4P8RWyippYVyyKE2sk5/p1qPQru/wyRmVCZgRRk6l6oaEXxKXw5zJHJqSCfNDzuoRpk
4MTpB0ARSYzOdAho8Aj1BfkgNJ0LOUlUgCsGNEkKlzyokMZNDDDxtW1Gu3xjJP4U6JDVyKQpBSPQ
uBdMFQ65xZZ6By8nNBN5+2B2TCGOGumE1tuhmJrNIGQeCw5unqpB8XZBzoGR//qS1Je0FO20RjsJ
hRh8zrLVrhn6YCvqBlRJ6mHuTcNLQZd37ZU0F7gUC6cfCdJHJEnuoFhvWbabQb+E1Qs9JPKOF5Op
lkcDMJWe+AEIfgHxZ3XEpJIOo3lv3GcIvjKm0T14cLN370qF/coVjOsahrK6tcRmjFaWQdDrCkr5
PnqOjFxaLoL3iQV39VlsJfLRs+C3FWNnYqi7iugj03r0c7Om9w86YiFYXflNxc7wtsEaEBOJrXap
/36DELjLdQnXCeiKRRVKGHoEsmQMIeiHF1C8SBQWUm93IwJDOoU44E0/xVA7E+VRxV8xafWH2shV
rJWCm1g6FR16CFRnW5wVjII6Djzv9ig3ReD3z6pGH506jsskCztgY3oFWZ+HJWOYga2oHHbq/47N
3yeewlyQUTtKkObGuPPDpbrGXEsolZk6t1OsnKfVohgsrt1m5AgoIzl2+XyCxGs2ZRWdp/1+LJ4M
T+HP8ROkGJUktDT+uE5cyUAah5dUCgcOjHZIZHyv7YB81zmr6s/H+BO+WvmtOUFoDdwXFA7TF//5
qlzgvai0mWQkYWiq1ighkO8qgbgh7dfnKcD9bDQ49gAM1TyPMtTrXrNZz2drjyzeo/jZ7V6Ct2QJ
CtzPWz3GYoyzc9A2UvzaGcPZu1QVd5HJ38dNXt5UzKJ+pwdreYy981TolHkbhmeEiOLK+YcrTIfr
eL6Pd41mNGwl6q0ZYPBKVzrNH5plqDPXHpBZB9illUCGGnZVcA4tetUdC0GQGAoNlltg7y7OC81t
BY/m8/iqua3zsUe1jDfqyeDml1hbxAb8Ka77pxTr+OOXF0Xv4ZPIuIJvqMfYFUX/8cfa1cckKgPQ
U0BUhe6AE0KBwqpB4NAXgJw9/8xrUWh++OeCVNFRJ1XNIhcomLUmnZ5Ie03GQD4ivSQL1f8eLb4Y
b/OvZ4UaNORTKq7anGwmUVIJOPqlw89EX4otUNfzxNA7I/qho6uRi/ERl8whna0PnCoPHnvU3tl5
CwD4K+kXX+zlAyJTt7PY7BZeoM9k9YBtcqszb64lnx2DtrTODaSg6uBnLWK5Fu14b0G/jKo/B3dr
q0+OfCw30zYGNqlJTuD5pGfqT4c7DachHK0+SY86Nm7nqGJxRpWC2N0UnJzI/pNEO014WW6GLfgx
noj3BfNZCvjNWZXzPRG2NoQNytCqoDFHNaSwgHy8KG5Z6SPbu2nkz0XuKWFk0kZE9XGaWUv4O4cb
vFOIqMMgdagDDPkVT0GmvgbVSVVCVPbwU40jAMMF5QZ0XbFkSk1AZVYw8JpM6ysZmjQ0mYI2UeZ/
uopEoOrA8OdaekYKTca51Zc15G3h1LjQcub54nD/gy80YB0VUYVmAOBEyc7gPYlweBifA+/X0wFN
4y2usMbmKqnu9UEsCelC875kehUdyWsCXhY+5IOccR2WUpMdinQkf2QdIO2UI62/eVqp97PacM19
tDuZhMuenbEYiTwa/k80+bsq0u1Q+YX5hdiaJTWrjw9m8jTf3p5LY+nuMSolGDFYMyvFtFxoWrBt
qiOgw2MZ9ziUMiJz9s3CmVk0d+tnx20cpiSTDCDNNquFZaXrhTAVv0ovgwD7AC4t8W7yYAT4iLpZ
zRqcKbnSVaKW2ZPK7VgPeSoPaxeYnoIrXCd2UKd/SUGD5Zm2atRtTuj4e9oBYVGzLjJc0wWLwnkJ
LkoYAZp7L4X6idDW5pvGL62OsCpTMhNUecCtj+25gqxjeHXvzKi4t8iDJiWOYPdG3dX6FQhGboC3
dicgD0V7sX4Xs4HeNOPbEjV5eO8x/QKAL3vbNS4XMMPSDAwgxrJT7vI5/Gh/JqluGNwYVdmAVPzM
YFIRi7wbiFGzIUmwAWbAApSVJymJ7IgEz3VyljnHX5PJI9WDPoeK2cH6LXv5lPD2Ziv5JC9a9m/2
nPjHnVD+U0BRPRW7l+MtZULpNe92u0j10iDw19YQEBfA7hAGz0MxiwjULg4rZ1jKg+dQFDjHC6cE
TUM6D2jjk8ArBCMdh4j7ZaG9tfOfJsSIY7W1TuCEnnZNq58tixbR+VOvf/I9g+T6K9E+qyM/3y8s
SgGbL6fvykxYIB9JLdDIA6cBDZdAfXYZwVm+kd9WMd1gJIeZUhemZgRnLnnkXSYeOld5O4ct5phX
6Jop99MK3wibGOCVldv2WdcJpSCqKOC7uNFuoBx8QamjNDJng0ld5a6upeH4faUzjRd36mN53cwW
iNCcpVyEN+66U9IExoEYgLNQxVPggSV4pdXEbm1FJpFjmNvZ3ewNnBHfStquc0MInIOc96NB9W4X
4c9t4019SvaW/ostAdM+07rii+qwFKr1mlyq63pAgVJ/q8WiaJ6g7bBh8u98xxoVIkYSdkNxG8Bg
oXxiAhW2KrKTMY2UFwQpIklDb9hNATG88zAapw+2wqkUG5zZuXvjE9ISyLdJLBcTvzQyn7tsAaIK
6bmW/13uArQ+22ygVlEs+J+RgV40gjd8hdM7PGah+Icf4+jJWlS4EfFotBkYG5LVtuI6v1KIEUEc
VoYxLWsHF9wBIE6zWbhoyNK3QjXxNaNH7jON6L2+2tzXRo0WlF08siSNpUJlmhB20aQHee5kuby+
iVXNv0Fdeb6nTfqeBDigzWWATIF6lgE5AXesmbWykj3Y+h/6wOe81sUDaHyjhCGGLiWxN4UWTol8
LNhCA+frpUI5at/YX7XSsK3u/rfZF8hBiiIDE2sH21TZj5Hi8coTHXvVf2gdBy/bAigtV+e9HkKh
Iua1cFQKv8jQyZ1pdKeAOjlMELHbFUoXu1g5+JdWsvrb1LccpTJ5iU/8n2ZwUCtmyebb6G5nO2/d
0HTU++EJF6rKfyxPqnIq65YLHQDZ3GmjAEMT6/tKpvo87o0eVe1cXDJC+/IUXcBqCs7c5rRhysKI
VNnqA7tbX2/1GAaH2VeiJP5/4xcPe/iEa+yYEe/e7D4pPLFniWb0inBT2TN/NNvB+T1iOW479aUq
0elI07WJP75qhSGomWZy1tQDQ71N8q5VEcIZh2GneQjpfWP/bK8Xfup9qXY02EVTEmyccOFHbOOI
ZpBqi7cN6s1kpNi2gtgslPag5wnx1TCqYioMxj4DD8Xlg018dZRuVs1d9OyunAL8Mr5mHUhW/Coi
30KurLjqBhljDQi16YkGb/61qGP1QBVlVMOe+z5dvPW+aSjn4p8j3DSQo+kq2NatKqaN3RTcVI3v
J3e8G3FWROBs1RtWk4sDzRvAnqyNWQwAF/FC7QHIlD0xdaG94g0+Wvzi57j5ePY3F3CxcQ3lizq7
AHLf3gXR3A4qhr2LHlpvUjZc409XX03w2Lx3eFS5MFYh7EYSNbnpzj6bJSOs1PvrxaOnYRkEuxDx
FHLIubLXD+gnJ20MXER174tny61ZQBUuVx+9/4RqSxLY9VBhGacyQxwDLN5ZfqhK2rjJtSkoeGoB
HRwkkI/riDNhwAUcWrLM4mhp2zsHXu64lrqO1ZTJ/FOQvtfe4YfchY9Bs0Hy70uGWO/HNpn2nNd8
HHS2hgMVzoCacbAnmsrC4NVXrScKzSxzMIbh6ilR3rcrxg6QoFO3zJnFb60sFm8zU6vxy66NACvF
9SJjiarh/ewsPYpHuzaJsBAz0HpwKQoj81DeHyHbgQZkP/aS/2xmRqcGEeWtIUKlEQG0xLcOiW2f
vEuMwMWrT0k4aWY4KZ2vmjFhhP3VhP6wU+k3b2TemBm1lC+muJBfFqnm8Z3/hlgYuMiY9myJCOc/
y0EpLWkRVvUeo/rKKd3h2rg9RIj9ObV/q6RgFcgmpLvOTB+JHWT0KFDg0tSyZXmF+j1jFq4SHBXd
z0b2C105VLQb1/FOQlihjl3CHEmKpG+QsSiXgmCu1tjoMLXW2RPfF595njqopWBhC9ItLPDbpYr1
uCjHnKfz5HYjnOCFRNT8d2sxhKXsLaEfkTunMauEh0LGWlRdWHBEMsOkSAXHh0w8c/LmTNV0zT/l
TD3H7CJ5UsZcG2D0dKqhTFHjzwVybnNNWJdRs53R4BEAJvfsMDkRZUeCvf23SZKOUGj4ekNQHYoF
n1ytWUV0SqqmqNZ4WBfRsMFF/+JzeBv8vm6pmcP4/blYL+CHUsmnIQC0QouG9mu2h7hgcnnTqXnL
RTnXpOI/sdIJa5VVDtZ4dHM9wcOQ9SIaiNct7yTKD+kkna5oFKJrbf7vReqdcu5yN1Yp1suUwN6g
3dNt6Jxr0523KfwXoVRSGyNbfpHRRWGBwX9tYxYrKajxwtXTtb58RmXHiGybpYogMZjh0YKJDMai
pK6zF8+19xhocw56hS5HE2THZruIFjQtVKK3RREf1IldMrf31POz0/QsVFJX6qHfddFNa1JomKby
zKR1R13TSdvheKsshHrsIv9O8m+wHT6t+5kY1edkuLsBch4exnZ2kVvLn+euOa9qQ0TVcVWk0Xqe
9h+A6U1dGg/Wj4T1DQFL5LVmJvuQ04/MMskY97iyi8UZ/UwFhU8o/EiSDW2hmgNd9TyiW1NoIBFi
kz9o2CwDqxiM011VblAE/y+KF16fVjVzCvxPce34eAY+MZZTl533KuT6r2JeBptv9F062200ZneO
sqryuYbBavX98M1Q70PXhE9H45dpc4XbVtoRN1lIU/8ETmBjKR0zR/z2g6SjCzHtOtwh7P6DjJD6
cIZw4kFOOrnaGTlesgL3vBdSBo+FEtA1u0NU2eC0o//6t5jzPa64fmZCJ9QwSEsUgdz8ZG+8xxAr
2A4mBlDWjX8KlV69RWDio9PkKuxkNazQwRG3w1kJKHWodKe2ygOyjb03yLSvt68bWGoUh06eWMQP
/T1CKFzb9j9KSw7WAWX/s2UK+HvYrzI1/Pyxc/UvHChaI+Kr6pgbXridtzqeyT3KJpq4n7TfJcNH
btI8pWvgkNcH6YNssWj/SD6uFyGH5kZI7Xmnrcpn/VmT7dmX0ycOJzkMtfw0oixK5Uq1QEVy/8bK
k7b40rIqlR4s/lswFg6Pb6o7mGTYDetfUeKFZeYwaBXRxHwyYwffvb/IcD4v/qCz2pBVWdYGzakp
nfzul/HvTY0znYHETwx0EjcpjGsHXprzLg09b2idXQUmP2epBUiyfFnpE9vy6NPqv1wMbub8z3I+
vm+cAZJY5WEXwN22e+cx/oiNJNsTHGXTs95DrYwqPnSJmO9kzyyN/LXFj5QYhCqv8yGYYi51zfDP
WzjU/DhRvW45EnFlA53euSUfzTKwoC4YAwvwhhEYPyssUWUyr+si/9w1BwijNDFAMv/1si2FSEdc
Hgi+vEU2L55mE249xGo7teRw3k3xlSY+De/jVmIqJ4U2TaK4Chsmg9jCeJtwjWlEXLK0z9Op1fyu
8omsmYgmxqtbZ3Fs9Zv+FSR4tkIELOgBXAvr16vY06tkCRSt6KdhDWl+7wQmedACy6t9GYx8hng8
X6mVyrvP1+LR352ZppDsXIXUL8k/PWus28KtQBa1F5+Soo6vz3PwBqh/PFzYaCZ41pnyT8XM0N6i
N3TPk4zYlbOOFnC81CYt8vRYQ9aj8Cbz+Oo+ZC3h+MH81CkTSYYcsVzTmHzJekEl5mdGzT5WEKwK
Zj6ob2BOhp4t1fVGgF3VR3eviB3vbmcJiX9pUpAtC2RHoRr39rvHj94ktB8S1o05t8FcWoF1y4Xz
KhyISr1ZzahgbB6Cboji2pKps8fnm7wYYRCva9yFny1X5K4ynHhM3qorPfqW3YlUvaKT79fH6FR9
1NjZbJijqa/77dAjWraWA3cDnMwo6gwA9wvL4sU5DAAZqSftqTnqrkQMSa+drPRJ5hChUh3dzxgu
URaUkwrR+tmMJ6aj6ArtBcXpmp12iwggIpnREt6JtRgzAIEi+eq5N5b3b0xJtAjEC6FCE2nksyx+
Nu8Ho5eeg2CcuROGnkDy2/NR6p6cKCPnYOmrremDqMu+EsILYyu/cyKDFeyRRzuZMrYoXOWvAW79
8ZgbpVmcP+NvUl4lyOLQhfe2N7sXY5ZAQPhpO0kcbzLJvIBmbD0H9KlTJcPKDzcPuVVh6QT//nyq
MC4JM1wmnb5Ifh3ehQp/MNLMYKOGA8OC4YS5XIPQC4grlBjgU8ydB0uWDinkbeID5bM68wS4sfC9
Y+HHdZbl7/5Z3uJcSKcDnD4zuBwVjxe7oc6Y+r07Pou+3z76BpMR7zOmc06CnzGR2Y+L+fcBX62j
keCPPUf+dOzWJ4sAiHYVNs/wK/fTmmaFl/VZtbVfb05VMNPDSrdbGqpEy6d7GRh2eeuBCYb784+J
0jJaE1tkruSdqU8DzHPt1jpCRPbILtX4Hfs+nplG+AY65GlXmYZJUhHZV0trxjzuoBLIMwEnjUV1
SUi5MyZePbvYlMZUNZ3ugjpvpQwedih0BMbWgPeqaaQCCJGX1J3e64HNMpDTsUC/dt0bylU8pgbr
75GAVDWX4SGDpUjc8HgueMrYQQGM7JI1yF9emdpZntlijiFZfd1sx+1KGC77z03+8mCll5rZRs7W
n6A82xih3GmmvyIBim8SZg928bmbakotMSroUYKyYigAFHIyv4fBOl9cq3/JA6CreBnaFsd1Dstf
s/Q7MDUfbMqyUhKG+a9BTcOpNELeDTZedH35pcSiz67weQHDdJg2+TwvFWc9dSgRm4GnpEPHQiXf
2AjBf2HdX/MkgIuRm5CrWk/dVfu7sXScQ1GxSdvYyAnFXJpXemgCVwNlWDgXzeQ4l4KHsVzBmSac
XplKNcnaPaa26+cUQLf5P6OMP+mqWtCMf4/fu2Ngie5KCgk9Nd9Q93WxXnjkoxjxkAcel8RtrTaK
PcbkYRvU4a5ZHr+ZxMWF6uDJvG4urbf97qq1rIf1AksuI5aRMUiBZ8AIVM67nh3tCNzNKI+SIO5s
6vKJ+dUNOBCc9CDyl/jPg6fVsgNmOuGH7ChNCdCTwJ5Bh7iubkgudwy1nXk5iSi4tWDD7qk1rXY7
VrxJxeYqkWk/UkSs6iHHk8tXzgeXtv9sZ9oXqaPWKLXij24iAHHy4Sd/2nUGcTipK7agqHCcfm5z
NrUuJOXlT3ie53oE9UZkwNPW3RGqD6+uDweaTj/WJqXMRA79ORgmLOQ+TpC6CQRQV1c4ddCCqcDL
WbYE1FVFdk351MY19jlJkyrS4QrfXAAUaRe99jH1aEzMTil84LgCdtgjdv/Qb2TgdDH3zSWf9bU+
HO36Pu4fFmbyCcYQeKSa8nLtGc8lyevW6bgPYr3ublakIFVkK2/Gq5wXwSlrJ2368rRTggEbHR++
jr/wZGdzYhNnr2lkKqW/fQ8lmiyBwozsANPKqUJVpGFpSqLzry1HbGnczJ2uIF5GN1FDvTtPQ8h3
NPrll1zEa/7mPfdPU2G4Vg8JE8cSnfwd3IL0ySsBLVlS8RL+1AsjJtIIb6GPBLMQKvtAaosrzrJ5
WH9YWuU6Sp+dofji68CkSyPImt4LX8H/gw5a/tk+XkUr+Tw3W81Eg7ZDvL/+beb+YBIXmoBkTDsl
qSO8HYFoDzKXvyFR8AIqhrbz2ZTP0Gh7ZfuhQwlcK6iw4/2RXnmuxkt3+xICs5aVS1/LwStxnVW3
E6uF9znNmF8FV6a2pkmy3ZWfjIF0bxB+io5g4IwXMhkGq1TC0BrI71afluRGPWEznymSdDqaEnkB
hXSPlq2wz0WkgbuRiiEsORzMYqeurHGFtuhop+fjs2Ec5N+kOQIzXCfSY8MtFWus1sAJ4UICMb82
GmCY5zsDTnt/WgVFMY4pVlZmy08GG5GwTUsC5TNn8pQJOiJF9X3x7p+Vx5b5dhhDxvOcij9Ausot
czePRh4UCug/mShkCVtgR+pqViFGgw4a2Dnc5l0SSN8U7PJC6njsgiKABZuwNawW6hkcHxgtyKB3
0yYu45YV+TPrVWK7/ezjjeaiqbgn/Tge/iyvQV25OqikptZpKkTsHgKQ1hro7b7UmmFQcyc3B6NN
+DFskgV6cFgAjc64HifYop8N3gBWmeJoOiAtgB7Vhn2Kym5/rgEILH8Vclv05ejx23ggOK3/brG1
aDTaemOgzk3mojRgMcwUPMky4fY65pml0yARamJKtvRe31WW/qINVsK0V8iy9ZvXxjCsNs7+vtkF
MmSRmm+5yevEWUzvBFwTgBviL29guyep7HbORMe1kDWWHzkheUyIylZzFmsnt+kHyCbFrNbHMWNd
FlSWWoNn+jLfRxWiKJzA4/fGgbFqaMTwTEa7yPybDwtCHOm3NT1w2KW6K6xLBC872R9u4rhkzRdT
kfadxKECjJn1CC4sOjyz0oPQSG5hgixIjjCh3hijkriF/i9COY7TR/SibMmMea9UWJxYrYxRhjxR
gRKyQ3uECc3efGimEStCCvOoyMjQsrkho5xaAbQPCTkjI5iUEmtUaB8nt1MuLtwCo/0YyN1DcrqR
nMvVedDCBvOO9u3/C1NCRWIfs6KSz1ch5GdKrcg+ddUu+Kbnng31bnIuqkJ6DCQHOmLRqzxv/KaL
4WYxPBhGqfh3QQyeFewpZmT5VvL1I8T9RJzmQNcVVSiQrtivWgsWL+AIzwB4c/ErFWO7hot6udyc
KvAtcnvscTtQdBOX43OVlexVPSvjNw2mhM4TjWioeIX65UniKmqG1tLa3SMyKYBAvIGV69Wbln6q
IKyMBaDUiDl0eD9vxjNE70SgbW3D6dCnvTJ0A/DJ130WxIzo/G+Y/GNkYu5IAGxbfKFZXJMattRW
o4JX/Nl9TdLLWh0FTuQ/SJ+TpprfpvbIvikFDOIBcd/GLPzqXYdmfv7jzf25CsA/Y9RdO/hn4442
k8yanWZgcdibZzFSc+cvSvwEJcX8fP02cKGZ0Dmi5ulQ+3o9uF70XuTFdGXOKPkJ9QU7PYXYL/On
i0R+p866WXmahshiuk2AAsHEiNbcG1uk2a5fiAGCusxU38OydsQKkdLGFIb9atlgqH8jymCgcYjp
rN92XQtELwLUBmQOj2WfNi0uZDHZJ6idb4CJdWrlkr4YB4YjZWwwm1V51ggOOHdoXYBWFmfi35w8
BwieyAVPZar1oStqbMRrG7OHYz+fRbPgP9rnP/XOl3JGUwP8wahLdT2s7SilfEAYT/dMHd72Ohxo
mo5lICtJewgcNM8m6dkKnk1LAuGqsWwzV0N2JNzcXSVAMM3AESj7tgBO+3OhsotYTs8M2L7x1dA3
HTJGuzL16VMo66fX7X/utQGH2FjdoruH/fxuQ6Tgh6p6TaxxDCzNb32Fh/MXMTX1BHnW9GnzHw25
7scZCwSyt1SQfGKYTNVxpwZDJpmjT3d/hmI3t6sdx1Mhfzg59IknCkP2wHkEOeS3Zh++4bKZUm3/
MMiTIMr0h6CJ0Jvyis7BqwN26Aqpsr2PcYBFn7MuGFwTqXGzxSBaL62+wD0m+d2i2VUHtDiSzoQe
9wSD2bRTScWSI1qK9jfXMEgRRtLblnYHsoIQohWe/ssch+uQ3fTQUOTEj6JNbb309wyo1KXxR9UL
n3aOY16ELYn7T6k8DTNNXemvERr8RCRYmCeXCq3NRox3UxVoRd4G++Tamc+qrA46v4F5R9/O+PKc
YKSv2VCIcGoq01tD3OWmriTpVcx2PcKlt+ddMfVMUBqpA3BG+KRlMWW/iCLzL4C2DNe56lyTAYOS
T0fUMAM/39NHO7kK1Z5UaUeox6h4cuLpA0Y17MEpQipev/W+3BsLu+aF3Qmu58qbQ1krVy9BVh5G
tyG7w2rQ0p8KAuxYB1Utc2J4ClKb0NEQY2ipsAb2o2t6r1DFHdXnI1gmyBsmZ7FpJRCl/nGSlm6i
HPHmHGVQsl1yGPceB4j15skHl9mnVaHOl2F5zstyKYJybblfBxAct6vue2vddsWkxit0o7wzoKRU
ucFQOxaW+MY6qa3fZyq0dB1igyeURTNUzdpnYvqQ8VgNBFaXzuXEaFVPh4Kd/Grl78sBwO9lSQ31
WNbWZ8uIALkJ/LH0OrBXKggU/+Ewen3YLllZ/UDPx04cwLBSiYHFRsBhfDQo9McPUN2TCTkyKWWB
tQpGIY+8pjaMaSsddu0R926gCABilc1yNKjzNZkaDtQJXinSIHUybOh10FI4j+ffQwTkJBwlTBNa
vocXQAT0NdYTz3JB501yNts+X48kDybUS2r2s8nxSXiAgrMdGBffTKETxPdeWoDlhoi/Spi22flp
tZY128bqLmgVMxyRx4NxqyfOyKzF0IsS6wodFGxgEZZuCwaDkJBvh1CSwu37uWNdr6lFFiaP1HHo
rSTDDHC7NVKdEBCdNwVhwDO92GUlN5yMWGJaAsiRvFmORnxyNQRw81OE4z2LmbFVkFA3eZ0ZIctT
gQtYZaZuGu/fcB1x4Ox6o0Rer+DYiPd8TQtvm/9/HiNq9TqX2K0S3LFBJsLT+O3FGsBB48s1S15e
ndkFmhDEgqBqNzogpwEIhcU5S1LK2m7Lc669jnaWXC7XMTVv8cMiBdwhEsLzV1RJXkUjwdxgCgso
WOITJa+ikdZEQJDeTV6500+vEKqYa5Z+IvPvi3xkB1gD3yFOgc50HFhXF2D+20zowb+1ClDbCOeh
PBumiBQVGglumhOzcaF07tmxlDWZoMkiQd+J7zEBvJJgSqx9Ct7Gl48vwyktHtYjK3h6h/O7zdgF
u02tv3GnCN1d5249lR5jFZUIkddGFrXoIKBjsXRhZ+M5LS6aAeq7G7SPhr2kFK0bt8b0JaRHzTSg
ZNeESDXIK6iPSWjtgVgKHp7kWeTNeRLaknxX2cH4JYP0x66Xt3qYjEKVao25/Ul7ztRzth0Gm0Rt
MyzfpLYoKilvgUMN2SHQCZ/NgGSYCFn/ppA4z6mZHXiSxn3h4BkQl2+JIPivZ7W76q/g/3NjAR/l
G0oLd6OfpCmrUKjCLn2YO+wF5RNA2/IastK69vhp1jw7ae9gf2al9BdyEwzwyrBqewR8eRW5+khL
S6jaZaAxUHEhnLLeFO+Te/6GVI8ADlRmNHzIbSzFbpdT/OgEN0QCuh5mqZbqv5ROhh3Hq5R3zSCZ
FV2jvmmIW9lcFDfjRaLtfkGMazaVMf5AXuBcXjTxnMuX3knoosiyIbWNrR1jvYSVLOGUFhIecMzw
rCEh4JMyJQZNLxJwCmhTPz95UbjTEBEFtpY5Y8LOYg1CRplkYf1caHYo7ZXvZevHhCLkyX2hoClt
7BFeosK+nuHMPZv1iI+1+PN/UMC6jb3/X3eUueIVn7oPIBpb3OapsCQwnGJ36ZJpsNFSXBcXEDmi
oolORlsdBFWUDX2lEhWCBPrI7bMPpPvcy7vg9xPpkwYx1qx9QBhBRzbJ7HackAw+bsHdZruqhe6D
evSzz8uQkx187FpzkXovtmyC5qZvJ+wCMBXVGWFq03fUhb6u5NRnFrt0sKnW8O0ZGBOUEiktt0xt
Sn3gtLMzqoL0xLgIgwbhfdfB9jBlzG/Y/LiWQuMNrO0aYe9NDsGeayax8Wmbk40CeenPMwVC5Ao/
5fqskNeac8G9jhinS8lWCSwYN/ReGr7pa/ywZPYjxvuEkTY+3BjSWtYRN92M0TdZa3UQQGAHzlNg
mgT3e+vV4CI2CHCd7KJc/KmhBmze5igJkexiJDbccCnBW2vFiHJPqb+dCzHn91pV8nQ8Idga6O5f
i6cEeAMuyPYPGsfx6ZVh8Yd3yOf7Pfj3mutGliaN+WSvyrZs8+7KI7WVWbSIPlUXPkOcncgwRnkT
+VT2p975itKWtBc0TD9GKwF4Uj/BxFyAPLCzT+1Eto8uuWNHv4O90AKW8KW7+1VKI1VDC8kb/qao
8G6g9hpf83e2YZ72nfXXlqfEq4pd591nrn70G6W4rMGEFC7FcZ2TVAcG2DkKMctn2NigdIXsxYV6
Dr56rCQ4hnCf8zfwaSQEIwqzlAwAVQdRd/sOiggG5/rXGESK3yRpx6lUSjN8oAmv2jzEJ32fVMYn
cyz5NDpeVOOylMUTrg7NOCbN3a+0uVu4KUsFol6Ko6Q+ZLVGELE+UNoUBRx6y5nsBVRr+midlhH9
qR/ca5SCvB33noQknFqimDNXQYgbaSRuaGf9dVaGrGoGOQsGnOTO4Ce0gYJ7G/+WSlLEre7GrHC/
cR5eoD7M39oK6LlwRqKVdf0UNrFKnrtwQH3jQkYrbfUV54bY8TxVTH6fmhxIC32GQ/XVdndOqxME
Uc87hWrnZrFF3fk3+6B1LNqOReilq7+UKAhzNV2VUtR4o6GaECEGPy4GuifXNRl2irI27H9ydI6f
1EpjmrCir77MkHb8FRUrJwoCXmD/kf5aTtA/rshh1EXU7LTf+g95mEQeFKzyUGgRKDTNttSr7xyh
s+uVMF755beuxl1/X8Ru3N4POPkoHsd4Uoke0hCAWJIwshkfhn13X9r6Io1s6qn74y8omVHnR0jh
ac0qcbX4Qm7oXv8kBLnCLjehJHSWkNR3CwfcdHW9msU0d4so/rtkgt+Spvza/I3cExQS8Zw0DIre
x0POFb6W6NNlSOf771gBDiXroBmbH41ps2JoNcLXNbTuIP4WLjn55lWu5CPEElmLP/W/X18f27yw
h38J8t0DPYdWFKTwwHVc97uPl7MQD0rPqkomEkGLMZO1kgSxe0QHA/1tOE7NQ/CTIRl6c6DPLJbA
Hana3TlJU/NHGRwu46zrHm1KbvJmPYrCdVAlc/5lma4umqk+Lc/Qn115bS9JsM3/g0QyZ5CpMtn6
w0TSxCqQD0Tp0m8+7QrGILpCWJmVb+fUVVv78Om6jFwLQAcUBaXCSJw8ey5tBtQS/1p9raxAIAEn
6U63aATi59GTyo41/5LJqw5tGk/MccUjZjmagVkMpIaA3easaIpzhnBfP0z/EgJHJ4WPovq6qMne
nPShyaYGIs6NiHKB2t8R6iH3OouFBSnQyuylOImWNkVTMw4sKVl1NXG8ngHyCMEpvLLxmbJamyCh
v6DAc0Z1ljAjC/udF6nJmGHNTjE1ScngDLmxKsp3q+Dtgv967XN8XrzY7zCfjzmhjWj+SGPG3yXU
ZDHEK6m34SqoABYw29X1SMkFdPaMKUKu6E85QXDTPSyJxaJME9LRwSkNYIX3E3JT9WaBeTR882CB
e64D3fkrFJ+82hR65T6kPT4flS4p4eRKwla8pcK355ftZvKhTuCqZnChh6MVjLi7gHjKE/8P+LNx
2ydl+bvR+1CGTEFf8xgJ3E7PUfmw9fqsLF5Tf5rkAgmM/U0pw6LwyItRxVxb38SwIzsOdjZxxlkw
FyWugrzaccaaor3PMmYjDndEIiuRCiokC8B4fjlHEGmC9Hhlhj/BwZNTJH6veFhan5pY6R5Nc3jm
MiccpX9FV4nMJR7atrgrpPYH6Cr5xXo8a4JKya9ZsnfWP8LiZRYBC4c7/dzHHfCDv03d6WHlhvB4
WQf6aoIrjEyJp7zdDjFPKA6tov2MRXHjrx1NScS/7fzzTbx2mY5JWxgMrJRMixWDO362Tirb82PM
DRh/NSOcZ1twouKFkdXax0Pem61hwhR5T8eYLYgo+dqLFvlMEYPcJh/4K4Du29CU6AkiLXwEGv5+
cpW8NnEwVK6/oaHHzwWi4oWO+29IalqsoDJeMumYwkF+eFaCESgfTtvE+v7aUmR0AYxTJD0SeQxc
BLSPHHzB71zsxl43ljon1PvP1Z/hYZa5KEgycehPzM+li5QFavKIn+oi5/6YRNDXIPjvZTTepyTQ
BtMfpAbYlmm4raca35Qsay81chvA9XkDCLl+FWYojbJtILdjugsHnwAph7nlHLq3YiDKH4B0hIzp
FRq8vImFCF5RBMPKgV/mRfks9jwxe1bHaFb/Ibq2V4Slxh9UIr6+dBowMXISRMZdfKmyeQV6VT2e
DVSGX0yxXC1Ln9jWuc1Coqm6IzlHC5iYYd294GlIvj9pTlbrOL333gtfu2ji35AXlznyaXyUgJJH
bkCRBpH8klFh3Qv4sAgpuUrn1wD1FjvMeJ4qScwCxhNUQJofTDbiEZHQCSZQTBYBqgEPVcB6Ogag
PPQOhx22DusWePCgnyjx+eu90oVm7uZTr/1vfdeUkM/FZiDyfV87nHYK1kO+2ha1qDURO8uOKLdj
5KduD9Ive0aZNJEr5TEiG6k8/EJoGC8N34zlZVyy2GATcJd/nXU3hqgAJx7Hu4Iu+e/VDMXdBqMV
xPmp1IFkT7dRJGDKD/br+7nFGNd7dnL1NESfQ6ZcVgqjk9aVyHjLtKEj0QpF4ajrqs7+fkRYTq04
suiZG9hgcivdbw+4mjrd28r/gd9q13pRstSC9QYk00K/AclqzqrvtMUusc+XB3Fui2yn73hComzX
uVIZ2yI1c0SukF9dESZlFXPg4K7vbEtCuebRe2uraGONSitEUeGUCAF9Rfhn387DY5Ss23twoTMN
OwGMHK0LxJ/hVCgRs5rvJ5OA+UTupQJF8FCkEMngDCnFf76CN5GZKb2WawpK6faWp1lMdAUH7RaK
Bdp4hE2+Ws+sku6ez2nq+t5kWUeUigmM3mag/lzMwlsD/0vlt96HdALEN3mLOXA8IDTxvE73uxMx
kieCwqOnM7H9NOK10/othJwHf7FLaT58PPPanpeIrma5WzuPkBL2K82fIFKIsGCwWzRO+AjcqxlJ
Ra1w1f2HqVhSlnAiVLLsgLK1G/FCdoceeGta1vv3Y66LLgoXY3dTtwpJdALVUvHMt6qfyQ/jlE0n
X73VKH0ylqqR4fh0f2s7SsBCn4vVSBkG80nQ76Gi89s+UjNaSrtzGGPmTDmZevHV3djJHRkOnjMM
IH2eLgJRwt0mbGBE0hnEoM3IDaviSQvwJFQ4yLX936bRKjByY123Wcm2Dm7e7OBe96aoHe+ZrY/E
5Q3KpWGtxYwm5BBc/RvwtX+3ruMRVJrT9uCBkAd1kGpjLHiJCCXCZ8FECsWK8JI3hWzNBUGSauET
6JfIaa/2ByQBwvSUurA2ZQcJuvCHT5xFRD3jcR5CQPx1pbwE2p8CCgbAIBysggC2LR77ogWyqgli
YRBU44EvlZdAeLC1iPbQaotXR1ssyyUENrx7PUv8CsYRSBtpXrTDSfDnPUI7QxjCiG45dBvR6/S1
0MAAfENh5FqBAnVy154V4C20wbqwi/1MulVDD8IqVGl9EBxuN6NVEW9KWV0v6R/uh0l7WlHbMdi6
eDk6TD/mwRrg4H95eJXO4fr9Y9pdROdEBd/96yuadrQGiQhWaHc2B51Prbh1YmTnyp/zdX6vj9mh
Qizl8MxLWeE/HQbQ+ZummxwrVC6yhA/pVBUrNUMUqSDRL9X4edJAtLjfVkP0QBncAThHL/LutvgZ
yuORp9ToPPaTvU9O1aRgVwA9m7qBeM0Eb5hLwz2WuDV8e88uhNP2s4trl2wABdlj0ZI+ty60lTXB
FfTqEmBJGd/Imj7JNDG75OFR55u5YHhKG95eCslFVeSQg0+iCIB7LTfQ1/EvPUypAl2aZML+AbgV
fJs4+0b1OrMasdUvkvQTlcv/d3C3nlyG+MB2a30ewEl88b+cyC02gHVKa0m417tkajzJY9p7ozM5
XJCEBapyNlUgLEFlt8EScWQ2HfAxB14tDKEcdFHPGQhsFTVKb/ufHAownRTALR3e0I8O/0IktRNB
ZoTGKIe+YjfUITrr/N3J4edQSnfrONjlE4/PMm9U9/romQJaLzZB6+oeKns3+5KJlrMFCNwQ2rJ/
bJDzudvoFcfkEa/KC24zGIaRSghJk58fXRCD5P7dRewUtdnCNv/6x/kXht+hq9S7pFT9ArkUKZtp
y9hl9wY424lkJlyM6wCh8NkNlQdWTQm3nz38fHc+nE26kqt5+uH6I6ZHBUazmiCmB8QxJ7G2Kkrt
OEPU37s8UnLtwY140cQ1j2tpfPuntoKeszD/G4kWbY8jzg4hSd263a/W1aAgATW5rjzW4LVp7XAq
g7Edu7vgS6e7bibsegLljsQPeXL5wV2A19wOHLYwhz1s50c6yY4d7M4fvswzabz5rrpNLedPQoC8
VbXbmGJhcir8JyIHQjrDF6wkJkj0QzmWCwshZLI0fWlU8Bz+bqJXSfL2tQSmFyrqJDRsqwjpII0O
dxfphiJKN8VXN5RID/8IVoLtjVvGYo4kyTbPc8aKcLr947wbf4T/J7o825+AexuZGfDqFfOt8b4v
USvNxHA3FLIwEPNe5ehGJ6z7ZnKbKvPUz0Kr3O07ZDJ5AeWdmOYUNsg1taRnw/OpXRRPeAX7/qr5
WkxC0XIz9mobkQEuwmR4lcTYztbA2yF7R4AW5O+t69OdIn1mEM0OzP5VaUJQLlEkLNawZbkIPyTm
52TV4i+nhWGNez2q4W238IBDMIpCxMyk0/5xDhv1U7y++9vqG6N7VOU8AMl5J4NZmRHExN9oMoBX
iF4AW0i5C+SbnloCquJTKqOLtPsvX5dQc3hGbSu+lJLfc3rV1QVjFQDbvDgoMhzI4r3FyG0JQlzu
tXR4xR8Rss953GmDwa6h73dubjtJtz2W45R6nDy9fg4um3O+Mb5z/gYnnYR7SZPBe+AWdqCWXPfr
nCmSmKPtnj0ufhDvEh8c6BiwyRG7Kb4g6jpiQ/aSoc3qELkJ6JusG3hPpBgCXWeC85Ub2QYpY11r
S3NlLQlkn0X1Sgq2ZWqEW+h3y1+5LcwK6JT2llvd66aNXR6adcQJGl3+AjfaxABnsl/rQ3EwN52b
2b6r+67l0K/41OYydkCgdcFf8EVoZHsznbeLGXm+t25u1Wh7mEYcfC3d0tUQXgnon89H96afJvvL
H9PJEfO+duwf6awOjQ4VPmFq0hD2/55W0m1kZHL9dnEZyjIGqfF3Y1UBt/TSv/O6CZHQRHvnILdD
QBxinZEZwVaN2CEJ4wIjb6kLXKUFh6m4z7j4RRZzuczlifBUo/NCHXKQid89G0G5Hr7T3kQVqLEe
LxhaF/BeNRverhsqOrjBMhcWwSmTrC8ZEq2a78hYjeT5tX3XGYV8dEwLXFoH3EV2w/Uoi4tRIgWY
iarxSkuWPRdjw7Zn5pr68jpicwbr9frFRBa+tv6+zM0zmSVRtLpN3jrFLvKhWzIl1Acwscn6ngGa
m5kfH0bK8jIBPB3MPFc4cxvWaIb3ymhh0lSJISVrPWzLIqtKNn3vFIm3v1J37hFavS4keyj3M7Gv
QwHDfwgZWzhI+c50aIuhjB3f2x7h3QI+pDJVFJUBdH9UW2I4qZHB6rMdAbYK/ZhHfys8EcfI/24U
V5hY/XHxMfdLxjnCI3OdVj0RkQG1O5IN1qKpdC0/ye6lKsdCS16G3mdnSVMBpb1WCYwKrW6awqGu
b73UJNdiN4tI/dASDJNi19DRMRZgGHIOLQCud+RINils25WOdp8VCkAOS5Ta/sBMWxDv/qcY880Q
25rYK0kORcVtN+Pi3tCdwDfKAwY5v+bvH6La9N/V1vkQFo7rIZ1TwPxnZSXf2cJUNwVjGFifSPHQ
0X0Da98Mscwfi1DJ81kqjdobY4MNEKhh9KaHXRuRbs+Y2pt7n2ogYP427hROcCLHavxJstR1yPoN
KKpWCt0lsBak0KqfXcWnGig7y/E/nLHowlbHh+iEka6tU/TyImsgAUDSfAOhXPxQEz2i7a2pzekP
EXmycWMOUtyImVHWhHqJQ5lHX/TF9S1XXJA/IDoquu9LPo1CvumBmAp5Cupgc7VEhPBIqNjUMkRg
O/V63SHao0cZszB+ZxM4g7+cyKs89A/dzKXR8h+WJ9Ml/QCtGyKNH9A7jdc14NC9u1gJV/WWSXpn
QvyPyi5o+6e6WIf9tbratvjISMTPedWHrvJDTEjKFsBl2QvHTWEW1q16+/9NvBa54XsLNVkUkcYZ
tS5QX0iLDxdODsipkNENRI2RGclg1kABZu+Jm44IN4CJdZefLJMwHdJlM00GLlU3Oq3cgVRIBQXZ
ZJLYk48PAB2UOhQ5u+VRDB1coSHTPRJ2Fj6gkPGLLWZTr+ONYoveyBwsittg9HLmitk/zc1jKIEI
ZE8J+l/+g4LsaI8SSsyyJnNIRiQeG9GlRsTsaPWAZeMv7ZpSwZ521cTM9CVsdLfmThtoD1zVBD2P
vPrSSqR32g8AfH+AIr0yp79OrPMW1NthmZkCQ4Qb1dpP8eY9LdVA23rZwZxz23gba6ssoWMD09Th
/TlFiYw+diDLT7d3pZy+qD4U7UlUlKI0s3JHvjihmSh51ajVLQMypay57Jku+ZO3r2aTN+ELjRqf
fI3J+yZ3MTFeCbuvfLVEV8ltcPeywMaCJZJj9HKaDxsW28e2n6lhdlu61fSEA0Shg1X16JX7XaAg
AV1/2FAkFyfWeT2hPS3kKqBPUHssVn/q7yRrkyUmyx7dsbx1O5ghr1HOYUDFb+rGUWy4s2RlUlTK
0my5DbtShyvMZP7TFpc4bgvsju8eDWgL8LENKZMeNbQn1VVt7HwqY9X1dWyTdUnC4nibPigzqesX
kq4Mm9Z2kDGGP25gFATFQ3zTBnRYk04kQh1Y/x1Lih0SFbYGBLgH6PVxYI/IKB8th99Et8JhUdLv
V0joAQgqFUnT8/03AdRpVHOOHXXML/NmLs8BA1w3t4uuq4jodNOyRG0FgZR6hzn3SZIKzr6HWCkW
MY/+vtNIUG3W7E+R+hPfSXoBuyiZh77ewXG0szh27Lkh+BVQ7T+rSDObllTbqzHql04Hqbd0lsi8
CsnOZH7bLvqLBANNECAEZqP+STOH0xxs+6LOS2gH20ESP7xJn2i4TQZma95K07eWmMMLjDsk2Bqy
DIwNsARPt9cL0viKYsf1qHl27Fp3a7rD4JZ734TIZgLaSh7TXbRxFl1jpiMjzJKuodSllGv86hKO
oIIeooqjLG61zYz6ojSTiuDPZ23gez6qxKFw/SvlyBTuKfLray9ja2ceFFInMvOeVNxcQ/d9EuI9
oO580Kq3p21EoVqatf4g0PhB28QZVTN9xIuVe68reTmj4/znqw5cIhEFm1YWEOHEhmOjca48wZjS
yDgS0Z5gPs3aOKbkIk0limKnNOcteEFa6XxIK0hxdi3+XbU2dTsxOZP9M0I9YIZYSuNT7WZ+LA5I
gtdQoR1ma8rgc1UvLh2FL2XQ6KufufooDaF5GcHs5jIQifAvPgx1GFhXDpBQGMZCxhRj8QoflzHh
3GweLNplc1Nh8p38ME6SEGvvkLmwI85TKk7pEghCBgCSt9ZfZvoL4iWrFsU/3dOM60EWyWq3WRKJ
rDP46PvH9FQXvRao/1hict68382Ul6Ia/MFdQsQULsE5ZjEQ+SA8shdvnKe4/3DabQ2R8sLDmoa9
bmD948n2HUv0ETBFkemg/wJc6SSyf6YQF35i2zhbfJjKjJCOlSX0hCJkAtP3IeP2XJjSTg2LzU8/
17xqkO9YRNLu+nj5UskvAbffns3r5+KuZFrEvEo5hzAEyV3tuA0/p86hQ/d9Z4tR2qxRWcnO7vSb
zw4/WMpqbwd6SFpVETiAXHuISO1tvWg+YmvEVePa0KeuZ0+Fqsdu15Cutw4gcX7WDWQv1FSP4W/Y
p+6gSBWqFV2JW/KRTQr9LnRi8Dtd+fZeIlzllYaKV6jJ+z8gUDXRgodUORITh9oOVBDWVpCmtOMU
qA3cq2kasU7KiNJBREFxAsyjCrVUZhG8KrBLpS+Vb6Drj/0kHTR/pnUIluogcGWI1nAgmPrpQ7eV
7S814RNLdQ96UF9GcRnrEOOS3a5OaWl/gzTDVzE58guwo5QxFHtdekfrL7Palv5FqQ6iuXtDAYv3
3xcnSSzB8rDUmk8OR+3+Lw+qjmqMQF/wnhkiCPguGMxcM40pD+PeUOxP3HkdSRxp//VtMZLmhQEO
yRdxlQNz1xgJhb7Fuz+oxf+GlbREIq2yo4HcQlXUm/f00HFOiZ+ojy/re2q2G05sbqAvra1RRPAJ
feXGIEoJ0wp6tyFY4OkwvMDZ2dX7l0IBnP3k2S0Z2Pl+0WdoTkvpQQy0R9PdiBR9yglBDCNHEPcr
UAM4wX49syPYMGFhsly5cuEhxwc9Z1yH7LAx2tBsi+KqyWsMNRZJmVESUZ6i7mH5N5XkwNVtkdLP
0e4fJ/HHHycYOQf6/tcTDWInScwGQ18Y6Kb0dIC0WPZT/gSRSUkGWiyqjMTUr4wkYX8WiaUQnesw
OGY6xdaNkzmN+Xr6d6hm2fU6nwfHiL+4Ax0dfdmZXLsT4Ajsoc88876WMTNX9MOONo7JDE9mE2A9
vdfT1kk+qAW014Kf48whAwkn2sgTwAVUM06R80fq3FV5gxyVUdRSbJSybJqKzhPa5G4tZfvWvZm5
/UPynQvWN4Z4NqXlpLWNvsQoKx5B1OrTOgQj96oksG74oGAWxS6IEBVkJDSOU5RouKWgoYjRcAjd
5L0ppLWXm2y0XkqO4UzYJY4+tUxsQV52sLGXFlyX0SZ/MW0nNA80uFaNYKfxwDigdqouuGQAsaOZ
2GpfJ+GnNoGxuEjHrpsxdcTEZi1zjioY5K4QKacchxEBM5WHe5Ia+pXV6tauNP3iautQGW39GJLV
TO4DrHcgAMtNkVo4SgBI8E44uNwa0nETqKpIDktbMmicxWHIgswVG5yUxSQK/APv8uOW+kyTLBT+
Yku4K7tprykQNLQSrl0NnlF+iLEA4d4x+PkP53F3i5KBBRTeMx0wnfJmaAVz1hxE8qfqie3iDaaO
QzjYXIfbVj0pKIJKAZ5YDJ7g4lqLV6Hs5a2Ma4NVe5NfDsG+HfOXVSjAC2rPNJSxBMI9ndIqyaBi
l0vx5ioYB+xajTxYy0WmC2rsoIkPs1d7G1TcRfMxOkEBxzU/kMkh7Fze8twjRIIHUIQeglkdDH2r
7S9NeAGhhe3aKiL/28VGxmcuj/gxHsTG2SoxC18iLQ1e6ZQkzhisKDvds4mt1hchHZ01roz98Zxi
FEbcQW3N4kFcKnXbR4nMwAHc/yfR1nmIzjwCe12515CbY1GJrcDVyMQddxYEHAJeWLRO+MU2viOQ
UreNA1TCT9bS5GJ/OKKvUiGzRRsrcJMHGZLL41/VP9bvtWr4qTBeSPPygQgUESkx3F/Zx9BOn5Ja
uR171XlkFLctIs5lyyTOuc4tx6sdMmt/aaO3NVAKDRLn8QzIE4hsOklgYNbykx9MwEf3YLrIA7ok
fHpOALK5NWP3dR974T7xiiK+LBiSXNhvzo2kmJD5/0N0+6BB69s8VwoiUjiARWtq7/jM/Mm17sOm
EmMoQPw1FKbKcgaS2xbQE1kBQOEdaFvURlFcJKdLoaFnKlGPsOiYb5gg6/KGYPrzXyfIRk7JkLoA
ffXy4lGLOZrJP/kyf3a9Hg48mLZWmh3cGW/1RqN6MmZnEUJLhNkO+DnNjLpVhrNS7caMQnawD5vX
7ZRHnLBGOgCoLG+tIY3QKzNBlxuvsGmseR34qp75Y8KsXuPkOts75d8hyqmXVNFG6sPhupWbkHTW
FKLXZpkdlW8mVntCzZhgCxj8fDvDHin8X54g9PXuj3xsjHsLxqmWKE7h6goa5PrcgxL4DVUuu0EN
BZ5MUBDtMBsUdxG7HEU3ZneeyhFTnv53aKOwN86WwSvxqUZ3KM3dIfTkeHF3PAjMIWI2Jg6d/hbF
UiCYiWes4UAbJRqg5Q/WdBRqkO7sepjWMqZkno0fJrlY6LTVHItaSUjrkfk6Bk5+GfcgUTfrXxh0
pIsck4qDsxl0VRpBwhE4XfgEZ57SzgptyE8UqzqwU+1qS09/qcR0/KBmwMzV6OPzP7PEJdeMVRrj
r+VFTAJ1ZlEyOgugSiW380jUYereShiIGX1h3zuvGqOLEsNQrN5hcwQ0mO9WRlU5J/0oACvaR/16
GZQpc2YDKTX2XND/V/T6w4OMVTOaFW4knPZAPYHI/ZvIeUw5Z7LsRpbxT9BhY/lrA+9wXSiP9pZX
pM7p+t5PVBd8JSqx2D6WgiOroMrIzERRI7Fiv8TfqyHQo2etMvxed6FCbchkXYKk/H5qYtiNWOKr
Zd79ZK1LjLadfDkmTbMjuEuPY5LHMX03zzLILp0mQtJALdYd6EY4D0JfpDIBBN2PQyYqDE/vIdLa
m1n8h+C7ZVgNJ2Pd8srruJ/vcvKCNzddlayYdhJJAj0Ij7HltYZD5LHbFBAofBKUt4addhM13Yvk
0SPSHuKqdl9/n7pf2B6OKz8/gQqMKLpNsz86SQrd9ayk4QF9QTHuXO2i2X5kgeYI8G+a1NpvpiI0
NZga696Kt1TQd0eJxm4lqcQYiVKqCsEuxzIpAQEU/oE3Tx4pnWalR29TBw4OITXAKVoW85DFIJMN
Z4zWVrjq6cNJW+kbzHNhmD2VbL6I2A1ft0tWI2e3xw4vEvioQpjjiNBB80pmshfCSDNl72n+WBgn
AOM74eUluT1F8NKMRK2MtHF+VHc0sDVUXXlagsWz4AXhsiJ6/hx994T5yfTseWQ8s4m2gtrUuXAl
3yep1I8Unzn1CaQ+9EDzyFlbuLKKz+QOQJEtw3HN6Xai1X8zH7eO4gzmnVXkZUfpYzlpEEoq93G8
EvFRy32jpSi9Pqhh3ThLLjvBdR/2LbHLa2x6NaSMeFv47DVtWwa0eYB4+nJgB9mDg0Qnnebdgppy
k+PjbepNczzKCnT9m8IY9qWoObWogqeOFWrywe0hNLAwbYKtsl0L3GbppTliI/85T2bN1tiFdrTJ
2wQgnHDu155BleA4ISKZ0yIAr5s9imL9FxRXf5AY9so/1ywZ7ezbkHvQf8m32EzJMChnaj1OSjix
iT98HabYAqCzVLmR/npsJu5N2EwlquJd3CtP33YQs/qrmYL3xlewDn/y4qXIVXVUyyhxmFD8wcrh
cQnYtshZHN24XOIpap3huXOO8yqr3sa/SYrYukaD02aZ5GSFpM/lIGUmmQIKzl2b2KltACJqhbfN
ipWAYqe/NjGfTaRCLlfLoNPTqFFkWHG+9iPWfeQJhv24S/rWc8vRPDUDwYpT1cMFmdjKuJDTRl53
6wS2HWaTmTHA8NrXoI3qv0Amck+OES7LODKago5loibX1jJwHzsVl4/gx1mwx4bBldaKwFu+QGEx
8867O3lMIQX3P85ceDZw6ZTjsu5XbIPd/ka335J0trek+d9G7XbiYmcgug65y6yKgnQ9aEgHtDyG
lcalw9QGK+dFpLSfxaz+4HItY1N15I++XP2PLQxyut751XqYOZGVapnlE2iKAU/kcn7zjPB5x0v9
XEGy+7UDj/VRZaTd4Ou43m6EmNdzdCVY5ydID36eGZKToelr220aUldR+LVt4iF4aU7rrySFgxbo
kNdLSO+Vr1U/nGnA8DOe3KyjSwqqdAwqZ3Ffz8re/gVL4VKE36IVQCJzKAcD4Yg+SKmyVzuYGIUx
F7OuY14mOV4r5jIntVMzwA2VlGFKE4LBkGM9Nh+MATbT7uFzOX5pk0+1IeBxgG9e+e6RJYeDHi6p
UM+1bYxL5wS7rPR90c1DG1A2T7jfugbtXU6IyncLzs/v/0svJv7Jot00hOklqTzaCBqFHm+M8O2R
nafUi1EyTQhrDJ2TU3QV/RwvbjYAabx/CJr03/4oSfoelcoETBvuA4j7Pr2NZp+/32hvR5HakEG+
koqjcpeDVEd01j83NHs2MKIDqyf+/u05gqMc8d4er38WO1T5hp+5X9e5lqXsloK2AWIVXBkxba/2
0YTVTWSB/l+b/xbZHLmFsZ6CIgvFiAOtjZXXXwUYcdK3CLImyxrYzmP24w/I3vtdCXSSWiG/3D0A
yiJQBevKu+oZJdX4+B4YhlfTWJFqFJTPPGVYiRiiX5umsPAqdt9fW4jxSZcJrHfsp95sWLPuiKrU
iCR3pRUa3/o0jMM1KDkGjxB+lfJ1qxiuQG/5La/w3n0EIKaQi58RjYZDY8JQavHOAz5yu48wiRWu
vRmGCTSKQ7NLFqwldqBSvtWJG9Fi6JSbvCUb9ooBvvbg+79E7xIcmWGe4GU5LOPJq/9nSi933754
o9kCwbzHoo5LYLoo3w3LiKRbY1OcgPsYTNPDHRv4pBA/6sQiAXI+seOMBY9Kc/JwQG4PAZufrgjU
bjj2vpJbtmnNIAra7KIm2DSAHxcqUYcEAzjACxtQ8LAD3EZLBUxfYqRB35+U5PzPaU2bgClCycOw
mzIrWItV9J3gLH9vBD/caX+ojv4/Wpd7BxNLAzIiLWeUrqTMOtUsT5ZgnAdE82NR50x8CJbQbiEY
3jXVkcu+E9vIk0geOCBY7WgkFoEb/vF8ptU7AdEpDMx3OqVdzCmGUKgIpdYC82u02/C6m1oNw9Bd
5A5Cfs9gSQLXOsi2Qxg2VCBJZmA5y5Sw1VXHbOR1GKiyA23EGCCyBMbeyJ4edIWwH4AtWPNkWQy+
Oom5VbGNWuh4Hb8aTtMIADIYGEBTpFzFxvyBQwx1tBnAsY6XTQP+fJWjWn2pYANqbGJcvccxzLjC
oh4rUDM1ranRy2XRx7eUSufBHcqI0CWBh6Eyf12sVMfdUFuk7Pan+CGkcyh4V2rgQie2x20Du3lX
jWfDHG4uZ1DhZ7+u3kz/8jLs8prt669j4GTpkG8Sx/bd0VpWcAy8ioibZGg9+RDjYlGSNvGzQj1h
YtQ1mWGpQafncdQwhRlXi4cS2EcTSMswaADpNztg5BL4logS9DmRoR/3ltMYcwzQXXBMulWxH+bm
HEiBj9Ofn074EfxPUTOReHwB/qn997nKuP3D/S9CNbL27GThdv+MFAWvXiPIfnw4AVbVZIeqc4IZ
FZN+neW4fv1F1sw97ZuIovNm1UzUdiHs2aaGHu9ocV97Y4Wn1ezxnNALA1gAR2JDNzde/VsvkcaZ
8PIo2hl1401OlwhZGPZpGO7FKS0qdr7ThyTMfaCiNDMMecK1JlUejjjL5lbZXCHtC5A0xRq61uWG
DwTTpprpNpRNNsyXoiQ8ehz1atJ9diLhOzGFnJeaHiHeAu3ACHQQ48hR7nKWLwFK81CW/YQFXNyM
Ggt0jwaQn7s9sp7apqhsPWNZq6CsUnMIThZAakuDMZhFquHKDFnJfp4LYr4DtdbR+pPsYki+Y/sq
bUtmIGAQvazmEf+uHV9T4u7U3Az3alewhn1bNn4W04BpYkXQvArVhPCzuWTPJ0dvsEz6WdKn1Ar0
HRshFZglVk323maVn7JcwwP9BhG5u5ycTImimuDc+uBxMF7LQCAV9amWBvcU4m9S8HwLZ5s76V2B
fp/S9DAtUxhhJ4xn6WFnBYopMg3HXIUG/K6NDo1mJXGdgaM84NhHJZJhcOVVj3AX2BBFE903WYY0
LBqlbc2ZK1eRHRuksG5tIVha6JXzYygxoc0RkgNgNPzlbXyDeoAlb/CqeNeMpWyhonU01pC7MNJZ
JF9ajxiWVWwaUYgyokkz7dkp0Dl7zS0pHjKmtDTF8276XIW2wFj0io+zIwhO8UuxaOcHxTo5D0OM
Q+/nL9pfkLcLEYYOzP6lgGGwB0sltYnROKHVxwtyl+OJEPhTM7FuO/jwv6JjXUjG5D9MtzkSgzAg
WU6/nNHA/uXZnUVw2LMuY2UGtrfcXzlH76+k4t8/jkrJBlOVoh2NS87fL2xzXkEemWMLoYGlTLmA
BQLX4JQZWOi4ILeXi8Jtfi4Wu6COYUgKWfNKV3tR+Wnj7cH4zuRFWY0gxNP5EaB33+aXxdh1TwgO
qxtIPpJs+nfDyw3tQJhBw/dmmyLfIzNRJsFgj41nbuAXEvQvLB5XLI5IQkbsKnYtG/a9lAZ3J2mc
oH8rGGYTXwmu0JAbdu9lF6rQ1N1WCRTPqo+abW0iFt8sqiipJJMBlznLO3gfsAci08hlrgVui89v
S8bADiQ5wTsE34F9THOgG5Sjofa491I46u41Q4g7dXgGDb63MVXMUlHhokhVauShGiIjcERdQfCl
eRYnxgtl4MBYNYifvLFyb+/7OGsGd1ECWGygm5RLjPo5+FhP6ffUK8L1xr1TDMqWqlLDRRwn5sof
xKGBMu/beB55dED7l9KF21oOP4uMt5I2cmlleiNbbm/j+DowixtXJ5JJkcrIkHIg/uN1PucRvh3M
m436VgmduQlDwAxB7skWhItKeJcQ2hHDGAOPj1PT4Ovp/7n9fViwXhEGl8mV1lk2CceoRbaYZlqD
rBtMh1HB9VVxNC01JEpp7v2MCN8MVOfMzffsOH/CVJP11OLLRfuqYaj3WeVL2SVxpsN3stgJOneM
RWX4PESn+7lp9NrC/2fBESkfkt0ce2SQaB2OD8Wl+ifiqNgMhCKFWivMloCkxfOfUSKhcZ0lOJuh
BX+usyg/xSV5dyer5n+SWWoa5DrAKj8EaZPfw43DPvMbA5wLGsEolX4J8xPEGwdSOS4CNp8AmrlY
BLPfqEBw72JTaPg0V8ZctL+5+39g35zIR0ByZRNUyv4oyn2qrcrnvISH5139UqtWUxdxTYxv40HU
cissKODKvhOJkru0vjV3GdOHrNL7iKJgMGb7DKXWNjhOeyfI38J0shz1hHT3gglkEYMXZVb+rjjQ
f+WumCjmUUmaxPKVN2Y36Nz8jGl4k6gToEybm1/fiEpc6zIoEWia3ngpuZcSBuATTwz4nzLT94y5
90M0SCtZAlsyllCbokFkAdXqsJhb7kjcC6QBh8Qponzoofox11VwqzCeOo0vBLanQfBBV4Ny4TdP
bGge1O0RbjGIcJnMtxMnvRDPefhuLpInHlMtP8apHBhtSSG8oPWnAkcOg+Tzq+2hSQTWtjGD2Txi
wAE0wfommPkTLABNgn7l4Enqiwqx11zem5VgcNMneh3V+g8pO2hvgwwnftHMjNaGCq9G4iqJ8sdv
5ND7IUY5MrGgtJ9k/kpMO//3IQMg2aEqSVsw9SezIgEoqr6ohDxgqdKPkEQDIMxOAAYe8QPJiVsz
b9l95HQp34H3PCITQfcl6o3vTTxAi/y8UoPI21DI6re5cprfmPOqMst3aDRXtOIUMT099OSO/Ab7
iV+yKgxoyDNftxpuwZpWDxaXfVv8LAjvSKxeSJG7UU+OF2G3fc74Dc9KnMWXJeacbVEYxJphIGjc
6Xoft3WG9Ri2r/yCdsVxhsz88FF1QpMmtiPVCSN+DwvxZ0peQeUadeQItukc6L2pxfoLzHztOxRv
Ip2d7YUyr6LDifmis5Iluc2QpmbNyIw6Eo2er3YxFQF+DVLEobxbwVKHkjoUPaY2/WQG7sv1LFnI
yUQ2eFq4cq4j8hIgTvbS7IiKTjaJ0EVnbnwOrNien37nRLnwdmJwFphmkttZ01xiNGrUIT1YINPt
07Zhh66MpFqNEHs+OAXIfAwauIBddMXnavMd7vjuoP1wvCdCk90k3if4R6gvtOHC3+/voWzggR9p
h7h072lqrCwGNvU1u6KcIIZXjeuAu90oBhnuB1jYHsScODdN/rV58bGLZcOyfY6VfKk5QmgT1I6H
gqhn/lBahRCxheRKWhHSOup5eYdPxUpebr2MJmmsT/G0jWO6PZjmitxP4WUPzM+oHplVQpjl1byJ
qMs4eNUJsF641JolsW0zg2IobHI0ykpjFgwwsgn4r9S562RY28vzcIsix/LJkAA7xJaL++Q1BSJp
vp8kIatYfH/MxmXxj5/9TZALWNVA2S3JAhG0NwEk1B+Jm3J4vQpxa1yGAlfvwpdFuIKc0mO+0ya/
kqpeNHvYdSh7eNdiRG5bvoIQOmquhvipPJJhWhDMxva1rHLKDN9z406Pcq5cMfURwYN0y9mxacdK
pAcM5FLqe0+LkUD2maID9Gs4Qd3tJz7aFI0HUjcoKj52M5PI69sv9hoXp+jqeUZDOY2nR349lHns
tVwB2IHL4FwlFa1KmLl13v6pbkyz25EqXGEl2i0Mx52EPfS/r7JG8Tt9n5CTfPgBsUmR2FHodFNW
NJKfPA5+7wJfUZkbQ4zE1VaOw6ZJ3M5VwDH4CSciEr+yKKljGN5oa/rRg/ZCxUHerojLptiWbX37
4O6p9TNUaDPPcEtewdRtMe0iBguJ3c8zh/+KZoHIUL4Km0GnpgJeeiSM86UWMAHGoGv/ytFmspjh
E8aUrZoK5h5GoXFfexc2LouEdCTon5MFJUa9KUJXOEaKXlO5bG36pPB8sTg27kUPnY0VhbPu/HUB
IanMB+wj0157DTRwxNoUaEUgzAv15OmAt10tx1Qnpa/9NsyzliBW+pRVUI+BVOX/NUIk7H4C8OZp
zcP/xDrMUA6VeFd1iBw07TJ+qzaSe9Z/DH3b6/RrZPSv11tTYGRo6B6JxlQuaFMwv+UZhUFfpR0k
Zm8YnrP24BzOpeTYhEOa+1dgm0PWRQVB6/UD0giGG6awfU3WoECht9IhLhBXR/mjIjg/iIClowDz
x4wZsAEDxx7X6rU7PmEtD/2AE1zjIbDVeEVRs/JvBuXCJc7/hGhrQklLpq7tSUed6PWPNwD7d0f3
P9A4w2b3y8oQuGNwLoXaW+njPyji0Qah0Vw5gd8lzeDBN5bmIFbIXL//tyMenLzOmOS4rwbupRCW
fHUS1RilhHk8mBNnFP5vEWDBB32i0YuYl3WYDS/mUKV/K+7VhwbkgbjaI25657NBvsPqfL7xs0pV
HziZNjxt1F/I5JSW0IXtH6pDNAVK+JhO2Cfd+mmJ/F5j6iGT2GhUivQ3JTgk4Cc35S4jb4/gmssn
nlFoFB90V63GO9tXiopYchi9ctuTdXlu9nFzJyaz5RCcLJJw9r5xaB7EXva1ZDtLPQxF06yO1Aod
5uxfBb67gURMwVt0++sRrKuFelgRYnGo3lPZ6zU+Xte3OmhEOuJdTFXDxXpzcrfdU+u8lujxXX/T
DhwiWqPE0dBbYFCWehQRV9N+wapuprb4N7yrSKm7FOEX0Q+e65xmaV8CpaZdaC6+yiDOf6q6JE7A
0gnTTPgrJLpvna4tkLdwNulwvxiZ7GcliFvulq4sR0Kz1N/9QdQaODda4RjEbp5eMU2pBEF1blps
NAzcpXRruMvGlyY22eRuAQPmEAbs1GkiPTbBi8uZoZINH8VBEaApbDbGdUBUfYlmubxN1kjOWb2N
Vd0i7IPSm6HWnq0Yms9ML96N3Th1ppqMYaYM38EJ4qBvEnyOPll20GQRcghbGjiQxs/WFrx1JbqG
2DcGabXiZp+Iiyh9AUycXN39S69VuJs20ajdltbxRJdfizepvv5ZWuIMYBlqOACEUvHGPgVs5Km7
2DhKMwK0XPbwXYAUI1OhRECS7TK81xjJW2jWiG1RpAx/erExlq+wlSt39dA9PHdexoYFbNcfDSrl
DEFb7UivG+v9mSL5csYHKR1UCJ9r/Sus4w6DucSdKsAMhjpacNZjVAWg+m5np/DVvSVEei3J9Fq0
XscfoDiDj8TX+GpHkawp6afSQQPoYC4Q3UjbU30ck17FAJ3KYLMEg9tqFrl4zm/DrCa3yybSetDe
zRj/lIr3TNWEnbH2O9XPEiVvnn07eLuh5iqZGTJbxO8sObqyj3UQHc4ZTtbyNlmOa3X+QoJ+e+/D
UMzM+HxHNMoxW6myJB3X51xe2jtQN3a/rHHxAWei+H/YVgVdkwfSnNZqGUFuQN0n9nK1yas4eQDu
KHJ/bYHqt0dgaOrRlC+y3PLEGsTQB5XFvRmUSGaW/gE1SgM+7NvT5dP7a8l2wAkCmqL4V344T9IZ
CxdP77aZI2uChOiV6/VrN7BDdIXHQsXp0U0R+T70toDeRPSm55x0DVHXueAAM5QhH5I5gWtiif7L
PG30yArmLZF7In2fkymF67jhXY15+I17sK6PAJ4Y9wYYbiQF+GBFbEQV9ygHThe/eH6ye7VoDsJ9
jpG0XDXm9XEeHZLwWBEZzkLeL5fUK6wr1Kff8RK3argvodQeExVM1pujbKbEPPWPS4zMniK8bWuz
vWATvxvr+ROH5WUTc3HXWxyUccT6SB+ISct9RkzM6sTLAQ4Di6QeDJuxVPNhRNQkN6lxEE1MT8Ie
WFMB++3NiD5YkuB+v0WOT3/5jBlpWgpNElr0dasTofyRlXxs8vL7ixN3FHtAoGwTZScsXY9MtTrS
0cKSj7oefawauB5Ek0DzPUBX0JmvtxWSocbr00uq+WczgAOblhRyOTwvHwPi/0HAR3Jxf4xv3xAw
UK+Hflnj1MJdLfCLfT77/NyH/XfwsiUQVieoi9oX2/uRCl27jx9S/asX3bVdlmkYBi8sQ8FP73/O
lN7YNta4IbkEzQBwoTPkdYf6yeRl5ZOQxcAHwNjehVPvXlog8YRQW63A5RSXNQOpRDBn+jTtbXcv
DyZXD4NfFcZv5g4p4RwUHsBXXAFDblUPF0xsXCdtyHNBhBJByqQC3IbTUx10kr15mGmmfXy3/eY4
8bR0oy1GchsVQu0DSa2A1yPxZ8XsFczTcEB3C4vLDI8ZoxeEL7sLRUbUVVhiDmqkmTjy7bnblCZg
sy+yLDUXxgyE/fwwbky6HPzG+Nm1G1zfkbDKfAbeSXLsaq3frNWFgjg7tcvGyFJFqbzys2a9HShB
hLfAtwGkr0AN0nE69KmPIRItW3YoSKyWfc7yx3T72hP9lQ9ZUS5lGpzlnAPRf9/kzBR4pyk/fr9J
N1xkTiy87N1fkibKqUbGEcU55FkRpWhLyPkM+PL6JeyfFFkggTvNhnaQMfQLq8HExZVlPeeD5FKk
nvuCKp+FL9X/4ZA6ji8yf6ufzknoIzMoKzBKJN+Vzjqjjg68RaB2Acacwj9REsNfPHYAQDjum/ZI
PedQ7zXunQy83N/Zrz5j1zF0ivrVk27qioJJeXecNFwulwdfE/V3xl8/ryFImTEaVMuHdz6Y2/94
j7/3l9BTKkvKhfkL4pKnACDUf8Q37JKnZgVCTRrHKV9zn5NfdyGj2JpjWf996WVD3Mpdw0S03Y5V
ooZEbPOpcp5c9ugdXxmnNSnsFqYd3Efk0Lc7juHsYvhTmE1KjXvYeIWs03WnmMQcFyL/3p9y76//
lN8s6KSGxGxjBek0+54NZzMJpY77LOM/ctxMBjN6Gg21TFkfj6cFFMB9eg4Ir6xTHPjmSbFLAAFC
Q6OiBhFu/+8t+nU0R5Xw+2Bb1zxoFg9n+Ffx2t8pe41y2RChLHGTj7zsYajXx6kZA7lC2cjpVe55
OvGr9895mZNNOo68EiD/4fVUlT/3Z1Q0o3Lf0gktgCwE4NNBf1ekNHV7i+ZNo+oRFK103XKa3sQb
twwaIzXiScA2/uf+g/g+HLpXyzcA+Ev/4emjCLwA2nXz2z/+r4C5ZUotjvwJMIRzSZT1rGrtCZOz
uMUSYP6EZu98EcIOFiznppE9oLVY8s3aQfpNdfraYunVXi2g5aZm4Y/RU2GvnvN5fh2PQXOiBOrp
2rhpIfw7znOHQhvmeU2SawQ26LEVu4jHhWDoY8fEYCyfOSC0m9aDRrzL1bdHBzRl4kYVnY0aTD5D
zUERRsV61Jf/2aPjDP2anJGuJziQQWGiEid+ohblC+JzBCZaT+3yntG1Yvs6nKqpraZk+racNnJI
ztaMzmACSoqPLtj6Z74fBFLv6laAMYx3G9ds97DqMGiH5RpKvvm/q2Il6wYCqVtYTd/J9UpAlQ+H
Ll9PzcwuxfYfVyu0b8xhJxubYdKA+r7vPKVA6qd39pF2ucV2ZRR+mz3DQCzfEmvz+FbbaPozzZWj
Hl5WoFkB7JJ2VJQHcJbdeRVzuZXAZhOgOtvO+m6hFX1sz4CEBEaJrfMmVSs45ke3TF0/lAK7L1pn
zRd9QBizA0f4PfxDBOrCreY6Kne3g6fBQ3agDULFnVuYqMA4a+2E+MeyG42K9G86bhdyN4qYpVXE
LhZYW7D8ote75rhRW1IJnSeSl0bv+2JeAwjvLoewonz6WMuN7qAFlAQXcnIkBaIxf1ffTEUiuXHT
4czpTAehTmhb4vaeWjL1/7hfxnm1h3eH8kNgFOQGo5Njd0L6MMGpdkAUTmXyMSCtSyDuIPVy0KUz
L/XxAP/XYQ0ZCZ818i9WiLrApfSWP9JGu3991FfOJkAzaHFRKjqFNqlTV6X0k8jgmHRe4sguixsT
qYZ+1GT6L/OMIKMRbTvSwdBdIBLG3FxBLUKjJ4fgxaAcpxSQpr3VxI+SS1vLvuGJ9hkQKJJx2Sz9
6VpNCX+efEslHvFI+fL/7OG3KXj22F0xmG2itZmt32VaKr0xqDP1zQs6loUetrydZJ5vaidhr7GU
mxBNWSklzefH2d4uGiJdZfk6vRKxVWSTv0+6wSElY6mUVxSrLagFf4bcnBJA7VvHXr3RhzsrJooN
qv+fRskcXmZJlJtDngGs6N4+Par81m0c5kX70JV5Rc1V7LWuVp+L78s8IGO0xD+g9WBm2HY3Gaov
gt2RfxYdbX7xnSOIgbarRbl7oOxEM3ct7DA7+nG5Fl5emFJPxkV6ujFlulVPTqh5I2iQyVmfUjS4
Dln6xjSpQigwVu3aPWMHu6Dw0u994k42IOc/vwuA4WbiPoyvFTy9j/x7K8/LgTMGT+UP5bA25Yk3
3TsCHvzdWwskVfzILHViW8abBl0Vyag+kpUmUkLyGD0FJQKpF6X7E8VZnwjTvYkNa0ucU4ky5AkP
0ZVJ2ZOTFSJFskLZpkj884TnW0nqPySuT6aHlQfhgFbEKWfOQzfk2GxIFeErpvXbOUYqgkXvhlH3
7gr+NhX3NIzxjSHDgZyBoNTC5z3ZM1j0wwvc9MM0du+zQXICvAT3cDHj8AF8eEYGRBJjp+orcmZJ
BvV/6i5Zjlzh02ECyjcJFIIFjHeeWIQnmg42IxmFD5gqTejhtzqOBLfTkdNe23Jxsxo/QXvT0GnF
lqEmOKF/+1jBQssYEEVl4TWW1ZuIuGBGfltUr9gXS7B/TU84AO+OBiQXvDze5gkpU52o1a9wwS3D
Pvr3i3dkTf13Cj9J8EwcWjSR3hgioFkmN773LrIyrZwHjiKWXXzCSkLtUumBDN36Jzmt7CxkrAFq
ApmYBhcQHg///YcBuRuml4SKo5OVPsAT4cn/EIrENtjEzZFjTsXCEWvbIFo9gjZbbOegy65ven/T
3eL/bykSQTlEs79ESk4DZf3r1rRs/n2uKsCD/UnwT+cdPjFEtbx8a/2F9hrIv2WbBoMu+0BFclDA
wxsUUi7IOoH+/7hL95bi/Bp4McToDuUjVU729LZUuemQN+ltAc0pXsT3eewyL5kPndsNwKVeLNNX
R3dbJQ9vRAsvnssK2BxOU2Y8GMYuT0b6J5Gaw3EhsQ1clGopc0ef2KodPNKjF2ooPtWsDBpx1nfC
0QNfecdDBC7rmO7R5a1vUGsNqcfQf2TtMinx2XsGwZk8F3XJgkcMtAsv0gxfkgyvHuTvc+yAflZ1
XI3AnwoH5zlouH9T6xP2UWhdlMHAkz+sEV6MtWqO8Zmaztc8ZuKbiiwbZkiV6xyEi/fLsX9Dfk8d
Nm6rZOh/yjLxAI5VRA71sI8PSXZH1Kv62sM4f+jM5bdGU9PlmcXg8hX7c4fqLk1jFRa9sOFkjUFw
/BMbTrIexAzy3BtrvJ2ACtqZfVAQytHbufCx5Vu79t2M8JYEV1dPsJtDm861Gzck8GVIqEu2zNdn
UtyNe7ZQEUjcdV8J/rlMZ5nM9QROH/3RdnsCqJH/8x5AQPsOflF6WnblCdYvS838MAuJ0pqKMGgQ
01Gz9CbCYCihjsdBlhBdGXaYiAUkZw2vTTYsJA06njQDI5U4yRqn0KNgrLZ4P6DE5KAcreQlL6Kr
EHbLY1SXCW1AZ9pO8dQdHCLoS6DXkT6z2g19i8qQPpjbwDN7s5mNKVcj4iHVVPDIORMifbFR+ZhA
GQp2rsfLBomXg95mTpQISjrZhC7q4fC/zMVYZMKfoGehYE+ytk26uzx7wEW3Bh7M3WrBf5US//sI
EhcdHx47BKXHboeIy1RkMtfevftD59QpUuwQXS2L83Edy8caHW1Ij0w76l/XHrsDEt87ANuHl4z7
S1XLEWP+ZH1Hxe7DHO/DE5F2gYeBiQsIbGmLl67FX37jNqhN0NWJqPf8f/Pnx1A4VrUKirUrhn/o
DmXze3zpodrrF+TtzBNLLNtu6vKwn+MeZAa0qx7dI/06MMhNxyPVWSFVty1TkLP9opxJFOR0192e
3zSqET5hAz8qKSwLnwNMCobBkg6ynjAE2KIDZ3x6PlLhcDVvrg34n6PZEWpUiA5ZkLTEPc6BIhtA
nRt1SvcRbSkT5uUzDGNKUHrHo2gEYCosw+vEyJ90GkSVpYObpVciQUKnnMzckBJypyE39Xmj8ICn
k3h3cadr53Mah3bG/x76oXks6mxV7KVq+lJZw2rqa5B28mFdXa46A7DFRGlc9pEgL2ABHPhCtTYy
6JKaSG7Z/Jhz44jvNidvhA/fHoHV8oyaCC67IW242oWdQulhzcGDrKmllEG/ijN7wn0qXNZf1Vsv
ZNDBJ6/OllcnQmvSrZAQG0O2PaFk+h1bjXyPcM1teEYi/NKzd4PcDFGGHULO6yLl/7H3q4oNBmWa
a7iYS6L5SApa6rpxIr/tTANNtiQ84qPJqIgFBOdLz/LhVpT4GvRXeoltYaLNGIKofxQ7Pk8j5MVQ
4IuYYJCBOncTZeuooqCslpU4LmWZoMr9bi1qvmjOp4erZQOCPptxncaxoJ1rITco5sYMUnhmKEkg
E/K7ms/E6YZM/NkMtI80r/xzX2JEt8Pqn+aEdkkfy9HsCd194sueXcB8Qj6aIyKchOS9XBhnQZqZ
APUASQfTr1hO9Yt4dS1r8zbpU2E10FdFU5L6QGeYX+asJ4dFmYqJLz9a+RJpoqOLboDrPM7eguRP
xq/Cr+SfsZ1rXFm/E0G1wFM2w6vrsD3h4+zjuJmcsNsUeasegzIRK0eYLTdRDKxNcgx68BNQHkq2
8OdSULfUxZ1GQlrFtneBqAx0XTLgrsjD3u/bkTg+heyZNSe+lgCX36BOADE8Wo3tEuQfmH3bt9kh
zykec/Duy6QIjzaPLT1JrryntJf1yEugMobbsVOh+83fvuiU4q+guasz/y1XdPY/3xmlDVQWZFEI
gpSuybfmE67J8P2axmhUv2Ns/ItQQ62Tz4kO7uGvwzN9sWyhSVDpLyS+vVWgkcY6MbfTJmg8d527
owvtOLq+TwvfsH4ryH03fmc8PX1tcRQs5Xn3fQv2F5K+VjBvMH2rEg6XUQdEgqhjeWKQldoVBLOt
Ta08Mn+lwcmMvxjIjZTO41px78i46yJfQY4J9Xkrbq14BEyXuH9c9xDslJ9jgpEafITWyl19VFEM
IMXeEzels9z+9xgoYBK0CpwMYCI2RYt6K+pP9pU3FcFI8E2G4v1xrm+QqE9abBY5RHMCqLYT46ND
tTdypnl0kP8aAhUTRXNz+Fy+7j9y0rG85dCCe1Vv2/ihhx9fly4hKD24FAL0VSaicvzTo5ugFKO8
Q6e3aynVvBZKiuTKTznKCuftR/Xzw8Wfm896NjBhOYTk88Lq2hKm1BQqiBl4QgvbWyTmHol/R68m
5AfV7LSr/3E26IM6tHlaealWdI62pkCS/uh71j8b9r7KY6prqNuJkPTa+i5XfbzOu0NZWkLtZCry
Epf881hxzPubJSWorXsS4Xf2QDUBIrSBi2qqhajcAe7wt8OVzXZJnkIu0ke/veb/OSR2JEeXofBv
U7VeZSB7LVEWSefP1B+VrRN4gQePj3sbSnCYRHvFwaZ+9U5CyzKXwJibMITeTJ/7XQvUFJD7ia3+
R1V2TeK1zk5BOIosPBTtUTLPCIv3Op3AEFdmKxTqC2h3i5PlM6+W/irDneyS2WMPvTNhoJN5XEjc
RBS0AWuzYuWvR490rPa6Vk+pb1aRNEu9ezoPdHco3AgAyxAZAJHat2rXmF2io4XsWfnk73caA2wy
NZP+F9tOjYCAWlHBUk/9ag2kALBAY/LpreZM9tGwgBeHIXrp1tLvqPW9RqaOAV3aOdzaJv7fCyaj
J2LzCOysP2xR330Zox2B6m4+yTob5pIbzR1L+T4IUQZH1kjwPVqs21WBbLQmLxx61zSZJA2cPfiy
Bg4PJG1JWscfPRSHzQYIqxuOeAHPo/AqI6V+XnsJ7byVgvMNXXrYodnji57jgFG2An4gakeWk3yn
/FHOBDsdAOyMWcGig4q17o9GpSi12nATHa+gJn2CElmlbn9MNKsEs/V312vxGoE8AvNwkxwaZX5s
eJ2DA/h1J4b47YOOkT8Pz8McRVbXMPWBKjhNdZo9zRtJjo7vTWB+DxsezgEHmi9zxTEBlNQvu1cx
zEqIDmxeCvxbLoq9Boe7OXZXMA71jhix2X9fEjD9Hj1DcocioL1meNUyFpE2AFJa+sreoafvhwVu
MTDQCum7kMSwJeBT1ix5qvYYWfOJNMpwDpEY+fzrqx4hHJ51HlM4nAfwGjQTpLMraEd6xToiBYRn
pPchLXzubhz9gtsmEcvxVxoO0+cTQTYQTIxzmrSW1Rwg7JL3SRxFoWylf5CCSFT97JxJj9bkWoNy
ipUq6jMXwR5RZ/AAQNcOpJyqRrzC6/P1VXm5vZIL2/sLkf/elOuSQt41uyJ9ZFTbGb00i6LLRaCp
l72UbqfQ0VJM4HFDBQYrsgSCLjInbK5tjNPKhZWohm8U7x1xW6tk1f7UBptpduhDvrJjs8zwFwWH
9j3+d3p4KFziD+YWo/ee/+eVpC3cKl9uNOoyX2cFt5DNtQ0czdQesBhXfClvnpCzUiid0/lMHiha
5FT/d7itFpjphBpjgxpk06PEJqAMHAb85RQmgjMJhzlDNuwgH4lkMmbnSPwdDC5mPm7/ouTsi57i
xH6TjXmJD9veNM3h4wBqiEmd/LQdQ8Tuje6p+aq/AXJaMnIqrsaK1AuikMXksyj8U+gOffLodsRu
Q3/SV0wxoN3ZgnvU3uXIXntHKoXgtN2wqBtZulApFi7AdgYq5vwLx0fwSD2HmTAwd9E4WA8S3f0T
BY8SrUImfO+PqK3ivhxkiEru36RmGX3fxApy0JbBaURLPQR9sw2D0RV5AVwysI/qJRbdCiQJvfpz
5fEXA4vXfSN7ny9OGdg/DHUt+IR3GcAmhZ8zkEzyuCG26pI6e093RXSguWj5ICrJBWomW3p0KPgx
xrehaFWl7hn++Ya1XKSOKqZwboWerP7BBEhKvKCwzrrT3upgDvk6CGOLijSfx1cXuqUfsoV9aWXO
jIr+LROcyFuRXaRdiEhGi3acHofT+gkeM5is/7q648+f35KiaduAYTaEHEUS7RTobl0JdYAZg+VR
xIittbV3yZYBxPVB4t8LRZHL/lNrGoIa2c0TjA0EGu/ZOH2GQCycfm9h9yw8ftj1n/tkGl3IIJPN
tDeg1ODJtzF9/+gUtfjcsckVdHYx0BRXg2/+g9S1tzeUd1lxX+UB+YwU797uQzhWywFh8RbgU3HJ
lCvMwqxHIZub8mcIRp8TQPVjfEuoKJFgy0KQxYt3uAl+K3hYvf2UJLH0eH0DZ6q/oOoMU/n6Ky+w
JXWIf9A05WrPG0mYWm9AWn9au+OE4qYM4upR45GFTo5rJZVmac+XczKFWZ67nbMB/DZ9zK7K4RVl
SjKr94HuZ3gf8NC1bVZlqTonombuPVZ4plOKMn5nVJji61UICGbm8i30HacOLY+VknX8VsR2iaHT
vdOBm/U9SEPa5BD6flFr+PYHNw4WCZiJTg1/x/5ULpCB40aUOLqj11vU05c5ekmpvb1GPJ1D0QwK
Ob5IViXtwp62u3cZwgHLNM/FhJmaJlTKFq6xrDmjvoZKN48/eXHt9ArXrzQTdmDo9kQ+mQf9j1oE
tFbq5n7jxSd2u+YzNwCMTMlLxSrBA+DsKY2uomOFjm0zn89yyr02GwX/b4xgKfx1aiQvsMRq4XDx
BIJtG/dK1QWIN/lytwwpbusLJ7ff3UdChNRF4DLkeAXvSjXx1FsvkQNpZXV8CrTlTLq8uTALYnZD
dAq+4/g0fSrglauUkqcPUcd8h0mJhKCC1QZPpcGxGRhOdBC4un4uKSBLCjIUx1+cWoULdkSi+FJu
/UBMrsAN5gLF1dWPReySvxuANiwnu7Eqi+ZPtwD03P124HQn8r2LoRvZe5y00XN/xgJ5mPN8nri1
kvyJEUUChbhqdO9kT1KsQ13XfNAoNPlxjBF1PkotbnACR+hI+BhVgiuggS5na8NSImmDfY4QKrb0
W4YqpebUE0b3LRDPhqRy6bYtqIE5YO5qgobc8OjzzFzbC1tHzzv/KMMRIWfBLnf0ftHUQhQHUXAP
F/XIEc48tV0MZKJXCJOy1YOodaYX0pyaQKjVjQHgD1XqLtztxEsq8w70aCi3dzrRoytUsx9/yUoO
/gxnM+ahlJDnu7vWpZgeEa0k7XVqaZrudDjyL+MlhkdkoJMCpSI/FPBkate12uQgp/xxxGfLDqDF
HC3rnVcajaMma3fAhoQ33iUrOE3QfOHPWLMVnn3eGF3TsvTrPJNGOHGeSbhsaqNcTWLmQfpUozI5
0gO9OFMJr2G5zVBDGxO8RSxdT/BJ3fbXE6lkvwuB8AR0y3QRKUiq09TRQNuHql7JGZ+v7IVTBiwX
WU0qXMGo1P00JmpRV/ZMk/dsDzMvotukiPKvtia+iv5LMTNzRDRlGtbVAJGAEiG94pPjh/w4u/zz
lvGKPzce5u+a3bHTbcefO+q2K+kpT1EH/Gpf/xxDLjMN76S8EzOwkvTvYMcNs3qUpJeGeQHOO7lA
+ocZxw8vIwSBE+n8Zz4HTb/vyjrhPqHyODIIwStqnTQ6PBFZe+nZE0n3Us0924yTNl4ouNonwQei
KZrmxd6SCR1WYswXYRqvErbGpAU5I7pvWiZQeNed5sYtbteLrNpvnAc8myU0IT+JyA8rbNwny20H
ymJWGsznEX6OOFwastnn5FQG4a0GYAuYgJHL/7pPuxbNBOIVh8zF+Dk5dOd1BdtK1Qm58viYmRDB
nT59v/DbVkTD+HbYwPflhvBeZ8NN3oPPDDemIg/N/DwpzZwLUCzV1GcvxJRSyZ0YjlcUDDPLCkBx
nMzMp7nNtQzWIsYXMnMslj/WkGQ1i/4bcWi2VnhHwW7qGMPztkwkZ92vIIc1RiV141cHFFZedQ2e
kn69iOkqLXSg79FTOtJBobN3rav/V/oH0IU+s9CTXzFiMhI5m6Liyj6tU7tuFrriHHMGMN2YE4Q2
K+n1L/tBRGp8PFnJCgt0C8GYrogHxe3Pwo/VV40jcKtdeCwSkF0LSoeoNFCkOgCVZitECaOQFllJ
6nVjETvzRkvpsmH3IqZiV+fweCQoejCwRH+DuIWyYL3e55SOGjudJX8Dh9CbNV+TA37lnrT6+bp4
mlazUfMbmUJSsJns5R3se3YajOu3NBil9x/LfKuCsjdsftuOKxWso9CAWDWJz6k0aqlorRlx4tlz
sIbl+as2WgLgh1oDiqPAYtB4NZGWbomtB/ej5VRwllwgW1blohiP6eJ5tJUtliECAt1aMIxs4myb
+ymssPllowX4jX5UTJV6eMQ4kNZSHe65n8xQP6A/iBptFa0Zi7LqqzQWu9doqNMeJPSeQPVjt/Jw
flmid7WAoFIH5Kh5gjau7YuP3gD2p4N64kKc9xZf88QlXHB2g4j0R7u3uC2jdsW3/EAnpgOngpoV
2dt5ak97xHxj6vOVYcRSwCjRxcNUj/iikD+7kHGh3hfOFiE09YJt+xqzsSkqmBwIFe8tU+JiFYZ1
WKzwZZTZ7P+jHRZX5US5DqMPIW7FGD6oYejP8kLz+WEq36Tussf/7MFDAmtgJc2RfNjqhVfPHUZ8
nH6UHMx+mk3Yrk+qvpEilkyFZnxM4za2CZU0KVX+wNNue8cJ3TZ2Q7uGD+3dLKM8ER1UUfGh7wm8
ze3BPYYbHqIwCtFX/Hwsh7Z7WwFq1br4SXntJ5NHbHVWLqEAd63cxMSLIiUZXSWtXMlylGLAaFNx
6a530N6kitUxat3KLtRBMgJBTrxDHJA47bA8xNbTSBZEaizzuUq7++wwGMofI0BFXdteoLORH+u3
HxJeJKqM38wkOVaYe4XG5bjVaGyzwlLKguJaFs22aoSQD6iREuedeVrINRo/maOr1auyhIt0hxJA
C5aWvj1WEuMS0hIBb//jz4O83rPCzwFDpRZP8IblugFVYEqtPn6MQLHBMbeTRiU7m+msAcMJC75e
SZeOsJA1GrNWI+j08olKUqxb6Y8Bc/jgEXR9yGO367RKv8UqljtgdDfFbQnmpIIc8mdD4U2K1PL6
OHGfAOzQi1vxFUqOjTtv0Xvoweh5nRSYBXZQKj/BTdoswnMmxBritt6VUS6xQUPMFcgyXfSSFnlL
eHD3CXDJaYi1Qru04aFFBd9f1j2jwtSZVJJfpj13ioXTkscPKafjJFcPvmbQrdCnM7O1da/stNgy
p15YcgK2SCXDLgMysr2d6shldb3TY1Prt3ZnPG7/gP6xcjIMhleXvbpAgqejh6U26AQ0gJenT4se
DmTAVAk376NPn1Viy1jzwiLipUOYeFmTJEXaZbkI7pU+Edojr1/b6Lrkw+F9ciJzKpBmrO33A3B7
tsdFILpa1c7cjPM09+N91FKGfoSF/JcrFjUWYir2iR/xsNRiVgvUOuu9FjpnZj9+Hii76s1WsV5z
jowLpBewNnrBroDTlqnkBRzLhXu4wIrLJrCLWSi3NZnB+ihlfP77xEc1oF4B9TZIeuawf3cKGKK3
QGvA+LadO/mH9+0LwDtpdm6/x5vjt2btRrbtHfgk9J226AUNhxnIbnwrbtR6r1lH2iAUDa/HcSre
mBrxv32COGQP9eGMHU43FDesk8+OPfQV577u80RZTsyghooApYHEWRc4+4kFx8b9DvdzhKVv+44N
m1z33xP7SdH2LxNVY6nJqMmmEJfEzmnzCl8U8z/nuUwWgYzCoMdX2yOFsOHZiileX3i7aKvwtISN
uHd6imWRnCDRGfJQjPYOUCLAmtKxRyTPV0q2k0sQAX0uV1yD5DlrWMH7P/X0QbhbZYa5422lZuDV
YBoSx6aLwArW65EicQFn52ex1gCOBEwBhWoLCMJwUyBEW2ElAO09SlM0mkKcTG1E/MVJS+b1kgnc
k6dwyyjKBxjiORsKVmbjc/05+yJz8/zISYTxDjwgC9yKA1J7TMANFdbo89FJDvdI/lzL37237u+A
VXiui5aML7daWXU2LaCaWKq3d5+yujBYd8NKhqnhkz9QivrV74TyO8cgH0R6rg45otNv9dLmubNg
LSBA4s83LSEmkDjW/RMQ1s/RxCjnzJSFnfmyvOVbXixXeet/xevzRYV1fRrQTP+tOg33YCrr9I/9
MUGIeAkJOlnmdTKHexxrfTVjoJnEEI/Tb1zX8hgYaPO6utWG7WheG1vfc2mVSvLorXin8TrbU/32
umbo4enV4XPWx96sErkFCfJhSfhL0fNQfLyduOxZD4Q8fx1Pdxyyz/DZDHWF5kCcIWF3D39Cr8GR
JUBq75TajHH66zvcCLPtVvoaw8a0JVBcp9ZOanYpPAUsvXn4arshLszGJEbl0PEEkvcUWzn/Kw/n
hRq4bSi+vR8173eGfbk8GRgh3Go1sXfyR8LD/CuGwqjxPVK6Vsgsof5J2YRmHJ586AnPm/X5WAgl
Or+gnOwPNGwzaQ4XVX93eg3weIAikqL9VnX0xaiHTOtm1LTJEF88YN/82ati6PyOWHrSHdcnYdXq
k+CF2AKDOsUIZLjlwSWyankPLJwmF9Kh//35elfGpGu+h3ZJocQ4X0+3H3v2XqFN+tIgAf3mYeh7
TT+9YMgYKnPx0drJEhz9WmYqjWUbayWfHxedAtVoNI55yJFAQIi3o3gWM0qDEU7aGyOiuB3vZTi/
c3S0SF+5Y0m/f8AlEV8paRdf7mGKZtEIHsVtvdKo+yR4ozR5+RmLuTqNF5cdnebbvT18MGkgO9NS
I81aUAUWtGqoArJBNm5FSFaGLYd1Jt5UqSum8wVvzRNsg/1rlYt9BYHTktA91bXzXGtWZOgwmoca
h0DXXdgfI97V2SZhyYxLGVCrjrI312tPGHYbhj9l9Q35r5hrlX4dvVtvgj44rDLy93T1PJAqaHeA
BSN21wFiRgDVR2awVfbyBkRjpIhE63Psb+GZaxvAqnk7jIsar8XqXV6EC+KPUlP+gLgthekATJkp
SV6dIB+/FDKCWBu+Qdzxiz5HUrEupt/wuzoyTyDwCSlS+SZiMKrN1iUaqqcBUun2wd3J+AGmRVi2
TAxpwEt1md219hHjcy6lm8fy5hAgTATuveaY9uLrdXb+5uAso1foUFtk7ZZQWEHVdXlYH0Js7RCd
qc+fc4wbrmsUXIOaBdY5PI3OfMXp15mpeXMYCwPZYwocOCQjqRuUTI6qMr0NwAVt0CwOA31l5VAg
Qc3cLuV0XrQnJ2LR39+HcbGDo9wBBHzEQyuLbblUWwN0Iava3gqz7eclrdaIf5FTlPVuNbu/K4nQ
bbOc7Q/RCeN7hmPKrp1Bfn1ZsF0eHmr6076KbwsaKpP9sF5Zze6YPN50euYnGdqLrxfnCHW/Xl+k
Snq0XzjI2g0qZQIKqAef2WZqX12ApKxJv3ESsuFUKB8FHR5ddB7vVRtdKomAJFbtu/OEkHILxLft
/APGV65hWATVowQrCNbBODsTchj5M03yunokaFcC78ycXHUB8xWcazVNNzmXuyqmOGwWL7QW6oFA
/+2sUYfZTZ6d+kUubSh/5iVIuX0PriZIXnvVMwyWeyyL8Vwrzgx6RnQt/62HlMgYLBs6H8BbQyBb
6gBg6ywwtJ4TR6SovaYHLk5HoNeH2ozAgIgridNnWSju1YHxa7L5tonFog3g8pMaEpBnrsYdAvX6
eGDO2fmmKxy+L7N018Bl446zfux/rIBN9o7uuxezPmedQMxHGtr0aqzMo510LOzwVbvx/TjUhWms
sniOEIrSUL40hLUuaMvJQb7fUFsttjOA1dmm8d7dThbiMscTLj5lC+HSbMkQvx8KSlW8ncFFQ3yL
RFHt+1aX2oQ6OPfahlMkUj5DnEXUzpKTDyeVdJkKpTKb2508pHTU81MVGMwAZ1NKLdqswzj/F97U
HZxoTPWcxKrgqOPrcw5jfAL5SgMRB2LjUrzpX5W5iIpRtEWpO3DKl0AOFJ/ms4Pp4X0CFRSbZge9
WMt2Ri6fuLu4hr0xBup5tRtg2ZPh0P888Ggc26OayEyWgclBcCFT7HeWi/WAGdYtEDpWRbGBhXE5
Ih6gEblCb8epgVWmwZNi1m/nQQJHo/J61RrvPJWHHZe0bxF33C1cXsO2HFgHP1WX09Dq4UNckeQF
cC3FyO8HCsC7LjVdTNf1hL8/mx2TPDybZH/RypYaDnC2yFGRe0ChE2Ow1n4sHtPt3yxI+GlNLdT6
CoL+YQXtuKz1MNX4tLI/7Lq4dMSsrotZ2xEQHiSWspZjbGkaG/8X5ajvrM/OjMJtPN/aibpn1O62
Uo++0quqzR4LwH7V+ZFFiMVRp56Q7bcsrtpyS5cO5sy62TQ0951NODSKOVngEHmob5wfgNFhlQCu
DHA45EWp5Li+aCO1iqoT54oPMxo83iUHat2LHfWhJaA6S9r+qD4gh1u/2oxVTIEvdLCz9mwqsPju
XUr4RIC+QzQcDqN6hSLLG1OH2mm/X6FyE8NGzHorPKpJWJPRVuwtYpvZ2wiffaOiJ7dw61eXiTbM
HUJ2K6LhwIBH0G28cYk7YCMB6LcEtiGbk4XuEvCAx4Pi/2HcyKIA7fFVhtukYJr8giEgtOMZMbCq
y2bb7C8hMu3PV+vYjzamkMf55M8YkUSY7ciDmtVgiySpHxgSbvts4YJTO+T5R8Vjq+RT+SA3W7+N
FFyDXLFnEFRh5dZoCbofx3nW0fEwgXHJ+WARqReFRtYkXp3PwOdnRV6p8dVpRq3LjpCkQobmqrjf
loh0FiebICs/kJtWlxqVi1bQF7JWiysiNr+RIDgxwzkNoj6i09TDoQPQUCiRvc2DXD4srmgvq/xx
m1e0YciCuvKKn2fRpXcGKbVYCfKb+HoELGdAt3A1jsydMqWBnT4M353GTFMycpyjCkKQWT1FEF5W
+LR5yWfQglyv9HbkdZnbBfdPen68HpGR5XgDfDVZ0GP2McXmEBg3oWyQtMDPi3gm99XbE2ANhYjl
Q/4KeMF4UiR1fkM7WLy2j9oyIohuVC2n0qBYtXbtbEhy+o7oW09eJ0Lsr7r3EgAollLnW1N7Sjds
ZvrRW0T7h5TV1GSD+e3Xw/+8ZJFn/fsqigyUPON8tuAKbFVgdWG7TvqRKw6FKgZg8SEqMQ9wivVh
DWer3IbkOUsYVO2id1XXqZsF88Hw5lnI7fJvQjiEI7Rz/MjFfAUnDSIiFAN93KuhiEhdjHBHTB4a
ANLGNR0TFNjccjZmTzwA5ns43wy2ysjLMBWqumKpxIbjNQSqrOG9j8E5rfyqF6kLVwLZfiIAU1Qt
CfODhnG9He9kqLkn/nET4cuw63GUAji15gVwPYdvsh7YH7IqgQyv29ZClvYwaKfMgAY1y2pJ0uaI
XWc6tVt5VCVR6Knk77kOoJXSsQMJuv59TAooX2i4T7Ha8TZg8QXYKUf4pG0Dhkh9/uDwvwVfd1fq
jCZUXny21iearGQ4IxxIVdv9IApL6KRRGSRiaSKrq48DINLj/f/+JAUQCqyRNTK2TOrWaqYohwn1
5Mcw9c/2s0PyHFmDsKOFpN2dAQEVFHZo2mmS7CDdyyt9AlHN7Y9HbGSE9qRzI73AGV6orfE5olZ6
PYDhybTthIFJJ4S2TAa+cBgNo4hToGX6NeOIslbpwk6oSsa/ETFea1pxWV61mfQkTLiDwo2IcWqV
52zVoXpWEcJFpE3x1kgTcRYB1yE3xUV5AIJfH/E9A44TqYRbu/UkXsKyxMsvyXZ6Wd+EcixDH+O5
UDnM7Mfcl+vijazG7ioY4bojZij3LiWkOWOjiJ21zikCqCQlmaGfxS7AyXV8dqQelskTidqE7wKg
hs0uNyy43vWW3lx6uII/SP0Mrcch4yk0VopnIzhUY1Ua6HmNlkIGD4jGa/7CgrjzIYgGfp5P7aJ/
aL/+CjRPn4YOBZ1uSbHILnht11O/nT6pkRkDor1s+nhvY0AwerX6at4Af/QHa1cqumY8hNBpHG6l
WGesbEInbO0fGHqTzdFvSQPMor2pNvnY9GIJ+/xk/IDFsIxCaSdzjyT/UtESwZneyxBL9Mwf6Y6p
3zF0Ww2gOipxGT0Qh4d+baRCY05iDTpb44ZOI8cI4GdHGXxqMxcg528ZEwrD+qwPvcyWgZAJMHeW
eIlgAZE83IUw6KB/dwB63sS6SzAiRg7iWA4atDLlYpmcvCdcOsYT5C8Scgm9OQe91hGLkBYx90Dt
11h4e8Ovj3bDszoCJXFxdVojPOWszLwoj9sLMDCDr+4NF316NHGvsZEY270pSjhTQldLMKtyuzR+
QjMFDvum3wCqVM8wLRXbqrW54roPKP2ZohliqyenPmLi08dVKpfAe9y2pAXz0gB3a7ijSlIN1MYK
z4cX20nc3jJK+lHUvE3RIczWGVSbbLW5YgsFBgIT1ebNmBnDHP81cHkan3AVMm9ZRscQ/oiETtL5
PUD97TZ10n/Wj5GCe0FNTBXvUNgHwxsh9FBM9ncx9Ckr4Ti15DIYfvoOdK8P6jn/W3T2zT2s1xE3
0mmHbdEb2ejdOAVc9lHBAsiqtRQmG1ivJY6/7ryrkK9fHWwr50Zv3aejdCV96xBIfPN5g6wfUbZp
prdjYC35NZT/QG1fk+eLtgTurNKW1PmSkWl3d+JBbs3q+Nc7tSTsg80BsFB7yBg8/jfqldJYciON
zKSDxQZKKbaRye2LJk8CNclW5aLwQl7Dh5kykoXJWx7Yu6xU22dxvTXFw/6MXxjsFsZXsuA4bU+P
cztno8qP3yAjyajALtacrhbNvuHAPNNWxpPYNEwgmuOGzOI++T8cE3u+t2Q+QihalfYtS3UD9ijc
VQZeoa+gQEVjVXTKHUbIuSWLfmsK4ASrYJc4n7nMIyR8PKACw/aqzCu3cowUOvEYriqhPZMKWKXW
hQn95ZOnBAa7RfX7bUHrmbcj5YKz6fxCIN8cXgUDqZvCdM4vWua6G/EqjiBCRahKGv5Pvzje+qN7
37lt+fNvIsO8VI/rfJZaK6374LiruPlF4eKE8mmSNm/e/O2Qcj7HJIgPuis1rYkHgV9UCsuWxSUe
dNjs3V1sGTIpgRvJvrb8xURpln+ULkOMp2CPIvrFiuvlXFTHG+nlsPdjyJlnDMihoHfWRbfZfIXD
V5/bbzQMtPwFWrFMnC/mMRUZ5RnHfSNusS0mEGDFmsiN6424toqdNfrwTxcskS793quOdQKXts8n
TCWQ0k84Sbr1zE+qnQdsxp+QAAV8RhWMYcWnOnOvtxl2MADSwqcKDiCJJCFCh3sAauTvCVBtyUHS
x0b28ea76E1knMWUuqH5JNRxoS75zj2DFpUTCVlQTIWOJZjdVEbXdFnWoutq36O6k1eo5LeMcboe
NyE3lMFeZ551OCBExNoKrr2y2m4E7oabEno3qJd8rKz7vegqWOuk3JkSrwtLUeDgDUlIehSAF/qm
CbcFuilNMNxw+9ETJl0NH+a4c6yB59TnQO2eDGE22WMMBWFSBj+9qVzgd6QbpFe4GSrwLQiCBRxN
f2ctshhiCCXsnpjRRtdmv4DFWdxL8EVn0uKPI6pUlK7KB3fEJbpPETyRZn563F5o1djkC9djBVQn
Xjp7qUITJMpeMfjblMa/kE14wbX9HQexOHo5QRDuoijL9kaVYcPii6hiYPPmyGFqBuiKyPkD03LM
JvhPk7Q/DeWwcCng+OH8mq5pQFwwypFEvrhDvxyPDWwdSLc9SehCCQXT/I3XnA5ynYmzhmhc1ocK
0dCzNX/ntJPDHDD1AeJYKfvRP7pa6chBpeP0R8EMcOU/IfczAGt57Kxy1E7YTgIA6PUAXXESZwjO
KHEwGG3ytoX+oZwxf+K9IurwO5CVpPMJ22qn8kBKLo8PVXktKc/0FJ2K1JXzgY0ihozyB/H0Q5c2
zcBaFcfb16cVgb7WOhUMlit5caYnePCT36fkvgYWGTNe3SXMvyuZSFrPnLn0kj5650kO3rxbhNHi
YSlu+RYrID81Fl8y/QAuJHh3vT9A2QAKuhk12C2tCq+oxpkmWEHnZ82CZ28BmQjf4zzq5xJu6loF
Ec2Zq4VCFu4tgXsLTf8+miCepUWZD/0N8sKSCk4c6xoD5u+4dz3aKaVfW0sDha/hSeusG2Vnjjjo
IYM9nG3RohqGwcW9FbR8wWJcM1M6h4ryHLTCZOwuuyPnp2kqdZDgR/FajXS5kg1thlkQ0kXl/81H
PHIGWmEmKy63xuY0S8fUlpdP3eQBk0APUi6AzbanGgfhnGzoUeW85RHBaKJ+NdsTVVNqbEXhDXm5
7/y261XQBp9Okjrxi876uFEQVB/DLW5ZK3UWdWAiPJ8K2toTrX2RzlcqhkKd+pgOKho2Qm3WwMgO
yYPSNyI6BeO6/MoVE3qzJ2IoGyz8ADZk2iMFNRfJTtC/X3KPWuRFQRXXxLPKNZKS6lj/Sw6N6/dQ
rHuvEUf/RBl0tB5vTZC3+rOWU9jY+F68I3IwGCGYLgZp9E7FeesSNVyJ7fUVzCked1s+LS9x1zn+
kajVCZE+F5HKQEKK8lNqNVZTsmRcxOSUNH1eRvS5GqcTgzu/1nfkJm7K3Pv7KvCk2WazxZubzTvV
IjO3A4FVcbxZpACCB8NvCcT6MSz3s1HEhrg7t8FCUrrQKCFdVPqm+uxPOBpC/pS8Ba1JiAm/pqoF
b7SFy8x3lrCfL/kna4rTkb6vqLtJ/LmBaP6y7xJ1W/SQ2QQMX04X/mbnoye/eEODA5nKZPmgK9Kb
9I7H4Xd9pEzAeTwVMqhTXDyuLgzjKd1LkhQ10sMsn3mZee4kkpfSrjt+h9nq9ekGJmTmjXmc01d2
NU3dnDuFoeC7rXlw2kvRVcwbXUkH/5D7Bf7KuexWe8T4wHJVvIsy0ogd1Y0xnbSblIk+WOTKv+OP
oi6Qs9Hbc7/REH6GqYmpTA/O/cZCs3AoW26XQmpkLMxJ/nWPynFNtHj4OUoPZb3afgQHA4v2kJrC
v/HIGfrqSp8+4v38Osx3GCqjkjfpYsyJXmx0NiptOs8/fZRkm6r0oaqVrkqr+vDlwpr8guQAMWz+
jSrV7/VNRQ/hhkwxtZCj48cJEOaZwdJ8AMKNZDDlm6xOQGFolbeeyKON8b0EKlodtEeRiuta0Q/z
0VCfvj1EQsBLNRg8W2JTq++sk/EUPKSX4DB1efoYiW+pPYubZKXR5KtU4SRg3EQxpRnDiqCOh+qO
PYzJfshtVMzDx7t5u9x0td2vkLM9uXP+MLsj7fP/iAuqjCZm9K99ZDBc+I4yIw6zZ33gkG0YGXpo
FrdlyC8GSf1Ki86ucYRQnwo9v3OJiVq6HgWd1UuQsZ9FwppeyDpWjIw+uBfQMRB4wCcgt8EKKIiy
la/sCW8b485G02nvzNK7ATqYb8IbaeF2Jacr3K5V8+zseXUs8Q7lYCdJFNPwrYXahQ6ZX6BOUpMm
PDa9PRgzk+slpSP6vGq8jeELDUQdp0hfv88l2kDA+9cpPk4ooU5iEoNKiI4X5XSrO0560dEBOqwP
UWpz9mAAxwq1w9x6gZuz9fO380Rb+fFFQEDAQwW04pUNKM5PykGvSyFyXkqAh8mrHuFEf584Oja0
b65T4Y88E/dd8kUBj0QVOntKTAdb5DZ+8JIVg7hwkPDxP9znxwCLPuXNETfJ2dwJvbLO0xV9UavT
A4rvuytsniQeBN2EIWXnwTwlaa2doDpFx+IK6s6UijRSXtmCuRPvSj5V9pAMt154BCEfB6iDODlX
oRvXC4E/rdmvtuW4dA/9uvJ1FS0y9rKW7a0hxB8+nA6fkGQijctKHNl8NoYeZLyHNwtIQ2rbMpt6
AiQkOlOOItEVpzw3l5wIZIpbkDWqsJjGAdP3xOMiT1fvqF1fEB0WbF1GoAWKDIx/nPQhxSRRbxVw
A+qyy1g52e4MZesG7I86IIDep8jXzIqXpv+96H/GdBU2crFu/FAAPzuuWgJcDKN2+hJghRWSGtIf
6NMTUtAVdY+xJh0tDefLjfkExUEd8Ssk41qWWHtOw2seLlZPY/ujnmW5Q0PyDw3i48N0UzErx3Lb
/D3AOylzs0W8QzxJwLjPYmhEpCWrvTONbXr71eve/NnYCwEmXMUyFmT0Vm5DRwJ/7TXdaWBd7CtH
qsRmlGk9EEw+E2BzHFMg1PDv7MQ7YZxbBMJgu7w1R+zHjSUvPB8fQeKD+EnWsXf/diSObbH+4h6O
5R2ix/5tOD4UxAMgFBFodx1LLf1Xqu2lfVwpA/K3u3qYGCeIsXpobSWyZpMVrTZOyWdD/kvq6Zf9
O/o6ATXOVJdRLNuKA1vZR1CXioCIW4a1n/bGxIwagn+XWCCO8Axq9DmtzmpZ1sYA79MRaYMyMGky
DlyyMP9yZKMCoYAGMUdYYFufV1HRlbIE36Ry8Z2DN57W34WbLFfOOQ18vY9EfOabYgtaB6ahMTBE
7/N43/D+RDAauZF6ZrfepuePPOnc/Es/HiPjwAfQgVr5aPFqZqZ3Emd1ABqIh24DsLJ+IJYxH5cJ
vlB8TNtZlLyA7IdbB7+bzVkopjL8bl5lPajgN5HWWsiOga8U9CP6lDbfC8Yoj/pklBOWrq3VsbIO
JOIaYCZd+eOxAjpAYpaCERKTJOCLwM5LojxoyoihUxySbuK3TToih6A2/cwidp4xfqdaG+dW4JXK
hmcL8eF5+33P28k/3c8dV5z9W79yYpK/fVTA5tOjH4xwwAVawgOCYF1Gu5Gil1giKr3o95c9KtPh
71tLPPkrFVTholhr9gtsVbizXSYd22ZpIHSS6KC1aPmt/dyWGW4OP+yd2ik6AzOTFcZwKcveOF0I
Lxrhqb7OLAYVozetdhnGSnbhV2+TtYoge12WDb1fjW77TpATv/SR5JaSqodVQ5grPQ7CJwCNejY3
xYN+TtuRpesGYpxPikxZsbA+SOmb25ywc8aH0CqZVIvp001ysHU6KXXfOSXVgJdHqLGcvpIv77J0
+jigNHfYP1EwbCNFYDOqSsdWARNoUJfc4v4IPCXH4FpDldzno2ehKxzTkquqDs3BHULY0PIBwON4
S0IZgYAIaKsP2jDATTTcC+B5QxRzYfua2gRWiQaJYX8sx6TNnXbSZZ9ei0rwzgVNGIAhxi25F5fJ
IsWuHhuEq2oW0L+jnP1uRGVDa7borlIv34bwARr8oeuFajPxk5qLtgjgeaMFKW5cd2zoU52ApL0R
KTYGv7uxrrd7VY0L4FJsN7IAhFjgaoAEECsmSGXkhERMnXlWRczLgTR+SWKHChu4GrYUM4I/hgCQ
8PLRn3+2ymR6TLB8JNX2OrS6g2u0kI3xbW8H519LovE1God6nYBuaLnFC12You8Y3/ZvfT+g5AEI
SFSBVKAVKlAFxwyHj0bPiy1hvNb0LmLNI74jB5SFxJGPf0LdPXVHJ23oEg/7CX1atX4B5UHbgtOU
QGSNIVbYnZvNmoxQMlHNhN03wdl2zURlsO/zJYgRHwkcqisDM6M/DdTq+jz9tU9hXcEmqndP8mXd
NKzSq7IX0jqp7KWy5J1eH+mG26Op6nWVNeSg3WZAZYNytriQ9ZKQc+Hd/EcjhmAK3K2TQGU6W4g0
CH1w8qlqm1ITMtTp6z+mxJlT0hxoBl5iX4rgrcUVWVgQaoRMZ6tPpJ14ZPyydLGt7hqW8CwFp/YW
jFb+JJT7xJlJCEw0vhkHy6IM+in+aYqSdTxQqDfoOL5oHif938piQrkvMA+2mLHBzgDrBQ+RMxwm
8Cl2POW1Ki1HDNn+n9HOe3514NV9QHDXynfYibRX/jd4KWePAlSAIrNzhzEXjYUHlOdudTRdV6S/
EAX7jPyqlEEbQTUe/54ihUkyemD1Y+j8aI2K4PWuuRwCFwRCeY3OpLUpb+T6hXL3l2NzjbfJy1SW
iQAMcT/fH/k+IG6ManYWWgPGQbrpbLKH03sMxNS6yIvYKnWvUIcAOhzNJQbx7RZB5Rg9iMkVLAI3
wu+upZ3RTx21xuKwxeuhNmDnnWo7PzvOTVn9V66jf+QD14cXzRNw3xU0ro98gDcAueHIX85XYtZV
M2LqTecqelhcBOZafNHAijtw8O8rR7UW8yLH2xxY2Zf0RfR8uiIhtKK6tMp5n7sd63B/yQ8ToRIU
hjE/Xa22DxInM3sqg1tIoFvEcnUXc0NARuooLtHEo4/gWELHpwjTVjaoDd04/CPn+9eF2KCk01O2
878xev2bMYp1xS/LbuaulTuPD3pxz2RtIqAywDu4OQbbPrZcswW9YK/ozPBqWcZQRDm9IVpduhcN
M80Sa/M/tt3lL+slYouEkXMUXpOeMIGjPAXCKQNLTiEA0VPYfVhO5qC5dYk1DmhG29NbXL327LV0
rwRN+NHwjjUr3calX/LvbORYGgtI42ePaxpXKQLhVzjuvE0dTwEIvUOKARww1Km9PaQhq4AgVy4n
/C+QWUR8JWBNZSwe5//fzp1Bcvg7/BsNrf40c4EB2Vobnzl0d9YErUa8/LeKM1+facbeKE++hNTk
l95Qy1QOZJbRpjxJPoIiVa1u4UW9UAQ5zFtc4Cw84Pfvv3FuUv/um+bTQ+cHJr/hDHNUT+F+Agqo
tidSYiBgf+jFawfxmZql5ZXLw2Xbhz2BqHz9PW0pHKEB3I89sdYYz99RS56TDYBbgRgPWJnQnEnp
3RF7vflzQHH1vIdLquhzCf98kg2f2gyKnDbZ+RuIHcXIhGsObDb9zipj/1GdDD2g1I37JQJBZjL1
1b0lRIII5X32Az8lXMQeITr4e7QXNen7coPUrUqqzhmNhaAO7sj5cv+qeerUmFoaStuHx0Dzzp03
xBly/5Kq7l2fKrjeJ5ccKK94JCi52lyZXqN7r4QKrIBVTMLmUZlDDl7/VA8JGslA1ZvHI5+TNb0z
mcMdzhZzIOCpODpof7ElS1FuR420Tg6+JwQgAl/X1Hq6+tUvafpndHBLlVT1VMiJk8s3jH/WBH80
9db3g4agoAstyPMiU/CnEBPddrLsQfsJ4RxzPfHz7LWfnB8Od+L0NU+uuIxFkKnlK2l9Nx6zW8vT
W1ONaL3So9NJZqY+cn3Ih3vcDXBV0vhQXIl+Azh2QaXozRPm+MQ1fZoCtfmO/NwH0VTb4e/dVWUG
NBbk+saouSMVjxEfyAtlBsKbb6Y9ULDLlLM1ldz2ncDfrWDZTpnPoguTuV3zf/OUG7uzMu8QtVTJ
9BP4BouW3flX3bo3Il8Qixcn92r11SGMOA8RE41VFyEheG0hLJQqjeyZ4zUrIGtvU/4uz1u7tCV+
KgYOl8BzLMgZdTglllKEQ3Hy/oBUBWhBzDkEMQ1luDvjjJUeXX7+WOyNPRVfIOPV65kr2hE4p4aC
ViLza3vrb9pSBru6dj9Sr0psj+vOFdrz3/fqZR9Cn6iMs2aN7DrCBA0S+gCrEriwG59t5MrQx3W/
zBgVN/WnKvIRgixwfswi5GdqAKRN7NObEtIwdboxQO/3mrzbQ+1BVK9+ER7kJS4w7Us0W423rlfv
uiiKx1v4GIK/dIVPasbwWIhsCDF9vm8ug/B3unePDM0oWSdN4ip0G5khepBmWfLwN4t91rIJpFkl
PgyqQfbzu5APHS11Ua4uUZLg3NsoY2UwB4UWkraKVC+AvZcm6QC0T/08gw25q065vjjHhvbK/9Gv
Mcwg36e6g3P9yBVmMLQDHZdxFRKJv+Bf6x1AAKh6RjwJs7PdXtN0fbqcXmlMLzXkM/Ydls/2pxg4
XAP92jNYgBZ9PwPAaxNwK5T2P3rYbRhr7efYXglXK4b2NsoePA451ZcQuWWR/FYN8pVUB6EH92Ec
4QxAEdbc7+ZWFCNslHqg8s+c22ZK9+0H77IGPO/5evVdmdRZ75if1imO+oLdeeTZF7NC9WBwZGzS
TCU3A2KMmP0XbfCj6zll+V29PPZjSZ/9NBHHaof+z+zJBlKvcet0vAUekBHaiXh1/KtSdZyZ5FlQ
OBkWEWsn4qAWCuPBxXLLJzqSjsfRPrz2vXmet2+FYWj1qT2bZSKT9IsWYL8gfDTf10e/IhQtwHMh
fTOpVs8IftT1gchhKWeibqYcXsysUDqfgj24u6LhEm9rRQJu6uJQ05MMl0Id8+eKcNwq5Yt711y8
rq2uR5kSWE55rjDy8HPo6iyI6W3xfh27uo+s1W3fDKb8zN8JDreBDf4yncCZ7cHrIwXYb1hVjNRJ
FlKo4fF0QWh3OO/2bj3iixpyX15vgdZkB2GsOPf6iPWKGsenrgpjjj1i+Oz8il6hUrX/FFlTUwn4
MOiY8fx1BpwDKKJmUrcB/gxmxuAycPpEoxm8su6i16oh6qdv5pxEWXUgdVQBwgidjiuYixZdltRt
n92lPiNGfq1Fl+VXJEJFFri+Hb4Iybptp1zN8quFNWa3G3IFQoH/MqWzQrLxVCcTc/IcywFJZ9b3
ek/gPQu6jYASV5UGS4XFrBykXHDhQRRlOBet8sbzoCRTTtM4mB+sVVHGndkDPtmqbDsntLdesYWW
pY3tfQs3YVEiGHCEgKcb2uDNodjJqxwUkBFkoKjQ/S0CA+HhJYj73YTBPZaYanK5w15pS84hYghO
6elC95k1ejyZ/mtvKGzbufAk0GXi0H9yihfqLxjqsQDjDaHX1BX1+rVsI9796I33oyMjsRD/+fmj
lf2V2/3uV5jAuGevEKHs4fBHJu0J4ttYkh3LnqT3QJuFdVs541OHeRxLBORigHoLurT+7Ya6pzVx
4qjOZLOocYW+AX/X/txSxTxI/q9bR/pM7EH3giunGz/x58iUBEHKKc1pUxuhdh5xnNF60dUDKuGl
DuqnyREHxl71oRPTy9I87+EweKZUngXgBxa1GjbfEaaZqxl0NdU1wCIyttM9GEQ6fDQFSEdcToN+
jZR23iKkeXvxjPx9OqYcJ81U3QPYlzhIutw/AZ/CIsogWAqfs8WZ6XJGd2Ya1fZHWH1t3qokwvOY
wkpPH+OiAhGJsI5BId796C8W1HmDxEL9RoHdAmSRCyQTtkzxnY8KAMakQGjE66Kbej9BqmUOuOeI
d/98yMlPdzUtaCev/8szF5OHLxqTCiXVm8t00jzbX0SmHN8RVfvMGQKoS3XRh9xc4xPuy193vd3W
Utka2QYL3byrkYFAw5aotCQrkrg3KCDwpJ6i9vUndVHbseeBXEcYN1pwsZTpGG/IBWbibG84xx42
DRpuGMESGmmcY8EQ2EiklJa1vOjcdSMDPCSymHo8CmQ55oresoURUxof4ZzgPabYVtRllJ0MCxfl
oSYcwtApvLn61Q0TJojaIV1+ZNgSpxECzKi/k0sJ9OD8E18Ager8rFs4HiVEH7zfGGKVHeBCuq9W
vlPGs/hxy/ex/zr9d0SrC3N2sfovuilKm+qyNCxHgqyqfBPDKpMZD7YKEjYGxzT3aYl4yAeoXtA2
fvgH0iKO3iU0Yck8l8jb1LSJHTEhu0jmBP+8hXrsuDJo/SuFCGFCSPKUbz1o1x5Xcngf5/ZWmZr/
1Rs00kNvkP5dNSqjeT8GZzlIp8bVWIsMIWFRShqWAtQit70SL1St+St1DAhj9CAqrAeuUfC0cppl
wsK1FRaLCkFTBI6/gvHdeNdrwZOU9XN06cPQhZr1rgBdw8XrSsERLuv1myP9fId0X9QW7+XJtfAd
bQKD1WWI4V0gvyLbOy5L4yeb+dt8ZbileRwUgYXOLkhhJ8OBTV02H+8X1QRqXpzr2gTzNB1mxdki
NYRw9tVzY8v4N36THcwY5J+PYU+NYRuV40ZH/bPstQuJcmkJMjhbGMahteLOSqWFnRqqrqIDgzm7
OYVRkt/3l3vdwGsi+RozYgwpJQy2vAEv67fbsY0Jx20hXi+mZIJGInAVgiIKgdwxPqj2N81ekyd0
y1MmRoRZfsrIh54rFshun5qGqfDi//tYXV1M1trgia8yb4f0P2k2NLZQUboPUGiOEd0+zVxqQ2f9
MvqhUTK4MkZU2fEGIp1UqbxHov1XeXYt3bkYMPlOwtLq0V7+sCPjWZoJoapqPxXdA3P34mFP4KoI
whaR5ymQ7FNnSxcoIaK2fablb48UgOXKf5TBNzN7Hqpsyvta7jHKH4ZXeChjzLQrCCIoK1D1M/9v
N0XW7D2l7AqR7LG6AAlEM57tXljbM7Axh0cBlWUK7KNocPRl6HPA43q4PhvhwtmRqtknBDn6Uu8P
fTXKEJUv54swWCQWl8balyOV+auOjqLtdy4vzzvV3g5A9VntQNOBlymSx408jO8OvexYm0I79ppH
SgVzoXK/DeLp52+iSQq8MaH2t37ykZJKYX4xR+gh8HiSJYfLgV1sbgS5HAmJEwUW3kU8zccQJHiu
luGEuNL1WRM87eIiB1MUuHaxInU35NCGb5JkoLhiFKaRzdrC/1+mpxHbi7HhpY4JeBcrlG6ZtgcS
dvvItqWxH5wTe+DAEJU1Kt5ShwkepAWFSxeEmfy6r9gk3ZMDA059PE5pzaGUJV1Nu9U2wY5Kmj22
s7mjG2r+3Szgp/1OhiXGZ0F7X/7qR59LPgEcFv3nsZFu/CtYYAe8+VQ/8ZjmHPkzB6hny+nPcfvs
cYyyPeGRFQv0NuF/v6qImZoUXbZbc2SHWUpiRfitsZnoJsHH7QvvKp+43+1NUStptLIIArRopuLk
KodZMVMPqwkHTpBin5zRg1zBUjZHX/GCoRL0scmeR96ftlpWl0Ki+r/OrK7vRKV0LhUsf/PBnJZp
TuiFVczpK2UDIPcDKgnjVGYzMoHrja9hT3a0NmcsN4UszPQ/Ie9ehpe7AslUXafgZpr9piOmKBTN
dXz30hyQc71/ftzPdv8/YjoKA3ar1pF6P/hl1sWqmXNk6WC0cvgkKoPKDv5mNeFq/TDywPwZFR/F
YC9r3W4ttCF329UVl4pES91+wyd05wi18WbHt2GvXgzaXL/eB1WZUj3RATnzXg5zqgvv0vOIz2Eb
ufhadb0pwPbhzoU8Dwn/hsvNzp5LBshPUkj5HLSmDvCm+vL27P1dRq8M94+msPlTBEf+xHP7ClLO
x/UTheoDDptLCUgRJLZum88YmAznyWawShU3NmTYaVxQ1HonsA4MVyrso2qeKKk05YVojuVn0cRo
03hitoJ25wfxnV25eqKvydP8GFt0w3xgjddOtjhREHh4kooY7ciYFieHrdNZGPMK0xiGqVm7iLB/
4mdRGtDEx0rezd5ke8wUiXN7ekEtmYAxCljTO4XYOmod3xYE/DgNVXNVJBeYycoT4I33HWVyNJVL
pVgJqQZPeJJW/m4oRtzPnB6yYM/s5HvoEd7JDB28MF3/GQpyCaVz6qRoJefq9337GmdIALsGzH5r
+TDKxVsSfZB/FdHSWameV5t0glMqV1Vor64FwyTt/GhsLxxqQcSbWG83lX5tDEpwlwCYbjHTyOp7
ZGtCP1LvpCQVylNunFckNx66UO+LzfaVoyQBS5GOTRNxWdzJhBMGFxsWQNz5PVVZyYLdWDz/pHmd
CS2f5ydNO5wKiHToSCNQQGc4zVNDwtp0jNY7pT1KEsYwG0omkiDx6rMdYJQHJZsbqbTEzwyhxLoy
OMWMGSpXDaDRn18Nfel77EJlhACn6pbkHacaAkswoGmtYzyvwGSHEvWWCs3HkDxgDrA0YRxmOLCr
D7hLnlEum9zy3ccPrYcHfQy6bFnATjz6xVtoNKs8wH1kXSstWhNexq/wLx/84+MasytvvqR+rpNJ
Yb2wteFLMI0OS3JiPL0LwICT64Q5a3LyMEKi/3Yh8AsFZIWzBe9S5IJizWcuybAirvqoI/my2vUx
lKMxibR4vATH/QXbWAM4jX5BHlC4ApHp9wRJnc7DzmfcVMKvC0QhDlHiZOYu3qNVz1iadhKUCwDq
SJY9EDywkOVu6GdAJnU9mp257lErkMcTWd6qrzeZkaWZ+aRbL6Sch3/225FvcNVn9qBQE6gnri9W
ppGEO+QNO+EFpVk35+5maOORxA2b5Kubra+d2iRqgJV6lkux5S9r7NzX8IeXLCC5ota/rmNaJs1I
tn50CoYjK6FjLHrsa3UrjByrkoFgb0uhS6qRZHiFKGE6bWtO+3VlHS3bUqr6hrXyaTDbqNFTSyWo
f+vrU4mAP6cHDigWHLKp4XaK/r/vUOpURIq9zcctL0bWXC/4mJ9z91rapgYQ8i5AHM66Ej7wQyH7
GdUOHSm+jOCYQ/+vosy4fGIR61XwqtNygLsK5EAml+Jx50Vej9sZS3T5KLfKvvSyFGCBg1PZtGm6
i0RF/XqnxgtyJnezP9CkbEXQJBJ+euR6JN2vS1JzuLDuIRnB1rlfzDVnTxPp78DKGV3PZqjaP6kL
CTeMa9FmWHNqR6UxPf8ckHTeF4IqGVqUev/vC7XLZSWcGyZbjgJOTeBkmqULez1Qy9TMYFkmzHks
pUP9Y4hJy/9YnuQ0SQnyNpsAlhLYyiwXeRWGsUJFsjJyA/Lb1WWbLXC3iBH9g6SyTUsvhnw3Zte5
b6hLS6x6C3889T2D4R04fB98gYYwzI+YmgTanKXvQ0zuKWPXAW6/KHToU5/ldcu//Zh9PCo96ky+
2gjfW54o609OE0pElXGzyT2C49LhYnFdiyviXLcRWsW2OiEKS7iTVX/CJFtriXiEoG8e6rAgSkuO
YLOteRQggKGpvlssjT48g1vjmCfc0ei1MyMp8ohK4xVuJdlEaxTXK4vhohjXADnlQkaB6+mXS7FM
1fo3GzZnjKP39QVoaYe9HS7TJRSuZGsRmh+s/axJB/xNlfFlcPD0d6g+fLKJLs/F0pdQXhdzI64E
Sp8IJZHrzf2Pi39F/vMUsJGMLQroMobi37XTOqG0tO+6aMnWVMI7+ATsgN8s4Y4fP1N6MKAqZ5hy
k473SI52muMH6+HaYIJShOw5pL0MoTbGeZPWklcJBH1zm91aodwK36v0wIoZDy/xMlbbMVacmpz4
tCKlqAIfFFCrh7qPK+FSHFmLJLOHt3nf7SLEemu8/ob1+n33YXJndsv6J//JFkzU62cgdRhDXqke
9YuoJztA8T5PnQBBd0f0j6xxnIerE3hSfj0wnZIdRs/SsvchvfR8oO6u9AxEBMs/Ex8Z4TA2bkzd
T0crJS4ztasteAJrnwn/vPo6HVW4JRxLwqMQvRN5M+SgRCEKR/472ZHa89gL8Zj5/HOD2X6hdl3T
+yFwCGruBlBF4Ky44blbgvEdyponzOi5ty1pQLy30/6f5X4C0oKZAJ7465WreAkhBHIXIfyTaI+o
L3zm1gGA0IeZ1xHlBQKGoUJhK9BKN8Pma0BbXLAUFyBexY+lgba3eAaqb0C6gQAea2yHNm1PGG91
yz0fgl2tRygxChL3IstmKeF9ZJk8GUeUrmR9rp6eIxkWyXa0Kzmym2kycPZyoABj9ejBdv3x+hBH
b/Ug6FSHcQcnYVn451cxad0xADrGz7Mf/cw4Ovmm1LAhq0JYqBqtzePuht9oxFF43iHf9v1kSFVp
r8lCcv4L+/AHRXvmiRNyEUVs4rM1n3rtLgMXjWPd+r52KxxaQf0ykPcrYAqQOIh9x68ktjUl3sdw
AJyBCZhI5wKzwKqmW5egCp3CpY1z/iHGBGAMEF2mnmS7seS4KaBh8HYI5bVEpEncrKBGjR9An6B1
CHBd1RmnqRvKTU5zM50xkDWRVsiBfZeWNQtPLe7sRz2+DWOy2cC2duhn0CCWK0VkXI/5pip4WH7w
i9vwlh9q27omMO3p4EEdEcQTn4+jz/x0y83+aoQQq/3zMpmIs2lCQn009LZpCPAoFKJUpq+iLZF5
CNCbnN2ceZaIjcVVFLqXkM/2VORIJhZjAXkj6RyB8zLaiKfbbz+B7Fkq5LoBuo0XzkTo+en3OK96
+esnwzfYq0Tizz4K+/okjRt90Zd6cMaY7aVNj6VxUPBrfImttQtBvoFLEMkB6wzPh+Ngj4FdrEHp
6GjNY/ETX84qt8sksDBHklB5vX6+q0b9It59LWutH/OI1XFoWAMmGo3dXHZjwueh9FHtO/LkR4E9
IptqxUgLWpNf1PX+sUJ605VaZ+5o5iC+AWSoK9Xwn2Fxv7XWdK1jGFXFGxfoflygipdywaIMG2oU
2pq+2OteoNIWQn4EFNXHSyK/nv9JZ4rDnYfaGSqAkv44LlEGCv7zFlGL6bKbQutej4d23mo/4rte
UPEvckInu15ZR4/SegFvkXExayk6Dq1q8dpChBD3erZ8z6bQz1N6lkfDdaoPMV0Xste1jXgKIx8T
TSd+wxitithjfxT3RvsvxGQ4+QBeBftTDYcPcEGHWlEZS22wiW9AGZOXs1ub9+VZthEfx56MCrqh
MLtPif7YKeH1/6zEtNrmy6WYemzljrNKP0pgHIFKJKAGnaf5+PgzuYS89iSZ+g8yX5zvGZ3BNwzO
HSOLWaIEorgNpw65yk+VnDpYIfc9sdOrMDQngtbaF/b11/nvfcZLDChA1F2kgW1eW4kFPuKm3Hx5
5A+yg7WgazSwqcg72wPRw5k+1/o3b7ahkyv/QzLLp5reI54ecDb5kOvMAoM37EAvQ3VBmTbut76Q
cGrdblIuE3ovhhksq9qSh62WflCqCtUqrYyjGkYahrIof1o9s75iOhult4rvr7l5UQ0+9v9M+zBM
UEXXKth5KRYGwKrslkC7Nuc/XLcCh6DJmC/5EwO3MHcLvLV/SBNAPIlojsO32cviyCh5tUkuT1JO
PSkonKS4mk7AGoFY2t2Qv/JMm9kBwDWMmE4dh/CQWVAj6BT4zqjTmnoujpJACbYs5JrG5EosePki
MxQlECvQrJHGCZmirQLPZ0gJkLfgIKQtJAX9Nl83mmyElEUk3XyiTRrm8yGREN/MEWhyVU3oO99w
DfPyjK0BZ7Ck1cjwhAq4bU7Dm6EGOWsIrGOysBLRqdzVlDyMYZ3PK21KLZcXE1aP8bCd5u1YF6am
HeB1kU04uQRUI2S7KNWzQJKyrwYK/VOoUIMjRFt9+uUQNPL8LJZ8iZ53f0W+T0R+GRimZCTxZjez
1XVNLuhJa88DN6uBwEppsPW4deejJcjdNLBl6jwwSdM66AhqUDyW38H4PD3r5XizmSU2+91Ktdif
MaKhXDRzqmIWkqZjVRfHYhpHAAqT+LVw1lQL1REhOtLUwM/7FZd66WliDMIh+jiPA6SvdBFsR3wd
eP61j0NxozTeNVp4SbfS56NhhAH1s17a/HjqBOP8sT9lj3fi4ugE6y2wmRunTaERwM7pl4/kCyp7
kFl6v+6kRID1dyFEppvz1Y0NFMShZb1VcUrXthjo3u/7VxnHvM8fss4vma2bYvhJyvtJJK+3ScMR
ETX6SXD2MHE72h//E+JPH20NI4Qb2Q5cj0Oy0RrVcoElMnNFILQLl3T+ZT7oqc4W5NFo4EKpB6X2
x7NcypFAFdGr7nTCyDlboEUWoYtYgHzHuJR3FwkDLboPSQvPoE6MLEgRdCico/gObnQN34Z8ZwBW
kA63vGBfObg6MQueox8YskWcKy7FAAoRFpr4hRkLHqYM+GHlneOF4IwbT+5/XNO+Udxa8qplp05K
vyT28Rr4PP0vGuHGrwfpafpIxjFxpO6zFS1gHxrCkl1W+gC51hVZj4aKCzMqQHy3xnOgNBqyG8M5
cQ2qCXUZ7aHU14WXH7qNdJ11iVHtgEkBkVI4BqOcdLQDt7e4beo+Oxw/XFoGJnSEl6FchLBUqhY9
3XSADHoSEoWK6DTxlNV/hk5rvPOsOeRrvD06YAKqPUivOuMAR+Ogy1innktzhWPR/0hkH0PynU2p
xYPYIsURny2Nb39p3vzUePr2mvHmaBW95zE/dZ91vSX/sHR/ah11hdlQeQal+SinKXRyc2u+12/e
pbTJcyjK7SQ7k63HSL6Aa6h2IUclKHdKGHD51i874tQ0kIZiyhD17Qd1FLE8gDgj+B4Y4Nqgg3bw
LEMgoHSRR3HBFf9ZNxj94bgVcu+YjexneUyFLpX/vlQiWyvF2um/VpnKuYs4XrxwD3/J7I5/Av3u
HVQG1dl/jHugSkC69SW3UkSX8xea7kMZv0eZCmzj+ByOmfV/MJZYO2mK0M8jXrp/PMF90VBKl7Tm
8KWCDCcpxga1zKzlS7KdH8F1ovZroLbzn6CR1K66wZvIcn+G6aBJMh0u+lDCVXVsfV62PIlXbocA
nY35UCRJcT1xMvIZNbVs2h0YeiEbefyF+8EmEvI1H84YaZquxmC43+PKIIsBwBG+95/JonNa/h10
N2Paw1o96qmqWOsCO4OPYGkRqrxmDBt0vzHLx1svE7k0PGpXQtwMCjJGhuvtnKIBWmzbOI1NL4JH
zcwXA855mIS+whMwvASSKvWtTk1cBD24JHS4dSuIVzHrTgDPOvDUCWMzeRVR/iUv5qkUZb0l7w3b
MEzsRcB5k64cAzjH56Q3WyOZ4cnUEe2repp19kFWdxSbwiRou7sdJvSy5RYGzOMYYbdXRtwx5kB+
ki4RxEnLuVE59/UMm1bEDaqFcxB17Nr3IG8U3Snnv/uSwwGL4myIEiNN6bTfDbT9B4y+sJU6swLa
wyjMjVjPmitIHv/1U6b9a0kOKf354cTmozfL8H/QmEZYHWRyKLD7EELMpLz9sqPjZ05YF4vZO6+o
ydwWaWeSTvD6letFpCE0qudtmc7CkB+IbOMasr7Bt6TRSItVo5HImpP70XXrdMSuQPVKD7HjpNIN
Wyd8TRh5OVUvyVDpAT93uaZiqoTETWBpWHEgrcG0lbMULZYpjstxIbona6+uJ5U6mfR8it4nXpmi
FKh3ryFaOLkLxX8RL9jw2UeFq4YH2Q9X4lisfxKF8h5lAPL4SKHk44X3/EPXYmehVVz1yws7EMDi
kEULdyxuBnDDg+Fa7+lfmI/1NgSDCl2rKsZZEyqGxKEelFEDc5fWxVZIAN0QdXBb/SvIXAz6yLZW
LZ7aaCdSJ/cTS8biWVZ5DnX6Tq0TuNZIoHKr4NNziy64J7FLLFhrKRrhHAIyNC3w5iku3WHnpzWz
5Lz/p7h14J9BcgOfwDsxx/ZP5/KwtyTr5C0Gda3qQPDMYNhl/PhoQyf6C+4tztq1XPo0XYwyQ/iC
Xs5vfBWPtlhQzKH2N7gdhatgDqc53hBWBlY5rB+/qJSg2cc1xOrT8/eIOomDlJApl9B5a/0Dp/EF
ayI1blXafn8zWNXMLY4s2hJW55/zYDdmlalhuvX6dJ53+w1Z0dS5jhbZ+WkfK/fJQ4IrLM+RShWH
CHinzQoxOzvtbVQKuh/AkgCYRizddTeoeMPvwz0iBchS5MKcJTRy3pC5ep71qY8Aqyh0QnzEp1b3
BMKFUMUhSxJ30f56wfdmJC1CnFNbd+Xn5PyBYvObPFbsfwp8XAMqIwwmkNROFtkn5nqwZD0btgEm
itH4g7FkcyDe9ug/noSPAtus2re9p5sU9vzoCpqAs+rcde0LgFAwgS7wO9VSvJX5WE8WB5OhO71c
tEckkNMlEcgN6k2UP8D3ajBC6pUQ6Lt0oo5NroqdV6em/U+9F0C9tmPJ21wGig8BPuAgIPkq+rX0
r52Cw/0n6KV0YlpUHk0t6TQSj/E5PqX8T0T630b63u4kpwp/l73Vb7Jy/b61i8WjrS4/6xi+xOa8
15dsXQL7KDKXhcZ6OF2/Ub2lan2vteA0i+5KYNMIZtKAyHAk59scOZDyuFXZAD8mELqBhF34mHiP
zsTL/WYyu+b7iDf7qpwi09mtSeaDUFq1WJ8i0omhW5g6lXnQTZYfbHV1vXXPPwt/Jvd1198Nmz3t
e9q/CvMDakPf/DLVd1ESi1LmR98JqCpDVBQT4OO5pKkSpMuxQ0pVbm6TYc8tes4vjGoPLsktDx+T
nT+HTqxrdyqLj3lw1OHFvcDS8AxgWu8zoPQ5DF0YCBoLEi5dwBG3K48uOmf2Mv36Y7Ihuqx+1JC+
I36LUIvRnsEaN98eRIUtRWMlfDRLZ7Apxg6zxM7fEi08bCjyqHet0Q1vOw3zecYhQ941sZ1KLDTJ
Gbvtb78f2am8WedJTIcMWkrjg9gw/dBDf0hwrQC2En5+2j0x0Nm7tR5zfnGpuBGyZBuo0maCGOHT
fjLS14VHeWUMB311IwCQCs6rQAdI/tcd/klxxMhqmFRnt/C8AAAHMsoFp8P23ViRNWr7ARE/k8gE
UYgAM6gWVJGBWjb60tFaMOulr3KYQmmegXdiF98Fl33q5AbWI17m+G0S2FJeDaJLeUrphAUHFlPM
s3gdb0iPVdC7GvK3RSEsoyxcWWmV/E4y3gNJXuync8USRon2FlKwX0IBonnd46gtGjE5ubTUO4g8
yg9whZzoi8CGGtwj+Hy1euRyqloIJM8RNiJGpzOtmL9wdNh1jd5RGVzmFGF2Q6lN62ZN6sr4P51E
FHGdg1Gng4QvvR4lglHaP8pfVQhkTDJ6iyffYYMTlxJxaIce97LzmyF8OO0uc8dGVH/+VuBBDb7t
N8GOmLDOJedxMXZcqeNedDGnWO3h/VcDfpVYBNBzu+uZJw8TYcprsHO/Tum8MWc4y9lSM7bsUIY7
QkRFM0j7PCTbiFwyQxYw4ySS24H2ywRYbOtp0gOVaLZXvAl9kc9tSEltTJshYvvU6CxNI+onMSDd
TP+lIMLnVY1UmB2SIy8szy4NSdRj20Mm+7GpnokYiAsbkiEKE5u76OFD6XgxRRgICNYh8r5K68HK
gY4Wb2qvXnePJcr0g8cTRpV4rjLCftW/OK8FM1Y8cWjHy0dkJLD/LuKxiPK3ZEhcNVq4oDVPDs8q
pOG0D6hCyle/B3RtY5Y2sPtyG04ocW2SCcfHahQDNpI+kUpnOYtdHm9/CZPWGQTQ4u1yQyESHEjz
4FG6eLU/EJksvLJpFqwNs4mf2Q+in/zGdX0fJl1AoT2qhER99y2mIUW6NFKJWaHvCOstNJNaiCPr
//QfdzlgQayiCqgdx5FZsIIpOdA+QoexqnIWGUDnx31D3VsR7GUYOSHNjULzRSAMpjIp1JMfVC3w
Jkq0s2fMFWZZiHxGD2x7J+R6KquFPInTxqV7ojiAH5G6JyhCtVx4abiwF8IJyggr3LaVk+8O2y5V
e3NJ5TSoKJ/7LN++8aq6QniIs7XZw/3UU/GDzueN3lqjxlrEnNqSKrceiIJhAQ1igqJq+T2H5DN9
DI+EaalzuZbJW97r4iFtIVpxYTEPFdAOIGXfKShvxiu1fRkVUZHy+XGe3pfIraYORLuSPFh4GvnG
98sZs6sVkfcZfbOCvS+gjv/2kZBDy7dsr6aTVR+PX8FUXGlxVR+cIE7VxES+w0h3JMbEI4aEwo/O
3WewOntyVID4GRfRlrwslJCFOXq4jIN78OGP0mJA+L0zXrN4VgTIuAuik0UGxJ0MbD4sF80AiEDS
Itp9GQmoOd8OvOIbcfcvyJ6YGMlWsF7xgi0/WV2KmIxEMzkxkVpFT4+IKePoyFJWOqcP/dMg+/SS
NpgEMa3IRumjM3JBGmCYjde675KfmdItMJmpcB5iJ+m7BquwRa65LlOv4G62mB4yBFT6UJHsOnP4
ixOTLvd1H1RUAbvCr+4wv9DxUr6pRWGXuVdn2+473Ewt51n0/OzBbk3dyUCsz2Gp71Stq77dGABe
7s8gyKsqGGCEWigHI+dUYpR+5KeJptT9lWODcg6COHaaapDEoV6Ho6uJhKzJ3yg6giBMQx22YpVW
vVHUGk/xvqP/joQJNsF2mPVZ51SYLg0GIng8d3/U4QHFr65PH90n4JCqrQrbsmcD3QCygnmOtwS3
jHwsK0p9EnoYN7UGtJnVX2RpngZ4dCdQAXYK9UMOTHh+ZTe1q4/8VQZJgk0K8VHLUvqFTWSlsEGV
zOaF3tZm/SLSe5VewtUB6VOal6/aMGVW9/9PnSynnTqPI5SKgMfyJENZvuxkEE2Xyh6gxB5K0qe5
q8mC0CPSbIx/p5/0aG/mIx3GwwRAhYbz5HnaysQOIclgH3ke8IKcr5EYKq+iXor3B6V3bVAb9Fbj
oJ9E64gSahVejSP3sVyXBMS34Bx8et/Dt0tz3wYsSlgOAcPmJ0KMtHidZqYDzPy+W65KeE+BzQWu
6y0ysHSXN3j6U4nx+/9JJqR5HCGjLsskvMVO2XAwhvkZhj4VBkPIBMQEME8RNeD816FRp22f1HUP
xa5L8eoypTMyMUYZwQB4WTtsYcsqUmujt18pNsZuXggynRWvJFMtf1PEBAjKFH7Z70P29LphBrVb
IhxKqhmYktkY21auFyHrtoNegNDha0wRsOX3PZBVw7/+WcYibDWSizH8FwA9rv3jo/GFpSpzgQ2r
ahuRnk+X5t8LT2s3FSAlT/utCyxvDTcp1ZMFx8VFCDtf+OTSCeQuL3weM1iOCmDfbGrJFU+5dwb1
0CSkCAAt4FsbWCH1P+zwl8MJSQhoie8BtPU7V+b1mO/68z8WNm2E+B6qG1H1yUUN/r1cMk24htLM
Wbk/Ue9brsO1B48/6qzR9r5KoAmy7YQ4ItByKBqII1FJKicRio/4AbUP9VfewB/aQ/vongiyoijo
RzeFJLOEu1lkeT0UGgG7z+owoBqtWJjNW3n6WX94riOejgX/eOR/FSH/mzaKQLTL/3KCTigl2214
1v2Wqa2/4yvCQdtZxXgmfbLEbN4ezPNpMlKWWEg/hijeUNDfQW9pUkIcGEdGaVi4M/TBztEVNivc
bSc/LrNi4jDy7ykITC/Eil7GFvwcctceZiuPNtwYe5kXuzx0hslb5uaMm6AtSgelRr+8GMeyOhMi
j5d6lPVCWfTQlkRI2XDA9XblhiNiuNT/02htqmiRIuCtcLODPwBM0y3YrN2nbAyPhXMzf7THqefJ
DLBeHNarCWMqilYN6wQ6tafisFKbH9fJ3vaRx9cHK8e3jRH3Fxhr8QOD2jYlbP2GQKNy3wyO1gwJ
HoyQZV552BC37UgpVym6Ge+V5FbTHOloFlxYGdY+TiQD9/5CZPSk9F2j4fpLbd/icxgVLxj8ZeEG
DN56Rt8TrH46DcJOdDq01hzGkr8576BYNO0qJdIKy0b5pBQCAwpBUeLfKU0LCzMG+q66Jgxzfi7t
gzfyQlWmKBl6cOB24vN+KApMh73SKg2GPiT0vD3xBoaN1hfNKk806gmWbfNcDaLUaEoQxDUZACUI
irmTznB7IYXclePUS2D2EqoG35h9csIMaP7eWwVIJceCCyJEh3U5lgpqAB/ZTgtpzDD8CgvP4Q3S
mcPrE5ipTHW9jhqvskpMl8Y+iI8qsW7Dxbkd20cqccHxHd512B4p2uLVM1qzCUlP7nZ/WOiz5QJQ
fqR1pHPV98Z211rsDHFA5guhWXOaiU0JkzVtCIn68lVE8Jof2ihIZulm00u8Un1k8/RmziyK4WZo
J7X+aFRo6b0FuiUQnZljdeysv9aJfbdUZsAmwNtEbIweCNSciDvE14PcXvvOVdcpxiCYYIJo3jXV
hkaU1cess/csnzAtznj0W5A7pHtNoAU+T039NN6wbP2XhbehZZ01RSESmF0UDe6Mz6Mf6wWhZgWv
PPs7edxdncJgyc7xxS2rWBMBydOw/AkfgmgLxqXmGTfumF3WSjm25Bs0mpwUMEUu71XqjjTkeNTV
CdCvQGnPvKPcX7CUWe+LtYDBoXIucwUb1vLbjJYfdiGxjF65lJZ5m4OVG70mfY9M5fNCPlRa/lwv
pG2MG3Pj3lfKnLx8wu/ieOhEM2cW11umwH+fDooNv+ai4ixXmGsyTwTVxOZ9X2FvVfqvjARpDl6L
ET9IaI7B5amQhHF1vRJiGAr8FWkt51Gz1Yt4A2YSRu7VJ6NGZ9nEzU8nzEktWQU2+4LbIfm7t1VX
qtxD3lQRC+GE7s3j8G7Ydr4A8ddJQjlTobvoULN7nNKXCAbjEfe8uE4gOvKssaMcZFVheKtVB5uA
Qpclb86h4CBxgCZ7UAodwnh2k5TyhQBuooT2dUdz+JF6guJGbTP0l8A7LGQgRd9jmNm6Rxd4ErTM
vpeWm0Fob910KSrz0KIHcO8Z+AcL+K6JEJJbHzzWMSc+9c6nTpxVq0R3h7BQXq5iSakgHPx9FSyP
LfybeKQpS0BxFe46p0FuC0umRbDJYmrF6/tgITSSCR+xJrO5iqoZT5Qmo4ahPBcZizmIk8JK77aP
+DH7Z4oyPoYR3HkQsq5cOq4PQ/EamK/9ojVQX7bQO46pz1ce0Ia2n0LQQMgWzom/ZekJsYtL613F
u4stLGy+eXt7bjGU7EhJla3CqY+8Dysq30OpjgaPk9x7+jp9u1D4RoOTR8NZRn3x1HZptiePIQAE
wSaD4QVwiaTRHMl4I+hVH30fe0sP75rSmaSWjlPxgMsB775L1bMRSgvp4Yx6o9vvO6SCkhbE/X0C
EgmyxU2R09iV5Qm/nW92SVeKu6F16JIr3lLMjucT376/Y+j+Hut8Yo8qlvxidUCLzgp7KplfEcKz
xHAzTso1M+HxCOiFIHKLLXv2O7jgxOOLpd8iqxd0el8vco1Q04wgoHoKD2Ri4+3PHhMYLTwbrYOC
f81IsxkKu7V8WmU02stc6Xn77ECEUaTuIhAqlPX9ugtqnfcVwawa+JIEOZn7tgdwWZWtcxJG/EKw
bZmjReLUdDzqDqJemAcGO4IhGbnNXYUn7ZUP160JBvMB9SGKaYCT5jVlIIawRLmzIE8RVFZmMSJX
jKgLLe+fVsVwUSIfMyADCXbzB9bGF05FT3m2UG1+ktCiilOlZvlEugm+lZfCYIzzXgjnaNtnK2yP
P7v1CJr0T846uC3Ryw2ga8ztXDp1EznCNvcB2jqhJWWvuR/bN9ZBgGPNJYZ9EzlGDZVS5jtHGnEI
7dYR8boqnUAlnaWuDCa86KJKrG8VlnO+q6X0iXnOAEUe7yutz+Kf+0NOtSQ6rC6dxwHPaDTQMFny
8ALTky3e6794B5/g5TBodV52Ws5VV3UxmFOYlw01sYGQAUKUtQA8mVCFJCWWl3TgwqPh0la/Pz14
uP+a59MAfmHc9byN/O5Ip1uZlGaFp0or684Z1vEfINEVQmFLsorNnAYWq7MnFD2a3Y1qtAoRrhvj
gVeATEARXqNLXNLkibCixLL34natRduzzI4wvyWR0rU3UF3LrFUIlAGTLtqIyU5AujrcpGAuz63s
Tt5dQvQ6Q2jzKjR/EUI0ymMfJQ5aYPnKO58Ffci4EfXYr8yJrgPBWHwhvNB6UYWEStFX8gJaxhYY
h9WaYRDosZzygJPUPDWbWwrnvECAzmUqvaJDmI8gwbof66cwZKGCQuMfBQIHXpigF92gl0GYeC9d
/gH9pCl0TJQsD11RuK2RdszuqqhlbwBt99THluikWkr1MZzcnFnSMxLjoQ5aCsnuoSOxHxNTtQ46
pdON1i2hob31lP43vJYKxvqGR71YnKRySd7j9bmO8m1cEinglkB5ItLT15XhFv6rbfQzmIdmS5m3
OxvSoZNeiqlGxyodm4JTq4u1Po2QcZWj3JwTehuHMq9bLdB8gz30ktkcSvezcqcy7myGYpp17j6O
NhRu/5CiWGSo+gnFhV3AWzLTKbSd3kdWkmURhdqgGLgmznIy/AN3sEKMGMO5QNi46Ol/SS1THcK3
Dhp5bpfAnxu1PO862k+A5wn/bAIIW408KpJNKgHhLog0AQL2fURW9opp9i7Sp6Q3uyNMT5idYhOZ
e6OjhQTxSKP7Gs1nya0paMlNAP6EWd/gbnxi9dN0zXVvL2cd/UFO00ylfxRGVHZqVUV4eqoIrM9g
WeYc6bxQAgqC5+Imzrhg/FO9Zi/0eQEzNnVVE7+AV0jeK8c3zH9kXJyz8cXsT9poOnVrY1o3JK2h
26pbGWVgJM+MT6zMSMtqG6otP/C6MQEsofxTTyAOrD0AEu7qxBk3WeJc93n0z5r9QkL9tkalDbHP
/NcSNd3nGupiGfDdzU5tTj+vrd5DavphIIg4L6qabieIvR6BuHdPU6fhMopLjmrOhHIvy1SEbhbs
4EIar7/BdkojgrtQUR783u0hrrwjnf/bBr1Gv6cc7rI3CumYNwQv75dV+I2Ep8ug2ZYsTA4cLzqt
rM0LuBDM4pbVeci08v0CyFVkkIBNLCo/o937DPx3p7N1hdNF1ZQcBgyqvR5wF8Gku7zE1C2xbPWM
0XN08hTpZ2QW4MeCBF4kuB3McN1+/+Yglld28WUoszE9Y7Qa1MjLPqbwrgYOxma6BVl6CwmwrCa6
3nPuz3vVg0+NqAlPKXrCPdhZgLONWxMruCQav5JUxWjKL4VzKym1kMphlZAun1s1u2XbiAXjpOx4
kNABW9NRvaG/Dw1oHrdWqUj8EGXsp+eKTO04kkMJ40udSjGuwG+Swp/J7lexIWryV5z/SVRROMf8
1H3g/3x2wCsUgqknpyYBoLow6oZF+UNLTxCFxchWFeahO+XIX3+RMWeGfvZQ/VzadEr1WX0t23+r
EsNPTO8z0R0He/tV6R6edpvN0Ar5MGRQv5jL2c0UPRgACE85k4U9yysdliJT/A8lJ3ET4LQbA2I3
oePBoPrrawIz6+1CSjARL1dSqhzJiLgEeRgBGtXlkgY09CDGYem0f1HrakSHSCRV6FWqUxY9IzoQ
F8KSqpy2XUhR82MXp/IA7aPHUS5D23cnOWkdRk0hevUrG+pm0wxu71vZU/2GEfnRqz6hbgWiseag
J8wCVZQRh0mGsU6xF6jfnI+j6F5LujYI01xzPrecgOh6n+s9PM3jMVAtxJwoz8I/uEebouw2qck5
KED6mGqfSxEVfR1fKXKHEWhFeSJVaFo6CnlD2mylPy/ghUZZPnrgYiEbGHqITUxRNxr/RD4OXL91
44QURcTmKGMZPbZ3gT9lrfemvwCkHBHQMyfGb3sbxZqEJs+vRaZYynxfWXi3chMEJK74r1mIZJtW
0/LmnIaY6nWCLsZGTr+cZdQ67yzbDBiVgIwpseaTJAoAGwcdbWYJEhb9REaDAsTT52W8Q84/oS9Z
2vQAY/qFUnqg/ZaRhtgHB/y8G7yuOeFqj7vtB/uXRQihObEKsrlLultZh4xRda6+JXiEuOHpcMu9
y9y3NeBHqqxJOIxu66V4oKUacy6GrTRBRArNNBhcjJdEeYmUGZHNvN+HDuEHy4zWS9/UAMRNbDiK
y9Z6CW38pbzglaLhDqJwsd0x/7qAmwjuCeeXQPduCI+IxqGyjWIXbGgBFOk8agoZyvCgG3R0iRdk
Em50kGH5IDONicwc+VzoZHnBWgLKAcvkFnYq0g8SGZY87Pot5/2sWAhBhqu7IIunHPyZyQudqBgf
XrXYp5+H5mI9AuWZ7a7MYQ810pa5I7tmcXeFBLuuVrCRhuhZx7zwz4KaobNvGnW2XrL8Wu84GiE5
wh2M4QbTcrhaWmfEAgTmKEnKGCtwKonixLmYX5PRfpGLDbAnY4erYoulWOoJi9L+0W9TXDRkXyvZ
DMr0K/Ip1fJS6zW3rebdKQbWPgsLxz1IZNjJOAZxi/AGjF7U1aK6at6rJVUqJD4l0jYwFIk4yMH9
KUC6hlJukwsyw3lEkXlmWlFtU6p1GjG6ebg1C6GwKL0hCi+ic/S7FJCSAL+I8t4q2nNOaAiJxGHF
JfkD6BTy2fLNq0XB6dO7Om/TxHhVTwH5awEyoVbmrQdMzryQbJJNB7Q/EyBAI99/ow5he3kQjfIu
ytWW2tEEuh7vYyT4XMoBSOVhZWu+bG0yNqGdE6R3K4Dj76xSc9s1hs/imNiAZs/ahMynpZskCkwi
Mwi1zMAy4EqL+Ps6DStyEtpslThbHPySpxLNc7FH75RX/FGmMzhEUuqIXHO33ALjRNE4yTGyvIDn
3Es+tzwNTQH8LjfcZxD/sUZVwOnTeQ85mLg/F2Pm6cs9IYLWPdgSUFgyeWN1qc6amsuV/grrjeT1
IX+CdXOoU7Un0gA/Rfd9KCjZUDZP1gpXsiFrvtXQ12Ue91H62MWTCzObimCeCt63TfRgmX/4o5mJ
Ei3vvTD/SrebVbHqQw28kYsm7Tg7AQNiX168KtRL3Wa0y4rXxi6fPuXj9YZVJJosdwXiQ9I5zsnV
jDCyMKp66fMJsDa00hWBL30uA+6xQTK71TgVqd4LsgJDLv3fuuSHmg+vAklXQmDfsdcTnx4JGs4b
luxkvuNcSE8losZsq2EU+pv05u5ADK40FunqeopeGTmplC7y2RGhlOo7WvZclQzwMShjCdTSO64e
Jd6dr3euQaSIGI6zCdlbinJLryRvrTP2vdbG76zViwE76ptUZsgImpUwI3+i50GGjxzcJoXMVLsU
gxUDFHrOEZ4fuA3XXIaRC+CYn6ODjK77Q4UPTL5CQ3iqI9NM6NJRzlbK68LB+nMzOCYO6cNdwbMJ
Esur7pCwup8pFfP4ybqTJa68w6oDFX+6HGD7vsZi/DGkx0dLIJU/7dbkkSUPXx9gsFVIzfKnkT+G
WtC3/9I+cHXPMaDFiQyFKXY6Pm5mTB72irH4DkzK6I5B3DNnSpc95TpMiuLMMcB06z/EzFJPcXRq
j0m4wPBGNw3p/92fY9GkqeZ4U8k04EbRMHDq8n6T7nCsYCUp8jek+V6AaUoMzUuyBbxygpMFhTxI
FuWUdreuraK+qIBwEygnEHRY8f2j9vBkLjM3YJgrHl2fS46RvNo4td/u4HiD1Cx+zirEFC3Nw7ez
s528VKtojfxQqTWIK4ix8Ux74WdXGoc8nr5nXsAGg0RPOnDxsCbrv2VlrlP+i6Xpj3sN63G525WA
8LswYuO6s2QU1hOCwHy2mWnQ9ek/0avRiydgJZGfFMan93GOpvU8clRfWuwNNCF+1dLxIioUdLHt
lNBoqUhTKBRztZS0o1BYu/i27skLmtqhBTXvM/r04Ilx3ZSmcyWt2swKjGcq2aF0VgJGNK3yb4db
OPPlLA6l6cAQf7V+y31OTKOmrHipXqE/z5q+kl3CHR05IwvfkILk5tKhV5DI9+jfNybDn1s4ojPN
jcXz251IgVd69m73LEUWjYrrBO0CBt3Hnx6y5r7T68BOFEBXC2BBVXszDeZpVcglvHYobuekd1bB
VE1FcwDTLR5A6DVdZ+VnfPttfOV4C6TCkgjFs0Cp/aXcoSBbCJt/7t2keD9m5L2VQQMNGGscNPHX
utKr4hjhMKNsdddkYb7noDuMXL+2YjHklBDybnxGYu9ngzfnfqnf1Q7qE0Q/bMSFlpJwvy0eIDUC
AgWe2/RF38kmS3joF07uQR1/1BxOjxo1XQDb5Z3KVItEsuawkbwPjFsSPoSt9Jbsm2SwmPxuL8CK
gfvsBkGD60OJ7i933qx78HSv1hPIoaTye027JQ2+vIIs14Hx207hpO6jenBU2T/Oig2ac+4Fikzm
k21epremqg44ykfRtmtwrr37XWDdiLdcy6W4/TLRtgsVmXbCrr9yvnDLEhKjKxfqLJk/Cul6fPRk
SmYllyA8Uq0Yy9rQWHt7x6PN8fPnVzZ9qMg4HtBt4pZ4Iyo4iNSdt2OlFWxCirjrh0yx6nAlqTNK
kU4+kdewZ9lhPCElkOtoHr8OoSX9o79WGJssSr2mAeYjZGtALhn2j+1Tno3zkrG5t4rcZQ1AqhbU
HDnzJyT8TbvQcnL10Wau4wv2AuEUNmoINwNcuKmOQGtdayODZ85B+1drVMH7AHvMMcNw7z3UZ0oI
Hw831mAoXzlidQ8Up6Ysjst21BsSrQoMV/Y9IjM8ZaOn0LlmOpQCXzUdoR+fG3HfYmJaKsHa0JZ+
QSPoYC+iRri/qIdO1yhyiAwHX32GjTWMbNCnjHvNuWnSoTulUrwirD3xDZSBg124dh4X5WSbVGqy
AzycAeq65D0PQJACb+lW871G1dYdUvbeenHc7Gd4koCeSeAtDy24v6KZ23f13tRXLlW590/W0EaR
mLyFI874BIq6DLJv3SgxGlqWrV8i4GzoiCH6uq2I3lstEIiCKX4PW8BZXz9bD4pzmcnBx33RpStR
YIHThIzofaGbI7SsUYR7L6aDxrKlx0EBSn5l29rzMMMqwNaM/RCUasPTf35McgsYAbRyDKbV58Sc
oUiPkPWSdDRZkSn5RIRv1/dfo29Rd+oTTPcICQleDezlzhXPGX/b1fKT1SBiZptnsLykVKZCTCpa
swxCLflI09+1e8agC630OCrRGHV0L+W00On8sLYqaodBV+/qO8iZ8EevCGESoQ+Cw6u1M1S2W8+m
9bz70xBrj0FPk75u29tR3yx8ubmLe/v5AcxGl8ZjYUtBzy1SUeXvodugN1XWadigjt9rk/qNuitx
gYF1uaf6fTLEHTnD5m6RTHUAUjJc9fzXujUKej0i2dbtY2/4xvf2vnXQtUxtfYUJFLYJKkJMdPXw
WKOrlheH8RMvJK72TuOaq2UKsBodBwJyqGtvRb81cf0yTACVHL1V44cXAAawB1/fi3iR4hYjobZP
t0YyI33v0WAYIo6+Ddp4jPyIGRQ/KehozsfNGlWMBu7KVIWQUtaAY9kosonnAvw1l3q23Xhk5/J1
trPBF1aQ/3/LH+BoL2ck2frnHkaW1JE6McyGB49aEY1WclvW9bMuUy+t/tTRaCkyilK+342L/nV4
/VdRN/5wxZjhCygFzk2a1uHFvN3X4CqtR5WqswErejCVvWzF3LZ0xCyXrWhTzK6tbPx/W3HMr/V8
6649sTGOx2SGTN+4sRLMxiSnp7/oZYuEoBKs0ge/rXWqtqf+45/IQUf5/Dpb1b/Lhwxce5cJbTvb
woOGpdJfRyl4/vZ5YmR0RLc05jMqs5NaCUcer9GWnYZK/D28nxJrEqPXzDOTYxN5xfO43Vx8zQvB
22zteBiRdOvne71WX5w35fnOVBB0HkALLYvhgGzEfiQs5YJHU0U5Gxpc4IbLRBO66JmqrtBYz/X6
WPLSt74nHvh1nXnN5EPzUfHn4KiUJem4s4mF7sBQpLhtfd4OEOaroqlLPTm/VbXotmPNQD84KV3U
54qqw4/7250m9sR9ZSYd/zIq7TVUCsZoN0s2jekKttj3e8Wf0hHYRic4gt6UwCT4qk132zpSoDOf
ky+hNbfACs1toZNlI4tAQnmGIydl1KbHNEqpvbp+6YPfBnsrd5Vbrqzrm+5jjx5WsLTIPxv6Adn3
uFDPlPIdNuAUTpc7BxtYLy/zJLoo9PTl7K6cmwYQvTPUtJFTa7g/t4GxT2K5k4HUmtnAkh1zWNAH
zxDHoOAKVMumBjpjc7gU5uhVEmNoBisZ6PDZDsV2h4+CFGeRymnCD2SPJbehSncaQtC8El8TewRf
ceL8pYy/uFfY+rMykJ0xcUlvPYM4xH5OO/nCmsa6qDUDIBQzvt7cymWNtqSDFOiaZ0z5iTFHcr4n
losp2CGSf+/gEKPt2/QpPvhYQIT91WiSAwZjKBb7aFy4p9myfSLMGEOkEFrnCKK16o5JH1CynoGX
o8e3JpSmJailOQz+krMprbjywKH9GI5ZlKVRyiSUCKr5PFqZq2xbva6AJvDv6rbwArcvKvkPVcTG
vw/J+kFlTpNXqEltI5X2b4q9rTBPUCHWChaZoUwQDXQNYSBQwvHt5dOMJXTe8vaSpKOnomeCwZmy
cHT1TsftSVdEZfqFxNaMSQE6Sp45qQAEBUPTgmsY+beuZLY2EgPoaKDy+ekVphRhi0H4f04JWbUa
jssxADcWhOhftBv+7Pb5qm+eoJ56YdbzZoxncHeNKMd50lCs/XXNgsAvc6KVvRFK7zg+iHRboCbs
oTgVRXw7NjxGbvyQWfdrSMti8tE3x2e/hP70ceBV2eeZ6fnDk80Al59aAxx6arCg5O7V2nR7/mMk
jZ32d8EKVqvNUnS6/mwF4kstw/Hdr1en9zC7TRTLTAdiYoFV8zDRp6vMjDc7wkgGJOqKpL+thQPO
6IvbBdL06sS7GaiOh9QjoUXSiR1ZXr/gIfB7jxjqBQkurOTn0ChamvVOvgDOrK/uGwF5Ax5doM01
D7wWyXL1JEpAp8vNnETE+NlXq8A/zU6NDbVSZj+p+eajaLFgPWtmNUVfdBnny+a095S+XRMNLZTW
2Dk9QB2RRHhGB0VxrfRmeNjIHe9Xh5dLX027i3gby0gqnpU35yERPlDoeqEmsw9fSUIJg0tlXohJ
J7I8X0r96DYWpzmqlfXNZuujSiZO5j4bLyzoEPC9mSeXFjtGWunxElthdrjMqlZlbybmjQfVW1eu
aUJprXO8MrA4NZHGUhrZvt+KpvH1yc+HNlTuBctI9ctB3A6yDG6Bule27Qrs6IaQY+hYHc2IfyLQ
t88ti1JBJ5tkVGpaDFONpAAbRlfg4AXK6YRoeMAODLQLd9WjHhmC7y+VmSpSNFzMt8SlwYhiILPz
843ra6GMvliHpkfiC1kTsuIJhjGrvWDJzkuNUr3hl3H38KHnahDrTpv2kvAyxS7aT9K5veJruskg
/n2WVpjwfPnlm6BSsDt5eLJkQx2BzdFxs6EG5AymeJU94IAB0mG1Zi2mC4oFNa+YUAL++Gjm70+i
S5mjn0xwEqmkm96+O8w3nM+X1FIuUsrjb3JgaNEP+EaqwKrv2NHgnheXti53MyTnyAXKqxZtM3wO
DckQHqb/F6+qAisUm5aBKE+hSo7qPhWqeO9WvZzh+mwbi2rF7kA0VGzdKlVzP/wkZ0X3rDrXl6z3
dq2Ngj1K43+LSgHWLbRERG5ucsaEVuFlZSoIvZvq5RbLo9EHe63g69YqJzjyr83a6qTccWGlcRKu
ChpOARj8UMk9VqlL1+4+nscMCZxSPKlBID/Hv544at5BUC5TJxpAUuhLOolfHbjyYPQ32jyCXHLy
lQBdNhyU/9D/XG7MapSPbdzmot3EmvbMHH5QSY4O6kRPZXttK9XmpcJSRR327cVPiCjIlFmenxtZ
TzBiDTvg96GpeDOKGafVrZ1rPT4opTfh04sW3mJsAvb9MBDbiUqL//nttXbBSptGmjm4GPKY/3V9
f3lZTRmU26fLRZzqqlY60GfhiY6y3nispe6IAnz5sO2IS5RKgKlhCGA0wyyWL08YmVXsawp8oIWA
pXPM7XXBNBOCJKc0A8AYYmMeVeWK5FQDH3HlhMO27+faiGASeLmq1VsjkKdekmxqU+E7o5du+4o5
L8HcEg/rW54qVJ6CnKInndGQ73JpNzn7t1ESGzgGY/hRsrBXssf9mAkJro+jj3x6WJtxHG/z9658
2d5ig0cckED5lnwUZKIjTdVK3ZwenrkSGp8DK11P4D3bmfUuJzQYannn9GRpChpmvX2oTAOiXl2q
07MMcFDooDFEWJERgXJamX81tHTP/l5c5G+zNksdNBRhfbR/ygqaaDbe2W5E9b0gHWYOgSTrBwhW
I6RDW6I01RHH0bok8gXyUMC61i2KwjIWbNBnjIGzXGC+vKuY5HuHRTSvv1RayKZtH0FCVl7wCX18
s/2O3DUGlfvpJx97N8cw9H4M5eXtNhJxa4BDxn4uKHsRZJ79ZCxnYEClGO4N71jEbAsP9MxmwV6I
tzIYHJbcXFDcV1nbb/p2Q7FR/Qt/MAUSn4OKf9Tn/qIjJVJEN4PzzMJ4VbOO3uCGYP7UEqBKu8cO
fJqw7hDmLXIVY2dMkfUyWoS6GUKPnPqc7O5+D9o32ShJmubGlwA/qgK8Y3jTfK8mGsHgT+wa/yaE
/OaK/P894aUG8KQWyNMS+qs3ZIgX9SyJ7Y9qrKbatRSLQhiML5sCq38yyouvw5NTkrRI/I933vQE
9NSoP4q860hE4iQJNI5RjdouU3266LRP/S2GiGXSdgRAyBKY03OlJfmWdAiwOIYqhY5EdhMCpnpm
xoBB4HqLwZcptV1zF8CucCSB8wNGu5uwNquYhM/l9MTicXlaCvZXNMGMir2oDnIM0TvtaugBlHCl
Gf0u3VXAYUCFcSUGVulZvwef5gayOk11Pu3rNGO1n+zdssCWikrzc9ocyCkZhK5hdZT2NMmmyjJV
bwZnnH3hGUkSEROf5W/N0krajPNcdiq1YELqr+M8WzKimMeLYQ31QdLI/ydv08wVHSIF8f9IUxNI
6/ZeOjOQydBraFgggY28Ui6qv/Ico9FTGpmZ/jXLej3gxdIraf936ZgABovB0Btqsg6CTL8U/WDC
c8JtdHRivP8ncHDEfsYvWqPU8XymalTeyi7UKEyMgp9maiF+bBNjQe0znMNBP16FT7kTH30G3DP1
+0ER/uD9lgD575mILuj3a7LaGA7JsPe6lXYpMYAJ4OCQ2xenPK/slo4hLsfRIwa1UVn/gsXoa/VD
QEzuqoye5joI0oMipdskPPzj6Ywscf3G+a/98UsnRA+BcGp5Y1Gxpf9d0tKpmQBgEuabxTIYE2Nf
jVcN1FvoNh4Y5gb+BTeYy9ovb64KimLGeFfoSpZj9Q9gccEnCn+ELOw0TvG61ggVtqN8sxIhADDL
c1wZriROsnnJsQmG+srQs1hhFjW7gusx2LXH260z/zzZNZuJ+2qCeUArF0+1EgZTM6eQh+vy8mOX
0cGLo/erB4/Om6BOlSe9Apg9ZEtyF77NfUuC1+2MDwDCSl/TyoDmBs3jvYuSN85MqgCmLYO16/0E
tZizukXZOZ5aFl2seCPvFofcE37nxUp3gK50mS1BM//3mXLFTs3FrIfo2mujFkezB444HtwO6FHS
qF8mOIMMbmlJ5JpgK25EoN6WBk6Lg493oR/VIfXDY4h5QREnUvlEzv+wMK9Cx8V+3+yaBLzLlGDM
KrybYOdId4wNzwgE+D1myecwu1hyxAuyfUmRcXW8eHjrvA+9uUxO87wToOEnG+RBMjzsgWDx0TV5
GdSxYsz1nylJFBfyncEDAMZJ+XKlIo96XO20UkkzG6c/puC5UKV4NnTl3eSsbwzmKLo+O/dGorYq
eCfmN6d3gJjLwlENND7qHTwBIgJIEwXucdkoBHjDT+tZKGhTOghwO60dDHmwKrgE3Mf8guEmkEZ8
ZvHZpiQTo5haHDRiOl1rtfuzpHQ7W3y1wbl1fpgUC1o8iofUU2Xsbzcna4h6/DyxFWSVVU+h9pDG
yIoJnbBDlJCQmItobmpTUKDQQFPEbU4z8nu3YGy3NF5Frri6r91yTgHLg2+Ui05+EQrnD8tQQC1b
G8i/a1gqjwfnfXNBm5EO/Yp0WAy1H1Zz3KvUiUHErZePR3+RHg+xpJysPJMFfN7uHHd4cyGdfnPS
1jlFCKMZEGaviVKHeAvvwxYOCs8pPIMOp4wQPfPEnhNlUZly2+wRxaZBebbQgJDdFqAxsTDCLhVP
BcrgMpHTT9TLYX6GvDgzG5BBmSgjKCXSWeoFdRFfczD3EsbfQLjMPlWV8Q4fXW3RBisw3WDh+hQv
kwb88kRINXdoI5RGntEULyFIOeSvvAqSCM9wgBbeWHG1nZoR5NPMeW2Tm3aJBFi76HrgG0McfeRg
Po+YmF8MBqvYH18Wl1A8MIw6tAfrDWNA9yCC8npNTOdoEjunv8l0Z1DBO1bVfc2Q9RfBsRFXcD2m
+i7ObNHpcmytp7exe/1kaq4OKrg6bu72q9KlwvsHtz7CHkVOWkW6jbY6UnDoX66JoBWlAVMrg34e
xqnaZe86CYZdCL1kbDgOpibM7v81WNKVMef7JqH8YoFhehLvnyAVvEseZvEXNO6ByEBcpaxwMrzA
amsFmUPOWUid8qsmv9r+ohmmemtqsnwNRpo5fC7v92kkHocbXSVPb8JoWgzWjQH98RfLp1w+rTaO
H6wpgnt9n/0eRpTBDbI8wIKVzMV9JO3VCit94xM47iwSm5Wwp2LDms8WTTtysH/DGYWc2HXiVkhK
ez2OYWIENEWFCTdwTKLW1HrbPHBnULKpWgbsUpJGPFTsiqJFYmky7Xj7XOGJ3c4b46+cvXXLXZ5J
No1ON83nG2dS7COCdNcjyQ0CvLN61QoaRmBmOZ9eZb3SIGw1NUgg1otg3r99rGCdVnecSqiiZtb+
Xvx68L0XNDh+E1hpe0hWxg4QVYhWv95sORFaMj+ned7L2yXWZ4tXuhVwTAv11MSTEQJ1SC5EVVwf
Il3z4Q46UODWu+70BeUjnZpUoBb6zdcSFk45tzoJHR3n6tiaV/I+Mls9vLzgFoKEzYNqx3BSsjjf
mBmMJkE2wc1xffhG9YRcJCoxHrKgLqTbcXRbIvIoYWwn5P9CM7OG7hvOz47AGSgCcKjMzij3oPGy
LdIEDundM59TZ0hwyURpUpy1mHnLYEF/II/YFjICePXTwqK2zQLmo3jmlug3y7EmbMFdYHg7NNle
pIzJXRyVkw8iRxhos7MNuirJBLvoWrG6bYuQwkVcro4x/t6aJW2VT0J7TIrnfpRsqeKwn9qlkdmj
IcPqqMzg8JnnPwvOWScn0xmIe5Q9A2W11EHNj4q31+QmFLnG1acbZqfARuVAFLJS9hAI5zhUK5kz
RTgWv9zQ7sVCddKU3c7lPX8gMfQrwAGh0VH8qh8rBAj6hfsFV8bZX4D+QyBCX053RSGx5AdcDK+Z
ULFJdtePmcfDcQ4wA2lkjiOaSmz8BFw2iWjYYIsV2vzwbPPzb1yXJuleQRcTPhcZTAZA6P6R0AZw
MLMhYhq14rUPGGmS+waVVVEXBIovojMcOIjf+khehIJUL2etD958sqxJyl3EaRbrNahKVRByyYsB
flIBGacmVNoIhywMeyYmXiXmFE70CBRyLpNhk795ONg8OKugp3csXj0dboA4sYT4zHdE1HPKSRvj
xhbmI6zL8Cuf5S5+rojfPDvqnq+5lDk1+pt+DwUUYq2869kzpQ6ZrZL+1ZEagSOY6JfvWue/4O1x
PlIsD1KgSWUykLQ9aDEttCzGhMAyjz9+/rEBU4oqr2yWyT5hWtODfrk0fmg/j0iApQ+rPAq5hACj
w0rWn1DdxyLZGoKwT6utFgQCKDzU3Q+ejKqp1JosCPTfe4bkP5/ILadP5oBb+1hea2dfQZh+dokP
bSZ8EWNZGeBE+QSiL4wTbh2zsWhlWzliiNigaiVnmrEyXo0JC6tiYrUMhfDyhQCHhHtZqujiXH+p
EBLuNc35VDIwwjz9C0VlfOvhFuhFQ4Mm6fTR4V9CPTBGy3B/kDbRZa/y3ngg5Uy5xEf6Db62JuAJ
m+dpN+f6dL5RsXmtAiAC/Py8pNg2NaCtzMqPtsPPhbpHhsp/OhcAEIv+3CdmfVa2RdvmtwwfrawE
Vf6qbVCd4UNxHN5oNxcFu+4qQRU1HWeK1XRKIclf1ZAf5a/lxjTJJwB64s02hV9r9l/LZIkFmpx+
saf414LKqO8xzyIS8JZqcTKcXm+TvyOUgTW3D633pR8oaku7avsM9WJby3S9Udt/El4a8W5rrXMr
IZ4Du3hwq9Rsae6AMkw9c1yrBYh8Ucci+cp6FJPsR/n5t0OE7wzuHrXqsJcO2ZTUK+LUSyHDrsZV
DppmKwb5xkrgkUo6AGMARKh2XjZFO5dmkeuNbthfqHuz7nbS35S1gtok0NlHaMQLhH1wkGHr+Qpc
A991C/weLk1sbtpYqu1izlZJnmzHyRTPL/c9gcmUxeWl8Zo0kg67wtAVKC02vSGHeWfzUSr1Hti6
eBBhZTpik+SqrPXpOBn+NE+nCWyAkz8YW6gkVBONEl0B1OJTMlqhyQjtHbJDbfpUDu0RzAxIgveD
QTx+xSmGHK+VGybXIek8qNwBl/e7zNxAbhUZifmMiV7W5EzSauwQw/OsmbeRzuaYdxtOUe9b6fFX
wqXnDfbNYc/9K561bNwvthDbrRM3JoSutQW8s8Y9mG68OG4+oKmStZdvH1YVc4GzoNKQrQA18IQX
z7j8s/tSnDui3Xq5pp5ik93dw1x0EdzJlQs9spZ71TZ6ajxztfYu08G47DVmSlO7jBfALLNAyXgN
/o8vkH/qevb+9DVqmU/Oncioktz4LndmLVG4YHAZyczs5R38KcbuErV2gR93QLNxQnzhkoKvYnUX
slTS3+CJVh8fIluYC8aHpoCNun4DxwIYcccRW22UjEsw8yTfWGxciavnGer6gDD/LLyePaoncvTY
3XG4PY3CWGZwEShUrPtEabvD+cz1kIPcxyqNFcX8/lNwnJEhL63OkLXhqk2gUjrWwwZwshBMuLQJ
AvQzzteHoPZMiFp6ziIouXAJRuakjjNPwQkmRerAAPpo+LBg1fs9CFTQyTWOnVUWsSEk1IgLEGa3
8wEsHAv3R65dT5rbNL0In5mCTFJ9RUzzi7Y34KJsvV58GdlQLNhKioUt5W/DUFcde8+Hw3IA/G9A
JrVcLAEAXnZZBEkXRM6qWTleF8+HsbMC4Tg1Yfecgdy17NiJLJrWo7rMGEbBBTtzfuMi5BWEprY5
jBL37og6pbrFeMzo/sLjO3HC7bdmb4dKsnpj2YGLRolpaARpaKR8BEpk4I6BMs8sOmg9CRe4RyCb
QaP5ppeQt3luh0Xb0L5OMz1/YaW8ObvBCdVSXQ10+lVAKZ+APwe+p9wuKRLgi6bD46jDlc1UReVy
0ueYqcMWbTDkt0BYRGo/qWwLtC+AuWadZHD4YOVQNZlKlfMc59ulq48aAUyPwzQSMXdmDW55a6k/
O1fKfEvqAbr1n8CuBjYiGgyr1PNNfdHQVToPmcfMOOiQQkc3qDIpLpOrG2s8IbAf4xK9zfAgnrY8
8KSC2pxeSO5ZMi1/g9cOtaF+ImKmO7efXgbXG3O2AyL3cMenLcGAZBTUmnpXFFRfmcKwldEwinaz
/p4foPVSV2GpPVaG70nIcvhtMe/C2DUO00X9Zel0ufTFmm07xNL3mA5GjHePMhErAjLSc0mJ2Diu
ehPEnS7wvHjt5IFnZiK4fQmvsmhGq75hx/VAngbX0jl1DMrJGZi1PUh9iqzFQghSSSwyOjwdpkQ+
riL9amAlAjoIU1uF3hHljIEQBvhCO4T8isrgJberXGg3qdVaJ2m5eqF66zWiw5kbPx4IjMgVmMhX
uQx+kvy52NQbMAIJzzG0JQdQd0OuKqdOKEAAzJjIqXGl42cAw3pou6EafCjRp1028yhbeWEJ5jQz
iGxFAjHQRz7nyXYzRtNTm1dPyXD4+78scK352g+Vvkpa5caaXdejvKvsMGTr+PxVGKfZHpy2k2z5
xiO6QqCFmwNAqaqCBBWrHL+LMt3kLq/elWnuGwMR0O2ZtWXRP35He2qfU7F48WGIk+IfkdSxwnQz
K7dvw+ByCCOuJDrGs6tB8Ib+IQQlt9spBpif78WjCAUDoRTsv+6indmht9+S3xfeAeVJ5JE7IN5s
oCWeq6SWsv9Hpr2FAAMuhkXdsrGJYZ9fQTb5eYk6i+tZkh/cOn0quU+JvT+yB8bRFuqYov7acE7t
CfYAEKXULYXmAs+YhhgP5rzwEajsTqT0JcJwHSiZYdwEMjfLxb4w9Mc1Z5MTLnV8Bt7fKsYhSOHB
yPJXj/aSub4t89asN6vXjbht5Q20Gv/HggFp5QFW1/doldtAFjds8fapLxvSrDpt2OMgRcJ0TSS3
hT6ac9WcOHZUZQHifZbfz84ImRqB0x0RRHaCe4c8DWVHSQQf7M06qIxP0h7O3wUCSyTMEtk5l+Ql
UEhbEZXuqcF9FL2zd3/1H46xo03no+m/J1+pwHEwPUmbAbVl0KDA3DEfY0Oog5QhdhfioHZ32bFa
ZNOOsP2KJT1MpxezEdgVzegIB3nPZ77krfQrAjySzGYrFPVD8uFkzr/E14aLuqGPScXXDa0oQ5jM
/iE/ufqJpc3ew0v17DI5Ryi391GfvdFpkzQlnjChn9hUgYI87Eh25yu5aOjIWhKGv2xfFnu72ny5
5uJIYCXNBfo+WXQmIaZB12hjxV/0/OhkWL5S8rmndGjJQfs31hNatH9DXri15CBtuVOK9Ru7/8yy
5QDyE7Ag29KchJMV4gcuiUnLAlBC8D2nIGdm9ROcH44DdbWpXKKmcaZCFaNWWvcJ3q5OmmbovkNJ
cF26MSGhLV1fh7xKNiQ0vq035DZXwPu1JVewEZqngfpB64Jffr0zTr7rzkIr6y8fiDoYgMHnt6be
5U8/rLldK1FhWT87cURpuDObtJOgcv70C1TNBIh3WaKBKDpWxmc4+kaNJ8ZCjlBlmtXFlMkQ86SB
7uqM2YVJNPG81p5aLepGDnz3N6wiQlQaUFSk6fpKLFsLSdQ11ec/H1qOscdLaoMy4lNZfnNDy+iL
uqVanIxsjfZ4FeBYDP1ij20n8Gy6qw21dz/Qpj+ts3B2F+JvdPgP2blsQfOrLDARMxSXHUSngBek
Pzo3Is62PtdMUHXVD27OX0SSgN3kmcKnpNP/7B709YQ5W2k20dNLUJN4oebUnfvCscpW31wt0DqV
mCaa5nUjw53YM04zemaRzXe9DdO9kRKE+AIqTopzBCz1mj4GnndsWNas64vZLIsUbtDSMVEpkPNP
9ANVdOqUWns2555ruOOJ/j4xugn2uR4d8nC5EhHV+Rthi2mcDorTsGKrFBjjpf8T4DWYsMha8psr
O4ljMAnp62DB1AYNS3J07dreNM3kXfiUkCc788OQUF/ALtbPZvp0JbKWbiJIhJbO9Oty9L4qDqxp
T9G2m/fVdcbSndqV8HS8mAEqNlGp+o5lcEjJyuPV13G4ZVlXQTtDm/4FItuQ+tz3hMSJvqjE//gp
DhxDdNZqMrA0iOqFpGApvM7Hrl8jAPhGb8R/3n677AL4fziIEUDeyjkHZuk5PwxEMlqU8jorVcgB
R8MQzeaYjRU0h4sTjXY/tWv/qZuy9efzH1wS0U/6bflt9UcHLrYB4JYzRERBmnWD5vVN5iEDxSWv
MI2zjUdLT8WbwTafbNH+hTP+jM55OWijtvykDGW5lh9t6ZUzGaRyZcXJh1pdDRDt8PChus99w163
PDX6rBdhlopm7xNlbd2vofG7keezHm7vCTGrpvQpOxuvjBxOyilxcYy0+5+SlRad1mdahNOZs120
KAd6JM15ZTDBK1TMNhKcPQtbs/0uKBuPjtPp7xhR5dVTc2052c9O3DzWqBz6fwC0peAH4Q0p9xf5
7eO7VGT0TX8mw20bF4TQpze1Wldq+1AISyZwO/QRR2+j6OgoesWnUAOQpsS0pnCVO2Ea8qfX9LhG
4LxppWfQBA5Ua8PULXpzkNHnmTLGfthVZSsR2CeqHPAr9Ovl8qE1SdYdyd9PpmF2Pd4987zqFGW7
7SCBvB2Ie/oSuALRpLuUeNmgmCFM/k+2vOe3s8toYymNYUpGhIQAlwolPM86VkiyxvaQUmCW292x
XebZlXAz82M/H9hlmHFVGDOtmEoQk6BiL/KTIcz7WjOl7sDhYDOTM/3GF+qh0aqzJkKpMvmaEB4H
vdOCRHDt/cRBopZqtgKzRJUYVxWPgbtylppCjfYy1d5TIn2YIUcFRfXGXr7vo4r1ZGYX0ZB9mTl3
bCfYZIAoITmxlkh53uB+UJeJ67YbHzxlNHRTbqvVALmoU2hUiBrIiu2EJ7q+bPYf4kOZHQopPXnc
pTzQ7t1IYxlrA1bxBqgLtL3K+BZurf94fLSSEj/wzLlevhrh7oDudhkBzZ5vRzIg/xeuH2H3lYv+
lytVsMFhCcvaa2/Q5Bzzdf/iUZOvVy0NX4Zb8X/N1Z0ayS5Wum6L5pU+Bzej6gMnJzPIj8olcY+C
W2AQQhEzRN1F7uygAgTWJdw3QImC+H07w4WxOAVWyLvHFOyfamNeO7GH2rT5kyqUajUSfsM8l/J3
IQczWpbkn6+VqFwNCUlU7ZTmjs5EDRpJFqbKTsuZ5C195NUMlDYnhrCxAWxAs4jzohvLH8u7cyum
YBdSCqi9PCIJKRdhIoFsMhM93jg+SST3lypQ1Tc+shPim0AiQU1M7zl+l80ILN2Y8Padwwc1QNP5
zF8F2bfU6PdkRc5drF/HUujnWmD5kJdaPLaaxbUtTBjwf7bxNX4uizCPwJYezdAzBIEjJK8dHKAW
GyCnCrUGkIvLaDIL/7QeItxkDmTLQ4xPuUeY0OchbtBIkrGZtHBoAXupwa3/LtKSBELO84zKyLlL
22E803+X4xfYhboNwHzrqGY588zq+7XJ8W2797mPBOCyeBkUwg9w7uA0gNwt7lW174Ck7uu8QGsj
Tm9Hsi2g0HWJLZmGdwOlhBrkgffijGvcG0y+MxLk3J6BSB61Fp/FCGLJNgT5SQNGnQksTD+3lfhb
FSQ2FowPOg9plgEKUvxSJB10tSdvRzPGeCs9c1LFXXkNaonFqJwE0a8VJYrHvKkD6j30EEsiqKMN
scKUAsAHv+80lqWV9NQMSIOPfFXq1jIi3p7pKt8F6B3gK38jPiDqc8yyYLN7BW1acs0IXBdL8wiE
ekcYqOwj2J683bunvS75xRSglaMA2XFuxrmSiEOOi9ge6lOulf1E5hiRGZpbqrE5F+28pynq+6Xd
3ovt4jblWL8YaCfPIuPQeZCPNmlCclgoYCVnHBCkjOmkGvferDzV3oct+v/1nH1vbA24dJ/z/toP
v69vRsUcFLSm/LfyX0LNXho4UJo0wW3mc5rX/r06eKnbNklnz8FamblmBe4CUIg8NTOqyli+7XX8
/VjCHauWlpQPjyclySuD2wvMv6PpG3xUVDCkwl+pxQIenuBPyXt4SYfbqR7LUFB42l3IZBqOOr06
q5ss78TYPwKUGf2eU5aopTuM+f5EKgyeUHiC+18hi5D9V/RN/N52oHHmFUBZxNTD3XmrZOBsP/xF
yafTsCiZyHrLZ4M8JpLILExC3SPh2bop1swgKNDakqefjudl4EianRsat8vd4QmXanW7oYJJhcB/
PinAxl+FPaD5szZYnvxI9qahKexB/WPyd+zKxGSaLCmwcHew8J4UZrbpFXWbs4FwKk3skbn52ub3
c1PSUaAu8ZkvBN20p29lq4wNVTKMTeNCpfMA9XbyvlwCPBHd2M4UGkdUTWNfpkGG4iDcsWoYeIYJ
htopJOre+EjIcBG+TUbXruVIHxkc0rvV6PLoGOg1RqhKv1zKP5rqReGZ0IZVVYz++JDTneOEtgWy
jZAVbNz0H4HBNw2YJbfJY/66bGaLZjSEGI3v+WrpEIBASm2axnrhjjD0eHR/6LxnqngG+/AcEYC+
JZlCov2/HTkvyem2xBg/XG9tUWfpQXM3kpd6yI/0Hm0Kijlos9k8Lf1QgSutWVSayGdpe6/SAhS0
H+9p/SVIulcDjlRtmM/x3gBfx65K0Bcvng6KaV4DC+rGtcdiER1y4mviSu4Q/NsTdfijSEzvYg2N
aEqliGW3AhGQGh395r5QiF59BMNTd5+UAgJIIMaY2RgqZU3jIxsz1xDxKKxmHfKpmHT61FZKgy8u
nzAhk3WfQ2GI9AAH/YOFWLpuufxnL72kJ3cpDZPTBzwOWfnq6Xh0tANjuYlWzvEZ4Mm0xbntxB+R
+ONb3Fv7JrKh42ye8CAOneE//gLGA9Sk9CjhCDOcnSUBsSqB7TwQEE8aNRgau4Fpr0b17hAQs3T1
8M4ZQm5fV0jerKbY3fbl8Rgy9tb7z6RlHkZKEqIPs9gR4arz6t8hd2itPvtWOvJWyVr3NE9E+onP
5u+GaBxmS8zhMvDoNctHUVxANMP9AWcR3HlVlHh2OzDL3Zz36nDSBF6PsDMDD59ZwNzh8FoEcrgm
T5k5TGcr0wyFfiM27/RB78m8jRC7fusAmDVjCMwTFzFin+UBWPw6Gk5YNQnDwDF7hQaUNhm2+lJ8
I/Jvjx04xeHotEzrSRQcWQRKbJG6ecIhdfNz3JC6TR6k4rZeRoNZuJKaiGbbId1SJH30s7z462T0
3LWB1ZXT2yOfvBOsEka0VCKk2k22ukXWdQ/M/DL9jJAxEmrbjyaqZ6Hu2ExSg4fWCX51G6e6IvPd
Hu1ygYjs4PmPZvsYq4QJUsh6u6BKvHFmTrRM8YTW89Pv99CZThW1xwEF0KVN6ZZsWSZUGVcil+5S
D/ZWkZH+Rv0u86zp9kj4xYQqT0HuCDGR1NEsA97QdP5s1w37jGWSdHdY4PqPjE9H/kauurO4NUhs
sDDQGvYOjEywGhlDEtI3ZgAOVPKUVtl0PPtqF03GKvK4yiRebBwMJgiHt3bOF7UwdxQvB2sW68G0
+sI5H4AQDyEwEIqqpGSsK3ghYMWmveRHt+xDLtqZgBiqOmXbAowCQC5rpSHp1DkYsbf9xoUrNpM8
zhj8PbZewxYRNwkIzGNir7H8zmpQmmHwxvNOvBhb8FEsAe3rcltkU8N9MzenFdw8tVUEvc7RpIdA
6ignWSdBxfi8j7wEQRuaHsahZrgpw0QQ7DlSR/Hr+zDT8UP/KQkvZMlBCqpntpTim+FCGwompNzn
xkiqaNS16jlTGUmQYVe8jNlcrOynJcWWFyRnn+nQPsZKZk9I82ni1Bb2G2fczSBuVYtDX+CMwnlL
yQGgRwS0fnkQgOIGyCM3Y79sPgvRYXxoMwLCFV/qCbLo5BqNXnAa7xq1d+Nj/UgHLRC6bKSDUTG7
QqDDyZT7ZkWeorH8KndblbCZKTAPTfzhi/ub4Sx4R3dKC5aCSnZ55K0RaTJR19BB5pr5jSvk6jCO
kBm7PzuxCCuoPSdEDImtw6Ch6ErMw6E1G+cgo69XnElcqRao3JxfiQQx5nKTyhVOF6g0+0AfC4vl
Ksr45jm42091zdaZNCimpqP8bVYXVdfDyCUXfa/UrqibXUegWIY+Ch10ex9y9nURxCgQEmcTYLQy
vRXdhc4I6JU+mzdtJENKiKmrWnIUhlW1B7Z8wXX5FiV35b5HaQjNoKsYzENabygTxAF971Su2Zn3
cqbApmvbVA31IJvexZxTeN0ajP3IHfhH1eYXV5FNasxMpZiCn0+bkEddTfSSxHDNir9zqJB8X8ON
MwQyczjemQ15nDca/P+wjw4HV1NbagH+TusoAPx3wJClm4X9P+TyU8n06T2YV82wUBGlSeUknyR0
pLCdgagJ2Ii/4OthtcROo/AQOD8e20k9K8GzWgUsMK13xK3/W5HGrPEuiXQQLCFM6o2Ti0U/bHMU
N+4mAcj3iZ9VIVlChuE7GbBCB+R769yEb/3lzXsrtHAyyhLZltQQYw/2yMIACfHOwedBEXOSoygx
kIDtcY2pJrP2ySC3Dlf2YjCwg5sQiKMXO8PiTigdYgDuz22KGKVSN+4f7Y7DsSKV7T5dc5hD1nSf
fcFDIF0TPApyu+y5MqPj8qcivE0d0fN37zkdCZtlR/LYzCRc+eI1QK17/jsFTbbXxV2NJHj1+KcJ
VDZlp73IF0jT9ITmBH298hSkZlwXSBBdS02f9eFxW9/XamKisQ5pkrcRV6nE2T4dlr22zaTGQln1
FZDSiTD26LcEnlg8b/XeXgjz/7xHUxNOLtjREgixBnIL1wpgEeFNsjFQ4SBrW/5X5TlfP5pE9Ndc
POGrbl4I39QAS/FOPfdftfHjvuvFtg/vdIzmZJh34SLudrapThy9MUB0HVj4VSjy1WQ2XRGUK7x3
aMeoGkYKJAxdf/ITrc1UYn/Oy9/dyAiAr4iYE48CY/eUyQeBwDGMZlmpteJnJOCV/JbJuuLhi78N
eCmRBB7DMbltyED+I6xTIEncTqgM4FDJvjCiHcFvu8SHJrnQv0w4+BjGpz6a/fQIlnxkrCS0iCJ8
YdbOiIcAS7gDE5efJtAWtKHV1LTXzHics0tGRaXExS8e0MSqdD9TW7xL6vR0jzhzhJ1j+uvraqa4
qorjDSi53rx0XxKxBWTEqfOJQNffI62iqAOLna0E6CZrI2PP/kWtoCFwBRYIVSibli1GFgYYMxl2
p+hJXB9nfKolRdH9Ia/T53BRs2+pEv2d/xvgVJVH1y41fKBVf8cZamp1ygOq6ddHblLPBPrWuFBl
bFkYAvQJQaDbXp0F8/bvuw7crqrv5mxvQjBaG375byzRqTYsL8Qa2Oe1fHB/J/qAvOxCcIqJAFal
i1GP0lNvC6dwUbiDKMgWcHFtFooJULGP6bO3rJCQ/cbGTcbmLDmqGIfPnUYCJyznlqOkHQmSucjH
FR6PEG6+PwvrWuUWXNe+yUzIHnp3zH0xpgpw8a8Qmd8wQvYvhy6Ia9+aJ6iNctO1mCaZDm1pfQTN
y4lXipmXWqmN5o6ubyzo86hWfI1qrR5QcgxLjlJq3nCPFRrDrJgZ15wtXzOGzgiJjo1RfKjBinZQ
f7ZVM9ABk10cMEWiOYA8eUlbXNulB57sArCPTIXzCXjT++UGNH32No9F6FJ7VSUabmw3gx2hIcLz
qeiqaIbOrxLx02K1RULobUdmW1vEjn/1RUI94iyC5reoNhtXGUNT/aVqeAkOg2IRf0JYrdnSLjoH
Jp72z+4GsCi2G5QqCSoiDQrIDYxnekv1slyRMg8ohfnNJt6Dl8PQWdn9h0YoThxSWulikAVvXLiw
e1Bov+LJ62QZBzijAQzVgpqriUWqSUMihuCcl6qIZFuTywmrLJ8l02+7GfuhoUv+Uw3key4MRtrh
TjJKKvnGztSWqeN7zZ0/wVrsBkX/GMwIftJIjHTwj91dHkvtgpyGuP1JzwcnU9q1RoWub4fpFdye
Y7BoM+/AWtLHHoq6hb+0aL6Az4KsO7J7ciJ9+cSfLNzIo4/pswXkH/d4vqnQAKdSkdrgbh5+SJ1m
LeQvJTKMK1hpdHBFV6K68oXzJUZyekg61MVLgYVOwYfQCuR4P3YjQnlFWI3t7MScIjp+R3eeaOH2
ger+YzK/6lWM7wldS6zkkoOdvqc40iyUg0v1ZcVfT+a2GU9neot/Ll/MOPl6n9IbhwlUyBx245fg
hq/NKuh8sQwxqK/n79YYR7QEGiAmhxrVGMUN6El7m5sX1jbkw5ePmt27bC7WpGm2Np4L8i+mgkPX
pSPIKGweytU+LH6l83+nUWwMhwdQ/aCpkA1kFh3M3JuVP4gcQL59ik3eB3PJZsMfi+RcTQW0G9Bd
EPBBIov2x1estXSnzSIZd1giSB5/gPnBsGl0LqFL4gOBVqfT/lKHUEQOgE/6H92t2Oehxa0Tjl8J
bB2AMT/FEDP0UmUnZ+5VHjBcHWaDfw4iA4bFUGyUZ9UxjOV2SNEOVIK8MdHLKzl6A+JegQgmkS6Y
INPox9grNy/eut/thqccRL7AUtxf+Am+0kZeXEVvF1oYPGCpoZGOLfpz55XJbd4mP8Olw2I1bpZN
PCHQiaBES/YGJYf7wATyDMD9oBvY7a7K3hfQW/4UR3dQQxLTy7el5ecb0S4VzzAASHXRxhjtJkki
6BgW2krA85Sc4/qtv/eqqABCe5IY+4Gn93uUKNtXe74xDtZ10qcc4TyUnT2XFSaYaXACzEQJV7oU
wyYoEpI2qcJ1PODHQDTmN+8tYRz/YUW/PFv9MjS8Wk2L77ioM8dmmZFyR5K/o8WmERs/ywDA9dbV
iz3K4WKDiVZG8YmFxduqiLr87RbcaPtsKZqYt+dqxudmUSE9Rc5+Qcp6rUa/CAgGYqZOfBrG6bkY
P1IbkxqJeowkz+Ol13aEn0XOBWyrAJz/BphbP7Xqng89jyJXd8R9ATCyByyFB4EJKllk5X5IK9rP
Sf5ocSd9CrtNKOp+BuOFhPD3JcXPM5iiqTTOeekd5W+9nxrd30/aHwByrwXDZMTgqjY+FetO2JOz
UY/FmfYp8AXXb+2NonTm95EVZ+qUSZmw4fgB7WOpF0MlOagkhNC3QMNB/kDfI3Feg5I2oqMcMfb4
nyuqAFuG7puR/LYrVXQhBkCtU7EtCUVibPLAa0P+aGspihPrHakH39rTZXYHF2nB+asv/O4qArtw
SQSF0Fg633RoVdiffusirEcvbSbNpeemnk1snqMJefX1CqbPMmAxVvB+avrWFKM+EoknAK5Cy3ez
GgheXnSALq+GNHOrKNqLplf+2xAFa/CcP4igssYhO7Wxi1lSCscNsWOeOE8ZCxbbVmm6YjL+I93l
yvQzcaEMbWsCeUOvKwLvntDaY+43z47HHUvuRnHCmt05sCgkS35AtwSthjQIQWK6S2eKC2MkM/3s
NKE3VKAY86IkZHFrhhGEgSlkAj47fDVb5/dFq9VYBMQvMNnAl6X1p2orxQbBWMHQN1hstm0GsM9D
pkInhjMu4O7kJ3cEh96t06SZROuxnZw0vyvpTRsxLgaf9aI7wGIsG+emlfnv8CM/IB95bWLhQfEK
yvwHB9sgAr2m/S9L9tqvcBN9sfQ2K4sTBRDOWIYc+EyMyNH3GFjETYF2Y/H8c/r6ega/upEivurl
m3vWRDzQ4szl04YIoWN5pANDJ5S2NmZCTWxVGnJokyIaVlfp+zES+0XtdOsqnd8rCWvfX+hryCv8
wuP83oiwlfO3mfn1b/2zLx1H1zoLTupKkR+WR6Z13XKtjmybFGdCDnu24QdtX4wC/IuMEMucowGX
7SUdDqZ2r3T2lHex4RTAAUuXbe5rrxbjYU8aRduCmaqpY0B0CgtQtmrnm7eUCN3NSahxaFIzsQNv
xK9Q0/OWFL6aHiIUZp2AFGnqssHF8PgMY/RfV5V9sgfsur/n/cN5qUI1DnOHJeg6Iyo7TGjO71v/
AJHLwlVf95iR3ygP+YtYXrPXL67rLL4A+NXKOl/xR6/C7TyxGN+E9n7ZAmUk+4siBUJrSAuvVxgp
d6+P4vj4p6r0tiIIanseSOdinZw6NO4+wE/miJ7WlTT2zR5VbIW6iaYnZwAxDpczoobH7Bh0h0p7
LhL68W5DO2BdAVleZo+MajKf3wZ4lsTZxUIJlvufBFB8bwruTBnBErgruKd5eFuNRr1l/tjcbsG+
45XPlRHpVhBwBIwNmrJgI3NI9EWg+ZpnpOvgjFJIH0uGpykvtPuFzv2aaJqgWVS/cZCielM5/Y1J
MBnscj0iCGKmuRMl3u1qdN03C1g8+V3Z39lOvOUlp7eUQMo7R8d7/JD4cJ+PHe1tj4Rl4qH8sSP8
mT2J1SIggyR+Ko9RsO52J8kh138UK4zsR685leQp0B07k4B9H8VOqL+c1w1DwA5rzY9FKinY8t9y
fAtxkAK3XhLqMCl0cyZItAT8uQn4mYgxlXX8T1i6Fp6t4flOKvYWIgM9ANP3qKNFTSLxMIRETb6P
qBcTWkrnzHm4Pd90OgQcyti15+IENAJr3Wwvlbdk4R7Rw8bBVDTUgRiP9hJXByHqLvsOGHL4+hbX
WZBJEec7RwbjzOBMCfu91A/O4dFdEU/O5KXj39syVc2oIF0namNKy1bhCTqlnzdbefOiaY9r41ht
2M8ry4FW/Au4GWwpNWoO1xIexnYbRJzzycBCsJbN5ei0tHzw43IEVPJCSr68pYRo0ZWjdTCSBZf3
Lr5bzudVFnDXoLbKRM/n5sHkzDRWFEEqsibQnoLvuzoEIcKie9lPOW/hH/gePnMzoyZW8mMMDSER
K8W3dmtVzpFHFr6XubwqLgB2xPmM3XihQk9U2XnLMwCKzA/vuVsvEKSt8ElvrEe/6p6wq0u6mufA
VGtQNNK+N5Znri1UmhIGk9w5SYxEFHN60ztiu8cgJgSeHSclEgX2ILPoUjO8x6jzSC2ku9KiOjEW
LEfzRMDFYdmf5LorGJWM80wL8Aj3lbN4cSej8g86MCG0WwHR0ZlT1O3azjC1Stz+g7oef8HVU72U
rubN1sUYkZbXONL7aH5vEHWpuT6uYejBuDptHtLAOcbSxZKBQOJzAYp7OSe8IkISU1sUAj7JoSvd
dtz1d7MGZ6qcFR0kyaxdmilbQbyo3Rz3ZTfNGF/IWgmxoG9fWsqnABdV6KWqrX1wxqWvEPDx66Fv
PAl0MsMn7Exyq6WvHC4UYxeCib4FGGNrcOvo28++wPsSSOHpOgZOnQpQ5wOcAZcSEzhidA7mk8Ef
gR1bM/tz/MZpssvxfs6eFb0fqdpkFdtrUPbcrRiq/p4/vH/PDGVk/d7VjLgvD5M11+D4v4wuGH5F
cSP9covZswnU4P38lZYU6L1cIC99KsXbJoaTFONlw7kyKTunYTiROntCyCNbOKwylyXC24e9m+0J
kvwVkC9o08xUL9Osk7LNMMMjCxLR55is0ZB1Ba+K7YZymN0ILi7KMqr3YySW+MaIAmYdkDtuAJOn
aTGJwE4Jbt4NCDj4oggQyQg/rKKObBggRmKefzSPiGpesaxW3QCa2d65j7lLUj8PNcXAsxjrg60s
DVix2/kfBF1vovseIcdRz5DuDtFPed+zZdABgPg/FTWr7BzhoxzUjlHT3JCctKQLtafLa4xissLr
Xbjqg4CoJuuMYurHOuYS4Lg1/mNTLJOyT07ufuJoqWAFhm4oI40eSHktS9oF0PLNKyGd7hXycOXR
1JIWnbxXB9aB0uOD7MY3AgCEglRO29s9zrLQ7K+iqHSew/b13eKR6ICuK3+YkkrWSQct47k9X4jn
r1lUUebbN+xDCehou7hFmr8KI4e49TYVm0M6Wc/2lZV2svpBTeZh58IOJUDQyoe54IZAoEOlfBE2
T9wVWqeZBqo94QSYShzOln3o95sgu9NGYLOU0VzjjoouoKtxp60yuRL+ALMErwVZNbY/ihYlh6PG
Z4t6FhP4vfDkhWUhKM7sg5xS0++LX/Z8W5rgsHS633/AE4eQx4PYkJCJlNN4eMDSJpXBpJBV+o3X
CnajEuz7P5E6DFCc9oqnlbp8lONQmP/SPWe/Ibcq5C9BWy7SmMe5D1YTRw+x5htGzNVQEzDAebVv
8hGGY3I00CUR5tj9wVbvqpOb101FNQIeRp4AC3P65LzY3REs7r4D6J50cQDMKV2YjEaUkX37C/OH
d9sHABfylulEF1JLcAq2M41C5BjrAzAF7Tv9amPe0w/OKtKg5Gbdkkgj9P8GNlLJqJ5fEMk/htqO
RuO3Sye8BDqe6KseKdS8uJy0g8HS+Bv9pKwPLwNumbjonLWEzVqqJvdJddSv4wGyNUZUlgVrA7NC
bXBbu56oe6W691IdwY6fp9sQpv7m7HtaDUPN9o1+FitaOCoJC5ZKJAP4NdwOB4piJ9BydgjeY2c3
pNeJ00xL8GxphO/Sf5AVzxEleOeHCHMFwIGFuDm1nJQ/19v51RWuQUzAWMDWxf/IzVl/AIjZh2L/
LEm5ku1UU9mBC7gL9QnemZXLi7V7qBJUEIrtuM3d7Ti8zImm5STZ+S5LLOtj11Dz4gnDaBRQMUoC
K0Z0ljc39agakXS6vJd8296ZcAedML8k+q6z81TNVkB1oTZKp0qNxuphInYfdLoMsL2BXD/c4YlF
M/ofUhyVcMfcWj/g7YBm53RKbxx4/2b0XQk89nBXL2KaOFbvnv/gS4m8KzMfEJ+jQES/TMsY0hhV
GRbYFUaZafeExpCSFGqTLOS09LAgk189uPllchcwgMlL9S81OsSxIz5OITCb4SnjYVKVDho0L6o7
ZItKX+PtpZ0+HeWT4eoX7CTNtHIPW+H4AMFFc+jhyO9/0hDHeDd+Nd1tuDX96V/mntnCGsbbUM0W
fU+tfcuvXwk+OFgMv7+LlG4N7joVcpkq/8m7K1fpJRcCP8hvx2Ukh35WCZvX1lbsR9CX82If3Ij6
y7+FTHpQigglqW/ctWXHv7eL9e9YQimPEtmQHXO/+Pew7wW9Ekp8bnuqLEJAfduqlZd/sGy9ilDs
Qvwy+YXkgKfijhHo48QPchP4h6oMekQp3g4XwLnloXuW51pwHqYCBTmF2A4AtHAo5Hfj6LIRILpX
I72Y6cQkEkVd/wqtEAgN7j+j4x1pmNdJNoWK2ga2Tgf55aPD1V2JLChOhF46KMaqvy5jA6DYM3Ub
UYJtjKGIKiJXdg7eLlJ+b6Az5ZvUZPIzyIKOkE/ppRQv7JYiLcw0om615WqIHIm64A+yoWbrRGaC
SOG5ddPmYeWLhDOaJyn2ymv/NNxpr53qTZC8nZmLrgWBXdl0PWdE5oJciUJQ7zPnX/O1/BNmXfGx
BcxI3infLVJ96vCKkha/DTyRDc4pWdvyLid7B0GPERdeQxV0Y4ob5jhtBl1mY2uPSeBtoTIm28Xp
d3XhgRDELo11A40XGdmfrEvHQsY2bN2NKWX11YgNSjWWtRfU7z7QOBvm2twGchEXdxW+o3+1ImEY
GkfJU9RKzqSy3VOuybrvwIlDefQ6i/nQM8jYsgQ+AqQKDBRmfoYOBWrBSm7Rw/siTslpnjL8oX/8
gNu6UCDAyZPI3Sk+4HsJG26YJ88lFIOBkdYcxHHm4zDYWRDrfpdLUT24U+71A6kc6rxIHmfHxQoW
plV6uSXWhtSiwGu+svTtcHdwhKVO8zHxVygFzPGE+4RvE2Si8ff3DLVPBG11QuHSVayjIFl/B9/1
U52IxpNOCjj1JHEPOrrDTIRT6cUQaY1uKB/l9pJm866TSn3EyT69U9QytMxZUEYpsrZX23p+K+Ua
arnuZyBZdN7PhE4eh6MttpIzOdQJBJTlr2Dr/ZtoiKehWpwpwrLjbGjCFBpW3hDXbRi0RDknUajI
HywIrRvVZuTbM4R/zAhe++3ZrFe4uhXBPz2t4gYpZhGhauhh2uidMbyvv9qOHt7NjSA2LytmxaeY
63Sxpy18AOLEQn9e3LB4LH62GEZc2B2vQ5xQuvZsSZnStdaIK1lAvSx7n2Kbi4lYGxzOy1q9U3Ys
SQooQWevTZimB77lqqjkaletkbOGcTPI/VFmzb/AE8XKvEev++TBTy6vq686KT4Zz11HJdVysBDf
Lcpg9TRDBQVAWwgsB4Pmj0rJvP9YX8TQM13oSC18mZ01yLoBTxzygpL/BMGYqHzmX35qStkSkxY7
UeL2KZ6FtVhNksVDvBWBUF+Qb2R606x6uLJQ99xTIB6nd1hnLaQhnFpU6trxxmdkJv6yB30QmCga
DfsHcnFnVu3Bu+1ukJpjBTLmrEfTYS8ZsoUUvfM2JycqT3OJ9DcXK8epxff2yWhvnGC1GPzui6af
6Fd5lxQks/+KRe035TLfV2ltQyu2TfJcmvTValQxiPKcykVPAxND9Jcnr44E3Njg3YbWWg00mUi2
yq0csJfGfeTJkr3zQhnkideDhLho3nyc2oFJWbdAdIjvbEOc1mNLbC+md5WgwJ+8zYMWKawOZ4iI
MOqYaIhqelumUqOFaWwXockxX/r/2/WEXrhNDmBjcMtf01L9UQ0Gzx0gM8HIXrynqmfg++Ax9LCH
T2+6eAxCEyCPAR8yF+FC3p1RnXXUUrtKofzdzsXV+TWZXjTbeCEL7FZNDsbgxhX4rD+197KjC1kR
3NZm7lyS/4RixuobWPP07bg37jywwDTnG9eRZXTziESYU3wVe+cGun+d45hL/gsvkaMR5o0IC5Tz
fF9mcaBVX8rTAWpn9MmqGFP/OBZ4p7nGvemavmj5ljpY+t2BCNYA3CkiNTJ9gGZtReCHACvtv2eQ
82BPEZ/eueYH/72Re7v2VhCSVRMEPFzKnpzmNgTF/76x1tpbVjVxTRSqZdn6yMWu9wws0z7Yybmb
6AvdHeRT9kVL2Eg65059U9Ro7oxW9wYFuyh7p0mjFuVLL8DZXn/fSy+y4dD1oRpVtYlwScKfZ2cq
HpHy83F12KvIpt0hKPUqQ6uCikx7OxYh1yZrafJJXhNBT2KFUwH9t4YcD9/4THqk/XLu9mBhHuvt
uHmge+JXMGUMTC43/k58E2EJMVeHgjUN5PQRoy9wINX+x64tx5oZO5OrTLYd9ucXUkJWoFIPtNvx
9As7wO13u4TtO51mzlicGHZUT6vL3+0qKImi/KnmI/FS5dGowyXai0e0mm8Ipp6TRTR6anS9o2KK
N4xrjf6taEWPQvEaL5YEF+vSwFxiQTUtrPWhtxcblxSOUInYh4rQvOmu0hbyVJXtox2lvG0nLTIV
e65Pnf2ecRUp9RTYfrGOUbJmtnVbPaxT1BUD5ru6NZkPEIq3l81I9OLcvWnhtuJQATBtHWbZU1gS
RxhW1OdwFCKxBaS7uVJT5uaYZhKFSO+W52DG9ya8x5iMlKCOBq8Qc5nddo5yeeUoriL1ZbTDoJ6E
FKbbeNkEC/PEtDpKzxzh+D4QD7vZgwQedQ3pu2hJIIGxHPRkL0s9axNFWCxxZdRJcTTPDaelxaux
RH7a1LnCi7sfknId2kD/4IOGyCMWTxAU3g4qufhRWz2g6ywCtqIDJc/4lzVlxy9Fr5YyT/tKGCKr
ouknx1auf79IKDSsm0Ua64FbRVsMAwGayvIkFoSs5ABLRC58jS68KFtKUt/srFVfdokhyxr32lpK
BNY+DWnyM/1chKbpTMYQy2yUHSyeImjd4czY76Vp4DonVZqc+hb/Cy3zuT0JalwfjZrPKbYpoY0/
sQmqOS9IaQ39eT9woaD7yvE9LyxRSor0q/neMgeH6/bg9riUIdukQSunRGvWYGhkmu93Vi5+SDWO
OKTBpChq/JdehMu65cNyi/l1wHSk+tANA0TANgfpZ8D/cAwrdr6waBc8qgxYbsJrqNGcMpJThOEZ
XALu3Rj3eau9utPauUj6ZlS9EVh5YlkjB0uf0i8yzuTpopj9LoOONVhLDWqUrbMVHCPuYarrZ1CX
w12OaWcIixoPs+hEdgIDGNobUiAEYjJPOkvdykeUuT9WunZmVZKsp/nDbNkpXV0/me+WwRJojMdS
Pg1uE7ms534uJaII9b+COLx+lrGnPnFJ+1BB4TTFbAC1tKK7926cRursnpyLB8oOgcaFWuARgCIe
kfM7LcfXt+yMy9Y7krar+4NDePjfPa2/4lM6mgB68Af5SiyOtyMsn0ib1I2l339XfCOnKdWIdLkK
qZBRTOh+l33lF+qQIrELFGmwSI9M6XHzn4ye87YN4ifH07B/0SpRWZ+fZoZzjjihPJMfnpoKlB8+
KRg/FBxlg73+kxKiEpolnMEEj7R3AeOudYYfwsMA0CheS+zMIjwKJy0Dl3UOxmtIFzwLO3bU1CmO
qCtOF+AUi2G3UC8QhxR3t0IW9heZBFySPpnJBZ4k5g7fLzqObuSCoU2cNtsAcxGmLghhK0B+vno3
ppUvfH7/wntwCaalnisv2SjaznUSPxWoOFiEK/mkxG9JTYuhjpGOC+lmtLdp9LSk38w2oc+vooTm
FAzlt62IATATrnQMZ2PoBklE6SVJAk/bFo3QzBxPTO+g+Q9wwJsHGO7C3Vq06to8XvtBCli0RjXh
Us8MTSNMOxSwLYGs1HYzzP8ZfKQaNsONugsN25zVzdFUlQzSdlrTz2bzUEaos+H05q3D3hyB/Keu
ijBo2zihUWd2pGVozsqOJfs82utjpiI/goEjxBeQ684/Gt+FpvoE+FqBuSsFi0yRDn6qvHnkqrrZ
bSgGyA7KocXx6ymyy+Zic9YuC93vBT2PKNnv4N8SMcIpYNis6NglsZrUET9oN022AR1sQDtOC+YX
fo+GXlXlw8Ps50mGlf3OkS0fenbe1foblkquEqhOA2KEgdSYuD6gyX5p072n4gFJ9BlNKbc3N2+w
rEAXCl72vus0BEvGFw5enN7s8Tt8gGeEkIIgxl6Yhc3MkWS6JaQ5f/SJ+koZz6PNW0x1Dv7riKuE
YrFJcXMQU0vs/FuKbCDlWX1IBgAEwB9P3aKGgfuvogbAmpwTxHqLWsv+/TogKwPQe+9KafwfKOxe
5Vzx0qwjp6whTNjNcyE0n2aKtBp7ZG84zO7ilANCDJI302+EMt5v1qGFyRYTjNwFCghUa+z8//IQ
T0Qb2KM8sTmnH/cIfjXknauHFKNjvsCUH76voQkRy72Kf7p57MkiSHNjtSyeRC206jMH1JOJQKd+
kK0EPmckKwzQ+irHcAom2QSjhcQCLQrc6wimunjs8csAE2vlbePGgQ0ev/4PD5o5aYY76ST0Sg7e
WbVnJ2jgFOPSxsISDcmKBi3VPl+iFllXQt/usTwjeGxJfXoly+nvpAmUZwaUqT+Sx59UMZgCgfWa
D/8IeBv12vmVMGp/3s8WRE5MHDJ0Y7jda6x3Vlt5ZV1CiKYR38V8l1A0wqNI9uTbcf+Tv7reSIFn
wevS1ckEbFS7YsKbtDl4YjSp7lhDG1E4RS8uY92uB/GWl0rmZKbw+vj+HqXZfSD6ncP6jxpAbnsH
Eyv0ikfHTpbQbRBU2uQRtDyE1x7YWlnug3cJcgI3QEdo/qrGUPoMaLdcFvNUepKe9HP5YliTeXCp
5XJWbb+ozuNJVla+QJLVRG4mymtzc9X77j+5dnrzLUja6hb7J5ixTQ0Cc7DqfSO5Feyfz6ohc72V
kcMVkwtarlzv+9R2+6M03W5Q784rcDbPixQ5UZEXYvHKCLVpIfq6qjec1xmlG/+McPy3HJJd74qu
/AcUWHqzUtA7JREzv/dB4cSArqcV59mRlGijwjzjX1B6gVV62Pg5I6e4yBB2SEUSR0P/9NAg2KHE
n8dvIHosy9eadwr8wIK4mp9AxQTGC3ePuNOV3WL512R13nT8bNV2PhHCyGglDQZxZL5mm1QrUZNg
PE9JZWmmsT9tkkhrx2tcNwHk5bFJEKLcfbp9QQHiTVULPWF0hG4P2XgZ82uFKU+wt+BHXRhcXTXy
s1qacgYmnuOB3uDH3nn62rGm3iTVesxF/mTXVNM+cjN/CoMHGL0m6wFopvmwPwzRCSRKIh5SkdsC
5InOtxua7IsrrjqmNLkN76pfYg/F19U+JVha7JFzbc8KW40qwHYxIBezCv1lwn7OJSQ/oFtlNHsD
BuSHiE3HSmbUorj+dHqqrQ8IV4P2rY6fu+LakOvK0XUWRM8qUYfJKUcG44bizjNDBp9TEDSNGV8r
fTlKVzjcHJgLAZUj1yOQsgJZxNvrbdHtT0d/7VDqe6Yyw7gqMgQiie4nIeSm/GPkBOkZR8saaPQn
itdHyB72RO2wVCTrdSTcAM/Rb+AbhkjPfVqQ5acLmpRwLTdDTbtX+XBiyxQcuWyBeUovtpE97JZ+
iUKq4R8b+Xkfme8xpNW5DFkoABcpDi/p68HVAHgAuTxnDJY03CTB4yGDWw0V9a0809ofkOAqt5jg
ba+5LoB7IRZlRL2q/Ro50EcDdpOsajkLV92XNt/zpoQoBnFM/iubleHj1i3lMfsjk5Aedp4ZHziL
zlu25tIKSHJX1dFIWStrkSyAPzRpe4IlvLCwWFDp3Y9+mujLJ0G3Q6HCVB69XxyF88kRo8Y0Nmef
qmj3uLsGMPJ3r/JH3iVNrumLvxWoiomh0Ff1aG3Oru7Suj2CKaUzbOi9HmCyEgGqk+FOGjHsmWeZ
glY9GLmFD8tFw8MwWEllHPcXl30lYVYXiU6g7c5Qwpt58n0K2RJVj8zRM8+pt2MdVdSBZ6aeDvi4
1QkoejBPk3NEY3ix5ZhgUIQgq17Xtl/LSkcn0R9Godvrh832aafH8sF0V+9Bfoo29MRmrGF0wE9Y
6yeoG/GkIaFBTVF9AsofW3tQeumNsZ4GdcccceyZ5PrvzlpzSZ42gZf3cSrXE7c2PTLYwG7FOenG
aQs9ByXTDhsyrDNAbZTEj1EQbsO+bns9gpXNZVmyDxp5k7QZU0Mh4g/r9DH8jbRVe263epdf3F3v
HV5TchaZRmumYWJxhC9hN0RD4GpS6rfvqVonOCANRUx9e0IsfslS3618pYAnjuqnHbqg9bzhPNL+
RTLwEMPlLjMtGpIiOPj740B8XNofO1QiHNR2yr+Qsws7Ik2ZheO/iS5JwATh4StK2LpVePyCs0K8
Wol/EhlbE/Ymgo97+X1C54Cs87dFFHmBtDtgb35FJIZE4elE/oLjeJLjB82tD9H2z1gcbNF08owi
3Qel2WOjEaIsYu55nbEd+6JlA3yMp2koWK17mKnB0cT7jr7Pjn4rwcA2nlCSKfPsPMjOLv902EYo
xije9qKR/MKOg+OLLiqFCo9wSA2GbEjCxmW7Y0z/NamxWfqNTIS5pfckQCXEOj2Ekdbwu3RaGOFw
nBR6Hb6Ss0u0H4JavBudDGBvEX1ovGeQVj87Mhe/V+jSST+Mjnj+HIztx+c140MZrfp+HBd0zvCI
WVcvaV5EwOxntE3pkb5C3Y2eMjOoCJnlCEWIGzXgnTPYnHGXeN5OVLUoeTgCSZ99LqvqaLaoLReF
YrLumHkLXR6N9wCjPnk9aAtVfhaz0rQY1kCeYMv4Rt3TCiPqGqGXuQfB98iAjuY0DiEYPv5SdGz2
69CjkQZufORiNskQERPUSxDu95FOgnhbeCksu5FirhVIotlDtY9cpl8Zz2pggHEbUcIgAlkar9AF
KlXKdFPSilUOw2njO2eQ7ZO06bFHLb/9ml3kLLOKJKMysz2HByvNJZV+AF15rpW8yHgdiCd5BqJz
T6tt2itGPEt8AloJIYA6ONjd1xJ+zJDe0LAl81Jq9DvSNWXrnLFRuq6AHLDyS9pAVkD3y1nRSFnh
xL5+V3l6oQvwAv+K9OhPptQbwo0scCcnfVU8Cg5f0szBcsvH/YG4lCUeoW9biZdvXDyPMiYHaSOG
Ezn6WErhJRv5F2BXgrNx/mOUwSYIHE3OvZtqrWyEHl35OjQmhIBYZ8z2nBBFiY9oHDp5iNLopmtg
kgQk9AayuBJT+lZO/OWSqIYztQ5xFO5zKNqfB+milAySmRje1PcuwwF+rFeMmXEbQvO466FnX7+C
QrjyyxaHV07LbU71cOdvZBmoggAQTBOpYHr90KJIfsmFUZaUaeveXAJ7ueLcKwtiH44d1OJS/Tul
QyaPTl5mg34LrS8KaWcay/j+w2nfS786/mvBokq8tI8JXGRD1g6Xvf8ZCECum9qFoadG50bdMr4p
gcSB4p4gZ8ld/lEM/jmsEcwV0f3saB5l73oRCLBFi3+EWKgu7g3Bujfli4csyG7TgUJSjd2bJ3Ky
sUmwneLsAX3P5lOOEGisVaDLlFuVa3kKNP8Ol/Gw7Amy6NRgUi5pcPXtONFINQ3c/dKSmzwObMTR
sI21FoCCDdh/zqLTWVEKkF0K3STeb9egGUVnWCO/ZUvbb1cLmPYCnsp9RWWatgm1x3oL2VqqKq7R
yv6MG+iRPgUbdZcLw+ZCEwKMYRx79u7TICIpNbgTnb0TLqlQi2+kAMDRuRyI5fiFb8L2nLmbdMvK
YK8hu5nBCSqpZ+hZrGaDiNsKwk6eXIiA9dkxct4wB1lFrX/AVLMcPbWBmcy375+1B7zo+2tVmfZP
qwnRbEALr9PiTBR65jEMENxXabl1ZogNskX6qMiJSYSWlgko4CGsQNv6OPLF4yeVxhvXlUTzhDch
nCv4KBkU8RObfeq2AVu9pOStPEc2uOCME3cWfUT+tMZXOg16Qq7rbkdD3hV2eG2vfaldwGyJCpux
nFNPbO2L7C03rkBR6I3hXJRSYVPyUvq2LaEcHzwsJIMrIfIE0Bmr/r+Zq7n2qOB5DlT2YOKAuNKY
SkpAqgUw3eJDzcF6VLVyzlGWu4RA8eweX9lIliHkbLIfNJxu9JjAX0kCFjqGhi2BhzwJEAC1O197
a//fTi4Im+Y7ze7EHVrWNyc6t96HQpFDqw9uLDem0fL0dzzatDRPrvmuBh14G7oXgsbQ0R3i5eS8
UWe/MD5GfMbhJfkbaYFZ/z5FDP1tr1ZhsZ1gTdaZtKtu0RLh+W8UJSUsSylURYq1zJ5y+1haC9KZ
J4Z/yORExgJnalC0q1ED+yn9p3eT7an2ijLLC8UJeg7SjJQKKvMi5dcvFPqAEmrTNlj8OcGpJoiJ
Hkzv61qc/vL+GTYZXedOhpsYUBBz/Qg96kXUp8zZsUid6I1xzq47v6BYyZHQ53xqZBI1sHH3hWlJ
LtiZltRBoDxn9Lu83dNGrLz3tubuFfygoAT1BMMBl0kEDaVjUCtaTXsiHsKsTo8srCSg0G+/Sp78
peDuWkutp8P9BBXSeT1gmzY9tVGdWZV3+an5iISddYHOWOFj8AG/F/R6ppzHOOcn8hcP9JQqThWt
h7HmU7LpsBtc/8UbZDNMS21CP3fp/oAAEfaoJRHkx2xZV33buskIIT18FeKvS4kziLF4Q6Bgw1/H
JbE5RVEBp8qzc7rxeqKbKgs/+PfMYYu37rpa5XfBYYri16BkihclJ3fP8i0Bmm2HhRSV2QwhUurj
Urg6zh4Rwh5Lqs83jKFLtsWqLuzJOHogyUVWIwCWll3BAGB+Co3CWAXto8blGTDHk4tmsEZLxn85
hBNsIHFH+PT4Jw3IrQ4JDRGFQU93xI4aTQr4qxtXegxetOKdcMSvnAblY9UVWduCHMAgr2lg+GiM
AykdiR2x+enjd32c2aURs+dIhCWY10BAkMDG1NCkOqnNMTdPctCnxMi2oyZYt2kNNRpnEQd1D7nN
SGZd8nc/jT1qahTArsbMOrqbEFvYcL2DFy3QcNNA2FQtrjccPspgLCSU5B26jPo2Cxwb2DKCSisB
2By0r54vKOf1+TaovNSWHgHoCNWvyJK4Y212pyoDKnZAu3ftDHffludt3ZM8/YACv20onn/wZanJ
Izxp5o+Jy+mw5DIi1W8ndSHGq2ZohdwBW12hR5VdL52YEvTg5DUtvs1XslfyoFQQHlFITlK4pu7a
yrmtePoUv7oHZAzchZx/lWGNnkcIxWs/bw51nvDitlkquar5kkTiN4HsYPvwOupd+IsprCeFNj/q
zBmy7UBxUpPIhHVR/lYqdoyVzOExKH7hzk6tstWoWBsjWhi9SvuUbY37HfF9/EsvAOcSO05m2D0+
H/k6cyEEop9R2vBgTYwL4c7g1Lj+RSxDpuNGKVKcbt1SkbU4+J1NJdNPJc3vH1ysbSvN17w67lRR
Z0A4Y1qBrJBkfSnsSWBLkt6QdzrMlwc7TrLHCrt15y2l9yDmUJ4j7RFwpMVIe6RPtntJcyhnxUvC
ju4xuINdvopJHySCCkvtCBeFsHoeT5eZYKDXxtIU7xISZHMVKfRWzNmejM/LHQrLpGIqzn7UiqoQ
PqAesUxiseDMLDaJkC1WvbFR1JOOZ9Ki+r/pDqXoczjIWedZy7Q1dMb7n4fRHENOndNWIO8FjX8q
3Akxf+yD+sLS+a41zUgV4Rr8gPlZlcAYDwJm/68sQm+HTcLrJ8uRfETagr62FktUG96wNJhC3L3X
ixmxJ5BXqkKQs68UKGm6Ym1ODOAIucM6YdB7JC14dpn6pFOinvbMgGVfby5L7/RmkrVER2Efj64h
qUrBaNuF1K4SalP04hsvbEm1JK6Opk8FprOhfMQoNoC4r7Zr+pN50HnZaMvJXARVXes5Fzzh6NPI
X2oNKEGM0AIrWF+JSGPSTSiyRiiOfcWIZUWNgnDHhjZUncVGFQNbMsxRjEZMHv9ekQ91XF1q7npS
GciGxfpx1mPLYHZyNE8poI6aiNk/GgWAeVztAeu4Ia/9fD/9pGgFwfLCddESLmWJPA5UBQvLxUQD
82qoczcyXTpNChCGweT6LL5AJ7xI82YUa8JrT/TDFIssD8wfA3BWNnx8DrXmEfon2rG7AryYqasv
hwTInoaHUiI9HjhJIW94UPUd5wMS7tb8BC/3h5F4D6Og7l5RHs3J45Xqa7g36ACCMgYJk5ZaXLhG
2FK/LyA8tINbzlDp22lpHakkNDfXK6pa4eIxPb/fr4osqLpUq+zVFX+gDj6baK07FPzaFEYjjRiM
JpdUykOnEYHEw70WZ6xQYcDEmiMEhRRNLItKrpssNeZh3uNDlgEFFqwdLYeWcILLBxtfgMEa26P+
nxxZxZK2VKSEvh5SbZKrykL44l6IvvRxgAzvKTvE6NyLJZGnVLYFNliQIMq5um3tig5KFiYjSdir
EibFl4YIfLwAvN+7kHUSg90/xcm0+jZRlobbToWZ0yQFhE/N53OECQhBRifWso9YVGWdwQhy3amF
IUjClr2os078XVUnBV3GyQJwcNpHufDdnw6tfyqjnKm5+dsrOxQn8pGz+PhD9l4hsJln1u1xeAZV
IU1KXJl6Ab8rCBtY/+2N1Sgwg1Y4rHHuFTCivCeQpPG8bK03dONYp1fcClnJjLsorPDRf1moDJs5
JIzmDIZrZcaGYXnBe9fCWoPFAQHFsqU8VgaB3pfdKG0T1M0ZCfg/6BTdyWbW48Jg77OjfyjVrCQl
rEMnJjLo0UoNVDBEItQNYUB7CLCeywvSWK9FYbRCLdmO46ZzwPS1dy3Asy57Ey9GTk46kVTcuiOm
u1nVI5XsZzgg0koGPo/3p7SZ4IxiD4LiqhgX+6Q4l+99u0GbrrTNP/X1ChBUEmZrA/nGwT2b2Blf
MFAlKTvbkYzw3O/RK2eLmM5gUcfaADIe6NBJ91/+U/WylmJLAlf2yxsde9wIkSknw5vmIJKkE6Ny
WlNVSWWgQwS4OIA3f9joJoF6pyY3mLensE6MU/J5dCTyst+DmPqTTdnvPxIuJ3OKjkyxL2Ge5ljo
d7240924iCPckbkjhlPcG3aCFbFIZ0NNJy580xIt7gwCes7DkMJGQHwuho6h2CKOoCUt7u0xbIxJ
q7boX4Z42Z/vJ+Y4UyE430R5Ww08HD9RXGTy5SBEQqeYx/Tg2o0JOwQLc0wZf2lJgogJr1GxttVf
Twg2nLLTmx+eaiIjWeD3CWZ5AqhfgSmUVsM/BF4yCQ5MhXJaLMblJv5EkvEwvHm3j51k2TwuWiEn
HoDMKKce4bGUb0b5iAM28mrIyFAaY7KqrJcmq1ZGmkyaHM9v3zOQggi7NSvPlOsIA6XoQDus7Kyp
iGeQBPH4sOql+LOc4ooQjzvoFpFH3xDmS+D9IIbUekebtait9r+vASMhvUQ1n8ghWrAx6sev8xJ/
GEKl8MRUwys1cbZ+bnJWeGkDKBhLZlt5QZNRATt6XCGUIpU6duIH6/Atooh05luAWOLlSmbdkOuo
AAFpNf4IZ/QQYTQs9ygtGn2+hA5sNYjCIV66gYmYsjXznWJwerVAkUczcbrUz1eqpUp0kbQxhzME
MpJ/Miy/Kmt7P9fpcs4afqX9/q1aInInAO2rtVnC93YhOpspDh8S36NIw9siMwNMUmPlGaNkmmmz
zHfciG7BhLvHDWMUQIq/O5VItq5Obxe66xUgv7ldT82IvX/ktbERuvxyZaRZFsJKqohuLYwmRwj1
2Z0RXlZAnZ/GY7VSV0yw32TiaffpYEKpBPAGOnyFMaOIVN3WnOP3aBovj4O/FhH96fDc+KBr25Ys
2T+aOLf17+w1oYk3MveakpbSjo0ZdqaMXzlAWSyT2seXZ5n/pGaKWzKLP2MjE6eR1kqFX8t3RL3y
7ObZ50af9PN8Q/GjwezQImXRb1S/4tnRH9OsUd08UYnOr1ZAL/tS8OutzwRk3W4/Cvp7Fd/WRAwk
sWWuO1bL71xHYz7T0cwlwMA615/bGUElik8pBAPMgZsXfUjOUqvqUBMs9RcNqngiM5wJFqw8jMPw
wsU7JoNFXSzHyANzcFL01siWtCxsSC86JgOaz/xTum90TDmLKVVmwEXr5NtUvSAVq/ankQdVCn9C
d753We2SGSYlhI5yS3LMGZ0p0sH0iBavMmk0tbI7HuMZx2HY9f3JjFMXslwomOsMh1Ip5guf9IIq
/YkDIK2ZaPHoLrmVNN1/YofrjnU8EE9JY+/p/YC8tcmHrx1q7Ptw1boRDclv81Hy/hr17BMzFl6U
5Gkrj1EjAdI7V3iU2MM5LHDhuyuLho6okk+X78oe7qERSDIvuukSAleOMlos5mvPcCEgyMPkrr/w
DIryN3Oud8LC4g1SxMTASttdYoXHepTqNf7jDAkbdWNCi5qbD7U7OVF7ELqT4832RvFvHOf8GcaH
m+0mPiclRVa1B0zBl2Aih51HxUv/Z/NF/vLsAMhOAMr9HGULWbbYVMuLoG+OeaC5fm7LaeHIJN32
jg/yrACKsAhtFYTKfHmY57HQ94VLrqfe3XSmc+qteye1FH8y3Nyj3amrNIdwvEjBAXs9Ph5O0D4N
vruXZyz59lISLxZ7hOLW5JfUwRKZQD6D4A4dZQVcvfpMul3s/G3OuwZ0cS/rdTEK7oQ8iNBsDOT9
QfXIWXDU6HaH0uCCfhAO34U4qwyL2W1+zJGOpvPtaWtQ/jTS2/YSAGxlVra3CKLtdcNDennx43zp
RPkHqW5TtHRliIs0posGo+VwLo4pYvjr6pbOUDDd0WXFu4MjwNIt+DQvfzmkUZqaq7w9oS+39+Pp
Z69FqDNaCYaJWWsa3yHUXPXa5Z6YABO00HrmZVcc4WU5BVJv/8Fr36r0/+fKznF7z66ZktBd6IGQ
vbYmvsgaEWup6d5zmfRIctKYrOo0WcEIsEDBixaq7c1ABDqmA7ztsc9FEMKcak83s0U1wvkJ4P9m
Vf4l989Ln3gErGZGk5a+yo54HXoeQI7GgBW6hx/1CL4aNhjWBLVTCJX9HGNlnAE3ofdg/OLcqzyB
G/jiVb5lALgWNRvhB1jzeoZkS5z/dW2qCF7fT1VAswTb3G5KuXb0K64spd+zOOct4Ht7/hAE0HcB
wh8CWjETh6SAXKMnuqBQqTccjSlHWvcMm34cQOC3mwltBqkxEYb52Z8vhzU+4WMAMcnIPHHCHJ9H
AwKoXxL51qNPnkepBcxr4SUaIEy2vFhIpudvIlk1JaG/WFwrB3moTRBTFtcDd++4MopAAQHyb4TL
hVCttW8XKYnkztVfjjYfUzmWz1pDSAPxx/rLNhBixolhNqBzm7feYizY0i8D4gK2fajaunKT01lb
OcK4cZQODuL9aB62tDtXiTLgnO7irzN8MYZNTWFC48CB3UnR5aiukHsh4N5qcF5ztPv1W//mN1o0
G/odxMYM8YJNwVcEgUUCiXmxQLWthKG7bXqCekIrAYpxpGVXGTJdbqRvs3q+44sBdJMZcHgb+TD+
6vZPq9RCWHs/CTKebbK0FZgSLkuH3QlTKUXykjUPfyNqTI34eMbcPxjnrdBU12vz7kR+jA+n7Wb0
uqSsuLgjrZD3KJJRwLc9+UMm+yBevtTMk7r435lqlqLmzC8WLWT4ZLYgqi9QE7fs5pdp8xM5c407
AneZU66R/JednGS3PlZrtaLAgOyEbDPWDXWtRTT11Vt8CNSGCC0JXZujqsKv+E5w0fJ63wY9AUz2
hrQTvo8/l5zAViLfyWlqmrHSvF/tilnUZsYLYw4gneO1vXKCah8tIsBYnwewgx3Rk/Bynd+tvjiK
f4+M1qL5UY51ghg00ZFn0iySdUrauCPSvS7la1M4wLBz4mjsgiqZFAzNZYseSGmx/VqV95ROsQZ6
nl7XbihPPldvHVFBgMKHOmchf4tvBhfu5FCHFVtJSgGI8nMzPJ/Nkbwo9HNCH/YIu1PbMNfV/lE3
sCw8RBNyd79Z8VHE+coWSmrRe7oclVDAAsQDh/Mhe//f84e10wubBsTtxDPC/8Bhvck3xbJ2bEZP
16pqXggDlYnM/neQO0Q1M5Hwk5j/6/hRjCur3HSOH3DCSrS5I4YUhqy5Ncf3fGNtdC6ro74jfW67
yt6UQspVBCtveU5IYwvTWzE1SqqKUwAz+1yiuU1qZaE5AU+ZQRdpWDtchXIgLn1Xkl0i0JHsPr51
020LMugIWmtWe07o1RjjYanYe2O+BalEnX98iaqr1vO/WZV04Tqqn4gyQ7/rV2W3BfKZDyZwzHal
XrVxAF26sy99k4S4kI75UdJ/sOxSLu53FLmP9Dq5W+ZJAFFXnvWlblcUEARPFU+blsSEVncbJIsj
e9EUG/OJUPBJsBUGe3LnWnjWkzrFwKUAoY86xcZbGdFkpZaJhS4eyCx+zeFgCI66FR9Xc+G/Rc8E
82FkGfNGVALqmzci3gFphlQ9reueGeEAyLz9fvdrgotTO/a6MWp3XJNS4Y6mKLe47IB4TGMLofTV
2DuWInhhYrrBFqj4VccnfCXr5AVEGyDaLDFQEPJ4qx/lBZN7pugZALlJwSTx6BqiVRWSfseZSYgo
4+HVQx//eimRDGjypfpF6Nh6YgvrDnI06MmbPevAxccg0fyavjogaG/Qa16c+DeAWJrx514zeLpI
FBf9r0TNGJ+HFFJWW+IUfGdUICcgH1in56yVdvPkVpRBrqTdMl+pQF34vR2Tn16VPcPs7B3Uj7ya
LoYB8JWO0+Vi73ESfeYyNpuHW8QzBgJ92Er3u/175Kb7vH5a9lHdcq0Pu3h1zhRfj0n5ouxdFSkm
r6kWGDXnjalrXwHqoXSS7uM46zWzqwkvGiHRYtqE9MoCyIjLBshZWuojQrzqiHNWxZohYA3nD0h0
pGkazhl6fzl8d9z6caZioRCBIAkZem5/pSGK069DxacBV0QFwL0okzOmjBWfZkJriWWUA/9pXy/9
4h+vas/xo6hM1nshDWf4QOjzEK7SJuWg7fiLScLdyxIxQv0DEvtwp7VOInHMXJStWMeCvT+8lP1v
24nVdxTZfKYP8/0Dc8117iMMHVy1tBkHoBHvs9194QWi90V6EZ32F5tzrc+bHaLKdkvIUYNcXB+A
hSHofg2yLQdk02nR7ZCi7v2CbTtDxq2oP7QCeJQNTFYDsXjkLsitelDkyZXotRDB46p8A3leCU4l
5MCWz6lTvqXKIc4WMekSfEDlyHWBVAbdukjBItcArTb1LeOnF+KZIHvC0F2iY4Gef+ObJvjeODsy
pup4KUGWMZo6PNt/aiuAOve6MkQEDkpysamqfld/LjwXfBBzKFGt2E9kLDr4jdcnlpJTCYa5Wm5j
VeaZwL/On9cJX0LbdaUFWtUImFZ0jdCjqR+dENjr1JjDNObNLwUJKhkyHcCubKp1a5g7SBwlydLL
PylDS1qYw+O9uGMgtDRmYSUfe22lwEdoj99b0ydRZVYtYH/zU6rUcB5WfYWtX7XNfacczVUi1mzI
FGc9+njipzPzrNn2mwunSq8jyCP20tzL+f7n+yMspVczfwiMIlvD9jrYb5dC1y28eonG/qK1KBo8
GQNqLGXhL/2Yzr3Arl6pckttMzp/iv4kHhu1wU4qB6WQXWjFcnI0cJpurwHTzwtAHSoARLfnKUZ1
p1ooStrZL+SAy9YU9K5wavWI5nue+zlI7pkZ0VSHwkG888Fc7gizfURymDwUgN1sy3C3ZiRCr76d
XiqzAUYL+VqofeGaNbJC2tQZVAX8EaDUkep3iVBG3McEFsMfTsTsxv10JdYV0aqTLkxCOhI2mM2C
fisshscO4RbZxq5vfcOpG9ofQmJa2BShuTlUmsjyo2EwbDWU1yKfTSDfQLpm0Ym9b1lyt6L62EVJ
6AbTtyfQlHY3WpuxpQX0VydlU5CNeOXEwDdgeriWUZM4VG45TB4631oaHzz+gUkXe4ahvvJy3cp+
zSzKAirdM6osGCA4fNaQSfKX7GLukxBMzniZZZhvnNF5PuwrvGzy4BPZpY4nUsr/IYwxyKuYk1zA
jIl8R2Fk3MWywkFwONq+7+N3zv3Loy9Yi/2oPKijPQbIt4tYzAkpWg3xRFSxYoHGtWdOjgLLIshp
MDfErCS/GvIYg4lVqyXMNcgYlYarmcHJIW7ncij+5H7mrqE0amhg6m117bJQQJOmKnjFd1iysBDY
M940AXxt0o4NJCXWtqtmxpehdSsy4bFdybCRtBsn/kNqJ4rp/y2Me7R8+f8lQfPv3PKpDVWPjmiR
mOXkKDTx7iZuB60q9MoUb1uilBsUiF+xjljDR2i3d2UUImql1foOxmjquDstZC+3a2SBbL7Pozog
fV2ayiWCBtkqGviWFxHJZrygSpHqpKMWc33V2d7vCyGnquhFjEQmzw3EffJsZ8fFBCuQCzf75OMU
p2SvDF7RMBOaA7M+vqukVZ+JrFm6FuyUZtzZJgLYLCgdn32sdfSaF1RGntba2wqEIcXo5bUgGHeN
GvMqi1ayLK0T8KH3xu6nu/XqICSak6ANaC4MOS4SwfXSTZmtM8BY/TZ/AF36LqPQDyfMS+rlCT82
LaBG2P/onjHZwIoiugc6/UYxQ4WPHcXWXjSPprcp9lPpbTymcBM3bDK0WQ/+nHGwqfxZvT+n62t5
Ns6aE1pmME0s/xmfzfAt/P4Q+XF7/ElX6ckOgllrySKn0nfJeRDuLnC1cn0F6iETN4xJY3Oxo2Vq
J6NTFrtGYh9Jge1xGWQJct2G/tat0VvDRgKAb9GypFy9tbRiZKNAlD9QqE90PrJ5pIEkQOtH7vVK
rNjJcMh7Qcy2WygWqeNeyUr2hOTilZuooZksm29MyCXnAOU0OvOfujKOWKynWW/ZJGQKzBoUJ2Aq
SncasxcKcCf2k6SYSrAgyS83dyFvlOqS4qG7Anu8C+hOMn3QCub8wY0tN0DGc8K1fmtW1LdvX80w
73B5m5Ut5Wmydf/5eXX73KvzJ7vqbC4JY/AXQoBeLbQcITPQA81bn4XT4swzVSSDE7qaP2PH5z31
E1XWe7s00gJFzKbHa/p5tCYX+XMSu24o5lhxFoIs2XClcVrr4xeSEbbQpfTJOZ9Ke7xFt+nkT9IQ
kzguOj3tNw/Uq1yd2btfeSahpC593cRgls2mhGp4ZJrlyw6Jjwar3WEZ7aZMwr6pZrEZyeM9j5ZD
LFP57Anmsx2rPD/NkbuG4l6VnkDCtSPNlRwO+0GrdGoduHIrvSqk9eXoRf52je45OIxg50/PzajY
glDoEiYhyv8OOlf7MPwqtKVc3ut3Is2tVKlVRHv1lTwLLGeeC3yL2lDPVBaSyrCGQjSoDnlsxpIB
JsYxVT9vT+5BdK9OjqeZoNayz8QUXzUQ6y+HXPQ6fJSxdLuENgQAZr83lA2BZvd6oxfDpnM9lmPA
cnvXBjUd4YAgeVQuUg7NjKxCvK6eswO5X8HMpHuVRXn0xAcs36hFlbR+BVjIminOtG0g74Xl9VgK
L7yj6niBFcpHXrztixpXtJyQdK9bkyfc0jDsJxxv+gCNXVRW7GCmyHbQEPMD5cXvT5f3uvkFlIeM
MwaCfKUgpn9ceR3JfX0lGlWUDS1ZvNvQVZuqwjvyKBxduBHhhztvAwlWz39IE12TsFWkv1QujZLv
3utIKeZ42gnc97mIkaDZIO30QCnqQk025R34WxtLAH0C/ivmbxwvLLxflhguv9UiisFIQs3UShx6
YH1Jc9vsRLnm7kUp0ssY7XKJWvjNp1vg7tvjslNHQpeliFpZJCK8ZoZ54uuFSMOH62sNSQFe4i1j
TDdKPmJjQmV0ZThgaYcKYepflzmTcHECmx2LSIGCE9dRaDZHScnCPz7qSU++R3Oq9kVXODTQEKL+
8mxpW2NX3O2Vbv6HTR0evb4udxj7CjzWxGAjl9NLMw9vaZlBG0SNoxxXLihewMQB++5wH3EeMqPS
/CKbQDAdAN8BWTqookCH4vvUMzEHVmYrbdO8puPoVnGf8CKfLrnOZ9HQzzuXJuCvcH0JV0M/VWwW
SU0pkYghQ6XGY/4WWW7v3YgoANyv0fC7nROrt936BEQHQkWZcfLpU4FpLBdsJ+bxftXG3QqVf2JZ
3/6uK8vck8CNJDb1hp+yfGlKG3Yqo/iVpRSmqx+uWjg2B1BJBnHdXuG2Sj8VgQv3Sxmax277S99i
Y30wWClDcIYNnYGiOIJEI6EH1Mz9nwDmDTQ/IxuMcBL0Ti5ZpqjluydC9HdFJula7yuezLqZvp7X
Sf0biPnmm4XiFa1fHB3hks4Bh/ZNYGhRVY/vwa5AR5cAFSS7zkyFj9GIogomYV7vL/U4qdzPVeGm
wD9V9N8qOQZdwyo9S96y0dWGfjVB8FfY4guTmbplRHezPg1RI3GvBk8zoxqq6fAnW4VZjEi8Sstd
4Zw1DC24V1aui6B43Gce+NUrJOSgYYEv7AUyfCimz4ipVROGtyarA+s8lldnqbMZZ8hqbtyu0Jcv
dGT6i671MgbVxBASQD4md9sKrQHPbaM7w9JgH6r76KsUBa/5j5LI9CvejdmXFoI79BFoOBx5Urph
ZeaJ4JdyXwmJzXF7gU21HoZte176VQm7oDuGK2fAz5avRTiamSlZgC5Vw2lq/5dca6IAu7ftQgeS
DxztcDca9TEd64B+mXKAVfSFPh+lrHEYPPBlVAa+Clco7DLCDKZt5lIQLhwSL1abSP5Abx0RTBac
sIiIPrxrp7j0PHBWkUXsPZKug6dAfl9ovRRcmKhfSxXWvAY25kadXf1acfhAf0Ho4xYQIj7Fq0OO
PqnUPL+xn0vCz+qVxeZD+e7AOcKaqavZO0gEAcwPnfk2i1D6dO7PEq3gANbL4rBIrtGpeG9edowd
Iy9j18b0yqHZbaAK7gXcbo5BCyjmaAls/ETL4MS+3++hcMRchpIgfLjgi2B+YoOb7lxwEvcgxvNx
jz/iqDNkzYcMZ/WsXU4SjPb90e3YmFQ9dRIK1lm12Zm3pnpdFRNAAiWcGxFYr0EWot4sWokffJJv
jxv/MwAf59Kwb8meQDEJSjqTtNPCvb3Ne+NyNP+RiSbO6wxQSl2rKeYgyPEQdikcKFwTvftPNt7T
EHrnh4YNEFKsP9aZRDk4DmNkFZw1B3J8RnmdcQVZVno02zDln761pmXV5McChULKNxeI06h6oy/y
m2l6nTcIqbuLCvw8WBuLp06O0IkpfVPfnezZ3fxl0zYsaRonoqj3ZSrnpnJHy26Tm9Hw936OAzRW
8l/zSa2+CIqsyLytfslnO3YToO2IN6e7CyYhYIqae34lUdPKGs45sHjVIAiejju/a3gdPS4K+cGK
wRTmdrAIb0q7mqRJkvMZHGVfHOSVulP/hJTnO+7oAj+yk+UsysG9w+HXaLnZYzA+3/P7OQgJQieq
7IAwofoz+DXYylZ/EjEVEJvfiLGV6XcEWIj+Sg81Ch+oyBHGuFPOXzWmKkyc1cYZmKyHBhB0NtKJ
mZoiBc1kBqMmVzEeSa313uFljwK+rS3w6fWkT0FClSjjUbt3m1pkOb2CLWy5wHZjlJA3rFCnA7OH
BtZur6CxlYxUB6cz0TeW0Ik50d5yKwial4hj7Uo4b/hes5jtk/l1q0YLquG1g0qa+iYVLLwz8QpY
CI8XRKa1nj87zzYjZNZiNqe1n2RMcMuNJ/gB8Vu2gjJ87BkQl1zmgApwCiBx7igxld3hvv145glD
EHktV0xWFLW33DTF1ecWE8qyUCvzlYjNaAusP/dqMkcVr/ddjQUGMaY6NreWzroLWhY4s+kXng5W
mbfiZJgorup8XCrkoXdeKkx71ujMVBe4M4HnPnoIc/ARH1Pf6GyNTXUkpR09nni+YpyzfsrbPohX
I/WbreipX7xdryWi/7pYGDyP/M8rOPnsYGLIgUNrzfbU7cPn9VmGlV9xq71NdkEefo+t7xNt29JC
5ADkXsDBJ0lhe54V4TZr/vnMHzxqASghj12ZaA3asmzlGW/3OzfQf+oP9QfH9qLLsrEYuTbxMHPv
pfjrh5AwwXDGbgjga7AuXr3thzTygig65XOG4S02ED6TII0Npa5OCvIqmw4+jkc7ZmmtJXsexNl6
yMWjntl8Qf1MGMJW54jHjwePG5GIhNVQiFuy6M+DHnnJ87LNaw4ONcQB0C9TuQvP8tQvlnoTVBwL
U6Gypo9QurnI9DCttgFe74/aSBAhOXE3jJAnSx/0rw1+KValObFR5b3gkfFgRjuZiBX1u4lKLkVj
mwbYPnvm0wE4IQiXOvOI8SH8Q14rgfd7jLPKW08H9l5TmEUsYOIt2F/4caSbQkjwAKqlsgL6WF26
vTG3tXXgkieRsNzXh11VZudH68X0U3mRMnWY1R80a3wovETr0EHc0R9vM/bG7lvKIXw01pMW+hDF
qskpnV14dU+X2LNomo1Ulz860cKzc6aOQKfk2e4Yz8ccSJW9emMPbOfAAahsYDW+RVnl84u7deA4
WZuk/wD28tYleqObOHAA0mR/wW12cW03naIPTohSb5aKtNY+298dtyw9YnaDYV/jtOweU0jxcF0T
491pEYMeppYVI4KgvYBie5Ih+ehb1leiLwcYcRgsddo8AnPWikxIXnzci3wHiKd4vpgEBHrFpUoE
ZzRxCx2toS4soPRQRJBNd7FJrBo4wK9xPbCsRoOOniBYGxhofJjTr742D2U7OIvr2kbB+p+0ydcL
O0iVnETilT4UYYwwGPKnFhG7IxwSOhpnnX8sv3UljGBOmyPdjQBGNfyrYCu/kEzt0qCTSL3AfPLq
5mWXR29lh3MnuIEb39bHd/4YSi0b6dVlc01tXBSFKpNKE31ayWwXWRFqJJth4MrSMFs/X72x7fVV
nvAEATUjaiIMtxF2g4cMQ+gbDi8ro9XQt82xuxVHlDYt30bbowoJxsWdzgaQEZ1u0YfjpaBg8+Qj
pBal7wsTt5iVFEpmLUdbW7a0wYvGCSHOriJ2zWvad7L36UTytMSAYQEzMkOppLt7K4aLWUYhmxXl
LP4QRYbaztugxBcF/BaACkF4/FkqaFgKf+jn+kQbLAMSQNwqma4KQX0SY9jsCPrPPEUwbafVn9M4
Mr3d/eSQuQoORiJyISax2xUcU0zDE4AJ03b4f50wXHhdR0gjwSYDLdn0cPU8bzDidiflijyMOi+i
+4zqIyzqmYM4EyKjoapAPSb+N/h/HWGSn8XhiBCaAbdB0HKEQVO9dMA2xx88lTvwJ7eAnF/uq8CX
E9IMY6kePk9Otxz1rPR/5sCysf8YZFvEsqsfn9v4DjjF6HsQwuLqsfopJgSprahfpAgeq5Ruy5GR
HuSAxFW78TMW4FK/J8wXntsvoMhQ6izXtiK2PK8svFu2Q4hcE1RCqBqQG1Wcn+8IB6NPT/AegTa8
7wbHVr/cece3H5W+fxZzYFjL79rT2Pdk548fQ1u/jlQOUUKx+PCbO3UsnpcUtWN+6KqO74nTVx0T
rkfdNEno9mcksBwoUWJs/A47Lj4r9Umy9npUWkF6Mo0eOq2NLLzIwRxkKVfwaFEQOFwMEzt/3vUh
JOztcLxC2vjzYu5lp7lyRzUEFif+s/LbcrgTwuxOKgyctDeGhmnfZEOtIxLl/7Cd+4Bn2M+yLdfl
ZorVnYKWFLNCAhUtgodXTfHSHM+oBL1Z+cxGtpRlPqx9wUtABwKhhBwo/b4XqUyv4j58DQVH08YR
qaitDJulyEM/kqUox7OWFpqSXDh1CS5BY2khT0R7NB9rCCR8mcO953Qb4cRjNNJZKbYuMb9c38LF
mokf1xlEje2UEJOiVdzux84Kt2wKqv2tsHntmPyU2UBKH2FBiy0uuM4NHsa5OtW0a1+JcU49sdDF
hgfewZSROTD7q8zpErPTJ32Epry3G2bB50p6YObTgBAr94YEpldlBd/mRhbifJwwlgDz/EJbwhUH
QWPsgJP13E3RQZoGBngyFu6GLm3/2IkhcfZ9rBNBCSNvijcSXFxTVwraN4MSmt+p4itwy5XStdfC
f/kJyid8pnzFJ9c5C4POvfsCuWVa2yP9pQNH0lHcE1vVPzEn8QkiD60GgknscnrqAHdCB/bYfru3
gyurboFvxAc3eihu377HkUoUa1XbNTp7HjcbhZbR2AXKKvkpj2L4sBIxjjBiEF78KzzGxnJWH0cc
6JWQ1ICj1vPIMrFZx90WonBlbfnV9yqmzo3lBr3unq6pJPxmf4ut9fnZoPWH8EHscVMdZD+QUWoY
xsGScRcCSFh4SF0yXi/6ix7zdKzkd3LdAPr5zv1CjRVUNThvTfsghopM1g7Ev4lVtJxbQVez1lL4
QAXjJ+mDJCWt6cDaAXuBdj1MCkzGVO2tydh522XNflQ3bup2cTFdMF4rxuZmwcdkJgt7rc+P/IIt
Br7SzzUXaXg+brs2vECHn+fPbJOYIpOzhKMVoIYXkSh+j/TCgpIfpnt4DAjvpCSBIxng8dgsoZq/
Ce5nX+ETgn2W7Af6wLSZ+4QlIEyL9EK6L4PYjinLN60aWmr4UwP2jh7wpxKHWfPgunckMBBROGZ3
BFTHWmI3ysHG+1NYsFtuO2FqO/GKF1jheYuanJ7yBtVd0SrfAhqz8xekX0LkIw6lxNJKOGSrE4+j
4FDAaFppQw5o1QgB2cYrSqEb35A6cBDkCAQ6VzW+NoOCeRkVJNU2J5iBvTikxs8J37MefzhuRDGh
VAyH0vfYbUqh8O0hi9E7jWLgA1DdG+dFqvGUmtcGd8mMa3nnhy/FRZ8LykKgkOJ/nEyEMywR4t8Y
qb0fyR9LdX3wMdeWhjzmO2dmrtPda97nWvuOjkAp44bQuQb5WdCZFqcjXisPBunAi/qd7hzgCp4c
VFt3bOr3vXX0T0lSJUhUxs8qZiCkPTA3Ukl//crX0mZJ7ZSrbdmapU1WKVEP+0wKrPK1k5JaSY4u
xYe3OMis930wi7MnzPw3nHuIBU4Db/MuHOSXQgW4yBuRt2YEk55CMRqFQYZVUmcbmEqdqnIhi+VA
Vt3e14ndLQd/9zm9JlXu4oiFBo8eId2SwcBra+tG0PhcT81EZl62bhOqqPlIbi+7AYHqbGa59wey
ZI/Ay0Y7CC52SadcA9gdZ820I387su4V4GC93pqQzF4xF4dJI7G+aqmBCh80pm1XMONWl91uGhrT
+SNIbMS8QBIjl17evQt/OuW8SqQHEAm1ywxQSciydsWGXd2TysVaW419amxXBi/F5TLyFm4s07J4
+g2RyHU4G/MRQbwwdss0u/EORnTIIfiPWLvE/pg575F9UbNnydV5rGuHIGATrw18LKQYZr5DguX9
gHYL2LVFaTv15kQwhHxUMs4dqQFh1Htuyj3mXE5ye+s1Yeh7kqyN/YF3St/Et13yOajQCUfEGeq6
+0gQWdvJohD5QXbyIjs1y0ZF9BtDb6esJEbdDws3D/tjapYXmUb0OD7or2cOcgrvs5sYUyK+aB2d
DWG9ZmMfZBtXaiyPe/xSSTtDught2KqQ1yjEoQJdBhB2KEYYufiV1fLOrj8cFZ7+FNNWEBHDXOks
MK+idsayymIA+mpD3pmQ+ejYAlil1GK45Tx+JLqQLtkyBcilCZD3E+3+8PkV7717mChwEs/yPyqh
IkoXDFZwtq8gPepJqNtBXEWsGk/kJl6WuZOes9NBMezcks0XDC0U+aF5LRb2A/i95KF4PoQKSwWC
YGqIcUYAj00P4gkobTLknFVSmIU9Xamwh2zryDGav0L9jABhLcS7bH2lsy2YeqOAuI0eOa8OlBGq
2sxexdg8UPCpwHkDVrVKk5xTofkkh5ZTt3F16Io9+29UF7W/lPpaapcYPzoZSUWz5wpQnonMkiDL
4ryP9lo6KCSot6m7R0zL3xm+UWdTcjLE+2ecbV7FKPBHxAGlZ4kb+PXVIndC92zPFyj/aUu2UmCJ
gi7Zgzb+4HIGGfHm72Vrxr08r49h86NKje/sJmjzzQBGvrFtJbu5YWSlMWqY48Hvu/KRAjieghRT
+YrWfRtMCEpIO+VTGwt7dxFyre5U0MT4gnaoOPdZgLR5WDGPBgP9T8bkZo9bQ5KtL+4dvSPoLT1o
8pU2FUe6wwqrRxyDRndl8yN6pLU9nrH0z80OIrffnU7k5+TPiPQJOixTqUICDiRQrfFx1fasINFT
9AxXqgdpMz71Jl9qY0Eww49Rh9QZ+wgoshYQ1ftON1TSeZy419ZJVnQ6wkpXeyD7YWhtZGkXx5h4
4s8IxZ2eegGSxLGnQANhwzrPpOplA5RgbH4GaNt/mx8FrK40YCBKv86Ei6Mph3B6d6NBWcW7/LZ6
RJtcTQykMQ5jq3w9K6Meo2dG3T3AtPKx8xfendYJTBDEZSL39h4nYaLM11qhAvJyTjUmxnLPSIn8
OQ++trPgF/ne2raOCPbKzGypaS5V4dqvpnBGaXqyVuuXxRdosMD92pNdkfV0y42Hay/EdNVn/VvD
Ti21I3g1G0maPQybsQ/Qm+WqWx/mImWaGCxMlrdGcqxmHlLpbFir6ZjnBWK0i7vNCwZfD8nKolsU
kfe/gkZd/CcLTasAj+5R3+v8BkL7e7iMxZMHd1zwMwtV3LPYj95RTawnFaKuI36+yHyKqHvQcxIj
dhxZANmo60nnm9NBESwmfZOMURx/gfMAxyOgG+LJcv1YK5+uphf34FgcwRzEnbkxieE5cs2nIoMJ
Ml4Sb7Ioyi8WHxDeL62rzHGR96OK7IZ6LyS9fTxwlWhZOQOPQDArgOZjEtB9lB5Sl8PMVHqKfUbu
V+QjYuotJnhJ3fMAtVpv+3cNYxFdbHMvAo16zG8J4l+FIr02M1rYMjVvlxLn5gSHV2oLpLNqdCJs
1k2WVOBgqnAqrHqtDU9eqGAXKh7nspoOff9ALT+3hJk//hkVp4p4R/fm6mCt3MpUX7AU0peQ0dyp
Lyer0x+2ZH1ibh234NweP1tkCd/YoDFdMeaMN/a6/UEZjQKHuqHzPI4eBbxfxZOYNjwQ51oBu0RQ
8OdLHVECSgBmnjKRP0wioB4XAwiy1hxgDaH+1cIUupQNpTKhMRDjaf8LMnsLO8f4z14y8ljvMKCf
ONRSaU0JAFnmSLJcmAln0sm2ckI2w0JX0j2CtUiXp6lo3i+O2Z94oFAG4N8T/LcrKB1VJ+A9vBHS
tXxxhlL70QalehNLKmwymro/bS3VIyvdkiwuuEyPtEDIFU54hYe0B/CEldLrFIVoyYfpDjyXZ0Nj
hbEDDsXdJA0bt6qDy8sHNqioOj8fw/9HRkw0M6CzZPeSkDD2+Q9Wsz4inODx8UFzQ/0eSwzHfdbU
pMBZL+KDEi4xjRLD451SHBr+RNH1Nd2ht+yi8/YzQd/0dZ444G2z8TJswT1NODTUByky8doq3xxm
xD822ZJsQQaxlMRRDb+SWOAN+SkiABDseuWjxdcw/qJTZLEZJfhM38Fa5yXD/tgxKRQFb0D3snAT
UFZzrfGf0g5zju3xA/4tDF2LaAsNrg3zAkrzpbpQA/J9HYVAyzeSW8vBk5/d7MufcT8uYVx6ZUZY
hzjdiWR90pkWQGKVN70njXl1u13Jsq/14Aebo51ld+0Fa1K9sQHy87ZG8TMFzkr9QSpDXss3liGr
+rq1BLqS1u/60ShJ5IhD7ePjfBP36G8QK2KFBcZVCEqe0XSOuWdQng9KptmOLhI83NN5qXa/P1Eu
vAItbGZs60ozdWGTg8BN4aACr1NyVav7IX3WhCV9htAWAHJJEJu5p/6HXHitbx23wTg2IXAaP3wD
agHvUM0Y50i/uTUMP8C7RWD0jD9uZuqlxoc+nPz6DEU26XQC+dOcTs3K2Iv7ReIjRaUKIvMJMT/t
wycBCIq/vSK8iB6OEC/h5vR380tfYdsD9PbVv1kX1OJt6QkBnW6hpvGyVC4Ak9KWojVjxXxopQ6D
+PH1PS/BXHoD+vkUy8vmZmrXTKNsR6bmqqDcujFd6zH9OFxTTo6jd7fo/5UVX+t6qOCy1e0lj0OP
wGtkVECe/a9wW/va4dskmllQ8jNOGHSHAz2Qw3rF3KcVOkBiy0XRiC5fVRuZrNn3nKfpWO5+hcOv
fz3wP6n+qlJ9FohznlOyd5dG/ktUcE5KM6aem5I/9nIFWJygYOJzAKM0r/IkbCf4+QkQOkF/tJcl
xwoHKVh1Cth6pzXzLdQwd0N3S16iQAj6IO4plPTBLT+Oh98d6NbY8eO2KxYdx2JT+zitcguCnUXe
ZSiYOXc0gyFwYjxNmPt3chxa/Jxw0NgLLcQ2bRP04kqhASfl/W88ovevPs6yc/RD2YEiLu9+Pv7A
JXnJ8dK/aR8KY47nOjdJ11aDYq5LLF3DYzk1rhAPDeZ6Y3V4dAtkKePwugLjUQxX8tTbo0E3kEkM
dLHKBQQljvaqoOoL+vteUBMKOf7aduUZMuRhMa94RnppsJbtWWWCqyjxu+OEWG8vSCYbc6QE9qCG
yLrjtPacov36jpNmy8MOm/JbWFzOyy5ZkKRWJqnC2RFY7Y27PXNyb061+2ILXkIUWVYSEZRc+93a
kxuvJA5owrlOVfQab9/JK+MA44aGWY7bQRp04o+tsPvUTB+Atajhy5JKOPnZ5REvnaq2XH2vzvsW
aaR6EVe4Me4UmuYxLI6JiqUfvKzC6UTQeKGTSErJ9ePa2cKXjth0b4wEQhDkRbVIxDg7AOlLTCoR
4fkAgmHO4snOTSEXEhCRxfE5MUMiiY2F+vzEOrmVN/uZdfFtBX3s0O9CgPXArflXigLi0VcQVZsI
CYP3E/qUsENlI8YpO9/8EenwPMWb5y1wsnyXc9fgyD0hclUsp3DyZQNDgzzqPUG1rQ9ZHEySatI5
JtMA+MO51hXIAZ60yyzAgrR68s1U2Bc2fwukSMuiyJcwBS4aMCqI5z0BnqVdKfuGkQvA/TpBAl2+
69Pcq12+jWZEcpxFvHehBRIlvCFNPWxXtVOSqSdoGPR2EwDlenNdd+ZckfQFxl2xlezzupMVB0vi
maWwJ1aY1VUlImgH30exAel8nEgQjTZO0/vMfyiE7IfMR5Bb/ZtnCjaC9e7WSwmqHO1AINric6Ku
oiLtBJfzJGVCuKvmdkrUN/0JYmadSKxcTvwUytw44i4Zkv5u/uIRfhZBWUmlL1hH+VS2SdZhe4Hf
Kh3MbNFbPXzZBN2BKEgs4IsjiqHAbE7mTHjPQmClrZBpzFSLVeSLq5FUwymnfbu4in92ZfnHixmm
ehdTecV3GPCoaUaZhSiGRCvzuYVBKyd5wMQKQgFlc1DrO+gJMXUUAhEhmjkOPtPAInofI98M7Hpe
i5wnOdJTpklIJMrs6Vge8T7ZMKW+osThhCw5GLeAVH1lN0k+XmNGLHuMAn9KIq0zBkdpveL7DjwR
dPkr1+kwfsweZ+h/fszmL13Dnt6OMf95L4Rm0VSOQoRYMKFuHANvkCMB07u/JlCiX7QBYo3suIhD
6RpeMjZ9Zd1BoBSD/WLOYvybM36EWcCmy7Mqcx4GADbFTjTroHiqaddf7AM9UrBik6KH/ZV0YOo4
1XOw28LJx2EYos4oPge8Y8pGhZbGkK1Ia0RC0ANzyJO+6Nf8joJPZHkIMEh0vr7cVoU6nwq7KLqJ
rMG2bpcQbgB73mejYV79XNkUM00tyfT9bh8vkXWbV+fQ0OP8ulbhDwQ9YGM/grPnWYoYsxDJkDBf
Ay5pCFVw3160BYZWZC2OVuZdKwaPodcgdPQV/1FtYQ6OmVPCx/lugQTQienTJrQlcD6IyEsLpIGy
FnY3O301KwiQjlfYHz2DXETrXCCuRJesrM307jNjgd/HOI633k+Odc/fRmTRnVsksxdhRG1d9TO3
cqwLEKe0QcRQY+js/wtU4Q/WPgtrWl2CH+Z7d124XESkO40sot2UcDFWkRijzqd/sFBRXZd5YehE
A2OA1EOtv0gxxdmZvSZXryorWJS7OF/eieGn/yuSu+29ElDyhan91iupCJAbSIVlx5GiVvey5XnF
kvdKP54JIS8NHciw8GpkFD1UgByltYOtdjuf70RQExEsKx9yyzY+fWM2uiEGqaHFGI1ia7UneWJ0
EEp+CEcyivkjf8MbFWNWkos/MpaRuhNMuKbXSXvKQ+0XaLON8N27eV9TaAu+sn+VPddGfySn108D
PotC9qp0PJmzvxdvid8uBRNkqtAWwVmJ1Kpei10ssy9j9aBDTqaQMOivEaW9sTHPwHcQ47xpxDvR
kEd7Eb4RDioHQshZ7pYlQ1IJznU24grIWeKY+pEGxkfDbpJfSX4fuqaFf5djc3vExAEZKmQuafk5
zF+/Ybm0Is1AQvr2N23/HI97f4VAS4aqq9ukWVc7UXZpjPjBttcasHZRvT+1TYqqQ4jSpFLE4AOJ
WM6gURReM/s0Hy7FZ4jPOEPPlkAyZAYeXn+c+2s+HkEC4qx4GtAQzB6bIXmUUinWtrxQiPidcAFm
ZqVLGHucfo6uDBdTOrG4lBMCnfMxyaHkY1tcgL+QB3UrT+IAQAZF4nrhwEFBpAEJ3zjDypfjqBOE
1Yw0s/SX5QOI9zlBAs4gTa5J725jhxs8pgVY00nRKYILZN2V/1IgmmqRQa35zGmmBbE2920hj/An
0pvR5PJLPwjHOFnVxI8v1zh7m3P8EB4Om/7G0o3VfdgsFRpV3uo4cU1hJq1qGCe0YNx1MSyMe7YG
Ru0hOfpU7B57FrkZtNMRlOH8gNdFvTxmdC13NIOOpCyyrN9s6sNckfqT00s4M/akdG3N8P9tVezZ
Bgln1WQ1ocPhbKfqKoOqwyigYf+RdIpisxfXtQwLLoa+1p6tLeT7Ua+VlNRGOZxY3JcWpPGX7xcm
oy7e2oD5N87RFMkwfqMrudtypOH/Rc0mXS6j/yJf6jEBm4Z//p6z+F92RXXdLYgEutwgyQ0HgM9L
y7Fo1EJGZ6tbiU+7J9N6Gc0QLeq1P5ajbzc8cZYSPVI5qOwZCpnBv86kEKRNmkAQxkuT6mQxUELg
dPEnsH/ousgVlPwEux3azF6NiLwoLh8+3sXjzvb5coGgkMvBzmQwAbcr3JIvZmC0Lm6WRj2DfcTH
qNKqZM7FW5r6U2a+vlh0e3fO5nTud0e7+VB5nz/GxoRfarPisY5tTsrrsLAfbcs1l2/Fa/jwCQMJ
lku6pXNgAH/mYyW0w7ol5UCMqugrZDpdQ2eGqaJlsp0wq/FdkeQxWgvRGZMvl/eL5XwktZ2+zVZw
Ey7UgqLcYGAowbnrqNjTxDzYJe/WFshk4z+/5R0VK/w0++aq3JV9BrRnaozB/33rAzoLAjOSqZTX
GKiLcDG2/SnlOqJ9vRHMkZ+DLqzK4vRU2O1sIjKkVKuT/VafISdy4zTrMrn0IpWDwz1xaUjq0zRV
MCH5lrGyRoU/N2u/khgbMm9n3Xz786fXGhvF6eULJtj56q2yDBAu6uSUuQk/FhSS7vIO9BeDDQTU
1OuauzeqJf86EiI+KGqfR96o6Epo6L/PMHvrD3GJipGVt4XVQBS+q8x3/cR97d+dzh+NVf/Fts28
NxFV7pVLAAjZ501QZuGyIXaK5GC8BYkDafryAW5MAKf4+8f/02Yydh+VGPxGyZBfG5LN0NYzOyva
1Czh1VhVGFnaaa7qFC7f47Bp9DGJ+qvKRYi01XK6HdPoiKtnmcCt6QyFqUBVD6yAqoZYZAzJs4yp
/nosD4SNQe7NL+18x6AW773rQJikaZG1XQqtExnz23R+Z/ix7I0TwlThQF7jQgUNKF30V4nTZq/x
BComhD0ozmYyaMwyUzfdC4b76iVkZAuMaiE9LyiTwqxoNVWwfa4Beg8BzwHzW8c6LyMgEnd6M0LX
Q9l+K2mcFPVqBU4Kn9ukABSq0zx3JYtd9FgKSnjsQDK1ONsX4zVCzCoP/sNpgQpxDcVsbOlZ9XGl
Nyfc86zd8jW5+gohp7FpxLoV2T1wHKMLWA46DYnprTkOJigqpcykEZJg/5bWq+35QWRHI4nl5kG8
jIKlpN6G9wkzTYtRQyDkNToZrWYnpWJHZdM0fhYNocUMRgITxSlUS48o4PWeeFLk0C4OlHiIE+x+
/avbWbWl/P7UPynzb6qemmDPMa1N8Iea+nfISspeVOQ3x1axN5PL3o3cI10TZgvCb2/S0CZWXUt9
iJ02zGUKUtVo+5qmxspRqz1fTxtbQDRmszAtR62quAUXx7YW91ZEWK7+C/jcycu2B/XQFt80N8DL
aTxWwkGYaxSdp+svAxH80e8dr4PVBpy6AoK/Ny9fxLzwh7Yo0j5g3tEjxZ4AbP+EMKeYupwwkGxI
z/0fDLYnh3EJ363iyXaZmXbYaIUlH/ncgz0NQ1b+tZV9MgEgzy1s4U89TAKVEYd2ExwkKUQO7IVV
dlo+49IDYQHTdGVePkd++C9XjAXmbSEEtIn8wEr/zie+2TfqHVmWEIziEQDiCPZjmH1HktbwvTLT
2OPEovI9iuK2jIomHTv608U7PQ8AuXQgGwkvjXdhZN0a2Pln0oaJr6pAZqA0Xe5BEnCWssCAr4dl
DJu5fBaREiqXFduk11SENaJw87KkAL1mKiUpl37e7h0ZZsXlO4z+cq7iS3v6e9m0x+SzsM9IvlSE
gKIh/1OXDWQFS3DirYCGec1RNXqay//9rJqKmL1TjXf/o1oLemu8+k4HDSqbHqmu5dyo/TeVu4NF
Y5t2MtWYODmF9mDdNWmYuqzXn6kDArKNRb2dFt85kOzDsnpPzZcvtxSea2cg1zuo/+GhBvQB/A0G
XnLYBHx9j3hLyP3KFpgYWoeKBI3irEUBbbLrvprRuKCcxAxHiQdcRhd3HrsAylErJ8zVttqYSgyw
TXXrjH996JBRxgczCj888JpnKMFWOSA+xrh3PvRT6gfy2p2i9l9k1ZcOJC/ij521gRLA0+GoUe9m
vgxQA5um1rw/BAuQDaGuzQoTRk2+PBuskK8Euv4FV2rM7uxNFbC1aZUPsbUzF94hinbKAXUimpGG
j/+PNxHlg/CUa2AXrOlP1iFr7IkguAasqSYfUo7M0dpqiUM9v74lKBUF6QsmCbLoCnc02ECVAdV8
dJ/ESOVPJMn2lfdQiFHx547t4icUt7Lu3ZHqFymV9x/EiNRn525vL4w3ro/TsouY1vH16IeAQQa/
/O5KC2KG5tXaj4kBLoWV6Ef1pQRfaabVPuHJQaO3z2wtobPdK881YElxu6AshbH6W1WEGCL4lynf
AAdok9FXBGwde8LcajuYv/zEThW8Uj67ISlh1LFIVVNsVP6B5G1bnrNj3zvLF23lcvQ3cP5JzLxQ
tK5ZZPHNDwIyhhDyaufEFX9qSYdH/X55/Y0oGxjYLo6p0H0QPOyYyQicmGPpIhTcSeQVPy51VDep
kKgmoHPlAiPW2h39femeYb9QZ4Zx8F4mShtdtvTfdxxC6bKf3AQp4GADaufVHDOTtLIniBrCMq1g
6mms0NDtvaGixdmNKdtWit7j9oqsLlnyGwcPcf6EZbteGs00o6i0ttNhbrkbMRb/f/m4LCBFIhel
lSeOYP2ftPfOIR4+GkZKrFLAKkegOUiLH2rH7iXnMNW3ei2NPPO2zfBrvDvs7TtF5j4Imk9ASwzl
4Czy5tfJy78d5iW0BLTOMtOb266i2VZtPtHGZmc9a+zNJYU6j86sxlwNvbC86nJFyUIcjLT0bQKX
CxDP9kZot+HJJFr8MZDAojMX7UnXB2E4qkLpjepapPOrrzECsP1qqhl4Dz6DmuesvuZAsnYuexTB
r9x5sLIpgnkjF4/lxUwK+7iN2tmqbsqPOZSTaL+btLSYz36lvsmAudbSB99dlYMmAhyzlbQ6CNyf
2CpvapQWGQUtq6hH1EOVqUKAeBsB47cDqW8SZzkK8R+3ATXPkPFb3hTj85YHfvN3XoMuB8yGhsWm
4EIQRGnNZ9ZZ27MxdrD9I6jiuC3jTaAsOImC0xpSDYkRYPE8jaDbJ2PgVjpWKKxM1hbxlCu11X05
fVou2lvAdwFHaLrtSVPOw+EJqryssAeLJSOA2B8zQboBmxNwDqWVRzT+NUjqi3RmCwxKkTFf6zvd
gmegrs0cuHN59oZTM/9Pfhd/hJdfnkxTIZKlksPF6JZUdFC+Ec/gsZkTME/rqjaiHPuDbiKqY+5c
1Zb1QC8FaUPmJyzS6aThq+uIw3eHSkxvbl+rRyMaGGJ+0UaHtfX4HemX8Ihfq7S7K6hBhj3Rob+B
awgHI8bbFYhjzTPGNHAF3v2h0FcR8ECg7Nf2WPCQL+5kX92OzaK31y14jRgtbd+nKrWnfMr2Hc5A
OJtgfP2QX8nrC+RsSZ4jaVHSVYNpPbn90vUzMzpqdpqj3pcTDvhbcH5rsSUCR4F8Qak0nt3S9dwo
WjMebd+wrqN7GLt8rU7E++9/eruVeJgzAQNgbDbVTPuar9tTCeBf/ltSxlw6eQmNy6RC44wU1Fza
IeGTdjQQumQzUsRjbn15UAqMJoPLVk2NMwgLd6nekIiMm7W/GfzTtEBNh4LMbuBuyqErmcnHeI2j
IxxKPiIC170qJMj4aU/p6nFPEwQ6YTq0BONRBT8dbRmvnn8f+ikfao1hE2gLfAb/Ugq12R0sIs1p
a1SRFqv3wmiCPlPh5aHmGDwN5das63RkdG7kJNnYLA8w3vzHSl0rLFkhtPw78Rlw3j1Uzc6Ohe0b
KbqcfSB39f85nHeFMmG8NRSzRcA+FzaTGV76FtQWiLXQjyAX0e39p0/lBgwrOb8qtWKIYzYlDtbr
YZiI2dFbL14bkdq5M3cvB6NWZoj41Gd22P0aFQTPic0d6VKGh9HtBmmDrUGwHVnNxIN0OTSfwSdg
CF7GUW/Ci/Y3mWXVDpRg3i96Rx0SfTWURH98l8pYX7RM4b6NjnIRyh9XfzpMJ9vVdaRmA0QmYCi+
VEW736iIxPJ5+hMYwJDLEEbdGDsRlacy4rZY2tktKZN1Ntwmt6v4H50Ts9fDxmb6LyoKeVqMnENu
8wwGScgrAsmwL8wVcmS6GA7WW8oZEPhXFZoON0WR+RPin0T2A9E305oxKgpR7ZDJyAVNefYIKnH3
RyQs+9I0VLs9K/ml5vuvt2ztHMAQwp2PqyJRi57+iVkvMtsngAn5FbY5GDUC1itEUvLd73c8lu2Y
aZ9TTh+UW031LRiCt/jnjxy+t2Ajt3xI6K4S8B7LVzEsMZwg+v7tL/a+Oqk3JOU/qOfqtgrAkP7d
1rGYikrVtHntJMK3HbeO4t97S7yDCTh8KbxOcgc9atoGFuBnPTiGHDzYVpyQU2hnuvRBvxhVKaKz
SyZy6LFnpHRMmyeNGxDLJDWQrshem7UGpBtWuczxTAIz2nsNpwQCKifgQC/DaNptbQX3L1KM7GXM
OirV0nTznxrr0Bo+eR7FASZSce/0GXhOXo38e6ZoDl3kQG4DrO5U2ZQ1a+Vu7tmmlPIE4tUukklb
As6TPj72L+/aByrMZvs5dOGeLIEatu2bvlDe5tB6GW2WBQsIZAIjUQPVOhKLwxzBi3FhLU36VWbR
/gJQyGLLXmZtlWW452IJNNImdQ0KjIwyYtWNOe3b4qR52hm4rImTku66w5jWX1ftgxF46dz0KVzK
hpd2iozJya0/C6hfq1SB2TxxGHMxZ1eqXtLk8pHjKikzRyRdb7Q9ZnBjj2USvtgOU5mthafg52CS
7lpj7gnDiIf5p7mAN/KwQ+A+mRj2cHnFLuuYITYZz/u+f2X8Jqdjlf7FLSqLOhfJ3NA5g+x4EOt3
0ulyt6y18qqtspBkQGdwUiIPCNxpKuhx4LcaYvbgqxARQvyi071jPCLl6sSAnrgSuGgWp3tOPHiM
/L1/Jxj0I6JepwEMfYsNpulFDv2lTdjeCjA6nCe31NSFBinzy22JdcmQDADSNakxpMlisw0v0QdX
GpvOkE1AAQc/gUNFyu7Y4Rwjpy2whv9HNM7WIfWMiFwT2fEjn6VWP+z9Y+myBhII528XFklRMwbE
+f3d9uQ15EvmS3ozrrEDDKEXObrSdkgwfm+YQbqZDhIKGWuFlHnh1eBjKIDB3+3vRcRGqpfOKbm9
2ku7TcKkhck9/hQ8rMQ4EqD1M8QWnF8kJyBEZCBU5PG944vRDSmn7V2ZcDH587980Sl7Puo/GODA
9x4o7C8UcXzoqlzt+X2LhxktzLPbCSeAbQo985cxrFLNZpAYPiUVjEyTLkJwvOTM1/NYoSfKn2kE
3MB1dY90gZkyN91P7ZjBc5mn6bGsxEO3YkAc5jKu7Uh6aITfM/ZBCgCK9onV5wypfk3DIpyaenWP
ETTEKBPBQ9Vbyo/SjHusgMrfSGSLBY0+TqIfHKNuuuFkfi6q17dsL4bShMjJh+HD/yWMokax2SXq
X3htnPznDbIQIvv1d+pc3RGxPmAfevHkbhpgU4CPvnCSJgAn9R7wuu72lF5v/I5taKu0g/lstSti
JxdqwR6hvSIPfO0dzvUXWEiYUO81GsKz9cutVLB8KRuvQznPGOcmHO5BiY1tMEfKjim46WXi4sjB
SOHj3uvMqllOPbjkw1K8nUEWod1vv2uhcd5UIXOwQePDOs6OIxZcIz+Xb5RgvyT9g5r68AZeHEg9
k4UFwLB4aZtepFrlaMSsl0QmRoiLBjJTHX64Xei8NeX40+A/J1vBqdB2IKsbNpRlTCSTEjJXFjgw
HHcejpHXGy5RqKgZsspr8r4lGaMnH2AJUPYxZlBxeLa7Ob/877NTeQcykjnR5kCO04CqHzFBEpJk
1OIm/gfqrJ+o6V21sqK5PcDpR5vXv+Pbr/nDCfWRrJRd9l0AAYnzxdNBztfMDHPVUsBE/sQgxGHi
6g6mK4X+PGvV9uzl3AwWk/WsPSVPr8EKFF1bY+Bnc+MlzyYlfPHubXuv0bKt0i2lE6dfqxD5nxMj
ypaYexvsMi2Oqb5Ml2i2Hp39tBInALeD6SbUj9rW715MJ/Q1OvAlgmrgX1dM22TCSPwRCUCqD3RS
8UJG0DXUI7JozdytDcldUKBj7gqdeuVGKtg2PnAxdwDqvV9rc2PPb19asw5mKYDhpt8DfajZdjvX
2NGQO29r6vsGUzBfSYJfDISF1gbULOWMphFW1Jo0UBl4b4NwudkyEOgqHpSS9LKHUVy6SCddQ4+Y
iUxqt7BNZR8DMSGZh2skOil1q2zaN8i/p7upoIi+/I63ew0/06sSyGUPg0pbYbjzT3sV9EjcT1Ld
UWYgymWEiIm0CV3aSGwBhSg5QJEWchasF7leSZxgYf03I0rsm80+8dMAFazylniFkUS9sE3f7EMG
SDC6YkyiBqePGWiZ4qkYL0s/Kp9j0XbMZ+v7zKtivrZhfuJ4RhqPXA4zMuDmahRbYh/NZXZMiRRK
nNjmbztY6F+aaOL/6ETo2Hv12k3qzeGEtuA13BF6qs4rIj/iHAVSXo5jsiQdpC2EzFQG+LaK/sUs
rUSrKPIY+rz+gQNWy7H+ku2CvVQnw7+foJBWox5dAH0k/HO5kYE5ripOles7+Mg9Bp54NMAt07m2
6iXSqxpDmYkhpeUc3Eczmq21lF4m432zt1rWya3OoC5CYfrhKAdOSlYqgtT/aC7/eYGlGGnNThew
cmpTO1dNFwZOdLSoUIquCL6RP2G0gk90hSN2Mo25aZ70upT7e1r/W12SlCLZ5kVdESeJV6GyfhWy
axAHvXkMfx4Blo38FAVQ7bd2+t1KscBG5L7uHKIBekd4dLDW3XIisGDbGlz6ikMSJd5tMVL1qI2X
6ZFxMEziY7U+Mjjgzx70Dj8dZd9Z2S1FD6x6RXJJ0iVxL2cZS3gT0hjOkeMHZDpq/mUWZaY3/WWF
vbJ7VFzSNuvZBozdOKbjRBP76zKbew9gnoEODloakfylwupsrQhRXd8fT5uok48EQOyNt1D4s2vY
tIV0mX5l+YEJ55Kiz5r3/39i7RtNiZB9RUZu/0fUx45cx5vRfQTDFMdowhqks51+vY0Ze6C7f9/r
tlqOSCjPZ4Vb8b1zfl1VI/srHfcebjNcgkMGxvgaYOuwdjmUOJAxY4gz75lBHc91H+7eK66kk8VB
hrDfkuRlrCl4kaQ1XfmUXpns790kvTnpHQSKv580X00GkeFyzKkxrd6UXq5E6ibcBEnJVJGwg0vU
8DMhtHiix3+EO84xNCGHZNlJTinbQvEa/oiQVIxILRUXQHhOVZkLJQ6NOOT60WgjS5yGWsjd88K5
sb/pPbiX60iM9OHKMLFJDbTqUN98+5jU7d9VEI5kW/XSyq1b0nJ9ghBNQ/IBa13jlAQAt/wWwLDR
jwX2/mOqKOeGv7/o23o0zU667uihT7ccwWKs0uozcHrTJ+dhaoP40qkOimhYf/uEntOt2ciZZEHv
ByGKgFHibvpJlLseC2xey53jt1KWcLij2pp5wCjOhGPIsYY7jDST5DxsuV2jRRZ1qunEeXH+WKMp
8v78tgg3PeNTS5Y9qD2LDCVAFbI8Hffn13eOV4uUGvjMJoWUBtksQyHue+j2e07AFkEajAQCnwtg
scqq6N3Fzq8Bm8p/E+uLIILlp2byluvQBeax6GeVbMF28zw8oUJR4SEeszO5zY57WIvHHSdfkGFO
GHVQVHeXYBKehXm2A287vnk7La11JL8L1FHsqIJsZ/Dw9mOzFJNL8yCtLfolS1EXUc1RBrq9YKLt
Wt6cAY5xW1Vf3CxWICJGvhgRmLERAW9uM24WG3cIjAF0lq6zkBfiGfY1/gFHl0yo+P+qxVhCWCbi
f9R0uBm8m2dfaApW3Iz05/f3Iy1NzIxoKePo9Y9wcPQAqEL3E//QrPR7++19rB2s986rzlkw+w5z
XAKfG1PJnJAcYiN/8naVjMUINojsvQHm1u+AhqS2un78sx+Bz9god/oN4uuQwj3aP5WKtGugYULm
ELPzP9MOVVfQvPaJG1SrFII67pCy2wFcUaARLtiGjOQXuwEhJbuODHBqQFFJOGHp1gPciY9I7Ybo
/IPEKDSASqs8NxtOS56vLiIyp1U7T2cRwyaNSMe+VOIQU2dqvWQM4sU0LJqtd0fHpHCgZPii4ejx
knuQiyY0CfJ9io7MWZxL21LTCjCrlre6vU1fvD5Kyhu6qYsNFAOQco70BuoRuXMSCbycoF0sDKk1
pELPXjZrym8D/3BtaH3RRlhCLOGpQ/A3zShY0W9Yz13zYo2IGwKsbapS1d8jREz7r1IKKnOx7oS3
nDrg7H9forqWtkJ4wqS9ysWFn1BkB9Tw6OlCj1IcAAHeL6tMQMJPLDvwmNUkMlkqZGPjMmnngLwD
fYol6WqcY0NPd3yW6af7GtTMxQKzjfZmocNgvZO5VfbsTPcpF75JwoZaHniDa1TR0Dxw9PE45WLZ
VrA/YfH8Zy0Wt8mifZWU6SsdpoBi8WLpv9DMaYGvFdjvIkHk44x6Z8cuwXRP7Drkmeh97jgNwDNW
2g8w0N33WZ4zHQVFu+ZuPsYAePgGX1KjkY5hRR4DHyPi+J7hdOZdZ7eqWeFHOmR7kkD38zLF9UpF
uBSkPoJInr8cWEm7lkt/rRQSilX6jmaOmv9Qz2QDlWkzXCpQnRkoROy51mrMh4i+6MWlcqrvrFOb
7li6PiavFfF5NNXqsLG/KX9f2wwhtS4zaTQUj5mRtrzz42aoukRSh7rQm7IwvUZaJWYjFlPwojZr
JHRADT01atIgVRIuvuzVhJ3lbMBAAxsOnfEkXMpKATwUXifh7VjarF9Y3uITkUsBGKBV5Sjc1Yip
6GpvgXLEnHxBhUlNglxZDJrEBVNQOBB1kwiql7HZcQ2Q32mkvuFOu4NjfQL2rhcABrGPqA4Nit4n
nPeHkzmQ32K0H9hmHxLQKAMydaM7THDB2BH28bA6J0ziE00ZgfSr5uCn0h7nr75Vk/2eSUeggiIg
/QA+NEHGXyCI5SdsibmxVijRGOx1A6pVSpT3UGFlIdOoanDTuABUZaPW8U3MOcelvCdu6GJpZaSo
NHn96k5/rMpFfcWucFtoqeEv4wgfGl/XPO/2z5OB14WwGgnC0UcDmGBlnePqURrDpK+RQUB+5NNq
ekiQZb4SyIe/RMaVbR6+q9DUnDzXUb2THuJaHRwzFKgwisf5yu/8NS2SlQl3vlauRGmaqPptxQ2N
2jG98d5coJ6Jmct1CdkusA4jnoA5ZqQCRku+wGt/YVqvZTxrtwvNvgjf8jXTFqL6wYlBt+nbmkiT
LUoqYt/Bpn+dWCUILLfD6/MDZSb5efohcGJOEY6UumQDPZthjjiwbfjFnACcZo/ZBH9bk8jWtcan
eWFUsL3dhwLXPjr2Npim55UauIdN0UWAalfJ/Vm54H8m6lfUx6Ojvbs6/QuyeXMomlY9gbtaqQ07
n+FOMm2KuGWTQgTdPcLwz1B2i6ai/u4TJ6Ym2OZJpszTM00UUqPEuBgoWB9hQXaF9AgaHPN00AJF
Bg9Tw6mAPxAA4MKiBD4aVkamYJ+CketdL66l/qwjCGHIxDhGwwjSDZ/iU4R7W11OprtTmHhvHw85
WKljfpzoYoxrWsfLQxTeddbXojFHHeHFgWDkAGgHqMJvKpNlAEVtOcPuBRt76KkuXssSqALimCRk
oYCaRs8xmgsOAY2uarVA1jhes9RBbcBNl21qrST7y6vEgqAcSupsdaBuZYey7gRSvrsAPFS0LlPW
EW2l+tkg9p0TvQFfDKvHo+YHyBc0vjnbVvfe3Pe5QXSWNjQ2fkcvLx95Rmek15Q9wRWw79cdyNpS
O+aMPFhNThF2pYhgQDpcCNwG+QeQUIgdCzKATi+gE8ylFIZCGgBQ45o7cQopNQ3nsn9MqCsSpMqO
YkTAoFcdFiQQ06ydGgw1xm3FxGil0h2qlhMCnnGCUm3puWbcXDw+iwDC8Q3fr/+NG/yrlLmyw6ol
eWYwpoCShQ5lFPtWRSRAnQTJ2kvTdfzveQCtTfhxU4m/ri5lBKATXZjOqNWbQznSxJJgEOyOHYpV
BTongo7I9ciaQ7a2gj8POZ5sMjpOZORzBoMr8mITakiUdkSbg2VmR72/ufqSdCuD89EIV0s/X7GZ
oYFV8dvrvUzhtYUTECuFmJkTBkxsXt/w1tOXEiinuBBxFit9cf+FZShUmrHe+IUWq/PxD7oX2xX1
tckQ4JOtcOOXfCQQXrKaCBmGgRFovf135FLmOdnJP1/ScD12NJWR/aOaTnP88Xe6as2T3Npyet/7
XZs4hA1ciINY2TIJ9CjixHCbdp5CSicXx11ICF+Dwg57VGf9wUI9kNNGhBWDPfEFOL3rKHxyFkew
NQ9zODynzOM/FD2HyE0meVCf9Fe2u4PzTWI0nNpBEnvG4zcxvjx/K7D497s3iPrp7DH9t4pDf4+7
7+NOcg9ZeEslCqnpv+Gd3jzFOPz89M47uGrTdrbUtA3/plgJgDyl+45T74VVp7Es1w7JBoIVAeJo
T+SGzbpmDorsJR/MmdMyqSzAFAea8IPlxeQfmaIr6+2s8hnsxGOzqfph+CGmMg8r8XjEJtPDvGaH
YN1qhW0z2sfIwGGx4jwYNEw2WEHz6/QfM0XEdKB5cXg0Chx7QJ6fb7UxXiMzqlCqZsdB5rQv5Y2R
3UrlbBVAzwOrgzq+o0FKbStn5XLq0vr6NhvTXI5wSacCo5Hpg3+CwcGnIuryzK4YzN2icyIUaURs
ZSFLwEvxCsiXCFCBUhAlyu5zJ1XLPgNEEj/Syy1E19FQSnjMXLnnAh5RGCtQQHp4cWWLQMyhUZ22
oolAxrNLfxnCx75xOgC1+KzzT0Zu9XXuiSJhuu2v6K3L+r8Ejo089cwT+N1NT+MSV6uWL7DVsjMI
sBLb1bmAXh5Zwi3y7zjVmm62BueOL/EGVAyKxSXtPMLxAv7DPu/9YrwDct3bE23QyPGzpbc5AqJr
+VxQXtcic868nR3gCcz9zYkwf1BJoUmhYBzP7zKexQOA2Q5BJ1rP3dsQLOKCMjQYrfRco1jfX5Qo
J/fTSy5TD1fW/8mVtX3x1v4dAIZxxVfU9INYOI3+t2lX+CPIObR2g/xiRtehj7pJSHoXBKPKeH1E
q1DPodkICPwK/kPDycv3NPo9pXxQ/dP44ioyJeLaURL2yS/iSpDrkhQHWJIksdud3o3uAj+tlqkb
8UTZqSJOLluAb5qLYgb82CfjAV7qAlHHVtUiGnAxWuojb6cMcb5n6dP18wmUIFKZsyoQ+3HQT5np
Z7u5G9OOA7+jX4VxGWARWXV4/HEN7gJs/6os9u8H0nX/ixK1x/BIsyg86rj4KrufAzDQwy/W+EqY
ZSzcYncZW+0sDMaYOfHBJKqvl3NFA7iFXvQer/NR+pa4hyD+tLHeGAoyjBHoHFGM8I9J+iXBHmv7
V4jvzCvLymYgJx8TuDsdRv17uGCA6N0PuDVmTUCyG/OeGTXYBD39HfuLmny4Lgx5TC7Pzq5A7bNe
6bsyo8QCiImepbq+caGAOs+76o8qewGSabyoOFoX6H+0uFhzx9YPOtsUcduHxHgzFGP7AXC3QonY
2NNpK0kWDKPI/F8Rj1XwHa2EFvhh0xQbtmA7VLLKfv1fke+pFVqvBlUjFF8Y5xjc4+iBx4Akg6PC
ozs1K4SgQ9mguB3vhWIeGS/6jLDrqdJS00AWGfl6ZH/qLUo+IwpCBTj2zjzKq3evRIMm7bFxndO9
irbKYc/iHM8OYjNBfs6FEBmYlp4eVfEMG4g/vmmz/4IOeLx9waAgpCew3VEUgrjM1QaXGzbA8dG+
5/tD6zO/cIKoT3vhCJDrQ4SPHnapsimeHaIvDsKY1uD7DcjYg7AqCI+6jEtuKmWfywBR8TARgOun
cjAayeipxHsX+tW5dnrWmsi38kHUkYvSsuomU58rvYYi26Ykg2UYL63V5Xi3PX7ebKya2L2xiMKM
6i96ddCiEQWZXNwhtoIQ+ZU55U0rozUssvFaSiq0GvS7EVaXGsQbBsmEwuvNU/tJxZfly5gclkxN
SiGOuZgFFPAVd8ReVAloaT13GFV4G25j83MGaiSwVDuL95v55PFBLtYA04OTMmtZ1hjMPd8wDMw4
Zj25R1yLyHv6iiaLvOA/jV/Brv/of5AbOubriWj1KCqpFydksn0NzplzjcwSYmBVcjyOl3TsyY3b
sJ6WXrh9giUWOkQkgM9kDCsPMstft/guWxq/qQ8ArU4JAJ7Q2927pivhQxmZjmg34OdILReQTFHG
F5Hu9h6TiFJi8sr3qT3aITL3QzUeI8GaTCW5WUPE1lWf/vFGuz+z+Tz5OJLBi86F48aq2hZ6O4GW
6iZv6OCfc5KNHeVMQFOzboitHHZw3q8q8qQsJJ4Ir3f5yjhzrB25/WKpnqbd5t+rZP4HQUG3DI+F
CdqUH4i+aZC+zyojemm5V282LC5U2SWwq62sAcxwaM081Wznzza0CRLayQfMZWi2vdODumDf3p2q
K4Q1p6KWJAQntFeAc2eTjpYzdDS3qTj+rfitbHBqwto+4q3KtDRiNUk6pwZZCZG5EbXSqevWZ1zt
3qi+5aBv/H6T7V7PhQLe1UB5Pa/TJLrOwUFOiwaFlzRSION9X3P071hpEvEpTnNAbrn/bxmUCW/y
3Xpi+B1DLJjCUW1gyXKIKiqHCX5PkYq84dQKFWBv9yzp1o3rsZyzNt/1YFo3nK9wOCWy0X2WclVh
7+nuUIHgx922CCYL23/1UxDsBJ/OWdsRr76/y00++od7XduRKCgRv3/BLR6eHqrm/BLZp7L06QXl
2u4Ii4VpOroSQ1IPXy4iRFPEu6MR4KekxA0tHbtkkKJwL7H5j+xNfNlnNEkQPcOmWhmiVt0Lec/r
g7ykmRYQ/lxVi68Ur+EPhqcqNxyoHJkHexzHSHtyMGiUrOssTLQ1sWesPq+Yj4NfOwSufSGsd3rx
gVEy55zBUQ96wcstrUwBISXJTr4hzjz65PK7bUvAWC9Vxbt93hL5hRV/XaTFsKOxhku9PLx8SSNp
JS9i1jNS1+WVx0YQ18gm1KPaUJSUwNGcgSYYyPvyqRkak4o3IS9iA3NA8yIWV9Jlqm+aaUNv89Lr
tOC3Irmvf3SYXrWy5mbWh5b4KfYsNoNYHn9zsEzysZCds754/Cj3YcGgxnrfNqdP7aQxqGqdypw7
V0R+Qu1zbyS99dPBWkQt5nZ4SkaFB7bIpaat83hIFwFhQDtvT14N2gGyMLZeI1SCyRXkJIj0xgZr
hQRlyHFQ7CPFmRNycxqH84awd5CeQfCcXnvCM9wgIQsgdTzv5yJ51cawDaAYzU88ZTmk96Npjl2q
oG8nqIa4NXlhwfc9VvhiDGcNxG+2F74z0yIdCF/Nn3G4R8c3hMP2MKEkiquXQPnMPfrJIgMyHszH
bVsfsiifwPrZ4yf2sz5JZAuZ++vBFsyq2UuhQEaLRws6Jaf7PMhJ3jW3w622b6OFDUtcd1yuTdS/
XPsRq4pxmkMNRdhuo+DkkTSZQUWDKq6H5cR4OcHUYWZDmjeysDPf9HelfBAP/K0cZ4srJC0wf9tf
gICy7Cysqdlh98C5oc5p83aPWvW33wTgFbn23FRcns83ggi2VrBbw2PCgX6zpiRzyUzG+ja6ZzVs
tBaza7Gpl0WKHqIb3J/XDMSKCIB1hPkswiWx0MLmE8aBe6f0nOmkhICeI0t7utmJ86k6nTFbMe76
h59Fyn1CRF4qqVJb9hVdQSrk32opi6/k6HdjNAg02JcnkDHq0Xz7T2PYIX+RrGNuI3/3hOCuaxbq
4drRrRV3t4HdntKpeTgMQj0FCSFExCKOgSeui7A6/la293H5tflE46jOEU2HM2X7hh+lEt530zx0
Auuuoo4yDgDgNoAUyQFh00ZwF6Gkt9JKr/DvOAbtj696NChcQmHRbkFvVIOVUlVUVU2fMevUVbrZ
CLuWdzlRLBIcm2fFOwlyFIMYE1EtVqwWEg66Qu2nEEQow87MNygsfJseIf8bF+U5sbOqPjdQWhKv
XB39OMRYFU95ftUv019bQr0dl8Nhzd6AR8F8W6LHTRqER6enE3AUb1mY6fvlmswxtuH2BcHs/bfo
Rvlt/YUYiXwauVvhRI7Pi4aNTzsoTpWZVVZFCkD6F/rFLV6K2RTDhtE4MYzYuEBbsBe2m/7ESaQ/
GPXLZk0Hv8FDPXnXZdu+2KfB/FGnr5X89q3HyDe8boBvflBSjxhothgO2rO28t4dTRzjJTuzrfrl
euDJ3jiWCVlyXCNSlLPXI/vjhpq4Ni5WzWJtY6l2R8bFpixteen8iDlhnaItQSDjHXOZ6IK2VdZo
1z7Y6dJwacGCDJ6cx2rioqEx6zcWltGXxp6i24vRxYw7vdigyciJ+s45N9qxelNt81klIaW4XICP
YEDfjdTVQahRplZtS9ftRt8FC7zlBcoBydhXNcS6DxsJvln2I8DvxF17drCiS80LpGXH+eif0Chk
UdhHh+w7VHl4aUuJOBvwfKKXyQlTp8Jju6qDOLDDseyOn9Twgze6zJzPO3/BCxWauiMoh9KjB7pN
OS3HRInvQju3LleSJw4tg3t7qpcOApvdrX6yhSf7O/6tfDKC4B6ImDl/00x3cuYws72OxOThVR4h
xeHqy+bia6ZfXnek1vHb+CbH+uSqEnhnViWUsY2IayW6XdctKnxhlot+USaEOsAx3k6ld5CDMlfQ
qhpv/nGntBJ9SN1zWbvI7UcDYz4uUvXXPrT247r/xE612IK+B9Qube504WuQH8vGEfpxTxYG48W9
THxoPnu0Cgi5rqXTIVx8FhcSPbnQCJ5tEzz5qBitsdCEVFYrONAQ2i2i5zMetHi6KAZfjkuSbLqw
JI+6aGzfXB5F0oUd2TZI+dLkxq2ex6MRVV79nsFIqIerp/zO9TgrS8pXH9dxVjk/+KT6vuTYbY17
xn2Tukfph0ArKvC1sl+vn7DJhN3sZCna2aTT/VR1gYEII7/8gAVN7qkwaSlZExkyT/kK8N8sZjsL
sBDtYCQmSzd5euxEgyoIN0Oftdwljrn3iBV6CkqRNARjl8qV6A3d/YANtDgu9rM5G2L8YeU+ss3o
lRhqfcyJNqQOx0aAX3YWAR+kZFRTk3a/QlPMHE09VErEkAVffhkF1a2/Zarzfg/6sda/8pWhNM9O
jB4/5uToK9gRx2pcSFQT5XpCl3A39OLKwz6zXsPgBeiRzhdcUQG5LOirdUROTi1tVFP9n7/M/9JV
oJnZV6Pc3Xj2S7sXpqx4waorzpnYFAKyMTELPYCYhQwwHZiYEYnO0VPJoUX0LxNu6ld6fXkIQbyw
1qnNtIt2a4zzCZjm/Ocu+hre0gecqEtCc37cyBOcKNBRnBv/Ew1pN3MDGmUtcUJhrU01o8ESkcQ3
kTWPWq7yiLtpF23mFyAOCAJEKr3xqhqZReYndkCdYD7BwM8t7MiajYULMEwyafdbLlywSCWJOr1K
klGWIHXEvCeWCyRWSELdKmssg2bjZXtRddWzseg4hWxas5tA5Lj3ASzCjLQA1Y+xJN3wqwKNjah2
K5OKoEdD7Dizsb1vLaAmgFSBgsrlUyJbTlgO4FSZy0wc6ACKD0WjzJxDBRjhfo7vNHYkvJ9TPuun
yHGNs/nGljDC7lReRS7+9JIKXwg8gWVNrGnqkjyohqkrDZguzZ9S7vAz54wSH4NceYLUpqW7pkSI
yiqUU/Cwjcq/7ABtemPj9j+qObG01li6vpVGSeK/72oBV0ABlcSj4pdDFCl3S5iBu6CcgnRfB20a
/ZzVNRMl3Vt/BGnRaleMcIx1+41nYtsXTG2HQ6ViwzfAbcBBOiW2nCDcJP/ww0z6RGFoNCG8ck36
AuxAG3MgWxQTWOPK4v7QcrsWfH7lEd4x7yynLHHszjOtHSId6oM4BPlDOdaOs/6to1V5ML5Ggs89
HtJzD7zx0gbL+JvgpESr9QvbSZmKamSwO6GRCO9IZVP9Gj02dKinAdRM/ZrRFK3XBnvd+tE0mCAl
C8In7bYM2g9rQ9X7R1i4vsUQ2mC5QXlc05Nxv5TpJjaeIYkjdtFhe4Kb+oizwjIx9IIXLYQmGpcQ
VYufKRjophoBn7H4IRBZU/1yXoLd3qJQtASNWaNOLfHJxMLnZyASWfTLk6yJ18RfXM5Wp1awgYJd
583y11RGmuGVomiJLOA+hxkSNHGzOATjPo7qq4/+RZfRiHIlDucQRqDfyDceZ2G7jKYWtLChe3MH
2HtegKIZ5iwwRTex1+i/BAJIjTVL9zC37hbv19nhBHd80osm9GHy0vqvYrDsI/N6HNcZODKN+UYL
7jpLP0u70liqovL6yAP67gUekvIQ07YASvU8os3bqLp/4bVw/2KX75g4OcDIY015zUzDNfuEnJgq
sq4EhZegA9ZI4mp6yawDnEHQSnK+fw/S3033bxJAbOKjYIr/UNZWr0kdKXsgeSEuugEerLgCaN+Z
GO8S20EbIdikZyF7GA1C/7iQAtlXcKcp43VTEmwqw/LH29KOyC+ahf6ZCLaGN1w9yuguw/hgQh3H
LCJQVGkUxPgY6pTb4Nb4QYVs+I3QgWAJ+6WCx4T4eA3U2wUl5pAVfqpCSxDe5jgoNUayIxe0/UpI
TtyBRljwgVHragVBD6wC2rraNQ+DeS95JWBkAr6xOtqLQxnnex94m+ixR+e7Zq6S/GTh9ZAv8CtF
d75RgRsyMao6tS4TWRfWGSC0/6mLsVv4O+EoNoaO07nG/S1E+30LhKJ4AW0fowruQBAZuUAdWQaN
JMlshOCrhNbvWt5A//uzmRZzU1d6RNQWbxCeDtOyLpc3d6MPR/J07guW8DuHh/oC20Dm1FPVbP6D
l/xYaApQRxlFnLaakHmXGVZRIK9iY16XIs0l+zGLjZtiGJtadqV/1iAhhUmvpBesf993lYdlDoS7
xWD5EZ2pihhNOw1537xaVVgVK7lorBC+qWqYWM9uYvIrHm/RlwYzrQOkwE1UFx7SUGp6QXUiw/yn
uxUhTpuYJ2CVyW46iazoRu3Vb2eqFB5P1E/yE3iVcUgYT6Ny9FWpOiyPxPtfT3WSAsNQcV3k7fK5
poDP9AA7cjuarDFxpyFLWTo5c0FglLL7B9NSej1vLl6AaQhGqMaG53+rjjbPeW6mP4W1QgWNZmgy
NbdfpC7BUbPT2+2B9Sf98NOPFl9V8iSIDK+AMH8EhXDZGjf3li8V7N+a4XZsiEiGsfj6RE3De8Kd
UMifzUFeUkL+z2nfzVrLVltZVP4dHFOojpvLvG9nSKUEEFd/snhPNP7q1BIzSv2zgLaOYTgnT26I
sVrOaMCiZADNSbRJlueKDOurq9tz1KZz7LFarzkHsGdeWtktXPLFvK+f01TzjZBpp5H8MvQNg2+3
WL/8WrD3YIOt8vT6mE5iKeDJwjRaq+G/5E/suHMv/HAEZZv4D3aAyD7yBP/z5yXM1YVhaVnuW7Hs
DI/1TM7e6CpzKyRFUfgIrFzG1D7AB6v6eV88K7sWPXC8Pp8+e4CPUzgc4LR4ebcuSgXcgn9WmjfR
Ts1WVk3vjKEviGkW6XGNdg4SScfy1L2FuI0KmUIflyW0Kkv8h3M7d2m0ZB7/L0523asHFa0MkSQI
HLkpHgDo3qsMCCODwOs2Ee7we5bhtoAv8ybfm3/LLLHPShtTJ8vaNWXotwJrJXiWrQxL99UQp6gm
MLlJFoPgrJ/gDamG8FwymmSv/c93ZR4wCJSru2vMX0OeZzHjL/cefWXHpV9GMmgVqEUG67/znWHo
h/puX/bpmnY6/PGDvfZWJriN5nIUEv5LW7QLZqtllAZ+kXvXc/tllNwuo8QKmz4/9OwVdwmFMQ4G
KGKN0m20p9CS/8dvyNtZtgW//cqglmzepb5I0hOne3uFiM9DjTefUYoMLXo3stzhVG3i9u78jiqn
gmvBq/fpHt527fCIdoxQtS4eDzugoml9RzvDXUyAjWg/H+n6vMbchIrvKa9OPL3kkEVjLK5T3hFI
2I303D1Rw6PBpmo8VRc8CBrK/IGu0Va0/ijdZrmJ0cBSlV6OVLmO/Id6gIcCuoNEvyRCJt0QtE9U
c/nSzoUKWA0fvD11SpiI7UKFL1nHfh5cHV3jwli4LgE1XE2M1bmyO2J0sN40bIRQAaewtRWcwddK
8VvIST1R1DDT2nSD9ozJX2E3zh61RanOArL3xz9ODBZfBuRiUy6iIutzgGBrSvxZFoNZpBoXWfGy
sGLKgG5psVHrSzM3/gZXAVn6RHCd8Lh1IRGHWL+f5Io/X1BSPac7nHO2Q39ipyq0fvSf396IxfVh
2lXJo16PfqRrAsvYpdT4bzxlRMjzVz9/iKB+Pc8habqRd2p2ySRKpH4YtLW8c1OVfnmQfEerOfoq
CkbdOz3WPq4qAmuQntJY+vWLd/bdVxIQe47VwyEKzOK9oFY4AkfyFL8C6fr9vNU+eNFR0+lWB+HJ
kgv5ECZZnJBIaDL/qdGTXM/JVXxuB+ST34AII0bZOlv4dCET8jbA2bw+IlTSTNJhzRsQ3nRrehb+
y5FFj19wONyb5xiCnT6fY6RYnViWNtZnHreuILC6Q3N/Y5lNO5ydwup398pZ9ap45aet5z+nsqRU
DIdg15VNDokKtUrVNMISPnpHjEPoRVpspUuoHYEEi3umDcJNo1eO4CrhGvHA4bg7HM4H8WuEKC2/
Vh8MHqr2Ov8dQs31mJH0ZYLdxAHkPg/cTPRYZM+2YCpdiE+sZ8O0RJMLTLOLRC15QVw+tlgNbbtx
6/itSLqxTfuZJpjwQbkUU8vEoEEBVeNYBCG/8pCsitWA8tbHJV1Wj6RMPUteqBI5G0YHRYHWOL8c
DxgjLPnwmq0kQgfZ36M4UiparSKj1Zwchv0zlHaIOMiqqIdcO8IxzsNOWehNLvXsfntPkBC3VTno
xc32phEuRh8ttREqN86IV8OzxvmQX9RZoZdOurVGfQcnyeJot6+ljz2rowRfWFp0ymeqdA3ABpI5
qUdb+QHR/fLnjhHX3HWK6o2MxfELy2EAV6iDu+2Kp3SSj+6yvFGBq+E0DiYSSKRNAD1Nq9wIxITp
GFBrOWzHu+GR4Y3WmYujBSvQpJS/Otfve4ET41R4979PkT9Jjlgfxq8aGEzgAdeGUjfayt/jdyIi
95q4HVAN11Q9qvCE4qoVkwWJfKEPjimaZq0fs4nIzu0b0CpSZ/YmaaXbEGIoKcn/Ori2fGUPywuX
69b7Wib4315OwsNysPPbPmwIDk2VlGyLjhAQ6Sygwm9N7FjhDasdrt+pH6bZRvwI/0uNs5xAy0/5
3CLwJA+JsP9atcI3qVMNcA5I/TPSVCguO9SJg0FpTvi7eBPxzMV/1yEzybzTSH0/g/Zx9azOJTo/
7efZ+vBy2vBoPo22tGf/lrlDkSarpgAV04RR7t7eMvAfylFQnXUAUecKEfDZMWnVN61DhJaQXM4s
nxehjBuFQ8rGSTPuI6bp1MJ5ref6WsZMWQo2EruwSP+A0M9vNfsKRSqMeEqmZq8LSTZOJlqf0MFD
X+MSRfdL2gkxpzXUE5aQ5v9GVWyTLeRuqSab37Zu2jO09FdpgBjBOIJZrz1MJUVbS4V0xvAyj277
RgfsXHWW7k84f6yhnukE3ME9Gm1bpsEwXTUj/qeFAzZMI8Ddz9+fZGEYDoJYF0ftYvuTB2Tx0026
LH5Tm+DSE9kCrvhEW1GFWjL69qyE4+C2xUEST26wPcQ0mBRgCw9a5zE5d28DSHSJjnYco/gd3d1O
+ZGWJOdszYK3D1SGTBBDoo+858+RsqvLCvgnD68Q26q8QGhiW/nRhqey8ea+Hl/qi7UlEhcAaPyD
62+qP5WHvLa5D5Qx2T3sxbmsbIhKav5Ag2nbHD4WpdiPO87vf9mY5EcNtRMJ6blTLwvPgmPXm9tZ
6otGiLmEEPlfa1BsRiUJJSgkLQy4UDwKyu4s8WXfyFWnCNeT54mTeXKFQ9E6hOZZy4CA0MijE5OF
hm5FHi7NUgFkCcTeOprcSK9zTLi2bGlIGb+F0j1ThJKSX5BoCw4T1ggnyb1f1uqpruKyMC+Nvvqe
s7Q+82O5JtEN+MiiBAaUO5cm5wxoqIauLV6UGUgku+ZPb65gOVmbP3Fqy7ZlI7GrnialLV8IjYxw
lk002r75VnzoHx+5FallKhVcUTfImJWxJ6+wrINDg0/nkmCNiFYB9xyDdBVzWrgDmvonqkgtQHaf
sdK0TdTlUMU3pOHTAwBE5KSytPRVmjL/9KP0E8ygCMtxi0GSyjhGLDJEmncuAnWuqxmcJK8DXWLj
7xg9JVjpm6JKx4+29b0E33Is81EzWIQV9K9etptlD/hovTPFYjGFkjmwwg1C7mO46gseBsyFOV/C
4swkpDKDxf6cySGNHRhpY42uj/jWTIOR4RTKnpOWIggiSpvtTnC5pUJm+8JO0ESNW1CzG4ajuovG
+hddsufTPjqpcOeuTG49RVe5PYPBCDz0rTDB+/SyGqcj8tIbNQ/qmTLK4u5Yf4WDkmcf+KzMRpHl
abMPSVAvzmT2c0pUHtnlul5+5J1prtYFRdTjY6VKEwqtzGzClHwE5NNGYk2omlVHV4rULE0vBQgF
fJd/HnezMoJXFkctmsfPrJQkNRlnKKi1chJjXHXh/oCzvrIDRowlAIN2mK0bDXZIg/nnZQj1pmT5
nx7eW8apjYPwVbKZc52EnU+ts7ciaJdEIs6kqatdMxm+RChD7NOWhH9r+A+KZJhkbAQ1ISxA4WC+
Df+vQ9i+s3h8j55HoKvuANxEakQ0m6GrLTg7iB4CjqkuDCf/2UEDJ3NLv1ymOKH3up0sRgMFfIHd
7Jdzt8Ws10pTNAgbr8WHZjCigIKpR5KAIGM8/szqCDpOv2Z1wW56TB4LKQSVlaqOsQUdEQEAoO41
psjunfZBF4q07DIqlWWnkzQRl5nneV2Sp32ZXHBKx2uIzplmQAUCGcp3xfWjnZRslJN1rAIhgiy3
NDhLo5bPzZQ2qnYIAS1f4Gx3XwzhWBUWrIgR3fiOHEefOB0psZQdOur9et+oJKmHDvlOkZgcHC2w
lFcIti/4RTBF6xJ9yCbpV5wfxhZIgbdRhXCcIvVdePYcIMrDSOwEarjV/RViTci7KCei5rNdcwyy
ZSPoJs2kgLSM3txAky9ied/k4pqMkr2MVDrocnA0e1AJFGn0FPwTyttjHTiJuvlKPGLtEO4sy4W9
bt3UvSmMbRiB77DWbfrHs9aQw1i0mj/YKnWSaEgQke1UIRSxh29OGMfp7svmuRh5MV9jKzWpg0W3
LXJ9jeNfoyqFk/LQOoHjmJ6+F0C0C1ouZyK9B2LVr4Qfw0UQXYQxYBQhXogY4giRoqJ9ZZIvK+g4
cad02KPEcB6dokd3VGdN8GW72eiQkilthF1P0WVima8RPJGitcK+SS5z8aSfNCNNOGsY7B/9gNO2
0rLJ7MpFmXLXSVpS6EMS53ex4QC5MyWdGDbGFwrDQ6MK8Q+W14+swpCPjekEmjcJAlZgt/687Vhj
25+SKdHMeDyx6ot+KQutXNEm9DLZSElFvO3BRF++LqaSP7QsG3+AyVqBIjDZUgQl4epk+5vKkMCe
FzV/u8Je+gyiJ/3k75qGtmqqbIYuKTrqt/Yaz3w0IynKt1fSHWLsSUTGrv8OyxulYXFc5H8oqSNp
6NncBB+7oMpIMstQg3qnqSLEA/MaqWfoYfZGGULkM8vkW0iDXGhivqyTbpsQTAONfiDwutLVrsK8
ymoNMwtBXXJd0J4I+J/2zhXw1I7nTOOwJlsh7y+diUB8JAyUOzwBN90S8J6i+tNOeBvmk0nFI9eK
jo2vB24nW+Y/o1HhDEvXXUg+rD6zKhoe/6EcFhAD3hoZ6zLkVNxuueOh/giBZlxaIjcKeNfI8FVf
O+UvWqZDZE9QnIwul9X8znXN1njbfXnMpFxxvLlfGoOB6imSCC0HjmKeqUfVVwhwlB5k4Lh5yPCw
LdCBLcWdLuJemMWQXnOT9cM5J3W/LFGhMyCUnUChfEpwyW2gIGyg+8La3zO00ApSTfbek8Wo2I4c
yPp3y4I32sy2a5C4Cc2SHC8iYBpI5Zj8jSsCcN9P26vecbYG7Bj8LDApG6Vrdruq73h5HoIs9mby
mC7ivj1K9lb0re5C0giecL/f1Kx5c7o3erbWTQmnC2Z5/8L/I8naCGf0JH2cw/W/lx3dchoJK5T+
j0fXbqlomuAQAm4+/90pDyzcP1nmTXPI5zdEYBI7UoWGp3uTs4rQlbOTLfrXiKL4zuKLo9WLUeTi
VL6+a0xhGlKyyoSw7fpelDItzMsw9TX+ZTWS9O3GTsB8Sof15u/zBa3ZiDnImSB2tfon/K0RtXQS
x0hvibYMrhULX5j7iKB01kcl3e6z303untGNKKTnPBu7NcfE02um3XWTRbXuVKovsl6s7HzYuGhz
EmQYdoA0dxE8q7bLGF47q3QnYAVSM0/td58oxPXZDKBUaZYy/KYXXfMf3Af7lB7XbtKK80MFpmBX
BCqgIsEPoI1h9+4z5v4zODh2K4mHp/drv4VL1qVUfksRZuR/R1HXM0gWqliqMhCs7wH+17pR+deV
iw/NW8rWBJd5tYOZVsDgMqDsI4sPNeAHstQr70Uoqj3i47JD1rLeWzGxzMnYiXxBCif0aCAE+jwe
g69hWtHXxfrSHM90fmi7QDn/q2iXXTHJNN+a8xqqXCnPsys/FmZNaV8+z2RNDJIPMdnqkZr3koLX
bAWznlf7NIhG+wG4Ib6DcVvMBmekLj4r0J6D6zziQq0ku4xaM2NwUefqkOFnZ0soVF/BKF5jz3vJ
iSjgMF02UUOG8TIzRXI0wv14+JPwlG7spYCAMR8Nf/5H1PNjtjRkZmFZOQ8wbvsDSqLcDslweC8n
zB95ivRpMNEN2ZNZcxyylIrLAALvaehj7/nyZEfZmKzw/40sB1o6a/EzGjOvwQIpsPjb32cMa1+d
sbNzQ2SMbJ7RzCpxTOTqo5MD0oqt+YdbZYhgXWkwZ7VP52s/WeS2wrY5h1Kq4YLvJFvkPdhSmPx7
RURFSw6n7mr+voDCXNnZBu/mo5FN2/mXP+v+IjOncs/zS1j7rtmCF0oAv314SebZS0O06GagbgHa
VZ+Ss+DeCH6bCaXxuMU3xtvHznyufhswbfc7woL9fl1KJEUqKSynue+RJHjdHhE3FswECue/Oabf
yKGIwVW76jmu6TtNWzMY643gpu0AC/vo0lGabmohdTHgY5bJwiVYhotYCbfAO6Gk8UozbJ4aU8dZ
+XzSjFB2cls9cjrbeJsLRsklpwn55b6hGh4r0lwpnVafoB3Auev1rcUZvKmUl04zBaBqB/QNWGr6
ch5MK0MFj9NyoYuzouBJ+dj5zBK2tcCh9jS7hMsZX1Yw0CfJJfl4z/V6bu8F47PorOMtHfsZUXVW
h/qAxH9iwbMcoj59TxDdFsgdGcOAa1O/6UBsNIO2n12P4xTQeeREAZE5lDdgq1MQAxcHjvaWzkB4
LDWlfFL3cqd3stC15HTCG1d9ayfgfjCE9ZVkVOcOgfFZZGEJELxx+oyZT69WAXJtE0S5s+jU/+8N
u/xV+P6s3n6CsaY9ZKeYsFnaGMgopqKiMBg4K3BjGoP5WMpfpYz5Z5RBs+U1KRrhFOZ+I9JAyZRY
Ccrox1ZEMRuWC6xQ2zZwSCyTUs/7T4c3K28t/u+bSbv0G/Daq3ZeW+zx91sCuQg+VL1h/JBzzZ2l
9F8Qxn3roDo0epI78JpkUHkk9ZgkflIjkde5VnrOcA5paO0REEqfLep0LeJsEGU3VdGbWioJH1Ca
nEZJ567QXbdd7tfmPpQpJsodc6Zh2T3pjlupetAFEZMb/JTxedeXauCM2bwSXxShBtbd0JtVzYRM
HG5veYfoY9SOFsSBQxaKhFzk3FULvbBShMiaelRzpq5T0sLxhwCUvU6zbKsXwd9u4dfS2A6wN71R
NzLI9IrywDxfK4CJqonN/BxwKs5njSNLZkbG2KnytE8SYmTLhSyMxsjRjgiF4rlhcnE6tAIc4nUa
4WNUFS0g8RKT/xjSOfhzho9ZgInATy3iuTfKWfHRyxgCMRmEFUabYfb85Mx05TlXu6OYPD9TNEv6
OJiXMRnD9SsgAryHHu9e+WPRRtaZ5W0hj0lVoyJVWa1TIGqtS3WBUvAWvSvVMxI9PWiJ9ou91yJ1
tRt8hFKlxTggFFl/A8jGJWusScuhmyuIgSp6y0rBwUUV/4kiexmNezem2/jVM89OqxMzKIFiRvUu
6aDVOoqc+6XncyNmk5dS7SMrbf3wGsEEQB+s48C/cgzfzONVPAMRXs6Zs6BQ/qrIlY/4yVEQaXp9
Z1YgX2Ij5TV+AwZk0vxtJq9jw6oTjcmCpXvHGhnFlgpPc/r8gPSHcqzyf1uNqfCkG59d3XSVGT4b
nNQvmVWoRMl5023+6vA8UtDw1nnbjTNR/MyrYN0V28hqgEFr49/bQi+6kvSSITrngRD0zx9ASrSO
JHyymm2smg7nioIeffv197yqtyTT7kkV0d+GFQNZQ0tiHtB7XAmEon+OpuijOkmfwSOhfnykMOag
SyzrGp1UP360zGyGT1//LpM7/BwJnqD1P0T6pJqrBrmDhewzlRG7QMPK7JrG1eZkczzpaSYP5Sd2
s0IK6nIFRy7LtecQ0Ehp4fl4DpASQtWMROvl/daquDGMUvuSfOS/yvd5tqqJWKFswlw1nK+UomP9
L6DwABRRVU/fFXY4FX9WbkNKa4eoLXg10fuvA2p1lZhrspFkOg0LmWskC8woqT0FJp+tc6ystu34
Tzh8lCdMwFD/W8IuhpPfA0k1JOtJ3GLOyY8o7vfbVqEjmMPKcOzjY3yXmuQmLKl1Nl6ON9fqi7R5
b663XVfkcpEXuDWCixIU81J5I9PZ4BCBw/+9B8AusZzBgP8u0Gd+zxyaAGukLaMkZBitrJyBJ1hX
ALSsydyBoRnpZTgxyQlOUQAhwEdmF0odffKM+D1A2tQ4K4i+Hl+E64BTSVs9SUPOtazy1jd8Pmjp
JJGDn+3E6UjoNlEPgC/vGa3r8GvoYv+nmJLXuKhxwocw/fqKKcEizJd0dAnINMzQT/FA3xKLIzyd
8zr6frwoRQhccPjynngSnL2kSNNWS/W9AU0xnlakWpuHYiMbEeBNimGx3rkUDR3w2Him/6vNWbSF
CWEZgzYsllTlz+AVUYIpi08kYLcNeHevATCtCkdxScDj7VRI3MzGbkGuhEbh7r36BbezlKM/iUJN
Z6yUMPan8vxX86SaHKx8DJHM1MfRYAwVPqoSL2oaXvdeDLUydZonwRz9Zb1qTufbC8AiuiHOfMSo
UWAK/CgX6w38D50fnRRwXlELJf5t+Iov/WmMRYyZW5IxH5fnuLSm6Y1rIWwFiCNnMwHlnGpi1dx1
dwT1hAGbyzyoxwndSRSIhluNlVGB+00X2gQRSQY+TovzTdQsWDtSR+KEYIL4F18K+vvIzmmyVC0h
lRebsPsACI0fR2/92S9bcHMaMcbXjox83/3Dxap8pa1t2rHdcXJdO30ymT6d/lJLyX+Pw/EXcLVy
Lle0sFTuE69t9kvpvPapnqYUjn8NXaYIwgqukTqndAymHP0N4sqB1qax3ArKQ/BWho3jlBxoGJDe
KZsS8MDjsuZ8lcw+3UTTT0scf0AdTsFGSHE5yNFoBSg22G12wCe6lDXPBdjVmwhV101HI2rdFn1b
lxHlAJXFniSJvWAi7vX4VMEbGUn3Z81qw1Cw4armoTfJh3JAe521tlI1mZkfJCbgV0BbMAK+eAc3
FXnjjF4LlifNL9wVkT7S9Rh8Twdn5w2sthfzKiAns3gVjQUgPFb+BGZBtC5KOhlg69tGsflmZo0a
4sPVNS20R5dc3SIBGwBwsukn7bQOgZkJPXMLXf1r1QC9bhEmM8Mb44MHjgG27BHJk0Vuo26N7eLf
hQGBLKcS5U8ek8GOZaO2wm+AhnBTlgo6SrcsExQvxAKlZlsoq9aVYEjckggz5bhuh6m80TMYiWhm
gWpEu5l5s45KvkF2s2GYVAJrEucYq4SGF6ELUAUjhdVIIoasmZgDucbUQOeFJstgghOds9pmyh92
w/CLUbe6vmmWr59rIgmyZcTxEVCq3VBIUkowVu98seJxGw4Ys0mTGc1QgigKAWI1T4hyTcedC9rl
vowST958xYJm+S4IFDtVWBeOZMdzktZDKN/hrTJEizjDsxXGrnA977G9oDLY2mOjirZH7qzoizlk
o5kVRu+gA66+jGG/MGNJaqsAQBGHTIwqD8u+k9GEoCdZlroY5FwmPw67sych2Z14dIZMNuJMDhW/
hukfIctjmRtH1/j0KFalkBxjvFpuNFX6Xv3g25BvsJHxcS85O/reBPyocUsvDRc1nimtu0+UH6vu
Dkmqb0FkSDVcRYaruWPfA9a0f51qj/3sMaMQ+/ISz/SPSH3/RZesRQMICPixlwQbGZ7EowmRqwdK
UEZDxGiDewZeiPBBEuyimh9ORSTocCrVtF4kZCx7t/pUjSKgJTiztVfI0NJSvSImLmFik53CF6BZ
hJjnlh5+7Zcibl1zJyx4prj6pCSA0Fxiy0/qU3RoPz1BFzQfIXZ7c8lrgcVZfAnhE5FC9E9PREER
q75n2CBpHKgjylDWo1NybHSr+cjTMfoCQucqOyOwqvIm3env3IfLn7T82mVy9mCvFBKvFIWiTiUz
OqialFVdm73ApWGEKv3tHW+nEv99v5wqAzSfVgbdSm+grpPJZ5sMoqqt7C7Zt8mwSQ3xJOuuw7OM
KwhfX47TUhEzIon5ZbuQVakc9y3qjfZEyF4OLycZKtDxmbrU4o/7fl8nX9J0ZKG75248O2sTfaV9
rxPkNrFafOO9lKcOZ3fsVoALcbMIB/2nkty15R6LZVgITQDRrIiw0kev2qfHv71f6Vg5da4OkcLT
XrF7joanApSnywHoBqOc/srL1OlCguSFG4ZOnzXaL2lgNMklCYPURwc1lSykriNnV+D3PElDV73R
LlB8uPBj0bZIkLJ4o8kpT2VurRPCZTNNr/7YHd1AoM5qVDMZS2KdOdbM0SCW+JbvzhbgyXC7o5BB
JGUmpbfIC+aBgrf0qZoX7s+Ut0rCOuRgvKwjaWJ1V1SXTZ30QCnZVtAcn75kMPK6S19O95wdSyFE
NTZU6n6Nelc9mKT2EPrfc93/oLwRtldcfKWWFcv4FBfkQDrise6cIjSCZ/zukoN7oLzYMiCSWxCF
7PbKKTh1VfrAKJYDuH3kD2N+J+Ku5fL8d3VBK5uCKY57/E+Fva3juZKHsMbVT0K73OK9T+U5TgDO
wWLs4SFYLgyoL6yy3p6pVswwHy1EkdwE41R+ktehEiBbfJ6S2yQl76UMWh8PFWASqztMkKd+cMVT
kKHg8Fi2+iE22hBjP975eTubZSvCHRs03FeZgARuFZwhfFDtFLZND4o0FTQhxtck6nL7DRDpeY0B
Z4SX0dxzZV3rpSUJIAONjR9kL8hewbWNfQycJNUpWtwSI0kZsVuUzav4y9miaF/UIq/BfL8U6f2k
ei22t0tUYCBf3s3u4S4oTxVVMf8TnthYUy3MVMkc/p9p9c5cZyssnZLM+XPjolbqecBUIAhZuDqy
jQFH3ktv54y5mUnN+Ngyuvzf4BnLD2MRbNFmW4Szdk5G6m9adW1SdoFZRvLIFD0odgmZv7yV5qJ7
6t6cfIZfd9hg0ySlqMQwPlM49eOb+qwUrBAIbQYFeDBDMlV3NBTL3hP+pIJFHgXY0Z+piQegIMdi
skvZMxBhFwz/S1fBILy5XPRDzkNd+Mizl9JiDHJwFET8rG7heQU2OjPPV3Cho5w4k0WqqbhuMmt0
BT5AnMBy5cfU/z+LUUF/vSrj04Ii8m+sAE1cno6FglsD0hklr7fGgxqbz3Vj3LCvqbOG5L+54OLs
rPP1dMcFL+JyXmiK/cOLyWtDtcKDveZCiM1EK7+cSy65DBubpeBqDfaneixSz+pndSSZjlyNWcln
RKY/zxGtE3lJivrTha4m93r3ugLExAW0+13nOg30VRZfx7aDiutkHmFGNOgCzgeCSouFa68awbdA
Bv17FkoR8lFZl7nA7RyhK9b5coOp1/O4+GcS1i8fY7nbz8qD4gWeFzNTtH5YztgEi5xCyG6HRyce
t7PjT5kPogIIEcGhSYZnMJWF5oVlKArDE8l2hwiKS/B2fD+SvxEjLRyhUO8L9dn+pXHTIx5Us4dr
50gKwyt+LmMdLp/IzEU0EZqK7oKat7peq4Ss5jyuXXvD6F+levw9VRpVIhq5cB6es+Hx0Gr/pNtS
MiONQOvrxBAg4ZYqFLk5IsVfCbC0MSBNW3aXC/i5ukd3SjdTWZy1L5LKo56aav1wk2+6qs77dkca
fvjQgepWMB2bnyLMBU60ngvCVSeKVoXZbL2OY0DBui7xiuHAv6K8cSMNBbDtDcwfo/I7tMX4B1RG
yM2p6eutuUWVm4YX1wXpYg+ZFfzWuf/9sewXYSZ9bFBnu3lmvbpzTq2xsxlIo+53u7m0QP11c2kO
9bT1oHJdltv+qbbZg8HSQ/tTvRKtzJP/ZgEk112OiWvr6VtPSQRmwONlr9ISx13+tYII6SxScvDB
zmwnqUsBPyGty9L80w+x+59TPeafAU/Hhdxyzxhf00eDy/vJw6ghldvmBcvGxVPLHsj3aDOgfV9b
8SSbd/nStgo6FdTqHfiqws83885C9+365lpegUNn8uPe+QpUEaEydbMZKLRvsgq5aT2JfgD7w+dA
UV1Z+IsC5c4sPOBU/s1FLD/0hLHtgnBehGuxXOUMk6lBNiWuiObH7x6+Sj3w2GlVQtVhl16tXG8O
P999gijpjTD7EU8HmsktAkImXxbY9xSz1v5CC21BkhWexVDq+2GoQOFlrUmWBiRysk+oXC/OZxuX
fpU/nfBCw3A+R7AHehTU+PZew3uDCHBp8HZQc94dqsZLbXtWxa9nqBSO/64wxnZ/pzoQ8y3epx+M
hYf0ZVUPVRJV/QnK+bLUWNjcDGqp3y+27b7Y2Lz45k8Kw3D2O/X8w6kv6XVK/QTyxk4pZJhgk/6F
hVUqCCDW4Ho5tl7idVAglWeGhrFUzzYx+rtSIq3cIk4oJekohiF4LnGbyRkmNwBhjLlhbG4m4hCd
ydM2ljffbK+NE2xI3ObaMzUoj9fW1G1YK3e4YHPVa+R+XdOrOA0Ff4cJjqgdOwNp//l9vaaglXEk
hyYY/wq1FgvBpZtMYxek0YzX71fTWKuwdw2bPJM9hXWPkjOmwNsjtpNoewCI+Uco+c60Qri5oNDu
lIRAgdFUNcKmXB4PfxqFYkkY8nKXJLP5bEvji3aWoWf8Wq10KvWNoVeyRKyA68gOF+cTRhisMPvR
QDm9uT2Hgd4fF0vkAdnLUihTFFIAAVgfBOZpF2+E9AKXJeofOD1mDxS/4WAKUkC5Prv42UIp+b7u
POLvUtPobP68xdoduZXJA0YvweDms6iL1i8stvb8XlmLkWuuzfRkYmAWcWmsDxtMYhsRAVizSkxy
6UKoJ1IWhUts5yC7OTCzXgUNgDNb8wkKJV8A69ALsC7Y8uF8I6Djr4sH4ZOOyj3lTnMzcvOL0FpM
JkZImfGJZCHMI3fwcWGlqzmRHr3CYEX2LPb91aeIQtHzNap7me0EVYKLOMqHDcLhaQxQNdzrrSIW
PbjpookcN82jWAEWVvyuxhQ5wLtUQopljCytzP1vcGkzKogjdTBK6dfsfwtsJ2KDaOgKV6C+M4fH
Lk8v9yM5TtoMwbLGR8KIkjvn4PTPsMvQ0RM1+MfKr0DUg6QBIi/blqlJSaTF1FeqBAwWC3x786rk
54C0jqVFeZlz8gBpxwGrA6JVn6lB/Dwoc8nefQep4pDgXC7NYACzy09weFua39WGGs1R9mNlrkEP
8GfF03tdtJU1DGLFQhsX3u5Co44hscqSU8iexDTlhfyYOgS2Lz6rOfOA6vowHfmTFEv+Z/A+dSiW
QybnykWbPFhA5rM3FajvzzwsD5FX51O1JvFfwBvddT1fcBzgMOOnGzP23mj32Z0EHlbvZcSTR0Tn
aXeePbxxZM2gRjCIZ16Cd6DX7J99u3yD3tjfhOGebIUOpn9MAITn7LB29+7gLBZlBTh4SiYFtMNf
UXkLnjgOf6taWrHZnSb0nZsjTpux88Lbx7xgm9s3Hzo88kcWyi7AT9GcKYr9KtdcbNNIyBhXLNeA
aOtT6qauZ9sTiiMN83Zvn5qLydh2gpYsfSKii+XNK7Z7CK0ow5CyFlIv6DwNBoLtsPxJFsWaWp2O
DFEBvaoupajZhMjxa9Ql1p8KdirUYvyXaq8ZT0pvaz9qYbICu6qVuYXSgQePEftD0fpXENwNGZPP
XEO9Itvz1d1t45WNOqPe6Ht3pSc8PIG0vebfCjKojLb3lvfZZaz0jChpm6Fy+xmVe013rvzJin1d
9KS4ZvqkeeGrkRSb1IHuGv0g0NUNQCSDKNdOXvo4fHcgek2hR49TnEtWKG/edF5uEBK/b2sezyDZ
BCwurLYbgYuFaiUcblPaBDv4eDND4jS/tYRUGpbJ3bkBGswd79SqY1LuL7Ni9hyhS1lh8J4zuoy8
AwavtucLfTCUjnmnVNBe0a3XppRksyfO73hKd/Gm8pElO5+saztlFJFQYaoMvk5xbgRdDRyP4iWM
wlFHCNhvY/MudZMU9Qt6fqayJWG5vyH2qKBXLkkrQvfuuFHNF1RqK1lfcYsuTp0Q6tPTZ7a1zghX
gN9doOvv0W5nOsxlNEWV7cjInr6UQ0WJWCP0eKFmOmrx1qNtUv1keYWSzU8HPEjecfVgovy3WNmK
+5ogF2743t8sSyT6O+YR7rqWujF2yFXpwZ4y1cjxsl+Qg0SF4f1QJkQoR/e86ygpomibQ6OFQR27
fJkldfeuHsl9zSKQnw57kxEHVR6ittPHwjLeQy5ucRlGNMNqkQULnAYik2nmQbg0MkRk4cXX9gtq
+3lJTyCiCJpDNd0lIhB5hjyRU4DQcj7DZeh7eCNjeYPUJofjxZ0+1flJwGvjTHRGGUKR/yvwNtjI
2FIJ/vqdZmFPTUe05417nOs09XVt8vo+NvyiDwqwRuDckPsdu5tgPv2fipgYNE/IO/+9FvX+Pa1D
X7Q2+A1uw63yk79/+Iy3cSMPwLtNthX1i+6bq18DYQlEbRFp1CFeF6yMf+J37+LPUoFyU0MQQ0a9
iRYLhlmQMzyLuKViSOUdplb0ih6RGzf3nz53lY/RkO/eqBJmCkxVoUXqrvf/t0Y+5HtnVP6ZRnu1
WKhSe1n2EYcj64EfcOgD3vIObYWbz70CaqnacxeX9mp5ZrFjkpFusVq3ikKS2WeJHAoR4iJh/Pui
Mjjof6z7JXjxl8Ri7nFwJj9qq39r5melGpTP10oAa1eq+LztETxsUqJRU3PDq0IJa61AvI+OY93z
4G6iYOvQU9rKClj2Et4F7jQ5x1vmSZd8v5gKUViNVwm5kc66FUuS3AXblr626c/6SEc09IQOI88L
IPp9k7uSgqq4Ap4sJv/be7EClXSRGiIGCJ0YBTkn0Czzrnv6v9mtQBMDuLNZuB1QmCpmw2yKfdFx
/L3jhQFkCSmoHspx+boJUfQL7aP5qFya7lk1CYFl/o2giSQrO+nfR7DHyVd6A5nDbg/0LhOuOxW4
S4lrcPbMt7QoN3EFURVzG7e3eGPmggj+Wa0c80TqWSKDY4iNZLFTGBzMzFWmpQoTYuj5YBuD9AG6
O8rX/0l/pi6QCumGkPlobsZBJaKLhnOESo4hjQHSmbfk4FdX+jL4mSU+yltaLFfP3jnQ0coGNB5n
7e8LOhpLfCIX3MYv6JeEJkPVxNfNNzg/ViaHyRYLdBesNJ7DQoFHXYCn6ZtWGs3duyOrbiHaS15u
iCaKgvsk+Fl1X3OAXFOziMHxlnKabTWSQWWKpyGw0Z/NW4UVoIgOXRIiVk0o7FkAQqBRduG2en+5
ji225lScwRF44I6NuVDDO1GuYXEfERwBjprTwfujkHBHXn1Xix8codyC9Vqh1asXL7EI9BxKvt//
S2Zk2BRv2Oc1nbn1clDPxQce75aifNRoph6um3MgI03MD+7RX2UF8V+h1OZ1yVmZITQtVKIw1IJY
b2WgGvTekSH+CiauVdYlCruYjUtXKoOjJqcYyN71gvbHh2Hm5Ym+azCHF3bOdWGYh97JeatVvWZP
WiFXB9PMmZHRsXhcevC0t3NwGk+exeHYBe60bEeXGhX3i8NMNZcp2lQqq5y0/zHhYuqKiz33iiej
fDcfXNSleHfTYVB4hlMA2SpQAaQ/DrF6aqiLZFH8M2Bx4BuO9dzhVutBKeNfL3RYfmAZ8j7dyug3
WkteHAJyGBDAiY8NnCyZLbZ4MPEZGifqn18RcCC1rLWnVdIqK+tN13MeQvhonFBOl2fFRn1duPNc
IIdWTn5DdXvabvSu8hJKlXN0fPkZO/Aw0KQH5szby+1IhG9UcSxS9HBZSYh5lQCk/Qk/4mt1k3vG
rqRxqe0wqX93IhWED7UtjH//eaWcSBOJpwXawtWdZL9rPOHJTeS2wn7PdRFgPUoiPi4X9DNChSVP
zBh6A2Uffs+71gaODsXbX8fXqZ1uvCx2psns4gpPAZTM1u+t6GaMGbWkWERVq9C2rxZAxpF/+AS9
4+thi3xCOeeCyZYNahRfXDzwSARZnkj68RYCJ3SzUqcC37AEa39cPaYvQku6nNTM3VmWr2oYi0sL
mPJlHRXoWgmbTjBjGARSX6V4ZHQSu/8a0jumhLTlFRcX6GI4n9ClZqetiSQ8fAvvqPAjJco9wQgH
Vnp2QWlJkvx/fvR5bf67BwMlkoGmAhM9lydNQVGbYruE94rDkd+3IdfBhE4bip0ufFPwvziHnFW6
1Faj8Gk0bDX4fwT8kNlKBlCoMx2xbTviCCcmWPBdY35hjc32BfuPz+HeM1LrfltuoL55Gtgoxyas
fljb2mxsAX1rYgdB5IY1X/eAWYaaPZoMOjikznRnU/AA+o0gonXO+sYBr0pHX25Mv81SnFCjZm85
5IGCdhoHEL70x4SNImSQUHFSRUKtkSsnFYhomk6W4Wr7XMma0lIhUkTlh2bqgKtPX4cqZVynxQXE
tuRYzcFIVeYQmVxEE5cghMCLKHvFbydK9MWFGLe56erlJISrl9C31Q4G2FYhzztjmZOvzXwX3FW5
ER+4LI9beGId1ogGn7aCu62GfSch7VEzcLi/7LAvmxTz7BNz679H9/Yh88HstqtjJy77OGaUeIof
4eIC+4J4cptNXJyZ7kOpLVvkSYAV0RrZkYFCjjC1T8wZCuC9f6Y0Vq+FhLt11rQmPvWAlv+lOtQd
VOa93d2h4CEsF6B50iWqrfg4qrW2ywj1tRhfm5J0/+xOLql2GOsb2rXKBZP8roJJj1qSQZkh5CWa
Udv+E8ngNOAhm0/lvIgcfVqvVG1+9chBih4gTOtNuV0h829gE3AusiJYKIlmD1bPFa0dtWfOM4Yk
JBGzk1ITYF3xo3+1gpDEK5VgUy3yT05ONDbzVnPU24TSEOnecBSrD3ljFEovKnIvFo25y1uMzdGe
eTz8QuqkE8MEq22q16/FWgPblqMQw5q/enjBjI26PBJPrtMvGh+aUrQr0/xcw2gFSN9KNu+GAbIG
b/0N73RT79PhFEOxqCh+ZXBaFHDfZRATdTj+tljq3ZKm2hzzDuFxD2RaFOQ35/WBVuVsL/zAqMsf
zjNxC8C8qZkg2e8PCdx3mV+VL08toxj8EtWZjyrco3Xt+cXau4LtqG88S7snegTmVC1QNxYBOQA8
4BlqUWFJrJL2wP8m65KUZCu2ZHMTga1AvhzFeVCsj6kFTlhdTZydUyEtuMidqm74Ij4vsDaggpVf
YUhrWyPHzNBUPFtK7Qqw5ILMCQ+GRokuel0fmKTVVXBGtdHjVVusV0C6o2qPshggSmv5laKptkO+
olLdvx8wHkwkmqBYJZaUefnHOYpMM+bi3zjDRKb9EGM6W/F3VhdM94zXX3aD/q/J+huZCJlY62Bw
4zSn4ynrjlU0y+hu3YME1Pa+iB1R2bf/97TdCwrrq5sbbDdaIZNEI4jjR4EaUunfMIwfC4rXSAMz
2l1MHcJ4fUvQ7RWFQ/NYqe4KxY2hu2tmhzdfrGffuiRDlXOmQkbWzoYt6yn8UNG1rXBe9pZaCjGS
ldUV0M69w/vNG9U3IPKQzLoa8t8k0NBBhLni/BdXArENlD2gHIapcBbNbjzHLhhJK5cV1eksXM48
TJoVd4QHUbzKnrUYrWEZpWetZo0TJOuK/vpBgVHEpETcDm214WOvYvDKRWddQ08H+9MaHJ6gAPPw
rsOUBKHmiciSFq4kF7CWMzGG5IC4hUvHIShDZZxGOeyhvogx87Ww7TZFaC+H0qGkuAoYNVJH1f7Z
g3T2dwk9LAoT3fGsFFMmzzT0zF3tGrKK0RbXdkJHNAnuU9xpv+/EP9df7dYTWD7rAwUBCMMUx5yy
zwsOqLPSibINytYBf3QGGciOgyfByCwClzuMLFiuXTVTfW14ouTaygUXbGsLd8C0gvRx96yXio62
4Hiom6hTaGVYO13G1wZgMSF7ot7OTjRFNY0C2ZLVtZoX9dwMpEsFtacw47WnVeM+hfcy4uMISrOc
CMSRMNHp/TxjpzihND5BmOinn/uXqMFNFOQdaQqSV7gVpV1Y0qaAUsXx7z0+H2k2rf9cVAeHJh2o
Snmhd6ey+eaxQfvhdc1LJV1xtUXKTB9VeSD7iKaJSA/wJwl7e2T3zptYiLoNxLtW5J+CQKsEW1qJ
gbMOUtCnLfcN9X5ZwjWeC538K1Ilha8F2WFpc59xYCRHvabWpPyNLR0i2LcmivdhjVkkF6LIPeVC
tX7e0JMAumZp37TwGZFVr9H86hkAo7ibpOWyqfxEf/PDxLH5rZ4zmps1Q9HmCUZ9EEJhZCNXAeFH
6nPJVJyb75J8fUFAyss4fXvyjZOYX6G7MOLbup6TVfu347fft2tFibwTngNA8sAfTDdGdJJAYm16
Jqmks2g2+eRX9jyBF9uGpowi6JC/ZNMR7bOh4qquAlMMCfIXDrIsn7+ecOlOyBISctUTlS7vKT02
KRvzJS4U6GapKppO7KmZbBTcULGrzhi2/qpsgGWa+SgHZ80Dmw4mwBn7Xn3Ziuilr0MCL7xm3hKS
wJH64NMoN7KPBcoSDUa2uGIRFuwW0QambuoF9mkgmvX9ou2YrEAUzXOhqJ4MNm9iVr+wodVegZFb
Vzk5Vy6EEW2t/inCcHgFaKpBw3ft5jThyfZ2CuviTqoObv7Jfq2THkCvPmdQFYvvSWKz3z+Vj2ii
04VRqLX8LUttYHSaO9AbTRIEAGzSE/h+RTsi7YPoJrFRyNg2lyY4OInnntMeGywjAX6dqmJXB7bn
BxIlaV7T1+w6Z2K9mMIkT9apkRJ56e8O3s3wJ9mtOyon/RUAYBBgiSItuSQ/CQfmFdmwu3NbCz8E
m4NBrG+dTs+7nRfnYdrQi1qG2djaVSFzD8khtmwNYIdssLvqQrWU4gGfLXySYUu4CJj5a9TJ58UF
RHWXJ4j3ExeJS0gtMDUUcKCT2BBiiz7jBP7IvjmPPLNBAvMVI+kaH02kV9Qbf4nucnbhkYvxEeIO
XTc3p061DYfvvEU3XZVD6El1m+COxIR+4g0vaenJtn1U7G7exT5WVhHpclZhj/5lAVj/hjwitFcf
KWRrolyKiQOPMw448nY7TLwGu9yivpPRPRO3p75eIEbZqmnCToQClWlqmLJzPk4riiiT/OU+W10X
f/RTVRz4K5Rl6VmOJDA/zuXDGULQQKwaKjOUi6jWi+Ov/Hs4okXU/jLvFzsD3jmp1jqLPfN5sJjL
OmL2ozriepQPm4EpbGQexAmSRsyjQJ7RJA4SHtU4cgZ8HxWqHsO2i86FEQ4yFVOe93MqNNUbhUV3
AuIV/ikY30+dm8R7IU0TJp3KlwjvSB070ARskqnb2qXwXoaxB4vPuiRVyv95rQXsDWih75MSGfFk
uDHcrZCzB4BWMoMT8Eo3634FhqqnBp4JNJDc3Q4F9wMRMwj3Y9/hrg2y//DXhpkAl1SX3SDoSeXX
ZvrlQToPgDiQ1UfXVkiUQnsihD1T1K2rXmekmVVTYjJ1Yy8lLZqrD8BhKod8qiXNBAaGYTgfmDjf
blb+zKP398YXsXZsUJ0kR0VkTESGM4Jlr3jZrt9rcCGaYMFpUl3A9ukyUJBy3o9GtvKBHXMzuSWZ
fimysyADkABTcG8U//6W6ir4Fl09lJ/ddNRLtPvVJmVKDh1Weq2WvUK8tCmd+BEHaOw2cbNWGZbI
PZhg963L2D+5xJAwvT3Z55I/rGShv6fb6jiA29hVso/wfjEQDjOfVQIRX1fhsKkMuwzB9GoZtHBj
Iii2OrZ0bACiYABxkTvVJ+MQfmzxZtzbR2qFhM8cSLXfaEAhdEySyMd2neNywSvIPgd2QC8mX2V0
2Ma6RVtr/y3ewl0l159u/3ggDHvLfK9KCnVvh3oPOT8+d0SQON3yStiwFx4bQdHoIYYwbLXOS5hF
hWLjZeKj7cIN7NlUzEMlmTOeSrhAWCaNJ2Ng9hwYLYZatZunmWJTJYiceO5EZlWwSHJQhuKsQ57+
ZBR4bHE7Zb73qCGADdjKPGTLsi2Pu22xtRClqgrhU1g6WFGOXd8fogQoTjpHwctcd4gNgk6+D9Ee
CUTodT9d053wPGDdsExKpXD1AO05VrjaVg93ZotDZzIg9/TeQDwZ9eNtuX2HU3/Sg4n3w6zmCT9h
aSrYRtpg6MA3Nqm3O6dSIFnfiAmZjnvUL15ToXfKfoADVndJMm6+M1Nf30sm333k/t/fHd9SD3oP
X8AiPw/p76vF61tLpONrGFu40d9JIdnfN1H5a0+IBERKMLv7tPDpBLw4k9R7pT0QUIBGJS2/adE9
BFsiQ4QEWcZWnBuj7/oaf5rHwKXHlAAm2XAqxCq0AUkMDhZApNTmjJatHU9NYqc9GSzLFPgf69Ri
jK9EPzpxtKdx+1lWwPC/3LgKtF1rPoXWITHML6bD0Q7CbluyoMAME8TeE+QrIpZRyUDCFq/C3em3
GOG/iwfbbn/pR3U3oOA2zb+4SUUV3srNRvIsAwNOcmHvpNltF2i2VUgJn9V5rQKowiFdULRjLxex
EYlG1BTsjFHIygTiJ8zavKYwgG8Bg5c5S+oY9MLcA9tYkuqw3azsFekbxag2q1UBxOJd+2p6WyAd
o5FbRy7ftO3EUIMze4EKckz6PTJ+mSsjWeBwKFel80ZWC9n6fKluk0BZtrr1qAlxHOmd4PCd3f6l
1zp60sEJ68FphM2V103ZsvI/nkx5hiq7CmZWvrja6VaxpIHDcFWk9XcrkkQSBV1tkfyyc5o/C7xB
8Y8vuoW/NjuzJSVzJ0yIpgBQmS8e0UW4/aXVdvPiCF75didUUJGFBxEK1qdbSUPiahj+MxkriwEB
lwkLuQTyG2ksO2M2dbhXhdemqIgtB3VRcMkcG//jEIQIfqT1gooZwMlmVI/quf4rx2vRXjQ23M6M
DBZjG+aYZJVpj84EinRVTWoJhCKPgjFaSP2J9SSGIHcY7rjB5AJWg6NQsHqSw0L2Ccrd5NLpzD/9
MmFLtcWQ0ZDdcvN+6bCN2L2mot+kvEHZTVeWFPjcW6pab1fTIwbx7tlSwoGFzvfar6Jc2qE0+R3Y
ds5Mq1zTeaV88KXBQNg96yOtJl3BfadWu6tdqXT+moowBaC0H0h2jYlXhVJRsTC2bdx6cbccO3wa
lpIiI9qPshPEsLKNR4LU7OgqY+JlKj4w3nY9VYYYU4XDv1TzZSmDJrXoqHPuNtMFGBNiwsJ1Y/LX
U4v3YaUBi0NQ7rUOgPP7qM78D0f2qg19gggOM/JaZiMp3svHotFxISM8X6/gQZMkaXMSDWyf1CQ8
6Eo+53pjCqxKZCixCdaO+jcDZopu+LQcjIeeYGM13+JZxzB0nkf6CqleXBwWflEl2MiraQu2ru7m
rlwPWaXkTCo2kgv8L54q7N0Vr984uhD/YB4lb23iu0tifJF+R5c9SqmjMvd5DaciOHwZwb5jn8fc
XGPl6Lpxd81QSTRmQtyPG32rftxjSGej67g6DFjTzFHVA3FMTzp7V2WPG0DcaTZMaZq9Tdat4Qm3
BXlhS+ItvPqUdvDmYcATSHHS0I+8asKSyvi8gm8NbdiSLnO5mQJlDoxEfNSZfc3Cc8WIy7tasAV8
NKT4lsCjLwnZLzSe8dC7shO/amgTFYxyFa5qdue8fj5VrvWvTJSbGjdBsWJP5XJY+yUBQPlEEua4
Pg46r7NA2GD0Bf0b6Ru0a9WSTz4uiVFbbfhDvezUSuHPLyfRKqhLQRfr4odEOYqfGj9zJlOiCp7O
rXC6wMYKV3a3jc8A1f9ROi25l4E4RQBAowC6ciLiNOcinjmugIOnsc5VTz/nWIknHsw89MTiKogA
s5UNtGRb/4a5bfxJasfyTGfx2PKVAN9hzx3+rFY4ro7E3jIumFGl/32YrkeIpzFg15YjYwci/FKZ
mfzV7YIhSFhVdFKwhVncIWuShJXYL9mGj3tA0n+crShJ1/gV3m4Rli2AlqB1sx5r1yVtCcLBvO8I
0kSn3Imhc8jPcQnyNPWFydZ/pLf6s5NKYetj7ksVNd/KNR/9b2oqaN9pvJ5itgjGQ7usDhC4/7St
0RWHejy/7HvOI9Gkayh8hzljYgTbiQKayADCeVMicIo18+0XUOpvZynUDlukGqOff1O4aPPhklLF
NTSi0yCyYDEGgtG4xhsRzSv4m0pwuNNtwbXGQuVdoBuUfKlFvbgNFLII3VS7NW9EES7zcVQ15I5V
AqWdOAh6CWXpHUHyeBEQBpFmjISuaO7tGWeSNhYInmgq02VFwhb/TKgzURMn5eewX7NCzKK9/Nsj
1i9nmJu5MtCpDDk0MjLpgpkpm2nLUucdFczH2/1+0NqD2ppbT3sDgfZybSTo/tBF/17Eb8F/KcHg
Kaz5UVhLpv1gitcjd9YdJrfwBuGhGECTJE0ChLKlQub+NjfF9tn8xVA1PJYAk5pit7AufnTWEDDv
7X294d5PuAXrQJTWa/eYgflgOTQhPvqvwuBKB4aRxgfD7A7wtxCjYT+oEYhdGU/8rdXMPWKNGaLa
KFJb0pXlEUkEZ6SrRy9VETdVvEpxF/M4DA8DSXBbCsGkiu+3BJg0+aGv9KKIF5cTU2nPcOQRbRle
Agb/T+uVy9+Ohm49w0xgW5tqZiTbdv9YcKwz56BtmmisSAaR9nqcDgm90z88kK0VbPmb80JnItfo
c2P0cb5I0fX9cVXUGJFCPND5OVZvruIAMStfuspQfvsEh04r7AaUAQA60Qcn2DZsBiS/HWE5vCU3
s7kTD3b9yahJiwh22+dt4W5fOaiShSdkA/ChbwfdoLdtFrGBhZGhFCGSfMvTqh/k01ZnCRasK9OH
/86Hya3YVaJftnmlSTypYUodpUvAwW8XQpyEAeH1lXajKrwrlWha2ZNlxkx/WXVWlPcOVgrQRB/B
qf3KHk/Y7qnBgmfv3+b789bzQKtgYE7cWPt4rZIjGbGr0PCvLXJoWcp8/YZLlrLVIYHXrpDi1K8D
DX56JsqbOWlW0vH4It3EZmzbC1vIpYXLa2+8O0i/0uGMgortIJtp7P2n5EYaVUgMXXd2xQLee/Nk
5g3IGEW3y4NXmU/hYiJd8AV8+POungCVdVYQA6GFojNWopDz66md8CaM+TWOJE75aGaPqh5Y8V4H
fYhxgIUSoDvNHtGcx/Md7AINn1oGQVdGq/sCo9ln+7ZFpfb448J0aCViTub6PFJeJHgre7KiuZBY
PNg/ABIrWembNFuJbJzh3tTuYBW7oBzrDtX0mNOlmpGgG6eBSBRh5lNM25R8rbtdAZIYSIxcX6sI
AB3Lsme+7xRu9sh17OJJ691IB6pUKbqISgZOto6SIKIjwROv6wgmmG4qisguGMF8EcEhqiMOM1M4
ncxDsInMGNX7rsPRo2bMihEPun+CoxoxIEzel837RlT/Qj6LskKPqZAtJ/mV/DCDmUe2K5UkL157
tk+seoZcn0s2XcsxeCUoPqXfPz8Cqj/C2n7W9VfmYIv0p0edd/dmrNQ7oq2/8y6MsuZw9J1RmcDY
tzVnfoZpvFIvmChzSep2Hu6OFXK+MmXA4MRMWg1SgrG2UTiiDWet1/Rxj+n9+GoIulXXWJRWUAXY
wZwK6RnJObdniP32DlbnmNWbwdggSvR125DdorbuXRxFlopja3QL7CL4BFUObE5l//2jX64TYBup
d8loMXkSpcgCo/VX1cQ7tNdwzA6OaI1DH6Tf+i81y7IKMhw8iZb5Wow/OwVfBHtRT4vb55tgAqZH
uvSBmHehVEOhEkeIvXkKkKKkBjp5/cDiX2VcLVSrDx54jaU301BDl6CrO6hrHzdrf0puXhOO3boh
8SbVnrEN+hK4yudre7FuDp7fte6IFowJfchkpph4zGPI3maVXWyzrcUBm6KkJtzlONzhsNX4OqYG
pnz+HvdbsA2x2TY1s8sw4ZWWXAc0k2gv/k/bjZ6VpsjFsrqWkE31aThXtOQO8fYYjky/zSzs1pTn
sxN2tOYDMaCjntOxed1roHuCckJf9CYmV+DdvPNi5PtsLTTsWMMBk4fLywxRxnNSpO57ug7xUEOw
zPoOec2/THoTsY6m4z2Mq2m1Xfmeg9ie2IT8Osqqri3v+pMEC/H/iC5Xce8mbkw8FUKotAMmLEN9
o2ohcqQ2EPR1vCvo8+EaX7fjxlLRpP299FY1NOam5OqIu23hhQ4ZR7YQg4awCXCL6hhsoiTsLj+P
4prXT6+39ItBKZzhmzSXZ301ZFCb66DyfrEQWowUjV8dPdjvh0LTMG195kGxD3NgGZeJHNZVTwUz
TOM2QcuXrKJzC7nk3hyBkKaPpRFWHA3ozQvazaSY+EPFjvDYEjQVjhJBYfkkpztKxM8UuDhD8iK1
STREotA4ntn4GzjfISwodVnN8OpjV5WVZ1JtINpIV4TFdXlOZsq/L+cvlHTrQXatKuqgmzEfn+xW
HDChOmlmqSxWMYyqWM97hnowCZ+6mX68kXcIBinNBlrAVmiivatiIp4eZDZCxDzhF1EZH1L/chHT
A7r8hD1wUleBiwFNA5V7HiIU+7Ysqn7WOMn2igRp7dx5Fsdn/Ts9V8hgR1PVKeiwJwGTsZB1dBYW
NZErIteoffBWZUwI422hdU6S8uHj4sj3tNJMeyoc5NY2c2vT4WOqFBONAT29X4yC72Wxn6dBqomG
cKaLa2Kh+Q42qA4J/VRgbNTI9NwO8fxF0sYgRZGOUqT5GY75gfpCIT/gExLoldACPrYTWDUCXgKA
sd9X65Pgt+VaVnpayS3O93PMmVTFhIqgS8IeCyaxX4Z4EkiJ0Vi6KCmXGxZcqCdsj8G8CcNM/GQL
m6si+S+QJKXYGAxoNM1nbRgfR67OuBcjHazp7w6rx+iMQYJ06AElHKP+8fjcv37lEKDVrsxXP+9f
0c9Fh0kQQjlWidVC0z0INwRSylX9QRi8bJdStPvVdryuzlzoWH+y6BCTRxnql/OY4hFfZlJjeHeX
iZEog1jImz+qvZOFuH8t/7FcHvW7rBbo4t+ptC2aBD+LVunygdWBnizm6Nbr9C110tcsRd+UyHCL
wXvT+lEqGU+kbhkyKMkbJctpTm4YTZYlnuRSDFkTaXdvWOCkp18PYNp2thN9k5A0OCj7qtybdeqb
jyoMuFa4K1KQkF9tyNIJTaG+cHC2TuIDFF/WR2Sq4UbRaY3MPGfNysYhGLedUteqOYZF7s8Wzi/b
ohz7Jb1WHUNQlHdGA8APc8+nE/29vca10H6BXR96EPgjm65F+zarb7FhzBF4+eDO5XqZSckUZ5Kk
wz3LszYTpJ85BB24bTLOxqXC4ITXR00raYotGEbcndo5UfE/qS3QjDC/qDXsOpsxqeBDzkLsEMA1
DLZ+KTByrFI7I3ms9FQt7aMyfHmsdomLrtvgrLnvJ2UtDL0v2DO8WVmV+jvYjjpbzshhMN2kzn8n
Ab359SzFhYkRCvSSAMG6naJe6MAwD+hEgm+SLoyj6ruvRsPUeBEpRMfwtGNgICoYGeXiQT8ZrqQn
+lmHGR1M1eXJj1Yc4gBL+7aHlHYQCNiOQtHmZwxvpTnoZHqaYB/HZgsBZJ8StXQksUQZ7J/xboLt
+d+/9a9KiEHpV/Htm72j1xqOT7xekIHC2BpMsjGYFt8vYWAaD8PWUiCWuuBRjKFkeW9Ju9gNcfdd
/+jQzyeVeRycMw2JKRWxQEGgkIBN5RN9iwHkySjEGZNWNPkgxt/VwdG6IfpOP5/X6IDfXhw3q4t/
f7VuRj4kLFOu1kADCVrsoUpmTMOb4VA9G/44CmoolXB9UgLLFwKE+45XKlibBZXHUljyC0pebCvq
7+d3sHwLFylXfUHJdxLYHHadpFXk0D/OuqIu3Qv6RLPHMwZ+PkKVZKCya5Ac0m4rfPrsYz9xQMZJ
75MYPd7YzWzUQOMNyWls/6sE5HZZdpExud0VLShJDbLeiobMR9IQ8hIKd13vpVtH3jMruJFPACkK
9J1JJbqE0LVsSxwCouE4t1GgaehYjcTTUGpdaVnxKVvr3ywB69KAEZkfhl1xU9Pzkhr9JdTz6/KM
iOrHt9wT9+RYXmECZSuXEhJgLszauc6oZND0uwUey39C+Bwr4G+q0hCLI8EbueAfX/ssYFsZ3xwo
f+ZxuE5foGy5SUD55xHihOJPSI8nmL82uAJHaqDCjtmsbMScAyjuLsvZKm1sFdw8DBQJbeEUKGp2
8/P0OluEJVxyYl962NXITZm+0sipLMoQ0cCQY4uzMbzSVqOrvmkAYfJpPHPvW2czkHM9qTS9XRxL
7ekVtIxOWqOyBCe/3/Gx2epl84ZZvY9DahGbijzD1MurTuGHIGBipdOIxjv6AxzEbNu9phtRLzd3
utkRl2FahnKx4IKYhU+l42xTPvuN6MYFu3C2qEvQBXqmBZHUMHS2T716iCIMUbM1bNuAoMyUI19P
IIBxZ7x6ky8vTgTJkOEwT9ycnuNnfS9Z5VXV+Wf5+xHRafHla236wMEVqDYWyQIgyDmDTEUDHVH6
IqMPdfyUjICxvSO25pT4LI46UGbdOikU2MBO9+wOuzr+BGQXEYgXRWlpXzUtCbXNNjnY7el+ddeW
nKD/hiccehvpp7ZKIKv4znl2/UaTmncK65Hiy9kOl85W785WuttQD87o2oNG4urAn76OyNVsmtdd
rcLu6WdF/YYbPzCaQPbnuzYdchjw8ATYxsJLQEFzWvkj5+B7223FUysyIlDRGC8iG9zWl7h7E5t1
f1AwQlapXWM8GnA1JMip+LQEscapLKKwNp0Lt+xzvm3SQc/LPHLhyeSdlVrJaPSKRxHFPRMx7h1F
nn8uKS7kENe0Tp9rU9NsZbLuQVEzN1DXro26ZKAcQpVmhR8Wv83D6NasXZmufDP3yjAxa+1Nb789
v5Ttsz/DkR+6e3/aDVn/nqyWtOwTTQaSUjU/HXS2j9I6XgvKkKpPvSDUNLyVQfON9V8hrYLcGMI6
juQ4Ih612GzhHMcW+ciIMpXYh+gq/sn8DRYuI6JtP8VvWXDeEyXWDj7bFAsGqMbvhDWOwB5Lf8rT
5nwQ6tHDYT81HWHTw3JQKtzfmo1h4p/d4lItVmdSb0kPD5s+MwLnSaE3tcx0lXCuM/4CSe2JB7jd
enKfRKKgDO1sURavSyoU4BT9l3KtKFGbyhbZgoyZd1LpVmT3Wk1+CJtjP3XmYtcWZcpheC8AGF+J
mmH838wjJS8vG5jo8ApaLua3Wg4mLDG5hd2jEFNmY1EhiwzgyrXwjBFjPsDGKRuZ1sJcz5e2gfao
7VvuvP4BgDrhKqMEKmbBhmHWLTPHFCayqzZ/ECaOK5hm2hpz0zAADmg8dOyNbuQlz6mQMbk1LbEc
ApOrjKLg+ZyRX2b5Gk7TuPqnNWGGLY0TkhVT2X+U6kvyFuMfQEamtxB0m4y+TIGuxsmZz9LPu+Vq
XDms6czxI0tzhEhXm2hAgl1qpOnCZTgnZ23IYPeGsQkTAyQfnE8xt/Cxmz/zH1/uDNJh3BsVHtsx
dqA7dPFVp0pWKU3GISNb41sj2boLLVXpvYpy4Yo8jhdXNCLt9g7SnC1V+3DVkI6UbE7ee1j8bTK2
NIEcXioiIBkeR2R3UfKPE7nr3dP287K0m3HIupvShr1ms2CWPXtxKWULIeqyRx0/5aoawtoFD666
Vq0G9oot75FBpCNyxpv+HHSIBnbAuP6OXXQAMgcDH7MnppG6IgpOYGXHxAoGDA+qETcNDHScxwid
z01yf6Sh4aXd1JK8w3eTYi3DLeq6v7nBcFnknmEZW2q6De1CGor/3SdtmYUqeJg8yiAILa9TBWRj
8COkID4P+PTK1xRrQBpCLsYxqT2UNNO5plAGNbMGllgRE08h6I3XMnfl7gzxMQ2WYOqUcGzttALb
1+5qvW2EWIKF3F1KW3OQctjHgm2Bi5l0n9fSVoAN1iScbkiTEqFI9ESfvnw7NEZZlRQuMPfPRMoO
Z2sBIgJUyhkdtzVJ1zOo3tQ7PxIuWl4WlOxI2AA8xQX347TTUsdIOWE/ZMVxRyYxBvFMeGCyjy3e
21lWmYzM/Pf+lJnR4zmLWD2mE+gesEC+ulKqnueOJW5a2SSCYxGZPq50oGuu/fj46RFqDRSGCHep
uC5rU/OX6fatcyDaFYCIK67zfaH1DSSaSWRvax+X8192SnEtxCFOtE+0LgRxVVGFakZG9qXIFMJI
Un7Kx1Gk1sy5YR4TO2swo2mSS49XCIMBIB+zmX1uZyVs90/VhM2LCBoF3JGJfKX34L8tLbvdRpaQ
9MTCT8Yn4doaVV/g8GUptKIxioAsXjjL7RGPIVWFxbtZ8s8Gg7+/hYr69hcZ/EeXzv6GcHz7OOWA
d8BvIl/i4ep+r68mDyx6IMdQKroStXu0wg96UjfBVEQqxHx65i1GpSsCdPun0dKoaxqkU1uea1N3
TlQnY7DzpyN99yy8yc/mzyNj+QTlWUoYcz0VlYbeyxUD4pLHr0fZnvCd8z8wKy6PvqUKRJ/SNyON
p8co5OJdvh3DUjvKONzrW1oh2+NTmadxllyhZ/J6MHdB2KfwuUS33XEDJmHlDJjNrrphWtF6ngGq
In8/mS+/yJScrtCGlMZVxNQUVYM9IUGKGbUCaS0j0N0fIpxmm2fQHBDZ39ipqK8+4IHJFlpUxYkt
RdOXNDSy57nXdTFeDaFM5geZ2NenKlGtbaKTuwe+huGRj9JeFMiTLUmFP5rrGYrLYCCDY4LhPs5z
hoD02AI2qZwfEjB81QUOrlFBhTit2BkFzJThRb0wR1/A+4ou/ItQh5fqhAEQ+AgH10+FRLezOmTM
9L02ti9AuSsg6QOxWYTzT1UopuPj4OokIrmMCkti6GthsM7LoXrZap2qA86JJkQPOgvbWMcocJBe
nu/2Nur10vpvPA1WhG53KvxCTysfxp4g8lm2Sayf0uQegOhM6snpFFXOjMrntqjVeRTSueZxjcx6
/xRvPcpfg1QKk0w4+M/L5ElPzoDCxEhtXneFefMHFKtMhnjuPiyRu0pslqk2HXEB317X+TdRgz8i
cvv2eCGDgMkRYcsOwSI9kjAaHST3UrZvOYxkzXRPfMaUE2BG4TlDHhEGjzXHzTdEdOv9ths189zh
TPl0nFcv+YO3S/VGSEUKx6apEM69/sb8+dCDB7lL6eFFyiQrkLeoiMrxmOUcn7KF9U8aMNetQq4W
b4/30zh0873DIXec+yt4wfktQF0dARI71Qh64wsvNNe40ZwBMFXeB7F8fjGX5Zv33cNp0gtKI1rA
vxsob5uFOwt9cJzdWXgVAyKWNbEwguMD9STJBBMsoqFhgTvpzNhB4S23a4aClImKroi5XxzZ+m1v
nffYOOdny1k+29AddzBz9wCuvOL5kCk16UZ5egv5GtCfcObTinqJ+JOsHSngRvS63/W0p/Rh/E5u
4IvtNJ6wq6TFq9qHAYuRgMaE6xamrXclTOffwOl6WBUHSiLdeNAFAhBoUHghxP0JEdwwXSNLfwG6
1pacwzCQnuVywJZtvJl/KtrvCwwcKWEntl32vWuc0jaUT9Pit4O3Hknu6Oa90Xr95FeYyC4HbASd
Ja2lEG+0vF0oPV6ofvjWhd370GFYEy2hOqxrO3tc6z/VCDAhAnNmBSoC3MJP2sr2z4dJrsQzfGCz
14Whz4L7yRW6nnnqpS5nfVKHOx1yN+tdOUhpttS6ttTxDdYexzBdGX/Cezyw6eWubTvdHq9nH0E7
Nad4oCW2TlXZQDEjW9KLCQJOfYJ8YN6ed+hblx4N7huounNvTrNsVn6AcUMu/QEYGVywh3z9iQxI
DKTi2soQSiIK5nAgi01rAPfWs10vd3Iq1YkBkkFguFEMak2jo5DAcfHQI7M43RdEH3FZIfr6bncs
3fB3YDtWHpsrvrGUsCQ0RB+YUDgESv3wsMQZcZeSKiSBeOS0gz37Ry7vG+WWON4zOdqAH3deApXq
gyYH8IjyofXLhkCtyF+gVxHFW7YWLyAMMi7Zx/xahHf/cwp0QSGbnyXKloo95k80i2LcAnJKgCU/
NmeHJrGihcmdp6SkNbR8SCD4mN3Swr2PGGACKGOuSf1kVV2+C+fxT7jjg63jkGM5x4d38uWdsQJ5
JDxp8wHc0+psSNLFEUtolmMAUWFfomcOE1n/2tv2/Ndv4iYgvym4PIjhcQGRwvX9YZG/+frGEdzn
Q8RfW6HgXBUZXO19cuKPjLta0DzaQ8VibAjyN/4a9UsfnY3cRi7FAO9gIHSSktC39N0hN7wPbJ7V
SWMlC7AACi328LRMWMXMK/kzNOM287zVmP+aHbSe0Zc4UMhV9zcJ3z4sW/cq856slpvoPR8XrRf7
X+AwtjxZecuF6zkdrhOtTd7oB3uBVfVpzs5TbR45R/2Gz0r1ypcwhTpiYllhgVslGf5O8owpCBVX
A738DpPwOK90dPrHRWSdgq54uZsUgQuYCAGOA6iU7zT66h5uwAE85xX+94nm3nDLIRyrIRU5OUPq
v6PBkdFRQFaS0SkACbkAKcnLa6OY8rzqYQKKH9Qrr7IuKRHex7SFUyB+nWdYY17vOBnbJZ65c3s0
6wOe4WlcKlzcYUZ9vcD9ND0al0CtweOsG3/sgGIMSG6ZnS9ILZgSWz3NiNYirravsl8OrgtqehQ4
+mtb/iabdBV/hldRSleu7Mn5exDwpu9ZtRHrT+93kr4mA36VXu6lgFjUuR+lMrkGfS/YTgkTH93F
KNJdDz1oj3/iQkoqLobs6fcS5IenN5LUjZjWLGP3jDH4K7XsEDugM7tj3nd3RTd9gk4pYOOajfa+
DqCi22BDt7xAz909dUwIts2MkUHDoHd6hnuFCtGadjlHjP1yXiAYpmbjC+EOHc9VJOF/4JV6hZzr
4PQbozkrsdKO7l2bpb1t7V8YuCh6EeWEiIS0+fhPdX0zwV6YblVD6ZOrmv6cmJt0gpVYIVlaaaHL
LzYT8IvSFCtQOaVGs7uYz7fAa3iq1FICygxyNkebiyf70aLd6FoQ4D/DOOzmmMAOH6zcnSo8hmtJ
+hAefzzJPtv9JUETMz8YExOR0oHcGVz1yxvNkUaX40jgb+kQ24Dc2fhOTkwyS9a9hMWOoyxWsJ/q
HYeHthw4vwJVhfW0L0XraiMyin0vKQAsByL0im033NghjEjsgMrBQnACEnlZXGM6xIC4M569btLO
U5iezwTUnetachnuCj7TGGGd5gwkcBSQtes4m8A72wGhd1ebCVtpx3SYh9mMSUloUYdDSh9qRv1F
PmB0nqZLHDRlrcmo6eZJrGLpqtGkJEC5IUskAwMzTlT7NqwnM72haJ0Bsqy/p5KSglBtWjySKNPk
niWx89SnZSFk3defoeHKE5z83xGi+0YVq5PAGH6KGukDTjf8w79ED/hWxlhQueog9fFNgaAPiifB
NuIA2ahyPtRpBa+feXKXAlZeC/Ldjpy01mbZqXqySBRoY8SIVfDsO3OqcP9xWMb2XQ+5RM7LVjND
yJ5gQ3dYwbAWsf19X9DWeAA2KRbtqdmBSLffOIkikKW7UuLgBPdKJfF5GTHBKlLqzn6N2fBc1Hfe
9UfIR+WpCfonxItFNqM+OmPae8sJFu68dvfCXMKj1saNEGiGfDDZu8Wn9ZJVuvIzpXONKdE8pA+c
6EkUF8ExE0UVZ5IXNYkl251uJ/wSV5GYPmAz0XGip3VkMRTT+sHNSdI2H/lZ4cC2qZRq1Eqp1sgN
YRRwxbu6F9SLM9v49R9zF3FoFFMhL1I1G2XZZZmJPnJtHE+Oc2NVKFxR/zqr4c1VHnKxuKCy9ACN
XZ359PGKH1ewT9jJpfHhejutzaL4HLpgSsj15RsxL8CsYvGvsVcJyxCMscVwZs9CbadbsbwzxjPL
rN874EnN5L/1Gyp5RvCSf2pxS/TYfy//ub2VcWL6ufOcBf5hbrLVfHtKwzHucD1ZMNj0BkeNt9ji
L/BWmlTETKXNBvIomoIo8A9B/veEfLYEhlDz3Gd3/LhYOti+Wnye9GF7iWDfh9sKZorFASBa5blS
F09/Zwf50x+ofz6udLUF04ilGhv+464Igsb3ENf9KynsDWkXjvn2MO5SP5LetwzI4SRb25YI+k8P
RC2ongueAOC25R++mKB3OJbW7BCFi15jUB9jLahGmo/kZ0qtkRZXEzQfOSSPF668AueH4wNPoUZ2
/1CQBCmUpqAIoYnJuv0QXajgzfnIMk1r4zqLhmMOIhcI5U3PFkQfVXng4gff4yOI0sd1ksreDxQf
zI6BgkqP6xR475KRDaCJgUxiGpm07joEYWse0HV1YoQnHgEiorsUhqrskoC47HydXGD3OeREtzsi
uX0xe2eb93iiC2NxGpMqTbrnqrKcgVm+xFlqtODhBzfNtQ4J1yyYkF2gwxVt2CSXscEgIEthRB+1
9VhW/oNtk/mmZp0/30e4veXejNT7JJJXpEgDuhA9iF2evU0IxIMsQd3U02p0viiZux629teLTnHK
XLkwhbDlRhFbPHB6zjfytDqnwZLsusIdrmmMwOkgWq4FzDCN72Wduj6Hd/EANISN/DUFa4724QRz
0TcAmgYjomMBWk2fk4dq9oVZxq6qRPMV7g+aLYhtLPRCIfjVThCxjzBY8fzcCWikUzYk9KDziu8q
ALJDjJxFjxUzUR69BdNpDYelKPUzLT5UjXIH5mUNpVOQ/dbGJY2GS+P0gybTcn7gkAgP8+9afA/e
Us+7TcZXRrnTFOGQPltevjltQIghzyzyPpV1SHpUALwGqDEY9iHz4tHKU/a/lqCWmXCmrE9kTagX
pWoBsC5/8RBVxKcn3/nahdOYciOz5rBHqa/WKqyEd7sgAxdKJLlLIBBkJ0kxP+I06W8Q1xAH9HAE
LagyoRZH/1dZRLWe4PMjC14xScBRSjnK0UuYPSBu3zE7h2vYEN9i5PI/6gbEUyaPlNN+F+5e+6N/
TkYcdaypqKugPwZ6bofSpAsXhe9bdwp5JLHbC3j7pGjK1awH9OQmeL3wex1Bxf8tKbAbt3fqK1jA
JeAy36AMC3VRlBPLTKUwzmdr4T2BiyRxUqKclxlJbInT3xskbAtHEHT3NDzVGlhmHErLr4eRSh3c
+tr6aWSnaxoA7G07FBslgkRZ4nxDpgxxfSZc/n79WPMGwOkGHRzSZGhS0Mz6dOObV/Ryj4gVwR54
KBaEkahtwNiabJC3FK7MwY3jJai0B/Pw5xv8j76/RJd+DVko49BJrvo3wuizDzfspkP+PWvcZ7zA
3yV1Jm7A8dqFo89urQZsg5vhP6KiwhYvZnemiDefIx/wezllNN8QTbSE2bc80ogZAsYoWUZLG1/Y
TArtE/gZkfxbHFxWdWNbdCQegRBLszmHtgESxIahw6K92Bf50BbxF5yJ3DfbUXTdwXjafv/E4Ype
X2oT1guUin2bnqv5lu7noA/F4pqklLvajAZ8TzATzSQ9Ss08Tq1Lt94mSntV+C0InCdAkwkZuF1a
SkTPFkC3z5kAh36Q5xKRiIoG2dIQFjFZw81eYgM2GgKCdJpztbdeaGSlRZ6k3EuvL1Y1VjTmmz7s
teZCQXMPGzT8ELyCTcwCoz7qwO0zKbL2ddl1j+VdGEkwrp/lso2Py2hu0Xp4J92G6WnOYABCiGQK
zctUxvkBGaP3JteFKz1MD7nttVuKbtGTfWdg3W1Fv42P/YyusX6VYmKMlxtnuywb95W9NqgoewY+
1DNKZ7iJOb93xdIveTfk4eDjuOb9J+o87dAosiy6P+KqcLHGr6TwkXlk2u5lBIQER/6yrMyHVngn
KqwdLCBxg2/8Zi3b3OE2EEouWyk9l713oK5LVEGULZRot1VKsEu1C4H6oGKNRV37LzD9fartxt5+
s0Opkeomy3coGT/YgkeG8JrsdHwF4yNIBVQmr99RVIXpXC6SmN95p5slh8OHxIwCUp2dtUiORedF
McEh6aeQIBuMs7NgwCKHBUAgOQQ5BABOXAahSn+cmLArGrnwOLt3g51bvL9Y1btxyJzCiLOTJtyq
BVFrEUhir+k2nz3Q/ZFBXdSh3FioQf4rsRxDbrZbP4CnTcRcj66iFlxqxU9ko/VTj8GIoc+DWPbE
as5HpcIlE7cTHIbs6sPbqIRQ8Qnpf3zbXBU3RkMXUBkzjWxTtsi860Q3clyLldZkRr6s/7QhbfTw
UX3ERTdXN6DsaVtu0FCTVKGSOK/nXx38n9mxt+S8EdD1i3fiinEBO7bZDrIPk6jpT4LpMF/KK4Pa
LFLta2Bj8Fsr3HYFF8/3SdXtwHUzcYJEOPmO/h/laK5lmqsNihyULDx7afg4072topPaaVlWef4w
/rlNaqgPI+2TH/Py7bBK6+/APwtl4fXEVai2bOIcZlkxFS4/9ZhAeV6ddckSkbab2nmVt07dzXtv
zy2tek1N+JDiIfHwgeCGAYcdgAwMsMZBdfje9xeStsWqEpHKdhSaKuXZS+1dd+SHpk/1I4PHuGNW
9tx64xljSNoJMf6foz27J5iUo0KnPfCsIsvz+rurc1akTZb0Zaf30cPnYipWR6y12nVgo/0aInCi
pFsOrWy/vzXFGc+16LFU+2Yeq4EPYVcb5LKursTCC9Sup3mqPgC6I2piHkYkw8v3KSlQiCafevuh
EMVMZlqhPoPqt0bc18uAO5D3amJLki+sB2SFAMZ9Rp8LK8JtNNl98QFErlJzLcJ59la25ExkT9Vp
EQRET9bZIRjZf5kCEHpRP5GLhGeXGBm1d+Zbc3sgf6rpxEFbW+KmpuIxFwPvY0NaVqov7qDO9r/r
sC6RLOefqiA0MLIu2aLRvh/ga3XT96F6C4O+DzCYKmeZzAf74mTLZagGTYhvHskGoa+8KUq70f3o
YnmSldbyEJ52TToiiQJPO7qtkxOuXqv0orqOuzX5lyBGujWdZkRXVcukgjOysIbujfAaWCG7J52y
HJOGmAkUjlWlXXPDWBirqHbZJieCQe+UhVsloIr58V90XAmpwN8aEbvMlJb8tVFYjJh8M5OXtkbN
ieRr8E4Jp3iN9Ie71OCvQ00ktnSLJx0bCFNoebatNlgthPjO+nfaMl0m3FoZbh0CB/sthFD/+/rq
I+9ZMk26+ISKlflAJIAf7AqK6plPBp6HdjQXh2+v0rlSMHjMZe6UdQlAx5TVyar430GayXSNAlSh
DlbgwJEM/wa/5WiHDBopZznese9QV8ZNRObInzHEd8ySp7nIrol+6sGyEqb1zQ2koL3w6VU8HACV
hEOnCNNQfZurWzS7mZvjyfGInITkz+O9Vcz1pLi7ygZP8JoEGl32JtuQQ9qPosoDez1gzdhgAktF
FQ7wOldPHmd/vR5LPC82XQhIoJHOgfc1msMyr4YG48MMDwztCPe1sOfaHqjY/0iqjhv34dDjuC8G
wB2e+UAE8qIXvIjfRNfT829Ofgm1xlgns6G6CbwX0uxsAJ8JwMv2+muy6b1rl9It39lfCA5zjwqC
90zHI7v0rlaAPfo7AdT3CxgWB2Am8us0VlicAx8f9JeBxWiT6iFPJjB4DHM4KBA8xM18bnhe2sva
2osAlYs9xfkpdVCJKfGcAxwDvD/mq7O0LXrN+ToxiimmkIfEWtNoxNXvVUVvRwWEBj2+D8+PsbF6
gRAKS3aXqJrSEI+5TpzahjIpfnK7cP0SR48e2pqVQUY8oEwVmnfgCG/c70p4WlQQvWnCrygr2EAg
QuzQ6j8kmtOd5pfvwkvVEwiocCsUsv7e9nq9ZT1kpXSIxAZTjunnudgHx7XLiOC7nQFhroQABlS4
sUymswyNoAN+7Qe5+v5DUEGzqvAAz4GZEE1MezhosPU9gv+2dx/rHwy79AIlKn+u9Csvo3B/06vS
LFpCj2WAdWO2dGeTF2e/QjrBBhlWAoDtes5L25U6mK1rqdTRk5k+vbDT3aUZkXJWxHUbqlR8k5Sq
P+K0CQvfxQoNcUi5D2IpvwJsGMvP5GMk85+7TyysnFdVWOioYtl0vlL0qBQwJlPGX+eSF+JbCthL
ZKcT15RkTMZY4iO+3/QqPaLQuZRnVAaOL4s4+Rv6aM+WX7qU6D51WzEBuw8fZcU5wwK1JH9U6TRc
5rJAiiVNyxr/9PXvgcQI9cy3Cg8PNDiAIjGgGXl466AsmSckNaEw6HAu7oQh+B7UMQ/G8Cq3R3Kg
rALT6VUJRjS9L39kEcEGasTQ3qBglgtTX5EEt6Cm7spn4o/hD4NduCqcXYzCMT1+y+EOGJHlAZKq
fRQAJBRS1S3fDw0Z0snzaKTi/wJibprGTxIimbhX9RciJHdIjfm5qwfQvv+PYdPuqxZylwdUzZeS
X3C0MkJzqD18g7OrVX+Yl3Ccin8b/Eq3KI0USNC1lNCfeZUrkzli3BUFbmwBfD5LDDDiVi6GmsRg
okRDIEUo4im1u7yy5KgFc2ueZ9Ln+0GgQNBjvo/McrnRUVPj0/ZAoGUqMO4CSksGc7U67XGmsE76
gcgJk40smxT6KjGBzjlSt/9fs/mb0++QkyYv8CPpSfSR0Ns0A+jKOXN2d90hsC7DYFb13uV3mIjd
ePiREx5Sp/kfGjb4mZWZt4dY34wywiRvrOz6a3cDcHWMSRZzY0YqmQkpND7j6xBzdvCsEg7ffGZg
ejVFUAxxiwOD9EjMgajsIPg7A7EQGltOtGtHZ+5DWSIwsVB8bZfriI8e8aCaUPG89SSR2xo5NCfU
lsV7dNXUmr0qj++baeYWSW8jt//mELikS0T0ZaQjxJa1c3AKzouCPTVZsidAK/BofFqAbagKulOx
H9gQqq41LIGcuuGhcsrdA0l+8FdpnxtceAv7/I/iZrOJKUpZ8yJG1yPM5qzMDO3rrbLyxDK6HCgI
y0ExG//JM/oN/y7Js7d2pGkHZ5bFCe4pFz4GfMe1Eq2GEUAeV4Oa+ykeVc1OcPVK8ChWqdMSSPnE
iyZj3NweC+ikC0sfzt7FxxbRjhLhmq6T3dynKpYVvTXI2WhQQl+VapiFDeHiUomNDaPO78LfxHDz
HFihS2WVS8HikHGqcCrR4yyfQALwyApZePl+F+Y7oQEQDvzLja7RGTsMz0mh8zrW6tMz3XMtAYDq
kI/wH4gY4ogqIMORXCYHGvgfYnKsmGP5j2mUxbfP6m0d1VPEswbtXgDFVZRzdoLbpDvBEwtKRgIv
bDd+h48RrIAJYqjD1Qi+3fMm3y7fKAF/hoXongkaxDb0Mw63lXS4P11oP2WV6Dr55PZbL6MyXnuu
kqk3yRKE5ua28eH8REqbf3e6oZl0Q3YbdC5Lcz5Z6Sut3WxF4FbA4/6UXBWxeoasA8jk3Q+s5dZ5
7VUsvhjLlKHGkyc07Z+9G0+4JUIVqVGyN83hDfv5+biqBdWLv8FeUJqXUdwoMq9uZSEkiVsL2MXy
AaitIshaZj+abFp70X31p1R0KpEGh38WoKK1eFcfbV1qPKpwgNVC2BeZM9pv2FbuPpsc+SuxsFAT
omDc/UIwoLQq0NxHCRhjameRFLr1hNfcYg0gHciykWCY5MgmYZHe0ZZt+4+hdZQxS6DgJPKIyBoC
HkL8OqhZtAj8YpkgWBYbEr1so7P1U4RZ3ajsl1RCyt1jgoDdDTsOcAbQRKBYboXi4beLZQJ0BqRK
PwIW+oQPlwxP+Kb0yo+HXXiTOHGSrUXLNfONnzVBSsRVLxY0CWBFLcldvYEQZFP67ag/BZLllitJ
xJSiu+QwOzt0nFtuUJDunVAFQV+bUu8/E7N58koKGU5nrJB05l8MCtF+j2p675+V7WEqgJvPialZ
PZZZWOQBEHyyE3tiKBghu5onXPW0ps+ukbyz0Bw0cOoBYZ6FDzko39s5SB6+BqJGl3ajk/ub6L/r
2+JXT3pe0sUf6N1Wy9di12BF3X4Gq4L6j5qVE9DICvo0lX03ikPz5YiRVhScWvQlTrSr7xEIsioY
zGNh/APQqvGjXfEkn8s9EM231BBr87NPlRhpCP8YjrCmhNANZxcTK7rbszZbl2xIhL2/nmkNh2Ht
lk17a5SW9kFUOlqkyzaVqikZnVNWIKEb/U+k7rnDnQHC05rmp+kuKy8GsKZOcYG1/gbnIMyz773U
jGqHljijLSBuwCADQxtoP93qd2bxrqGzBWe9pPzX+8nfowG/LNjyqbOIaNlx31dYaye/UujPKJvE
qvAkTefOsVsowVHD8ucP3ViE7ZVuwMHuyCoJ3F6EUWClW2ehhegBsiBOStgh6h1+JgwAiJ3z2LR5
X2og1KnLhH8YsZqj0aH6purVgInGiZlwfUARJQEy/TkHulDgt48c192lud/y4pTc9bcLvbCArKaJ
a9fnBr699ZykZXS75vI6aIFcfWElhn5LzlzKl/1a3n62KT1lIOdBZsUwuXxmVRLKOeDVblmoEhk6
sCgRTViAYPk9c3tqh61q3ZCZ0zmfYF6slbOPg7MARfvj+9EBC4ZidcitrhkYLWfROjdpAwmP4cSS
RLOUptWuwcWLRzEiK6VXNNmKkbHkx6nKq8/e1WQ+In4XAi6yNkSxNTHts0erxjMNOY9bO98TtBFP
aGwvaZEFY2lOlfwwhPOrhWX3mx1t5Ix7TVGTWKZ70k0dJf6SvrHyll+DM/Zwfo77NoejjadVTVC/
xiZk1iby7KMGxganWg2at2AoIm3G+SmiFvMyc8ehrStr3IgjL5wN6IHDTSciqWK5gEOVhzEO44V+
froE1/rEM5w48RPM31M7xnh4V5RHmjmvGzyhxn/ezwCkJhhBRVVo69Kb8VlhBTXUteJrlYoZesIB
3VrhmxMvFj/DG1yhqCtHWvORufCjsB1oY1oXeRl0+TDiEUSJ3Jddf9yx7igxB5DZnS8iwDGkknmm
fs2cB4EZZk6S3Xxe6foTN+2SaUvknPPv1ZKiC72Mvcl1gRbNhHits2EoEC7xYbGSUvWPZUxlOpn8
LQzgOLLx9ncmmRn94Ys6uMkMd6OaqQR+bfyp3apuM5jCDL04jyN87+B8lqTslDPKIUcgNguaQx5p
jWDe2IEyEbpGRw6cT0F6I5spxd5K+EWRHBanzEAXI2K8cVcK2ETXyGIS/SzJY+hlqhkq9V9Vqg27
3mm94yhshFTAD4XYqN+nca2Ht6gexb2k2uHXwHwvvv3IncrTS3gOSFIAdMErdwjpUDWr5MBnvf6i
qrOcfxLfCOQMF3bPtRYZsdPrBxBOje4Gnu/riAUri0hYW/clSWpaVujzpSntyQf4MniUVnmGoZNV
nd4zHcyqY9rKtSUIt7SngkLOKABGuyPatntuKPflOPhpYBGduG9QV+6UOVQwe9BLenSrb7yb0EbT
5f0ereeuZQYLeR+QPySDeILaRG2PktOo5At/BvOF8d+94iYYlweQNNLK6PiFnM7qJm4v0yFLKPF0
EzVT9XRQOvyIRiP+KAQkfaCcsZokab/U9bvbgzbuFeedypAFaoUeZ1nBt9wK3dSwrWsgA4aHgHRy
okvN9uCfle1ERbUO2U0YA0GYYObButJPSNPgfAoAYxjKVHgQte9R9rbyOvJ5HrtNtSwEY6Wo6X3V
LCkPccKJyq2U2wKvub8uuicbH3Xlqq3W/Msu42NjYbfUSyfw3CWJzbHtx0e8c94rY5Fu5609Go7D
jssWAD0Pbu4j8EWbK72XRKoTiQhMFmor9bn7E9uymzDsnPBDpYkS9Ul5eYYNE1d0ogIV7kGuFdoa
RHJDFeGk4Ygyh3HO9gQYPIOcDh0HORwwUZUJojo2uw1PYU66nCtMohoLv4QGT0lXe5x0dn/iqsQh
LVtRh2QTO9bXCOdcEQvoho45G9wfmTNr1IPkutPSegfmT5PSbzgEBRN9u8RNuHf5+/sSHA4GMZVk
OeXP/5aeC8FD0HXDZMayA0lnrgxuv6i28xXwpKPIfDvJxrbA6RVBijyhzY37lP5QJfnS2ZVP8RbB
VCyY6EcUhbB5y3KL6ouHPPJEDACmEcnE4WSOjTY2ArafPQCOpxIzQ+KLh6hwy0QQUri5cckVzKZn
/eUOD25I8eniqp02pAMlgeVivOwvVEb2pCdFyZPI67YbkT+RcfCiHFZUS4zwoM+UrSi31NoWloqE
rEI/owA2XhqLQJXUS73WB12evB4Dn/GNfa++NKvk0s/ADeGfjvhO2kQZ32Q1EtBECVjXcnJSWcvD
qDlsxjPUsUII7CGtjrMT6EP+F3En0HhcgmIXqzw6VQagb2AzCZ8P9BCNSjc6Fa2QQcaYaTH47YhK
++CRxP1xich4yc559/CZI9hXjEpbVK5dw6rZGhccal9H2sAFocwHgSYPF5+SY5oTdElwdZKrGEDU
itavn+4bCf0cRQzgJkXpuGgLlZ80tC53jiXKHHHQazpWjCM3UZeOpyrU4J826naWfDl9aTCM4qyp
YOKcLOmJLyhKBWQXH0pVM2I258YMafJWx8u4h9Wr6SoLgMCMaunoM0jw5/5Qoed8Ls2EhAZTodHh
X21J4WRSPxoOHa4kL3+YjjDNroQjp7RyO2L4FKl/UMYSKHGoS1rR/2JCFCZPoTvWVl4HIc3AR6rK
66H+EzrCt5Ofk1Jfa2/HE7Rj/dpkPHbYKCO3Vt9xVNHEUM8x+rccy8giujQn/5IofAIHY96+WE82
TTA2oVKVjxTYuOxFfCOXcuFuQSA1nEiKiVyFg8Iv3B7Nl1B/cZPHGMhJ7PIIfNwNveOkBw0yO3cb
seUUecFngJUHz468mPOz3cX7JHDUh7drtERp3QuNqiVCCsa008ta4Yp9f+nKU6SrIQQpD+wdK7HH
zLqOy269Cxlmoo355/einZyGyHs3JVTimFG2bHHCs41/iMyHyBhMz3TFT/iIdycgzTHGVKNc2F2p
oYT6tbLmRMwC5PXtYLQd/pRwQxvI2dyqFNTHelYYNA6CEbLr2wDqoIKmI7DQiaChZOSSTsMxPW2Y
BBy62NsYBjJcPtcb0sma8NwQ/R7pLVdSXA3oUr8eASrAKlMldLFsL8hYIyle0/xvgRbStRQnrZ/D
CIrIr4O2oTIteI5CjmPfEA2TehleA6GpGAbLJZpk6wNuu3ghhSSLlwI/E4Z+xSVufCeRMvQAcxX4
dxNHSabiCcwgMKnDJU7Iqq1Vt1oPS80pni+zRer7VCWus+qw1dhwas7RpkLLFPaG+41Rar9PKjT5
Emk9zpFO2FtPMgmwRhIANlRuhRcCi5jvdyGDDO2zessYMFYPs8zIaKr35j0mHphiQodmPkskrFXh
6jHrjgkBKbFhu+n/C7EGqGO7WFtfgBvpF5eiGw8138M3iInXy9H1gNXhLjZYEUYa0C+dTOe+Zb+p
kEEBNHxmJZsRaUSRDHIIgFPpodWnSpRClG7sRRmsS0/FJZcsZ5DzfVbWByCTn+ZETkeZ/ZZCjskK
79B5nITmhOgBp2O24ZWMzTZBbqA2inyhH/rfE0xPMyrnVqo3Hsrvao/rCTggYxONZ0ZehvblFG40
SwhpPS0BP6GdX+e6vS84uLEUU1TeOuSXwcOjCrL5P5jom7UVUlt/X2O7ehk2RkjGmbE/HQZzRuao
ttuoSZLyz5LzxbOIfNzQ8FmUJXR26aa1XZ1yBU0CCq6d6ATwdWubHfpYcj/7IU5o0aSK3srHEuoN
R2WPnMXM/jBoo58VextpAvB5i3NBhTWF7lvOdTAIbCClb+EUa9B5faLAzTaFa5sYujiNbzYoAD3K
qvKHLwOll4w6eCKgRsUodxM/pxdJi6sXiG40Ctztn8v5oi12CM37L+BFSpNcp4ZHyvTDe17g1C+F
bjhuHbAbO4mPFkZERVoUxKAs+awIH25WY7AjDbUPrrvqwYZt6lCnXPwp+xUFxHmFb17JgTUFSRmN
He2Te4gaGhyxIHEjbvwDiM6AalQMc9FCbRtGu22SXVQjZI7l28t1NXjAQpDiI5cVhUTH4q0P7+uW
tOD1FGcJ63Ebu+ZGiI5KWyOBQlX1EqWmIY2LDyJzD4QgVWbLkhHGJdzJ10tUDu79NApcv6BzmVv8
V5SKorBlc1yWzAkp8RK7Tz76ztDsB/WOdwxXO7cWEBwyyz5iR/A5KynRicj5ZZdT+wXWVdNe+U1r
vBbgM4EjpzGFM/sgLOLMiHzepqWR0Ksi4titVAJs3PWkw/ouhq+A1l1xFB3fA21zL4r4EE5CN2ye
ZpFsR6ucBFj0TS50n5oI/KPOz/3b7MYtHO/G2Gpw6nfxakqHQ1djoCWM80JSe3bQ0CTKj50hB5xA
OfgC3T++VQc8Ps+iAK/POMVhc4qFN1UhU9BTvKHyRbhSSW0++pS+F4rQJWCv2DvThhcF+Uty1Hq1
tfTvx218xnJ6rSCcCZ3RLGBlI5ur766TDvWRr901FbLNnmJUoRdyMvw96X8JWlTyWprBACoci/sE
4XkTv7RdiE898wSpDy51L/KlLRTJa/w7lMk2IqdH1h1eRmWZDQN/9WLI3vodRsJiFg+PFgLnNoFF
y6JfYI+JKB3bOlSqH3WYVIE0ScuDHk3VafOzlu4EwFB/8bD0ko5VSchg8u8gkij1RsTZinONyzcR
iQfYl/Yo9eNwtVUnSbf1Gy6OW0i3lusnpKQQkQvhp5QqwLxzWOsUlkiYW5K3//ZY7aN91GXMOApc
gGpC1mQb5mmXege92kaCUvGdjw0goQmn8g5WQT0w8xBsYOxNKKsuyrjmA0nH728qiwBGaG8CQhoj
JBdMLEBCNfwbUv+K35mJK2Gi/HU+MwNSuuXU2UUTcNY/r/QDxBrm2d1rWDenUrrLm71cFOeF4IhB
ZqVPgob3tuciL4mZNk18ZU/OsEK3yvTYi7SCno70vANYKm2C6GLjDYwc8aR0Fpc8ADSGang3zMhn
DlyFlo2cSbP3FNbjvAKTYu8fC30O9VWvUW4mB5vc5wXszTwaOe+ulaMaeQ3pZha8oAVY2eTE1KoQ
PpJY/Vwe0XQTk/0Mo1nfgOk1jmEdkxZ1rRA8K9N1vNRSKwLq0FusL7fQdmqXDaxuEY1APR6EFyZu
Ais+Wrc1oN7RJg8TkBdf5UnWJJS5dAhwmSu4ZuiUBtsCavEpoUo8r3caEkVF++wFWgzJQsFtGdYE
DIiKK179Op6wo71fV8osPm0kHn8p9gVVKAY67r+HZmLZtmFNYUCqRs9aCrhq5PhFtk/zePylDoPo
MEdt68s7OFLHuUpiBYnr8MlnTCDmBw432JWelEskRjqvm30ou5TpWCFsqH5Duiqblh4IPiHIyGRa
K78WNPTXbpG/r3G8kfeZPDax/HNuWgxmb+tCY03oYdwebbSzpKDsNgPlF/RWEuup9BSgvWXbXXQp
2V1oefya6aOjBGOXa/9n1WAgSK1XX7x0ziw5j/631qzY+O2WEDpL08/CKWKLDco5OaV/YaEGXRCi
++f3PDH7Pzl0zRtBcJuKBYXvtYTVAXEuQ0FCnzDZWcN/begT81oxpj0WQNM0z0Aw5uJy32wxGKsI
TCQJtUjybRjPXZKeuBZlNYBB7TKnGmosixhdZ1AEzItAaLtRssucFNxYDLTeAZmU9UtgBfMfK2rL
XjtaspC0fLKGkhDf6OpF99LHsXOGTswpSNI/jG1FaVtXFz69uHQqBRNoQr3nMflzANAfooS7nb5k
2Xh0JDyPovv5BUvDJMtZRTi7suJD06hmuLMk74pim6fYaEuS12dAbyTOPv2NNUa+dP/GCyTNtDpY
ZuIgLsp41ArOJ+fIav5w5e55av12wUcf3bcYbC6oCHd4DP66cErOImY9PebvHN9tG4weLlNIUZ0Q
OA2QX4bjRHPer8eAiGSbJu3kb6rr+TrrQN58aIvWK/fgh9KWy970dQxIbJJAoRna4+3W0GGiMIE6
wkHpntbrpUSFbRv5zPdfcgm+ep6xfsWybHeX3rDJJ3tf8BFau27NNqtWHhETKyes2tohv4dvKcHg
4mY2yrKq1somvYdGIoQqZeCxAd+QmTKJst9TdHDszKulGxpvT9jMn18yrCW5pddm8fhrxXxLrIuA
RkUXUPAaETh41Fg/9E7JkRGDiW0s+ILClXZ7aox3ssY5vW5RnsZbjvr1UevF6DYgg7DNor4Tny5a
9KpJ8kvgl+ZfXacz2Zls63S3Ct3mPEP/gsorG8iGYsJ4cymnliVY9n5mDtb604HtMRA7btIxnAzJ
52xYgyTuMJsMg+OnRH3aWWS+VnMN9F5EnUTu+whx11DwU0Vc5HUI5OqQTQ4+NgQts5RnvO+tVrf9
IFYz+cfkeJ/hm5kVYIrSQ+dW/xdbpXiliD+0HU9sqj+5y7fqC8A+JzTlw7xFUo2hwzQMw6mEgJv4
ZTOLckuTOULOVeNtJLL2t9iqnhBytfjr2X3CsG8yxqDJStoQLGj3eT+pYnnf9nGWhYchXvg9upUW
MMWe38hHqY0mcUEfiIRaA59WOGm8IlQ5AoWl+5CjmukysiUfcpj9pPEAtgeYBBj3k5GvmBe+rKPc
52eEeHl12aOL2QmTs8ndvbEp2xJ/xDwZIU1ydyJjdv04bKldDfk0X3qdLeC8xdLzaDhzyUh40+ii
KuBeZ1Go1mYOu6RU3kFKDOPuBhY/9Nf00Epnzxn/WcK23YM74FoI0Ko9dwBKkxAct+yeHw6gjPQu
g/epKAfVJzjeZMjui5FoL7EnDplxUNtkqqykgjk8hF0YuF9bVT+EV+assQYJBWjCh3R6FYitN7X4
WXn3YsfQgWVtCzVQDOldpPkSVa5eQrdvLU9Y6occRp11u2n0T7ta3i6VkorrSkJdNMMzjjOE648a
mFVnNR3tpwWIcFjcwPteWivUIeDJ5VNNRkSWWgzAlBSGrNMiw9ktIHDk9yeob5qhPKw7TuO+Rrmm
KHqS2Wo6B1/vI2L9OhLJWac3r8zIjmVmA0qWJwZpallcE7MdIfr7PiBfWc4Jeq9Eot0dK/EOS27D
jJD6S+ASpZdMnI++9WHRFyehgXn5tzSTPn+oERgmdBjDAgc5nGTI7L9WxOHWUY51LulHAZmLRL3n
hX6VTp9RjVo5fH3ddZHUSdwRZ4SRJV1uK3nnyzMJE1EBNGcXDVNh+Wc5pA0zk6ISf4LVeC884OXW
eDYSKxxZmg6vcwQBgYLJrK82C2fpXd5yOMlglpVi20tMYoe+3pBpF+ExQxOMCAdy3ATLa5oHTcE4
/f02YHH2wRzgfnL1XaKJMgULVBYYX/y3vhtZbG6NNGCb852rIJ+dU9RbER40JvJ8b1tMG9FGJQ0G
YD8mhJjhEwsSsI8mbHdGzrOoUsxAjSae5pDnhGR1/1Soi6I1e1uth6ryHkMPtzuYqHvVk3ClBn0N
gDQEFHIMOrYoKQoW6OZnsyxpZaclT1E7N21XFKS1SG+4+e9iTBM8/AtP27ChUzU23xNgXZfQaNm8
DZaTj08i3MYm9cGsueJWpthWkzftTeVS4ixS+Lrf6B2iWVqh6YXwE37knttbsRbiY5wRHpcgHN5D
xx32w8Ki5Ui77ltEbVWrx+iHZPO4ixB7zQXN8fjNWkHRKUJQFdSR4fcM8VbXob16h0ga7BTT1ves
O21W1UDKYvOkZSVX76/j0oF3l1TQOCvfhVuf65QlZT1Fh/qcImB4CUGeYHe2tLcYr5zUhQB5y6F1
ouJCj0anri7qbSrpdOhwItW5wJI77pr3TWJRFHVFOnBFDDNuuIY4DFjyq3bIAOh35XH8WP7UwT0n
C54U+XvN/WaF565HPaMGd9gmuoaRy34I9eU4Zt0X01cK4mNIZjcAORzDxBHEyIZwWnNiBG2UZiXc
N6ObTUqLFZSXvse7qKDHpkjhciasAnhjqMFYfTS40D2UDettCB4ymprqmdsVJT8WVQe+C/6APxIP
PT5qMK/hd6BiR6iV3ym0WqpOEBuyEQt7DfAiCO6HeEWkFzVYcoVVziagrTeMk84rjR4Y9yYoyZu5
nB8WT7gQLJtlshE8B/hLJTh1PG/SmEcSUXHg8ToXkOLUIrryT1Dnu42rDtrB7jzpO3NNWqnDLw1x
LWbECYdRlE1Ba7uuhBfPSGam1OMrknp6gYJQ4hq7Nur9xcrOf1gRaw/8EuMWfZY+QfmaybZAeY+w
hibKhazpNBHSpWv+P518UnXDybS4KmhV69bLqNb1nYuvUqpVRTLZTzRCbjcmcaVkTgkAFVGmKIBJ
GV7Wjus/7AHICjrNfclgBUCNO25d2xaqCUBI28ksvFfsAHCHiysVAdHLB0NMfnROBPODu1A7xrud
YFhYbptvF4rzLBPXLoElm1iZh9zcGFtfdgSXjmhv8At1jwDm0N7ZXOb3dNUJwFY5D67NIwI2L8P3
rH/OHWEcB3sg6dFfueMrgU30vmNW7AhoM9kT92E5BboPnsSOgWpJAddEeJ4lZP3eFFnapJ3Or2oC
k8G7sWRoqn3MHsUbdYFDPkyHa4s1SzFRGDYJx9AifohNbqFhjkcfZGxaaxeKDH5RtDGIgBarn9tF
XBO28I7K81bDxAgmLU3WT95q2gL8oXQoDKzCJADKM33pg/xMM76Hlk7jZFFsh4G46jY/RGfIkPoB
9KyxmSsMjy6ewHU6g16YXyQsmTC/VPS1nsinNHzqQUU3zwwsKfIHUN/yY98ruvC/QZ1tzRPbjJKn
ZhrAo3Ju4zilY3kuuwzlTag4i0seAbs112w3pLMp2BDNNi1Mm/eqh7tb6p6Ps8yWIK/iAgks/HYs
avlo4mEMHy0RwDFD50ghQKpKDync8smPefPr77sJSDbEZ4JYLwBEIkZUui7zivIPwlcclNRv/7L8
bXs+jcOxBa00ICbZGMWvTBLBKwtePQoNempfqvsn6bYStZ80krTdU3+vnRh3+AFHMCxBk/pyhcjA
I5Hjj0Co/D/enWrwsS0PhspWB3LySoMbW0yiZ7gHJQkfJAHVpLaOz55JHh6JiA9suQWs38JztsL7
a95vAIZhmuCs2IH+njpac5IwBXKmUYMR9sOdCVIhcDQz98Tkcb/PZaLP53MCqrc8bwzqeYsXYOyU
YYAX8b5fC0ekCrpqovWjYPV5rxto/xms/iN8RemQvHG3AyhirH7JLQhYSvh94E4LamgOVDLCnmIv
5HsPqY8gzM/PB9cYl/Zw7DExUp2dDgEDLL+9hb6Ph9u2hEDavF9JO1DDJ10uMhF8qeR5n8ThUNSv
2XZNwdFteXweMXFPPcFTGdzpzO1v94TfX79PYB3LnO957Ak5J0weR+d/cxKRu+753FACkOTKzUhJ
ZrevB6AztxE5nt0epAt9m4DdxVAj8FD6Um9xPP3clAVKylvZZp6bvSWzzJZVcc3bjY8ZMYfb5P2+
b9Ie3gXf1qyeyMtl6WmYmP+6WJYqjQpnAfEjsdV1sjAEBjjp9Z5BeeNCVBBn72cEMOqKzmPl1nLE
D5kwArZtXgrH0USnEpUeGf+YIXqnzjqffPCXTJdA00chhmxr2wBGgsjse9+o6S1AQ3dxtG5lYd1N
5yOQanRJnLIHRUdBSYifgWURgnTdK3uY5w3H/d3NtC+Dske5Z/UHnIGOlxA/MAH87xvEGLh5WZ2U
IZt9daGw1hlT+JEmMD/xJpnHYtaFroo1doSnbUGQUFq+gmQXqc1SaQ4wAiFukeMlmbBDcJe7ZX+0
tdqcOWox0r0ALgnSWyEGCPC16O455IG0i+JxvddoEY4ju/GO6mJQKHkLhXxz22Hl1/QVP2rB5WUv
EOo6tFJA9SmQIoHFmOxBuPWLDEWYH8Livg9rj1e/mHiIB+NMop4zaGc9KXoIznowlNyedV3dVuyO
Z+51SjLwkx+bcjL5ltH238hTZX/kT8EhvD0A7a1ufVxNJJLF0fldQmDms5+o8qpGscpG6i50/Odk
/rMq5rpLVmWYF9sdUNYB1s+6V13L8LZvn7G1pRXJCkWt22Vx7d4Pc1AWQ0BEB6U8crV5nBn4IJqj
mKY9KWsvWI4116E3G9Be7aHOrbYy7A8sYR22FtduoTptuFBVmYLSD/q1jAPQ+9QiRCJa6/4ChCiD
62wyzagYuBTuHStMefHg31u7vuxjdwU0mjLqLB/t62NdGHyjfu7yb5+xkmEo5Jr2spxPWFWh2iRH
igfGBJKnHR7Xh/tV2NUPDz9VttboqDFMxnSHDoQycnwOA43nIrTKfuV535xLFa3HhB3W9u6IdgAt
fc1rqhNDmReiwRIGSd96MLd7a9f8BwKUen2FYi1d7qe3EzdSvYTfSbCmGZhPatDq1EZEoriekEXI
8g2kDZR0KSC7b43Tg95ZNUfuhRdv2QBo0xCsa6hxi7WX3eiVd3ZqoOExVzV1mJP4eYxmkZVVj0FP
36NCHR+qwizvfdIT7W5zmmXX8m44i/Y10ukLagLwwY8ErY4WE+GXv6Mi4jmMjlpZIq6V5RIX/7jx
OFFXr6AFB0K79DKOg7bvCdm2Ae/QUZhKwqALLUkAcWWwZOeBvNp64B/5UtYvUzMDUIJPLdLyxshB
rbMz6g+/NgXWP6bSH0wNiPYKa6vZf6HRwbsloLEX+GieBBSOd/pGYQxyIqtlj52I0OmLykBlM+jn
sCGFcoMHAa8h5fvVdeIW/lIEonlwMLJ6rNXRhX/E7PmqYO8J329m2LqPczy3IYqkm6oLG2lhGdAW
9H0eIdlNWNplfvFeF2VD4NKqswnUpsSJOCAQqbgYRdhWQ18wx9ecCCe+DpY68EBgJ7mQNiDgU/fg
YUOKheQEe6gCoG+TNSKC2kKTBtcyWSGw03zWh2tW4CSsqsmbuR5qBnWx/d6Hnm6rPFM1agbH4yjU
1ZNkapt7tFqEY43F0Y8C+R0+w1/TYpmQuZoI+HPIerx4m4ij/W3dBQJUZB/5SWchfol3htrDSxFR
DXDjCasTmuWFnBK5e2T7VP/d6mRfwTnxsMgAX65eB5M0b5ebBZtTXHc2kEz/5/1CpmpBs4D91tNj
IXThC6sytPBrQNNKEtBWrjkKWyPpGhpxHZZzmj/ECvdmiiV3/u8zgOKvs9ATpEh/XMNrfD5tWYSe
t8Or9v47/7jDZwwExYkFADYwSPXXyHeUDpJo7zoHy1sGYpD/JysUn8iJKnTzTUtb89QSEQ6ZqJbc
fJhO/F0RQN4+0Ol0m+dfpXqcHLd1MY81igDNHLFMdVA8clGPL62GF4W6RqzpyFTwshDa7R27diqh
SC5+H8VUgbAV55SSQ3U78mYbi2KqLlIdzVeqSJxf7KQbOJo1l6OcNQwwWoQ5BT0TJiydzfx2x29o
eI/PznKlZ0W+vKxscUoau8Fnhuh0oIREo6OPCRWN+jjUcRlXnC+9Ut2BkFpEKDdeohDekXDn85uL
p/OmIpRtZZyU8Fq5GyTxo9zw1DDesFOCXzVuxp4kRA9fEjjGJQLpi7QsOuiBMwk/owU2vm0tRXv3
4eV3JiQ4X7gH6hcQDMts7+5lnCwTGRbhjBN1uoHBVPZ8fH2UFP3Q+aXbwTo81ESKC2Gh/1AdhkpR
xKqSjUH/XJbRY4FZnww0j+gMSy2BwZvcUlfE/djKn+Wqg519gNMa+rdjDLR3tkeGKrbYtuMvjTqd
zW7SHatySAkvDpeTcHPH2JgeN/MFnECFoRXWbmHgqAoksmFrHAG+iGmkc0CybqXg5FbMlRjsHaI5
ZQo2tyZ7qdAE2uAQpDXrGiBm9UzERiO74iwaBo7OXUH/jwN1AT/VP6a1zU62v9ggla3T2NQxZJeA
SSFpaWQUk6uG95Ofjr2Yj7l0G7ph/JFByQC2sWTDVfRcs7stT3GASvl1G/rrPj3RE6C5aEGwtnR5
GM1DLVuDXLnEWELau6jdBHbpTgrvbyAykkS8cm9Yz94DMrSyH3q0qRT7aV1MWvgXZNCvYbpR/zXP
NAhBr+XWqEUvoXCICtyCrJ2cHaRz4jGdMb0NyAeH38M+BnXmJyOGLsaYwkUwE9jce0Hui5l5GO3C
aCf9OA1MbYPuU7DaZ4VHOr51N5Po3jZhX3OFv+5iJJlLvZ67KzdsAr6Jng3EbiYhDfA4xIzYmOlR
Py7kRkAtMhC+XAW3iTDGW6La5q9Mf/N9dk7rqvuLYlUv6L89xPS24bpJgNri1A/kqtIr56VyzlHS
SFtZj0dQIL1JaEoqKKHCPpbybz5WIsOCvrqKZ5TZOvc0ZyKd+m50agFU1VrXg3taHd+9zvsoWoAa
kGMXZVL6BQBiHJ4yhHgzM6OcIgVPV5owDok9GRJQ1mcsWng7wqyjNBzNbNKwwizPVp0VbOimY1Yg
4nFDl9CfDzWOtAFGPvq9TtVM8+EwZdDpP1NZhXtKDv81IIrSSPtMaCv766XhvfkCZoTFEUqQi3uz
IxJWOt7cKVTJTPCWGcDoqoWhRnARKBe9CO+JlLD2ZP0hfgcrLJpJse2Ebg+jqrt/ArbSJ93BpVjU
DFYTDCFpvrbZSIVZSRfI/VFQWpbnT4MAL9A4TjVnJvjx2glM2pt8k3m4Fza+1xGBvYz6QzSkUh94
/9sdwEPRgQIGh9rm14Cb+UOlN/5mdPuFjHK+QEGxuXX1N1OGFfjnk11oPtvdPtPZkrln4TuUaPoK
+ZqZIVgDeaRx9KbwVU9JJcqkYHgjsTH8cjX9637nVgAyzvQkSyKcd/Tmx1R6fOy9bK3VHLyfPcq9
KYItBixNMNEXaWR/h7RhxOWeayg+jhrxAO/kv7dHVPaccQ73kd2b6yXBChMnt/5k1LiNjrxXE0g7
MLF9KYtCwqsH9u/ngf1OStcjlLZBTb34fmsuSL2onSTIGZpHTf9E+YCyZqOAkVOcOmWdB6nVQRJI
DHuoL8xgLPjh2BJxFnwk8rM2CLu9x0dzPcVmBHllzOLh82WxiT3olOarqTzVWvuOs67ZVcVuIeSR
5rEDodXS8f1VuD9CFSro3BQtMoOc3VgvoWMBf9jnAsrubFLjcXL9BqyPA48HqfRl3bA9zyP7vlNd
hdHbjcPJZWLR4RWFXH7C6lS8ALVKMJAwrSL/ocA4CFlqcwBER+hIMtWJ38KKPSyZdjLa0btw4Pn/
aFZ47luEu2vIk05ymaT8yB+168F/Akj2Wp7tNk2MuxwcDoAWCsHg4R1cQSqfjHrD1n1jcjh9p0v4
LVZXaddmqFUwQq8wNieo6fY7/6Rgpa/4YFT7oAXDoixqtatyP/02P64wv7/C/2v6lJ6kj9UbTtC9
9mWRwbuWIr5F+VhFbqneG6SeBrqR1a/ZJJMS+j56rkGIhL5QP4IKZ8fpX/HXS1o7KPF+Pxkw1aYs
6+qmoiCTOQXorrBu+gy6caARjGTPw4r0LE15nRFvpJGNfoFPkJz0kr/xj9fL4dEpbc7yyctFjMHl
Te8PKyW2NwCyh9CIB/KT1rbwXboaUSggCJV6YfM4WqeXs08/1dnu2N73pUFSIXLNnoeolo4Khghs
fjhCxDhAdC8Nb8HU3T5Sft4/ClBWDyHYUxYYTzisXljug3KET5wIC3dI0ySyWds/RzJxk5EJFj1a
HE6Y84MTJKVv327V00CBmtstUF4Jfi+W52Nk9rsdlVvDgmJ4Vv8rlJglL92LQBR/nEIya/jYi34B
VpzgTVRAb3A4U2pe5xoMbVcKeaWrwABQ9ZeOCfuToXwi1aOq0TPsTA0UKvMwAj/rzpX2+g61S8gk
YAHUn1s0fPRdCQAWjYvKOf5Vl/Ab7h/efGaVrQzIr/qjaRWX6zF5cmVOBhSqi4BcWXA+8VGgNJX2
u1atXDyKgTMlQimsrc7XR7CaSAuIqlzBRsZUYktaRWsUEprDRvX7818q7NPzlYTKrjD3qEVva1Ci
tU2+ykxezcRR0kiYngMv+A4J6F8ppC3R/dDLdPDWDint/KivHPFVXCDDoHEQ9od9KRCFi1Ac709+
d6TEx4IB22lzJPybSpEBRxy4SG4swripB4W9bLOZuvtfgg2WbvSMrfnlbt9vVWDPsy1sA0wA6jh3
qRQ+F326OlYKUuUU1xSFXUXTW/xIHtYKC+U2JWIWrNXg84E6vehGizOp6Wjqm4cI6vy2yeM8rJSv
IgELvJxg+UWoEBDuh6kvrDWCHc4+rYl06woZzPtfcV4hSJr8RjWBEsVhythUUMyHbG/2fvE7eerU
ZuGwTUr4g9/fWjzSlVBGIeHIqCFUlPAxg81b9H76Jc6iYlLM9RpBUu1OpNofE7HM5GJbvqH/FEBP
TQM2EK7+0tipG4bKJyU6Dm9bbnhOjMsxKwS0KJS4K/y6rCti67UMuPVtoQoHotAMmIvOnbWYlCq1
geNllteHwOa3HDBvzbWhuu4faYP2vG9nbnIlatD8rRYyAVFz921B2hbJtkkKAqNLkMgrXV7GRp1r
qMzBpexi8F5akuhRQsOpnWXJplVwsL60JXdwMgisc5HmSHBfiHSz0M6QJ4pzFbQLmlnlbiMzD0KT
CQkBF2kyfuvj+78BT76ICnRCWTiFTAwOjAAGMMpkaIgF387eqNyE1ym7HT5d8dzVGn3zX4othF3c
ZuA8q3Wpfkmyf0SFLUtRv9CvRccWrWC++shJuQ8IH5J/pCfQyKBtWXcjSoyacZ/piIgGZ+NjFpgU
eDqk79QGir2K/groZS05GTRY8ID/DMING2yaTgun/trxueVScNehR60rteb2Z1BEKOoie8YY3ctv
PIFkJRVocl7D4hO8A7Fe3bg1zVeXVIKHz+sbC2n1ATSJnx3KTOSdt8CGgbiK9VDhWVkgsdCZ7Niq
66VRyrSTWxWn14XUUD5w3pAnBPKSqgmwnLFeTcXjSZsqJNoGNu6RbyPMXrEnh0F/qRQC8mBglI5X
kBl43npZPLB/nlmKTKIPB5DVbOslmrk5caOjot8v5m1XstoKoJBMi62FMhxmoX67peoqhNRJe8s8
0TQYTsbqw5KybAjuCwiBO2/0E5OS8Vk1nHe5ijbU7lmr8U0lGt99LkfHxVPJdmkfhwrW75NqWvr3
58nkYfVDvyixqqgi8NuP0gjJ76rGpMLfdt3+eKn9b+/4a5CXMtWfq86Oo0iVoZpdk8/fsa4l/FEe
3ZnYh4ybKxa9UR+Idq+BS8aRAtoftiav2Kro6CO+o8oNG9/1mc44XTEdO0JfP+wZjj/rq/iv9fhh
KP9yLDphdUk97blejRcF0k7tVldUzeymEdUha38lKYiq405/OPoE+R+U7mgibq/09R94VMFUydy1
463i+iSh45NYxHqGBHKS70Lb7NX3dgkHykEo4OjeZQRO8iP0fkIo4EAU9MsP/RkIbxIB/QFZ+yqR
iT5g1lwG93tmPFlPuiQcO3eV+rIY1EF8rbGHW8NK1r9vrZQLN7EHhOMtvk/ZXUQ5f9PCMIiKLEWI
s0cu9GJdxLjp2Qq6Btm8HUkUtH5sBOuwgaqgkV6VDDIaEUPM1X+Brv0Xeq23KJM79UsKz2d83D+N
s6BObv9CKPtJ0J1Fvd847HQ6Vtxupoeutju7qIY9FYDZgr22y+UaIUGnXt8dyhFIoK/e7p4tL2Wz
lpIqVgE4eQbWq6Zfmvt4loRYahBQkGgwMCBSry6L2JuJR3TX8lA/mOff4suC+su3JFZQ+CmII3G7
pzjlV9SsQtEo4mt3HZnIt67as1OG5Iv1Pyi1/hac9gzn6bZhSlsD/j7IwbEDZqGggq0441bmeHur
LpKPyzSo2P87uxHCa/lCzZU/cpB/8avUq+9fu+8tbJxB1rO+W9cdXie/jwVcjH4pWAHWyv7FeUxu
basB/649k7gQGTVNav77JaMr5R+A1PUNHeTYwdUpWY1ehxda5ng1pQZtWZMLP4TeQ5HsbXXWe9Gm
wKJtdvZS2YSbIWA25JE3qXqOgOvCSB73sZAyiiaeXct9KNd5R6f7jzhJvoK7UMGGugru8H1lasSF
lzZBrRy9IgRHARbRUxnZUuoohK8NC/7UbQ8KBI5OcYbwBQWRC8g+ussh20H7XZhHtkSe/OaIXZvb
yrMGsUPUJ59BTPfGxz97/QZaWOtKEOChmtPXwNtgqBRLG3LnGefEMuXzfPw2EoFgfoFI4JMbu7vx
EnMgKHWiAiQ++m35ZLqCRedfdheqcR89hLBZInJziFkRSx3xOqvTFqMu4ju4K3JLwVcSazGGHO4D
WD9cmj7HdLpqThhE3e1RRPj4K4FnIS+PAwX5tkHjWYr97UgscHywszS/efI53Vr5oiPgjaiyvI6x
G6CLXZo7m5+fdVdoNv8EpWd8b1E0/2C52MaOJvy4tGijRSxgWI0xdZm3aMndCpYCY8XOJKto4kg7
hgScJ+V9lCN886u9ZJgbnittdNFThU0vhQeeYJ8dI4WiQOpoIEfzTTIaY7fBDIT0+Upqx3DYPlMC
uzzrv0Xd7lOvMiPSPNlcP1o5xArsGYJziuEkNiWBuw9lA2uH+GYW3zu3JCKsE1FLuYzdKsHpSrA4
nbjzSqEdWtprJPsI/t+donWC0jeYuha6MqJy19eAkwLbS8ao5N/mlto0L/nu/syFz77A/R3seHtn
aqk6ojWpzAb8VFVRavYCJa8P0ZCRDPpayliD+BbpV8biP8u8dIKuoGlAchPeNNgd5dVGBxX0QPkF
Rzx6Y0AE6m2t5JZnjVhRAZ5vP+yv551uM+vMvtI/33nzoOr8BPOSUGVCMDBPdXCtXLPm0h+VmKyk
6HN3VxHVrUq6tEp9treOh87miiVO2j99LTIOAsDRukWnVYY0UGNbdqY0nFK41kaFCHdFBGS++Tbs
VYdNx1FDEeUQ71F9yyGgwCTbYj9orS1WIsY9ILO02qU0TVbmrcUvfPRvv5BGU0YbYXtA07wHX2dZ
zJKqtcWvjAt49eM6LiFz8SI+u8C4ivlv0zvLKovbpa1T/CwpSLftqKv1lLy82xLqCB7aaBO5C8bo
Pn+wl/i/QKva4Yd9Tp+iXgy9oNoWcZFI4ROeHgq2R6AthyAwsD6FgT84WJGAHmeqFMKC6+z/K4/0
wDfPDbkL9vHVSRljCSr1BCV+Jc9qfzLXrnz8d5+JUwTiBcIUPfqnN2yjKgRg950JHovPcTiW/NuE
S48+RXbfRzcAmC+kma2Po72G7BSHKhNMtcNSaAXhOlglPcotFF8xA7HO/But97QSeVl4yONMELHC
wtc1dviZ28EU1MsgjumPduIuiTY+9aVZzFVLxq3EUs7cGDUOKYpkD5shbhgQnah5410FX+BR5J/Y
FnYzO7blMO6+e3RmcKJhs+xLlEEvzEdG3bYrPWZK1orr5UOaRfQMsHnQw2Z3eQLl6JHmqFM53W2/
WUo7CIQ/5qwBQNFNMYgLqgrXl8ZRx9mBptu5Zf94DlLojiTMh+lWP88OUyHuTMi+Qgs4nXf6BDos
bluns/m9weM5c8FivWIasMe+ePcwpB/AY8G8p6ApWVqiWO2lrt70+CrLbMQ2TZJa/6QLeZFF8Sqs
b+9NTul4N6Cb522vmqU4T8WmZW/0rOqWzhL2ufG0srvJwbx88MAdtEfwj75FrMrOaKG9axsoPxsn
ClLyjmfrYEKinAIHxjxqxIBXEp9v4SI02NCp0bFolXT+qZ+9oHVrkNMIjpygbvp8CKw9vLWsp8X3
FRxbFttlI3RHgK2jdCEjXtxAJxpHsIbgj1OJuEq3CT+M7G1semt2qupFkRvu9LD8an+6ClSphIM7
ASqzVGQ58COHtqaDqXeT6a5T2sGafUjh6uci1TxTk9m5Wc0VdC4Dj44kedozYED/ey7QdOZmRGQa
mnD/unumRok0XikAtaBDjy6dL5BuqPmELyAikHBER6S0cUao+PcA3MXhto2ibyPVWo/KaV5YUnaW
sfRDJMs2W6MkyVX+ezmq4Cdl5l9KJ6V8WM5U38CRaFKVf5awD2f3h/ovpdonfIBUUY4+VbCnXIdJ
eSW/hFJldcoQoFvz+NGDkWUyi/ipPZiiuB6bWXgB48JPmYe4dyWTFMCv22Rle2uupZSclxERojGt
NI6JvsuyYG0aqvUIJWYWDtXSD+Ik1xFk+C4QgodelQEEQWGqu+Ll6Jr8EjbwQ6u1HLbBSVB4WEiH
A1t0ez2QZbYFy2L/Fyu7RIGORdJy6x1aMRAhm/naIrolYrwGb02iISYU87ehm01aZz5JlUCFwLYr
2hahZF6WYX/36SVA4guQED+x48dbf1FIGM68l3VJ4yAoAcAfdPEGKgK6o6zazvNKbSCzD9/qHUgR
uVsli+y0U2wn2lLKYbIz6Jn5T/QIuXPtH1ZvG2eKUsGlih3kDry+GOsR6CMFrEsvDWYg9xSYVxHX
8UIeAYq6JSqbYHsPxM11wbZuga4r37TLxut5gn9OMX/XfrneybiInW0500v0gwocRn2sswxMJpqH
mV1l1uEcHvnNUgAE0CzlhhUQlHsniV/DghhnFhO+Ee3gl3Ji1bTgO/ToQKZoxpb844L5hF1T7IRM
mqdtKIbQZiI1X+p+XmWh1UtOvrgNC365oS6dOelu8EF3hYT1OdImT6WjtFhWXIb/k28q2g3I9d9V
CNV8Larrp3DNY1aqcFKgcQy26aeD7K0MoqyTGbnNR0cuN6DtNFIy0wacwoGd7VMzK0Klww7qN41+
OEN4b7Q3Mw7vtyfa7Iefa7kaUckpPYG6bJXzgiOeLkWX/JNAUhIv7zB6rN10ysm4HOuf11EEUOXC
29Q+EIQ/Xxg/cMVSgBz9x+qPT0VhbOkUnfSVGUgvlZuAuXnqv/Z5NyJN+HDi7mRazDMA5RC9dKPW
lJSx1bFqEepN5N895yk01krzI5rFCLuZE6FBHgkijf/t8xy/of53cX0mAXpRkoUCgcSox65CB/m/
9lLoEA76j3DSc/sRqb2XDHisO0hwSMGYx/tgNrO25gAiuyMIpphVtn8Zsqh6cHLK0HzYnwnpquJj
qVhKUN/mtNfLic8/obyKaLiP+mrd28bTi7iB5B/4KBpg9n04vxgPsdUWcWakFZC0SifxGZ9Rd7BR
IUsu3gUxp74gxnIfgjhPGzwGXFanDpwis+k5Y/CMLqBmzacfzOIfJzxqyCGtEsgmPxgG2/yNoGM4
lgWXoc8nYONrf9co8R9RHHuXVJE3KfIY4qWE8m/DE04OMlnBfZvkyri8aX8zb9jQmAocgVfy7lai
8UqgLHSA/SXdSg0XkHbGiuJuPgh7h3daVo3BBkHFlYLioMn52cLo7OlTQuiDHGh1oX5AIT8NyQZ9
StL1cxMkD7Ffi1JdiBOJa+6Jkpc67GVDq/76xdL+kCB12962TzHDTCChQBG0L7OrQdVus7cCWki9
xBH+l+D7KanrOgewEbB1jVYNoumaXL2ta9Cu4wI2opBkBIq+6lWbHNXcbZJMw3GFLsO5egTtuc2V
vpe+gphBzaRpZTdFp0F8/ifHcUDYIWHJGhOJvpYwIwtINqmfgzU9f0IcA9UOO3EEvbAzVvRsLJx8
z83q7AGXwrojTmeHzSXlAamnSrOMuGeVvMPgw2HM7dBX3l6Ma7MhCvvcr6sjF0gXoqLepMsI60SQ
+8+ZhXeCWGBSFveCdviiUd/N63n4vq6U880P8Egp9vM2QCKH78xBmUQfBgrBZLHikBZlYeMhHdSx
g8HnZNIjhA9TCp/t6mG3QCmJQIZ07jnzFo/SYRw5HYyUBtTc02CF6/L6cLyoETAqN89jqVqd0xTf
ep2quFhWnLJHyN0mPyxfsoXBU3nZUG1ph9vFtNXetacnWwOU5I9xdrXtHDszPvKZv/XccSs1+8E3
S0t5Fm7EwQyalYip2j5CKXed7QJAbxchJUKfXiS4mB6nVDclAZWBa262sSpJFHFhcheh/uESTR+7
HPtpI5mJqNyVyZKPCUHGIqX056JKy9ZHKOuBTaZCfIF9y1fiBUhYKkm6+baxat/4vcMfC1LgRVpY
K72+MVhnt28Qmy1qZWZ/zWFgNpYnqOIxhlsndeiMbifduvf/b+2/nER52lT7mgMv6el8O+iTRT/v
umjEyLD7rfIqpt0IRUU1x3rFFgG3ZQ2ptJmWfMwqnEP22hHTH5lpMlVPJOkUr13E/XSJYt46XB10
zCZdZCH3JMz0kdW0vdQpomjbwruuzuJEmLcKdVjq/RUZEwvIkOONL8J+eCVRXg48zTADqcLPi+2j
P7E4A3jESBv7sqTXJnBzAyblYU/SlVVfu71bY6YtJibZNdT0kmXG+C3lXTGE5+z8NO8p3KW9qDfJ
IyjYlNJle3nnsqrqCnxkNKxdRTVFlJ75E55pB4gD8a0fz9qaJON/OIA0zX7VVKanFN6OXyJkXrJv
2uCHt+duSMCse0OOhDml6VR45c78mXRNScnEgt+lO7r7KhAuKtAFUDylqkc18wJeVdX2I9Bxn9is
9ZNjHP5U+GmRE1p0W6NPihmCRddqTk4YR0xNzNMdsi+m/X9oPma1Y91NpCoze7cILaT0nbhhY29f
kAnDDWLDQ2JrQPwAFdW6YBRJPxxuo8A2HiztERTRJSkdJkqxNEU49m4/UoMJSTSZOoSuQjJgzAjy
rcZFCdi6Vq50EjLlwSLSwKiwIv+QZbTaosx6Cua5C7LloyMmStVJVO0iMiVHGNMT1uGadad+vB74
jTIKJYaIPORAeYQ+nV4kQncI5S5kyp0Cz9qGarFuIV3OMTxO17CD/+xEd8xkO8Zl4QSipU7fVwMp
7SihzwQhEM6Afw5ddj11c+EZpZ3Qbu1AwhUyc9gPowTNAJsICFn7tczu+37aLvxV/pm2SGVtZ/V8
g8mBhUh3PA5r+ocefPHlT5z7pr03fgXINu/jq4LR2/dAy7FOfODXs0+wdH2iD6IDgBr1WCxPcIJP
7W6wBfkbrBcPw/m8XBnQStfMOgKaT0wC9L8+bLxy/U8rlZMoPFYY8sbCxlDmG4YwBJkclof2rjKR
NAmI2sRrS4XrGl3JhH5NkrW0OlauM1OruTvYi95Bx4Lszk6ZpGFrRAYb4vczYdggFj3V162iMhBH
tTxJB//xVQbCbpwvyqkJCxdeQJqW6X6TWk5DtK/6O1LHKk+2Fz8SxfETeZ5NrOyM1vBgFP3rkcm4
SDG1SOBGniaJ4AzQX+Ai8affkp1DBUOoDQw63T0Z9uhEtMNR4xRvp4HmrNTI2w+KfSsb9HQuPYFN
twSDA8cAyHFzbiDZUyWs2d5WqK46ChGn4sU6uDU/WD9pajPuphohO60VJuBLg4zXJr7sUXHkOX96
ebsGYLmyNKwxRyyC4GgwdnerLC1/+5/OL2tvC0sVi+jGfpcJD4UbvkdMDblzZ/0PnMK771Q6t5bI
W29jlyTir94BYLHJ7DswbgAQVZ7kiM5VF19Thf6RO0D/j7fbbuT0IrPFGmmrsCXZoY8BlTyPzG3Z
g53jMXqmBekttwQw/zBMbq9ElmlN5tsIlPxek4EJo3afLBCZC2WVYUMQTmXClQqz2g1ix5hatBCz
R8WJTmp1maRrDHow/6a0kS8q3Ao5ci0m2Esyh+82XPuZCjU/OxNUC4tjgvv+CP7a5lmqyc2IxRIH
hoB/uk51/jqC+qnQL8IetPtSs4XkfwePPW1OzFBMI9G0zd/UIUIoUKaDRNdOkyNBXo1ODeZXGzxP
NoIh5xIqrjsjTHe7IgdmI19SCGdhcPMKC/dZ4Wo7tZJ000LKzFuA7GwoE13gu8qua7xUVd/g0wa1
qCqOvQcnSKFTWIEz3xKZ7BH3V5ar4/fvtKiqr7KLd9LSTRHrBBESWr4YTPyYVdurA7RehPCd2xUU
pOy2ua1p+nkHaS1eU0N+tq1EhfJ82DwwgZPbx6mMTHigZB8EGuVs73N/g9/g/l1npxWB6dJFjFYy
YTjqVoqmxNehb1Eqi4hfb2bwFv5IHgd+hJyboIj+oC6DAvUwXT1p9ulDQL4sM0cx8DDMaZLzOMid
LKV87l8BVphiAdbLZQmJlUfw568A1QPCb/TGX7QSyCmeaE5O1rlCm3DogQ9BTSfgDXuuF509W42w
uCcmjyLrIiGoY/FeLuFeTRS2cDL2FId59Hw/aSSN3AMIVAlP6x4fkjaGM8UXgHkD0UyWGyIQtRyk
HJHi4EG9HwW3t5esIxFosLogwSFu92eLFSGhY+RmeEExqjwJL0DRvO7fWuwHa9iJZZ+3z98tpsHl
bh93W8uZF0v4FLNaONASBb9PjF0HMlWy+P9d2bxxqS5Bn0C7rezY/WFipLygp7knTWFmPqLWn42e
ky+ARIoFtf2JLiwGMRNg2labwaHF920rWnHQzfBzgvlYKc3IV+T1VUrwPNCVN/v1FcjlMzTOQwFq
Cf2Ed4EgGZOv7xUIfRFZieQKMvRONcI+NXnyunV6xBzf+RHNUPyYhFPcBdHVc0BIo9Sj7HELe5Z3
H7pxhqsj2rRPj2tkWP9c+yRGghJvMIguEhM8Us9GpKljvodJPVMkNhJTzi04Ih/mW7pbvUEk/+7s
lJZkeOmmASHBC6/kgao9mu78MbPWT3FV08NOsLGZxLUUr7/fZPpvD5JL+tC5ktzbsYIHvBbKBdDv
SxaQijcHyXujtyxY2R4yaQ0kTjMh3hMcV+GW24xUD7rkoYsxUgaMFpEnt1CBAUoPB8pPnL47l2K3
tdG+89VIDbQLCLImq/Xp6ohsAFtvpXFXPQ30jFp45mvu8F5uGsc8Ia1BVbkrDKPaF5Ik4PYVJ9F/
7u0iseNqQERD9UdzYz86A0DnmXkNA/Lf8SuKQ4O2sr3PyA06IXBJg39WbVcA02daDSChn0Gdhyxj
WRwIhLAr79fIuwe7PMl2/9gnfoMhmi1JoplcHSqk/OhJwqTY5s5hi5W8uxR3QgfsN2YFjJY9QRXp
kSkqpfCK7JKN7HvOf80rKjlDQvWl1iss/jbrtVa/XYVurfTDL1mwrCqyHnY95/NAsL1lQ8U3WrvS
uKwHSpilwfNBQsugZc+325KB8BUtroZy42adHlUNMyse5uM80KinT8jsAiTuuGsIQlgIWnTXY6tW
Mk+7JoMNAd1VgQBTf/nPcIru1jIE4U0Rzrb56+eJy1287auKrbTZBB7H/AF96uTsCTkQR5F4waH6
N+P5CvHRf6q54UQw4d5R1rOqWfQpX+3yMH8P6aU8k5mG/1or1zWe77GvB1/cfwIBbVTzLueFFWGD
BcUCbhzKyKiLsgEYlhIEX26uTJU7PXfxhgqaiaTscoL2an4GKRt0gjPPSqCgO6IxTix0sw6DoNpM
oRa9HuueSIKMDuUyEG6Bj7t8nrDJWqO2RiRs6PujG5a8qU+BR/ckLzn1g0eE+mo1g3BB+vei5lyj
vfjodA7J37sDWB52IR1vfyngEpNuSjAVxO7XQcscFEw7ohu6pGBX3E1gcJa8xdEHD1fCwO1zt/zP
V2Wq6ZEx8DCJq9y9GMSAmFexPklOdXy2uUYprwmpNylNfA0Y/u2Ewmhmpur71Dfq9fCOeMFFFXgh
lyJZJqiY7GjOE+FpRY/Ro5Td9AqxwkVufh5J7XiQJ1NjOZWayPenIH3GvYh9acb1Ce8efjXiNrIm
ku9LNJywEKMF5twSOCxVHkv/CMsVKAFovJYNG9PU8rhmdRiuQ2NfTWz8Pt3cZDH82UidRcx7MwqB
BEOK/B1hkW+nU1ooqQREpIYmF60tJc2ZxdviacB13tJjmdXBi3we/4l7QuoPSVTEwCnJYf+cU8Dc
FsYGNCBubys+vhibYgbRWM31ujdS3v7+1H9mgaY2N271+iuzf6d7EIWM2D9sQpQcISz6oolqSaQ3
9yRXJOlFxKZSXuV9NrWXZMOlIiov3kisUhTw3w220V6Dg9rpOPng3rJjUncKP16oonieaV4y0HCA
zvj25P96edWhCX8006zbQXdjsIT34KQgj1tzCAdyAfzJslkbkF9cp1aOEN6jopF8XwzXT07KuaFO
crtvV7KI54f0UzCXuWJLwFPQXnk2E3s242RuYuyzM4dzlQSoi1+vPpVBMP6pEjnFio1n9PPaeucV
6ka+twQsvZul6+oKvj5TKgcMQW7a1vmFLmzed+Yol1FDH/yLgbQe6Y+OyR/p8WRa6GnszHykEkYh
a5Bltp2BFnCznaRGR5YpS0EOkQlylLCS4gfPk1GDBWbQX+/QQNE31x/kk0jdtJiu+kPvyvdSDRU+
kWIJyZJEJNg6ZYdbDGy3Sw6KaBcGfxCteS/Y9G04vBDbC/7GQBfaUBthfQoVKY9JIPOOpyF77O2g
ktirIO2+AbrbF3jswZpyzqgHsV1e45tZnVpVBGPkd5isR1bn6v3jCdw6nG8OtNYHkdFW3bjlBZG0
M3zSMJd2FnmoE3w/c3yp+tcjsVQcsdAEsqnK8JjRuTsrSw/+Iq2T/nQQGZZM7I5WSw3vkh7a0fiY
yju6CsFubpbxE9TtFeaScAuGQDuWK3bS9ViPmMUAXxozTuoI1l6M1nxWTcmH5jHDahVNB3k10YJd
+V6MPA3HLZPUnftLOUO5qCTaldf8Cw/9wLeZawzNpHevUDHiRtaBXDAfrUR2K/RNd7sgkn0yyqQE
GJJvnEsQ2NN0oViKtVWHjTaawXFPNouv5vg9lAneGdfK9wVO3+RlNNH1UIPeJDV9rFQkohiDgb/i
csGNSuVoa0aIAM/97YIyAInl7fgJsEOAMabqGSSIkjsrEMl2Bi0kGveh+XkAE9+MXcGZLZ7ILvVK
TaV+t6PnvcygA/Yv0A7MjvGP37J/RnWxSHpJ/3K0t+leM3l8GjCPYTfZO7e8rDQ/QhuBPBbA0XT3
sMY5bXaywC7ojARHVFpq+LRCadck/gtdU3+PGe1f54I41dKCA84MyUbhL5xuW1Db28SOCYgxCrrP
Pgd2xfpuKcDr1Aop/3G4Tl2VVA9yQYIMZL5YKMU+ZgJToKwXNYW1D8iRDy3wsyMjNSc3RLBP1ajM
jxIGmL4r3yO3n7ffo7y3F4F6Qppg9Ne6lPCSgmt7KNB000cH3HmRoPTfuJUzjseINGE2hj5gFd4N
0blZyG5hRbYFjkbgcXtfJGLWTwdCrcur3+HWa8SswPpxO8ikpuGwyTw9Hjnmi5xKAuYzdWgFUZUj
Cueo7rySR+wJAyHIOkFtLC//wqEVqa7EAYjERlJdlzwXSE7YIMeYaWmsZtVZyHpcjrFItF/V9vdf
ODW+zyPJa12LUl2hWJ/MveXilZyh6mBW2oNnuXLvIFZoIpjUwYGwUrSDjgX1SB8AFtEiyNlyjacl
PNwOMdjjZJ5jLl0lyhBKR2/vHCqP5NOuTaz1Josgi/o1t1unjh2BLlaK2QyDodN/UlDfYb7zbmxu
3a8fgvD+/vWeq4b9KPhodtLXmBPWl60PlHnDoVf2Vr5K4S/WiNEuyBeRHJe4MHJ34DR3AnA+eTDT
gEojEcxtt98dIBbWYA5ApYw5dKY7tyyFGjwjJI/MG2at4xV8OoIZzv7h0XOcER34M8wiwPOUfmRV
sfRpvVIS7TbSH2Wa8Kn5y80AI0YQn9L+ArygdWquyIFbPzYh26V5r2hV7aLF43sFXAlXqah1rQ9R
hfLvJoFdEnr3mvObftoGzg7LSCwyWEGqpy7CGxocbF0m9TVjTtDKHtc0E0rlNEdUTxam/HfrtygQ
GKCcQ3dMH+dEXA6LirVELMcG8hJtwzZ2EOghwdLxowwpyeRoqoTNJCZl4v7J368nARd+4aPPL2k3
PeIcO09sMFCIELwDE0rP0cqddH96xqevyGZI6NMwZ0BDXodEgMs/0yjrL6O8DgmgS102YCYyDWeM
Iov1A+b3KcVpiUwhsR54s9bkHtaYmqFcec7nsZOiPCLMr5fyHhZjrQ0pbcTCqfmWbHNLgCKxV1AJ
UheLvHrKkk11jYprLcJ0ezQHEGPHV3QpWAbZR9o790dOYeZtKSrX2JDnv2/OZlMlPdsL39DmP7UG
Qso6hTZ4Pfx4YUh2z5xG2XLdqLbR36ZsZ2SwjQxPb1Wmf1oY7wobeVxEdTRTVntX9gFMdTXDrYqU
T+1FtoOXEJzEy38voIefCem4yzi83fGt3UuqWXgHxz5P7TvMAS6QMJDPqFe/MMzu0TX7Ly/aOurm
T2YhXXULX48xKD44nQUidgf8mbRrvnIe5soR6GjugBayvhi1HMOcKDEBrPtuPIg3hYzYadUyw604
ItI/0ft1HPkUrbe6Cxa/aZJiPEEEu+B887AEhw4MvkXhCUGP597JREgMHdXH2kR75IGauOZ0nZEl
YX8mhsvFL2HM5wU2Ae/yTs33bktG9tCs/2M+76yo7o17w4vESCA8wUqRYRmvz7CafKfWelPadoyR
XGPmfD75BnJWTf6wjTdzmh5jxJtb3kAKKSPK8bubaZTgz4zcn8MOC6KWSDJLWYIMPRGH13mBhjxB
OINrhIUPpX2TJF1pJ6ahK/0+X/sjxFmYEu/QO2cQCx4k01lb4cnHB9Sc0h/fEHceqf2RQRTs7BC6
esPR0cv4GjcxS/XK6DoevRjf1Mo/jcWhdlEYWorfqD5GUnsnhWR0C67AM/RLuO51qYV3ZD4vC85I
/0TzWUHyJQTW/y5t1HXJXqgLqUZTGRdFCQFi/Hnvy/IJ6vxfY3OtNqcQN+6GJ4VMmHVDC01/QPZ7
umLZt5Bqx7bYeBhVyT2XSMjw7GG0zc9w3Q3cI5wDje3xcTIQ/CLEOrrci/kldGd1+HP7cn/udY32
EwBoij3rrtGS/5o+FVQ+CFLrUlNGr05Rfbj5gSGje15ahnCpEFpDXHOXdN3MDfV8Vukj67LzJHNz
TDsWIzBVHvwypxwUWpmYvqXlmVR+lyBwOB/OcxqZuyyCnoJsFDiFIYCHE/o//mAY7PxvET0V5JUI
TcK4oXUkyNCKmp0V694pkvRRDx5ymrxqmktfO1HdMmjQi8lHlMI6oQcwrJkxw9SyusMsEPCQcGH8
7yVKe4UM/tMqaQic+73i7jDgfQgOpBKiNu6lHFMz4XWRUC70F2nDXYQElnPqd9Cl06TbC1Cig87z
tx4k1Zrj6RZHhy7ASgD3yfqSG+3Tlx80u8pbiQpWQRthN8MUxhLHSNAaVepT2a1n4kcpMxiWeOgR
g4EpO9ByY+B8u0VMMS2SSOaLi88TLHLS1GeIeBFITZBn6nau1CmdRXTC/4FcOZVkDh9Pfn4gGVPW
bg5OUpEzPmwROnOZlkIMTama2SNCQbUYqcadDbEpurXDCh6TZ1rPVSdlOg4a2z9q6Ton9g9/+PDG
fj9xdTmbbWV0jTBz9Xnb8lg79CNzBKOkiKwxXxgcZn5eh+Mk5fLuXMtpGOmU0bgwF0qHEi7cng65
zOiYwMTzGbizXU6n8w4+op94E5fHkwHm08BzU092fRKkuplFVaVW55YNZQm4cj4HjCrgS3b/beHc
XVYDFcfEUgwQ8hbf61Qt9fZeO243vnbdsyDa0Zb0lDFWsfTivRfeiL4PM1oUseodNZ9eKQgVnAOW
pZ0gZ8rfH6VDceCkA6fLTBiRwHSqZqmUfRIWFNUHeIKNVZ7NsxLxDtfMneFJjVk7BQDN/QqxND9Y
mli1wn/vawp7RT9Nrqdt6Y4IypVo2kcVDjvRvibZkKx7fXoM7rSsuLB2NPDxnTLfAf+GTGVEMXwf
Vzm4+UqvIzXtFXKrjfzR5Mlep+I7gPX2HGZfGsxZRXv3+chKwxvjvrm6qA7inEsyCLO8AwNPLPdt
H+ZiGJXMeOAjrl7cRa+Q7vQ+a+xS383O0LQGyXXnIEWhNxaJ1oE/cvtLnaSwkNGGXPfYS3eiM3Y6
paiH5NWxPhSrXXVSJPJMzRRUAKFaR6gooxv4wE7xGejMUPPHI63Jj4PUMu5DMIlp4lHylNhXdK62
drTn2OufRAb1e/af6PixqvmdT7E9EEZo/rh3Brc5bMnHNLGA3XRVnpT9Mb0UjYKn1lZ9kqIHw1w0
HsGHbr80LD4FkGw3rzWiOknsPsIw5d6dVAaujMWi8u++IBe01fDc+vl7r6KlNh+HyPm0KlJvmCZ9
+Xmr2rHNO/RfekTe1RBds8XiAqhqzKrnfdk2cwSUqJB1699pVn/f0IEMp+dOo4GiMcywy4XIHzqs
TCdHtGJ/u1RFj8vXPDujlRpEyTAOeN9tk5BlhoZafzaoctj6wD3Yk6QjTjJAfOdamhN5eqLhMqPI
7f9LwwVofJyKAZaKvplZUVxBdd3ZVG3gHxq178qj05CfaTgOYV8mELugMdeIMofwFdhFR11GU2Id
w/O2CqbhXLm9Vb5Bwlu/8yhA2Daysp+itaqhtcq6GbZq50VLnfU2mKiOOEV8rINDHjF4qebb/eSx
4U8n+Hl4UgFEqgVRIJMD3FWrI6/ia8hSQy466FpZqUBHnFMiez25QzYo7kGRyitFG89Eizg6sv35
YCRZnHxtYjY+6cVS0jCXxUT57PFsNbc6WLb5TasTLisS/uKv+d+KY/bvoQ2OutZXG19+BL4ibRU2
OQogRSrOtyWqwS+Mn4OfZk52xuiocLC6RZSkQb/FUBlIxYomECkAHh9Utb7l2Y5re3uJ+DnGV/s8
JxIzENvF/20Q7pfpaJ26oUIcx9jP/7VDDDrE+FCyR1gXXvhBDHgpyYgvfCIaAzRrM3pyqlOtDj4a
9ArARxcnIhD/XYlC4Avbd8+OfWwLsfI/UV7NJzqCpOvFpeZAL2zSbSVK4v4DgI3mDtq4kIKPLvaY
za/Hm/HO/qwYroQeBNVVDBxvEf0kj2i4Wa+f5wZsv8NwjZ8C3yFseUzck4MXoa7v6SMnvUnG7WiF
mpQgy2zwSCu9MDmOMQohtGqqdxprzeCxeomEo3k2Lz2ZVgKcbK149W/A0aO1t7Ft40geLEp7WiM9
6nQX7vTu7DeOjzrZ6nXGiYhcr/gDgrbd0KdhT9/s4uyNpoV4h0SUzLDkja+cL0NF4LJjU7b6+LbU
OlpXESLUQzm5bNjxR9lsuUt7WolRMfixtzY7w5Vqz6f1aKBy7Hd1iV451wTc/Dq7wPrfj7Ex5sUV
Lau1xGH7rQt391/Hf3h9DLEnVxlz4jlbsCxUkZgxrJZ3mz0o+gIMGwyWooEi9+0jEU7zUWhJL0Os
1SZ5k0gUZlLigqPwoo8sIhbfWaNoyVJ8pq1DOgjLorku3Saxt3CdYWqkXRaRBJCblTZVZjuEYCIb
pdMa6oPpkom64ASk8lhTncBIGCkcNNUGz1FXSQrLEk1kRHDuShqDkYPosyg8AtN8mjgSeVBGpQGN
H4Uh0ABcN0wPq8+ykop2zRsUCehCOWyM4Sycrn8mrJBLzJaQ9A1Bg8W+EsXvVLjIDp0N4YXHlekB
lHwJBuX8ANqHb7vj6IIpZgsP9Y5rozidNpxoOe5Q0U1TzGDSAPidr641ju3XVwkQqK4Xx7j2PMsJ
Kr6wsgbwmbbM9p8Qc5DS4iMopq55aIpf8D4sgO9dCjgef9y5Zk+YDukoOrk8CLrtYVZwTGbsFJxi
33U1nYO4WSqnfDFJItr2imQ7fkSu23CsvoXzkC78ToDtLv+fbzraqI8VO4JTBPyt2SYawZm9hfzR
1/FAFob4PLiC1zBMbya3JfR01fV7ApEYvf8xc1ohyxnzmN1cF3qKjpE05uGaCmLZnaiJ9N6ZwgAt
7E10pmWSWYjRF3d7mQ76AbOyuW194Yb1nWgR/UduzkqSMPcRhYdMr7/6EHG0QJ4DUGTbvAWqJ6eu
8pPsbrMEs2eR8f6jBQt3Z5/doqrjBI+nUEG8p15hKRQLfJxvh/mlLpldziIB/8CWjDPcipBMFhTz
B0/18AG3fZrB8qOI9H2yiEMHGCv4z4kD/a665QLiS797F/XdGMj4HIeLLiqTNDeQXl+VQ9ppHFTw
U4dMXhXisFV+lBdWHKIz00B/MxtGwXonsBGnQ/u3wyrFC6bFanNEQ9oBoUjEa/mVJE7P+KFj0HKW
sS4eada5kAbkOdXeKBMz/f2aBeBm1Ip74aAfQmewkK/EdQHjQ223VA/C/qXmxZ2Ie+xTUPCnOC2f
KoLEmR1pkXkJy2F8DSA6R6GJ2R57WWCfhv5/gbqyWxsjp6Q0OoZCVC4DMYR3++pd1yHBrfaZfa9J
QYGFV6iZ9qtleSqHS6qBiEq3r6VJ3jiNqJrtVthj5d6Rvu9PLNw1SEAF/wAMi0NzmFjcVTUlRfBt
ZaaQNY62FEZXrgt7MSxfSAGg+ao+6AlV+uTaR13TLE7c8CXipcSv7SxJUiIOLABnQWbFcB5lWN2d
lj+OVCZDUIQK0A9i2mMSYzqaD4jnU4z6URrtKIwhsgHdj826yPrrMhXR1F0a7B2O4446qG0TujTi
/0Pw7Xhmwq5zaYCBzT6uyVsJ05motTUM5UarRhWYVbwLMVqxRZlfXi/9Uq9r/7FKYJsqucAx99cu
rAEGB+EorT5MNnnpdv2njAlRkZUcES004RpL9vmb1YiFyXiy1svrkGzOjtcrO9WY77QhdfR1KBQJ
W0X4ldVMUPE/i7gM2VgDVk3asURP2ol/XjVFtx5m+gGlg71fFi8stwDU3Cz0iFhpHwx5HEDLu/Bb
ulzfmtWXAMOvUBIKmkN4mRN9fpq77t0j6Wnsrab2bK2by9ToxPEE8/5ATiy8RB2DH1BPaT/AtvNq
ILMVUSLfdbYqi7C4JF0it70KH8FRxmK3CnCsP9pOFFKgv5S47TkG6JJb2LmQkMDFSePsa0xOfKh2
UoQMeq862cUXbWHPcDP5Lv1c9lmy4N+ohui1gacs4i86JgoVTWhtTYTy9vAFI1Zi9QIB/dh3H6FU
K3kA0vGsOmJ8lt0PD1tnhyJPxaWCm29o+7PlPon1enUI2Iy7xOiggmq5/DYUS5XRCIqQv4ly4FXV
Da/4W44uZumPGFsAagsi5P+Z0bsg/s9CV4RYxpMmTsvvmMUpv52DstayOqgLGW3Sx5Mr4b22zqDH
3lRD4+vx4XJYz6oJFpfP8QUoAJNszm5jJsC6C7AvFckXaimu6qiJGKcJPDum59dB9+78tpA6cGoT
YB4geNQ2MptjGdHPcZvBBgtPnw+9m6WKF4xG7urdIWCue/En+azXfz4MoGw5weNlAQrVDULx+0NL
vBXdsJRsl980R948EmMl00hX0ymmJ+hM7v+lZHY76Jka/eMgziCBuBboLFuXuD+1fbymN/6E++T7
ZVCQ3XfGrAhaUkdy9pD5oOB4lRiQpWC6aKd+LPu5Gq6NnoAfhyJuHSyJQzMYffYzdwextFT/csPa
fCBxlBJEVYb4feqkFCtgEUGSp+Va81mJen2LWXVEhQuby0fXq+Jxsd1/UdwrsS/7JZefYOyGI8Yf
ps/+zBRzTB4oZvNwYqI6owhm2qoxLNyA2xTOZOBz7ax5gZUv1aYPsCZIvFCAMkj4c050jNlw99VF
NWdHyL9flkbMUxcHp3BsFfK8k7AYs16XCzD7FvJH7Awaq4HzyBHqeM710b8/D61ahlVS6bPvJSB5
jUE3E28y21T/JgTZPexP79K+cgGhTpRXd1TMhzJeYxnv3MK1nZ9P+rRFVSvl4WrAUDek91+90Yx9
1ssq1SVVxZPKzUyCC/gp15Mu68R/UbggxkLNfMTOkLRyeO0URP6KbQgWIbyXyV96ufjJtfnK0Y9C
zFqYQx6LkHOaV/yIX5batWm6UgHB89mS4EXteW6q43VJmswp8CzEwYEtYdad4c0/Xp1RZzRDSAZa
jSeZMns8V0KtgcSIvNSgPX45lzUH8SutI3uABUS9mXoJdpDJSjdzDn9stZcn6uZa3zDvOOiFxIia
7/uX++LkGSjEpzDvsmr6AqvAZpei6d9mcyjtSx6o+7L8RQpW74PkrG6e/Mp/iye+7hcIhxQPvDOJ
toOKODtYE4huiwvv0OD4PLy/VA5C9kEOLcC8RawwZiz3RZyrna/Lm9e7xDeu41wEs4xsTSZ4r88e
HJ8ATXGl9RgPUyHvMOTx/l0MHzMNyhX4HVFIhqY+sO2eq9i5wLMaXwyPZGTtkTLbA62sokrthV+a
kektJ2bkpQpwUHF3h1vJgNRqz6YkCY5PWSsFTkrUlrZqr49IxzCxP2ZYOnjDWE7rkmzehVJG9UUf
6WYN3dCTPb0QnGfMbF9zNNxMQUI83O8UdpeFVDPiIUqjdnVzYZoroOFcNP+3nzKVwPF8eDxSuw7x
sulq+urPWtO7QY3LTFgBQQIp9XwRsileCbsQzgwQA0rG7FpLeNOUAWfODkzP4cBUbJAlerqcZaSN
i/TYp7Gw+N+cvNl2iy6U5sWGf+fcQYcKub5472rLX1neU6nAsD/Rkq8WucacrafOwd8QlJLwkRFi
qI29Q7d5/tjERGTgKaUg/EHWiXJHkJuHt8tv87X5Fv+N88FMNhfVRIkukzHnfrCe8JimD06zNn+O
xV3arOYlW/JDd0SnhDtTpFmj4GyC8UflHqJmeEMfZF3zDrQn2QTS92U6MejMU5S1nOKm8vk6iZNn
H2kExkRKVV4a61jw7NBMyAWfUqKRd9e+3v9ciJIjg/key3UIYGUjU7jrq82jxUSYadSOsTKFchRr
trfzsB6olHyhBxmyjA4uxMDoZhtOc244lGkl5z/8wkQzoy5q2FzYQfyPMWCvFunaq/9Gm5ZfTDJh
aSbaSoG9nSwhEJUt4y87pE5RlcPN0WKo5sS0m5V82WWrLivsbY/XPzGjiRZX36RKWlXYOHCE1x3N
rAs8XpGaZkF0A7PSAOMXAJrv+0z0kKPL7TXRk9qBqwZ41c0TAtyxI8dwfAQwaELxBMQoqPH55Z/6
9HwZ/4LlyalnjTztUQwIzTojYa/8h9sdKzSnQXJRPoyScaTQqrEeW/cpsLCNS/gWyvbmrafrXlSo
IJ35axinmp2yqD4/ZDHOdDZ7VENxemCUCJLo9JQcY21XpBo1ix+WNNYXuNUCPbt96sdllegWMvJY
A9xCsUyL9cF/hunk/xk7Hk42ns6ypV1knYnZtJZmO/6V8cbyROtGJTFnpTaiR0JleGdL+i+Eib17
o4G4l9IGnBsb9o5nLzBR2WZlDNY49xXs2BeB05V2jZI7B3h3AX0VLap8u4nMiovpLMzXiIZPFRFv
e3cGrUsHti+s6Y/RHYglgeXCn0xxTKGKIBALG9eapnlgxCZhf/OSlU+Dyh5bIa9u2SrpxaIaoB1r
uxma2kUuBvjczoNDpy2u5H9m/uSFJ617lIzMxtzeGMzy5dhsob3UGDh9a1crMDNOV64YPLyPrY7h
CNfN11S3jBCytqsZ5uxPyswe+4oq1lWG7agM543HN77S6e/seBv+Qk64pZ3DLDJCOm/tPpTR53lX
xIkUMJY6ECQROvBpnPHJJvy61ivohw0cFRQqHsUWCEgYdgofGatw8PpXNUEo9oXbOgJ3CD+gU/tg
qd8bD47VCITMJw5pOEZFml3agHFHQO/LfHONWHfaUOeYL3tXlZHwIW5thfgWycX4qGL92TcAdtVF
byKzMw08iCTpqoHwrIhUudyjMd14zmV8Nmg1unexsXp3dXECO7w99oPbspdsBkNKUWzsaIRwN5Dn
rv+uZEzTHSKnyVsRlIINhUO42shB3A3pqXNLTVKbGZ63Lk0+92wpBhzBqCqVPNX46kahCQu9nQdE
JN50k+acKL+DTJ0SVvXWIRWWxox7L/xC3alXtRPZrT3p+SgQalbzkmy0AFy1k9T9Z2u6SBgtew8N
l5MYVlJvnHSaqXyhUy4okmvb6EJxiEmVvvcgm5qj5IMTzPZ6xE6jKEyAmTlnZjueTVGU/lao8OXp
Sp6Rgk7Y5Nb/LJmb4pkr2IvEzDQ2Ia8LB+lh082iBOiSuonuveoQWDqJGlOn/zk8oNLVOEZzwTWX
74/5Et6UnWqiEOM74xQKLvJ3H6mQo/SAXX9XjCRzfhs8rihL0eRaHOQWMvrSWO5dmvBMh5Lt7lyk
sl+/v8aH3aC03hgn3HLt+XGTzwuuYzQtnTupkXtw42CqcWztXgJgPfUNK9mUS11hEjopnWUy64Xd
9TGNofJJRkjaGp4wKZc5zfl390OvxLhMdJopC2BCRkOVBDVrtAPBM1gVwWwVHmzizW3mLuc1AxXs
B2N+HwPAM42Gt3wEXpR4IK6szAO8+JMFrBO7Xzzj8u94a55RySqHE83WgLuhX89/ziIWgOC23dDV
bNcleQao2VzCZCfq+1fBk6+T1TU+exYg/xQ2jQ9Zwf2812Z1pw5Abw6tedNk0nir7okOpljPwVe2
vqUlkdMreLwWqnap9h2rR+17GDuvwytIoZOo4EDMhRyzs+ghRwhAue3iEvdeWnda6s0hN5uhK64U
3SU/R+ztcu9RVYGE5IgecE/dU9YsXYhQoabJtR9DlTWxyaTMjzpl/K1IehV/vArlciIS49DStUwZ
ruwgWmnKET8P/whL1CqLay06JKo27yF5oSf9RBo33Hc6dgDK9CR/M93q/DixWJBmZ51AY9kIirzX
knZ9RwkRcK0jmVoN2ve7Bne2UnUBbmSsQvt/nIEFnX40cwdeATE/rfsSRJ32t/oSGivH1P4c2gwK
uLrU+gxDRuWe9RI7Op2i0VG3suEhYrwlEixbceZXQCxKqlc4PV5yKaMVoKa5RVD6WUrUI56YiagB
Y35MmeNSLpzYc7h4YE8mmIHJ8O4tnG4UqJqjFk8DfcVNMRoxPbHikb1gJtm2IsMJHZnH6SQLsE5o
6sUPgH8fkjn9hLeDyNv18pWzdF489iTqLVlPSp165mVLQ3ye7JJDxFGii3isTOUAsunuJHpwc/aS
TsP0S/id4nQDbpdm2U91saJ+8IGrodYQ/cDBlbEtJR0zObbERZ7tOspNXYyXSRc+5A9/04Bv8lKS
eLya1wk7r88f7+06bvZIuIC5yEJA2SvnbUR3qxv6U08XYvpUPebfrZQ9ocY0WKfwpiL/Zg+K5rm0
CdkQasCTmTRWOpAOjYw0CCjtDVdlM1vz5BYXYnL3011pnPdhdtetRSv+bta29Q+Tde3B8GSREM96
G1g7RNii7jcpXO6cZlUnBEzs9MZEKX0SdKxKxYmS0FA8JXwo2rBqzvHqLMWyGRTPbqd0OCRiozl9
fuTR+lko1jrG80+AxvOapSzLLuPReNuYYNioy6V/ItKu99p0F4JoHIjr19rtG6knhpUhGZXddl9I
a70S/v0TaTSfLIk4s8hnCgX0/fnfK9X2ek8tuEhR3ONvKHTpi92/kf/os2dzqyDOQVl80jFbG6+H
Vk8xrb+jeAmqhncWasypEmYvsGGBNXmr8+vJbYXPClfYtqiahRNwbJCCWfntsuB9Rl4PdWLelY5M
zy0BjrdBlNQIKQ+Ggabl6nLjUB1wchjj2D0eu3mIkUcRA3TdwyOFifHs1iTr5irBEzqwdW1J0M2G
+gaZWrpeRzVnr6frO5fqLUJk7r41NetxcAnu8i9swrJeO3bQsh0F8cP4ZmIlzxm1jeKO8W6b0564
rNsUynKB3Iyz0hHvqDAOFThQz8Yx/GhjxfX/kDdjjMdhpX9PH0MbBIZm9D5zUzvYYUJRNFGcmrvY
4KE2++885a57iGQfkpsXh6a8qVBNpZkezf0lAbyBBtjVb9IIWaf2TKrIB6pGX0+RILrcPbDHMgnN
o8Q5/P4XpQ1kxnB6SCHeRHAaledOqfsSH5TkGXJUg5I5A73AMwuQapf5MiUuhI3Vo3ITPlhDSB9O
Pco3oaIlKIFx5OwKc+QZ/TZ3PnuvCilYOLIUqhlYw/D41A8PiYwSnPs7oujpKOLHPapVvV/wDWJN
/Ccy6yqQxT54z+tO7Ja/YNwtSHHF9+w8CpTE+KQfSOhHl5f5s0IjCmM7gEZC9IZFq3lYRsJ08BvT
uk+C/YwQt7emvYtD3dvf8C0jd7KrPpvuCKwgG14dnFT7UJskn6ZIKcqruXWvzbXiZZnhagXAm2Yh
tiaiYXIcKGUrDbYKH7h3b18TbMVVQIqfJ06UUPNql9iXbL/zJH5h/nuvANtn4pmNbpoSl1U1guPB
Jt+OnESykIom8hb0XQEn2PXG7Aoft56hci6uswZD0t+9VeGp7Ge77K/UR9AH/78TgVs35F6K5C6B
FUsV9IKDwKtYVNb5pFbB8+CvHFuZMMVGOcvbKak70SI33MQvH0PVVpriXrH98d8PW0mDh9T0BPrV
aDXAS4Tt3GPIgQAmqeH1uKsHuJh6dnl3/7Q8D3fNAhHuohdauyqHP1+Noq9fb8wNFFIDERE/V5x+
KI1VaI6lrT7d58fbMwon8PMTRW3vNhu7qrb0HjZ3GtNGrTGkcNrt9dm4vK8iXQH3hRmpPaTLNi99
yPl1K+0hArZsYDyKYkRuqd6AhiJe64jN2Qyg1ChgH9DzGb8jGx7Rg92Q6SU7Jhmsl3vGKwDzHp0J
ZC7G9/rHv4V4a+/qKvwBaehjvBoajrB1Y4py5g2pslk11dQkrxG/QM8M/RKpBKRVh22qS6lGU5hO
MeX77+2g/9wJCbwPcqGGf1r3yy2MgpYg5Wl2zqfaIcp176Vlf7fA2ZW9Xkqf7S1AZ7BtmTpAJvjf
EP4UpjtlF/rd+V17IGw5XBJjyJVNx7WTtO3eKsiauBJMpMhddQjENC0A39/ID1jRLOCw6lnU9/fk
/O2f8a9z+ClEIWL3T+m48lsNpw6IEmOdFISe6zqQGwu3TAF24ptMRPDJsEaVTRJPcfocDVyRoyVC
RW1y6YinN/tzcDKakZoYpAZkhE/XY/fJMzM4kjE2IVMxOIs+L+DXQVNZcqtb2NHQ/FNUQmslMlOt
1cQrrQ4M3VX9xj68G67w0vxcFA2eDe5mT0529vJDQ2BJtSkj0CLfytSUL52k/P3TtcywA0PvAtcV
G6qchjGswQjXEy+14++93A+9cW98JcfSjEZdhusG2tlggBkguQ2qlTTi0UnyvJ2+24qQwl/zp9ef
EX40Y8WVwGYg/wV3S22rWvxYr8JS2/vhayv6WBofPjnd0qtm2JFW8+hIMNKl2Ka1pHMybs1N3WHB
o8b1Q9x1BYjlTcbBazKoN3sAnO2eyxFfJOirgZT1dk8gaqWyJCYgvky6/xTmToxkmI1m9ZuzTWob
0GJMkKOdmy7nUzVQtwcFpDkuu7mTUxePjTIBXzOP+K3FfzMbbVATWFvPs1/E9RECGUdwHraNtx2W
L50xsoqM/Nqh+QPtn+K4xQtyjZRqisiu9X1VIN2AHQvhykiMQiSGlZoYYwhkCI5fnP2yHIg0fEDc
LiWeolmjsQWT9vjJfa71j7l2u/EV9FGhxr2GEBiRZS18/ZHLU8Ry35IFaUQ4Q0+sD4kIqYxswyf/
4s1a0tMRBkL5tClzX8Asiyhcgu+eWgO9iE5PlA4TTxuoZ9OS1+mj8j3FDB4RaBQWOwF7SCdzgMur
ofqdK7wOa54IpwAvUkkqQq4hqPuIPPum1mYdIpusk49MPzkAdhvP5CPeW+pOQ09wnWKQhvkwOIdN
2Ml3Ax3QAn5XQhrnVVP7tsJMLd9UKyLUp76wea7xXn7ob0G+hY31OEcdaL57m1KJPdyfiUHL5K3D
gnCofnattLmB8U0i3Rx8UAXYXAnSGE0f6sZR3WWrcz1NgrT8SGsOzHUbgv0Hc57Bb/cMWBcnW+pq
gYOebnt3CMXDlUhgZ5+skqM/YiubY6xELpI3tbs4C/PRCY267+Y/sNIQgPa60ltgOloNWaY4ccfL
aoiErswhEU6pAM6Pd58qrFjohndJ3dYlBSaN571ud1cCAYaf6dZyYiDwOoNXTfOXCsm1wUINWg/h
fvErCmm2/557cRY5+ivdBvP7yyUNbqoFCTPmmBC+KasGHKizQwKlp2P7f0F6OmL7QDS2e7b/Xe0a
cPEiYhLdX7tXwzZsahCKl39mI6NcocnfrH6sFMXG42f0PWraqgRwgYwXjac/i8y48E9EOIQw71Hr
46sRQpt6GBFzlmMqj1DDYhVLBQZ3vYmPUHzVehrotpzggsoF7ghC5d6495XspenJ8tXtj36hv3+t
sNYvsql8QZ3UTwZJKaCLpGxc2R+XrzNcSXQDZZcgAGwM/8cNLKzqpbLN2ULRky3qd3uc+Lq7ji7S
3OSvTPy+di9uKnt7vn3Q5v2tkahizg/Authdpr4FztVlaXsKO1565gqNn86xmK8p81giaSpKQmuQ
Ywl62KYrS41Y3r9SYTNNafOcAqAKe04SVaLk6aqWes7ioi3hY77s79EuY7uNydpvxqO+/yZXYdEp
6OiT7f83EkEmQj4WjEBhyVCwuYjs516o9NzWeF7guGg9Ti+WQrkW2kje1pWvYGniZrY0OxIDcHIk
/sO+inS64nFNrfRMwsf/oxrRua6Gnc1iWQ5KInwfRFSLyT/VqsatvbIOL1oxzB8pBnrOb2j1fQQy
B9n1aBY2U8PuMVdEntqW3b5638g1BNJkKbNWqKxss03rNcrWPdop3KSErwTUHNyKt2Vt8I4K9Sek
+ck5hMjEQOn2utxXFER5TbcYot82B6VVdyRhZUo/HxhZXLlr3NAnV8w1jVzqQVM+0MRSCoCzdl9y
sj+qdbkhOuUi4MHouc6FLqPkKFWkyDdHLIfN6YItxAg8CQzd5ZvALcVfLdo8qUsqz5CjGKoli9rB
vGY6BRbL6znDcZnoRWchQOXDd/4Zb5+C8AWc/Fq26m6Npo3pBwcBW3Jr7nqppgupAcZBwRHsjTaL
LTg2jd5sYKLsRwBRbGTeMjVJMMgXsgtstbUTt4GveSd4m4hjusqzmGHGTCbwg4UMpHLBBTys0DwM
MCueZw/6VXoJIdtpsKYAq+8iu2ZvJeulKnhm30u31QGxH7J/Z7fjUQ26brSlZNq1XWMawi16DHs7
sir30t/KSRhe7J8Dgpwsuuv8Gn1xqPc0HhawJULoHso6jpe3tRXXkVpLvz1Z/cpIczI3fzwFWwlU
5BiLJr7/5kmjqKidX4+OnxVPAdcEWC5HP+6PGAomVATayy+ZA7VfKFdB6CRNGQOs8y7iqvf/we9f
PvtTrbE8M/6/RZeUUswv7K7hql2E5HPPQDnqBY1qJYVEL/10pOnXf0vHinYdktqYXYJlKkPz6Cgd
u+IR6bZbixywy5kyQtkTpGIbrGiJgY9PobZ7OaKWI7pmVswZ9l3SZRmBxpEfT8T2ptJSXm1GE6Ko
bMjkpUADnbaMet9EYLnfcDzqcFkU7L74r43PKjc7qUTEqmoJzYviEUtZCwZx6nbDcghXX0qK4Znx
ASpu8Zs33vxAiiyTcYYU2bwL7njb0RIXYiwbONP0A5TmWgv7+bqBO3A559L/CeCLtkyoiHM5ZGaf
FzcJ4X7j4ojJEqgr9tWi4akpfW7jdCEhbH06COhW/nz4G25Di6+XRe8Qle1m0F3is/Y8At9Lx8Ld
m2QKtBKYs1FJM37q8Ckh+CUsXPhi7Ll/ruWosvxuVr437ZOl9vS7odlW0KeyYFf9xlDhVo5z7sAL
r7DsV+MuTLHguMsA8bU8t2xToCYdoZNYc03+BPf0AQ2aQ5Mgr3y+DtPKin+RZud9rt9hhh4C9Yta
wZ4ggbVZfZm4j1iIy5R1femluaHlBHf+kwzi5LGvMrjvDlfx/vKCxn9lS/yo+MYyPzo0wFaqAxPm
HMeWoDsYsPNn/nZM8QmaE3By/neR5bNApWgSCD7vZco9wG/pvS78Pe6CU0aGeFRfPNdQrr2oiZHt
DjYh7p0nMkakyu0xjl1M5+973hsuHWyvJDoOf3AMnho0hPzHQsXQ/4L2cuoylB0STRjlZKZxz6aa
sgjrSiZq4UISKPJ077jWGkNpB1udv3KDDKx+YhSkOcWsWVyU3SoMiJsTDbheRSlF5Fi7SvZ8McE7
A4gOyoZ+xT0nbPdLXBCMngP5tDb92MDwO0rNyQPjX6Y42mOrP8PrzKHEZ97Az6hBXGKN30w4QAIX
P/6Mfutoo3FVbAAUjCjjT5ZOvgHYXlw5b83K8yzozlpZ3oatL0t2z2j6W17vzlKJRMzoQ8EGihBB
hZv55UyT4sm41ccb+mPUmx0z2M/6F4Nw5LmYBl779LkBucC5Ef/pRYB1KZ+tkKzTjIwFpG9uzq8F
aKMtCKmJXm1oA+gDnI9q9iSWsaq859MgMdMxiALkNNgXf/8QkkV1HjPQMIHGyuqgQvhfO6Mu/7SB
c17ZiO9XGHvB4/GlVo4mvw4Kx+USvG7JM9PYECa3LSxyuU1+xMU2Hltlh9lLCWB/Ap464t+TYhxd
yJqbEDpouzkdSBq3H6bbn9vv+VhjUtcIELWlJ8/Boyb5LJc+qMzo0i8J38cyMJGgZy2RN43OV4LR
eLfjCdAz+xKKCdbnQAudirpp34bjWy9XBBtDw+qU7GSE/xBEugiyjgABqGfbYihUsAhEbiamcYsv
oW8CFPCCY7Vpx+G/2vXo/uI2wdjK9Wh9SdtA8wLW/5YyuT9kfjLwG9aWwbaBIe5O/z53rmJyBMhY
MwHsehMWw8bgjWkQR8nX+RYNmt1CrmqN/9TuJuge+oYe3i9+K1xzYd49V08uPj6MP3ibyHJ34LDs
iwVquVgJw8ChHd05tTEfTkn9p5tVKPkvELqVWJw3wmsEE2ayvkUfDsmBdzq+cyVGfH4/TGL7ytVF
wLfmQQ1g/e2g/5SggxdVlDl3p4CguL9k4mawHgA3GQdHDplEuBQq4R/W4hb4FsNguHwf+uDE9nf4
5jiJV0kCqgcBe2uFInnAFsxWRWdiYwPHZw0L5xb6ieNEtPrev9yKQcKP2hLqxy5k8FmhcoyJlrvf
OC8QrI60BwDjt8r7Tvpq7lrRfJ8HvYfn1ehOIyFcWwa+v+y7yDONogTqbTWQ2jbLinRoZ+a+JLpa
sVjy3S5TA8QcqGmCgz7n8D204eh32mtLmH4ujnuXfNt/XkZlq2SDBCX/AwEPcwbB3h6QyY3aC8sW
32zQG8BBvZCLajgx6Pv+iTvh/u71m1SBIE5V8Gusj+xaHLlkI2GWAzTFMVEWaTWBAl6Svb6kncOu
wzB8M/o/Vblgcad3bXLuszwqpPIFAzZRvSBXsJSYnN8ycym+TYkHCb+HjpZ9Uv5pSp94iWOE37Lm
Wxxn457xF70nJ3MMuvTEDF2bghN97oBgL3sZAmw1UMAnwg9FOXw8qgenOHqGZcYTeBUztbJmgD09
PdAmI6Z519M7VMKujarQkm2vI2vC2I1mWIq8T3Uqp3WqyQx4a8xLUogpzqQc89YTwbmwT7rGPUsQ
wzuiQuhrLZ23E5+PF/9n++iO/F35HRcl165VsApyCTWoLPep1f4BrtHMzjRfPOUcXdsKyv2Htuyx
E7Lqg14VW4lK5DxcpNHf2W6OndjU8E4mRXRkyFNesEXluUpVZinnzKb4lgDzhl2TxUl7Y1ocbjRt
IlCXyDT9iF+3/fFWkFuQXzZ2EscZagsEW5m7ikyvdK400lTqD13u5HWw5s5bVVWXj+DAFKA0vi5+
O/DMwtXU2UE1DVJmYtWg4uaTkL7RrAuMj5xwbcPLw5CdBlo67lGfO1X1iisuLN7jkBKmRbILvnk4
fjwVJ7PZDjyneq4Mazk4tXQUsNVjaSAQ81aQI/A7jgJkkSWxHo9fHt/cSW74iDaJiDZWWzx/E8a6
iKAhsx9KTOOiHygJYLI3qHFGDkluZMT1O3mdYRNbO44JOIDrVXahRjnG+6yPtomts+8HzY8JLHy/
i8qHpDqSRoAqxjG1Vcq/UiFSSug820u2u+5ObiD1Mygeu9mTK9HpCLfr6YsWXys5jYhth49TKtCF
yBdLHLwF48j1Oean/4fvJ9YPjy/Cqlz6d08bIDMy3EAfDBf4vWzBZotno73DTjFlC2+NMZZrSTPH
WRRQwomXZ3M8C8EOjyDc1z3qz90bY4/VQ3naYkzv1salorThSEm3sFDDiDNE5+Ckeu7wHSsjcQZi
RxWjx98bidsP99yKacZP4qbleDlXTLaP6YH+2/kPuODweqcrhcqkEZzhz8hA8emtu8GZtLD88YCu
rdy3R3PaukAIRJnH3NzcPVyG84Ea9pHDYhBG+tZ2eJfgdGyLzyoemxwf91HOy5bSjacee6wtZLSZ
eL9ACwQv14qgDObT6X4q6HmkgfAoCcZ8WjOw7SopfFwGIf9Y0BIUSUnMZPc0bJgE+sRjhrmDsFth
dgsiA6KaCOq/l1s/deLy1XKwWoI/19wVW/HXuD8FLyFJb37vq8vQmHQUioUy63heFVwRrkK4uy9+
bG20MprS2iSJb6C3Nb/7MjNh5l/j2VX1276KciliABTUAiXai0Vo9JnDAEAof9abCBjpPQKgmdl3
98LMxVEIMV3vJwt6GHVzT7OrVZUvAPDurisyNM979SwS5/8+CoUSqySeQKI2PKuLSG4LxYWiMa/e
oUrx7oAn3FgLIFPnQFoO/SOaxZEx4NxkVIq5D1+ziR7KVhYJgSSIeTEkct5Ezx+fjp+2+y3r3o44
05preVVryCqFWhhrQ5/pIqMk+msRNvjQx6sfR62hZQtPQdE46hwkyI5dsAy6f4Mp4TlGQfQ4KRPr
ZNxdsPbHSdAKrhEKtPZT5MEW5+R+qqQ69kPfB5otCFhjdhTM91FpBI5n6t2zrQPdnggW0BXHedM5
2Grs0hrzsoS6rYExSB2uApEQ2+ZvYX6VHGGZO9Ch3/PC4bf+mkrTNEiDfw5fBNnJV+CSwTCXdHW3
oQ4ZdW9js5kzNKTPZrXxqs9drPd2sYac9u5Gq1TkyLkZl1DHyEwJj/RW6Ii6sUAmer44qEl+/mGa
FIk4sSxDdvUx4ovmmhhUMZYME1DUpmt8f7HMP5wNbWLigxvFnN+uYhRaGfta2CzJf+lUa0meRh7j
2ojAloBn4iy44hy7Qa4lqurlwlHk6s4ygx365ieXWwiaBGVznPQ1K9ZgMPgtY56nxvbdB3UwFqsD
ANiQ2++LFoYShVy8SQjO/HkyMEwhYAUkRlpfaeKq0GXm6+l7od5V4E3OI2Px9CGyzybpUvEodKz4
gLxJnsOt3OZulIqvkkYzAiBQgD232pQBkrkHHUccFtts1iakvSU8k6u3gAT+d71yAnm6Ih7BnPQc
qw8jtmucGRM9XcMSs2/W2GNRSecPj+mEhJ/4lwWyI0TLF3SJXX2Kuqp1YDTbeGqgxV0Lwgr4Fjdo
U18k0hEWFllj/5PFJ8ZSLXUq/w2+Ylzi/OeK++p5xQ8yZbW/kpZ4Dm26ghDZlX53lyYekAN+EGil
AUnAliblmpWNivWgS7zpfqKr5kVSzfm9FV6yd5kvb4xt60vQzPCmqFXaAFiY6kX+9VYO5upKM00g
iH7DuUT2hWtkir4lrTtVn6b5accBWXeWaUABGrFCE4ph8z2qwbZ+BWFAsQlpQnqBlZimJmketcuW
GvrBgv7wRBx3P8gWIJIHsqf9u1SlberlZSfVwhWgmlJTwEm4Jl9gdMzg/njD+W+ElLzkHLfKsDiU
evCuVB9lLsvwOo5eDroZp9QnWAXn0bFsZ+3gAgMEGFoPqJBqDp5ehmjcpzFdodthPf5YRkwQclD2
l0lnVjkjpxVaWE25luKgv15G45sTXr1oloSbSXmVfIuegsx8blhbmQwVzSYfFiqFnKC7/V9gsB2s
k7lAkAaq2q4fHXrAUUAwiNkeeTjWxk1hWJqgoMVh+VaSLDcWmLcActJIItkR9jEzsqyJhqTa2cNX
JlfGS+cZm1ni05ssYSPQLFlgALu3qOIm4uNWI7Wmnuqly+luhOLmT1UTcndfVYlhfzpqCGiBAPGL
Ec0sRUnhW+2BFsVk/xiXNugmYiT8CaBqasf2WeQI3EArMtn26/7xhiC4EsAkS+kY21oOCeF8H8xX
yYyf6qyCpzc6Mb5HIyFj3+kI/jiGQA5/Tf957EhUqjyAWP19FjQ8xxaVyJV/aAb4XTz8kfSXJ8Rh
B4wfdTNPLTs2Dxx9l2V34b2tacQBFG/VgBQkp4S8g1Ni+DIrqRh8SRALIeMMdmVRlMMlczi+aBsv
ftTpNiQStkqw2zuNr1E+G6GNkBSqjWANAvXr+lsxr4zlNbJfdT9oCe4ywxgcJiVBAJh6L7n60yhz
XObAIQmdUcJOTy3q6p+IABIOiCoaH8ZzqFqrWrhpqBesdZm2bSnOiodO5xXiAnus4iDIiulbdLlq
uriJu9cGlctUsbFgRUR6Tj87pXZXFouHVRUUu3EEnWxK6ATV5Pb9VrRFAwWz7RLKj6OQaGKR711D
d6/1D4ohPc9/N/PSKpXJtV7PpVjjgMWPbQf75RYTUCJCvxcHeFZiDPNu60sji0nJHNIesMTQvLUr
Np9RZbwEbuaGGXgxX+UWY4Ph+tmhZno3iUHrITeyJj0F5rw8anygtv/z9dfo3l7OOZ2iDTs79bos
5Dl+e6Cn7Rg0ly46h43tinDD2UuaPCKUDOo3BSdbW2Iv3HFilmx7AoS+wUbzvbZpKn0YxZ7H3krC
2wyEhnFXTLn4wRtrM6KJjVQeSwsIOGN/7XWB9iWg+/ddj9DFLj+kbDiTzwEwHMnHN3NVZMO+DlAa
rHt/qTIVQv0FGPQBUqsgb0d2Vii3WazLV/umGjG2+GnRy63X2QeUsHa6jFDFEW1UOH1QJCtJd741
di7h6LaSG3NkRTGen5ztfru4NAwB3xPR+4VTF6FHcZAdRwKEe7W3vAtNSArakXQksonpwqRjo45N
TTUXvgRfa92pqBPZ7C3oP9jXiGCBmLi0sr81nGrZ+OE+gP5LjE3Yc0xRFxRb4Z3bQP7MSdze6ASm
7LJbM+/pk0mfhE2XoGWdI91bx1+MZacaKrQS6bUw9mRHF86WyJ9ayMUT+0mITUe94ZeFGRBz8ilQ
T/7ciEtcCjijZzwDmrcM4in8LEopPErK9z2YckX0S/H4SpIJC3NLOg8t/63KH8Q9qynBXuMDrtnb
I6hkKdi40Sh0qDE1wfuqkZT4a7T9bSXGHQC8nKMU/nl0jlJ5VCRjBbUveR3pnJjtttt41WZ1aRFG
xb8MgjI0K5JpgGx8TNAHzgnlpFVTIykiugUMHCRcs/MuCKpFiOxBrnqycAJhCL9jTu7T4ZUKKUk1
l1OKZdTez6K/WILMWwZSNkgqC/krilOOpv0qu9Y0dTi86gDTaR2qA94pPb5KM6ieeff6L1bmfYfC
oMs4SEItI+okQfEyTowo9nwFwGmRz5FqmNP+gkZRoKs0ox+dl4oaDRFEPeyrPER32LVHwstRysDW
COtybbapd9DOvZJncVvK91PHk2M2OWDp2iZCLzs5Aq6VXkgD8dVYwz/BWG4vMdTwZgZCaz2Qdfrf
D80SU5L67kHaEW51Jrjou1xarqE3i/IPk68Ab5AXXdpEXRGcJ0zA/6quVMdfOnYKnLrI4bpQ6rzC
egfZCUZF1Mnx3Ef09PDeZFx52wBibOzyWf/Nsuc7uiUlFOljN8MrkmBocoJZ8rB0KQHgO+9F8eiq
/SxQDgWBkElDwA++6xrb95WPCArJA8zVvbOZj/bK3iOOPIQZKVOfnZXPb9Q19QjTzFHLuWyC9aU+
J5PoFmx61eY2aAN9noFkT+/fmI8czDBNtM6eHnIHTo6/6ubSHROKaYJb2b6cL6dZfbaMPsCwLHa2
eI7bbFECdylx/6Su+qOHom88mavjH+lMq7909NNEs9hrRniyr4y8fphs/8/bErNWYuz/rAVMzr3a
QKFMHXnjuO8SjHkYjLSwbcHQvvvLe8j1NDITtX6K64+PPLL0N9JOTqFuD3mVYvCI1KhTPEhcprfG
Vwn6Co4e7Gm775la7sjb+fJviXg9WaUte3E2PF8KFeweEhHpFRxi8KIRIx/eZ7m51r+XhGiCRjhZ
4mCNJjoxl4bWP4MR5v5PQD+BIKjHA6XOwROrV3Q5wN3AwCLbREMQ825A9mmMqoJIFR7r4tr5q0rI
emGdZr+6zyjkiDyROV0SbWvSaOljLpcE9A1Nlt1JnaiqG9t6eBEfwJMRrlDNI2RAcB9unHabc04Y
A1qPPctMX8rncdXrSSdqkcB9Xi78xBTFYT9t8D0N4g1N2o5ehrXYrjQdjAQBsYmb9HfIRu1XTJqR
U9w59SOTzT/p3j8pKZBK5LQ2DQaR/VlnnyYqKY2N/1JPULRGcW4amENX3ineAUsTpAAPF43Ibkgm
PVOHXfgEaVd3td+flzr2jkns6wkdHUulMSahihPt7CyrxoStiu2isjJlkbUvx4lnhVdDeBOGvYXh
UzOTwmr8SuutAF6Rl9WEdJTrdakJKsUanQolIrKtxamSOYR92JrjeptP06xn6pI/GFNLHOk7sur7
ITb15PVq0Cb+IOnOyZxnMy7XbYBj++zCA2EGsoktz33WKg+3jvCruSjOFFiP8ifNeLWbAriRAMaE
rvQ25liHygcIoVDxNdQPAz8/txsQjZSL6cMjdhD46I3cUuYCPAuFYQj03mcjEQJfs2HIrNv8N5V8
hi0Cvs4Yr+tq7dmg+eyHE4NJtbTk0usT8xNF6I9hyQL/Zz8biYaRBiGXSA9H7U5GViZAwFiiWaUS
mNZ34+nRTWXUloil70gdHrUcalB4PpGKjwmtB9eOVlo+fH40s5QmAvq9YI6JWeAheK9DPNir0p1l
AAzB8lbBWOrnB6emMEWYLd/SjkxCyzTwDTynVRyoQqi29F76ZUlx+XdON/fDfLJASjM6qd6FSCcM
qtCNOr4QPeNFJygrenJkiL2RNIJV6NriDrU6IlIgVCeycqgU04fL512TiLqeb0ynrTerUSTXrHNI
DhxA82Ovo4vwOUfU3L6mamzXBrfAAhN7C3QblQyY+p9oMk+AKWdsC3kplqmJ0oQE1aOiAAZ/lKkC
Q5Vu0hcGKkqNMEPT2yqXceHJuqSlHQLRU1C8Snl24Qo0Srp280eNZ+T7HeVowuQyJ/989UKOwqs4
kdWhGiN79446bVIrFnr/eFzs0NZrYgKAoStVt5fIFt1lgsPj2EczOByRSLKRbXCwcdhA5sztBkfy
67GKq6C/j8v4Ne3WqrWd5mTfq0ZDorB/eNPNbTbaqNr+9J956m8n35DOsvb5oAOiTGt6UKw73rW3
GlPKNUrM+GBD9Jtb8XP3dNoY4W90pfGD0tUOt93VSi5OuplEWL7QH1kzKT4tev957IQhucsO5MhX
QyoomgVJjXOMDX2+b3OjZ56fBhD3phNIuUuRLzrGHu70dvQXEYlnI8zopthMFMPenAPG+/uO74qb
oNNRuWK4nSUYYbQ88lAAFinGbBQmuHWsZ+ICTGiP/Fj/hOASXJlBekcyz3mkb/gYfQAnFlgWifeG
DtpI3vrdFPSAOftZKg1+WUsnyGYxuxGQvKRNoSvO9SQVUK1stUJWKo06XUm4UWadrGlufTVmL3es
rfvJCeqrWW16lemUJ02TtU0c2hLFZT+PaSTBTf+veiFQOofr9PK8Gyia+DWyONH4qjWnGlBKPCsM
eJd/jxtXZhstZMgU9JInC5bMLYIqze12WFkJYdZHEZHIqHuXX/GMS1J+3j1+tSPcCWQ2kLDksmaD
Neg84McTnsrk4D3/RL9hhxPJwDpJwhQ83nixJs9vfIYqIiyqzAWResuhVMqdpkdLiSP9uuGfUMD+
/nIKoTplcl59mKnnbs3dC8sOtjJYam6DeFWis3lULYtZhhPKqy4vJ+8sUHfSzNewjNXlDtGBu1cK
wml0ueWdNmykin41DHut6s0ZBv3FgI1ypnLB1biSdKFXWT5SzLaU6vKHpZlwPp1BmpJPdxn7/6uc
+mXU6yo0TJfhIP/H7hSR7xGK375P5yi166JPDBy2aCScgndl/aXv/GhzwypkjABGE24hUL5xKt97
ZTgsNhUyFY3XjoAcOUBEhKi/K5BpKMb2+zkptNKZiL1y8X3KEeLWC6GqapVazZjGXgC2OgOoSnJT
5b+W9g/GGaCcgioQzOxv2kklCqdJnPwCiZCnPfboL1PrwXhjQo1sSiEYMWvjO5Hv3AARMN67gRge
J1K/JzXPLywkNx00x6miKyW4R1/0WBGgQuan9dveQvJsMsqXjJuHKE9RMWkqJ6icZalytB0Lml2S
Xvk6jaTgZZF5h3Ttx4YU4YjlCTSNtAV68i0l44ANTLgPKvmCI4TQp4R3OCvaQW7AgNf53dHzMEkq
bVB9u483l/s397et1kWkK+ZYohzBEfntRfoPLhsOOHyLHlVNjYeN1Q/kQnmjcuU0kVf4NhOme6Gr
xVYBfanK7QTUqAITvF4gzHrrbLrAhrixTAx2mNbFA8vIs2nnJUKEa5wcUpKtYmt0eSLhtnocX8H5
bzcVei+jJ+Lb5+W90Hj44s/WKBRASYYN3+WVBcaOGW90gfzA2BEKOLGpgZQC9Da6vjiBQ2sk4qPi
qsGs2xWTggRLUqte0mDHcgI75ZQ2VdeWP7F61WF+mL8ZKFo2q7MBwdnLNtABCGszTqvnapC7QZj/
aUdEtQ1AtG8+KwWnKSEijgRPxbJ01acNbhbDqXbBuJkNSWAFJq5Alor4RCgkq9C8VljnfwbVS+c8
gpYWPEN51D9QDfQ5ZTeADNmjqSsXzoC9BKpSGgvCAtx4Y6jYTpBPYtm7QQhCeSppMX/HwBZucbLc
BSl82LJVO46uf9ru4esRgevV9eZFVlJNKcUcaRz7GZkxQWoTU+HTCWuNzv+Wpd+R+da18nr+OjCK
tRhaWLcs2GsZwJNWX75hWIhNY8gq3h11SlSNPgOrom5ERZfydoPY4db1kmQDsRW6JqtLb91fxHBw
I3HJ75f+plF3syrlembjrxKGIxN2Q2TM7m7+dT532H7ZENsZlSHGEUnnT3geFRkPxHM8t0O6JMYb
p1ohWe1hqTJggato5Xogld+Qk03Wv4qeMyjp/TjGaesbbjedzSgTAOc9rC7qGmwXuaPSVY0pIv9G
fl3MV6nionhXSKKAsNxAQcJRGMANAB2WZUslXrT/GKSERX7I754eMwYZtKWt7u6eE0h9yJvM2uUk
L8sOWr9/JhTBe/I0DJS40vDZwE89fA2uK3xZAKXbjezciIjO5qy0P0UyZVmnDHFPbwKDxWZsb3TP
gKAFbz398OEgvZuq2ns7+Egf4EdX0zYGWzGOa3zHRK2aFLHi3ImvcbajUa3T0kZSzAicMpj1BLkX
ledeCLcLNMT29BJLk99RCRBH0fwTdJgNXCC//9sYut/Wmoltp5NceDfaS3Ahx3uzVrAnShHurEVZ
uuVglm0EHwZzzMQ4GMGWNHQOPMQ+yf7MsM/ZLleJ4Gf0rZtO+7gEqdduNqewoUi11YkFgFSEIN89
MbTmoMklCy3VSK3lblAWrEnQ+hFTobGjQ9f1649nY/hlixYHklkMcQ9hnNzhNr5f/uOLjJdfSEAv
Q3SX07tI8YEXz6IDuBIO1yYD/EnDnhQ3+Pxcw+0aSot+iPRJKqNiOQRlP2zQ/84HlyqQHPkEg/GA
tFOileqJvruo6+yNw8SG/tkiMg6z+70k1ClMrwA92f+/vBv9H6cGxc5e3lVLMv355HM/w9hs5JSt
newEAsEJtTSyV0VBRrKoDXsJy6TNPAf6OoobDZoVByC/Pl9Z8d+OrCbikFhnte21oI2lfH9zlWlb
s9wBJhJB1x8N3clDwhX5/NY1lva3U/lBhsuOkFTPQ60ageChu2XbrlKWbTyUfpZrAy2KpnOF1Amp
qF/QMSV6+4vdlDsrsduj4X1lCHUoGV6WRQFpQh9C8Dch8WZ7vjH9rJ0Ui22lLnRMIXqh8xDMCO3j
p2IIWNvJR1i4zEx2AYDhVn/de0rXV/usiJNMngwuz8byiqm6qR1uFhQYUtp7rQR2UFAYar8IbXjd
rvRH7ivnfWO7Lx9UsrXR90yx7EAgmOma+hvE0YiKKM85JjY9+LG84CQuJzZW8pMVevAudKEDKcGU
a+x7YIuQLPoVH8xLFNFLeiFpj5AGuCS8d3IVwbga2WZjSw9PPLBo73q+PXjPz8IgIa2FyM25bWBS
N2QOGQ/CVHGWZOO0b2ySdM+SCrzRYr/fuALtUiPo5idcFMY2GvRRvE0aXPQa0ds9dfRbzKqYDCe+
uMuUiRsUy6Duf7YacXN9AdzydfJTIktsmnzGiVYGbj/cK7FkIgtPdwwA4hHj+u3BUVPBInIXY3JI
fJKetFtuK4zQq9E3Gb4Nl3y8pTR87wS72SwMaDcijYAJ+TjMPl/QW19mI938yaqsgfqZ5ollQTST
M8aoLHK3gWPYvIclZjDrhXZCGlybLKYm+/MfCl24+l+jDo6vdpFW7oxWTLlU4HvNUXhCqxoXZgkt
FRlVyIRmPgrEqYfAbdnFl5dwikpfWgEPvB86fwq2jUr5GCAPSJXZRVw/1XkJRgCPyLhKOckNjTNI
JzDibNDgI8bCVsWZF+8N+F7y/F13fTjWSEiY6pBj2MVTctA4jJYcHkPTCriBBY0RF5tGd8VehoKy
KbG2Q4X//3QFUU7pbcQ2QgAIa2ks6acMGSrdh4aPHi0ANQrmf1XZc2TSUPuNf5Lc3AmJVu2cWp7e
ur9TriDIckpSrmQw78rySUs9g/6rGzaczdCYAxOXLuYUPYZV7rDRfde4WFWfld/ouJXyVk5uduhR
UM7brb8ULn3GQVuyuB6hNfcDR5+lgnL2HWMk03iOuGLeAXRWcEsVkD4vI2Mi1zLiSxAM9TcdwOL7
we/zwOBm4i5zh6b/TOMK4zpXF0HZLjqF830SkmSKEWOPA2BldlyCF25Vd7rAdWw5QQdGdeLEN3TR
yIuzWBbB+y9/IMtJdYA7kebHhDoKsrln1Luxj60pnkK+/qS30kCo9RpNyUw5HajfYOKdLVHzj9+n
LgGfJzIdt+LGGXE9ynyxQG5y7oqIEvTjM7LQl0S9Xmi1UkB/G5xP06X923ja3mVMXQ6xTA6+x+qD
JFOtkyIAFyWH63nw3hVFA4AAFGR/GjdgkB/XwvIautNW+Dxi0ZwcAN8W7OXroSamxerP7q+HvqwP
RJkkJRV6/ywwbppIYASmZIK7p7yrVCA88BMKLA2hqIIYmYGncJ3uYQrL4Mbk3v2H1I0GEBu+mEAU
s2nZapOA/3Zp4WjE9EMIHGdvGsK3dAo88Q8HDf9jd4UyhKIe1DXWfjtfMX1HroYfHKa39gG28Wyx
Y2j3IMui1ARBNPyjnYI2sT4oNpHAILrzpXa5sHrcz7Unu/vCB51KzQOeYoBFu6Q1oWYxyYqMYfeH
X5R7/8cy0gV9VRrrIJ9mkp6kh95MeiufQDDWfhYxbUccloVPMNfZqOdYnLlSA2/ZzER0ue8239Hu
LGPxwfVOPpqjyJDt56d4cvxD+Nm2lVj8jBge1er4YxkYFOHmmTNwMLJl6wQVVXqqBbKwjqqqq1nw
vdJuznEdbMIe9Q2r4Shb7VzN5/wzpOZzaueOeeOdha1RBh/0/lSPezuZRpFO8seOrX3TuEm57+sA
8lsZuMwY6cEOTntaxUGxUUEO6MkXPH6zlaNOlAcoWdluvrOVPL0lh2j1scS+STHWam4EAf6t/MUx
SIA9t8NZJtBnkrBeHbh+cDAkBIIP5LOsU8PUsE2oNn9UajSxyGdyVzQIaRyUeGanDGPoEK5RBuOM
Ko04jQC33Fk55muC9J+60AxYF3We/Rez9OtwJt56IwiEvB+pIZHho85VD7IFllnjdS7DnJdhwpYi
62V79rfstsWgN8wQakBJF4I1dIJVk48fCs7j8ivp7ucuyG8MYbIX6MKKcpPT+ksMvdeJA7csfmmZ
UpycpN3FS7OnnHDTvnnAuXWlKhVCwJID3CzV6r5nUEztUII7Ks/laQox0JOFzC4RFMb/4WDJrxJw
zlh78UenYbPOwV9Qxnwm0OPcY9Z/EBJqpI8OSxZo2EQqL7dfes7bhiuVO4nKEIlYiNlg2Tsrz9pm
/A9IWLdda6Kp8qMm430hWRgakS72mcjED7jLkT+A+xaShAzolxFrs4QF8sV2WHTKroJMA3zE4a7L
do2jqU1Yq57yjNNBIilry8gSRkgrBGkBO5UbIfZAxxsOCUHjh2BjT7VQnAepEu5CIJQQdgcuUyiO
GFiHXfLEiAarv5E3y1+S1l25jOHjL+RfJfDji1oFj7vIBtcyvRSxDMwKzeSXLTYbGkIT2VtmjqXY
PVbdzZI+MeSUzUNL3Q63acaLvOiM1X3pRHW52vn7tgglAMeLFXCE2MAGQ2EDuCnfrN9B1E6eRwe6
lDJC0dVRWOGJVEMPI2aERin4z2YCovB6COAkVyQ+c6NxPnW8FnKkKidY+HZxXklPilzRB1RkZwQ9
AzjscKD4gkPr46LtJ1LunJVahS90vZGiUOgqAmr6FU1b/RFIC5QtgXQsNNEDp4O05cNSEAzEVHxz
gUp2j+pZpF14vUPGndye3ZrxsRRaKyaQ7n9yTkD4B3MWS9KdpgAfBB1p50MQwtaEzZGenvTSrCfy
n1hWRQYKLq3qlcFawLi5MMm0rNEnJgvAW7nfvqhL3kK47QOVc7bt/KYEIDb2ZRxgOPsvxMt916nC
LR9F4tYJ/1D2tgnj3ow318w5y4MlsuM/cn9MfVZfVNAbI0ZmuNHDzJ9mOAntHLtKCX1KJTWeerV2
o+67bJWuwL1GI2BQJZHvhtesnDRmsfjL5HnUQDbQ73St3faCuCNQK2vtZbO8Nbj7SBlrAaPOuPq0
jDodFQnHvJdY5ZvLNaxK8d3LSThtAkgZ9kE9VkVKwipaM8XJOZfQCG7pTZkLsEb25Xj/LYtOkYWs
CAcW9apSPc5c3GsX4ehQvZvMpLh/8US0UqXZKfUATMZ8l8T2cISxadjqbp/710dONbC/8YhaNIrV
HzhdN+b9GYhctmvC755rpco9qdF+vNd2LvcH2bWkeZ1gSDEW7uZ5Yg/0NkSGO86ZGFgpxrfSSuBB
EJCwB2fQSvcvnWC5CRTLTjTHTlanG74LnRbgYZPrJKetkGpbrK/R4eMEeuQ5Nr10ee9bvRAfijc5
Skd3tcRqWeSELFWKgfWK8nngIyTi0krYxEyT8TUC461dVmBs9Y8HYr1rb66olW6NTqBPf9zeaqJa
SmaTzUrl/73sAZzi0G/u1qSgjl/MWjJy/gjYWPXfrNbVdu8U3+qskssC6EvkxUCr4k2Wn1vgwHWj
Uzst4lg6RIkjZ+IickDs+N/W6k2lQYfPkG6LvASTb7+BoiOad6TOQOf/Yj48INiCTquP9zVckiP2
jZewrtVi73R9+J5IhLoGij/1KBXVl+xuEvbL0hYtVx+TGaDSh92pGxP0gdflNuL102zI7qQwWPiv
vVzTUb/Q8FrCplwD81YohaSJUDURoMR4FzsyqBDx+taUq8c7c8Mxy66pSaJEZt4L3KzpSUYfPpxD
pCMCzwAycFE32FNJQDFpX6QN/jvTPXW90PkyisW/dgTy7rp12OqkkQERkcM7mubSqmvNBeKDlnRI
S1X8JpIa+qucmSuqC6ukrGHqfb69Vs9SrDLr2/EW7RDZc3ySN18Q4Xf1tNWRsknHo150qpnqgYc0
PZODB01y5uGAsVQxaY+EIQLS2fngEn4MjzuT9qHGzledHykt+WGO0Ta18C8LdILnB97ZRT6PgAjl
oo+HGr9aLw8dg81IbT2drW02IK2nw2f2p1inxes8idef90bQCc9K7YywqexVWYSke51iic374PZY
yjtttJ1ZpAZbxKmH8IV56rBWImVw6A0v9aLUq6KkVWlhPQCb8RnlPCkgRWJWC6HNSSPwfBKX0zpq
+B5HqdYa7cOG9HZpGlQZrpIvVpWICsxhPeU87E+29AFdoJME5gIRyvniMEkwoJY/HkwqdVmBlOMu
y2EidM3HHL3DJfnd072hMa2XllNK+tZXrE8G6kU9DNbxO1cQDTAHgloavdiYoYfjuzhZ6Y6EwsFd
s99XoQMBMu1LFo6ZqGrZ2U/mInfWZLlWbRu4n6Ihfgaeszt5B2A+QbMhQeodyx1xbps7Mab2xjPB
DGOlFu6ziRKXs1GHp39v0OV940Oa466ZxQu9d3tS417IJrhazLe8cB61u73A5DyItz+4rbtiaHCH
FeAfLTeWkMqE/5+r/Gg93iY5PPYOFpWOi4ym8l+u8oBi3zjosquW89PoZW3wNxu6VKb+BijBZ/PA
1T3ggw9WtSpJ7DGBlDejsABhBRmtP4t+yWGoY+jNJY/PLxNkwEDDUMGMbX2iJaCV+GFCot+RsE59
8AfhfBE68a/KrGmnWWPW2CrMTOsuuVgn41mtof7q+eBqYF1R49PRA8uKNUKAY2q65KyyeO7H7Lbp
iMinHyuiObvh0P9Fvjx5K3juP/JVmb8qAMSBz8QQkYJ8Fsn9iZqEkCPx7XpFHvZv2huVgGZlWkMb
20sSXoXKVgCO3h14+XC85cormOQWsoKvKf6ziGFdTWHaDdIkK98QQcvnWC1JW9OhNwVNPPdSpvSi
FJ/BM6jmCyqGyaHD4m2wBpuevZ5VIhYlq1yEjjQy+1IhXleQiFMEIl9B2mdfp/BI/ascBcZTYqEz
d+9j4JGUC9bpSHwZBngqSby4xWw5WD+02o+RXqICDHa0yCNZeXmXHa1tBnO8OOYQXBxZvCOlXB5u
wYBP6zjJYl/AvvmqK6+NyKYJ61wuNaTluS0BJ13+HojJPl+ZseMp9P0mXEvyrFhN/2Nvdj8Xs86D
HBfbqqr4zoWqfCS8hO0Jz3ek6g2PGYVNgOy07k6ZSGul34oxJYAKLztN3LIY5P5F+MFySg8TlKKw
kYnv5WSf95ooSn7fGKGpdWPjVfbgTdYE9j+1KusGgwVwpvwK1nHFLq9446klokCSTOtrKYx2RZbf
Yxgejz3ySGv8kAE4rBwmypxQJaT5wWLxSMWKyAQHx3uFNSLsIt7fXrnabt0SbIqjZZ3EvW9rskTO
lxWJGYw3cXq1+6hvuLawSw5YbdOlfwroGOdGOJhdsHmohi8RCD22jBY6z2yaH2XRP57RQV08MMe8
/+oOTu+tVVucYidLkG0gEx36r1GbQRSlKFX/dsPDNMoadEuWJ9wtz0L6Nxpm4zvzdHdL1igiHbbv
x0DOZj9UGZYVSTCyv0DjciGqbrLUWV8Ffd5btP3grggNk/OzZJyTFIY/UR01whpFsAPMMh/IgK3J
1zD265yDVqeSag9hz5a1KLA8+KFyWVQiT8ajrTew8MCn/BTIRsJEbBcKlcWRkQvLJlj82zhmaSS9
mI9KGom6927OZ7kBZL/5WxcNdbsRT4OgKSiV5K4VEfLEmH76md5D1zZ0jGTLs5DiZvYUXNT2lmSe
L77/WHNkXDfKZwJ8uqZ+ELGhUhqn0rXX+4NJszhAmTFdjJ4KUYLeaJKRbU729W0Po7oetk6qGcmX
CWRenuUBigUwS0fyPHBLZ7arnrLX4eH6BVfJ6yCS9yMBOKBdVAitnH2RrZzJ5WKfmllnl+SHHcAR
7gVWBUfrOanZ5XJeTxqnMTrObdY00IRvl6ebQya3kwPUck7GC9EeNaAMYNb7Q5Tizch97yH3MkTd
CkJVoahsW/o7AiOWPb6vJENZXGypcPGCD4jMoQ/NLRHnSH6C7fUE4cAXaWOefvF7NYM16K3mTBYk
vwnrA9tqVpn5ZPT/wHeoD+2UHgVyLkc0Tq/LXENYEU+/fCPfPOf1UNeNHOYw25wGT8Qep7ldWJkZ
2Hg5quEb20pQzmN3DoSkk+Xhs3XnJxfso9+yeqbJQVRMKwGieAuq2CDtNnQsRW+nsXuK1IVB+7R5
vBXCuRdTkDi96lBglZqe5Q8TpgP5tXo+4n9jIz2NyVBoE89iyNAkKPNXNOk4b3VXc3E6ee2wrNL9
dLVhyFN8fiLiXLjfVRzYUgKhdwPC7Fn+R5X+gBGhGkr/ZB6JDMsCgvVIuM0dC82Pe4anV4IkOzOI
aDuSZWGIQiNEumMbPUqplr1A4YLlIwLzcIR007UsT5/8ScuZ69zhnFOOJG52kp1ogDAyz5ORbdr3
P1aze1sm345i6+Blft4uHIryrr/ftifqGgcdl6ElZ8qsQwK+wmHB3J63jKg2TvEwVisdH5IyR0rn
A63vuGhZMi7nHcOxcY1qbWEvHt0TwrRvHsEcXHnuyHqptPftE7ifeGD4s8RsCOv64T099suXvGxk
B7DjWlfgWdgNL0NsC8OqmEivgcPjz95KCrGQqabvDAcY98+qoFexZN4QPVfa+CIqcji4V9UoaTQW
7nE69E+dzfgXTfO34rEjdowDBTBvObT/0GEhNa+Jv0wyGgPGREyGWw/QN0TO+jnUDH2amirlCDLy
YQ1W2g5twqhNiggmFtyhOr0o+aYX4Z2Iq7DV3buCPTLjuE8MjgCquQBCcl+/kKWToj9aTjqgUzgx
V4yaLFGu1IVMBnPhQN81Xq2Z0TDU02SN5gkHre36/f/jeYmwfdhNfzcxhCGoHcdgIhkS2wzgBMnI
wff1OU3HhbhzDSoaTUJmRIpSJHhXJ9A1BzeaPL3kCFacujdNnF22oPe5rgMkvS2ToMh7wdzyQxXj
7aXeOE/ugxJVqkGPzG3eUAdEH4MoTxZn2MqHY2pb/cRXm8IK481Bc74OvmRqODsd+SwjqB+eChFQ
cHrYxkfxWAnFoFqLw5S2vO2EE4eGjjO+D6QPslitYYHQvzmURy3f7/NdvVK+Jpv+W/OC7899m9pr
P6ViH/Z8eRYzCtt/XDkMJhMiBzMGJA7k5fsaa/oB4E3lg5Zt424gU5Gu4OyhkfSrtpECkeeUUWe4
oxfVtwyOxZbqqLRFj644z1aN5kvi/mXjMPFVZ+gZ7e+LMx8ALilXsQtH9TtdRYvglRWNKlx53EMQ
gCFl5WmMInWjUS9v1xaCntlsKU8ujRYb2+/GBJXPN7sYN5BwULayQMdYaKgIv8O2qEpyUdBaCTku
iqB309LJitCwpz77vKJmCJbrdRl3CAjP/BKxpwWwzNQGt1jW8XrVcsjLJzV/0YgGZLp3WPl3seXr
JsIRF9jMeIrztRaWIZXp0ZL8xLU3HDwFlouMF3ahPLUeqgNKklC2kSTuvZpWKvru3gt5dbctUM0x
/iqt7phjOJ/Qt+iY5VJTt7QnWniaa88wiAhZBEa0UQDXbQWJp6m/zKU0oVyE6FIlu0R/4Qxf5bHK
NuS5cB/GPa52/f2/4GYJ5Fl6E6Q9EM8dnJQkn0mJvOdFfu1NLis//gQ3zBXg0hXKQDHx+EblMEkF
smc7uiXfTFkL9Nhgib7+TDIXeJ4yHBwwpLvp8/UeDZ8C+xn5dqkR4U/pWKQAMq52FWCPi1WVibaZ
l8iH77vE0Vo9BKWLqaR35/aGgY8vxNhXw54I6C2RtTo1i1TZbUGJzhEhJ5F4r7hv7YMPTZPm6dZd
1Al6Kyw6/GQrk7mb0q+dReSTKvt8LVu86cQCvMimojAH+gDLgmP4hhzM80TlfjSlCePEpQuOmwFe
ad0tdeGEKycJyUoAGUFzsn0aZ1Cg6vBh3Wtjvfa8XuNEuChGafN/qyJ6z3OAs4P7vDAXNfJenkw2
ztCp5oqQltRHb0aIgUd4bO6D/P9FQe3FWkFi+yAH6BMGwjYrGuVunr9GylupXbuVvdLCWQROb5pf
gYkpMeWpHK3eU48go6cvH5klCL/vz5mBVVCkvIf4SaO7X8uB7Lptp3vuSJdtt3j5mls7r0N1Kz6T
jQq4h18pMvbmQs714jNWxyuTtgdNlJtjZBxruDyLSqL0Et2VVQ3PCdEjjKRROOGe7w9MSLapa+X5
y4Vq3opVu6JVmqpSqlNiu6juH+bcDg5Tna+Set78hUkC5Ttl2pNSDRYs+G4dwdoB0VmgdhksDJIb
q2Mhrx8JlNDTshkoiA/AYxgkeN1Hi7KFHfcArrXxWGlK+a5vG91mZa4h6BrQKwm5mTAiiDTqKXiJ
zBzwiHMamsQTsQtN6JLS6Fo7tnht6qqKpRWAm79RQi9uNUEp1SzRLfqHQnMmntdQbI2pBgig3ndH
oR2ab4s+ucEJpdvpkUaXmREdk5UNvvpxK3l9BUi3y4wFfTe+tsaFNAm3I0kaLM7KO0FVyPONUNMW
+rtRxulzHc3B6ft0gWG8cdnM/d6wwNsAJ+ey8R3/5J0Og+9U381Hex18zIpLoQ0613cCx5MkJUN4
GyW7p7ON5f6aLODSuQOL16DnnTBfbVzhxJiRbkT88AOZhse3Jb483zxEO3R9k3BHcQa1XpqV74Ys
pmhnuRqWsnXMtZrOkOc9e2cIYS6qOTyS71vvQuxNX3TOMEgVqAAlAlEp8W4eMYASHqE4D8kN/4P6
d0BngPQ9nEj/IPVxmdF5bS3dzd/suc7eGQX5EVDBG48xbMwSDhfA+OaFuNW/YGlwFBbpBMWvsmlZ
h1X8+TRC12VDwchzbTUUfNoNiwcLMDYqX6s+jlcaNHJWKGnCuRm6tXvdQFYi6x3JqXzvsyXCJbcM
KBhy+RBxzseppxYZ0QfQ3UH1xj/KqN0RiGlPZG5lYTcXUjwr1/EL0iIGK1TTDLwX4hSDoTUT+Hq+
H7gMr2Aag+wvLqjngU2zxcrHdRzMWDAZ6SfusiRWxeB3wBoSydjeCGN4iFDBHUEC4WfF3TK3DVXa
ysqGuPUSV20EgVy1TGJZObBF51T+W9nkK9lcYMGlOfoyAwbDkZC67YRAnSbaQxWkiMFN/sGCY7wL
O/BFv5iXxjFud+VHCVAc6hoJvbN84XuKFxbq8H4xRWV77sg8scd677NBHLVQdIi/9VUKq2ITootP
X4zRMeOl5X+ojlJxOcydH9C8HWHoZSiOFuuquqBGO/lxXzCAtBlUAC32HoNuwxBOh1pDnOub7Kq/
TXernv4D54VJNf73+4cG1gpTx3SHcSrAUUqnoYjpFuEZRfMpNxfMqKwKlgTL6iePywXQud3LmdIr
a/PwBbEDJPtFc+ZYD3FU4nD2dm/QFruiD+e5th4e+N77K3jULXLq+KG7j6gjeMJaC/vG0NbhdnxC
RdJxkz7OJnIqqATNr3IEfanWRG0BCljQD7cNmyoa8wQyh1CIuopaYnugy6tHdTRm5hiHajqTw0sR
Fq74TozsXRqGfTxcTCdTeEaIEptOaoml/ge/plUbpvIYe5nggb+vtHb+fBZ0VvWBKPOp3VGJ+1aF
FyZm/aTA9eRQNtDzVu1rNwcSLJflPbQb1Tp0gskqbiuGTYwBAFpYPz6v4hWBUWURmN56WMWXPZFI
AlNHBbBLm7MYK0F4zNMSflZZjt/5oMj1OFa+sQHaQUPQ5HW21OmcTUFMBOsMdjSt+HLJZdcuzJpi
mc324XIuRa5/zAI/vLGVMHvo3NOxPTATd9wG2MMMSkH+/xA52YsG4L0jcEn9+KZEq9zJtmGX1ocH
/7JN3VaNXe5g/1yqVWz6rn03WJbaOMntNQCWVd42KJuKiBr4K8Mk7Ix518yeN+2J/7MeTdhPy0h1
EFXYVxg/zy4SlzkzO9MZxgt/vuOwD1i17miX2JqLHtTymIjzHV0dRDItX6ZXzh2gRCVa1CHR2Hik
KqEeQeYICt3BtahRR+z5EXwfTYV15xPvZrT9QbOChLL1LCG1CgtXt+FiZy2wukCG7FTOzEoP7A0V
LIDUHCOKRzp7dIJ7e1mGnKujwaTHygZTT3MpLjo8/09niZi8t1grpdZEGnCl9cMBo6sdo7yKw3VP
EQ87Sm7GBouwTZL3ck0Gl7uI+ABf4Dg3Hz7o1rdj2DpzbFJ2aNUpTUPK++XQAAwJsKPqL9yfZYOq
wXLgRVWe02+gj1QQUVz/Z6T39DwU7eOMaNSSFC/HRHt/3yhpC8EbU36ppChtZtobYxvLlzXrirWn
QxpS6VL6SevWMkrHUjZeDkuqeoqm0vjDUiFOyAiumaixyGhsdUgdQ6ueZEL1j3sHh7UoU1S8iTFI
XJbBAFMg5ifWWoutNtkymw3btZOZgfqADvbbzHjVyyYlRUfOjyLCSxLLAbWufpMSNh+yP2DNphgj
tPq5wwfoaYIqNma2cKTY4tyrjtHTD75u9BiVnUlvjK+oWURI8+0t/hQapddfJNiEYJgVHMBSD4Gw
SGjJwTeOB0StLIZBE401YrQJT+DlP5Ww6cQFkqRwwfBnvLiJFW+EZpv6WDREwj+jHo/nt7hJNFZh
z6PJh9qLwr4hzQvvupL/uIFjjnu6DPnaAbz5S+bauV8Udx9mqlSlz6RzNexEQDeI5/TtzqGeHp/T
ucN0BtkahEBCKB/9PN1VCDoaaNeNKbdToSKiyX4eNK2qAeHa20cshmDIrgEWDLSUI3MKO3v8rpOT
CFAL4GW1wLnj9ysRcF2sXgMDbTb3KvOuGOHalQXu3+u6Z9Un3WQAscp7gUx7mERmZfCWcN7d7EBd
VSQTrjxtPKpVqsQPiJb5iyo4YajWxcEuMVX8r/wpGKJqumlR7edM+nKNrX7ZrbMO9Vwtg8ws2Wa+
Im/b++tg/7Fc3SdQdiHZuWFCpeJ3EsgyUgSptR6Dwdo1FEsaEabQR5bdXBQJDQiPWcvzI8QzxYrY
jlLq1CjWijLz+73HBdssszvJBTwLc7jtnAPTQ2TKgZMVfXpeXX5NCUk/dtQIfMIRlLnlF8gi/2xo
lOzf3hqO2JBlWx45tropAuJBFjUmoQHCrsZygpUIfUl1MiqCl0ezqxEQ0Ye/wQwmnp9PVH8DyLdc
3Ddu4/XdaYDmt5CCyMz1qqU9u+sAB9Lh/fv6eom8e2CS9C2eCMyIhuYobIxMIWjCvAOAvrOPr8rM
z0oLsnliGijka1+cLvDZAaxOxhs8eX4PbmzXVqpi7CR7DOOQDK76vjzWD0kleCPtiz0j3dUu7n7w
6vlTaBdT2Rip7qXr0u9bGyFzECB1vD8rxs3nTriAGRQSjt+dta3gRspqLT7e1Crnwnl/BA0Vp3LN
7vbHBcOHqGzw5LDwXufnk33fBSeBu+Dpl5eo3xowhQrkbrN7Nf+xg3qSJFtsaOwcKmyWPCH5ZnvM
gXVkdbnps5eW0nQJokPM25JZ6iayPASeW1jQUl/Nrcgjeu0D9l0RnNIGLrfs4mDZeX48JdBD9P02
ewnhm385eZvroZqHG7nPDtfbDIReSQZKDj94GU1PGocOS6ieYN+g0KnfanzQuA9p4IQ7+qZhzN4O
mRr/uLgNXO2P+9ktNhl+Y0LDMZHCSLhTeDKJ+PJk+BX+o621R95GQeSmvQxR4JE8xs5uMnf/SIO/
OcSQLcjxpRQ4JcA7ScPiDEM68GGLfrNy768OkGT7MDmWvBjwpF9qTbGrYMwLSK4dH5VLIsEtRof8
SmCHhEo87hhI09L+oK3CWcILmLyhy8srF880cv7PvimnKg9uJVTl+hdjvI7Bt0qjJNLeLgKHfr+K
snE03paTzC8IG1bKPLvfDXtXslyZufgZ6TPTek8ac8oXl6MyPnwDctU6fVOHMwtN2YXrwajUAl4E
skD7HOSctCLY2unMPA2v/XeYh3p+FfXFJgQoRBdck5hkeXIEQV1IswImsMsiU4T74hXRR7bwIGGG
IbZKcJce8qj1Onin0PzjoQwi4B07KO6kS/xoHSeh3J8bE6ovatKVI3R5Pqh3Kc6nQgL7HDTPURky
6JE5zhinYiVq6swIFroSn0NMuGdhWu4RQLNcjqp8xGpuFQyyXPg0UblzMW2qy58UvmXGT1hojBcb
myOa+5mUsu9nxL9s3nXiYOiNVyWG+xDPpOUq9e1FStItv4QTomFtdANPHIoMXXro0nMUnGcoAxNl
BfcNE/CoWwNGNnj/TI60l1U3WsxijURSSJJvWc+T+nTnQ+Q5WYlw2Q67q4NEzv2zcY/kRj1zXtqH
OxrmZBOJLiVPBxlXTmvtfnrP2Ud7LudcUMfwNuUlGPR0ToBgy7IIRQ7DtTXEeUeJSRaVFXy3Kfpc
DYSM4uT1KOF+JB0S7rPQrNtyKWmn/wMlJAmn+Cu9aJ8YsQtUjdSmaACUzR8ahMf/3EIA1iV4gatt
UsrgmMVLFqyljRjFCTKgtYBdtW3fvyfocgUlPUzugPNm/DWOm+3BBot95L6+EWepFuGcf3cmJY6m
yM8tofXW6R+l+FH1BlnmEMI76tpcsyk/Rw2o4n1NhchrSqzLs1pAqhBRDtjgkTszHIjHF4assdlp
iWVTqIqmVGa39ysCGQX5gch2OvKhoCF99aAjC6F+vYjDHh0PH224PhmZWs+eVe8GfNab1iE2m2oa
/mrthNHp71hlr+WgXnEd9cHsuO0BXEQB/YHO7UwQPFJ03NYpZUbboUxJd76oPNqXTCKjcQOWNU8b
BJDuxhOUzIsHPXsKVz5+hMyWf1F9LL4Lty1nWKFl04uOpqEbLaGPrToSmhQIrQnLrhZRQiVcJ//g
J8uPVNpLh+3570+32MnVJP7Dibyx1rYo1QM3PhUioHpwIEQ8RXoZgtgVwtmQutTkBsZturRHjFfs
kgc6Xng12PCdzK+OH2pzCayXeCAo2zM12mRu8rp8sWsjgaexZL50ZnGAcUzlqhaB0bS3UTZGBY46
TX/f3agc5KwxtmhpcZBo6nXvTN5K0BSo2GnfPR4NVjJlhny9pgpdpRbgJxRUGZOte21wn0i8PzSn
CPonqHFSulOpT+MLM7u59WyhhNPv7/+SbcHNCJAM3w5z9RI9TTxYs2LIQ5hSrJXSRP8EBQT+DuDj
tBqd3wtSSnA2CCEZ/lYTrjfaUlsmgwUIxhuQMTYIDG3HgjolOKYpMPxjbYuwk8BKA8xPVoT2Q3kP
u+nW3jfEgYWoafGq5/SyqbxFSLgOPh53D3z1NBIWfwXbr9melEOOI2fvgFEc80KX3ePkCloZYUxz
gOevyX4oeIWVGk8DmiPJQ3DyjQmJJ/+odyPJS5Gjg0XmulQd3GP584egjmdlfaqwfj+G61+LIqKS
BIwkRUT+jR75j5jtgcPd5+btCw/Jc4X8e4dWWUnlMHVtxPwTEHV36GXMeTNKIPGDd6APFekVtdoD
DAM9/ituv9k8ruaE8BcKnMU1eQmVI5qHcKJnCXhnr/mVgzNDs3vWvy8tRwXaUHjw0AeMJgZFj+58
3OrWFzYcXdRjIwbXewytz6FkWZei/zqeQd0obqqsKa0rOm52/8v257oUkm+K+sWZz+Ol3gMF1dVG
dmJiIYLObf9nZXwZrp0zUbfmV4oydrYcSx9ErpLnZR96haAGG7uxwDWyYrC0/XW8yuFELihvEUHv
r7QOXaiwm4++UuOOtN5yGhkNUruWMYANAR4B8GbCZq2z5MtG8loMyXmTT2OKHevzCbK5ZLW4WToT
lkt4TM64uwkjcp6YFGly2MO3qXY816fEFp7JixNjvlFXkBPz8yPJhngyJPDp1mjtRw7Gb9zCfAZb
wZBEnlR7eUlYVV198oClqVbQQUkWDIUEM73qHQ3/Or+cXkMiFSUr0SEf5Jr2DvRHmJo/3pZm0ZDZ
D2241LHfX3cEO5n/j2487InAnXlSNyo0q/NjFlK2EN7XVXAhCHivwVzvn+0dj5L1+PFarsolkayY
Dc8wlvXVCYkONTG9sZK9HtpGQYtrZJwhskJ9W2mV0/vrJSiiiJPRQMF6uldSFXB39kYMXLcSZCl0
99wiafuoXKV/adL9qlCsB839NX9Y3rK2H5/TRm1eag6fGVv6Kpo0Is+VmtVOuvy5/maPYDpVWNlQ
7YEEOxCGDyoR8/N2dlEyti13gd3KOYTneXmfBIeHFcQC19ciGgObD7N/PwysLqSJZwUK1hTOg3U3
aq8MOPkwcMBHmgMzEI0vR4934lMtrBTOHNeNYNCOd3fbNLQQX3ylH1PMzD4+lnkt/4s/8lPy5qxp
Vk5SFGa28IipCH9ZNQs19D/VipznfvP4Qlo7Mm+FDQZdSOwMX2luIEY/vPmqw1u3QPHPZrEwWl20
nslvQVLzWx6X2Tm3UD3zOw6S5Gw9WEXkRmR9NCOA2VXEEvDC5fOXixuplGTOEY7chl/M7a5FggTa
9M3ZB+J5GRPz1vCvDSNbuVH66cRvWicSeQiJYmAZEzcYVSkILdJT9KOsDwIQXY//TXksGBwUvWHk
pq5wFsaoc7hXK2ETL0z2EDg0LTHYKPzNGuWkUZrrkerylW34rhnfYkUpIieLDTLON4ogmfPuacAN
3LUsD46V8AYMsCLeoCQDd/n8ec5D67ZwjvLgpVmDLbEsy/E1nLBFcZ1Od5HLvtYMUWzhf02d73kg
mbPZcKha77smxexpl2soL3EfMPAGryp4wKfRyn09v4oyvm3qW9+TTRytBHFS6Dfqj4CwrR8XiOOk
PVHHyHQfSUhiP+LOZ6voS6KNprJIlGIceYSuXrI2+vColy5zLM9a8ylZpJlEFXnLozoIXnKXASS1
nIyL0s05W+SL6MJ2+Po/i0YhETOKx0UX3ryV+8b0IAoTOKUcP8k59Rifg3d6SdQzk2U7nOTIB/4N
LLzPvZHUQ34Yg7JOhuIiDoMBWf58NzfZQkw1AmRFpoEMwKL6sA/TGcZmgJPiCB+cLwr5UQJZEpdT
w+Z8SoysoOW69tVYSu4SgVu9Vbx11NPyjuaYw+D0qjQqWwqT2+fchZTl9WvvfdVlpG7VUOnbPSNy
5b6wXs0Jilzkthz574Nv6DcQ1tjYzPepDKDVMLRoJ3cZ6ez80svY3qPZ6IIxxDNEbibhDubuZrWk
oJD/SkdoQtqENIyGQ9g2whjv1d8wRfMhTWzEfXZh+9hDenkIbZ0ksHLVNenNtox0O5giqe5zXj3V
RtMR71RFreTQKOOSQerF6FwzQfblNIUn5PHANk+LbjEknYU8pW0d+ElzUHks8odKrwgJl03Sx42t
BL8mRJMXqaIWgOmX7h3tpJqVIKrABcEcyyXu0rWyD0NFiHfgFIBztvSzOJOCc3WY2IAjNPaEIv/5
3NNiFRlSf7/MrnC5I/lIJ0OE1u/YzX10qBkaaKcqiJK2XYgtOGigHyg1p0IQ38mhuLAmz3r7UW25
QAF+Aa7qbowSgGjJLuvaWo1vbAkOyOk2RvSOJqpJP+1wNkU/ai46Ofd6GW6xirbADxWhY0hbcIO+
mYs2qT1FAEro8NNcVULYoR1CFjEc/QdJSWR5+bdB6NBAyiEFRC0GH4LaqSS0Vflm2kteQ0IO9YsB
k2LUvsH6HhVPzXLcTN5dwWcqwtKnf0snN/gQw7oQOPuPHSzW8YG+YM6IIH4KqhR49HU/e7Zs3Y6k
o0hk2icJT8p3cZqPi/S/zuScEn0+QHrogXWBUmFuHX59RrH2dDEe+BUcyJBBVMEF9LtEJkdZLDVb
KtYrEHskZ8sCP/HZhagUKrXuPsQx6HAPkSShmgr0MWV04nSdz9oFTJvwdq8hqivHZxX8osejwm9h
CsBbwp/gOAQybpQlW8kGcJ1T1iFqPLgHROZ391qbMcGpWqnwe4bEJMqfrBwY+4FTIhV1yHWXnRZI
10DxO52EeAzPCmAxWdbo2f+RPTJrAoVXhavM0aADjCo4qBmx7uSW4TzhS5hP7ooJFQpobKuPckRg
w+OlJgld4Ihx6HUWARyJ0aZcbTqLM5ertXVlCEzwlW+D0w2ZmIlQyTJCsBSR8f3n/RUB/cvLR7Ea
SxRyCZdeqwQ0RGl2nGi2f5QfJ5kocooCFRBeLRX5C/A8rSXnduVWBXBnQ9Aq9AUeR907V8QB87yt
9BjKQoNWgG/zx0sSNTxDSxT24N+KAqfDZNN0jdtZyJla5qOpUmPsvUCBu/4xzkw9L+FLgSl4U/aD
z2ZjUvoi3Z/4OO2jOAHbMBrdp6XM6qAho4eRt1vLr3MoZV7D3NEQQO2GfBTFV5B69vtJkRI65cSH
62cFLiRp85kRZEYKYOVa1hI4XUHpfZTkFrNaKEljir3SDuOiQ1QfeOzuCF0F98Swp29KntfaX513
jh3lPTUbl/ngh3REkG+u2c42qu0eu+kx6M3L+CqpvFcr/BlQdYUFvEe4wHRXt/DnAOiKJ/Z0RvaY
PeVNEzVgf+oq2utU4+jFFSJYQYy3h0/keimkbc4YgrpgHO6pC52cTjS/CppWdzfsAVyFJTq3D1KC
1YuH5FCB2Ep2ZJa3s1af5HxcXpHJ+m5QMjcm/vGjSZ7VHtCINTL0LtNi0xnFhDNA1CVv/Daa7fPG
HCo19enF8rk+oGCSQpbvQ0DnpyJtr0e+dVDBV4XpT2Fq921l4qelzbU1IZVAbH7Beg8WQxkbnXfd
8BkRLZmset5FWVwdy9yF/IDNFoSK/r3zGRbPWbUnxb9FKQpN6w+TNKeizoJW4pWwlP93OvF0/E1Y
Jl/4ny7bMstL/6DU5Fwnp6wRbwz9IAaJIqk4ME6I1qEL6JH/lf30DTByjDS3SIeIqsw7INpFta1z
0pq3mHWdcjC380ItVil9vtpnaheN0OQzoo/R16t6U3Z25Vms/DLhEmwUvsuLHfG8vhFd+GL7HR15
kpIVF4YBK9fjXarEdUNKw12Y2SCJDkHHZL4klGLRmjQ471Pmdp1n4HUNHMS4/6cCJ/aZpGzSohOm
iLmy/F+FqelXCn84h0CXGZw9YNSxYhq4bXhhXgocxaQ+PsySbL0Q4KDqs8os/9BiRkTtQR2Md6yQ
efp6r2uaNVon9fmq0XXyu2hf6dG5pdKso2Wdq0WicX+4i++4hNDZ1AoHQNbaasyEl9AeG2GN6AUr
CbIIxdfKgljN6HPCX4VmCgU4yvuACZC1neq4gbngumNKKgyQKqSN/7nd5Cp6Hizr1gu3vVB+VusV
yRegV5pWY2aGL6D23BM7xv2HR1WME4YL6Nzp1Wln93F4YdXV4piyxEIG5WXpiuHVw/pRyq16N3A2
bVaV3Nd897En8lwI+NUvFSXTQCaBG6fayXM3JQwYDbvY6KdzKRA7/hQkb17XT535gzRX+1AvikLV
Z39WzJO/JtMPjFdizx8o+I7SDAALHIJJEfhuhZEt9vB7VWqCeBY4sES+JvVIXxBQF0EOG02S0+n0
JavN/6w7OIV3A/CELIDDq2dgGXOw8uNB1tE48mV4YqeWgNyDct3Qjz4F43KQ98RWYppSxOKAPXYf
FPqpiZpG9xy7CCJeFSv7rdeAgx71fDHy7xJGdE4pNs+KrYqJjHFMCJVxWYeHCL0PRRsBoVJ0dBsI
tBKZvxmdgHBzFFBER58bcr8jzurNt6I6L0Mcnf6q+9sTBDdl25vv1wT2AHcdS81voeHckBfcibU4
4P9D2piZysMJbcfzP1huQ+VQR4DcaK9ji+91RGsOFhpEmeBkeoVpanw1fDJOSrsqhVD79dntJMEu
iQm6Kwm+BaOlj0boiFsHbqQsXpIb2DWPg3C2gVqU7JTGzP7ei2VCgkGVif4jeZSxti/PrHnF5a0w
/Bf0wWhUNY/a8jRm+CxeTn1yXCfYU4fbDOghEfaTtGVdiYZ7aSjTkWLLQ1Y8lRiU16EhTxfJwljD
dzuAWh/+7leM1jIvOnWE0ED1tdQNltnY0FHXaW6psdbvbh21XwW+zbGJgJyden3OyvJpVSBcKgos
JUfPKWinx3Au/djySih6kXIOFzR8q6aFINWdqgebVsQtrRDLMNFyMFQ9mLCubeeuZGXS7Tv0/lbW
Xl8dYBvBl/973ZF9tkwV/FYUsHjmS/k1qKtsVjL36QQ1qxKBoss6ILMs09XZTUIYazETKR7vTxzU
1EDHG8kkEJZ6UxZHMAug9+TL30k1VwYxlmasbtdfFLcDASZ9kjRDQz+OEbhLAqj9g9HajG/GHab8
zP+DspnlUmkjtz6k8ZiR29RghdNRP5/+QQ9BYco9z/4MJln7yGfqV8oU+Y3KRoZhvZZZu2Q8Cfs5
winmrodveVd0exOMs2Aal1K+TE3BeDoK8yD5xWtp+kPnmXfIngPIoYG+ghPsokjctk1nZ9eOim09
eK2pN5SRT/oSKa6B/Y1Qko+wwLNGcu21m2tJyaBEkWqqAVMR8/ZQoM23i32pVq4cmegyqfZrPGGr
NQbNW7T0RFZFfoq3cT6RKnilxfWmONFmA38uNkuQKfonNtaxLO5tN7d+p+ss5rV4EWjA4anE3eL5
vjOjDX5bVHDF+pkvegpRMwuH+mIKZrI3pcRhgtYDXdXmHH4AiFplHbIRZnWyRJTKOL/zL/ialEqk
vYVbyP4eT5ICO0p+S+cRULzoH8vA6V7MJCyxO8cJTh0/oaP+z1nJWBkVkLv5AQNYfmDKfVy3XtAD
RVC63JU1eFZa6B9dhpdw45a48zFsXZlOdgYRzlSqSL5ghTdBmxL8htF5q1VgiY+zepS1tpkX1vqq
pPAnfOGpr9CfS2Hu5v6y8T9VwF77dOWpYAYS5GSfu3c/4j+1SN7Ca9oOXx5S8DrcOl+ASEqcZUl1
DSmNypsHRfUEMPDARFxuERhSuvVarwkfjsBDqLxU3yT3FLxzwPQFeyghVV/OVkKiru3by+Me5DKG
xWx/c/Vn1YJWk1eg0j8YPVI12Wtn6Nw6SBbkLgXvBpwC6G3MYodQck0FmzdA75MKKDZ+XJqaUI3N
JrjqBPoomEMoyBwNAkuuU8oYWuzX1gjYdWi+XPHwl1cZ9CT341mQ4C+WTpAFDeKf6YKcYomb9r0w
TjEnv/bocj0LfKCSl3yARxGfbeCzJjWMBh8PYydam+KbfjoXQwFUWK99HBI9gA5XT7yF+IseZ+W6
51Ae21EA6XeMbQh/pBFyjGbFtPBqKpAOZFLnVKd3FExqr/mgWLqGHQla/cvTe+YQ08a4wmZD/GhQ
UItuZjdeXrbsD2Mgr61X30DOGzmGXOo6aopcw3eYB/cXcNYOQitS+Y1OdrRCwRJW8YfxshIA8JE/
kp57ETrolqPjveZTh8VyPOxaJ2lhY7sxZmb+v2R+VJMqsaKZ9y2qbqLSPVPw3uQvAvXOVxoT7rF2
ypB4yWood1MK6j4ntj6HfkoZQgmwHkC2NcMOoaVS41DVDfuUyCbdXQzq/5Ut9g4zdIDJGCZTB8ml
Le4jqFxdQXQZuRuwn7997L5uRvhMK7BjkaI4QPf1VXW5QVz56lLazhtuzfLoeC+a6cwzFfshnXLZ
9k82JRIKfN+4sYwstrx2PW30UzPEhfdrAbl9ITmLoOTRZymJtKtho2ld3Q2RfdXI3avOOnMkLiLb
F7EGiAFzw3++A5HacU3Cj6X7khgKcbOHTt7nHfsdM1DNVhpmwu+lNiD6MkPq17GrnpP1K8t6BXbu
zFFCzC+99xcBqOE0oe76QePtZVBa3EWN5m0KKXku3ddIl8rpr0ByLZK1H4s212beOmebC+doOOXH
07FQa43FXXDIPh5CAY6JVvvq8cnNGD0yS5ENnUZI4Cth9Br4KbaqqVmA4q/6iSxbpWc6kM9/5TKp
0TFempHZqO1PDoBimCHp2cnWhxLUfJpiFn3BPIjNs5ELSsqDYg1+DxU5/jPNZBfwhqOKZkjfiYqe
EdygdvWrC1Paki1P237ND095mZ3iXdwQwZ00OYonbFxLUHDDcJ+z1Gkej8Lc5rkYEqUyQ66g5FzS
2uZC3T93FqK7Wwf8hPLdKv0B+SjTMOKOpugrjXXv8El4SZS/IlhmSAwM1zlrRMcDsfdpbPY/r6p7
rvpp+fNQ0JETErUXSRqg5gn4YapG11dQVbOdbxiXmoBTdAZcXBoCZghJ29g9rYgNmvL4+Asw6tuc
7zsRVj2/jY+obe/cok/6RrUi+4vkgAbabKhep2tmK6wyBPATMuOH88xImwmx9RbxhcEnYOlhfLgF
3C4+O/QX2BKo3eAWrQicXh8h8HgP+ISPtkEj6JIcdLonv+sbJw4tIputSg0QclHrniGSyjwK3r+7
tdspOUC0jxSOw40c8QlbGfB20vpKYxtiyS/0vxO6G7Pb+6TwgMe4JJ/kpwqkkUagHsJkFhvjVMBL
IJgWapJwn/OCFwbjBqFADqUHbLUQeqKmJdZZE6k91yeU/HYmm+RaxZgGCltkNY0yvXz337p2L9No
X1EfXdCQFgHgfmoGm7O60VMjibTxYxHPB6ZlPknNPbCYaSyuOjxTH6x1iCleVZNYLWP1HcsUMxjR
clG/ycoLMWbMBhi++vi9PtcsfxljpV45WdlCDNi6pKDe2zj0cTYmiejBij+fJpoKg22PAMIcgDmd
xFl3TVN5yiChNK986/vOmBL9PtpBWWyLmSVebqwc6evxBv/elZQNQW18+xaLNZwn0BOOb1NzN9Cd
/RV3OwiLfJh99aEnblwVnpP2+7HM7A6f1sEBxG4/msAmmFBzExhtBv6knPzMwpwlhuGQTvI/cwhM
bLSQmNEKTw6a/w3SHV7KKifipR0PFspsJjlpg3Hr85t8boVaz1yNr8uD5knsRkGdPBpPKpk8i9hB
i/NBcccwxF52in1QsOnOnS6LrHGUaL2p5amaeakTgwuyd7W3ju5+O5m9XN0VIz+tsQ6OXEf1Um2K
CQ3M9NhsrXKEaKa59InEN4wSFQ/h789xnbkQ+yjZ7tKbLpXQ7Cuv645+zUWm0DVWGhjIYntSz86b
COWElHN7vGP/LL6CuXkuuskML9Hk3F44r5m7qoGrSorbbwbosD36m4FweKVOxy8VHd2yafadP0lp
rkLbQFl7fr4C0MF9bAT4FptLs2yB6HjBxj9nicI74EzVogCmv/K9J75KRKqc+aCa+zd7nHyBnx9z
NATHUkgE6Pr1u3QqCbYTZtbW7F2RyPMF3Is1N1C6yWELMZyJyrgB+vfpoS+8QVsZH2TVvsMbtHww
MK9ZygbMjq6JUfT3TR09D0M5xc7EJK7QAyPxOIA7PvPhvmU4zyf6vApEat+FxHkkjaD/qgHeldTa
TLwbdJ4DyyLSq4WZu3CTm4Hyxz7HJREEqamkxyXHPgHAivy1oEOMY+pXYDIlYdNCeI54kQlHO0l1
iRK3NoDR/MfbET9FmoRmJUvwtZWZXsHC5DfwDVlcxq1TUn10XaT9osXPi5iPbQAq4RtYzsYDpai0
Qwnwhm+7S+5tuNZFalLK3ak8kME0iaKX51f6Mo1sT2/NpKQHe1yUvqx1iC2CcSheLXq8s2VGhuJL
N1Zwsxmxft8dU6RaOnkym+iHjc4y2AAHT/N81fIVinv+o0X+Z4++DQF4Z9lh6rjrzjphwM1HJXOS
4WA8A2GDPrX6nCQpc7HqgIOL9b6z3UY00uQfIumqS1jLH/oygqe29o4oOdfcEmtADIOvsqir+OFu
lmlwtzETnmOyYf5F8vokuRBD/TwgCv/vKPWz0pQCcZIM6z2Cw4c2FXLj4xyV34uiiPS93UeEI8Oh
2MnHR8lcX/35FVXly7L7d1tCSygHY3QGTXjR3Io2sbReKttp8D/ZBn3vrQAaWFFrR9zxjq9dGHOQ
idLk35vDDgDaZMC2hmgGuEd1Svhchu3Pkvlc7HpIL0gj0fIDV2bMAu7mjqvpVvoV2CfPznUlU9iO
Nm75m4RJYQYNaRA+9KzILbtkDSpwc+cia7wp52TweCzij0iSV/G/LZ1hEi0VWOiQ047xVk1oDndR
uXtJVxZx5gZLBSbWNJ9fRdd9GZLfuX8awoPgKyZdMWtb2IMZyyurHexLsVxJZF/h4E9wljQj2ute
9UddQYg60XR8NWATcrhlHTTr3WYRi9LDbxEqcQusjPqhJ/617hvCrY2JLysod/ka9GpO3CxenJgG
U5ATeLq8dQnO2q+OHRY49jNe+9Fl0QbsvlaqrM4e4QE+gP+Wsr3ermRLomvVPkWzPieN6//E3gNL
Br/GIw4szKPqkoJgfHe/cPIDxS3COp+o0RH2dy952iiXocp+T2LeGQ36Ziu8thv3RLSQt47hhl6r
67J+UH4oNps53rIRZOGJxdBzTS1T8t32kOdHYEqig+4Kv3p+9oQSqild+LGOxUm9yixGc/0LkFaV
f6tJ4c+qM5jT3y4jQmqzGUc6v25njjJ/3DNFXkM3qXxrbUsTbZ1xNbvODpecfNWiDh/RGE/d+hrq
Uy1pMCcR105sL+bm5zrdhV3i+EKa/6sxx0sMdmwjjGw1r2ISJjYrHBuJX1C9a7f46L1swgcKKZ9F
90zds2dWaRVW+HQHFXQLCwYOMw1BBXQiREDWPMvaJYw5MvzpN6oHVLjLxCqw8GVgkLao+cZYxAxo
Ky/n8KG/69pyEXEvRGLW0bnSzazQfC83LBHomz/BfBbi//9s1NIIaL1+ULiRzZbQcjbDatVnT8+K
Yy44PIrOaWonbySeRKSaKdl30nRfS9poLCiGR8M6Kf4X4YEy3VR8H7RGpwnywnG873rpBpPQV1x7
gD8ymrs/cGBBz90p5D6K+209yBALxPrYmYQmT+IhnsmRnOLIqGcWV6QioHjLYdng4P9JOATIrqk9
WkdOOW7rtrqWL8NLXyVVJllMInMDhTZ5RnDsMskhtHejVmRFJonzrGUp8SbqsJU/N/o6DZxjmNsu
f34VQLAtyB1RKQZ8lDeZfU3rkH0oZtZCP1NIrQoIykTXicdmwZLmgYvGBwOeVa+0WYEMScUbo+Vf
ZGdDAUGmMawJGBysYoH0SeHTQA1+THbS4yqexrZFA/gaI0mGkeLRKurBn39xRgYn4X0YiOJJHzWD
EMIcrkhMWLjXl8rmXoAIRYbBQaVlh29ElByC/di1Qse8lKLWF/UwYwxk/bjEVjlYdYPyVNbeqhll
DROhbcOXUYR0JBxbKVA7Ih54cLR4b/tq+0FVjWoKukPLOwJiAFr0V8hz2HC1CGHO4jNxFTU6xGE4
f4udFvcriW9HK7yebwzPzD/ZupXtmqJewgwrbow8d1RwW0V+xWjZRqKLjcqqe5voXxBMxzbHEEHT
l1DrFKy9/pxgBZYsbIGqOtmuJE2MTYwjaHIsYmk9FB6ovOCBJywhJGDhN8w/pSb4etTbNTQE8FrX
AUZbz3oN3cTMgmM7YiePBlqJMIO69KZ2KHUkSrv1fXu/1Fr2riMV9bnuBSO2HUEQK/WnY0SjwKuD
P8QEFoQs2BeBW9nYK6wUwJGWLjvK9OfmXCg7r/Bu1w7sHDVvGnzrBhr4tDBuyG8uaGWAa/SuJGB0
rPZGc8W5kw3kjSTYR7AdyIXr/o+2x06QCkAaA84PdSlLTlYoEnjq8oYPBxxKY/7YChnv6zA30VD3
y1sOdvFuZinky4T1lOp6TsJ17LACCDYowaBi550ZAUgmr15oUPZhxpOWvHDvsGpBNK1GgOGa+msK
1nEGycEbUQh6A72lk9+FSE08NqvR8GMtcB1WwjTR3I+668whXNldsUF5OkUSPd68PbuaJjKnwXVx
D+ihUJFHA/vLcBaLuJsVN1i/7pWb12Z4j0n5A2tZhOEpu5z50WozGpGkRyYhRemu1OYqqB8CMJ2R
AV8IeOHczvh5iupVzHlExAa92bXO45J2fWi7eA7Prfgk9Mkb8hgnii2fS/1Y245wlXDHz6IBP3Zu
gdHelFKZKBNITLIKgModqLljB2tZjESsJZZQcK3qix+3DMVUpwQy8vvDO8T4I8J3tN+LzIzv6OHX
KZZWC2FfxXibSwdTycE7/jBIigwKhnRdVjZpxyyPEecU4Fna4bLsZ1k6TBUJo9qmgI6DsW1y+1J9
7Wd4pmp6cjiYaQg/K63HoRGxOKlRky5Fy+/Ry7LU90NOxtunO/ivCNPoiBlWN7NoAnI98cneuaQN
Y8XfR9ezG6miCCvkXdVBiwrD7wA0piCBY0yI4iGG4yfXl83UaUs/IbuZaw24rFsOH+TIcFIAjINe
kTLL+5kMHKebfdzbJX3sG3utWPXmUPTNC36rwRW56fJWuKz1BqgkbdNa3mBEx6OahZ2uX8OF0tXA
pKzF6ypoco95R5iQa2HpD7QziXlKu+KqtnZLDJoa8bzOXS3+2tlVKhUKN+kN0romr3FmbyGYxdze
o9rEjhvHN2Qjrgfb+IIpAGSPMXwshW/gpUWoIojA6JyKuek2NFt5y1xpNIm5KcJWV3KXuXhR+ikp
kRTfFue3rTWhEkyHsQDD32Nx6tjrEtIJ8LC2LWUnu4i4vqk8aS5IsJlMFwsjLqCNcsb4GaVMOCww
YfD7gpGSo1IBYRWDt2rA6JlUq8KObt2hbScwcr7YW5HG1vpKQrgN2tJfHKZVMwKPFF6FWOjhdwJH
eVpdoA/6pEQS+u7KmhOD7wPuY2W7je2AKhS+rj/t0QdLhNrLt+U6t+ozHc0EgHhXZcQgOpWFX21U
JL/JzFVf9yGTWNDcIbiPMbQSHtKaaGkx+sz+uiYUNFNppCksPcJO3rasLBAJGwZ/9hlvWShibR2R
M1Z/k6+nwKcVL9lR1JPvyvE4ohGjroYwhh0W3se1MoUDcAVOZSW20/YGnr9Y+bC/Hmr3vbK95KGK
8ZgzgtWS3aUt1lfTsKsMIQz/utMVHIUh4M31Zyl+2t8ld1mG5vLT7MYv1O6werqyssi0Igjs2FFF
nF0AEpIWPSUSCfmfhkapYT/Wk7POM6QZA3gaZ+VxEi/a8KJnLj+R/08PyZo3N7qLZI6yekT2UWHM
Dl+4dwLBWr8Wz8nvhSD7+SP9Q2+7B05Hzh+Omg5zah3kLlrxuTjE7MfPajwR9VI3NA3FasNAxYiS
qMsJ7VrM31eSGl5NKykOWEYbc0dU4kb+u5gNNjA5mdlfuQk8/0xP0qcNs/8nvc+xcWw0RKNZijCb
a/s0PbkdQhRQJHLFnqpsTtEebcacTysc6dSGhMjqIpYUKqB/G1QxwAJe08oTR27QfsJCL+ovflhi
v0ORqDhlGv0SWDjIjWq6+EdRqgAWJOTOmippyVwul2V0zLZoRggDXRMC7gB4JIi2tY7iZBuk0Xgp
T9NWjY7MM97iHL+lqVOS33R0zLH43VDGw7GO2i0uHm8PGIiZ1uhcjX2T83uhgWboPGnQAXbfwq+m
7f3bxonfyXKXQEdtL7qJwNFOYv1huQgQAsM4eZKH5EkeodHn6yv93I5Zb13O2poey3JYquYFC+83
6NM9HYtLnn/1X5PXNl7H1K3oaFBR9cAQjTlgwy39bjC8qJUkwzaubzi/s+3joJhBdcVJ6gCX3is8
GUd3KU2my9ZOHowZAqBxcW2raLNUfAcnMMQKYM4fUkRSbQQnSnQVDndlLqhI1ygDyC3C5Umjcdke
WOmZ/MlpfZs0YZEBsy6cbC0tAqjd8VNCqNZL6te0mJP9GTePAMPB/ikKKK1IGkGvCqAYn3voUBSX
qHCArzli0NWUzO33nRoOcIAMJvYchtv8GtKgSsVHcE7F9q06yZLYHokLfMB+Ydj7Ll+dKOj61OIF
4uR+pCfmvQZp8ZxYrQu/doWtOrRUR24B3QGhIMs4+mesgdR9EvTh6ulaR3Pdd+Z0+Zn0bqezWHss
ZCGyJzrt5B3UR4x+upRCmmeuRklQXPR7S8EBDm8HIP/M8qy4y/q+jXjPHbXASwG5MIbXLcuUSXq8
OtOjSD+TAeiVaCdRvderaxPSflnnqya5JF0OktALpZusbVyqgz5fWWhgGTuvD1WJNltyxR2FucV0
OHg+OWL23VlAcAIXwKqq05p95ODrLtpgD0HmK+z0d0jt5Fi8ryMNYEBjM8d7HoADXrgV7NsU+pS9
lB1dTVfXRKgKbRpzpsIpBjNsxlyjmGEo8lptd3Sl8XnIWZ+X3YlClsx96xwB/ru6xoN6ovNYztON
Wf34ERdUpdU67HUMFDD2jQz6ccPa7sKID6Kg2hskszjnWFzjx3SMW5cpsbn7oemurLzhFnlftIwR
V0rFOKeOgoalYIGH4eUYoBmbu/npTdMQu+H3Qh0PxS07YFrETiF2o4GcMoazYqGJX5wJIi1HLG67
lglXZThOHaxj90UyOB/RVuupj4XhTXihFtU1YRgCaLJfNuzTN1xswzFHVCs0gTmzjT3ULRGyJ8Bz
3D/P2HSKGuDfjGYwGM5gqZqVibDih0o2F9Om6TCcqrDFM0Qf2zOX1SZ76wdPAoqHkXjYq+OZJL7y
01PgJRcjqzSYiv5QucoUyYaLSZ39DigDKF0f98PQpxO8Q16ymGUogmNZW3PPIq4F4uPhsrJWEOLp
9JSD0cTdse5rzr8X/b9OSqybatrNa1EptOPeJFpkZmN0I0Pf/GHogBjyua8TL8xdgfggQ4SPpNZp
Aju4lPsMUlzB5DWQhIrSbIKdLL0wfWKVRqLVNeTFPeW0Rji8QaPcoiVhnfvLqrQJbDWCyAw3bD3C
1OW41v8VoP2cRlqKAHp4HzGQnYjvBnWu7RpGdXRAvlQXQA6ZIsFjag0KoFzoFPbfkzkXwr+WfdZ/
P0PirGcmEM2vDrSywA8Zy1pltbsayaX9dfigQlo0jAhnS7OAYthB8ff85dlVIqdFrqBXd5CsCYUg
+GCdwPNxVe+haVFL0xaESAOERjMjFZcc05HA0xCYaqanHer99KK5tqR3DqWyNLgPvxHcSMIEi8K2
23rwJfsCA/7j/fRe5WwNftlzEV5OMjuq9nwkf7/uXlATtbfsl8ZXEcJauWyZX4doslTMfnwbDzCC
U4nBUFsFdsZkQIHAvW5oi4575VOsWfp27+Fg6jxXhbz5WdYOYDvLPpi4LYnOOIFAxMYXwM3rdgiR
SjLwExfXaXpVE5py5G7ikITIjQ+N0iAlPkqnpZb9jRGfQosg45AZvaLILQhTRXIy6aSmXl7gz6tJ
ar+xFPRopBoU64UTM8cT7/2ow3VF3a39qf/Emai3BhbwNsPa92xVuf9AAeYOSEe+df+VeH2KnzWl
Imjt7h30MXWmXcLvjIeoHA/NRIGxJPrsqrP8aqsCs5NprLebEGupFtEpnREVt5akUj7o0DWuTjxp
UZWcnV+c7nRsIpxY9CuaL0L1FtbvXH/Al5IMpW7zR0TABJjEns1BXep4svMHZs80ofMNgD01rmUX
WcqQ6eTEMts626tpyXe9gOycknibqznReywo+12M81qbsm25hah9oVSpqWnpOMxB35vrZd3xGFub
YhwiXt3FlW+hGSlPwexiFg6PtCLAcr39IAelFQ/1scz1nmY+c9kTzB5lGeBgs+df051wtZp1m/eW
JmkRhKVOEfhjlnp3e64Fv7J1k1h1Wm70b2oFWjuvX0Nnr3xWgy2oCFWwhQnww50+Q4oz//f3X9eL
2LDeOBBagLKx17eBUJH2/2Km/uoYlat6Rg7I5mdWBCqdJm8KvVdRbxtd5xc4HlaJWAmTfDxIz4VU
Trl4l+3DjbjyliYMR4agxpJhtyt7i9s4G2lgiemUHKd9M9YYxDqsp2VznUUuE+cONU5SPGtZ2dAo
tqTSqOy8AVHv2XtuZ3oTSuGh+mliwBZOCSJDRW5u9zzUfOqambAb4WAAewG7W1pVsUR89wAt2gKy
b43RBvk9VyC/xcTBm3k9UmJCAwRiQh3yTYlkoCRhVLIVCbq+XB0IRoS1erSO/Gg0pfjEleO0XmCn
1FiB+coArDGGRoEG5/OpBTNKBqQ28l+f2gdkhA69iMi/NsElMP6Qf/xRa+u/pzoeDVdUU/Sts8E1
yykSOcGRlBznMSxfIITY0W2ccrLOUiEbawoZNw0FA+Zv5LXrStpucCU5dIKZbTNlFvzj1XfkhaPq
dGBcfS3yOTLFrgb1ZCXWwhIQCjBx5uTYkrIBsa1kmYvmVhHT6hOmI4XszUSQ/rQ5hTpNBE2b7XZp
pi9Z+uoh6xbNRKtpA3lxqV0DQyp1HqNKnHYPza23sYhLAZWVd3j2a+wx+75YrjI5pu4/HuNuxSPr
zckpf/DSNxks/udyEiwgDA9P+D9ghx0XuYa+2KrCyMDXDxQLPweUDSnvsvh7OqdHsJsTkQizh3dr
h5IgV6BL8jOny+Z7WiX1t+O/UuOBbuJh95KBFQq+3sPe01Uiljinw77ccMajaI3AoZF337RD6ulL
LNMoG11LijrM1q9xKrJ/RycLsyHYt/SyvVMxpdk6uCAupXXrctjHTbOVRBgT6zE696szko2Er3qa
hjRVv1YpgmfOolnPeq7ZMxyH0vmrTaabt0RC9sPc3eyQ8KGnjp2bVGQrNiI7Y20iVw820GwzpqLq
qeMq5y3LXadI0XSeS+6XSQq1xg8XB2mGKRaFEtHteKeZC4jWn/G8HAMmJTJPRpBPhIERgeg081Ga
/762mG883y05+DcNWBGekh3xezCASzCL9oLCXNo3DvTffViucJIDw8x7a5tWoqNKkuuF7H+o/Lq0
nyRt2kbWriFoJAHhgfCexaCwVtbEUoMs1MROPV/RRfyOmT63+qnmyDO+r3maTq2dwcKLpN8uKs7j
yUnDDVwGWpXvm/OPH0G1LSy6sp3BydH8zPCm9nhrZ6XT8xxRb2Xhiuiip3M2PiDyLA7LVAseoVeP
mQkfSKWsYHiAP0xquK+omPl67VN/UVd7mngvpUZUZqcpy9at/rDhWauEswJUzgExVBczXuX9uwNz
cQw4k+8XPmNE5sQ9eqao7xomiB2j/h0hVJNcwt4g+8ScpDviMO1wrSodRGbN5zx1dChDU536eLxj
CKBFddFI5pkaErK0TZKQYsDuoKf236jEJOiOAg0Az6gQe/CLttfxiK6l+Eg72m7XoBXHKTv5MXeo
L8doRa+HkRmkE8YLE7kVJDY3VuQ498Wh4xxr7HJ03I5nmISW27AkO6haMhaYlzKcayMx5paVjIVA
6fjR9xMxRTYlPFZlq7O8lx3y4lngK8mau2AwSz2/up5xcFHMs8FWQykc9RFSRzbMqZjH5JL2emxb
bJbyEIW9DMQuBnYlHLi1TAztMlr0Q5m67qbHvFd9I73H2ayJu2RJz3hOwRR/zgZYE89yoR20vw+d
7lHV6DnCzmo0OxbklDvcZM5aOw8tX6opIUYJbxL/i58eXDaWA2t9ZmKAcPwvyLXHki/PIo635i1C
hCJouCjVqY3vXMY6f2162HURVN9RcjDYOoKCTdoeEZjc6yQQJTRZr5Irbb28cxUmmHILmdW0gdNM
HBsOTvjq1VQEsKgqoM9NEDvkkH5bwbgVmGAR6xHmSx9wQL8pwMi3DqvN4jS8lth85n8TIHAbZM+8
qYQIk7j+PChx+JQHqTZukZb9Dl/NDdxLL8kHM/D8TBFZpltS11Cxk+l9waogcGaRsig1DhpJXca+
BRwypVXRegVs8+0llYf41WeaevN8FS+q80JkLM1nqnxK1EW03LREhaDBkgPnJIm7FqBFpLNFRdR4
XSOTJGZm0lxLdGs5eKda1JpDR989N1HkQ8QF4BZ06vPkS4sazvBidX7lDKKitjitoc61mIDQlVyh
RRBSYPPtPbavbjC+HaW+jgXZvzTLb3DhKxic0xvQhrcvm73d3/mVRSxufN/+gEbXv8xqVOv5FfOS
KCvquHwWUunT+0/JGXm/UaKSuAN2fIr2vXK/etKNSvLH8dh2YuCyGncWg6OxXHhOnKHaRX8i8iVo
J/Txo4J6uNVzzMHerto9jBrAV7xbTlU7GN7bLS897XDBdET/OZn4vTn6AAaWZQUD1m6+DphUdgAP
20/xY0u8Ui96134F53mBzrD7QqPPX2CxuRlD7XryQjAmW9K05uj2oGnUQ/l+ZZ1SBTWuokYRBms5
DqRL2oAy+NrGMncW8rix95puvluBWlkkSdOnJh+lISqlIDCJILCXZOmZCP3pKWDuv82gXZju3tMj
zOia/1uBxaM8SnzePGOse2AA19PayhkLr6UMAzU9+ZXsFqH9zOHJW4pQQzGh3kFmV3VherNs5jZl
qEdzKe7qcRTyKW03cfgm9AIK1mwvWU+U+aqBNDos/Me+mHOzAzOZhExzCNHMkRlTOMQcfpk04org
VQKKfc+P5sexGsNkIzs7+Tx5RvEGyY19y79beUGEgVrGXu69n4IMsGD/xSdwtQXZHy0plRrXSEL6
IQcp1G2Ga09wyqRR3VGSMEhkH5eSFHe8ge0YlrW50vZB2Qps/SxxJ15tDn3r9lJYzSQPCn5yt+iQ
EXk8E5hgQwTn7FM8/WARR8LNt/NOligS3Xdz3liyky5flp8HH/jyh8PNTcNcqUaJcXcWKQqbP7Yo
j7yaHhsCh4XAB1kqKJ1CIlrUaSWgrslsxGkf3SIP0EIz2I3916X6VdaqjLDWzCdPGYaW37mIZVvZ
k4pAfAPPF58/uscG5NOrjxQQi74UKTz0VHyzBvzgmV3PmHctdjnYb0wKOp2HpC9wUiDG1186ZB2r
xJmod3YMdQM8OtO58wTnzJaA3lGcmr+2U/F3V7Dkg2YOI7ix4JcJR7USf4VNDwPRX6bxGNoe4A9R
JNCRfhP7DAl8BeH09ps6tOz2UnIy7JBX08KH19zEp9NuiTbFZpy/M7oaDS9iVWYIBM6MgKkulCVc
IJS9sGVyxIjedESoY2oN+9svCmG4MwySznO7aK8cwFBzwuH8xZmKFlg8rKiqJyk4tPHS9lB7kBdR
e4iRlQjSW3UTNb7kCBHvXDqzLQDLvSbNg6RvJZGJdLujmi2rooiDHh6+mfMPCmYfMXAPQNMgT1es
YHMO4ZNIdTHZuONhmlwORFBCj8HFim6xYMvj/MPjmisJwbZfZAx9XDXweq1S+jkIYR/DyVhJoooV
UcDQwcKld3YE8EDV/Ws3wfxtIrpGc7JSJLOV6xau4J8Q4kMG/4gzzbiCelV3J88SNfa2Xrd+Ro1Z
kVfY+TMTsqr8Ud0jCiw+4VRHd3CZ7ewvhUJRHSxBG38eLO4FF1+5Z7iDEQ47fSbc10TQgkOuNKJU
ftUsHxlmjPZ/VQnCumC6VAltgP6JKgPQD1ayz9dSdxTOQT0q8Z7jF4zNmd0JGiOYkTKDFgpepFqG
xGkbPRZ5ZUv7+gMhKbF0/kgQzBawHgZL9BjtBBp+1d7p7AW2K7DLwu9yvA8Z8ir63fmS5riLLLWB
5PldT02fh8bmSlE2+PpkXziPicWw726G64NntwPA3EIYscvkY7bed1zrSNMsKwTnZ+Lzb6LWdHHg
qzfyBarzGpVJ9XtepHmpoT3yyEv+MnCQ6ByufsbFc12vX219LjTxS7WtKinRYrDV6YsQdVD/lA9S
FYlv6zAGu+9ncy89uwytsffdSPeYne+yaejsP8yA7+c43spUKzcs5/GeGSVpSzzug16l1eb84YRf
pdYqXgg6MuL7K7geAbgGfVrTNmaC3voDjgRuDH3FCJ3pzf/aGHfAe87CH9TIoDYTZbQ4ZuR+/vUC
VODvELhfOMSx37PZDGbxir+3g95bhxQn3FvlUKTgr95xcF3tc2pBpuRlOBSqVQjc1GKEcW5nUrgR
C3Oiu+NMo8b3tCPibG2nDUfjeUrKugeyNIhYQqCH+WDIuGzIP1VG1yjuxZdib8Stk+s6b+aVbl1X
/A4BwLIFvH1IzR+iAe1H9wC/iixU4DnSDA+mRu904ZevKt9TwdiAe0wRIvWe4za0FtXGGdeaW2Py
dANphoDWGT/7Xgw4pHMB5r4KEveUzg9skLcYGyVOJ7hNPL20Z1k9cE4cZEDsUOJtUmImrF+V9gCn
7644+1YYNhajO5uOXCqTzUQCQF1gXQatelqhYHymVEC6nUczrwGgrqJdl5PuDqznbfgDz8TWLGH0
MH6AdEBcodmDCPHB2140B9YnpYaX+D5Fz20xXszGpOfOJTp9jpUM0JMpxA2cvNLRzohOZyihlFRv
oF5xy5BuyPkWbrpM1mLHOlFyNtRUUq4SUFuYbLwh87E7vVT+24OsU0prn29QL09hY+/mqPN+ahxN
LVT3vFBV8dwcgZgohHdHfY3Cy+VaCFzm19JIcBPvz5ixgs1AIViU88KA6A6GNet4InXcinDxF2+S
00ZIL40RCpbB+LaJt2tfqNPdw5+ykwXX/JV2Oc5xKaoNz3bDuxr8wI8FDpdPGfpRfoDchzb4sDqF
6m0AP+DQt3iU7rwUjUYAMAwkcFFrX3CvlfrMeWB0h4fV+u9Z3yg9mYECHS3dBPzeAmCQXaimvpn4
//lmID8EB4Cy1i9/raVsLIBQUOj6RHZwr5riUTKGC+g5P7SyZoAT0ojuJBcWkak2Nv25eJ6WBIJH
5PJfJ/mw54oV4HTYTHOYdhF2nNA2xXnsnqRoMbEWSX/U8hpIb3JNDFQm6BYQpzyC8HyJI4iXF/BE
GmCfLWshOTHEMSGr9ZUgq8x4Vt95h3Ze4T8IvL8xrlrdB+SbpXK1sRit2WsgwlhsNyrOPYJOvmzi
WqAOQpFlzAPSbwcLIP+yIfeo7U/twZDEt9GSNRpEOb7B41yYe+uhQJa5F3L7avOPvKXDgzfOVT0u
wRMULVP4EqXN/AaBZlVx2qqcxm83Tx6r0ugn8TxdajomDGe3rhP1jeS+Q1a29NbWwVqP3tAocFm1
Dyat/SHAfXrQPPiPa9kj9MHbwD5VVpn4mtgcyZJoMY+JqXacti9TCZsoZpSzBAehyETyRzm2fJ6J
MPY9zjsNAB3XOBjxgGIjVa92syOGL1IOg/RBA+Gb/lyPH5YKMVh0MFI1HkGntTTnkuvD6blKXmos
/ql7awOnqKgHKHSmiAfVItDB1wGUzReQ2/nrXlW0uFzCGPTbc+ClX2IY0+M6yKPWx+OoSAEQRsh1
AS6nK+jKc10LYca99ou8QY3pvMFpLYVyo+VliQiHlMeW1053wJPS5uXrpHoWOWyxz68b4Kx5G87L
6+SRV8RWZneLU1C4lI5YOx3trySynLSlN3kQiZlYSMMKq6IuuW+lytbeGOlvwGntGP86nZK83WP8
JcZ30Y7EhyakrTeYrWLExNeREAQDLGPrMDf2zBgZDnC8ECaM6iExEAQHjAp++7OF6cnTbFtJDJss
79N8ERSIqMX3y7+/yNJdwIHdvXOLq+c6y8YWEA22rgznayh7C9jqbxGKi4wqfNjkUoKjOUdXzcS/
CqlYUbKhb73+hKc+vXbi6bLhHyIkvc/+0xeTOAXAldyQU6kNoUEC5lmQBfiK5DJzsg+IVU4T1FOW
5QOot2VSXKu/yQ/X8aynh7NTW4d1zwxf+vJR7lvU3GYPZtjf+WKMcQpZcKWKscijsZEZPgbvQDxt
gwouBumsQacaYvNVQEFio2Mfl3Mc6IrY6BwRyerVbISHpLA1RFsTvBE6aRGZytSKqhDvpgsaSJhD
PvX8g3ynNoKzEAF4PNQzvkG7a2dxXe3TzTshwtOx2gpkb2NLCNMK7xrAAnT/6uBWR7OZxiK3pXnU
hAK7lT6c4HZ1XLzDq50ub7iQaUTatPQPJfoZ9YsHaPKLEhO5MGqS/vDBb9uzf55YTWRyIyIVS1aU
3e8uaTSKYepqk4+4hTNIqeid4xPMNi3hu2EqQSO/4LnYHxB1ewYzYBtfm6nOcJTYlqTxR8xdk/Ae
iVlL0PeQ1M26xExvg+JGWa1DcnFbRyggPFWGSw6+mXbIrzf01YfYOXeN+Q++pcfltXpOEDs8uSDz
VY0rUdT+PiLymOmr09fXK/kqi6dk7NBLkk+H3xtnAAcbR9zmvavwJTvYvh8Hdu0w8nUQ/GQfnT27
PQXlTqXg6DFVJolJCBnbYQhf6SvLgVOS0Hud27aEqQRWCsSII7C7QF1nqpymw73rynvo4SYORknJ
ABrYj360ksyNGnbWDoYmNJbhdiy4FI/9nvvynBn3WZKCPOW/PdKksrbFP74y9h79Oun2wyeKI/BP
qADKL2ng01sB07qvAUb/B04neR/5vPjZl8EWpCnqmYp2HKQNY7590LHMBSpJh0jrMSUX+HXIglWm
rZHYsBNsBFDlUfESuRmjroAAmbqQmTLMEPzWIs9mx+okXhOucgXnV0m7oi8DGNHISKyJh5GaTJzW
lVuKaTxhGy+hx1koq8UF2oRHiuNNFhpHOJ1cHjcRHnQjsVr7MrBfVuHnxRh5jMCTreKklAty3srJ
4PP7vau5rgxdurfyMS7tX2sj4+4mfkLfr2aLBHymucXxC6XofL4rTZUBt3rkFf6zqufm8CZcBM4B
e8V6k65TF1yMYPI+1G/nnflmoJV0dlAbDwUUo9w+edVAHFe9MpGZQo1dG5QGM4fqgTJ5gU3lRDND
bQOds88+TxnvjiBkOx1CrQ6hnT4ff0WNcnN+svpywZyX9sk3xftlDOyLfRwUsx0QMBbwxVEK0KPO
RSq54Ic6Mk5Gp1BMm85u+9D3JJ0HfQu+efYTQgvF+uyX66xiSah5xbk9s0K9SF9Gd1V4RWUZ58Lx
CIfS3Vl983lI9dE+WlJ8D0jAGPOmcGVK7KLnm4EVBim9Fi0LC5O4sj1Ef9Hk6u3X2tZ1X3paZXIH
k0rbMSMnh3b+KW9TAPTZ9I8BhPkFP63gLHuow39Oydm6fapBo6tPPd339SXd/GXqNnXBSgruHKvl
/9SPatwpumnyLGKbN+fV7lSeg5qQuM681E0wOe0lQLUtorEv1ZZTz60eP3i5LFG1GU2fZy7bwdZT
E2n7hvXCqH9LXFO411a/S3I/U2vKqCR0Oiyql1iKR6TBk3EFG+JjGpjppIpcRxqnVGPwWtdM3Jxc
1UKrkvhFnsgc/cXwTwLFmlrBHmlGKHlgmE1nMWmuwftyGltUILp8BBUbKE6IheRXdKjxeRj6kAuI
GAmiDpEa/xz7MNu1s7tm+6s8OLmLSAoy14UDb0RwMT8BGb8XfPqWY/WMKiqIex58dpmN6wAqSLAz
ItzqN/7kjzobTGU/xFn22Lp+Rl0BosFZW4UjgTPgAc2C70eJX3RkVi7VI3/aOwMn4X8k+2vgqId8
Ln/IO3Mqze7SrnUzSBe2pZ1DjBNAiSID4KkvVTQuGxWrK53qz5YhlZCKb3DnqHSrYtUIs8Hynyyu
8NE6pafiE0l/fKlPiQ/keAUCJiHIViAcSwuH2qBkdlzZHXyVcK2VpujrBd+DCX9K7vWA6PgjR5kz
iLQhkf0kG5rbkP31vtLDS894a5U1bLf/UH2JAc7I2Al2ohk7elmxUWFv/WU3VRzNRq7Y5CBhZYNs
pE/7LJ3BormSiUDm9w7u8q2KpuSBgzUJr4ClGRGAaZQWX0rkbgzCvC7OsNNJ1qVjHWLSQTPPEiiF
tkgZoxf8WEWZl3LH4MRGAFvVjcLSN9w3XPlQKO0+I1d3Mbj27tOaOiOyHa+JCQu/4m4uYFHhIbwM
FvrcMjL+9enlGyuTg1JywdpbjNXTREdsO2pnSljyjV6JVMhTtAf8tEtvFmxhFEsDAn+/r/Y179pz
9zBUtcZJfqijU6nuuacuIgEzwsD7vfClwJpqjxIp+jjg3aa88p80I8UaF+FNTIR2yr61PQR4H9y9
92d0nQq/FhqV020LU3GG5PfqQVKzS8zQWYbvOcbbFOAiydU9cRf2IWEKOHhwGq6C9Hn3R0TWA5ee
jqznogTBWQXCqAmGLXEG8FpViSeRYcoui+5PtKwCqySqxEgiyFs2+E1wpA5zbFvwQGwfSaYd+a4s
zlB9nK/fWsMyJjyz1gUe7Qss66UNitYc01inJWF2aLw2ple/BXCnPjFbWRwF22pJnzHbAq5G2QRQ
R4s97kNlpHul5ekcou8pUtpBWYkBgJIiv0JEK2Imv/a8sbvDe6p5ToIU8uXnyX0l3DN9qEU900sd
tSltygPEQHyCJ/ZJGkw8Lqx8LpjoQC8EMBqbRzZ0b5XbPynxvGP7W6VUioJpMuXr7f6CTY4cFI1B
MWFMTzZN7xLW74fcapC5Smh3z4/qZ5ZHfZJu6nnEeuPOcfn/1xHqNgmA6X6MOa42t8wFXLRTYRaV
lxwnMNwVkMW0lXLgefWHYOVTQeLvXHzM5/vr/mGXX7UoCOh2mD/5OHBQNQe28dc9Wg50VmDr5ZRq
oq2ZL9QspqYHsTfXjc58TxUv/QB+lLjO7s39vIEhcdwVzBrK7rDusunQaCQi+3HZASsZoTjevQ3L
Cb2h6ZF6ocj+R5IFCboNXgUhe4wEey/jEAejUggQRXP74vLmiPoYQhgE/QBfYLXavMjcbL+GYI5x
IiHAV2M6JN7cFyb7hpgOtgxdJfBMcWo+QVK49v1jF93RQibofr1f24FV46PUahdB2ACEa+fm0Fxd
AlxF/MMiVBCSV7G3X5r5+JRZ8Eyx/JUFaXPNZWhHwpP+BzD8GOK3Y8JnbXtgJSpdtB62+4QeV42A
XYqOEfnBD0tKPqixba+aVFAIP2rODvNoIo3SXxdq4y9RrHZ6jdj7dEPspplq1Y3NoDsyevmYu7NB
GnNkU67NRP7O2xhvpEHNNEFEMehoBc9kt1ZdbZNciqglM+fINYlEJKenW0Twbv8MGfgtduGLdMVY
TEuImQF0zgzaWEpyHeR1jgyCKPBx4DWdCX6GHLomaMEN9Oqi0m1gLY0tpTlrUC4WjDHZN8VohyXk
/0gmywp4HhzSY7AJKEmuiAFAi0tprSr9n/KamjzOj52UFFRs3ixFaY37fg1mfK7jmvFlLHd/Me9J
CgkOwyKkUIMqWq3qLfaXTeB+dqgMmAG7reKxCBqV7xFs5nM6QMnJyOsg1RZMHeTFXWGnjvfzu8Sx
Z7O9BYQxiWxLxFUoyY8jsD7C3mvAdZ9n6hWGjLZxFKYBvYg54kR+ewWDOXxH620khkAcNmIqUPTX
5GH0ruM0wC4jh0pQMNn3/AtdogIc3cxaXW71ajSeVVIfQhEAZb+YqIthWuqLDM1NBeDFefzXBL02
V3W/Ku/CMefF1v6ByG7pyBJCVHpLg4a5p8l6pj9HLSFyDO4qQYiqtemIwVUkK2DcvSiXNQJMd8Xh
sAN06ensV+MzBViYAcIqjHVk0/CNKZVL4OF7AB8/X1iAxWDdvDOgdWyfjMqNWqXxgQwq8brudIWA
gcrYSOWcqXXsY1Yv3jsNuOBh281X3z7lCnFvRIbeOJwv+GuTEABmnzAp2GEQzKtPtKOGIIfBFzda
1NJgvGlQyjY8r9VvNI2Pk9e5b0t3S6hf16SyaaqbcsJ3wiwGaCVNfM8tGfavA7rT4RKPSzWF8U6s
g6swLH2WCtPd/TxShiTt14t87YzGG4XLgX3gT+bsvyOkeqHns0TfhETfk9tL6WdXZWLw/P35B0P3
6dS8d201T+E2QDQEeJ9GIipx79gaqUeS7LgzhtobjhhiqSyMjFisevHtPkjsP3tSZRbPpr0l5YfR
LNdnAZ5xlaIB7DuGcY/ORo6ZandLB/uzgQWIbO3Wy+XqrRZs5xzcODKVcqxUGfOUvnSJYe2YB2r/
YH5DTLazFEXHKG6pbjFBa3SwoPyxebc02IPFN6JySbQUWVQc1gVqZ4ZUEsHJnSwgoNn1dj4bB55x
Av6PC1MFfEWiw5O8+qEDPBlQRER4IjJ0up32of9YYGzHRzECQUlZMKNCsW5d7xc8bSzRs+iVXJnY
9/fr1b5fKEZKGf/GiCba+XkfMHI5bHQ3NPZXWMq9L2zveCoQDWZO/RnBgGuzIsB7a8oeOkJI+UXA
KaKcAN7La07ykUoiynsSqxQ2X1DTPvkqOG//TVdggW66G6xLOJMxzDXLjrVQwRbWXRFhrRUTYxRx
Pbt+pC1muR4AbPLIe+zd/8yLkxcEC4Jv6bop2MlsnsGbBCsn9oqRk+/vdtMZR1j4Z21E7zOOBscq
aj7FYPYD9Or+6e0bRbOlVE86bEbePWPzUK2ct7KnhVbubmJYlWKViuQBgBpufnajHWs3wjGlRN2U
FkOJ8u1jj++stGDD5pbZt6SJTB/QmENrHsSgt4EwZHJjELFe1WE9bvDxS6YoLi1QtQGFtPO1/btn
AAqfw/ni36+Zp9hbUN63z6kXixCH8T5sfnSMKt0IvfGcOBQyDCwCWp4O6vV9HCCoCVEcUC/jV37x
k8HjjLvfcsSXKn6Mm/1pW6kC6KEq3nhwHly1KvYjVxkqNQzRpxgB30Ps4c2Z0olOEJnAI6qJuLT3
yR3yVlNNhHhHNhpRH/DOM/05ncpkFlJP+S+PwHOkMm329VQHzS9TLsm7gBOMC2zZlQsWvOgyWJHs
eQASunOWz1Ol+CfbZ+sOF/Qb7a61C9z2sMn4rpUW6LCjwwGvRf6P1It3/JeEWgCY0ydKKRjxzL2R
Rm82ai19JYFgDtv6BO8p3uYDOzO3f0ZTm6mM0XFztJ+qOMzSlT9zhLyqvhb3N9nwJ6gxy1gJKB1q
hYtA8dTZ2prAtIT8GjrJBQ1S2bHIt9rrwRfhdq4lEaQvikyLSJ77jB+jcwIB3uOlvI3sdwVsuJwp
RrqvNEJ8dSLtXjg3heLOrklwuagHQvXorpcF0enOL3Exd+bhgZ+c2XKrNZfWdGTDW6wCzVu9jxPH
wOA13tcdVu4JujJlADqRxAyr2I9cZTKe25+tlSa7LxoBuw6kqVekRnsZ4kz31gFpa7qUsw1xMllg
L+mxFEvMrCj0/Ok7Lk6S6ByKUKWEoPnoZv5DV5Wer0uxbMl0eGR7tEjXzJ9qNdIINZo6RIAfH7Ne
sWbEgl/+0ZkRT0FiBW7meG44f5tXi67MgErDcGe4PphkS1VnylpaWp/ZY4adnYARYNnO3tNYpGJE
F15l+GjUY9TGmsuOp70S3o4kLFnJDMMzTgLjX36uFPMbHW4mNQIV+SUoVUnLLJoPE4GbC3XVKxww
LY8sBeO1sFxBWRquFW2cdGY4QQofV/SUQ2+nqsWXUi3s13C76q1AWNcIesbLw6YoXpjP4qaOL2+J
JoHpDGRGFlDPUNRjgMqYFl50ioxdml89gDRTCZjXuZp1dZ/zQeBhsaJnltVCMTjs+d3gu7aCydoY
gKwhExpvjL4dBBx0sK+HnYztTqAWuNpg68qGo0OHGHwAaCAqWlKi5ZKL0llIdDCrSfLf3w1dAaGk
r0vC0ngdqCfoiECgz8MgfmN53gB31LWocN2zDCliMwDMW8JEiZ2dFK6BKuGdkZruF1YwfVlyV5V9
Qn8TpAw4xyZC7ulnMBzO7ozLpFyVlcLT9GRSJk0KAyJzq1L7iZLIR5alMyXCxxaH+dIte7EJa0pJ
x3Sy0/DvT+2U9oR7wIM6P/pl7pbjIqF6TfmGiAqTrCDKLrplx8Nj1gb1AgJTwdmO/eTVbuznV4Rz
b7CAsytFxHzFMH1++fnOvOSjuyQbUUZhIvcenhKHjRph2+MQBDHk0whi3o2ws7v3b3id88IivDeO
2Z1n42k2w36WUTfowzgw3yf7Gjbmh7Na3kLIqU7ym1KJLXupcenKHmT91t2U8hCrQkMlaWds6orw
NOzYA5sL9HjP6M84rleyTQXocM6WOeut0Xub+vK10x+TEt9YOu8QJdYOF0xwayxqrLLx/R3ieu0B
MP1qThSDV8FLuU0IpW8QAEpFxQg964CLanOgKyF7VNrOc3X3OpcgLFU7DwEHbBGZnXDKg2XPRmRJ
34Y9164VU+CqTbzW0ex6KAmLqIznyS7uvDbHsnPr9RLMAZOgX7V/f0fCUtD/OnHMgRi5dP2PBCmG
xrQKA+K3HWi0iUqyjvu2Ycin1JZYAQKVLNAYfoSYAbnqqlgbx1URldTt2MZZSTPbzJaFbAwygmEI
wSr2Si90f7C1HFzt91G/oifvfar6Nu+nXJmex0sx6772gnPN/OXIKlozgLs+N9qCg/IBaGR5P1wW
S9zp2Zs79oT/sTZvqLW1ea/iRu9tKlS734WsqWHI7MncJ2A6zOcxvGsQXywRvmFPUe6xzLMrF+D6
o+SWMxdDG+CC7vt5KKuehgO5XyB2raMKJEJg4wrT2d+E+VX7zIDcpBsN4B8dG+5XJeVe2kN19sfN
68urRFepRDfzqcPUJ4MaWhw/p0Kp/uYJOZ7umEmTbk3EpNIghOCm9xvEKhj0DZXzU/FeXGX3GRtq
K1z5C89U5cD2/p3Pa1oarpFXROoNF1OcrWMKaWgYHxtiP9w41fO5rq5wpJJADZZC7w0oNzU1iaQg
VmXgJdr0h6MkMvicqX133LipIvfqouDu6ZYrW05L2Jc4ZfgMhMGOkl+zkw+URv8wczNvmpceZA8U
4sRQ0Ba8+1JuINHkfpdJP5h0wMNhlrTV+zZsIi/hSG/W+L/3JJZVmYBH0AFq3MxnB+40rsyX/reG
uDdMiQhV7ALJAvrgORQEsoljznnCPkF+ncQ1ajXFXr5zxXvIGp5CiTY3ZFYhIXb4giSLjmVJgvtA
m4J2M0k/JE27CuTrvgXHXVcm5Ve7laT7p/+9zyAqI7MPvsrMlAvMJpkMoiRW50D7NKEg7+t1lTbq
3HIjcHBVCStmnt+YKpdjeTxjPtQh117Eu6EUZP80YZDOScGSZU4uRn29GL6w6QngB6LLS9m1TQxv
NAY5xn20XYls6Nj4yZhspHZDUfbGOg0MKqnJO5+rNTBh5D5AgfgQnPnmGzZVz+jR0DpI3G4F5UXp
cf/zW7opi9nmfI5XAb68YIqnu2WmoWlaIR17E3Vt3zJK/9bce+bcywLSBRiz9HYZMFHH4ZCOAKsA
tJDyMncZIux/4H+f2D70sHmgoffHFNi3wQx7qIS06gppAuSpbpTl31heypiCiBqjg1+znuzSj4Hq
uLRNtDacwaefUeuRISQbHE3Nhz+bNQqB+sR1U/dkpqKwOR7DItPIojJSKLoMJPojGnxmFGkWY1Dr
kgTW3mYljnAS81oMrjFdAvfwkJxWRf3RXfEAqATaMA0dElzX++VyCQY13vARpA4o3iZ1ux45z3Ed
yL3bQ2hEj9ggTD2beLK7RtmTYyKcCD303SIk26HMVm/7HYHXa1+BzoMEBe7e10iGRXaI4JHe6J2F
kslZZqOQshe9Ubp9L1xiNbJnK5GE9Y1STBPOWJ3qGdf/Adjjyh8GHeXTIbi9QCRv9frjUwn21qA6
6PL/xs11E1Bn/TMOBCGTqfsSUzioZc7/eF7nei/eMZcezCrhE67M6Im6S1lo4TDMr1awcnHUKefR
A6TFLivpKjZhbhWyXRCgh/da/LCwNb0zwDYaEQ+d9IB6Cof2DjMt3hH0wqBw2j7f2NP8PBvHu1vk
xz+PFZUu8GWUUuvVRHQQhqfFyrEXTnZkdIpcqqtzoy8JZllpzlGoVWP6tj9xKe3POa+4AAyTvj/8
2gG3E2dT+5W1G1NV4iNsG0GqSYgdrH13oGcVWRj1vwmXH3+tlavdvpMN6xHku+okv4o8yFHIZMlh
NAMfz8sX6XIbWc2G9fpi9Ba8iwmt5bo9AnyQcl7jZZBFYJD9SOexBGSy1fyw4IWwwUReJ6SjdO+C
WIYn7+dskQszhEPCrRr1wWypvCZS4Z/iuPlANdsBCkfM+/Rbd08xH00m9hQIHhDRXiXCy7IBUuMd
CIyoNEis/PvckRoAwlGAG6iXcgCR9GVQBeLtMVgzQTcVXf+s4B+kSEdb4haRU3VKA8DXVvW93KLH
+t5NZhRIxvHVdLGNwdTMPc7knAD4Pik/Mj1PWJL7QqSr0Fll8w7drMWE14vPR2+j1KLlAATkxjtq
awK1JSSRIF8LZgFh03WFON4gWaevx8/CpZymxgeZII7vljiyK1ufavfLwBGMP5HarbKQVaUmpQqv
nkjOsKHQm7CV4fDoi/s5rKxRlCUhxy+GIlfMGUvYNQbSZm2VxDYQN9/oUTDQF0tPOy3FZuOrAjkI
/uzNACi5hjpZ1MeMdBbUDiMxeRGtcfdOZ4vElU4ANjuyTtxaNcHq21XtkIC1ZbCzYJP0blf3jGzV
E3Fq+F87fnuPx1Gg8nqMvO42rhc+9Di1upk9InfSlDMQ3FZsK7B7SPf0SWrr3K2eiY+dPdoLqZfE
Q3L5ibtgx+PT7P7iIh7Y8Iemwk2DL4wz0/unNLDTQ3OdUbLX1wndTAyYCuVTKC0TVHnxAAnb1VUu
fTOjywGqmb9Th1K6Z1wwHPcPK+uAS+Nml86r0vZqWNOH8T1yxkVldB9WrZBFyb3S+V0dxvTDxcki
GpJdGuw49lW8gnApdV1WbO5GRAagad3eWplaE+8gcHYIW6m+KX84nikd84fAo6SJf6ioNCRAufyC
Bfy1eLpEwSVkmtuPlPxBH9jf0y/fCrsNVAdeQzINm3LnYtTM1mIKq7RoDr1mjGK74O6ED4PVWOed
qay/Lopa9dqnckjAw+VHirb6N/sdYTATx6zHisjf9IdBEPq+e9bVHlJVjFVnNBFZHqEGAria4WHE
jxH9n4VW9E07QWELrbbdfAGpiHFj+z4LTTUT3sXq47thmXBEyiJTNPhyKTOXYoQ27xG1tVmSKi+m
zhN9rM/tFC8Xy6Yj1W4ljbf3DRZ4tk2t1pj8Z+mi6g2lRG1sMt19auS7f1G1KomslXfsBgviN4+q
axL2nY29TzAFaUwYjL9IrgPKI4TLZYznxOssHHq2eICNdaqpOXEYtlaU6Kq0W1lgmTzp2c6de/nQ
Bb99rtrDD+BUxl5zjlFpammrTb9NCh2CIpKGLTvgmMevPCjMu+WKWvbP9KqrN5eTPW+24JY06nco
WHJFWvnM7i0fohg6B2sfON/52XnvyXUl+v7Zra78asq1UZcA+yge4hrHaWJJm8j+DQyrzKlNgk7T
4qWJW27OLhQ+L2Z3JfsrlynRx58MKBgn0fUTrDnK/TR310PTI/fp9Yc3/tD39Q5YxZMOzv99qBwJ
RX6SAMcbiTWKOYo0nxW8XJkDGVO2g/xhLo64V/BuSy8WMTe2gfeXVspuHMnyKkKVZGPB7acWwfhY
pnN6ePpUp0mPTbqmqm0YUQcPkRl0eDgqWK52hGRHKJjDkscrgcAwKM/e+O0spn0wZTSMjsWPO3Ue
8v7nT0//vHoxTiB6F4DErKZ3polvd7EjdfTGHQAjUQnW7+yt3nR+8pn/clhokiggv9lUHDXdqo0j
5DRnSLOYjPVWLjBgrRJJMcx2eSNXkNVi+yDHUfTeUI2Ta4VO5IyZHxQxDj8YXUwL6y/sJBazdGwU
e9AjWgPAsVZ0aRxN8fSKLILKRjdsTpj/sgueK46wyX0Sgk4fdVWA4HMUeEyyKz5WGSdZwkz/v75C
/ucaiTx3sJVZnzhWTWdWEEb54V5yWsljaf5uy5yUfNFpSXLqt1G9TRDrRZywjF5y+/t7FJLmshs5
CU9W+EBMGtFjw5O8+VU1bynAFCll87Gwxi0+LBIIMPYdEZr8uYbQzj+/S6bg/xJ9JEXJvoSP7Zcj
pC01eBkkOXkAyvr6KTI0ltXpcPoykFlx+9Ewn1BFqMPgOZJThTdQGz6Cme1nTREesLC0w7bd4Y1u
31cMKvlOXjM+1jCaOL722RLbJr/CpDpNlFJOZRuxc5b3BGrgGU0Os3Qh5TdQe3Qyn+LzPWwmXpHw
3v9aQBJ/V7IKu5lmpq4mK0sqB5xIFbUI2ksRUm3ZzYBynioIQew2iJIjjMj/vuD78yLd6BVyRBYc
v2AMZHJrbl8bG1DGLVZWUkGXIaDkBQibDdIKgKLfuAglZEF0SVE8fVbF8Rix3a0MeMJGMORVBMFD
pJtS6uCjTRQy+nBlIeEUz2QoTcWuxP/BnuqEK/uUQRQNmG0EZ4MZo0cnPpimf2G2MuNR5lfSSaRB
DTeTRXKzR678vdXvg+LiSa44jQzJi1Pr0SwlUYEzg4wVAcuu1AW3390qgLzLZORVS79wCipU79Ta
xl1djdzlKGBHMKtS+u0C3JJo4HLDBdh4d9O+6q5FtKe4WEgWCj0MUIW4ijjdVBVlbQTYc4Tw8zr4
YqIz09/DNafBuxkIc/7sV60ItpXpTqRiBeZKzG7S2k+HAJ2yXXRWRK+Nh4abNu5JaFQkBwNpgOag
ZMYU9trLtaEN/GrqjgBn2fkGkClIAyW86i6E9K7g4L38ioO6P8DP9s9TXEhnG0pqTvyuRsnxs/At
C1t8NycvFZc+rMP4Dv3zB96GygsouME//3f0YHOehVv2FRD8XnFi/ootHXHDKpzBCFfEtPUNalCN
Bj6SvXba0rTOU/UFOwQufjK64sHY0fRuD8aICEuyOhquQ6i+dzFMjjfaqT0J6a0hBl5IUT+Uxdp2
5icirvplLnAn3DJ2yFfbuKfhGh1KwhP77DcxY4PiLvtg38uj7VJ9zo6PtCHQmhcuVn2V51LqIcsL
ZUWdkhMGAtbsyDDnrK00X3lHnFm2skLUCWVpoX3A+6d6X3r85rAviLiOH3F8qVk3s3f9FQpSC0Kp
mTj4mNh2nhmx+2MBxPfKR3zMuvGWOzXwKsmZh/pRj1QylGWV/kqwdlB6VzxcnPum5KmfvkSqDEAg
vAnl1V3LWFFJMBYvy+pB9srrEGrWMlBya9kp08v6t6S7H7qkBYeMn9iZ3J2o5gIOeu6Y9PzE5KIi
DnLNttOxMVrg25dWkR+2sdoH7GB49/bGVJe4oyz+4ZUizCZMrSScxxwnebxEWLinm1CnBNFGjrlD
QBPu3+tWeylcQ+dOp9kmg3XtcQJ9XGNBYC/rohsYQqtwF/ZrhF+dHcpZ0tbI2CCkWkF4M1ftBaXZ
SKqmrS/bD2+3wEO5rtycIx/CN1JIaQYqmqAWstEmkX//kQ3VxuCRTNIlsJD7T0/8zsicwemQX/Cc
TeC/8+BmPH6khNQsHA7MQtnwXWJzO5gLc68IYPodLEKy73PehYv6jOTmU+XbUpt31IeYnnELITL5
Vr0dH7xzBuYmgLl9IBu9Sj0qwT/0Qmy9y8CCNWaAPeNuU8hjV5CPIvyfmbbNv3UTvSZiOk7yxbRX
iKiGbO/1hDkObkA8GkF+5S8eNQAqNa2I01MxmM7xFzTL5+GzhT98Z9UzO3e1XhJ32PRtQIgWdKeJ
PEbVsmuhcAD3Da5eRx9+DZfQJXQNmwgxz3SsykxVA7IDnBf9yh9xxd8rC70ynd9dfa9wU+BXro4l
GpRymlQr6AHBlM+72dEet7wdLhLz+xoa0cDnLwCUbHFLwFeCNJhvIXSxkguSxQtm0cIb+0x1tEYz
M9W0zhEWMHeDis0Sex0m/BVyoKxeOmm2D7dV4mXARkP6jMDLfjjilTgSWTdL/KzqrAnGetUJ0n4O
krbLcAEQEdW49wUfgeB/dLC0lYZGrSQUbRj2HhP53hb3/x88tXjbEH+pwmFMC91H1X0npq27WhDN
dNOrNu0MGsXnQb9nPQ20JH9Sg7t5qsAEDiGmyQsKpqMgYPM3lLe1ZdfvLcxIff/3gRJRhE/tCsWN
a0SymJpCSGedeIH5x/k7NJMZqB3g4uDLuWzI1y91j5TgAyQwB96vAz2GZ5p1oxbwBpqCz4G+5Hlo
3ke/wzr815Ceu1PZiDpS+Efjs5npsVVA04tiEkLXFcIamIFQTj7kf9VTa9iDkJiKYEk0KybE6RLL
nlWcjSgwxtCw8Ip9vrPPoedL3tlKzc9x/eG1CBkX1XcEB1lLgJcDlQPqMsPrpnHM95Kz8fvjgo5s
wrzuUWxrHBGUA2+viF7TJ7sSMJ3CjD/8hUBQ0C+CUN7GYbmGm5a7/mfCX7eKs3B0gN2i/acQ8dqj
UYU3Wf9TkAh4KLWQQ52XE3kC24XM77uIgx5Df4pocvwN2HFHDHsReBK8//eF3dWrYk4QeHe8I5jy
xqx44yQG6HBSUJw9CHgipyEdQUoud418mJi5suMVqer0OY81Udpg9r69VsZPkTm3lXK57T8mHzAo
jSP39Tcbxdcwg+Le4IwrrYrwavZ1WhKUigHaloAWYMjCh0SL11cvdpVweyRZWXQdjHoidJOau+03
HlExIPyU6lhvFxfm0XxjlRfyPn6Xrn4niYiIWHzBnO0enAQETuCbJ4bpCznbq7tnpwTb1mjqGcS7
LXbJtB6LuCDUdDbpNouWEQFtTFm/F54fh2tSgSuFuvGvxX6zJEX4Dk8EbfBIpB5Jm0SHWq8bQ6fq
80pUKZOHWaqgocYcdkolJIv0WcOZ8GrVxipWCN7MYXFhS+Lwl0y9Qhj7UyQnRUnnCvG6lXN4Shyg
KiQJ+iuWGutm/165P03cj5suvWuy9ZN7DHtCB8i0jOiqScW3/Xy9vD9eLMAYs39J3s8/zdNoLgK4
oq/aYnb2galGXtfg5fiozmpI4xcCXG4EV6C99eSnvA6QgrOeNtKuIdFQ/uHbp8AvuH76Y+EYDHnT
RM4ki7C0HzBWQAFsK/yJQv3MEyyRjjvQxWKuV5cHrwdpYnuZr0AnOY1IV4MVqsXRDWcs+ZImatxY
Llgvgm4KLN2tGLtFXZR99EuZRkjUE79rvoaQ6yuktN3LH0g+bcbFrzXkvgkz4sPDrnXiBr8P2Fb6
S0MxbLJsM4TahVzFP3BFhzqkxRhbuviyCucOdRdS5xeKz5vSjd8utcZd4tq1CrtuHjifJLVL1mPc
Ahk0bug2LfRgFTWNrcTwz+A1DhMAlL6EpEDcZwy7pKv5vF7I03e9OIPAhG39AZYAP6Jx1OHRV0eH
o8pDlOXHc6IbwkZoCD3Kdl1pFiwmbFRvKd0C8nCM+pXqRPH1YXUbeds+l0WNHw422zlpdHqc3iAz
0YysXFTDmAWA5Qm9Uj33QB27r93apcpOvOiJZhWjnFlZZbQIoEm4n36WS2XLSJLtKqa7ZPRxQERp
tD6WZOEkstsxMMY93MTo0fblsbc8IhBCXhBg9LcCIqrjHGK4FmpfGrUqKYjFBokuNkimi4mBKHN/
L0JWyiR1zPzzBP8h2bMyt1jTOwDJt0K6L8PfgUiX1bY7fuBnvWEeRCrZVJ2nYUCsAI+jc2opI/nT
WVc+njYneXr5iVLF6V9hZ1hIBf7W3EokDQskpRlEtdQemLU92eVNaWAWxVW4nWaTyu5f7lKjib/q
qHesGJ9BNCrfinIV6OgwsG8XAo026YcbxdAtTWIxSqdeQvuZjE/qkDxvLAta3QKJut3ytQ5yh0/8
lwDB7VrQEHb1YZ9uLgql3QGvc0BEzT4KafGFjLWQtLKilHBhbpc13RcnXkujPUmMxr6ixvN6yYai
SMdqsgBatJ5M0pmGZVzMub9mvm+8JlwUrlJoV2EwmGzWeM2U5MaXp9kDq3zc3IBmt/eCkGz9h2DT
7dwr1aki0ZGAMSQu7l2MQ3hWPRmZHslOE9YYsb46KxhsQGOV5UONLWOECDPjBm8A0bMkVE3mnwKz
VQ1r3O7WWd3aYz6DkXWOYQPDYlQbPpAsvEtvGzQqL4WTiLwOv/Zxc2j8dkDm8mkPUV/963dnh3oS
zkCcwPEhBQ//5iPauWt8PuTmB9L2lCqK8A3fV4GfiFPvmftUmF4SbY6DfZcbdBZlVBwKYWaVU0eJ
gvMfoJejHedID6vX4laApwYI0tm78Si5UGGqirQOTh3W4rNz0T96q3aYzXNLPb0RxA3le7gfDT+0
KKyepEqcfMH3gl03Cq+bbgzZU6RK9+PjOjFpySRGL1xqbw978CZv+QH9btVt3zPCjYpV1y8ZTYhH
kMFzvwCrx42a87KKh9wGEQtVaGd79RZzYDRTildTjSSpOZ6phfFKzb1iqxzx11k1qbxwpiAemjSG
aePHw/ak9KXvAqYR4ytgVorA7LMDfRWve6BfnrYrFiWEb3wvAUhgiXWDerT8UInX2CR7LFgDFQav
uOUvPmA1xwcqyS+tQUHOhQBrKhQDlKxJfOsIgIBjAmPrmWw+rETnlHQOVHmHS2+Hut+4XO5UXjI5
DHGUFSY5oDlNoVXHNhnbHW75BZqY0BLD5mMmGD69d8wCNYF327gVhE5EgEGIE9vT9l6odP6JICvP
g7PGtuOEHq1Ry+2PLZ9whH5vISLuSlrqXFNptJccwZA0UmIVACg/sAicC2zKUmUxkE/fOjkdrPxa
W1mqLbhqBufOqQpS1ew2ExqGGJF4fe2Uc6kj03q3dCkGyZkrinYHhD+IaBYx4ZXyvmEUbM9TAlly
A7qQZVPWYBOqhJ2zMgOGz6P1BMJwvQSkZpsl4DrBSRxlq2tv7dKelhbA8DRXZgCT+xcoVek+cuix
SNDKULZI3vTFPXMFp3aISOE1sobEFyBQv+7gsTk1so61EaMBC1OG21gtZEfY14lzC+/slAQ3K7Dj
a9JswvsNWz6p8j7z+yC9B82NE9NxgO00OEp0jAuQd0oJm3C60Aa4itCOD1/3KIYxMiml+EdGNeuy
Fp+wh0RziU05lcnV0AhA10Dm1+nZh9AapR8P5xdQoa873rUAClGCvfDF8/kq0HAOMTMPB11m0szL
jkHOD10ZmJJk92ehBQT0koMpkl/mOBPLUtt4Mc1xFzdGN5uUcYdS5HTo5OVFvn1eQtwGlWdwbZ5t
8H3+IXcdTtEnxby19IfmudkPMXKa5Q830bPE12Q+sDzAtfr+zNQDjgWSFRgoSzK1ezSCr3qK4Kgo
DglyHFxkVzaHT1o8delac3xXIIUVmUW04wo2IpAfLl6iTc5uyKwAdHBC268oIGxH5Xy2k0eIDVQv
GQkRNraAz64CCI9TMBE7XbXiWjgQHj+c9Vfiw9jmVHCRwhYPdV8YjUnjuGu5MIgIophHbteERNj9
gw6jT5piuHJ9cXL639hdMGe3FdeztzcCmbPx+V261cgoLzbBGhUjlkWru6zzBM28unz48UhGlSaw
Pz0+YzeBu9v0xWf9rzbg7Gni0sO3Uj9sqNNSNroYpAv4FUd0I/qFHaDdPG/2CEI6xEir3ZaGWz5s
RtSD4GXWaYLuMMVciA2y+zQWEgRkZye8svhu6inwazz16n/uIW7GeDiITH3Ku2IJxe2taj1zGYf4
GthdEt5WEVm2ZyOSrCDk66xcECLjA4mCIPcp9D3VNyX+GJERbLqgTyq0RQNN9pbxoi0VtM+h3mE6
88HkYzB92luXfWLxhtp/9srM78B5bbJIHRY/UahoFoXCzVCqcqPuQ486JYDzSurUmTREs9UQ7WR5
KEmcsSJ2aU374b/Ggs+sN+o38xgTxoJDHZu4GSir1z4cBkA8YNu01IaYysO5R6dxi9I1SAsRoL9W
hu6jxU0k4K6HMqr1g7pzEydkSWFBOg1gluCyQxWSaJFCyFdSHHZGCFRUDeA+CMTYPE/zhgSJA6SE
SCL/nKbYEF32dxMMWan3F7dh9WHhLJprcU8YDorVnAGiik459NOon5LqaSZeUh99dMKtrWQMhykn
ciGIfrGQV4yRaz4jAMgz8ZLqPBuCLrv0fO42GqikCZuPMkItAgGvl/5eZI1F6nFL/8qfzhLuevY2
TW/qve2q3EsN3CVtL0aNrUO/kGhkf8V3ap66GNV61egWDTo3SYfywV1X406vkcO1bCBUoueCyjBO
Mddh42J72vR9f5pWWL0wM+o2DeOwmtiqfQdUaxJCAe5mpE0/oCfpnUroYw8432sXOdVeWFfucsQk
2211tRUdPsXMKKhJOCAp4tKpbC3vMM4/6YzpFir8d95/E0kDiK0HWMujzcdbvO9bZBklcjglKPgY
Tn8l5VsB9kbEl+JH0coekgUgHV8hKISMb0uKTzcU0EAFBw2UbEjWiiJB5hXYDSp9+QgrfKU2j7P8
6xGxXhskkPwhfRj+0kNc/4q41z0k1yi+p84y5wq43fk9oYyeuwP0TM/2ph6g7fy5UrqlpioaeIqp
OPTJbctUh6yNTVqwK7l97MbOx0ZFHdn8K4jjLhoRr9fXIzamIfY5jOmSwWYyYrgcKWnN0xNVKbS2
k9FQmp9yVQPUZ89VjoT4TWW3Yxje6xeh++G71n3MJWleKlMJttDx2fbtOUtM9jVhj+qBEqnT5Qgr
2eox8ytVlLhhAhf6YG3c+TBluOk6D9hYAirQL9nRk5jqR/y9Uh35XgSptbJowJX+McYJm58NDpNP
4Fjz6IZIo2+U3Ss7BZVMLEIUBKND2mKkJj8oX89EILEPD5QDySBug68kU74wLtEy6/X3kH/taBYi
ORk0Vo1ybMsO8EgNJmLIXRBiypTfyrcENgLopBofQ6z6/TiAwOAdGvcU5X0OhZbOOiB2ZwhlY6ey
aU7CSg47WulNW/UCizUOQBfn7drZtGucn2HgY0wOF9v1IHd4m+LpkuRRlIAPLAEPZEvD8Sxd2N18
3DD2wMVsGI04om1z9zwEeGqqK55tuQ9ZOm1WyY5NDeVjtUB1SQiFEFpQEoZAIw9aXttqNafbDF8R
rzfj94bzMHMMGJhN6lZU/kTI5HzpbKB7G2b4N8wzVH+trxmx2UFnbztvMni9/c3GfAXboWGAB9dk
34XDR9BvqN9kUOrwvduT67Uh7xT9Ydj+79eb4j+9tEZS53KwVtZeD/676913mTfnmbkT7LcOiyQe
8Atk/QKzFXUoEQMxmEQ+JB50hh9rxEPd0qf8ROMpmylbbdWyiZOM/FBFJdSj6wY/R3VlZnhFm4o0
enm6dp/e3CuesAlBZbtHiOTUmwbNK8i6AQsY65MHIQRudHxAVRgScj4bTH/ALtDr8JnkbioUl5Aj
grsAyhZ878xno498CEf+kMVqLjNDFAyPWN/Ys7pH0ugSQVjITYp5kiQnj/NJ1S00QD3Qjs3DzB7y
AbXklUjmHAwe6Z/90L+IDaSY7RvOKLBYjxV8q46Gqy7pf2gxR4LRFD7UflSO5UNpKZJkev5irWIK
Yx6kjy6+QRgYiuzoCMmYkIaOuPTgKM2ahnDjWLTn9lBIgDBz7ksygZA3yi5OTORDM/jx+f54g0kA
fz+3/DPKbVWIR+kTgtxc05xzibUuYK0DO7M1T6gUfAjPAc9LVurU93oIpPerW98AoFuew5mqQ3jM
POFcEPJ7fgNDWmYTNkIwL7OaffdN5o1GN2mhfPf8MfvdMeSNqvb4h/ilXqoutfbxdYPGyK+bRZXd
Oc0hUdiLPqawSDtPZi77wrbakVfMgvAkamlb3WhQwUsBNql8+31lx5Tk4MwDjbqdAz+wfEmmCsjE
urPOeIuOhRg3eyn9XT7YYEoHrON8u2l4SYrCUO3UeM9GCUHsH3KjQlTbLGJH9XZmVxjP4MLjyW3W
MLG1UQbsAleLZ/265VZVxAChhkh88hPwYlz/oXeRpbk5pkEEoO18QFIXAiIW4UGs3PJYqW4/gGMR
j8LwCONnFzYuATxr7isjyxvmXYkbZF6LQXA0TqY32a5S7gJIJ+SBUaaffovE7z3QR9DakNVTSpFu
X6RITORUi5NQSmvdMVZ7OES+qsB2DCn9yeqOxa3S+ZmESXrSGCm2sEn+57yXi14kSWQPa8puSku5
2qF6Iil5EixHgSFpQMnZySz0opLf9f7tJx7wwQBdKsT2zaP9/tT+Vdk6J4tdKEvk+nGdDPfc4IOh
/2QsWWWri2notbkIUchg9DE1brLea5o+q/RCtKi1OH/j7jSNXhkBHDMZuKCVfJzf2gwnUFXpYmd7
3E/3pWApE5Tbur7OPEvBV+ohJtwRh0076NFBK5bP+Q3WRk9vl2kuX6IQjScs2CwByw5CG7ni37O7
vKkhr48YVLzV3jr3wRfxdZXHNkgHD1E84VRVCxCmjz6ZDiyZRCMAw5+yO9Ysvz7uQYj/GOBacX5q
mJpuyuFzATPJ6ClWIv149o37UNd7m8RQnjq/ejSDH0ff4Nopf/3U6jU7yEAyz/n9DnddPN6dtX7N
0tGemM6qH/Io3h+KOoZ5LSXNX6IFEXU1x8nG/UTGtAQWoOVb7yCDAl4V0Ou5wnEZqjxLIvt2hbBk
I+gCxyNbZQ9mHBfpmXrUnnNzk9W+or/lcoAnpXsRRbo5nlKry1rDVxvqM2ZluBRaL5FsEQn15J0E
+ZRfAFlSupsfP1PJRX70cKG0zDJ6E9uo7+jTzU2z197eXQla5FcsyJxAjSCuNFYdhq96rp4lqvDb
XwV9qrmvvaZhpWxRgwJhqZ06YCen3BjLMEXgj779s+mVdyZDQ0FVf9b0y4L5PBUj5AZ3bL/YvOvL
VD2mZ+nEmmlLj5C1YPVEccszU9tzzSE9RL4iZ/qpqa7zko9ZC9pK41WUaSafbUzdmhWdtjegjk3G
t+Ith/349wuKLcOk6YXDyC+SirNMFHGfjLAd9Jjmk/k7JmQlbOgyw33kN9jDq7ltZbfyXxW1VNPs
6pla/xdLQi88lH06leISHAnQtdFAay/4TCybUwj816P/KtvJrugS7HFwS/hoGT8gvjUUDonFd8Nf
L+L/DejOWf5AEM2TKO+741UPHkvcGotKE/FaWQe74rsQBTFtuyTXWLXO6gEngJ7acDXotwF54fNd
IEJ3jUfu87kJhJ59RX94XEzWlryRXhoL2HsegRzSIYQ2z11gxAzsWsoPmBFhEm7lgVMEDSfo0cWc
eMmG3K1+rOexVDwqG6Bs7cntoCkMuepddo0n9NonBRQCykBfQTMlXJzB6uTpPu8HFgDTk+tqDo78
yPJ45Qb90FgFOEsuSi+KgkL6eSDdWgXJX3eDjZWD/QoNeB7ToE8XhgLNyoAxMZTYcTopLdVeISHc
ywB2+FfYFpqcI7RaFm6UAxVivlToLivoY1tLToUzi/MZZPJGPsrJlja8pBaSXYUz7FHmEv7bQURI
UB82wr2A1qpGUocXsz+D1hd7qHSw+UUKto6Al9c14EWguQn5vUbAeahFFtMEIcUDBq8IkxnF5vrF
VWqjc6TZ2Mj934Ge6rJ4EvP+BuDV+xuN6ijovvTBXmKra7A5C4uh80Lg/pOSHeYm6BJFliOlJOj6
x1QNmMABPHvXU6jlAziL0NjuOD9y8CfIu74480F1zAey7GZOICiyM4nbLPkkKCENP7gZ7fpQZBC0
9vycwB1jUTI41j/wL4EwR0tdXVgumgdbtb7YJgKUpa5iZL+ClktR8qtpyq+PYVAJ+UooJ13tzCA+
JpANPKH1spKYqQEO3ZLfu4LlWp5v/4TulOa81sBUWomik7WtLCbfVDkhUg+2tcQtGjXMh1uqCWrx
mEzxiLFMRXTK6dIqVVAu0lejwedygrj4F8hds6lXdN5c0fihvJFHYAPI9ZVuwXs1mvULt9nk1F+G
yvQXvpdzPsCltNWKHLfq+8nNDaAExFYe81rQ5QevYHlryIMRjuI9qGSpYb3g/mi7HctMME7R22JS
dw33wToajcElhnCentQ8sW6VM9S44OL/xxGnvNNyBxybM2H5Ka4+b7oDLcAYLT48Pw/znEziVqfh
s51Qlk3HgioDKQtsYjMIDKlQKwvXzdWuNVw5YPZNW2XCqqQRWeKx/gS3A99a4fGY6QbDqu+/Wmq8
42B9ZaplrVt6o/+AKiFV1syx7fhMDB1TeTCMus/Q4JF3Xs4YEvLFnw5/Maf/owZh5fdjtA9Jvd6H
p8BmrffT2BL5FHGiHqw5Fv+zf5f8RmaiEi4yiEqmjKI8lA7OOT8JxQF/jFUToee+E6xHf48FkmF0
9SO5RGRY2IWWhHOnSOzV6JpYLD0b16q9Q3Gk4A0sRwD42NU/EUymvSbD4tHQEatcFin1fSGb9/kV
6OCBOcXg20rvyGw8QrvKu+W0ti62lqb8cYPAzfMXkTT876WiN578XLe8ps45xNzgaV3kUcLsQgY1
VjiQAV9VBGC+smS/gc/g4iiZoVcnqJqRZWZ6ceaDaore+r2Il3Jsgh1KLH0pTe7jgMRU8GSz6n7j
LBHm043MmukiRKVqKhAjjkKsJnxBMYY+q0Rmvhp+H56TfIwzQtQsLd8mmtd1hsxmj3h+dRlr73Qv
jKwsxxK9ON1R3RVJ9D5VLeLues6u1dA+i6F+14Fct+sgAXrFSWQZFoeNhGVjcumx/woNEp0iXq4J
+5k03feWZ1z0Cu8A16k+BtmLJgt9ONIK0+D3TPjkhZxXbcHfqm0saWURfu6N/VverHyzWz11Bni+
TtBjFBVfV6/iJ6+o/K2i8PpyRQxtcC4XIfDgl/1ZyG6XtzFg2c+sVkODABiX8+vRyb49CwIBBMTp
2gBLTbDpvlATgcZcyf8R1wkqAaTMGy4VlkMaAEeL3lLqttyhHJhZ3y+ad8ppqJuLbwDya8S6sEgT
YSXlf3HlQJoYAMcRTEAEJ3IEjK3Vv2OlTT0sKTGak698r/cVjGe17Ml+DSaep7bF4E6eYGcqvUwl
jVvEmBN6EDiFpVicyB4UF3hejIUFjeniRsvO1xBghE4zISlSK6/tl0+t8o7ZimM0mEyWKgLUsH0W
cts/ttUBWq+Dki2W9dfPiBSqs+8md1LSkLhtMUBfbsKj68tzxdTujCygnhq7W9kuZF+I//8YC4L1
IVHZ52hKFGtt6AArTjJCfVyE+lvFRVy7JJvUO50p7E2EIyVmTY68UtBXIHceIzF65ZAz1cZkTHj+
fQHDX1dyHrrrz/DlFg0ffJlK0X3Tt6zNBY1ByK8CsHpcgdpiGlk1RDZdts1AhkPCGhpZwA5Z3onD
JpqxyT6YLKlSS8/Te+1Ub3q1w7S92f4jzxwqbLBnTxAzl5xHsTSKK+QrbgSlJBClDpx3xQR0PiZ4
mOHgpDHBTwx2krzup0ENdmPh/vIXMRh0tqov9jFe4RmozrY+55/4TsIhRueOpvzSyF7C22fS5cje
AheiyLxs9e2nhZKhxuagpgUpf8F1NgAHaOrG4LMPspy2bhSKsl79453C6Rxi4Zo7s8I1Tl5Kna6K
ieUA/HEh0Yre/IHL/2DkiuaBm1JMCPUob4n+qnFNncfam/f7AnICLb/fnDpN6yPLjZ07FqEHmMaK
ekQ94IkNtWmJ73vogc0BJTarfdKJlbBuuOOZLmn7yTwjdlTiexrVVcKrer9iciTuuHGqm8z6ZIVW
O+c/c7V89zxWTM70toyWfDJHz8sYdmGuMd8BS9rCxS5WZKbJE8ZROBE595GD59bFcEGGdSYAZJ41
RpNn4M/fz69AAn8iPpoDI1g6ZSXM2DhdVSq7v5k+s2vSi9T9XtOAkvivpAYXkQIHcTOq8g3PIDc5
pJrSysKnpmbPHqBSjGYWsaF31pLOPlC9UQUhvrF9XxQeAhvspTtMaA3Lkm/KMPcbhc7AhfnomhZo
T/dQmrvWgWrxHj6Y9F5gda6yO6uHwdrS6vPRZ53P9PuBW/6RX84Wt+vUPf8G/dsXbkEO6pGb9AD8
nlApVZXDNYz0jBAYtz7tUddfRQRJfknbmVCdSqEneheavNXWMwCLivvNEisHU0MWiCrI76xuCCkF
NlTEjhATwAxhPn97maHV3BGdfk6+wco9VDYTtApp8dpkeLlDkAbdFVSLooxxUYgVx7P8amKk1fTk
UeLk9ySI4QzRHzlvRPzmFxPhLKEXjJGeziHliIZyuz16OwHMC8p4IbRYQGq/gyHkemEZT0iGLb8W
p6NsPoOC8Te+gqCrZQi3JJz2SrBEJbbvOfO/9djUCa+P+lD3AlBrXorY0ShbNMRA4LW1ELOXqAX/
H3aSgMtQhp3S24pekX02e6+jD9Aavx1zTdtN2r5dKunowYofRhtPtRujuxAB+bnwL6egDGEtucB9
rZnxhHZUjhprrZF9RZM6DzTNZkqFiWAK9W6NaesV1ozxfbO3KMl4UKFzhmEC2CGQ1dytVMgBW81x
cTMDsJi3uBXTp0d0dhix1TW6OLsfH0xM1N2Afloz+H0ZADIZ55Fg0AjI6jDy1Z6q8Qihp25YXkLI
PLCdm/v0xF/xlJGt4ZG6AXAbLLF+m/zYryQ6BYJBd7YBwwK8zoLPgGvfNM9nS/IyyKKO2Y6+T9WV
frzNlNynVTI0SCMnsLX5eEFdoMYpiLOLPdlzQS+l+U7JKMKDE0nvvybm+WXem0X+i+4wF2zX4ga1
GoHBDD3pq/U54aAONsOgWpSi04ePseqshfXEgCKUMG9IaSfsdBgkHCfsE8khOysXKnF3RYXGL1ti
ejrelGnHEoVKMjHymCTzApZe8C3Rzk51okhYcT6ZEw3lS1lljoNnIqmnh5gjHICHalXvEe7fUK+3
XbdKeL/UM8Rw9L+yB4PM+hqm9V6ZJD3yPfW7vWsHb0BAXbPPPxv/e8x5y6nIOFedXb9iXk9VTVF7
1Xg2yPYaNzRiSWCCptQNSopB/AHKpxBcjyYYj3ctIJyktL0Zw3/cHRvVJ+g9g4AAmHLgVVEbOL0g
raZw0SWuobRabk4jEDKh9gIGoU+LlvJcAVx/xYTOxNR1qlUgtN8PHEgtblXCnlY7LdKk2Lg3kDX6
GyFfGkfmrPBWjKMrydYQiqsB8N17kFPP8MsH3txcB1/BlOiRquyB1zkBIeKezt+79vX7jl4bVqbT
B87jzb3fV8S+nAEh8VUEbZXH10AoLBemu59j3sUZaferHJTWmJAa+E/RWnh35+DT6+D3kBg8/Zx5
lyRvqajJ7V85jqS83u18JYU69iDIOly06rpC53OauGPQlvNTUheCZtvzqDZ3SZLRRqSsdNbUkbI/
JHCtniVWoH9u8+8y3r37+FuoGu5UrgQKTFb1s0yZK7J1tn6KLXWvsAh/5BJstkcAR2F47sr1aJVD
lhMV/fuBRYPGrHGzKW6weVCR2HtH6zs9FK0DE1cBv4ae+YwhlZtXrGN0lK3IU2FTeFZxCVSa8J2B
EceyCH4zp8/PgQIVTsbrRNrwPpgAsGt6Yrfk09pJO+mh1BNt5Xw4mPHkcnx4diSQPCafG4sZ0sLa
6oJ+iLYVgPgwiz9Mb/7pPXm24sUglwgLRfkI6CeJEICYZHi5jp6B5AZV4J++rYVDt7T/PswNIy5T
UtOoB7rEseALt41qMEwb8mzStNK6GoE7WPzxjC+NwQMADdTKlOYc5DVnon1fXumMtJDWEHkrkCop
EUp9MrZqSH7AIMrG8ImZSGsqaN5+HnvSt/yZibHwsvTasYZQlfj3/nLMBTav5g2vtSVKPoyB27pg
APgFqpyTr4tLRxtphFnMPRARwVDTjLaFI0dKsnf1Bs8/uArN1mry9I8McmUmxFeuBNkP/j4e2g+Z
/thB20pZ7euaDz68ZHQ27AcGj846xQB9AKggT0lpF1hMK5I6oEOA6ako8dRR6yZZQ7fXIejvGVmd
eD5rrTBKgvkmjaMMul9hTCNPnvhNvKSQ3NXfmaKYZxvZ0Dy1JwPI4QK48kOBMvv2rCorrdEC8ev3
v1w/7u+6Bh90ADdQr5mhBofiT95M+h4B//Pv0VHmDhE4C0IhsBBEZSocinOprHh5PwIKJ7p+GpX2
4zCHR6RdWDWuMQoFbk+2fxsViFJ2L6BzkH+jsD/bpB1ERU5HTGJNzrmsF5YqiNPgd3DcD+lr5C+z
J0hJ1bka8upp8wx2+21oQEqamkZRoH+7Xf0VIVrgpDGzsCZDlMLy0sP1nbfcyq3jEwKPRgccZdCW
5hoMDEGNOM0yOAzafr0mrbGKKtquOTsdjAUs5W7mpSIAeA3nVb6kd1GV4Jbfc2RHoe52thR+g/k0
o9hGr3WUYAp4PngoqeTlKYfwu+i2s/BVf2zPHaQElGwl9LOnI2I7EqrLn0kNVh32X+jSgNy5B1ZT
z4OY3LNP/5nUcBEsIWZE+wYZx9uf260DW3lAEyPuZc4JON271wfhsbJt8EuuhwkR80KV4yJqz+lg
HeKQbeF0FYW3rSnU31WSzAEG0yvAbGifACDbFSbY/ZiVJqvitNZW5qMcnwK7/HoWR6an21kHOWSf
H1H+CzB7VLYegsZsAmF5QfEnGXYMu9qK2Ienp5bv2NtDg4UjI4ZBt/furUxjmX/FxXjG3U4hU81v
oEIqMu9hfVu0IxYY3ER+ZjWziksZ3d+zdWBBxFPFJYXz6pWCCVtImnftMCCC/x1gGc4ttF3kRwzg
2tf0GI5MKUHFHgXK/CrrIB6IFHnkub4Quo8+yZ/nDJ6zJf23y20eBEJtTAdr9srX48seuDRGA4yY
/iW1t0XWA4ooBQHOcIh/9orh1mQMgJbopUgXtlKToXeUpQkG/YopLKYQ2AxFTph6BfIaCeTZZRdH
8Z3kYWXIg9JtZKMjGJVilZEU1aBs11oOGp6OTFyq8Ci5iRRDQrAl3E2on5qShYEB9oFbTnW/+QnQ
/yAowTRGD1czZMp33X0p5P0TF7rFqQrOYmhEnLS7KI6zeKNlTXXPB7PYHYRwbVFLAROZ4PdVEXGB
pAbO4bG9uP84hooi7BRS4/0GxdskgEtwZUVA3t1Gb8eo0E9qABzG6l1Qy3xfjeALvfQsqp5+mtIj
ec0vN7OsPo+X2Ty4fWkdHSByJKFcuEvBpoyZLn2GGZrpQwBip3RqPQJ5sUAF5sQVAeOLzHjYpsmE
OgKAvOWiL36Id1MoGh5k0cATvYQ3qIKYC8qa9EkWmhP99du1gd+Jmnsn/Bg+XshaIwAprC/s23ni
3GpJJMXO2Cn6EzBT90Cki1vcKNXqySmFuMXoSp0sX67Lzx19w5pQReyLknPqAe7XN08RrgJ/81Nr
IpYyFXpkQlJQnZoovxD/dcX7K+8f1+RyMs0ZWzJNJ4ttKO+0wfnMvVwv2FohPIwyMo5jwA1iwJVk
WwSVjUqyUXJ3XkTdpNdZOSI6nk0OojFK9pOPGhuV3jQ7q6S9yznylQ30fp+LVH3SlLgLt57BFZW6
DU50Ig46FCf1p/tMtJ9E5Bj9jVgoYNtcXjyA1X2lgrEmCki3kSyxY4dYZYg/JtXqFiOiYzJnknwD
gN20ZonMhNrtsTg1kyy2wixpZOznTDF2rVf1IYsD5L2siWGSMMhqL6/kXj8KgYCh2p+fds8NfRo3
lYkihCzl7HnyC+tQJ4Befl8vhkToQFRY4RUkwNMeKyZIplhk8FUg4IlV1uiFLIH33XVM7Ut9JvMp
CrJhetvHDFTQstxuMKf5QqEbzVUFEpT1mtKj5WbqiCkD/9/6ToY2KFkEqdc/nDuob6pRXt73Xxab
s2Half9CRSX/Wf+awrbkQQdqGLe6W7WAZalk8hokgCajZe2ISzrOlMdoQhWiX80IoWEBvJtvQ9L0
gLAs8I3x/qUKnS93hZOm2dyBWs5xSGeOHxUBfsDP23B2k8l/YeZ/RC+LT7htUGbQ3yIjj2O5YJVv
Z3M3rEdhUfkspSCyCQip5fMlCvW1inlaOZ6CCPcPV9ukR7I+kh15MkU0MTrma/XLLhUD+eO1rw6x
8PrXONCuGrV62k37AycHbA3kdo+WT+wryxsQLphxkDKJJT3/atIJmIj9LZLCfWn+wwQ/a6R1HQZR
HAjU4d4u79OLqMbfCk5fbLIkPESLNDucwSma2GSUpWShf+zRme9e9NJ0CfPEnEEsHP8DFx99SH83
g/Kd+8FrhxoeU7XQMamdb1I7B1S+KWNBfsGBGopsuDYcx4CZ8Fin7vDjY7+fM2jtsX4cAvUggqiI
M3q9f6oOqIPsYP82XpV+IvkkMbXOYW9G0VT70N2hFPHwQUpPS1nleoSruQkhFNja7T/qFcfOmQry
pca2nLqEV9TU6esFVgQlcP4xoyfioIBOCvRHqTBGObvmwPh341pTTyCAQ9ymvKhf9voyMBu0JAAu
r4ceFTJBMF/nKoda29kA7Yrl0H/eA6rp8sc7j9xWcMm0KFNzDADoPK/CkR9oCy9jXry4joLLrWCZ
7zXByIROTHdVP6iOb9muZzCcadwR8wLRrOZ+h73Tek5O3mUV9OUNphBUmTfYZkJiKZGLNWzq8A5g
Q9wYaS2GyXOuZ1NfG4XnHyDkhZmo3cEKoK/trPazCQFbqoXdUvPRx8u/fjBIDOP4rpxXO7trh5kn
0+Nf2qDeTdLGuuTz5OarcyuZL9INh7VZSzPFLaTAXqpT551xsUOwhlsTDgcuy6enb/aUcD0qwIGT
ydpZR8OW+xQnDRDSb9bw1FX1SPNjRvFpObmH6e7xguXh3o35YFMdWzXni2IUHjHXW2P4nY1bTGlA
an0uSeOg4OOekiHXar1CUkvzO3IqRnJsH2kO3hceXlpCSvdWZrxbYotWDK7eVCUAVu5a8kRRQLiP
zAb9BNeOA9RLyJDDJk0gw7dJQdHMyiQfRu71EhNJnXvMndZFE+ZW2fek5sbBpYIXtOYEEzWtcjkC
hZbDJvxOyQWnBkx0wThS6Lt6qj6xZ8CqdfojwCLSNaP9yF3XO2qduZvLz5kn3KHBYLKRb1dfYiUM
Ij7V1fRNTr4+pLpDFic9rFn4YJhXPF4Ur64ILk1nawA6Fiza03zoWXZuWLpnkbAaB5ceuxtfZu/N
oKMnwkqMQLjH/c5ESCcKI6sITeGc0nanGzWwqINOUk/qD8zUUHAlv86zJ1JCtDDMTZcyw6iioa/E
O/YGD6s+AtB0RbXn6Q12sSF56jKMa+cOkBntyZYHpQ7rg0iyk0txzEmDiRPe31fY44dnfummyx/Z
jr4iZZzT+K9vUJbh/XmSpABTjDLUM0K2OSacMNy053amdDIfRCpgEjkIKNsAseDaATUtEON+5naG
EF/qK/oh0wV6VF/Vg7ByhjhLbzenYW81gNiVjIFG1wP0MWsPJ+tmDIYpcBpN+cKoIgoLIfolMWLv
voKhyxlg3wFEwx+o+65FYsIyS0E2A4nA7kPksX5oH82IiZ3EP2e/NwSYJRDx0eOEdMF/0dWnQskJ
1YyOfwrB2fmE/CYw33ebfh3LpLK6YgFFvH8PCOeHsHB1iVxwUO4RnKWOEym74WwUkI574CPDgNhe
bamLBZgnarN7JrwFVt2UkgXqntPYEGdDkjK9gAvI/DPv71um5w/iVPsHKQa1Dw174V4oyrdnn3vg
PMwbzy0xql51FdgSJvOvnqX0DBOVzNShN7e72uqtWXJt3GaE8NDrprH7KyRNRd22qPMbGv00dJTz
DNwKKWNgM5bODjqbp+Ax92jfVejSjB5x+HDumg5yI83DimAMvl+L3TB7YfgsxaYb4TU+/Nqe3obc
joGU9p2+kLgIoO1jzHGFCS85uUXW6cWPi8ateDXZao5PTiGTKYtYjnqZxOo4MyRqZxVMjb9WYILU
2239g5q2kmQtfCHKcnduZtFoGPyK2r/bZB30cOUdZgva0WL/UCYSYCqFYs4zgKZmP21LUIvdyUG/
MkRElmKADzehOsPPXJmhFWNmFsO1WQc8eU+i6EAKZjrkYF/wg8J8CDH5enMWcB0mapU8gp1svNGC
wl8pbs47jSu3D7F8z74mfk/5jCMAdFFP9m3ZQACIIESu2vPAbSR/nfTnQF4mfnQ2EJnfxAs5Cn8X
dultGMrMQ20kleUuz5iVxKXqToWsk/s6a6ppwwKVeoGG2IVcBe0IYRGSPgmcu6Go6YG2/RSxBRZO
Cc2muKgvtT930dunXiHIFNYp3LJ2RgzAAfxr+0NAUHt3JbIMrrO38ZAKedx491/jgFhaOprMz2AH
Rw6UKEo77AujQCblNO+yX7XI1OGvk4Rr6JBidkHWABrmoy2wBVIAhTCqiH7lfwAoN3uJx8lBKJlt
PmgmRpAttub2F3mkDABJFdt7ddPxv55nGKi1Hl8irIKrpqJLsaRkJ1RKQfnoVQHJCeo6ePWShfMa
u1eAvRUwYGVFPx/xmQQ+5hlXvRMuAWMJ3QDy5Rfut5zmiYEG3ZMfMPbITqdMqJS3iBr0T+0pZLus
7I2lnes26zQ9hIqYsEurTnjRz0UXaewi3qD+Agh5PbNfRIqYwErV0M+qM0tWbvwaaoTG4qddUa25
FE71QrWqxnNrIoMqrf6393uznw3bhOGT2jsII4T0hOxOjhhHsOr/Ttw3LbwiFcq4vA8Ivi5IFFbs
E6OOp4qnn7baZneDQJQsZc3nkKcLSyTlly6jG2gdppembwmb/VLn2bt+rMp8Q2cai11QkgJav1eB
SZEmTG+KEqeH7NWYmMHfnBH3YWBKUqeieveUV7YmvhkDcgc3cK3STF2EQ2PQs0iK9JT9SKDOd+/4
AZ8CyNbqet+zQ/snpy+PEeO5frVrP6DON0RHD8w9Nf96t1WTLQ4LqOFeapoAx4qduaYuB1JlcxpB
ZBv7nmObGOzy3tQx1BCFFyJjEDz4hmJ5/3A535h3ryCoSoG6TtB/4xbDzrYMKV1K1doRj4Nmn47w
Xsn2Dsvk9lSZahkbwFpwwQwBzXTbM7oh+Vmwl7sVYGm2o6Pz970tX9dTW2c7Rpi5J0nyFNBQ+Vtp
9rkgPozdWjEMeAwrDgviUPUZ/HhMsIZhEFt7C452yhW4jw+97QNF+0E39v5JSpUeFMyjbAOYpmm6
FEv71d9NZT6ZJUYKA9Kq1duFo99vRf7R5wCJdEO62k1oyx501SD52yDjqrHzj81CJdn0RcHoofQA
eIClNPIxER6GY7nozReMDs1DXa+lksGTYOR50zeyn/tGf59ct1H1sgsJ5UBgn4GMfiVmaxhk0xTl
hIYJFl2LeydzpLh393O2oGAxzWYvNKAiX3b9l/u105HIeEY7d6CCjISywa4+4VJUjr6qeefmh0k/
aaypBzIFXPGmJZEcBF47mccfO/3RP+6+fcGX4PyqSva3/2qTG12+w+2vOz4bD1otQmXcTgaK7b3j
JFmRm8pjjnrJLdSLm4qWOPx28Av79IYffoWaGKARXkuqqevuZ5B5STU1i/koljO0mGgTx9H7guIy
QK5XIhPaoVjvWSs69NJA/8rzYBsc9GeyD/vANCPP07RBV/1afkPkXxb0CqtiwYKe6odOiAtLM/Ir
BzOcB2b3NfS37VRvJxY2eDPZzH7KhsJo3kMF0VR10aaUlokAQOdyI7bSRN98wVJjvOaLnuwkNPdJ
/SJ3uG54YsCtmzSEH0BOsRNeBaRDeaJIvCSelrStP+NuH4+NQzFKkWkzhhrpgae/SgoBwZQtY52p
oDYWCyTzYxXjZ8k5/RlzEtWOZfU3MB2bQfzP6sY/QICiBfPc6VmXUwiR8o2tivCgcMmjvdfaYHO+
C4d7ZfUzVWPpwbQUS42dmQofwzC+oT5OewQ2Bmg6I5Km2L4YgpUSotIz5js1hgv2LgerI137ajyl
tNcRCLsIbatnZaVZngtWDom0jsQ5TjsBCnJevTMpomBlZdpRc21TxbdpeJCaIYtik2NddPBQj5G6
/qhBgud1fL5IAZs8MDojuy+xqLlMmqrY9Ut3bhO12dMIaPy9DFat7cQLOqdkaSKiCmMdm+h/hsHK
CFPzKMIHZCMMXyzT35wuj7zZmKMV+R9BjCHbhZEXfw9EjEB29wgQpaA96NOS3bwUyWaF9A53VB2x
Rkwv5kul2NNf2CV843U4hXauGAiyHp/EezTH7WM/UPmXBJtG4Sy3hx9aU8v9dJzyeYMhpMhnvKmn
S5ZVyh/Y9Ki6yPSd0tZ923gdiFu01honsRlRl0A9B+cOhxXyAlkrhHpViPA7aMroMOpv6iidZRcw
/Ch8EhLXQslZDx86arb0RrYUqLltoU3GvjpVQdtuiJs6JBL/y20dmsekJS7YW7gA6Z0EtiewU6LJ
tQqLLXv73GmjanDNmvdF3YXz2K5pIarEUOWhwKD7TXdynv1P+giIt151ddMnIziYQmVOPlsRJFjU
GgQ7QU7qHAmPJdBIqVWshCdmAWd1KMWXPiYr/+SdgUufpXX6yvBcuGIaemxgHpBfGBqmrp6jwS1y
1uaWEWlq39ArZp2tgLfvu/gbMvD4DKKxQThzOroIXqk0oTRNY33Yg3QT2LHmYXqkO9Nh89PB7AFv
4PqQ9Q5DpVmJPvoY52zQLk13BSImNsy9BeiDCndBTSDKT5/QrDUKykZAn6bs5SiFcHlQ+u8aHkg8
QgJdxqqLOdomxHNDavL1P0UoB/Wn0KB88eXgUdKVvfTc2U1n6UZY0WDs5p5lRjjmezEWG1ViH/09
GIHD7dfiwK9TlhoPZckPHsmXTelY4AUYU9gj9tbqpvzbF1odmAqrY4rhTErX0wC602Vc/lsHesA+
M3K4ZgnSBCrG9YmOHTNHYbNlWpUaVbK4fSyDB2bB7/9N9xrF/nZstxCYM4fe7fzUM1YQ5LmcyoTa
8azsyyV9IxSpP06xhU9H6KUj8Mxfo7LVt10FlzK6RrhBCs+tvtdQP4YPuGxajetJDu/xbcxaYQPB
MgN9okMVrAcgR9tSIste90dEoo7XcKrKPp0jaEBRW96TOBI+f0LEZAbNRtIyQhuA/11/w6s41UVP
fgYVyoAw24KOAYf8evpH/KsVxXNC6pCq5ouxNZU3yHBpBAVZTCjXeyNGSx61I+smFn7tLWsehJFo
R8MkOyqp2lCdrdkMjBLRrfwgDa6iHytOnzgfyuK6Vab38lrYYi/uWQWKulx5hynkiPy5KpRUOXzr
5c8kZHTTlP5lQNcatj9iA09lVnLGodpPNCRHsfD/jlG6+suLUewVGn9W0cNAYLKTCi6ZTl+QaXpp
NFv+2dgjlu3z0lrOEazdIXQ0KEZtuExaqX7TZh34PXdc1xmeM/Smpq8V3pSG6SKhE79EbyXz9d5O
p+NWi9IJlCgXoAfUuzMRvA2V/n/Sj/4jvaziTSKn82dhVcfBbomHT35/76bbcG2w1mEJ99rl7IAg
IRiWUdkVYhoGafik0ivKdX13gO4K9RIT04u/yzCyf0nYuTNea5R+B41mmaM9LywsR4fGSBE8mUT4
eRKrk9YaihUx+t9zzLmrzH2DoOfaefQqcD4ZQVtTurfVzfjch5QDnor0zbGQs4A6WB0BWMEkmx/k
Qws7UcQf9KzyRkbZZxV14G5nWzoX+HEy9AAjy05jFDtd1D0Zjku1dpSX46NivPY/3ugyMrlvOliO
YRXShiRJLahA2wh+siKiNriaatjx2I0s3IPRGQa76rVKS0MknvZBcKJWTN9UowNvRWEtdxdt04mZ
HE87maFbqoT+rhXQ6IYTB7N5nU4lGAYmqrYwQjrQfJV6GCqkHjbggR9iwRoXg90acH+/7C6JRUnH
PuwpkoZq305S8LbQ+RNtBmkM39UqDJCHGl4x1A582rnM3TtIAA+pq+WJXFjyiXyYJv/VFJDINKT+
pPCqLY0mlnv3exR9irFGjfIQockcTY951WF4b6Z+4ARJtoL3Mw9VYAisc9R07ZHiig3lr7gEElA+
hf5By9QqEsk/Ok1rP3kn11g5sCO9AoV5nUC1XjXbPWsbj7Vus1fGlabUCJLPs4NOL14AMhXP5b12
gLZmAWSvdCRRGqfTkVs47aj35pf9vJS8BnZgw0sIslbqKKGc4JSwB9eJyQNVpQkhPRFrtAerZkCg
ONfv7YX5bOIOpO8ofp9b8Row3sg3cGWw6lwfzlk5KPjywBM1Li7mn360vK7bxbxo8GYqFWUYauMy
5y0/+tuDpI2OreLHrhFS3QIgFNcW9D+HFDJCTXGWjIz23RpuzRKKtmxGWgu8LwvXCaJfj9QBwKef
Fo+7DZHLljLlrlUAwugmHmAeAzTK6r8CqyiGXQ83k/pai4iz9ZRh7CnE44m8/gMrTFS894yxZ9vD
h57+LZT2UidnZR7U7IJ8mY2NrWOOZDxK7VBvB0R7GncL4LrTgYH2W3RfXIxCKSGZ9izHazVpVkp4
xtVVxI0+X9CfvjRAVD5oQIFPXfUIyipPFD6cQNBtdl/2oBJvyedoqZMRC/xUpOK1N23svxHHTGDa
lFnMFXBX/NSbNOxXE7FmkahMO2mJjlJrwaersFga0oyYA250EFS+W/esV+1aF4ZvDXkkaZFo3OIG
mwKXOPFC2wiuS7h6r2oIyJLs3mdE4NUmzwG5Y3BV4qhU0oMqmHrpG5jYtQwyaG9wZdUcaMHf4a8k
T5MZE7rjenkycVsCqFGFDjg1u73baYmSrT4QQhlHQtVb3wiLWqRSaOGjQ75yxlRTtxD557teR/LJ
U1Ew1xDqk12fxIRdwOG9foSlIUF3SJHGFzofo3+60mAZjtZgkjspHjUORO8wdh10FtQ3RWVUGjWp
jfdNtcEcCaPB07+xmyxrGVtDi+R7tX37Jgs/TABX2HAV/AjePRERRSR3icSSMQOBh4GLi8MV+oSg
preZ/Ab+kRNdOA/cwOFrasE/SW863mXuJSwU3c04nkH9mVKkRiP5M17u8wWbK9APg2Nc+liu9A65
4PC3AFIcu8ea36VlQbJT3jvPRvxJOTrYBZhRLy6qgl5R38gZB2VfftIkjpanGyDk0OO4cqgLIZa2
Se6+RASpA1nptbOolwbcAQNrhjEmHnLsf6js4568ZyNbt1anqb+qyFLH8AnN8iOCtqAPK8TMww+m
in41m4sFRNY6LvCxzPsbZS4nD3vaLu97DXRpbnqZq25zYG31rJoqi5SKXiKD9L4HtQmu8oPihL5D
XeGfIAEs8vSxZCTy8Axuc8Nlv9c3m0cHc0Rsq4a/kTigYF1huVOi8gu9jIc0foTpYMlJm6c311Fh
C9taqrHMqR8o3eZujLsnVWlI1atBzk1Mr6ROTrK0VleAIi1nwCZq++bo+iJbO3+NI3N89x5DIPGS
suLeqR0jDgN3gLmy8B/icQu/iXmN9pcPF/C8wfbkcL7Xsw2jxOE2xeidrh4smFu98rOWWeJnM6ei
TLLRJ+pKkXsze1e+WNxErQjKFelFbklPh8ylYbeBnK3g5wr87QX8nQw0PwKtB043CKnkvghdigZz
Iu4Dv4I9o+XMoqQlQSeBlSqxrn2mVnJluPqBeAgEAkCGBBSaloQXkS24f8bK285UVqkqNumRA+LL
C4NV4z9tnDyk2zMJLAOmWKJ97Lv4E26bqkmz7F1F/HcvLk6Khvjb0suyfvKZEDGVppB7BRUclERf
OMVdvjKgeet93d9p8jnyAEU0ve0Fkh+hkoyVwi49ttu9SQA2tcuZbF1z8LLTR1626CEtMh0oZug1
qw/xtHWzf5ZOTG4QxIm7pyWnVC7W/60wHIp9/N1x9TsAWM+EFFK196FG0wSCySAdg2f+7WmdrKYi
M/kE5c28YuHC5UDYTymmpZ2UlB408K4irUAUd6QBIJ79PkrjAE/E9JcJqV7/MIfj2s5GUFbuW9Zf
To6UPknbQ6DzxurV4WqF9S/Cl0BcDBhWQTuBdorFlOFFk4Mvq0onMjlnRpgwgA7C9FvtvBHK5JLP
CEZ2rcr62Aibzkshr7R1OceoYPDDjKFht5u4DDpgdDodpeDpfwLvGg2HiA1AhikiolszUUivwOp1
Qu5g/RqBVmEg0oAUo73ZoN07aM1p2ABApADUXsshYBH7itghEoS1BrxU99wwaw/GZRJU4u1362NC
Ol8K7ynNUdH/jb08V3nF/JOniPOO+TekVdEpXPXMzYKNzwcrWTuIII7n4lv50n8m3maEpgAlNIBN
dDnUSYZ7dIBkHKcNaw1VgQf7ajyaDbOAog+IK0vbs79Otf3UPbg5ZslzmdysStmgKzTp0jNbh5y3
Kaxz7GjWn+T0wcCfH+tfkx+hUW9Ngf6zDNT4l4NHw+jl/u+nVP8jsH54IarX5lEJyURDOgb1eCzz
Z9GmsO3Ok96sLWMxX2qg2XbhdtlnXreeHMF3U+4MIrakawEfOFKA5pBJg0zy+TSiH7hW0Msmjutx
OmPoUoTCmUqCYX0kZPs6IK3TbIhL+YZUzj7SlLePoPMQpBVPZaoRrcG6XCu4ff53zfKdh/pa7J0D
ccg/jDXlPfvfLyetpvCAVBnDfRyieWphslm/9WlFJo50mVhhsGKFqKpLhZ6t0C/E+zBw3LCgUlBd
na3CCWrnUEExJGRjO3AWgxqQ/YpQAisIwChl5eyr665pZ9D3fGvOTw3w8eo0Kv586As6Tv4E8SA4
0E4tVsTn226TmZXhyhKz4krD6YwzLs1ZTmRHhGjjoLnBu4pQvJ5etqWaQ++FI3IHA+IiZ2LE3Q8S
auDCdpKwERmAj7vES9GUD9xNlMUe67PEE7oLM2WsQQy0eLVL12zSEFiiw5TR8jq/Eb/peDMt8NUv
vF9bGbNzQ9q95Ak5gFVWdqKWGAANqU6A6aTqwTKAHcLTCMEPZ8bjo+L3UXTjtf7aFx31lcLouJ2B
EJ4Ur3yUlMIM6IcrCCb3ZKds8RYqXFBpaZ+ODDZUYfetmWhKiMXUANZwNWMPoPw+vUmBcT2AxqL9
homiG2p8wBKQN3he0gs6/UmqhAA01lM7twxqCkuqqbxY2aRniteEIummepH0joYwulG9UfrMpLKG
xK53Um3viDP0gatmfaAw7iECVuvyo+OrLbvOSY5s4xGo2ZY+rpPVl+13DWBnuiJrfnEqBJOysW0z
DqQQBSJriB2JRktG2e7YYaAxl0UyXDUA9g0B64n78xendI2A5FA1lbPCiEkeLjW0SfxmJKf4nfJI
pZsZPuGWCKPcn7VaI7h9MtH8PmmSFTK+ytbBza/4eP+v62c9dhWadQq066DUED9YBsXJ9fL57g4A
4CYlZA6QPm4tGAGEOQ5zEbnJ5jzep/Z5bS3srif7IY+6xrJMms8y5vASsxst0FVHVJkjpNHuXKTO
5/0+8S+wytV8U2G0P7pmWDBEBuQneTc8anYHoxpWeiso3la/P89qhXMwePHskiBLzOk/FL8Qml25
faq4+eZcdXJ0yD7LSaxiFpicehtk4IIX+KStqDjJSbMUGAUWMyY5uKDpLy2Mnwt7QohNQSDtspA5
suzE5Vyx1E2H+SSnL5lmdfbcO+M1AgrQFuwmrWi86RMNBNbY6efCYwazxXp60gMmGIvOXnQwnRnz
iSgEXog6nG/9U3QBEpgqGH/hqmIPf3715DxP7+UVeJxjiz5CC4LN2I1CLt719jFNmuSlb2wJ2KRC
FjtIRFziJbvTHnW0rZuoeIwGdBZ9buXGnd6475JTiW+iwjSnH8xegsOSOcquZLwpP5s3PDPQmRcZ
EKLs+BYRBvLwxBCcD5NKcgtSKZMEWTUEAfdGFVtu6MWn0oOFnW2nIcjW9wXa/C90Rgh9fqFuD1cf
ENMS+zYozA1evQ62chq11MNNB5eEPYVLwLSTRGlUYJauoV2mZsqORkKamEE5CvDfoZPNbEJ4GsS0
aZSJd6dHj5AWyNeFqmPRZVX2sL6t+pkLNfNaoC1HtZtEK14/e2svNKDbiP/3xME6VBTBMKoblhr1
YHvNey4ClPQOzLCdz1JbVWt0JI3vI9UYoGggJTBGhxarUBIm0N3rU65qJp+kSoGURt8nOc7+incD
51uxQgUnhWq4L1yagMXPF/pK4CeqnERpWfobVtjcmF+bR1RPwxq3NJpRUrqsYAKP6tZRC5ZFg+oq
RVLUf4jIFZogaVXjuQB6kahLuV7jNNHXMJU3XD3n7TbNwcNm9aBu51f1rmair1tlz+ELPEI8xxf9
fLQn/a7M0ocBPqy1AngRemMLp46ibOGqPEQsQk9YOWmAqvfPaAlE0oIcdUulR2dMcswphzgm9qm8
QIHhmGLd40nYlPd875Drkol3Ij8DgsVtooZiVsYxO9G38U+jaC9tVtFphFxlmfnOax9B7yjePanA
bI36uvCFX9Xe4qttIEM8HGMEnr+jocCa0amQWzF0wG6pFfMOfwbOE6gco9DkoBlAAXeg+fmhvd22
0BUf+8nhuWsl4WBk8iIiMkg0NWEJYc/g2XTYg4yjyHiyfWGn0DSoIdbFh0aYGZ3AjtD/OHWgslOD
/Bp4TzY+HgXYRQFXNPDbVluAGvXw0CVoEHpRC64+BWGy2t0XHvFfyXH7h/BenX/xaMJ4DJfs3yx/
/F7OaReyWUTwYbvr+inaq8LJeLMNjvm/l9N9BbpqhulaRDY/zPgOCkQ/1XGXGA2CC2MFyW9mgmL1
KYEY/WuNKrm32+E4DXYmkC+ej2LI/PTFv76Oxn8uwYx0/O4jU9i/wAPT8onmAacRWS6j6hzGpSB4
UicNdvfp/74ptcE+Hnxo1lSntt8Gtp+0MbcoOQsJrgNo4EXYMzByUiPvn/zR8VGLJ3C75qN0Wben
doFFtya3xvsektuF2HIqUwcV6bbjsOhtt5XKDH9VlaknILGyGR07MUviSzsAGCiSgDuNxkJDeEB3
FQwF8tGWVcZa7MDDjVyzPish/TrW/l+hOhtQaAEPdeuD8sz1P6riSc7veZki7EQf7uzGvlJTSH34
IgelV7BvVi3bo1lUOCmLsQEDXaGRztR9DR6zgWmqS5tURnQu/gnrUbYRFZM9MpypQAuwPtN6m47j
IcD1xpaW2twQ0mdS33+TFZhIltSPGN/gYxZCG3nm+rLae8x/N79X3ey/fNAhjWwniZ8lVVzIIzGQ
Jxyt/KRLVoIkuWKX0xEcMdnNCfZ2UGT/hn+7De72LgT/cnQ+xGBgXk+3b0rLKqTUG2fOTdC196MM
lKYkO2cPtWWr1a9Ucez3wNrIKyLOYqVhgIfNBGFb01sqih84+Wi+9sL0zJsz/MZM0mvpVcAZHQc4
6YevEtC17Y0hm1fgYtWa9VwdkAz8KRfprsf9LzojlzC4Zpy0MUtojD33XSEiSeNTf/BNpRKrhgBQ
e3unjrw1qAhn4apvmPdzX51ypaEZKDKXSQZfgzPN5UZVZEznE5qx8SO87sG1sAgEcNwV7sPIHkvP
tnVbWkShLLcMh8ET1cau8ccrWkevcTYM0ASmfhmgK7P8UefCIb+w9n5vpEyaKaEnIH3rhGep2zHJ
sVklmPCe3Dg3KazgLYbcrHrsVFKYLWkcYKoCZaMLkV1dLh5vI9B0hzz2oEwFdjOprEYSsBvH5e/y
SuHqe+0oaVZjkBxHgDeVnjDi9Qs4gUVbQBVc/4Nv2CYWNDZOCLUa6q0/b/33QJk+VhmfiXlUnd4E
wNmlQZ4dALVxM8M1hsgA6SYXrttKcdLxG9Qu7OhLs6o0L1q1MJi20SZ4k7p27x/O5FevdLUSByGP
rBL7UWLPpQrqftwFai0pQNxcrp6LkgI7M5muyLl/EJd7I6jih/ymez79JS/8S5r26ZTcGgt/PeFV
pi6dO4v2a1QBcA/fNp9h+3i2hTU4Hct83GJOepseTMsALG5Hvs6PMoqy/VP5Mi2nnPxVOcsu492/
u5l1tP8VOuPB6/oIRFdPOTQWgv/XBM4OVHSf1MMcGoojU3zX0BRJbl5UNvxGyHIY8O7GolhGVayL
VLnajrTmwfHjjl2gdzC8a9z2fk+mbM3HBsd1z5IyEvfavYkLspCr5HZbWDhX3oRL4YNx/x1IRgRg
JeYSx1yzVygRjHnTLFKooUdPRW4yMRL3gtV4CdB5dBnDi/VVPbgRJXNTldXVI4IIX0mtUhiFTQC9
UecaQxxJW461kA+e/glbt/ILAe/eadM256LX6N7DPNBgtpGQ7G4Pt4dKMg4O28MS/khR10c784pr
cBO0e5B+md8Zv/kCU02SRhWzA1P7QEn53rX4XO38GLF4ic4ak7K3JR7OrCqONXfY5GFrKoE1pFoq
RG5kkOeVuJpFFW3AMAYngPruYUACBUi+xs95XtKzfYtddxVuGAVrvzH6yu9WHUtg8S2/SRQQbHMi
oQ31b4VFesB5VcLNurB6NGN7zDdodBpV5TEYCfHsWHqfoMplisJ5oQ4tw7h3qNNOXXEOE70D83fu
5/DkopPsOyl3NbbS0RP665QNZMsnpLBpGUmd1X6bv4zIgGH8jEJCzyPRX7eYrnB+QB8A9Q6npzCd
9UCtQIM3Pv0Z1SVOFKPEMqlewLkHEedKYFT2CU7zVVeb2dqhSca4xPf57kFut6+X1GdXEZVYGpwx
DT7sN3gLuNqJGlm08lFSS8WWf8XJVTTVWcXoT+b4f91OWYtpNEwUiTVXHGGuTmcVXr8Tl9T9fB5T
yKtHfV5GJ+Ai9IEaZO2zY+Nzu/rZnRcnF2YL6wF1yeXsjJhpz98cwCeiavCaBgsCsaEkLjP4Gmnn
XX0XYuOduBcL0Ifv9nEhBQkFc8U3fb60aZ20cK8sVC/KP3JpLG8UoOsM2D2Pg5G0XjITrD+Y91jD
9xcgnQPCEwOaqkK5baWJHZKQJfbiEcRDKk63GEgkfXTkVxnvpqvW49Bnl9xfUhziJD0unAu9KFUa
TLW0KZNzfOoMc80feYnk+FuvOXDjxiXJEqIdEk48F5B2o2y7qhUy3/0Srthyf/t0GFH1LjoUln2b
oSAPhMCSbKKcWsqo6n3OrGFm43MEXcaUagf13ohDCWkBDrnOSpDCtHjefDyo63H/AcLm5oCKsU64
EcqMybp1fscXxta4+RHRmIrYZ3LlOOTpuTVth2t4whQ4zEpjwSEPrYbWCzRL9CQUd+zrffGDCAx5
ROmWYI0rNy+WsSJy2vKQMBadSlQ+DWFr5QSBqd1gdAjHNE5fo5UimJmSf15sw1Z3/1i/a7NFljNl
wa5W+5ZMNG2biZgGnwIR32W2E2dg8IRbN2HAufN6YjNAmm5vPCgGOWySoftLFFostdF4D8j4jFIR
B5/IapUcLLN+htf+J56KcdeHVTrQTjfINydyfxH+8keKSa1LjO6eDD6asH/SuV1OxqzLrhw5FhkP
Ylt12MF85mE1fKQP/RcUyGZZw0S1YIaJYfPR8kT9Jeqm+JYWFkMhbe6BK2HNxIKTMY2LiDNJRp7Z
wm+advyXeZKaY4PvGpgB4/5TKakplSkpuF7Z/rL+sQ6mjQXM52EOUV4fT7pN9djTVlzapFTvlIek
YB+ZFGY6rqiycVNEwWihJoZCiUOUwL0aU51m/j6YC7fjxEYDAstqbcpmiBDn2kjJdnUhkvUhoxvc
5UyFHO4Bja/++IsNDyHPH0MOdEJLuvRr526zK9dxf/xDtVAqWfF8oOba6v7DbMgHXz9JLWPVCOgr
rZ7zqbEXZ4LhOlgLllk5Wx+1fi3XJNlWiReMQf+grz7YA0l59Ul4DhEbxCplAnH047f4bVV2pZbj
ssKc6dIlAmxCH4qagyZiUOOEtx3m67NB0zcXUAOIq/Wcdns/vZJAHnyAmlaNx835LTdKqeVfReC4
laK1zb+nRuH9vGtydMjBWP6SBkpEMSKchrRel3ypd7ryybgXc2qvVjLhvtfAcY8q0fr3lU5Sgqxn
xD8UDTG2Efx57/Q/cClr9p+kcIJ4Ly0HREdbMqKsZ4GbgkIO2NhE4rEVCenfIAq6jssk1+CiqeEm
MsOzcS+jmllVUb4Pt2BAYr1+d3KIZkaajH9qupkx97qtLMZlBxxEbD+db2xFKuvm07oYDl9hjMfV
0kPBOHtXTe6N6Qc2P6BqTAcmkQbFcrd39KyjLXvQwbuthTvf42d6Own1AnshU0lwa8vxloGHdGJx
7JOXgyebzCKHVMPStebNVm8C8AGIMkfvjXnjumH6u7/WZEX5AFblcY5rI/0lC/4/jLa1kN2WkMpL
qhurOMdT2AZGKd1Bxtrc7dHONBlJ1DaXGpOSCsoUfbbiASUaEA+D4U2Uv73z0SuRrrDZ1Urmie5u
e8nNRZYiJdgnYZcvQ2r+CnvK5t5fgIOhOAhWPUi8Zxxy1WOy62BQgafztbQnFCZgpO5dstLIAGBi
b64aemRmkYnTClbvbOwbEoZPURRAbDPv0Q4xHT58E8ICxrUqLJta/NL6SXcvC31cGpPW6mcoVDe/
ie9uzzhaTzU0/D+kkdBWs926PadXRWczKbo1Xjn1083iKQpnRh2ycmNJ8LQj4RkuKj9HXOUH2v9m
ccV0kdXq5nQwv0yw24oShov778ZikxcfucdTKQZCxt84w3C+2cdu3WSggGkAGjvTQpx6OBvEUf3u
FArcFnOa2blwLnPz5P23bOMmMP4MbCurzpj+pj3qTISnH9No+7ZPrndst+GRrrUoNikRdJqLLVay
u0Mmaro/ldXdKjSWtW8x7so3Smj0DJuGqvqz9wmxqbA8Wm2WILQbhlPqupA2vvkKWiLEOFsxLdeX
x0eYc4ZQyxlgW3RC9sTJaI4B8NLMrNm32xA5JB0wKvrM4WYxL4mDq9gas0NqxGFMKey+hNHtu33A
NjPTdvuegJItV7g8R6LarX/yePpoUJm05binNcq6iT9+bb5ELEcn9hLZB7TwAlcSodteke2Zi373
ukS3afg9L2ZFR1RvE0U5jprSb4VzgjdGhhKVhlTZGceNAACqAH7Sz08cO7OYMT1FuaBlM26e/8Ke
NtRqRSlxuShmPmMz3SDaxjBzIgI07NebCv407gAG6tXNVa20sx3/3qjv8YoKmqO4uKGHWsaJK+HG
wLdXIXiO8Pnowfre65sgTjnZIh9dgnzehxklxkWw2xYn6DGaRjTwg/Whuy9DZnzrGQC7GFh19PbR
nR0QJxG4uzvahuRNg0AWCjBN20VvSbW7IRnhVyr7qKmY5jigV77u0hOQVxlwqkv9uRp5lPWFT1fm
3hVc6j1d3L0qd5T/T4q1l6gQJIUspNMluRMafTLbzz+OV09kyisvfh5WKYp7nErHpNMnTRJW9PhE
nw2DkqI7AaIX8cD77wu8C3wfVBQdeGdm6XT+ZHu/IX7kp2GHvM1OU1kF0DBv+wQno/jTgA74ChHW
bbgZs6EbHA7i20lL8J2XdMcZJMzkDgBj26UmC156iHAPPVNK5dCtszpvkzj6ngDUgmfHfolrTzbN
bVvGms0a2jhiRtMk1OolDGPFGPM11c8x6u20uiTf2uXVEuxz5KDub5UGCba4fou5cS1UL9WYI+qS
ipU/cbV6z80fygateZhoG9CH5+Ag1FjpGKMsz2ftQTir4rFVw5fhsPz5+6GKCVl4HrcrJljqfMF1
lAMmWF2QmiFNQK0tjvLgEb+jZKIVRSvwDqcKyxWa4HpEZ7yunwQ3QKeA8mLccE7JjiQscF+T+vk3
OPIJwr6j94vsP6/iTzwcZhsuPEAIjv/U2/jhvQTjxEWULokVc/L2hSYvqi/3puyU/j/OF5MRN5GH
r9El4MJRTeD6ZhEOTQ8x+hdSnle5DnND1j+KHYKCNMLhbnoPN+YVf+KyDuSmCh+jdvy+PQ8BUNa/
ZLGDNQGDVyErTp06JirEUcTfy9ODJWzGBiGUv/C1nxgcZWU06gCoafETi0moTpayl7g5Ap9rKCcP
VjHdFM6n5Ahvfs0e6N5pr+Pt9FZeNJeAJoI1iQrkB7e3RBCfHGdj24aVVJ6W/sjqoUUf6SDbwnJB
iN0a0fIhZ3LdwecJanGztJXo45Gw8SPaZKrHWQNHbuw55a1cJHyuQ5dGTXLt6WVT6eoWsvTAUZpC
1BcmQ2LAd6YMGewYHfz6klNfWWm6qbyK/Kzpn/H3KvimlfACMKPpyw/OCBRz1IBwRB0RJHbqRwHu
TxLqEnpPY0zRdwP5ckstA4jiHUY5sTfxg0oQBo1Wk3yktZbPCRbc/6YPlRWyPq28F0JjzqiAtyzH
Ahtzp/a6sNmkxtiaLcsLBpcExOP7DSfL+nO2txAEJ9SAnsewLSd9Gu7U/Vm47cPntzZAs9xxKF73
NQj8YH8TWBbggTAaHpeoSa1AmQTCQ3xky5KrGego7VkhuAZyvBjVqPKXJny8XIG6RkbrRi3BgSgO
yf9UoPAc4HH0ylIM+DZFris7O/zTw8ojPR0whMK9mXoTAyVXoKT3+75Q2DXAsA5NbsVIiLynnV+t
MUnJhhq4oW73gtwTTP5zdHsSlM0eryJ4DhrHmEsBsWV0/HmZFzzmC58RTHw86nGihHWY6Zl0u0gj
VrYp7UAEDjLQis3y51P00L/BjbXoPk+nhV3SZL/tfu5tJRv0DfHWbPWxpNzVYIX00PbRWLUsiv0+
E1ddF9B/ODdBGPPEX11wC40Sa/AYrOTDb6HyZQ6ixhwwB3l9UM6PB9ZgdOnQrxrK8FRohbS7ur0k
xRPxbKbNpvVvhzWo/Cpi7Hm55eLhj0BkMvwlls044I1Kc4g5AD3aGFW4nj5gRHW6WybIChZVV9Pt
KmztWSvs0VFzXwiYzrPfSusTbgzO+3oSkFGAmIOlla5aIAGJTNruDPxAf85qznZLAptCgB8GqwM6
y7rD8+abS0V96Vpolji6HtUCmlP7gV6/NFf7UsiXx8NJAL3yVJqPfGra/NnXOEPnt+mx6wKVGkVr
JAgT/26YKWf82GJ8465I3avqYt0sDmzRtlDZiHDX0fPTKGfjgdPlXTG2syxsM4QGhbnsxG2AR5GE
+OPrQNtUE13kDBcjcOi9mVKjBBE3XIgcWlrJxwBHZLTxXZHVH3cPKlBH0tf6Fy5SyteW4ZELj2m8
Z1QOdJNdbgkJLw/01mws5pHBoqLDCEnLM646A+hVaFtXxKV+6fU4bQuQ1BSbQS3mqUOWEnqT4/q+
1YjYD4B+tp7wFybU+wBpN1ENe4DrXWO2znI/Z2WsAvoqrBPp7sXqGYuNPhKDHW2Ia/382KeVzLG2
/ayii6dWj48TEhqSNulj4wIjFtBLjf+mi9MHJQ1Bi7o8u0Re/K11q+bvJjbD+mYD2oMAR4kDBODr
PJk0fgxdLUjGx7cKEcmqBxyV3PT5y6sgdumI1neB50HgvFRg1fbKbV/+zaJ/sOnGojVx0ahu4FlS
bwuLJHigCfQGthd2MNIojo6ugQZk0hNlDWrps3PnBiruSMlHN3f6l3yrGqwxeYwoDym5tTkQA5Ip
mTkgk6AKpzwvZzL8YBY3vxpAXyJ3xfnDmM/lNyAz9gvZZ7YHQaDp7k1Lxe0s7f4MQz4doQV/hdlM
+Lzj7mr636eUsQU5zlOW1zp+ovSR/Sa5ks139/Zh7DYl0cSGjSatF7voyeZ5KHPSOeBHjuzdVTy9
GyEZNPcORc7pMq8zT7I3T8+Uwu+fBDGOxXFdno5Mh1afktrlnFfej3WlpNNsuyPieAPyZyIog7P/
PVBIeoutHK+xkuKII3r+roBG7oxHHgop6aislpQOPQpP1jubgxq8KvV1Ei4340wAZUdE3w5NvLTG
zKUv+ag7RelBWNfTtQGvl+E9Quh8iC2jC1WM32Kq0kwQpuTzxvW3kRuoiymByRR1REMfZd7y3v2R
W49TH/0k1AmWL1hI1iawCbiRFp7PAcXGZ3witKLtoVgIQPs0xo5PV9oVqZXugmtnYaW9L2n7YSqM
V63aKxP69YLpeEusJvptRt7tV+0flWFBnThI3c5DOWWM3JylLiaUwEpwwvP9oU2f2u96IZ9iUGkt
vXq1alIYIChLSoVmCDgLyNxD0VpOZGkTzU6EsvTcBBQf0YBZ84TYmL0Vl1Z+wsAka5lXDxycdIw7
EhGw2+64AmmZc9RLz0WiYUxpViEHZ7p/7J/f4j6DKIjUN3KRD9hrCCwtpJPP3c2+OOxuj7kchaai
u0MXW9sNQAnDxYjiYL9hjN68lubJmn0lOwtqTraAjWy9uoKFyca1y72qxVRT013yRxglxR/7V0eT
xnVu3p627+yWw/odyDQLvE5Q4GbWS0XsTYpyJHLrPu4vJQ3d1S47ngWDWeqimMqh7/FoS0GNUKvt
1FcT/expUqD8x1RrPGEQP/eg/LCTFIXc7Due3+cOIBQ7eeQ5MYdCrNn4B9vIsRJUmTBUqS7SrtBq
/7teAh4tyyZJ3ulprEpaFFNbML3kV+WK0GrFNR19g+n5QwlBBcEfniJKai2PlDScADxwZ8lQLf8u
xLWS0c3gwwDz+itxKQrJMD8MCk/VI+w132HEnbZpf/sanUE8ZMiO7ljNBp/2ohWUr2GPvW0TPzhE
5+i8p9ws7JkTg/q9klIM36KLWlZvy/NBJMVZKGF1U1wm3YOKwZmowBJ9iGCvy72J4z57P6XNuF5/
zqWA+HApiepAC7K8283eeQsoBBMrnmE2Rpf7CajE13s9HXfHQGJYVgq1H7VijNUY61hZAxb5/ZUY
x3nOfINA0BYY5QC24bAPH96nLzV4rVm6JB659p+nBacPYF+DNOfeyzYKEdEQel73zrjC76vsjKVM
r1xH8Ht4EQpyCiBh7Vvz0fv4vxZAsWTAcYLsvQB4yGPtA/yre4gW+EiILHO3J9NbZItwoRmkV/no
jArIabQBwfgu/6UXt/v5vVVxCSPZu6x1bc12Su2zs89w7DbJf16XcAsGHynBcXjWIrZQFJMtGjbn
MfF5ZbhLu0z00E/S6z+0L5SaVX/EzaDNNLqKY5uPvv1zemIL+shaLzhBa+VpPcNsP6N83NWAgsAq
UMfi0k2/+bmzSSldFDi1bsHinOs5O2/9I3QPWIPPabJ7QUv8akmjub6ycVMhp0TvphGE7PUbtsEc
FiY3dSppoHpZ2NKlWz3hDWKwAL+f8LRfduaPe1fP/tRRAI5qy39kghc5A4PqEYt0Tpse6E+ct1L6
LdpyWu9GLNzjtJ9CvqM4JNJPdvmc0hLXGP9FXjXyBQPTBDsip9yeExPt8ii6TUXGlGiVw4rIzxbv
UjU4Xv6wlGaW67SL/Nud72fWupZaZ/UU+Q62mzH/oHgUufvt2HglM7JMjFzjvQBcL5b9praxyuqZ
A0m3BKQT9QYkvdR4OHN9zdO8lDr0/HFShg3rrJ0TgKcBhulFRrQQRAK53dIdmjBcGYKjh0rTdEPK
OjC6XdOgMMYb5I808iQVGT5IKt1/1nQ9Z2ncvHjJPGhNBJ1AdGplqyy5k360ow02gahOB2IVD5Bz
wUxd7EJr3yL++egnl6bIrLQFaRdKLVtmmP3dRam5t+IgxlyBZhkyf4kEpXUZXtrgra+rrf+ntsfq
P45QdAparIW2SeZbH/OqxxeSR5rxpd1esgcYFUD74qe0Ve+wQfp9u93u0rrktX3e6vHIPjjQBUJg
6uMqlcRqPUBHsEi7lnG2x2KTfY6j0+DqrbxX1ZlqprEHiNL/wUEWRJceQZ9U3aV13JQFJamFpS0o
HH6X/gqmp0Rk2z7jXcsNbykF6t/3kNSSxDPB4TqdmYshCBEsgo85YNonndWQXepLLzwPAexkaZXN
6rMrGYiT0wHGb+C5FDzPkx7G3zQu/G3MHaK6pgflv2r6Vj5hs7SrwK2Dwccn+WbMvIPhFAQs1fVP
w2NJnJTlSAPGNost2WTR/31SHjOe34v9FooOFiIfhVZBUOHIPCK1r4tDCi7HnrwY/MtuLXN2au1q
tzOwjD7TkB/qrf2vKFPhDkdBKkV3QXbypeBZwozTvfWTkVARytAXDkllcJCE87Jb0ZjsUy2l8qby
BALWNfnR9X+omBPHIK2jf4FSwTf4p2AqJsaOS7dL4B2AegYN5TwXOSJIWIZ+HJi5wxNZUqYF2qCP
RnP+u/FGRRAw0wfW/6vn9bJZdoZpaFkwOuIOZCuzQijTA4TJaRoeBwNj/VIL5nE804kR9uWMj3kw
QBw8nEaZm552sgThhY2QdBDHw/UxSaBWqwhjt+QnnyQ1Gn2kfzu4dFmRE8KbPXDSR5oM0NiN/cwt
Qxejblt0Jix3QkbJsdpRNPSKOZZKkrHB+dIoctVV9DwhlJDvb1JSFjQiJNRU1vAPOWNXLhvFFiB0
hm7E5b0CZtTI16uiO0Qw3rfwyIcibWkaAJaWmrec5hS6UD0T3w2eXl2Yi8kDlbO502/H6n54BsDb
MTZ9+WpqOnO1R+8WBfrm1NF3oYThyy7ULffz7XptRezYbtR1kyWRHQa5Rje3E926xVa2mGmdMW2L
fLoQnCpLEod92G69yxfwFGNhZFnHP+l0hkVuKj2n8kF0bk64FWWvSUz4lbuK6rtxXE92ZK6gpWAX
P5RU00lXRcd1ceCK6dx1Zn7/R5qF84kZvK0aCdpVxw0ViuuvkVQxlyL//f2PCqbmBWmtJjAbhuXd
iZPbPCJmjvfzaR4my8fK0dSHDqI64HKGtJc5COvnTUp5jR7bWPxLkmezQ8Wdi6y6cViO8WN2Gc0s
YhYqXsYaQCD4ncT8WNRjB5qGqo5g98qaKEh+AlXKHVgUveYIFoIGpiKf9O1A+UXJjsLnqvpYa5UP
DGl03k5lYHACkL/1U8kluLJqfhZSvT9PPbdzAP7uIlZxnOjn0ItkiM8AU1wfNjMbtee42JweIdwk
lAsv05Cw+EnTZzmxqe3nWZ56yqvmxgIaZDndTMRtahRyqmn/hZLGWSG4p+lBHCLaD5Z3uw/MWd0s
H1zXE6hkIUknTSJMM78IxRXzcbNqzlPzbiSVxFDUO6UOjxAsmBuUeSbCRKwF6mECfUSu6K1MtE31
SUrhRcDc2kvq2R5pSyTgnrRqQLlLyFIzsoTrdMyZOt4lVQv72HXWtaiaGSbcznPCCg0YSCT5vM1p
Z4iMQr2nEio7qm8BWbnaL6JoJawS+fR6KqVGensYbg7Z+nU0RimKpaxg1QY9rPDgSmWQJPMVHkAK
0fHoL/gV+IUBqfWzUDI4e2L7qjX7nYLO6D54S+/x+PUrlzYMjptGwhGm9xyUEfxnB/uZPg4bcpuD
efzQv3LVM2jranncG3NTEpPjFgnWHmW3PH9fFV57bOtZQpk1+bCnwU/HE7QZ6NJu8j2lsHNb4b2c
Ht//b0OQ4nVEmwmQPtXbnkn7sofSCcVaxKKLIvD3h8y7wqMCgDohyR3zbEsPCZtQFyIK2CghHJr1
8oWxeHryj6W/zZBCYp6gCCizsPhIOSjjuJa6zMMq5jCJGRbY3IMagLoZGSp/h2h5WDcD3wu4SZ+z
4XYC/hHKidwMKTWgo3gvkw0oiXEK2C7eGq3YICRVS4rhbTmcOKXh4u0o9FbDt8B/MrNnAe0/P7gt
be/p3TGffSU+GPlrfXpwfPkn2Fafr5fEmy67gWQ/GLPjuRexfeiEuqCti6wnmNapp6ClEsgTrByN
qTy6spARDJdJgtkzmoPx09aZsIi1juciZoC5mrVAgrE5JBJPf/s7Pi+2mgb9tM6gdmrkzSAPRgQ0
XTubObsGwQqxQ+dbEudIC9N6JeaWENqGdKsTqcBYIijycQavJqstURv9Ki5Nmr+m4elbokKE5mrd
ClB02JQoN590dG4h8zzFaQs23Gp/7o24Hr8PWHWb6xk47bFJFzwqsktXYoX0upl7pDF+SZ+Rrhx8
6lYr6nPhcT/zHZ0jUoZMQcBpkVpOWpwezLPZnHT4KBgQZPkMa3dJEcre6SvoOFnUde/sNEjY7N9R
eUT6TDEuBPKjWvniBpfbPOWmqR76/kWDlptYYDXVxAO9o/rlaVJtFhgOZVT4Z+9/ypcHUWVYPzpV
WOqWTO8K417J6qz+7qSmLLylT3eZBFEXwDh9VKU+Eyw3edKOTpgvwcL86jLR6oI5xW5xVZk611Rw
xKL3MfhbDP0/eBFYO9T4d2PNMKLccqMXfusazwtiys0+kyMNWAQUYLUnnfEhNkzYKYSPK+NF0NIp
msm7y3GE2rwGtaJYQnf+pVJ71nbRHr6+pLpX3Mui3j5vzmAhKNhzEKuZ9Rliflie3MeD6EWW2XGg
rTg/LjLpRKQ7S5J+PIpuP7i+uAs7SvGLG8Ytj31Ekh9xqDZAOUdHeVpUkCLYk8FoBW8idXwkrAhh
2MimRYb9Ah08E0OLiDZs3w8B006i4g2J6Ri15y0o0Mb3gdmSBNNYN0WmJR9ZNNLGXhoNTAVRAEOv
oQOLdYCv5cQRPdmc7dH6qRZEIlYXgSfbz0FmX3vCp5Q80235m5bs//iGvVicdI68ZxGWGdsa53Ze
NIwROWZ+4yxCRLZZmMhucVmczqndsWJi3sZeToi7wc9Jm36V+VO4aewVXlpzhXXmPhKFunWpqZ4U
BoDBcZMCDg/ZLbb5A2uvyxR8e9dKYFg54RNHh93gPhj7KL6On7towBWs9ESQJ037IQB9w7rDZ8Hb
2IR55AgzJiuQTuukXndGKltQ7Ofn3+Sq5tVzToThe4QvR05IEErcyiwcMaWc3u8aiakrXuGySLKM
zP54reu0m2KuyD7y5JVCCiAIKnrxwlHs2Z87yMPWuOQWFKgi6a9gILejlF5/Pm7VcwKFRwehaQCH
81gPE6+sG9xNuoY3A5MqsEh11L/hflwxleeIj1aQbxJ8K6AznMn3GZAlZ8Nr8XBulGv/aLu1YX4q
aJvQ09n+6ZgcOk7tVmc5cwmvByalA5L0ae+cTGnNHN/diCaTqbG166S5CQ0Nhy4yJsyGVBOlNRJu
mnP/znVkApkS3ejAL4WQgfxQC2uIspxQEOCzXdkJX/4cdPF7Scx/dXlSD5YDXpI7TMSABUScEOGk
EQIKJcm1s/PJlmDHSK6nKi53JQkLxWmJspqN9d4mnTotaEzZZ1ml/7Sl7V90L8ouuPOnwysl1kqc
OiRxcoPUmsGPAo7F7FFDfCbW81lje69KZIdZOtJqurYGyOvCMF0qYxF2cQVu/hGC7J/6bmL7+sa0
vbiqVsjVPQLlCl3xetIe/lFFbpZAsCazdNiUB0E18O7+RAm8v+/sbGGX7FClr42NYVB6Kn1JX6nd
oca/l54oqjPHr0r8aMoWmEnL87J+TVMz4M9xxTOtkUdd7VHiVqDj5qAlAxRxRZMBhRLlwbrlfVtv
TU/oZb7UB9f0eeZpQKUDsk5tnZaVQAN/B1dUEF066BqZ9RLCHulYL5wJUyMt54xWXj51RcesDofu
4HbbuI+k+7XHX2u08flfoCB1ipwJiUM7KW3JtIrI474QK5qz2Rx0MbzQzfGZuNy6Hkq91obPDu9Q
iR5t1+29ZY8/zKMTgzKACZp6YkTvuNOLSy2RKve0wgNrOCjJRbdGn8VCky5pUQfQZ/LZEMzs0ZEx
7Ls6zpw144p44SrFyH1vgEj2nbf77GLm5xPjRdyc4zhol/NH3z84QQ9rPxlNCmIPdHh+5jCtSldG
DaMaApms1iDoKOl/SB+PIs06HH1sHmxSwbCS1BHmIz0udkunjisGhYW2Jy8pr78qzu0VYeSV2wb+
c6fgsIZI3CH85JXifRRW6JO8LLkcEe+fJDJQCtwC441eUMVMhkTek7XSPajNHFOO/LDQUB77OfTL
fXhDiIZv3A3o/m97URF8cBJ2LBwPxtGXOVwNKYitkRC75MyxliR9uBFyQl0eRkyIEeJ/icuB/5A8
fh/HrHsfwxsGFzsbNEcERDbXrgd04r0YTYFJtY8S8hkp+71PoQ19o8rccoW+qMSpy7odsmgfFeAq
IXQVOMCySFOXwbtCO0QGsshnSLKWkCL2sf6Q3U8srrSsJtDHlgY6lCKoNg5PeTJKBawn+RaCitIB
d47Yf4nKAhXW1BIN0dR49B2OLYGk7sYR+AfMOE4T9xI3bXb7PNQPMOzJQ2u99MAYRu+DUXlMziEz
kE2t+ylMf4ck692K9P8ZX4+ZAtq6fzF0QN43KRrFxtA5yyKe0n4JdhAM1JXUSyGVq1syWtpsUq+A
iIIfVZJPr5/HrYIgqRZpK0DHCEiLhQoJ6b5q6FJKk4xq3kdOqYeKG6ZSFBLZHoC3B+z/DeiRjYeK
RtZsy2s0V/6nUgTucILk98rViMzkEtcMDdUgy4UJDid5bZ1GTIXewkckzalXbFX6jzWSy0wW45IK
LLdNZTSaBeyoJsT5r0WT94uJsDP48uxp7ug+KCEHbJOAOZ4A5DpLf6Mhgvn+hj4ViH3pSFUsV38N
mw5ZLLfr5T2h+1AK3hI0UOVMlASX3OSsXiRhhEBt9pOTuSasNzfySg7doHVXBnhSVptBghWcRIol
A16NPGw54GMivVzzabzo6mgSId7sWBv9EpkJtfPhnyMOv65RuFer8rcM3HDTv4XuMbE5VAUmdfUY
A11SNoRvqevmlT/mryhcVvBbBoomvw7xmvR7+ZWDvlTmDWiMXMbzlSYrWgspx5pIMPHjhd6swfeE
z9rmp0WhrxNyVZoicwgWYwUq3BhaKD1nDc3Z8iw9TuPG33g9WeV0DuGur4AIKY5ZogSL2mPD23ME
i9Rnic2SC8NrCAROcW3FbVQ/UMdhkk2uiv2NXgUCQ5zM+KIVT19/ZXeW0jmdLYIwgiVrjWVpfLua
F5HnlKKCrjFruelj+IPcMhe5aI4oIYmbV2goh8MjxZ2kDEBsTvkzNgirS9mTDZc3D+jTpBKTAwv5
6hFlIP3d48YNrkunZ5pf+C3/qlAnczfkCZirCUjq+0cXlvQWQgVx21E34zW4tlw9d6P6YMzmsEiR
33ENQJB5bv2J05JGGfZWL1At6gQfJCKqBHTnFcfrqVE2q0jZ+wvl+QLvYY6Vhbr8eOUhXTLhKH/K
OlxX8YQCp1yWnVAaHxA/DPVzzp9aO4NJlEJaE2w1/doZjSJ5yBGeSF4MZzmNT4kmK14wNCN5k7aC
Cf9J90295iNWdtEyVBiSnMCy6oMI8X+hZJ0StrAJQNbs89vyxote2+uYGsCAW7XMwHKxXiplRbKj
drnUGFxwa0RT2CfFGRypkFhaF2hUdo/Y0wHzf3C0Dg2N5c8U6/NUEvgUWKt3KggVSqZ8NQ2ImhJI
FpyhFljszrnnf3763LJjtxn02oz7ENAa4/1X5BO5dfL7Fq7T99RnOhR8Is86TVJQRsFTfXu7rUYe
FcetLkhz/8hvcSckGhGoz9sY4fe+h9KKpyYvuk6mgipE89Xsyvmvom/IpDapnyNZnxnV4XASQVIq
bdWX1Y8zQZDRNHRL/mDYrO4lL8v1YBgX8e4Z1YR2x3jcllyUDTr4yE7060a3GGps0m3J/NdvTFbv
WZBgboIWP+xkH6t7OWySdJeHcIXOG8GRmlUwm8YJ4k8LbG98TCmmvFqhl76Trew+qmLQ1J2Kfgol
BWDc24QeuLbaFuj3DMLv5aMZjXV0bf4bAy4b4SZjwV2m+WnQMN/AaSbaxEvNVG5LQkC6ipIQ4aWL
RrltMu9/ZYsW200v/OhvpRgFQzun7gqjka4oX7A+AUd2SI8sxdUxDjLkh+sD3Ypm5tTb+uABEJVB
R6fkqrol7PuE0WDl7Pq5F+c5fHDlU8oA0YFMRCHWaKI1swRT+wgEYbd+4R7hPt7CCkHOINDebljx
mEOvkuTPzgTMa5/CsioMdrpzOro0F/bexayGG0FQcBIIPcgZ1iLW12NESXOgSSLe0Rr8Ysgbt4jt
XheCKSWYezJDOAlDXn8//iV3st+neBSbpVRgBufmvkBI66rZha+/4D5GlgLMkBcVMU7ICA6cdb2h
dOttg55NU1yQme+3KA7lG/zB/p6ktxO2XpTi5lQuUIotEeE8tyedJw/Su1arwC2S62OREr7zA/DJ
W0eK8V+I07ZDFuIYG7MXoFARDlQvHY16vuUFcCEuOdHWBlLP+1QiUt9gXQHkZrbtpf0Ypj2iggq9
MpOte+ViivgTKZMa2o2KJTJu8MUmnbCiGN2zbvy1arrcObWZtj4o6dba7trUM7hLne2txcenAY0F
glUn/8qkDtCp5xxaeVxiUFhrnXOy6c50Wh+2KquanG87cuPZwewmLNDE779SqFuppkMObVD/wNtj
Qdok4QIcsgOpYK03ZUfDrcw4IGVJwKk67MDA0EwPt9eZGI44lXWRuY8wcUNfm27O4KGsTJxcQuzH
/sCYPs0KSANNpNsaRJ00SwzsI2jXs2BFo+KKmIRvx3GMs4XyckYTEKqoBkBRvQwyOmn4d0+3oT3K
lolIdBRs7vOP1hEtViaT9KWfQ0nmcM5oNybwsECiL7QW1Qk9t52mAogHRUHT0cCoMbRNv93DN8YI
QmZXCqRefTiGkakmQibruBLc8ngku+/aPjT8NzNCMYyaLru2bzveN6WxCl69eeGnB+tyOUANadTS
7iVH5NzXqbOIoiixEYSy1kiA1C90gG9JY4TakaRGVROZpY6B3rfZJ/BAnVxWwjxSVKZvKSLUfb8K
bpYbFIVk1cstBa5cxVH+fKWdYvpUFDdUkh9L4m369MyyuyxS1ZBZavnRmcMPgUEMg3T2ZSBG/8hH
BTmACqlMZ3+60CqzogApdouaoXHs/0Q8v+LJ1n0iGUKjromaoZyyPmRDzBsFsJTkbD61pHQT75TA
o50yaKB02xWtCW/sDr6KbYtocSK27LWThPMycLQMp6OVfG0hehaQkn20Y1RfgdeqGTLEpnZKjUCR
YrwbZeRPy/N4arsp/GnIdlEwaKsY1OZtpu23rxifij46tsP2vwraEK6jK7gxRRvczz0petFbC9uv
1qQnx+Teoj4U3PLPIc6KkAJ+IYDw1i2By0cK5HzSpc/rI747Q5UpK3FDeZeaVTVyxSmW1PM5xcSm
JfJPVqFPrtNC9GcxpTPOtQcv4IMsd/sjXMRYHcj9tkE4G7vryK5IfJ8I+nbgTOQeab4hrBvDJ9vR
oqG0U2p7L/Kc9RPd3KC10BLkqgCE9n2vP8D3wxgONPogRbb5FGqf2KEDqaZU9vWb3QQSeLG4HSPX
KwFeO1PfEzTw4pxCcP+BiDTyDhzt33fyP1691C7wzt0menIDJHQD2gzNE3z4jL9a4pp0Rhzvg75E
Q8YPNhKrt+ZoTBPBxBTTj1OCD0YnzV1jSCMbBfb+vqdj7EuF6XgjQZU5yI+Gyk4FJzJcFTRazbm7
0PhZM1vK3Yc3Lhk2DJ8nEBnGQO6I1x05V5lKRlAqLepKNqgOP+ESse+G76A11aCG9p+Y11LhXfAm
WOMscdqAewYIL5N+KcrjJ8AX85j7wdRsgAhQgb7a3N7gmgsj6ZDquMUf016VILbBOPVdtldqjewA
LUo4lioKxeBu505yu1ZsEn6x5lpOmUax521hSIIDfzwtrTXhLA/YrwpEipA0/r5tGPBiKF4ofkPc
3Pzf8ZUMroSstqMiNrWgNRO9Rd8VCKWeKTZ5vRkS/1w0RFroNBvLcod520/Zk2lHVsA50HHGdGTS
nyAPm+QkSIqQya/A965Vh9yPpdw9ou47NEU3t1/tTZ41IzJhJMGzWLgNtVUiL30ThyaoJPeCwqda
e1NgdY3peZpCkjyAbMAmfmTz9hykll4dc61cEscXNkIq3jFNetuJEC8unLYdQLB7rqxMc0D+01ku
phDwNSrYirjHRskqX4M5SZRIzUq5tV/PIrmXFiiX8EqMcVazTdwfuWd41GH7CVn611W+W4/apv5f
LqA+0UOnXRRyxr1EXQb2e6QqQoDRz9OJ2zxwSpP/hE3eUaPxWDRU/hjFgJLJ9UjgfakicQKPIqJV
+I9uMUrd5hxv/c5k+cVgsfoMp5iBvSu3bFaMwFgbdTFezPuy5bvGzYAyD79YIh1GUa2Xj948maXW
mw/ZVllLEvFStdkkpjGpSbDsnU+PNdFkUa/r8luSlaJs9PLn+8zqcKioclXD+KwC06vefnH/Z43E
J3qxcs88HTYa3/GtcyIQuMxqskTwMt30MXS8ZtwvHXpYAEQIck8re8NNsuuSIwC0Hp7a/Hc+J0DB
aWofClPTFWaBm/SJCi7/Ka0gccX76YQ/Y2AJHpSj6B6yVLGwQfRHx+KDrLQnC998AxYcZud8C0vQ
6F0urj5JhFNNSlXU7LXoH2LwyC9hEpscLMry8mZAYYnC2gdfEes58sW8V3c2/wwfcCAj/oogAc9N
viVdj6hb38JibaO45Z/guHxbMEYNYUIloHdWJLMCwjyeOoja5vjtvDPqRaRygEZ4SIj44pgNEOt0
WkGcc8yWYBkCenYWXYToE7K+QnYHkCxPDqcWcSPRFzYDqPDLOvSHEk7QT6ifc8MzU1tS1P2dDDUE
UkdbytdVJvHdBlIXk3+Oe/26nc8F/NQH6evGFJ9syRc6GmZsHUjLd6AmXdS4hlv3mMXkHMgLNhA4
ZiuR+z1e6kQK/XHeVcCjaQkzVOZOivowzu4IQLDH8YrRbAWNLJvGZW1anNxQk53zDiM0xpkF7HzH
6Monf/2yhIdVNB1I7+AW5CrXUP8wU+0uMLD5cKQDaJF92/H/J22DlPKVTmZteBfGazltHhXuXKk8
V9SRgS3SUBeWxZPNt34uEZgUQ7WORwbQhihckrxjwuT7ftwURyK2R/E3XWUD64lE6/75yrAtrqyy
u32vLyd2GugE0MOk545HtaSSNlJwtNbvfy6N9CuDI41Lg6q91dzz6hKULGwm8U5N2TomSn3B8C+v
BJFtG1zGp7cqmogL7zoZtycFyAAE1ABDQoND8DuA8NGzdlOIyxwlYyrEtD2R31M2p1cNWjhf/+VT
DPYnLJXZcjWUU00o6in3FCmGXlkYdFUUQIyxgIeXxotynknQiRkUKVCwuAJzt6aE/IXC7Z5Rpzzj
cmqPphGcSO4/jhGsjr3HtAaIWdCetVHttA1QSGURLnf6H/AuJ6k76fgD1c5fmCa548NBbflObTVf
4V+eIFEWhqNJg1vA3nNilDX82yjz94K4RIlseEiGAj4NpR1/+H+r0bPEmc16KmapasWWETeSdAxW
EttC5EBGYR6XVvdo/fstnQdf4pfBjbLIxw+hbNGvitJkor3cON5yQMld3MmGByK/BfnwPwKZPwm9
9lNUC1+7K89uv04cXujcEwxyZL4FzAo16cY4j23PigKslIi2q6gxZ8VD4Q0gb+2Wl7zjyoP2cz+l
6gtxXyphhPQdsDtueTFYS2kg+xEDw+/m4Ojwy34uQF87Im5Q0ou3Lzr3aebTXfexDu6peB8Mb0Gx
zA1lolrCj+L6HxjFaEsO+Pc4+xRGjhEPZMjFGLH/mgjQTMTOKCdpuc1JzAJWQg4gRaP1OZVPxPzD
MDYp5olgldCX3YHAtgjpiJyf9/xjb70sFVuHRxfCN1WRiEw1ly/aF6wVKsCJCEYfcQtNMJYao741
ZSEnbTDg+E6ylrI8YAcou80mpzfljypUdTwO4clMSbcjWnkmQC+54eshuzyVNMTgogSmPHUEaErW
LMuaQw8dcWgB2t38AuDYsYWK6XNTwOqlfboDgQHhAVKZj2kArs7/hGLWDUPgUGgfYuaEahxQgemi
Oc4+Ry5CNpsxWF8ugTtvDMSf3FIGTmvMyCVJGOx2aEJjCdDPM0YiNuzj030jDAw2cvj5PVaAj+YZ
RIYO2ItM6UWQD+cn+s2t5M0bUEncXoQ14QGLQUGf4lFv6rJbAn9jZVUAiDD0snZyUiyQK6H06wIU
zBqsLf+GJY5NsedcnpFCcLZupFzcxLC+g02jc3aAWBzO2lCZl2Sqx8fhF2kw6Q4CxevFvMIX5Ipc
vgijq/CNZmGjtC8k/mTFDCqOibsJp9TNRlpHJArcJ2+VSCdwGPH/63onE21D9DCR3kVaJ8js/rTz
9z1PZAG1gW32kNZiF8HabnlGxnoD4a0AyDWtR75xRzLdWR2Z+849gb9zuNfnMxiBEvU64im2sofc
mJJGxXpApNS7qvLemV6OKngfXTP+4E4OeSih7c3RfNN9HnQdsa6e8c1cVLeeQlABL3QoNhl+T3Dz
xHIJJ4vYD5b0TGA6c9A5Gr0QQnCDYGv5fVlYK0hgP09AXGZqFy8dJ0fOpE/wzy/iUBzqd3ciAA1c
OL5WnE5/RKF0zdqYDVogOmOx81GG5OkAN4rCBHEI+F0QmtCwOcnLPFsC8DIZ69NGS1D65LVEh6dv
uUzU/bEgvPQNjBq0uoNzS4hgnxVl4MJrgMCL7dCcb+gKDwgpu5Ij753gohOZfjBdxzoT3mD2E8PC
rBdjA8+b9AFIGMCOOMLzLr0MCiJ2qm4obBCUoMUmcTkbt09XxLYh9BH4duLCZ/njJ2YDanYJm+QU
rn3Z1j/Z4naldYpKpp8OtpGi7IAbsfEK61oQwLUo7WVSYB9HcXpeNjhD26Qo4fgKLeuMHuu7EM/b
8T0kDK5paOQKIEQcF4WoviZTi5cFfKWKM8i9FMuS1YBhk/CCK4OUUt1xl+8hsXccv4VUc0aPGlao
Lc/oqkvylZhAKGqZYomXgxlJ8ZGa3y1vpUNnczHC0MdSTwpj/YFc+F35z01Rg830TF0xmEVqkPrK
Pe+VUAu0BQU2h0Ilz3CZQeb2TETgYCRwYgrG2Px7w/UcSY2tjojvaCFWt6GJe1yWFckKbZjlqqbs
iLgab4/hurJHcXWk1mYiDz6LX0asZ7qMr51TcRqqPjFyEPs1HJ+hWkHslhvz/yTO+BMVQntkWXlz
d3t4d4inWUw/ihncdSV6isQQ2VVrHASIHlGnS+tsxujoPrRXpAYQ9bzX1C1FYiSz/xXgLDcVFUZG
/cdSyZvxVILaesIgie0oASWxE+xcveB62ouBxJeWsEr2hxAJeahxts6Iwt2xCydNfHJC5U+p/Haj
n7vFZv4EUlNDUc8faN8yDssqNH80yniu0s9UHjmKjUMbZuMRNbSkGOIbzAxidfsdY3CRyuPmR9+T
bo+owxLuwmI1LwrwHP+t4+d786o5Kth09DpSmkoAL+taa3iJa+VQzyi5+enyH42TQDJhsT7BSnDl
xuIHG0T8iQ7m98AE+wfPRxm5JFhOxD/5uNljFPfn6o18QkLCmZAlwDQrWaC3mZld/0bImnmw7kZ/
+B8CHIJfZMJP3unRahaahZDZNj21ZW1SpwKfQUofQqamApFV8NL1/HyUyP2biptpuGlt7lIiX2KO
KOm/h147t2F7hylkYz1HO/CHYQ+0+4forJPyzt8AsuB/ch8fMuG9TgMCqViHwBiC7HL2pFv6fmiK
EIRE7iWcrJ2nk9zPCTAhzCcakdQ9gth6HQyYIdqmFNWtPP5kQtZmblUzGFrMO4jBmpvqHWuZnBmK
6JkCKZb/4IXYP098X1dxc0iYLs0k/kttLFIBLry0O/EI6veDv69bbO5hS6RfCEEIXcjs0VrDbM24
QpQfm5U+ZdleVioZez9kHLJu/6yEIwMGKmWc8qhOrbzDHSuLVLVrhVG8gRqXERzqou4oeED21DAM
xLfISR87qS/QoJbJHMN7FzAjMUmbGIB59rpBCsaXhOpW+YA5NuSSPwa+skJFb5tRJbjYBgBckTbA
3h0EnfyxevDY+pdL3lBKZQz8EDza+zw+oH8t53JUHh4x55UCAuL9VaJbYvEQwg2gJf0OMZZ3WKsQ
6xM7minv5iGzoeKwn9SRMQ2vDmR/NkTftK+yiKtLlRHCo2c5rFBYLWWf700B5yna8FAtAoChDtFu
7IkWq+X+br7ziEX1AMiblgaImlxbizbvI+snPX0EgpchGJCeGLhglZUCTynjzwjXxmcuALc2QTLH
PMC06KJ/v6+FhILDHS8DoHrMR7zMu01wSB+KEaoMNTg0/z+orkEsijPjtJ81nPmqCWLm+o5Qecl5
ev/1Lo0UxOXxICITUPiE6ZcHBFJVbCfG3PUpC8V3ojTGH12uV4xjLFR7XOTyy1GWLEj7VdMi5hTe
cNcKSl87+wuddTLlzYbV27zoo34NBpmaTwaFt5RaQn74YQBmqT2nes+qbkLGS9O2VnsJzq1Et3oH
/0mlxM1x+rBoC96ow67VRSHt09ZACtDTtdP2kTV7B6NjVnOY6ANwXyC2t2HC+WwiE48pTzCYzjgs
vtcxwyfxj2rlbCdWUeDIr3dYWvIF1ro8g/6Uk7Lt0COd3d4WePypfg8OwkPrSVEfyEFpj+jGZAmt
s+6lEFvxmC/lsT+DgSKFhNpXDbXmTwuX2JfAoE1dswto1v4hmjLrlxSVnxmYI7MA1FSoQZXK2GoA
Wb/jGdZZnEa9G5EEOjg/AEQfqpUlJp3vQVJArRqTeqNYeHFpWl/gaWh3/8Chq/W+x4m296uk02lG
8CBqpgGKqUjtv/Xg2Ydu4uxmJ/Q6nAfV2TZnNdTo7EDR/z4FqmPtVqXDh5YZ8aWp8Y1KtlBzskpJ
kx57SWLv2CuJHSkt7oRe7ut2PZvUDGVJ9BcyWjSj6hGQXh0/N+Sa98N7uTbmGk68WoU3MDoYJ0Bx
luYB6t6LLjM0uDdA88OP1UL2vN7taZAncDZMfEWhLv3sd2oKAAJWpRPJ1bgPBi8sfisJmwoQmw+Q
BPSx9B73mVOEgl68gCEoa24tVJnoXOe0mFbeuKjGBrXQyBDbY6LjQ3tFmhbce9sREbFupZRsjOag
1WsdQk39NXyN8I3b+LiakPLPH6WRQDZUOZgYUlXjdmYr6uLgX7XVbfZ87O2FeUgwM7ze8pDGuBBr
HdsRF7e7/hSolNCNj5y7cAaOjHc0CJ2+wjv272u64yRY4sAYDGUC5W+tl0nbIbnL5i+myQQKqZG0
i5ZzU9X/DP/A6fmFVPda4lxhRZu3/PrdcxAFdgrJ/6X/rDHtrLCRsuvopvRWA9MH5+5GUEy1jg/a
oR4Oz3N/iUYxhzepKjTy7QKCZiGQGtmDX+/YGDTNh+I+vD96+4sfwYdHz7gcnb3lwmaURVKOG/No
0jPZjOxWFYQl2y6yK+G1TyDSRzkFbJtRAP1diyK++1pP52IdeZ2lyhhFdyZ7vblCPHkGrImGPNx+
8bEkBUxPCLwVinA0zX9UOuDCKVXEsBAnU4sAfxhoH1TzEG2t6CfBLL8nRQl/bPu3yWPjGusVJozw
0KjpGqYwNVAkgmN4SwoEfbrbLKRIRBZXHYbROohhVzxykfcVETmRHXrLPzPsKELZ/1Rz+IO5PEhp
w6ADLzIUk4ml6JXGrmCZlNtDZ+YaJqB2b1pO6yUjvrmedso+KWjJDMdysGv9dXQAl5AO8XCZm0AO
Ecml78aRMEMJEwEClMSCjnUME9xlbNJw4gcN0OTn4q9Lq3RnUF65PKSHWCb6dByTn1QuABCAF4dM
qxPchoAD4POJxOxpVKMumlPZbdd6L0cS2dUPsiXkAbbeRXg+XzsxRDpU0JuwRT2cuoeHgpaTZcHf
H7dTMVIMOd4JOdpoYenCQ0I4DMr+1CHLY/GI8nNptwUqX0hZHPx2qcYyo1e2cDcPwuGrKed1Wpel
mke/YMh+nHXD6CScPwzb7R86F/22IjTp+qbMU7USfSkK8vFj55l6B9BdoMXyW7com/rKbSnpS37m
8vv3Xj9wfuzXekqxMAWi0Ar75GqqVNgj3pNZlN9awsprLUSSnJqUY/8GoYno3BrwdeGkqVqUn+6D
4aFQRuzkod8ke+ekntOphMq0elQQQTeSRPHAidk1RjHkI7Jb7TDG8v2QQ75PYJcI8YtTgVSF/5OM
8N/LcL2a4qp4KOENPP4n3zmHu3Lh66A6sGHOatB+p7jKu8KyjzhSzViUa8eN7Tzn+t1FeepSCmM+
nlwVI1zy5SeBsiqvEg26YO/lsdoZg59uvwg1QxYYW1j8MoQlIJPaae8NvJX3BaDJ0XWhnoRzjTKC
aFI0Pcz0aLXqnEpkRR/goqevrHDh2a89tVNhNJrY2tcR7kza+GcNYhb01b+XKOOuOY9EHVPMywag
FgOfc0Y/n6dMFHPMnzZVR/P1hEEahxg3Tzu3dpkcI2EZcZDhgFIZSZx/u3D7lhv7dtpRcPsfcVRw
21NQEWyAVpJoHsIhCvkm2ETJlxPF+55AqcKN/CH3JJtPaFWsbCcdm6bLTzFMhvHzQXREeWPfO5lH
xVmct340BbcvQFSED6/6nVO1gV5G8F0hmxmvKBgKMvdr3xxX7TrRipXawOSMuOduxbtBTo3BQn9Z
KFf87QKDOzz4u1AM/4OfVh71hgR44+MvIJcgBzBQGzuj/oHNY4jS7I7yMoNPZ0Iqdp//TeWuKzRZ
fa8Z2GYguBqMBOexqfMGd6gVTvFSneHboP71uKrSoFJJdPnVUNIQuJmTd0PxVE+JlD3X4doeNUJM
00V22aqWtQ7ikq9J6rAHOrol3dSONtLBrUamhLuHiB2DKTz35DQejfv4RRvjbUhApzmaH1NNdY+q
YTahkOKJE0dp6jlyptZ5CTvvvSITfyL7TyUIVDq3e6TDqDMTpDVAM0aTNljYScB8oOcWha+Ononz
Jtemyn8GU944uBU046BEByi2DMXeKQiUej3Oifu6jQoXQ3gKdwDw4gmqlEVPEsTD5o/5gbjnhOBd
aiIvC6wKIHYpV/XYBb+oFA9POvYAZEyIwsJL+13QHwsahuvyVWaz98udPT9+rPbjN4EiU/6IxOfB
lHJFvCmjvcFSch1a6Q4Jmbse7soGctLaTl65849JFOgx1v8B3eN7X/lQ8tOrFIxbSTFjLm9CGDCG
AyJrIF5cjki/Orozoir67/TwxS7rZ68LdSfBPpZyTOLtA/vWX9hhlDhaVSo6JuWFeiDO9cQ6qOsR
rjBRXHAoiwu1PT/P4xE0/jVZTkdsu80lYWwMIJ1VNtzaZmwJdMoaiK2MtWXDDKNb7N7eU1Ww31h2
uB+6TNfT2fbpSDFX7K6J8rilOCfe1+ETWOLg+V8FT57AOEa0ucG6yicCOAq2vGYTtaLK9C94O9HA
5iQmxgT4clRD6UVc0mPOgkpEF7G8KnGnJV62BpglkRou9aGw3vItIPu8HEkvg7iJ2ibYeRP1S708
uq50PDFVYtXzYZfIh/oaNibKXrO6zCFRAYcEkyX9WsfwnPZvDCxt1Ryy/yQiJYPRct6K82mKeddZ
YC+XIZfcLRRdQy+FikC791CX+iKGXdfvp3urFCScgC4laj+bM0O262aV/20nv2UaInj9F+xA+rl/
1hPqa4V8C3YMElf3x8upglX3T3efNoDH99WqfEO8kAb6UEc0170BP/1U6pit7igvNbh5YZWz9SXs
ApxK4rHdpeq3eNaZ4IaZpSeAqsDUcJKcwBrcUzuMDVhdP8jrtxtdVmA3Yo1aamvHPG7+U7w4Lqq6
Z0LK2Y+nMBSdMCF9TvAGEqplpxsOTjaB3NQDEynG1HrzZHhp8oDnk2WajCVgK66IhfnRZCtp4ViS
ddZbqMGgfeQ8dVhdAc4T1HQBtl5Z4S/joafW/cVsBXmPQlfVn9lDUuhoVZEynMgK3wnAzGELztVv
4q+wyilmWpu6uwfQspIB9JDjJqg1/D5FLWwpgSnhF8r88KSRs9k09xQCFqWHecEmg2Mij2E4s4zK
43RP1YDD4xX5vjJmGoy6XCLwmNKfJE149DJZoAFkbM+naRSXNzwrIGA8/LbiI3Bn8E+1daWzdTKi
dctnVyBTWrQmWgZFIPpjpYOmwmuhIs0mfyfIvujWPR6IKBXOy+A6e9XBXKXNYoq7dhfmA6Edh10W
+OD8FRWQpevyY+8bW2+LmDtMhPxSC9E0LvmfXWyS78qC2jrKP+az+2FPmIZY3BAw6A1W5uRVaDTy
hHMjlgR20WEARUvlnRyLBxVJRhxAYPuYa/bhv05uA1MSKeId8F/w2FZQD9CfGRvvU2o5c5Zevuq3
y/+H+dX/HoqLD/lwsI2Zha39UjYSYlCvYx3VHR4Hp/Y1RGc9jRlLZ7kABTJI454zniySrzDZNNSx
6ZOnFCzqIAfAT0/QV2zxdmD03G5OimSwL+22glq4e7bwMgHDnP/pbrdC32cSr5DPsCuoEqN5WmsO
iUsiCHlEqL8jq/b5GJsurad0wodHWKWvd7HhwwYYHiLM4cr/N/hrZaHEzTCevAhJxzRv6u01z2Wc
2dbWgWZTE8oKxJBG5CrXOCxeA4ixKR5thOVOOKUkrg/sj0wfN+QM+qkEWyIe+pDcT09tAkhZaRbF
6uKkDgOlPeBL0MT+CdCy53mE6cAk01kqUIkKpr4fv7babYWU2InZHZFzKar8Z2DnEQIXPGei6gSl
ureMSWBkNz3VndQ+chASc/O/8mWAOLUtPidIyVHhAsByE1lM4Lf8g0Bd4ZA36Y9uIZSxebatp9DB
dFUQV+4iNpdbM5JkS73O76nhQfV/MT4G95NXuPa8cfuLP5I3liWlEP8sgPV7B68Ci2gxlxuJbC0x
VCJZCsYewrOlceabfWE0MB78gIUIqDF9aJN8ef5NBPSrUqpkWCp6ODqRqi0sLg11vSoxnBWIYfiz
Y4S/odTYOOoK75FX6X8W/XX5+a4UsCKA2sYFGoQuo8NVBAN+qopqLtTR7ZGWIewRQ1x/CkamOQVz
xXevly14824zzTQJ73mqHEUonPtQEp03eadpQkdcIfZ4yji59b5gP+NIRJhddWB/oArsSIYHyY98
NWY/Zbx31prxEE6rIbDZymAiTySmkpgjpR4n79HcwzN7rbn2rBmb3vLLjJTOmdDfdIRqDiIGV5Ud
NguM6zIMz73OGpLeM3FMU32OH8p2EOlfteNFXZJS55kl8hvqs+Kd+BBTu2J16MHYRbElZfrcwpKs
aHhwWu4IJWfDwo9YLp3yrxPiNBXsqs4YbyImV58arCNCZtZ2E7Y+slImtyrfVj4tWGppRv6Tesq1
9fsYCEba5021BC8Dh4YNUMSwRGzfo62lhR5MVepTLlskFOqMCvpRQWD6gntJJZKzAtcYH4Vjoux1
2o2mJkm+GbxuhkqI4UdX8t4IACRihUl1nYuFJc84Ut7gMk+zflob1J01BIIahof82zULyEcmjq2N
cacPI401F5OFmQXIyWhsTXdqMrEo6fsMC+RG4uZ/2VMHuyFTnGorCqvV2a/eI8vMKnyxZMLzLUkp
hMuOb+ObXDRIs1/ZkEoDZm7wzewXjBjUQHzmRRrENRT1fC3+QZ9wrK+qmZkpJvg80AZEzGLiHxLr
Fp9dytn1nDJ7nKrQfdK64ZeJ3npThzpnAE2+wf83RrotCh+fJSIdiWjSWij66aGaCtiyFCS0QV+y
/3BDvTpuuUYhrLSTxKviNtoqYloaohNt20R1vD6v2ShdYHmbinnHaY2VlapDNs1fnPFK8d/utFaO
FL+Q7iAlQzg/PKygFWVXUmHO5SKN6ici0FNyCOq09VU8gQLu398DHGfK+jxne8OOCu9Dct/PHheU
e709NvJ7pgUy7y3q/d84mH6qIWrN029povIwKetyvcxXac75M+pcPOyzOyXw3joj9lieKG53cwmW
27zxH2X1OHBYUi18ladTsPFfGU5EsNOrT8D6KIpgmwgvkYrOR3rFaw7xwY9ijldGqRJbfRFe53wn
4iIYbGLv5E5bVCsz3qTavFqpU4fsUBJUoHuPyE/dgBt5ZPgEswoDmV76DHPQuDesnVMlZLwDzMSt
fZ9k5CbNf+7Fohy1XUmtJWSNh8rjxByPw1pQDR9TIIL704KIpDgbQgKWZCVf6gvWCqoL71YVPQgY
sEjTOFuKiRiVZkYa5a8+6l9UNHEKH7uSwk/FKeNN8cvdgQ/kRTj8HM9r1MLQVDlCEUzN7nMKsCxc
hPB1NLQsUw19P6w+v7A01qROulx9W9ALpj3Hvk9fomD3H7UtKabEvTTppOOvK/BmJuNmn3WO/4Qh
t7azEJaSvhelAzveJMsPA6+Jjye5sfpkrukc/WBHLYgk5rjyhxpTR3S24iydOjj8ZcIDP971FZEW
pk+k5ighJxHrNcLf34VlEIrR5p3tEINS9WK+q5ZXcGWN8yuf0aw/M3vRXSUMR2LIDT5gUAKE12CR
v29pfY5Mb7Frs5eQcSLvKHZTFgm4yRJYnd3cym1DT5zf8y2l+oRK+jl0s6tObxD/5yftrAx6j6Ai
HUAJOcf+G7Rlvq+yZ0t4kclMZnOwg9qz0dJad5rAXHK1uUZINOMZPK7/BYmgJqcmtZYosi0DRM8Q
Ys7rXmz/+5wsvgfttvm7kG4lgk0TbY8Wno5nHjImn4SHtxEjbrTAV8wCDE7BBD9surYhh6YfzLnw
jCx0iSRimBmL5nk1Eh9Xk+UBRB3pJl8VkHqLSZ/s+2CGsb8NzX+F1FSaB0jjlPBrM+5cUkcXkhCh
PmtySwt4tTgEAZsSXpFLuCCr+MQ4dnjdEz4+2OpawA/LszWsphfVDnYWuqS9Mgm9o1pDnEwEXpDQ
AYJ2HfnNMGJC63NMHFBLQ4+lbaolm9DCqHbKGwMJdPwgW/9jWBeS80/sWN4bZrHcf4Wd2PAYDbzx
BnLPJUtgn/0H4hRL5Ts9B2Y0EdVhV1eeuVYBMHlWtftLfvWb61Js2tWvuOpc9mV/tw1SQizHx9f2
DI2Gasue1NzY7mukgVyNvwZJL0FTRHGqTCDpXBwPZinIROhgT7+a7fbkUffl/ZozVLNfC95FRMlb
5Olyb9iTX2j9qqcHxS0pjaDbNR6XNcJCH9RqDZ6vGcDxmAX+Hiti+w84G+z6e7Mve8O1fnJ1VWE9
kLCNNQ+Aojjg4CXLHEsrToCF7nt9W8RhrOSA9B+DMmfFlTH5vDHNFnAsGJ7SSG7OsBDz5QJyNhgS
O/WeTGvagg9jHOqtK2M4MHSs2bZx5jL0Yz+pDeabe2t4MvSZhI9OvaoJWE1rXTcFRbN/EeMSxmzR
AxbVX2IqzGw8RdzL35ntg6iR4bt5bn3pAzGIxHO4o4T0YBnLp/jehoLcH8iuVM3C6AR/v419wE//
FbN5liZFU4zSjfhijkiDnV2RPOXEtxzWC0em4820SaXFX7BpGTn8VpPB8q+EY/Qe1GEd7kwDiQmY
9IITdkyQMZBi9mch76sc8d0PpIYQIFGdU+qn9QpHw2MlhUvU1KVtRE6eKFlDLP4i1NGUWlhZr9zU
sHBa0wiUK8eXjG73xbDyl2IYRWSZqZqv0qWlY8gc/NcxNOnTgs8ZbZQQs2JI3StJSsBeUBE0lYgb
zfMGUA10saihA4Re1CsaBoLo+LKbsad0TlM50ULVZMFLmRWydHV/Ez0DkQ8HZoudj1I8hvYHnNNi
yDx1qTUaMtELrU06gyJZMtvd1ytNqvWIdTB5YW1rlu3dKGrzQQ+YCJiMsLWRVGQns/Zojetgt6O9
R+OapHpYqo1opUxNIM7ccS9BwkYEPjX3/qmXg2JpK56To0QOrOwLnACBlcSTAKEElbP2xoqCvMC3
vN+c4kJLbXZBAI5wb5kRXk+cGyYBjUrG/7HtAGqMXOjuqr1xNTPtBEIWDS4vkBgnQrCJs1szuuEk
gsFOn9FjgPxpKZfGFiGWSczn+dDUJiNWhrVOPehl3T/Gkp/neB0W7YcUR/+B1tFrThenXjkmWf4p
Xx0SJI8GIGilIb0I7jp6QZgiI2+xYWSxd2IWd4Le3B8cb/hLbInRI/g7lB2OMjRYs0euGEkAdnta
J2ifOmaPqdWCNwRNwljk0lcM15pvBNrMIWjLr16jBcgHHglkLvtH7JnD4U38O0GsA9tE+svofGTe
A3+JPdmmzhYKDaAMHDyxVr8/0HHJ8WGPheHg6jX6Xeb5wwH8LUxxZ2k5KoQlCWuwrPrDgjCzxYZ6
Q7fvB3ecx10rA8YtlHEmazhRt/o9Pey/2B+y0OixElwVHvi07l05TTMYE2vmabJ5/vxr9y5IS2jy
KEGgeClKlMPvNmw7JCiw7ONN25OZT7B6xwLcA/vO5GeyZ3dm8V5Pp/3A4o5C0Sx5kHmuMB+hu9+h
Cf5T8sNPO1Sd9z1eD95qEve+9rwQHhFLWgX0LE1BfNLnkoJvJWuaFzoGo2DEGfO0Q7Xz0Lzi0VqP
SGJsavkSZhMa1kIyYP8HR4GjE2ASoFdq2sBE2J8e9NV4DNLPQMZDj5u3u7ZVdZS02TRuj5Rx2QbM
AKzP99GaHOWPebgMxyVdcFVDZGQKFSMk5ukCY72iedO5w56/KWB9BLMUxHuXmu67vLDBmhmbJ3S4
CFZpVxagAkNu/skaBoTzKg2jr0nAjkIrjOd5ujGtwoyfP6hE9J1lkT/VnNPo4OEDhLTcDWP7JRN3
5Pen0uO68xF8oMHHUfWL9kMCy9BWdLEalrkrCQpLOtUiYjOFiWnxq7q6wxxgHPTIcav2T11Qw1en
y/5NxTHvBcnlgxTW57LNR4zih9mis/odS2S8H+k1qGP504c4TUV2K/0NPs/B0I1fCzSQobDtS1ZC
Os809IOVQdnWJE95ob2iEUpr0u9bjq7gy8SNE7rHdqwqpx+yemEP2BA39RzrRsjX96/2zrJaYGPZ
wSYJsgaYH1KJgtaSghxlBV3AcPfvC9RpBL8KUNtMpdv/YyKYQOj43VSqoT461VMqBQ4ZFpW3IO/2
FX3kUCRKNLkVSDjQVWYDpMHWyhgNYE23SbEmQw1oHzncn1Z5VgiM/za8Y9/c+K1CEfepP+PQi0p9
4awRNkz4SyILoA7fDAsroWAiMsgS408Ko6nBAqKFsXO+yvgcggsMyH7E05mu1/kxU36bgvB+MSmx
2dK5P0KFwBp6n7yT+TBqtHSboG50bYyGl6J8Z1BeM7EKYcYceaT0zDyxHabT9rKavkRx7fcIbn20
/xcRmulm6tpm1IzDiAMdrS6KCKnC8HF2oZ1w4D0ZpKimIP3etfswEw0ZGFiYMptnlgyOKLfKwlfH
auSHA//6MVrTityxDaCOCYzMOyljwpAuhhnVQwGUBxZOdi/dQhzImQYpPXdxeckd9y1LMBYv+XOZ
ewlQKBcg7GvpQjcD1DOgttgBOVLEyzHRxSbiORJwjXyyyNRQY/rUc0i1Em5Q1nUCt19rO7+dAkP9
kUm8kyjVcBa8aHUHfvplIuN8gJQ4T1n17jDwuN5Vm5Wepuv73QiF63UEWtPFyDkB7swx9QpDPUoR
ldhs9t75RB1igBwJMkglygcEkXxWn7IiYuURNtKDupMnNo2Mdr3zmlzo8jPCX/Z1y7H+ZC0HAson
wWjBXCbw/mmYunLqzJDAoWhgBEyX86tC6A7V5KFLsPzIWPv1RhZ8Kp2wk31AnYcR7OUBUVMFJRmo
MkseZWqvq5IJnTdSVINbCeWxE5JPxL+1+awXxJVi3kV+zq98RLvvJS0d7HbkRVW/49+2//vsPs5k
/aUNInAtbKPgXz/TtERpssTttnZn5sla1gxN9tGbsttwtZAWKTxmbbvbxEnwt9mpM4oPLS/+8hTm
KF7IWm4ySwfa+FCJjLXRJtx9uZ0IsOWcy50NFCOPjKdiJTWhR/STETvyAA1WmUNW2sm/FC9W5xF1
SYzAGgvXPjR9t4daX2DJBU9KeTrhvyJ4THPwa+FC9gBrMg43/tPLk+Lb5Q3RFAy8QZ/FNXHig9C4
0F/beS7dikdPKEF1lGk7aekKytXyYqjATz57V41mTplbqMoj8v3BcEqGxGjFlpjygnFyFyq54jWZ
J+alJpWaal7FRBOXC9Ohed+7VuzGgQUrVOyfrX+/7805GMxjkIrzrICIXliXpL3yM5zsHHDv8rrr
IRjSRWoSuhSQ1cvk0ZYSh4SNZDdyqxa20ixmEMg4f6uy1JvLR+6LPf7W1Tq8Ye2no25oERcX1r+S
kIK8nRHg86mNEyKjuUM0jzJ055YVucvmKmnk9tjx8aS+za/tmxadxVD8Kuyda5Rvn1tLkJ0ooDOu
M1EwFq7hV2KaYC4uv69gbwrwDNRB+/W5wJDFhLIcRleKRPE0lqIw17NpyCANg3zczldFtSYZ1gQ2
D/I1y2hbRiwL59KMIQKgYmHo4fYINOQ4fSM4vwn+eo5RKI3Y9AwvwEdVU990upBzeuoIn1sV7y/u
kFlh6idHdZXFhSh7CaKXBEW7iyDfOVyeWtqC6N+gkI4j2vEvz8B/8l3nE4I6k9kLzZkTGa35e+Sv
2YbPwngGdhN5TOm3oWiawsBVUyqx3ZI38PxXDEs558rOJWZM3/42tajklvSQUa0KLfOuvkmeiRPR
mld7av7ZcBkUdH1FCE+KuW91w2SoJ6aTj84nSb3knDGukva5Mubpw9BIloG8/njLdZ41OzTy071W
7kFLlok9tWP1zeZGSF+eJDmlxJdezRa+PftZ0qGERKYEPcCL0AMONNjFhFXAYtk3EYjSYX9m3E3y
6/Ipnw+NHCRR2hfi6KBP2SmNl3I+8Bju6yawfTTcefrCP05iNDFBWJijY9Dcg9NwrRlCvW1u8I2O
AOdkPsSFd2ZnqELBP5FG+4mo0O5wMZoL4tlIQR9RoS+NNyLX9LyoBnYBLE8+oekqzjXnsVFBQFtV
l7IfLRl5XgCBu4i6oqyUuuaUX4RlrEryXJ6DN3adOwdTYVdBfG0x+w2woOLcvrsuMAIYVVC+DciZ
bYWxfbJ/NCDGtYunox79YLvBqmjSHm7vad2PUSz7Xx/9SG2X6b/CioKurMMT9bPVQR9RkONV7ved
e5TTtFD04nV5Geq52M3Nr6RMcV27yP3ndFwUbATnVMfZRIP6xStuEMu1KgKYByKvqrJHfb/xQ9af
iaP4WSMornYM5cjXXpNT2z7+fcALzFJBZf8I87tD9SGgOWi8qLJCmXxUz4R60PLM3sj3NgKA0nz1
szrgm2VDBejxvPf+HqPNLzoOLqtfl1jNCpHFekaFjUSIGS1g9EbT15ki0wcumIJItoCASkevVM/w
eLx3FFVNIHL1qkkjxXyQQo7PtTFaOXU8UR6KMUbvM7vmpACdl6C55oiUcRmWCa0z0+tmwGb/UiWk
sEx06/abVAf2PJqG35nCK/wg+Ym9lw0tzgq10OLEU2fEI+L6KPo3pQPAifwlo//RUhJPH8dNniE4
7gH0MukweTTOOMcDOJnqF1Gz1ugxoKwYJyIcp8kOZJBvonlsSI+Ad/qkpCoqNtQ9pzAKmhzEtIIh
8UqkHDGtpmhjbGMQybsSkg5dmmHb540q2ldsEHPx6OK+ceelgrXDU0TRPV4qsqwUQSxQCRPdb+M/
p0kR/zmw+GDQZL6376H13/sGvSx6lEAModkHosx3UfOpcdxq4EEk/ICimmY5hwqIpdxYqqjWg/cc
lQ9PNcwb0gq+A90bW28Xed2ZVzZqfTDeOqpRP0F/qTHSdhnKOqC8BLIuv6LZMUThIq43K5suvyQc
qYzVuxIhdN/Uhz7Q099mG/hMraA8nQV+w73gua76sEYhgYco++nVvPEDkMQ+FrygVvytB0o9pesT
OUEfGx5OudQSviaXZHRLWDap/j8/WNL2wdb2jdqOe+3xA/bxW3l2Wz3XegSIfgGROAyk2nOh4E03
VKsV/zvTBO4QpJD0m6wmcXb5IL/6G/47qvESmG7gDzQ38pzeOpULTTzSDSoM19yGxOKFq4CrDbs5
DBPm19AJ81V+AVqV1J5MrTRRW1T8HWXseGRENrBn8SzUVFZLQSQVo2Grr9LNEnwmo1txH0xPjsBO
3QcSmji85sUIrermga0qysrvn6MNHPTWv0ltKIVIrAHC3WANH3jvH5PiPwnMuU1pP0DMp5IPeDQQ
vrEKz658HxhoNdNmuYbNVV3VLCyh3hhevCgw8HK4cVP683cQg3q8RzxH3kJM8pyVpNSHym0B+oLi
SYgvxnrwsx2LqH3gA3fb0aqBcW+3BIsMiHKOL/yyZ9TKzmjlE4dhoYSd6FNu7WwQ1VG6fb1YJDiY
omqS1SG6YWDK4B6KxgAcljylE1uOVt9riRheAJ+xYKFzlGLZWpAqZR4x5t2PtUyh5lNHKKDc0uHC
cqg8YAgrXVKvVnwJDMywPrST9SrlZ17gqSd59UziVRSyiCASKn4rJ91zY1sRww8yr0h26InzTe5w
J+c0vzmaLtc3BvywnFi9/ugQNNLx97PVQk7u7z06Syy5I10hhvAmU3fN10TXzJe0U/N8rJ7fakT/
ZBf3Vv0cZ8bfLrekChbqM9y6XDa8XneQ4Gg3l0YaWqDFPksQmMDDB0OrU/nLH9fNTyYd7r18XVs8
yu7KXkr886hbuJ44+USbBqKPZ3QLSoawbPVR+5Cdf7HKuM3LQP8rja06TR5Fjk6ChgbUrFMjF10H
yQA6JpkoyBELrWqqJyaECwTtX1JIw0/xyO3QwS+SHlJmm1XY2YhC8pkPy1DoCrUmCj8P6IAsVe1E
hTqFEjfOOJNnTK57PFLs8q0fkA8qMoEkWrEKDcNC8Dl168TsCRFKxAqHfVLls5CSQz7c1LSH/upQ
ew3IahamXTlTgheXKFDkNql6mZsSgrEG5TS7hFurs+7rFciEBaIVB7NJHnVBBefNdOknyBafVOdG
dbro7zkIsToBXlMufidrBeOw1t8U4OKHP3QH/xjZtWJoY+5SbWXT8sxgq45zh5h5cTv/+v4h1rMb
dRlniyocJWftk1QiW+2e7kJMMTcQ63fsGVuaAMcvliPH42BPGu0I7YJwwyflSf4GUWgwhl+03SCH
Fb1+S99n2rjCAt6ny/JnEHE++eHh9DTJWzChkzMwPSU8Vko1uzmWZU5xQqBjNxoS4U7sga4vRHop
tuBQQsADEEJjnB1/adWiNM3ofwgbFiiAiG2y4/oeIYiTt0DazsP3Rhy3wT1ccVqMc7FNHire3VXJ
xn/l0ZqkkcE6ZtLRSD+N24U3xim2B6Et+yXTMs0zcJSFwuq9bpeiVn5osuWoJXKZXpEeBSobmq4+
5XJqppGUhM/zCZ2gxradqD5vNv0dMgpPxRVXIc0G2auGFwFXZdVELg/LUCP07DFtYGi1wfq9karK
eDB3ToYyCPJfX5TgL5kJYKWYlOk+em0rhyHIvOOR68A5cPJNhjuf/8r4+ivzWBnCJB4ajVvwswP1
y6dDL80I9jQFdC8sTRVZPZKWo2eD3S+ROAsaj4iCGzmtoKmWMGAPRhp+iYCICqZO5wa5ZoAVrp7E
fanTlVg161ne1JW2X76udM58YP2yU/f0Jjulj+WtYOxcBYYISXsSNfUL7j6dvjAK2F+AnbWbbDCz
HnFlj7/TRxGVy/xRReGTus+g7pYe3hrn12Diu/96+O6mZwhyb+2TsVNRQ1iQPWzULi8mrrsrjAUN
ZaOreChzKFNGszcInIh+xriTlcXdaJmeLaLc0HK7PiEIQNmB9RLg07Ui1bhJpSh2WkzSj14yoby/
90uWid2vUkKswRKuo9DLfke3qwZ/DaTMvzTipHEIMOGDk9twuzEHJRqBdO3lss4sU74c+hak3k4v
5pzxBenAnbvl10Hb/8ZOnCwFVJ5to2PwMygCmoCf+abU/uPQyCLjj3dmXY+6idDm5lqOI7OHNAtC
7JyQvJ5WIN+t8tbXkkSS+HUrRm+xY9HbXLBYTs1yKWFlCN56OgmlxxoVw3cuUCDFl1Lh5KXpqzN2
dTKcTTDS+vwsHnHWSjA2GLTk+96bfJ3ksHqafaxMfpvWsGJhBkJmXwdgx6LbBz1le7sCmknpZSYp
riwzr6nuAhz4OgQiaQo7k9ykse8O6Yf/GPvRMXOLl5sRpY/jpHGmWdsKgaqpazEFG6DAq7eTPAwQ
wp0N6VuhgzywyfkW43gWhbwAg9mBHSWJHbyFhpGV/hRd0H/EjlavowE6b0STqlHTHmrL+6XCSxoS
p8+eqLgVdtQSAa4u5acekozu2+aSXZQFsEjvtzaoHDC8yaxxC3TUzCCLW51l7SkHBnKBxqe+iuu1
zbDqBI0LtB0U8pWkBXxpIenYwout8iGObIeUvW1LlRQta6GjnLGClk+EibbW2Sc0klj3aFNm7Aiq
UWTczvlRfp4O5aqotzrGIAjK157PNB5P4AxcdrpR81z3lgpoeXZwRhLQ7p1wWB9a+VdRXHKC/1tg
kezfxlKXW27zXKWZ3M6EMXeOkwq2xGae+XnNutIZ8LjFBzxSbIQ8uNKfeADP/FaGbhu4UtUGWvRr
QSr5rFivu3ZrGoqO2X1RyRBLn6vjNPXi2ikm+lrN6o2gfR3fnBAlbQvYtHI26CO3hOz4p7QLYUXK
hWrKhBn/A3waKU3z80cvsht0OPFw1jFbgiTtoxTpum91ZLnO7Gtrb1Qk8HxELSmAw9ForLirrLlI
im/sFrQOYz/o/WboCNGrYo99UwrQ/6aImz0PdYFNWduk4u+W396YhKvunL2RU5j1WwFCaIQ0j2ev
LEn9WSo36F1f0S82N9Iw5BU3xzyBv9v6pFSSYIPH5fvFKJpJmY++olBhckvDFcotblFAM5PsWtE4
2q7JKKNbs/ZNIeVO2EQFGpaAj6wfI5tv2VkOtwM9DtShqFv4l0eS8X13c4/OQPDuNJycKlg3JWGD
wGXPMivPOzuG09RwVAun/eBHcRNYkt8xIKGannTxJLGaE4XdoL7VZOIOq6jGbmb7Xo/+tufcfuCm
7wJyQGu3wHtqinm7cvPmV951yBAFOMFxKsrLR3k0p6eLxvf8NQbCOO8Y46k+I2DD7aQoQdJZQ9+F
MRT5aRM0JIijvra5dYZpqt44CQGREfghPWXu9b1hzEe+VX8Pm/rU5lRX9A2uUP0VcrlpAG6EtFn9
3KSWREPhwtcqiNJoqqVeAFoZLJCAOpFV39BR15RKO7+4iAGERWSiV+Cf+kFyr/Lhs3w4/f9vtcC2
pi6OIzVjJmccGrt8Y+6xAwH7RfNz8FMn4e0W3jKr1CGW4obOuaa+mM1Apx+hZLukwnNWntZd1h+c
GpLduwsvq9eL8MUp6kEgpkerDTC/+jy4zCpof4f9hnfMCLWQZU6w0GiOVTDmHAwmO79Lk/4rjVNm
4Hdse9oIgynptm3VSszDStNlr4YdE8AtQXrgYJ+fZYwQaaa0wWj1rHnv7aPhLSB2cYjiM/Ka2TP8
4lTiOeJXz46CHKtrRcz1Ig9xLatfohAhqvFcaucLzbiOYXpHE8UPsIcA7cej52nDCANzccvyvQjz
0SS+A/zzzyHjowDvGZBl/OqiVYO5PDMGwmxv9VjbKJSL2QL130fTaOCE04edSHv1s4chSvmWP8FX
zAS2lgAW+kSNnz3UD1CkIslxUlLx3BLYS8JQi2P3Ni6JRcKf26GDm3P/k/IbvJToZmYSXf+7wUgA
TiahN8QB1PM+2DG1bwCj33A/iDLT80u1JOYsqESqQkhfSfmJr5SNaTDjeaOw548UBU320TufELsu
xijlojgdAFd8l+C0h0jBwfiJL/0vf3ywuKledds3/dPBlUsPtKSNPFdFf9mZWKEzpwMJYXNUvoR9
k6KsMwELiEs4HxOZkrvuVfh9QTqko3WYWGcWDltGpXjpEI/XjYxbBBGnexhb8RWY4w+6VODvLZGh
HDeh67GhEm9ic5ZvNaeuzU4Dbwoae/U2Sg8hGkUpwt8UM17ajwOzWtC8KikO+lo4YhvmK+BzGFY1
Nzor+6pM8/I906rCtzlOfmFr9l43udiip2c+GEfCMR7sey3yOFVrUdnjCQfwGn2+WejcLHPNq0tq
QnoUmMQ4swhxvlTzRmKTDT6jiYEAhv0PDSZccP9NaNGoVYXK8qBY3q1wcMsnnf597F3Rh0IXbklC
7oa+TKzg/gKJiqyCTUPDYrM6mEbzgbFETfzEa/P6BYQrpcETlO3TqFdjX3nzmUqGg4RXTWEQmzMq
9xn5Y2aPCDQcVFgFvO69MXaYB9+W8kFH2d3OIn4MYxXeTAZW585ja5998hiJhsk0UJ+huQoNiPYS
LrauZXtS4qo/7twU9T9VOY21SftmZ5dqvPAjDrMVF2ZS+Fe2o1UoziL4QYeud3Q+C5C04Z2/q+5E
YYkDHnBp2JFJvjrGcmvL6m478lcfHrelqs+dXsNX49yAkgmL96w5RMFLsAh3iwJpO6OBaIWFrPCE
KU6V6moUSV5SrnqE2DCAgKVbNvZgkCtiEmu0L6L9x2vZtzgYGI1GZcpjPVAQZjL5iSUzK8e038eH
RVz6uDt8islPAfw/U9tDCAd9/iYZ3hjMCN58VZgMTm694qVFNLr0w0nqNlIQcCi+yWacB9BSiOAC
7+ts8NABxwS8OIcQIqycVWHelM2txdRTJoTtAG1Ca2+e1WcA9SIS0qnNp8V7jGudOHuzST1mdDnh
tEEQTBH/TRYnpHKNigtWioJRv0Pyjh0LFNFS7KqyK8qD6ZD8B2fcwNFNxsAIiRWYIGNLlHJY8ZAm
pInBv1ePe84FjW0OzbXeYTXMAxmDQRI8McXhVvp1GhQCnSHIxG0y2P5aGi5yCQNUCdzHteKQy23A
YoB8POuI5pPktGxj1NdnisMVUdfXAIHBMNyEt6PrwgweAtg56ivtioyDHdrMsgq+K8fpTvnspR2r
d5G4PLFYOym0Sa379Lw5b/vD3QoCwB36A7QkB/eJTYLzcd49mSSAs2j6cVN86i6MT8crRPVphs+b
taVEq+9Smz3pMwNEMx3+1bQtatpZFiKVSenvaioRvOW8Y+TyZwEq/VwsdGGhCZA0A/D4B2JX+Ovu
4N4anCd9uJZWIVF9q2rqpnhN+IosVyeZnLUi7rDOTzwKJ3zo/FMC0DsDYOyQs9WE3WWkV6IxP6Kj
5rS6U+BjE7Ky76PqHLGS8fd6w7GQ9Lxq7nRgC20AHm+G4SBqBj2ikp0FTRAhccJ5HY7/YGJWDrcK
7ErVSY1gxhjTmvWslwHmT4VmfVugyzglwcn6IVvC/JmWzpyJiOujKE7UJREziUmOJDemLE4R/xz8
zVK3QQ0fZEEaUfv/wUhXQZHAhE7rzPh+ZxD9EUwDyXUVskTdresdFJRfwdaZehpLduBE4+5KKbnn
95fj2VUxd2lxG4sCkMUqofq3lMm/nf7gVPkw8l8oRJhhwwj43KbfFiIsnIZJm6qRz04YuDR75sWB
Pm1QoeBWaheBCU+5uakGB14eQ3N+hDMTwqamQ0Bx2aInjCDqoH3BdyCurYRVyjpe4n6j5qwetkPN
ZCAx3QuujujpiBmPrPrkZaVGpBFVGSN7ZQieKpRWstT8yNcbDGh45870ST0pQ+AMPMBDgQCsykbR
NgNAqbfAuC7xv++kzOkMUgEtG1l8K1Ob0gRnyMrxNKRX9+09+KyaLWAIoiufuRR/C6iplOG3ez6D
VxbPubOUGYxnysZAuouOiexEto0uKNo1DoUUSF/02vkWyNeu3/3y5SWDAftryeSNONoYAmNJkWbf
AaEJCng6KnWYs6wszbBgx9k5huj4KeFUD/nlwU07dynIjQEyDItw2+F7G2x5Ff8XSJUcUyfLNddg
rIngnjmEsC4Ls+NXBkJR1sGFgZgnHyOoJPmpWFdsgdl89ecWFvAHs+Is0Gc36QlXRojnZp6/UqOU
qyyKDw0qDP4WB4c9/A6bni7+xOx+zHs1poqVD94/h957TKr5Xy2HL6pwWtGDBTNe+XSWpOqFgaED
hwCcJE98zZSthA4VRmYl5cuhMl1SFqSatOI1yIZhL3FkTO8B6M2BduYJI0Vd8kL6TivjlSXSEiSW
h4h7LfsarNsZOredOfQHybPYvJAsieYv5CSBdHxwxPbzh8kawuxxAxNCvMpigID7SFa78Qjn9v3+
BeVg6CMPta559UKY/5p37uXLhcauQ8AmENF8bK6p9M/t+VP6tih6oXcQbtIEBZ0vaMldxIrKJfbR
noDrvumVvAlGFAB2cBlNABtPviZryEtsN7u4+ZwKahRYN7C8q6vo57GQSl6cRnKrijMMvsUbEwib
JOgEYjoG6G1A42Oufrx+h2onMIqaX4IdIHaUqW9jxOyii3grk5BAP2iZx9WSLDgsUevpkodi7TVD
ul3GVWucqKAUsWjpdGL0yWMEA8EJWWbluhLHGmBPvM14iSNa8DW8LAKPGzt1OD1fPbay2dR7L58F
6mL3YRqNyzLYxQNm+QFzuB11SkOtRQSzfySIX0RPbTdU1c5MSVyXRkgAfGeH0nmbeTkXqopmrRan
GnMgTIe4RIeU8zK0XPKWQxI6EPUsKaZYshm7narGUuE2l3rBY5sJZjr+j3yc8VSd7VT23jEa2D1T
3EySDY8DgFiyTyCES622h2hHEzOQHrr4ydm3hmqhIW6jjgYhrzkjTEjYFzZynK4nxQM86bCrvr9i
RVsOzAVPl/wO0RI2rWX/ZAs7Pjv6OcsgJh8vuxmiAURxutznJkwbp4Ed4M/qWhSVnfThTJRFDiRS
RdzXmvhVQ2FOkOTR3S1ZPW6rLeES7oFI5x0ILtEUOEf5d+3CApoGW3u3/NkzchC14pyEWHTEdIvC
qV43jdelFOG0yI5FjDDUNs7kvJP06N2WMWdsdFkFlGinSwLYlBw67EfvLzvPtjOagVz/ywFkKSrC
aTnPEmirES+BmJbSCHVcO9gCIqheekRz10qnhUAe84TJDPECx6WRKjWBKIOMjyEMPr/CfPJJN1lA
MG2wxYUynWIJbeIpd532b/PYn+radI4dnweNrtWyPZxSQlNMoljTNruBkN5NciBR+j0yYwnEXcew
k/oPWBMMWdwwaFafNpNhXCCbsJiErS/YuTcv0LJsDGFELY6FkUmbWeYM26uPKPb/LFympxggpmlX
SXsoZZDSu4ZlM93lZ00KQ3Vk/H4vZNjNSpR87+jFc6vXPP3qt72Q1vabkciG6Iboz5udi1VLqys1
YSCJ9e2oT+hHx+BVnWSnp/73wSqcGQ4YZKrOLfzHNoCGDN55k9OHQKrqDUJ9KbyniPXqj+ju0IXf
SYKIUelLxu0q15DnhHIn6g/XpQmzx2wuRvNq7GvZbVIK0t3l0tSsWO1QIMO+jIK6Yjm+CuCiNEFr
YCBNRqZSzXBLflxV0dxJhHh3MwySj0TuJ8kwnm4NsIP0CmmwhArbR77tRVqzC+3Q9M3oqnuIXOck
2HFpH4HXCqSC8RDAsaIRWwpTvxx75+y+1aBVUiyqWmy65fnqMHgDi43wsNwnUVDqNnO4GAUP1UVg
luExzM/t7iaT8tpV9JOIPaQ2FEDKHAoyDaDbPLQgcQ1DimXSZuqWsKmnG3xovmz8FQr3+zRi0wAF
HWZXzYGRyHZx0b9Pnf6k+UA9NRha56jkMTuWdUq+0Q5plm0I4Sw0IIPjF4HblV45AjaEJoO23Oc3
l3gGPEV6KHTOb2LMPvJV4mirAV25p/AvmjG/Y04xaOEHASyFhm/KBO8abb0RCFP9F1HFEBCLdyOc
ES18/56nHRRD3lYzuFWs/2FVNlHNg4r38E7EW2VFDs5uXbxkmH9plV7OLM8YxHU5Jw6GoO/u/E+r
LSOBWS92ATSYeDUZ4UaPDwHpuDOlBwidbJykwixB2CZO/xRacaHg3N5SH/AOQ9AQV+cCatcfbZTv
S8fFKyzhH45qKdnWN4uhrlJItVvGBqkG38VlUQZtOt5YV3k36TWZD8OkqXQj42rHOD2rLZAPrwv4
HVESzG1q2GiwVGz9kaN+v0ApzJzH4FZKpYHYKrUi0P5prv4Fnwslwx2wCCeWXLWcaFZbKE/xqNYf
Wxv7C+eBmAkS/h9mWt5qJc6X7oWJQRnGuyyWH9HUWU41DGcfMHubwQyz7ticlfmlDFPVzYSks6BD
GYo0h8msHr4W3GwPLlpzIFjqBddeJbahXi/pX93ejpp3rOcikbkMnhqkUVz8V4x165azrEv7eJys
Gvc8q1YaxZUauq/MihYfE1X25TBrtwXYK8G1R66PacDm5Y9k/henVY+FOn/2gawDbTLWk7e8GXFe
Sg8gmPBA+XRD21Opzw0KVnn0AztgAxlqDFGEBKBJRvCarBT1PgDSFHdDvk1qPHg+uVTE+wGa7UMR
4LOJhRkLCk9b2eAkSYAcPqf3XcVIf0g030NMYSUl6f7hNFHI3CSduMW2pCwqxfnVQoW/3iqEgV1y
agYM/jBtHRKKvjW7AjWGmrEgOa5uJwkNG6V89AqY3Vp0JyLd+W8bkPQN5XQOt/7pBaAPdb9B6Jtd
k9Z4Nlmfi5xEPuYdq/HBDrAvwYS6KBHwqdTNkfj0JsGLBw7RAIAo8LmUX6tP+WeDJfqhgvJkmLsG
0v1pGK+Zs1RLGgSEeFI8bUOOy0VX3M9ncCNvR4mKmDdJ+YgpnSjfci2WyB/HHZwf4aWx5jQUJsyL
pC+JkTUeZXpSzLAsrH2jjg0pV5sU012xir9Q3lDhV4UP75rQ2rlSPWTZPM9Ur8iDk/GNw4Q0WDok
m1l+A64JALac/4T8mvk6Y6jGFf2Dh2fW7WIWlj64DqqusupVoBBVNGrWuyLjfqaPuwc268VOxttD
SrMW7rBbno0eszh/y+907kGDYJHaetsfSs2pU3VJ2hZe9b6hLIX6NeYOAgDCxbXFzd3I7QAdPEhS
AXXf3JwlCdVMHsvtZ/iCdNy/T7R45psapOxIeYP9GP7xXjxvq7dXYUl+ICe8gl8RAojJbrTcPNBJ
01b97voXGn6pQGkHa2BfQWzCvU/mJJq6CEDV8rEmjQ177oLIVGoXoKwESepvg25zglZlmRWvHhYE
asXR1tvK8UVPb/dZxj1QN8QuFTQ5qBoBBYO3BJDyt4o8giXlgtLeTyc+hQpothkCpNBLu0R6O0p8
WQwlSeIB6zgIGE8jl5ytBy9cqLgVX+EUZPeTnBcIBNJbnDjG11DIR9CdIVrmDkBIMjH9hknyupU5
gVUj68TOjfcOqbRzV9SCuUTcmFhVJ1a+kfOBf1bN0X1fZXs5aeaNJ3DsMuB3N7X5t445ZF/0az3n
BF2IytGwVI1FGPi1U6+NkWl1RCeyQcYHX4fQszPcNZOXhuYXKr2Q//gfZQgiMApiX1iW7fzQJDl8
TrqoWO1H4Ys4YgCdXm9yLtwJruJj/DJIh2PeFGbdV6Kd0zoX2wyDizua4ZyDtJWDEJIUul29IIHt
IdM3y0JehFmU9HPk3l8mr/uWnLBy8qT8qAZ69JOB5a72Pbbtxm1QvJXI+VmDviTYNbfT2Qe+w2hC
bByvnhLPdSG+gjHLY79y97xK9LfBFMtlFnmnmumS2OGqF/oM2eb0/P6bhskRQJn8fjNIkabZaazo
EVPIK7XC23bWDxCXchFG748BeQ5GaWn5cjADxJxFsN0YgyCvDnGXUYtj8wfqBTK4yZN5DgJH5XOe
83c7YKm0XfmptQfEpLG1/NtJ5wDkkd8Oj0sFCVsxoM39AYmN5Pek/8qCa3pYmvx9qGn5Gez6uJvr
RTFzLGYtzzegHUCESBjbWaocmc0QRYfRj8jX2XKBaD56BI0Q60ImjCnrwsrBKSMLcWupQH6LZS4k
3/jYlckxg7pu2dUqifWnJaRgNN/DJe+tqb226PE9jsSM96gxD72JyeOnMvy8UQUiLdKUl5MzSlQh
AXcHTCvrzCfGnFz/TrOLvF9ZcurYP64OUfxQirkfOevz2t1tSrOIHy86zHpgq/EYjRUc+dywObKL
01mjLjzSJ9pNFdo97MjcCpa5xEcDIIgR3NUjOK6OJ0t7pbRMKS5ImcxL0MoLdHr67yckEi5mhlDG
N/de2LNpCiMEJJJ04TmxhgoRJXgybXvNWQTrW7TVgok88xdhIn3i6Mqt/KcimK5h5tDmJzW8gdux
DDfUyhwKdiOHjLbysMGlsSOSXowVQdqvhXP+0HxjeX5Fvz/MzU2MMdPqKYBQNeo882v0GKTmaaov
MtsMXrqAG9P4fIu6ute3GTTqHDEGaIZG/tJJkzzgLSo9BFw5HFykRZPYYPXn56oFslQ7A4G3oJJV
dl6du/lulOdx3dqKeF7MhXV8IVRJaUMiabKLwil52MXtZFCBWC4/cY3tuX815r8RgOIas0PkL3I+
QsyIei/7BotsOO44TxSviRq0HH88QocSIPpUpvkwjJLjv9ydY7K7itVkPS/OnhK8nhBLhPAtY86p
YCpQFR/FXNVrxDLs9ERXyphIGh0uRMKaxfHHLw18YeKbwV0+qnuQFhev70w+yZXWszZe5hjPjTkj
/XeB9PiWQtdVU/9gwNHU+r0Eh8zWziD2OUBUYEzozl+h5mfIo9HNzSqpxR0tMTUCzIjqnYSgD9sR
ra2ZgWETTK7ER/GXluWx58yAV8kCTRYVSP+HXmIEViG/Pm2XjhuPyI9LHfCsLI3T0+o8rF9uBWJQ
vH/JzNzOj/0DTXUMLVcDjA4drPJRCN7tDd+x3hc4fVRrOu44ep/keDJ6C1gMwhKShEUA+wWFD+7u
03/Pzzlk9C5/BfzXKJG1WFjuespkQjjbafJrQCVQXm8sdom4OSwmLee/JBUlwvO9jJIcpDk7kcGw
x/9DoKVPJJW8mGBFOVH5TZaUYhwsMy9gUivLIHcFNpaCOHNr96VWDROj2/GWf4PgEMw+bPEmt8xa
bdoAtDN01aySjMnHkO11IPRxKe9ZnaNrpV8DOF02/Jy3+f9vq3rl+/edEgSKKRO/7+EhClS2C0Pz
mqQ5rtzRluxEJJ8EeHG4VSUDIOTKAbpOuGF2NHuvAQo0YSEcPu2ERC4FWWIei/q6sBIa23sh3oyZ
9oTSqbe1ha/IUr3LvAsWZcZy0QrGzS5vxoswazwP5haMesORXu2KfPSLg9opSMIYrQLwwva71XA1
AmYIEPbRGZHnZKkXt3tasYJC0hVN8f+qW/uL/G8ztMqnU8PeW3e9V4Dv+hJrcgO8iLj2xItsC2+1
0gcDGmE11a0VVvUs+089Yk++j7k8bHdN4pkgYeOdIhWdGHs87l19Y9X0V/69Ek4xzpPQkpUygieu
yliGfW63xvVITKt/V/qpZCHGz1NANQn7fL5+0YI8kOCBFTGTy7oFrE66cW4lWMfrd5j5jtPqhL9T
9ZLwMvn6Vaii65jk3L9LSgPq8a1ZJhaZLuXKDi+YLn1eO9eXuuh6FGMrVwzOScmtuub5mqxERK0z
SLk2FoOtiTMymSfzCd5UvznRgH6nh8ICs0pxymhj1kYGpfLwZjIvAQIHCRkkHFCfbZIQqLCJTZZZ
4ihiwdl1Pupm9X/hY03IJ1M1OtJcP5AsrgxpKdyFuzT0kYIbwJ64+XUX/gf1YT5tgTxNTeH7mGNU
TwisUxSdvBmwHOE72X1pj/QS4Ll7mUFYbccmTZGlX9sC0GPKhAlO8zzJwlkbYsgTJTBR18xeP+K/
hMpsHMu2pfQWKcNEbVYchQZt+R0TEa5Htbwgg3iQirAKUKZw+ZcAExFnhQjilQxbOf1XPWEFj/15
v9Xy0AxecCx+R6to8+ltp3ADGOqa2qAwRpvly5nob+SwecyFSBiBa9Dt2s7gfHFy0MIrOP2aUgLs
rC8h2m+8ntUQDQ1HksiftkMYw5sHKSQYL8lMuolfMgcs8PxaYLNsgzqRQssIt19CCHKRF58ZhKAm
4juDuL91X6chup4k266OTCO3orkUyku+73lsHbn5Wvb2o1SL0sQidjfnPBnjY/gZuZp1pAa/6XtT
TypbRQ/XNDyiuMS6MlWhgCpxl51avRTIBDK7ywjxVZc8j8JGB+UFlQeci//pFeTPut3xjqIoLVZF
DB/yzu/MxblH/b5blgrG6/Ril2ftNq6m1QywZu/CvjLy0QkmHgIixS221kDR/hs+znm+gpaTI9lN
A5rbmlmWW9xhmRW5WwTyqg+V+72xwSLLu8eVQjHoPfLy7aaj86POarQlcOoDYDf+KbrOdVddyCuv
oeGY+41zwV/yhTCyi51PTeXeE153AcGHsohln1QE/O0wqvFKlYGnZsIuxbKSGWPH3mpYERqP6MgO
m1rxBkUSdiucJpXgqfrQd6FNiA1qKKYNz3brwe6VmQVdjjZClqU0001K7P28D4uZUT8oz64LX3jU
QZ2ZrvT68A/8ta/z4OHM0Jo8qmNZ2p3PPbOPHL6oZkmxZYsyi0VnQ2kW6R6MyA5EizfqnANyEX+5
Dc8xFSXEO2C3xGNuezoo58Q7XcRZaowEaHbOJmxigIrJcXBqxE+stVFxqT7SVTJ1BTCZWqpeTQBa
jcmgwFXETukNLCqQ9mPkHuVsZ6++m3GD4BiWunP7IONsI/2pcWo97wUdsaZCIvD4Pb0B/GKR4wfP
Nrqst8CJRcd2Xt/1CE6UNUb6Tuc0vHzJKbZyzs7VdQpmOzodBnEkfNZuc0g5JbdTV4dZbWcrVHE6
2kWPeLGHum8z8g80o9Hbq4pm8IlTqzAH55P0UL9K4l8mA9eA2pW3D9pKJtvQdQZecddbAd09ZKdD
/1Z45PpE5KNOSCKcbubPwO7h5nHPajFFlOv4JYWAnneFuM3AUM2pbfPFN+7Obf5I0m/30M0CynrJ
pAVhOzCqrNj2jJUNejXOtsxoDLE9nr9eoGjwQSQV/dnXlua3b71iGLQDOQC/NokGFfl9LzqmO2jD
l2Lo8Ws7De/iJeUmYXJlh1z8OUM4Sj4T+qmSKit5o2rAhNiOs0HWVsga2M5AHoMZUlkWtGfli1Jq
d67Q9NPcD8/eIWUKzItqQkl6BqzhhUFiDGrdSZXc1Uv7mI6J8Sn32oz708qeL53dh91Sst9hxsQ7
StqPGWpBS1wHVzswL+UqxV7ADXqEWnzd+V18QDjk/8/gICokHaYrI3y4CXytMCd6FhniTa47a+Kx
VSjiBZLEg41/i5Wei3R5nWN903GE0a7H8MzY2EMwxD2G7VfIcNF+lwpuCPpN9wB9HqgPEwp5Yu9a
m+ZsXVOfZZOIwZN70mbMjfEbj1YSIGy5XC4yO7INysDs/MSabj/AqA5Mx+zipWPM6EFH4h+LM6ap
cfv/nQ7D4f7EY5gTopWBz2ltMIz7EfXo+fxARiKSPOuks9KfNuMla9z1HK7lOtZ+UelkHElsx2s8
SNEfueKXdbMRU2E9zOlMCEZptYCeq6mkSmJNk/BGzsBSQy4Ww/6E3ZQuZjB8wmKxfif88g9c4ZeK
g5kXyNG34pijqnpKTL8xMIcqqAq7pTXWaSz+Zbu34EuDEDiaPA0AtuBD5axvgL0MRslAsg/T9NxE
sgHxRG+OCfknHBDmyOyQZC9GP0iNw2slycQRyLYpw+Bw+X/Yhp4mE/f905TqucTmTwpFiKA+xAGq
vbJUToBXsXauM3iNDceNLbGrMwAGcj+tVRicIRjpqtkV+icKtJbr+Tkl0wOmhcP7ImFvPe9ozWwh
P1Hp54ENScppzwZDyZBaA/XMHOZTmhQFTcp5Ags6WQ5zI+khNog0D5Bcp4swPwohxq7CC8X2524f
iI0MC7TVTmXH2dHIV25MGCAjXq1X8Rgg75MX4bj6seaWWXfUic9raVOCZ9cftWjeCge4AYTc6Wv2
Ok9Dq18vwTZTGujBUyWNwNa/NsvBBlduTXSzHnYWMDxj/aKF48jC7+e5QCbc1LwPX19YMC0laqst
x9+hAfQWUvxTaHxqgblctigxMK1K28k37ZDF/vWMRaiJcKnceQm3G6+PUFWwUK1xnfrtknH/VLvw
6xpmwy9vpyBiD5MauudT8otLEwITqqLhTgZ0pzY194cFahIoeeXaC7Z/g29t/Tmgzg4RuLWQRS4P
R4qLAE6ikFyvk0yBGJriw2F6z10izY2AyUXqIa4Os/AH4UwT7C1gqYt9e7KMVgL0x0MrS3xnGJrp
k9Exi5sCG+ISIsc+LntlHyBLomjuxA7KWJyUdUkgzx2tpzjVTk98iCMjxFgLMbOznEHc3vq/p1Bb
ZjTZIaVyG7ENl5CZp9aOnxu+k07SLKfyQLgYRv4eGcSCKZl66Qq5hvHn9pSsKAA0Wzc0/QZJqWjE
XAvfVVVsCBS39bgx/IlgmCABHQyTe++DB+vWwufzqufz3y7wkyMdaaflrYnE4rap0mF9aw+Xu+oS
BpUjmKSXEV8x9QUvKDlm0peSdufxYsP1V92qJPAGXcHe92m+uxG/i3+bkN7hHrF5t57V3mVo+QPg
QxGgCckDnwGSYQXEhBn1if6YjCFjvDtcSJUF2X01Xmr3sKRkqCcoz9QfWR2NMJKDc9qsGTrUGKqp
vwtZN8LyBRhVslQV91xP9dC0KID8qcfOGjYI8WHDfMMWmDasGtBmwj2EfbTo1f4M/HdTDLgcrn6f
0yFXSgnYfwoCdHj0ChalZti+blxYW+WT2kIZh5jKvn0puEJoMK8ov52GzdJ4H7FanekReT/MALP9
+e/K4zypOnPUpy//WCeN/3UDYdH3Dh7d39ZRAQCv4lyOyuQz7AQOQSkkJXbfoMNvqwnzsiBfGkoZ
13VCfnnOHldUwZU9BDsS/zfn60qdH+snCg2QP7614lO9vBkpBbt+5r9sft4tXZTqKzHiWrTkM1aE
vGdt1giaP7vdhXccr6TvOU3pbNfl0+bi8LkjrkausubHzKwGq/IPLkqZfNUUeeMoOwZolUbIwuw0
5zzB3R9+gCWzZut2eyiBoTrMOJKArT3SzXJt6ZXzl+KE+sdnDNzH2wiKwDPHvOHl2aifJxVBiezd
58Q3TO2ofEWEw2pejVW9IQ5UyMG29W3xUPCvpuP0RywTR4iN//SqWdGteCRCQ8jQRccnmm1Z5IA6
IvTSGzrwYgaUkvJt2ijgWUKN6kYpI0fw9JVRgZVh/L3/C5qi2imM4J4se4e033SLFsWewn2NgJ/G
rFTuxwiZ7Inefk0YBJlCtwRNRXceB+V/kSpjL+BXExMUBUDdFg8iQ+IvFc3AnpNoSVQH/76L9xIN
KRh/LdzwtwzA/t2nzU+eFfg90fUllaTsUkOH0eH6TbRHpIVKHktOIKGYhAQKv3ImKaKsiiyU11rm
n3cno5uMhG0tuM7NiolrQitZOIAw3rtrQJJdXKFH33gYNabiDmqbfVkVCIdpdV5vFvNEvvyW+ci5
pXjPh5XJ85hvTwkkXSov6KawH6vs9gy8VG+4wQHlzbLsE2zjURM8Fbi6f0hg3l0sHcJuDyfn+IX6
Ig+9HZcvKeh0VEcndkYQYes9rqyD2dUr0YHQqJla13a6/rhDlbw0n1DDxuVoWAbk7hWYjLIEArH7
jLWnjWX3xQ/bQAHLZ+AXJ8tYG04suqoalXJ3pdXKF5DRYr8RpG3uoeEYnBtLAMZQn9+IY5NgKjZI
7xxPxw0zaUtFVHVcLsm6ZVEvkVO5IxSBP9EGedL1AV55IH1OPaah9/9NcLjPZgOrYxJcAbiV7N8L
4LdLHUL2MguFVcCjLnYKTV6ZWg7bK5Fq0UjQuZtLQOvNSjb9SJ7ZUwH5zkLXaMQ02LTmNWUBtxNc
6cDPUlsrs5aSiGfpQrqdLCO+d3EpnzCzpiASboU48BvXfUak+ia4U8dmC2Yr+fstPSILJWbbt6A4
UsWpMM+Jrt1tO+fo1wFL2kn+CNx8bjsgc/uMEzAZy0Ub3w8V3ifgAskFyeWwlRKbDPvNj1+q2H9M
nsF91DDHAUevRluZV3FXw9UK/rV5IQadPboH4MFQnXgAD2T2uoQvDc+bfMpy1tMRYuf7EjtweoUf
MtNVM+nxDQWezYRikpPS1mZjbJBBqiAJCAVYdi2mjcXCg9P1Nu9Aay9IBFOLLT+TAWZChGJqno+a
Uusi0YiMhUuNmONc1q6WkYPSq7xsy75OizG25GN23dpB0e0dNjS4lvGd/gqHmeuvZZfKaV42j476
IljN57mClR3Kh+daHNRwQ4DWqCHILi0/3QXUQBPlPwVZzroGnNb1+mvpl7qdfBwmvi+PSe7FRNA8
JURaMLZXyTPFYqxrExLHQG/RdzOxR4fOgIj71+XKNVT0vUlrL//GxfKc81HoHS4ovqm5lMkNiEZV
DR3f5UhSL+juVqM+SJuRB7H8oitWE2xexPUq1kk9NA+1hxZcoILKpS81m9XEedsKubJiwf+cWXjV
gkxcU54vLV+Ukr76y1oGKcSjEG1mfqxpxXPkRnAI0yd649Et7rQx2RHw7ruvmb+SXX0hWzNYJQl1
j5OmvRJ0I3nOIk1z6loVZagm8pBgDHJXcwBDxqHndFqsZlcPuvOrE0XmpGLFNTyPmzM+k9HGiwRG
N4t8aI4wwp+xqQ/xmZR4hJ5SmIg+eY90Xf9eRaDt0B/4vljRL18O4gT5g/KN1R0dSsDJY9qwcyHG
2K5c4Hb8vUCSii36umdGuzwJmCm7/Rn4OUvZKGDahSyW2LiP7YZZo/SiwwhJXJFsoYL9h2bUiqBI
7Cda7c5N7mhmNs02Ya0YLosgkKwAV/9A+ke74RQtI1NTu6L+nRhrPSZF9doMyurjtvAMd9Ng2tOH
hS6qiwsRc41VL3T1kz4PnC4apQPJvFarRmhWfw7C0N7S6B5orittCYHojbqXWyFGH21wjhp5U1cQ
q/oyRCa0E9RzNVZ+OuQdOTjJ+MnMC3f2CP7HxjOwdbUKDaIHfddc+2cgP7sioAtLQeU6UFQaHt2q
rvWnJiEskWyc1wgiTclOrt5I0Ly1lzL9JjxVpSezghoj3F6AObA1sKDcj3VMTPVekZymP8CGhOrh
Vx3ZeutqrRYIPuZuYV2SJE+dnBEaXrl3YBicsQBwqTeTW9b9w+tpqoc2LMDP1UuAfSTiaXZvBhtx
M+m54pV+Z0AYKqvwlb8+zg9TFctf4osJUSHAZXyXmzLCIboZJ90lEyoS1QkC6Mt1WtG3sH6noBTM
7AklvKE8HJEuZvOyzDBld1G/ebQEvuPoIVYIJMV3lpOcfVbHNlyevHJh3S5wgaatr0fn0L5qNh5q
HO3gdL2c4LCNLodI2eQbzmZeohnFpcljqt9ZxaRZ1EzkqeFU7HCVegHSQUU5HSZeO9fvyjK5nXvG
iawzYw1IoRQFQCBvbqr6MdHRyn7swxqF3j9rV0WZ1bbLPSfPoAFdkuc8suOfowpuusnQ1AEMOQ0t
LB/kXoyD+GfLuNoDu7ODr9Lxd+g+IVepeSbCq0+wh+IoPrj3LIKOCpVPKvWxLJ7P2SgltTGTn6sF
XrZlG9S4ytOpe6y3Js7N4i1S3k7PVW4Hap6ubQvKA4Qd3h0oViaIUJHXyLeW1ypGcq+DtgrFJrqL
uklP2rAOUly1pkYamahX3snrX0earrdQJLlXiRnh3/wl1ifTW0zu7zXEdATlfnCw7lme+ooDb9pc
alAPOlLMyVWgmF27lRuS/hAUiZ0QhqfimR3rUBn7Eas3jGyDAvN3brYAEZ2VLejkWh8Wfk+ogAG4
cmV0gEhLHuHI56QB7oXkkO4R+4TAeogeza7R3isGQ3mkRM+GQI7ZpTWzLfrCH0xr6jjuxMaZn8BE
pF2YfE2VVe8xVycD9VOr3bGYohNVaSX6dirw1PMfBt21um3h/2xyNprPgkLjSofzzOMmjace45MB
V9DdH5n3RGKo+m/rDEhuIUj6Q9Di50F0bo92DOrQ5UMKQ1aNxp8kLRKZ/Pauvt7oBLCKyQXzPNxg
y0u/2WjzT1GxQwbb/rCkjapJCVf+J4xTdOHEha3nxoJZ9V/hnjjBMzLnapdcEO8BXDBPeXCEl0vx
XXP8RFG234ajgDakxy+kbFkZ+ZaWMyVToKP3kDk+6JbrSIW8GZ+5mT18qn4OgcYuF4Q1yGo4ESS7
gxPG/4KAgRhlw4hbUIeojOhDOZ7s/CM+MR5ITRwR37WSChg0UxHFhBm8HFSznYyq8kFv/20qBwbg
BW+jzkXf2eNb7qwbRDCSwiWlPWVn9/AyjzQLB4lU86VMyqcByyDClf1NNZ5c/7/M4liUkXfYYwi+
3eJS50DLpUwFT+VjR+kdmkr9LqmdWIWEtfCd3QNYBFzCjPlid4Y/OpQDfNu0bF8sjEWCxEQ64rXD
GRxdTNI3zjSQwfFwoBwzGOZY5ex0NikeU5ZHzT/zGa+2bSMyXeG7UAByiP412lAsXzqRetaww3f8
u/cl1j0pjdso4s+bTa89FyD4OW6//eUnntPzaflblZdRW02h9B5jQib/thEY9IO7FYs0Y92yULQ2
4L27GlFZOBa69BbJ+3spNIA6iGS7duSb0XOKkdDnUwslQkVWxDbLlGjn5OwFoB7OVIzGozaMW8ZB
JVpgZnnJpQsXQLHJGl99CUTdFPdr1BelhQrZsmixJjAR5V+bM/Aw2E8I4LJKn9bw5e+QoTPtER0o
/PIAddBnXXYVhG/18kWvz+FneIDkidQWaCo97s5FycJyox1InnwxLYDLftb2f9ycbLJ/b3Xls8My
AwW7+iWapKTE8SuevrXG3RtiPejq6Von5VdzLOESbgoAtsBYKx2mJHe1qzOC9hhehGFmKqgrmvnv
JEdtXFkFp/24s7RnCp2Ar3B93YTmxwU5LiH+LVnhGjM7/JCT8j4/KCxhcqocuZGbDj/KdHC6CqNq
iR/ouBWW+geDlA47Azb9md376We8Su5+S8kDr56j1XqUsRLgzOyBqB4NCwPeQHwPmZBYHa7o/x8g
0yPpu9XtdpaFssodBr4EU/fENDBnamL2qR0otJWzQqf2zLa3NfP3RF+J7/3auhqCaVT1Wy7jLbqO
BP5qyKquaiMTCRirWWjrXY58Ya3jiWRSJgCC9o9h/6efRIzMIMKDvgEbqq7fxdM0czOU7izNgvrB
nes3z59j47YK+8qDYyWn2cNBfpFK6UlYUmDOHCzBgLmfCa5fVCBsJ5ww6iqbfU2MCHOGVmefqVK1
tJPKd7YI2JUS8WymBGAaUmKFABNqI/wJhJkw1Yy0/LkUKiiWLZNlziodK9KEvzXsXVXzqoS49f3C
8Kj33rsIa38da0SZvgt8YwjM8LPuxLs6m4dY00DxLFiJPDgZkLgET6RHHpbkkwi+3LNNbvL5/5Uu
0I9/G3hzknKdSYTGcUqXx8xfWyvHzR3pnVEAJu8zJDvVIU8fqjGRu1EqtOTDUp8xeQT1SpE5gqQL
A00jjdGIuhcSjzAypHE7fYFb9+csaHbGywNfgy8QZa6U5X5AV1WQqePwXUnM2mtyc4eYpoYx5u71
GKlSCeNljRLEUvKNIBomOX+shdJp8ND9vTn1WGLaR0MRsV9w9PSXXyuwFIWDBC4MaL5Jjd/FOkhN
XfLFqsu4OWXyiwGdve8gUZk13VfUFfN2sTBiRhQrzOMAC8Qr9gOuafQjxKErjvzH+oTvAjGw0oCH
IOUpyZL1+RsINAbXCYqUhroYAjWmjgbT7FvmsOjCzqrGyp6dwgE7CkB5bwwDSi2fra2lXqJojKrw
FN2C7J1Bs09mJmckDLvnKFZ+DZJu5YGX2oLTQ1RCANR5C1TTwLj0fk1qjlikUWb+BzjWU0DNhF9e
NZEx1HlXsT3tydrxu6sUjcrewnKwGb6xqfSTal5Cgyxzs66C4fZkIhoXeU5SamXPh6wN6ciNVPCL
Ly1/sVs5GZe+ruZQW/hbgE7ErHHJNl0SVhoFVYDF65yUk9ML+g+n2CWVbjlLdeQaD5DKpbyayPFV
RipG4sZ0x8XUM5B/2jp4kTSH4MSNb6+YcP9FyGap7jzEStkkssc7MhM2jEwJNewxGgG+cMQIPp39
tCopNicXl5c5GqFXWgItB0U7qEI1gWjj2aLJJKcoAVg1iUv0OWV9FbwHCTq4G+aVFAGtVicqDkbb
58dyXqPEh8Z5FTDL5vnOTao8NjWt/AuWXHaTxmmyjpMg7UOSl4897/5eJZTPbZGRmRnKGhv6eKAP
zZ+vZN5RN/ho0BGmwzBhWWDJjxFHpbvi9Qo0M5sKPXQC671JDsqq0Zs2QWdF6HL43NcVR3XE4SH6
tGTESUt3iuGRR1PGNAVgyhsAgYTX2hzzH2zSN+rd3jjv0C3UrDtixOY+IU24t5Mpkt64YEaBZQ8N
FQYSQke4I10ihGazV2BA/QunLUwnsshTk22xbZEeLVXri+iLdJREJZ0Q8K9UKisogWpv0p1wlvxI
K7T0TciaoxsTtuvFpRebBjpc2/WniCIECVB7LN0hRczubqCdiIbHcs3UU+nfbGNzlHzcUEmbCAHx
e6ecEOoLlNFkyZbgjaRPowNlsUk2mP+XKHFqlk/3BggjTtnehcCb9iUTLfDb4CYNayotYVPMjwxI
LJyzBY6AXM9jCvx/HvSIXpbzgbu/lW00VygHqSDhyl+fCKf/pokL9zPnzq8am4Mws3Ja8bTdClzE
ydww5lQgamVuRqqxIhWHEGigCbfE1lPSolX7wTp77g3UeLBLuKx4HEUbhJQMLnR1puZLGg5WHoVw
AABwAc+EGeHwO4pGUuIbDy55xcSgKGdfk5gFS4opwq8aCxOghxwtpoWfkcEwQ6WGsH7cTtPTnq2v
RpHrmQA+8xjgL7dwpPdRU/gaAzTUjy+z4mGnCgrctGKtT/QOA0qim2hSUSrJolkIkFL9i5ZYA/xl
ZMIDCuwUbn3lYoMfEEiU5qgvUK/k1cSklGyvsccqLUWZpmcu7IdMPSdUbPKAkZKvXKS0PF7319QY
naAZDdVdhdeOX9o6buS3JMhJsb/hUX7sZOhv4VJeOm8HmNM5j6k2mWOxdTB9l2NO8nMz7AHccXmb
shDabIzzcfd0Wyz4bLGvq8qHvde3v4mLYj1QEf07GZf2MCQ0kscQLXQJ7bHJGTNCGyOJXtCWqzdM
34gu0d/iwMvKV1bx5ikv/rR476V5EPuLCvW9Ps+7B81ej+cIw7AKh+ZrmQg3iICIY5oY/z8e98Jj
SWwTaww5fROfi+xVmEnXI4BG/OpInEtG2fXUqNKBl0+/El02mDzY8GCNgJFVZtYkwFFx20aZD07+
Sz92oykuuFkaEKnqOSj7ykaEdk+YB7nZa4ltUkhbZ15IoRpIldTG8YYtaqZpMdqRFHKr6lDwx6ik
9C4UUhCuAb8dVlWwZ0BKJ0oLN4khptBE5ERE14OK4RvLpHMHu0dl/WcAurZD5PRNdoZP+u+CukEQ
hBIcocS+4CBuZNsn4623cTa2QHePYfPAtEN35VDcpe+CI8JZHYmdWGpBhrepcVTn20VndbsYooMh
HaHLdeuYqkKIImn+87XMJTmL9E6VXvHnXjW0RxB1K0CIyFdgfb4mbUO9h4pR9Q22pKeP3TTWVD51
lB1HN4dJzfX4vPWEzy8e5U25Tb1BW2S4o0HFNSBQZ3856Jzx2qY3Z9YyltLjju/hSUK9uBhhKC2E
4WrosiRLlDIvbSw3jVtVkkYYcv0kG/Py4DJc03RC387NM9NGAgGPQ711geyQPl8+vnYClrauVvVU
4mDRiPDTIfq1jiTRqT4hu3gDgSJH2Gx36hCY7+0sx1SEM6D5beuzh5duBIQMTblfLvBdY5J/FDAf
ImC/EuwQG3JBlOK1Q6mNLkcbVBoozfS9GNeU93I3OIPX84PUA/ctSISC+ND8e6+vsIlQzhCP5cIO
aJ9pD90nyvOY0t+WIS/UKMBGL3hUG9KzgoI99didV5wSe9ggAmI+md4Yt1grLep47otPuTXNFu9g
r381pFyvDaaG7YlqdV0ncvqQ2bN6ZZ8h7BOPuvWuLZIsY8jdpTgCnK4XBq3U7YI/YCcVJ9CEP8Qn
zBDBYv2vnTflVgFBDjgzrutzXdMu4+4vhsgUTzzZK8thypjWSdYyMFBjm29OE3oDlelQUXF20eA2
0tlrCPyuuPx0/fslRpcwEaBz/TboUIoAq9Kno5Ab6XqGC8LYCT8xUdRprUK3FIrIBU3VQLe61w5E
Sa8uhtI6J26XyPgoRLy8jLIWKgEyCmr9OmjNVJPsH0i0o/s00jy8rNg1yEgFioZIcxCS/SHqDeZm
vm69wGiR6RdtcCBIAyitCi2sNE10IiZUUItr3Tgo60xpJi3MjTHXXcsDKEDd7aK28kZIRXAq4g3W
n0Ipc1YbF/P6xaimtxNGvemaAO/eKsmtwtpJOZIM6V+nA1HqxHBYd6UgWLiX3j+ibCnwtV80at/q
X5al74UKBByUooFpmpgYeMCdPgF9dGi3Ju/zwx8OhF7xONJcNKRX6TEUZltaN1W7VNh2Xj/MsSVo
DU4Hn3qFp2Uw5maJo3u8/AD2nz+6RZ5dPvfrtM7YnSE7lCiiLqpga4p2Xf1hj03+4U0I8ht0pE7Y
FLbIGBEBGKZdl44yV6mX6gY1lfbA5JEMuwQt/PHpppD2/7jCG+tudUulf5f34UU3DaQmrYOqGURZ
p7mkmefc26jDuB8sz0WyoNKdm7V+pPGMya3bC/0oKn71eDtFSPyBFCG/YX32bM5CsWL1zUHNOU5v
sK2dDsCg+kyyLhtL6ahkfWvYoh+e/VUVSd2GMRFBgVKjbtn8Jxlnx1VFBL+9G3JADpYZVmdr6K/Y
blPFGhFyuyhRMNaOcgdIyLBq3kA/+lRzyU6l1gahfT1/46XZlBYnRTYoifPNP+4SvjEDXcrnkVxr
ejQ//ho7+T0Ac0kFrdeFOP7MVmJvcr/M+0i2iWy9z8PCs9g4bCETmcZOZCVNJqWjhSqapje0gAwD
ssS1a0nL9PagiOYnEw4czLPXf0aTIAi2V+2oiDNPQpU/KVg6NnYYJjGEaosZ0le6nT7C4fVGvlTe
RmFMCGhnvavBuer0nTkNBfPCrCPvqsuIMQmUNAwqEmxg1f5O2SkQw7dzaI/XDYKKI2qkfiUHE4l/
lurzpsNfEZi0qaHkaaNv3sQJQFVeL6oulF0gFVLadh2vmk7f+LLOxfR3f6VIMifrrasrVvrMwuxj
oiO3MFEGKk7lasYzoEd91uU5SHCnSBgWbvzaQHn2zVoi6Fvwp7U19vqbDZlClPXqK1FMf790QBcV
+CXcgbh3mee4FOqDJj4A4rqggU+b9WXgaSLQUrHXilfsNU5GTFwLjDe9mXh/bgKPiiaM2wLlWZwl
Dpm8AaypYxpdBg9Tat7FMiOI298NT9Jluqv48MFoGokobTjwTyEf/MXgPaC5p0IjYHRCSWVo4miM
08lbYUoWWpzYe49h6Iz1yLbeCfgSHd3kbBpkXs/IWR1S4V1N+hm/zktmuFmIiom7U62ldU6Vnkax
7aLKOGCdBMxC1BuUuZAbw2qq75rOwU0ZGMfcnv44XVCgiOMce7zGDRSXShaWaNFgy0NzyLovXVln
al1o/hLc4jQPkaJ68oCxYok/yPFjsQn8rRzYNmdTuGUdeHc+9urnRnR1pMEdQfiqNx067jbb0cYE
7zxYLurbeFfJpRoQ24RlSp4NWXkOOqG/IPivRcy9EJlPOzMOEkrmbPRLTibcQbOPfswmTr9ov6mr
y1F24GBKmuB6EDmdnkY9FrHgUAS801gj5SblO5GOOv2pIyukRhUS3OwVesEEYQNNf/uLIX885geE
ZrN+eKd8zTm9ai74E/VpFoXjXOuqT+CpSil+aYaqub2ea8OKlYWW0R2Is0mw0Q2Ij0vviSQs+Env
bIPsggkpN+kN0J7ns1aj6UWoq7YcJdB0SmE3XAwc4KzWeYfHsfSjw+iBCZlYTA4Jowd/pqzCDq+a
IshoWxtiOxxFC5353eK8s0wOkYpmMlKOATxpcM0P4sLAank18OmbS63PE44lxpuh7785fxYWkYyS
LEMe7TSpEbERY1vnk25Em4mSG72nT6SgfhDp0fINZwCEt1qCkRpLcg7DmVqiMNUWCOp/gvQreZbt
jLRdcdgPllvm9yro2ke4eGiZobq0w8ocLQcdmWqmUbtu6HSncO+Bf8X3wVebudo8MRSTBxwK2GBY
hGztL2vIiYIzMlvTli5J8rRxH+/IeG+fS4QGZ5Iah7SqD/y/D8IiRJLv/kjA3IqG7yGCYGPedNFQ
4U4UejA/i62yiddIPHGBWlWP2AVbusiX1JTZXjtwQNMSMQ5Eju5FnZGwHlsCl4YEqYIdKSY/QTgB
KxlEuGkxAS8HmQhD3UANJUvirBLmmk/lm2K0xdCV5wG8g4SsF5NE12ZO+PLP53IvTNzEg0R3dBYs
lqcu10kQDcUEmXsM7fjNe9yDkPHfFjhwhdHIJxPuKi+3yzS4zk6e6l8zzsN2FBlFUCIdSVT0JatN
vyxxaNxra9lb+vvjPcBU+Aa12dZ/RMwIbCUW6La42GMHluXkACeDH0ujvrLU21RtGgKtpgJCEjil
NBad8HZED2gJ0mURRhzC2eO/47/UPYnrPOar5NjYcMDQXMDSREiwTGCJuaepgMHxPhJjQxvwrRJW
b2XYHDL2Vvxd+GRZFLNCNFLYQ47MZ6Scg4hoBc8VpG3V5RA+gNAjDtcmNDQXAov3YpmxhwaxULrA
wnGD513A/QjRZPGoGd3TK3yRBxnlxRxMAs3taIMh36HByERF79qaYDXxQ+XSa2m35r5mfmKjdIr8
92gWkdvABzjwLJShe3WevL5fW74/3aqLnXkW7NoqaMvG3s9Bbg7Je9jls/g6m/W+mZlD2KS3ttmM
Z5fP5pYVXlpWyzX2vws1d1ROJkmISNtbaWlhJWKKVF41lQjzs5KjFY2rr1Bj0S8cyKqHkg6zCXlj
oJ6TGFSa2bUMBuTw7JycTjbzm/5y9TNs9qsm1BIepRDyIv26C9RMHL1nH2Q4b6nxJGJBiE5/KHaL
SMPW8iFEmPXVm/6bduVpXELTuWoAlP4BWdMywWStn8fptFcU0S12urD4Eykhc/nVUlwFITFnchq+
ogs2VQWoscvFeBoTjdtZoA1wZpQ82lXS4K7XyCuIcqZNRXe6cSU3DbfPMoToSE+aU6okaKvM2uvD
0ngD2WHPAfX87iA2l6LPYEQOCmUNkaN80OY/SFLNUp308q4ZCxk6zIKidCB+Sb0hKKkYu2oXCZXb
ISRyvz7IL4WjDW9xyxfYPYVTkTAhv9Ellp1k4NCW+po2KuWqJomaN+79V+bI7dAG6kvJ0hlwkEt4
olFpSKtBnfm5JGrb9fItUDQhQivSQSzssPMyMFSXJFDLK5E7xlA25gv8aJ3CTXHI5hVcCTnMEaIQ
PEUmFTofPItr07a1KW58tmQJ9939HULPoOmfyIYNWimWpNmzsy2XctTQgSOtO8E/lLbfmBajcGQM
X7WC3EVV8h/V0/uyq6DT4JbSG4+4JGrR4gZmkNJknerk1CRgGIXQisADLkJW1QKhS26weQK9B5HU
3TzylJow1UXd6wEys0oosdes0aAKpgHs+se/AcKMyhrjJ9J6bmWvkn/q0fsUvHQRnLXdbnTOkpmR
zx6zh7aUmYibcO7A7GuA6mTrjyRN3nA2FVRMkSjGHKCAavDIuQrmQZwZ4/HCtr884IR5q5Bx3J4D
GdmPEFJ2EEWYQ30uHXcRCQN22DRV9csqFMHTLVPjLqOSyH382P4ncB767wYoy5pjCJqmey48UoD8
0tUTwc+BjmDAIsklexdesr6szK7SLWiEKriLJbk4tPOoWjQVcLTp+flVmfjremPFaMU1RzEOFOi4
UCVooF1z4/KdXdE3AE/f6dl3kO09Om+tmnJVUPuRrU6mAEOk1D37THx3ZF5t1ShfaiW8jxEiBEaA
7l4uBbVNE2XVVvXqIqGHUl/GEyb8K2ZuN36HY3trOdBKQOxSXR9Cn6MUhSl/4X+h1kvrdUr2Q6n5
tFIu9Jt3sjfBJzv4EdFE99LAeM5V3RtrNp795aI3JxCXDF3zqqtQSlEw5RhfREAKO2ocHAUCkjvh
R0ZqzBAkSVrflNGE+cS9p1+2b8tb2icZhOzwPQPG0VUHIn/IJxrZSlLInnNRyJzFZEO8c04Ng77D
MxFqH2m5CuSgoLA+3jyGxTxvqHR3xT9LSILfQWq/deCz68Q285zd5YR/1tuynEMfA3ZPzLIi7aWj
T9Exj5xMh1cvjHx+zbZRiNwsNocGlGAusPjj/5Q0g0pV/k8Qv8j7ATBl6LmJ7a9WwTqYdOQsQk78
dgRMY9aLEWXlw/MWcI3FwRTeQ1hoNEHIF4jB5dEDoYN0rbjaE92952Abywa3LF/7cD2cnaD5YJEG
33tZYoixI/PPKLYZT29wQXa85ipojltZ+WxhF344LmbX0MdLa5HH4QG4uS9F5xdZHEEeQtvxl3EK
iotr+drv6p2NDocBXXiarJ9x4Mg9P8Wl345XvgR8PJG7tKpKPTDWwplKObt3yE54Hm2gyx1PUm6p
0oyJuaW4SflhHE1IobX+8yk10oI/qev3xWPhTXgJbfVY1SaUDXcY8apsTcUiTXSAxe/n5X4/U52Q
LQCVST6LhUeEDDpgxp/Xpy0pLHENt3arvyu8J2DwUIoByOCTSgdY/O2R0sleDasdzuHIEvCWHyif
t0eaLY5fPScKNwWYLIH5AmX1NNevy9GHHr2bDHRgc7GU7y9JWVJ21+OzTeUyBMft6IullYw1z6Cy
GRMWYXxPx7RSUV4+X1kBq2jUQOzhpgH4WMHGWJPYwJFNP+scvzxvg3BgQOPRyOJWVflUyqvBZFiZ
gTP5dXMsnGyZsXET9hqB5DNSPEvCiGw0L424czpl8I21ehWtc6EucvahFcTKoopybKiUfSojXi/1
mF1YQ4hwBOxCxGTUyRWs5aauKc9FlriODYuVJNdZV9+KoNIKPVuk4PqAZZZ2M0wsCD7jh5JUI8qe
usjro5j/BzNSEr2TwLVcGvQFvUwjiBsE4Stwa+IhONcl00TvRLN6lj78HMK4YJMzPtbdMq8TIT0L
wcrgq4nvC+Afu/HfV+SjcvWffgfcjE1IvAZvgVgFbYju1P2Lc2iWn+EN1jLjpjMmQ1k/VQgQBaSE
diRHwmkgiQSyzebUqijZPpBy+RCmWlXCxVsEtagSUM+278219e6zSIdGpqvRPVOnu62AHsAhYtFi
v6xsXNLQ9dk/JiCQF2sanFrLzhqt2JKg2HLk6GHHYVWVjyjedjMFiFG3U9XQxQ1JE/T29jm9pUl4
WDUwVSkIQHULS8lfgQOSZSfIoCvQsZcv7TsVyVYgGhazy6KRKy3f90lCyG7RSmNVOdQ26pplydYe
/gbQ8mpgWBhuydAcyLaIBRfM6ZcaY+6xvesbBsnSg7BZduF1lpahjXHXHqlWGdrqdgaDfo+tkonU
Zlj8kNDvoa13izbeo76YrxPycIqdDCVqlQKWu41YcgDy7N3hpWrX8WKgjC3I68ShMZrXR6Wwzawk
z02ffF0KNtr6yi46Td1h8zDHheT0SBqNL8plZGnaYkWsXkQpyFTdk6lxMGqgGGEJquCT6tEhI4yd
2xyzOzGHfo9wMzB+oauN6Lnou3vX66BwKQwwzSDI7SIMc0k91rI8XUxuC9+PQ6LilhaqkTVlqvUB
VbfvwznFOwVbz+mh3OJaywbjpHgOzZmC6s45PsdnTXDKakUi7bwiebHsHMOdOuPMNIQpYZ2VMhme
rJKeaQmDlt8SYpZ7M0z+MRwvlyHuBPrRgu+fpSlNTjhl7megNYLEgMy4oH94zRpPcZzQPe/2IufM
TP5LDZZYgil4YfSYWl65M0c05vo1aZx718AixZxLv4SwPkpnKEkordDlMdo3dVKTxcFX/Ii0xqkz
bbsDRC6zcD+GHXzaNslawJal1WEybE5DIOTNBFa/OMRDi5dHdi5mxxY1tgoihYBKXu81VJldAvVy
u3KcrcTtozc6/9k3yqAPq7pWPxmxiXN6XSJYIvsf6yYOjs1zwXm0MrJZCLxJhdHPEhxgAwM904R8
DE9jbmwgwiuocSwVyr7+0WH62UfI0btlOsy3UqbSrJg0UI1G21BKl6jejTJZB9c7dLAeKaOhAwur
lbtnlQ2YuR5v17JenAqJP/Cu5Qzte94SxrTz+Ne/3+NouJ2ThYlh/XokOul/H1O01ITERik3m06c
4YchHLc/qYaPVnmQ/KRc3iOnp9wUsn/CHyAEqqbeovI2hyhf8YnFPWBWtR6tB1QJF96/wGpe/hdU
KnMzjySzbour2XV9MnwqKXXTaqDb1NgMzzgBuYNF/0WEZnL/c6xFLftJVYTZ+p0v4Qq5KlS89DhH
TRiqInO4jHuQihnItlybi6vzSP4fvFknX81mva+4u+jeQ3Zss5x7id7N9i3rJQ2M742zXgTH91mC
AmTIilXAzB0ihcpe6JSZvau2a3uoIM6WfpnqzpgWDFT1KmWon/LHsuza2ttP14ueRqJ6tu9IC4Q6
jCB1e0A/fmj/QnpnDyz81Akse/B5Q6M9DE12N5k74p5Fi6cwtWbLdRTdZS4xUqjaWz0CA86ixeqQ
kY5Esj5A5RmO0Tr/12gTtcOW/4cu1M5ZvbYUcOtQJZVvLQlvgg7UJeRmJ9+eiyfyKYkM8G4kvg/F
/tfwP8WJydr7NCfEScaIu9lmS2gXQSVwZC88PseEfR/JbeI2uNTV6XeclUQPvyYpgUSrZfo2JXK6
nbYZGgN6q//xT/D91irYKtygm4KILwHFzVdvHxvUsq22hIIx0EY/mthRCOobhQvVbliBAMXxjH8K
zWR6LXnYKKzdD75H0GOlz8NF1dcWmig3cDL4LOqFG9H6FMB29K/BV2vHAjYp6a2d6bNQV/dTGogu
iUNIBbd6oXsc5Fm/9vOiULcoO+9KR4100ZUUFLQ7mX4mm1beGXdPlz4jDTtWsM3IrqgkN6TMmGbu
mPC/UjY31A7aYYxvSMj91rr5KwNQJ+aS07D/fN7D8G7haRiKdLuVSGFOClF7LOGMYFkgJtZ5VRw0
LO3xyOYJh6qmBnQ0WYCSBkmQp6WUU3iXRNEUzzGbTYBgFnZnz7rAuYGHyori4lyTOKQ3vibiP7O+
cWtjBJRLVz5CHyJ23dR92OkGHJPq0EHeOjyH9YpmYW7VhaaKCDGVhsaF/TTq8LPWqMw55m5zIATN
w6z5JB5iiRnvMYLJeqjZH3+fFYD80Lwj+NMzLEQYGfPuJqPs1dRNsgabVpS0E1x9VvQnvXLoGrIz
yMrkmLJoHjty8ASNVVFUX8qfTDRpz9i+5DIBZbepvSJBwPSy6XN5zohrpTUOXiU4eIU7B5yfNxLN
kbOw7Kd8Dp1UR3wJS/Bt/tOp0Ir3KMRw7w8l1Skr04BEeBFLkKqU5KkNd4X8xgxSH126S5CqRGcp
cIFVZuyedWVMob36TG63ZTb6T5ofEReTxH8VlaWgyLDIrt5IZ7sv582ZdfcSmYaxPqoH/SyaApTx
aBKlIDVqywbJinwkPufBf0gN1pxNhIEm/k4R6+RRSVjBNPcoFTszh0IWvyDvUq2GTLTqoOobNwDS
qQPbeg7R3pmOtUJwv808bWZlN9dms+1og3iYe55//8lZxMkDLVq1SI8SMhzKfqhv/sfxI0sMgScq
4N7ogB2AdzPhXPtBW0Jv6TxM6SEYXtdpCLncdh/+CY9jXpPnJH64pQh3qfRuzApscEV5TZNLKO01
gy62xr0cqbVDGpIspv8qqWCTvtWkle549EL0ug53gGVWpTbGPZ9vyfrgQ6htIdrGDTaeR96am3Zj
tm0v3/dsOa95UKBpXOKrTtWY9M7AaqJ0l3s3EqTz0PGuuRBuPKhPiPkvxii5DwIaNVN+nE6tgkzS
vTOiHDGNZdz9HA+9JQrAdgZq2k9/0pDIXzbxc34pAcjF8MpENHMHNkMew1FcisfqaEGF3208Eo7Y
BCE8iyJzbyI6YMYSLYnjGUIdl9shX+/I/lOVA59NolU27owEL5e6G8KDtcM4hp0OVYoIKibV6J1G
9RyrpRIlLWxTdsuSsTOXq/mQWW4fSb6SQpfSEjz9jHFtFvId7y8JdWKfPE7hy7Ezu4ROIlYCZr1X
AnOv0/tKFoCEpwujf8fcYL3LId7PZV+LKV98OXru5NF2uVsobJdZYRjr/iDbgcBd2XyR1By9jbZo
YhKjsAftAlunmJams5cYvq42j5NjYmXVN8wZe9muJuhxM6Sdm+vegTiqonx9crSIfrr0QXB6wRNQ
mU9/CwfvCe1QXjxMuRPGRyanWyjLEUS8ptCyur7pm8u/l9nU1ZSnUnJ/zeeny0bi8Y+ZCRcy+ply
5me0qBO3hNpqIVBTpy6EMylxtdq6lC/JyQyo6+U+CPqh275HgfrERPY5zUmwtbNJT2ZXaM4OxqMW
Y8l1BsUxgU/BeL8lL9JMHLJ6kQynHP4Wz07JYC1i/Cf37HicRTBk7OdfhlYb7wGI5a0CIlHqhvnL
XjHk3+EaZXQ5+WDzNnJ3LNAmwvm8d+dUN5Cw1ssvBaspvlychU8I5+fS1jlHjLm4N8C9SdTC6FoP
U+LplDUX1mOTyFrvEEel7SmvK/MATFhjGV1GQoG2lSeTdwF21JN1lx3yxvqenxHU0MXjli8onWPX
nEqMk+s2rvx/4OY9pD8rLwVZ1KL/2ZqKumjzWNkoHG8NI8Jp4XPKHxXl/RMEkSweVEawF9/65tU5
gkrSZxdUvITOIfFxSCMm9XjG5QOJXlvS1AOSAMW/IDlB9hXOkqtVtGeZ4MwhhCXfXbJZKlLqUL9L
z5jJTMTwJ7yXyzI502x1hN9EMQqMpZRncW5r8qwTyLBJu43HM16rrGr3i66Xr+fWr7pHufYjOqFb
bSUQRy+2yzy1I+iYAfTFON7R9EmE7uSPLW5d05NllTUv2J3KZ0Rv8gUtj5c/Vb06f51ZPn2pNY+u
paIUSWWha4kklJTGfZ95HMmfyMFehxc0ZmnPDR4kGveplU7al12TRw+kDQAwGVGjKSSl32vqSMzB
NIapFlt7TBfc9XmxkV2hZP39iYU0MHKnEURQ4sUHEVPMjSfoNDFjXsDQPSzASa6nodUaj49DTh2n
9vFtzT+mDSqB/LzWDgAz31GgWu8YmH6eIlX+6eje7HF1T9i6mrhaIQ8lok9n91yfTXOopba4xpI1
D8L2W203nh22thlKu5xzhzpOUs2RFKhyP6pcT3001r0JZcDIrRyIeZtRpsOAPIIi5HuVb4qEGPdE
yg8co9iCJEE0/JiJbPAOvAaDBiUTkkkkaAD6CggCnXFA/C8VGgIIVVHFJehnan+J8C8VIuSjZ5DR
rO0+eumKtNih6ybOXR6SNbGeqmvYe024xF83gtw+aw4OmsE2KLgQho/M6IeCXRoNvh8OL9PiMuUz
t57o+K8beGQtrG8Vf2QOeyZVsjQNNcSjclbT0zfXcaOCAsBIYaPQG6aAyd5HZOeQ87Cqxzxq4yK3
58oK0arKgL5iq41av591bL0QcrR7ygn4ktIalKYO837Obxsl+WdFtfaNEBvXPHYHpAFd9gR0UQqL
o5QTLY8m50SNlWcnHYVMUh8Vz1SO3OVuTwe7J2GMq3wnqp468giTBXSl8qdlHtql9wleU14YNR2U
EdPDceac9DlgWacKG6jB5DPTsVDPVZ3DgpR3DKkvDoKMBiFyjgL5cDy//PlWkLh4Ml59jyz0a6GM
po5Kgj2H5DzshyLFroaj3lY7hE+anbBMc5Vjorjliw95obBGIU9vda3yB/82Kkt+8ooQAi8guIOF
8Ds94Fx58cE463SVxw2EyiS+cZW9KTriuJKnGA9lHs18HTRfQ9IrpFGhi6G2YNQ0a/GHXjX6RtL2
tMAtLOyI7S7WoYuTIKZ0dSX/g+2iIS0JLLe0GOBhWOQp5HgrukBUe9Kv1Ib6rGN22JzKTvWkPDYM
byGXxRrkM/To81bGNynlYkWwQMr8h9j2f/2qgmRxmjyyFtvdSZt+pYSFjPpPlSdupyf0lDmUHT1i
Ivra8lrE/xw16KPPUhC7Spkpa1qi4Nq4URaXFMv7+uEjANJB5F9Ei0c0OL+mOe1OfVMj0P1DmoZM
0ZKPBR67PZtlVsodHy4XR5graS4PM4w/UlZJO6btL0BeiPSvs+jqq/HXnBul8MybAPndkWlLu6WX
EL1tcCLJDxxBXEbfLPm13InKuht56jpnKespUwHsfKxG1nJx0rsfaDb5ji5QLAdMzDVJ+Lx90TT+
IdxfXtkfB3G8ZN5QiajyKbR4k/ZEQ6DbhsbypkfReZCXoZ2JdQXWDPQH/XkdMhy9eZkeUrMkogR3
5FS0HXe9WsrbrfP3P1kfVOUcobNNX4tnaY+STl39X9Hz6dFP1Pi5FoXvDULmOxRpehIeOiuOvfvM
b6Mdjn5f+w+maHxPAB7s2RvHyGNEJdl1a3yYFd817l8VXwDvOMNS/wFplFe7X+s/gJFVE8pplHZ7
EvTk+9gb3LgrSG6l6DcefDgCMDMBr6Bj85OteFT76+WsQO6eoUBoJ721eqUCKTqIYwF8nfUSu5Mr
c57xwuvRMc7lLvU1HtUJ2LCQOCUztdLihTXx4zXNj2UM/wHJ/7eXXRbtqMTdeDCp24cDkgq4gS1p
0xyfytueYe+n+IpXA1ogrOezSKAg2OWKokA86axhlnjFb/IKzFbXBzC9FRWu6Pag0cztmlXvm8EE
ZANOXnaDFUmJEywGypUidoBMX1Jj+vl5nQyKTxT4PVo5xyANc3lsEvuVyafF1gNAedRGkW39EUFa
rIt1NFWpM4nxUP/jOqcOhcKGjrR34MR+VCv3QmiodzvXVsdUQYkkr8NjiQYcmXrZk+Aq2T3CpJSr
ac89ynXLziHS79p/j3pNq26a31Ho9NczPRy18qfol6RuEkyHl2BA8zEJOYG97+alzwoEm5btkygq
7bcNbR1QgRxlbc0eTZ6eobHbP+5nOhkDZo+EIc7ntaDNA5yKA1cClSNxUSJwtWcKgysRiK70CFA/
6RvlJZXZ+mM9PCpoO567b6rBhQz9pHfcWsN0/P0lfnQFVXN6cBV9fhWC6IjNSgrA41POlpCdmp/k
EVl5CsgT9VBofY9cHCX7jaNR0yUeQ35U6FnVXg4b3YgedZlYlaHDDRZXV8pJy72VHSfEGR8k+PXK
gKq+sosDP2fenLEf8SNUt24hz4u4QIAx/+xAFoQ0beF7WGtzM79pz2TpIKwpNHu+xsj2RcEmWWMH
09N+jxJ0VIQ5NRbSMG6Y5D5dDQM/5k4Zqe4OgUaX5qG7bJwJGl04ugMe7XMw2K0S36Hj2Z1yKPiO
FzH4A0cSL6jgakxrRw6cIZmZ5mZt68INy+HvZqawQ9rehHrccPnxcPoxPQdqmCjoAE15i7QyuSrn
3a33GnPtgZvlW0mxNWe0jB/CurKVPumKyW/B+SXQnZDxPSFP6YBLoqEDFzHfToIyXyqC3/FjyeKG
Cwz38G60XVVyKRdEaPH2LSWrO426TZPfOnrkye2CQ/+G7wjHPwo3hT1/qA1smkE5mapyOMlzc8jE
6RLIaMbGbQf35kor4ZIcvZi05tfczJvwx3pI7x/0XHzoR9pzEQO+C0cOZP20bJRM87JzfIZ3bwn0
+7SVwAIz+fH+DH/QxUm2WX1W+ydgXxSRxVq+Ujk4XIEzjXdMPULFAPMX4ZSbypzYYUmUYvMLPBxB
LASiIQdGZ5UvdUS+E3q7WA/7vCLHxVLXejvOQPQh9Ph9eZ80Gny52k+Zh21p13B5SFKFfesLV89N
djf7HqHEg67KAZSUp6kp/Bo2Lb5kPRAkepvO66OXY6aQgCizBLjly8MmSljrzCM0zkIu9bP3FPuA
1pbqbtOqAcL5QXKAiFej9SFnZD2NdkrqxsFoEEREHOfsWahg5s9OISVAgy2g0n6rGgTTY4dsGBE8
+m03NvuOOFe6LNbVCu+gW2A5tSVJz+D2A2GXVuwQXXHvAsV9RE31WdRITRH51RNp4NZvENclKNKF
ub0To/V1N6t/izwSv9zku7j7svxoYBu5Jnl7uw5wjEUlZ0/1k6jplf6K265Gje27P3cy3RifLqBk
XE09UuKLDjOSxE+EGbVvJIGBgthzaeR7PkMuBExUCLuYj9h+X+9RaT2WndlFgLSWTa657mjLyusG
wuRQtoYPqZIskIFi1IH06cZqAhCO1AExP0dv153u+AbD2Y/ip9WHAwg9NcreztnxRDPk0JB7dOp/
lVYonYTpsQF8gFxi3Lz85lYrv4lkDYfzfbJzkQDRFk1Hx6A13hldh3vNEH6sWeIndH+k4LfGTEtm
/r6kw0Jk2b6BG2bvaEScWu9DoglYAErXwJblS55uo2kwdMY+09SqGO6GEt+WlPKvgVytsh2gLi31
9mq7z55/MvV2ikmXFfUqQ6fZph6PdRS3rEeqZAh6HnGWp/BB+bI296tSN6dczFxVXGa+9jtE7zvn
LETA5f7rYWUltdtv2Qo0ZSkQR9xw7/iM05ZtI+Qh2e9MSuBJS2+rKgSevTOLYuHlxHOwGaOuWibq
2NSOXg9V2onj9ibmyS/G/InG00FzOPpOfeNP2/oE/vev/VwsNUEhlgV8qO4tkLt8sOyg7j7A5e3t
aj6yAOacGnDLBXQtMzfOOnVSMNuDNSXj63OSkSAZqAB2A9B5wsts9BSMs1NY20kk+wc5AP8hQ1tS
rsOpf+x9khe7QXbXfxXkTz0oJ4hasob2+B8cWe9YxVfcSpRhFkj+2zKBeZv8tJ6atvwWTmPmNMVF
uoBr4XKC8vO24Ae136zIp+NdqCm0qwembX+MwCPbxXrCmhaCrjRYnvxfm1ehMMcxFSt8mys6Wep7
VMnk3EoNtlBkKy7dByBkN5Z0ZTB7i/naj+ikEvay86fUOfrtG6bcEC8kyXRnWvO4XIDva3Uvj710
4q6rS5BsedrxHEXJLNmyF4x4GIzU8AN4mRwX0y66dN55eRPAf9QoXW7JMqZJYjSiq6XCzeyQzpUf
GWE1J7Ut+SaEx81Uy5bOzZFFRBwArCwzupwFn0PbMZKn8Lpg+czpYMumza6IgW84jd4TDzeGVXa3
ljz9yo4UnAnRb9Wep3m6fX0NoRac4dZ0+Lz5UUvIYr5FlsjTsgPjn4mBqDku4rWVZKohD5EBtZZU
T2Hit65KZpVn7xogiOEWG4aU1jfdOxDfgRZhYRmfBYkdm3TT4OCwzHUbJRQ8wA4KrdnuBW+n0eKG
yEEidwtcITerqU6cXh04+s+Ar9lF+jOCTfLgp0bamyX49b7lbHIH0wdrgGj7U2ylJDuTWFrUOw/k
7YM3aflc/i3IKF7C/uQQ68pFQpOPNQqD+zVesFjB4xJjtU8Qz+GbdTje+8Jw03d0OiYH1zHyCazQ
Wvp2I8EYDwCFZhxy0HdGliid3fSb147WLo5g8+Uen/6oNeiKs9+IqRW4MtmqxLJuykySObt38t5Y
2XKQbZyCEGigr94jA2pKn9QLLt2egI4lo5ieG0lvgWvUXaMt2JJDGWmJEvBBxqkoX5Df4haY1sTY
FdMQflpkgn9mBbrM1qgTsSTEdWX5S6CkbQ8cMJXHgvYv1mLEcPaiQNttA10B14EsAsmcowQ74RGv
wE1NaJWPZhEd/NROCrzBSSX1+OSxPaCWpCgx1rRHbYxKPNY3Dn7DwBAvuZIQGWqVEoVh3+MzCm8j
toAjAXAiNYbXTJaoP1U4zeOwObp7dDsrvltoXfOadnMM4MAOIn28f1YKPL1XaX7Vr+WHQnSrwwvU
0akIaxJbLAYLNmu+cwXVcocgRAmNfDPxGP0fjAf70Y1SbJAcdhO24rDwKTSCwxC0Njufdu1ci4LJ
ywVLSzKGbygIvPzMYl1IU50JrebHWyEuUGkaEY8QpVYhyftwtCCV1D3Wx/Qk0gpeLT7yuoDm22pW
B9lrtWpCBbT9GGc2jgMC6+6QZV9N++xNpv/FEDuAt0gO2vSK5BAtCfhDREnkL1av23UPr7W/DvA1
+TkhosALn7wJlPOkQmzSQRy3KQMH5JcbL9h9PQE6d9t91CNFATfdckDb2IHoHuZLeP5HNDb2XA+z
33xyKP+Dx8hhNOvVgT/jIoKIzEGpzXIe84cr2OM/ffhcYdwW7MyjnvWP1kpq0TN6wcy5eH59wKAL
PULp+CiJcEuVfXQ0gqyEvUb2Amulej+61MOyr9WrbJVq5bTSy4asK6n11s8vCYZdg+mLuLy2Xvqp
rpXtgbh9AmH1StrOb6ptA0NeSR/7Fbtg/46J7CKwM+JOFMnQu+url4+tZkHOBonUmTpX0BEFnUDa
f9/dbh+P+bi04fmtSbt1JFlAMtPkE9Sx20izsBp1IsU3pE99L+Rv4pJIQ8PcEER301vh6qDej81G
BmR0rfh1l28R9Dzt9qeqKo6k2rXlj5dUrGQMfAKgylhBhqEgA7beK4gonSeXccAVyJho7KBI0Hhn
xMQdah1LxKMWQ+9cNvM7/dcEzwvdtvoqyOkJuG0KvMVyKahj4YjM2nA5NwsFf48BUbwNtugvhbKK
RN2cPiBzn7BbyqY8uUP7mE/tCp1sn86qRksWtKKDDWAcMPEG6ZrVmyNZgu8LLYE1MOyEV6k53fhe
tw5a/BfMvQSZ68JUC+37iB+0WduPXlzAYkH9pMiFHCfQgVWESh9lhTJlTycUzJyzbCrizlxDso+Y
OB0IBnZxbMGz31qdH7Fs++RLcuIdpALTyXYc+UUcAHPHV63A6Q0ugXquFx/JjazIfkk62fCNzfAR
hysd2izwE+LLM3eHHmxBcxQYhjhN47CLHVeUJQwCSgn/UNY+GqpfXqyfuEhh9q+O0TYT71Qb053i
HKO/ZnauY3YvtEqH1oEK2FOrL5kIbzPZYmrG8lmrshlyw54Uw5XlfYPvSpsasIYKFkaJBDq6kqt5
dRWzpcozrD3kIp5TMlRAE86BmX+ZSJPAGzcIsF+WGfZJLUnqsCj7UOG6X8K6GDOTVzpC+WgsX2Ov
UBHg+FZzTtXVyPTyooTGwQp0xG21LAZ3ioSZc8TZquzM163CEZTZ/eYKK65JcuGfx05MneI3eRb8
xNQXnAB5Jv4fUbNXiD/wcpkyoMdMbjf51G065GIV/vqxmoJ3s/pxtElobrMolG43Y1GFFJYfbk8/
XBvZcVyv26FA6EN6WCBwBGXLn8+r1AId7TIBms4XhuklNvtHpgJjNK5VH2OcfbGSTIIJVgFlBt2h
kIRiy2gmpGvB8MKAwbMDcxASeQF2uPHn9XShFpFgh/Lz8SHWe2X9S2a0BPUlQ+d5yVO7YlAQLIbJ
JYoBg7TLHzLjMoY9/LBaPL/+o37VvoPfHZOsbQDmhhdrte+fpkFJff1aoDRL5tO3jQjRDeOrB/Z/
jFMrMEti0iJ9hmQHh0GHtWDAYq/Scbnq59epJGrkKqvlmRbPH6LAHGeFoz0ebN2wSRC0Lx2feSgn
4Rn0RjIqD6hJqQteCwY/r1nurZ6cp695juI2rxRoiaTJjuXpLVd/YAIAL+9iwAWJeyEZwS43HPIH
wPdBWgCci95QCPlSM4upAKNcKeDFroFiAeXV0dCjwCB4byHS9i+GetVWJeZm1rUXuEnvDwZHss89
tuk2NA44kVr6KMK5hZh7LIGiXSg17uqlQCjK5r7LQy6U/amQw0Ya2mcpVSIVvPznr+8CI7N18ygB
FkrGT2OccbWbT1F2K/y4yRBcOz453+dXTx3rZdeGyuSVuZU0yCa8E5qjKWLzmpx67NeswT5uRVBa
mZ4NB+m/eBVgorhqicB9jLNZBvo/m162u0ARNouRNJHGf6bllYjrUC7uoVbmTamvSXpUfwQZXFj3
9ZEcbK0vL0FrOHrQa8Zto36aM2ONeqeNZR8qRaY+63eHQhEaf0mjqcd+5T4P+SPNt+PEfnsMX9nn
/cutXkpFAZjMhXjEn3Y/JjoiT0FQJuNWh/EiraIWc0GsdTDfJlfHjXrA/lUxwM/PEXW51R7QHeGi
KIpusaCtR++rQ5o8dKUgazhfqsGpK/M6bIb62RQMTgZp09bQVBQLeNcHUl8sUojhk/FNdKKkMQD4
Rtxs6y5DkUNuyMM6V98czpSTfOgN7UdJSfc7/Fp/2KPJIG0t+Cr/tN266cxptKLTgOINkawwTbJX
D8vGtbWmMU26PHyVwAGGAAjXsSE6TyiKARcGkVDAaVNwEBkIrLg+VWms5QcXJtflf0JjbBBegcBw
D4zf0BaWtSuRa18sx0b7BSudL7wxPxYc+4WhaDGndgccRY3kpQfgdX7G+iH4UJPb53L7JkOncM5D
n6Yf5NSSJOl3h6/CTNXOEjvj5o/bjgPTYJ/ZjhXpd1qLn3T4o8nLMcJH2zkXnjuBjWCD95uAIB9e
Bqt2eswbF10/w1xo89Qo3uFrlJuH5Y1Jrbe7p2poY5uXFLDBdNQam5dQDrhxIOUIcUiZKXFovkBH
7L3yr10uytu3yLULXsECQVLedbwndB26l+2C1a97ffOP7IQQMSc9zF6LLXWK2jJJs3XU+RY5WbUd
3pmbvQOTnwX07jf+KLlD/l2q3+0FKogR80Ed7tMOU6vneDabDh/MQrLBnss/swN5JrM+pyFndMtj
JqNAfvuoVWyz6OMw9x3z81PE+Upr/uiELWQDarVgORo83R65K3AbDCQbCHZXX+XQf2YqRjrDqPWQ
fjDNwyyOOs8rHrFg2d88Hj8q4Rim/MFlFDLZSJfZL3XR7XfxbyvKzDDPdJjAuDI5HEWde5P5SWL0
QEGtShd3GDNAYMI2k2Pck6ws0XLy09xndjBC3g9X4jiZAZ0I83vejjPKHa5Wc38Xxs58fFJRtbqv
gwAE3aft01eoleBeYJXT55MOUyeJsJaXwoTmep3Muvv5wMU1o/BWJgSSfQgbo6mZoRdSdGhYjvB6
HkozBF+ogIBuVBQ2W6wdziL5KwixziLUEi+nsUqkvy9rl6E9VxdLdDQE6vvpuoTuWVFPOuyQ3O4v
x5d5XzKhx1YApi+Z/gCwKmu/QuI/cQnXzXtaN8N6q3Cwdd3AnnWszXks/wKK1YHGzXH/rWfbw95S
Kj81mePtqbbfb6TCP06WzTFnjB+kuo5K562vyKRoKmrLWMlVWR8olNKsTl3yR0hP0c2z7HPSJwFQ
caNJ6ilIgIy+Rpil7kB+IosP7+Joba3iXjG6sSy+oEZKTT2VxL+E9fTWOfSzKGdkBLYBqTb0BqCc
SjAVZ0f44QuSgPvVsOd8QHIz827pOK4BBZCLZqoE+PvtoWzlLjFyaHWmn02LV89WNdBbVkXH7akm
+i4Qic+r+dTsG6p/iGfiV58hPxG2aQxrt8YLaASko6lV8UREC1XQmTe5E+02VED83wy9Mm0vMs7I
0tvfmTU5Jzh49+LS9ExTzVNcyChLHzCxEO02zQjUpohbmDUR+Nbzwd6JG4wvwAxk8ZEin8EVk6H4
ISQWE74dXMFVdDighB9wAffYyvQ/XhSJw9XA3Whiok8Y3xf+S72D1kNfNyR90icREjCPjRMsBe4+
ALvCh2j57/de2e11k4ge5MzgC0IMISmJ7khDINqHKx5sJlU2YuoOhdV4zx11aif6SMZ/7eow/2iP
W+7IEFBg/owFImErYcOA9CH7U0ih3ENpG8B2hlx1SDbsmzxLaB2OXqFJNO7OR2qZSwBzcvwqtkZJ
YP2ODs88kSnWztCbqM56SCMX70iadrgZ4J9oMa1ycao+DyPFOLzvvkIRw3CTNjWLmCJyZaGh17GW
cT2nSEkpr4zexSfugH/nWZ4V4Dbm9Sa+XYIMwYfSiWHRQ+ElmNqR5j2jj0fHuMsEd5mKccXUv6Lm
d4NnQcUKp/j3SqJ3pJWGjLuYLi+VYQIOpWNDM0H0/p1HWf8XPyOEzC3WRWhJ6hZJjeckNXoWZcTz
eVjPCPtjBrD+9RVAOrOcTGERz8LL9oObVeAFernOSzyVI5cnZw3eD54MrpzUfZGZRcIs2BlikcnB
bMXyukxnBN48rOcviF2rpyax/VHYOjci6xuUTG6wP0+JkOQMzTeOOnPD/YdVtMxFjub6EdjhD6i/
5iOOeIZnhyRvQZBstdgAetPqKkrQuDwnVeenjB3aI21XwEeEKH8JKmhba4JbNVPSP0okQV5Sd4Pu
xAfbH4Rxh8ZdfyJkbB0/vfYryDrvYZ3LlS9NC+oZHLY2y304u014rSzcmKwhhDLYL4Of1Qzacj1b
On+jtVbHYQb84S+mZA6LugpBOVD+afuW0BJ29VwgijGFKpeoDa1k7gKofB0L+WOnbP0K0PTUnC4K
AgrJsRruCD9KR8KTlakwcaLFz9L7bSf495dCGZIkXG8RlPPH5yErq7UH49YJjRPgRDia9xPIXrtk
A8tLfoS7rLpb7kGP3B26GTOuRoGHmxhjJkein8Ul8tVfn9PvQ3NXXJcEADOO1M1ObEllCOT9diZg
DgszhvRfGDnQMJ/juUYCmkkb5sWXdc9dmNrp13OBiHfwHt8Vq60RMPcV3aTz9PJl3C6jFzou/xQt
8ICXLW+qpkroAzTXefURy9DOsM/+hsQrAUN+dFZxFcWbiLZBZJquPLxVKTA4G+vwSq0gjDspgzYV
KpdxkXOAC7Xd1sNa9pabnzXDRsMhfDzyrINzcbkLx/cFJbYSmmmCVdbjdMI8IBa4hjf2j8Fysy0b
AoFdgegk/hHLO5ObB02sydyZp1JUQmelCYxufJVVxi/Xzgi+lIr3aphMDC/CIweXmOCrGKKjWcWC
cWYAWABYjLp03uTb/ypwiNl4gvEdNOok8c0woklM0FPMnSQeNAM0Oj+c8G6/wmqRANthqrRQ6cBb
GvehceIsKhyPY4/Er3muU4T2ntKZSCYGgrCpPZvG5R8e9bB2nmQg2clpk7vUZc7EeWkh8OdOqdAo
rwxJtpbSfcSvSiz9LTeI8ecTo+nB9b2JDK/5sHXhK3yMlYnkMEIlz73dIPxyh7c94VwR68/pyP5s
SsBwVpoLDn6PxpVbMMsz2DdLtImH0FjAJ1xpfa/nu7x840dyEXhEk57O4RAMWlzdRIo1+U7DUiVC
Bbr+eRwAYu2Eq4ykeXaR04HTBRAl3F5MPcWQGlYwhnr5NL3tLhz7VAkA4QfhJtNjivmkfufy48tC
heTNE/2Bcq6Q4AkdWfMry6SQ7+imBv4XkfONM1NWOwfphvjwKdKImkejryMsK3sDpMSQerebzwNv
HPOB7INBL+kBGqHGlHjujNtrIvru2H0cxAU4fa/Nlka6LiQCBqT6F+c8sce+6vxPTIDovR5cBINO
UHsKFUYX7aRN8b5ngTIJvPBbCJaL93wpymBifyxVwLYzeUF2TD46k2tEqefflRSxR1xIR9YEmSsJ
9PqlC8tSdrabQyPB3ivCtcpBNAYXJbPR+tTOD8bx0fRRud4vU5EvYFVpdfr2kPL2b+38AtQpZK8J
McRuKm53TIFMBtnjHbi4z06v563Eb5Ap++DBarXhQYlbr8t5fios2Jn2z5km8mc2aOhpG+9VJVne
p99wgIRMMkiUY6SvJJ55W0UtGQHqL66r2zBf/dYVe5M/1lMQV2M8n4QV5n0I32AD7YZwVevpyDfa
m1N5EngVoObGhEhuHCysZH8rX92W9stgEzGCwAR4NdhUfJWqE+ns1Q4zeNxsPM59YZzT7o71SQva
m1s4F7YihwtNw74YTi9pwKQy8AdRreCVJkLG9Aj/lTsqMzwjMAr5+PiDjUm8+xLIEBRwx0OX2n7i
xbUDUBfPu2cvjJAxpKqyvlEZqeFa7PaV4UILfYnFr28bZQIWbnR3SZ1rMOsp93LIHJLkX9mLFtrs
6Bf0xH2IIpEEYc4nKLTnJUmbP1qiYcDXBEdKEoVYJ47l4H/fGFvdvlLJtfx8PdbXMhsmX1I2p8Zi
j4l08rmBpjw7YtQW2jHZFzexTybxOigxTJ07Y74vsUgybAUIm069OTKdH2YZxDynAY8TuPGZRTv/
UlJR39W7Ynqa6BPOY3qhdiF5M5Sor3w+KiPoiKOjxDIGl+8v5ai7GiE3eWF6MOVpHOtO5gd4KLc/
T5Z+dO6QZo9GvG7CJpWfuPOvuG1Pm3RJip/GTMFO29tVFaKDNAA069HEbw6K6wcItB/kiNXDA0Vk
1Lm9XRHrJIIt1JI8Tb/a1JX+0HjVr7m4OAieDiLU1Y5unz/NlHZOMD1KO1oWEHaivM8OGFvb+X8P
LWAMxAJyuHzECSGqkdTlcfY7vyMvefVuHx3Zoe/db/kemGSv+S1JWas/3tuhOVYfDK18yoFxrYqh
YgmItEsdwd51Hha7NQ7fqOlg7dKed0PFvVahFH9hJAR+iE53bfOlM8ms4W+5TvS4i5soQgtlX6Ym
Zzrr90yMj6MlBtS1uIH7B15juRDSwZEfsgU+Jsay2KgF/20WITW2RxOPx9KZROu7vRe7DuSecnUe
iGHSS7g8UvO6cd5sOVJbcsE2TZfl5LXMdxrteW4cBgHaXOvOzeDC0prpyZLlMUoUiYORWs4rsvwG
RYrrA+ClWzLlCDjOk6dKky63QFeMAtGA85p3C1Cj35wUC6eGoxs+AOSIYmyWRyO3GuDr1q0GoPma
3B/QOCLC0JZg78k1mCKLQLixIdB6/ODZcTRSf6UuVq9kCBzl6mSHhmVrKtTGh+oX++UQ43FNy1pG
zKZKPKRpDzLNpIBnb6zsEg1/Lw2/bxVjDkjdo43Nt07WFeCBUO/qFBwkTF241hdyOA2cUZP6wML/
i7bL/VeHTXPhPxptFOqRFjrZQ8opNZ8zyAAUOH767rPu65WPlop6n6V+N+ohN5n8qwIBoL28RAKd
m+DYeNEfYN8PO4SLM1czycAiUMHv1E3A5FmlDCn9PMuvPH1iBty2KYHxwAamWs980PvMta+PlOzc
otVUzHySTS4YYanvinzfiEHoT66qE/Io6NucZH5aad4lKoDLHtdXQrRQ9EO1eC5h6EPsRMyjJzWp
xkQJ49fnVytBJq6nLdPvhSxZ66JZfnY8lEaPgcSfxomX+rhFAk4r7QUQ0CPNtpFltSQUdbu6oT9u
25rENX07M/qc33mAKKPlsSFN1ERgDJcpXKP+rqBza/diiBjnEuqh/5eGvCHc+Wf1Z5wlFPFBl5Y2
+Uy+QR6Zfjvvq8ruG//NNyEB/vs0pnJRt5EIQP6Nn9N//kDR5OseAoyqzVGhVhZg5pMwMzDxDxf+
+sw858M47ZA2Jg8FM5RX49P2DeDoIuQhcMIVeSDU+UL+MuOTUO/U8s5xeHStHhCJMOnE5ypnVbJH
p6XQbHY3P3LbfHPPwgFkVQBmHcbyshY4ZuUamjv65P/RxUxC1+DrHIo3RDUeOpoe+Ez/RXcC3Lgj
1Tl8jucr5z8OTIrXmNfTBCn/z8mRVPyx3o2Q25kJTJnzqNbCZlQaLJbLBq1i32z+uwjLbmW51Mt5
cwL/7a09he+H1nciT6ifbGhsffmh4GuLLblThGKiU3FF5iDCS8LzT/OBuvuZj3GgYshbGkLlJCr0
cAMjYiUJL1cWHKmKMG5nzzvg31/PwOrU4CG5tJm/By2uvnWDnwu95mtlE85oUd84SlL59XtV1YIu
Lyww6a214Xvmfa+1Xuey56xoaYSHdlcYwW/dEGi6y9CTIb7Gj/7vPA1pM2hAEmzW1lzBqVebPbx0
y/EfwP60Lk2ovnn/pSE/croqdKwpE9EiUKsu9ZpEuAecknoI/3hmT3PJ7u1uSb0iCTuVxNypKiQJ
IaailX1AQXkTSMEbSucLoEfyYOd3vHvDcgnJLb/7vC3SSkuIRi6Mx3mmaerIgt5GMt7tCKbo508u
yYBwETvq/6ZdJu7SswYpR7+dZFreReI/NZB6arARATHAavKGidaMV5Lo8VU6X80/uj16MMDydOho
jrzKWogBg9ysM41a9SczidpaYMOx3Ll/p/UJmBTA17wWhZ19eHUG3PV/cM1kAnd/XiHLfVLaqXVn
xonCtu8xbuqD/yZxiSXBaypc4plpfzy2aKblwLDRPEFilpCQZYZi+KTNyXF+D2Iv3tqjtQc0h8/z
GLDq4I4i0F/syMmW5XS6UTQiYgFPPb4trQPxO6H4HfMS0RgMROjrk+xWmpCzFmHMxadtbWnArqF0
J/X18ffa39DLqYrIoztjYDzkUCjR6MjYqE0HbOmMTjfASMHgLE9KOcBiz79MApLHzQKhguaBYZzT
exfc4RtJeTxVXc8nVWZ3901luzEGwhxl9IDSCu6zf2fkvMPQGPGmXLh3Cm8Y5pTKsD+Tsb0NnniS
eTdEnMHk1rtXv/9jZwHDUR6Mboxc4ksd5peQtr+fcTNJqB7Ia1ugwhmUbdIAqUcku9n5jROxFIJK
Yj40xPtLLGq1b7AEaOwQ0GKvsYFVarPN0vPNXQ+/fhRtde2CXdSmC5trPSVO3UN9uwEEsM+5o2AH
Y1RCebk432lZBx0LZV2kNQE22WaADzw/dh70kfOhX72q8Yx7ZpePznud42I8aJll4ThK6we+ZMz4
NgpKvjX8G7QzR7SNyAkDAsO+/D6k3B4n1034iYieSDjI0DwcpB3e3RkyM3mRXFHT5qSqKD+QVNup
Q6FLIfyYap6QXf3ngoh96axixIgvOHlGO3gnvqg/beFQnb0y1CIgQw+r9cUeHkXJkrG4qHNqVj5J
0gHeZkSDpHZEG/xmClUlIiC6JO0SwM8kazPuraoyG2C477yVSTkZj7vbzC2qA1+4ZpUvJgbNCHHA
0EFhepRg/4RVuHCHIHFiTqfKY7Qog96uPdkW1iU4KY0Je69IvvA4YZrnHFLnKZaE8OMO3+Ug0KYH
NpAsbsOZcprV5bo1/bndu5JoHIVmZIp4Q+T7Cyg4+dIuY4cie+2XJQUatzIFtOQjBgy1jQPCGikf
5I+DVF+M7fYTfH3QspFkNU55jWfjPlrSPd2erqZf1tq9sgZ7kS589JwYWOmGV4HA3TJQdqJ5Ybmq
XDn2ERemMSXpcpbBp74SlbxXamX0TDjvWEOVfbwirX8uIrf6ap5aqEVQo0BpjDI/z02JbeO+zvBC
1fX3tvZ1DtxhMG32rQTUaM5W2FrnnWaRccZsbbouSnzGMeZ2foaej9Fyxmre5Byqul/XTWJJ2LRM
Zpdn0l4/mZkgKUeYOACkzHSsvbIh1zE/6bhRohelNNiKNI12Q4iVoiymynLPuopDSjjPR+He2T/a
iqZHh0/BzRAU2Ak6nW7OYeiram1Nn5Pc4VwVo1PGgxTX23gH0Y0IK825KNJP0lYpIHdALC+uHGkB
eWXRrSp6FQ628WlM7Ds9/hzw+5JeIkrFUcT8NMvnkWL+Opjw6ABV1hh8BetOhOhLIEQcbx1FJLaw
HO7wer/Y5tkxNGhldPWZzPeAi2wEDbRX+XxFmWq+Vv3wVL0SYXBfxfJ4Czs0p7fPCd0KUZflZqJw
sCJFd/bzs7XFutzabk6e29PozgiA+awQIzRwtu9j0+jnXrm2Uvz6/iKhi/jD6Rd46g9piEZkUYWN
m8asvXUlLaf+h4+2O0MQB4DWsWDJNPCAdl1d84jVEg0V8jpUZuu/1GgBeoM8WCMvshT2ELwdpaMq
jUKVrJVAxKyoyKhiy9O3ti3KwZZLnAgZZrPJrqb4D17J//ZcTI4/ZlxkkLrqy7ZPwURuChPIoxkH
UMMcRJvyx84hT37xxe78+F7+fX5osOKrEe386isjdF2e+OfEA8wYEmBo8BT9W9oaUe3geW+zhDR+
xPYoaYIPJMoE7DWMI/AFQU07uh2rvx5ijNn1YqBjuDsQ1YD5//D9ukqXEqyGwsAr3ffZ5Qg9Vwa+
Kv5lQs0T8EJRtv1KPJeYw0GoBjuudnYhY7HnWCIfQo2FLPbhtQvDvrboiIR+L6TlL3FTRxVDGAQw
fCFwbk3mbP+q+O0cWyljmWSCHGByJOQr3fk5A1npSQHgVcyyklbbHlcdrKlD1ZeERqIBorBwGbh6
71TecmEYZW4NFr4rlqIbdUACg6Od0UG/M6+uULqU2V8C3X4KdMmkAIm2zVktrO2EIr1HN+p7IcJJ
a3fwECbQuvwSZS3EcAsjVKgVfXrpuRBqfsamHSUhBL1cVwjI8Qfoj7MGCT8z5M1BQjPMqADDmmiJ
o0XkTgVLKgsNak2gI4XwuCC5d9fDR6eIGxRD4OHBGCOJZ3giNeVlnKj+iB3xP1Feyy3S+Qd/y6Jn
ZKTrMa9tRV3NDFD52LH031QXmunKOEYbGOSDuZkIfyM3cZ4EakP4MdIkfkiZHXQR9d+Vlvco9g+y
+Vlde5Lcp4T2y1pUBpdC4B2sCL/0t6ScG+mbgusuSzEk5Q/je4ib0BHi/yL2oNqTI0JQg7CMe0Xc
/w6UsmXa44m/VuukZtOkNauX/L7uD+WhCCxYl8ui1TAxEiNfi5uzYpFuGvwEZmsI0yNv2yJ4R75P
rosk50H4Lx96n5f1BISTi6xugn/4wzNG2RnXQZywUgtstXtiZZyHiljnlG9LOJwp1k+lNM0ZYO/5
LiBZY32fWHd9I+g5T4OpysmSo+rDzQG2sHmWKUJQsepZG3Wgy+3VN3Zq78txqG6yTjwKGdRdDyR+
kp5mcHg7+Azv/IoUwGiCZq/k8LvJB3zxHa26DlZMVF39O2wodKgEJ+mtgWtN5/E66b83cXXNz4X9
4rdodmkUATPrNQsf9dhKyz9+CxYbTI5bhtcCUmoQD78Z32grUsW2xoZSF1f9n3ysP7aEjaN7FIvH
DzRZF1wP/1ciqLnW2xMUKaGX+SPD1Q2PvB/Xz3G6s+4rUt8PzeI5hxYrdBItq81soAsik79Sv91Z
XkeNa7UzQgudqwGgL5Yt9ty5/Uzmsc2f/bRejzGNBlg97u0H42kmkJUR1ONp0Q9X5TSxEptx8KfR
WS5MCbI7lQW9Y02S9oKaY6MCY7s86lEvJCnhFldYQXjwL3pAxkDxKVzSIvDyvL5eGYSp6RZJNVKw
+iKvCYby38+kqVWHPkI97Bbkub9P57GGF4NvdVyb1oD5tXW+eV3gqBO4wlo46is0f67hefcv0SKv
sTr6CmivYXeXdW31LqMiYmQ303Q+9fSRATi1zdEcrsLEk+w82qmxCEidX2MIV8gXzNKTbiGlRhdq
cfN4/CaxPJRYRPXW6ruCXeRIhJizWGGUIIfnL58Ke1OYaGa35qNO+03/qg/lm+gNxGQX4VsApAXw
mIOQ74dZdkHYH5Tk2C5LyKFyCstiF6lYv6IfwD0isWmdUTsGg6JwFft9D/5VVsX+GUH8Q2Sy7kYx
Gt5CjwhVQehwih83mHGr6QJrRNF8GKuHNG4fJlFugGQGxXZB75ZiyucwjUAcHqF37VMa0i2F2MgG
MUUxw+U+NNW/YreRfjAxCtLfFFc8yPnoxUmu8OWoNBaXvSe+2AgrA/yD39xqgS2XD31POV0Iy2p/
KM9bWAqqOd53oiOcrLhbvqShhE+L2+kWqkHxYML0hkZu5DLX/T8G80lxUSAwkOYn/Racjofa8Hzz
Fs7Oazd1rGcwC/6H65qMNoiRHDFdRTo79o41kHk0bDAi/BTRsxzDRy4XiAIaZ6uqE+lVStL+rfsL
MYZc+PXtQNlWzjGL9W4sywEdpZpifxKu4gWQ/hkaJ2OKIjqDm644UTWTdYdXAmRHOTtmQqSinRWE
/H0c0gsOstVmnHnSBiB/p2iLr0/WSaScmNrVNC2XUJpO+C6erfEYOewko8nDUeg+7OoG9ceecvzr
AS0A8EYIdjQbyGpQF/LCywAFiiUapW/nzuUBkeWQqbXzAydLDnZSm3017FWuMxK8ZIUDv29Jb+NZ
WWujeMk09lzo1RJ3ctzWw11+R8+TPGkSfcQaYlYfE65KLx+AJfqHTnUylgGACbN/66Vy76MOK7MK
7L0dLTLrjojLKSo3t9uX0RmYebQyevO+WfxpOuDFzkstnPpgVV4z7p13XgeRjUM+/jr6kWRKNtYe
67qrMAhoDy2jspWWbTFnN08rg73LCtfEHtsHlxh2/9DL8VhP5kTpDfI41jM7PdHx15Ld+Akn39MV
bcefA+QgP0EryvP+tqoTXhTKhS6KwFdx1xiMhmJ7Ikhnmk00im3nd4pQw6qD8Ifbqow7XqOivKC8
y31pVVXrDJ0ika08Mjhh6hqRs6j7YIKCIyR6VsQVVe1Df3a12fS3CmDEpS25xqhilxlDB6GLGAcF
vaMMYhA9gmviUWtAcHBYWs00FV4dWh91Fx8aNIBUCTvKMBbqZvmoijJFPezqxa65LJGO9Mepa91Z
wEuMhDckAy2luKUaiZQLpaxuCyhaECBDx9Uj/W9z7y5asTWtaAda/71SUh5qody/bNA2nGsaNT9V
uMjhzdJLVPpVlbbTLW6OZqdcZuPweu0uIaBiEXhyTTFUaEkk+58+Ws1qfYGfAo53Pc6jMHJRcyaz
QnnkEF0gs09kpRiCwgI5ipy4Kofd8v4jCknZD3TA6nm3k1NPDpeIZtaikIuDiHpp2KcvD1L/vX2l
fHOfspwIMRXvMXjomMjq+qBYbaAFtTXquj1uq7FoCUQoPF1tP2kIkikKKLSRRK+X21ejLCnINj9H
uspVBRFgwxZ63tA1lZ+3LZxOmNZiXrFYEgfl/nEktf5urB1Mt4+i6ukqPOh81FpMoUjGiuYG6THq
R9GytDA5+OA5RnDeMb7fLl28+DT1SOL5AfKk4SHNkyYkOgUBq08dPRjFh3o9NQYVNn9T39LSmdgy
Ps7C6BmuRp9sZCYQrM1T18bXeg0DI1BVRIOgjd3W1Ws3qbg8RUQFRmYmAnI3upqKSYd2YuJ09kw3
cr6zHTv3JU6WsYq5spalpgfZO3x/eou3L+y15Ir8DyOlJVrHqE48sOoOJnphEtmdRWNoxn0O0fcF
1Fx1pPyDCN2awrSBmcyc68YScrVhtw/11clVyg9cmAQjYKIIULbx7Cb1zz1USA+SSGi//C21soDf
z6p25pS88QYmVAGshEZlcm+ut2G/RMErgYdLruSXPgWOohB92+mPph8T+g85dL5Z1vTdyBKxRCBZ
8Ol7z+vGfj5ukMFNuNN8kzc4xm2E+xt9uQAc5lQAbY3nHZwl606M2zCnfeOx2zKFg4mnJjuCqs6x
2D2ZPXcU2XTPAAyHQbf39n/9+HrU0fH2100PvLobvWcZW1xFdk/SBofQAdvyGxEIfujjKfie72Th
JnQShKPYXTzCDpODpERGJfmnfb5FoRS5xHrMaquI2z7yrBBsSc7gFEz9FrjrdFz/rZ5r/lZNshbY
AHyYm7RGOoL58OZCxBhPtr+dpmGhIhWt8/Enyz0ApobKJqb0tlYW6TpyMhcUFrGg5ymDA92yZNsE
Mjo3d6mWQCYLdDSMT0qNMGO0d5tfk4L/KtCnrnTmDivlxtySug8twa5/m/huFccJyemj04LGZ1Dg
A4HXsWvB6/6EHT6FQf5U9wCgiWXOyCcLo5krrDXDpAdmp/kluVHJwrxVl7dHLIYVqUhca8NSffzD
QmZ7NQjMRIpAGz8imghK6gpDGwIfl5qCQmSIwPgtFakajZxlHj+hqAIh9565YIn2K4ZNq7mjoeFq
KX6M29apYtKqsuQifV706XR2wHZgVbHmrnAtzJVnKH64pRY81a8tpJIiKwZvah5hv1McjmK9h1va
afEdbCUIVJmZ9a6Mmqyc3UUp40FbaqPOh7cVsQxdpceaswGfJt8DuUFy9EEjSFZTFbLT/dUZELOW
H0mgei0W6GV0LEBvggOxvIuNEoQRMD6iqIkTfQO1F1tWg6QPx4aeZUfDCnwKKl1eUMbV/txfTgeA
uJZFXsVg44EBgLq8hblp5bmURrDzUc+csbbcnIuet4y9EaM9bFPe3NX6+aYJ863qBQ2PJvu50FOZ
qRjGhCEd4kRlzaXrcw+5mjZf37t0GLKZjsMyDmd1hAISfHn2wAtoNMwPkPFZTe6+YsSK/59DRDp7
nx+UU/lTxnw+7M3ggmI33Pqlta2JDgQiBeb6xH17JgbCuFa7Z4DQxDLcfPNJr0AXY3DqqosNKpTZ
ULWmx5oBFUYP3OABzPT8POA8Ozh1ge30ZXaeFWKESgKQuorYrh9rqHZwCGQYxv1cx3Pis1dNIxWY
pW9v+06VrodsFFBEWeYRZ1WErfnRRUsO7X/A6Krt/I2qlX/pEuxnSoR8gexuLj4Y8MP+LWMyED4t
98Sic9JNRj9CQ71Oa9I4JaxNbJz15g2mfNHiOucdlhvYi2tIn7C/xtnrdidGOudtSZg4r5MxZNWt
8ykkLAudnCbdXFGBH2togKgfLgqXEqHvm+ROcoIyCc+bfnO81moKgFFhb6nMMwbsU2A/6AbCeHO2
jiW9rBzg6NAaM5RXmgKDM/Dsn8Ij7zxAuoagU5N/lwK1p/CjN/rtXWF7EE7S4eSrZpLCm3Sn8Z9y
vdiJkciMcd+SM6mYw1vXfDDOUFmB8yaAas+Xgry7pDayYCAQ1Jz3GCjw7p5Cl9sF8YD5eJ7C8gN6
oRfp4BWI6wHyGnoXLKNGDiLZEhS9cJXnd6CFNi7VNKPMA6ROhJdCwzaqJUzfNZW11nfucQX6MC08
BfnwVyFvvcSgQyV6voU9j1SialQMc6fF+DhppOnGRqiaxacmLtfNTItoir2tvn+ZQmgLnQ265NZF
GT7WXvV+nA0wg92rHh/TzEc2q043YVmxIZ9TURfMjk4JTcb3aiyMLOQ6MxfPmqa47O+wqStkqd/a
Stl5XOI/Z2KgCbRvpozvLMWcOHnS0X2ZHcNX9PFHcVQUveinsftQ5PfyxVJMUXoob2/2FRJovbEj
OVrY9JCepSq84sME6GSsBmzXo+xCc9oEZGDizoGc59GTmfHOmndgIwg5amxYy6Ogc9T0lzdnNuq6
OHuTOzL7QSbYVCc7kqQJEHvB5CLuHZEHHwovSAgiXNCriWKoWIVsHimMQnNHvyLhjbFuIy8Lse+g
GNgNo+ecFk/RVIKOMl7vO0k1rd0ZfumVx9utDNw+9Kj96YKZNIFYU5855+XzZFS8DRN9Zdxz9NL1
KY4u52Vvy399n/1+bEP0nL8Faxm24LEtFPeGQxMb3/4THNGv/OE2DEBJyB+lpoo+YIou+awvXXWI
Kuf0Q2YJcRBIRK4uRM+RVQrwpDsW0Rge14aTjNY8zeZEDF8whCBjUT46xFO8Swn8uudNnRFUYS8G
1INIu94Xy7smER1cLrOTO/uFxNE1x7L+C6MmjX+KgCiqrq8qtUy+eY3ZxnXNHhXuAOoeTJYaMdeQ
pWHO2oemLp4WjjhfjVs2A9whWSq3UPMMamYGD+YHm8ntM0QbcttXpFhEhqAwIh22HGcb2QzC3pdQ
YtnLiQLezMvOC0FivZrwJqcCpeHoCqEwnfNMlEwyDrfDjVA/FverwDt+lKUq+HCumv9fM32wYMhR
THE5EA5on28rAF5TszYwM241yLFCRcLU+z6rrwiOR+a5zj6TO317E/GTNmS8KLYYrzGAf+3wMUeg
B2Qox0tjNLLf3cx41DD6grgHznLsxEt+E3bI3Yyuu79IuQ+W3PbEgN32DPnodJBqrk3L3FtKtEFq
+SiMCLABFB4wO3FKHeXTl0lbP02agNsE+5TLIMsd60u3mGPFHF3DELhLTKz5qzWgIvFDCdA+TzDY
FCFYzQqTZNQgjsBh+iDSCXzsH2f9/M35gYgI4Q2Gq5PEfMu0N1U5qIkZLU7bpIFwWWboku7hPOm6
zmRzsGQx4icrMvGv9y/IFB158y6Mvx06g647xOuI18CPIJBR+/pBYK9ZJjIB/9YF+yZ+GAdH0s6N
c0CAM/TpGY12+UFj2fDg/PCS2AdVPA9tNyk97jViB3uw/SyrP6QChYewRB7tyViFld7Un5p2tlUG
+AY87tl5PxsL6QENL25DVorCxYU1hF3bxGj5VG75It6RqbN1nN6p4+2NniQJiZPLpaatMXVP2EwM
fi5Q0JwnoUi5XKwQv3S2+Yg3ep4I7B8fYsmS2tIcR5du1jBmKIJrw0rkJ8+QtLt3ZzHIrZ7Y67zF
m7JehTx8sYZa5NfjOeXCoHDJsDX5/DnGSavUV1fNHCohxqVb4223as1AZbRqgNabnDYju80kk77Y
eK4VB2CdN7Cdbhv4QryV4XcY6exylFC/iQAdUt086yZc5LDN5TjDIxWiLq6/Iu5XK0AiqbKRn0bR
8qPR7t/+Db+3QVrVhlub0RajeObt7GhHaQJSVFtnJYc5jH2lWWmnmMV6lxF2+W2W8wMPkF5VSbCZ
Gzcj78j9hJ1QCTteqCyH+CA9BCto691IUMFx3dz2keLMJy84rCRzLzSHnfGDMqDtNEjV/LhsN8SE
sz23a3M3tch1MsCz/BudYxrWQ9Q+U3hGkd3kitCvaMEeXo66C69Vi1i/D4fPi0cjI4sdrQOLflbG
+2kVRK1msiiOh5nye8EgN/BT5hKxQD7sknWjhHRYGP0vDyyhlNp6ncWugMRn/KhgyZODyFHBWQJx
RoiXlNtiavKemwx7S972Zo7wjlq4vF7xeoZqRaIjBXn7ThxYXqg/6PN+L2vjqOXEW0tjy3kjZWd5
JRJ7h5ldSkC983/cd8WExlvRSdjuTMPvSZlrsKNP3uEHIJ6FLveO5klP4e2Cv+uMlgZg3urGZ4De
xQhz07hFnavw+YpESvwojQxUBI6jEAvCNhks3b0JL5lukxPLg/bLEtSMMAsyULCUkNa7Gc73xXHQ
VauP9Ci3NKUNW1yPOmlUhH9FaaBXGaxnn9nJ+Ff1NUsIL8cPi+J12T7Nk2H0Ozo9bapYw7lOzayN
TFpDeQinhwm0ICMrh6KQTapvHOHPIzSVND7KPw6zS9VJE0+6e0b4Go/b6OvAze2hlAp97e/+fuo6
pxOklSAXHBp3bnWsMgXhxZiV7T+/l+JIvzeJJW5AN9J49DujLhdtclzJO0vL8Ugg1seg86Wy0Due
02kJ2fN/L822CqNIvTzCIl8SgNSP+c9iUFXqIZ1mzAgTImFDbkK/JxZKvbkac5yfIlBwjfCizuPC
/KdnK2Pbtfq8ENxATJPijbY7I3j2ktikfUnzozn3o9TYX6ia41KbYrzSvsoxparOGi68EMrCiPR0
Io0i2o77jcIm4q4jN7NAzaQj0xYTb5W/RSsDd1G5cndEpR6LsaSDFlB4iAUIvn59XjyRI1fkOYsz
nDDZX7SfBjcBKgnvakKCs3QBgxewcDlJgg1f2SWkHC5xHw85y1lTDpnn2Dm6hprea5a4IRLZM13U
RIQ/SsMfKg88mGNVjbMvLn3wAk6JyE4iGO6TAJuX+ztLALmPpUHRDvjdC92/FkyWiqvWMiA+9/Mu
VIvEeGxNl2c3OyjHzJLVug57RmV573BmctgPQSRBK774SeIC0e7OQIpo3uGxtjvpV4RU2P7QzYXA
7VQP/wa7q3B/ZF6+bEy0PqEgpSoMb1ieyT3za5wxoycuNRSu03jmDqW/DBMm7VX6bEBXJ7jMo16B
OdpBC3ZTuRzdkvnoceiNEHS6wJVJ0RC3PZcuLo83/2O2LRUvVHTecbbkrYzRb9ZZNgCyKNm1K0Ne
Ml1NdyNPha2TNEwGmIF8Q70UBt42nQpK6CpcNLYwK9/25DZX6ttN6PChr4/CVAImPzQz3nkYE2O6
jKNMh9W7uXzCMZLxwe9+FMAxHBLV1SInEB4AoNaqtfSKP3g1u87Jjj3S5lsdtJ4Pe1zJeN4kFofX
B/F56/vnL/qhpOoIGWLv/5q/t9D0XRClN3P3RggHW9FLRqtD6bL0tLqgIQbIhRMumgSjoRjFxINV
Hh19Shuv6E/q8hN5qio+y9iYo/Uct2hZQ6ixfuzoX6GL4f7U0tM6/0OdWPam8FL5is8AHhdj3xS/
4Io8npSSFWstc9OZyojnAU1X7H5vPL7GrQvwtxc1a7/HF+ALwVsvpvkN1+Jlhdnm+ljmwjtWyctt
M60wDwId2OCRX1b2K8b4ePyz/58KynF7JvFEGpY9DHwMk5MRmw0AhuHDZY3k6Q/H582CbOpowg3P
p3P49qN02W/BW0zMCBITk7M6IGcNd5c4IHWZsyR9hlXy90pdHFG27rBozmlSrPmt5raKO0CD3PXc
Vx9lcvZcrSU1leKf/KW87N0hbaM2Ba3vTaQUnHKlyAhD6wiwXdosckb2uej9Uj8vwdsS7YDObtSE
o/OViH9T/1BSgv1lMUjQ4IyxehqE+tCaK6LglNdM4WWpoAjbuGgVkHyComXTPq1kYNGmPAarUiwY
qmZNFGxVSf+w62NKJNizVrPPMfxLqXMOugCkLq4fGWQjan4/101ETlz4pGGgv120xH13ahj45FRm
GshZ00RXlnuAKUqpl57KZRqgteXPDEc0KUpq1ksZzunnAuVlRgEOw7CDaiYEOkRZgQOAf4YBLdcf
QKeXkMIjK02noV1h2C1xgmpofs28lF2aUkLvgmAi0wRuDe/qcsAJpbOMIRhPTeMtvMvcl05i+S6+
QYLnIQczX32EadD7eso947H/hcgut8OjOKCbl87/VTG8BdA1yYFLQ3gcIsIqSwmBpcCAKdYYlrZh
mvVqufHETeM7HR1E0WYK4vSPsWGqRa3ptnUGrFEaAReTdxDdfAqzjmGBiYfRDS0Nz4rQYFI5hwwZ
IimZcu/+b42sXy4GPlJnQQI+id7PHSptCsHZ3dB3/2eWKhZ4f7tp1qrgu4t4Qoo7nB4KVIIBu5G+
/1M4cKfeVkBZitGUI/v16qi2CqfAc7TMF7iItlLRTxgPrSzC+aigMwVE7mbmxo/M4WsXqIY7tiyr
iOCVr32+OV+grWobtfMkuzqydbepz53NMkl33KHSydY1i3arsXjiq+oEHiju3Dv1RytSKjm/be6S
uh2V3/GPCBBKdso2W3ih2JnvvmRjB7q7JUR8uL/sCQ2M/k14lnxx6xaUYLSOx16HJQOrRNQPCnVx
BgsE7Ero0dTU4Rj/e9e4W2EE3WQE0J7DhQB9xpdAqtwlIHuxjZ4FqRPrgC4VPsAuw8SlI6vFlBW7
56VZ7ogFnIsZzOFw3BlpHnCBILJVFgHHrTrkgmwiWEn+JJHDmWjr2AB3zT8KcDobQ4fUa1sipoj3
TZgma9xXtN6woeh0crTQO03nSCoRxn0WT7g+rRfCxPEtjJv5F+4mmG4+tiZFG+nQq1Qae61g9rSZ
e/XT3bLOJxcKS5jnorweeT1uBEbFi+P2DFOdf3MTJz3w9G6/se9jf1dUvnCn2QlPJRDkQ92GsR76
KeqWHEtC6eQo+K5w36eWjM5Z1Uk8pDVbavLfk5xKQ7DpuCUvoJ9DDcB6f1g7NcfgnDEvWyebp5R2
cRtq+y2UAx6O3rjPlguHkykRSVY59KYLMmgBvAKo9swXYuKakOIgq/1VjKP4tcEMY0A9yOjXPI9u
0yINgGilcK2S5jndZYiuBg5WAWqcAfBBzFBXfoSESs8QN1HeqO2jpRgLWT+NMq4mKi7WUynuVIRA
rd8ABqmAn17Ny3Ne0odfij4mTvquDujYmxuZ8IGPShBmqmmIrxZuwBStSn23YzIuAXh590sk8MWO
1KJYlfes9m6kfydDySdRMC5K2LuATgGm4CKrceLIxo/ouXIc3NqsETpfgDp81hqNhKx6lRIgGuon
Ai1yi01XDttpJEIIkzbQbcSrBie+AYjrB6q/GNcFVx+zPfDK+M9XEyyuhvsW9okR9qZg9To36dO+
kBR36zuNO6Yekrt7yBRuzWcv7Uym3KDQumxFmFdxqhU+agulN1JA7foaHZixWWVqpK1F87D+PlA1
8qaypyFGbDjVQsGzRoVHX20kwKyw7FkBkvDZaF8X5thm/fI/4FRzDFUIhxOpEqIUMZze6Eq5cDjv
/GtkO228k9nU3ET6WOvBoWnWEIvruwSVOcjxpkJb5CjaEsqdcCtO42548jfUGkg9GR/ep21BtBDN
waeINTvZ8sBJL7Nf4GhJoPCKkVdWSNWixuR3cmIXZVUMGl01/e5zuP5STx0x7HRbGqNzy8Hlresj
XmtaSZguM6q/zD6Efdfje8GORCLzUzc8sD+CK7vNFol6L5omxT88nWBISrD+Sm4fQAh/fX5cFndr
herfdZ+F4D22U6mXN5tbGaM7jG9zmhiO12FT4cXO5QthwK6CfxO3/PvhpA7eiZko686hb44n3aPm
K3VSe8ag5ARmeVUhy8c3PO7hNDamMG/yjbFEOY09zOnM0GX4yPeoiv4n2ifSqFvcnkLN9ivV5pOs
EbkY2aef+c1w743fS+Y2BuQBDBDzIvTnct++llwKgf8pP8h0XbhjBXOB2jbwa59fnnYwJsbM/nd5
vqBrUYqzXsYOUMjfYWKB2iYhYwhKru42R+0V124MsDVpEzZMI6s+T2WsCpE6HJLM4ccZ13m2Bp28
2FSnX6bpOdIT36TbkvlmfgPIEN5xTuur6ncS8NYmxQ/rzAtYArNNnGVmmXtJ4waac40dnj3+gOLA
Mh5J7Jr2no1vAxBB7QpHyUWEB+ueZaL1xY3R33t59BXXN//tMvkeRaGh4fBf2nHUl/oaa1qoB7KB
0ocJ5xEa6mTVT1m+TA8r9hRAgTg1hlj27SBXCDczgM54gSJ/Jc7T4hibLu6Ilixe91N/BF51qLhZ
eVizhBffyD1RKJkIvs6pmqUZo4YZc6HOIGv4A0QjmlmYL7SbR4vbW5JAm/0Fne9HHmVpYYdgh43u
VCnNf6av1fVD7nskc6wBLfyB4koMgBvrkej0kI/e2zDAyQe7gymisP3l5YUFQGoiptt90fGfLOsa
5grUB6M1pkeXxoy34TleYfjjxzjnFD01zmhKHFtaVluv8+TdxYT1PuyXBGtt6Rd/g29zL9WU9FQO
Fl7JxzVL1MLUZKVbY2RAipmeknN8Ri+QD8Uzdj0zpTDwmi+xEXj6crsXETLLZogNGzYWyllvuwty
T/P6PZWFno7Fu6VsE1G64a8QftTVyE0Rjo0KPSMWOWUSrFJ7Jd3RXSVe4ckd9CVymAvofEJ/l4IF
c060lQbDfn6Z5gbt5wihso7BSAWqZ93lRCZEezmeuZcPrLFXp0dCVWN8rtKGkbsQOC3SJybqlZxl
BoaKJYq66ySCKp9iifFaJ9+Cd09K7uWxvD2Qya47FUGaARZmMO4OyzYR/9brFMjbnZMM/f7beif8
+Iv0q7PBzW/m++q+enHkcC5Jets4Aysk1dr4hWSm3YSrOpIUCUNKOiY+W2URmbz6rh3njsC+ufYl
hJCQUbhnPcai8wL8EeRXyLaclcpKBW03viK/ThlNV3KOtvGavekDTBaErVkoQ8/8UZKds1RlpdgW
Ik9ElaT9iLmhbPmX3DVXGuMG/Wbw75YhFObgSzPvhH7RZGopUt07JxUKTObyuJHccMAxmcvoz48N
n/kBe+idjEdhrkXL7+KVb6BGQmsmLl+lkOxVjVdMZX1TrYdCDE4kvHCbWPxltKzkahLsEH6RBHQ+
Fs5oxB9ko5YPtYWeQLMBwE+MilN8Pe66yWzZgVvIMW72uFnNkwfnJCGKEH5QgQniduTw6B5ewlH1
w/eU2glVNVczX1nqpsDhGtk3LHgjwIA0U/wL8Xw3vyFp5qALP2eMLE3P4pEYgJAmZbOrI8VNQ+D3
yh8pCZ48OjFGwTUtY0zYJ2ph+nLrR1oZFLyy8hDYuTV1wZPF6JoyMMCtMe54Po+S/UVt2DhyRZJt
6NJbaLkRthRJSQqI0mtVGt/pEWCDltrQ9MTBi0xaFwMo/BvSSN5MB/0HIAM+16B/CzC5dDgAqo+H
O6DSAoJ3MxplZMJJ7nPZRl+i4XMuH0GIuLitfnZN7Z/K3MwsB+LHnaId0Pz0Q+TS00dIapaGWvre
awKdP1LEmtrNpqdLliFQ3UXW+SeFHr49R4KdRIP6Bx3sMHNCt69VhA2mxg3GCN05VgkfLJVwMOO5
nO6ILx5aRuXbL51SRC2Ex+sH0Se8f0bd6ZCvCrfc8UTdDxy7nV5vL+xEQvax2zF+M/bAodyi6MDA
fHtvsVHrTN+YpreKBHpXOgkWb/gXtoE5dkgaOhQPtponCyTPq4mV2k/wfdF7uOpqlRuKdo2q62ee
RPZanQqCdKKSC/9LdpYZvupcPdS5kn8uXQYrr+fHxNBhX5PodFcSAMzfZu8+eqrxkTRmlv4dqkXR
kkqcm5CbaJkw8Zrshk+zRtcEMWqdflUc5JsBgfNBLAdSth8rLkpL4hlj0DCoFu0MUEZRQg67NcGk
S+h2Tybk2dUUB+rnP/hvSfh+CORqMV7R90paPZadNnJabC7Nh/Oib0BuakLHr4wRJuDnL1iOT1BN
QsCzV131PU3jaaGLnqmwHPZ61Pps2yUjO1hRrxUdcgoUmJa9QhboQI0u1tY8dqp2rD1VheTVf+Tx
wyiffp40Q803Yst/21j4r+PKUWZrtKyzbFtnVpthGKkam4Yyw/UIfTu+xh+frEnFGoNoVRyO2hGd
hWQIai+9vFIZLifL07ObmDxtigIr6rF7rXjOYJSa7njrRDPCJF+Vi7mbLiR0qSHxUPAsTu6Vk90l
RaLeV36S1XFcUENo0ma3luJbufj+HHKqzjWbM6ks/nOlam0K0d0ZWFnAm2R9Llp+JQF1MDimTZvF
mVFMMzkDJqsL/4aHQiffyqyF2eFp3Ih2Qwns4pBM4xBmUCWyOGT8G4/EY67ahqrSYjlVb3MCY4D/
9uz5uj6dWnA6S6NbHnf9TVUlB/Y2QqaHx5LO9k8VHHRGqJULHrzeC76+fvwN+QA3aboIs/15b6TQ
+KBedwBHbfpZiNqkvcPw+QWDR0cXgOIK8Ah8/SZWfwv7wZRw9MSoWuou2ZrfFMgsu5D2Pmlk428B
bybNddtgIEf8E+4AR6WbWULd2oOaYkmbo0lXhODF9986ZjUa21eVf7xhkhvBLIm0Xph/Y4QO9W18
cKHrCN9zusXejabIbDrQwagDI+aE+wZfaApaiWJQGhTytsmJt7MucQi0SCt+FVlgZJ13L7IIVrEa
g2BEn4ymEIU3/acqtWIj54YaxmsH+ZdjbhNVzFDhN78GGoX8n61klA4dW7iD7wiqN2NceRVTcYwp
w33FUZv1CRBJFxUZDkBv6Vb0iN+Ikut38JYaWIk1liflccX9KaxTy9tKlF6kfP/MARI/lWg9AuEU
sg+iAyBbmiSvTOAx12Gj9OMu3XK3t+ZzyDKjWTSwilFXbi9nWKyHZShVzoPLiBfrm/GAIp8cKtkI
IrZ4blt4h11h0xzG0RnLCe2k+Szi4bPK6UQEN2uGmGK57Xp1Ho+o0k3BAxWoT0n2LRZwCcHdplcT
r3si5YbQ1rOkRIOGpis/R+llXFD/mS2mukylHDTUjLKv51lmCMpR8/EYCm/hKdNkVkYt16KlePMf
gWrHpPi9xWBucyNTd4UDvwC4uCvGAxiCUtKNsBc/0l8nyndlg4y+kNegROFNtriUDWfsSS66VOPb
z/f6GFcwYV5UqwJbpYBUK44GqGxLCadiHUfbgo6Yv/iVyEUPXvKr5AWpAyXP7EXhK73Tw6U98tO6
BhBumWazjHbCv+MqK8bTawj/3SICXoOy6POzSPOiZKz/gXy4jZzxDluCBOMbcQ3NhBisIpxPwk0H
svdlU0c5+A8h/WaqG3YoaIe1mPqeXZm5VhagsKIPjOkrhOFrcWIrRPPckC0cNymumT8vzxxY0BuY
kQZGuBQUmTuA8WEE7W2JIcYFJRbVRLsxKgIpCZbmhEUx68rTgWu9MTvHQVT418G5ngldlYG8BQjT
aaTecckZhcSbIoO9TbdSp5++hYoh9S/C6VQpWqtzYL81Ta1EPnntZpcM5iuSXkkLd3kaLerHLHFd
0qvat8d9y8ioaKDbdo0wTlzOEIE5mHJovFR2T1t6iB0qtyIMHsqjpgMsRkB9yoy9TC8zfEbg4wmd
s2t7q46DU8lApUpKe/1nnWQoCTV85Oje70YJdabzAa7DNsvh8rwT/SjavcsM+8heQwJQuPHcm/mB
NvAeX6gauLF0dDrV/pn5kEi4wJqmzj0K5VJX0Ds469mPn7qAd9NVF72AxJmgOCWhMIMlNbBkACV9
dGkJWucUXN0evT7UjBP90yhYQMKIsmOMjse1cp7h9GROnQuuhK4QZLfgi+/Cu+MAKul/LSFBjFxv
hdB0DXRC4ZzdO+q+5nHRb0/6PfDWeKaRTtl5XY9xSUTGWVKkdGpDXX+XvmMCIjqQbW6G9ZyxuBC2
bNqIARkBY5e7qcuDJ1/d3UqPgjBS6eT9M4rMqBUggCUEC7LZ1FaohGZxxO472YoP6YrpGiTg23Va
mWUkmNgrH/BhnSQiJUv8yZTIbtfWduAij0r1ZsZXWvf3X+LBciY/Kl+hXHflo4I+hpCF3KtGySkg
VHLCN5oMkoTaYNpVTigJsd84xox8p9JGXtp6S+ZbP01BDU784Wg+DJ7au1eGGyz7vQaFefsry+JL
y54IyNnseAcJ+fMKVYKKk/4uqMW4ub+oCtwPiUxKcMfTIOBn9N5FD+s6tiSS0pLPwpuP6zUU6ZIn
pP203TbNJBSqlbnfVrn686QoEXF0k14tDwlbT/CkpHFwSKmU4PUcYzXaSFxCYt5BAO5XjHzrzw56
n55DTCW8axXqsjr5PL3ffrb9JG5Cdfc/B3NZfqZ2efxUJb5mDrIczzzeu1AUfN2FfVHrx0jwDh3u
XEV7lVCbovDxnFjSXTn+rXi8gwVXz1GAAd7E6NOLqbwD3hw2Matl4E2rzy++qytLV5japzz7oD5u
lHlXeZ7S+h0Zp3fzZabJ86UlxQL9YZW9QA1t308X1QpgOctXktiFuryDl+dcDv+ECd0u+U7uedoV
wNKPDMu00qtkfI0p+JgIGZ85HxuZSmNTNoPrj40V480ia8sOh0R18dfPwIGvnNVwpQZgC1qq91xk
LXb+6bVhSGVEC9fYmQe/QfFkXhMmrxH2Y3ouVfyiGl5SA0PsNfUx1Lp52T18Jy8gCtj0LaBDUNpr
U8A312TKRTbyZr0xanrFivvNk1A5tnjVKY0wE53wm42mbQrf06yAV0fwkDj9t/Ekx7MxW7t9bFwD
alDji/HE+i1IIV5Ixp3Xj+g4I/CEQP/kibR1jHOzxkQHyZUNQdYrKqNX37yndyDX4Jj8rkOEP9yz
kRX53KwW3dVz9OAqAOsquoOymBlSZIZvvMc5EhVcr4WeY5ncwnDAKnwxcYRJJl+slzBPf82CUQYA
wdNUESPHVnGxj169M9e9HNx8SnQfm3Mk8ueezTRYq5MZColv+ILuJiK55zYHc0wZLz7bx1VFnXs7
sSfVNKWUs1UHBvIWKGGTurJiElGC281W83AJAlfzCgs0gqzkTc540Qyer+HvgzoT8C41Ednti69g
OF0jEzlW2Fex+PtiJiVv8ANDKPYmVQL/ILZy3sDZpQwGUpQLrUj6EQAhcFroH76L1XxVeY84JmNw
hRFwqMdb0QJ5KAO/fYiVX6+DH5GOkN+k8yQm0wjlmQyWHXSv7mv/EhzgUrB5X8Ss90AO+BcRFXac
0nJ+sWeLGqGQNsw6YgL9l2obs3zbbfdYqd65qgHqJhKHw3Lqvl+uS07xP82aXwiAFvnxE1VudZYs
/REQowVttOc1orwPEZ9GiuHOW1Wcq1X8ersSCnQu2kg9ZiTtUG5/BPxI7wC4cxLO2cNSIo2eLzd+
SAA8kOYCPVXzNtuXT1t2bF9CNgsiO9hu1c3BhSv9itWaBbQPW6cNcdy60AT637TInBkhsty7tDaJ
K5PuMJmrLwjo5xvlLnbE7jPNVip4FZeafbgnEDer/f7VtbdXDc7yQ8sK4xfC0z9IbsHrgDFc/uEd
FVXK/OWhy/Tx93ShsVBn+o9JllAFO4uchN9s3+6LG1YEsDARUU9TKVDD/PUkvYQBTkB3/i9/w2OJ
e8qhRcS2WUS810ZrFyAtrGrFShcCUG/iJsIw81ZUCmbSUJ+JQGLO4Ti0zuyhoCvq1j/tG5R6LiIZ
oqiNgvVYMTw1ZRdSJoc58YKZUp/sPw7T5VHEeKm165T8PfC7JWaP0Rz36KiKnkMgMwY/TdW/s90I
RC/HpOv9MicM7sVW+f4qvp5uG95ams11IMfnJN+hSvtFYf/UuTBdNVu7eHgSwFjRgFOv84pXI7MC
VbwfQ85+aUUnXarW6l38Vk4KiKn/0qanKTS3UgaBagNfl6PQjW55uDjJavOXDGtd7TM64qyFGYwh
Yr3xPkmRKB3VYdUCM1suzYHN6OyzQW3Db0Du0OBfUVTUUrhgmvzd30AjDwRTQakyKzDxtzWwNVjL
5VvyFwjxqO/QJGqNPJ9y6TZxhfIgIb2WXxff7DyPIMraNxzqWVIzPZFizDg9qBd6WkgDYVRmqGic
pYWhpLJdloFyi6SEnWpWC7fh3Br9Txg33tF+p00R2nSdjP6BTtx36xqEc73bKNKUBhvHd+2HE2WK
ehf/Yy2Xd+E2LK9IzHmNPrbuR4Ya1GveudhkBsIJuP3ALZHgPMhUWpEKGe58W5Hwb9gsGM5el4FS
JjXLgH4+P0qZFvLKp7/tLU5NHq1ilSUdPgYRKHuSB0GdOwYJJx2jcvkckwZxw2AgiRJKc+9BPPOV
rusb2oeMJ5q/P7WIKcTxnTgNMQM9KTNqaSJWvdrKJv5p1aW4G8sdAGRIMFtemDFQeIKR/l7CAiZU
qFWhuTQNjA3ITyY+8AnC8foaiwxa2cNRKH1cU7lLkkFOjHPi1nVaDksoq1j67P8rc8zUN51NMFAB
ib7iSADvdFnG/PyQuD6mGs8v///reZrgE0uL5pXML7TptYLgZjgvF9HxbAKHoHYugxsHPxuUGovK
ZQfxliwMgscK8rSfUlkhgk+/GlqjnbM+zRCxBDiBRa8xqCox3c3RvHhZeQq6IwAZBw3PoTWMrvk6
W8qTHubMSp5c3CKWukEXtRC7X3gVXt+XNr4Y9aNuq98EH5nO40LtlrOdKPvGGpFKsnk51V3rwBmT
pwYjHNT9c84LNMCkgw7+wnDPlI+o+Vv8aZrBj303gYEPpX304b7deXL3fWd0jPo6rT/AHgCs/Mz5
SFWszsiIB01kt1v13A6bq6CZviE9OPmf52p5+21Y8hb2oTHsHGN+lOvsc/V14/QCtLI4W9Exei3F
DV9vgFEfHnSmaPNXyxnunmW87BmFA5iE/PNdylEKg4rMwXUOyO6bFXUxA15p/llz6qWJOK3JFEq1
YVqr4y6B80yMJ4ImeVRVxThEkiZAVcc4SKbt5NLR8zJIkMzy2684UEVbz1ACLjK/ip1Xf/N8mImw
j8Xe0HWZ7hk3E0L1fyyXZfO2r981aixvtfdZtxKjber6naxttP8QHpw7ATNrRqIOlf8Pbjr4AShi
6ZDHhDY1OdMDjN5DBtjUMD6tB1R35UD+1dk/6SOIbrtxJOyn4E7yJof1d+z8yyK+5/pB8M05cq8H
RgR25t0MOpkeYlT1WLNrOswIeDtIX0yTI5UhXEgyy3ohebiAatCuU+4hEg6B+mRGR/eANZyJNKyC
8pq4dYivb27H9uOWJAmc8yp86Wg/9UXNu6FiuhdLgsyyz8fUHWniEPjXJK3nYATk4opO9dtrTnz4
uhNlDC/DO5voC2lEu9sPWzc6H4lrZgZHVL5xTAbCT2V8cXe/nQrd0n5D3jMbCwo+VlIeaO6rNIMe
J4X6BFx9h5N4fvg0502WNjTjcX9faJRAMJ3VsmlPx0TbaQhnF9EL1dT3Tv0GNqffqTUaes1s9XSs
CiW2BEyz4T3suC06gaxDuw4bybDqgczB+g2SuuFBfb8d8bzULypGDMM4aGPlrLBwFW0Ah5HEECpA
tU4oqSxaqUFK2LtfnfXhLEVjInhU9xfvJ+wpn2B5IcF82MZJ49jxqwDkP8J2ukHBuhQNjIhavoAy
oY3zA6bykefPI1KBcmo9NGk2VSfG4h/M4D8erlo/JzN6GQFQiNVOr2z8+ob9li0nNcMh5RtU9EuJ
/f83B6bt4ytDjydKoZbLlX0t/JJNARJNPvO121I5V1wKChrAJPr8idNM2y091cPAuA4Bg6imZdFL
4ePiX3HABHMAm0Q6t0HLax0r36QNJkemZMldFKy6ZHlSupStLPNt3Tnm7Y4QMpjUxZE4dp3bsfWt
su/h/BTF8QtlUXjtQMMrGFmTQXAlkbJtLNOEpXPIjgWTJbg1BppyvFrfOy13GHAp/Yh1I+OdiLil
wET39ekIfhd+363qzH2iqGMSyOe3Bm096OBSN5S9XRiAaE/AKzztrxTpiHBRucMLh+LiIy77q6F9
kNwmmEoZ5U9z2DGsFTKzWIt2jMsUlswvizVGyRY+5+xgit0VBozZAW2nFv3JfU1WrvHhoQVbrDDo
whMY/HHg8kVOE3tWjM+PQXrn1KSfOGv17v6q3l074BQkMqORTUMTVtmoqydRScMrZW/Jvfm2LTta
jFtnqUie0viiF9edK6gmD/pj4RCkhIqkcdFoNyBFhg1eZRiuzSYx2d3C16Ir1dOjBwh2SrPdk3np
hebcRXoH/swbmApe79adfmJ9KGus1ps0ircj6uVjYMKnyVMZdCLQ3chFoqGDfViroUfM3a6D3SJX
xUO8FlyBB+M0R0b7iXHNaNSoc93vYV+7yNU5d/VXDWD6h0RXMzOOFfxoYeawmG6df9rK+tfbw7LF
apVV0CgfuKtn5g8O8xbI12nYyD9TySOW2FutoMHcMaXxl8NRBUSA2DlmVhHYrnJOo6Px4m0wQLDb
JOqE/rQORm0xK21me3HzC0k5LFhse9bUlWmKAfJHKMVNc4Ef+yHrV5mURalhaAxZjpjOgsNiveTQ
s0PacUy5l/+Mc6pHp7Ry+hMBzt5auQf5w/Wn86MXdFQbRvNn9iJQMdJ7WGfleM6b8Opm7H5GD9hg
smqhLzWVVLyXAFVokrLh6bHhyOkT9+40zumyneOtbks2EZ/G9OvEGnyySSJ+s4UXNxmdiZWx5fAv
DB0PQHKCNBRG6HnRA6GXWW8pCS0NMaa/ZfVsTiVZXd6tqD/KZPEFFRc2ZPuLNHJ4lpkiBTZxNfmX
/saWzjB37pnrmVvlpskCEW+gHQfNOmZW4p63K8lhdyw5/8FmVfZtOM+eUeiZQswWKpLkj3ws4iS5
EPc9+R/dxV63XLmGkHcF9J2Hm7SbEYbD8UQPhZ4rzPcfNLWdchc7n/KgiZtL2iptzNgZor2GweDI
9WU9Ps29se5Q8cBJc4BjwkZMrxKccuvYvHqy/jzvVOBxSYpMpGCbf6mv3SsKzyxWL31bg9n1wHHa
IXx0mGoYKXCUeH14YBkFsojPw5sl15A8iR1VmIKl8ZwZw5i6tIkXsJI1stsW2ezgpG0Z1D+iDyNl
GBPKwwSEinzUikOIXs9VGIm2oM8u+HPqGZJcKyq4XZSOm4qTuKJy7R6aMGmWlRwf8E2JUB0QzKQB
2b4o/ntQo9iDQVG32gc4QfHRanxj9wpGq3RgB31x1AcuW2dsjO6OBz7oWXK6zj1Y3fOv7YQ1+aD4
pQemA2OOqKTLLwasbo0Wrn1NE+S8ExM8a4iRMwXGfWPQj2bqqfSC5V2gHY8Q57cvm2wmLANXKYJx
ElKzP+7RHNR9DJjSQktzOYMKPlpTBqbHd7Oyfk60hii1Puu5028TXer+WTcvhMzwiMtOxAFuAUg4
5bPm2aBgft0OudeMgxhY7ePfKPYr98iJpV0/3nzURlYcuz2F41KClHyQPHS+Z0MOd3Gmy0Yf9jX9
MRC4e+1vrgj25LSvgIdLuqaHbqitfiTcQfnSdaJuJhXNCeQcvwURoKHuhmi9sHyTr5fpx71siomR
qT8ghTlMJWSY7PP42b5J8gZJQWSmawssTsPuQpurPwI/Kiw7bU3z65uiFXnCfSonpsS+8/2jXof0
fRdlNx2reubTYRvwGXS5xxBJhYE7epf+M7ZfCin0pTD1lO71p2+AZ4/75cb0xriBohK6veQmYiNC
zYJ/nIWxGotqAiNa54C+UZr6aEYS9uD8xs3M7JaR2Hu4PaLTIa2WXo/bGMB04MjppGtPVss1WvPC
eFuN73sR9wlGK8QBXhtF3XnFdZRV9WnlMPNBD2Zjh5zOlImU2TKdXAatfEk60olTGKL8VVoYFsUq
9R/Gt+zkSD+Q5Niip9f7s3MAkrCpD/C38rmYEGK2hZb1OD+F6F1Ud0bl71TNKqFQiCgZNFQbWQsz
2GvRIzgI95/4OQIE37S2Bjr4n4Xu7wqTJIygvQfLfkDTSgGb2YBjSOc1Qro8ga7hpcYG2JFOe0I8
Qh9dWXbumq+tuXoDQpDYWd+HMyaVpl+hshPt43FmBIXvtLSBz0iU2L6XuhnUb+o4SIjKznK0Zlzf
2L18HqPeIYOsQXn4ttHEXu2ISFzH6b7FKSRryEfjCGgqOD12JziAAJnZGoUIzCGPVVAFwrblC97y
sX5FkQeLO8AhCqfJIvrTubEC9QnOiTJKYET7h0rpPzeoRANFuIbpb7p013VNAN/U/2XwGifva0Px
Sw6GnktBtsYi8biu9lUBtuxP1/ninXibhls4VlL4UqNfggsKAfqTzRnGlBn50ZyBU3QCinLCzJ1B
L9NFR4Z1TG40vf54dxCXOtVBo+KJtrI7PFp9MXa7m+UQfxj4GhH6zm0i2BsCkjQMFqNG7LvQn/k1
5nQwMiBmb3aQKT8OsKxoYuA+DIVCU+vG8kq+zPjA4MaOOO2o9c9hma2URlbV7taw4sIHEhUNd0iR
d5kNO/r40JMCqflZVqz8AtHpddKZTfArmLR9k2S06DYeL+9s6cw61y2AbXY7q+si20Q37gDk/byi
GVKnWqZWAO5rufoLpn2R78uQj7APvA4NJpPqK7lrNZySNJGho3Vl3AE70Ub0ZpfJ8+LPEwD9MIYe
wuX92DestlENhrSih4GhU0RhlH/uHBlxP9S0zkwZQQ/OT9G/JRq+jEKSKUC3fKpkKua+F5nUDfS4
r72UUvPk5pxKzTi5Ho4AW82ixaajdOv2RGk2f8ZTlIMcBbb/vLZfaZMFLC+BMIrYgddl4FEb1nv9
ZsdleZVXNJ5+h+0kqCvXydXlVY+tmBDOwZ6AaWhUeX9FdHC5eF9bkqeBCaCOGTYMm2G7Bb1JHMIS
bgofxZX0woyzDmd1I0hB+JWrGhYf04eJTXbuwk8o+lEkvQlOBPZn5T3NaDAjRSGCmDDg1q/hqS8D
sh4pCyWzlzRZW3loVZk0vudaaZXedOFzav+VLcd9ewrRbWaHUeBea0wPcfz7u1qjafjgNDc22N9w
1Em6MBkoSUqwQkk+aTkcG/GiT3AH5ypuUWJlagxgSWSNalaFePg/FHj/obz9DK2XWAoz1rPYtzKV
12mwl+G3hIqgaFcElcbjVgh3UZCIvLgDEz//Y6ySO5pGsIS95Fopq2wKWjez8G139pHwMEvAFgru
g2jsNFx/WQLzhOfDoRWW0G61dzSUwZ/35kXdHgsd6fxHw5z1PzsX8mj9i5IgX2zmhWHfo96PSU60
l7tvEbLHZ00A2deIzW6O8VzeqQA+/qsAFv2CEhgk/rwGroCNnE3WnuoTSd+5gwlyd6HDqo3Tk0JQ
TP6S5ITJjiU1vuoHnjRtWtZk/nvZnuTdTXgbYSnPs1GxIcv1l+EsKvW2dq5IFJEQ9ercVwMrZOHX
wieGzmzkt+zXUt8muEGu1Pd5Cq5O5vSYbthI++/C7mvdmMuat6xOUbgFVH5cc2Xhy2/gYpf/yTCV
wT9QmP3N6WohKf5lGaF8VR8f/EtV7g+ynlI+o+AWFxe2eL1N5i/5BF0CUKP3WnxEq4CdASVikl1J
AwicG2/8YYNiT8lj938Mu1r1JKfmg8YRh15CbDejY/yxxQTa3mRLDBVuz3xBbhOGIYdzssYDdwLK
w7ydGcUPSCndv72womeatHRdsV3jIHk5m54raE38FsODIWGJndvEvSc1LzHOPhwUnfgIqI3JdtFL
nXjII+unxBlttFqwaC6fie/2sf0t/Av9uNco8lK/vmzSNc7tNhITRf186z+D9NVz0WoECRoFn6i2
WyFLXh7Nx7Khe7nsAkoOmDYejxsnh8PPui2P1pfmN6MFpw1N33qCk6vl3ZRF1SEQOeg4+RxCoS7t
PjvTlyF5P2nYrGrAcbkWyf60n3CHvXfPCINersTvZjXXv3WR9XivxRnMhMkULcTvsX06FdRMMIF9
cGaLKB71ShJlDDI4S3Wux5170vONZ7VlB/64YcTfHA2b5tCWizwczqM3FbKomsGp+7iF3BJqGO8w
/7J+hvQZVTQ/WosbFVCc/ROisrNvwNvTo0G0wqHQ8qybhfU71gyc2Vz+DiMMvfFoXi2iJqUwhUGA
Jbj9Ljou5Dr+w6GLd40gCWzAQlv3G/qNgDr2VBgARZflz2xratoLd9etEPQAuwYuPhlBil/n5if1
pbvckbhTNuhC6vj+uCgE0KsDYWQ4vCrRrXs5nrNImIE0C2Jxbgz7cTL+aqSdcLaHzDvAi4V9k8YO
/3UqlX5RNMhB8oiH3zcyRZS02X4tkHrIplSx++zC0dseBrh/KVwnJQ3VHaYw3mfN3mGLJz/ybk/T
7952USBjtpe8fycBhuPLyhdNkG1WxXceKst0Huh8KFIqZOtJEY60TyBR1Q5UjCTKgT3ssQG0/h1O
lhL1cl/r1ZwJEpv2P/4C0hnhnfHOQ+wWZRDOrsbsqtPYm1WPrNGmWQenfJTxqqScfDepjUig3Nbn
kYxI3+Zg06hhaAgvOBt9FChePsWWwtO5IMRpr8tzkKKVtxfbn0kb1ZmvbfGk/uLqyN8GcYQQY4AY
vq58dqh4uaoyjivrwJNwc/Gf3mRaYQ+PQQYon+e7IZKqgxHTivQX/UdxUXCxo0qrwKGEcfZ/KRVS
wa+mR/j2rtdKo40kCNOrABFe0Om33VOEzklb9LAWu+hEGOURglOmljtumfqCznW0c08gwgmqLx7g
tyQMlDxclKLm65LM0HU73GQL7DopomTRmJxq5Y5aFhj1LsRP4t0FVkQvRwKHcUpo3ylPRjRPXOuy
gdIDZxToeCBrcQWcoqbSkwc8xuPNH2t8eqipD+G7l4Vb0cMozALWHbqWIo2504S+aeNvRFQ1IHOi
BNn3DDs2xUzTAzHqBIomAYhFVA2fMuvkbwumAxgi3mxTWFVSkDP6A1WHXhgpLOjke4BG4tlzBlHn
ddXPiv7JHD14MKS4e76qHctIx+i2p+Dqr7r71+c5LHkeScsHIPXaWg/9GXDLhZL3LnXjjusM3ZtD
tCGzKWnz2Bd1+83+08is1puE/3JYAwnKgMkklIjrP5FnfToBiIVFoGoyzfB3yq4lHpOUhAnktDP8
gLlKw+tGWYxv8EUltbuKIMVAZR993nbKZoyNEVCCooAgFrGgOvtKF3icENgRdCGZ5HQj83ZyAZEU
KQFMO32E4gEa9hXAMufoPFt0z0oUBZkVepdklPgI+20AcX4dapO6PHHjAK7DbdAldfhwUBUXPUO8
xUs391I3diJEcU3cGyyitI4lt+yPQKzohpllcPqtZSy0hEhYE0AiBf4CCZlNU1zcwyIqm5VlVwOD
yJE4x44x75O2rSPfdrak08oLkBgA36Z8qcd7tUr/HahTyXOTwzS19gDX5SfgVwTnT3vBbnSE2xFL
GQK4nHvuMzPqrmw/VciHv9ggrf2B6jVkXWQXT39zw1YrD4VP9neaCM9qp3HhItcwzlVq9PU1+cbG
YEahw5AQSx3PncCkk6f2I7fTjHau/pkCWuU4fgBvAUeWbjMMcCF0NJoOy9mDr2EVS/LH+u7/Weut
2xamQsQy9oRbzivBwKXHYbPiYR1JBGei48NevDOy/BANHhwJDfIrwXuvPyo3Vovkq+u6yaiod3KO
optX0XdV8h+xgAvnVMTi85jX7o3rSQ/+T2O/rGyMVaEIjeJYOCHK14b2lbaL0VgPWhRTeQPSD7Qg
P0v7Krf9kLggM/mxRHkiqnfwTzTe9vBtsyEHZfa0ixIy3UXSLv7iPICJZ5eNpme74Re5iRQEkFHN
yo86+GXl85eYWhnDvV5R5TCEsm5alQKXes0/G30FB+khfFIZ5Q3hYG1gVvalSmIuHjCk7OvyvMDD
T7Q4dJTYRxmQwdpuCVCEIT8zj12T/p1CdMlYDobv+GdhTRp2TuswXp6setIsk3lMyHklbps78v1U
PlhpKzPWrOhaMAsknZyn54QIpp8yhZsm4wtQrDE+Db1fgu34nE56gWzmFG4U6eZT/czHv3cInTfO
bh++XQyQV7EaSdbpScQPoIXLX/qG32xMiB13ZcX6mVYjJ/YIwNLC9MyG8IkbsEKQ9WBmhdo6RIBP
96jtRv0L49v0yRHf8sPwZJmTHjUrDO+F702x45SJ+hDjNd3cJFjcIwFhUd8EJtVQ1rt3LyhTgfGc
3KrYgBcrnLcRKM0TjXtGdxvMU5nehGbod8yEj2tjf2nGHuT2pURo/8YKrRBdre6FPQwDyFBskutL
gJR7cK0KBOjqjJpxdsKxnBwLHRKKnBNaMnSC/fejHIh0WV9FnutwR1UEAWeVDr/5z/Mr2Muzg5Ls
ut6w0r5JZf/khYznNnJABkVWOPqDyPeFPljWfi0uGqD+sFm8iAL2Hu2wS6tZT2h0dj+NCLsULE+Y
fJnDFuqokJEIRDKzEd0JxHnzf5rSQ+2Ue9kRA+hWtCp00iIQ8XvA9MIl99/z4jq219x10NfwL5nr
8xKz7l0tq8CIGS57Uuzs6JGORKnFkLFnoIgOrolYtfjwBDQsT6GsZ1tOogKcRtujEsX3ztgIw8J9
jMBCIBvMwmTJEvF+/5yVqjvlYvfL9iQ39sDWCU4gSM1k0t/NGCfKQFYKEpA2EEa7wFH8zKxgAieV
tMIwWJ3b6DApK0zOvMrx4CfzY1YxSIOEaNG/lFTjViFLbC0GT/gFmtolAdrMK0hNh1yshzH0GhWt
3U9tcHYxVzsUDWK9nxwdkXYVHN9ZP3KwH2EEVO4npYW4fotCAkx3Zt0KyCXeuflwp7AmwXGOt7g8
CjzXra1QK4UehxnannHxKv0/yutYvI/4aAjfS3QlE/wvywecSxdZzmXfRHiHUhn1hKKHaIGvDBPV
sn4bKxwpXkfl5XjLcJjKbDGpKnkLzbRjB6YrKS12rrO1XB4fhYJaBUHXJAbNfNsdxWOBisSa8tJk
q84eS7UxNJfwRh/AX5GOGxSNnWSaR8eB0QiSNNJ9IS8MjsTlMzPyWUmsxjx9EITUQ4wArXF4V1aM
8UksaAi8WlRGUzD+9cJ1AAHiXZiBqkrEXncbUJ1S5CbxYGP+vGYA6KpCNL+6QXzdOLzfvZezCaDo
TaZd4Ro4hth7ijVlVSt8/Z4NmENaMz05GksUHHzGzZG3u2vT70VLLqE9t2+N5S1Kyj8wiasr4WUv
9GdFMT3vKI7g7NUGeJiSpaDlbMqGWgJUsEN8TvEHfWf8G0h1wtLSmF4jmABljhbdXkbHdE96scw/
C77Qo8tmAtpJRlRO064doSwR1WoT8Fu+xhHKMzpJT1Lhh76mN8H/RooSS56tTnfAU6xtAQR0PoH4
gM1+lR3v2LuWL9sU3plG/q7Xz5o/fNB/jy1scn+3p4v/UwKPyECK9QOWfmSBXJhPlJUsongkX15j
ShtxvDRqOhyPtBgxkrn+e2jx3TjntIrPayhszEN+eL/R7OULsLHwVWfsY4tapbV8iMizdZN1Ahz+
bRRtLjuabsuTWwIP7gOMo/+mvpsaQSz1Q7TnggkIhZ6+GCtNP3EoQA08qJNa62Uv7qJc/SxI0z/U
R0ISuc91CLl8QVrcDjzqnyYEl4q3SYTikxevvbxtv8NMme+G0gP3ZobPzFVR7dwLBSAeJRFcuMD8
oSC1U2lHB2IXxiz5xYOtH29JTOuCJrGPEQ+f7nGb7UAn9B18VqllyCWF79P69Zm1/nZicfvZYvv1
umxJWRre4j54feNRGBWN3Fnn8JAgwUweeo/z+Rb+bivNR4IKyn3AfQoNtRw/kW5+q79R1E4lvxgd
4TgeIS2b3xG61uFLchqb12/xULl5xYd9/Nr8gcl6kpzqSAX1ykBmEFTWd+YLzvw6xtOj5aev5NEI
gPTKDAWEefPKZq7n7BJCFDaRdbgfonqkpQsI1KjZkIi9K8X9APa7LOMy7/OQDAuOiI+Ijee8kCvo
T6/k5hbv+LGUK0CmV3x7BQEI9hbOmVi0tqxC8BO8V+nA9M6AvPW2xv+wMYRPIY7/PLNQ8wO/Rnly
seDpx/SVNn34oNhu/ncx8t6+0Hq9zcdur8ttPuZD/vJOZo19X61Xtg3VgAZdLboVSVY7UrG4Nq8D
Gk8EYMPx/5wZGMe91yoAhQH0WW4/Ms7vAwkXie0wZXpzRjmYDHHTnU4AKmDMa7zKfC3zrkJTIrry
QtGEmmH6tlrRc2oTUGbCyjp3t4Pstwcr8k42FFEzrO3g0shJcM+hWzN1PWRcoXqmAtYVGzY7wLDT
PfKa3x6BD3FujyWC8NBmbz4AVh098TbGn6A0dTLm3JzzaJcWjkHCLgctzjPaUOemdNWxHc+rLQIr
Ez95M/qH4RaxaKXpbY91K3F/fdQyLxtxTRKjO5kEias4wBOim9iDOV2aHBLcH8PkXYAIn54Pw2jG
d4k0dGy9hJiXVrIuqH8LXxf9hp83atRPwLRrntjq1P52X5N71DvA0RwWcEMQs3vi+JsY9Gm/KTqp
vchb5FOCgZJXj0Kiw2ZC4DrLCxol0ofXmTiQ+lYbra3c0V9OjWMr1YNiBceabktXzN0FKyEsK4SR
zntv6nedl5HGR+0OsS54rxJ+hFVnaUTQBQw9OZAnFzdiKZuMfnLaVxVPkds6gKCN0MCHYAbUAkG8
d4T29OTLdEHQWFQDydRMkkae5IreWT7AInKTM+8btmFcI8t4hUS08X4A76XV+bDPmdnQmdldn+GP
hCwzwJdY5li+Kj3KbaRxTataQbxEF6m6c6/lx4Y3VH1QwZVymVesWRrk5p24NXEDyX17s3YdiFgq
C709tnMD2eDYItduXcvZ/x6OmdFKguTfUV2y+ICFP7QS2Gs9lTjaUQIdvLqq/39lrZb5OlCX7REh
1wsdufO9KP6+kGjRAxMyNGa9wPRStTxpqK5z7nTgbq9XS2OiIk1pExtnO6ykbXQ6ZPBxlAHCVajB
S5V2c9RxcxCeCbY0uoO9++lEXeImlIK9d/j93NLt7TVszXjcwY720iKmqiKDQwx47qh/O7DPHTtO
PYt2UymGsMHkkwuAlql7rBXhtOpykAvNicONsHPT/WZ2BxMri7BpHsMzDdmqkAuP4KL2asXwCLxY
mGyXDBUk3h7OTTJKUOk7BFnzQ7UH5hGa0qFAS5KMxLClmPEf0W6Q+E7lLv8Bd6QzwtsBbOQxdqVk
oVvEHPGh0Jj/oONeUgwha54AoSUQnDzedGFGNys1vGc9zuNt/RFGtUkZ2FVcZSF/URN+EFzxw1F7
idKvxbHtI/dkTszbpUIODbBDeQHJpmg4sbEGlsJUukK13ivR9OUTfPVmP5EcgigptWYrk9ejxuto
ynjp7YTYFMiQ+lBFfN0lNpGEz7rceMT0bHtVCvf9/cRlubzAX4L7EAJrqWs1KV9A3WsyUWXXTCod
3NGD5X/mIotOMwofd0r/JUCI+vobzTR8lemRN/pHOhKzNPayBJ6rI4rWAycLwVWv/4SecYDIf3Ib
lw9iJQDRCtI3GhZoC28tov0EiSX9/egjfYOFSJZPZc6oF/vril/eXSSaqunY9TkMHsLS5BHrWjtP
JMlXd1W6/J0K/TlquWxo4+ZZC+t49XgLkK/NkIh8SG7xjoiSwYBy0cjZlrvmJPbVoC04oZqmwaUH
IAxSZwD9q66mMqLKNXaKDZUBooA/ezUcfbCjb+MG+gG0rCkWGvMbB8SErYdfDG6stvZahHngNqhn
E6HaGXwaA70TmSwdshrNwflMAjJRLLOASfTcsP1X2DeA2yuWg2wT/nXhndq4n+prNSLipgJmv/qy
Vo+s1YrMUZ5PDW/1xQop4rz34Uass9laGy/S9G6IjkCr7h+/gbT2349XGhEHOuhBQ0ppgIEcb8KY
9tRnO+X3bpljW8RuuSexbB2m08plgs78JGZRSJzGylQextqLFMK8+fVyA0Re1C0+n6WiFWIFqrC9
xi2TUlNA0G5w0C2AWvJrtoPwPCxEALHfmBxFCaLgntYDKbJin7XNAt+h/zRlRIjE9V/3/YZ4cRk6
G5qsUIlTYLY68G5zRPe/u3DEYn3rQJItGV3a4axcwJlCB01PWZGYpeRQVvXeIoCxNFCCmkl0k5PS
kL3ACmWWKzLmqtTQyplkEoGC90tglAjTyyoNsvjMVEujibYfeYfR69Bl24akg5vGkzx+oKDQ2+wI
Lw0HZLxE8Rw4gzO/XzehpSNR3r9pLOWwXaw7+Nf0CJIY/UxydfC0nLzWigt3+WlLxABoLGbqjKw9
IsC71Yr5dZ8J8rB/sw6kdUjfp2MKALnVVBKbFDJQp4oGtjT5rEsASnJWyT+v71yF5vVA4gt5ke4q
Zx2DifipOIvpGCSsu4123jB6wDQv49ZS8xL+Be3G4ZNPGjoEeR48rQJRigvf9+TrdppLKIte1+Po
uf2vSruS5Ksu1dnAiLa++o7cZcaxtKPju+1HGvOFEr8rK7D2UIF5NDWwArmgAkoKD3AVrcH8luLD
/neGHFuMfOhiOd2fdef4prKzlarc8yg2eEermqM0P3b80/l8GwtaQyJZ80+YbxS4oIKBOQNhL2mu
NnNsmmikXUSFqZyTFjIhRk2zQuBQspAGRACCpuz2Sck36e/gaIyuTukPzct27H+8Z9CiBM4exz6O
98RBagT4PE/LeGQtjGkSqvnnuHBVK92N2Cp3BW4nezEim6Q0MqtoUsj7uIfZgWmNiPdNzyoH/k9C
iWg+lfOD7MqQe6qQBJcjKEEcSc2Tm2B9HCREmnngMhtFB+2OJHiDAF1CEbPcKvzRm/YA+CbgNUmf
9ucV+OY55yIoiE6XrbsKlpKARAwdD9Kh7HyTuWN4eJA6HlwQZ/HM02VaO44n+gyfqBwwPsTN0S9v
FnjfdsHQ5ew5uaVmryCoo26j2okeIWuzzlKa9FcTMwFgIgWxlEWNS3LMjXHxIGXGB3L70G74HdYv
LYegCvUvJib3kVJHxC4mtA+gRneB5BBFK8/voYC7e0J7u1WT7q8sAezu+GgJjTNSSl3+Wf4GunHU
5Mu9xXGzMBVPIvwAb50rLCLno+/za8IuKBHLuEO73LSrQSpD5HjH4YBwsCnOHKjstl2twc7EbWps
AtpSmDINTh+wuU2Ck4GOsIRP2rq9F0SUH7671QzAUMEnTgWq0Hfd0c9WrexTAvfDkFFcbH3+xoDw
lcM2TuYkKYJRK8Hkb4s4A8GgF0MBkBaTaWpSm01SpZNX6E4wR14VGW7cy5Q4Ffh6IMsCtEzgbe7q
u0+n7HNQuyjgy80SKJ9TinJiCYVTdbKjBUzBqQlL+RrPLZLxn1zei6+Z1DoK5RHRlhjnftot09mx
EvphIrngOGIMsi73sPgVsipe2m/fvlf48mYKpngrRJ2Gp2ZkduCoQYFWuDRAvpIJ1AlqEPsk+woU
cwoAEOQRqUtiYN1DJDvP+3LX52k4ZFSNytHLAB7HG69ykdOWKHmNj1x06/T7iRUsWR56Qh/XPw/f
MzA2f42NLfvju/E8eDiPoD6FEvbhphPCo0PlSq1QR4SciVcYVzunBbuFunFD4oA2A+5Ue5U4x+ie
oCFWWo8N86e10KhfhzpS+yEAJspYRZmiXeofjOU+8vsaoh13u05eYFaQw+lU0Z/DWONJlG9+5duo
NqGvfoGGvdh4FZtOH4ar9BaH/FRKv9WG0oQ3hNVcfvSgyaJUI8VHQ1oCvfiaWKlhDjadlcdzJwE7
pwMgCNIo5MOgZesabvInrtKqA7SwDyIyk8VWTRrkgjPmopqY/kcVYPf/ivqaCTsn0lQXhXOGo2GS
4YEmu25sLR9LEfE7y6cLR/80HCYQNa3hYjG3fmr31vRMS35JX4i3sUn9K7xeuab8lgYU36axP/XK
Hen+VtiOLzCObAqc7dfVd2w78VCAIGzAf7xYzqMdoAiV+SwBOGVUfspZAPAVqtN62lqZsME+wLc1
6Che2Tu28KF+tjt7fsgSH1LtoTWLuzUdyeciXLzxA5iioJd5xrMtitGaOW8Bh/BtPQAtsou++EtW
hi0fzEcjy0hSVt8115JbOyv8J7NWbz4lHEd9UiV8nD9pKpf9PpxV9Wzk1YDH2YTm5NtnsvfhqBI4
iLiGbRuzILpGWovjzP6rx3KpsAKE0y6oK+BxxnoH0hIET976bwFdOjjPaS96iOxdRIsT6pJdXOAe
1yHQR/ImjgeNyiAItr0Ph+qJn0BsWCu05HnN8WcS8zePY02ADryzVUTWUimRMJPcwn59UO8o8s94
QjXGR9j8YtyVI1I/b3XkCPx9EbsKlwW0FV5osNAn+AC+9THvT4MgTzW6n03/sC77HGGHFGGJld6R
WdBZfcu1LUz6pF/334KrT4AZwU46kPzfVknDehfKy+a07xaQqSj1/kSlGJW9t/ZzifYGyGCZKsnO
GDAx2i8gEqbgNN/PR72qZVSSXO9jw3PG4T1eUHiq9JWJ1zJoUGnhi4d3zrvnlHVDeUysqaARzTvs
CqE5xuej1kPg9ePUjFrQ+ZxejyV/4DF+CEQuAGNB5LG5tbmQLYZQ4Fn6GLSZPYIodK0Hw42yxMhd
o8UU4SGUqKdRzeE38EcgBc5+ukbRtGwSdWO1jbwYyqTOptjPB+RAOULwUCAxHcMwZbd3eNwUMkXa
y3CSHgm/sxVdJGjx4doK4Oale/2xegO+4neTMPSDgCN/+ZT59GHBiT7ZNTgeCcFxulCN+7LxaHs8
GLADfpmjY3tk6zR5tg6Dy8tBPxfzqjE7CDVkferae/JcJbehoodeBBoTOR71KGQckCg+Rcmf8u0S
UQF79SKbK/02VGUrAKB5srgf5OT5ttI1NIs6kH0nUxkiY+06zjfh/xPjJSyvJQ3zsky6A60QUlMP
CmyvD3QEU1qLyOCd5lZxmnL/WJDWtVcoi9jLUY7nP1baNV7h0a1BfbSlGQsmzAHjoF88Pb18HQID
RyMocNSqKaNzdjLYV5eLTDmoBzQa4K4L1ia90pGS+3kFD+Fq8LvDB8xKbaoaDb4uVo4DUdjzp1Fv
iMRNShuei27fgvknjZULiTJt94CItI/jSdi0m1IAO8B0S+4Lp98ePk3m4/YBFRq/roZEM67queVs
vpNlQyP2NkIKU9TMfxXI7ysrXOxJNtH4zHkMJEW0uEzX21eOa92J1Qoh+WQSXP5+LK/6pdeZ4rUn
OGn5gdcY1TonzJfOzPpDzSqHx6Wiu27mXRL+5QEMHQpm2SeY4wOJ49gpza8UINdY6pIHU78oEj57
cwPfWFSbQaZej2+3j6pk7DwLMFhIcG4Ro4TK4UHXbSiG40Oj2i2JcFZgtlhDW8nxT79ti4n7o+UP
oDOO+KQ4T6IZ7haJAOBMhAOLBkxnV8wMQjRErOGJPk5tk+mcUZm8kNAmS1jjDCW97A7h6QnFVbii
Pr7Ic0Py5688Q/x24/5fyNzqkY5nh0EqyJc57/t+ChnfMu4Rl9OL6mUqfYp5ornJElhXc4lP+u3x
w4J5P/NwXa6/+zbpp6fFB8fR9d0NZTMb4itkGj1jHt/FbZmbSBnbEyboSrvmTtSrNOU/5Lw0+DK9
UOJhc854DKmnDdfxDMAPvfh93j7Y4G58c91W/+OesK2EmOJNtIwLwpHwgopgoR2xqRxbTFlG0RyT
JoVl7yUKNhdYzZHo9kfTeSgNJv3qRO8cCWweofqhnHVziS5jDQ3vW7qNpdc7Ds8aIDg7zcRd/D2f
Pk5QIOGyTUq+RK9YJUYqLF2OSvsUTswBvjDmh1//X4s4S50y78/lZGLCV2x+5BzHP1Hl3w+3aOth
3LtrQsMmo6K+AsdwuRxr/biWGD6IgjtD3GNs3+kSLC6wRu6bKilI2xNfWQklGmILYLJKivYASoGw
eOws9J7pLL9v0AfeiHrCURKdZ9hTfIMtGkdYYh/LAY9geqlZBPshiS+yysxZXuHOL0REan5Mv7Jk
6iioxRk9ddEw1a4/BrSgI6wBbunongG4qFRQYEYLe1r+64SOfdqcX+jzMqul7fArh3/A2tZ4B/CL
GYQTlJ3afdKDhTqcHxcve1fO91eMFJrdR/rJjKXJVFMoNyAGzPpER1GZo3DRNdlzWx2/RILuUnpM
1e9+cZZui8SVP8AzeXoIEiv3xImwRDJm5spuol05YanqAUN01y0wUe4kjVPAXLcBwE2wDa9IkAC2
rade/lEuxWfdMBb/IN7YhOmSYqb7R1VdXTTKw7JQjrq1yxP1x5aBCKoAY/Nz422nV2y6ybPdwLdd
AVdzRlXtLhPxLzFL+kHJCiYI0JjktuLGeOM6vfWgiXleuMOtoWHGMkHZBqzbKCs5+Q6zGimot23r
3mMQlT6Ji9kYeOmXJzL9rSRFBohPvYtcQd9+9mAtfmBDu8XDeMJujULattFNVMwJYNbzpdEi+FVB
LbdqIVZvkBvyOeX8B1/rNTZbHGDRdazOnFiRZDOVV6gtWE6tGBt7+Czkv9pcjwEhDcG2KH88osjd
Vs4Ic9HWcIic7IIFL2Vt/7WBZ5wzYYB6+PG6iC590OkE+phpK4I6jP8UQdV/yfbwSeptxWc/bz09
wsWLV6mhbMjdYbiSnkaRlSFOWX67pfRXhg1H5Gox+2CNeNmedECjfOhDliEidYvtvam4HgxPvtuc
UZByFxjOswpioqLV3URzmyhfB/5PfAWyh97h7TmC7Zcp1Waw2mRXJjl5ywhBGQm5sDogUMLrpwnH
ARLtWNL8dK46T99S2uyHAtPEzLmKC61cDBNSv+OMDZ2ICi20Bl3h6/IUFhUFmMiInywuB/dVjVEh
99lveC8H6kE2uEtueh6Qptu650jK6rLu1Qrb5Lcq37GyKV9LGJ1ydJ7wpIJwyNLbm962qrAQszLv
3ml9OMSZfDqLXmiYbgT5UsRn9Bo4bx4x0zxb+Cv3dmJY0ccNQrzGgsMsmTGouQ55x7OmwC8mYafg
dJ1bj0U5ZbHeUaw37h+RM+15SnAxjt6m6ukjPZxM0N0UGrkMr/vw1q9Ux6D2nTIVnhXAiIW0m/xo
234L3q71hCFr/Zj4uE/Nd3KXhI/Ey2zp7cAYDurWoQTcA9Sh8JcNk5GgMMwzLynpYlBCUfOynXzz
cMb4/o2n+m9XosETSHwWhW/1l5Git2+5Mfysdp4Pdvi50kxjmHf8C6d8b0iXhLt4DZxZXC1REHEM
F6wXooNJchUKI6yNtRTUwCMxvKcPE1B7cuDCM1e3Xa2ZTiHS1QVUE2Uplzr8f2QzZFnxDI6nnd/c
0DBYd3qWAPfB6uXeg0OlHrxrWJiNEaD22SHUdwqoLpbIwq+YaMsF6Xd/mF/U9wuKw9xLiWetSnMq
aNCZVcAdgZSWRxERC7kvXEbymIgKXk1ru7qVPUVY2cuZLB+kir9TCH7bDVv1LReL0aRd11zbDze0
UJM/iRKa6zyC7tZ+WEPCxDfzr9o02Lhh0Z6byTnc4ZwQ0mFzfyetAavDWVSuj0BeVu0BjRloWAwU
/JH0O9yei89eKbkY7mN8xloU4JILqTJ4MNfi0Na0mGRz88T+hhVQxIJQo41UwGBe5RzaP0bt5GF8
x0N1Z3ldqFRJ6dUtGN6PcyfMImf4lau4vOtkaO7M9khjxCDYbL1fqZxnAKr73hrE9+84UYsCkQNA
kvfu0FA09L3dwYgxtIKQvIZYk1Fuw/FCCPQB+VP8twO7hvglLBL56QFFt1J/d7Lb+Aa/ZarTf7Fz
rhMwFCQR42MgnjpL/4r9PqSERKefmkYlAygm5Jylq4yeCegLC+yU8sEn7Dv6U5gzlxpqVlePIpT4
6zZ20CCMRrbVDiBJFGvl2CtcWXRBtQ2RwHlxR2KDkCD5ngcNzjJq61hHo0xfhyWhX5/Q3lDDuMXM
eqaNBEE2cGhZ/0Rw+hzhjZKQh4fVm05q+0ecDsTCxDEJK1qCzsMxSRNQMX4F9oNVVMIX/viAsnrj
gmWXnMlqAuSDxBLZQkUwdFw0xpVP1Eo1af//g7BQ8YL3KfycYR2GaQBBZ22Fdy+gxe5G0DAAaYsh
Odm8W3jlaaL8NaZcxhZJYz8FIJ7uilg8eGRqUZvHFAnITSdYvooNxAwJUhOlkfmoJkxGyXViJWJq
k6GY9DyvTMC71coaBT16O1b3nJ9wzgRHMxuAukuGeZtXHYBxVTQYIlT/1hxSzOMp4XCJ5JQcjngt
Yx0GFveouFLLP0/T5a/DWQ8KhgE2Men7+kMrMTCb/r2X5pXI6eVpsl/4Oyzayhd9vmIXP7zA4HBQ
cXZQkFqNlhe3W/9SVfaZ43O5ki6JslUMvQMWmbcve2MPSs3I4z0RKgRij/HhMOktHgvWLAq1jo7Y
h8GQxGUJwnVkcoFnLaYa/B7jqCqRnzxVsxTN22R/dDNHg9akI6YEwKKR8O2XFYelEAwTYnPwqCnU
EA89wwhQP0H2hfTj7cDm0AZ7hAd1m/iumiLxuDPCzmD9ZxENN1oA7RW8sjLMlCIXVQoAVEoMtoCg
zgtT7k1U6gG5vXni2gk3axVTdatbyUdWhtFOZ7+FJzLjXxhukoBwRXPzE59iE04zLzOxB9rfVdt1
zJDJuetMzTTuORB4TVdl7E25bkrrMdHqaMs2jGCPZ1spFZL+mlciFVM5gLcpYisWSkfe/8bNtg15
WwHEpJOA7Fwu/wa3y+ydqyMO3ZMGbFG9rVxisOOQk+OVNFHyfwCjgUuma9yO+eDzuQQmKqekM2Th
NdD++lxVGzbBOALeEsujQhlEMEqRThk6fLR0yPDcxW2bC9DLg1i2x/8BtabfGK8YqtmKU0DWOVv3
uO2/lefUef94bX0uru5rpvHwCkHTwERKKBMUq3Mq+N2hXYuQ6Wn86/j+IUkdpmLOpVS1LDDX5KpJ
M07RiTDbrEyVAIWTqJYddDK64eLOqwv74/A81YaA/lHiju4hK+TNcDvBaXtX0qpQW1Hm186DBUIe
NT23dQ1k/RtgWwsr1smwfwPm2bMOi1hJbpYxWjVx8OoRTPJRLyilBStrydIeLGIqRmnePGZyUury
HqVjyVR560v+O2h/nA67CwxUH/i7L8r2pupROztPkEknhZ4oBChMWCDDntiTC8TAOAx3H4aL7otH
fUeXPlpGXqogxZe28lgM/ZuCLKxDRwwBb2yhoa0axuVPIyw6zE9FyhrzEJpTlkP/P3BdOJ5kIBP/
mRTlS3ok5nE3MVj6dJANpjRnJGBIVjYbcpY6Nqj/q/Gy3VLeIvNNkNihjfrWXhLYiIWZqobNS7sW
7u0ruZENt/+QX8QK0JN1YBWc2Lh0dRSx4ezye2fYJ7GKKwQzgqVQ/h3Sz/b6zGw8JnSdNafJVaja
R9sSHZOteFgZSEDSjsTivduCThoqaIbDIVSQfC7lVzhVNBgsSpQqtFg/pZtuhvIMJbjzXcttFiQ3
K5IC2mEzNk5ZzkM56ZppFsXDiJeVzI+xyY85TV+TVN24NoFRG9bEcxJDIxdFHwkU7p6KdGk6lYOc
pQq233IqZrt4mGtDRmeDpuLNAiK5e0RTGvjTL3NInrIIlBuRtcIDenk6Q8gAOx2+1YqDPioRez85
0QnNnn9dVbgXReThzw6/x09CVisl96bnI0Qn+V6TjXQV0BQlTnk8PIE+8nMN2yavew8wa52bwLMv
dktR1oP7nXbVhK6c6HMEF/VezEJenWIzwtkIBql0JaFCqq2ITtpZHUYnp6O+ygiobzqxmicCv04H
/RAqroNs/LG/FlKaGyB0VLDlxvwXPIdV32AvBcaqBrQtCc5NNaWjs9+VJB5eMZPuJDwbu+g1n7SE
nZVU9OSrCfpO+k4Q9y36QD4QwPSvaCgXnFHmtoR/Bb00ItJICF0rZ0atNJORg2YerOAykkycF6cv
JQL8v4pOp9hYvY5A93IzSJ1cwH2XVMLpc4Tpp7Ugd83CjdCTGEZC1tzH4oFDkIQFjUd0C9RAONce
eiUNJiuDCSMwW93uf49GYZqclUPtDE7m4IE2c43ss6pRVk/Rk04nOBR2Md0PhFT6inrFyJ+a6Opk
qU4puFMnn1MMV/lEoVbyKW/1f7Hwca2cVcT1WqFdJ4qydXL3nLsnUIMf+sGOBjSwNsfcIxHOmIqJ
rxN2S8nIqJcTlYKWrEW7FzMZSDN7XD3bIaVk09qOkrkmmbCc8Jy3wN/e62jxJtzbDHX8yk+fwBaz
7NpRZDvoIivkWfb8BN20drERk4P4CcLQGyHwCXF/zQFUe9bPqG5b5s5mqOF2yvsNNNRCT4srp+I8
kicLyW22i+o/1qk1Z4RgOq+FduLjcTvhsUgZXowRKkEpiRuEn6HkHfYPdBeVRqK71rElJGEiJKCL
z25Lp9MAJxHN+RCrpN35MTpN7s1bzHynAVaT3ng4vljZfeKU9viadzNIU0sYCeotRJlousn4awml
J9LwMgeiL0c7kHeTOZZPWghXbpPM3zsL4/V3LSUc01YslKIvZkHQRF//QoIY52rbeUBtcfx18JDn
SxYktkq+TKIAvd25tKyCjqYcl8p4OhHMH9IGUMDrDsxJ8NG9kC08RJEHP2vGHw0E1qZTV/uAsfaS
SwRGA1rgctpl1RQ+540pHsXhQSfDLwixy0A9GE29Xs0EHWzTix2pjhjqurWdfAP5D0nsOLlmAFKm
c+kbVKa+RY+KdlsAIvc0LCOjViZXEuXTG896zAhkxk71tQxpKQsQJJDtrMGQ4AV0LvJPz9wS7WjU
bp4CQN0Ac9i81YMTkkXGF1WolKJpdF0lqQ624O98B+dv/nCGq1a+ST3qrxw8YFxccYI23F3Zur7Q
auB1ihXn0eQxvDwHugD4Qd1HEHQ98yNW1isZGQ5pPSqOKiKjzN4Q6SLpLHYiCwJ3HB/SVQxMLQpS
KOG0oOGo+eOwJOGYBny6PWI9VgoERfM1tOkBvznjaS+DbFOlyRbQbUcWYvgoDur04c14vC/OvVRt
d1FcBrUiA5PVKFJp0A0d8W+hvntfjRIjYNQtgHB18Y8MQ9ecMmq/MlIhMC4W9ELI73GwCxJd0Phw
57u9xZNvpe9vO8V0mIxWZA59W2lxZfWxdZ/759LYOEU+ggmTNpuxRPlttouTn8Qw1SAsnAe3mruQ
ME2yyO633zXWjTbQnhnPCxYcAw9EzaJHCOrgZPGIlu38kJeRyFpM7NGOIODAgI6JmwZbaQnIim8c
m+SQFBxuteghuKS9ovfVl3OJFi/zufu25qPstb4If9DAxpKdWRkndRelfgKcWwbWBsxOi8pYOCYb
hJq1ukDQ9JmFnxCglyXp4b8M5cdRNhA2es3lLeZMEfNPiu3kEFP0LSE13niXCOwJXbK09RqKkbR/
wZX7TbOXijhwibTKayXa6HAek/Op7iQxBgYpsv72SdQw88Fm+WgdSSN8ZkYGDUywOQSFblgVkio0
PrraDWCmN3r89NhLxTv/VSB5srGlvroJOjOzNfsIvyZsKhnEi2sqCMwZX2bp89RLexkKhpwJDev1
khJyY6+vvq19Jr8PPFo+Ka1ayz/rkBhiFEfSdMwj7Nvu9D+HOWjNty7SpDjrI2lFgePwwt5GOMfW
D3oDuis5uAqve53INWt9CadH5RiaXpVPfh10shG8c/6dgi9fUfMaLkD88WWfpEpmIYLoqpMwxRFs
RaCXiL0X5Hitt6+Qc0rhrwxbP0fbCt8DdeRmHAmLiPWdEusnlSiSQyvMQ8Td6+rfwYnDlrNd7nF+
jy1IQA+gjcBLFdPk5Q6x98s7o0/sKsLavnlqIV3qNaZixUmpSD9s8RlNBxDZTllprhzenYKKTQb0
D9fSNVOb4okUBL8s62+FbGBV9ji0L/+zzDVC3Rv8/MsKSA3L5/E06MDejBIwAMczIWBFn1jakMNO
XAV+V5zLRL/rvIv8y0EtDs/P+bBk/ha3wLVTUiTNtFNBiurNekaE0oCLITDkA8xLZJqUb2GxlNIG
lWGtJFI5P4797eNmoDp4ILwReNg1uC9W4l1n8isQpHAqvvVqW5+KdVSZ4TdYPjI/hbseA5AWcosD
TkQWdGmJj17qMKQ5lcDUyJumijLBFX9GJ9IfBIaPCYNOWFnHKxj6PyphCncAvrM+irSGGMkKu7p2
yRKIHAdBHFCujg9kz+RJUbuwLlHRf4iMDAl3Y9UKh0A9N6IbGKixe44oVgwV8vhoNZu19RYlkEj8
P38UKbM9MVedezc3cE++e57N06IIQ+cuBwErjZwgvTouZj7A5/chnKa559JWGcV1aJGL+oJbtuVx
tWP3eW/TubnC8zuZ5pI/6TFFg5OxSDgCuJfHg3cC48z4X4oa0vKDsMAkzgmfuxUMNtN1bry5wfEV
DdR0sZqohR09rvfnPeog/5kNtdkrMQFtsstdI1JZ3ueCdJDG1zPa1Y4/io6mmlCavgfzLziEBSsg
V3Wv86N2lbD798uHCQrpA4krXiTkFdMroUVDFMkQ2C/sCknG3C6FnV+FcIHSr3bbjeIaQ5kg3hXI
RKoanzPXywi2IQjGsHjSJAzxTmXJsCALeguZhfLS7FysD23IejZamI+9OvyjwOP3sqrH0sAImd7K
T36yj0y3eBQbwQ5wA1Tll91152s9YhW8+ct3nOD7dWO0ivwMJj2yCODREnJ1QlpBiXS8X0IKggow
kAS4uPQTYSRmYoy50dxn+EBXEBeJjDKjX3NFeoT/enl9dtL8RNWDB46t46/0jtfz099ldDnUDrUX
L0bhzoXVfytfyNSJ73ne2URKNjm0AqUE4AZGHslBHDKj289z/BAljBVn0QhMW+XF64EJkMJEUx0t
XkoFgSnNCne6g0B2Seh42finGaBUq0QazzZwtLC0hVoYDgMvu4BMYqQnVc6sAp1yeStBaKnmsR/+
eP5KxqyNRQ5Ef5J++JCY7w/+pY46DaWObWtoRkBKe2jOXZ/bDhSdegs5CZaXhfE2lFRkIWQsybIb
76KHts3pFEBkcB8bocEUl8RNp/ZbVPYKlEi8dQ72ceMWWd1C+jHfus6KFkvuBJjhuWbhCvzTm01k
D66GZB0IStSDjHZtGOZK09F3EJVfrPlRtJzPmeSsZEH14u3FUHZkOVksfg9eU2MhZ/p25eI8jbYI
rchqATSPURgRJky9xeXbBQ+2fuO1eJYx1a0lMfskR5WRIg4eOBmTydeOUOoOsRYL7FDWEjZw1INz
v6NfsAnzwmrmuiz5VX5QSOmhldxJio6ewJtb8EPstsGBnYT0koqy++uY69mCqtnBSsGCXSOoMf6M
sH5GJDBOJK41Rb6/7LLm9Sq1o5D7zuRCe1/+E3Vlz23dcdt3QxRdaCBBZGiR6iiiBh4/7A+HPrc8
WeSGX2O7r/z8rmCJhpiCUmHZ/HqYtEMv/EYbejIRNUEgzMj45TO/QrvP5+mC1sL/8PQ3FMBN+tim
kJCLirW5Iui2s6O3J1hHMRqyHQ0CmNI88J/u+f2YIOqgokAZAquPbw3BrzPMTZVqGScF56UjmsFi
Gt1W9LtwuSdMnG0bRfrJJ1WiB4U3Mxfl30pLw3Yg1MC8NVfa4sglpgNluuoRQUrww+09sca/0Sut
8RJK4A9dSCGa4SgFvHR1ZUOZWvCcTMiLUT6nd1M5g2fPnZ0Z/Kvhl121ekhR5JjPWilV+vER9FeS
RCRuKDJhw4ReRtb/92F8yoRqonH9AmTuxlL472LTgy4ieBZPQ4ui1CiIl9nCoeJ6fbQtXDm1XFFS
aRd8/6D/hbQfMU8N/zhtlli4fcWJlwd2IiveWyBrsB/vcwaa86/tcZ6hrIaPVdGiI3EAMpHkTFHb
pPLBDSjWtzlex6cbqC5N5fWA1WEqIeqLtL9J1usUCK4Lv/bOuQy/fejsjxvYHYHKTcdjCtxHRAqB
VFxkc1HU/d2x4GwyYIhKLySzxB1py/co2hrJtIlednapgQamI4TYARl3e9S458EsVkAfaukOLU9h
yxfGIw81wUsKFo8X95iA5gt2yRS/Qa1W7goxmMcsJitZL94GYv0fRuTkTenAz82tjAzKeKDcOofp
bIzz5+eoMp4WB7SK5fPgxLjJ1kt+gKpBlyzIPM2eO2W3vACf0DQ91cwr2n09ZYieqcH81lVyYa+o
W90Q/g1NsBrYLf99d1UqIAeAIHJ8Y6wOVRYyMa9ngZi/SneJ1sid/TD5m4T1xc0AzuVdaMHnI2+h
XZYp6XRhYTn9Nc0kd6p45FOZFDRX8CRNXIYEagvReXgOBKS4VGdVT5p/o2PGmUqzZc7X13XB+UWh
ReOeqv0EsbGtjztUIRLi2oqeX5eUjVelt6p2pTs3GITlb9G6DjA9ujYrEvKwL2m4AYluWYSS9jdk
ycG4g62LezI693znu083bt6a3rnbIAINBbufzejuqJyU8Y8vW1UTCIVSZAL2Ei3hPX8BqeZjmSab
gT6ujQzD1nm7K+YaJRVj6g+mMwPgQ7+uuDQ/Hi4TQXO9cHSpuauxesZA1KSHA9QBl4eLT+zJRkLL
UXSLUGcAwkm2pf/HTMfc6jSAEy4FOaVa3B2bBR/SLFzxwYWvDR4MfMejh8sno+55Q97zchKeMvmM
ZtxOZFoeNHwhK5lfxm22tckzjb7OixOzJ7wjJ63535XUYV1MVHbKqQKb5CpsJa6ux1E0+sfBnzvk
Xx1uSZIhxqVgSkbL21+Ts6KjkjLl423HRLXMooZtMUzUvifs/vabPk5MlICFz+yX4cJbv9Jv38mV
RZxrHGgMUqYkcDmAyuUZGXYn1NUkoO0pKNXvL2Jy4WEo0+NuV1X3n0GEJ2qoIeNkCwXgu9cSoCN2
IGsNTsQzJ5ANAQIXntaKuTsLgAWm428zmUkBzsIWsN2qUCW8GQKSWCz9KWw5jERJYpGY0rdHqloa
QcOWS+MW3v3ym6H8QDAx76ytKoAzOpO7y2hwQuwNt3ph/kLoc4A/IS0fGLVIgrKXqAAsSAPb5Wbd
lqergrFtnKA6ohvW0X7/XhsFGwqZqaOd0Hhpd4Eq9+2hYy2KnxJOQgli/z5vWzjy1UNf1RdP/Ntu
unFDkpIBmIWPXKgtJvjHG77tfUzMnhk10vimKGPfogkHU7Lmj6aJlttC5h4/qlJcPXZZ3B/PfAfA
HLW+FEwxw1SzgWKhCNSp8gP0/u0pwjRR4Hg6/YqVaYc1kTqBW5eneMeijRtfw9HLiv68cK/iONuI
ljPuy94YXFdWpyqSsu8Lbz3wPOwT4rcSaQmVq4vb+7WRlqaQMQMi8RxN8jP7ZU0mwmgGqEFyU3wc
HYu1H+1q3CK9oOf1kgVcWsYirGS6/bAZluuGOz9OGC1tsUTyNs/ltbDfqmjcMru6hgwliZrjrkoL
1XRFc8rBiOp2sJUZ+a12WTCTxn//qMJhc+UbjCHVEa32hnKFCnCo7u2B2lbRICDWcXZxkN9VfWd1
2qrSBpxmPnyHCTAJe2XqMumCuqAavJ/4jLU07GeuGSxKxt06yhdTLMYKQQ08kiUnqnlw7sjpsZk5
i/EtZOCVC1IRcGB5l+S8ucaC63yQIqrKVe8I2vkWRLrBA257Eo1/QLaNVDi0I5nfLudXC4agzQsO
wxSlCdlr5K3Q2s1AzaceDj7SVuoOVh/tHsJmeaLRs1TdvPjVNbW5XwKSw52y47zgPCPpdrdpFVjo
11QtrwURecFKJDyiwCgmDqgi9jFs1Bp8/rl6m5Pjl1LEXfGEZKa81gunKUT8FtQ3qK4xQhoI8OFJ
XKt2KCXdtHfPuDKrHIXyf9fcMOY1LwptLrEU2JEGF9vdKu4++pH6H0T27Ss6YnijLIU15cpYc7rs
7wVwOyp8hAFabf9YWJCA4h0iaY3UP+K62xvPIvZhHKK2EiK4gbKnbOgd5YoJUSUcMshold4/STrB
HcRJbrl7vQNbKWH4zUqrrByifEbtmnZgV1FV353V0xKvKU/zCzpa+E//zlMeN8D68IGbl+Fxhuw9
wBn/8tnXeuoQxtZxK5rTwO7AqVpFLivgIUYRB72Nnd/Wd52NSgH5gZW5Rzdvrj+wRVMEGVtYStIT
psnO4eSg3fDelTU7ZiLfuvG7z4Sy4LM33AlVVlpYvdgs9rKCuAq7vW3PIIekVyraT50nTs6Bddvq
XKD56W7UwJc8lzcQfSPDiT6odqsO2v8HGUJOxLM13UijFGdVy8biToyH4X1BNHkt99nx9UujlwPi
T/tBSw9fXVPpFZKYB+59fE96e+InFDe+BId2fGuFItDmQNVLCrJ31diOH/kZUtyNXChnH6buF4Z0
lpBOj3UxLhSwQlBHtK6du+0U4reuPKcIjK2AnsdovTq7EKM3zw/k/tuu/eqB84al4LJCUsDfkbzh
lqTT79Ow4JBqwC85iWUocvFdBS31yMrvhodEt9yQjLfZOyXmNZi+bR0+ctU4OVDkPelnw5mfh8pT
p9DHCEN7uyiy7CvhlNlwXxta8al5ISYezPvoNfrCmJFzetpv4hd+TQFT2lLCUV27GIGRTL5l7ZAn
M9MIlZrw/hOI+QkNnH3GcASz+TZJIzybbaZIgln7mcFBuhsqeW/CFvWvFs4w4yFqlQfMga2t1nNi
rHSISMiWXmEQV2r74TKNj/qG0ZtAbrMkFZYOHLUqz0kIETUoNLTzh+I9qlMDvstsnp1yCeDNGxmD
Xgize4u2mhC6QWXjlckruOc+SCFK2pWbBpq6t0BhRSLtHruLFgu1EPR5OwTJOXoEMlA9ER9FEFoT
dAQlXb2b9uv/k9t1ILpLsDHlyGgBwbZnAXLnxTi8G0YajQ69buLGyRpfJvd8Wvcg7Vnba9ENXgJ4
oFqOywOyD4hBj7k90iGTHfr1wEvJK0pHakmtOXkO6x/TTpFvkJ9pTLlvIpb3qN+hkkBi591SZ1/T
hnuZRvPY8fBqgZ/gnO4tVfz68hlM9xw287YmRKVdmhk9gr7eKITw/X6gdthgfUeawRCxKwMsqGab
E/vCljr8Kf5iPV0GrvjSR4OZy6o+VoV1glne7a1waYumivEIhTlM9mi+hIXrZdGvn75Fcee0pfG2
CVE+DALiTbVb2XVTD1+L2Parg+5Z4BEUXWLTMx4/t2lRSeb1oJF5Jbwc0uCStOjybp6CplAiXFEi
S3Gpbo7Moj5ko8vshzMlDGTuNnH/h3RwijS6gXRFirbM12I3sU4DPLOJgsWRD85I+zyo+295diai
oU7NS5JBZzfJ8BkLNUrh1xQtXYkiDwsG7paFYdyhb6So9v97LniqfGGyvT4dEPk/r0mPm08mNvn7
RYUxZ8LIwAmH88Lv0aZ4aV6N9A1OqVsmnIY6QxPhe8SUjjTkb0kd/sGp13sABHowhl4nDEpnmk52
MeXc/QJin3XPS2YIXP+eqL9h87BFzxtoD1dTm5wRCcKulcfTEToqaKU6OdRzN1hb7NykdUdvQYsb
n3txBLSyiwxENK5C5H19fjMdggO1KAc64k418jYAWiFGatRMmG+3FJokOqwZYrdOpA4ra2mdWtLs
+KaIr0M+tqhcX/8FPLnA0dKW++8ItZ2G2p9NrJoc+EYGndjYDBHY6d723GjxUZSdC/hQH7q/1U6s
ucqakoTv08UROv5CtwLKl0V0wTihUBoC5huteKbcUYmR4nsqRSGIlWrOQ//zQiRmpK6TI+ZArKk8
mNoWWb3mycpDwf39CoBSZddRokKW7jDMqQ3YVSfNsAcsfF1wWqPJ30+ZgmR4b7/JEEHvg9LYLZnP
0AX6o6zWwZgw5hTBIl18A7AyPFQRbaC0owV7iubP1JNVnQ4Z5i6QVTNouyVfUCDL+Ff4ThOdEC3c
ylbbvISt60fc7o4MC5g6Be4yg5QRi93GK0KTO1wnyVmW4L1dWHrPTMcUYKrMtOWsi3lEaqX/Mr9n
P6rVX2uSQhPJA0kNes9pEVilkYROdNpsrHjX2xaOMLZlKDckY2XyNendWDUjnGwSfhD54HIrTrnK
pNfsh6GTLe93MUjNIyfmI9z1t1JwHCqzjkWoRJ9vHDRMtAHB3XUWZaU2ObOyY6hS9gsC8NNik/KJ
CC4vc12DtWr8qyO6+SrQBbx9uG3A1ZrJRVP3B7siId/6LkvC6HeUgeSJYSSd76w333KpGcK6fs1I
mv+T/q23jzBjWAMS7xKI5d5jI7h2kNqKNU5+AyFXnE9vYZTIIaHWKAERp8I2xMpGCwfhMUcmDF8N
lm9R3kNp+fmiuelUySOmOPZVYFrkz4qLP6o0UdCdzOwGTjW6hOdqdYuLkoXIWs/KdC//eE3CCYgB
1Yer++KXS8n0HYAkDhDX1ZB3H6//8qBCKzjtBP4rVfLMg2FhomIg9/O0fuJ2Qu3rMmw667VbY7Wo
ABP/pqp5V1HWzPIwOZ+Sd40rz6PvfS85iYwvBlal4GoXP/0JA+1DhNEAZnxKFkts9x2ltuTPLfoN
BN2uD4wSjNMcA+fGt/wgpHe7UoQ47054SXom6kEOrBVs2Otr9voNix175qsvxFgtSVozUcqBdql+
WH/pMW5HjJ4+Mgqy7drxvNNB89/sSGN6HXRRbpi9Bt4VA8++4klddqyGHVxk+Bd6wVTFdPV+ceNq
nJ5kpZBl3fgYiDB7gkDK5a4OaexSCqZcf6mDiC3uldUC3UAKLzJ5iYFmZKBFfc75pfARTbWpWErV
2ReXs7pcSO4aodZCHXH2B5ZXyrqpMGDTnwcUjFl7Dlw3PMCG4NRxHdbouWAK3n3mHBcdD8+F1xqC
V0xXq3LmhMSo79QgwCCwWwhHL3GeUbqzshtg996kQ8R6AZpEwWf77DhBxwInogqpVgGN0PIK9pok
hOYAFAjHjsl2/cwiGmPGlV6Qd9zGwMymdosw19jI6CdpoIVFGLrQe6qg8n+uQKtyPTyFVOy1C1ab
3xuLcNTLHqj1Ik3/545cXsza2XrvwbQ9o1L4Ls6/6w1wDcCwBOo5Iu7RYPVwJc9bDC3iABNrlmtR
lYFJCm7x0Rgi6ZFMcp27+3lNqxAJoB90phQgAWGgLNCb07wJpNUpcfiP/n2Q22vmijLScyMu18p8
5zkc2yPZvp/ToGW4xIcULGAhe5N/41Cs19+w7s6owTtPrrTzp/Thnq9qMeOmvnIY7EvBcPakzbUK
xvRU/2O7enVW+Izc71y0ekOaGcJTVByz7n6l6LNsjtZrD1pxKxQuhr03p4/ALr8MyJzsyyl7F7mU
Zi4OEekrWxc81g/Eo9zWGxa4OuBJuyd3lkaulAKkVtkql0yYyrW2nW/dDRdQOh/pdexax+CwzCve
njP0skm7148ZDKgnSU5JmzP8wkp9vRNHjJEaML0xCODpcTBURG5KoD1WEWbMu16rf9PFg0l7/0ym
siT3/lYpOUXEPC2/UTSg8tyPR7sjkb3/SBXjo7hQsvfaGSPmkJ6ridn8rXFQbqzsvtv9MsVd7kzn
WeDm8qyasJ06MzZKKokxJqvat3hFcag7dpgAcfq49Apm2PGr/uQtcF07MmMCdRT+v1DZqRDzu4lW
Hgex43YADiz9gWFkR3hHLo40t27P/jekSCtzDiGxGxwTVIJgHu/lGN85L/saMB2cjmQhykJYjHKz
zObQHX0D8JWXlM+PHe1pwfTWwlr0mNhhWHs5OfEIIIs7k8eRCDbXAiws3b8he6R8pXvT02Kcu/Ht
68rc/uD/4Kn9tmGUXh3/uRde9bfvmGmz979Bi60E7npIaUysM/d4LNX/aI1LOWzEvvLCYzrMz7jr
mAs61lvNDBRkOlcgzBtKrW7/XzvRRC2q/S5iosawfRhbxVnT5VK8isrKhYkBDbqzJREqnKMkmRw4
ezJ1u0M5Oz8PXyLH5WxpHbUDJFnyI0KWghgGBpXbzfw7YiHPbBXKypyPlLHIqDCov51lCxaRLXov
Dmv61QXW4NCfrT07yIVXfqVpAWh88jTiFK9F7NvNtkzgV43/SqgdzJMvgYf6fOUE24QptOuawz8N
O5n371jxgrrhZfpkoSi9n2RzA4EorXe5TfZ4iGNJw+Pxs3+ubCsvYfzawJkkA6EgNg7i0WLXgd2q
HmFCBCzW6KOLx4Tv6Q0cSbbkMW9K9LVnFJZ+gVNKmzKAN/mj4St9x19LKA5U8XzF6LbTZQCN0tc1
I65VSVFJvcVjaFxUA2bEVWPOiJ0UIr26twXNpthvCJl60DvOEe49ZmQwoAJsciSECSGdf6vz08H7
W0loNUnmVaMz8w0lVkgEACIL5eIAvDv5khMy3o3ByrUBoJ8+GmZq2RDalkRYoh55URA3AJCJ8IPq
h1FHSz4eXdtD9Wow2egQRQ3QZYOytneSykPRMw69ZVPfL0G88mybFrxibi+ukE+muyT76K0T+qVB
kFXg8rZZcwo4263VpExGHjHyDhkHK4AR/AgFD+N3sAkifadDWj/dtOY2rBYk+HVN+cz94AWWOAJB
a5SkdqMkXCIFeHXGcQndnomyUtAvZqMKA2ghLhHW06cK0rddA9M1sW0MDoy2H1/5AmbIskb/2T2R
XpqtDL5xiiTf0m5eFcHThrh0Mz+IQ9ukmq/BSRRg3RtUmvyLOeD/hqpSSOcJrjDbi/SGncduWJwE
4tLj9Jb1W1xpWt10vSkMSs0RDUUuv0l480MRGAfeqAlobuKoNtsMZM+MTCBYnmcHxrkfTwJfF4MT
pQuyzcLClmuFnUUB/H/RmYWZ9BMcYMSHQs0rT8M4IWk/s5T9rtkXQFgL4Y4NNhMeOg6nMHYWmO16
jFZGB5bdiNEhApVrK+zArJo4wG1pDCM6mI/DwZn3Q27+aBMYEPFSNWqkJfw4Avr9WEySzSy0EOFL
pMOhsCRp2dQU8oSzZdk+VSX6l4BvEwMrJDmv5+jLWVWaWi2fT1mzbDFATsO5lFs2Igs0Vs28Fv8v
KoYvvCjS367IdiyPfw86JP+xtrKez7IAhuUkg+QYUTZm+H7wnknItpKiDmi4qozRQlOl3lrcfJvI
IHgh0ivCuK+5wE0U2TkrsTv8sIY0ksR0ICkr5G9r1vrR3KP0lAIcUenabf7J00olf8aSPCzD2/Hi
pK3Yin3G/h+mxdHJUMlF9/QqEsi6q+yatiRhAyenQ361HvlOyi0XgzB52dQeOBNwbk3JY2tD2hXq
w9WTZtEpi4ebMvMOthdmFANGj3rczNTcjuOtrnKkgJ+5nSYs8johjYBj4zu39W6n7n1f08VoL5Ih
eJYyw+AKd9az+xFjZwNZU843kIAY+Ks5zVY/1pSTefZes0lHKbaNI9O506ooKgBfEE8iY0XJYZ2Y
W3PC1yxpTafKWu6M3UzZsvJChsj0zhABj3GbU4qJahrTBM/Fa6YYM3maQ508Yu/B99ckW6yTpgPr
Tf4TqIHbpbDwvSvm2OFvXSEyMlDrq3OBKl9KxrhN5vdoy3d6Gfne6Hd2vZ2wI3DIXnEdL1PunnNX
PtuA/vCnjWXU5NoAPObjZ9eQP/LpLhSyV8aDIpKIMC6+/isT/0cBV3O6B2ebSofoa/4Ku3zaNOY1
2chjhZyUYvp6PUFOUAwNgE5mPh4cpEblgtyiHRoMXhExkUyAg2VMygtJRc066B17T1uXHZCi9SNo
BFgVAI1Yn49Fz172uXrS2WrwzMldBl/weR4yXhjBatVHCocjwUqxSkxTfuO3xAMxQnA4QIaW/RKS
65TZv/PeHA+YsscD2MDSlrxzqLsxl8cFWv6CE9y3kpz7hYQYJKs3CmxwhGIHS6zzm8N3W9Bkuqfe
AuVbv6uaz88TumXDGqPoXZQoU5Nx9oXHZmMSS9Ulq7QnypT8+b7qJl9z2ufh1L/+PF9lcnbE5Ct0
SqYgqsylGwvF3eKW5TVSsNIVdDRn4On5IcwEbjYXmOINofjfCRbYpECRm8pwumt5VuVaY1ow6FXO
m9MpI6R69zE+JuDqs+QHlfbzHfw3vs+Nt4w/vM14RbGgO6+LzFx/eyqLIBcqw1m0jXc3qhTz6eR3
zg9Ckl6wGf7XnZsmQ9Jg9XzK69Bz7cIA5LVD9jW0SA+Q8ESn/Q9GUQlb8RzxVSTumctPDfSa7gFL
h8LKu5qkN8iPzoEFBK6RJBzUQlBU84G0YrX/QXYBjM3yFbWO/KuyzPK1f6oO1nyHRg856PrgYb5f
VZPdUq3SwNN15m2ZN2S1rwPWQdFX24QyO4UOKGCm8AkThiwvmwU69uokvobA7/1cudhF0DRuKb0X
/d8sDi5NIpX+bZL3ZU7BNPJcbEp68cDptfWqS+eAyRQlfEZDPVFSaIhfSrhXWINZ91Ns6uhs3f4b
SjxjG+Ct46y1ybMXinpIWeHhNvuU/iLjFvGVWi9Up24EKFfginTlojzJz5QXX4bMwh1S2eCzD2Ey
tgTdn6Ba9HTdGHlglAHe0dJlJ2B4L3qS74SbcE9KxnW1/GeuQilzAH24MruigkQhvg6+0IHCF3Gz
V+AhwTO2eNua4IEACV0uyDpCXRIenBToI71+D7jOA//onCQ8l6FdJVQrzH+AKzTxgfwkJoTUxL8W
GFceRfiMrvP/gKFfsXie0XGZK0iftC31U9RKtSvLn4cAKr1tZ0WxvTGJV4/tHmmVHe1jZn3yh239
ZmxH6oKRukLZVPz7ju9cenrbegmbYbe8TM/0SKpiIzIEyQLnzP8pboBTPcwWyFAgyJpT0le98Chl
/9l1BBglMojHEzVfZoX9BVNLobxlBiLRY02LFq92cwo2XpHY2que8HtMcv5Fb5+NamkWBEIZFpWE
E63GlLB+OalfWSOWh3Qvuw4OTy36ghGTh/gGMEQ0V41OwUEV7y+NWLv5REs5MeL6uS1wRTKWYgJ8
O/wThCG+x/vQJE/+MnJ6XVUrhpT6bCI1yhStRy9xUsKJkAOG15Dtna6Tphnv7NAqVmRmijF/sVCf
jH8oW9LDL+7pvIH3kl6iYcitHhNs4SbtgrZTEhiQOEW6iYguG75hGlwUvECYjPCnFbr4zZDH61+M
m9WRdCoq/F3YtS7dMOLEfFfpmmHc3HxFDWiqhUbx43kXWBhSNT1q/jhDePXqbQvy6LwU2K50o/Wa
hF7FTVS+KH+mFW5axwtbT2yLZRJqGlNqD0Rtt8VbkUOeB7dmLiDRczSDn3mWeSI3/MGzkHBnhKdR
3o2uCuAo3yjUklrT7mO/XVLpFLPbt5t4H0oS0zUEh2DWonqED5OLEdVNlMoLvxKBP/QAVCyiNebK
yND0tj5j27lRowlmbEnuf6OpFtEkHwzk1gO3BdttYhEotJTw034zWm0dgzRX14nubcHV6Be1m1fG
feACjDBIwHNSe5CG38nOc7HDZWOySmUeSRYcZM7K64efpSDhKP1F6xyBibmZCUM8gC1j3r2VUD0Q
88razYxZ18aL5k1bCL+HF7I3+mI9H+5axrH+ZrfhPcE7HDFQ/HYS8qfbDZ7U2PsdoOqx+CeXXS14
KT5BvlTwYcQ0MeLmbLyfGFFg07evKOIzPE3w7hnIhwD05llxoLNTBrUqKc1toT9+VMrieXO+WR96
SUBZv5x+foibNjhwGO9WeXEDmlC3HK7VXOmJo6wc/ENWnZJt4FyfRabu6w+a7Z5pU8coFqw7LtEC
vWJB0fRHqPbaUxDmplpDWIewNzgZDhpzbY4YMi0y3eznChIQL+XRgSU2KOfb70whUWziYhTDYjLy
oJKkwH5ExldYj4J2UZzl+c6pGxTBDy8jq8p7VDTHJJ0pXWvsMkJs8z7wTnbi7h6tJzh29/181uUw
nd+ENbO2W/FhhH7iTxu2LOXTdQ1jnQ/XKefBURNbhSBWo35cN76PBqJHaZ2QlorXw3b4P/yqKxeT
NxrkNSW4cjVwNKXQ2cGb1XL+ypd6KHev93xUmTK5n9dVwaUuzeqHWo2Jj/iap1ve6slK3d5NmRXW
FgL3+s3v8iPNRaHP16JqAs+g2F6V360zbixCd0NtKVLdT3vkQsLooW1egwZOSsXqW3YLVBrl8TsI
9vMc0AHl67GGL6Q0b5nQ8dHXxFvdzRBrGmNghS3nhha9+guP98WTUfSV+EbZQ8fBUZAwl6zbmQ3R
qHok0gMteelnfLeDrDOEMK6nWgjX+Yq8fM3hhNqmkIJy2BoVgKVtaktq75gHwiaRxCN0vhb3Lgai
pCTqTDP/c23LhUbAWcUCca61tNRZrKQno54e5kgsOuO9T/mZ4kax6ZcdVSmpbGLYMvfyEK40hTIx
PKc6nxMzth2xLYXWzyHAIbMQj8gqvK0JTJPOZRZ6Iw+5pIA++fj5puh97Tv9+I/72Au+4mDrj1yw
8WnTlDjgazH6PC6+rUVSUZqNn16+YX3BsleqI+mG8yJT7vg7Dg3Qynjfo6dOqOMTTSWDEW83zSh+
smzs9A1IgXnnR5Wv0MKxYeY08ld6Nge2wrbJ0B+QQxG37Bb+gEXbPg7RQMdTN9EUKcAYFaH13cF0
6jwT5LAhWcWKFWALxuvvSgX0fS8hOtLiFxu1dhbdIvThGQ1wiuYObqCXyEL5wO21sbHetuODFK98
+CuPUDYy9snVC5wbRwq14ipd3Bi+hswaVVkVjN818FzbK6TBgLaA6gqW1c9Na0aXxp800jvSwxuw
GhFq9eIGQN7fm1asyid+dYB//m7SPsPajmKgZwEWE9z3Odr3Kgo1028kpmPPGn7Js3bz0ZNv7BNH
KPNMhZXch+IaZHhCFT7KCLLkIvqr2IHuhtV88tspDj22rpvVYSYzaMAlkyZLqKcWmbHOIdiaa/3Q
1S7JWdV/ReQ4FhHMQ8eiK5b6DAlZfpzfAa604E4Oyx6hlVkAbtxg9SEMVLPmgYDIHaBp6UZKcjtG
1c+VE+SNJ1eOFNFCade6SWBTrgiq0nYicX05z6JrxWeaCHHjlmNNbv42Bx7dsBJciCxW0id2UdK3
wyRN0CXJdHqxEMXqe6Yru2XGnjiqEClVHGhcwLkcEvL+43Db9IiiWbQdba4K+KaTCVnEnIsuBVV4
uYJiqmZ17n7OQq7Mm+5d+X6Qr4kg0zGb5kc+mgLppjxLiRM1XWlIV2PmIMeTAtikvZpVq6IJ9lrt
elBTPtArhEGBUErWVN6sOmpkRAXNq+w+3qcr57GbPil+sfLBctl6V1Q9HAx/Ixmec0gy2MKnN5KE
5S+Kq7Iwpi98r9nW06ocq2wuH/Z0xbf16J0F+sOVOdRc7p7P7MhGNiNH4ESOdnvRtIjHCkleq7k5
VS6XJPMjB40giIx6K53x/nLENibVlCNPKfIFQb2ql+kEEpLuVDj7T96U+G2/GqYMT5rTa7g4q8BS
Oef5FWknr0i1H7fTRbxcAG0OJpCfVwTV0ApjN9OlvCgjjlxvhZSYPPUa8kKk2/1jAFl2GhabcMQ4
pKPJJ+8DfOG4Uu9a8O7wA+InuHp0NOcvTbjDZIhLtwd5cJKSZSHoH3a3gLjPSEZsJMWSpUlGvfWK
v5DeK1gwHwWrKaIePbjceFpxMsugHX8IIkRmZmtoszrO4mMC/SzvrypF/4uBGmrHJaQihCUla0xh
H1EfeV4UUi+nJPkRmIVS8Z8Y4J/gWUZK5nB97vBgpij8uztdqXA1pIni5lTpS1pWnh6NcZgV3otc
aQ+FmARTVAdOp/WXkipY2/qLegoOyHu192ztSiobyf51GJRZddhmI7tKO1NMgc85WKPFsSNCM4Ys
MpwSDHmOInFQXcuFxsq2/hHU7sPrJcGbaZ2LY2xl3oZk3EmwWbODBe2/O6ewSsXlfIlHhz05QNrj
xEZL2q7wiDUdse9BRZNNSBmRIVwhN0i7GIxksrp5MNnManJvxdcF2C7gj7KtOeAv+ImDaap9zNfq
8ZFMmpUUjCjS6dLdbOkic00ziQA3pec/mVak7VKDhwZUjzALtSkF6956RzMw3owdLub43iZWWTnv
F9KCOV2v8lDMHFcyASPCrz15tKmbGSEXGpcflnMZgmCupglQfe+lYl3a0rjN3BSghs5UZPkYBa1D
v9noAQNfU+QtsSVo2yjq+WA28qD8dmRJjQ39OT6g2Ysj0+XlE+IDDT8sRS7Pgt//tBQMGHPsCbSg
PgKpvVBgtnixfnFryXvp3EteOjpD/yXPXM0KSbmqCt6VGX4lP+4cMq2UNV6JGbLz75+vZcZgK6u1
xv2dQo7SBro5QpHP+qBGugEmeE6k0Hwfkp2D8+ENcO5yyX7s7MO+iy+5ZU//Pcl553h5Yxw+nM6l
EM41V55hTK8BNNJmE7UoSUXpu+ab0ntIbRAdRw5ZRTsGfnb3MQjUF/R22DoxRJzY9WO5bC3QuUyN
fzpmNuQblxF/5r+SNUNErYlc9SYP1hJ1tfcTKvG6UrL6UT/igHXVd3CncmS3uwef0/wExjZqyPNc
j/zozGlvRiDANENv/jdE4xRnQ6kEQZJ32yJGiLUFvR9L5C+QXEV7mY3VfaqhiBW0TCbG+W4Q4/85
HdfR+drd2aTBRx+1UDkbJXB9bPEo3Zt9qIMj4fKOMinYp7lGN7fL+ObfSCICsnpsI3iXkKCPQqNi
lnl8uOfGl8rOwVUlKYKW7P47CenEO2gJjgGsYi7XhiJo4drVwFGDM4hwrgE/n8VonV0V2gXfBqAm
Fcf9LApc/CywPOFqfVDhDQc9ltuo9HxPmnSeSN0ZYvqoCJmZy8zKuzLdpNVOk8Wa9WIreturycul
bxjacWfXJpjf2YJqe9nNHswxilUtbmNbPP8ghla91z26CH1LklTgSGpZU7IG4Wyfg0UjN3M8j3D4
Z/Y96sVKrmfRtQcvVUjCSpobPWmkpMOqNbOw8mU9Ny1pCG5al6yl1R1ckcBRhlhk02b+tizdOeND
NSfnsBOWhVegl8qI0HtUwyvQaJnGhskl3uaNzJAOpmU+ffcGkH8v7gFL9MQa6r3bbLXQk0/czwaZ
jxvUweBZZpIqgYzFg0TI+DKcV0AJoC7tm3/U/4Ro/XDuhpWPioow/WsEPDt/5wy8ULvdRwZto3as
CULgM4nJTVW2JlkK4arV4/sOtF8PKgHucQroJnJctpxWq6BcPOo4g2hOeouxx38LtuXkaeeuGpcI
cjE/JOAKKEzWdRxuoCPNevxf++82TiDY125eVfJdQROoH8TmHGg7cj91UIU1/vRfgLg2HjX7Q/rs
xDcWA+uMhm/JOL+fpi/SB0Nidu6x6i/uR8+1FVygfhWPjvVjLTBnOerU6AmXAUTa3L59wbDYgpoi
xPYCySvmrMP5tut9CE6c9XTxAjfvZGiWy0l8BUJ7AWjmOe5KjfjdhCV1bZt/gmxgfJN5MBbHqdSb
QcZA6x3eqkMeVJJunbLTtOEYtDa642KgDCUFRDi4IuOpR7TzCsQjp6fR84c1hWa8YXUM+03Hr3lS
D6RCmPc+/oCeF4Q4QMv3V8MV/H2OHFhoHH7xeh18UzFtkwQRl0QaAGdSkOZ9JaaOkMt9IJU6dErW
DMlJY+7BGEcC8+it1GnXvoBcadnCM54KSfVVJh9BVKQ1x2b7g3nhDYBPv8qdCulqCkG7a7US745x
WFLNHt/hgIicEnsV41ULl8caXDh++zh+gZYGO8513NMLHGdCfN0rgNMuFBa7veG9gH5291JGzUO/
xflRKHX3IemCGZ97w0/zsVxiT7BrW/aGqLbIKk9WoRHgHOmzRBbCctMw7AbNkhKXit9jling1WCS
fDijNs9Bjpr5vSS2tIBfhq5QHz8QGnW+Pd21o3AI7dNvCFlcGvgCkPw5e3/1jJktfWjbV3v1zqKF
9qa0MXF1fqE2PIZaOAF7qxQq9bNYiIORw5fqViq28W9Cwhu1OK3MnBreuJX4AHnGWFHANNCZwwwT
F1xgNOyrvrrr4oHsXz4dYJ8KAkCrFGBPfd5n41I7iIXDcdTOqDEWMUCx+2RIh/2+2GyFDHgl92hx
EW15s5SdWFH5T5vjrr82Vl33n902FTpi3wLGQpsYjn41sCbk+i9bNub8QbXIrLl6J/VwcEvcrehr
POmvaF2LWwjdo+xDw1rLpgb8fD/xZ3d4Cbab8qVbtppHm2RDcO/vEFhu7MTdI529TGgdzNt18ABI
sGYgTc/iFP5h1BhhfglRecqKlhDSFaFtYIqw3F10yV5RCaZw7vjRfth33lO8XreA4HVi9az4u9TD
tU/9b2JcZD6+kOGF7hPXvI0GKm1W9yLInWYvSRd5qu8owZ3AOJAjIZvz9Z9Q9sBpdjeP7o8rlsW+
Z9opJWfy8TcPFa2C60vY2DuiQt2/rT9+jODVQcZ8hD87infPPcLQsz9YpsjYJOYP8nlu/7WNu5o6
6bgcNdzrpklh6F0YlFioZzKyNeRQWtmy5chhSJRPV0X/B6vO9bAhb59ClK1tv3252VShpU8NDhV/
W1GHZDf+VfPoRMQp870gRZS0MhK4MdGMdRsufA0jQgiAztDomkLKfQo4qVrswEKfzVvvvwDo+ytN
YQ7X088iuzVd7w97580ChmDgPr4R6VdCppCUrpFura5djZ23CRbUK5/KA7IZzXWxQfX7qQXVlAVZ
CaKRn5HkaeqvBH38mwYiixNL28/CwzIPN0DD/c65BAzG1eED3l6QEmDU5t3+vsIqtLANYMXgpKoy
EzCQ4olayXQw7gbMexEWCZDP+P8ir22S0VjOQUMcx4sqGx9j/mh1RB4m3pn6669B25JXgjbWxNA3
tKrpDrL+HBxsPaw2it2NKc3vq+/Gh8lA1mUVFgYKoPb+9vRddvvsuoBt5ZwkYs4+EX3/AlXnaY55
p6FyNNFkEZPVPQhU1dRy2demrZTXLg7C4szaNZiS8yQmbUccyHGfCu+wGjC2Lqe288RNpX9RkAv1
NpE11k/NKHqBYKjjAhc4Mr0UEr1MpGqJTuWKG3agdRUymW4TAPgw3MY4qD8GbgvcIAGvB6fMFv/G
2v/Ji5sQYR5iLhGs4oAzbMkpYi6A1Zv+q7dd+uqKVctQpgNBugR1mqlncxuQvB7ZT4CrnrsCMFI+
H0AZWCvNmyQPtkHVKLMCBewPfCW1tL4yaFOGrUPshc9B40yVGlcKsmCsoGRMbqx94bYsUPOJC2Pv
N+KN1H+cVoxE/6fLoZtUQ3LjTP0qnxYUpIfsVFWIY/3bk0POwPsLgLnmvytQi83phBYHVDbHkXRQ
zNiVl5sCvmMsF6Vtb7sT+TVvmTLRF9hbe7Pp4h3Kq1VGCo6zj32jyXswr3HU/fsZUHce2fFrMQJ0
CeVpV3f9YQDtuoEO+lJOoONwV8EZYi4tjDLx0YRmVxzed/WQuH9pappZhfcGDlGYHSR90QP3pWBD
HJ8GnUzkXs8ZAy690BBDyUxVoUq8fXBuHUIjQBcDQ92uxPp30fY2bSajCc8w7h8kk89HDLIWQKqA
CEl7yB4SPhab3H96oUipssgImPbLDq0GvoTM+N2Oh9bosQ2SdqfNrmYji8OR9/hr5GFEELr0cHAE
sO/GE+nkwsoeUDjOhXGbE4xPL85IB5BhQp9396jwqSZVnM3tZWzTVGHFu6a0TnAA5aGFe9NbiQJa
gphPRUaNROAK7hf4+tvU6w11YBeuqnQFEXeTd4RDhsKoWxEUcSYrft2qRzSousS1tkmAi3Ib5jCU
xJdIycR1McxyT94Mp6aoEIG1taSeGZSGTPQXAMC+jolUQObFrmWYNCr4XFo65wu8gWfaLqOX9teZ
w4gXHZ3F8acY/9OdntwItSUlJ/2SUdfZc7QJ5up6VSKHYqy+HRCslTDY3n8o6AuV7qBnxJqTZcNl
oM/gKtOB7WuRE/veZvKGOansFyHbv1RXyk2tqEgbNItZo8C7RBstt7Oi39HM2l+kdhTHGggFA8oQ
a+WtU4g44gdgdq/tqiP26XDHu52SHdc8d7d719l9X4kGmuElN5P5nZKDhDeQBXBb0PiiXm0cenVH
6gbZxq3WI5pMKKEwbi4sD+KbSr0hMm02R9TR6tpQFT+nUJzEYtKSvq3E7Y8/gnehqLTiq+z5IIt6
KWZSYD6wQlyckg6yOjhssKTi6P+ov+02Ic3J0ScW3KPfPZrnUDwJR3O/cJiEdN/9dv8vYr0sANap
/G/guL1F2YaJLYGjnX3wxGpTM6uzH9OKkzM1W50PwcSDXzevFyDOVUMo+EXmf4lSFYrCAO4JCVFQ
VjpTBpiexmMujHJo1BeXm5rZP5ufXY2oMyif09Wu1Sg3s5gPgQUFne3GbtF+J3onH/atZs3RVxDj
qFYNyObeIAhz6UT6zvtuCYBbqhO0v6K1ycjVE0pCjPdexeVaJjsPWlgUd3GdySOqdAWGdjo/9NCK
qgIKWNuq3pVY//gK4mzQPF4ITRVfY45v7dCq+mQDMzl5mnOBJJZdepnqdNe1yH5njl7NHwO75Keh
/G45m1/6rLKginSuD7jdjhfWwHyw/s8dA0c5pAYyegRQRtLPM2nr5UCJhs4YLU6TtxLLfBSHYK9G
Rtx2EXU6wr8DhsTjEfRM/EGop+KdTqLMG/qIQeXmNkOWFIO2sUxJIwRuC5DlEbKZeXxz2ukpNzYV
l+9PDjvzBH0spCPdNCiRKuCC4rQvxWxFzw3u9h0oxlzuRXu/lurRR4DuUtfCtvDmh9yB9tiVL+pg
Rp3JgWQAi54a8bSzLZ3jATnnmN5ngWUwopfvh0BIXBGMUMv8DXYXGxB7yl+xRDVChYdSUQdD+vRu
iPA8p2icKNKRe4JkrvwYKH57nrP1reozjr+5D3SNgT1AmXgHNFi3JV7E50mjeJ02kyRU/zythyjn
qqkd+sL/4iLCT6/cH6Qi+bR0Yi5OTp4JTHGHLzOG0G5M/+aiKiXXYdsjoOBZAJn3bERYwfWUaHVH
UBnRdRQqSRuOwV2NURAIrbngUeygTE0kTNqh52AJwGTetISZMKsgNMVKJQamAgaVlnmNkaWRbQaN
sqy9Gydii3i25R+VnoSu8T+mRh1iDkgeE35Fxr/PX/CN9xU+6ZV7mepky2X5vh+FZgpbqfwCNoFS
6JSJ5B1lRjks6o/O230HB+aQRYGWI1D55NVhXi7bThH31GoW+Aqb1kRnVl0lyibTuHvUATAuMWBj
iSXdGvWKJxYu0Ttd957SAidwWVUJoFWJzq3mL8GtyJZquy3SicCkQInq+PnZbWBrTMBvgxxNsGdr
9QJvtr9CAiEdDxRuE7b4Thtpti2CK+NCzZvAy8f/7CWVwrT7qWvYHfPu3fKYY3wOens5/kunDgUB
glZliEos2G0jRJsg5y4jv2xHAeC0HBviJUvCK/PsYj0U/XlgFborJ31OS4dG8uKSnPTP+9kP0UGs
0sm8OerMp19J27H0AoZuIMwQyAnWGuBl8RNY/L/x31SuyyYiK5781ACjSBMp/y8NIwx0MCiyLPL6
bvSVNhFFc7FzFAdAhU12/+HQROsolhaSDv76Q4IUM3qcWx8dU39QOvgH2pC8bYtDjgE42D8D7Z+2
sP6UFlU/EcN9PzgXWhG0HpxUoFRGUyftxLi+x61eYp04s+r+Owkfs0sVwsq29WF6K5ryL1rjiFZp
ted+mVQbIMXG4R0X/L2OODmu+W2rqj186IMCckoX9Z2rZLPgJpWZ4IF7mOWDuFU/sZmWOykz5mW4
LZDys7Dl+u2kjqnbP+29IEwW+p7KuFEeIs9WPVHhUw6HdQluwfw7y2lV0f39GiBTbKo0KLDd3SZp
2U2/SxtbhTVLLGvHIbcIGWqPLfIwvGX3giWpzAt5hc+Eb8kWZEvfF2vpOdfOzYJfYFprOeVZpI/r
on9/5r6LwTO4mmnj/iYnIWelt/6cxGa7xJJnQHXAdWZfL0BWZ3KcRaHN1/87rtGD+fqY9sRDKbmO
rrntBwvBSftugGSWFUpPzsHYeGFHyKPP6OxbGK0Niq69+XERe+XR8z2QHVr4qXsSgBVnp3cpniYp
EL8GIAmgdebSqGjGelr5aaPR8sbvFwEIG980tyR9KakPcN8d3rnMj1q0KEO5YhOYVXwHVZN2ZDH6
FhdXItuPC+C5mF4u1728pYzGzViwjIsDRPyiQ+6X3Xo/EaHcwe8bldxjoN60FMPIddvsjVDT4ep1
9+C0NySDqtGr2TWH/WjYcF6L7BKZv2AVJVDc7u7qeKt0HtWX4LasRVUkEg2CggVdVhi/3hRLdkj9
/gSktULbxtoFbAwx0Tw24OmZGIM5K0hwjQEbaOKWiJ76fYapPh+eGo+dXQu8WlFJ9kxJ3m1q6tBG
xsZAvimqDuwS1jp2QWAsogPCTfLMtKAJGDTSqckJqzJ766I4UDtNQSNvPgylpB4jjZ7hQZumI4Kk
t9bP1j4+tHIrCegkrIfXQlEU8DLEshUjTHsDHjZnAJM5B7r4GmPqPQjyUxs3PagJ18QU1qzes7hZ
bQZXakSdZA0BlpethCjZfLrUNaORpOwblFK7BjOKsEvX8dHDMU+swga3HY0Bg642rd98VrCRfQjj
JiESKIuXwPKcMpOF8vbr0j6iTwIuKkhy9mjwvqCv9MSJUL9D2ba0LqiTOcAgQrmXYARVVmzb31hg
FnyCu7rznT23LKRVhMwZqBTltOHLFrYKDmNZbFkWaHKRJo2Ffh8icrsHalqjJ9MaOyWrcXT96SAG
HPkauUZkOBlU2Sq5Nw+E6bYqqmqBjFY5uzf9G/WziY6w8Pf/l+vgSKEQK6L1yWqKJSnowr+EJDi9
zzVCtYuJ4fGaIkNOJ+GwjJwHdEO3ZXZ62ab6+0+z4f0aVpSR+M2JybhI+o/9EQ+lH5WXA25FdJvm
xwOFlZGBkZU9bNA2+v7BCkS6g6q0054f0Pfn3sS1EIGAD7lPQuSXb0bWwfBo0B3jtTZF1OgwZAGi
VmAI6XltdZ/i2CiTclCpW/lL/rpSFmu4arWMfnqQTN4dxL4ZKjs457X8ARU/TQKHk/VGfYFvQ1ww
jfFAF4eC3r/QhP0Pa2JGKxwPIomIpdnxpU5csLXWcSZAILsuYB4+gGdMWALdDS335JxsdbcwKFiO
/byXeBRbv6fixhyNK+pRPfdnaSJKKXbMQvlm615+rGz83a+omKVd0CxzatiMOWVw3OpB8MNjDkUL
Jwu/4mcBwFLUYdBhFIEpVoWBJtwXVMlYC+eV/93DeNPIfDWo0O72f0a/1HGsgdgOZyyvxAvaCK6v
BsjWXA4g/4Lygn27CcanfsvmuXsQriOB0x23WAOrLtj3/CzzpMUeOB5ORsZOVpN72xcp90yua4Ag
pfiZqMa5zmBDeMmJdRxtI0KUGgVkYUEBoiyGOUqiHc0VEde5iNL0O+5K+x6EY6JRG2w/z/Qq82VZ
Z7fKBNO3aeu0ilMxcz2x7xQQItDR0o/n9s1CJgnoEn1v7sh2qW5Hv/qT7eDiaQOcOhsh0JK0V0Ts
HXbOdjxVNetxPxL9w3BOaaSz3zklFK9KK7ZkTqZ62+E3vAqGmaQSJ4YjaRCAMV1rVzbddtWgtW9q
btvXkWtExOgoGHEX4y7wiUaWDlFdpkDEuhQxcXCsDTZRjE7zg9UG3DJ/0Kf4s4dzDRwqL3KNJb80
7G7hyFNEAOKSywSq1jszG46KJg8Nk8oiom/hphpUtCo4XY584guch5i75K+AfsVNwWLycbNZjKYJ
z+7njirnpKMlVfzHq44yLZXSHj6UE981HyTFanj+ub/+G5+BTfWpevm54HL4hpiUzG6i6kt+lyvQ
x2ETmwdvrDcYTa9ulfwRZuqQmaH6ufTF+No/higQzkUAB4Das2fSvwp1fa35lIJ9FmWfGz5u9q3E
+ssnV8LZbZDpAFVHDC2QpiW3vxE46WSFkYBzd1PdM/T+9eMNXYV+gilkvEkzszHnEjdkwUk9ZVRt
+Z3k+GznQDS6BPjj3bjDwdnt+Sx3h5GLMhYA8mQtb6mOhR1vzpVPenZJ5sIRqd6bTzSXX7a7SwTE
DKyBdaGjwS+ZYP06V590sKQ11KIKwv9C4lKZz+J7+AZgno7SdZ8oHyazrxbNJ3FSrEDptd2b3Dmo
gYNRcHjyfaj9iGVdPKIL2HEt+PVV0ZKa8YU7IAInGrGLTwn734v0rCc7atAJWY9+//32NlafBInQ
Fypz8x1OVQU87u/MMhvx0k/MOOLa5rF89nfYyAtyGwB0H04gcjHQJY54xh8UKowY2pJCkV7NHt4W
9QFc/9CcnWnlSmf4IEUti6BmZAk2vkaKT6U1OrpRRFhiJWI98WEJQ2KrX03pTe9dcWBz35sO2WBJ
mUjhoZppwiaNqlTT9TZ1VUAoOVEmsskWIYR4F01kNrrIbzF5/KDmtDNJlYrkt/LV6JVfOZgRhPVR
yZursJnMpn5bb8Sce5Jotksf0mRemqfokQMhdZTv8/jh/DfKBUQ7m/MDa+OHEXRMzGAevcMK0WO6
bGcedmVwwnk1Wure68fGf/R0FGBKnNjSXxra6NNimbKpyu6oIeH95t9qs/YFaMGh1hrD2Jecn15T
Wlyq89FSajISFcAcVoFumerqHy7nNRZaj/EpIV7ZXq/AcVdIYJ0rj6zdepG7gl0FR60z8+Hf3Pc5
MTXaYSfn6+l5MF8GecyDGc1NUVnuim0w7VjvbxYk30Qy1PycFCuqmvXWNwZiIU/0dciXAxGfI0O/
X57Q7H84Vz+YFRj8812KMy3OP6Q5MsJSBLWgHdhCipBCCu6CY1Szs+9PLiW3oLYva2u0Iyyz5zaA
YyUzffmX/spbl9+C4NFfYLa88bSpD8fBr4ejvm/jqvddgXUPZSOQPNdQN50iS/+fdLoZq2IM9Bn0
olV4mip1jt3IR17jfKj2WBBS0oR0Rp4qp5nDydvJ+g8+2gK53Ln9Wrc+tCKGCrqmyDYPuBq4cYDH
hIjoC0mPC4WtCeTUBk5DCGxJWVpBjD7GseXESREWHJE0VP/7xal0Y4q5tKUHTrTZcORGdfbW6WvV
qwaI11BfhC8LxV2rsh3QgIkZEuvtMsRhWz82XgHTkplPOOE8qaIHWOPqvYSFkqqEDAuj0O87BTUx
zVdTS9TIdZVEH4Phkir3f1uLxqLDXcvy7v2LiYpHcRWfKkfEcUgRwim5LyqOoWeIQn7F5INSXst1
FXSNazkE3FiVLk3fEYkl/3mHFiNSBNdfn5F9jKD++dmk7WkhyRTZ7oVKV4n9hXU6cSoZnZQPJHlF
J/2EZMMVJyjiB+tyLSW7WA1RKAfddDa7gq/RaEr3Ej6e8xet1iuzw7N8erruNByDZLitjF4i+FIu
mF9mmpqiBKbe3V4WeGOH0z6S1mrHJ+g3LlaoLAKgF0DOK8wAxlppvHF8dVIFNMO2XbLQwW4Ea8IR
6KkDNoZlX8LxE1yqv0mm+M8TORPDRBAGkoMdDQU9p5Py72rhVibjV49By9MSpK7I+CpUp7gPNPfl
4fPt0n2b3Xxu1Bfv+iBvv9sRz92K5xx/5oeVHmclwprIyjWDpbqxRON7bwrBdj4yuSXVjMShbm8Q
LA0vVSkmotFu5+VC+q9+x6uhSuM1G//IBBK84pFcg4mnguqFAwzE85qoWt923gsD+HMtt4223stJ
ebgnFMbJN1dhmTDfRAq775M2q+aAZOqzvieJDHPcMrjgJZnoNWiTfqHyF8Bo+G14DvmiBdvDPl+M
T6QVnoJuWCIxpxMaCIZmEUBWAhyk+tjtH+m/DYMl+vMJ/qvtLGiod9WbT1FSHC18L3GeD2R13skg
XkKQz2WIOtw3xQfVro7+AXhKguBpmYCderIoRb7jcYTcUcuk26ZACtxS+cwe0F/cZLxw8veOMDZJ
l4ipukQYonh5AE9eXfUU/zUJh13sD5NFM3MfZFSXAb9i0pLvZfstxhUULZ00bxqs3ijPpHNCuD98
bsPJTOpGop0vskJdoyF7A8cLp+cVfUqqXE1Lw4q21gc97wseQWgrxoQqZyGFiHKIDBuxNUZev3Vj
oGB33U2CPHYm4tvwmV5EnX9Gdaa+sTAqelyi3/9113/F8+wrH0ALLYu2l//C9bIlXrNE/zKFUJ6w
AJNyhlU6/PP5h5lANZiEQJjTN0aWE6GmX7LjsX/lILry9T79QyxiHKd33Ol5PQCy2cZ6xAdv6G+B
grSC/MEtBlxiF3ImwxCPHSOj2QAKPpbzpXJUMaGz9maqRke/D5d27ymYYNMpaw1GHGPcdJqfZCZN
PMMXud+pcTxQTgq4e66QtV3Ni30L4rez0ng+FG4/dKOv0x7wbvg16sd1WYzk6mLXBp5C5W2tICiv
RlEo9B5fJzmpiDZhRrNTz/ZmqC1hB9uVL+5R94BkDk3M83BwJ2RcgobtpTkORFrHEi5wKAZV+QJs
j4Klemly82djWz5GdBKOtIG0R+/0rdlm/1p0uR6KxjJEuKsrG9rtmg4gMZI32a+RrhC9QuzdFARe
Gx/MofCMNnu63mRqPlDLLe63e4PgIRnkb1GDMb3Yn8WFXpCzDIW/CacI190LMemUw5GePRVpRi1X
CmGJaxI8zbBC0DvsUEP3ljprp8Yts2u/AbNrjWJ+CgPDlLQAp3qRTf0Gk+y+6W3lFmWhB5VSHwLr
uOiAn5QCnfv268igxBpwDXPnewVFYQsvcD1lAZ2pwV6R8QV222PsDWFMPRqFzU8yWNsFW5Ouzv1u
VMWfERRgd8embWcXbECZzvcqK3oNRnmtjKbaF6/2NpX++xxfROx2OqWXIMUqkUektlQMxdlFrr1R
m6sG31wVF2950Iv9evaDGeXpxjZZvyq6W0h7SHawsQJYdtmAaRdS6yGzi6cARWTfPLDDuqfg5VvX
S9od1jdXP9JEAmntv5JWWwBuj2rYvUMKYcEeZV2dFItKZozQUueMOlg5/ycUwkmD6vTOnRGpSPrh
oukrLzrpY5aptx9oj53HfMjjesHR2nWyt45BdWmFRv9reFMZ4p5FC19k5i8FR8VKWXUbeRVlvjjY
KK8dEPqNmVq4+SDXWK/GU55HwuqZOJHX+xJ4YFKCh9OnJylAxpw7iFKC6XiIcbEpEydSo1xeit3M
Gbl86GKQpyoryJ5T5aXLO3zOIjpU8wYsE7hx565vdnfrEVpGqzb0RzUdmzCycCpTn0FWzFWFvu4l
4UGEurKrL47eJthuwY2VGOaYEHybk+yFbpIBujnMSVkjqldepCukvOUjxoVK+WcNP4SQyjVsAd4/
KBmtCh94VylSmVVfZs8CEtd3UbqT25XDDT5MMfL8AcJ1sAR+ik483Rcjbf2oB+QP/Jd3MQdiyyC6
OzXkgVP/x5khMNWJuRPXiVYqIK+uunDT8vwHhqouEf+erFEF6nRhZ+YHG+hm4ug0eeHYDnHNzs06
+NFnsgeNcOl78HlkTTWsFudmbETJxGpr3jwxd3rUObjvRwzS60OjqqgGBglTsg+cW3Yh4xpZ1d6F
NzgLu0Lzr1i7tUoHblaDA0wzGZCZSwb5Sd5lBNgpjYP8eMp1Ul9XH4WOsiABA0/KymN3MDLrxjpv
wXMn5cU/+EdHidaCkNerRqNkndJ7LXk11QR34bHfRZ3SgREXsaZ9zama0LMweaaqj4wCD+l5ONtI
upr1ojm18ZSO648rGZ2tUmqFLAIfs2R44FEWUgsDOqehe2nIqIQ/BsYbgOovk+FwJMDFHuFm3WNt
axjTpZ/6KgacK+FR1pnUwLPMawA0+DCl6uC6WFQ8T0rN3SGSiUUcezLQdLwuwZ0Tl0/apRVqvBJ1
z4NO/0KTSGUQfQEgOEKd7yjm3tnGP0QkRltzwDnD/Arpv+ranE1DSRVklQRsnAAGVX3sPscBhgO/
YdqbuzpdYWfqwh2aBQZd3y6bDe9WFRQSkjhc0xne1EA6/C1YL5sBhRlx91iszkrnraXALV9IVI16
OVN/5pZvWGGelqlQZR68on8lpL30Ops1X7VLVFl6Z7RADEgRztqUJFDM4R1Wj14Ttc/HChQYkwfO
7FELF0BLIOywevluWLy+yPw4ROKDfQtFY+lq6UlIGCUGROpd9ai9R30Eh6KyOcZlN5FB4hTuLGUC
jL3igU8zjNZUGLW7qny6U2oqMAr1ycjdpoX2NOrpcEVTc8B30Ti/bNfCakNOR4VHApVhuZdg9vLn
NemVPv8VwKMj4JAnIL3ejfCRzVYMU0/g077AdeadWbA5aIZiWnNlo5f8CI+fIfUZpGnFTlk0aEVE
OHjMyt9JZ7R3JpUx7kxMiHICcyTRjMKsV40fYO/qyVm2hh1XV6Cr/u9iJQFv445gvM58RBbQQtY6
bWAkGszCITaYFiWZ0BqtRK0ftWoaXX/vK1/dBv/jY8Rebc0FVlHiGa1MzMW0HO3ReYUC53tL/zzx
lI9UpvB8OAH2BiKpQw6N39vXke5QqH3xknk7f1W9+2M6lfozQgi4ewCEL4bPTr+rs71ALKZDe4Qm
F55X2cF4Ht88r14riRURp07fSS108etqQKUPEDfU5gJ8HS/UkPwmR4zLQ5KQRZMTE7Q1YlLVOXny
dZK5RiAuhgjuvpkJogXzfW2nBV4qLHG/pqo/rF5uBRJ9jn+hIstu8CGnlADVxy8xtoIUvAqCB2H1
PVVvfmyC087GmIf6DStOVKDNY/OQk4z3Qd3gcavb5jYXYP1EJ7RM/Od/OvdBlgULjUsWgetyABsW
yddQMZdoh5FM9coOy3JHRJZG8aydFAoSEjOYPRVSCTzV64In24S6C7aBL9eUclg7Yxa8FPKMJ36U
fM5bGLtyZwhxaklWRASmCjkgW3BhHzOfDo7lhsK1HeZQ8g5+G0tYrAMgAGqaotNWRGcXBwxbRy3U
UcgAwbKWYzQyhv/Dj5GGFNw1OWbpF75DqlSFPH8Wfz6L3BiXfuICJZX65tx6Kt3nK+EvcsyzdFAg
YxcnCwJbGWIHkUsPxA4LkuxFVWrpxEyINZ7YJJwvnaRmTAU5vScLOJZfBNu0IIzJuE0DVxaFXKKi
TQHCc2gdv9HT5H/aaL6hnBywgfbCUzcRGwVfKp+bJxJokmXBy2iONjCq2gq9PcLADh/jzWVTwAMY
9Sv5TPm9m7fhcqRAbE2AoLGpq9B1eIWhLQzzQ2QtNrXSdy940nOMW1BGx/qANk5GR9ruN2Y7UuUX
Kj0RIa8JWgqheG1RG1xm4VlvSbynnvTBQl12gM+KHcK90+mthE+UawhWI4SzAGNEJ87jNoEMO7ks
OFRUQ5WA/OMS7l1sKRYU7LGNfve5QIpTIgUJaQ03n5dBFkEr3KkoYvNa8I8ibsK4Mvof1kI16/VP
pVt40vayfzDVqgWBvCTnvw3PVeSSP+go+XNnqVhd+OKh+jB1cN71j4K7mrLCq1fs0PhVA+ZEqk8R
rmImAhb81qoGEpemZR2b3QDGtUZiBKs5LzqAdHbyF+bEkapdp4sArbZ2Zp9oypTOCp9ATBrMD0J2
hEIcsnK8/jUFf7kWSCacR0KLtOIOw3CKN5aCx6z7FYZHfYGDiRPc5e1OlsnG0pAGElaAQaZUBLcy
d5FlsIb8r8R/pt8arxoibyYK3qBfKMob3LspqcGYg4kq/mRlIjKbzVBF8zE+dIJJVCqWE23Xul6Y
0+NLTTMW9rHdL3RyAnJjWtMh8winhcsj+L0YaQT53UKFs2+R/go1X0uzkh05nwOcHl69WtogkDMc
bjdEZnEqjt0GS7f62pt5HE7MqNX4G2ePeFB/b1z3/XPJxa5VzJGKdzqfKuKA7FwWixISGMqMT4UD
4HEGnnn7q53Y1j+jZeoS/lRqz1neV5SoK6Uw+oLHycmYfl6pSVGWfd8l4IIJSZyn5gb5JLadPwFV
58NYyAXlOe63gEP4NvpuXyavQ/SfUPAWy77WTjePslDTT8vIaYAmCMESFu1pPKnYjO8LGFQpLb5o
GXEGGXfnNMYUMpuWwzEMjzw4akOdTEnywhB02wralMv/dl4sHSA/SsvwyD2HMt569+XXwmS3QSkS
3BBKoZnUX3RnXJ1cP3h/yOIREUcY4G53U3xjIXN1I6hjroS6Vki6lzKGKiUvUt0ARwPtROyd4DLU
gNaP29GeXHnooMZrJvujZTmskWNvz7F0dwgGU+jcG3CLDtrSWmheevadbx6KQX30UesH+V63yXR7
eFg4kGhr6aVqxgUIHkAkMfZiEDiSgMSE1WO3s0jyYh+zSCSScR1PcT5c+OtWVYxzpQj1blPbAxmG
5oR1NPsMN7Put2OzrO9x6n9GUfMSFdxHswDkiLtYphQBCR38PrUaLTMlZXEs0gYoKx3vj9OIZ/om
J8EU6GXJ6+XGL6RqgXpmlJ7gDt95EYhveMi1q+GqNcTtbf9maVadheOWBV6V8o4ncaxJFRMENPqt
na55c2m7aM/9UQb504PGtxItHCL3jY7VOQP8qDGGUTUKKU3kVK4kOge1sUvyUIgSIZdpIV02scYG
oxJHcKrDpF1ab//33dQgPWr6na7rTsXl9+kBBxCf7d9hBaDgVKdVua7hMz7Zg9PPyzV7MHzNltPC
0CGFVFm8ILIsOUu62d2IHp22XswXzD6hvsSS2y91oDfQW34JtGWAc3L/VcqUZwhHgKYFCMHvEZKR
FLJsCGvfZSPB990i0h/XowXnsFq5n9xxtxCQ+zIMBlwbhh27nMBiih5jBiRGLDLewVw+1swfISXg
WqYgOHXj21qPvSQ8d6imfahm6cj+0s1Opn6HUmpkKoWw4r5I46fFL/1t9SC0XQtADJPm+BW5vJ8S
8dp1DpqA9aJUed4e/rkDsCaWGS7nwLs4QiJ8vIv7RbKXmcy3qrqOSF5csi9jC/qs41jV2gyTXTF/
e9jKxLnRiJxBbU54KTLu5ghfbqa8pChtD1puyGgl+ON8+XI3vQizk7Vad0s9O8ABTqf8kn8uwN5D
K1hnRli7n4dN1fWyRZZ29EzbkAxtrcfPuogIykWCMXDugMsD3mZt71G6zVcXJCe5Bd6kwsbDKcV9
I05izalggae8tGRlcQKDzKYjrReMs9oVhJOB/vNoNpLs1mSxfIf4Aqu4cZygkWYDrsZ3Woc87XrS
JXhY5PcO7M7fyxxRNCl3dGI2ts+nAEoUsS7fhp5PkSCBoeT9PGcm0TLQrxb0e5B+C1fq0b5qmm+X
idiZDXUuu0bJ3SFZbSGCBjr6Urv8clCZTQKeKjmXcXv4kFyKPgFgqdfa9/tWcL2WSl/8awt3OfKA
rlupa12/JQoB9qExZFLrtaVP9DtUVob2D7bEyfs5vwU5sZRh19pd0zT3jGOKtnH+NwhbmpgSNGHf
jSxsE3SBOTweykc87GGs+eTpxHt3MQSNelM1aXlc1T48G/s6pOxCdjRWe/RntEiINIrVdbgU1aNR
31EoOQeGG4AWiiLmt9zFXHkSJ+EGtFwr4jt7VdwJu4pZiPWoqETYwM6oivaONzFXgYlNxz1YrYoO
qRNE/wVbffIzoxZ12fBFXGMM5zGyPt3NJs3OdFR+EkjDij4cXpopi0HSrFP2BNoGziAIIk65ZIVm
nvK8INoeBQlOrzwHmpZaYZ9PmjHeK5RAFpZ7cGiUJ1H2JqPRPZhYi9XGwuJoPRg/uePohukzwXgx
8oe+B9jWX5PWXMHeU/ES+Z6rY6qRftaxt8b86hqFuyv+wUF8N27xRqedRa6QMA+RdNQ2Lnt5DeUZ
aH/Mgb1FHNJlGwgQ0goGcJw/e7yE6OF1zOHF8vBSfgvE50D9XteGY+cJ3Z8J9Lj7zjJOJ2xhs8xt
wT5Q5QAgMkMhAUeBJziAGKvAte2iuEdwaSCnKeC0mYyrSnnkSlFLjV68TAxc8YktVYzp/JTcUqE6
FyMSYZG+Lo6cDWcHsAjNhOLt8V7WcOEbWoY50yuC5yrp0C2t8IZVmUSCb7JWmxR15V8UBCnp0zXt
FpuaBt5XN1SsUrOy0tq8goaNp68v92rq78D4g6DILA31ZFkmT9V28k6FAUYAosKZJMBxW/oN2X7w
6WY18c+nHRS4dASl8oHOA3X9fhKDBrPBtsrozTB9jG8s47L8w2o88NDUdZRmqSaQtOCYxu4kSQXO
W9FefvOEaq4BowNBa+Q4Dl8JLaXXsIbqlRZ/JjIYBzjtfCecvWA5aFNJo2eNsLcjHv0SR5Ef3A3k
ezbno24NITiU3ZNKfSiDzdpPmMTH+gaov2WKwsAqm6OLi9TCw9S80uqoGsLAmW3wxayAw7LjRjTn
cq42FG4QOn/6qoAMymrfZVp0zEs7CfJhUwV9tpi91Li9jFBoRrE8iHIWRZZO1zDG1t9In4VKol8c
k1SSiZ7cVewIByudUvZgZGftPFpPTqZVcbBtqAMVu3sS3g7RgRGUVzNP3jYpNOB14vUDGPsutqyN
l9KNOgKukpri32weF+rRXR1rx9ERoQB5EJ3pQVe0la4pdyMcOkIzNoRkHvJ0UBlN0xVjRv6OTtjq
qUPYP1NhtqPbXfnqOkjUqqyO4Kq2zhgm/evL1tHPTRUqjNZrcgc/Q70a4lxiCCqp09RvFxyVsNQz
OHM77IrmqDthmEwmYFvcJinN9i4jQlRH8yZRCG08pWaMlj3oZ2rxGwskotOWUdkkkszkXV0G0ESL
9/oefkIB7aceb5G3Ng+kc5p+LRCkW8HHRmBepPlUbMfhrnlbPCGHS+2hs3/7ZbNoVB/s8DDbOQan
5p3EYtYMUzHPKxUQ5nyYMNTvX2gAGrQPZnbuAJdMKxgz4vsPItCsnKAzV9Mvfa7xlm7QG5Y1Z8vz
puEwG7hkwB0KLqiQ/1o/lWsy+NL580WYkoXRDfZNZGrtM/EUrKEngnxNVH5hvAGzXO8cvb+jmSwT
avmBuQ5mcgv5wF/lwzbtDhC9vU30YgxXnsjV+aBfY+DEwMyev9b5+2qer5wCA8JxcurbJyTXwq8+
asoo7DAAP3PMX3tUy+EkYdZgVlDN74uwdzt+XaaMmAN5xBd+9pz7aRjVhsxl7zUrv1KiVkvvSyb9
nKHoMn/qioWNPj0kPX4+QNrvz/xwIiX2MA8bvFWFPf7vGGSRThBraBPU2X2foGOeetuVmJj1d9A7
M1jum0OkyDcooFrEkt4U1OxraVzVfi11TflLZp1Ue11PrOlxa2jLFNvh4t6+aTXAFb40t7gGvYKD
ejauW+uiUTtoV2TR/Cot3c00QM4y3VgbOOuWIuFOBqSGWmXAvTJ+iHNeLfar82Rj/+vq6te+AHcG
sH5oTjLKjglwQcmCmaRIYrci40DYFIM3RT80+x+1ARgAAgZCxUl9I9WMjFRKO5xAV3sl+GTKH1ci
vdNhmxgWmJ+YurV7mb/olc5tZN2GNjDi3vU+HXLE/o9TCWM+K0TbLp8oL8Ohu3/2VRQr06ChkRLn
Fg6UHldJvpuAwJtzaz7yU0LvINtRClY7hRRyiylaWqh7EE0p5GddFrgsg2J4IiSO+U1B7nMCtOZm
9zoUkpZj4XIkunNjhs8614H05SBx62o8Q64D1Zssi4ESJEmSheFhSAVzo6GeVVBUdLkEu8MfKPsC
jo2W8Ltf5jEuCntjvG5lHvPj2XHr2FWULByRcZyjEodo2c8JZ0h/wVbl9dJ2BMfEgW7sThpwuen5
T0f9aXSdV81C0NX+Li1EbhWei0XkPTU1xaG5E+RfUt2tbA+Q3L/NrZikkl7ZBBFT39dRXHF+tSWD
sM9RpUL9+veUVGlftn1FurdSvsXlFyvtsjgBlOEtpickcYNa7KctiiSm1J1qZERCO3bgGOWiK4Vd
CDFmMKbKIS7WBpBggK2iEnIHkYMytd2CJUH9b+dpqhwuaSXWxQVYku6qm0eqWe60KNphqv7yxKSh
bczo7aribweO4SQFCJPFjMCgh/xQ4aOui6i1vYTT5+ewNxZIbRzI1kUrOQ07vmSBQ9kjFLVzENNI
Bza+iUbufq8rPDP4kL6qT9TDwc+DUDW8mh+am6BCCv1sTqlV+GNrRjPllMBX8R5WCKVB+qZegn6r
W/RqgEt5g+jAlTK3luVRcMDjZfYzwLpmgGbXD9wwL6PqoCDcrNGCh+ik1fnmWr9XNElQBnX2NA51
k6P8JUlpYJ2v7wj8jORiUCgnjGzEv7bT5c7inWMt9ALlOfk8yXK0d9/+WuPZ/viw89IqHY4jubk5
+PO0HVyVKVJiw1NC1RWdluj36ouyC05COiRBXpauXn9H/gcfSdSYm9wzbEiM/7pICNa1K9brqUto
T4XPKbHS5fD0SWeQnxX9oDroB5KpzWpcDwW2LsuwYvn/p5nZUvz/mEVP+ysWE97KoVe/kdXj2Pmg
eWaTqA7TvY0Z1OR3eCJdXrbUhTmwDatYR888z+v1thXuCX9tWK8iMUF1quqBakkzLPvBqe9Cno4d
VQka3Lme4hfqiHIEedSufEhy79II+QQAcbmSmbI3ht/GLKrkAHi98/jMP2OGmQqm3wPbbFsA59mp
LHzNXDrRjx3pKAVgHuil50iGZrDbezz5YTVpO86uW1wh9JwUnCcbSWbctiKFzG0tnNWoR6EVTcfN
IQJm6nfcgSg35+BQOS7sp//Q+mPBbrtRT/V9tHBjtT44WOf2TVCWEyEYMku+kLooL8q60ZuNSuIb
bHjAhFrdNXoyBc7ShGX4RG2q/qdRemycfmqPayPEZ4o1DVG1HMuPngX/hTaTr9vKeMjbElFcTI6o
5OMbhcq1Wbh+B3u6ij9OIRENxAxgUAEIdQAUk0+fU7K2j/fxS6azQfZ7wGOggn032622DB9/rTfV
ezY1x/kmPCCurWqXtCZ42XjkkGJRAOSyeIh2EgsJ6sppl1inhWWz+QgFPEtlnDd/lb111/Nouxxu
eeJEtwKpoThgKoOxzhJaGjwjCicBDj/s3U7N0hhvEv6Jq3F8ioXfoBWowOFDNqqmPMkB4DGXHX5Q
tu55A0DNRtJDmm2q6qIUrAabVzmrMXrxb6sV0RpzRMDuVeGhiddL8gvQiqL9pcHxjd30hsWM+jhK
PQ791wqk9Os3hwnfsJJtBY1u0t1U3O3ChKFbbc9pgQwmiv+z4+RXUX81aTFZgDqBGAmR7HbpD5lt
lq6hH33KnEbI5eIlXWt/9nYF/P7Yaf3XuVz0i34/S4m/PUlzdUZpLSmevGYHBRoBRcDBKqSGaeLE
4h6Cz7loh0pEzWPWB3b4y83b8klFdD7KilsBd53WJcV6qlfxm1xNCLjMW3wp2WEJsbglFIWzY4Vy
sF/lVmM/C1I+y1pWzE9LA4dK0Q75bL8gQ97e9to7qzCe1x2vtpbhM8MLLb8ntkKBLlEmBbnJngyx
LkWFP1EEdX7GZ711K16e6CnqStHvcXyZb/1wafjq8y7BQflaUgUSXLGTQjOqjyEw3k5ex/IJLJYa
cWPYrsd8palkA9az9mWbiWoFZ4F7ZAOUlzAvr5xs52vAY39SWjrlnyZjHZTVfT8tVHt5ZUGK0u+y
XJz4P46DtP5mkr318J+r8gRAwwlSf+OlaklK7ryKntAPHKpTCm5IIbB08faT8ToKGrWyh4j/mTHz
0J4raYM1EogtkJC5MLUnxl020YWymO98GmTDSsILR+bPrVXmyRXAS3H3AhF9m3TYq2C/es+tj+Zb
+g+VWOelc+ryrhP/il7BsXepncVEplVMZEAyBFFOPfXIpz0LFQ9+Xthh0jCoDO//JylRE5bJBE8z
22AVFG0PqbPoQ97RCo0UlzcEejyn4/ZYJAIsav0Z/l2SciqqbQvtxz+KMkU9lJvSr9mRkilFzVVj
Hc2h0y9FGtEOyjWrIRjiS4+ZkoblkvD0ZZwGnIC6Tlh/NGIxnWie6sAxmsUsHUXJ0iPPY5PwjZzp
HzHSSJ20N+qdAAJqR9SrBpfq/n8KcNn7j/m1LMrJz0M8oP3HEHY7SjgpfHl+B/M9v4oQtFubrQSG
BR/VGAqutZI2Ou8dcSnteJpd0w/7mkeKtjpUJUqIN/RMjm2cCeGUm2Krs4okQzoHixx6HtFe10bT
8miZ+FvQQBJ+PzYNhebebNHFNtqo2amIIh5aoDv+ZHl1M+EBg/z9EgRvnAWDpmm4pSYWbZ0h0Al1
6TzZ1QMl7k+hK//KunOGjGgw7E+MDQ92WQIOO4hPt2UoHuQBlEWTyFOPnbQxkXnrX4OVy9EBBK6h
tLtCSejYEyzzvP0t5z4MzH2MmRueXNWD8PmVv4UCZHjE+ybkSwH/hMEz7c3WJPKhg+nVOWw+2nvi
N4Q25YRVX/si5CTqVEhtzg9nN3QnCwNFb9UGOfi3XK297qxG3bwR89roXA8B64UdeWCZP5RZsVwA
33rC23LQccwB2ISUnCWmmoPYeiRwk0C16f0cCjqYMet/uuZpFKeRJ/PdZfz9550QhkIqziSfCrxh
6bedb+EzdbfqAcs6ppWZI21giGPyFq4ZPxBQoXtoFF/52PJQdkxr8oP7vSHdX27tZ1kY8rseuE2Y
TmIpu2Fv1HvKAuNM9hRzQUOL8YovmZ9lhiAmUrgo0z0XSDviAmyPHGwgMgQ5NSxqB7q4eHyImdCV
HvKgO+ysq/NALuusUGykcpYiMGEtM1bPn/4+1ov6O3EjGjkpC4GlyI846dqA7BF53eSRyDXTP0GQ
YOtyguUrnsrRL/SguvcIB7qxvrdrhRjtJOqMJ3HtIiYO7k8LK0T57vr/JkuIzS5Jl7NU91esi12B
OmLPVkGqta7pTYT5LAS/IOn4ASoyZF6G71CRd96us0kPsmIpTBIjbbTWf40BDDCM1bbTUWQkxrha
G/+YAheUYtV2pHfJdjUMxLt8tOV+/lJpLUxnBg3bP5Gz6CnoOSIUVQKg5nHgq56X0/nyvm1fkXxS
4RH6zFBFGB/TdmqIYEoLNca3vLNtx7/MWgLvdd/y9qE6zxPM1BgmuzwZXKBq6gXExAYcZAhZswU2
WsJYTAYHlZs4TlOTR7W9tZo+9kdhBX+2oKXbDVq9MI/tjJdzmxdwLIb+nG5aBHxyGHRh6p2rsag+
QliM373sEUZCiWBA//hxod2OslqnF/N4sarp7zDRmqkA6Y9jm+/eRhv9YW9601/1BV+Z6diI6DcF
+uk6rmclLPsErZyPeJ8bUaIllOLiVpMOFG7+9mvYyuptChiFMELFGYPmWCqIVkIBAIdVdyqYLMcE
VD6Zd4V0NNB7/nz8rAsqu8ZAH7NUt7QvVvvo9LDC8odgpFP/bcm49ml7BVJx1rMlLa+ggwxl+Mqs
5jENAo5gSG1pIN5hX0cfiwd6+8sZb6BZZw3TJ5F8hps5WxqnpeEid6GmOezcJwmS1wnUXIuVWtAz
DuTa9fvFqfGI1G3VMe4bU2vv4dBzMKKP4DHUdUVFKjYdYAXoypFP3jXr9/2e2IgES5GF4OBk44Z/
fPr4QuRxgkC29W3Pn+WsMeT1DYIGJ5INyhJL6ebke5l7lqvSVfin/BhI7BnT6m+qA0sJrid97gpz
UlFR8iAtVd1j2yBUnA5HXcKjPNo8zUdqrp9w3agGDHIki5t+soRwZ/Mrv2a5JZ4v55ON5Jk4y0ov
Gk2kihlu0Z0TJGHK//knUmVYL1UFAESpmBeFr38xFFynYRoeXY+oZywzWRk+BroKPlIrLuYBFcIC
SYid8TRYScX3iaduoiez6slK2w+EDq3o9yHVuvWCEtDxz0PntT0nkbwTwbSxmUxt0pJp9D+pkFbE
lJ1aQD90rMPvElX9lSHDIB+UXBRT0M74RTzmc59r18HRwiAYk5bf4kWYL4tDeg2QwqT5LF7W3q+c
oUsuSjcF5bbdidWQbDRpq+3guA1J18RbIfKd5JiAu/UkSXVntGwkKXd2L7COK6HrRsGmVmy8Vtqw
5IoNpNDlvo/rsL2hrsdTrIqhIuCRwc2GCjnVlEelEdNInw2fEZRSpc7UB+WpMjnCmAdUZShbvDqg
OWuTAD1twI6u108epULVxYy7HwYiygizBmcGyWCoMo7RDsrQAxanp2cHTJldKz1T5c6khoLrhahP
hQE/NC8HgwwhzUdCaoUU1YSFrEuGa7EHQkPjM4IFhdHJqTtbV/wZnGnHRIyDD3gT0CQAttrSTNRG
/hq54VeKXBzi08o1CXty8TVD2RX3RC1cfUqC7XTa8qe2y8tfT1XFrk0bMS5WZWsA3Q6WjPOAum0a
5GDy0lLYQhGaIDqX9sqv1WcawgUS5s5n96Ej4+FzDTp6RUrxrP9euyxUYROszenrCBlolT+Xy2cz
eY7mpoTATJbt1CFYNMulThL4HZNNaYGDoC+QtWi/9HZxPQDOI+tNbarJ3j83F7f3AMhwLqZPZ5IZ
qlDvj+EU4Taxd3nSe0A8QVBZoF3jVrp8fadsmMc2jxsL+NJTkrPQX+TP8tyYEh8TMk6ymbAg7te2
wNJimm6PMVmOyfyUGR/C+8ot9Nfs4einExpmprmoPKf008bcnyjL2BSqryyVoytf2kSl8tJBtWjX
1nEzRxyG83JBapxx91zk+aN1DVml7OleO02cz8ASZb613rJr3KAdr0hfXmd9Nkm8Qf19/8yn618P
aDVbT0uEvrIPaRRRTcvJ3CoCNVJkbdORAyZImmgbXk4NeGqSjOFSR1mJjTtSg7H7zkFYJJ2P6h8O
eI+ujoUqAycuZcbfW23lOT0TtdLSkrviY5Ajh0jlRg55bGgC3+iVJcctPD379llNkUcOW9c6oUzT
JZRTYF8ktHyIlcetEgk85w0gP/LTq2xmgNJRGIBg8TRAzxQbix0ynEOUIowjEyuFRajgen8tLA+Y
mnVC/qvuKMnqcyXEzfHrbr6aAkcly686ypf3hONrAa5nmP0edYOzk7mmqt5QAe+odTf5jUFk9RFA
wG4FDy3A/xu9QaE8RTuTGvQB1lvMjzTlP9GveqhztZUnI0ILnJY1Rsxk6TJHk0gYhVMIq7p9t/35
+LAkjaDGcCo8VZHesUqT2X7qegebxJRckyDjZmpmL/CvZxZ05Dw8XbGmzoPjbp9pimSp/dti/ijC
7+6KdODBi1oy7FVkYEfUMDlZ+CAO764mCclm5Y3ht/H1MN+DOEcSG6wR/+YlfMdkbiDddQVZdvCe
jWwQPWdtt0Kcgys8D1JwONJfTBsmWiNvb2EJr6JhMe8UV5eysGpR/1Z0sg9Fhx9C8QhP/qF3n/5b
Oa8lc5Ctn6HnGfpS2so729uhrQjCjDWEg90HojOOcvrvYyyP7/nY2RxACMkp1qYOzXAATjgWWjWz
nMMlVf+ae34x8KcmyyP0Rzmlj334Jo0QGCG6kQDlHIBx8Ihm+bDUJRU4GFOWG1xnxdrEz7DuPhjf
Iv0Rtv9+1OhYpgQXCXooOVaKGQ6j3zrvz4Zyle+8G461MvKadLHDcvAHb3f8zg04cCBBYG92arXV
rO5tTsLN5W/UEoACsuXO74riYjYLEU6vgAQdEPfuplAGo/He/40SzniXHoN4TLNsskFTTwn5LuGK
48wSvJjKSDs8IaRnP83Jf69FzmKVjO7MYG/U26El/DiGObKlhGrK0abcjQdUhDN807V6tio0mHf7
Ao7nIQ4AXq11AQFk53/VcggWWjTiqMgGiki6iyW8ybCCgi0ac9evh0cN7+gd4EjhuahL6eOoUiGn
Q8zdRaoxWQuhtksmYLjWYMtXq3v/NZPmG8oZ4YONiAKofwrGWfqP/f6ofg8accMYoT0H+VfccYYm
1oIVV3DToJAr6mkHHx0BlRdufs7nMYpGAbSwqXokJOa6Cf6RWLtn33PMplgaEoKCkeyzsA/qGCdX
mUEdwww99dpTCwNjiaQgdBL+vbGOQO/K9dEIIZVTrwUpeqKhctorp1B4+LOdCDg5ntzxoWICj0Sp
YD9Dybnt1zWaONHGXWoPaIEiVD9lG6yqNsxaoK5GLsvUxA0vEcrtNafSWKBnkxH1P4HV6+nmL/FU
oALfkQd801YXwbwIPw4j317Tsksq+s9OltaNYvcuoas/5xWvMD6vysPUWEZkofuiOOg+huQhdLeH
GrbHQDSjInJfHVdQdFplFzg4fIjwmbrwzA8VzUljUlcJN9VAxSx50fsqH9cett9+p6Tag0Lt9vgd
j/pfoD1c9CE4DAhjP3Yq6r6MxCezPcdiYymR8MZ7Wl1qgzuEKuDj1Uo5HGgLwF4t0ZTHyohrjOYz
SNav1F6g+aL2VEpSHkwgu1cNkfy6gMToB5rQ+KazefP8PCmwdsgBJ6kbfMRsr5n640FBlnZ/MS+l
gsnXX9M1xDUub3SFO1AMMXTVBikavMHcZIbXjg/8zXc8MOAn3yI0G/UcERZFjy7mgyrY5KB7BhEC
pHqpaE6vKgUAjzD4jkRpLXJNoOUTERQc+a06aFDckU0ueJcmpjZYYhm5x69KrL7oM6YHUKG2KQtW
FLUcMcO4M6Jjv7PTxDHwKarVt/I87tY5FzfbLDcUMPu6w9ODeQND9OelceJLpVF3pU74MbVLjTGp
en1/1dPRP024ApeEsuLt/lZdi6CdVsZiEC2mvSQwZQtok2uN7K3AaJlBrAzVg57PxH4y0onPY8Zp
FgNcNrm8K3jrjjGPIzER8fKqQj9mC7Pwm0+/JLYH7P7Oe8kxk24dT0YYXL8n6H45Ms9SkWAaQdT6
Dvlw4Q05YsW7o5Jbv8k/0Ssfu1blG+Sv3rie9B3Ytzni6Vbqo7UFMnsjc06iJU+VQ2bZWqczP+Gj
07Kh8WDZOFf4mjpkoHEjn4rn6Ydm/ER0KZc7mogY2xU7ks4qNVU0avq7x9L3/LVb3K3Yw5U0ULNB
sJtpiLGpFcc1oij+l8IYzGHKfy/+fc2CtpjDWHtBGrjEuN9SUX0dOp4agJ8g3wxZ22puRAkuY1DV
xALzcyHDvIOLdtC4HTmSSkURzeSCk4hvth8SEkKUaEEDjarFDUt/fM7P12/Ak8k8jdJDUVVb7kah
98rYVS3q+hr8vtALWPf7+37eonuR0XaQjqIwHvCZxUkgQP2tLr0Za9My2QuV5/dVHXF6qjl7BC70
ZjeXZYK5BvZLHkTknf7Z3ynanDSkmPz1skwcvdjBbUxxM71LwsLoiThEl+yu6VuLR2cInFUCLpwQ
Pge6DbceRG5C5SR7XvcP8igMFOA0P+CymVMorUA9GYzCPZ7wRnrkSch8phenyyPAV7o2QlSbFXM9
Cmn9Hpb5ymfEndX+0lbcbMzOuHrK/v7ZVPAWE8GIUGaXhMmT6TXrGGClWFnDYyfoe1CadITSKS3E
BJhct9RupknpjZQCoNmtzrd2vYWojZnaAud3dScteECSH5DnDxrPWOfF7n0uQXPdjhSJaqnB+Kk9
Qxc2o0GNr2HyNbj8+G/goGOJByNV3R84gcjNcpsgtzegPKcOuYfj5gRo6qNXsPnU9QGMujD4jywj
qyLw/k1v6spv7nsx+fQCWGDcV9NbmNVDii8OqO7iG/pf0fX5pgtQSIG7u2KiX2JoCl9ERsOcL99n
cyUkZA6OtHcFJJT33lrsft7cSAPbSw8Lk/MZV7BfhpTU7LVjsqWElirZkpFXGJaTIem7AKMPvomO
32O4//OTXqVHC+/cqZnEap3gKNj9howpnbC6VTjukPLfwETTUU6iDrNgGbIQQwIf53RJ8gj9H6KJ
dmxuUHfHJkkh427XKMKDEp8GJh0g2+50mMIL6nySN55Yv3bXkxOseRSC6Vwa5AXmnU7HQTGHVNvG
OvvAhUmL9ecQ9WEt/UJBTqbwdjv55VcM7m6fMxzvByO2zJxltmbOLAYyrydO8h4sj2mZSiiWvozj
gNPhGM3GFPWwV99V9gT6yHY8xXN+lUwy165pa2VGTFCPNUaGfKhS+7cOsBLIYKU8ogv83q6b7J1X
eO2dC18Uw8oBi2HYJU7ppkPJucw8JKTzMSZrJPEO/ee99wgbOUTkJtoONv1rNfjYvtuBnzZJwobZ
qzgg6tk4Woa+6nptEWpmmdpeGdeKoKL2bVcNg0LYm+MEOpmNlO57Qj22cpf44EJoPRDUD7VEJZcc
qr8135WRl0Go2CpsvfdbfG2IVgZzDeUuygvEEhv6znxo59SBIq9lSvtvJ19hLttjahgixgaxvQ6U
6/l2hFlt/56Ah7feVt+30x7HWU+xQjxaHf/h50AihVrd7oM5w0DHs05JRjYCUZdAMh1xAECfqSy8
tmIKS5bH2+1Al3wbOTYoTP1tGKfjWVWoPQxqyww298+RpCSAuU8A6m7IMUPAoktlK8Mf2NRK/3kX
8AemHE7CiJ4o7QLVkbrXLB55nR9Pr2Hrgb7yKRUvEfU5eJkbjsXssuntqWcmD69q4VdFaSpvcC6x
LxVUB1CVxbdeIbCv2X5VB+uAg8zq8G/2u9pvdf0E1EhTgT4L11C01PZLZrFLJVxOmFGbPELc9wUZ
CTOQgHS0D8eXq/dBW71wQm02JTbpW1UU4//GWKSfVXWsCLiPB0YrP6agI2Z6nrmNTL6AK0AgouI+
K6Ks1dtXhPeo17wJuAepeAS27LkMgYjURjsgTqDNs4TPsjWQJJ3GtDKha/ispJW2jO1CKmMuWBpR
mHgwSB7GX3yvjaN2MqDu3iptolfTROvxGTS045+SeYV5iTvvhlkgbKbLF+fRg9HS+mWRIVgygmDZ
+7FOPacY3DpHcHNACrNNaTgw4nkc0PmQFqyIL3nLv6gNQdmv3R9bOGZbfCcNRNzFxzxENpfmHdog
WaH6/9BWBy4eOXBbTB6kYZkomsm8rd9BTOn2Yh1fAPktRuy71T478FJRUIoHcxS2GMh+hA98bed4
ZAuW9fy40Qzs+agriuDUaabPbuf+YDITNkD6W7u48Sfee3KSSy5pib4kd6qPtOVmXy9GqUCbXfB/
N9yjCDOtmjuew9TXkVQ35AeSQvX9wuaQxDhzSZ4xRfAqWPj1hS0ZEzxkptdqa3oPMm37jCeod+w6
FNRZkUZ51bi4wGT4TwUjPhg3a3zkjnv6e9VeJs01xafJvN6qJtzyEhEU28HvXYZZpy16HgdUfAnm
cYdnfFHdX2/n0jXJn6WKJIgmAFio0VyMFZY3gDeKBsa6fKPvtadCVxSVFBhPINzNPquZc/HtQX3R
WI/2gRZeKXfhR8ydi+W3Z98oiStidglyeS8YI7/JU6BFVKkJrf3HacvWSrEOB/6rhlLNCed4V+/t
iCaA/VJxyPwWNz3yORs84zCU1QCyuSaU/lAfp75GhckFSbs7BTFy2PIZeeu8b44eA0VNLyB90Qco
d8BldlFBDVM//aX8AedJO0VIgalQd2SJaRWVVXngitg9VrP0qEP/vm/sANbiKJhRGEYQpphG2Ior
Ze/Rt/DOO1wEhsewauveH7PwSXYzsnB5LGAd159EEOEImDwUpLkhufayJSWFBOGB7kwJU3ZDDzVS
XXfEFCHynWqi1G1OIG1sZC5dKvakkoKOi0vIkZbqUUNQZYnpuUXTDtNG4V1IKAtnv9Vmu1UR9+Ci
LXHrrUAHJx9G9iEcYaKPlZtrwqxjmh7yhhP7Ieb6uTwiAcCOJOEhv3bCtMdi2JjRO1Uc/vmH0qqK
ds5zyYYEzFmIhk2UcBvBmFF+WUVwaiAA4fOjnI493vsM4l0M66RPb8KHXsSXzcx3u3Iv1VRLj/vv
1WTUzkleX8XrkD+KBLrbcj+GIRKdnRq1C7nZ+8nigMFO0nUIJ+c4dZBcYb/OE8bXWBVErti3RzlZ
VZm5WgLpnQkJAI/DfNfzQ6jt/pKdBtaSLWkq6IYT877L5S/TJ+qxL2UCDRcwGCam5yHNSnqIAhUH
IQwLIBmVhWlANB4PccjDjqDa6c+eyp9IyMh85hPmiWqFdl4d6Oh+KFLiBu8/h6DZ8EeihG7yZ9t4
GQUvSblWOU0gZ2CVrXCqhVeb+qRuClqhC7H13VoRmZlXKa2cNYeUxKm41Temy0SQqxMKSI1O1UeE
Anr4J07gPmKbJI/l/3hdKa6DND3AliKopTYTGYW6FdfNBMVxuGPjS8Qrjf8Ky1x0aZd1rwvsLjLT
qcSOdQiuUnW/ja7RYSrspnFSmyExDvE0Op8Rc4iAotw+tTXOYBQCaSUZi+SgRaqvBrgenVQleaMy
EN+6nE2wRUIftQFF8Li0odkScUWlJwkQWeOAbcZSDigchGjTxr3pqn22yqU6DcKcRoHSUv+Pquej
4cr22L5s8Qq9Eptp3UjwcWAkOwWiqj1wXFh1iF8gldlXF86yLBhB5/3rXSlBAbuIyNOFg59z/xJi
30hv2INQxWyfBt9lw8asyyfKANRT9ottY3JjL/++Q/VxWpgtJjvzlP8veAB7zDYTyqPZjDTDuagW
WSsNdNllOLnE5p3Q2gi7ewafXczC2uOuqC6slQTkCsExzJ8HuncXWSIyDpU+rwGTRWv1TxiBpZJw
72cNxDEIMMPwV6xz0Uc5d29tnmmn4xw1inNof6sPj2pAHWeMLU4c0o6sWr8jOaqByn5pJJJsOLOG
5L2TrvSWYTfiT8Ylk6UjhSjYZkt2p1NL+/QEt1OKFVwCSQ/p4KdSxFAQV0buuHgAFW81oaLx+rTn
4RG1ijLyFFxrjss9KP0ZX2s16VE6V5KGifK1B/1FMFxuxzPE5Gk4FfeU0yErjWnw8+FACi3Yuu8s
lQh3rYCfgyHpFgz6M3gwUgQ9SGK57wJjJ/CjWsR5MBRei8B0EfvV6mlK0bExC5kFkLtXsiMSfU/P
sFAJvcG4nvac7zaWv5hPBPm3ma+1bn/bYOElPDJ/A0aF8DC0CxVPCyVQyuPlYdQwTDVTtiSGh3zF
oUXNBGa0D3E2ikXgN6UPAR9jRrJr4WZOapuANBrQc31FiB1sAKzel4OZn2h0TsbnjdfNAi8ILr+J
f/4pWp6vp2HbYuHrgdvs3L9myJKAHyCNCEcp5HJF+J/AHEuQBJROt15dQXFIsKMZ0RQ+cygMxXyE
jmmyRJ4KPgS7dnEzJZiFxjT6Q1axTKPxExvyAiKf9hYQApo6kSNMy6kHGiwpnZDKvgbaF+M6FDe3
aXibrr7pc7OH2tKR8/+m71YUsEAo04Yqk9+5vL2gp6Nkjk5pKHwKkJc+dsgapWW80/U9RxXYFquM
4VwwcrPFlwuRi2Er1TG6hL3bsMl+ZmVaqZhoaqSB8PD5q31wM50ufRrROkNjWWLcGtO55g885556
2uSPXlXCJs4c4VQcHtp4Y8CvhUxXWP7Zm1y3xh3xvW45wMFQ/zoxnOMwJw/AUCGpRy3o2nVWcqG4
A4cN2wQngtLcVdHf8/aY5OZtoGnc/YF39ABESab8//NDIoU5qBa2mS0hwIpUhJYlJCYmgpPbOzKG
548Rpn8u5m9QR1dkuxZs4Hd2dF4zECHtlJlOeOYKbbuwFzTEbRdU4CM0+6hpvRcBr+xOZoTNtcJK
QL46/BFTnxFwcczBYJcq6UMTMBfWJrdNjHEWMKvzOdy0zOMAPPNGchTKe0Byv3WZG9RH8V4G1Khs
u7HcGT+0nMTRvXzChvsYlNA+n6Wss8OdIbzpp/aqcU4GklMXTthwYW9F4UWNtmHy06oVfOZqLW+7
2i+Ks++W1Tzpls8LtdjXWPdxTfRfLao8ZX3+CFESgMAl7sHPtmN2ztadTbkwcUWUBR+0wGtUWye9
hTT6eLeWrRstACg3+jtt/yqWlz/gZ0XLZ6kXhIXOrhY2UxyXlJNxTZaiHlur9megbc7cvOAKsGt8
4uNSRe2RDfEJTSB4UmKiq0eZcGbFbjzKxAmt6m2u/ZijsS2W9Bah7OacV82+gPZAkD5GZ9a1xe3p
omuvV0o5ZUUA7enK+mgsX4HPStI9oiU6xbcD/XPn9Lxf18Qwdl1uGYrqVqClP1ZS2Ngje1z+ZrAp
21e2LV3QAZmd7K9D5xmu11wS5ekVXdpMriLpdbRIFeEtd+alPz02QczDE9BKjYUMEErnIRaFs28Z
ka0D9/Ofl+6lAjYXLuzpKWoy/cQSq/0dTzUsTKNNjbO5Uswj7JtMMqk+Pe3DGCiY5Nhqe8RvHycv
jevctjWDxQYC9OH1/sg70clNT6ROjQ73UUQlZSYeL9I0FyUImxpxUIftCySU06F/Lqg1CZtmaVE7
Av9EjbzuWmsjDqlS2w4YdSgVMozCj2ST8lzFtPaj4BdDuhaI0rD5EFWhy1ZXuvWTtmRxSbYvbbko
o3bSwhsxHt2duMHVvaEIixGC+NYT6/H9qlsF+QaZi4IL7BiW9NRV5kzysdwxFKlG1KLx5eykN2X6
hAIiQbaKuL+23IlbGcxiMEqaeluLgy8vZJOO7dm6DOdrY8pzQ+k91IOwcVnRLZdZbcJgU3yG4m+E
cBMGmBAPfoxelmHv6ra8yhSmwqnCYUn+zo1i6nn05ZYQGq8NrPhFYksL/qJXvhU503Qzj0ZrEljy
xoUxaye7mBp5Q2e6CxzX3R64SWoY7fSzMFAheuKNC9J9faho06W6jraw80NhLUxi41BSThAdV9oF
IftzpKhMPGqrFtnO/UZXsxxgA6zBYJV/OdpNw86HMvsUhpgYNd6Y8Q2FZ8N/TOKVuquW1Cngnlec
1XM/dvPFbYosKrygUvy/C+biAyG9FEQNjmBqnVLGCMGa7bUe0qm2l4rZnRxDs5EjoUCpVYQhxj3b
5IoCCva/n4cQKij25xHSx6Ea5TMjXhX2Nu2JwBIil/6hF79/HxYzVQvWu6dnc+J/GLLoI1oW8Lhk
diyr0O4qtom4v1SdFGypx7xEl1119j9WovIH+26AZzt2U2YSkc90MleWPL5mHLfjZA2rr1tLK9CQ
qLoSVXoNGavq1DawK5chkakQzk+LErZHc5c9TwkpdFPabWmCCzcUBGRRmLYqvYQ6L44LyRQ8pElt
qAZ8lDAmwOykan+DnrgxZxKpKt0ytVTdnnso6pNK3WShwrq77fysRqjwLUZqTg9mM9CihK2uX0eL
ya4PSI0SzKTnTb4k4PL+DMmyZEhCDWAwJ6jrMmHGAzZEzV4C7KDRmXdHSPtuA9h2oFsHXQlCEKGe
Bx5iAu/hEtPBpxgEp7Pta1uYVfDj+maV5c75XrYvGUtxyxv5JDm4qRgFtjCq8lwV6Ll/6w78Wxof
BI2woKEbGuG5zU0zapC8cNI+1H4VikdSjOt6XAnA/NopB13a3Eb3Xcrs+WfhO7swY+0NStY2R2UA
RvSr7oGko5KLxiyOTnhR43LSlSTTHfF1zZPGTzgcBAV5NEHfpz2Ws8C5qBTPFUy3JGqmLkvUxI6K
pem4FZyUfthB9w76qKyqmpnhq7l9rnOet4AOsbWlBuUpZiedvk3j+CO0poFYlbmok4pK+pqQ3Xwt
aRbdZqMFhTp1CezcA7dtu8o/r2WNmjWMk4kRLtJNlc2BhQ1Jz+V97//CgW9yJGlTw6Qm4l6mhVKJ
y5UrvaLZ8VOTWkfZwFQaU9TczcopyNBUEz6nhE5DXfwA2ghzMHmbSWbS1mHB3pVt0GI60U6zS8Uy
FV8B3IZQQojZVbSznlLxsjyLjBlRz9Ki29gJttNKceoc60BRpfE2jIVcDAKjHJBybml2cUcV6wAo
aRZ8YG6j1bebz0ctFUbtNnEYzaVGntHpekDySUo2zEQkfo7qU64balMNd9bIv9HWs6KouLt4iu9U
TtQGWfKOkv6xRf6kweuFg/MDz5/FOWXq8FE3NfJVFw4D6x6b2NodV1KHucldonlCI0uMK2owoKQp
LulIe/MATpM+KuFY1bCfeuh3qLbuPIPIJ9Gfu44R9twl2pk8UP+Nwu86hZpnAwj35krpOQadEqUZ
qz9s24Dt12t37L5pVMIG8jPjUeORk5XCuC6uKlTehIRHoghxgPJIPv1zD7DYFXuZBaA5twEyeC67
NHXJT7gkAT3uD0y2swLTiYK+cSbdlg1UET8YBLnh6knmHpHDjNsszNatHyHPPp/jsxlGgNKs1Uin
qzXj+bMIX41bPUaFua6EQSpCmaWpWUlvzW/AYjg3hRXlzLMV1TKIJrwW1eAD3/GB5IRyrUSeG+pm
gqFWmBEuaoDcKY8Fe29nY/kO74PUGvoWa2oS+IfTwZERo9eY+uXHMmn/8LuNGNcyRiM4aYZm6ATE
H5fzvphHoUm++CP+CHCn94TizAzMUVxi/5lchtrXigusm/0MpR9eYzka1dNiqLBZh6OjjZtsyT87
jtvFT2fVGhP66QE6hg3fa8YwxpTLTk/25HwbMOKAr5smDHNJd4WWMCkllGdoppzs3E1VqgMcxCYy
W7GZ+zp3rDTSeNaBjo0tlF+pLTa0FC6dPBDaTlG8chqsC9crdB+W0frG8xaYWfIyG+RIkxChVhRn
ZFOCNBHbkL50Iqkd6H2s5EK9k58eIed4PSGf8FB114BaLVYDfTDT/cTHNZCBzQ5j2P857QJ3ENdn
SuKCKFppb8Q5vpW1wzGrisXvYQroM81edu3a037s+5aRqqNHJblBu8r8dnTdBxIY3z54ObFN+kIy
MLaVt+CJOMIhfjQcMS7hgadLg0EBHYugYx5k4o8izTjoGkie2QyYAZ8iWSw9DzLhmUU+dDlElc+Z
OEz/6pPkA0zk/qa2W+tGO3utO2HISkD/47+csiYiJGP464DaaebcqoApSq42ak5rqRu8J/Q5iW3A
Y1B8ZAi/aB/Ve3W+2Al3IahXPEkxgxX1AiT2afHWtes6JfaI25r/gRB4gRDuHfXjCZy79E9jBY1c
V68EkVochccvUGIY3RRBAO6a9jJpnhVpsNGhQEFMFzPX0bVzrfAVFrja0Z0EkjH8gWuthLBopC8C
mz1rM3Dq5CjE9LEXzO+fDnh+qFZcOVQpQmYyeG8uTPiSUT/Kz1btStqRfoxcoeufb+s7tsJIpqyx
SY+BuPw0nGOERVpFnu964d5ZWFBY0ZzLXB2I3BkapLq6cIAHZOYZSdwKXuoNd8dMF1nAVaXOBolz
ag6za4JxdvzBPt+Z4ymHPsxy9NtxUC+yrB9Bkjb11CH7v9CknIVe9QsvKUSmdESW93vF4oofasxk
1Nqg2gfUeMmD0xiz7l8byBa6GyS6nG1g9SDZECqb8CK0jjrfF7HKhavaOWH8fJZQSXBZ2Pr3QExi
x6JVXTM30GcqO2mV1056YCY1/1K8j77w6XN5erGqhbmpPzE7dP8MbJWMOdJ2G1Nnc10lDxjsq3Yy
TVk/1T3B+k15cyxELaMosly/y8B4G4p6uixKa6shw3xumr38F9FDM1j43FSEM9dTwVPgoTHEq1qB
EJFXAkg+SxF47p7kQviTWNCn8XNvMAaewnbLm7qv6gpPCWV4Q/bFgbTbqmGoioT7wOuJkMZBBSK1
1jKzaxoLxRM7M0RtKnBZgzC1CLCagH/q89OPk5aD1l/09ilB5aDYZWrGXikr5yhfeROWX6YCJWCL
Pbg8EygI+mWMeuANJnqFn07zVed121fTHV2gbWQ0FTSCSn8YhKMtaR3RbPytk1kh+heQo6+XFJSc
LE43MtPSGx5w+5czpau6izJQroWjOnQHujrOIuKaqUZuqXD0olxZFfMhedZGuni4k1DKxTr7I8On
e1BsVSb2IxURfhjMu7v6Yw2q7AfRCzhGv8+QwEIGXakkk5EEY2sjnibIjalbb4U6vSxJAl+4SGXh
vqFvPhcsABuqAw06BeRnUhQ62VoOxh3VZqJKtMoalXnYlroDDj6HrTAbNXhK8LlFFox/rAoonYTv
C1AorHQg6nG9VAKC57djay87LWzTf2skliySIOcUkYDMlDA8Bclf9kszzu01tAA7A22jdblCGMzB
znaDyjuhHinXDu9uuJcdGaSugIKqao4i4cQ/Qp6lHWifufxF/ILruKJAKPvNCdFb+pnpFepCHxwW
dzXr3NZ9h0h856EN/5fm5Fn5IWYDXWAPHza/vlbxhZcuvXaNPwUoxpJJ5iDAQsqEKHRbZWPXYNf5
CgNATn8KGEwoG0sAS9GS8S0jKtARcmODLH5IOVurl2S+8T86qSPZ2OtLL3KPIvhcdYM39fjtG/lG
tjFm2oHgwTGIgTjgvSh6O+JYXguz5h801Bl2U3Axi57l0hPd4zktlB3YhiluiowPf8ELs+XNtA9o
QLdFZJ+oKF93DcI+xqty/2mkgEOkaJGkEVhn7LuM1VbthygOFYppSLMwEoHsnOKAqC3dT4TocpF7
POaBgJLLmqIS11Ee4ZKLn055RMZcVoB2FuGYezTjZ/zeD30+fzrh5v344mmOboDFNdc52jgrrC3k
g7Em2n5htRzJSUnGRHykipL4xttppAqETnLRz8Lk7VffedJhAT7j9Mx24VkMtpBmW058LnPjok0N
6buDHiSPVzqSUHVJZr9T1Nsb+alzFzlxhUgaeuIvZmc2YUvyKs441++PBs4pTGKPhXb6WMp4fxnc
eVrqnerroFGcSRg9k32ITOw1Q+7M2GkT7GyTfKloyZv3JU99z1v6Cr7AUo46rgC3OOPmCcv/hR3t
IDI+h+zJ7XgMLW/CWCRQUCL4diIxjv4T8YqaNvt6jOEMz2RpqcoFYCGAd8zN3mhOqx8k5jrcS/ot
fte9LZ1dg5/f9ptdFqtB+X/572MBiZ+Mv1b/BdKV8knIRGLRCSW2SzgYhG78bonFv2j5WdHK8MoR
xaYPIWE88n1Xm/PT4CXfJ4tUnp02yiuxgsOA85aoPjb84CAzLqKdgznqSlcsjEsYgnNuxVjE2N5L
FZ1BP/lJuqVc5w0VA1QN32QwEZa8Mfjevw5zGIY6VnZrbOoxDbes25Ih+0VWPYUGWK+pXw281j5p
Q3M9RPA1Qwf4cptx1QvKVquyj7O+vLvNRmbe+8W9OXdJizvUcLlqqf7T3xNXrbMRLtQfTCF8Scuf
pqDHJ5z7SYLU/muGODafXs+0kmJ8R0OiPaEgbTSj2AXPrKwGqR4nE1D2377EZPxzta2dcJusQvQo
dLudhjAelwB/2MbO7og57X54oUZKxtXocody0cFOABSiMEmEVN1MrQ/Z1p8Jymh+jkN0bRc5xDhi
H9Xqx3iEJjE3BQt0eJ97DFJHZSU/N3+9i8LiYzk0zQoOOtCDiodPDbE3Oww7J1QMEUjWk6Sqc0KB
oXJG09Y3dZZsZXn8iX4eWtYgHrgZlJBCx2txxLn9yyO1zAnmtQe0XD3q6+5AodDfZy32Q6Ci6ENv
Lrpkw5gPJX/DQaP6SQf4P3xM2WYn+nvRbDRtSooxH/saBlciLJhWVDvz3UXhOOLHUE7+wA3rR6fF
fFPq4FoansJ4+V8F+Znpn6VZYXR3ZoDQm7dQQ3fy5YZiKd4sr3BeVW6iGaHcB1Q+YjzoxN0/tEZL
oIgd3PH7ox2/oOR4y0w3BoC71QFffFDVPVxUbWnOvRXNyopB/V8QR6RkVB1YRSmV29on6TRyd4Mw
079l5FVtSOPH5QVwrbZ3Ncugebg5f+eeCzEzC3w01oGXG7Bwbnr4tIFo5F3JYBn5gDGmGaf0XxKp
eaGpWVXXqlVEYhB5nnoRBR9dIV6Wo3TJLbGzD/bAD6O9Wx6o2izIHHSHMhelb7PFeL4ieW4R9noh
gHyWF1WdspxhzcM9nyAOeui6UkTXQI9A4Cnqw0Zfrw33y3pUnQrvwhGPrwUG7aetqWO5HdxWIfh/
LeH5pdVEvnWxkkmyUf3/ewC3z6wMeMnp8WT8+w232Zv44CsBoTW7f044x4Is++5V9qVJCYx/SJu3
vDAp+1ShbDcFGlwb/VruYFFPuSogMBh944FOmevvWAcnM/xrcwiRD/d4JNBB/ch/MsVCipMlR8xO
rIZ7nQRKxs1Vjf4QpjYjRHUa9MV+vGqDMNL/uwiXP/ReLCyVAyJ9Y8gv2CbKiT68zamEbq8l5PjK
uSem6uxMVatEtHLcgy6sLqRZ9K3zdNZSUehuCmEjJsO+yyBr/+fPHzEEAW8J3bjxM4k4uiYMBRNE
fzKhlZcKWQVame1s4gof1yxcUVh/zAzIgwXyFkbYBxeUtmVr/+y/gVy5SZRvWsz1j01wGVGSmmal
QlYmd0we8PCP/44Ex7jSvzNUyioOed5wb2OSFkO2G2fE6MzDQ040So3H68ogeRaWo3ZcPQ1Ccg19
dwA6B7naXAXw88Wt9qKETCxFBFPaCOpzO+44feTJ2o5wG7ZPpaePx3U15qmwQe9TDBtQwsgRsVeL
wl6l/vtnXq65bfo0cxV/xg60c27MRLBdM6wLmLArZIq4M+I5ywbM59O2VF9KN3uZow03y4+7CwYV
rmRa+kkT0brZ0rElUz9YGzVWNouurAzPMHS631Mo9TwuLspVyAaim3MzcqDXIhFAr2b1CmL12TKL
/116p+5bD1ILbvFb3wC7UDvm2+gHN1dHBDpytzEwHFk8Its3wNvZgxq4bQ9bd6uO1Lh4Z0vuGgUe
HnkMc0x5kvjVGDQk6cuJrhQE/QoNi6Tbo1Ipm47gdCs6Oa/zj0CC+TmFftKRtfd9kwuGoY4MoZEI
/Y7mh93MTbfs8nFpwh0cntZYpQh60OXffj0zqTEzngiWmZ8VmChRuBWpyA98TwFZWgFYS88pMVUF
AwPS/hWRjNROXirardFZcR+sDarPoriWcSizyXdsGv9VUhrJYqDCvlB9DV6lItC5c8pW6wgpTxBL
OVEdoSYnfedCpnHtOeras5/ELxC2uArxxA+Z0/8W99pymEzVrygu8eqZtq1jdXlQaqIWd1r3bXHS
uX1aHtDBnF6H2c4w4lUu59IxFYRi6UCcxQ/WL7oFEEQsnW4Tm5szMtm2HETj4Dv45f8OESnIGWEr
Raf3WDe9SJg+4fbYuT4N3P3c8BS9WYpqwseiUuUs70+CO2KR/Y8QHMWoN4DQYCE3W8/zfWB4M5Z6
OOyrMsLboJkGPCTN8TFEk0jwMSD/lopfgZVgIP/8xRBqNNfo0uvLEJgRW+tI8fC0ZZer0LJfQKNm
LbvuhkO226Bj2Wc2BqtvTW0oNwx9Ghbpe9DRSNbDKw3XyBkJtavfAdd3VCXn6Tc5ww5RmM8JwK/j
T5ntlisR0xP57f68CJEJzSu1IZ29iOLTBTUN3NRNxt33A5Ee8FzanIDguaZon+YCsdHbdiw+iTX/
KANRcwZZj4uZmtBQEhRi/UjZlp3/fubWiwJ9ZVCv5snzue7+cFcTAJcEJBsTjzH+iVG9G93BlKHt
cT7ji+d3WbZG6JihNztkVB/p3AzLrRLMdEKpH2VupYxnHlOKGrtSKuVp09RLVryYT9AN6uoy5QcC
Os6p3tqRTkaLZDT32Ftuh9ylUxjW9Wjmlwtjd2Xbicj3Zn6w2agTd+tCEHRs1vD3xe2K5HeZSpJS
Lr3MKlMbag0XKINr1Z792T8Zya6bUWWqEqbXMP/QlHDWcMaAwXF8I4mCdu/Vcz7JL9Flk+3N4lhX
pXXI9nkDnrfqzuCDvWfzCt5DWbQLNZuCfgX5guBiQwmUOCV3/mA17XjAbKMAvBMujlZLjxrSRGPE
wy6qX2q4L7z1GX4Qhipc2/DLmvP1g7ml6Cb+qojcHK96atBWUh3Qkx+nKVwT3xzh1cS9a9IdN3Us
Ua8U5kiGVMZCBz+IT43Gk5BEhSPe0bk59xYYeNWhooN83Y6mPNZTg29ErDDhr14sp41pmGGhXTV6
fqq0OGOIOyYe4F75JbibtVAjrkCdgylsamJXDIZahaXa22n8+RV7yN4hedrMAGSTZLghPyFa6p0f
AeoLghybaN6YM/l4pwQtFxZWFEDwMDMhmiygSx1G/nOyNgEH9f2aCcBAqDncheRIHPhGhX/Q81HE
7bU9oXpytuuMk9LKrfl5fsmwLi8rLNE2H+wjno+LpH0cpSMn2orRrVQIVKXJBBaoJG17Le0VxixW
e3tDM8e9sr5kYzr+RsHQsGEKc0e4td5hELZ/yzlud0ZXuyPCWi6epVnGwVO8q2UVO1b5l9yfwtf8
hd29amS1VNY75y+UOYoawVjAwrTN/uAskowz56vap3RzI39w0e9bOpmbbJV65IUlYMcUxarHGmvS
3E1ca10yPbmEYXw66o8f6goTbqwfuKiAJhsDneGgnmF4FnFqkHsCl/CflKHDDF09pjftyIYi6RX6
NB9BajqssXpBLefGuTM8evwhUIP4SgAkGkBdcJGnq2SGXYkjdLj//eGU9ZZiWeKhXPhyXtj1ef9H
RwdWUEgGKz+CozttlPvdM4SBFvfI9+0Kdo2DcYbPM7sfD5MiYNqyFg0sCiocpvdZLbPTcPB/wHHI
icLhOPL/BG3ygfsuWvBOYLPtvYb159PPkJ3AYaTO/M8Bac90bCEqtSwG3V6LBozVztfq0XiuQf4s
nYJWPR74XpZaIgAbu3BwJXe737q7aCjdlaBiSB4R4ktbd+Ovn4RdmZNuhCWakTY+cBGor3AZDAuE
GUxvwtOBXaqfjS6NPUOtA0Rx6crjaki4SZ9ND0WYnbJCK4Wg/UC4GVcxezz2nx/UC2B/12akrSPG
ByFHEwEZl/3+j9wph++vypO41A6xV+n/bo1tcreO+hU6XwVwPYam/zguotVz+XPccxXTfKoqJ86C
7fNR1TU+FrkrBzcmICwZ1R43zeKtpdkVcpH/bt6uOb5hay6ecUM5w1h5J3W45igFbtRfJjbGgQt0
NHTgt32L+b+QA2HXFBwicp2JLBzX9kNzYLHcgJHrSN/0Md8QmUGDdaN8Qv7WSYe7rf3yTSZoxeRy
/J+ObDg8wB75g4LKt4+gNxbyVNBUwdQsUmxzWeO+jmHwAfo01g8e31jGASPV4oTqhLSCIlSFvI9B
e+ICIPsFr3cDwhvW3oadaG0eA6fVCspEUWD+CHD/y0E4SQmdlwiHViXKA+zVhRhnwzGgNxqE7fcQ
EC3c7CKo3GSNEVUTv4EiSOykPsGTlaRyIM8sjfcDHe12eyUUgV3wQiWdGhN7a6L4JVLm/hjqgejK
j0EQKMagyXZzycgMwrk85FcWSJl3F3+Go/bWBTi9PqvvnGGzvIBdqr8Oy7Zr7EVP8C7R08kSnHUX
CFbLc3M5yKMd32734ToioUke+Rzi1ZVTf5e6JTpithi0UjS90+9iFbyO0yVLT0WCWeTI29JA+dkX
LU1/uVvBcq5hvQa8/o+qrcvtTtUjvEaixSyhQZaJwqFnyHpPniG5SJk2YKw56R0FLcBhz6Sgh1PV
za2pxxzM+zreiIY9Ow8vyvKuTYcy/AReqPK5dswg/c23ETKxHCLcBE6P4IgzguH9NamDI9jQFJ90
PuJ9NCKbai4UblLirXMEa8Lovty5H+YKptZxQbiym9pZvuOCysoOiAIGo2asuGi7QKhy7ucpZIA6
jSEIT9yKXa1N3zwga2hROJbchvtMLhUj/vOSSWoLBeIHqTxr6DhOMAzRKnJ5+NX6tIWCqPA7/h5y
82lZd0rvMPUC6loW7VIn3gHca6U+zgAM3CQgC+pfjpi07SYat+MmeXbBbxN8ptVjYMSfIQLRDU6E
ja8y9bdskAvL/p9tPMq9LozrMJsH9wWvZW9ImPkmASMDMaHSPaQAbfhd/oQP08AWTa2l0nXbtbuE
V0nDVikjvo3VdUgRblcISdo8KmCIbZv2nCvM7O5q62RRrU4s4nDcq8m5qgv1IlCj1tuPXpVSqD0t
iroIPz8KTmC+iI8H1xRzMUOOTIW0EplFV6EX9rfFSYCpIshOcIrot2Ha4uOoXwpT3E/f0hWjXL/R
3/qEj5ukFIROTE/fdN7cp9UIOnEpQPvfvNcnPWRddTttngSz1f2/sKeo2naw6ZJZVHG+Ux1NgPbC
yZhXXj/aWgkwbXx8NeE/uBJ2DWGR57zMnxv1baoxe/487HGpEWsc/RKdi4U02GM8/b4VLpddCJ/V
GkKMdY4nChnQuvwu/hUjKOWZocHL2MME7uJvkUyfANrbsoAC0vK6QgM+rIJ3tQbD7zYylmmMVquq
/tpPKJjXSKK3JRYBKrxA4I8ef1DqUgbwX+AXE06x7t7nZtmhZ/osQ8pwHYbA9jb8p6XJY/XP1Qss
t0PCS/qqE8Xz6xwrDuoppBvVL+7e+i8+dXVRYjAuCjsUH09gzmqRRRtQ7bt2AsSgPF+1gn2fp5z3
3vvpC8hxPrtt30k9at7CpocNyf43RgN0rc9euvh64kgafs7V8EilRT50283mR15kBd12MkTrrhvh
xi59HmZpWLosInbYM0HOL12TRXqAcWwqBcRXmCl0pYKfwGrffepKQL1pxAVNA6phpPj7tx+QSzHY
FDS5zZb+Wzib7AFa4DjXeZOd/pvRFZTLi1WjP2SR12TqGiRmspMPjM0E6E+6k2nFRXAjZcl7aWXf
JAcc6MvWG32GhqzyiiwKZBUykqsHwslQ2OXciE/tZnSQrxLrxTx54gEWm/kOQrWsJEOm3/89G2H9
M2kjClVPR0Nq4xk9sS905ilM4ZnlLNHzW2OID5YOJvaymoSRxG/wkzvbv2yt73Df03oarxXzkqaX
1lhibD6aYKZ9sVJrGGEh2ieSgPcWrahwhPw8T1mmHDn8GikyOgpHjD5R7ukh7NcISJVl/H/8Q66u
JuY5R9K/cTcURI2Y0/BZNvWZ0hb1ERS1zReUloZKjhuiGjqsz15ZA2Qq93ofHVCI3zDhaQG7dJ8w
PXypbnQ57OG4tgu2DhKYLz+EBt9NVGIAw+fIYHGO7GOw1EjPFZ23Hd964pz7l2dxnvRMgMr9AwGY
AcvARh7g6okGY7X0zlGg05zug6oSNPV39b2bGdI3bA3OzJ3Ybaa4UphmU8dPT3pHPs4DvR9wH00Y
TCcZ37t3mAg5Mr/QnAgepWgfycM/spOMN6wP1VPYEi/ASehQgg7UTkDLPU+XJ3Ly1k0Ygn1NYvYH
4NaDycOVKruoqYX1Bz/hhRlzfY/Qc8iSzmBOY1n0JI6Ue1jHmdk/y851eXDF1rxP58YfUgxAMh79
KqbBjC4SsYx1T3kKKaGnsNAkzn5mGylJHUZygH9ILzwmXEpLX719MAMHBCIffRXbb25NkddGSTAO
KaqjJLcMEuIitYw2MQYPMCNfHZGdeHpdGR6HMZBjKTZF1QqfQkHG6Sdvi9frK6Oadl77cBaW4uDq
Kb/KBwZpUBcEu9gJ1vV/EYuZo+Ctdq1nLlwO5sCIBGHwypPURtT2NE0B4roq8EPAgYrDS4HfRQoF
Ju+i0Z7ox1ViQp2sL2wmV3ZLvFuMNlDzX1oOab6CSaHWmKVO9GV1lBYILXgK6oVrwi4dYTKyohct
6xXNemaXM+cTlSE/aLPwey//l4zzC11/WOTNHDjsHKrQLAwB/c+6v8nh+VqGDRVM4+/A/4Awt76p
lNSoBGJoKq4+yVpfX7AtZ6Z2vq/IcRd2eu849w9sLWzF1DvY46fKlY2icwWB4CwnNk7bxJ3vGQTx
XQu9mwuHoFVijuQLiITjpQyzcPaR4OZwLRBvrdPQZf16gGgH5jpPVBNrm5sQIJs2pm9/9pFUbzI3
I0AyW1zGmrXcFD6tXxchw149tHPIwFTP+IgvIsxbGgf8VH3XA4wCWNe7R+3g7ZRL/3ONUi7MH+kz
XEFff9e2W4D7k06tGL+aNaG6hI+M8UiAiUGopFjGNMqR2kLSIP/ehrhoyqi1j8S6Nnx9HkYOkwwe
a7ZHaYyt00KDEPFFO91UmC7XYe+uuoSR8mOlHM9I3oY61TyVKpxyYx6rAf9IUfbpLTKjj2hI5Uxq
AlOODIHTCIgd3qv2i6A5HxIo5iyYHivTaFEyInF7GS96PNCKnvNJHi643BvpyOoKBzDfcvFr2k8x
R1IbRSH9KtvvKz3WerOONruAeG6dydlyMjisAJMwHUzSNRzo8VBwU5ZFbng3LxmoQFuu4h8jldKm
puzzh3oKklcSrFPqHFtbtbcKoOYfsxfLpEKPsoVRQVJq3DkRWm6C1tI3ecmnWZihSeKKJgpWpmyC
tHSd6icAUedMFp0uIemloacUJhjL3/sfaLIFMlYfrMZ+Lp3kd1g/q285pot3cD/H+glwyvPhBFTZ
1QwGSstDc0p1kLSxme81XjdQNqLRnH66+ogTdE6HJU6UqiWrggCb9bmNQuKptBPN6ruNr05aUMfc
CY1XsHqQzlMcTdegVvVPi9B+fM49wokB+wscYNG7xAZoVyUWnuV3P7vLT+iGbew834AAnjFo39SY
uMgO4VvwVSU5aerMDRJlZrZ9TH+uMo4agU6op72l+xYGgaoYEqNKw9CovI0XppCUHWzexfLvEv6b
LgcZ814G5zm7dEbvg1uYx7Wt3frsMgMFs5MNFsjs2UmbHuUToXhVcVr3ViieLscA79qBmEXsFuCr
Wj1cWG4CPBmiqQc80ghhve2yw+3Td5jkNXaPpYugqgfgGE4k1sBqPBXIPDhVbb+1vJ535G8Pq0Lj
oXQ7zeqaZC0L4psTW+dHrOZ6Pynfw1lx5S3yR3655wQ+Ny6lZ3S58QeXRibUXq29FyXCIcMC5Usa
v63Th5i95N8l7mFU66D3NfHhmXGokPPSY/E5Af4oTcLiPt2njb/4oCo3Z6aaOIOtEWZl4oFJcQQq
BVCpK65Gyp7NI+kepwBkISyi6Fz4ynZ5AkXeAIHQPJwnUs3KQJZE+OVQdpKpXd0+z+EYATLAOJs5
0a84SKjaTVlYh+KOJjSDRRjwohcTSxma3JYZJMPswJYmfO0f2f4/OTCUgUG/7ipJIwMr0a40OEli
ou0v1Y1hDeFSa5ab99zzccQmM4agfzDI+x3r7L4YmWOI44L/L1YDU7+f1WBHRtyR7w2L2FBY67Y5
4XD7kkmcyloAHwbKOL9Js29gq+WauFwvgbEFsdqXBOFQ1CNsg6QLyTaxGbvMoM0aukAWHDIH3Qza
Keguvc+HjPdQzB3GHQEJ6G2UXnjVTC1KIS8s9KiH74UjkBtsPUS4RXflSP13eE2l1KlF8l+gWDGA
nMmVxi7VMCsfaNyZGecPJqTuX2vsZOJM7GPe95taj8whmF8xGwH+2mNuJ51YTpAgGRmyUmfJvVS+
6qnUcAd/P5Ndrd+7tmD+hDGmyaESkRHceSNfliLqXv17hftgN7t6d3RDUEcdYzWe5+AcaF4cpaTZ
WyX9V9kP8lsIHWGYQ/irDuZg622Qk7dbJ1ty8/iHB+S32KmGSqIUQ2h8exqN1nQ6p7VicC6DHKZC
hDUs6iRKnlzhjkH5m6yNpRWfp/GzH1WLnb9XBtciMEej/SdEOdzNbXBfJ/9RjravFD/zV+EwVjGO
/O3j+7gTlaX8gIxfM6AXGQU60EGqmDsZOiYeq12N3bx7Y4LK393RX7GvkDP0P3WuAcrHsMbxlgic
DsORai0+0O/h/l9etxMw2qsRYstNxgOq4e9KBGNLjXGxIVAn0RavmzCfby0tllyFY80wTXDAjSja
liqI2IhCWHtfwa50vLYe+UKdJiLSK1h9Ajaaqsg/5LPKgAOZJQVSYXc+w1dMwPlgDs7oTNGB+tCM
7YIkYksrdaGyE4lmwEMJzICxkoxDNUmYmzw2vLIIpdS2OxG0RAk7UnqngrcO9ZMIE0M8B8a1ny1V
o8Ws4WI4A6sm3NmIcUPJuRgU2vydMGxPnX52sdXir8UoyBM8WmmyXo9l4jCfz6stSc3CzrrfhZEQ
CnQPrtm+Llo7KhZ080fxw6zhXb9JgujnH1+D5B00LSrnv/nyyik/Ea1HfUxNO72gEFGbm/mBdfPR
I3oI6fv2sjSsfDpa00XHwaL1g4fzOydFSUEGyTNnIXuj4UKgZBXWEt6WtkPovvY8XrwlYJ3PHnCR
8qjHzLw/toSQelSqx2CyDwoVf2luwkZs6Sl1eUVyYVunhL5kpnPDFFCELYTECKl3R+Ji4GnM04m1
WPVzUL0PKCPXnHlQROw5HM4mKAGu0YDjv2kA9JWAh5b09jAXDsRzzn44VQp49OrGXvd8rqdFr7WO
I7GN7rhVH4rlSriwth4pxiqKJWBn6uQ+fXambAC7mGFT9E6LHXmdGaRrMx3PF7puqWZV0pMNdYW2
pKQBgkc1UqAyDyVAJjDi424piWyJJfvu6GqEnWiQMGA5b/ZaGn5TYJBGTBHbLc4BUIBPDSv7mJUL
Omxr0t5sgEpN5VyrFYNPSDO01snI6nvkaIw6kyuO9rI49BD+VnuFXXCRp67dc276TBXMrd3jSpyW
oqv+d1JYGjTRiCSWGXUCRDxu7lpaxSfLI5013uBI7S2K7BDl8LhNIsnlGah9Q62iTABWD3fbxP1t
CWn1kpZe9Nb5L5OcAfXbvNvgwSMDlfP0Q0R1421pNQiSpwxvynUSuZMoBM1HAPOD6c24AGnNb26A
9WWd52Ww3bUvuZDHxfDve+r9mayxM5x61u27zLwA7iB+OynKg3u83Tt21eQgcCvs1+fnnFmR2km/
QN1rYtYqboZFHV1L1psIR8Vi4jxp/XbskmA27+pKnBcXRBCyV1tnxnEHbUgJE1e9tmjFmY3d1k8R
GYK8Dso+VG+6WG7/x4GPg81081ZN4PrCn5QdQ9OSIn77kcqoj69L/wOCl9/aUDSFyEwr7lEP57TO
gP3dDH9y8cDa4KV9G0V2uwwrjHblD/dG/Bik9hiFvBCFZUcoH7fEnEqiHRmS18PpEkhSvIXFI8st
GUY6/oxqg4gFKXw3cLXxxbXaEn75tPgmIj7HkhBesGrTl1Kqm9Wfau6P7G2N3kHjEXNvcosBGPbh
/Crg+YNIHzvlMJ8SgHjHnI7PS/gwYL4rwGS0BkK3IZRPwqHLY0LHJZQS639BhhCRAEdr3/BO9v+Z
89vtqg2eMh62+jcnzsk9A5xW/ttq0SeBpDi3CVvKXUFC/PVnwEGG0pQcgNV7ASJ7KFyAgufvXfLS
dkwi3Kt7YFqjLfhAEM2jB1H25tQQIyvXTEQG8KGYoMI+442N231b3Kg2YoCH9k302+jyLm5S1bLs
mjsyf1ddbCbEUfqapNTlRZrswIlgKA9MkNjmeHZSsxvw2+al2ST4iIpI3rhs6WCoFd4KR+s2BuHP
o3SGTUqsWqUE9ocITCcaljhiuieoH/VOVZrRqpYNcL5AgF8ou1mPJh3LcqXPYsOgYOBo4tqWIowN
SYXF7ZoZ4nIMEAo8lNiylVHISF/FMiTuaelJ788SKEot44QUeWCUirIStLt2xUi/c4evKK2docrc
FAMEAyo3HPVmgljiHF6nJPuduqxMKpGGZAHQFFle8S7bxzFnhjLHd3oPcf2tE5EWgVQGw7bc7/y0
GjtUyyZDM85yqTnxSnkfdwiofCIdLIT4JdJWqzdtOwZ3xsa03v4ysEyJO783EYIhPNF7MY5pCfND
vhvx1cfsutBVHrloJhb7ub+qY11oxFF6FLnxXe5w6vemr2zs77qUE/Wu3txXb0tn3DQh96ELxxbk
dFfQlgXGHTVHxf4H2lJH+Q0Hl+l9x0bQSeSyFf6VLOfIwO//Vjr8RZ/ZyU80eh+mK92SOZPn9fa9
OKZaRRi3F2mJZbphk/rp3mqrwdaQtiXC1luENabwJoBLBhGwvWuYBRAzbvwVUeGog3ICpKBOPXZz
3hIfvRRdebl8NHw617JImHbWvzss6Fbz0w5lVbprC4DrZCjR9kx0s1By+coYQa+gv79YTxdkjgpn
a9o+86u+f8HpJ2JXmPMcCx5WF++Sx9pX55hsGqMS2cxOo71ms/q1ddMVaLvPpf5kNj+BBzZzZfrd
rStbRM30+aBTdaczcX8kRwFeICvh8KiXJYHbHFqAZw9kKpQkNhlxJ5UysmqDw3Tn9hEX8y1yan/A
QZabN7i/2meRo6FJVrHgQqsMg36QMXQaGEv9Rp2BP7pKpsjWUX9NiH0t5Lslmm7TmHscSYM8Y/tx
roKBRygWglMBgTMjk9+GGHc2uM2ugcy0Eh2N8r/7rNhWPCuAVi0CCSmqyCW+CyCsgSCQqYGpHxs1
iANx49cnsIepoQvXrvLehTywngVRxZhSzKdL9GtsWCh3ZdTUjxLcshhp8dRFtaOg0ODfjNqwdfVd
jmmkCvG+jeMzHsKmm9WHuM/yRNTI9gDILhKV+h930ZOEZzvkjDiq4Am0miUI2lMcpVjTkywZrida
LPVuJJAYGFLrv9OVoMJplmy8zoYwJGvNmlMSi918bnesPqsXqh7DROpIn5WSCuAsdas5ZbvimuHx
ZmB8guJT/oNhI1h4biwHfWh9f9oQB8R+TTfQ2cwhHzASARlZDiw2aAJy4dQz8l6EtmbtuUSiXGsr
icvbmqGzMTqKjypASUs4dqri0O8sovLMhWJTtAdM2/E3qRFUXB/q8UdvIiLYKBAuw1cokZ+fH2Ww
T12Gb49ZysxDTUOmQYD5crW8zolDh00BBfQhcvlj0s6F7cPJMwWzr9u0K9KK5QrpdxVwGVBz4A5K
pUxIeHl8Qu4rxjTIbl3jOxAJu9WZUUQBF5t9m/ndrt2JnZrDPBnRpnnlqpgH+UTmO0Q6RNykz5Lo
Jf5Vk47hj3+4uVpZcWXnn77sp/B+qIT3KcQmcoG9r8f4roiUHxH0oWL/Ivo9bKnXjCYBRpZc/Tfv
UNNHyd6jNfPsZzE+CyYGnDSDTSwUPlY+VB0sKTvjtGZDqpIvMR1/luEj8tP5F/Qdas7uxYoHX/h7
SHriFt94F7XUz5MUHU1ZjlxevG4rdW8r3KyCM36G9afAOamapvkNjjOHKvXULX40SgX//XeO2Qwp
zdJMb79d7mGLOTVs5dFtmO5dHQCiBwE+1sN8e3EFn/QdasUy3UeJNoxrn26KcfofNY9KXKHsyqOO
j/Mm7KlQH6Uwx8xRDTJ8AlGBV2k2pUgtPBq6Lb1uNYVKE41zQFJSZe55Mt8ibnnuO03u37B/aUu4
oc52ylw+IoXXNC+Pl/SyAOfy88IFwNvs+ima3XtYBvfAItbMUJJ2Kuf5AfN/Bq/UrwMLBqYRVlX4
/10w9SGVKnoJnyLKJ1/Qf1ZpjlGr/mVNUGu3lKVbI7Hb9F0rwidY20DIz9tK3lymPZ98CjTTJAG1
7g27A50VpyJmf3V2cHuvsWf7g72QE8WLR2YY1GEcO99iGfHXqLCDc8orRFPLyx2fFSQCG35cv8jE
xygxEvAcj9oOeP0rhlsdhm0hZpvXtvi7Ih2KmjUZDO8dTgzLrZmTgo3FDp2CvU3qnNxNUUVa22Vl
8nukC4livQaNIzUbLjwsXYctbrZ1hKtwLZzd5qrubwDLPcIY+kDlI6t5UNUj3RnIQLBLtf/C+VPF
iTWa7IQedhbndyc7PXmG/sNJqPvKyzTGf04VwZz4PTbqJtbnO9oOnU1ExZWicfXtMz1VSDHt3AB8
aVEa8XQ3t5+Ch0540Jq5x9PXLsWYuVhrG5bfQFt39MPRJGu7j56WIi0W6WaSZZ6oJWufYms818iJ
I7tf2K9egFm0q6zgGfP+WAXYylhLu8OeyeZhXNizZThTLLs/ZgVcJYzLklw8UwdWuHw3VdgvtzD8
t5/LvIYUsl1bDfYA9AUYdJyhEKGDqL1ZCOpa+uRAsmjeWpmMFV/gQKQbQJh1KkjmMVGMfxLUuRAL
KGBaEbi5ekTRzF2ovXsHLqBGJLpn9i7wPohGRGOI0RGPIZQM+p/WU3HCosFalDX73IaBSNKdaL60
sgUR7+lDz9o9ZJ2f0FESP9+NNh7W0aSPwWwtwyk6UgGIEJ5XetG7aHRSkXdZ38J+Sz/UmBM+lW+G
BO7AurTgAqXvCTPOvp3gTuK/X3/cpRIabF5eXpzLYznTuZ+tCurA3vyG9D4fJYX0R1DAVCFohkR8
wb7X8ysSBY3JJLn+KQrBVEhK1RFMktB9EBWcXezmBCCFIVZv0cb/dV1lg3DoWIh+jhvKqvCHSLsI
lIaT8F2g8Kn/56paS8qiZOh5eluLN2AqgpK4j4xR5jNWOSF4QFYE1pJvA59E8/No0koQhO6K3HAQ
TvV6Lic/uXLbaetOKqsEbZ2PqbyeUwVrz011U78Ym8b8TXiq013T8cPgb8Q4ecKD2aDgJ1XryCpj
TBW7odtqaVuO3b4xGM+grnXm+QwVHw3RWSgZ4xuru98ldRhDFPKd3swhtsG1vB6yPsn+wK9/GMYA
uB7Ytb0KQ3L0txu9Ctb4xNffeJy/ADzfF9b27bho+C6mRZF+DGgtW8IzYxCWpUqChrWnSmp/8mp8
tHaifhdXK6dbo5KM4qYAQaphdvsr5juALz4ABRQeLBWvQPTDI8myUz7yHnL5Wj4kgl/zDW2Tlsi5
AXJ1EtQ1dmPCEi+VehzoLBgIGJbadra82Oyp9wPvRVRJKDqf95UxNfXoE7aeMLGKJAbX1OeYGqO9
o+mo7ufPnxBkXJ/wHLUwcUvUV1r6pl6/a5EToSX/UgMxMr8KP899IcPKWvnptU6SD8vWdVBuR959
cFkmWFPx+zeWAw+vOVQ2ILWBeDVbs0mEKH9ReVsiotu92+rfzdgjr+aElH6tetVutXoAP4aHidI2
upOgWlmGwWaVl2QOd7u1howbJb4TBIQYNdydPSg2Pg1A4nmXVuu/8vXsW5M1rS62cdHjtKZUQppY
2qAmsN8iNZEHSGA7cDbXK4Ktrc8oncl7ZdIjSRh7V+DO0EO7l94am3xP4Ebj+O3NFqqpOzeslvtU
KttLVHzzncb2JmUrKG/3dl/U7KYWr2CgjgKEevZEA0EHz5BnPSS/18MY+WH/FjVczKgfKAY5uIJs
SBektpf3Ji0EgQj2aX0E/q8sot63NQ6B5J9eRff4rBz8SVA+7Y7jT9O5xN2QCl/ZZhXnbEs+9uaZ
tLUejjAQZ9T9GR3ac4LRU365aGQVrtKxZ3xi1td92A90lFIj4q5NSgLqn0LCxcyPHL9p7qM+CU6v
5VBvsIEzFCkLgx5ZcsNzUwjGh6D9z/P4Hdk3PcO2a40oacR6dR5/+h7Sj/7xhpE1Gd4yeHYlClQW
5nG1dXxB13Wps8eiHonjUYf+XOT5HXsbSuo1iFHryzMJYK4Jx16V6RpGE7gjODCEvL/69AyhkqOq
XWTv7y39R8O9kMtHcHDAhUfKGdHJMoZBMFIQoQLNj/MMD4WOp/1MBDTWvPQXe/0HxRqnRkG5t4+2
SXXb4LQh/0iCCUf1O3iepf0IR6uPOLAu8Mu190FKRlzoMg7+Ac57x5+IM5GR7qPj1gR0svZ5l8Bs
sKBtsc4aWTl6PPbZo6LwK1AWZLVxiN/SZaVk6M3nFQwTLA2ifwtTYkZulbGsDABvC7mu7t0U4Tbs
XEmiYAkz0dwKTgUvx3Wvszfhc4xIMMaUS1dgeOzYLj5qzFA8Clw5/ag5oF9vgyxF5xUbgKoUc3+y
ja3u6lChyPS/oJoB0RV5eIGqegoONIWLzFAzrPwMNEIXYfH+cfIeQfqDAs9hW5ft4UpVGp46+Am/
bmUokRyRD4AEzHdJyac0uBMJ2oWF1s/efj01LhDi6o9o2Nt+EvAzGJcIHJih4/WaL9+vUdAuzZxP
K3k6oigInzEplnqYqgkpo0toHVHoEhD322jLds8DXprVVLUVwGXM+vMuFKbaOuwjhodEFzFh2NrA
L9x0EcVFFTwpAGoKycjX04L/5/I4bgWDwqyZwGVS6JpVwGwiWEAYN+JdhgUsL9t0B6yRalXBgP6n
Nv8V39z7R43hwrMKkIDWaoU3OTm85c35RDbZCWkrcMIXo5PftfHnoDpC/Cs9RXpNEKNw3DWgxA7c
HD+cy50OhO+CHo50vpyst1QmoFQVAPIlK5wlgpvyUyB2dyxzv/wXziXcN/RFYtdghX7izDm/2ka7
jOM0iu5v6MzGIxP4Vf7NS+KoED1ZvSPFr6+sxJA0wNR9kvZgfsNTkC/hZVoNjQ+6m/8FeOqc1mLs
1onlHoRzlc+xF29y9HWRUVuXccME2JCcxZK02/tA4+NeCGvRcapxBl5ASjt0QfcCuVED7GmLSYHM
/3U71TZJ2u9958MC75pbod2uY/WX5XRfmn3NHQJcCwmMKEFbOguWjo1yrDSpsU+1HawsTZSvGcXr
Lc7jNXMhnAJuaWlhssr1pKvsrKKJsYTvp+nWoWwTaZo6MxdreLqtUVi08sGsib9RpSlNYKiMdGjQ
VnW+l06murjEJ/KXSerrWaMncoF4D3HScap/b5tOUovN7ZH3KPUVc7P00pW8YD5MIbGcq8x2+WrN
d/jtCuJfe9pF3uTCpMNfB5gUTSeA9sAiwKVzgrpUNLEY1Y7GmxFfceyK6tTy+VOIHnXaTb06bsvd
F2IQVJgSplPF3jUPhcDFr6/BgPzO3nMBJC28W/r/goNqnu6MgHS1EQ5Uptnoaa00FJCPFEdfA8IR
A9NQ3bGPqB9qqnYcc98ndSoAmMTqYMgrgDG2RWYmF8+QkFVK/Z7aFKETb5ezg3hdmhP4iwrHxCLr
6qGEkbPFyHpNZQH3m6WtHNfp2oB/nTwTrDtyviIZhSet1Av1R9NMSPt6hNqVmIagOwRZY95YAdF2
+KSyc3FcZfYLmXwZbonqAg178FZXxY8T4hyrp0C6eQvdZZ6m5x40pmDXtAG/q3aIrhdO2MLDnF9S
TPb4FASqbxkd7BVmIFSRnThtlqg5I2F4KBJfjMNB0E17wo5Oz+bXZbJGKlH9iwYMoYdlre3tVc8a
dWhPZEkOELJTiCbVTGtcueviUgw9mqMFn7Vy1aEPOd8ESipYgO00IlGrEVJG3M3OG8UbQwF7bm5j
67BZ3I/4PbUpXNA6BgqY+IUXLj2MzZ/hUJzJAYF8XHGVe8gaaecj/f+Oc/3kDpoWC9FwAPb2D2DC
iqokMwsD+zJaszJuPJUzHc8sYLSiNCnuBjHW4WC3MUvgf5tOk7XjOeHbIBTcQCWhEf4nFmRaVyXi
XDpdaNPAuvqdhU5y0/rVYKVbdTZYg6WXm75SHtfv0QDEHg1L6C7ItgDeATL0Es8U65doirjn/nur
+vhPY9aQpLzwJ95X9AAv00QbrGl4tPKxSASsae7U0nGSYUZawrPQMQT8xMsLhrsDBGiTUc+VLYHw
Y+Td/DNv7a1a4ILsf9vJAJyZGoulgNoWTFA7M9AJmMetCd2MOP8vhPWTD71uKMJ2HC9I7WyDfYo0
qK4078MisK9crYw5PosU8JpRmJomikyWBJg7B/Lv5Zbmq/V3uJqxISzQBI2dFkVWonBn1r9QVJk1
9pwRl4YowUTmb8Y1nzzbyqHzMFf70tEAGe64h3/gdiEwexiH1za8akzqfhlMX1tUL6zl2T7iFM3x
wc7w1lK7P5vRo32vsM6smBm8slPzsdzO47txLs0C7xELyx84vdsUWvVCJalpUGoRShMwcgkDeZ45
UwK/B67lWTFnF0gl09V7aKlZFTp/6GmvZl1PphvbhuBHevY8lAr3VHSKzpm2w6mPqKddbC7E+VzF
obXkdIuK1t6heVBRDVhDRsmnEC6c1sudnn0cB7Ch+beVzOc7qvpweILTXyCNwYsdKAKaaIwXhhAF
yLG7DInyvzLe/IPDbigQHoEE2k8JltkJfGnnZhRgM3TmwUpJBpxdg0O8XRBg3w5qyDhv6zm/8HVA
ciUjzZ2pFsAMukX1wktfcN7Y6DqgU0N4i8ppwgEEqaiR4aP36783g8b+Jy9VXh8upsR+zrskj7la
ePbPRfprW9OEyOKbeitH74UFplScdUZaPbkiQKNHjFCKtWvQwdOzNIz2iyAuyG9ClhIcfjwQqp4Q
bS7aq4LReedUk16T/uDOi+h1qofy34mOjv6eIcOzwadZNLkH/zkW/2lcsu5/gDriy19+HYPc+xvq
uf/aqz3cudDJ0/uiRtBvgWkjS3oNy8/tkabxuCjoj14vkrhEVD0TUqjbK4wE0m77irUiprTZZheJ
KmzXtoCeQBvln18HiQbpd14TW55jghyFmex1tZR6GZy0DarnzR3tCZU8a4d0rLtFS34Sj1oPJUGv
tfjmphQUf3OF+3WghXd/CTG3D2dqy61xDhXDgPylq0pKXJGs79C7GDsks4lZQnyfNnACmf24nSJN
OqthN+QRTxoraSOi9HEoXNafCKEuEI9m2N8U8vcMXC/gDworlm9mL7s07ppsPI5UiqzTBCuynVkt
QI6ysbs+/aAtPabTCdBKKt4HcPXC7kRUkz8e0SwG9mx0/ykhQ0TJveHJUkG9M3fPh6wMKOtwTtVL
Aa78g3cJmhs6wOs2/77dI9/YTK1Pj41iJhaILN+8t3A5LzYWAH66guikHvX852DTvWNy0uPbTgbl
hwwJwjbXFSnaZC9ZecdON+Vo9gi+4AHbPZBAX7e4YBMuwPmuhZSkhHMIZgs2RvQfVCkn18MlhJcD
ntkTARp0iDnEgWpwYiQDKuIMNu7fXY3HT9wSqbQwp9o9+ErvgbAGsfKx6dIRCLTdjefFFp6UQjWZ
cbNjVtWqcfK/uTkv9Xz0KzNprPsz5R5lv53XbgfDj8lr3JVyWzCO3Fq6bOoFKUISBmLhdUCYMBNz
83YjmlbwiWQTo1So0stOXPlAcPO+kYfnpEcyGRQ/VXPvfAJPG/UX3wHgkW5P2IkXsMU0e5SQSmzf
dzZzzuHNKkvIjC7aCcVt5KIeHcelApraMs3y8IhWrdOBKFTQj+sOfO+17148YPAWA44TYn6JyglK
yqoq4N7a/Zb1JnmPyfzlLOyBBgJUxK1o7gbJJT13nyWsFIx15hhETtUbqdZQUvfqxHqQsAJBQCn0
N5BoJri0jk+xqVBrL7HD5HQODGMRmO0o00F6XW1xQQ8rMiAj2yAF6hKjx2uXmmuHdwBGgLZ44r+c
UiN/Bhkdozp1QlG919gatt77+hmgDii57ZLew7H4MIfLGEJ831pQJPWWj9ZdVmTtJYbNICAv4Gzx
8OI5HRJJhNHL4aqnq/xx87tAexBhUFRWHT6X/EItGEbcW9ldhOlqN2g/z6Qt+X4SdCRSYuWSQg4E
og4mpLoQyXr76yMVQRIlwxuHqGF+mPZGMqN0oT0JhG6WxCHg7k4zxMLgiJ+MSwgpAc4T6Fo2+WR5
xKsd46/pSmO5v7/OaR6XS4IrEZRlyilX/QNH9vVnNN4lXgSmxF1WsaIF3K3+UMU1wjJgOZWE0ISV
aqIO28tMRT0xJhkz7+UFPY3K6GWgkqQBRWnkPu4mjo6On51kIlXbcbX6jiBjbE83KUYKodVtPV2C
+9s9UtIR7MGdPWkWmxp+FiY/03GoB6TVSYM3WSvfocnNcdFI+iIzSE/d6aR4WHy5tAv4G7T9zwDu
25fmq1hYMVsEmmA7cXkQmKItsSQEjUny04HjAYLKOsvbyWETcQj7Xt8KsZEuIlbRC0j1qO7EdNgf
OlsNnf+q19V5acBMvj9GoRw8tb3+7eKSOd4MOZBpyyRh5cD7Qr8ShR7L1FXwe1RIh/mBb4QPoWU7
8Zjq4pELLbxOdz7dvk7sOgZot4VK188Vg1WJrbpOc59eSP6vstMTxFx14udj5AzIGP7suOd5scXe
c7aP0a7VAf3wzALiv5ribz5zIEhspH7z54auLzSWgk8CyF5S/HmTygAPLEGMTYgtn6gPMH80enc4
KJIzlvKcbFa34xo83IfESvV7BfmKe+bRPmsvUTZ4SH8DYRqzFPKZDJFF5GOvkJfAwO0wy/giM5qr
apLAWQa/CiJckorZbJbCWkY+leEOFshAPot1BXr4c/TRLYrHUJ9taHfnSrNFM9oPbInxyYtpHD4t
k0F7FmYtMZ2lCAtIAhFcHEY/JNkS4yMpOzn8oGrNlDnFCKRFcATkjS2emLFXH85zyPqleNjKr8bY
GtDjlXyMnUqGsTkK5h8lYUd2JyBGtLGvntWSm8NHTvLW1YkNmQkxW6ElnDcM7OuE2wZUg5PvLkl2
y+tzzs3fUEmlCCPEP4TqqEkppW0KL1IqpZoWZ9o8fTI5WYayKyN+U/YXZpHnkl/i/Vz4X7jC1wbJ
v52K3uFOHSpU0PP//tnynfNyDtOk+NMbByOb9CEGNs46Gl7eRL+UNWhYV+XUUTXL4PTEyCJkcHnj
2HCsZXN4hevjVmK+eiX/+xRxsu9yaahS7BS9xFzAXEGQJT69iWl6JQJlmFFbyueMUFrVHBO/K0Oj
dktw2yqbVHIL1Dc0D4vxlMyYWgNZmGxh70o/PP1uJOttgiHLM/LS37yBddGJKx198Y2jDS/vg24z
FnwAdunbpFXSNBLoi2WRkeJN/l4NGwUJry6wSXhrlNndxQv8nSTA00l7+vTfRpIR++1kYHQM8lpU
MHyGxCZW4vFvg4kLgOdpABK1sZvGZO6yGZ3GKHRawZwY3FzSMchlppJFfeApRKbVfYsU+gLyDaK8
BleJuO839ZZ/PbViR41kzPxE54ve4OP8infZ3XxOEJxCc3WqWM8GTme5OEEMPoPLx85JY2nDjY5q
zGdr0CCu6LL9ahUaw4jwL3V7qZ8YD7xe1fTp6/1sqSQghwrXRY8BC1TcXHbSgqcBKHHE7dTdCbyu
QL4gKQ12vyDP/ktSEqzy+4nQBMNpAPGnru9kSQbk/BL85xGXklDqqYXdv/cDjX9MONiiVpZAAWyD
tVoEZYwHfbC3UftPU3Tyu0yPvSlxxpiUNpTfWGlC1Owcmye9P7q7DmNbPy2p6GwEYV18GxDjvAfv
px/9B5dg0V1MbUyn2JBbiDoroeM3SRpgXVh6/tl2gyqoejhagGHgAs/9P//HUlSztFLeGcW85hW5
kmHjCDnTJ8WossTo6z5iIVdzmwpGHW8VCXF21Ma+nbM75GhlsVZTgvHrU7Jq+yvIqwA8vmq8L28L
9poJW9ycGO0ooL4pQV1/jiq7usBiNxcDR6L5uiN3REbOFfNVv77CBzcP9LpASmL/Dn214jct4rIK
dLlehfYOB+VL5fosTzUGDRt7YNkNISD6/Ip3UKhQUxS71Z/UxZI3HdJHkqz8JU1z5hCRRKiaA8zJ
SO+DRkGil2Vtxh5m7fNiNI+ufhIQ0nVKYAM8q9l+67bVLFKrrJO3TwrAGZcBW79zIcydHC/rQLFH
iqRdPrP/v+VoL9Q/5Obv4/3cCPLg+ns7J/liOos0HB1D0Dc+2ND/8OAV7tUambrSDyB1cdXZfNVu
0KRjY424vNZ9ELxk9HcMiTJSVD+nOhsT6IiGLQ055R4x56ybCfbHbOxSNlqUPlkAk/uxs7iQacEv
+2T6gA1IxvvcG1HxPrEy676LYI+YkxLj01NgY48adZelAGr32H9RzoP6E/x2eTYE4GsmkYX93Ag3
n9y9ebzgKMAR7wZHqfVrG2xsVJORo6DNq/cfLz2HBI2owjdR9lEACaFIfjEBHqLhCeuyemvYEAE6
LAs3pGya24slox+wJPXMGGvUdSALbLxRgaviCrl2l9eZ2nJ8SXXL4YYICDSEwYq9E+EuJN1A7Kns
mDQplJkHkF7sU5299S+7uh9LCjx7ENK1qGdJUpux31mSXn3PyRvXx3YbnQa8to62kndT5GEktoYm
vyf0Bkf6WNjEHRHr5nwNiJMluWsAvWdJ2y7PiKGhS+UkZSCTIt4889BcOeU472ACDK5a3ZGbtFT2
TAn6R11gRriPrse01y+0MkSjKEsrfQhUFzj0S+0+N0wpgIIktgoigNACaEBUetRURJHpBc4UNFu5
kPSyVCGUT+oBO1peGKiMFqSaawGaiqyYVqzAyQVHEGzUTVzLNoJB+Kg4QWRbJ52Ru67/LbgMndIA
q4hpE55wcr6/5v7RmS6EveD8v3K9t5x0TPL//uycGiZwjaKiEffyu5gIwUKAihH/KRdZQlns4u7v
qWd93/+y6Y0VRueVQg61QEhVDLgH3AS8ikdmqFJYR8NpELtTpZQaOBr2j1JJ55lxAHEoi6k5npYx
rXVHNiXXbJseM5azRd8C6QqLf6r6jnZEZROvQH/j5NRCsMZ5PvPZ0kFNyhOlYWe0xzfUBUv7Tosx
q2s3lNzr34UMVSZO4YHZ3RaSLkRAESPNr/sO1euGpNB2oCzHBVkZtuO8SnG9j7Is1/O6ER+z8IKH
9yEh9Fwk14++tDEgoRubOwb1NAZ3C6+P5LPADeFeCfTW1Dcdk8NoM9Ic/NYjLDeJRbXxUsZpXpMs
5+9lYa/qMsegPF4CxmDRoseu0pMkd3VGyzvExs6SD9pEs3EzBT67AfijHiOZF1ZLQAc9ahYQCinl
B5oOIJR1JGIeqLX69Sfmmby08I4EYjFGktVjBCQ+0g145tJBa2RZhYBBipN5YyEGkSfmjbJ3fEJ5
yb1WAsxHPoIeUGstcqIpEDnAIEE2hrRY2SwDXQZtKadHb3DIyZLyEeC+kcxFvde+gjTlYV3nvgog
mRV7NU1S6JPIFHbRF+Zy720Um46bBSsEhgQe4WKXYqvYYO5PqdcZYeGLNTuhY3ZG6SEdWHcMiLRD
BfIw3CTZ4/yBnI/G0/RS4ymRt58Y913mub+2o0jIDYXwtx0yyLWgpt0zd8xJG1AXBrtQ1ZN7Oe9v
RmCRIKal+Q3jROvUvR2efTukAwmRGFJiLkMWlTXO9XASCZyQVYUq8MxGglYbJfbyn+zteuIjrvwd
vZsxVb9GvuuWzL9olWhBj2sSMlV2igqLH631v0DzekHP7SsREiL8V1uxtoY3KlUGmHR/rfUNDBhY
kFr3vXAuALEzzg3jjeOyCtFK0Vp3rlZdiDjlXG7WqtB7Q8yCU9zShsFeTtcFps8rB9JbnPOwqljR
SuPvVMvJhdcFgywZ4tkC8rnotGLKWBJUAV+yvnnqwWxMeCg9MgbdND4KKj0ZSpBdmGYF0MpDaaf/
uA43oOtGgKhDwu85KoqAkxPmWWQCkl2z7goZVxQo1gt9IX11W8RZEIZloFFWe0vd+yR1qJ6kWnoN
ah99nqSJetqIqTYsNdgrEC1ewmsF0g+PGxQbVxSUbkg9Qe44H58J9pGnqsbux4cIr89Hm1ZOWAcw
z+pmN4o2kIJo5nQpLyJtkw4qURJLWftdV4bojaToCXMJcjdIghJ8FqsWg+2YwzrrPSwzZBP1JuZj
8gaNaj/zBwwwhpzmb/P54JA8H9JJqw5mms1K0jcRiNPkbn6RFZd44l0Nm9RHojS1dQAF4TTMcYxp
4LcmfOweE9+ZOrMb3o01zcBQOde8R6XAfcOB2fEH1wZKwyFw9sCBOV9nQxcGvswyFmHKrFI2sVO9
BHZyMXOrZxlX64laQS9zg8otOZHKx7F1jz+dJmRkuUh4CpfzwtDh1liJwHXUxAPrHugekQocVGe3
4qc6TupzZm8WdrEy8t07L5U4jU81h5RAwlJV1NP08i2ROm3ldYktxrJb/b57uGgFt52a777hVv4t
hOxXTVbPFwXijEPmeDHxctIKvwo1jALuuCe2tys/12X8YRThtMOLd6HcKRRDLgdf8kIXL8S2dQE+
ZBlPNcKH48XK537qoIPmtRMoeR5dD3Ra3dFTavSjcj2v5BcbyrkTeql+94TQeoed+LOi5E/29Skt
4nV4vb9lsQuYaMITxSp6iK9ubpQOyzo9yfEgEvcAQ7Xcq0dYcNYSpEplT4870BXEl2/m8tGDEaM+
vagvHZby1/QCcgDJgg2t+RaHaKHNkywmPvwOckXsiMgVkh3C+JrjweI5O0dMRaAKBVzsTNNzT20F
nF7Jr0dX1r7OrVAygbd7mKg2dO26OOR8B1QO7es8J/9iFfLDkCcS1kLc0PT6Uv7r6hH/wAwb1jgn
a8jZgJkRBABmczii3J0y4EV24W7FrvPfuKIcGk3H1eVEpH25aKRj7RzffkbMK8/t5Ik4ZMHrfyik
gOud8JS7H5VLzhELq91TS02nkd2AR9d+nD9yy70fgO0TUEhevmIdNxjapMAVj17CSsab6Y+9fyoT
5dvf7T/zQGYOa8QJY0OaoTLHoIfqMGE1h7hi/51SOl9FluB1vcjiHn1aeoywlYFh1l+hNGnqa2/t
SOB2PqqoJa+ii+m3/YFBdE6iyODu+8kMnBw14TAV/bNBUMa78QT4hEDSiPhdI2rzkCh+0bIO3cdL
dMrTvt+ofVhiztrehfOyKdB5FLbgopiyxBnoUeU9BwsFz50lSCHUGA6ABVEC59Xaztte6GhadVqm
4OvyTU9nOafK4dcDdNzCDtedzlK2IIjkY6OYANCUU20BLC8LDXox5JFUuNPKN6Z6gOWLBc/Hsb9p
PjutgYmCvGyNEGO2X/MvGq+C+1ZBBKAYUHV4dMnT1XdPxUShBif81wFKuz2tBx8sZEPhrR5xyh7x
opbhRQCY0ueZB1VZzboap5pFXRiQRM29UqCi77evbNiiMhEMFKfcwuh7Oj885wN3Yrx5Qf05iuvW
Z8m/AngrtQXkuolisz5XycnQb5jk09gibvLKmJHmorgvjOrQYRuZBT3DCtZbzrHm8PYGAvqKy+Yi
8ZsVt+rYfr6Ys0DaYeoq0em36US4W0qjO/IPO0Bw9UXbm5Al1OI0Y7FOaZmn7/kBB1Olq3XjfrGK
pFzsn/bFV7JxV13NilVJ73dGbuBuRIaFCGWfLdzMQ0jczxIu7RNvwgF8SLKEWAytAIrCEi2F+Cxj
+NecRBF/S/uRi8ghpPvUILv6xw1HXvqNNpcqM2gdWWObF9lScnI8Viw9H/RiWqjbKI+KY5N88Xzc
mZ8iiMJIHUypCpFbP0/fsVze/xqoxveZzpS73hDuCSIw4nwB42CbjDSCY79f0Lr0MMU6ZC491a1j
74hfJ149LwLyG5TAflZWrJqAB8LQRNXujw8B3JA/eoKDKndZcWQoyFBaMufODeLEh0uUJv42nvlg
Udn1IBhaFZnG4tlf3QlijpI/7t5RTb0SU5XjVB7nMHdEacOtX233ppjvHR1/xK9KNBpCKscCCaTD
AjVwG9GXCUm3SW5X1k3jWG+vMJb+KtYiPOwUshPl15D8klrKaS69Cw7ymv3MfLSXUEZXApvAGm0N
MlxoGfaDRCuSf2W78D61qyd7yLtXCkrbjDTbTr229Edp7YLCF53SoWuSFq+Ly8CTK/MCaboNYeBB
7D1U8GDo9sqh9MBlvMUA9/L6FLDKR2RsjD2U0s4cHI72X02tJ2P2VwyW+7Hf8mSTh7N+c3y10xil
Q5CjsFyiHRjLlBPHR0OR93bHOyf83t9abXxwDgQLuztYTgUGLpaMERIjn4+axztqmYcmSamzvlu/
qoLOlHFC+YRxsJzXMN2kJzFiDq3hw5f9xb6qpwGRUADKNSavPK+NvbneEjM/OSSbITPiQRBMGO6y
FwCYbg7fql0oYXeuYKtFEyK9u95Oj5CCa25x/wY1yFRZkqu2iBY5eLe2r/lYss4EPYI6mIUphfKN
HGV9dyXTWs+v4eQYe2k3TC/EvGKkGvbyvnHoXGZR+NuNnjD3fwq/qvlKJTBX2byD4wDEGi6l4rOV
mkaf3JT1lwDlFSoh0rQ3NqSr5uDohW4aD7HmxAxA/bmXu+fF6G8s70aloTy0odyPsaN5doI/xK7v
MzBoiRSMx5Sz4GJHIERAmIW3ELX4L+iivVdEXS02lSPXFUW9qaK/Kr2PoH0DRDEOn9zuCNJ5xG7u
feP8y7MGySQRE58U4fqfxYsUzcRqOJz1X30QGmIjFr1c2NKHPqW5ygbuonPqcWAUn5Y0ZyQmnQPL
CbQf5g0BR+o1NoRJwTcKR+kfdnF3h3bkCXmqQ/nHTEzWJqF0b+eou59o6Bh0re/xTqEaYgGWqpMo
i0SUgV2DM49lRY9tgiR/hdcR5fRNSf4jVUvpqplrkU22dD7XYuv26jGZe+Nzvi90R6nGJLmUwwbg
ldnvBVnEuigZSRLp7BVniylPpsKUCab/2lp9wyg9tAHwxavE326Gd8KT+wXuvk15RWiTTzdtSw4T
XptfjlehXdBtB4JUtL0LWvtSl7Tx8XQ9Y5HXFTKcZErtUYMu4+MZhbJa4pSsC9n4HPcYvWKiQbTw
bmMg3lqeskvpjHNHXrQWaXv03d29iSgywBFtK3ckOwYCNPeJdO4FLPJ37Phgzw4x/0ShPsiDA3Pk
9FUe4INUVkrmUSe3c9FvvukNkkWwFTauAdEsRMwcO7mEiPqodjdrO7zBcbwg1w1g8EABFfaZKKw6
TaWNZ6ZQ91bBXDeQM9ILOiugIUSbaFi7TVBMx5ERZZidxYUWk8sqKq6gTd15I6YtOcNaF5ZveOmf
WugyVRJ9iO7s5+6WNYKjuk0a+gj2OxbOTmwkjUwwGktvlbc4hCnmtXRlhalr4Jm6TZM1HOKRCpWZ
UtrwDnTalck8zEpZFb0/VxqqDVLZcVqOArPjegOlvBhpv5L+3iLZOZ85AJyLh0A8NWwJ7KCKXZZ6
TRapIFKz8GG4urS4lpZl23wMOXUfzeulLwXXgCIG4I/8O24zpMFuBA1jx4xm0IU7mrgHYvuvjFK5
Hga0vPRRtUnS/f60QoFvx+urbimz744hoaSGeV4wJV7XUH58KqBvDC9wtgxjqhbgw4kxhiRiMDtN
Xf6I1rtl7Urkgv60FGS9o5OVa66CdHZTnSTbaeZhRWh3jCQn1im4ufP7oiuYrVRxWCDuJLAtSOle
Vg40F4UDM81inOiWYtKZrMWyNAk0Ms7Y/0ZhtmLqH+AFMwuvkrLWGIilCKAlMYu8tnmNgrV6/JTL
Dm1KhY95BOumpyqJlQTM4vv0u3ka1GKM76W3cNPZvJaYUhhNL+qn+uIQByJMSY7tVn981or7gF/m
cX+DS392xGxA51r35DFjpV06asEr65u+crOlpCqdU6iqKbQF/qc5M897Efeb4SLkAVLely742X3/
JQTjyH1utiPn1jX3SNVJCFwOMWddoDhBcyKjv6nAZ+w+dmZUkBwAAN0POxUsxjHGIJfkO8osWJx+
dJDEv96bZNgwjQZOtKTrf43QHc/mPwRqvIONz3Jp4+1t7xuDq0/t5MMF/GPWPPqd7xBKlgxE9+bJ
acA3h45G0OXDgA9rOWGXASZ2n6McV7cFjIAVSm7sL9p4aCuyGNw7PzYbBH/pFM690gM5rRjgplwa
cdZjx8B+QN/n1YiT760h4bw6QAtGZcChfl/1s7z/VvDeyINcWOkWcCCKssdBGpZSctdMHQLLMSrw
TGDUzpHEPsBR8CWqCtigdZ0a+FUSK0Mav4j1+JnOMAMTyPe7IwjsXgt7mqQr/s+qhRILnR+13Hah
LvSkh/2/1g7iwWNhAXDFEca4G3MD7j0qyZhxEXOOkHSTDlnfA06OyDv/xDbEzY3Ov+NKMJlPnxLG
a4XbIPBGT4OrY7ePJL/Wub0HX0BDBzgDJnkXoFc/FnZwmq3W5etlXDLbZE+ISp8aQuZHrBm4SSLx
JbZud7CVJ5vKojFVtr3Dc+T/EdtvCCpSSj63jwlZDLP7BQCU4nZ3AXUU4XMvd6rRbY8eo15HzHlR
aB9IXq72MEjXp506/tK0RuClesJDyFpdlFx70+VqWRXKNz4qalAkATpzBEBmoe/jGh0QHl4zCvAz
HWXMS7+TH8cgRiOl5SqKp7AwJbvlbMriQVwY8RbZ7pd7FiFG+25/sKhPsLGyRHWNQdTJLtyG1hiF
f6PKKJLTXhAOxAKmHy/kDJTzdx4spTTobAyV6v8CKG+9fNcGwij1jDmXSjWJ+rfF4XYCoT+cWmKG
S2txCc+uDengzVWoTeaHjaffbKt/ICiIZ172iR/LtGeDABLBO7FcC9necqCAVpbrJVMikV98PS2+
3YoIxBsMkI+C/dcxIvmu1afgr10IKBGmpKU3uxX2JS1f71ZXWisMdN+eZnmhALjsZpd1QoviCYRz
InqKwOFo6ng7vsbZ3/W0rxLXr1QEboMBmFm57raMWolFTO6DCp710aNxEzzBrZi8FiUY4yBUONa+
2l2VidluyLffP9KATGDY4Gqykul7eEDGVvF+IP3pOoIyTJ5x7/KXShw6GZbRVedLYdVySSJMUDDQ
9+01gtTzUxQ0cXIuyGJbGyiPpwQqViEoyRw4UOErZCmGs4gSLmz81bfgYTcmKhdzLiyOTUHU3HUM
3jF77YmQeWVqyQU7Hq2/xsx+AmfxQrkjABSWqFdA0KD2WOzWZSp4ZDwnHZaTgDHevP1g2rKx1/PA
qXh7YomWKZL7ikkMSYS+z8qHeDuwNJN63uhekO0RBArdipFmhD1CQMFaVtGvpiQTsHsEF45U7oZV
QwuDA+kk3IgT5cyHHjq4FXIkAhBhtY8a6kWqGf6Op55TUXdY6Ah7dKAPVStZP1RR1k8cSapH+OHb
/uYtt7Ad7nWUVXuDwN9KZbn32qqUGWPidLFq9MIoTivPSHkLs3wN7VteG+LRac/O+ko9sj2/5HlE
froEIIBj+A72hKA5mSeQZ6TeRqNjhPzodDzYQ3z5n7xHkx+2iA8L/0HKQ0Fn+uaf6twXtu5M6UO9
bcwTMO2Evlyz947BS0tBYAhubSCjZC1Sh73dx7R4bjZkXxDFI3fFUoC1+3Fi/CDA54UJt8wz7cY7
WKHYJjKarP4v8WOF7Jt38AvjVCNVQrlb5EKTakrTvJSO0ceD85XWeWNaKSx4LVG2pEoXq0hqsruF
rkpW4KKTwQE19eZKhh6ZqLJNSjJqkDwczKIoMlYZxqFodkohq1Ibg99paZd39vDR01Rii6y/g60t
8xqGQUNb0es2Uyb8MDFE69Rl0YYytDp8DC52sB2JxrUD6ncVWoZ2xMYTCtYw3RvBUideG7K41K7h
07IV4aZOC4/qlVO0npEwX3YosCpiCTIHR8vfDaPgHbAIT+6PxjHhSlCvdbX6XCrv3UsfDYc0+Hva
R2yUwcC1RD3M1QgSuIJRzSdQRUZvYg81ZYKOV/kLSLOP0u7pZU3bbwuTeSA7CQj6SPsrlWDc7VVz
CfGuRTCvN7aOs9VvGyc6N0SUxeNNJ5Qsp0/m6MDmvnhYHhUFGVvf2TF3R7q4KYmYXmSHxYIBV2Lx
mtz6OaEatZyMj7XxMM9h6xSGjnZ4RcSVdlIUmLwSsgfmPRgRnUJUpnHx0K4gm3UTlmYKAK1Jv8HV
iz1gpmp60aq/H8bwNlW5OMD+Lgt8h2jdapXwlZ2RK0960PYH1NQM91ETC0uj4RKhFTXIkTy7Nrln
vJkNOXrJKzRbK3E2yiqrATXUUK1krPwuY7jDrgYxfyV9y8GLgoXWrDYU3KO3BK+P1lD4ZfUOH9px
VArmX2Y33o4bfpl2f2NEdaNI0Tx4QF1sH5zzdQLb9Ysp9rLaEC2qUfs2IxONriOvez/TYP49n+ut
WQDNe36VbA+CGeHY9KcStuterirl9yoeoYuFa02UZQdcLOFH0Qfoj7TxYHvSD2W5rPIPEJ63jqkp
JUx41smi25oNmZ4Tb4e7sYurhgMNZUY+OhhuZ0+6Xtu8Z0ZTY2Nj+8HvBtmjLHDYKReiMO3Cje+F
g9JG0LENbH83zCT0W+AK/6YVIgCscMOZontdOqn3YzTJPnFHZfzuAVT7ld5Z3moMR5v+h2dIAQY+
N4HChMDmXu9uvCZPU1n/QRKZC/RGQvtHAef5YPsaiGRhVxgvdUFJgvbp0sMMWihVJHmemV2eERit
drCwEVhXahbFFGm9wzy9L0gLMiWuzgoleEDrGfe9f5s3Fkc4GNKAV3dEyhE7A59wS0r6oaMAbD3u
7Fuly1zSLa9P56Hg6UZl83ZPOIsSm7IHOhi0FzAcW7lS7Z1rrdQHYJhROEfDHT99ON+dL8JRGMQB
9KP9ECw15BfxaHgIW9JwSD+zKK0ZJ70+JIyFYQr+/GMvwc2Lj+rxTYzFCmWvZM92bcEAvuylfCQk
CNHQ929ebMvO/VVt6MAR66UuWMVtzkPLmiW2z6yEeYLvMGmM8sBD4CORdyWPAPluufs+s6ISYGIe
2a8JWwbW1yKH4pbQ1aGTC3dFzfqGcB+MGA/8KT7+hdh0WstKM15WWwUqwqgG9nhlgQc8KVSLtCer
GKLIO9pmS1TIcZV3zStPQtGqigmQvz+HdC9Lpb8JA3K4SYLwJ0QCS0t83Kxm9+RGh95IrSclXOp8
ljuM8NYJwHtenJ12w7bdtZ/r0ICGSeSfNSY1jN+hBp6hR7sPfCiXGp2JMVa7d58lUgUuY/QiBVHy
YIOxHoiCZD2uqlkr+LAWgvcqJr04Q0FzVdwhcbe5ZRxG5hAPbHbk9NDjkmpScG5dB9G61b3XXyL4
xAG0xC+GtVbnaiKQIn1VIFPuMAJNL5NTmEhKF84Cf0GdM2BOH+Kjpn+nW68TN7uMXCbw3Z/bYxuw
mvAMXXfOe8h31kKMz2PvFDSd0Ds9E4Sv/uPqUM2Zqyiu0k9hB+1oejeL9YIlvjVXHtKVsAwDGPCz
G0vBiCY6w7eqty3NpfB1TkN7oWLLcCLFs+rzn2EzA3BkkoLlc0aLxm5lHaDXAjhStxzlZSSAmSH8
mOlvooWH0RpFNKHIJxE170ObZLMoW4IvaQ2J2TLbCt4WpfjOpwg2XwyS/ITuPB2yJuwhiJYQ8kW9
FrjNAl9Kw8V5t6+izzO3Ctf73VDuXAnOsK4Lypls2s9EoleBpMy1PNyCUGBbRGLcAcKQaXUr9v8p
GZeXD8LL9Ft79gqGzQC2gALicqzJ1IqwQDQayu4vbmx3rVeHKgVCF0DaB5H0yY1WW1utwkiORy4n
PdCOvGiU+lgpaGOIcKkxjIqR0z1x48zX+tLqESDUedzfY0YXwIM+WXS7PpDn19I4y7mPRzU5pPQI
SfqXUS5PnPa9mTpQ+m6JGmfYHed0Fj4xVPhf0PCgxYrKno0J16eYWA73uj3OYZ1nrVr8OniXmGGO
P2dB6p48mrPNGxBbU1rLziifSNAjUAg8dCqnuuYkQ9Dtf5U0d0Kd83DQHIqpsLaF4O5uwnPTcWoc
FaufuMwg9DcoJzvUpPVEqHhNf2qgihT3atnMgTA7KAATSTqE26bC2Aiy1HF1mPzgG3yKmqlloiOV
yzGk0c/mvKqzLTJPprUcT3p8vGT8TwNE2LR1vydD+/GX4OBnzC/5hcQAMTg8f0UNcftkmOs1qOKz
7oXIA8/CPyWV+8d9NAlIYQjy0nKS1RXt7UdX9rvsME7zBS9f3TK3Jj7Ht7Z5xR6AJD1j2hVWpzVS
CKSdqz/lc4KoImnJM/+UJobLMvvtmD8juaIF6UI2C7ICuMNaDG7dPUPyRm36X4J3pFWpn8d6/Y+o
RR0duDBA6kAQj465aHESi5TkRiaBouDQcMIzZoz2BnZcf9BKS7nbqbcCakOXNcr4t3bNmnCv5YkK
Iyf0io219CCm/zIYgBpon2qsII2cJSnRKQlKJQJ+H9yJ1mFE/ARMoSoecTUp0woPvly4T+BBdJBW
iutbZcmHDGw7/lOGAnjGZvwyHOtziTQGurArv8pKAOwOusNVQOjGEkvZX10E36T0zHOq2ON5U+Oy
zHlesZ4iLNdYl9nn6LV1IEzMZjYlCirxq+jRu5INjfX/spwpE6C6rWCjDctBSRT61N1/olTcDk+V
BqosX13XU11Oib8rrXT6pRC4Lu/Woq388rvE8crsk0DONrRa06dVBNndrbdxRpUwj2kvgMp9wycH
6SQBaSNdSORCt8OGrJg481JVXRYG16KYDZ9VUECDEQzwh2SO86fGp5Ot8OxO1Mua8NK6cGUGrGjA
iEcYdv/DxCUiKVj4qvLkcFkaFMkMkxyNgK1nFeOfL8QNJhw8235dtI3b7urlNoCeH2VfncQ1K0OH
msGv0Oj4MuGbMB1nWhwy35UVKjpVeXekcjUI+sP+hQzeSP27KGHepgaLnpegytbsULjGYue0Y/Uo
/JrQ10WQfTDIjWCL/vwTTnJMAVcevVYlH0cTLM6uTHLfVa2q9cCtx3h3zjlKQPFxSiop+9+REjXv
CE0rtx4+uZG/u6uybud2PYl8UbUZ1BYBi46efWsRIZmBJRYCSW1J6XCepBatltPWWgUxTnwlIiIe
IdlIStekdWl0/3OrMgRfM8m0haB2Y7JpagiNufyt8+nfRYLgkAwie/rZf4QL+DZd6zyRZg+vq0JG
JF79mLvAPWvM786FOBm5Obc19goQCPmXmChYufNTOXLDufTdoT3G++6TOCWqVlNmBKfhJSLx38vN
1kDNbe2bDmf8Z5avp14HGTbQ77/PNlhlXINy1480b0QC/utcaMkVN7JGwz2hwYtQGYBzxRhSY8av
BankkEyTuy1pGwkKkSWI/AqfjMN92zSR7sr2uYCb9TgJLxmAnhri7boBGNxnsS4O+Hdr4ABTxiWx
y6ovCclVZ27X6ao6H1+6bosyvjXqVhC1NBO2SxEwT9L9+H+inTuBuFZgBvA6xpUIiZHKBqL0jG8v
A5trzwHuDZuurJ+RIr8fKz+r2zi5gB1r6bpdNcvgAHjbWpTYmZkjZjCnqiWY4p/o3202LVQeR8ML
qeNlhxko/dPi93jztSc2TyDQTbF/6saiWQNutpWyFuY8mq5EmP90JY/5nIdLY4oE9VMr+Qsg0SBw
aRCB8m9AyRLxdygruUcw0Bq12XFVVCBJp1U03mppEIXesV3cSaHPpIH0JV6r/0cDEXw0XFVvj2NW
W0ffjDj9TAnYmEeUWoSlk08FCasN1u+mFtXbmAOv4syQZfQ5NFJ7uO7jyKWzUPD8wABlnyhHrsBi
Co5Chub2STxy3njyLWtm2u6AR9sJZ5idIMEp/jEqfFUHeDar9drIydeeSjhEnYKplke7vdWPI5r7
2B6BfthcSh2JydZZKwin8UWdO7+l/0AIVeoVIq/xcShSzeflNo7xNpCYsLHdBFOFCOIp7tf7SSNp
JJWidUAYwCrKAs3EPKCTJn9hB4KJTQh2aYxfSHGiYnvGGGNBBXRKW5lbuJC+TjLUn4+FnhNxNzqu
F+JK/RwO1192qq2UK7zg2TrYcQs2OijqpUlbe+SSDJzuPWn+6kzHGOwHVt3WoaMD1ZeelaTSvbH7
UfCUvbtIAMjobxGdscMZK3p+HVppd6r9k/CyXwk6XoAx15+ZsVcMYvnCKE27524Hokpg03VwPFVf
Asx4t7KUcHqFpzcKRIcrTq9t3zKq5ql7DHXDLZDceDWfG5pyL6xJ2eBkGHEuSGSWb9o/yo2ls7LI
obHw0IpTM9Ew25L8/H/AHAeRRMrpFF2HVYdTffPIb+KieqpEQC6QfPO1kOzRxskaCqCGK5uVDyxT
1obyY96lGIeI+RnjwUK4D9caU+aoJrHuTu88EA/asYA/64t+/kb5nua6L4d41y05am+Y0JFzRYRP
dGt5bSGYJp+kGewKmWwbkt/PSfaVnVUC+mT3pzdCqQ6WI1J3I4wiX3do9VRCOc0VbscVW5Iy1W0o
JLXYtvMqPy1wKit7SbZIJMvR5hF/XuB6vEQmnCPF8hiYRZC5uLvquPpiYHyJIxRbAYAHtIokmOOu
sImOqMZ49zQGhySESKAB5+Z/ahYRpPR3miJspTpuffESMrZJHSgoj2bm3lfY4R4UGIPeRZJe5onv
/eyFnvrL30k4R6utRGsISaYNJ12acnXE7SP/kxZ2Y9vDGeFYheUCcgWfF2IaLh6J/czWIHAeYCsT
APPaK19P08eXMHTG09lkBzpvR9w97zkdQOkz+qzqtp0B/Fhdph7tYPQsN2ozK8qxpUeKKRm/m/a9
UynMU/OFgzhzzcjIGID8JXYeuIOlzOKHDQc5A+buenl4oW1ff283EohAnX2O4U2wNN+NlRPFeTvr
KH1ZFjbcwBbLT3IGGz5bedwI5qke4am2ZTJK3wBMmYYzB+qrFNtPNwKnxnqZWQQpGg7Lde5xmhhf
Wq6nObrgXfcK4fqkp0DGkpD+7GUBNeKF0tJcJB2RhK6DX6DNXsLoOpukEn87PpnpUV/iU34jjf8y
kmwDVbtRZ5SLJF5J28ltMeIMgxz6y0Yr2gmFkRZ1RC7G1MeTD0V6Dl8ipu4B8H8HFCDO6kxDIwEk
za4WZ1IjQjhN03KhIUt2jLGi40YbxD0g5KeBZk70UqJtM874mU6bi1hUKnWD82GmID2R6OGPEn93
+UUsi/T9oy8VgRQzGeAS7RqzCVO6hNyqJ/Mmtf3qA/GQvL7aKSdlAomyvJxSAwcjqyuomHwKYSyt
guWFTzGj0OCRofKmCD80k865qyWNPZCZzPgfN1VFoRIhBTJI84CENiLLky0ibk05MJQ+BRMxfrKL
uvRNIQBc/PC+9GH7fsVN1PiSmr5X0fW2elMS9YuXa7l22ai88ISLlXshh+WfQVK64b99MCodJxfc
23GjgZ0p+3U2Tgb629xucjmKU16rYdrnZYnxn4cn+tk7kqtIDV+aKYrH52GWygaNDGFHNCFEzC+b
+yapvOcoJagRSeL6MyWpXc8/cYNSrli9Rj+jPxcZ22sBl96IJKlBkn11lF5plZwMgAmfpCKxXgTJ
sMwiw9w7p0v69+9I3gVZW+aqzzTNp3c2GiL3XdOOoTdQbRyW21jnnZdiLt95jJ+HRcUQ/OK+rsJn
B2ZnVunsPopFbhLpM7cWORznt6pA0gYYcEXNEsz8oQu22j9F1P5ft7eZ4m2WNp+UuLFOmBRiXzcZ
cDi4AfHJ/9hTDoAcpXBC9VbPhDGEOaqKPmeV1VcV9rNi4g47+3e/Jvk0rHxOh7LyroW6Ev5pMzyB
PhLz/q+TNl6U/CnEFEE1GW9SDa3/BZPpwHL69db95UZxx1GTzejg54WUCDg9L+svQIdjAc4J/mVG
eqH8sA6uu5DuMUnjJV4Ql0VTmPu65q0eNBDIPb6qH0Su2k2M7tDzEZJZc6FlQeIlQH5/SAMcsGsn
LTqr/QDSvKk4C9s/eRFncaREy3K7ay0dOfMTRgok1WxW39MpJXO7bj11FcqIdbNzF6HeemksUT0l
nnCCHIKaHjBlHZLtd1oQb3Lwrd4VOSq4xTVGWXMzvdJ+/2V/M/JIiVIk6iKf42ezytQc4lBZZmKC
Pc3jXnzVIpjrBzI6C9nvtr+Us6DSvf3y3lE2+NhlNvhzTq4o0Wjd6Yzge43qy4AmYAqr2kW5/uSk
CjD/kmiv5q7m13/FaS+DvRBRdRIsNTSv8EHQAzvaeWQRVebpdnN2VFdyY5GoIETdOKtaFY/Ouig7
e+gPqB3oIKgenEOs1UQq/NEgBuZe9G2yQv8hrlfluGLHGGPKQJNBe7rceYslRjE7yNoHo/fDCAhk
MeuZf4ELh3yB3pK6+9+fw/Xqtq65fdAffPxuYmPKaaLtczLkAjpLQ1AvRWhqDQCui7mJM8Dnzo6C
fG1EIgs08p8AlyLmyOkqBoqsB6fCxgpyrNEvglL8OFjuevxNRWejDoArqkg8f5G6VpZMMd/myxW2
4OeAc2cEl8DhnfJ8WdokV+h2Kj+ZzGFwGSdMQG0tiV3b6OuMTfGrcOfF7rpKWaUkmAtaZfg6YGgH
56gpl0rovPD89i6/b6U/zAuUo291sJ/Vx04RTgQjj5sivL198dcQLgtL0ho75xtTTLCPJ2fTcDwH
nw5RM/8Mj6M7tf3MnrW7HhnCJiFoK/uRXE9M/AS1Bcohr+GDPn3rcS+K3bCu7BxIuYIYhB0QU/tb
AzBGWSZYrGsMGrtSk/+ytEa6+dD1BJnDU+y4wIPFCD6p6qyOZfSyF4iJR1PKkvCawULIZBFVQm2Z
bGHpHxhWQlsx0QKwqNTLfla0xSI+9N85/61g7cicIXhLoUvdcJwIBGSurUUW/mUjwYAqrXDNvs2w
cO6KVBDnVedt2UWJFja1nj4fyX48FjOjD3sKuR52xsAHndxbC0rCQCysJyeIeusCqlPICzAt1K/e
GcYKvcf8+Aju8DuZJJ2I000Mb5mRqJD347Zjo2uwChlQ/SXQc3ehD/MPNF9w/cl71vDgZvcc2Fex
Hkyuu1pyiZWcbzOHBhP3QJpmorHGPkUECIBSMI3t9YWnhqs7mEPl5C6SsfIkMe9eODl3fmYFvsoj
rcHq9D7ryrXj/5AJznF8EHhEmuGjWqmhxtB398sUPvKzJ8OflLfzgiFDk4uKaP75RwFPY2Pyg1gn
I5PwUuH+35b3PxeTz7xYQTBa3PlDeddY64NgvSQCBu2KGFjKS7W9Kq+8MdKvZj0lySfUM+q2loN/
Q0yY8bVxVpL0Fcgg+2ykh76np6SEDgnUkY6QR2KFi1pGfxpE9JivwDnV5L3oG2y6X11TfEXCogrU
AvXMphtCrLhPvjDAA2tOx4rnuE77L6pchrgrsoYjRffoArnAdIedRClcSVTVltkNsv+xDBNo2uAg
SVpIY0hwxLcEEJkuQcMsyuDMm7sUzBi0WoziTUBxY3/XGsVEHdNVh7pjyo15xK7s8SZ6HJFGa/tU
3+Z7ic8JHLR8tANeK54sr7JG9ByFuOosutTZWZSkFx7Xu9L+N19aToPENII/2pUOAk9W1IQ0J+CT
q5Xo0aGiRMFcAZv/svqv7UlEkr7CAt6uxVxWhaMW5jYHEQRGOGQnvdjPDiu1e0i5SNvmNaty9R5A
rYxTRLNz5anvjvtUx0ZUbHrpxyZSHQbhVdOMjZR3+VJhBhQtuMtXggv3irDNAJ9su70QT9CDNL+V
3JrcCcq9rmfk2Uy8NZPsrpc3trqrReiykN3YnrTFrpD2nrx1OCjjzSb3HahJtXHBcoik1i8jVnhT
Ljw7RMGwmLIBrbz6Rg68aW+g3yMbK8+20ck/jgmiDmgDb+VvcgIHkX6mMulxrZVndIXStj9aPt8O
u91c0K/z2qgy52QqBO2/2EmRibIhRbfSTvwvV8o7xTo/xjm1Z/ghHU+Zr8ZQMQcU2YRv+Iu9qAwg
kMCvi0agA8sHzMgjr8+Dq/0VsUxkszL6zmsO5EN9NgzUX26bkzFuRo5xSKbby8OpKDF4/ZLj6EVG
1TqyZSCbf2e/ZjBbuGsJAkp2PLW7rboVW9/gqj0c6jVbGHDIVKo7x7GJsHsSnhRpvcAFFNQ3CAj/
CJzuOQzjDi7rq+6KX/r0Iy3SjIl5HnIReNQcLFwF1g/f5Y9TEskerASGDKTbkUiMfDlkp55F19i9
uziBgOk2ncLWwYwnnyfytu2PUKq843F5Faw9NAOAcWxVod2BeAfXk2CSSUzbcb554GgYrEqoTRZ/
4YKrxEbiIx3e8PuFLNn3QQIsFzuyuPfiico2YTjNvcquollF6WyWrLSQiNOeZWTiDnWoqh/IjvU5
YMdOQBfQfK0x4/NFz9JVCtpJl8gHK/u5Cr4pIYD+6XQf0/eQv5wMofOFoy+Q2nSkZQr9Z+UQDosn
3EukOEcxfGg+Ohilw/WkY1HXe53+aV31tQtDqm1CytVWT8xcLMe60ZysC/Y1GqnjKR6Rmx6ooTaF
DNR3t7Y3tP9bDt5YL7g9HhY0eEdvIfqR38eiNO8EVJJ+2ynaQ0Wgz1n0pjQKNIBPfrc8ygZ6tDWO
id1gXNjNTugxfsXm5t9KkMVaNV1+g2CtiSVpvD9vqohbRwTMbxl/TqRZYDEzpGaHQdmdgnQRGOqa
OcPTMrW3ALRwMJdk1AJAuVsxbwCbx77R8oecWGnAgDT8OxDgJppsejjFwsoQaR1Gu4fG/FFYkRzL
loeR+ZTRli1iHH231unoddKRWqX910NKzSIwNyYHxX0+raNTtPWks/EqS1AuT2nzu74dDWuOOBZI
bG0ovrtAZMXr7KBvWrfxcXSpTWc/P5GxzuKyrjYMpj5faheHqQEjJVUfVP+qlPGSSwH9dN9e8/VA
Eo9VkY7uY8SJOEUVmMii0lCIx9ptzjnZ0xtLfXq1nxkqrVzy0o9FEVWnFseCKxAd6cC9u+goEEhy
OT4lnKVb8AyiEgFFU42wprsVj8o5weIXKHFXxzKZ9imudZlOtmOhDiIJWdAOziEWNqPOaOAAFoEK
ig4kj+yfCCqGD8CaOwLhehwrofSP0q6vaYiEKnn8lDPO4zOqee04FWbctVqCfiQ4IGH6uPvH2Pks
rvaYAkX4bEY664xxy6dOYoBrR7embPgq1S1bjzsQFgS2ttN+R1ookSfypteDmxjB8oXi1/qqItPc
SmoD5Vo3l8RzSzCYLFX7GoECYIt2GwYmVqjC62HuKEozN8hH7BWl/rym3VyMSrU5caFbzp43/HKY
5m7HpdzNc/bhpH1blTWD2PyltGvgSif2wmZ+fZMo77d/yMoiXrQyTyEGUBadCmW1RJZs7HeaAQAy
mtWxzDYddmjzwABQlNfEPRPfn44/ibTsGUuPMVrrWc/81Ia/QDpviSDJTpsYgi6D55T7wj6h6O2x
Q5RgjO3gAIw95OTdnZ/J6ilgFwR8lENlEUMagRputgDcH5jDnSzdeM4XdR74BC1lYnnOldBY6cWr
fmqTSXgVp7DJzwTSFwRoF44N3Hg8KhpD4VHdwOVk7InvXjsx6erBF8JnnE9ERMtkfMFeChD3evAg
HSL4YzPLMzImHUp8fFkm7OtZF6keIRMb0VObGW7D9hoaRCs8uJcaI4b9vewjwDtIepzCoVjM4hS2
VYccCWlmXg1CDfk+h9G4QKwlU/TCMHpjkVjUpm04wX9DkkC/xgHAUKUhiNLOS83k/g5HnYuVPiXZ
8ZKGqZs7b+0IyHaVpfiFLE+wCgVFb1FkO3I13/vfFxR5pFwqj8W8EX/NKlomKEf8kyT2OHZFFH0w
F9BdqUoPCy9/Zb4z5PHdvHnlyTuCxFovH0IDDpZEMphPUEvriFUyNUmmjzjOyixRj4mSRB0jj30B
8Y6goLdRpD9chqnFQLio42ck8ViPrbwLM+xsjlscAKpPR2NqhYLF+4JeYCjmItf9oXU0PS/hhk1c
GadpqCmfXvmZgzpoPhewlzmHYJph4OQOh5EQBAvzrKcm9q4rTWKwvoDITD7uZ70V15W1yfwv43cW
CfFKRQupNmvzwN8y1Rt+a9YSJTmiiYsgOzHrTIApLz6XGLNAJyOBhQvcRaZq5iDPc4y8VHbDlmZL
2QTMR6f0LT1fcBNkbB1MHEoFgy33K0geX+NPGZDwHaTRf1L/TOjwamGjrRCvVEUSHBQiP/mFfQEe
16X48JIvq48/T4/h+xKyjzbBmV22B7r5AUdCAGDrQPXo4Nw/rlZng3lcebzxFoKkUELEBQWp++TI
VynLIe/um599EuVpDagIdTuWMKZDqdzLYqT13IZnzRIR4LipuQRMLCXDcQvFOuRDxqyiiaAAV6qL
rCee64z0gEz0paTkzp0eSg9Mdsberqif2nrx1vOuqRQi6M/cxv9Wjeb4dyXBN6DAlodAreVEoHo3
Nk4qtP4XEm1bJpOzqTcoiOsHLw9QcXieW3MoAbdRAnsQhEDDUFG+cyuQGPwTTJAJ+ww2BdAx0NwD
sjiyqS4V/yZxQaD8WOqGYctJHqZpgrCIFIw+MuZJx8WNetZ7thzqckOgfpApRliTFA59KIrLqEnA
XpGWQ4KyaIMjY93O89SZBYgfGmZlJRAGfJHmwq2dtNCM6Tdjg5wiXaLSAWz5mmA7J7JEsQ2x1n00
Oug+IJUoCXufjY9p3484FoM8gKNkfyXFzc7xVX4EyfzEsUWe2U55WISpCw4NDLO+g+g6vaO/7a76
HIqWzLcYXIEmLH/KS8lMuE7ryEImUOD1L5v+VeWAgFh8ASoCoVP4m3FG+P9mU7xa6WtE1GyiSX1B
U9AF+ZVFX8XUQLf5WnASlwhrORDd4lFPKt9lqoSj5IIIMK4WAYkey8uvm+zU9fdxycuPYJWK1uVq
wJSrBrtlxXk77nQPGqeKQ7VcgihmAStDakrnUZr3k631KTAxd18Guk3qp6v/NdW0dbmYRfuQW6js
ROEogo5V+7a087gAZ+rcd8UJGhoDzQL08MKVVV/UdTg3G+X9EvWHoTef0mwLGJATOF8D1Qjr/Qrl
RTqIZcGjwv7MT+73+rleYJc6FNAv7EIIupfi6ojiolsBzPK7bcrVKGdGyjIG3xgQBAVGMQNezhoP
fiPTyagr+5eZwqVraLc2RA1Y7isO+ns47goibm4H8yzNbLLEJrm8NEEZzgZKLpmHi3q8cW6LnjzU
6ZBitc7fk9nSC2N9IMvX6l6D8AmYJhQWLihSFALeQMhYEdWw9jzKKkvWdsDnJKYIL545j9s5J/Yu
3oA9BxrGMt4y478KsAmqBdfIw/xcATWIEN4yc7xHLu6CmW5SnlNUSYIAqxoouA4KJv3R2C5TLa+y
FPliSvbLJrqtnklnBwaQ9ckbZa+R8K2w9G7rQO0VRUBKbIhcK6I2gagPvrdxnrEqHAzrHLWsw8v7
QqwjUUgGx051yZSkjjHeEtJ9hQyESMP5P80gQ++lUN6YJ08xhgeQzZmjL9e2k+N3o+g4W/XIUM+G
YTZ0iKTQxB7SHBTkkGHUz28l61q5Dbh2YpBtetPK9nq4TtLMIJmc5tG+ULgNamWBnXK4bC/D8I5D
hYhqBXNke5GSRTiba/T2rbPMy0lRjsDHpIzarhf077HWRme9xBWbrGSBsWMFxqlwMCl0ch/ertGE
8efEixGQ3YyTMzpBjzpZOj+9qKAt1x0fsIihyODrO/GDHoIEs9ZKRKkk/AUBNnE/T7aOwgnkMfsa
hMJQgRSXu7la4dwumuN2ThV9i/GQDuvNmV6JPoCI2AKhPOlFGAFKLvMgbSEovx0ztM4vPbdq+qDO
Q2C989twkPUpU2KEgA7tAycH+KJOpGHI9M9Evk1W3L1k+BcYm7AzUS8K+coF5fcAzI7M5yMLZuu6
F1Apw0vA4Fb6xkqxxxDiwPSfONhzLH4e1YostB01zfKVJmKBiIOcXoVss08N+x00D7kwymCdWQYY
B2ZF5aChsJCrxR2NW/dPhVValZ9eZ6nQupOVktUVkz+NmMmeMQGtPq40Qve4HdtQxffVHo2GsrAQ
ExIV9ggLcfgFbs5/9Aww4ClY5V50Ea7uuNopUUIEwYpg2VZaFO0vJXHYfsPYUmsdJYyNfP+8z12T
pPV1xUWH83Ex5cbAlK65w83s4fZBl0LTT0moy2GeIhyAY9HjuoHnqKtTR2PHTgGNlTEMNhTtuqtw
lyuzD85iwlBi3rVzBPndW6Th1H8wvCOXJNf/zea++Nw+VBhloFYEkq4PjQOY/By4FhSSN0wKwUKG
8HIpHTBw4lsAIP1YP8x6gIQPcNLutvbRqSYKiQWMjPaIImQ3Ycaowvwt4RAx5EOxBkMc1Hkk6iIa
gIjeLMDX5MfKE0KqlUjiCuFOv9EAw0PWSPT8EWaM6blePAE3IYPZaDfPSwHx44HZCkg6v2kLnlTz
5WHsamevG7AXzabdU1OA1p8Vrb+/cVHFxzGEm/qZoPtq/HTHwVwqXdoheNEvFkqLIxuKsgVDK0ZZ
DGw9AuJxCPfM8lQfC+GAuS+egFuPBwpBBDezcvnZhkhOiXxhwxooCh5o1AQzXXJ3pEsxRkKDgDZ6
fFXppPqQbxNBGcUuLeXJ74lfLPJz9quZXidPdzYiT2zbFRygaFD2Pw+Y/1TEnNbnfgPgOUP//UA3
Bs0ZTT90dGdLoQ79xd4dFqaryYfPhmw3TrB0jtjEZEy+muAQc2M9y6HLCU6ExTmN0Hm0Lo8Ybxcg
qhFPLjJSAhafPAEjuBqXKduP8bwEj5leKHzLOxISBYlPXKd2b+qf1h2fkmDeXbYfeHoaQYyeHkza
+Pat9iRXHGuZQbbOO6BUa6D0YgQJg/N8oaiWOT5hyPvokO3JFLAnKDKpDr37u6dAFkBUSV64BS/G
EhPBYtN1rW1NZace8Idvzz/67YClRZbKQFdEoumKF6Z9NPORxDm+V1xdfKUHDRtfridt69Al4UnJ
72zn/8b8YNLNvvYUf9dZdleMs0k+Y5jLGqY5VkIBJC6h/QmIOZK2TjWgzFohnds3Ebiy9E3qZLjY
pR77rTrVi5xtjv83TZeHzNI0XT4vEBmU1RZrjACsCA9XhCzSN0dAUmQJdAna3xL13ky0UraAfzZx
gFrcKO+pGysAPb6AearkXApjBiL/7Ep0dgzcXbShBhfFxahIx4NueRFdfmc/SEuKIVc21YwbdBVp
kC86BqJGh8E1xNUg70BTCnaDZsHzJVn55cEkZ8vA0zc9G+kxJHz7wfIUs5U70efa3hPLBnQMavx9
+3cuiPwAEgDsOdGIleVr+Taas9MhHs2smbhmy/XQTuvbjSJvdGCyFOvNlcm4fLpMTLwa87BKZ5uF
52E3TuPUGSGOnPNXabY88jVnuIjKdT+wcC6LFtk4vVuqLkTgls5AVNirvH/OkgM7Fn7W9keOMyr4
OvGcaRwtZr/s/TLyhorZcvI4Ed0/f7ykMim72Cs1v1tpiIktBaScewIYILOA7GGqFbkHjWcj8aVf
xUEqYGBOHtNetR5TnrAU8jOAExmfgrcv65FYCrh0WPELVvfW7A3V1ciLpbpmpQF9GRIbkfVDeAB3
pwuSpQPHCBO9VV4cjnQp4yUWABnFLAkeBYDH2E97uCC+7YzrZsq5s7fnPa7945AjFb3uVari+CGf
/j/MYA540XpXzGeTt/ibwRYaKqfukscJA0Fb3xIP+UXJG7BTkzwSCMWh3o2jpUlejEcMYWLLZ657
KxtaA59Wwv3f80Qe9y5CPpRIRh/KnR6DwF/UoPRsDqMv0IK3afLO7ozh4MfwfORXKPx06UInZFN7
Do9IImhnsS7tIt3NB+PQCXbs4AwIpwzo8MY/I+rUpnbA6Cti1rkxkzii2ULu2WtwdJSD3XA/zT2R
HP84jmWxnYoViLTyyOCzjctlUJWxn8BQWZ2Rb0AMG/Lzo0HJYcvhLpYpP0Rp4iS4eEZNLi/0KYfR
qYqTWVxGhj5nfXsH2RcUI8AvIosJHPsXpcHkpoC2C6H8HrufOhTOF04kY7mfSlcYKp87MBJ5T+sF
LM4BG+fD1QfV4a1UUZE6U5co4d5/JOovC8M7mMqxleCVPArSJF03gWg4MXrPeGklUWEJU8t9a2BM
jsi612W2yrxi7kaUDrgWLCaGK/p6d9/D5x+wQpVnJhrKrAlEZ1+v07L8QM5BMC/odxz1MHu4PCFf
5ss7VLEEQf5fLi87e5uUHSypHpvctdxCNInoSqOHfSTgIStdbndFr89pxzsi48qmrahxR3UraZUI
tD3KlzgkytJtl2we0Y0H5be8AfQoA7Bm+CPmli40ZVM4CUKi9c+herCPBym8MUGZuSzdta11H3nl
2X9DNAe+Pd+ieG9/Q1s1U28vmckFFfWh7GNGru7o3C7paRF/MDl8TSZBZEGK0HUKIiQ54EHposoB
1xEvCOm0KkfC1psuvI4s229gFq0C+UwbojWW67mFUlMIr3WscOSaXpBI6830OieKP4uBYF9NrHbg
BDTvsRoer7ywhZ5+ZM+6gJQl97eP3Jgp+Ig9sp6s66Z+j7MVm6o3CBS9VOYanHWu9h+uiWqglML0
7nLQ01wfQZCVWyIGamB5pF5fr+Q2CwO9kSWsLMGHClSjZwUzs3PqpeLGCBUdEnSNSEW1yZX9FZpc
eYghRR5+0nX25DKMYaVgTBzcSlRerFOgu87Hg2Hq/sn/MRI7kql7tNOW7Kh3XajW5flCs+6Lr6O+
b8w5TWg9Sy2K+oTcQH4Zp3sXZr2lGz2hPsnTfE/zprNaUEEE/lE1Dr4F2wmQVQYLjlbgkiHiDwbL
gXMCiGeMGDcVj8X2XIoxWGDreFJNZexzU6oEhXtCuUP00e7ogY3YQR2MzcfAc1ppJ0qtDGso60Mi
KVsFBUf23pzL2R+apqd6nlqOrIiak/U3Tl3xMqOKy9lo13BxfVC3Tj1vGOzEfJoOjdE8/xcYSIDp
VrELIvb4o0WTr/avCdh2DeIDXrR6Gme3a1ctSdBbxKJIdYOTW9dbw5DbviXdNKGT4uuSi3bOgfxw
CH3658WcYMGObgnH6YyhPIFLJpeJEB0kVgOddxJUY9LkouVtow5UGFq3AcU9/BFoOC9pG7AIwf1l
OGkCFmCJWg5t0SdKwSZ4h9JS7F8JL0P05m23l4dk/4Mcx46p2TQQwo0nDV1E90Vcx2MJB9cn8sY8
CKybZfM9UK++ilRYk/1zoeRmMGv1NaZMje/3cLXZZQn9taCGQbPApmVw2/jkX5cVmpVUg9VHyWMS
OH1FDn8CbKOPhupxgzrMl/urUVegB1ba/CYNMhsj5EiRpJNaQGslV67nVOQ1niAjWm/UYTDIvjH0
8OToadM6tGOM5biL68hq/nvp0iH9wfKZWq6UOrrpRX5xqLVSpM8dlDFjTyCM6mxXObn0p2OC4nvs
fSKoLl0u3ZHL70g9RrU+SBtXeIjWpJOWN5s6G7Cn+jB52+9v8/CMs2kNMkA/0Ntfqw+yXBzoP0At
uIV9D0th0dEJTWgSSFEFDEQCWVFUlwqbmOgMwIRlU5C6xZ756nnsR2ZCuAZRsr16WxAuGKVsAAMt
KQWl4IwmIfv8pBloF0IuNLPTgBJt1acbp37x36C/N2DN9hD1r3W2xDlZMa9xNazeAxmUUb+whnbc
fnJ3wGmspb/39aUPht1EIriAWacUgsL2bek0VbPNaVgWMmirdXjNO6ko1PPgvXo1aT6+vGgquhx1
r8vZ8feX+SpNEmLgz5COrEilpxwmRgJ/U5INwSOto8M9YOAg/HHCiZB8+IzlVGWCOWtpGUwe0lRm
My7MgV+oFtidmpg1bJwnjYltwZvQxBQYvp9uAZS7habII/GoIQXaQQShz2JEtnKMxxcOVpMFLmVE
dW1+lfMwyAYFFcdxI1iDGbftHhUidDkFbk+pQ7tmTZGRfsp76hyBdfDEtNvBjfmUHx+OfgPLmXMH
f/PjIxNQj79zDy3txEHF0MwVvxIxp+b6EGe8++hEUgBqZ3k9l+zF8GlG0f+FUNv4g8mU7pdAtj8h
Q0uTgLhaG2DE0mQiL0cRJBcy+XB74HGXRJxvjCA+fMCuaZXRLAWO/yZlJX82SNO0zuX+T6zrYtmd
kgHeevjbicG+yVaeIxhTrpeHe59kSvkEU3DhHwAHQc3bQ8YzlRI8NIj8IFKtBq2oiHzyrAdI9cl5
7kd7Bj95jlKqaKT82Uy0WtL6krtiS9MMR0Gixe8DdXMtCjcTvc5cU2Bp8G+3elQA7YkWHEe8weDn
k07iP1TfaD/9569oRFRUmHJ5lPw4y68bdLQGqU0aDD/gFmcDDivtI7fiWmkBS19FrnXZeZXGJbMy
SIxz0DIlLW7zsi4oBy+eljwAEZRQXzKU1upAVqaycfasMHYD2sPmAlVNQayMPx9HbIBDrfleNEoe
rCFpQlSQA5cvji3NUkfSAIk4wPaVYnnm0AM1Ss5/30YrqK6uDofMcAD5kEV4KGWQAYwuRCNS9tVb
3iLLMR+hQ0HDTnTlRhlbEQ275zyJ91synFIF6BORHv7NnWD/7tybNgYKDY+54S+6plu3p3Hrk5Sd
cWxxrA1Xcrgc4SHPMfl//siDkpm237oy+Jty6BYQUXtIIBdoKf4PiavnAz3NFOm5RjqNEPGMrweY
cnVdhc8+8G89n6oMaSWi4MaDtA1dJw9dDNxKW/Lg1A7B6emeFv5KOc0xQ1iRLw6ANLe53WKrf7/z
31KRB/0XpyoUlBxy8dSYYMGO6OxWsM5T/0Tooj+k1MYmF/UyIsk0Dg/8vggINksnPs1w6AquRuop
sYpwgM1sdHwOkIMJDrEBLR6NQaFqMlkzFj8GTcjGrLrohImjJpGcARoa7BCC6xv5e+6BPsmPLdJJ
vRJ4B4qJCa3YzfdXr8YGJR1O1XPFEnXPdyZD4O/w2WcZizpdKxVancdg4MLggiJjSqbSVwyHvy5N
d+Rl+omu2MKAVAPuSrS26LQSop8vSIM1iQ+ZmeNwhG50Mb7GwaD7plwg3sn/ZDUUOaS8p+zvgLr6
esiXqKPHHf5qUbY9UAAJURzDiW+4gaEzhn9/jTkNRYgs5H0uYTHj/h+tc4lT4L1Pxhk6DowW5gDU
rU7o/X+dtgh6wAU6uBjJlKg0D3C0NwXP2aRqPvI4N+WjQzAmMw1kAgMP+Fp7pUARP2ugQ9OdNRoQ
GUTQlj6FiYn6miBbzgNMS+XW00tzFQjoe4LyDCTQHXLlyrg6Glr5Cjhypk1lNArhpUVSsA0HjWRW
5qRuPT/i/Q5+gerMhsmscFLJsliQOKsaIcIYRlxU2fiH22CYb83lTmQU9lthZ9gY/+4MML4KqyGh
s0uBHTqtW8CwWXxrgiPaahCMKSTKdR5YQ9Pn3y3tbfjk3lETMEKHc6LdBKkb3DekxVSlj0Bzad/X
TDw0yBsUjCwwTJZCdDMNQcmi2w2nJ8aqEwUxQYU6tT1BEs0IDa97C4gMTpxIJpNlEap2N7+mXfQB
R6bCSSEMXLvlkdZ7CIOnit8iAA/jOI/6Yb5Df9Tr/YagQS+0jJXHG0zoL8eiZ4NBzjYFnv6U/PdJ
JYzDeqRFyw0J47nn+7GEO2kAWCOYfdFGsYuJU9UFXBla86PzJxIZYckSsCyynJXoKcZBk/WvPH+J
dN97trDS2CiQrq6NaWpVzY0hdQDki87vGMbIT0XJu3pG0zlP5jYRYCpc4Klo7+iaQxybMoND3CHy
9x2gfOgffXY+0WP8dpXjLEg9L78q+qW9PG4pKO/OCzTgIxgT+Tds8+TznBMcnV6r7bpPPBkT2S0F
bIgGkJXZA718KH2HVvHGdpTf8TrHvp6wc6hTgVQwu3W4TPeZIflBzdrgFfYvfYuUcawze4RuTChr
hmfThtUEbjSw1IbBwaCR2ZpKZN41p04pVlSwZ6JJ4bRxIy06iIO1XBZ68uhnb1Epew+xfmOxEbwj
QHz+VEZ91XiewLpqacj56K5skXj8P1jkYPKF3IaRfn/KwRZNR8UOJofptBNW6diqyXRtIo8/AUNo
/GMHHWk/EfVvA/TCAio0doce7KahbFOUgOOBg/Gb0eVahlTbizmIuxaJ+YMl7LU3ENX5JIbzCuHg
5qxoLI5VruQ8UJqMKylnzhVyh+6vf77axO78YlgVEyuXL++YofCJF/wnYBn4WcMO8QKIVrgUEFpq
2LiWJmi+bQaL6XUTakhnHElUUxrNZ7fnlW3/sPxwSQ8w4+m5lPQw9CsAbvMR94paFY9qzcPeWLhz
AiTHoeraHrTvfkXi2Miha1mseTl6f6OpOVRPJv2KxdAIIkQt1D56dl10jD0sSXpVxlLrHQQtlXw5
GIzWMgj4c9A0LOK3Xe+ieqPAJtKj3A/cfXBWL25FTw5jcDJTKNeUwjWY5bMWZQunSSgjtoBK5+RA
Py2IWF0g9HXsBOOWP8Ey1qKa56vloyffeVET26+QUejJHVJG7chAtvruC/1SGt2goZwlXSzEhWTt
okmNR2PCP6E9zZZOKz0oO3ArvFnhTHiinttKMMcnL/m1ruH609wZdu93DmHB+RNgcMTMUEtEdlhW
5nxX8OXN/MgIdQaYreADjySNYu90S3ieTst7WbzgDiK0lZMIkgmYYNc7axfFeiFOAIS1081o+zFp
o2hkjjbtA3D7DNeLIvF7RONYS9++p3qx3rjUNidFvM4BuqNI0CnNP0VKMlD9RXCoGWgQfyiWFXMt
kMPhniVtcfgBQLebRbIrH2+LaA8/wgUujhjoPny9gGqAZMvPet201VCtymThmz1RsRaHZSpvPuHV
Gw0vkAtOZnmfL7fpyA0C8tCcYLNYCqtJVT5nkK0O5esuKxB31DtXML35eEMClnY4r/LJes+HGov0
5pBbPYkgPmCiwixr8sA/az6DMRiVowu0aPrQCZtVidijz3ULhvLleZK4M5y5VEp+WUjP1/XnF9B2
OlZa8dNDpwt9jLaIxwYCHfVzBk2TWDwCgrw/4U698HxS4UvXa38g8wYXq/0/mZWOXdg0sbHq7qre
Cg66MrE6EIeCPB4/Ms3eNR6VohVo4KI1vn9/UwuIMsuJco/B0SCzudRWHNgV55U87VQOm1ls112p
tZGB6D2gGtUKRrkuPiVzLZKpEk10p+9yBTxrOxpsvYIQIej4+4NiMxEFJNBipzpWchnCKPARGEme
ybkxfMeLfQViHftayYYSrcqnY3VqVt3YaevwARRwod3bNMD4nT/UAAqqYtBfrjXqZxhhkMXrFj+0
AqOIWNrAFmaAEnKOrn2Dpir5IYO4OBZItaNbugETNVFmT9Jr/nryoeGBNqUaOvzxMoTg/vTa/cCd
60sYHWMlDlaW3XqP8bYNeamGXetF2W4AN/cY2+LtbYC85eGwd1eobEqoathpWqKVrIfHd7MTbTcy
d8HFyUFLzTtcioQoUeWp/2QwJS01oYiBHNrSrHqJYpJF1C+uT135WV3CK+lP2sG9aWU6dUcduBQp
gYlnf+04RyAJwwEMAdMsHnyzMimw3lKSYk/ggVYIDI+4BgHlrERw1MouyXFg064tYJAmrO9xePGL
cYdEFwKGuQj2vcTcAR7Nl5q/qSK2p2wuyhRSkTlNWAZPuSK6FTKvs/48CwXKPeGC6roGEloKQ6Ru
JE5uZKsTaSNKAJSO9Jce6G9ZXBxcnDU4YPLhNFuVuoV5nu2LKu2qmmSXWtLJJ2MRQ6iz0WUNC+jK
3PT4r0Vc/ZqVkLyutae7w5rJO4OXp3DJOlJ7lmsgI3xLgrWUF99rkEgQGSqH53tsZwNXuhh9rnY5
iS5eRoAiFwm+ky1ILRLNGr+4ulSql1z9P6O2CyLd511kQSwmQQ+aXdw0z3MNvd1i5gFIOmzZbCsi
Wk+0ttEzYdIRt6v0rbMgAFVs96PQwY0qmpycxB9CBXWNVeEgLygCJbA78ZlO3opEtYL46Wlh3MH2
bFbidY29g8bGYeLc4bu1MOOo7O9CyColKEFFqjEo6nt6ktU84E4dHGx6RQzFpIrf92e+WFMkSiOX
p0jWUWT3ITOq0i6GbefiC7ctzrZ7LtvHt7KI3K4FUYBSZQznN3kEWg3H5y2MZob7Vxc81jeacs2k
Ug7eQn7HHmWGoF7L7vQsryWsf+gJBs9qf6TfMKynGtsuAZrTWQAALaMC9IQ7/ONvx5LP1eVbkbDJ
s5THkHXy6Rw36jFqowAE8zQhOEWz0tndK4rpHTPEovqAMOH4T+RWU+A3Fi4PaCxDrNf0P3BzgW6n
/MARMrkVSgW17EQJ+tuwjnCHiupmgLonOX2+Ps/jdQL/5aT45JGSB6Pb7mfzs1SIN/BxUV+fmaeC
BMLM1i1t7MkYe5KREQjJPLQX5psab1hHsyQDlFCacjtjfAHQmLH7BJD8o7Uw/na36EsPFAs6+ZkL
WdJBQCLA39SEAXw1Wmt9cYmBWpM2xQxT98BUFYjqDd2ufduF2csRVGP32BuHgyRDmYDySBV8IJkD
PMvbC6+12yHXd6P1bnLnBintVrOU7wbQA8pr/kVEOZ7z7hwe9Lts8IJV609aKLmLtwVZb/DM9w3T
B8aXBP4Vayjv+GUUgDm8ui6aO6/aDJ4jAbm3c5b+W+8gfOW+SH88lYhNQzIPaqxhQYyCb8kWBXRK
4LHvMAWnjxtDz/TI9G5eeSYyNgzllNLR3+X95ylfRLlUEaYOnFjxPb/X0NYPhqMWHttRVWclU2+T
L+IPM2uroBiYlX+2hzVNpXT8Lhe9PxouSwaDEcc45zSfVNQlJzAJy+T6PQH856efGIThvUtU7ryO
UrbRBMGDxtN9JMCgWdFzcNWkBpKIYcvpF6Omq/SH9TdbLfR9mLHjKNvnSgkJ6Xn1W3pmg2BuKEa7
SLl3Vblxx7apgbkm4J4G7G0hg7F/k3O3lWc4xRr7jQY78Vw+tf5EhbD4w6Gv6iW7C3O9CrN1RRa1
jFeP46eDWvcmPEfXaz5P5z7g2dPXqap2sREolYt6uKyH8dk9jId9SK5UNGiY3S4r8sGfhLJkBovE
qh2EbbSEVzWmzPGjv+PIt35YUA7WSIhq9mMwcPn0RypSHN3CFz4SjDtgT5CX1+EfatCOn7ibHCIh
HJHJbJ3BHOUYcsD+pBBvnPALQGSmQu2PPrf1RWHa/QGD2t/4FFZn5bKxM9f/Yr3vWMJSgkgGTVRa
IQGXvjTu6VFtYZwM5nzLKh/QxqGGG8l16hme8tvCT9SAE4ETysSAey1Z4gizdRvMXT+d1oolreT8
tm/T/rIWT8ExpyoIApzDvMSNVaWPlV2hLL3SYR3guE4vnkqX2QsO92qO96Jzgi/g7O+f0VxjjBtz
lODK9DKhvhsCdQeDucu7VDJjckAaoDg5rfqBp3Yf++3k8GwErNahaBgBTAKX/s+KKkcRgh0VNyHF
0ooVZX0aKSLHwkGECWtu27ClWNgKkvfQqyg8nTOoXYPRKkJY0RMbyuv94ot+UjdMv8p9cWAjlQq6
XYSRlm7V/G+NkR/8e5tFVwCM7kzmJO8gPUecg2U4QXszvSFvXziqs3B7HvOHuYuuS5k7nEWkmwL3
b4CtAMg7bcvzdpEQXAiWZnUnKXmdfLevbjypibwP3Tpme07qdclwTF6qdeirUP2m4J9V2iqBzFut
JSzoWXw5rklgd+22KkPLsnEl3NPF/2ksVBZZJVVf2iebEgN0UbJ+LtIFq9fprPOBVJptrWg1vo1/
scxUhB6c689OcsRSG1zA8ReIrc0hXb10bI5IUxQRzsfEjspGDre7YpKQR7jb8l9MHy/ijSBpG+f7
jm5nBuwgb5e2vWsG3OCh9prKzlGuvZCB9rUN7SI2mRv8etEwlO1GxWswo/9UVxoZn0jZ89BsMVT9
ItUbUGrCTHw6M2Nr8FItlcl2wJ/Xcb/n1LPi+Q4OPe3R+WKgTgAHfiZRLPejhbP4qJVVa3bqvdS1
diPSQfdiaHNhU6jH6PVZgqnL77jYk9ZoU52+vRltmoD8+mW+l+QBaH8tTvk/lpT5twlI8fVxJfw6
/C9xZCwhLU1KFUTRvXCEoTzvZGuDEMKXN5ST0494c47eMvSxtzERAOhge5DvvIpNb9O39qqM1iPh
DWFsCVvLoGLLqgzy8Q2ktE/P6qJO6lbM9nIO9C0pjoS02ZTF7UyrVkxX9Aff1936QtC2hn0G5llu
xpfSB0z841GYUiHydDVNGcbACDsjCRqZudhMjRMZ5ySV0bUf3ZCUABMZaH+q4Bz79VTtHATIZvEC
O1s0/+0CnIPk+7Xt9qqs2oluPLB22Rqfx7batyZAQ5lEh9hBNHnjT61xZ4WvFpQmxF9nETHFQ/5i
X3+6/kTkljxYmBvEGmqmXcwSUu97eKnOfyoZ7jfxaD7K5dPf8eZSW4q0al9jlTyZoo08JOx+ySc4
LtgLXOn/+ypCR/y0i4KgUGFxmEMRTto7aPQq4SRggK7dVv6bXxGBUbNbJQuV5054uCM5t20KxSBN
dSdrHKOC1OltvJ4g0Q3rI0ZkkRshKVPhjpKEp8SPUu8q1/8DpsUROvl7jkIuxrcbfleQcQm2wG0r
9WIwIirbTX9n3W6trilDFYEdLXmU6bm7G3Z+l6xdNFufU8iC5A/piRxZH44XKXRgDLe9b/BaNOsX
hfv2dsbHMH7PnckYtmqY9RCB57Z2GwGTcycQoXHJkBH+AixZH1PLRC1I2MtQWJRbTjlZgYHImLiU
T2U+bhkO2ZH/M12AFLvLScFGZHHinsp5NdKVIKgAD2GElLARXXqIdY3vHaWh/Vk3tx1mZCnpdzTp
EVTnFQx4m8SwcBM41VmeHqebWvESoilnsGTJYFcQ3m1F1BYbfhex7127na/d2sIMVwot1sgbmGeO
rGHXjoIRRm79Pjsa9k2HwX+3yfF/PAJBecSgricjza0ovemafwHK1h1TGDfkQ425yPs2w+KbZm+c
1je58AkFnPOVMqi7HL30yddAwQYE1FONv1aqSTjdMCoiIPmB0LIqCt6U/aIMEWNNhR76OnzYBHll
ffGhFDgk7Ok/pAm+q6T0VitaEPL2OpeLNhX9MUtWuemicq1Zux+veUZVBIwnIxjBJUl9Ib2uiZeM
kQwprHaIl+rIyFV9C4X7JCfaMzLsY8P62k6Ta6Q70Ns+Rz83nkPObCpeAITa2udUduVKWaKCVYaG
I5ZiCU6WQzhAikVm5y5XbLfyWV7edZvVU3PdnOJTGD3YHEBbLB1v8oAiePiDpW0IGC5zO675WErc
8Z1Nl1uY6uEMEdldcCXrAEBrSz7BpsXAWNEwGo+mYuAdaRMDPZ2VMBLNLoplO47p5vpCD4FoO5ql
4fa9rCwbjo8c7sMdYwMhTbGYGaz/lB53VCOGdhK0QrtCiX7DYcR/OslU9n9PjOYpZMoM+KD42B5x
J5rqdlbHRoRGho3XEw6jHumijdMQz/nuzaXImeeoeoaPwLSug1tDjTkHdTtJd25u20DfoaALCAod
9AmgyjKr6EWvdEsGx1OgWF7SWt7lO32Ppg7+dtfw5ZG+kb5a/CvnenJNw2JQBNBDQUQd7oZqijQK
9NARCkx53AB+75Q1S4QvA3Hfz1RI01ol4/CyeVfXqOq9AGbOdoOY/4ftyR3AEvisEBxCwzVb5zo0
a079FV4obA+mCUUjI0p7IjLdmS6k2feen9Z+9dsxbGrW2i57tnTxPLAjWTPBe9vsLHwLmtiDueSP
rBe04LQz02C8Tc9P4rvdYVB4CtccjmF/FRIhgTO68UzAa0Jc2092sK2KwOP8pd/rFPdPJF5LdZJN
HLcrGa3dtLIwVbTKtpEMkcYca6cVJe5ojq08kV6jvb59lT4ODl50pKDvtl6TLwEeZq09cQ0uTa4h
TbmuYt+ObSR7vE97N/1j4g46l2IhiXtHs39s39JEsgrnDklsjjGjpAitHK2HeMDbYMsG5d/P57Dg
bdWB7kkpdNHszeeXIVIBr5L93mCM6EjIL3Oq6G9laEdbRX5wk3KAo2xfsbQ0i9G325IIhzq8S/Fr
7gwm91eKFAIlJZ/ImrcmbUA82313UgyXX271rL0+8XjxQqWX33AFsgV7q+QeYkhz5EK3bjvxiKwd
jFqCmjsDJiDJoubThgYD5FCa8fFLDnpbPQXBoF+q30ZjMRAtoEx50g1CCCbiRviUnFogZcQu3Gkq
xGJyC08xhLzgOsHu7aXjS2vAmiJX+m000qUJuVZwdZ9YfJQycQ6wfyVjBCAIHKtPrML8dlgE75i1
Fc7rmYM4zdTLfSjTR1I0agiaqutzkzPxdFiRw98jhOauMduoIppH8g+eM+5Ii/d+FlGepuGBO/Ev
ZT72jux+am9QA1olENkW3vEoiq7tRm+u5Ol5RyYgVjpmd90vvLoC+wmgOv8LDwWNQuot3SfbciON
qWeYRU+At1O3EHak7EqGYI5NEkZtWS1VwJSigV3oI70gkobLnFeRWkFSDInN/odPJ0aCFA9G5GC+
JIysyQEkokFJXFk9xz4jxjYdH8L7yu1JkFHrCkqt+AeaDL8hrz06ZYGXcErUem9z4LKIq46nwuSX
RASLqKvFgl6NkOcEwbsKEYuj3qccdo+OBhoMZ9rAovBOIMLqRomAqc2Yxquu5uTi0/30wXtcBKEB
2ZLZfqEoAl/VNCleNcfnrQrJ7UGaLzfPuDj3klIGub8ZSw+khzUq+hHjwSpJuwv9ffqlFIhCxnnk
yzkDRaTLhclRh7GQUE2N6BSbgoSWfnL82BSYiIK6HpKcpzqWTAC2V1s0/XV9WFxPCJvp6O0fzAwa
4USDLy+ZennXTgB3KmJ6SBH/qce8Bb79WQyaECC+0t/U0GNRXFFc7zOzJ0C6uSd2qSQnBUSfPsVU
h5OEzfc3Fy4Odf4V75Vnkg51gJak6LKdSRx7JE/szRMF74fpD1oBPTLGrvlMcY3xWBDnLajj3jhL
V2pdjIwWJrRc526xEPpBVD3/VbK0DCNokGf7ZC55wC5136Ia3J4n3f6KbnkDw3pxbk4jKeEsdVOQ
mlEBPIRojqTvCX+miws65y9c5G/fLZQzB7ni1fGWkUyJ/lQ/KoDZS7ZXI1rSYGS3JDYCy1eLsAYU
UR/39q60ziAZq4qKHRM/KsOze8FCG3/n69q5c3V5I7gta2GdiOR+pYReyqC2b9oLrvLKV/VyuZ/4
BapXIitU695XCnJyYCqBClxR6Q8QEzV5YKRaY/u7k+huPjwCDgqSUoReIp/libABvQe+Q8i7S2Lb
uRlpQqXLcVIJ5hSZjEGquP6ivB00wYnvT2bPNa8+Uh60E1LmgQd/MmgF0wZ4NfG1qHv8HCfm72+H
10rUbys1m4MJFGaPTU+FMpwswOPLXmaggx5Vt3FfS4ncrH2zhd0SE3ufgAR5ckweOXJey4BPCaez
cAzG4vwxh2SAq+PqpZnVRXZ3Xax24KWsBmHrOKjlOkGNRGyzb3f80aTKdglgbOb+1j9cU7GoNhM4
mHM7XvDJ7WZyoBbw39h4FPVeAS8CO9TTEgUF6ezbfzLUInappZ58CwD5apf0etpQ6Rnlyg+fCNmI
YksPnLoAcGiHzyjhYVm8Pzsjzzft+FqnCsLOQLYx39rxSrMHl4BKapAe4mANalDBQ1aQp3uhITxB
laOaPzGPKRI/Qn32skpprHUwLi9EFHoorULpu971fYDRY8Dhh6rrEqAufJ22V2JNex4ZpX1H1gVR
QLBPBD83G2yAONCmTXdqcm71v0hUZFFgb4CN/D0GK8S70WrgxWNCaxB82OXoHbAp/UOdytcxY+b6
xbAdnXvrBdNgJsfv5so0BGSWC+oNv7KfECc42Bzv+VT6GsQu+uCSJRBhyoqWDxQqklQmhKOLZUb1
qFCPaPi7GKB/PJ3DHyZ+rDAtBdT+S+DNNh9nyOiFcfldQ5AJJWrzvueR8LbW6FIZQYtL3u8Kg3qf
TAw1lu9Bkp8Pw/MfZqWpyDajJywwDOS5CGozULfXgYGF2tZOcppZ5ySgYAyDEOy60VadpTmfCpgZ
sUrS90KJd1EYuaZX6JBS4pDHKNqj7j11nY3Ft3rWoqHIsgaAzwAeAS8aalcfbBC4IM8CFyq3aAQp
5Dtj+RthXO5Fh9qLahDN/ndbKaFTjihwRQT6dq/tcX+ys1oCIzwVwc5bdvID5DJrZTyP+ogP8KZJ
SvklZ7GhVv72vO8IkqUJA/K/gCczpDPayXY7lxW5dazLIm0bg0n86oQo0i+YQ6nHtoZ3QaeWYfar
j9vWmvmeO/jDFWoWXHhPP8T5cJ6JNByO7HERM/BwpTvcGxuGr+bKbBsqIY696+O1hgmYg3B55BCB
SrpjCQsHjdjYJrQr20NiUmYsxqNJTUQ3hZn1u9c9TXSHVeHOKYG4KvijCvil/IBdyS1KfMbiT+Gf
JfBukKygZ8QGpOZikqvMG7N5pp11jxLoMoJLcb0qAkXsd2HldjW/bkdZPJOsqYtZIgBZIFnA6bnL
lbZtZ5elJA2gcj31AppokEMmBI+mZXr9Uol9PK5R2OKUF8LtNCqXmwVmmLynhgqj4R8FGvG0nVZQ
lOcgoBYTzZ4Si786XMKRSLB+sNxFrLmtfvVWebWMklR6fbmuubf8k/SeZblxukk1jmzHya9p+3H+
i/OHqelctlU1If5Z1Nvqrz3Rw67dvTvtUpQBCPB43YL+/HteBt8VwOpIHXXAcKa2G6dpjZNYhRAT
Riq1BpIVVOEk6r3eVq93R3ZbzZAfdViDlHxDNmaMzQMbLIBnp2+fwnlDZmBIVIlauqjm1nca5DMJ
F7d8DiLIgmcszbGWcqj71d0bwKlnalMTgYq44me9xNO3DLpww5a3LV7fATIMrGQzAOUZTlzhCJzI
+9zXyBIPCuucg9187i6gGQp9nvEStAiFeRwqLKm5Oe5WKjUmfXQ10swGAVVZ/YbmrMcJdMLM3WxW
VdwU164scB803OZrFtDu46E7bpIhlgk+Hyi+XNhXk/JcTp/Sf7uJGScrUpq/zMWzZyZ9JlSRZoha
jqEfC4+JIALKdyZ7oPKtZYFIQFXBNIYrPsZUo3pVvkxWSois1o/NNWGPqV83FMkR5qXDfjDOj0wu
AWTHcrohHb7QdTpK2bSnk1Ax9PTnGg2zHMlRmuOLLtK7ZZGDw+p+xzQ2sL98d9qaLoZoUtFMNKRI
mK5jdxGBwv2/YiG1DEJsob53ojrmhdYtyU+0Uzkj9s9LW1ge0Y6A3EKY0omk6RakjdWBNuWFwnkn
oBwW0hVLqv3Ups8HCOcDBvXgzzRSB988pC2GbKATkBTcWwiTuxe2vP5zhQzVDGvx1h1Dh8LHbeMK
ZX2ZWtUAaAzr0kIkPMXKy/YmQYydQLNhBmtHmF4lmqB7JCzffd3L26cWs9Qn+kQWNwx2xbYpxfPr
58/5JbLntYUwttICfTYL4I+Zo5M4ebdZsLbmu40ABqdOHGnkzlgX+Kck2QoTbKxhsItiiXPcxvCw
+ztbhrPNSCHWqIrZyRFTfBQ7lhJuD3DnKIQB1siOLndGohj4ORLdgm9UoP5enbz78LcSkeR+7qdb
fAcJp349s9nXDg7i2zyRg3Dpyz+Z+WEgBwFCnfRkXvFMnlk3zEn1WYtTuZIf3TrB6IfIFT8j1HAu
uJL0GvVrwYaGzuKvalJINPFO6Lq9cibr/x0jJdX5ijrqRJgLYIKAKtcQWWGDUiva/ethc7vBW8h7
Agbc9/yHbgQaEGcu0R5RXRW/3djQ7KUGwxev4/FJwntoWzjqZf3iwX8/WhLjBMEm77fAqVcQfUjq
UtGKfuLg6vRgmT944iHAE0VefpiiKg7EDSGqeQ8hrtJSyd+b+s5khicYYz39xLomc0pLUsJEFQVP
k14SY4tW+tK6/V9mOVj3HObOZTi+uT6rPcZYwHumcdCw2W4+ZJwJwkFLiecFG/juLepT7HB5h3P5
deWUZsABglhWxBhzPX0MwYG8clKyWoxd1XVwL2WsX4l+fSl19ybYwQKOGbk5IwFor8M1apP/cDNR
ipLJw4755qYzvNKvA8xvF87xXGwxZMVp93BFWb3coxh/U7L1lvSO4zRjsdd+lBygBPcaVEUg5MYP
Igau8U6apWlJ99ZQjxZDVSC/Aom/1BGYyUwcRTYNvFp0bQkj2SlyKkQo6KRM77xEVRuf4HMfPydl
9VSJO/jg1KOq5FGfTFpPuatkDsHTev5zyObqeXWoRs6hSfXb4A6a9w0oFNEwMFa35aE5kicPxYbC
ibs1a+HslbgtAZCods7cjuS31Yiy/eRAIruJHExAIDeTahkZ8S0k5zkP5IU/5LCFGWpm6zVKATEF
KeaKv64xtKS2O7C9HqDzBG4PIxgqgCCT7FGmKaprq7k+qta9sAkZkKu9ykQbG2ATjmv9V50KqbUh
pKTgLF+24M47a7LcGJeKD2BGc1BxDyPKnYHGM1CF8rgG+UJe4tRJI03Ei3DRQqSKGLJmh/tbCum9
PhlPxzAdx0aMmLC5iMbCGRu6Ti9CG0U13QFi4492HosD5SPzTVIKQx6VYxDI0rv/pKOCVSzcNDDR
Sct/b4AxUg50vz78Hzd1KcLfnW8wofd8lKTA0/rJ0pZpdOmzxW8jFrHZ5z2OUpurq2Wb7Ev0gRH+
o2zLppytIsC00mI2CA/Ud7LrfqSDKBq6sND36/SwN3A3raBksjwYimwRTIL33lRDL7D+1B3oHA2U
PppbbLRrscL3laLGyJVKJe7S+2l+wnv2j8gk9P0OFmRAT7lopu+j+JhAwIFBAcPvS82ciIxwi1pj
U7PP1NyhpU17eGTuWvPexDvMhqAnWsYNE57r5CfVJfn+HG+momQMM833wsuZkekHRpr7NYEzh4iI
bAz5qXfppEe9l3TZOG9y5/LMOp8+NqVM8bT8foSQrKMwcVBrlf5CLCyHoyjgKzGSklfRHxnwxVfP
KgebheZoMyhQT//3JrM1mvAWL3sg4QGZL40QMXHsehwat069av6jxidEMAXdGi1Zr0+OMBDx1uNo
zYFveUSyJmn6r8NkkeO0ipC0S4QFZZJIYTWRHHlse9xX6uxQHQddoMztMtZQ5mF0fGgJEkimGaOG
xD+6N1L1JLrdzNWjPYVPCo00UElHXCqKcJhEQs5CJvUjJu3tKg7tKRsVBeqqHLn55FPIaq/GL0m8
qKFEqJOtfVC5UnVGLqKjKsAv+k0YwMKNdYFw0UEEKVoder+8Dcb721kWurWmvdLSKwEbEAKr20S4
gmRs7j2mC692r8gpgCJAgM6uf6CuUc1oIKXNQhBb7ROE7QWuAmMlHAICiVDLAV0QhYXkgNKxFcnE
Z09Yihh0kWs9WwLLzb/Dq0t8XkN8gKniG6PrqKWy7srpzdEGxI0+3dHlnLhvG5knWC9augjSiESq
QTTYoJnzA9gBF1P7+J058TYfpHrOKCFsx8ey8ixG22nMF08QxD+S9q5U5qGnWxaoU3mYdhhXPJt9
g5L0TtVAWgqSxHoH+PMNHnwg+iMUx9F6T/31XmwmlcK/m8rcCPnrQizK2m74vcO1FDS0lJ6kC63Y
w95lv/kVXc4k+SxOSSy0mFI2unIve/QBH5KT3TwkRx8XhkewCB5ubtuWKXBqi1JwyjtmYExjDoLC
Hdw+GGM/jTCAteRZl+TC/EsNklkjgloCxHJI2rRyx/ODKsYQlfsgLBWINfTmVmXJFhE9rSX5kVAK
w6YfmYzIcsoB4l0daFe6LpSR61yPQVOJu0PqtILp4pZ7eibT0ERo04NuKkS5qUHVjPaEF8I+Vqgv
I38QUWmbH9M7bg23RX4l40SZhdFqLnhRVYPBaub3budC2Kl5JFpWWHbIrd+UlLYhHmla4PmgUpMG
UjFwf5guFPwUrFC1DM1blzAo/x3NnPWR/Xs19B2+CGIAkgY7dOW6Ljh3wLx+UzUuS/J5t23xOh7m
6njD81iBXsZtrCAN645Psm1mVuuGQIXVASWt649WKZ4x7vhbVAD0tTt14kwhXYhcU4P1GXLz7JRC
1utN09Ijm9w5K4riin9RU6BjzeMlhEf/17qC9wZ/x4CnIksELZkr2cDlxKqfAzQ+vfq3IOOoRAHE
aZthTwPafU56ffP2dmgdoLlIre+YFCvjUd1doTHZr+Clzma1DUiQ9BReNTlWxkmhWAk+dVeg8MV1
rW4RdM6HzgLupGgyxCbUfQpiK8tOTfrW8vjcjo964Z0R/EHWMKHFB4Eoo4UwuoZlByQrpc8GlqIF
p2cvgXH0NeFGGgvkES+3MsDzh85e1V0Re0PGeBk4YJWoJSNR450rcBqSKbFRkVO3sLJiEJAfxaL/
fq5uZl46ViE89nqLSGL2jer7VPDWGPc/D2ibfjLWzjJKlvty/1xdyWNQQH6fhHBkvu3saL0UOIjj
6yD5zg5Ob61aA2NuBLAOEMxaxrB/DcnNkWyiOPRSsyla6lcuqs3RKmZZaLmuEwb9EYFN1JCJFoY9
Yx5unVQvt/s+yC+O4BLceDkatxQSZn7bbS7opx+EJ354WOxcYd0x/W9Ft6cAbvfY5VtlppXjoysl
BKDEkjbGFuNMgUQj7TTAGq6+fsHomjv9rPGqKAnyAoHHu86DuXVKyBJccWL+5hsV+rESqIb8zkUk
9XV0v9EqiC0obpWzP0yGjLMx1LV9ywFoVZI2rubdworZcI1GPqopBzx4NvRdhjlk7eu5kqIu82uW
OojJyvo3hmlHW6WVBT3V0KDJfxmQrFmS1wUOs/t5CBOf1a+k7uvUKbAgRFAgJp2nvN7htZ7a19Ms
nRemCqDj/ah4VWnk+14QUxMCsOuCR5CBTGFDlcv3FbHvs9wE+J2glDzJoPIAhcOWJBBXHxF2nWTR
Yfqmi8hUYOtsUsX78V9tVqZQmZo18ABaoA3tCDFTamcKBGceiQxRZhXcP3YQDaP30WE/262G9VnU
2EFrdwqDhwBE7i9atNcmX9clPrY/+1y/ZKzafn6NsYAl7Dc3hGv3ujC5YdMwMIVA+0O2dBzIeSFD
7k9kMoqv8lC7AbvVV4q4gFCvBhTLPUymitzBBTTqnn2s4+aB56+Xz5U8Sg405Qff2Cy9w9ME4raF
ZARhW1kGyZhROoKPn+e4XjKc3nv2O4UXbW8s+wk7/yBeqg9CcGLjACsSeg7zSXusNYJ6tUAxya9w
0o1qErLSPVW5GpqGrPnxdb11dAmuxtZ3gDQFQeymhBmBXRr/xtDXnADoyGYzGbF5gIAthrVO8n5z
PbRglkwrLeOjhUGgU+G9+uMxO006ADkPrjx8aQE3w4OGVYGaBy7aeXO6Ezv63g9udyg5O1Fr4tGD
QYXVv3cO08voQoMLLzo2p+F/KVg2wNVMD+JoAxis9lDPHcyRdGnsJp4Ct4BScCBzrkoLHu/YCnd+
2nOVQFpiJHtyheHtpI2eYpmYbQNGWqsiQWr1CLUIHDxh78dS3hJ5kWtX+XQ2kSzkzXZ1sBbe30Sl
vUn9xm/8FkA0ihMiAL0D0brTISZbbx5CP+MlUuWZwkOQ5SqeKYW3ocFXDUc2sV1dj6pTYr5Sx4WU
DQffONDrLYi8+/a20HkSqfn2bvkUmwza0vzxxnz4nxPeiNirvnLBh6eQ6DG02oDNqyxxaNXZbn9q
2Fg+n6ynrk212yVaj7iSbI2uCWaxmpqFCmwcqyFYhWXS7GGWNisXecDkWd80paSH9iSqtTyo7RDE
q9cNYn8vfSR4Ty+1C3OkKMxzK6rCohHJ9zco/Ci++ovf3AbaC0jJ4sUilCdiVqnwwodfs2wYHfL0
UHrEyTaDgHhYQfZEcfksdxn9lzVMmhfDQE22V8s/z+c3hUIEVYidauEbqZF+DbgzvutU1WNUPf+x
5G39VnVOgefkH832QXv7DlvdVf2OcXz16Loi7C9v5apw+0lmCRlolAFOFWRQjKVZGCWDGDD4WINp
Vol+W14eCgc55ljde5BGQJfy+It1pZn29cFK16xIwA2LuxDWyPVDdIo8mnLZf6dEVeKgfTGzJu8o
QzPS1h8G4FH7iI7MIgdS+Ms+h0SHphOyr3brYVJ3blDSNFRhTIXbLb3cDxXQ6bfJKK8nyGS2B2o1
EKS5ZU41t3B0wZr5i4K3wlbUtSYd6CwK41KcaGLRwVVZ33eWraqs0t0WybE3pir6Vu7Zun7A2gBM
J5wSABA8BU/nU7oEPieJ+aFFxwv61LVHvDRGfB7+vjDFgq1yThY4gkpmdP0X/2pmJtMx4/gPh7j/
rYRhCa0BoXs6PUoq/vwq0a4fidX76jypR6leUs7f2TCcYq/BcNzXWLraJ+gwD3cvnhHQYy1ZmRal
u0QgeqMK/95nqKvv1xuX/jfaeBcyGog2ekGqZ+85JY2IXs9JFk0kpvBILIhQiEkX7MHdSSRFs11k
rq8wIxpJo4lUhhUrawY6jTpeI/njRLAbDmJsidakyyz3BJ+N9Ug8iALNwNMGl7KpZiqmFZ6BDneV
GGGhzziuSwX7sVORL+fikk2fgKtic/pSlMBqjdfxctf9ZRQY1SiMUwiLQ/v/cjuXE0oEM4pyJA9x
52Ch7r7RJNROuuM11PpWKvj5N3prAFPo7qANXSrws8dcoj0kofHl5TE9Uek3ZGRRWG+g92baHWNf
Zlh2u0WXkz7chvEAXsbKdd8afXqv9BsAZDpe4JKeGCs1jXYxicKVqtGRZ+DoQSRN0es2LUBoHLFi
ydO3NjzeIK9vmngyS7C+YuCJcOorNHqvTyoIKfRqMrDRMYz/2VNTjCJnl0W/bqtn2U1cCGqZDYoM
SCjBz48PE8hi01GqWRdx5fC2RJ6eWvmipl+QflXUSkSlSINk2Ehqlu8nNaCcMXQCxPYT8OhUNdRx
SEY/FZIBEvkY/HafAKo1dnVpIjuU8GgHxRoVZEmahHTuZnp5Tf/fZr4d27n+nqyJmsRbFwoe2+fV
aS/78yWUcFDSosPLdnt24NLiMVYHvbILQ6JXYqMGXrEDDGbQ7PXq+x9xrM71WWxD33VAnzvD3N+j
ZisyPKxK2WOkaAV2y80Pz6Bk5LXARHcVelDVMO/wDYgSz1mmbp13Jo5x6K/QZbeydlPBCHo3YByf
PqH7P6NbUsCRsEmuDJ9iMCut2BgoQPUWikNhcNJ8hhMVVFot00DOvMhsZtlwMO0YBxid4tLz/0hy
cDRbj0y2jcafeI+5d61BTKgaQoxV5ExKuoMmekotCU0m+4YwWcZzZ3rQzfGXBJCc7E1yP3xxBc+6
9HK10TZ1PdSiIgiQxx57jBkAN5rJWluxKtV/B8xVvrdLIc1SbTLZ0Tbj7zJPIatS27CXTNjlKT7M
omMNh7shOyNOCV4c9u0OOQz2CJBY16V0Oaz5Ihkk5E9cTskI82R50N6e7zyzskw8KHTZ/C1IQiau
/cREEcTQZoRSl7+iHZ6QNYWlTYzIMsAH3ERAF8UNgknDZzx86kCHRyTuYhsymOXn2MeNtz5DlzZb
04usMpHqYPNObf8n+ymhXwz5ic7sFpd8fmcF+OvYlFiGXsZ8NyRC7XmAYoOQh98M5CVp25SKrwQ7
tFVKSjSUsWjx3Qtwxn8QHhRz23naKVwT2nHsxNGSlATbV+WUUdcfpTrmKFXVPj9uQEhrb4ScVAUt
RrCuCrIcJ2YwzHRfGbuWCa5/vWNqW4xzlxFl3WtrKliVWn55NLDGdcwzs46/0hXPyQrQF19Z9oFW
451udsuRc9HCQqeN9/oyPw7bTLWTA3eGyigk6IOgOlDLyiTL322/1sQJcb1VC5RzZrSQT68Rz81E
wuwRF4q8rDeL8/r1ANgEhL1MkqKStIiHRqn00XeuiKFfdphfykigV8jjxox84c1s8ZBbKh5MxO3O
jFcWmA0RWSGcH7ReMV6mlzK5TrVrELLVC25Z/cSupI2pZCUEs+oG/c8Yt2CEPZb9fGhDalfX9IZZ
VgHAitCyEtT4PGko67rr5CkUuyAWzW0j8qrfyskqg9P7iyja7NCeE4NNNZt/q51Gbu9uxYugfCGN
A5WDoBeZCbj8xDOkagsi6nHoocG73OsZL35TxVDqrPTBX7K0Ou/GsMapyOG58rUI449JzPDZ8KJd
DOI0LnarnRxjIysox81HzDdrWn+mDYAtsT4PFkPODT539cRpyK10favLfXWsz2KLOVPU+GuV9sEI
AqNekjeKusYGDlLZ0I0TJ1k3CY+xeH01442tOd63+dITG1SgmhM/QMOrKGg1ZZ17UPX6oTX9L3J+
93R3Ot8pnWw4E1HL+auhhNm1Nv9eDhWloXAuhHa9yOO8LO0CdV1yEGnxeHGuy69K/pXLO+K1E2hu
ls3ANl5vHwxFUPOS+qfaO4vQX5F0Py3Clebi22Cgxk9E1GRbbokSfT9+r82gi45XU0ca611EQmnU
OIUzjMaqHa3Oi8As25jgj6gaD30w7HhvlozrNJr3bxsY/iJWC6AAMiLm7uKWPbKjbfyN0Qj1Eqc+
B67ArByPqeEoPEnbS1ureyH3QsQFwsYOcvaG81n4gfKjghNStjnkwL7IhKbhMIS9Rl7dTvvf3Rhz
KsE1/s+MiFqIJ32NBkgR64oxstsoab/4LONI6Q9xSQlxAHYvcnNwmM8yC3vGZjPlNlDFBSxeubIh
AdC7qRtLObQOUREDW4rBwo3YD2/pp15ETLepiTxtuhdR/mpKyDINtu4fmJ0fmZRJCNHWs7Oe1hcM
aS+buw7mVjcik7utYlUq7VLL5nOZ3vygq3izfLQJRDrO37CwSMYqr9q3Gdn2mSjFdLMLmJVbpoKv
LnggCkw6cYrhqLxdIBS326id7qq91w+ruJHAUsPai9vasjC1w5F2u0s6DZhwFEpWi7S9Fpbvnkdy
WlzNTwF1ZrDFCd1gs1qNyfquyWEdCysjcIUYD29ZSH2f8iT7E/7jcOs81BNoZKgK7RDjY3gdhpPj
dV9kDZ4n66x6IEwT+N/Kv2SsqIF/+v75e1UgqVFSBioVH0yQJvCxEJvRkMc7qmesJcs9MQ3Z2kmq
VxwESrIkmLCZgLpyq7DyFaeqlNXlYmwEBt18uJjpkdBRe/KVVA7qg+oYX4xW2sZ9pXXZj64mculg
pcXGr8aRMEufIfkWwp4q7solyqn3mhfYPwvdwa0FAZwwdYfazMfWvwuNXfK84jgchuVYuT0gQhdl
Myd4kZnkS2LZgZ0jKdJfZ6ug4cv5n4Vqnnr2dXDyzFcYxOdLbmBo+S3yNzgMaaJkY0vESBBtAFvs
kNc4EzYSD6onykL9V53zyfzVyFQY2cNWWxwgywn8a6M7jmIL6sPPH9yCNmkU4X9h0iHdVfysAsSj
CJEJQ0n2oFUYHt2DCcjPNBx/oqmfy6ctrJzKe0zRFG/A72eG/iKduDfU1eX2RRsLKqBsMvgVrzZF
A1lOh8OEo7pPj9k4M4dVSd2QsVIKlmka2+pY9zxzZ1P87DKXOamnwUX7kaITMZUScDMeAqPG5QD9
sBZ92xEXTjLWWprz26uqKNnHi0NL+Tyf7gbsMETLhBwvPbGa6WSS/LIrsbSV8N0YpXH1V0z4cfBB
0+qbSOJo0fg5ENPUTd+K4nWFKgdRONpvFiKr+pfa4a6FEIoZ3ojMlZ7wu794FlAXsMS9qR77TMh3
+diXehqNsshF2MUJUl1d48TCPAaVRJ1AJzcHnZaFVrFcgUsgE/tlENS1rEpuxRpeGkTR/XG0vBum
5ytW4D0V0pN3BvNy/dVyg3PboP++TU5VzFR/PPIBRMbfLavhy93rFh1A0pmJkCOgPCGSWO16eait
BfBb2VXBhaSaj9R/HNd1CzcBa/DRy37f9GR1KvrqLZ56TFM1wzTlBsHYs+6P5T2h5NPQx+NDnBjp
YbgW7J9RWpuE2lQhzOnNP6ZJ7P4HAn1M89+NQYO9jn1E2ZQqc1wlE5Rb7kQG0XPFF/cBaCBMPiJ0
dCnBYM9nh6hjyb/cd2BJkw6XuypiSL13oJElSNa7yOhwP8/9PVGjX15Bi4bncnIHZxY94ega9T+Y
A1u/ANgk14eFUEDOkaTvMJaEKHRvnri9/CRpsNjBqg6pkGSRPK6v7DtsWTSNnzhAyMxqNmga1WCo
duWpjw8/Skspq1bJ5EDvTyR8fyr0XuCmiQzvbrW769aUKoMY3rzS89EtCcJjFnbEp1nW1l50+gbi
WnDMadGgUE5uiJAhbUezjc5AWooyeWiVcanmbXtEa2wz/Z84ko73pnlSr/owEOzX2dPt8xBPNnb9
Im2wbwyBJHznaF7fMhC39ARb+jsySYZiwi7Jd7uNvSKzg/GR4c/bv64h/o0YTlh1VZctIDC2iIVc
S25BfMhybnpkny2Fu2Yaemi8GLz18JZ+2zzuVvET4BeVCaNXdDyAJCYMOp7FDbyM2nxjsGVmPAwO
yhF1siqEXXFjMs3Am5ywbrM8Ro59MJlNhOKDXSEyTvFOETrqfpfHAdxQ0tAbeJzHqAjSqY3fPPdH
8XlV/H0XemlIS+D0mxQyTEwMas3EurfQL1tb7MkMFgihMkHLozklxvcJulcUOvXH59y5uy3qdO+l
CHPHREENZC07c1MfFZkHPUQmG4WVdcHVb7lh1ORdsq5OzIs17WQ+UmKSJSals+1skcNuwpka0ZRK
Pvb+lOW89f3gGLHPUu0Zs/lKN/9rNNfqU2MtIHL2utdXQMIiQG/V07mN4qeRFI1UBMUF3WbNuquA
+m0WIqxMx3PZbQzIcScV3LFJ9mYprpPAmftnc037/hvhZM0QlJY/Ta2MthD8zUmZLJz5FUnHFe7e
31FGL6Y85O4EuVqy5+VHfe7fgyb4NKL05dBmnFdx2xqp4Hdb/DDTa6CTciRzgsZes7wVyQbbnYQB
YuJw4Th8jCD6ZhK8y3fN8ERnk/k4D8B3VJ5qhzCWtyP2/BcsYRQ/UPONiyXSUZ+3bktbiMSSvh1d
EbsUZrTMrxqZDV3GOlyjEr3t4vY3vjoqDxMiueWRlzZta0A4ok/eabrKFmTqM1JVndIkK0ukKFRQ
FDHfD5Au5rbhWwyU+TfQPmjmMci+TXVAbY5jZ9ufM5fduj6pjtMrlYERmbrpSPafRUQZSdqnJrd/
TJsMJw+M4sMtJraubkWfWKLO964ToGoSDkPANHFbfEU366r6a5c11aLVFHe+XU6qWyqc1KJMby5h
M7cayxNfCSyC0wo/5a3J+kFNqtw8c0Cg/mnz/P8WXXoZ5VvEThAR4AFSFK3f08sFNmU8DOtQUzac
QqUN/OzZQWnfsbxMz0Rj+QvfcayLUHH3Np+D/5gJAvtI5xJpeEyaj+nTWU7ZFoO/IDuPlmcyBy8J
0WvDMH04gaPxm3WqfzK7GqZxSBUU7ev+RHgd5gnDa+pRzh93YWu8q9rnUABqlcfPHxYhGbilpms2
R8ktmpiXb7YOwVeXYD3bfH4qufN4skoF2GCocQIphSjyuBvVeWC56E/SOr89sjdR+SByDKSnQ+xW
aKiC/94mc5o53iDHjNOzEt46AX55Kh1x3Ey4pQqXza7q1lMCm5biJxByHif5w1lorHCJTevR1Q7x
DcWCL1HGLyWnqi53wF2mujsTsYIzgRGmO3ulm8qpjuiCV08ovkzCuXph2p1tbSXD1g6ktqA0inS+
iF7icKuHnMVSDvURbVVfpZucmInhVRdbCKSkoylXgqMJYb36FmL97pTgJXcOopAGzf1MzpwjyXqk
puD1eM+8cMB4iMXTB4YPKL04HiRxs0+eDc/87KiJcRIfgr/JxebsfC5raNHVqsPPeejdOyfjBOp4
E3G7iEfoqHaX6gtB4bTXTvhqgTw7p9sizmr6ouM4C0Yc9voI6+L/P0hktMiKN5xXJe8A2Tvs0ty7
Maq+xzlR+EPirrUclLyzauX5H1Od6gL9ydsuyABuZ8WFdxW5xbmQMHxaZRJGY/gZWIHHCaZ80nsV
fyjRT5dQYx2BfMzZk1uCDDcMBZHOyJuOkzk2AMhUBM20jqzwi+jha7SEDOXBoPrXh6pfKt4brbHc
ByjNnDv6SBfKScwsOvJisjb+7a3fIQ8KFKhFnV00aIhQU6MmUMyGYdgPNi8UOMxNWkMAbj7lvjSi
AR05FRasWI2QfffEoILfaoVFVbHVGPgPK/LbsStr9Qg/0nOZXtY7K7ls0JL3EzbsiamXCUtFeMlp
gP+I2DrkxCZy9XPeQlTOAQ6OvQtRTF8EEb+tvM2lBC3wjxDHTFQD3O9ETeEVCDKPwPyrEJzTmX/3
fr+/X15eQBWnba0NZETpiOF+k56ff54XVAjbopao+jK4prBR7rpyJkq25Mpj7fu/i/S1mj0KVh0B
nWI6x+mhbRq/FMJqgtdpnh4mrPFUDzjl6pDxQSL0sMbrYy54GASF1Bc9aq6WSi+EjONSXluC8Udp
sluvR4ZLmHJlLvpONZeDMBKvBqDFsOfi53kkKndwD9QwH7Eq9PdNcqI8OeQuFHFIl+yw11Y59qhU
3VmDlj//wBbsFDkShael7DSN1zWI1O5HH57mD6z2mC27XUhCRSLXvd8r42earwlt3yNVGiyMnjX8
MQkWoZ1vs1SaghBT01Fpn4P7kk4LKHh+cNnjQkA9PGWBZpCR84YovBW6FbqyovFna+4LsKyHX4/P
UrsZ028gW+Yg5A5vRtZhGS4+vwgNmxTXFLSYUKEYQcaYgzsXSOZM9z2TGZ6/Ue8iaDfzVhhu+n/7
N1Cv1XngHnbjBlSbSX5Kmm9sYwBE/AMHMwCVSa623hVSuiXbpkAeqavIuC7TdY1LlU9BbtvO4zRV
A2eAOFpqwzIW/iTuYnhU7AuRiZ2GrZNpXyxfPcSKS5X1UTa4di7yTyBMKbuBQ+REcvBXMYgsS5MH
h4UOwZ1Cy7tzFdSye/BlDCmCfliDEihUzxXiEuhJOnbEwXo9IsIUkLjhq6abQ9oJspP9BrPpVB7b
oq7oFTBWXEAyKAjfk+5f6QTrsHAHebChS+nHaU+fO98/x386jXRS6hiwsqezqveTcOzt5SNnago9
zPcim4OdXELMO63T+u7eJEbsAyVsPO9t54sdNE5hGeRF9JHV3ohXG6DNYCyds7u1aBFa5SkdH2U7
0fKUmzX7oMTk07Owau6xzw/ddubjv558CXcGrohgTfvha++ZGlpv3wAK90CJcz16xj3MlcNjKssJ
yd0F2u+R+NegFOwOJj+boDp4Lgjs9ij03uqiXg+0LafiWxOcXpA4IDEaMP74iyCC1HukrKyS/lwV
hJ+hJNBZ7nRUQjkzZMvFqkbqtPrrAsJvnBDO5w4NfNoa6Ktt8RrePo71do7PKcn7b5fvl+mAjTQv
IM+EaAC4i5gd488kbgRUvXmlhpoeCyAngThKmHJhFWqLPp2o12SnBSrWVDl08ZY+dSv1IoI7SnzM
8dFBx/H0IgQAQ/8x0E3K6r+cqdetz0ggUOv73JHmnhK7vgRpUiMnhe0f1Tw9SaUXUSULUreiyUCL
lLEiEsSJTHbiwVKFkaR/lXFkyyM58UmCDNz5RK1lfkZ0XTRvvej8dgOCVjjA+AuraMQVAvlSAytg
nqWKpW5ozEXQ5pB47UOrNreLsdhrtWos9whVln0/jcuxL+fEMkJ3Lvz2j5V77Ki0R/GX/+grkymU
6H0NDJKkUBGjslvlMACSkqhIDnQHzPGMANVEltiBaTuWSbtVmDDzFaxCTvyyotVvqFhjgXQnaXDF
Ngh+/inFMvdlk6tbmHbdAwRNY2Zt7xLVcxe5xdWapJ0WdNR0loC/5NX10wKl+pZRzdnywY1Lt8hV
epI903jTXHRhr80GiJOqpgSZS387fwKH6a4KSLQz7OqCoV6xoNS3m8Yf24p4KMaYwSw01hsXs7K5
4RtCSx2Uh7bZiC0CT9sWl4UDvosVlI9PnYG5uxh+mtkmeT5hLCoa/bnnFftsdz++xYgQDmwGevxs
gUEYjzu+8S6OyS6KsSGg8safqCcgtJSZOO/8+9jAjbDPEW3YRpVNuQObvh4x/R2t7US/8bEJp/xB
T5jAObssAqSa11Q38WL+AZRiiFxSGSxd1f3HT6U4OqG6miFZvstmacDtWRKEvcQ8q9PASRRtiIIH
dOEfYXepeq8Gv6z+EvWdNF23B+gfKK2XuSAKCIvHP/ynmK2Wt+XHlZUXP9BYMLEr1kZRpTAl7UXm
DzPAxVpYkTrzr4kWlIgjb9aFrsc+fg77btcT2ijRET+zMslR6hihJGsS/DdSoZuG4Xzsmc4MEMnt
p8SVhMDC8glXyDwpyRTbgOJTmaUmR19YBosu68ehHwxUp1p2FDrPl5Jzy1WHVQ6mzv6I1R0d3was
LqMOPRsHFf6kyAPsvHkiYOFcD9xgJTCxv1ZSFUtBdlhi3HiM8AEWZptqg0bPR+VI85dT6+4tV+pu
3FXXog64v1FEnqdo/gerr/Q8u3tifynDLwCcBmPn03rAKQvSmQ2NKYM685kjKAuRxi/LA6JFnjaY
37XcGulMvkc8yQJpCiCoOPTWYI+2rm6KKMkZVI97DqhRhD5chDaTUbWzftSe4+ffGb73b8YFkFlc
Zz6/NHlwPfvRQe/GqzK0pn+FuosVu0DlZgAFWtejEoE3YSzCPV3YKTlvBywQU89cF7iM/mpomB5J
qGy9jMnEPGUjZr0f7DHqUyIE+Wzg1qqtmU2ao1lAlAeA+408Egi/cx/U6pTstO0Aru0cBxLu+lyI
verbF9HPc83nRbPbr10SrvweCxHhlZSzvRGzKz+YoinwzTfat8ERErcNQx5jg/gtQOLEGXHwoT/3
i+Aa44/kHSg+ArF+g3fvHOMe7v8gW8XvGtfaMIkKijJ7vcO1hnUm5/TG7Uz7mfignbG1obT6WQlJ
4GXGvX6Qvy9SD3UYIpG5l0Vfse4WIzlSq0oIGrsl0AKOrELUsd8DqI52qJt/S4w1PAvR9a7D/JyT
dNXWcvPc/uiuXKx2YGtGWDz4ZuSd9Qng64sVuxpGh2nXDuSDbouJqnc6O5GgTOSdtwuqg9qzy/44
Qyq3pV+2q1WCeVNqrpG94SgwnguboOt1wjgW4+//q3H2MkyJpjjT7Nc1bUb5E392sF4UEeueVe/O
I0qkARzi2prvClYeg1FrVu5gZzv+rnb/268VufKZs7CRuaKU9RMMtntwUPx34uRha2yZAbJ4afMt
uFxKeYgFG5eTh+gBV000tAgiqzHioWzPwdjeQI32Y4v4xeQUHqk1SGbZHwvTkOlmSwGqHlIWxarv
pzKRSufxTNW0s9zBEuAOC6HlRvcHu8bTv4xkk/VWoMXDlKKjkMXit82JPF/S93fANFfTvr5+Va2I
J7YGjzo1WKnHk+o8CDGNQzNNWRtwNljSF4BijnXrFaXGHPRJ3rhcrMdIL/XMlVodY5roLPihmUyO
Yy4GnHvK10578dU6BktoI9UhF8aaVVMj7VqJ4+Lz7Gbb18Do/o/sS742jb4PgCWkFQGU5OH+TtBM
gvsuX/Vd4A176aIhAjWjzzq3oJ3aBTpmLQuPMNVshnGydV3nUrAfwbuNN1SS3TpIkYlF77sTqr4m
pIsN4A1ByI0hrqiyQKLYFx818BRZZOsszF51d0kOKzwnx9MrmS0NtXlbQhwG51DjaM17k8x05Cts
4TcvcVYuE4MJZwGieecTmNhvJRVJilttzMn/2/cN95J9illqttC+GxYsxN1gUCRb5HUIztt1pC54
0k9dsvGyvyvBj8MSIebrwdVmGmljA1meDcjvCeOPiOvGb6G1NMm1kEA5jTQW2WUOiKXicsTUNMcI
m6+SwudHrWG1ccc6liA+JiDWdy3r86Yuc6X4tj3viQOTygrREKBFllS8F1Q2CwlUTt5scIEcqRud
JGjqEGM1r685SYL7rAcM/pZ2m0smnLWv/IEFkhz6v1FCyyZY+v6J1Bg5ELz4FfCWoWbjwnwoQxNq
Rx/seBDaHSZ1g/J60tuEYhGaf0P5/iQTX8Z3SVYJIf4RPEuRLjJapJ+RNR3KXHPN1p71MhOI3QSc
DlUNrpeii31N6RDJ8yheyDDtSuR9BuzngOxzocYVnbke8vGHKJo1JSiQJrt4iZMEaDXlF3iSiQcg
7JFsmBZnvHTvVuk54V6VHFbrzKnniKIdZtLP4eUAeFENwt64pA2I3y8jFrYVB4cu+Rww+Xhcg5UR
AwUgQZO2XghdHY86gvHG75F5AhjOOKSwA54AAxd8C3wcLOocqOSxP6ahybxi4xX/TavinYtFTm4l
OKZt/g4+mNe3gXQauvEXS6xoHGmNy8gAhzOpWMVFtjV/J0eoHAF435blTjDgkIF6Dme3sKb0Q984
jVG8lkWquKwjSQi2sDSZmxaEZUvrVvyqI26/tzZ0JvdCF8VcxOKUXn3LuF8ooAh9/+QCFIbIPU34
GKpufif4uVS4JclC50GHS998VXzSiXCj3W+cyfAaMwXs0SRc+Ba+2GGgpo7ed8+FkifIH0MfZy18
e6KURet7IKhUeaMFNKZ+HnJCHAPbAp3M1frTIDwV5A7Y8Nwl4kJ0fBozUuVvvpQqQ8Mmvf7FE6LA
S1aiPN0nIBmqiDK246aUc6ItzPU/3FNmMw5uqIkeyNrleej+jdhpQgbLfBkmSESAuiabr0L3K9cM
3UpwI29w3QMWIFri2sv4E7xAaN/J3T0PcN3yXDaT6N0jU3puKZTXAhaghzqR/5TUdOSkvl010O+L
5bcZSgeG0q/GzqcaeSegt2aiMTOWrUtGtpSGNQVJ4v//yJ+yfNM7b9/3rYadnyIVTtko7cWYESaP
m5PfSsFosU1wFb0qgOlOIfbEkhyJghQ51muzGBKMnVzfqhfzhIN1sw5FUzUwaeBvDnmdUUEBcl9T
Ng64nfj+4vygiy4rf0k8bRG86SdOHkLEgfR+ZlusI0T/ySMQvXj03lJcrEQsRcS9izAqx/1MFQWD
wgFoOoG7V798UrZ9n9+2lMtP+vtVdiftpBjRbcgiFwAOrH50vYOjU1xjJmWQetnPvRNJbKAG6Ehb
yMhf0lBwGxJliRQPF6umwEXIt7Gqf6SLstNSGyV1dqiT4lEOFhGWaQ4Q0OnaQ+GxuBiS8umC1pWe
U1ln2kTmO5j3qbC7I/9IawCmuERhaScMkwbLKJj7IyFNUQdw8QkZMJ/pJg/BSn5/LUrXcgZN9Ug6
oTtPErfsg8Ms8hP85eBLHO+NKW0kcruJsH7k1NkBa5tCaiu83qN3IjMl6UAeVWDtR2NSeIzI+09y
8aeV8kre8Mg5bw/tmrrreHZsDYqQfkGM8TpX65+k5dygbxIm7l99JJuoJ/U/Gi3U3UeEioK3SKc5
ZwV4Ott3lYAiUNb7vYPNMxGL/u/9kD1F37DBCfB0zbzmnxvebl1ZUZh6Lr/08r3lMkRhUpurqi77
nU9ZEev1I9j4r2L8MxUPEiYpHt+tMZImkZwmxsF+GEWd147I+wPPMwVhh2JHvThUJ+D4CdZ2Q25e
hNpBJ2qiEH7i3/VKdsvS2z8E/jxAYYQJDBJc89TgOecGHNaiOPW/JSyov2PSFi6DBr7FTjL5D7sk
/ABLDBYawkoKWv2Ow4IsE5c3GRiwVzTdNnTlBE8fQPeuSMESq14iKye+9rG5/QA27+65bGpcf+75
XDPQLBQHvDTN/BLS7YjiFBHuv+pgPP9/2V0lcu+H0+c5DeVxaOb1X6LezHaRfAwE7csTGic0YO+Z
5Z5Er345du3D01HnVR6lOtbomzlyJL2qJVnLQT0ddu7SI9K0GPg7oo5kY5A8APbeg+jol467peV9
3AwH3lOSbCbijaG4hGrLVKbVdq7q/9f4LghTROk3unNfptXiMM48Bkfr8mQBeS1R2c4Qbq1Gzsgm
mjitR/AQrGNd026y5q7JxgEZUVH/OZJjbzW1b/dkJ2m0ww0pDoItOUOGpmTNx0Xe6a8b0HnVwFC3
tEwZAODXBQ5ql48/vKe5dRMhppaEP/5ZqOLgwuy+f8adsODM9uRL5PODAFB4/OuMwrXLRXOL6oGY
YE/WnXuR2mrtXtO1njmV0UlBZcKjzOiZ3jpOTVvDzQoD3Vxcmg7WCPQnXH2LHLnjwrQmBHQ6/zOR
VJ4tjDckeY+kuh48lRSQ0wgTWBkdCYr4bycIkiM82mpD9ExBNw4t/BJc/uZs2MQ1TBKPGrK/5sGK
iVverMtl2WmgCtuADXILmSJRx605aeJT/U6fPE7ffdvx+RJNnKNJ5ERvS2wlBNyMHCN5VaK+bPIF
jMfmlb+qUxj6jzcEaSDo/KU38j7ZFnNRCfTzQmpmYdG4bmNuosBhoryfXMU53WvUDnqj4rr0B1Bu
E0m/mpZwYzuTNnduCAh4cgHAvt8BxWOKY46TRLshmrAnTTtveOWImSNHoe9Xpm8RcbjpkN+p4AvH
IEN+t7RM56G/UZBEuQ3abUfJYJ0Ps4cjjiO3xcyuqzknXcqD7Kq8nCGeFOifgc/bPLuYNdv/1dM/
J/bJOL0edonytnIRA4gwIKKdMr8lvsWbHzMljdkMaQaunOwPrrt/o7tAy3z8u8awSbkPt5E3fAMM
RGgZN1u4KJ86DIXQ+vKTX2lBJVOR4asG9Lu0pS4jVAgNFrZ7hU29WScNQ5BGYEjgOllh1ok5kKZR
JBggR9G17R3UtQv5acCe2/ZJIEUqcuvlWs7CFxju9q7bNDv3cwt/Az5e6KsI3zrNpdSE/1PMwIRL
Qa5W82JG6XXvii9/xCJYulzDVWzxs9idIPHIOIDj7r9gwklWD6Dy6YBOfi3Qp54UNOqEJpJLIoqr
wJMVM6qQqFm0Zhl93JPfjyOSkMd6DMZP+Gfe5per+FKO8D08jZ0i+kQ6U3XYu2aIfIhbGmJwuJZB
lTjhgprkYOydVtylYuonP7S+odELxqCyXSa30Th64mCeg+nVP132/E1MSXc2lfV3YP8ToTEqL+hV
xjaMUHikeK+Ulh46m4PkNj4Md9wIn3avvSr2tg71JT3R9k2x8SD9gghqfU0PR6ncyZoUbhpphgXR
WiakG/fY9DnYnF1ILVZ5H6WK11xqNZRQdmoje0UFB914xk7uOLdfYirFRNN2EEl7lDwMtvq3BcY6
Vxverkul74yKnlDYp4KeDRZ+yJFtSMd4webu/ePgfTyVgteo/7CvPCLBUILIZmYYG+0uIztO+SHN
11BEPa0tFmY4QhOkgKswx2/Gua9ev3Dojqi+RNCFH29ksFh9oQfvlkIThUKdOIxI7Jh/Sacx+9BQ
tk8KleuRLHJlquPipJtPoIw8eUf/EYfucc8bLPCnna3xMaCkX5xkrL8Utx26AXcf4HtFDoAUvN8S
8r3+u3oVn3cgv8GFRc6EdcjBXQVTN3Tr8wV3cMbIoOkpuGfnrIL3cQ5+8FkSgWm3ugfWj1M25MXz
lNQjtMyOfFgJCcQ4+u5pDg6X62Ho0ZnZr45FyezVxy6IvsLD7uuM1PRd7KCITrYJkxOKDtY1xYLd
bB29Eqv+4kpndRWZxDtcf0yp26q7dne+ZVdzFNhhgCnsYzdDd+JnDQwLwN16hNJdeRNrIGupy6qv
v25rZ3JMhgQPKomd0fWsT1162TRrC2Q28vOujwqYaPghziNpLdPCFbWYz4nkSL9/I3U3CpoigjUG
7VmsyR2YpjSpHvMXbBkoCknV40XxcfeQrvH900DXevF9zCr2amcJTQ/4AaUWjcRaMCCxWnu2uEoJ
4FPYN3Xw5fqKTcc1zqcoTGHdTwNaovGNQo044oYYjX+oA8v5fptxBqbsnn+Z5FpSxLoy3Kl7+zUZ
6Db2dMz4RCHVfK5HfQ6fgAJ5JIYu7kGY0PYK3GI8TovO4IJztKWzWevV4dlJLdq1nP0pwHKq1vqp
4PTjZaICLBDCBXS1DbnT8t48iBBexT8u9ObWEnZ5hyezO2ZOg91yci3UATU1Q11pF4N1K4HnxiCX
PX8+VBLt6qd7XkwE3RTcz1stPEOmWPeVt2FeFCMR2dYQxZbwa8RvilAKNaT5jBxxMAiMFDPOZ3hg
7bWVVH24Rz5ODQ/ie8IP3fY+EvwjmTe6rFDAmke/MIB4sEjZlY50sbp6NEsNJlKkA7f0fwKBNXWp
+3o3KhQOU1CH3nAmnZTP9H2iiSyYiYF7gMb51hjaz86ig80hakDmpO8Z1PFpn0xeFjd0aF1BTW2h
gSLRz+4YpVuq27Lsqzesb2ITZUs2V+4AyEMi2Hrm1bVlwIzY698+2g5zNq4fYMoqkgSH60MAN5hb
a5ju8KmYNlN3NWJDUZBPce3R3cspHdNSCjHTpx7xEsKtSYSXUTGXxiZ2xNCNdEDCp+v6f+/yzPAM
Rm6hJFwuJuYhQsJ9qfaJz/nZb287stFm2CDFIKuRzFeNGwnYabkrC3T6m2HNXcWZPvuvbQn/epFm
GHk9sLDkP9F7DdAc15E72DmHvdX6Cef8SYJm/ES71DR8ZigMmVQ0D5xLu3ffvXWVCNKLv+WxJQXP
aI5ahGh/t/l2xTK8bKn3vI2ndX8Rd33U64h3uNkI6YBRXhsk0p+rG2uQbVnHe8DLrzBPIulc4r3O
Cv8vVl5VWqQUsODsBFZles8Do0wMmsU85sQQCY4/4uWayjFOJi5EjWmb0N/Vbgx6/L0kuYQr1L5L
p+1lAQdD3h+UN6LTj0EHf1tLnKVi8zNV8bwsihHU2DgZBx9xiSRUXVxEKrXsywwsdAG7XZ6RIuaQ
2hbykvoWZv9TehfdFVbQwvWRAQSzduE3rPHq5j++mSxfXVx9gj/FqZctgaLH69vUOXyM3619BCM/
mWUlQav0e5FvdTS23pnlvdZTY7z0Pq2e2my7Y+2KPXQq9PQxZLdpFNY8vSNtqnCAuIlDC2KdxvZ9
XihTqMAWg1Bv9sQ8TwLP86FXz6weHr0khIVPa3JbYqBgBBQpzTVq3wqtJddujN9lkTfpEWq3NUlg
xC6J3vyiS1o2P7xGFl1YlLUAtMSrQx3Whu0kOuxfsu3i6sx1eBqhufSRUOsH2mL6KJdDE12g+UEe
ALjiIYt2jKLvPwvHw58iIqzoFLg3nF/th8tZdovk3+jBnBkwyuqxhQu+xE/n77GKxOWwJs40GoLA
5dhlUKw3Qwlla6bYwnyXND9gO3Rv4zhnCnG5O/HkNcRq6iv5r1868Qb1U1dHcJ2VrV7Ex/YFhp1h
Xc7AHWvyNj8g3u8fMh+MKFYcRlXbgIHXYEsaBaSf2UfCsSnBb4MkXlmFsJatVpHx9RaPZaspSOaz
xeIB7FA68rvH8SuPtOL9kIMjrsq9tGXD7g43+glkqJAZt63Me2LgEUkWgGPFxRUfMJ8BNlN6pB/8
XO7V4LTSB2pXUqiNx8LCOBD2+TXYw5ezNW8VshR9ninsoNxQuR9TySlOjf0fI1rHZwtKxWAu899K
HpffUPa9w2EOTb6F+gSsrH04R22GYF7x5QXq45ebRtkWkYaJYwcNg1u3z2fFV+R0dM0xm6qP2NRH
xi5UGBfQtM92libt0L0GTjNqfavo0PKEnhZA5/mjJ/4f+DKHX3nSpC4ApAThAy7KbvvmDqMbrNFV
I1kyKgejqUQyI9rXFWH5W56paSHMgK6dGLHdC9YU7Hdu6+PIHUOrhaizCbugDYKr2UGH+Za6VhOJ
smATYcHxP+oHkVoS7yr2Zm8XPIw/8opvyHXu+jE4MaBYHx4NppyNc+zBjIeADoa8zOZXT3M0wa5k
nVw/UaclYw0xDH8NDzlf3u7kRjr6cNvXNnWPrHG/hBiU+fi52QsEBjGvqS3qjQfqlx4buNrbeRBf
hwhNeRzVvRO++o48FMwfhn3sLRalMX+HuY1tmRJkwlQ3C7Z2+lkFN6eTYjiokUGgiuj62DkX/fvP
R0eLrGaeWACM5nxoKdKh9zoCBOjW0afwWEbVCwHqc4bp8t9y1SAQMTEGLqAeKLSlP1dLZ1kkcTLz
2TrNT1OyRRRcwM6q+rd5SAU5a5fUsIujxI7L/eyYMKmSy7CsIkSEhJyoD4/Z1z4SPsStLHUqVE/q
uoZlnAR0DNtKHvWL3yRBnQpLNi4SOBzamMJQ3CpYqCF9cHnzBTf6LM8a60W/3jnQuXYiv//QH1vk
DqgmtbgnhkwJpY+KxUOik9a9CngKPPytLBWs/4VWw7Jv97w+QQOQ4l/xeeQYRceMOfrcsyCeDsEv
KLitm4duoaDhkVOECEriEVn8TyrGNvthtDJ/HKtGD1ueWQyPzvVBTmMWddli5C/dU9exdvwU7qCw
aTGgGlJw6/BX8i8yPzqZJ0KrsAm5sBTlfFgxPo2Qo+mUw9CkWQ0wuTd5n51dI4bTDiRXNBdd+Gdf
VsLXJRQL26kIRzSIBtlwI9rRlTddEZb3klo64df6flpUKFxhDA+4tur7Yqnk1YXs5rm0DWGjll40
9FbfV2be+lifasyBGaAcERxF7Gnfk2HBvVv+pBaTkH5NZ93fBx0+LQ7IVxx5HA8gpekvT81ApN0C
x/UWSYISrRPpIimu8a/iCnxuoTMS5zUTSzU/hzcjLKzozLwJi+7Ns8xaBR/7f0XFkTyRx1eiYKzp
2c+0iNrVTo2NkJu/iW5K3pMQ3BM7zeV2LPvTrN0nF73o/0u+vMJukgMg/+/lqiAzsGJ5cUu9Krqf
7b3EfcojqtlxEXnvyTv6c5kn4itsCSla5bMGEgn1RFe688yPAu1gmFgnRNE5//8FF7Wu1FlZoBXk
Q2MEnRt8dxs2u0hmw7EDYs/GV/xSD4AOsrhvdO9OkWfpLH2gHq7S/4DL6bx60Fo1Z5UnPqxGeAYp
blDHnydWlAd8O9BmpvEi0T9wtmfcGVO10wEMFCcFW20qMLwHvxQxMAs2StPVa4004bwWwNVRChIR
XVkayrxoEmyOQYOCZEpzSw0mX32K3QcU/UXMonxWcSG3qE7z35gu+9yEUKq9mH8yQnMYOZ0G8WDv
e4U+AQVnN+htgi5qC/3mD+MJmZgOd+q1uKJ9ashRAlE6nfhwdSXnrFBxouBseDaqWCMO4omzRTcg
kCuXW/oWSGfsMoAKoV5sRKU8SZ9vCoxBUF5NVLQKb+reMfG14WxgdWYkSit981n+PDsUeOPEj9Aq
kGDGTDzQJyNNZ1Ei3MTw+uv10U8cajR0thuY3UPcjxZgSeY0Hbrkes8yOBaQbtIFL4byodm55EwQ
GSHGzUpuTiSOWf9u4DlMNtBSYg1Q02rtLhI90P65faFizQdif2jbGt/OojPkp6fih9J5HYfUgNyd
ZFa52CgtMG/aOTu3MrJ+J2Qqd3HlqgjlmjD90kb4ah3MVSoc2UuHJGHg84Qhd4JFZAZ8F/9gScM7
fquamdVxHoETXUktGZR+an9YFhpZA8tC7zpzoK38sGxStGY7FYDZcqEzg6ppuQtIlj78oMgT8O6h
fQZOtYnrMIE9Rm+F7zK8e6MnUADwqWVHhHcVH9BexnFaw2r2MKEvfRItGHiJxWv0beqdhJRQcm3r
VRTMDOGkny0IY4m7ivhvLgB0GnlPDOri+qrvfgKLoJsyr2EK0XtWw64ewew1RJkRU3G0teH6+2DW
DQ35kOjgXFy6CTOOQeqMPHQJ6QAuwMQ6soAfwK4FiWTKoGNTDCPEXNiULOnMVEErQzH0d8APXhqE
LBb9+b8zwPMW3e5i/XvLbLZnHPQOYAdBqjAa9NFi2H4q2NzI0XFRMvyBHCphTViv9DznAOu1sMH4
kZ/En7CoCEYtoE2IgXhU0O85PuPCcBgNUkEPToi/nQzBF+hI0UYpZ2187XEUtpdpNIvkEz4g8tuY
WwoLpmQ5QcHyGsNYDtUBJeIKNuFh99+dJeE8QsWpMGhBDeNXX28gfZSre55zj/Bnj+bBVKCeV7dZ
SLjrNdClIKmw+6/9zEwIKt+jSDn5/Bd9u4t41LwypsIPmX95QK86Wo3bLsvvHRSLP0WesTy+Ld8X
nta0+JqZQZJIdCzasSRdGPeoCOO7BL/nZn39odL0SzJNhofTra+P4y9W3JKNSwlaymBywhAZ2INt
viBU+F0JL13tevNM1LF0IGbpzDCw+wFpioN8dbXrtNFZ/DWwf0N6mpE18SzEbC4ABHIB9GnD7OrY
lNADtwu/dQj/wd0nLNVJguMJaZpXlgANTpztxGoZc9oCUq6EX4vKzQXixoIyovLAKpFzQo2S8eqt
PZ6j3SKS75HJmR7dnYftPiIKKvcJfu7t10EKEE4TBPk1BdmXAEXsnBrvTU0ekW3RJwSCg8bpr012
wpA0aQdJFynHU70JEzw7mxhEuheCXOwg6dF13+2BDwJDJ+i6Da6jjzhRJLwkusBSXC4Q6b1N822J
7DsIrXVuRyIBC6gqyKdoH6McSmtpz/wr0bgSPw/5u3OPKlcmaHdpM/f9ew8mv/epJ/q2umyY4N2O
8HTRYZZ4g2WWYOR2AQAR/1Fk9dfi6qXmsdrmpexZmrf1G1PxQQvRnB5My1WYBSoTUsrh7rS674xx
tuztlhfDYHJJ5NbDTZyVznmZTa1CjEUYtHkxQdKqQuwVxj8Bw7QoCLhh3DV2AMW4jc1CJeaix4vu
kE67zx6amRY76Fnc9EGb7IWY3xOFdSSYrUqhNMzt+M9WC+urjZFQJDnu/NiYdvPsHTUHGrYogS6p
BKk/CYKbx038PUSgIqoFwfOQzVufrKPPwNYUSx8oJcuuSP2hV1kiiJ7DlyxmM8iDiJ3iuea+pL0e
xQNk7Ool0XBp0QWFd8SOUEWPb/sMu74Q1ikDmwVtKSs4CIg68/+l+EpL+MlhjagTr257245Gdfwq
KWWa1GjQQSU8KEQPc7tzG3cHvcEHb1E7jULO3HIdYq4+Mlm77vH6Av8YhkSZWkFCcyU0XIqY2EUT
4kImYC4GXIocDkdtQNagcebJMlum4E+a6NejDPrObQeBByzt01s+lgrg1d/ybLao+MzPkR04TsC/
Hk1cGGrlp+HscHE0N0NVMVTF3xyL4e8OWfqjgxNLcK0s9gKEQq020JeHlFtpZ8rnseRyjKfwIK5X
ZVUQ6Cm282kBBVW+DyBubRWTBh3MdZwTv6zMnvyTOs3i072idaKRXAM/BceJoOTU/n9M/dsGSoi6
1A7YSyN/vydDHS8BfaQ6FoEmv3QLjdj3/sTru/MK1fpoh/EeZmuEiY5IHBpvpv5NGEn6rcineipt
Cdj/2/IB6unmAq8jo4IShFetZOCVVeT92j1qcHM5MaOSO26UTA7/9BpCyDwSX6lkNj9yP63jZN0C
EiWruTzCPaiCYtm30CnecH2nozDSzyuQl0aE04vhexUXlnz3pmKFJbWC7unYYZ4dE9/IqNDWzwsB
xRZXbLw/rH/IyqaR8HsJx6X2MreYV7v6Mflgy5/6O/6btxvcibjeKYSjrwMtcCueaiTb+p0dQ19F
diBemv4TQZPH/LoJ7QebCyPcVT12fQpMOaWd/w8BaTg76sortlAi84TchIKKer+xTf5I83fToMHC
P/usQBAHU6sIBi8WcEAaV940gZVHcREbtJHdMn5ztcdylL06bYN9+ru6CEE7hWDJK2mfdZDA58M8
hmgCCVk4spn4ErnNdLwf/6tJkNAc/WecxCud4zUK949wGJ7XS9oEF05hk+YRiuO3u1sfRKxmYofj
rxr3LeXpxIq+a+WfAUMSxc1jyk+N5FNoJn6S+ZpoBi+PCQkQaHQyomy0EBVT22Z7tgsouK/yfa1D
6KRwVVRXOP/Ci6CcaERWyvzFV6/colxoWlZSpXNWiPOzgfOigVZVkCUwMFQlhP21EZERmBSIYu2P
8QjkN3Yc97/NOXnNvzPrZns7TQ6R+zTOBtBJ3AGWzYAvyrD2gyPvgM2tIbdtwYnkQUQCIea54Ez1
tEcEsrsm4BxNb+ht7AbFfemuxV/qN0gyS7NCWpzpmsfc2EyGZ6MiQASMLKlICOxFEQ1YyC33DCvh
Gy0vCVS59woGp5wLLpbhUKAoeF9wl+v5h4opTjstjHyxejeArXVl11APgqwtVejhGsdckI6/Dfor
gwqfCKa0thcPf9Y439pfGiPi/VerdSebRWsFLaI+uiDCh+/7FmFId2ed5ExBSwfRRD1WEbLgbC1U
JrTFYR0WAq91Zy/voudCjRb/6nCYAvsG32v3Td2AkcDoveIXTUNGFdBk/P2fROzz05qqLRJE08Ky
Le2ikhxDUmUd7nDrFENrk1LDvKY0yKuKjQs/cFTp64XEHr+H/ma+OqoZy5PVmGOvTKPHM3soa/PM
X0FPUYXFS/yE9XHcv5Z4OXy5PSPSLeP6freJEAuudrjaxpcOyc0d7uvzNaXqSgaFUebX+x9QBANH
+Yyb5w7SpypbxDR1f2nZCbB/HAXEWM3OGrMvNqUsjmNklLWBbCU2LNGHlFjR00KHEQg2ZW/SSyXB
jbyZNejhiXuAZIhc0VJTswKuRmZd5xanAcIkSy2Okqvt3kYjYS+Zp4vB9QeoIVoX3BF0P7rCq6L3
zuVj8EVJ9l0o/hKpL/0BKmHYQ6TMwWMFye1bICwfo5y/2jga4ifPuT7FUMvZLk3uapYJUK5prz+o
Z2tp8TRFdP/LMkxbfifl7ND5/EUbwzEn5y/eHAjrKIN/MvVXi1ycSSF2qeHt8/x4ZGx35XwR+haJ
6LgpKmdjM4aIEXG3KwssAsPAr5wQ/N/CaDmT5IpBirIy9sqQBmyFtmstAZ9yavfM2xcyKSSzD+y0
2HBpPnm74/yKlz0f9vN/g4wbrewmnZ3JmkBIdQkVnhSxGPPVwzW5ZI/YVIQdiUdEERMqyTlAEv1x
eBmouVKASk5Die/wUYqLpvoH97ArjUjWoUrxvw5Jc2USNVbDcEuQLSvD9vCAbQ2McA+M5Y6BXzqI
LGiKXE9IiI3H3h7s+pF3Kavf59dcHGfMEiPWgOLWLIKDFzC8XaMqfVih0r7bLGNVnGl+r9M5RN0q
/qlradABdrIFVFOIM8wYgUFhrtsUIxFaVt9348TE+KRm9gpWUnSJe6hDCH5MckxB8wQQFxNkm+l8
31WEGD0QCvT/FwmBxIs53fjxms1beeC4/HiarpH4UdLw8I7rW4W5cbJK0dxIt+WlTbZECDfGq5Gj
fRnoCKEyHcW7VQevikZ5lRCyJRwUdMR/Hjuo46jvOrm3SWpF85EFjpbsm643ObJrfEmpoqCMOjYC
lIRhBAclB/jgB6zfPrCu9ym7kOyGb9oNDy78KYnvrPefPUfrnAtJN0H6DwZDjhhcFBqnGtTT5LDM
r31xdruCFKsmApNN1hMDrxeHx7Ii+BrDIrgrBm4I7XNWD1kJLW8tfwbTwexHz2JnpDRZrdFe1AZq
df1fPDnTKjniBaxaDkiwJiCZdqR+s2mAF7tB5nsvls0LjBp2bcq6GwS253yip2CQaaJGyg6qJ0fd
/INkfOoTv+cELJzkDAD6/9Sl9FiXpccxeIiJoGtykiay5+DnPEvJd+nqjAuMmppFBTtF70Ibt/0Q
VIL79vp6LMlzbgFWjunQ5naavbzWXUJec/rung85l+zuA7BA7HHLptQu/pVgjwSh2EChnBAB83pj
HFys7j/z2dbt3ilBvxyXb9yVIkHGD21kaI/El8cyZGXlEu+LJwRcLFqo0kcfGOmVPgcq5qgHkQ9w
R2R21UhHWS3rQj9PCLNE75E5W8s16735WLZogZSBjM3Xo8rbe0U+Ff7+HMvGzZFICWbec8y0Lx20
LBIWNOKD210ny7CfNvjqQ5nF4NZl0ryVCVgA6hnJSSlf+O+KdijKOfU8wwhR3CUpnnyPIBLZ8Dbw
lnok6AARU5nyN9UNdRYvorux28oUs5YEbHy5X6CiEGG4g2xBhWxnBq5ulnGZ7I7fa65alqoSucYZ
HBdznyYdXGr0cjJw3E/FAfdxYgneyqZ1fAZhoyufysrO9F5QZEZm+k4wCntnaIc4tFHK8Cpbf0Wz
udR4QFBMF/3tnGjwpkvzdhfOsDDlcEnI4RyCGUa0yykAL+fWRAZkK8aSStQtjiMQRYdDmJOqK5BS
TFxEddz4AcMMmviYKzUfejeYSoWcFuw+Z8u7DLwoBkWHOEwZLOZYBQ4xsh8tSkODi02pBTZsb449
Y0DeJTk0jckyvFFSjzp3QmAwcThiqpy/Jb45xQP3u6qpnYwbDRj0M2kwGQPTdNgin7TRbYxWF+4u
09mihetdFZzkr5zDuL3+Fp/sUfXSuq9NSymCk9a88atpQoHDKPuhln4L9uKaYG95HR8RQ7gh2IN9
Zr608134TeJwS49K52sJLd/r3x1L6KwBmIxOWBBvU+0B05BAyvxAPHDw8k9BfTb+RhPKu3F6NylF
nTqtSbA/e2D56qC0BaMl/03oB+7qgkVjQ0MG5LXA377YJGcKluRPWNTo7OPOwVeZ+30s1wnD8XKQ
GnwJnxRQldFlleRoWV1qN8zlzc9cdy90yvWagwXYoS9Zvx3h802oYB7LX0rfGkRn9O9WvA6GgLTI
tvDBLSkwV1KoQn5L2oHTYnQZm5Ytrvkg4+nnDEviwt6MCVo3Nt7fcHm6crTPNX5mJQl+mkI5wUi8
CnhSJbgC16OWN9vVhyAfDH2FjtMe/tFmSGGdhC+z64s2ce5CtMvCr8iev7XsgvmVDbVBqQiEQ/eY
NKxrbmwSbNp7k+xvSUtRUpZDGTvYcNhttfC5ZvBWoUfaLeJdFWgEf9LGiBPBStJdqb+xHZss2eH9
w/f9gPsLW8IutrzSuCx8kReiaELd3pqpacdgF4aijY+dK/zu1vMbqGoUv7ZD/T7xGOpxJMuvrXtR
cfppy5/qCqFrRv0yVbcsODN6+L/bSUHddXqeWbc25RppW24cosF+E9dEIMVmyEO6IfX3FkjJojWr
aJhUZB9aA8jlnL2rdjWEBds8YszxWpUXwWHgIZQzdYu7rQEKtCySv61uEpO87M/QWyd6IHfxlBOQ
u3p9+zWtBihj1PHtQ0dHGflHT11zWozHjNx5pfS4FTxLyEPFSXLhCmDkWhBYQvdfizZY6lhV7duP
hTni9s/5UJobqxxtHLUPrJfjnRnTo+WD6PKE160GY/+/l9hOupdeDN3G3d2iCHql9Nb+O7Ng33yO
u6uOqX9NjS8SPUezLwPg9MkjrsIorDzeKt5LW5GSpNqgvy8aK/7bmaN6t8UuBEuLaXB1hRhz15iW
ttYP14b/vb7Y8hfIzPiUKNTRXS3oyaLfaRnns3tfmqUbceRPUr6y8F2CxVUcMBmg8dpgN7PHsUW3
dG2zJ42Ad9kyxvOCB6fvdUHrkr9FhEQVxgnGfM66EjxwE1BCSSVPf8gftBGhwRrRe3hEC8kl/QOb
7wRi9hEugqNT2LZ7b4JFDZXkL8n5Gl7UTxaNrp7FFp2F7S41ZlV6uf5ZzhmJpXtPzbwaCpvvdZeo
zyqYVgOZMSwb1x39vfTxL4nmqPBnyDUvP8mqw90hYbNGnKVEJFsHXZHnbfXRn7VNLEJA5ZdquBpW
eKYXdu9cZLVY1VquLy5CaQzinm6AJo9NW1xOB9sGUZI3V83iuvJ7fEGUHpARVtwpERLruM6SMYCO
9X/R67EUfUUYsq71yOYXu0bCAJVdc03EnfBkYMpgx1TqZA9/yNVrvoZcUwT+24tQDs+zVRVSbIob
3hb+9EmFkTC1ZyBv3VIEovYqD8VzxBflOdQ2Sfj+Qp0mOeGhGRmfVed6tR16YRErLal3KewbccDa
/d2fot1Xwc8e9h17utUsUBEVGWKjCRcxcmqF2pnym69tY2iRa27hs+SCtGnyWWK2XWabBiYPgk2R
VeTVsFPp8GrguDCfE5eGmT2qfz8DW2EVweNM8QQ2UuRjmag+9lKr1L5jcoi3DyemQclP8LLQt6k1
eC/+depreETH27GzVa64zfwHIv4N+U6ePGiYJ8LKLDUtk+djFsri37tQa6yhw7FIVGGMIiXKFWZO
swC1yaZlPylaMIsKsvUyKkQGCCF9n4eFG+I/gV186/SZ0YbgP2gMDNnDf850yxSVwxv8Fw5qK9eN
oeAgekJJCInpocVuMc/hw0aWxXJGGXQC3+aNtMntEBRdjAyviboboX/247NkSMVswQ1i4htr4G/T
P/DF7Gx9C9tzghwSlBLdvs1eMWBS0ElTV/zVL3KnC5rufAuafCWWi69cP4/yAIG82HbWtJv11v5i
xiYU7VO+BdqOzOeECRlazC7cFTewhbZ0jZN3Mzz3LCwnOAuhTyKYmt3MgjhOy2ACSz0lJ344cd4v
lPAOQJAPlvgeDWBUz6kS/UBj1YmSj+M5QfoaFiUzr+INpPfSQCJ6HZqqC0GRaztMukq4jcIfRxk8
4QHEq21ou91VkEeeEImARI0/gznafcYhg0d+qN1Oi0+eOXG6jxi02U3Hpy8s97/OjNg786sLiRH+
Mz5ouvtzyeUy/Pzw554260mrlkR+GTGnG6vD1he4n47YgNJvbOcMC3dmuIWMP0dxkDHi5pGzT2aR
S22GCP7DIsx4fE/zPC+NRGpD/ZeHD//HTa9JWf6TTU3IBdQcSH1EQA+4P45MiWM5qx9eCccMTruZ
1aZ7cfiMj1Q3OSWdJod4+OmuIBnSJUB5XCJlcsY+I4cPh9WueWTG2mOytfDgxHuDuIbSMVQnITtL
zBLo6K7tPKCDYONQZ81/7QN/TAsgKE8HdXuN/y5zoQ9MMDv1Wzp7N+HHTcyRqlT7IGxFFzkYWwU7
cRwMjci6P/qaSMY2VjwCR0nJp3A19mDhqEwfOKBRNjyr/OtjQwOVp2j6+VV9DrXIh7InmRLVUYvN
5omRFvoB2mB5vhwIt2vbU2mBnnoEmjJLPVSyjP6f58Y+6KzPF+r1npwnPDqW5kq8v5biSiZv4vgq
eY5b44Ydga0KY4FVDqUS2Yv8HINC/1LoX4y4ovjX9O7PR8ZdD8bWgKL0CRzhlzWEtrqDbrDLspzK
exi+6euIgxU36XsJdVpFBRohfsVhrX7shCzenY+z8hZOl0f2QbhNAV6Moc5agHK4PtSp39L//+fi
f0ezPbZsy9dE6aIzJs5fOD7pNC+j78eWCTpBoeSVHSzSoX2mMAo/ytGg5zp5pZZoK4+rkwUD9qOM
JhyGZ4ha6db+OUsPjh7mSNbIDqYitvRbaM6qeu30XS0gItm6IZtG1MEoGcmJWCHAXWzheuj0ZIDW
aim3zcrZha6xVPxkmW6glgJveZB6OJsNaOG9j0hOGeWC9mCYbGuT2cCpy/xqdz48RWxhfgq1VvV3
e0rb1w30NcD3HvNjQd69KaOt2MN67Z9KDVuHwIaWyFUGQ/9XYkydk1j0GuL5VzPjw3noYxAD8lbt
p0TaQafTyH/79TepfaMOx8lETc4gY1SaJEqNy6JR7WidGcE1/xJoGCT+xcOxKTjP7x8lRpIoGoWI
pYA1uFOE5V220TFYd87rngiEzqvenvdj16S98uVELmjoXd0ybHtXzCCPK/vme1FrrVwyFDxx9K5w
WN3FJ1iadFwEJsViMWWkcrNRbQaHI9V+rBwZ4BNDNpkPNES61zAfVDh/YH5mymgelgyH28J/VP96
xUwe6GhpbwVjOfdTbzvGaR7N9UupsspXB76UaBRkWBVokZTbYwFMfz7glFFgD1Fg1kYmMSmLqJjd
ZbR+1NN/rJ4uGSUz/cPgU4GtbI7Npo9ORlomE/UKXZoXtdZ3dllBJBGC5DSMXi8yHKHyxeYzeLvo
yskH1vEhIP2Pyj4V5+W94LFr379RLxjo2U1Ezxrd3v6+A8eD42ptl4/nnj53o/YJPhz7Hko174mE
ghrFWrXDPz3GPM9vtI2QKYrKkzHp8WsGthnizG9HMJPIF3U2aOYVywxkJ5vTaux/F24TVe7HmSz/
1unMKcxUAdTxmN4SK7j8FTW6/hsaAdNeO68+Gm3OOPwSYVo8fejwxOdS+Jlz9GdZbQkQCGDK+Ry3
9Y/zraXhHUNbeiYVX1BwvcsULDorfhW8MzrAI8nuQBEthCzEfstRInvkBVgB9hXHe0R+iHHoJ4d1
eK8T+AQZdcasg4I8wX4O6kF+kGd+wSDAYc4lcXeSzXJrdTqizm00C/woDUdpnMNjGgzYCiTNJ/bW
Od9SP3ns6X2Ix2hswEWLcU4gh5o64IGpESp9qOfI2WlA6Nh95GjbXFYbYN4esS1qvXSnYsahMf4A
JD3LUJX88q0msR2phMlSe0nZaxRuHp66qmRaTcQhN2ttEqi2PdS3KEl/8R8FHH6suAeGWj3f5fcC
jyRbdmBR9eY5qsq8KwjrENA9SKPLxDdvwN6B13b22nnXyZ09Z6O1sq4yCYB13fvJjTgfDvaZNHGx
iIg+4R1zWlXO42EcYg1XuG9k+GkObgecFSNzUrUjFL2dNiNsda3foTctoHptbw3pGFJB3PRhShIY
G1cEnqNrt9slzZvKYS/MAw+KposjpRmmm3tCztA/UOjLGKdv+agp9pIpuIwOV3Mml8M/XiD0IDYD
nkq1SuIabmpC4I8pA/7QB0WrZyGIgj65PYOY4IrbxI4xPrN4HEn1iujbSN+A0MN+QbjbPVbY8QIq
3woo14gfGu5VKBxpLXMCFXLGb+9kyroqRsO1NWb+eHSXGkPx9tFHai52kquqHw2UqwPoASEiKP3z
ov6bOxIJsSDsGshc2OmaCHUNiVFbwVmNT7Dr8Ag6YcAsTeqEQlE94yoGs5FkvFfrGWWtpCcELMiA
eKq1d8uJpHMSCMGnxiGMZBCDas2MeKjHTSZPK6P5W/UENs93obrr3iUvRpQ7FtFjbSOKlQh/xRhb
e9V4CCj9gGGGjyvzFg9Uv49lFGr0fAN395CL+7oaM399qtV9aPLJWwetuxJXs6aKiHrXh1+XuIdc
Ol9CpHUHQm2OU+gTZ2Fh1dSAoQfXPbQ1kgZSvJuN7VM0HoKTqNz/ucYxHd3KrJ2Gm5Q8AaiEMTI7
uDrxK0/72U+2VDyrYI9FXU1tbmEnty5R4UIGZlYKEzZb8mDD4p5iM3812Uy+m2g9W5wgS2wU8F/Q
RdDK/ptBlSxxVTFm46nwY8JGhHNiPMpFzhdjNSziNtncbiCOKPfW6ednGQibYkkzOme21xOS5Vmk
6yaZebv5gn9+UK0LvbeamuWGk6Dn3RFyevVRscxXp4U0lgySKHq/F9Hicn1omIbWzQnSmJHqOAfy
t6c0Q3/xxzuOZvTY2qN0QqT/TmYGazr9/72rxkk/ILiiijlHJG1VexbfjgQGPI2Nk5s0cN2mfOn+
TgRyc0fOw7qpkqDniVZ9E5741iI8NXrU5X+3j1CdGWVDQedj6NfP1OieiKyLBP7v4xYUx7PQKK0X
s8wCh7f1TpIKic2pXJy5F3ZFZbks/qJtnATJx4tvXnuTJdfoN0oY6MtgTm9o4OuFc8LYqoOHVDQ6
7WKnhWn7UiiqhZVxzRBtOLWCx0/BoFmz7u12D1poOWZ+Ub+BeNwFY3f13J8wY1LoVpsNHxWb6Ssw
tyzK3J3vpSnqiUIDeogRfDp/Q9rIU77lZOvFxOBZnZUHkbkxDLBiJ6ZmnEe9PTW2u3WcUubc6EaA
rM60S79FHTNeOZNkDlpwXKvAMweeoEQWlygJRrhukKXp8Tr7dpJ5nfnEQBgnniIrOB3pdKDdBRdx
gxuBtXCFdlYf0RJ94MAkh6ggQzuS9KmepVTYNF8kTHvawG2irKF2qMGC5/sWBHSVCgnf9HFfWmYq
Sv5S9l6W/4jKA64haHBM7E7eliEZ/sfVW8iS/x4SWLt6OEzCVD6cp7NcFUI/65hra5MUlFOW+zzm
/wSSLqVRGCwLoAXzW7nzBMbPJFP14sC3fQWptMn/70O2jcMAXdDeyPG1Y43fTnUaRjAfSKDUYSAV
UxMA3+IGmA1Bn4IyEU9hiSJOk+D8UxhaRdVxDfsAhHH+KfrOHAEh3pdgSHgy1I21Pd651YuV4nY2
XSxaz8ZRov87txIHMTaZkqJoC87MXFyv5YNGdM1xEqmqOcxZZH/2Cy+/K+2t5IKX3kEEN1BxRqG+
YMSvsZ+dLsXQYE1SfZnQr7+MvxLXW61LnAbwdW1dlZ3AWHaJScyC7s5aqUFlrcDLGqmHdqsX9Iz9
bnIouOAICW2w218WLuqihFszQFTxUJSdt1nV6aNdFN2fcwn+mwTYukK7VZxEnLvM781W0b1Ykp6Y
H9Jr1Ym90zGZfX7Sc3k96o4UNnWOj2o+Hlq5CCtowMc2sxKrw8ZFu7OqLxGo6S7mUshhYn7i7prM
k3NjpmymiDwPHt2RM8a7Ta8eHbV3y2LEptcC23mK4dWBwqE6v1RybT5F0sjvf6m2sxjC4guWxBD/
4r9XC2/b/n7c9NOMik3EZekFMmqurnqHEx2lod/IuBpqby5w9JgZamoh1oLR1APwDtSqLaJc3Zlk
/5Jb47aciepOYhT+TNFvVBv6IahPKw4nXdM4d6qr6jUWEwaTQk+GJdkQBc/Ir6WOA8Xkt9lhH+/h
LDiiQaE+dDmx+ykgxypMARD/iVzR7gHnYo0nEjTzw8MbIByrNrHe4r6l3Sgu/lDNWPXGtFZ0WGHq
eNR4nLv+XA3UmxWzF+CfTjgWhque/DHGqcR+2Q/QxJgioVRVx+H2Lqto8uxdwsXhCU4GXo2216kw
692eLSE1sPbYTBkV6YgYN6ESN0JCZJbS8fDNPYLNlf3c7K+Fg4sgQcMTScDZVsFvpIdNxoFQLnFn
C62ORb9bd0vEO5k4XDuzZlHYDjZRbiKo4dUtRZCPcAngmVWUYW0pSUC5J5AMPqfd2yq9kN0W3LXp
qTYNNCx3uEA/7ZLMgOKkXuYBuIPl9ypdPROW3EUjJbSBHO4XreAk399HolAI2vVkpp/q6RFVSh0K
AcAODIp5tjtoxF4MGOIuOUIpAXP5Q4FTMZrKfJo9tZPETXK6EUslvhDiX7gIyTXNXnBe10xTRHRZ
qk6fOS1PHAPDIPHUlpiXkyRHrpehIT17WmWnHg2EymFSxaWo7UvvR5rUA2fR87DJeJc943INQ6Mr
uGY3rLThmecpWUPVp7/rJ7n2lyTDzWxnF4RoI6Pq9k/o2A2rwzONqjsHuYgVEAdfK6l/iVO+GOkt
eLQ2K9v9t+x4i11NVqUM3i4fa5330choBUMpE+MQZN5Wb98jVGSsBfvy7fLw+5PVwhQM6CS2mo36
IA0FdVO5+/WGXa22UkMTEy3nTUJWic+7jgrCn7MTT5RJnf2o740Sxs2i5hgfDbZtmHcFNuV2PYea
frES6J3wH01rpsJTYPONRRyowGy7qCIBD55gA+iGPDZbVxyiTZPVpAPUO/gSIkq0Xavb+AqyZuaO
DhUCXbSrfuvlVyeLZYeamJaPI2zACHNVfKj4mNkW5Nw1MrL5W5LqKcBXu+lXNcTsKMuAqGuRRA+7
oO6f7u63BlNC5nTA265Udk9Z/81UGlp1JZjy3cyJPOP65cQbg9xQwOo2AvJCW9syA7hs/ebkS7yH
qhM8UMn/FT6Igy+ffUu2s0Ee+tYEmL/gmeAOxkUbMW4TVJpAKgAclDFGZSEjcMtxFPCNSNNIcoEr
2l3ROY3aH31USvB8rD9SwtILDmYh4AjQcpjzRbKzi7Xo7rsqrjxsfISZOtD1oQq21SsbenrSHLkj
daE658S+vpxAlI8bZn+Hgs8BGrQzXURTY1XuQKXu8z/B0Au1ug9UbRN6WgGjLDNjR3BaD1iP6TqQ
X9j1OiSK1kQdR7GJYGxDyi86cQVLLctfEL6K2Tqgjd4Kl1g2chJfmxwFK4c+2bkyNCGEoVwaRuR+
LzyMWeD/Itv2htWk0i/ltKKvaWI+FkTfSiNWyv1vYJrezcijam66m3OJs/v7Faoh2+Rlg2eVquMZ
BLDse8yLjvj+hLPAx3G61MKJdf/EsjblDO/EdmUk109yxx8qtukrXF8zv73rFMsyMRSONiBclfek
Ezj/lzHLMEnUBtszL/fn8z7m0ffJmGvx52NGxHQSejqpsV6DDDfsB83rFPgEXZwOtCeTDlVKembP
n3BbCVY/ca2L7ga+iYtgUREHOkjkF2ARDHjYXrv9R6RkuEASIBLUXD5BXA4H1o8biV8OOFfrEfSZ
RLTZ2UO9ouW5U6KyetqsScJjsvoMw9aLJLWUyPPjOpTu3+hgSiQjqpUEJzREVWG+nT6LhDP2+1aI
UJNf4SUVAEkVD8+nYfbI5frSse2iEXBkiCaVBXFWaORh2psPVpMGUUhN7Ph0Gt7gWfQw6VwT/P5f
7ri/sg/oLujEit6nSgbaq1BeR9yU3GlW7j6QCI7e+6TL2r2G7W/4CInM57wwriHXKMFl+EWEwYFx
21oSbIRianZhY6a6j6hLeGV8yWq1cm5MAq+3VYhIhlYXCL1nBqDqK4Wr/xAuj/TogRYpEKsut2hV
n+gRJdbUtUCmJLxbHAT7fm8bnIhxx5xKcKPz5AoGD3fA32UgmR6eiwMD882UO/HEiIXVocdKrgR2
vjzR97Nix+m4n86sBK2j7YdVIOgD1NmDonNi/mGnhuKFtkbUyMAlmgFss/Bt1Mo19L6l/xvtc6NC
DfpH+gEgLQZhucPuEYid/WrfqX82D8YMxnWaADUFV8fWvzWQJw/De/hcB8EB39RFHybPS35LSFDS
nwYaHKvwjSvwHByYhi958IpYEfV9Faw0y+WwMEoSA1wzSNt/sDp38Sb8X9vb70fZyKCbD+A/6VKM
KUqD0qjAC0KXtJTuxNXc1KHtPA2VZHSOQsBgUtVg0ISFf9CzcZYF0vMOdLUpjGqLRBcmumYgTYdG
xb4tbmzlS0wyiJivf5d5mfMX1Tua3Lzu6eK29HSPQzQb6TQDDTSNglk85tiY71tR5KxZ6MqugDhG
XS9qGRwtYUbE5mLxOAJd0Dh45KMejdZaiokvEK4LckbgK7coEyElVqanfE7qWa1fqGEq6Hes/Bhn
rnU6z1SwdTmmcZ0DbQc0nWRJsyj8HvSG5Qz8doSPoL9B2D6J0XIDjb4Skt1EuCP3zvIC3Bpdw2b+
/IYTEQ8uQG0eZwn8ssLk66d9pSv2TnsdfmZDp9QJLuDWJxWECqXrgvA9zk6psgr4op+a6lwU3aTX
rWVDUrIHnZE0BI4uvUNNsstbJ6EohbJfaJ70z5Qn7lmK+oZlaqWlJQ8bKSwM16EBu21QcNSVMpHd
L4B8vEXgL11QF/PsV+tn0YlRSmVEgP9roubQMziMamM25JwQkFBJvzsE0XlpkQTEMURHvc3yJiwY
45M/s5OBt47r4GcbIDVta1/D5WgEYCdpA53eWOi25wG3fCoRpSi0auR9AkrvUIaQn+DqASF8BwdZ
0uzT5WT6+DxPUDODWZykCp7jJdqzoyacAjuzVkiB7P4bGY9jJDFK/CC+Kv14Yu4uMylGhF1Va1Sv
M0ozECrpsHa61EGp+1HqzS4rTMpVpIgJQjEQqfJ+ASdQayiWGnR0Ea2XIM4J2qJ21bxS9y3WXUgS
rWZWWxwoIGU50VsxuCIfYTIo6UQjttiQadphAG1I/bxB1CGr0vMVnZy36fkY3pcJNVGFQrWXI2/u
VYLN6D3J2wIE6MAUzSyAqF9Dzv9WLQ9tO5qU8R07nQQWc71WdwFIQnQp6emvZLwvEP+43yLwPdBo
qp1Jqhw7FDPdLBTW3mtlL+HuIsY4vd7nzm5KhhL2Hb1iaIQOXHywnnaYqQUDjReKK9Gyq6CdteCI
U3SYHdaluSD1IX8isLoRFFHJa3n+sL/MdkjOOuu0STN9R0Q/e6IQuSYvPG3635RRE+syFWblm2JB
Nzzs1CYQZQ7GuUGTxTXcVkqt/LTsyE7JkzhBHzbfOFgf0xgqpmx2265dxRWYjQWKPwVaWEAvWMQH
IwNwxKo8EUyHp1o+QV9AHnDDRt/avmSgCk/6yyqAeLEfklWkFUxlRoD2Sp8YT/TkaB1Rbk0/S56T
RYzXtoeYvjpSneqavRATXfSeWJhCKnO8k+J03NBbUcKEBFl2fptBUmhiDLQ68LlVUAYxdkCy4qew
EeDvcoTeVZutdXyQH6RPkYpRbrz4HMJRbsmXETpMfUQT5SvrJbvPgKZoXkUmeDU44NRkbt5+PF74
8tq/h7pJoxUpBgHgvQBDOlihdyVSmt1KaudgXxbC0f9tUuefMFIoUrrtbgWh4NZT3mE9dZj9V3Yn
eM8sWkDCryjHd0JYIoEXusTCcoVfsI+jaI/kJibGgXwhBYHV7V0JxCH+jzhy68OM91RQ98qIYXCq
CYQ2zeHgqu58G5uVWhFvS6gX6IocDYe6WXMTDdToDDS8vDt3Xqy9DCtNOg1LJ2jXGj15v4NTdXgV
KLgr1qL2NDZjR8EZAAFPLZGDIXqLISTnJYKeb2o+Kgpu7xeFWPd17elT8nURCRq2wFutqPRuU+4j
+E2k1xf976UZxJ/2qbZ9ZyuK+N2GmE05v8etlL9D2KDGqVtjCwzYxZdKbX3sZ86YeoiY5V7n/GiS
4PnM5CvlqZIhCQNyj0sIKGF56liUMbDyV6eh+1R6teaNq+Hq65zn0/Lxj5Gl177Rsi5bDgXU2OGL
lwF1lDIKZywdXxqZaAJDRmn6GHONSAcbw7EXWddz1u1aJvhI/dB4JFyGj4nfZp7pqjCmq7s0ct3f
wFg8ywFD8Rjclz4r6xeVEHriKxArbljKRWC8j8JSKPla6VBQFEjH6Q1RQevm92z+tuod7Wz4QVha
xVmneAuIC1VK+Dwf5s8PgOliXqD1BtoC0la77VZf+AOcoi7Lc1uy3+bnv46rpPQ88jGQeY/QqqJ/
ncRN/UAMbK9xbLbu0TEhKXXHXxwd0Tbwk+pBvcoEFYMEVI1AeoL3vlQ6jy3AO4/XUCFcF4PCdPF7
LlN78bxIAZymmMUxAih81KvYX3YW4bUEb6zwRDHEhoWaRy+nxtQBldTWVO9yrYeT9G2ttxJoY4ji
7Yqj9NbIZxE1rVl7qCoOhvjSMyF8aNtLbU5/8WCDIK5XtlTXPgAUpQzm6TVXD7Xg3UrcC3C8ByT0
ZKS/gLMywS190rY5roGvqlFWbTTaBVQIGDTfG3klDRFFVpYrC3nXubrq9Uclei2itQOz6rHJZDPo
Hl1cs3PI8wfZT4Z3v1GwKjhHeJnC55xT1d+1lCgdFCR2OCSkL95RfRyhA6J6s3nV73BD66uDmINq
jt0tU9e8jU7FOBGt07ca0v/P98htjOABhX2K1wz5cu64Vrlp3rp+ROp3julbTwiUc+RgZcNd2FBg
bg+ROjuVnuCCORJyH1LwQcOeoHIutdXoREFatPLXVxOt03rmGsSoQD+DDqC+Tz6ykIAqGynXCsrz
8RVm3rum/djOMlnVMlqiiSYqupN4GjoUcEPGe5D2yDVWFg/81kNpcL7/sOQWDpbq23I4v/diZ+Eo
NYMcW+Y/TjEn3SOzUbsuj0W6QIcAzm3ONGNLmlU7h5cOeFcKwJF2/5ocX4SqPd/csZL69QntFjtg
bv+80Q7xtLkW1ajH1mp94tctj3mphVZ33zoEmRfMiWzRZASrq/nexT/BtXFHZcW0ZbXr4iEasTeq
azlEZFDbssrAaiQZfQu7d2c8br25j7rIL4Rxt4UHU42Eb0kCxpbjKmdU0UiEl2MEBKVwo4kR1Bso
CTh0NK0BDdZlgtXnilBRq5UbEaGb++ry9N2c7AL0Cj3u3A+JuepjDtCEuR9BG0VrOsynmO2EIBKw
kdjidPAwSHjFxMv99EBNdajFiXORgV5HuZdTOC3TtV7imjJqWRKfFDLXKNUJYbDFWiruq7Y03xs7
gB44pvjTpcx+tiXig7TVgseLfuZ9XKwpazcfonQFmWXumJxl8xeKxDtjx7l10M5lyGpiLyVndQkC
Zb8YXRgdpQeTozsjyMH2C9dOjYtYwJdo9px1aoRYo2HfEkCPlzPsy0sWpm6MkewgNXdWc07YO7Ql
GdEaMCOFyuLX0d4um/LN/MEEdrv/pgT8hZ4gkbYYpYcJd8ozaaq6pOvRbzWFUeX0qSmc6W+cn3Hd
/5o4tMUkHbK7J92AnW5BW6Pjs1lNZNiMxRqEEfN4CY2Kcg1yMCwd2csI4K/YA8OLHt2ycq188cYJ
rx9S0OGNyn0tkTk85RxB7l+uKfKE7rzGev6SICU3yrnjhgZNx2vahtLglGryEGpjFIs0uUbkeCiG
Eo4zvWakNIkK+MXQRDbopDSogq09nMBpGugLA5AjXhhhWlVagKubb0EXwIt0fTUSz+ch8/9d2Mk+
sPBc8ktCm3D+9oxImDFfzcd2Boh8F5CrIzS5+chAfSZ6V5ERhlia51x85xNbF4o3ktCGJCguEW4F
6EXICUiQG2aAbsRQ2dTg6BlLjeS5rT7qVEFSdUSUHGq3zbEUE/yfvizk+SFSYFT9cU3L9BpZKStE
SY7cOPMANvkhad31RumXQKSs7j+4hpFz/8jMusejiioDWFuo/eormA1DqcG8JEcNYEl3xNOJ6trn
m/Ojb6/GI6PR3vUFXwwBjmKSTsxhJoZOD2pyi3/KWCSZPgrcFFX2wFDbO8I+b4KBK4X1Jj+HNK8P
7nk4ZFT7+ZVXLQzUR8tTCgFcgyM2Npk2GRc80pMWKV7b6hyObSGLXVyBtiYzndADkrcOfspAx7DQ
GBlgvNYsO3PuEKit8QWWkm23qzmVlhR0mjklRdN6LOkgrNvcfmJuRTxDnzubr1SYYrzZA+aYwP/L
ihIOd7uTOBtVZPDoU8+BpVE/xb+aRKYB0TwA+596cWqrc/K0BUN+CRlBpw84OUD7VG5oD9EPPjQz
CxzGr/tE5njuZDzgbuUBjx3lvLtxkbzncj3vNR5pSVD5QBIPExxqJgZJzK1eRcXxPwUUtohNpmLX
wBZuaAmIBJrBkMXkZElVixwykeVC1IhgVqNmXU/xcf0GYE6jq5ziTh7pYKj1IwZvyNmrzEietHm/
g6RGYcd0x3j2iDaHRHl+8hn7hEDnuLABEWi5iaAemTp1DKjrGVTtsOXOJNZyl1FALLW25LsLaFbC
7+9xAkqWt3SSTttmkwAYNL5J9+Gsk44zOba7tFebrD7znYEDk6/gRYVLNzd91qOvnC1/FWOO6/rw
O7P3yansY2nU4POkvKIkTyvrlmE17gGbS+LhcwpQbHpjeZd2AbF1B4jZQ82fTyxrffgnRJil4fhE
Mz3tx5Aeqzo4NycCetRiXNo8dGwQNmUCeWoVGJevD08vXhhcXh9ch/C82DX9LgIgWlq2hmaLlvn+
1s0OUwSGGxaQfhn1HQgyyjRzUXuKTEfFnwHgGQn0W2KkJJo8q8x0YHh7W9qEX4r/ehfZfio/yGiz
ostp8LufmDc3I5z376S5pTmPhWjWc9UlaVNUyzT8HKEoto4rfEtQZu5lSrUVINXTlAwr0y++2vTu
BlLbwOtM74hJ85WwGYrpXMy0e6td+tV2VCSAuCb8nA1enIc1KBFpGgOdROWApzDrwB4ejjaE70sx
RQRViL7z83LY+CkmMOs2BcoAoKFCQmO2rBU+P886UV9INZkXLVyKbQZC/zz5n1es02igN6RqalMu
40JCSHBQSNio9CP0wUbQMywqqABQEqnpF2SJDMYl6Nbz6vRieepzJQyYUxNzyD+EcV6PDgsUxSQN
cpIlT4S8pXl8eiV/6K2tZjXzCBCZS1ReCDEg58CUUPOgTLX8LgD9xHvA1aSE9wS3gvZAcWYKu5su
1CE2RERXTD/G9dEk8OKgSlCIGDt0KhXBLkt6j6zBn6AgtPcFoV2UYRB7F5KWyahhnUJthvKyyGyk
g6dzvNzS3wJct1hxB6Y4xeIH9YCtHtmI+yW3nas4JG0JaxzLRGAzONhaMRo1GeWSKr9dsdGYV7h6
cYIodKTXdgi66QmQFBFmcKHXtNSHj8sW3zir2PtdJUPQN//23qUa9B3nq6uzjZkPUdfY7BhnJ6Aw
5Usb2BZ8Ga1OMx5k28CctwWAvn2MRtczw1aIWMKdnj9sJnSTG/rkwJkIOFmHdKw6U7O2X5dSqapn
X9O+gvVEyFrnwFKi/ls/7VbbKDha9R8UOm5l9vhLIRxj/eojSyxsemnpxhPIrI/KJLL1qLwmJsEb
5IPWqGJxQ/M0Ms+W1MsshwxrT29b3ZJp9LTa/dAYxAP+ToqLLPptsYyuVMLIfAdz7JAIdP1KUSGm
bIoXGyubjn5hWI/yPC0YRoA0FSRKdkjjY+tpSODRiBQIzmNof9b6lCyilHEwSUxe+MiiH3BlEwtZ
LM7FXX39cIWKHQk37WQwOmW7aMEsmXr2VKtYHg+5UyUpQNljdtGs+5VyLLYIPWUyxVOpx46AXem+
q9YgbmzwMX+eY4Dq//r8utkLwJB41ds0ATT0Rr/5S0hIX6t7wLJe9SXvdQithBP1XsIf653AaX9P
GhAO7tYVSnZJRsw8De6NFuLDR+25JvMlmFUj3rRuNmFoe2Rp7UsmJaGUVMHoYX/UF/bFapgaJj8C
Z3pPGMhfg8xjPhwmPiM06teFZ6yv8m9r+yg+9SEPKdsEE7Uw2iahns8iNAG00TgWoH7l3OAho378
/Xbl7o5f5fiJL57Sh0G+LHLPGDyQgRQRRVh+P00yI72o4+mWvEZ8BUg79yIRGpWWTfPfvlV8M7JR
KOqNhyeYwhc6uwUjiiU6hgMzMtwl9k0SJ56HEq1WvhVAO7S52MsDuRIeD8fFlxv5GvEk5tkcy/NB
aQdQkOLtHx47JLmk0VKgP/rDYapGdurypGSR0oqieWpVlixZGFbwGezZhMqE1RdXIQd1rhwqWtk5
+196wYQxaLKKwEGqRf1xwQ3yrzSMC9PtY83IwPGhIppySTtR7I0W5MbprmrErfjM0kUJj0oTR4eB
ZEdg24Ol6St20Ym74zbCC4zuk7QTXYg+BYG7vDN8cGrtCycAz9umLxg5yRzXxUY2uDfuwY811lC6
t9D80u5CVCxAF6eCO2E1Qh+E1DUTz7suRNzx+KJCJmH/iK9/cU8XoZ6AF3ExBXI/ITZXOubEFACa
rR+RqYjHy3Vp7Qp8+tNp10XBPqdG8ZrGK5c/Ctc26L6kvXvs1Ry+sAQCqHdILeSBN/2JeiMTaYV9
7LKzJ1TM/K/m3Ff0dmKuC/B4D3nX9rsPS5OOA9crMZx159J2tC/Itt69qUEKOwns/0GAo8VJ2lV9
+V5PD7j8rTytzheBpRpUHpwwmu6Uwv+pJfYkif7Ou63T3R+1/I/pYAbIkAP/DhOEL6sfXRYXGBBp
99Xz8SPBtyWnTtk1UQOoQs7cGNIsyo/V4Furp4URHhmRTigE9p18wrET0H1N7QfAIcIjN9BQ9aq0
0j9cBvrGAg72MQinFTzTzp/U0om69+ab8MzIdCr3gX8CboGpsBZuI9TUpi2clf9IIfiDIDmWiQXI
blUmrkR+cnzVp/UOhNaTXI+qZC1pGUUwNNCH5JIP35DOxqtNBX+QhppCh83746imwQb5LXlyWajO
GfYizkKcdfUXK7hi6iZmMfTTCY8C0Z5XWWKWt0vp9jbw5C3X0Bf0ZYonCtUHRsxGdzBOo0G7vxKT
nX9Nb9Y8ndFF4t92PzA1wHNUvKUShcuArMX+H4IB3DGjhyRNJ7TeOGJWXKO/ZOf0WQOplkElQ7Up
aYAXjzG0yFKfTqbdZF40FVhMom4NfAQTN0/U0i+LkeHOZQOceybBMLVQRMmAzS5+PtIVlztnES86
yK3Sos03VpaqPAx6LOhbKEMJIoGF9ud21p19KtFEIZvMFPzVYtnbGGIZEe2Ztvuwg580X6UrN3h1
nbheFHIUmK3XCpwvN3Sgnbz/0qiiyDNZeRF9Wyv0QfR3610Wff187U4VP7C2LpIdlgyrUfKdivX0
bpU5A4JsA3XTUWE57/jeAigP+Kuklkb+Ex/KmZlipP5Nhj/HbOlXICSjcjAvt5wq/Srqt2uAo0Id
Moe1MgJ+rJMmFwjMR+RSDasnoM0NlA6Jkdil3LKlzdJQCa6lqPiW/hinpocrW9weR7hty+Rwv+Qg
qEaicaMJNsau5coQSlAzfewNOuqVi8ZM3TflosvxKutraQCHEYnqY2KUnHkha7vduP4bFv5WH/wB
/Pw19+rjevWbZ8h0iX78MIMrLctH+M+gLy43swqVYf8NA2hk0DUbdxFSfS8zFDAD2zftFJFcjobY
gAXnLjTRYORv+YWMSRNBcGEqFxVvgMWikzK5wTsBEQkk1sbHaUKD2SqewKbgdGmivkNfvoR6Pfa/
vW87o7LBWDBvu8B9uK+jc5HHsoLj7LfxAv4A2P350VoqwGhUifPr73cbOGPfNI+pyXik1IRGoz7t
oIQVjluMbJVZpnD9+PevNwOn3LVd2/mU7/r9Jn7a/9Rl/GgBZ2L07VjXV/vQEkJXS75KCOmSs1AB
BbvLUTQUZ60oJRUTToMbpYrBseVY3PnOpLasAPQDKrVEoSZMpwNofOleLQ//Q7bhnkqGIUMkjkCL
QzUOvJOWasf4OHXPPfdjoJEa26zJpz1NbWwyuRXPYNmbloUSgMJ+pZW7Aii0+S92R+R0JL1Z8ifY
YaLfLXeR1VF9bPwWMflpXNkj+vSz4X8CHH8DabE/3Kulzg4UoPOTju3viPE8Q+iRfFOrLAydmVxh
fdM9KWg0rx7JIITrzsBWpM755ZZxpGcMFCypB1HOlepFzbLv4eXqVTCg57qssJdwthDNMJcMQEoY
ppzmbo9gxILodYQ1XriqyjAYhyX//xccN6D4mM3NOu4i1fuwkPyFiyJqydB15ThYyzOs5tpX2ENl
RZXgMuT3NYNRc1Tfem182QLDUjZxueFt7YgpGzfmUxeYSTUBvOP93H3SrFXCku0zSZGMiLqsS2cZ
2McnBGABOVjClvWnHlrnbJrSxHpAifgY4TcE97MIkOBHbzwsORCHkiWzZSPYaftt+0ea14IbIJuu
W8whEMougHDXvn7FD8cofJAOIcvGH1Wde8uIonLkOgTFzPxU0Wsw3m6WD0sf4711OIyFgi30QM5H
RHzOea2G+1acqiqrQJuXQ6Ec6nLZ9Zqr8kN9sY/kKyp/2zS4dBSuvwN2r/bTRzkscYNLyfqZml67
Wl43CMjskrVfwY2tXtV14GPllZkQ776fQSod+AYMPjf7QMZbvYTsiRfE7nVYUrHew0Itm6MkKaZM
A7dxnBGpsHddXA9YuJmK+AzHYUoPfy7wLng7S/y+6LFOm8FXev/LIDMCFSXMCp5QZ+59oPB/PHas
b0eEWT3ofKD6jLxvQMyyZdLkGuwlDBNS7kHVFqSFRs03lrOPjOosou+Q3ds0qn8gy1I33Hr2DJOZ
BnEaFDPGZ2bBJpzA3O3IrATgT4qxLvf827WSCroSpdbsTMbS80J1xVtst0j35xJFe5Jfq/IKzGOK
Q5GlDSneXl4fo+z/5w61069664wkEUeovjQ425DT72G/t845wX0mkb1qxS6nB4+nCK4R4vNeKtDg
/yTaxaTUBicBMwQ7UBYUlUSYzb/4u1MmbQSjSvBah3slOcUKmPKvR7I12lD/E58zgn6gNNEUtXtH
qAPb8D7z1X85nN83y8Sz67jEz+Scsjdt0HPCNHrKjJ0wqTB3aIsR0wO/DloLyx8eIE/41Ou9E6fb
W7xgFqNRoPnkQ5pVV44iYcKLPQvc0MvgJtcHRt1gEJBSBE4Br8mBrHfGKXSWSyDU4OBAGy3URV6j
22wlYJQr9z19KMKNLU1f3RH3pHu72UhfiOeT/Ez33z244iuh8PxZXNO6zJTia7J+f86s+ygDxTEz
nD/dHClW+DHQwpwRaHs4sPbXvSvqGlU0+rHxine/MKG7tYTeQ3JVjSUkVYZkPTJcYHMCHDb6WE03
qZPP3YhaxBfc1Xkmai1uyVayNMvmA1D8r3lVxTTMqn9GyGYMg//emoSwyzwLsu/PJv+N8to81c/B
fBeC0GCJlX3y839nm8hPacrUyFlNlsx+k1f3TQSLOCM3/xS+x/Zw/8Nq+8IhJRMhCKEhx2jsGw0b
+BYc7KxTQyffbtSDn+/a9o3YbmACrBbSOPllBNHyIUAvlBA7fRTUHhY4Um1PISw8DCB0cHTJ4mJt
toW3LLPPwO9YigAEvfUQ+gbUCK2ztS+VtPjj+WAm2OyabICEcmYpb+TJPDYt2t7hk0DWRnVOVzYS
+N/vV6xj/VDJCQ7Y9JwZlV0mVeVe6zT053IhTF4wXtsX4/ZZcNRQ+lJWSg0Lx+llASNDsED6Jd2c
eIy2HqHA0ltHQjYww5t44/wszX5IoCNAzewRSUXchcVWNUUoayyXFerKNG72wXwPu7FAPal+NICn
ry8ba/R9n3i0jPMYRhcG8TVbTqa3CH7WqW376AfeltQi+GYsh+qUDX8ZTuy+cWQXufuBwXV32gMe
onk0LubIHeXF03fIxtTTH97nH0lZSFJ+9k28FSaZPleIKl9ftMvZ8qz+c6kMTmUAC2wLyZeivwwA
/JQBkOI0HkpPdkMpHHoe3mZjs6tNtCv2LfVc9aSb4JPsAXDSN5Qav2Yzxz2MfCCzt4j1JaKZpfUp
TOCugxeXpB5jdXGpadt66rJ2I/k5QHGtcUUP1ccDoueZsZOFcQBPqe5PW0BhZrKyNSeDPz3kRVOJ
VXXYsG/cYrG04TYBzNAE2XSeHRm/VqN5FGlJZ7bnuKeVO4qnCboiAGA8ZM36Gx3vok42m/P9gYIv
tQHDuD8z3LZBuHk0puACLhh5uiEDrnDMK8yAqbeMBBlr42CAFzPDP5JPJbA8j9+jpcnMUX8eyqZF
Ymip68ZrRpVpHEGwcgock3gAtvfrNEZCXNURUDcvZXsp+iJbGgZ5IBzBwOLyIPK8ozrRSC3GKA0Q
V+iANf18BBdgf2z0qDicFzPXKw4hQbQn+eHM5Bzvs6JuW10X67nxYP1AMEpV5NhYe/7ObGvmsh9F
QyEMWuTfjUt/lbNpQEhnSBDa/1Y3+XnjHeRcu1PwO8VSLVl98ipL/R1TJE2YjQaA5jq0lKWFo8NF
sDmQHU9fdqAr3nkimQbLlaysmwlo93YFvVEM3pVyOklybCBOSF7bBnhjgXQZsdYk189adAA4LlQQ
pwmqJpB1E2xHeD/6vzA7GAbes6/CdOLl/aNo+1TfKqbE+dXOSmyrlURftJVnOnHxMvQO37QD1njC
PVj/0q8a8E+s7154wGzw9vWK3dfzT2TspIRMSDg5dcyBlErKhj0xsJ6jqWdK2NPUV2W301i1m7f0
dFEKTWgH78hjEuceZw0b/vQ8wKfAByUMivu7+0Hvr3C/yr93p2cOXGfPKA3jAS458TuGnBxqJ4rU
CmDzkUxL6YZrBlmGSL/zAhc2ux1U4YPd+pMoO04OWuhlQEch4B6Qw1Ll+9UmHCya7mMJkGRkT/Bv
IzxtzAlXsjhkQeScEvEVA/OqQQuD1kv268+ih5TgaQbWAEWJaqnUgnoOzXdUOoIUOU9Ecn2ko22N
le2rpjDKUU/gd0RL1vlAk/X2aWeTMlgUQcAZkCbXGQhowkE8X25nsYpBx/ZX0bJB/tc3tRgxzPRz
mSNvoeleIzSvUtew9RfhnwrknBPExtJswgQE0yb3BAS9YTuIBFshiariSk/OEvZnVLRADQNia2Sy
uXmdUkdcgxZV61XaJSDGYPsdPeSQEtmAg7apOUN0xbU7YnB/rIr9qDKpPQeBne0qB5x8nAOCY3I8
WCQcT2pvtKCRvaOJxV2kuKdQrptmKwR5T1VQCGbqxjPz0AZ9s5NyaWgr8Ok371oiIrhvyJ8kVM+V
5Kvzk5hq95iq9RhqWx587or7z7EwJIjlBAi7Vo5T9PpzmyxZ3V6QnrPutoC2N8Hf4XEC3vSGtFIC
K6PCXX84Vui6fGSRq95q8nqj66J9qwFXgAXyL8N8iWdA9NomQytDC0C85WjPJU+ps7aRJW90sdXH
u699yTUWKXVQzOikU+FmPUUp731eYBp4d3/r2VJhv9+GHfzfB9a27sfv84DeMpsKLYhFruZHLQg2
8jmy6wvtEcA6ECDj70aUaaf50+iHrQj+xP8Wbto2G5jnIEBcsptjCZVkCqxD/uNEkmjupWO261/U
sT8jM2rcaNNO0Dd2w2NT/jC5B5xm6glGiT22ITBiLrW2wxJQE9EAQK7TdarupLzgV5ncClQUtEWc
18ZaLGoj8xd+joE8YK+KpCYEOzfReFjzDAABThwJevyuRLzCNzLR01uyoIPDyaG5X3cMjJ8Vhny3
0eouL4CEFwNsy4vp5xvj7ibNEYN6HZAeJcNlcUPa5Xu9qEPvipc75o9Bn+ROQVZFRYs8GIxA/ezB
2Pb/d5cW5zrfC7hVgNkr7hQU29Fl1gYpYOiC9MJW/Iws0WwJrRTB/T64qJHyaZmlhbS/YENC+kGw
ndDnfOIvxAi/AIERrFKhIqaWqbihP7Cq4CSU8r8Be25tYO5nkBbzG1etHZrTICp7oMMWrYvo9g58
POD2uN/MiAo8dX2G96bZCv7quRPBIJIB2xij57hjvPpqPXxVuRtjUnVr2FZaaVl67jZSR+tmBeJI
grhqd5oMBot4yo3GqDCKfjs82PwLLl7H9aVtPryn+bKkcGvBqwrLWEN/FGJ24szjLCiupjGwm6jW
qZwcKrDex+mRKsHzW2VgTwGA+WMSy4y9XHvPe2Of4mwWhZA7sRII+q+JHQfhk6KM2daUbfY2sNvj
SaWz+Y75CbFumtzh7PTl5rBqdtYA7IVyywedZ+iLScWqdqij8hBkkw+9lKfPMlAF7wXN8aNnVkWR
H1/cpvXBxYpRjjgbZOTdv+Sfh/dfLluq3glNcjzfrGKabukXdvAWUdnBLjxqJpPFagDkhMeJkrtM
fWRaaaHg86tgxosWxPgpmse7O30nyLqzcnxOUlUETgVwSXCik6Jd7JYNfsIrmsMimjfRLdez5Uxp
Zc1DG7HXJRc1SdG2l4148PEPsTFpUVavBNoop2Z+/UIhdY1ldehR0RSwiNzZFxp7oexkY0a7d1oI
lTJXgBYwsRBZPcINqcWRQZFZNlqpj0GZYlaCOfdEtbA1mXKczdqUw5EgSVtAuHzqbQ9KKkF6y7+r
rFZqKgixsyoWOwiUvOlkagIV8DLvnQX8Z8xyBw4Ls5yvlsAtHIBepHGTqOZCkJsubx8nghYs1014
JKvGL1SUaiEWwGgx5oAgqgrKaudxYOvox8RxZb+xsWeksNrhkvrTHOfQ63N/PwZgx+Vj7BPvNqhU
AgVgKdNrsMmXRsNzB1hSoyua0Im7voC27A3PZaWkIxNWhjnTL6yfwsN0LC3qDPj4sg1fcV4iWQLG
n/0d50TxDu3NS2pVOQXWoebO346Nf1WCi9qi5tCvkWYCOwPOULDMjNC3QAiz6Uca3mF9HvkoBKxN
dzOaXvx//B3P4zX1yUzekDwimQoj5PvI61wX0NU174eeld82eNMFNs3ncxsGgRhJK2G6R67yAm6z
e+RJfNwxRP7xtMKwfobKA5DVCyWR/xisSc5isAkcgUfICRzKXBaDlzBtj4UsSByybBKVjHgXd4rQ
0y+OPAuvETTDyroasPUaxu+1MdKM68FQQes/HsFiYoTe7R2n4Doqr70GMbhybOrICHa2hE/JwbT3
xHqXyXJ9u5Ve707DJf33pl/xrz7I+WmacflIfIxpza1WDdyE7b4Jl40S677wCASpUg3V3C1vG442
z0H8M7k12/xCgx6lfhv7pBon7sNlGnE3UGOCGuWLhnXcQnF9VN4wIoB9Szb21tC6xzC98jDXsksx
L0FtTfKxaKReCKA3JVe37YTm/uCR/l5H8PWCk6J76hZmAmzkgMqdAV43g1+NT1gMEsTG0rhWD1TF
bN/d47s7Ik9cP/RxZxWrA7i9cSJahaynyhSPwfvAyH/8MhuhlkOeqcEp7rYrlRvUZEpBNn4ZX05Z
Sdxkb3E8mBU9rCxeu4bX9UsxZDx4R5pv8tzKt4mNPyisj5ktd7P5ko321XFjhhcttQ1/Jcmi8vx6
43iRBc2opNEBfgemRZdTGswk4e/u5jK2voI9JalwvMXUbHWHw1NtbMjhB6qiTYnzJoanH4K3jlpn
7bE+sBAik+xgf2ATyU/2XOlNKxKYK8vmLpD0ZhvgSb4YMyCUmHXijbTvmhHETer5LH6L6UvwUbwo
CVMTveihXFsYxDRYhDU7GGz7+QvfHvzBsxxCxyKi2HJH+llVLPcBImZVVt2GmC+wL327jNTtl0QT
eHAxL8tz6zROTc6BqQiBhMZyKrMcTnD4bKIbqWR7PB0U4dvkYX1h6VjJ4Bkr865hkm1GYXBgD+OU
ZT0GWdFOFSBxw8zyCLkFHxakJ+Ns55CIB+9/9RvL0nQWWRESJKmK0zZbVwyDJ/B6qaoVdxft8pdV
FAt3ez2Ljjpvv0d0HGrJh038D1fQ72eDR9Gql2iWioztXTkxZ4mzpUFPy1sTXJ20TinmRwKDfJHl
CfaTLuvGsv56Fa27Fce9lELmS5uU3KvwqDNXcuoje+jcz6SAc5MTw0M4Uw3ULD/Wttf28fO8D1/K
siZHuZ0yUZq72mMVMqOfeNYLukGZes/yAqcp6gRK6UwgyyRjkxUJ/XvIkpYfSAmlUJOxdkTOG5Kg
35ckTqJTOhdg+pa5bu/t7g8yCXrHKDvHtca6KXPUyHK9jt7NofNpkejB/fxSfBxWso3YJrTVf8Fm
tvd0EExZXzB2FBqylgVO7AskwFhGhXIsUQ+8l/uWUpzo14HiWv856bLZiwb7/YvR4c0vJqy+mpVR
SD2LFjSvwY8qBaRDeAwC8kOLT/mNWuPgCAHMVlsyHTi/hahCNM+vsJm8fcZWzVjhQeXQHmg8tV1g
5s85PBbSrLw/vZVegZYzG9JbPNlLjA3tBaAu6t9S8j2OJ+knJUbyvbUubnF4gH5a+e8sqeu/FMSq
r2pWzI7Q1neVLl5l6+YWQtre+NrD9++5h4Q2w6jDU6KgDeKE67/GEKf7E8J/MjvFvxU9pQ/9pgbz
7sVWxynFKo0lF3oYUIMcgQze/7ZUCTNcC6mdMckfX72OCRNSRCGF60k23zkce3+oNHXji0lg8bLQ
ZtLjB+4Z6+nDjQwisG6uXJpJPWUVVh4g6DMgp0ojxTDvx/M3CP18zbihOellOihGnn9vB+8F/GDi
+oCFgKxGpj31Mx+VUK4bBQq8QWFGuFtIwuaOQUFcogONFytsb83gs9cLgzcg2+eV5m57IXvrWsPB
d26ey+LctHz+vYFKgsDYXSuq4A2gIvyNrow/X+ykYkdpgMcwsJxUbY/E500Ond0jiru6MqHzdxuv
EDH99TMBPXKajukrA/CN+2TPcwXhUDUt0W2Jv7/GjFczFrWv8faRAzwqOu7NMq0GJRygBgSRfX7a
7fdxb5dmFfcgsLIRmN9//7wOJ998XnTkbfclpMVVoY9aOO1I0ObhgsikXN7waB1v+XR7l7CBvGqA
O5EWWFAjqxlSAAuwv22PvU5LNBIO/agyFXVJ2P7KT0noAH/2n0Z5bQr4e86FDx8mD4K1v5vTom1g
yWFTpnaoxxKxm36LAsVVLCHZIEtvfM/tnjWmcRu5cb0hIpzNcPpxERgxB98eS0pAjQz6urxLrcch
S5jd+iWKoVb2AlRIAHAwZJ+6g6QaXfL/zgPHpy6rjv+AQTIOq+L7pn84pRHNYmJhbdtfUh2Hyyr+
cL37aiD/+9hIccd8Yf8nQNPpL3Lgs65tfuQe6Eew3Z81sNRc7dgtn275+H3ib1+Hm6LufeXmovq0
ZzxN8nfovz1yM3IgZ12N+L9uBdRO0H38yuluDH7zktBytKVXwweqaIgJobDN3cAGAG5uy5MAPKIS
x5xPoB5DCs7VoV+8eO+VqnnrJ3RkY2IN5xrTy2Pd6fGiRhyeixTX6eHEUxSUaoVGlbJizn7EqoHz
O5Rz1vDeWXPgBxgtF4ehynOFgQIQ+MjfoQDtl4h5r3u7He2smFHZuJLwMliau6wBQEszOBc50G+i
bV3cINeG5ju1sCvD6gLLY4yRLwbpBstTzQWYNgRtq9FlTQQ8fM2wqeoiXqkpk4xgsAmqDvke5EGB
WlQvHGlQDHQ1djjLOllIQMyoc+N77RJv3d+qRkq1gW0bukaFfLLRP0ddqK56mo1xzS3OFo9VQ2NA
ELy16Fi84XEPJEkYXvEbKSQRa8lqYk33vSpWA+3YFf4H9WIZ+81sPUxsfMniFXi5ZW3lZbWA6GTb
teH9laG5H8hVdqgLDYaDKXPMmq8AO4vQ3EVp44NP7Zv1B9wB16uxm+ZdbwOYrHwa+Ppl5eWarUjF
OgisCoIeVD5d83Q5LlrA6YUhcIrAU/OKeyTiBM+GFrHbuLil6S5pO2/C1vc1/1+mu/Pj+ePj7dcF
ANdYUOF2Jcl16/LBmeQjEt2hrEw8YhWKigujeyj3oMNvfMglYHDh4sUC2aOQefCtaHzrsDXy9rb+
hRkdSwRGihf1r8KIcCq1woi+/zS0zBVzW5ivLotd9OSDtfp0uzN9amAa/qUWbqN9qVA58VCKhHtu
Q0fHGqNEmEjLQENsZ4CWsIJkpkU/dTeYTUr0VpSNNbevId2YWsGv08rHkp5wWpq+G1iIGju62P2b
Uf8M8+HSCfEcqe+6+MEqFu1M1NNiCuuIRFhm/7Nl4TDdMBVF3QxOYeTxRVuFJX5pfIh8ZVSJ6Alw
/bi4KH6zPtFY4PHZs/k1KKxzH/x+C5BrRxZYamV35vGvMJpU2G//GyT1uqC7TtzlsrMLk0zLKEoH
IkRTjuWKJcce4d6SG4GP7q5GGglBrd6Ie/EPWHmzCiVwV187aSNGm49SYE0TUY0wzPlQyi6C5LbS
d49qBvNaau0ZSisfrP3LMb9mZhlfY/nGxRZJW9YuCj8QQ7cnXu22h92lmMapcx55KlJlkwpXM0Oh
CY3JYpj9X1B53FGxPRR38I6PHfkg8YHlT45jKht6QkAUfUnq3fZyRZTkIPonnmPK09D1f530pIKi
vEvGO8Ti5eno6xxT1rSYL76ANNGbZcvnypPCA9INkMr9E3sVtXtu682eaPFLCwxZRhsmHBiEFOQ0
HlquuKN1rXKVcmDGU4xbm4BFi5V86uMYdwvB/MFpb1cxXAnq6LROpPivkEFK9yHGhNL8oLpoWBTT
u/OL+d9x/M5imVtfaASA0yuRnVadstbuPuIryYjAcjGvfUVtHXufi7BIY4UtqEWGlfhkfJBPJPRL
ek1sJyGMAlUi7uVcIL8CTWW0CRehAdbU7acqXDzthhh7xlDtATtw0oIhaY5JSo9y6kqSQENzV9X8
0i7rYKVG07MME0ocYZxESQteaVOGDYzu+lhFvfAzmP4Z4Bk/H0SNUzr9eRvExT7fQao77gVENAeG
pe4d8aaq36kkDylf8EoTwqhhJjW8xeH/2oXobLNiRYL1dq3SA567N2CyVhnnBz/MNlnfqEM9zgRE
ndTkQ7Gr9emxmFt7ZGSruwwzyryxvuNPdUbTtAZxmvUcr/OY+Bi3q4iCxRPTMw83YjYboGEOLQjN
OSGhJImaf7vPalErnma49ucq+D3wEuHKMcS05Hwhj+8jWICCp+QiUz8or8kjY0BWPoXjeICSe5ZR
P/zZ5/sM7dQU3qZEvIqqhAKHyBjJJRXLutMalx0/FfqI/8Fh/DEtMm+t0akVQjQzrD1+isGpkdGc
JNzdzV41AyCR4NiDUf0q6eWfL8efhJSqU1XQ1LTqCgeI5mVZtlkbOAIw7aF7LT2Ff5aMv69HWwFS
a12FqNNjYNFul8mwIsPkt/OHiADQfpWV67PXS9knV8WUKQ8hflpFBbYoLDnj4NCWlKykqxciKBq5
LS4SfpYSLesDSuxlN5gfIDiOmIscS0tlaSagotPrTwaOZZ6pH0Ts5QTiN3SkoOlL3hsUiDFVOurm
GSv0X39kpSs0zTOcrJYziU/JW01E+mjWx9/IThBayj1cJSrVI5Mg88Hvnz5mddW2vs0/Szq4h80Y
BOR0kdkfDBcklvJwmONdZbdMuzJoG3dSWCy7U8MqEpKb9SXPwlo0lr9HB/OQ3GZWyikzk6LyySmi
IUvlG98O77fLnUroX1fB2LEaWyh4aSNYTepi5FDyTIrT6RYmMRSVMrD428lzASbokHYVisnRr3sM
N1z1L9T4GNqS1eAAVI37zyskALkCMqTzJX+XtTd2lOIDAsyuPVFSTU1I5AeYKNZV9vj5pjuc3DVc
nuaiiUSrOMVToghQQ5qlCCM8cvDdcr4rixFzgPEbJelPpF2jb3x/0mARVuO4gIC6Y3Mpv22a4odk
7KaE4Pyij8BPvduU6aWdWxAd8RrWnlgrCy22GWzpwYwyD5q+OFg43yzSfAlFgb2AvOobHubvBraD
p5H66d85rCV/MfSEJYJskQ+8l9HzfwxLM+dXIWDWXRgR5lQgbNhdFqt+x0TSHTcU9XArmjs15RaE
8r3aF/dXK/P+xBd0WzBjh/m7t5Ge9adO7eWSJWNhF4Pn95SrgAiU2ukPVo7z8lekjjGICruiaTG3
RUVzJcJD2JtBCdsda+VKKO1btZ/LQB8vRT+JYJzAJtCCv5Qt37mJY0i1OqlXVZceYWm6mBYdcFxU
Cl3002aFpCLCWosV4kDEeHuaZG+l+g9nncI45vPrE/eqzzCNNAVQ7kWtsYhDDfaop2Cg/UfiX5ce
EeE6JT/UJLmaz1gFful1xuok//WnDQF4fD8gAOanhgQBMbgK7RvNAiVWDenjcnl4qqJadwu3ix8h
z3w7B3WJ+vmce8PsdOszBZBH4DkODgosL/zMVHDKWE8hPWVb9Mq4MKV3LpFjhtqWIit2stNXx2Jn
u1Kzbl50fwv6UCiegEZU8s1Hq2J3h+uCbehRd0xhwDmrm2sN4xwc16N4RMgsD5CWIIsf16P8Ilsh
d0ZvNPANqTJ0d0qJFlmkCzhouys7XQyUXKNZYLbSJO9xvBGyy6FVudcUP14qZmo5sb5cdc3axNDm
NzC8Boe/agVmahe3VTDlTE/uDcXllDP6zJVfUSYEz+4GfUtbg7sKisF1wi3uxvkWzTec+Hlu0qyH
jtU5nIgWtCBkq9RdhMrQ6SuwzINuOFrZSZ/+TnNnHXTHrMokR8a9E6mrugOU3LrdcpuPQeJ8IZ/R
gVaCwS4T8UpVMUhZ0LCfMHJWnXfxeNkEBUU7JWkyW/fKS1G0nLgSnGzjCCtWYTAwOFP4X79vQgWF
pun8djBO1nnPXTzrCwEwRH+YDQXrEXFv3IGsCGSQ9c+0y6RK7gG+4gPogxVexXze4+M0Q3nutnJq
/tAq6FZyr3t/41MpvJS5cJqN935KPoL3vXM61tkbnj3//k9788khMLqyrvL2QBzpLGpkgS6WFeDj
IUiTPqj+J1rmhp7Zs5giWZ0Iy/4rYDpYGpmdZhhunn7boJRd8I448ByA/IBdyYPPNFbze9BXAA6T
wacQ+z7lNW9X4Dx+ulLWd8zo1jV9mzC1UWy86GP2Y2+lI0R9HFtG22iJMuG42yk2KF605Bs1Xpq7
Z6sD659F0DATk9NC3PfWr0BNwL82I43gnYb6WqZLJttrCNGy2VZhfE11CFMbxJzHlmGyM4AMU1A8
4xcNaJw8HA9ptHmDYIXRftThiGkFBeIe70zJWuorrrSC6yzka+Eie93Nc/Wk38kwdbky3Er1bSHz
G6gybOwNC3At6nbxaY9IsB6tJDeN/yvsrs0CUDt/6aSCyLhktxjKoyz3B9WI2LzCJtDPnwd0vqVc
ap3Fd9OD0BdSzbVt8/aLZ6JtGVlDjjhfKpgt9Xlw+LQ+0hj6G08GH4ggJ5fz8Ok7r6NedFQEBdpC
1XsEzU6hEGnx/gZgQ1n82a+kzJaBuGE7CTYe4HhC5hbqEcfDQtCedhUjnOXacjUeS/YjhjI2y2k2
h0nRn/7AhbUltGbEn6BPMbxkCvtgE1T/bqoI/TDF1rQrVBByZctOGKP26KBpUBLoZ/GwNGLs0AMT
htOTPwyuI0wTbQaE9olIv35YhFoTg8ULujGKS7NxjmNVdycUWRFKrvUzSEc16yu0LuFIn3gZAb1l
C9L9mF5+MD9FYhK8XRpXYhuNbLiI+SOhPI+XAJGKyjVVcs5SkDygsfMBcpFRKq7WErNkznWiLFla
CHXB8YHDFc9anSiMrIuIROKyVqBhwhKsvd94PQGvwiFTnjp+Ap+zHUL1k54h99aPWDZZSG7Egn30
6+tk+kSkgJ9owSGPHrGDP4SYTDiAxnd2es97SLgdCtj5tmDB71Bwy4LgzdWmYjvCs+kyFQadWPVg
ghfsHBZIF16adbQPPxlUhJbytCGaxy/C1ukVBoqa7aqVLVHXBOoTGIh42j59t7C9bpAe/ds2R2TK
uWgISx06DkaFNF1ev0dZb6QS234mfQR7ZZK7VW3LhNEsm6Ph6q5eGf34XgP6xy33uKAP0VvWf09Z
WTZrwG8EIjhxW1f4HxzmJm3RBvSdM6wEuOvi1XKfZoSOpxbS5seJLBSXHSVTZ1YJmePise2RPw00
Bu88soCwbgJUAiuYzEBaBvJZ7h9aii7JqjPEpq0IKt0VRK08+ZZMtylCgKF+984kvmqk+gQdWTA8
FmS28fHjnSAUYsAHbpthqk4lVyV8D9uA2zOffdQ+AZSB8xB2M/7WdFbWS3ix5cDqJv2o95S6Dad2
X1stQN0+mlADeE1dO7w7/5BUVnQ3b/2Idv1XFdpW5H5wrfy3kjB87ykS6KZARRkpT7jYWBJi+l6P
/HdAiP/6ZZ9T9bjoYh8nEYD5WKkd0QJx9rKwq8daXiFeymNcSxwlQWREOybFNbMJj2QTgBZ+7Wg/
QgCskgbMQIkiM1RSbHaiiHRKxb5dPjtOobuhzd6fCxTygIZHW6L14NxJmPFItCvMcPKZehe0HK4X
cu/l9WkAQq+V5nAtZPZQlJKByyKn/k/NtpLUxK5k/NEE1j1a26thUFruSs8LYBjQr3p+UatPp48d
utoz5NqeCt/L/5FX99uYzBNMeD3zkZtwi/huKd7Ceh9asdsuZ3Cj/bCHzS530NQTwbpvGtcEqgt6
dbYYxJzhPWX5h5y8YKaUYVtayRjSqPcu26hWGSn/sDzKH5MPcituhyZ7hznAuyngN5fV22Cx6n4Y
qX0yrARsNRXua1TvKBZh/M9wlLnSL0bXVIQWeCn5a1zBeht4O+e7sEfkcwvzmS333Blp1zSM39Rn
HImWH35QcuVa/un+TTLNw2pc2u4tnSY+9P7b57cMN3RdDagnC3LTZXGh1uaDv6u8pJPc1guf17o+
Qe/qH8BsGRdjxEVSD8GD7enl6j6tYLxAhFSqX7YagxO0lz5SRZVqZGD7qtb+69t+sVafgEjtKFVO
mS/T+idVzGA8RHrQlQNMJOwiD/q/p8FYx5i8OSnqiC5z3HyK2zhanL2uVBkbf4LaORDnnx50vt7I
NJV+Ud9RuVPikUzEg0McTA/YuX1RT9qYGz7vmlBsDsFaamX6uYZ4BI038pYDCE9tXaS5UuF2PBmO
a4aTFobZ5JscIKaGjQFFrumcjMdA1JBTW3WCEevxOMtJdeztERxx7vwkfXdK4XLPhdG1ZogkUWec
S6Ws5qsrBYw2y+Dp6DE11UFTbuoz09GVL2MYT6RC/iTIQJ5Jej2ObJXJwjhlkzn40qZiTL1WoF3V
qRDYfaPBAcIopyQvAaNIKcNHa6Ow5fHNHCiIULOaEfKanFqIYfTbg2ilz50rkHZDHcmKTDIXkLNt
1e3NwxuvmDnGUFJtH4jt04pYt5WfxiJM/KuDWcXLnevMLsKYRvoJkEsgbzvH7Ep3HvkSWaeY322h
WZGhAnkWdUI87oTzVlL+u/QeGPpqYGtBC9Tn7u5vlAJaLV+oMKFJkJGQo2jiy8pnwg6uhSxC5rnx
bIXBNo65RZIF/jSQEZyggxw1vVLZHqTxRs3F/bmu8PPbpCUXOiRutWadW7olwrVu8VXVIoNl5R/m
C60jlXq/9vjYVXVzHblae7d7D9Q3+dpchJfBsylpMrjOM42xHYuY7PcwooD+4Qku+mRXQeIUN9CT
ZQRWy4x6jUmdnsiBBNGobDMRqCGPDBhM7csZwZkFkJQgdEVHpe7Sls2JfruHZSxTiOSsWTeZwe/U
GSPKEjYfIi6I/d/SITr5EOpeWi0oGNnAt7hgfFQ+/Iw3wiWtqge4A+YWJTa0T3W9JqKZZPFpckQa
FeaeWvhPt9JNrI9AsaLvu6fcFtTeQwhpWoj1eOUX7o6n/8lJGBETOa/oKd4whapHYt1ngk4mVzwe
xQq7uw82nu7Xf0fjUadObxwPvvzy9I3RnGuQrh22uKN1tIuLN0qKNnjyHqw3YKkz4l9ebvFpP/PK
tTUU5yT6i8xi0qz13LlyVfh9LzmES61mVEK3abbDiLj36rABfJXBzHx+L3y2fFwPw4QfTEjEYOPB
bb3ZFCKoXwbcYy/CKsT2W9jCMBCyxie12ZKaiQXXTEsu6OxSvP6nju86Wq75zFiPlTmykUbAw4zv
Tac5lpsFw2tOO1kN+3Yw46wZobkaU36mxo4UGiMRi1Q4jnS0Xn26xfSgVznELlPdjw04WjvDkfzo
WODgUdnrPRkCk48Pq5TSDexjcW7iIEsDblbkErZvx7VAwPhkVi717FMJbhaFp6f04SKxRchLba8z
O14lkaBgVXkbpam5xMzHv6KoOrybMjI+et0LoQubXMeHt1WNq7///+khnYV5ziwsxiBmE1GDGAeE
wJr038HSGdDuQwsm5+f/uxsqEUvmi7wnKOX6WeLePbX850gPFQGOh5tUPdSNLuXzHldWTcoY4A0k
wdbWMyjbnrreQqgXiTp2BqkD7vpVtGvCR6ceJLTA/qPkcU9wkVT3OD/Wi93965gMJo+FB25a9JKC
lpVt9qLCELez69N26l85RLriuHGBob4lVKwf9TVSteR+jiID1WNO+F4LKp0lLKsYCxOu6dxoV2Ln
plNSyPpnJqE3JDACKjgqCaJv0HwsAymKGQaeDJixOqXEpOvK1/A6H7TwHFB39vHw4raoA9PTc3Cj
Y11p9+kZwrmr4gDBlHYDRbcGt5Nt+VFOcgdlByiSFzZ8s9sm+vhwxg/wtbo6k5NdlsqhfdBSGJtl
RNGz4tu7zgR6tFk1fYA2/0tHHvveBhW1KmX2rWCrq6sPnIzKSVRjEiU62rYbYgaI1FkWnoK7bG1J
RX6y3wQs6W164XSnwhW8lYGEkRLfHd1djYGEvsHRpiddbHo5yU+2lMUaPTH6/HKo9c78c+RrWfdf
/rN8F3TII1SKjOqwRFS/bmoh0KzFqOWSyRj8Po7hefBGPIc1LWf41Ob8j4NBH/DQuXqbFC6EkufG
2a6AcgJkXSsr5rKE5hwnFsPkKXtn0kDi6bRhm4X36X7WA/Tu+SERiZSI5URcLqLuJvxeBQtzirkl
/uU2ydL8fLO1zgVMbdyKpWRtBDxm8Uiio6bxzChCbXdEofI7N9CAanornSkSvvJ3Humvruo7ke8v
6TKOaWVrTSVEiViUdDrV8V7MKq+ZDQWmkFk+j0+wLjWwjbSuD4cqJY8lCZ07b2J66b632POWbY4m
h0TiNOD0uktV6x0iIu6yCDDOlR4emiWJI799FkeIZ9qTEE0bSk9zh0wfAZQDK5HCfoc9JPFNjQ1F
/oMBrFXypRgt+0BFdAm3DqeWzavA3eE4GTLWRnWw3b/7tyyeYbPtbu7rVelAQYbiePxEUxEUYtZZ
KQjgW9RsbA7BSg3XK56mlvz5yyorH521zGmGNO+mhhN6YAHUNNfKyDzqbPIUzJOR+hV0Zf4HGH4y
spRPilnbeY+sBqkx+5o0wxyf5fKK92lmyLLeWvM72AJGQN5PF5TPkvx+8F5HXMY4aVvoGAwmY7MN
DQzbuZJLmC3LCPBwgZwKT2QRm1ReFqn19USV+C4EHEtbSW2z8XIZmJpSiiPI8f4gZCPGLd+72OPM
eTYvvkCXGG42QH+hbWMrQRKYQl/rAz0xDdFtnA9GQ6P5xocEC4MxPBZZCn+p1vOJyHGIypE8jexA
gNHstA0koJO2OqaxgJmxGVgJCHi++ksIrBX8Qn2XVkAkq3Pomjtf58W939xe49Ij5WtFSQ6Bg5ie
eqOo4UviKBlzk7KlZlK+gVKk278Ec5qS7OtlWt8omO5fi13tk1h74t8iKZmWd/5GWthpeiGhl8bg
AAnvWvKPXy5iZ3aDvizbrwJG9y8sTuigcHvcwd2u5FjQjEnrTwofrHUnfagXvINMk3EcDFJCi4Yt
UydBvwRPDk/9SSTJvCQ5Wz/JeilGe7KPby0cyaWvU1SGWYODI9+cZi668Q4sT1j40ABYggloi3SL
lL28MvSlqRm2efjQVCC8R/2gZE43fTCKeUDMLZHjC+bJApDkDOM8UEdQ+kHSNhbBiwVMZtYCGLmv
hmQkX1ynm0vdGLyPZPrLLElV2X0kiaTVof98+RpCOwxHaGmagnsaZJaQz9z4CRpJMpEZ7uJI/EkF
+u+JaxRCHgNyoRhCuQXj+iVhcgsiZHGeI4+xkMUpTy98RKEDB9XSkIbDtpGmexfHuFyE0TfHVeIh
dz4w6fTVvN+YyWZC6EEHu1zSpEmdtL+mci3vJlfKJ8yFyEpOVpxF42i54Ys6Ut2y00Eccek8NXlU
esrrU0uVkG1PloS2FJIpMgBU9YfmxAV+3Yc9ZTQRw3L0YHTpPqj+5xjv3mxbSsn/jUKpc99iFhtt
nEm9MWPMf5v4/d/nJZsfecShNhfQsugN8+NuuUw51kj1j0bR6ONvDELRHH/yVCtpbQcrIhbO5VXy
hT95QkmMHJHzG92d6t86mMknyqvuf0tWbwsV1g8cnbh3m0+qCY+i3Mrl6HNaUs4bVaBt/4U45Wxa
U0Xz2ZLSQF+Ey9SEs+cOUy+9iyyrZIFwWnpnbiMO7L1oZ01yoUP97e2YDcS/Hp8JY9P3+VI4th+Z
JlTyRbz9yWpK6jP7rQqAsbheFKpBweqIwTmDp5otyYNe3vLN7GBOqu7y/Z0YWnMujyIp4T23b0wm
s/YrEo8Qhtt4z3BbKetc2fc0Gqb0I+1jlMWdEAy5mQ7OndhWI+XbZRAzVReaa+1ndHVSXApXdVnm
T7ZCY8mmT6ZT80hRmteddcE6wmVvHblTPFV/G0jjKDRObXJpj1WM5P4ww8b+0hZsCLnamiQAa4F7
DXOOs0dB5oj0C6p+uz60fSXktwP028g7f75SMPcj2/uNYl2ZogzWxGYB00vBEOP/UjcRE9sIkptT
YN7G2EKsVkEsOUNJdCbwFx0fuEJrAU3iMNdu0h3ZMHrtUCr/gE8Rn3cgb4Jtf1W97jmPgcjweaqx
A5NACLcG1zEhCjIiJ4esX0jNfX0iksEnZcSy2HC4K+8mYb9efR0+h4WbWA5k0lA7Aa/hGa7IY7Ch
tl+m2+Dd8WgR7C8xSC04kDGOJoPdUVHZw8PsnK4wibFr5WbjujpEZu9/yk5/yVxRgLpRB5Oi7rPa
smn666RyDn+BdtMF2GXjbGI7704hm9BN6v4XYwKN8Gh5J55KCsvEimlgMtW3b0ZUmpx6Ha7lKkf4
COgKaUGp/oyAN3E6taa5M2ECu06A2yGqdPCVljW+P45/edxKF6Ib9Ce/cQzWaTxE7WQm6VjVPpt9
XhMxV4xDv5pXNsOCStFs8VieCtwubj/F/nRHf+Lzri9v6NtmbFePRIBCTGVeRotUmhtIvO18tPF9
hys4mYfz9/gH2FxCXCjdp5r1rSB8Tnj8LC0W5LCpIkjQkI5fD1KkhbPGk1deEpwEz3CFMzjsuwmJ
E3Ai+SXnS6lZkm1fLWYz2466NVSwZM5KKSFmxFqATC6xvk3efIM0gmJcrUncKQRdphtqb6XPa3eh
ujD4EXEd6mC/XP2H3oEAGWnBEqj3ryFAnYxOVN590vBdKSbfxIPsugnct7pnGAXF8OCIbFqDhWR+
k7DEIH7iAIcAmhDk7BiBt1QXpDNvIkOw+lQ+C1MZDdnqBP51IakJrUFS6k+7jdabM5pfFC6F6DMD
y8hlSznHSFp9Haah6eHhG48jkZR/H8Tvgqwz7nLsfLPsavpCjc2aCLDtLh6cK10/IRuqanhPXzaN
WK/kTmN4vTz7L8q2LsofFw0w+iu3EGnqa/TbJtJBAiveBwiDJfeiGc6Sqlb1/M0lY3g9ywAGwWa+
vbCK+XAjTBpXlW6UYDuFUrefuDfectVQZ+3tgu3Xuqr7Sp/87EB/v2O5ar4XQg9vZLLmfhj2gP+j
KVJQj3rtCeq/1zMyMdeh4NrKp70lWo2hHBddBloMecB+Fibh3GiaF/mVDA9kLnOWnSLvVYs0gqMT
QWXebNXNTVm2dpui4lcRXtfO7lAVDiTI0qItFSRnO+QF9oRyfOtoXzWYHMRHrb/p3ppfYO107kzO
x+j+rTqDznbdtWfKjsFdgGTw6GDQw9D8sVSrohJ7LB70o+J+0G3C86eqK+edxzB7UkfN9J7IIBdw
BRFMLFFv627HK5dkfBApVueGYIjiVikfM4wzch38TvNT8ur+kLHX5zWIgSBSOyMG3bErp2Eo/ciy
VBAvJNwmWmVCc9aat4X2XvPflBFcw0lQHwq40TU5w+XRR0WSE6zISAdFL7DAswmo5sc20H1g2AKS
nPTB01X1PEMe22k+EhXLOuoBLCSnjqMctq2TvUtAblikLRTG4e+ftYo/OxDKYOBA+/22Uptzg7qb
nE8L7hfpu43QvIGi1Klxl+LA1uRtXK8Z8slCh+IL3OV73CvHbuhnwljVYkBGu29TEIwoigrXmigT
ybY1wapE3YItbCaHOVhjyyHJDlcwsI3UmcG6D5RuJWYXcY7yzjY/MWr7wuPIn8azqzcG/049Pqbj
gRuxqRh4SiSTMcS2I4U72jeMGzL+nLjCc7V7aMTEJNNSrAtNNlobt/PVXjIdOoFPmlWwFd1X2xrs
3AygPyKxZDCP23pA0xrwAG/bnZucJwmA0TwwCPtFaC1pJJY74w5leF4R5ENVxgZw+t7CujV6EARF
OQhbNDmClH3es8nt9Z6UEcKAMNU+OrZJU7hL6yaHCdOSbwUBBFXupSxwLT+eVmFRHN8Qe92Y3xeS
VomMyKMjCkxSDqJ1y37xTMsZDinQ98hiOb6pEMU0+I5dIhR9OfLrx/bLlRClIUaUIR04lL7/9631
2OcSgEt5Hg1WNu0xvLAUcmgvjBnZDY356xD+3BbX2c2/xWysreyEnTn5ulSIO8K2tax9fTgcB8pD
fC6WbuF5zLohrra6uVHA4yHyvTsUYDRKAcZKqp3M6CPeKKgiPWGXKSB77/2U97JhGBVuIInlUuOY
1eXLQDDFvKkytnal6VdNy+Vgeg6vD4yw9fUfB8pnf0mNiG2R+0MzwKwc0UvDpop+9+ZipncTeIIr
t6Nsefte6yABJyepTDUN1+OLIGWsHISR1/HNPIVONQwIRvMwGgAxXqEAcbLzgs2QW40izHJKuxLV
tYmbNeShplkJ4Ks9DPGXb0W3ebIC3n98ckaxhHtWgvVjwGLvB5O8J0e8gBkbJVJ2hJpYJBlqWEkC
LbrORArkDvbv/0iBkE0q38FU7+zKY8OalCGy2bix7LVhw9vVPxjDTOTvcQVz/0wt4a7vi3nGf6k+
/C/xfVMtdKOIeN/AJ1N8u7a8w3tb18NGYlTd4qYbUymGjZ4fxujEvP7dAQmUb9k9/7LI3r+xzv20
VH6/YfTFXkpmSGDl7afPJDmsN9LMBm8A2AkUrlCiVgOiq+CrDk8BBuvFEj85Otkl3Q9g2NkHgDex
M32eCx+k8k10dYFbFyTh2ERxzfSGVQbkpsG98j+83dG8QOQv4D2kwVJyO2rMwrR5LaQ5r71I5/rK
/eXJSarQQ279a65WKGY0fM/vtWYXEO6gQ8cvPSSQzDZtAaMREV7R4hL52m+o6KPUwxF+Q3Ml/8is
ZuViZMeCHUc/GI8CCE+s3ySU3kR2kI4/1PyYOXQzDo6QKRBsqWEX6ahzJTRVkGR8EiLT3Fz0K4la
+cdQ9+dWVr2IFQnzSSm953mRmjP2CQ0LR/JCTND4YJbBnH0tAHKu/YrS10cN6dZcGhgLWsjtDeI2
atlBpTmfQtmCPYxQdNM6b2DDbquqCK4lJ9/4CTvEuWfFTRo0ni3NUFdTQKhf+1EoTqV2JIJnC6Ei
L5FFuN9IalZ1iBfy8sBBHQo6SOaQ5CkvPRCCz4z9qwI9G60urMlR5wfoTw10/sHMwEuz2W2IwE0T
ybF4hoCgcHFgTr5VjOoZj+ZP79PkCVsXRJy6usyRJuO97QYFesyAqMSKRmVzJ+OjhJ8svLDgxM9l
gY1STuAxz3Gh8PW9y+YHjboHIC2qKAl9zpF7emk+12hicKCUK5X9BPWQq8efCyb+xhOnlQcWsxJE
lgz3sSxnRDOzfkAka8ZAGC8MoMJwiT4TnBbCAEscSQuwIWG9/+OJ9Nvm/adGYJAhFt4TxTKLt4HZ
WHtKYcX3dpNFYUh+XFQBs/5LVCqL9Eq4LCw4lYNRKU7fCxnQKeso04sHeaKBja+O7bhrkwmJcxMb
q1ZIvmiopR7qnSRNnyu9McybXpQgOYasl94GuGoBg9QNE2fcty56PW0qmH2G6o/y3kOO38+Ixszf
4ye1IXjZiKjmoTmcWl+FXncyS9KON/vuVKzFsX4eFCLowduRTUn8ySsM5/BLJNsXLrtFzS7LpXEv
u6TotLjR0oEMT8Ar9scLEqjjJoS/pGhr5GI53TiKvRmJpZHP7GoTpiJWUGIvR6/1CiTdO3cvvedR
lmPULn8Inw8YIUWW5kvUmvVVdtq6KI8lKXrtA2uEBAZFjsD5gz+Ol9r43vUQ+HL2w9xqfB3V9pLA
/lfo+OmKuD/hY0L+KorMyg02bq3IBJPynEfDIddliVltPDbIisDC+JAP3oXQm+i26vWi35/XKKxp
xQJOrLQjDatzMNh6TzF+h5ezVMYCAli4SBSoV7b59zdYrSsNPTqXzswagJxwb8Neb2rExysoUvUO
zvnzldmTOLf+f+sRQ4UIyVpF2iVwiuGSJaKw7/MGeLlxgRTlKu+RQTyVGibLARIQEltLTSlANc2U
0GqBXpXoJ83bU3/VCFpG1G9oIsHA19lz9u0geRpdWyRm6mfddgB0VmQFlel96BD9/HbB1cFmhHdb
NFJFTmnyoaX4yXbG6yUs2KHlYO0IbqiFsftyBR2Cp/hhhdzvAk3JBim4Io9GME/PX4Ji1j/gC9h2
8j1iEXiooJus6BUyRbnyECs4UL9tJPDm7JkrUxBY5hXVfYylqwAB6EHLbzp8D/GwD3K8i3k+tKa7
+LylqI+42OlO6dofrC1dzNUggdY8YMIb0Kv0hyuj82ycqMkeonKv36OA8JxIcX0ozpETpuq10KMR
V9NxLNdesrqSkrpZ9WC/BG96h0Bq6ZoVKSIXthTPAWMwR2O5J/1kkLskXRLPTu8LcTZYi3qzzGJL
TIobEnmH2CHtvMikTxnZSoR+2Ahl84E+QuhL2xeFcz0H77NiyWfdCQJBpjz1cD5h8tTKc80LDluJ
YQcv8gUULyS+OwCAG5LDQderMrpuEcOkF5brhdcfHEvbMgFKEQXeyBLkUYQ90aOuCurGe3cdvPy7
ilrFfLcWUXBEM02uNlCtY4h0n6hf9zrw3c524yQ8sxiGUwSy4c7BACotLp17PSWHfEtppiB6EBN8
R7fOoZQ+KsanLcBXBaB3IZIvajeLq0c01NKZR32e1VthnAxFzAEyBMloaZedk6qM0CNCMiQouLb7
JEWg/HWvwR8Xx/tOnye9xCutkafj3hW+xuJe2g6uX6wPFo3APSiG29HsDcBz1TtgEthg/ScJpU+J
ed5Hu3Ml/8r7R1VRclu/28IgQIzWntGZFMNXu4L4dciNc6TjD8nzj+cX275PH+WqM9V6f5a7v0IE
wfeoyLM8exIavYV7WvfiHYVnNvEEsQ/CwsuQCnS/va+uqKSwZ+R3ylSnMdG/8LoRt0p6DXidBKaw
JHUPivhvQNg+lpyZ9mhPX3rTtH7NPC9Wumpl0l8I3JX+A1EBHxe93hChQw0jXkBfaXYjwHTgePx5
5h2QOUHiiMJYvwX/jeCwgi7WPHWZgo3S0qw5m7c/KogzSVDCQgFa0u1lT93hcdB6l6RVDVBuXbxK
meR27uEG+ZxiY6zRGlfLqEzuvE9458vWQQ9SQergZ1+UFQvoBAzpq4o7X5E1wmPHMvrPV9rv3Xgg
RvCWByhhuCKe6kQQcD4ZH+UGhYdoQjr4Z4qHcs99BLQs44A+PIbIMSGcnKTXbutXVvXD7pzFXur3
DWASnlfbTnjrdYQqevz9bCkskOqHe9tVR7pyHb4RFO41Gw0imRQKzKs2DwUOToAk1oAtpOWc0iUr
lCRn5dkVNj+aR6UTy4vUCOQqbXADRwmdjiMtJ5eqbGsWt9duQ/muqKCJPORQNBbKDBBdXofwh3EJ
fze5wnolYZJI7+THa5lp6/pKIZzdUrfLZac5wufU4nx/Jcmd8OJdnRoOBCyg0o9fIxqUxwaAMa6K
4OEk2/PHgAjeBRPNU5g/Fte4G46bp9KniPhq6AZWkLqGz4jRdrYJPGHZCKqTWTuIWlVjs8WiyAWx
fw1B5EfAHwZ5KRcZm2Jj0BmeRKRg69CNhWKO4X2PP/Dg062T26fYmVJBhDLQS6NGmDCwjRlg0dSm
A+0aHgm/GoKYnCvWpj01ZUTn+54h106B+bCE5V957peuZZ6NaWDCanu+7X5R1rf5FoX6h9utcYdz
PFy1c4Ly4Q6Yg5DmlT+6v4DXZXsh5ugPYl0VDTymM6DGtaBnw/bbnDckBZcBYpjzY00zcRH3XzTd
RNEQNpxfeo6wLVta5cO7CO9O4eqOhsNSYtIz1FyI336OnutctXWxFBH1k0UjUI7VNyQgIAmAtuNt
0ITkAm6h7zknTujlm+eOk3Q7VP+EEar7yfsjA8I/3/Jd5q7EMDT3SHzi2P2dbYPTLZFxF5Rp2dyN
mwkTkbgzrsIvszDHFRV15+ih+B2rSP9GZyRuIWoqDMkq/4vDUu4JRWHUEMWW9zdwqWxU3lwVE9mK
1/NEpCRXRSU5Vsx2MKyxT2oTPPKluBm8jOhUf+qkpSHOvoHoMb+lRLiutOy9UiNtl0O49S9sWwgj
rhDp/7rIqp3qyS+ztlK2HPTQ5O8iAEjWEL8iEDxcic4OLVVESdZuO1LhBgxGf834pkOIWNpXgMaQ
8XcBcDOQP2wYdX5ubfDeD6AedzDjRzTKI0JtNcbP0eNd60RoPpSsIk1Lcs5onK6XDdnYXRPkXzFf
tDIe6+xvk9QAIfIfCz9tQnws5u2Ueoz1LSA6oIfiTBsFKNXDcvLRyMCGrGW7VsSbiNcqfiHA0tP1
QXnYEfgKpQPYGIg4wnzgf7fHroYj32NUpqIMMjkkePBMGF61LIlOeejQ3Si9ZLV0PRH03rj+CNAL
jujf+DTBI7ZucWgKxAIlFZ5kwP/i9ZjvUGtlRS5G2uR/p/CRQb+DtIHUvI84RFvhm2tkg0Y5fl7B
r+aSTOzdfh4KHQBC6z64ZkOJ+2Wsmjkac6gfCgG6Xg6OMCGAxHJeoUtRN6MZSOnQboNwaoZtI/ja
/tPCkZqa0RK/YHVK9864Weh2tE6WyC9Jq/wxbufAm/u9pwYnS6ooYWkGJfQvHXDvbhDP41ne06KD
rZCUgh/hfjT+Hdr/H81QZtsWBv8cblKE2zcsK0m0OkxttUggKIRBUyNKT+DHSi4Xk8bX50d6YgsV
GsWziUs6ow4cJER9WmrfM+l0qmfrpyl5TlMN95FWRvx+z/korx2/YKPxRfBNqWTSyz5FNQQE/qRi
wedQOG7qEEfLw46nADnQnGPkaOM3jOdoO2KrS1wSG9/5veSk4f+vVQRkcdpBgqpvo9KdgjOItNms
Qg6N4o/sFT9Vd7hrtvYpRx7K8yd5bRTSxCiKGCK/6QGFRvM5f3xX+/Dbny8MwKBT2pwidvnOf3xP
xr0V/e5NTp8K6+Pa6dW02GtEJMT3MvzM5nHIqUe3ye/BXLd9KjyNOJBlf69XaExzfYZr805rpR5F
19mHRx2UjiVgM2Yh5YSYT8o61Vh7XeF5nr3LHjoGjmPEXFRGJ6H33TQ9lzdeMg7TPAqKYCkAVTY1
MEhQzKRhKqgbXBxY97nTIKlkEiqT3k58uFUcGGhsBELTJbCoqDIrsVQMWZKqOmpZ6//1MyTnKeYC
Vqip7+C9lawDzY+LQkCjJ2fUjJPfPNWjt+opy+YxBI0D34xVTl+DlLPB36CS9AcKyAnGaEWNLB54
N2NFE31p9j8NSrnWOPXOSuqSn9/qi4ovSU7d9jlC9YFsEw+ZUm7SCusu9lvDO9Kb3pXqYOubxodI
1UTmet+2SfkVml5ktuibOeW0FYrbOwfV7A3g/7zR4SjXnnL8aVTHB7axW+8Yh5NGCEVsIq9YQm4j
yJBzAy1OCDSwsCn/OJaUTbLdaxcYPVhN42q51oqNHWPZ+kFIOesckUbrf9SRgg/CXBNzoz1tanWl
4g1nRwPL2SB52lYbBBvl+Rkzs0NirYfSmaCyhg8JSey3JYqIgKOfXrU56jsaAEzATKXZ+WL2zMDD
gp2M5INesXY0i+vvMpS4bd4tgImQ7QYUg2CKh7DutB4xBQpFeTUqmmRPlEiIvZwPV/r0Wq7Se9eT
uJfnd5KSZUwh5Dy2pXQKjM3nh89vvO30xw94t4aliZL1RXFDrcLUvSQUwMMLgxfCZuVcLgloHyEN
JZgXqgYyC2fHtMB/3XyORTIYCpJRk44OBC85IVwE0/tyfxoqcdMDHghPyvgwws/w/ZHLgKGiVJYy
rwL0m57CT2CsPW/a7zxxUMI88IeyTnWlqtXEJPry+/ATqXqOWrZv3+hN082gnAH2BlpZLqM43p/B
CB26swYq+vvYg8rurwcfC6niTeESuGZi7IyVIiF+6nOiMQRlpj/jhoJyio2Y2Vscx8S5qUOURI35
XOjCsj7lFygPp2HnVJNtP9xEIS6vWnDgANHY2sHn6P7CqlyA0ZojfOnfUZTJ8KXDuPEYBJ3MdrTs
Mdd/nSGn2WfkN+oCt4NkvaddEErQWeuJGPv+clAz6YmsgkBDequK3Ds60cS0zlHPPPjc4leTiD+N
zk0FbBOmey6Ad4AoEc5tvu0LlXXX838V5v5Uso3B+g8EkDC+NfTr/w0v5pagOzZGLfXVXM4UvVhd
W4Pvei75gWmhDuctEZVUCgWrtxYtr/MprLVSgqIwhJAQrTneRUHkndkhZ6/VyhnBh0zAxFalMLXx
PHuhm4oUo9rxi5dfDfxvA/osmjNB7jfcEUlQcd+lMl8ZwLCgo+mcvDZ1AbKo7U0Vc+J8J+71i97H
W/6a52HqyDig1mQ+nVsSyFEppNnn99295L6F0r03RMLqJ0rLWy0JaFOuSsEotbIPsvnCSuwmZaPz
pvNMq6bknKBdOvd85Z/Xag337vIaDSlplqo168qZ3ECh2f3FKSzzLcwMyuho+pZGVpzilvKqahcX
tbFeVkHI8ffs5KVqKWHwQGGIQNrfd7Nvxf7Jvw+SNYVRTT0wdArCZ4ORV5hCHi3KFZu2yjCLhuLk
cn9aFjl+av6CIZg7jX3rfv7P2YW02n6zeYcUQu3m3Hw5ocwXb/yQSWPJjZu7lVmH46jTh8MQrQt9
cJH1N3V4eb7Rju3g2LKhCNX7Cl+coC37PvveH1ag8mnd91WornJpgvgL75qOhuQiUn7ID3qa4ofg
H8hmZ9T3moE7OJij9Y7+fkcdlMBd9mr1sOMihetCIHzzYFDeQUd5OI0QjfgGeKVIwn+cZPOK5KlK
a8usXOmRcVlLY8duc3FXcq/jg+XoVun9dwwnSwAnZ6ClHxEuxlatj7yCzNLcpMn/mEVGEXb0ci/H
gUyzmv0zw8DZFNN1vyv5E3hKVh9PPwBkzjQRqXu2aBGE36QVq9KmCkfZv5nkv/XfNHZjfiYLij9q
aY91SJZDniRwsSfq0iEIkKmg0jEdIpfaPsaZT/ScG1bLdmCXjENmi9zpe+J7bE5ta6/awfUODU9k
QnoVT+GqjucakRog843WxxQhnCOBTvziDLA7d2uCZJnOD6sox/h+Kn+mTWpItdJC2VUyxfFyIVsE
9sbi8OlFvZVmIPFevWLTYI03f1VcdsJr8Zzf5IvVDC9woWgEUpmpVZHNX2dQu0iM7k29cOhgaU33
V41830ic7fnX+bcpKUmI6ZrqAxQu70ZXsV4P0rfOQk1q2vJ4PRWqmX9lANmmRXfoAARZdSkcW2fO
1+RVpk3FX9JX92MZgIQSSG4jFtHYjs6kaNmIb1QYxhDf+QyUswFHjGVVE4oRkRSrK4UI1KOL4s5l
aehcJ+T5WUh4SN3cEBLBwh6yj10xmoq/ioUgWKMCaGoXlkmMbRnqUhFpC+ZV1rQFESZGcj4tE7um
7Ki9KNpxPAvVxF5xgnG6TawuVkh0aXOlHVDC4uxEHp4TCmGh/Iv6yVhqN5gp59jbK2tmEMtraNmw
bMa4Cq+HG5DaC3ttAs84s60K3j/A3v9Kr8oaSjXDMruyOBzWjVhFnj92EAMYaKJ2VjxPPTRxiL3F
d9jhaVBUz+nCUIeaZTPCXXQihlrqmk1DfCgbW2bDlJBbwy6jO1tsKkaO4/V9FENnb756xJ8HZJme
wr9vEB1OjFrggVEzRLLt6OZR4uZMn1dHmIEdO45ss8gW+x4IAWkpyhhVWtJ/KeDJN9FOZvAfwkKC
XZBBM3ub2lbjrFAE8rcCSdUZOOivn/TIeiyflIjjiaJ3XE0vKf/vn7zZRDasB7NuJblokX/d+uN2
r7CbzawS10dad8A8ORg5XLBiv1RlsC5Lw9D3dHh0bfHP6bSLXaNyw2pWht1u9rAIs2RP8n5DasIp
6D5HyVZk7bVuH05UV1OBvWvQFlCxqNERfw88dDn/EyjSO+mieo2sgUxeV+ztqSKqGwfO+ZyL4+OV
YyDCeyn6Bc9VHAcCI0Uxy5d1zLhVGXHAxtPFt1IgOofWx4GLeHnWH9xacu8e8joyUfP4ctcRcW6K
1Sj6YTySRgOicVM0S7bK8KorE4VRInFueOeEXXmTUBOMWmvgxyVzI5RmkMrqbLJPz8cXFrVtja2i
TKIEchzwKOJtVAlELTaBhgXM1sF6rFt5mfqMrGAU/gfIJUTprlVdW71P9/RTBiwrOwMLSOYq5K2S
e/P2r1nEwNX5h5Af3m/ZE1k3a/IA9EMT9tbk6sfMhzzcQ0FNdZoqPwF8VJtyWbiVFWnoXwsNLpja
ifROlMqBlwqW+h0nlXzy5+DExEGjrj6Ry/9WVBtEpaFqmp0PkjtRlOcoDQbrc8xP1CxVtqyt4KtC
F0tHmmNLndSgKoX3WR7+B1waiDsFDVUjM51vKb3BoNtaNc3pvt23LdEFAvsvKntT6lAA31Yn1E+S
78J1H1At77mL0yY+Yye9q1BvuyMcPE1D8X4TkKSVd6166szjxgFgTewWbDDSHQrYzBJvQP39asSF
KfFuV7iedcrj3+9Pm0LdsvNPb992x3zCs0iydawx3NBOOELSrFp4oSKxgIUR78pLheJhjBbH1XLs
kJYgxUydun7cuY/oukIZrTLCVOI3rodVRcC2wKZy9aPgXwNKf76YWdpEip46D+XJMQD8OcAvM0jO
iQxmz8TERlCx5/FtOWhnYo4dyn60jXpsjNb688Y/RXlXTjDUJVMkb3k1NVER1O5HTvQUz9tihucB
2il3HawjZXi3GhaxZ8B/PlQGC96OPFzXYZgCaLawzXaMlvS2M5snVsW6oJWKZD1CGrQCrV857gq6
5dyUPJfXHoOP0LF99Iwyd6IwqHkgFuNKv3UA0gnP0CFF+qjQrTGQp6EBGQ6qLqh/YC/x7idM6s5K
/B6ml8fmHFSNelW1DQmYqF7fZy6DhN4yb5ALRVnfdvr6gullivolP1XiU0UPTg3Rhc9jbp+CWdlj
2aJDAUCXi+veTdKmbnMCO1+lzXZ5sYZ8KpYuxt76tOJWRJtOE41Wi72U+Rg4WWdSQBmVGQJgRl3s
ShNIQHI0bCLs+p6NfGdBwcbh3h8AwMqpF+B/LFbpczppWtI8jdB9c4cgcwBeHV4RwnhSm4ZjfWpz
xuEp4v8H6IBlRbDK2tPqngkzNN4mk6xNMdVLtoE5av0yIHtKW+gzGJ94ebn3nxvoeAIWZvMROV2d
EKy+Lg+minBh6b4mE9w9bIEQp5JkZbsuO3CvaNZV63/87Qg79qMtSf+Y8MI+s4IWtKMkyj9/gQBk
bEOgIRbBiAhmqnZufzcnpFwgK1Q6bAYBzGsV3JEDiwyYiQmVbbuY6Bb7gT7IF7ohTp5q988AsUkP
H+B1hd96P5fAF1DHoRNd4jMlUuB4TkwBGDN1KinOrkvyzw6VLqPm29Ef/J16dSB2UjXVxoViK5s4
hjIjCLLaIcC0tfq5FCAvHIWpzqjR0FVLMambmpzdMM5+79ri4rPHVVnBZ/SpK2VseJ9bQ1FpxQ6B
DgPEYN1KRTGhfyfOFtoPbmlNWwoBAnW6+DN5/jHkLdAF0sqIGz7a8P+MmbW9pVMKfzT9zz02yp9V
ZXMCg42fj445R91oA0U2KVCcG0WmFNh5+KjsScfTcCbHh2dscg1xIN0khTxy4kXldcSpJSeqtO4k
TMUOk6OjDm7Ohg4AH7uUsozw6wP3lCMyJjmIs3iEWmp771j7zCEUPE0jaM+LQ/c4PJdxWbKLNjk4
RUYONRBdV0lkFlHYCsZE59M0HF4by5uMqrEiauR1+TpucB6xpX9uJ3d8RhDgXgMPysVgoByprBTU
w593l84QKf65OVyNemsZffRqU8Sgs1mW7rNK+7Jj3KOzljRnaSNYvkuVxtYL+zV9uMpcs46YLTqh
E8emPIjAcqqGOOtQWlvnLt63hVXNS/ANGoKUwhmJrRn+kCCrgO2u+KLG4vJkJS/yqfzqMkAl23Jr
qTtgPp8D/ZlpZgJyTVlVYSWOj3i2nqVKpmY47wjjpaz2CXtgxW21ruexnTMpM0Q4Ix9PG58vJLuw
bVa7F/Q0Tcah6PhUQsuPMLyRcokZPDZ4ptXZb1SbYuox8lyLEAKBDrUTfC1LVjo9sZSvAtQFXcvZ
LGxP+9wrXg+FOKRJL72V2zzxurs7NqsiS6eE7CT5wp59Yj0rEUQ9Uv6pe8U6n+PFt80qjEhv8pZE
lJ/K3bnLOfwDmPqknJvp8hDyD15pO5lQR5LqakH8D6o/VHNI68hhJPMO4NURO0spfqinKUvIKHOc
1VkYY2hpuAK3nbfPMIS3KJaEv0IEZ9nmdoja2PBwCsPguyNmlCcHF80x3vrNUgqW25EomcRxn3vp
qPMmLL6sU2VfbkDUjIpOkgfOyMLm/74RWBgcLZfmYhEOUJAssdYV4x9Ffsyh5xRC8S7bbgpbsoMg
/iCiig6bH517smjprIaLApfVuPAJR3sH5r5Zm5CDFSvpOzn2OGysmiRhfb2WcxXIWAZ0MXwd3ZFc
cP6+4qXpbPiab16YRY9gzugvzy47cpaemRnE4U9brUJeF5fUk/bAk1DjpUevxh3yCBsCzIkJDR1X
ax6S5mY1SgB5GBe1Gv3m65pg87ZLHY1tLy3W27G9LmYc5/+1WKZmIJ0WS63/zy77rqOw/e/dCOPc
iVIjcGikDmRvHkAuhzAhYvrN3Yfdca9p6CYYVqQmTqRbt+UpI7ziMBe2sD7KbkqElrgVV5j6LiUi
SVSy8QiGqffmlY/XF4JEMwsvvhYWvdbvMaRf6DS5khmrMg4054Xm+jMsyAi8m9yQ7Vn1jvs4LzZV
LmrLUl7A4sTxFm0/9syt4i2spAFLpl+DuktsrP8OeGbGrYeduHYkEs+w2I+Y8LBipPAZQGWyFR93
V63lM9sZ/nTfGQMSD+5jk7pV1oQCNMHCojDt1XlDqcfD3toTjPh2Dqw5Fuu6GH69Cm+fZbTzaQ4c
y1YhIdIlCKbBoLeyzhJ4Sh0VpjMFhPnn55eagEQAKrnMoXriuLieSfEKi5BgvuFqWi/BpA4665O1
ToYbLdYiZDqqbhKAz7KRFi8Rw31F9cdBcbc1I3m7yFJlezSYOc78DFO7kOdK10NNuQpmhFmNV+Py
/TgANX7g/AwgQRG0I6g4fJF8GdX5V2tgfMBKg4+nG/2wo58RqzZjcgxVDMFb30Ihw+2v2PBD7UjJ
N+HSSv8qgNF6U2kbvPPRP97I0VGSXPJeXTUNLQrr4UcCrFrJ3xHcvjrp4VBqyfOgOjfwz8GBeEIV
QNwmmcev1Xbkejj5YwBJpyvgRzfPgiKhlDujBBvNVxankYASMI/gfmTHV3hyemuUuKq4UovIewC5
tggb1ScoLrFSE5Q+C+k/27yght8nkSn/kldAcVi6iL1BgZwLp/sbKYHbPHzE6ChlUTWKJumnLor5
Snn93VNXvNmidZipvFDzjJ/sua5x1ervXm/OMkLdgV9LXCekRnnEp7p0ObJkuEc68ibNrtWkxMCz
U+E35nmsDupseC30Va3MZq+OSB2yzGIlwq8CPdJz8tmi9JD/JRiOVHxS4kCQ9bWRONBRIp1xRnW2
CUQZLXeWUpxadvCAk5uN5mD3WtVPn0q8kfOMoLULBeqwKu6/gocr6mJRzAPb++6lNxNXuRLDI8Az
GHgAW40NRNVsmWi0BqZkmPMukcZgSG/zE+QmUpD+nVYXKhwCrvjLfMErx1e44aGAMhSt3ufzArma
jUxpKwRzJlG1Btnaco9mjtp0UvnwCN9A6+5y8F6FfnLmK8Yynf19A8x1vVepyiBaUaAy6AMmbW4C
dyKoh+hDFLml/xCT1/yOD5Yd1FZXRsEIYBrjnldQ9WyzWkWkc7i56eFEiabZsUOitqi2++ZCNeRR
qeMpAWmurvsnvocKjZ2ZHlPODjDHPgY4CgFDb2LkWaw/7XFtZ+4E7Qxz3erhf+/s+zdi0rwVBD3f
erDOR20+qXEJkwuMLpMWbkwHbs7WO9CdP80GRBM83tPve/eIX2K7obZO2bRzWqJmlJPMPRCJRnkR
9Zn8emFBjGn95UfcY6lGmQdCxSg9urT948d2+VulGQmuOdlE/K+8+d4TNra54R2oYtCH37i8uHO+
SCt66BvzfZzs2eLfqqA0G7Q+H+Xd2hwtxTRh1lo8C+YPjnIgqLZThxyRop/Qc+Y1h8HZLaBSEvOZ
BUj9MO95YoK9+Chrm3Ho/qtwPV3lOc39WbGVTSVpoEqxtZHGj62+Op3BMLI/+rae7phaq9kunSLL
xRRmLRG+hLeFtJzU1ScOPjC1eJriY/ijqhJKHDU+e+OZ1SjCPMZLcNbDBXLjqoovFQYoxuXT0lOb
C7h4ilbuDM3Cx64WeFRWHyTgybb8djp3bD6kF2hhI0LfQxF/VQQHHI/E/VvxXVUijfc6lM9x+cW5
DLa66z1suoelf5RWuKz/Gqg8LjJn5IoyGy8mHAbRNfYcgpesQQ0Xs5vx3ek2EfljQvqXrLrWA7BQ
jVa7ZBTb4Xl/wa/h6dibI15EgOdF1o6OTRhaY8yukX77w2JabGGYAYLL7t2tw0IikmKCoR7NnZ27
qxGPRQQ2jl8eNQT1FhuK0rxu8FB+LHzOOThQRwEpGseL7gItx2toJZWr6oDLDN16AdMgMVZuXcqA
0V8jZxWJtwqZ+qhK9JIaF7YzNAwSmMRfBuuuwADnLFxWbM4HtSz+XQk4p8Bo61zeiDjqNRv8zx47
XNG3ufbdI/HnvlwekLKGQXpjvPZpDIFoowllNIzKo6pIi8mIR+XV5SRibQAyin5w3lM/tvkEUhsl
3UsFIiuq8luLpLpbygna7KjHiY157j1yiu5cn3wRWJ0DxbytOlAcuHQJ2bBznBzONbQNBBKN4Go5
2soFLxLZ49iuIV36G09pK63c6VKyfzZhjlbZO6+0aPynOvTC+iCTMiA3H63MLMvlQ2ZCTGpBBFHt
efK+lygptbPTXUG0yBU7kpw5XBfP2T1prDClxndNN0jSParv/6iavVpTcns85hI/i2sqL0g+Dd5P
IKn02ISMylKEgHQGyyXlDhfsWuyTFZn5xRkQmhmr7gqxcSR0vgN4JHoMz0qJW8jUvWFiKm62cnnu
tOBthenZTqMuA0LJtY6KXOMY/N8JGlKypLIztyLqka77z383STnV0XuEeOcFIVKOgsExNK2M+hWc
Px6Oy8WPeTp2hQyLIKGPq/slX4O+jJG05nfqmG9whjBPu0cC/LIeaYpKYuwfMaLS4yyci0NiV7Ex
2xXZeYxrIoUH8nGbzbU/rp5xxr1/Ez14maqUts4sOeMU57kMOHEH6JoRulIWrK8Juw5ShTMDF+KY
n6NsmWD6ETiNR7SVtTGB6HlC+MqCQdNFog59MLfN2+lVYFlXm70VzSoaNj7K7d5hMHeAOVdQz/o+
828BKV4si9ao5LwiTcYYrjsGzCHqqyFBp723d0Ro99N9hDTdea/lYBYP2fRqLsAL/BXPrTot6nb5
uIzrzanSWEUGBAmB4qosvQx0OdY4D7RJTRn4RsoicGO4Eb6bzJ0AMlVuHrks04Kki1RoAytbLB0D
wa+V1VE7G5/+IsWC78BuDulqnGGbdscj425AdQ6iSQzbgK5PaUfzTx5RhQkCdmZt8MBKqaT9BFNV
+clzRW4VVojrppIEVLHNLeu1jilAqXuniXM5koKgSxNEaMRKBeM7O1aPpgEhpikcuGo44Ew+2Knr
360abmzhYHgF3vU0eCj3NQ7IFsNGw/TXMqz9DDWPh1KEpIbmG36+yV7PdQxC/cvD5iETKAXn5YLB
TWxMS8yMCPP9kc+nJANSzC8yLhkEQdp6x2jL/UzNIM3nhvwl+aJYJX1F0HJ9mPImNI1sDAkOB8lr
y8iUskHosCaBEAjLlzM5SCUhA3naAFCNwKarpG6GasoKvL6c8tefd5NLq+QyctfXeS8W7As4SCRK
HfDBSLKs+SSN4DdGj/TG/iocCCvnRtY9kbR4ar2tRv2BU9w7SM6UJcZ8jyTwKJuIcV+cn50bKSUT
UOfg32KvP9F8u57bPstjvJulKBOrr7OXH2o4+D80V6SGAypMBHkSel1nTT1FaTysiUvKjZBUFb1K
7zKUDVW5obOCnxDEPBJmIg/V2PpWzgO0Bt/zn+0gtss0oFR87a1hC1MRoFiM6BXjxPLM4OWLr5DL
EmVjLND63vi3mGQmbImwbT8WRMS9Qt1Ve2+Fe6nZp1NTUPoM/m3Bn0hf+Ih8ItcZH0wtg+TE28xX
tgMHtXCp3XCexSSb1p91RbF1sVq3zYCV6aJIhhZbxLga/ynAa2fwXa4ENPDMie61LqMVhubR4Zes
WnZBms7Yy/ZljQ0t0MilVW6VrmTI/9WBIARxFSURLY+5VAbsOhgDgNLOQEyt87wOH2qL2Uiw5dmg
tEQ31PbQbuZNxhqnsRfGiaw5iksENeQiuSBBQjLB42HeAINoroICRKkMT1AHF9GFVo3uz9Ep2bG9
/0A9YCN8qr+p47jrWLd3LYx365cFScfDBmCEP+9qkO5J6rvlKdeeCRt2aDc/M06RcB+Smk0lHtmU
X3uXPiBlxoMiYd3O/MREQkBVN2duvSPZC7dTbm2dWCRYxZw/qFTvhdb1e3IKaUgFCnT6Pxv7yh9B
ReCHUTe5ygw3msCMfoe3ln/C48EzDsHmSBM//psps8X1N5zbEZf2oAXIemKXUcEJoDQ15kVancPl
kzv/OKE/P38F59yx+PG7SQqqpPvzP7aQ/0yLTQ9VU0lE+BZ8zx04FyrEE9h8jqjuv8THKynvHxLY
taJKyhCsYc5qB5UuyQTYgneV/7vJj43gPTjJXEIeqNzZNxDPmBXwaCmQhOlN/op/jySuu2Jpb63y
JLywMPD5q4UNBtMAzjSdYmYeYFgkaF++a26cqdoda/5E2ON480yk58LKpHaZi0ndJ94hq/O6jPOC
CfC82vDqs+35bhmGBCdk6pdDCG/oMWR+XZsCE2q1vmmIzZAEgu64KNHSrKccLst2YfU1V/YGghO2
j58dbF1RnY+WUP/RZ8aSsy/vF3CPWRXQIZ5L/ZbnQzzZCSNoz71r8amtTxYjzkQP7MPqeJ11fO2a
w0jyB8E/oCbMLEPUAtpY0SimW6QOW6P4o9jF5T9xp1YMZOgPb7BjV7InsfWIOtApsZp/8rrVSblu
2Krl8KEm2YU2DVTku4g8m4n3Zz6dBfFRkGZctAbKa28BgSuaI1s7A4XyF48rXAOXRFUZl+06Sg4o
PBrNvMJo+ZRHEL7IXJ6/DrwRnfP+0E0MrUK/rGYQd8IvrqdWMsAdfp2UYzV9sJYJDU9HpprVB78x
gZ/hWxNHge/Olg1y9PiXZrRdxsvkHtuXY/MJkCTG/daDXKuEQnf/Me7FHcL/qVUHASB/c9pceY0R
cp36re7qB1UE5qiW+bH5JIBiTejmJUQBqChkcsbmUnXzrRFPn25LCfgvWVnH8+FFVipAPG7wjIuE
6DBSc/Fh77Y7s6rfLioZUoTBK3/tC5QVLF7OCm+IrG9tOaZPQRyLqfVTUuj8SOn3YUBQ3O/lyvcX
7+Scb+aUylemGCQBGbHT4XuCA6x/ZSPQ2Xd82en07Il/TvZka0QWpa1VFzUhOvTTq/cr5Iy98bRC
1opSMwFLBeu7Vsu96KQuAiH8rVr7Fsisyc9uRk3pjj1MA45ipLLdkH+NyDmWygOmVEoz3Chn6DKf
LZK0DUklPFef8HU/vIliJnLoYtAfP7X+TwEBrL48RDWHxVcSQAY0/3WbgZ7vVRqw9kvihPHnguCi
3s7XKvet0Y1ktkUNFZHwvDGZTqXPkypxSuIdBaB3aBvkNb1tOVqOG9lX8cYjxibtojhqcCDy9ZaJ
e2ZKnwRhu0NJ6MmC3JHzmwLWaZAbdxQLmKs7TFOf+0Qgj2VVwEmVmOTGP8EyxXY7EAcHcFJq1Y4/
7p5i3NfSUxU//byGmCYVViueoGAQETPrvhqSDHw9X+JdZ4Dp/Z2K2balvheEwwQUCEyI2Wvk24x7
djrgi6rHdpvbRUEwHLRKsGf7RSaHHg/Cq8t0iPki8m4EIbxKJAew8GuZn9HFG84/nTDeoZI3uhpU
ph0yf4mFEpfWjJfu2A/jIh1zOHSKER9uH4NFYpGuUY0O22LBHGxLHwHqQruHWRfSguPMclpMxDlK
aSk5GXpT9KITKOQ7Rf1oSY4DYyKS1uB312NBxoLuafve0O/4txz/SVZ6mn8U7SurjymA4EA1LIER
fow5y/7ahqZp/hP620DJFLj9lj8CZq6WQZkrXZYxTe30460KWz1shYiN+uuVXOzPc0zK8fN1El+u
r+Hfs3jcRz92WI6a1NdsP0xR+7jyjKzd7VdT1DjScgP9FHl3vF508KYV6WnDK2qbET/7oD0CKSkQ
dW1Iz2izogXzfh6/Fk5W4d7qO+Veu6ppA+otp5w9nhcOy8/3eHlDiQlnOk9fm3LERixYIkGZiKn9
r0w29bV2WF0wckfrByZTLxUB5263WkF5n3vCeZRQ4wV+z7/Ip8Bwtkcssl9ExA2iw2dmgUV8Fhkg
DZQLAPRO5tE6wG+7Xjb810TqT22IdQXYRWdMr9J6TKLyk5H85QYj4cSqOjlyvBfdEagevNWdCBpt
1RftTaWWRWrwUKMoecWyGSpgcFwvz3gq1PHa+eAtIFIpocgdGjAkIQCzX2Ai2VSF3Lp5B/95gBDE
qXeXVnco726JgoCzmu1chDiQkhBSLE4vdGKYEqWkc3pHAhY3vGyKMFFH1qyBzXg6T6+wMPF7jQNm
IZ8wTIlfCU7Kist/39Y0aPWpoFe/XLhTXpYQ3iApIWTzIHOGXJYOe/FWVyeLnxjoWpNVnWjoxyzv
6zsFdyIcdA2ck8VP3JrcdEeo+SG0pZrKPT4rx0gFepTJpvjaikCVWjuvmjlShKA5qZg5m+CgR56w
w5FO3QeXX4bcHJirNBj/7LMBzJxKPv8n5Ift067v5ePIDdTMjIGZsE6Hwxcm6hADKz+kjaFczLql
78BUOdIQduZLm9iWDf/PCvkqnCeECTt7Uwpn9sdk9Wop3VTiLvQKYaS/XIbqjhXkdrrWi13Hp3PL
YsSdhoCbX5ziEI+M0CqyOKw81RgFEigkDNhZnqKcj9XG9RMbw/LLMkK+kdcLmZSepDu7WwwASNgN
JF0kf7ANDiqtsX/9/R730YB0MwufnO9Xuzu5F7Ko5wm3e1PnLawH4LZxp44Y+bmeb8WlpxWVNqiF
BhHjVjNWk234N8oAWYPYqlfTFXp0f2T2R6L2BZmH7mMprOEJUIKRnKphTdNO7gqYyFSY4px5BF8+
J70s/PHV8X3AUVmHiiMR3WBROgGoVIqHUcRtnVsLiTzDKA0KrF/Dk47vrgZlPyYV065G0EUTQNA2
tKYAGJUI3UyIIfHe4UXJ0/E0zH99OKmJxAq3CFIfyh1FiqyjwkT95XIXFWcux836lEbeCF5eu/Sc
ODGogd+i0D09qm81x9VUi+wz/oav38Vvm98FN6gCI1l7YTasrIm/mMpbEv9aYj2BFesRpfMg2ymb
4fk2OARgkQHtP7qErR2ADL61iFvGtKqbMAInDAFEdWsjYOL2RDftsx/6AW8w86kbCM/0ONXM6K4o
VicuDmM9acvnfIBaR9gaDmM1IfVSHXRiBcqWBnQFA2aIFZ9Iym7Trxx0B0Fbx6GnxVquJ4Mqa7F5
EzjBM3wqwL9MrTlEpYVzt5vAhbyBTK3dacWtFqT59Ohk1sVG18cv/oKTk7oxv4KfnjTEARxsJIIY
ZmcD6m2Yp/bg29uC5/bZUcsFdhqd/me5ljUZt1iO7rmvGPavE5cD6tHDDvGsdJYZjKuxkH+BL0pB
jdB4g3hVIv8UfT0mTKBoLN4BQmmJwOJ9k8NQS/T8fAm4O3howbYW9uAPgdL3zraKNDGu8nnyy9Fx
dryVmnXMK3sEjATceh8MJ7TqqTcdHxg76oVacHgm6zapU37p6t/2IYB2lb5+jwAKUHdGtKNa6fEs
1yZwU37xPg+bP8ggXp65TCwQlaMr7Q7j6YqTu4ymsV7CqyQPKH1NNcRDjXS0JeY3q2GanFp85KAP
k4fSve5/VHdZzmLhUj7yWf+xrK0/GX7tpvcMDOwlJR0agg0xcFE1PHxTKVJLJNvcInCEKO7VFA1f
MnmVvtortpYJjBtmSSmxakMJubfvZ123mG4II4ZcO5nYOAP53wAQVIFvaqEsNcpQc58HB+LnsvU/
6tTc0HEf4WN3zBaSQGAoj58VVATrarfUpYbHBntDO0K+OD1lvVUG1CssBx6wO0B0djg2LtE7/FLm
BosBhVlP9VL8ROHv4Oscoq5+fEyhicKaeTcTBI6DCUvae7MopFbcfGcmxdvdD0bKYOKd1NbrMJTd
lBuoLZrex2Mc7oA7ZCm5vPdflAWPrIRXW/MUhpdhL/RQIjp0oyjUhUGvvi3E0pD2B4gRIbcElTdV
A0uN3jAtauSBLJP4rBsN37l6BAob0gK6SrdRlgOae7YNwOd2iMdNjhdRTcIbOhLpebNW5EJCQr++
GTEsvuHA+yPGXG+73/InBK9h3OD7IheYMBIwwb9t8DWX28MBMyDXBlPt66DnPqYBTr+CWB2zkbl5
E4PwyYLAx6OioYUebgFfpuXb5G5SVJQryzlpTExwHYBOQXq5dhJG338isgW4kFuEy7b91S8Gdj1y
Eqr2XdTZU4Kv95gQpX5FHd1huHHroqUX7tuSzf2fc+4hMpd+5bMQe9IWUfGK97uXR1+NlZXb7wJ6
DOpFeJJz3Xt8GGVoDM80hGssnwGVF+jIvxYDEQVgWhuq9QB/4u35/OXbUu7VGluZgfoqouzqjCPE
YeO2716cCTjWVD605+FZy0/o8tMAL3zXukivRvrzpLICq00z65pmu7lxDJJ8Q6YC5OxOe2Kq3FAH
ezUh4zWnVBRTmUbzDUtTjCCwY35iY0MIt2ni7iN1cThilmVsd9jpqZC1vrONpQ1Z52nmt8FQnLhr
3+wUO9nwWc/EoeIILe7i+02AGM4NAXfriI/O3ZjOa2hLGivkALehQXjoONqidFs1wyhq82qKMHoA
CuqlKaiEGp3zuo7q/IKoX/VIGWt0xDfDL0u9bIEI6v4hrAdQSzx/pd1U/15vwD/OkD2z92DKbiXV
UrYW9OESU60WPUuVpVROifwcbcFqQRlfoEWbx9lnu0dLPcg0PINn9XJtzvKOGKdzR8VccRZD2dZl
fOZ6vYctZ9P6tOtmUcpR4LdPzBX5rsthQjvycKQFF3+z/MpcD8IkAajbCD9z8sM1abLE2kJuAvfz
cKdYjKPQ2shQueus5evzTYk8hefZyC2vLweukvUXmEZ56hChrI7xhDYG7fHkxc37iu5t9KiXqC6f
PW/M6aa9YrWa6docMo8o+CT8vWQSjwmgh84m0H8ZwOuTXGAJGX50c58ectRjRBB1baLHXRczrXyF
pGBsPa6jl+CNjV3qTjsXiAlIjgO0Fmu5mpbjvsO+EsPJrkEBsI1/ujJV/avkPkwiM7fqFnSqORfS
jbichKGfwv86s0wnwyKQCxgDAZuIReEEAWubasyp7W4DpnXZWzpAo9Es1o70l5K7cy3U+Sg7/rc5
kmXfd0+AYAP4RjkKoKz8K833oKWjEPTaXC9BOAFuBSabhzlpjUTZhoqyKdyQtoJwS/8DHMETAW1F
0Ok/x+B6Ct8GYLueApAktulEBz5G39YkzklZcXs4X/xM52TKBtKxSjovB4FcSQ+WeMhXENQPmCjW
baIlxVJ1g5W1xUaWT72MAZnAN+xAvaEy8FQho74lotGnaQBkypzON5uWfB0NgKdfB2B1k0dOxRtO
tlGTAl3mpjDPudRkwHV1iyM9PAWuED0dVvyteQmrNUK3F6teTnrB014s3//wSHw13+rxNlyKcixq
p/+liM+1aa5ubNv1iPMtxWqk/E7+bVqxXCqj/YyIxTrNNDSFNJYfFBfcG3VaF3Ch56S/mHCcPxP/
aE5fGpa0eNBL/b45+2TDQ9XTuawKMXUF4FgqaMBhsjAfSPwVbneWOa+LVnaHle2imSy0cual3IJl
R1nUKNiSUCiERbGH7M0NYB/J5LYs/aAwxRCidKp6y4tSuV9l27MiSfBrHKmSaTbjawZHluzVs4ms
qutMtVamMAiMHHgtS/iwgMdEIjm1XQ4dTp4n1IEQmOc4tN5mzntU/RE7yIRchzsBAxb3iooT7lRZ
KBX+y65OODNMUkdRZlFXc5LZ+T4uksMDMGfgfeE75DwRQLWIVjL7CjKCNAQV3amdJhqxNo8/wraQ
/dbnAXm1h+Ly450Czqa/AwWIeTg6S9EtHgfp9cA3NmG6tyZUuhBSs6meYKvMVbj1zR+JdPcQkLv5
1UYK4RJgV4xLuu3z9HkET2sy+A5NUN1/G9xEOiZfxdT2O/W1q4m3mQqrdcDF4y3WezlrMbMCcEhb
w3fgi1XEOhEuXX7eeqtOLrQq3fXIG05ZJdeZsshddtkTM2/xpuzMOjX77JCfgNcQzFwrYvbMukVR
ZMIliMCIH15oE5csQrONNch9KNySrwfhFM0KZdhssZDwkwPdWV8+Vn6KI7lItKBT8kEbIbiTY6+y
wx3CEvX9ha3ztFB/KqgUNQvX46jq5vuw63ZxmwPMMZ7aZQ0BT+2+b5x1PmF5R5nlEhqenSzggJH4
LGovJO5hl+7v1y5hwZ+T21n2asMGYWGOBR7elyyynE/rJ7d6of7nrtqH3JVAY3EaQm1rJAa12reR
AqoQqHkWJAYtgM73xipJ5qYJT1hcjc5OEh1BTbcIcL/4jJWpK7S2TLapL9wk/POTUIC8YIamjLt7
QnAy6UKL0rmLPFTtlcBm0jM3N69IjRC3OQnAtgs2nShoqz1LrD1FIyGvOWtU3sOqg/vlxuWq3Gzp
FyM1A/ghUHF3igXXnPChDkLW6DF/l22vBRgwXtZibMIh2csZp9QxVTW9nrDi1ut4zrGSzmwV4ls1
1Q0yJwf+NFDHDTADnVPiVcBCzGyvxfpQ7FKWwQBBvz/8dHkDn/M9kyNCaie3Y70JJtR1jtd+sQeW
/qtEEKfjYR1PPkOjlOLYLfpIr0FqGJRZHu/QhJZzGRELcjPRy+4oC54hof5912OgpjIDPi9jIk6K
ud+k7cvwFUBGHuKXC+b8sVOtrCQ08D/RIUmn4qS+NJIz0EB93f69U6Fop/IGMHNUBMlPHudkIfj7
k4MoUfSzENQgumt4qBXKpb874OIyelnAmLngGQsK0Da2Y7Shs1CuwleQVQtuP1B/fD/WqMsnCRkg
Pk2L46v2IenChARP4sNl3UL7fhS1WOCGdJRF9orlQcjPyEvken0f3K/L4vp+KaQgPcgHZ3phhKDn
wwnPQcc6xH1hkDx29ZwDt6iEqc19p1srJEjHYGmHutGGBpoydWLAi5lFj8gXMoI4wAc9xN7sybRc
wpOYLzcBQxeVeoMeD+FweTZAznJ1bektX8WCzBSHdLJLwyS0oWsFyZWxb0xGbVaaXpi1N6gkIh+j
ytObU+ZtpcateH1kaWxfU8xpJ5x7T+IFo9Pn2FBrpgJh1FMrlJF9HLRcUyOEBEkOgJjpKXdjToCZ
QFuwG1BUz+pXXNjknQzCfSIURVuDXok+YSANu3USPV8TKCdToPf6BedjZJ4nB4eOD7r5D5bzbvto
0m0ZpDj0YvFImvmOzZcII35IOoVKAgXtYOiHk0bjj1M7Uz9kjPLWATsdYueKNV2LIW/0g/Oymmq5
kYE3iKbqxmZe8/MDNcqum8JGkLzFBPRLvtxnxVPqXVRY3xqZ820WuEBONI2T8bYJ+aHABYxRpdGo
1aKORq3KGZMpg1rsbyTOZsXwSCmGYqyUkjnXiI8AaWP0CkhtAetbfmRB+CyzHUQw5k6S04vTXXCr
Lah6bDama7cJdVANJIfCwZO6sJIlI2hnFzFsoyo7BPJqO7urZSHnYNL+2yjfdLbmHKUjpmbInD2t
fXVq4nNs1F9jbGesMZde/6YPJGNMvzI5f9a4dvJhXJEAPNLdbbIVFiPCApkT/Xih4AZ4sB1AOni6
d0OtES+Irq7somxRSE3AjFJfFXO6DfuBNhq/8fK6ttT2P6CKXonP0YpezlCF61xrQIpwsjWTzy3m
P0xBvue5SDrcjc+G6bffyYf/x7YV97VIA0JJoYdaPg40DDJkAnI1OC+ugJakbyrJzmR30fhIUyRw
Dr0hwzC+B73Yg9/rDdQPzWSIAppAhr4N9uJ3KITjGYukZIL8MMZbJ7QCn1M155K9LcK1rkvXsS3E
zARmhXyD/Li2LrLm/NM6OWD3GJYyxA5NKazaWtnkHkw7VgBQb7VQUP0S2IZ4iy4fjbFG6SaX0Zsj
S7T2Aee0Hr8+d0XISxcJ41kwNqbw8Pvt7mGPIKcl1elQ86GoAvwOZatGOSDk/w+DXM4zKjkiXbxD
YE5VZ4O7D26jVOJdRJAr/C5rXWZENLGIXCDmgUFuq10hyEPojlgOFp32NP04PiDxjbg2Xi+2k+h4
3rdoCuAy2m97bWuUqLKZxAkjartn6fYhjq5Y+0smdt57teLTNPQQJgu4cy/d/93YKUauE4vjgJak
auijqG2UlyRLvoWpl9tD/dWTpcFt0QHckCPAhRcG7/jQfIXYhQseWQZnalC+BsF3BZdcUCmv1WBb
ztOQQpFw4k7g0dzz2iXf2e5dJPKZjfJAuxJ4jj3qKk39Ge/P/PKkjw5GwZM1C86h/NwXfzVZC20T
NOJq+zh0a5/axpWuE5juP7RA07QxC0xskLhbebfZym0mo9i/ZtEkBOmWmOWAIvox1nJvudksqCps
xCW059LEftkFpj7MWzmv7+IOhvoasetUO2ujJuahTYYsmA4Bv8Bwd5xf9nhjaQ/NrNipDlJosD1b
YCmsu1Q0VKXqTEtUeVQbcvG/Qmyhhn9lOQCNfc8+1IMmjTcCjkzi29iCvXRPyQshcKmsjKTMaSkv
I6E9MonC9+1963mEZtc0YV3yOjUOXxiChYhuI96IwnJY9SUwHoOR6XJlflkBONr6a8juBgzZS0dO
DsSoFJ2HVROgIn8rjGjCFH8RpxbbTdgSOATBof2UEW+U8Ib7A3SZZUYfX5BdlMYuvikdr/9pcPMn
sUJGYPT2LAZEaBBTu3kvMo/vmLZXEKtmKnLjOF62xHHDRBvBIQ13T/3DhURHy+paq7U363BbOf+k
0m0wvG8zGpEPIg0E5ijQLs/mOUWK1fVFFdbZo6AdUFvTTAfpaJevHsXw57aSJn8B4uDppedOwZRh
bZlNVLYD7aNLBo0DnCrppnMs7OBNNOD0OJXe76hEeix3nqOWhAgXDg+sYPlI8FY6LK3fWdO5GI+m
bKWUaToP4MuQ8Iz/cA0nNsDs5rlQsLn7UBI8c0W+NwHKvrQPWW5eTuPnK/q/jY2xPlHf5Q1fj+zt
yw1VXTEL7jFV2kKvza8JNp3GJIuL659wV0JihFsJcdz0e8h3s3NiUqz4PC++arDel34h/wN5bE6x
3N6WDsrIbnGdDb+8xzr70pN/GhrhaUqZaUhRGTtqEA+utlY+79vtWEGad3vPG+t11owNrXgnY+pA
s2+JfyPJQ7d1joDDJb4PVmvgMiJpLbu3qxRHus/cN9sE3pNOcxn67ZQ1moMQJmyTvPehL8Fq1ljC
9ln7D4YH24SSj7VKNNrNPAmX8a5yj36rnE4+SIm1MHnL1j67CwTWkD8eT9wUVdvENYjR1ZDFM4bn
+Gt6ZV2Gx6W60Cwf0LFsjnVED+z3F0vW9VDLDkCvD7wwk2BWUG777ILO+RguOJye2BpyeqPKlu7S
SwsBPFJXC+ErxJZ5R1jcUZ1ohdQc6rINL/Ukl5XmrQ18fdeAzr/c0LH1EHO2ydr4/13wxJuyMjx6
6MhaAA13iE7zwXJ3zDFm6KPtGGFcqu3iQx+NwcYav6LrEUzKS2sLm7sBMrUXjI0MNLrGiJ4DJLGL
HvybZuWkOxLsVBdJbWAg8GLcSfdw87CN/BMsfcHsCvIeNOtq0YC+UfWPazt9gi4zyAFny27d9aLb
5C+fOa5K7f5AoxfPcZy04WRAh0JazF9gaYjyR9yzhMTaPvCtFwofoRdLdimaWLsJ0R1Mwd6ZqF9r
vdZZH3wK9uTkfXVkDwIa2rOcddzkDEzD77qev/btdVvxyE4m2OsxCDk8RDQ7ewENdFQAwgkYBBPB
tkqj0LGwr4jCAOkcrAJX+gu0Kaov6nrYrsnpkuU6SdM1lIIqbmFqyp4/eySuO9z3+LaTytNyhny5
BZzs0VhNvPDRLzBgaWLtieBstBpCMSbqfICTx3wr8EDjKPVcGyxGqNPpVY4frxjTb0aUxIS+Lyt4
CQLIEwxAx950qM64HDzwzzuOpyb+9HBmvKsUoVA6UiN9CW9ImFfhJNN2IL1P4p9yImp8m16ZYi4a
T3lcWSTPfYPcgZ6es+eejpsioC9OVy/3AnTVhPTk7kxkpmoEBuyqIIhrv3Y7wIaV3RXDNSACTwKP
PEWs4W/tSI/IU4FAohSFbxVh5tkjqz7H8znp9XXGiuqnjmWwXCWmMCTc9JQLa/n9gzE5OKRzsPI6
k5jOkaqwPa0lskeNTw8hmOX1a+rGk0yD6e8TLuAioxVMVzDIU/JE6FD8FVpZBhNe2yZJ4hjmhImb
YFcjNM6bul4Kny0e+72gh5H2WwbaD0n//Clzngidco6MspmYr+O7t1OR0DOO3U9uwQvW9hiOu6Ns
K2/KmOQLxOEAggld+GBdqG4kBaQe3VHzzlkMWBzfQ6jk3XqKA37+D+Cv9Dl6oI4oOhNvnodZbOs0
4m9L86eLxAFrmz7L576rm/v1syiViSJwjxvAAfsMHIiKdgO3AfunuMuyVEMtre5o1w4K351Zo4nb
JFUNf43jxgrYf2xoef5DG5FtW0Gbdp+x/c1ELAIjh5hbVAMXEt81fNpX7MV4yJ0ZFAnwfNhBxIUo
7LmdqeYlb0JE8/OPWUpTcEdYPyNv3R2l7c4DnEkj+CqCeVKWeEZOdD15LViQ1+W+4UnVsNCaecI+
J6gnXjsP8pvBllAbR3746pk+LUFpB2PfyWHFA3y3mocWzDIB/EuUum98syClomsELD+bJB0ZWJXY
JMkmE3+rnA8xsu5H9zDpKE3A081XBRlHcmeWXerWpauZM8w4dYcHvo3qkHOr3NAwkwkAEgHWOjgM
MNW9ulbAl4RPDx1okb+Xn81T5Hm5OE6bDJAL7inl45eFgK9MVV/+Gu/mAnERqAbMrIOPnGnrWtht
JKiLUSE5vKJPHWdCQ02s6xiA0T6eckyEX0wGG6uk3A0tFUVOXtkwcuXNoLAj0dFFxviPTWFp8y6o
m5J7tI8954DQiMAZY4j07s1WAU3Bf8QbulzeRtQIBTlG+YBRgKnpVQ+0Z+5ftp1wnQoLUVTekqTP
qFx2c9Y0eirJ0hfB6vChdlwbP1fasfasbfsUrec5jR4EzgmjwSchqMURUC/m8IzX9tVz1baEnXy+
8YnI4ykT+LgHmmYv1fNaOSauH86lM224zapDoYg/QEAPWO955ApzXos7fWHcTs2OLU1YFK40xPMS
/jGelSnE73LQqPLT9RqyZYIfc9ZfQ0R9GQgzu3c9ey9njC0CB/4xUl9qiIXlOWQRJ+npnEvpMbaB
pEoThwt+fwhYPtYLsbXJFyiVSeICSZ2+vzlnpGx+1lmqWuu4JUPMLTdNIRxWoMzCapbQdy2Xf42A
bldY3QGSDJBJqkAjb/cy9g//zwXNg4u3ODwNTLIpHeW8x8XalfyDLmBVPqaM0w1XE6spfc4HvQMf
maZcdK0by27RRFQNwxjTWxFw5zpEa6QMEhkaoU5jyQsTZRLn52NvG5uahe7egTKN9KQPMlBp1F2I
4DkMblbZ1ko0hdahiPNDKJcVdSgnClS2CCWj+7GluXRiW8wDjnuaQZdahLckskpw84vkB5sNAuu1
IIoicbTR2g9c/UNKf2x4LiymSwt2QIs4wQtk2iQ1us/nZJmsg6vUofGUA6BSAJD9LIxAgdXC7db4
G19aVy1n8bBermVCBqUABK29v7q0XosFUcke7EfGprg8RM54K1JLed28DCpYlXaDViUmY8QilUpp
9q1pIK6R8B1p6EXndxC3U1SoHdRPMEG3b6wtN1sjMzucQAZPeFpjDn3fkqP5QtPUPinpJvdNLSwW
Ba1/h13nkbkZLeUGSAYBy/wzbz15xeLt0Uz4XNMsUAsMlYN7QhxP5XQ5oM+GnPGmbQu/QMHQl+2F
j65NRIl1KpvqOTf3mfd8gobYP1RqW4wYbLDHBfWLVmYLutNVnS370g0zSluGJzJDwQuiP7zkQDXS
ncDI+IGil3H9BtIylUiCBmOVhPM8//UxbuLlSwF7XSMUD7uYfWJy8HUyKHO1VGbTw4oK1GbotlzO
O6WSbm3OO6WE9uv03FBZvv32ni0iWX7CVJ0vRUZdB7k7DuXfNDWGr/i2on0mNaMjrnGqN27akF+P
/tWP8bZCKtieNj8oAoB1pFnsnEHkph5TVtFMkZHaApvlcEU8nDtehbEfNTXqQ1zsNIFiDy9h3NTQ
oiwKYjB9EkjhXoKeaypW9KIYo/ojK08EvO3O20sM5DefDcxlmR2FhSXDeO1Ns4ajwY2/66ME0CjF
ypSKoOWBY4SpVJrdc9+yzfriXp5f5Pr3xLQTEKcNPQJrNUoY/WKuyJiQUrETDCYb6xKMpOB6h3ov
kwYHw9tsllLovfkdoP3WDIhfV8E0kRi26lGDgpM09Auc8fW0wb9NUT1Rxq+CSJ/inRYzpGwFJV6t
1fuFNy3QeWGe1iQWQRxVN3YJAFgMLlECKzPqXLFlLG7mglgdpa3pZ4EFjecuU5TsjBtCEGhYNTiY
m7j2wB55zU9b+OVt6VFQJT3FS4kWnB76HKA2xMxXiOVuVnL198LhSULqW60dPbTujrBVwjdw/cjq
4wtf9mdIH4CvZxdYP+jd//T/2UOqgc9XetmaQVvenWKKzTYNXM48obtiG/TanSNobntePwoIQEwA
hZ8lzwDTXEtb5OSLaqShUkhm/LCCjLUIe9+T8J3KGDfq0CwQNVU7qDp3NRIvMk13rfCKDvG8JbPf
b+cI9lmwSuVd47eSJeax9kRgaBFHw9SBq7nrckk4NZv3hNNEcFwFetex1RdKUfe/nDpn5EJMKkJ9
yUyqO5fE827eiPb6lsNNbgbJFnZhKJVFDdDhPEUktDIDac+Zr/PZIoDI4DRl1+Lia9diNuvWd7rX
q+2tTCpnhxB2YVlueDvLbaOgn7N89hHuGw7iFMyT3MLqmOP3LPLtYPN9D0Z4HsqlgNqJpvlZ8fdv
UpykQ/owaK1CR4SX8WN6a4MhePt8knwwmqYvWKUhT+ZB/7fQQSHnvwSW0dbr+4uT/61R9pcUaQ7c
5n8VSNfqF0MSOR4FmcsLvJDiJ7HVqG9iEIr4btpTV8hBslBKDyePlur+BLdkpnKX8gCvkvNrBOWG
YHB0wFuWi0xdJw+bh27+3fFWQRkAMMJKEBMqYO1/TV4K/4XzPtMNL2Dz+prN6ScUpojH0gc+mTf9
K+vu9fZeohp+N3u8IJzMLESqM6zz89xgPb2TwUZa5dmL6bN3tHuAH9d/t3Rk+XURx9e3BlwI2rzE
KC2XhLTRCKzB5bdT4ngRL+SYhdgAdi/OL98enZk/zrnnjFSDHtGUHripN6f2CkNupqteRioN1lns
3be2kSsSlLdMUxvh5nnsMGzrpNhccnfuPfQBz+foJfssII1vnKcc42jjvllRm/7UlaL2vlUN+F6S
GUuXVaICVOPQlgllURPZ6JNbT2qkYeL6jaue/TLILDr9n2E3RBRpd44E6YLgBlLCjEwsgjlhSJ/y
8xWttUrnqs/SA4Nk/rAaDd/GDNeSMxc81/MvgxoQRrd9+BjFwvzygPGBtETfHTFOgFj/hcKlH6EM
3Yb6nqEzFQGRcNCkWoyb6JomkswlaQHww8/EhFRwiHdsYzJktYkRtvWCGFZICITjkpxiBaUUdpod
Qa8IXTVR1946RufIbSH7n6/0mokUREwBryzT2XJfckWCQRRJ2iLxkGe9g+7IzEGFz6J+p1Hi4czi
7MxPFLHkNRILhaxkAhuesYuTs2NEskrKoJ4DLzrMBrX2IUiO6n/oqdT9/o3mx9eRMh8qyPH9C/pB
C9JpabrierLBObUpSnh8EEeIO4lLGt0MKeV5eeLRlzjnA07PtXb/GwexL9SRA77wNZGaDbUgF7Ay
+lDYn+yiWSQZbVluQc66sOodv4dSqFJ35hEFfDwDPh9mfIsK9wNMNDbTtRC9lXV0AUPzmhJz8fsL
oCI+jN+ZLbK9y1bmgP0rrL/mMnP0PYqyn0bKcHbwRw7SwyWIuk5dutsEWt4b07/7NwWi0Bw+DvgS
qb+5m1vYzi5+5k6DlaMooFWZrTZT6AJuho3mLtcpFcOdkNxM6MzV9OF2HOYNkfpT44sQIvN/CyHw
ccttfhWu6bDEId29ixn+uzw1hABjMziB+xbekKTgXGXO7KkSfK4hrjO7zB6y+rulqVElfcl+rWci
z5xfCfNet5gkMu1LwJYWzIoTJqCwIvIZV5S0Fbd7l7EPsT7OVdkZm36k1/dN5KiKPgDZLrLZyjnT
CyVIkCAHob6jqe8xlz9QIPPcZbxuxGKk1TWaEgK4wQ050z1zkCFZoSJIE3dab9vLIzUwUSDipR37
Hdk+pjpd2A3OcTJjSkPD9a+pBqzl7rtkvYThKQsaCle2TPRe9Obgnvi7K9oiPPPTDwrl5FEDqAK9
SLW+4Z9VynG1G3Fb1bWUZ50+RgKmjNFerdRntPMldwol4aMkhY6IGxBMJGyF6/vOVP5DUncEvhxI
I1rAIO4gr0LuzffJuI4AZ4mqErByqBWbK7RJ5goZQRs+9MuebiaQqx5jkOYx5TIoRA5iNt/C8CaT
vlu5eBp8B9Da3khygqb4mK+ooOg9vP4xHtx7jUp0V7vnAU05EE1TvO3Eppx3PosaSWEyRFRUBaMt
nhVv0URwyBrJGy4CJswmvs6W7FotdSuleU+7/71cCArhqA6aYcKlHzN52Ew4XUj4u1OC31g39QGA
3M/odadt3iuxpwyIChlUU8urHKs04u8e8jiUL25SFBl4gT7QsNt7qbaXEf7fjDEIxuzItQN/fJoi
rqJUFz89dP+iDT/Mw5ZjvfCy2r0Q2XGUv4TKrkY91bkpBVp/DawQIiRb9t/3VOuZvpUP1rGgC9cf
SHTnSLbOdzfxxp7phXQD0kc19pacsntiFtZS2k5kTEuH4M50mtjxm0FJAa9LGhTFpOI+axhAOp0B
w7i8RSYDy4zOaXNllsf0OO2r9DjcqLvmNNK1rZVoTRx2XzHGrQR56ZJlxtdqzZ4R4t7aXm4lrgQa
oy1O0dFPtPUqwPilaDn9z01Gs7LYo0rEymGE+07snISHRFHsBns2Mj9N/CJCfoW+BknXKybzygn3
TnWtRNtljAs3fD0nPfMoY3TnzFyXCKOyq4fK8atRu5XMEDD7XDavwzJSFa7tTtMg72xuIx6EE3qz
M+QJQVpkEBqTA6z6/G2YSOBHqrM6cRC5hqMSsnzvmEfPmZB5bngm1MSTJK8CFuu2B6qxOqTB1/5K
jG837EQiLxmEwwy6eERMVgcobo8iYdF4wocwZXxoBbjXCSyz+ozDEokgKi8az9mD6n/NhyaS1TKq
+7no4A79LPhwzBSyqTaw0nGc6gS6MclxBrHZMZkb9LGfHQQ0WzHm7EGuntPrgFPifBPzhJwK5JNd
GbncGNNiit0INqQzExgoj3Iax9rQH1dDiMkH2NIEMJfCt2X3IJtVMdkUAS7ejyHJ91pt4Dnbwbfu
b/OeHOmJ0D+7feBknxA2VCJOSc8jyZZA01+QEB8YBSi1HqlRNLwqCQVFP+WMQ8hC+eIU7VGpbpRF
YHVBqTyJisXytQwD/skbPEq9CJ4dkFsuLdfxegJN0TDxKH2nVlXWxsKP4+b27qY2HiRaReh6F2pm
Ati9T6ONy01QVi8kP8P23JRtN0w9Zi8VwzeK/UoUgG2WT96+6YqYmmLdWqbZKuwmBt1/9jWq2Hhw
g0uYMY3mD9wtwU1apoHr37YDEPW6mDQf4BUD51qz2uAYac1kK7eQ3eZygRyr8BgBpdKN2vlV08mc
/iEcOdwkUsw917HwbCbfL36NcKqfLuXZZ6szYStCsH1RDB6jCWIRycqfq37ABaMVLAkuFI6cP2ly
s2eu2+o/lA31FCX/bR/d2M//iRnmf4M6vWVJoA54XBzQbLkrX5882pf8R2XlCgE9xZuQBm/0zohN
UzgOK3ptp3Ekg+42Z0Adecq9GzSOGyAoeDJ8k7t5EUrCFxeysF5hRA62+mF5AkOWG9iwRo9209oe
HPT5bGSbnDIsRuatU8k0fz1kwnG1bsAeN2rQYeYxY7U4TDg/q1UkrlKNjuRg8Qg9FL+XpGCW9owg
9JsoWujYwt5JPexR8reYNmtdWoZKDja8z25JfCxmXa3Cp4bXOzH6LiegzJrsQj0o/FWxdkE0+cpX
Ne8Sd0rRPRIbLoJ6sQkyDhpraRi+jJwuDz2HaXM/f/zPRVE6IIs7xnk8F5f2umFtLaXDYU69+mZE
e7beS6k8iOGXtUJXX2SHhOl81XEIknT7FqcsVDAOp3q8AbKpwYJtgtjgJgi6jNqDed47Ih28oePz
47dwMblVH4fr6KwTQQVI9By4yo6wtHNMxXHsrQ+r3CzOd8F3ebRWMehcnDnwJg1UCiY6OQpcBzrY
ByOJ/osfPS+8KFLJy7l3D4jzJk/3jxKZhsKYNy8QRlhNuSA8lTNJX+x3W6GNjOe6LTRUgLq4f8Cn
bsPJsCPp6Ur5AOaRvJJJrlJMYpbBayk7FPXysTn23dkCPa8fuGWZ5FRT1uQwgLJTXpnN6AWAP47X
OFtR7OKtP0ukxSTOWYaBt5xJTI2tUbdiJDXFVMPny3VLZXbb47Z85qqesz7gp0zf+8wdzvCWh4d1
oQBxLg/si0x3W4dZUZoVBNJuYwdOtuGBmKHHs/VhWV99NidQaC42ERirJPFQuLZg1MTxkiZSQ9ZA
rw+36SLHN69NlsQyubXL/yyxXZc1CbiGphDYo6GWV+u8FA8Sw1IFaCtlN+B8+4Lt+AUvdNJtex93
ELEUyN/WUFaN5uUkVUFfQ9LcpAyDJPTx/xyKZ+wZZH9xwND9KZXIpuIRfM01AY2d/F0WjWQpZjM2
yAfWYhfi/D1FwKiAnvYUK/X6QNkWZgaOGfLtfIjbDxG6i32cUH8SBjgSujhg+cpfytrD+7TnQ5GL
hpVUErH+t1ZzTZKqngc2jMA+gBxoubik5eFrE0wn78jiYUA6yVTy6rMhnYzMoYq6DiUVeSbWBK9r
ngEvDnBpInyvSTb4sToSbN82mDBeHCUOtgLx8TNUOX7QBjEB+oI00cyosUAIyak0KLcWjwzq2ZjM
QG1Eqk0elK2iE1C5vEGlOGuJ3/LoUld3fxSm3SsNvCqpAWZ1tRnu3glfUfnwFTaFge0OT3DYzR9z
A+q5JIlSe6NXsZ42rVTN/XBtQhUk4eJ90h7JKE8+eeh556P1aNt/jOmOvsO1RFxTOCmXRZt5oD/8
PQsnokzNMXveevHEbXUaggIp10LRwAAx+4OYhUaGngPs3wDlPOGRz6I5cpHB6DRoDZxA9QOo+Wr+
PC8RlI4gpL1vm1/KDW+FMDJXC9q4PWtHuoo0YX3dxjPhxJM4LM5BddrE/gU6CPJJXmziKhx/C4Rq
K9a26cD2j9mdAcZ69phFYTc3WN2yVCFbzUpXvGVuOO3vEos+KPsYUxz/5CYoy7GhyAWycwGvMTkB
4LWBKcjqKcylG010iNqa6Pc0TeVi17/6VtsJBZ2WMHwSJOcg07eL3b+xUezzZ/XVnlTYZ3sd5ySd
lK+q5fD8wZMdEgrC7x7i7TKd5dnnOqAwBbHA/AE9lhWh5cqWY+rZADFO+wUB8ZsdtT4oT/o+KtW0
C140/l5VJDM/c7K/rLoWjnmIanqnu25h6G5DNF3/t/BN4nMEYgZXMsGKC5rzZCNqQg4BywEpthbe
VbHedcjGq9Byg5V2tjeIVDmFpOkLlai2P9/z3otT8KqYWsv4f5lgCkFLFNljATRngdDJEUcbCmtH
8mPoU198UpXbIDIQlCoGGUyKs3PBPqKsjz7citMu+9nDG/VpfsFP18gd9yro07LvtWJDuPgmuZV0
APdiP4MTsPyOA93RcEZ45QCSAbLkuo1eV4HhwxI/CSFgZN8MUo3Da/QtSaSZS2MKMOh4b9fvFwlo
sUhBNy/ipEO+jzJQu5AxeftvtuUgXKl/yW+uJGRdOEmh20A9sKM+2T7EkTzWba9XAQK5fWWzuACA
OoFAiKOS++KTy3RdJKoQG25iUAsV6rbUMXg/wcoqqTFiP+uOKtSPJTddj9AuEDlg1/dkdRp2aLcs
xgx5AYBrI85T/Ym34bDnHE8NtUEFq1ArMspLJW9Kp4zCciBIFTiWVRiiY4FXg/edM0V9PRa0C5VH
4mCKMVpX3LfMSOwY6i9Bjl1sflXbbFixuW72xXoOpiOcTRMAh21eYT/u+otK/aleHGETSOPqP7Z6
wipley0vSysOZ0OOmSYV+1VqsPc96hrdIORuIPvbwrbs3byWta7pqwRwiaLa9bUX2SHXGmWpezli
fyDWmD5WK+CNmOYyJhRyYCtHHnM01Y0870wPOnrjd72UQQ25CtLpgFhAKu2mOFRXfxLe2EwGw41T
gtkOCyeQW1KOzHRYDLwO8PZgNT+dMq6WMLQGtChQ9UpHPrK3qMnPowD2Kx1tloUChVWKw9zXsGpv
bu1miKVWAF+2qho/XKBex2Jn6hVUIf9pyB2E8q8xQfR1+ZzSz4K7ClbTI/79QeuoaNrxB/epxrs9
LXPa05/KnQvjzNXpaFNCvxsbifaFM/GU1EYTP4FqF4KzaLY7onut1iSmBsUSYK2vkmX7h6rZRgr9
C7TGSwm/oT8+ZfU532wB+8kcyS/VbZNRlcX3IV9HfOHZHkuampLMsJAaThHgig42fao5rJDlSbU1
KfMHZkQviydKiVSQRK79eR0akT11w9d/+V/bWGuDFWPM411wtiBv1/r/qm+X5vLPqI8f/6BS7aTf
1ApdG6v+SybZs05ELgk3TkuQuusZerJtVnWGXVYe+Nnuj7BGp9viuBzvgLythYLj9TkBCrRPxDtN
v8/iY5W3XWgDPKVxsi5Oh7pnfkd6hU7cihb6KVPHvIo4XM/X4VYXTyo6ihN5CC+pP1iIveCMNyK9
+aCc8ACHGXUvRVLsx/5OQ6bpx+pHjVFxE9IJ5ubN9oXKqNjiscUJi8KGmxgEU00stKp2Ax9JHDSj
vCbXomlO7tfhSKJ2XYeDLBrnV4/ypv+D5Cn8JSaHsvyal1VJlytdVi1hivJdmZk3w2IfDqluJwrb
6fyuUZfrugm+Vuvntuv1gBwhXRXbuTK4yS7AfRb6LnC3mUE+XrGwYul5tFuvla5SmdGljP8R/pWT
WPSbzC5fLSRHnqS7ipZZajATwCeKshcSTCWlsu8hQLAmkgx+s/tjGbNn3TUor+IuyiKjiLcCHblk
0eMZUA7rUY++oHo52i95SpddF6P3w9D/uzzxoiKwrKiuaORrrmR+6MRNYI0B0uIhW+Y5rXdDkdIJ
H1laGhGvWjCtD7Q3S9RA4ALlfW/aqrhQie70WADPTlV9bs40zR2LYqKlHK2/Dv66QHhnjLCTiknL
gflPeYhGPKdkCukD0dw1ot0+s5t98Qp6Og16GtUvHkj576nY/gPCHs34cnmZ2OQQxTVXzFpW+OUd
8oks8/akhldPJh6uZ9bawaT5VdVbwlLwTXbZ/IWBF27lT5HQGDo1p+hufpOV89/yZ2e69VDyk3rH
HukVRtcA7FwlSVEZDTfVgfG3goqf4kpgSP/A39nzVBP4nr3Mp6os0cx5BG18RfDfD2QHZteMERSJ
puiCn6EyhfHUT7mCHP4NN4zSepGCQzVtt1ahm04YserJhYNY4O3/m2kkzSUiMVepn0V2DuIn450Q
9fyqq/xS1Am/cEo4ys9OOuQ5v8SfL6AgGQ5v9kr7c+bw+gZ/8K44G4VZ+WogcKMzGrs39pgh6w0v
qJWpq+kltwed17hntSCmsCkS2U0+sb/X250AXASoLHqLrwdx05nEuaEAx22wafd44y8GhLAmEdNP
3C4jrGQoCRnGJjcmdCM61zbWjsoazYoMOl2fub7LwVIzGFXUhO4XmjvkawEWwqtJlLKUwoEHXSII
dhj73QjnvlUAnD5bewRg53MHc0si2z6r2Iqp1a1FHR5xeXamZyZjD6LqCQd0FuI0/oct4B0/tv/T
HGWkV8EJ6an6+0uIoE0D+CDdnBu9oDMg1cFEb4ZWqs0h6ZyaCFa1G75jXsbm/kJmxk7VRtTKpKth
u4XvGKEdCPKwJXfFE22/VyaPblQPbCjjoc3XxeAl1/TFjPYBwEUvluk1FfF8lQwtBAeA6p/1gPYu
mUWj50ffOpbS+CULpHC/BcXstUJNHRO3z4JxFYfB9qFKObAR+rAkE13YOZVHIcZEnDc1pvxRjjnp
om2+HPkPGwXnqyUT342XyXOcdW6ydTcIxiYO4jrgHxnUNOLJ3lj7gPh8JFSAsEpq/98KlwcgUNyJ
RnU863Hq3pEcFz5TfE/5nkrnAZq/f8bCdK7f7udaY1GD8GGwdnAmJMP707qjH1bwaLA6Pk9QoGuW
LqztBhMvLcakEZLEBlptOSPweqR7veuFsPuo3Yn/O9Qg6CZpGcBYscphL+VtPsDGbozMIFCAN/YE
ZAmXpBbiwcCaVYeZd5/NzbufVuww3EPY63aZ9Ty2CZ/RTt6QW84wVyxS34eqzBAVBmYBXVIhwvV/
c/0ivZ2jM+kHZiwRadHEVeS3vONj2sdpsh/lg8u+ogNxPfc6PjT8mlxcs9Sf83ry9t9JHRrerumH
cWNySNPPqxngwaPBkQ4yyCd6zc71gb6WfaDLC4LiQuO/LXcdqovihbMRaWBc5MLYgfCYy3hG/6ib
VpPh7iRJx5qmuxE34kEsQvJzq4q3PcjM6Levm/oHoidSSRP8Se0+nUXvwmGkWX0BuMiGF8HkdlMM
Xl70V1iL9J3wsoP5IsnnxAR3sBVbOnVf66hGurYKTM0AIAK0QA801Sq/bmewDBFW9IFcc6xiGPHG
do0u3ytaw3NxxHze16QAv7z/ehmK90OvhTNXZz2JmrkOR4St9EmSXnJwwIgwgbNTS1eonxkzWTZ2
TGtsRWSZFWIVc932pICttqQtISUHeXGpTs+WXjT79EOgJ5kESGCYadyco0bvjGxJxgh6k2TPeZcx
g/mML5g2GxzYHukDo/LzYbyAa2nkiqH0LPQanc1JApca39+nJEo7LW0drHqWR2e7W0VAeFqLvcte
+OTeJSMhKQVLEoIBoUBTs1wy0Cz4mvoAaPDiA7JrmMZLNoa3XZcV3lok33eh0KTrW2c1B3BveUIx
Rmw35wvfrXtFXpmTKT5XaREOBKTVPxWJtx6ncW3oJ5sFzxenNOGtsUPD9Tg319uGN8vxEhmpdQjA
/jeK+QHLxPchzlKuhfnaKZi/W90JKQwqU3o+TsK86MHFY2veVG8IfK9wj0i+L0zIFh3o+zX5uFMY
pyMqfHLVYAuxjgLlQKCTl/w4gkwAkkw2U5c93omquIRIGhlMItBXgV/Ggj9s3kc4sk7JTIWoJW+d
RjGxQ6xAIepfJnMYxIT3gCOVt/Cz7/ejdb4xv1EgjfXYBfVFMggUwsMqQAmxt7A1m4LFb+AnnqWB
oBMAAeBBvOTX/hHI2lpWEfy9Vc4qoox1hxIH69CYD1a2ZcQD5sVUW1AaleFZKoDH5RVdpdLIDTaK
ula6ThVG4ArMDqyrjangG2ycrNkTupvrEHqewvLAyKP0suV0IzZYv9+Ztj2wtsYPJp35FX6C94x9
vVP3KtDaSa8KtwMAzN+XMIbfE5JHFK570ZBnbR2z7pDwYyeMoC1LzcWiQX/b83fpa970VcmYgQkR
3qlH/8JOWyzuEq9imWQRQSSy5wl71M3nmgQvNOVhf1+Afb3uC4aS+Htk30vFPMkCQLOx/k1DNoN4
jDsjeFdOB8Zfr25Q5FDQt6wjYPWUmNZ20pqmyzNK81OakHFXv0PXi3YZY3hsUJwng3oeo6o2FIKw
KN+9bXLpyhMEC7TLO/qCtxtLPM6X8/0CkciNkiRof5lHkcvpgqVityE6uUt3ILCj4DV3nz/7W7PB
jp1TRNml3xKkSQ1Kc/hmgW+A9Bnt315hblzzCE76XTo+Rvtq6PIaxh/n+8plo81vjDDU+M7PE4HV
NPXLD9b3pW3d3VhQ3jhGSemDh1Hlr2t2AXijR0UxdxPVnUI7xn9mDHj1fKl8DRLLJH4rkBg29wKF
rQjfNDPVcJvY38So91biJJrV4YzVtTbtiWz05BGInDVYwx1aJGwupm+dLrb8hNJau0omRm4TFj6w
e9Dy4kGl1xaHHFFuV05o+d0cS5MsLVgWdHqjJcfhYD3a7rxdjHZh89+w9x7JxdGNnAIgjnjYoIXG
kssMdbldQzdCm5wuWYfiriHQrn5I8V6pmdppJVDAc9nHgZ+mntObmqjrisGDvn+ARSGKeLVJWyNk
TYl00GBq9YGxqYn4OD9BLayglkI1s9P9slfY83lJVOnzV5+WXGSJ/QzVWLyyOot1Kpynpo2ZWVnL
Op+N+m06b00sxXmtCNUJGFsERlK/xV2FRsDVefCQUxHEO56j5h+5nAx2Bewq7bcGFyQ3f3vRKS5s
/jLF24x2/z3aHUiHYjnkZakv1XQdKBT77LcJrZ1ANJ7MF2Qxvbnc9bMVEBOK7zjqgkHT6SI/umiP
nHs6b1oaha28rEsHAtezwuxo1NaBFq1FUhTghQTxoDgKGfBOfiPGHe4MK78m1LvDYTJgpDxHIFI9
qtif58KsS9bC0f+MmNUfzTLwMspx1/engs9aClZ2dGCNGfQp8vgQmUHWsosuxDeqzXYbXvtTx0KB
GqIeYyT4vgQhvWHrT/eXYBAoUbqaeyrYI8m3HVBTCgjQZAcu2tgrPNtvdJd4Qmi9S2PRSphslYBF
5IwRUldpj2gUqYgueqnxi5tWJn/lq/Ze+s+StD/g0BWiW80nvUcODRMQ4dTAbETJJ3M08Gmpfxrl
jOJd/c6JHD9+5PseAH4zRNNHLi9Tv0gvkqhytnuM1ygpqwht66pcGCScL2bNNhWkwvSNgSCn1e4y
h+4qEOBIpMJ5SMO88OKXpQN2hAtCulaE+QVfOBJbxSEJ/wFeD4+2PWRB4W2IAUP7wAxUKQTQNEW+
UxjqwoPAAnspKngUA7vZx/yKj+h+xD56TaCdW7uPD9O2VE8hY10IT3piRWT7teaKqzV178EkBs+x
RKMGDxopahAbjotS67cag0wy/jGNmZh/nUHKAnP9A15d75a3CAeYoB3J/tPU5W7hBaIY37aMJ8jE
1nT2vMGLOx1keuPEgqoCzDg6SoAYOFjYMPa1V+fzoziQS3XgbHAAaopT++6uwdNf8H1HYuEtgxyi
f/GVbUonFjWULw4NvdnEs2Ss3G4ffIix44Bev7G64igL5LW4QoCSiuSmz2H0Zumz89xH6bqrv/Ft
9K8OJAsQ6DACRGAodjXvfGsF3B8W1Mj//MCk6MSWyRpYumQc9GDRSx73uRZQ99hu34xE9GPCKcS8
/M3dIGoLjkbPA4hhFxu3cr3MBPyVCTp55sfrwJsDcoWMAd/s+i1Bg4hc2gjNnOPBCqV19eL3Wkb+
5UXHR0JeqRFpDuiaq7mRc5tkS47gBIs21+i5/oPj+XC60WumpAFtZ+SG36vWXzTYY+dEpQyhgnKR
d1qguvJVhtbd9YXmKzaKywUBHBWmQ3UTWtMX+AprfalbE01Sexaepp6sEs0tYmioNCO78bPAQrGn
5JcS6XjC4gg7NPaqYBdW4zfpdpuScEMTIT/wVfjEKQCkGmOr5WMjbsAywVLE34avdVklo3hs5opD
xa+bSN+bgIUDcagBYnohKA7M/TzGN4/Lf1Bqce7P/qBUXyIU37JhHmTvZuf/s+NfVzuc/IdmUbYs
9uqJup2g3TaP+pGLWLDaYadmt6ZwGjRDimzojAOpohoP2UD7kWPFTDTAw4LWhpANI86AcsHylIwb
lL1599d959o8WJFgna/5N7GUsH7dTvsNHv7uzFDeJ6Ju/OmCWSLEUF4D9D4k5mGn5IpXfgQt2egx
fbnxMLzZatUhxy6bISEP37v4PPhgQbywx41LKaMhTtQ9fWIeqLqUxy0PIEY4Izywg+X3uXkjidov
p+e1cCn8rE593QZevD6UXUbkB8rIifDTyA8krT1eLvM8EP4DTAk0H27jwjvx2V2WCD5nsfWsDOyg
JJyltdnfzcfm20EBEGdWo9UiKex84YTdEbtZ1UmZx4nG7ZsEqdqU7dbHXSlEScJ2z/I49gOnc9ip
kyUynFQaRJAYLIcluO2awkC9DDxgk3tt0NSGzDlY3DelgYduNJ8sqMW/LwvFnY/p1hxaoq7rufHc
zqxMmGzAgZ2qgx0sFvVu7lqyspzrUIAba+291bRO+BkfFz2yBrwBpJXoNNeoRGS8w4kiW415pnYC
FYABkl1f2o4lSR02gcAxoUAMXNiz0pDRTmCVzp9ionFEIPA1eKCcoucpo+DeMy+YyvM/p+ux9wQb
tvosqq5Ufms8AYmvtoql4/EuKMd43udEssMakprkmKF7NXGqtGtYoF7xCoaf/OaQ6B0EqxPTzbXR
G+qgLzOC36ySAB2I7f2d6VUO/aLiIdEyRMT9u4O3QWqp9rix40nWFiCZTacunmxdOoAoUQtqubGQ
6GXYlvWZVYOsAb/vg3YQBjkCyvnJyaXELkHfvtEeNh7f5llaQRG5qYiViUarKBPe8Y2LrK8Lv++i
WRbQ/zAcC5446067eeGcPt8GgEjX9ucnlnk11Uf6r+LGNzfpP2ryzecGG33cZqnG+3EpDvR0GiBA
LirGUp8sPYBe44zEx7KeQUvDkQtC/b/gI08weHv5dUJKM1evYc2m6w8n0WKCICkXrZm0vBTW95RB
o1fojtyKY6wsjyOduMTqUbTX/hiVD5ssW8Uo8DG1mSREEniiv6xDnAThO9xsi9Yxycrbq7SCJrJE
W/JwWotS0oidPnc++IhtrQpZGgWkTVy4leDQ0iNpdeIwZ0JcxAMh9XJcS03Qw+wUSYlxkt6tauBg
Cj1usWe9G+BxrzwZmvbDsgbEtgoz3h6c6wCeIBlqKxtIe+/s6a5cPV9q4Gm7t1Nes2bAwE03/qaA
c5/IrjFJ9JIKfU8OIRxYcJAF9cz+BedWezyXWAlURVsHNPEEwceFW8fMdmOpnsz3FrY7GKLZfofa
gVx89zAaNbWt436Js+wirWHq0FDPsJC1ED3bQg2pSXU2XgmXNpWSGh5s+HV2qsu/A1CM6RmWbOHi
Hpke06J/w/ZriOC/a0eWR+Aw4nv+qplvVcAwdJYk+4CEB4z3TIM+1et9hiv01to9Lz7TAEwCmvQO
X0sjFlT3hM5Jsn/P0zoBI88ZvGRt9JcF4KkISmYj32PqBI0UWHvspkiwjS87dTcNFBuCDuCLQ8yU
HV9lxB5aiihHggf0iWG5NDZJ4dTkLti8HbmtFZcRE6OdrIKJ7mYMmMrYuO9uxnO8vKTAUc7LJqem
Q2zlNSO1nNbBQ2lHrmENJCFuKtXMNYK3mnhj87fD+6Y+DI4MzAp/MEbwSIbaRvXUzOFiDrWBDl3T
CvaewQRd8NhOjGVc63YUbDnnb1JA8yiQqyRHb9h39NP8Wm9lB4JvkzHserx5uJRZ8jOdTHVDYwfY
PC4WjE8oEYrxDFXDmIOPsVVk35UsMYXL+7ayMMNE5EUHlsZZtT+99i8BKmaANHfpgg4ppmKET3gM
6Yz3VDQ8KOuYURAusAl3qQlREJyZquJbJFx8cN60EBXjbQiK5Qz99cr1CHzNaK9yJhRGiRCEUM53
HWFrmW/edc0MYJ/qLlGRIfpyRO1JNc5xZwzn8vCONg4GvVV4uhoveXYanEROIMWFk2ADsTNDMmdt
0fZAmmKxVrAlK5uLeVmWz76AAdKwujJVz4Orq8/+ez80VN/Sm58XpNsGwd+3E22ybf5mym96YG4m
Hsghb+HJvcBerdWOAMYke9WumMKyKoq+8j7ybCco0Os86e2UwGdCbB4azwCN8dffgx1EysLS1k5s
ANZ6oWBcpPqF4zwpntupvw2aNQWnjacAiTWl2TLjD1rOx+dOU2GoeRNMYo2PjTpAiA6CXGtxkV7o
AKiQK3eI3/IdRKbb5DOwu0CkMB4NQ4wTBJQRsN/3snavormcVT70smNMEINNnF3kWA+Um1jdNf8w
ox/httL19JJI50rJ84nfqfGLzKg/6H6pgw7Zro5Y7gD3Md5//NxlHLFyxcIaRUlgdWZeQEncczwb
OfSg5oAid+CcGUppx48xeGHf5gHUT6xbUHBV10mGNZ8A7n/UDazc3iDmFG9GUWl3YGvHnvUllonO
f3XNDju8C5/oEi3s6+9spHht5ZnOL0zY3gaQBdkFqgjC5vdBWw2jm/drd9e0o7AeGeGnB2p2JnaS
OB43bl3K3Xjad6fFyb0q2IWo8EkHwd1/YreFrErUFQQiztyNW7ft0oIGkRc7lCM2NdEdvq6r8jhY
BiRXwMMcRg895bwuVSMy1sWTWRhYtlB67L7ZOEhfU6+25HFxTE9qmxfROUccb02QZuNomd9EGGyP
X8GfUfqsnc7LPA/4lxYyThQ6LoCmu4GYKZ/Q1DOBqZ34hNPWDNlTKMZTFbgjRwh2gGBOGzsMiphM
GxtBdC2VEG3mzCfCv3vtlyfuly7lukOoOS0R6pqR/bTbIpMXl5f9nAby2G0hIDl/CHItbJroCg3g
LwscVxG57283W2ycitRehlSK+AcyCZ2Dbq9dN2gZHz/4F289Y/52jW3in9HyElqfx7nRCMqZJY2e
9nDyVVbPgmsObZvnv29u2eIB6UB75Jd5G7SIO6GhUuAVnzrRLaJRdzlpH29BP3EnDZt04+VL7p1S
5TDgc0zXwT8KWq/H6WGzvpVCEn88p0muRTA5L5AS7J/kMblBNryyydrG3gvbYkl0lV7wHc+YSP0G
JAkhQtuHLbrtOTr+c2pEVLB5kijG0jofP+M1ZAoCed+nt9EmxNDWhBOGuJrdbrXe8V3j0VDlNfFW
/VieaTRwx4G9sBaN6L+mzsZNZ2QFoB1+ZqUhqcoUJEcxpoHJNs5PBRyZQdFvQjmYILMxl5jJh4NA
UwW3EhZ20mSPGL1gkYUId4VyBALZiNjcK4nhXwyJaxAj2nHeVNyUQctlIDWdWCoDk3gQH+yucdPp
RZnHem2/UUeE2SLSuHF/RpmJwb/WgwccS24X5EkX07CFeYbF/+iYb+OYMrPPGDdxt3sPagiD/AgZ
suiqIh+TIZyboNuVdxGNivAyHO4n6negMNNEFdI6UzkDtwnHjFo5eVwsky+5jSTGCCGO+O0Ssmdg
fdcGDz3/CUTPYpTJHXOcHOp/TmjuMPY2vq/+F99fmtpRqXrAxpO/ZNOoM/V0evVFxw7lr45Uqoji
C30pwIAVs7pBLhTtLIbNP1pBkpH30MmfGIrSHFiu79lnHRSJKsVaIA/HW8XR+4Um/l6NeRTE6Nta
6YBEeJTl/DMusQuK7H5cl8bhzlR5eTXLAwil1XJTiuXudjOYadZK6A1Gk1d88h6re4lYvg7alGyT
KUs65OdgyjElKoP8tpj4XH3ncb2STpeW3U+5jVEsWoUeLSRs2o7WyljgXK5C4+BbLKBqgOAqAKkH
ANlFCQfPTHmyJ+SZqwLp2/+83zlTdP3uUSQAZNTiSZkCBeIX6gaKXGatLuNHYPh3g0LJEcdagxyi
gx8jwcCkeZHl7aWwMvFBuOqbSI8Xw4NYeO7vqcT59pQaLDX0Kp/waa/hmFME2ckCBqP+krjqKgYU
9dxydj7jDTRDiyuCPSjH3BsU4zDjY6CQ3GETk/4IP/QsQMdDwhOyKhNJfCQlLVhs0ArBVfJkO0Jw
Khat+7hbk7YyYyZx09u3Y72P9okAALR4Qg/NvOYjbWwKlJ4wx2+536Sjy33pELJO26RGQMhkd3+9
k4e9kcjLNYFTgNn72lpSCbHA3djiCbUptCY0RnBw5VTe9qH7bHbB12T/VwEck/phjR7DLLZ/x5hz
QUyi28GEB6/V8UOfQjaqyKSkF/PeHxzXAbRvJiY39SXeSNrwZotSERKmIqIk9q6plL1yk1M0E3Gu
TSfd3wHG1jARVX4K9GiTPr0Kr4fGOAO1fpC4I20OduL4Sm3KZ2i02WBYQctfkt/y1+icq2SzPgGT
5fFQmi8Mse+wOwyrIfZqYK6EYJVaqfVJ8lH0kD+nos5mGhJBSOa/MaAf+f0ayZetdcUznnK9MY4d
hmKetiATUUy5FL1vNKOW3+xvwg2dPdy/byBHtjw7i2mDwhcaX5arYUrL4QfNeV+TaX6g1HlCWtrJ
6p+u0yIf2AyC5kPlK8/P19xxphxaYjKyrctDnVpYU4neWrgNjTXZ36LaFtID8pJQsuvffqJSjl6i
n9lzpZZ7SQEtf7Ym+Jl/GsAcyVyNYv80foji1JlVFsJeSIZ620mtoDtf1sEvzNfcWClDuMYC1KKP
GWBCU8iTom3YBKusttUsWzr1MCloXrNUp1bHwHwGcbaN58GvT9Q65qTBuf/CiQ3MD6F6adLb+lGN
m31y0WLRZAkbrnpiNPdKT31mEYvUrRdClM34dFPbfqy19W9OHU2sNzrEjn8tbSUCdh5lnn3OZQQh
MtCtbz6frcslrWWyAq9eJRxKRhuspMwqVTyaCgdwjfO60T84lBT3Tde+GzC1LwkD2f4VTALM4nfp
+r4zZOek94JPnTRWj5K+Mu2Dwh70oag9/lXv1W4KZ9d/eKV8oFVwbCeQh94LBnUteVTqxdebz04R
uB+DYYYW4MWuaVsN5ImoeKjqKA3hDHrSRVGE/spa18tZaTbNuouXFjZ5hVtcBRPs8tiJdFyQI9Ua
4NOEsSRybkaZfYLkqpPghZr1zFm2NYvBB99HNnmH/Z9kRzOEmcU2AlCEF1GHBgyf4fFPAjOKItge
xkj+GGul0DfmLBq75zoig8dxjnOydkxCNws5RjyQ8PXvnttsjrgGGNsCFMqQzA7S3u7jIts/7vC+
U+9GPqg2xqJ4Oa0sEyN6KZryanJce2nnLb9PtIlaZCaOdP3OcHOgdaPB6Uxr9VCEFZMj9K1jM5LX
HoyONCWdN+8GkKBVTWQIuEB2FbAEEHTHoLtDn6sC8arpIvImCzUrrXurHfVrPUCsJRr3xfG4+hnJ
gxzBptfLV6lymSycBXfE/yMLOCvQSeS+c+n9+4OnIK6kHYSmSPP1Rfzd9J5ZyUd4uiqogtk8IK4t
QPh2EzFnf42LjuZ90kAcYwqhAC0D4pGs0gI4kez5HB6gzJdvB/xViHMexxAuHm3VSzVrbyA7FE0y
gBoW+3fLcCb6vmmti7j1QPz7XrhdiTzLpGj10Nc7eaTB2IKZsUXQFEFrEyLl4I+DCjscwKm+MzFi
pJ+UH9818sLPZCP6+sP5pQ6Wv2Y2NBZmECMUkv/f5qI5EwP/rP3YS0yi0BSTDnH8905nlNIItw2i
ypwBcaJi3tXmmPG15Lsnykeu/cRbKl54pRrf3XXvMpZVb3X2AMhNk0GaIrD018VdB6PNEJFx/pWE
E/OUNDtioobngZB7Z0s2GnMXbYV/O831aX4xVyi8PbY3yQdnjP3rbsWgcUH3q03v/cP4womTuEXD
KrggsK8aQywa+Obp1M56vdQPOE0Afo4lqMOAxKLuYRPK/ghIeUS4+HB3WqHYp6urWfNwWWnOIiMK
hf28Xw+dDC4JO84kQwM+45TMq6DRaFkNlW5hNzT6/ZiyAoNPwQ+V3HsEySJDEewnngxJQfYP9cdc
FfY0rrVbmjhLA5SZhg2vKD9YC9zFRTFqqV4Heop9Jj+Po/woVdHWcp04sqoEVuPzVSyakecKjkKB
hDlb9v6AzKpmvt1f52baKH7hSwuaY7DHXZozXwXFgiD7wt+6ybEqhhK0G3/YfmmJJ+Wd0SmZGHLC
bWpL0k9cDeYEe73yaJCUZ1aTsXa6f3QoSp/0Vi1CkhQKPh7ZQhMyuxFjCASNvufjuIGcGFmnyHOi
cEKu3wd5Kth9xKU5KeI76MGToHkV3IkWuofjITIXJboqPP/5pYyxxFpmgI8vw31LWOFyT7hUdUNi
mPc8OepIG2CXyiT1o0PO9xVcZs6Mb8U6Rxq8UupvwiQCXCJF98xdwRqIWFaVhPIUzKUzImExtwVh
0aiN9z4IKHUYdvk2CMTk0x/zPP8mwWBLKS7KcgW9mXf2uyD8cEPV6UjH24LyiFGvrUfllJolexwX
GQgQjWACEM4aodnZH4OiVus4ylCjtWOJdO4qFoR0JtOZk//wxSzjTQ3OWu9ylLwJTZN5GcLnB2ya
i0noPNnJ/w3BJnKA9blPSytDdaEQVHtdJ2wBzlReVub5hH284jaJIu+VnH7toSx0kFU2xWebscg/
z5gmYzTVi8tDahp3gCL/Nf13HI4PtX3fLkgqmrtS/BkWia/b5977FyR+C9wXNXlopUHsewa5Fgr5
6QsK/7sn9NZi6ycMn7VvbHgfV4rj0OJY/HGzRHLU7FoPqYvgodnCv0WpLUdFeBcsZjCw2vooh2+z
r5wya323GZVVto4VtaKp60G1IIT/3IcGzaF1FKD26nda8ELfrELKgAP0LmDYsBYE4junRnZsbqi4
IsmAA69IZ9ePjirQi7QjgLxRMVuPVBHxya1awAJRrMa61WuN6vkngrH3KhNnPKEMhH2w+IjM63wl
DkYiUz5Cj2ipmNJdKwVBQ3Gt8mmRKym/SDqImIyWZUINdGwlQgMfIHiNBIDVOWOcvnqX1i/RxHvF
tJsia+LgMGFIx8XFiZK0nz3fVnHgOETgnRDbI/XvdsersZ3/kZcKX9F+iuJG2J0R12GhQs9QKcr9
rxDWHOLdWn2euKTYu26Zu2foHkSivCkiBEvvwYaawaHaE++zMKmly+XYP7kWrpkUiH0mFTYXHeSe
LKmjxNMeV+FtddL/rbnx/7TyLMcMIWe+s4feIFBoQXX1YzO6mx62209jD2bKoU73IKr25tktI67H
KSpYICOGjO0XQAm/jObduptiAaZMCHHqPylEIUgNPVS9proylBTz0Z65hponYezeOloPHMJXJsV0
IJA7rpenWFKnN90J94m09cT7w4o5//1NO3YTnt+qY6Ihf1OJVRLBWiwiplwJT4dZaBvCqB+Nu2zb
CzQkw1825Wm6x7YiHmGpv0rY5nrSlMlpJYlHDDmOt+SNbfJH/HUHbMzW6LjYe1AOhsdbGXeIUsCY
2I7yhIe4pmN3aGHRcrJJEEigHf/DQwWdIGPxvvpXNT/lt0eSYJwTW34Ed09JuVSgQAW2jc5OUkfp
aNYUSEU2oYTtAGVb/hTEbgXreh9eNOLrTaO+AL40hbQGW339r0xNndX1qblUizgxWbn6T7dmnfF6
AX6b9czaVzqvaUtNXIhiBsM7hFi1i3wYK8arKVpsWzRJAr7V4LUMpbfx758kkogJS3GeHwg4CSO+
wiX7lXHTzC0969GX591K9gWmqNusw7Kz3MGAKMW04nyQdDo8u8cFJpTmsPmyrJDZmLVFf1dmsQAz
zE0W0HDqqZ08mdBjaU/Xn0jjH48TDbRjcvstSRc6NcVwVsyCV8kYRCQ4gcmT/SGTC4YguXDtoZu7
9sZLIaa/OlLIK9PB3u1u7cJwPhpGaVWzxkQg/i/LB2LbsgtdAFzsuNlOAoVlGvIrT0dTomqeQZGT
z8Z5Egr4Nu8e8KAM0GSNIukQsoGmdKmQU6M+PEcxHLoa3MFvVKyIBTB8RdGZNbrlVt/l4awOh7s4
ABz2EmeRYeVfHm0052H6g3dl2NX16Bsi6Ti9dvkfRgVm6lYoVJe3IFf0Div3XtEZy5+OmBgJSHoJ
0L6VaLkAobUQg3tIcNj6L/Y3690Og0wf0XkXH1hhaAe12O9BQZUur5v6OqRi7Glql0HzV3nHWHMm
xbEX5t5NEdIsAF+aXmrVMHy7MlA4t6A0ZFhwkySYMdefpzdm0gG2Y43GkXS1DljKFesU7yrpj16o
eiFj5mdrxbrA0hHL75oF4Lco+If91HCNP6AlE2BmD7mWTI585bGoXSqS5p9FwjCLwgq492YpcqF1
r6brDL3JQgKUNPcoDYPGLTpxCm2GLM5v9JBM0LPZe6KvVrarRaQreDUTmPwuDMsY5BGf11mxqWDn
sD2hR9njJYg6cGjHt8+A9T663PAsxkjNvoHdjgIGy684liOZ4vx/aFEwhZyEjK5VQA3THdN/GqPp
KuobWhwyqGbRpPPUupW3JEsddVOsL/7asUHAhjskt6Ajfi6/GhPPyIUYvrsHAd9DDjLrCVaUFaYU
kXYeWFpHfifGsD76HTVqOR4SJ9FcuJ7o3fM/ctIsvlC6l4xLVuar7Dkf6zssy/PXACqc6PVDECh4
gja7xPq6Ujn6J/wRhUV2RtD/lCCtrPvaTCyzAZkUylU5pXgOSDTGJVMu6Tpm99mYG+T/sR4Vrp1F
7cseKWVjqBSfDhPdYpNF59NojXZOpdXUMjOtQyZ/XYmStH+lhU+tYjoc/hAj/kXEKxAUz+PnT2zM
SydQzA9Vl1xGAPjsSb3GnRWMDkcqFqszTrJcIiYB9fnV/NDcRenRfsUcATGKkyG9kMJGRAa5H/C6
p8sHUG4orGylq+PyuX74ZY+KESN4F5gkcs4yXq1bCsrHO++tnv2EvEmx7Oq0UyiF+CnWwVWRMJSz
MOq6FvV2c68akm0/v0qVZQM0rUFiM2VsDpu5BfbYNYe+j5sKpEq7K0/xfUKSvnlgqFbAL4Dx2nva
D1w4wqDIJrjAolpEnGskdJxkmfdjEC17Bglch9KWUMhFE3yHYfArUseVtwShxOn4ZbQpJi1OKgML
twY5YfLoIbEFG60cAkUsiq3VnXzrppsotwwXkhxcROwxezZAJDrWsYEEP4VXSFKC21oiTGqPw2Rk
HYlCNBbraZAo5Sl92jbc80iXbalxFD371kRAiCUvVV24zKknoSLhgCaQRX6fxd4fcbRzHVi4laT9
mSaQHXTBnXQ/7kf9hty4pI0oWB0vJKqnwKfLrWAjvI956ox11OKt8IQH54zQK+TS0U6yPe1+K5S9
vuv67/N8ez4qfHUB2CGN93E1Sf9EmeSfJObXe3GJ9vo4mlcyHG8q60gLcTxzvLfkI/zrsAIN1cEg
1SG5LUS9kBxRiDbLOU9JWLAO9x6l0fHSgWVQ1n2KalP7enf+M0ZFBzuJifklIoRmSMSHOwmGHaSZ
eKvMrfzo9IItvusK0U8y0CfH+M7j9SSNOTfFwrUIozNKGNgOK9laESumV0F8hZdhTUeMan2BWi8P
8h4HMEwO8Ugy8yNgV0VrrKUYRSf43hOmdrk+0jC7OSUwdpm65EadFrW3ufkOWX/bl0SVS33VcOEN
NJE7NDw0E8At9N6RRFAV2xXcVKyeZ0KlBkr6axNhudmFTemMMF7J27KSV+2LuEvPlnIt59DM/5TI
YjxvFFPFYJ5jnt/h4Zkh/60fVvDHRQ949iUsibjveTTKMN2qgoecflN0kYl08eIAH7VWAvJLZNEt
l2V6EQDuZ3GYhKHvGw6IBeHxRe7/NcXTVcCV/E2N2LobPEds2NhlQGa+0VKbYdcPpuURO5UPEzn/
U/5xzMRyeBbcXB9FVf3ZKveAcTEtvEsHlOmCOd4ta56NN5BD39jIYuvV7YRa01Gk6v9+ZMml/+7c
wWQ77hrWtjpGmxr4ma2jJi7dx83OOR/mjm6AIU+JNxi2q7Gg4CdoPh50GtQB+Ur3a+zsLuJd5vBZ
UXEJC8iLtsrMjoheCyoSZsp8sDjS7OuH6p80jgDMqh0YWPLnrVfFW0CPxzsc4bb7ugn2YaUl2+r3
21EHWrJhvjThkuxhmz/M5QivcdF0oyuVjo/NahDADZKPd7MQUEyuHgS6ZVVfoRy9eolZwHjFzNay
pcOjUNhhP5F5KgKRQRUBK+FgIpei6opbBD1a4dvzwnLFGyJmvULoTiIVc3k97dDBZSHUIJdPbpqU
3UjONNJYaSuIaDregSwfrzFWPiDwH6jDY719Ip1cBamqucbkcZUwawordbGZ5P003C5ieJBvd0h5
WOuKYmlVaDQl+UGr/2nfJAyoNl7IXg3GGP2aJjcl+WlukxlP4a+G/Rsa5jOaQA7Wa5GjpkHQT4X1
MNqTzysIPx2jVqsDU25Y4BylEA/FjK2i7W6EolParLTQVYoXmJJ6cbIIbYQdfofuAlonVEIPP98w
zWEDnFTpgwLOnNV8evzGm+aNA5XIN+043ZG2ZSHjrXV+n47hHJJFEgV4OxydVfWLD1aXrFnr7LDO
I28elUT5IYc9mha6n6+MpEGmsvM0qC25aDuxhQ0rqoZBv8hHkvHd0OQKWcEcarIu0kOegN7chX6T
L0Tj60j4khrdn+PTHXqA+BBemYQGclDhjgJf15M9sQOSmDz1nzT+ktrG8AMw8GwvLiR1ievKYtuT
Bgt8Ewx22vssCsMaQiGHqJjJmQ70A7XSqu2p2LN+pzSCt+HaxuAKHFn27vo7PxAIUlhHLbUlqfdY
QaCDDIH76ICydjhDhbeZha4dCfdJoFwZIaIpy0AYK5pLfUb5nS+yfkN/CzUGnsnh+gn0DilJVhRM
KlQDbPfav1BIXhkEyMfusB3ZTwlq4PIgsQzDMXv2YC71qLx/sHQPYewtOTMsryvOyMsEZI3mswK0
DX6ve8YUeJKI0zCySvznv5pZ6l1wOpH9pOlX3EEqKvadRyVPZQ6KSPcLac/Fg8ewVUfyuRN4tiuk
cDBRAyRP2vHdWRTurc8LI6R9KjsCEL/BAHndkawK9tbr8H0PWTvEGY0/uqnFhbFAFj/T9/GOs0S1
JJb0WzrrVldQhgelzQ0eUMjW2arDP0V27fC2DfHM2zREyd0pjBM23tf/ausIwxfa4Ry1tlU+Uw42
UsT7UnzQ/t0WMy169kl0jljP3OIjw28xnnWWGT/mkZH8MZqv3iD7RAf5ZXGolY/DUL91+/q0B04C
X29QFuc8Rkca5ExJN3EnKvdKqekaqBnbjZj+begicv1T2Owueh9Q5HEbiq8+MzEXCRGDFU89oOI6
0KFxhEfb9BNWhJUloHZY3xhRwKi2h2q+WpwJ4MEXLfPDEGfNqH1LkXsWQYksviYoRSIHtEhRwEe8
RS7KOSokoYRGHwtLFSQ50tMT1vyMZqVoL2wTd9QZZNaaLDLCLOzSANPek2vomOvBN3Wt0uumYWcB
kPHBYjV7eFeMAEhFSe3EH75wuOfV0xqwfGYRT4rEJ6guOyEHG73er8GTZVZv2ZC+Hgi7+vj78IU5
81WNJ/fT72PPjR6DtXEnmvKnSdyGbMZ+yx0xz4pDF3PpVvfwLTvRsrNH3Kbcb/LZ3rZ5Cqk5by3t
Xb1Dem30fLOUu7aOGg+3OnaN5CUzBqjPUEBElZELZpIq2zgfB1CoWMYShSbXbAS861G219JreSEf
jk1GVdQSeRR1pnunnAq9o5+NvEEx7pSXNeWM+uywDLShxYUhbWwutp9EMKMfVUTPZxixOwy8rrFp
Ah/Mcn4/IgL/Tk+XxsTTYKdMbfucdQ8DsZpayIxhVW8Pr3GVC6poSTqTJFuvZPTWb38lApaN7MWP
NMek2pwytI8NDYICOSFnq7H98zH8vYY52Xrj/VTtsEbnXdrWDG+a+PdHG1emykJwnWyYoLdhBRjA
yiN9aoTbNQRZ4RShmBX6HyORRMq8xB9xfdwzU1FOWu4QJQ4/kD6rNIzKGWr8RiUiKkhHwSz7tynZ
yTHNSFYKXFYJK4Vcc11OWBUn/O6o9/jfNJ66H9uBix5gGopMwj0i4qtAHqoUy5sNQXtaWat6GMtG
hq9Op/FTvS2kOol9poUj/dANNV0EkVO09UolQ/9C9NYbU79L/FxCk2EYXLoutwartI1pAfLy9WmC
KfbGpRf2MY0rIAuPtjhHqNCcIV1Ln1/8fxuZIgaH4scdpFdDu+Nx2vuYer0rat5+QsWU4QOGtPMI
v+f0oPdd7S6n5rIaatFt90MKHVpvrEejZZPLttB5ejrRK/CFkzcGxH5U7WALEYEp+DLIO9vmJ/8z
p4wvsyAcK693nlpvm30w4PwS+AHA7JDN7Lh2+V3psTXreLQp4pZjgP/t/Wp4N+jXCaxQixlfDoNz
lJQtnfE77O4jPDe3AF0HvU0RouGDTaeFi0w5E2gScOpJQrTquX5mIGIvawukld8GwvrcO+0FyfKT
9KN3FOYLzQhG8p9HdhqYd5Y5YiTGDec9K7A8/Nquv0bPXUaYrHDNnE9/PXhj8PASjg6bObQBLLsO
pC7lPEYdXERKX8YgjBuRlauAskAgmuDqFOvrhCZbnIEyJlWfmnQnMJ8oM/0wy2l/lAYdma/7bofP
5DSWu8V+eLH6GfNdqKxVM1Mg0OGnOVlszIXaOIJBY3EQSfHuRsIU2/b7LK04B93BTeYODyqzrUYL
N/D0yl1Dg38q3buXVLZxpFYCnee6VeX9q6y2FMi1+h1y4Y16QG4krMWvk/lQtlFnmKWQ0RmW0JcS
vmbLSxr4KVcxu6kifgva5v+CH274LoJoyENcO5TUClsLODuBmOH+AahXnHm+9y4bGAi2YzIzLeMQ
qm4Cr6TMhTB6KXDi0CaahtyKjwnDtUFyOUn7eb/jU61rwvGRQeWNubWY9R9++hoFnBywy1KntQ0Q
Dj9IuFrJaCE+spCOkpiXXgmPNOTuOGHwmtKqBYD8kfSFkJJFO9YfJWSUeNy0IETkSHQmojVwBYgX
ZagIvwV8K7ircFFmWL/F8GYPBbjLCkxaTJEAJYXs0lYNZiZvtVq+0uk7lcJHCXHr/KeyKIOP13kP
RkCMku+faaWF2mcpXUKscgR+eYbIV8Kh5M6BL0t17AL0FXPpUeOSPOvXSmxq3sTfKKDFnhg4qvDE
ny7IP7lCmAUY0Tm60t6vxemJWrdfZibob1JMgoDIRPQKPtjIPOm/k4tjLlF6hU71uj7vVopw/HB7
h/cIVPr4AE1M8UKO6/Fd/IhRfUEUjnXn59IwVNncdCz5kXA01WCwHMp6rV3vmFRout/O4IudosDr
jpQYhbfgb1X+dyVbFKX/JJo1M0rSpb8MF533Bz5Te+VpNl4uWp8bGUZYLzF5I2neu8MP0FtFEieZ
Vv5dJDpoO1M+oiSFPvDtBY0mujhodsi3s+txenaozjpyIw1K/B0owNZS1nT4RO7ZS9XBYC1b/4Vq
23+0Qq7kT1Zp3CuKwX6E0UcZPIhHZYvwYENZCfSRjpd3Da6WElX7xr1A7i16iDu5fsQwmhFS5wDa
+0tLGn8zctcjN/j9LMRehirKJmoc9mdPc0BtH2ZBvy4pIW7uaAqyjFG0mguLN2pl8tLVIQSNE8HY
AfHiVe80yvUPcabxuhc6wE6ELfYsEO/K3JTEned0EezyUZY6Wm1ILAkIqA0XbJ0ycc4VCr9vZD6K
QG18wbsNjcQQP62NXdNoqQJ9KN1R4TW7NulyuCkXhOJe6cyA1aCeXyZW9uau/7sX9iZZD2JtXxEr
MacohroZ6opCm4JzDiFIv6DLhO36sxcLdUDefi6lOJbKv53Ki2FgNpSkAHjDWd5E11FH0AoCUsZJ
Zer7iMW30BGviSTJsuOSuILXEVKDIxdEBhPa3ifWnAFrAHH2GdG2GY4V2tjoLJQ/lPzWm7EYAV7f
K9nszyr7dBcww0tTcLvkalhJLxA0PEsMZfOWYYOVxrbeuDep6EPx12S1zWh6Hl4id4gZ3TaSUixy
RU8Se5o3GANNGv3gfjvkLan2H76OIm0ZHfJkxcGHYSv/gjp3KZOfyV9OiHzo4H6Iof0susQJG4Ty
k/Jg2OBkO+g0H0cWLUw0gr5W6CRDUtPxbrc2F9g9PwvXC5f+Sq8u9kTchLiWBw3Mtj+LGj/X0XHX
6NpQLHmGErOq8T+8aJMNX/LAF+4VlR6RL6BHzT9lAQHZhm4/OCKJci2NVMt4C6NYu4Y6rHh57iSq
moDX7trqq/CxJBFNp4TwsLL3JnvgguR69tyKsOvgnLHZ4jsA1kSUJcCDqbwQ+Zw8wi7vkIrdKv7/
zZEVzuFOI4ilJvk4RZK/XOTpc3z76sJJBZnq+v1p/NWDsDLn+Jp630TgLMz7J7ZS+G/Bf4zrqZR0
K6hRtI/Jb+aYzyXa9yR8HUrH3k5kmk36xmUKQDNbZ3DX3uqC4pXWr759vz3wqR4ZZE63tD/uOxls
c3oVb/hnRxz5l7bqGr9CSO6v7Fv59X/YcUxfBZEXpMbB2uZxkVsvgOlpzEKrY7M9WohNqXWEmxzP
xaTaTGr30hFE5sg4kWtZO+fEiRbqGbtcjDBF2U3yZjm+IrfEJn//hDehFDnAZe5uO6UmTkOMTLIa
f32DHz08F8RdohO5Clx/7XnMGq5rBNaWeXxlTdnyWhfNJK1YyuzmQZirJKn75lkAgx8XM4bu5y+A
Y61NoD88aa+od5CwcnYH+11e8A++m1eN+cQkDKNARPqdz6v8yMtWDS2uppKSfuR0Dz86E7hwWpoH
rXdlHbLekjGGk7abUGw+4QKenAyKY/cyyrxbzFMstFYZ4d1zzWu/BkfXrseX1pA4D/IOAGfPpiQ0
so0I8MdOeZZKxYdyVtT6UCRka2+9WTug5t/F48eJf7sdGtj3jQvldGSdLDTelynhCI0pvy9JwsV0
BjEs0F9+bwhnFGwVzTavUcE67nwEvysXwq5JXwrz3QFhhkMaTnpbUfmBhipRh2MG4sXHiukBN7n0
GDpKa9T5IIG/OcAYxmeuFlktHBT5vuEydBbIb1TtSxbEVSj5TNs3f8sSQjvsaFcLXBCqkcKDlbXR
bpN3Y4m6TrJOKRM1bSzstfX2uA+Yg5Ec2S81bRRPGOQdb6TCItSh9A+2WKiikBReLYsiJxn8ZrZr
2aTf46Xf2b3SeURoI/Ak5g4Ebj8rT3QKzAHjMvWsEAiUEM27RWfuQ2pp4LfqOnd6BCfCG5jas0a9
oyx2Zxxbr/6/sOFO8k2lQ0iSCy4lQsfgMVQNNV4+z1j2rUAKY00DUHAHbqKcr4djv9qg//ovtJ8B
mDcvikcGUzt2ivxov6I8Q+ZVogJ2TM9Gt56fcPJlQjBBrsk/KyoH1OrsFBPIVoFWxYN5oR8E7PhT
9JTa9WAgdr6p9ThUdlCroQK0stao9YZawXb2XrTfPkQuaoubn0q2nlfhBZriaXWh5icXIJRxjmXU
6ydAQlc2qeXq2GEAGlmUQwl/5eIRDoECEzMiR5G5HpxZPO4ComkuhwzDGUPLBc5TV6PRHx8vxPvZ
bQjljyfgHLsI1nuyqBH0edbdNStDwtEz8X30YIuRwA1KdFIxYOhi1kR9FtYtHIioMWQABRlHvyI/
wMXMWMebcQzIYXLOP6NieqHp/ySYuSY7Qb+Xekpv969o6QnDcvHvMs+bz9pyPPXd1lX6eocw4vua
6ghkDsUeet9UsDzr3l9KoCLhDstTlWoH8eHoTjotdMTDLFz2y1jqls1EJzOXC4Vt0wl67sCoWAbW
48A8KpC0Kd+xOdQYPzwHjsBZprppmRXeMDv3YPk3grqG/tfNgNsd6Xbgfv47hfQS6vr0T8CzPB7v
7oxHiTN6tTggOKdtDKAXvAdEjaM8q2UeHwLGgPEbQpVITzk2hOb0vVA+QuE5Xo72sAUvZii24UbK
a2w40QV23al0sm8aDmQgG+hJ7Vp/WJc4cExHloiN+cCfR6kcnjWoapObY4lGqQP1RFIs6IRdRjJo
lOEeZuYw2SQ8bI/wBIf2QFamerHM+X9ivqG5Ba4oNQScBOeBp9W5wYaSrxjY/SDDeDWUMEVAX967
h4A/mbRPJFes9ZalManppoMm1wrjoOVAHCCDRzVuy/XFDHcsYtLsTwVpxV0s/NYYS2S60DeuQXiR
XSbjQ0UDZyXzRhUJ/6umU9fAcfszJgmk+pqM0x9D1Y+x7LybYBIqfHWxZkzHe2TlOj4LOE9NrZkA
kEt5eEAlf6IHg16xDUPtHeKINi7DIjVpZmIreeC06Xi17RSw7Ea7PVrtWYKrs/c4G5cafdy4HYK1
qWWixtYMgzNVgD0f2iq3xXNJAsOKjQfNX3sI/RdWxTNgKRBM6WW1u4lv/XS0t6riR0HdWLnun9eM
le8zLx/f/3yQjHW8pgQRfkD0JQmP4FpGACPZqQNAoSSr4Rhb9HKYpXN0TO8nBK0i4VOR9104wPR4
JV27H2zjGqnM0/Z159KYcc96kKB74dyTklAfIbNu/gvLTh+AD570ikrFBr1OWyPDepWi9pYNoilc
4KPDHMiQmEWeHGvFjIwf65EtZ3wxgRMAzNiOODCd0Dczu52mRPBk+AjSrBEH58HQXPmqw7SFuNNa
DVJgSljvpVIgh0ODQiO/IjCO3WIFxP7uxUXUjyoEfXYRaGtZBhRFJU1K0kaemBA3coxf8BYd3F2O
JvLUGzB/wfIy+irI+rRAXtZGnfCcVNNGgD5zhLisU30iclHSRjbWrWusKufH4QpSbjK62LDRNUOP
3H5zUk5BCleHZOU1xSnZb52Xs8RBXSulsxeLaUIUcBl6fcHhkaVDKJRalaCTkx/qORIir+HKz3N7
ILEQ7befmeUdSq1QafBwIHWCHeqIXD+NUVUzrkSEXTdOyPfxeH07DbsZ6i7Yfgo0g3cXj2hz9Jnq
aeupLC71IWxgnxEqyGX4+Cu1DD3gK453Rp/2YBu9Jd6zzdD9zMd12PhnEK2/qRjOY9XjOa1NyngN
EocYT42azZVHj7PdHp+iRCYGg0uo73NTdOf0YzUPf4Q98B6M7Q1JeLHDN/kI88g5F+CrS4HD4VYT
Qe5Vun3FfRL0oEfWuxo+PiZcgzOFVbW1OBxxrKMJwQHxPLDCwx+vR8Hp4vBbUv7Xo3MX+fpTYXBL
nGsf1ToQUfOmdLttAnhMLk3FezdTIzoN8cJHCJKhZlwqg8HjIjPHl2eOT8f/wUqY8wK2wz4DZ7Yg
ADfEn/NK3FKuEjhDYfTrntzlVsctBOqAuqmH7MH8qdx4gvEbu7NktHjzyVCNOMYOJJE890M/tfEJ
UBpn8J5fHaxUT8gckmGGBmJOaMAijeizC2ewux5F3Ec1uwSwMJzpOkEgBWW4DBcuz6LupAor/stl
sIyKo+rqsqQE8/fwDSmp7Ie3PnX+IuWd51U/KGkwtMQsrFBOMfn74HHUMlyWlyYWD1ww/0n9r9TV
AumKkI0s+5RF/nsistpQuIV2AcIYzyWqThch3iBlIDY7UBbxhj4iuFZHqBNwWWbXSBFOiTbK2NW0
oN8CqvMfoNlqOfyv1cPGpiGM0aJglfzo5hVcMzcjEQ0YvcFRwI9yRhG5ZbRsfty6pmIU0LrNBMEF
D6omqvSMFhkl/G2VYw2AkxjwbIn8/f804QUtODazF0dNBOQfnqR4F6kkyzKuemv2t3FyMAGyHCE3
6jyWvSZQBZfVMT5UGseEVzdWp6vbPH28A1sWaf2EUtd42KIL+6xLUHl4jZeE7Jj2vqEikMuuO2/x
uK5IEdcyDbGwJRyKhBvKfLPd+FJh+4ObYG16SfWHB3iFK2P9BHruIXjrhQ7VBbmUK9BR6lX7XEID
0ZombIK/scRGrxH+zL5UVpXjd8r70oiH52n1ZuPqeR/EmUpyAEKiRX4aEVjafTY/sELTGaYaBv9J
bkQs9ri92NHLd/+59Ml6Ab14f6ppRxuDpiPpxQkNG+Lrg6LsvJf3RBtO+JighqFSo0pfvGGUi2Rr
lP3FzNEDVPTZ46UEpLNIK6y5MgcWXMrnUmSONc8GyR8o4F0ikf9Pmzvu97NezleaX/kmjvLGUDT5
LxXucgiw7dvIif64r9WIGaYrxuAwNRS6SL3CEBLCFXwIWDqh5D4OCK0mMgtqcezOtNjux9jXvS02
5RcO07iuQ5ra7ir8uEBqhG+WPBu9WWC71vyyT9bRd3+BkaYkLbfj3WFYspxpwZiGryFPJMY834ge
UGPUdeJrc3WshQjQh9laeAcg013cN9/wnv7uSEk52t2sRtnRigmj8zDkrBFSiWZ6R+2s12XLm7FT
HFaF/Ew4AGa9CaDQAkpmFsJxfQnqkyjRE2jPR5vV5FYJaogSMnyry/uCRAPbny2hO6E9O4fRnHVn
FpsH9U5uINgTO5xpACbfeBTp0ig3Wl2p/DgA710IWkj27/haed6ZRaAzC7qZbtCNLDvEPcMQM+Dv
9Q9rlBip9Sb6VHTFHph6JrDf3pxC+m5NvFRqD1saa3C0Q2cwKGK76xlP+O+DX/sM1LQu8la2QB5W
fwfpvUG5SyIu7DNJjiuiR4do/FjIdkYYLBdk6tXtunqghch2181KoklLqaBMs9ZA+s5X1JD4QoO8
9tvqHBCfRN6XkEw7q7Lk9Coo7h/t9uSSa4+n832pXjtO3+oBRsaB1/ApYQV3pnmMZB2538za58Ej
pFk5q4+JtMCuxc/YCZ8PB1K5kIfQKaninKP2hv3Y7E3TtUuOPxt5RtSjOZcuSpCutXSZ139Jtx8B
HalsE7sSEK65B7Oo72raTT/NmTT6beMk1rxAFx/ArFU6MyyYvq8oT5cfr1oDvom0uYRt9K//IYdh
wWvcYn3MhRoAZmK7F7ANvZUiOkWIiXrQvcyG4oFIWbh0fiDseUestDxpDS2xI7MZBEFq5MsR0H/a
XyVqrz6cwMMU6HzizO69E4oikVf3tvqp40MpxSZonDrJNOuqZ8JrJX306E9N8F1izO3Zx/foyhba
HMF61cGTfQu8xeLEazGuYRSl6FlRyT6+Pythk7kskZk2ZxJmawokAhvvVrw1iR0OllL1kVUnSQ1a
ArYfVE48XIsa1lh5b0vuZplmG0+J1U7cY1fvxCD3spZYvBezHJxLvL1SmL9NCgm+sxUle1Hnrpj7
j5WX7lW0KEp0xIRh2z7sI6tMNtLoJvCvECeeIZYyoXD0/DSI5tQfuP2H9oEbNbd+4S4hJdDTXxD/
pw91Er+ytcBKdYTgefy3w9gH3s94DqXLaBzcFWbFZkNIe4oNRjgHqIFv640AXRY4d16EsfSMbk53
fq9ulG0yHdFWN0DjoZMdsrm5yVf0Ao/5I04hZjyvVT8j3dtMUcoJEwZxXK32Mu890+Ns6M8nIfFO
+QQPZG5DPyZ+cMCvaDTfRO9qA1YdRr8cdLYTuh7fs13P7lmztgBs+LTRKBoLjfn+GhV+NID+3TrT
wZVxoJJ4nztHUneqxTWsNAwbCUQGlZ2TCtadlg9WgU6U7jho9LaZVhSdDcvpwofDxQyJGiVkBzQJ
EiRxgn8VevikBlMM3NhE8/deI3avFUPln09T5lLJaS17IwsfLF3J4YQj0SEsz+IUsUbYrvgfzT4f
s3RQiVGSPMKUcBqyOTQPyq+K4Kp4fuYozPQMLK470BIQdMfqDURNErU3EQxbowtoJ6CbBJYCs2Ig
g7706w4NuputqEec+dJ4rKpqgD92V3iSSu0hEW+NoYK439QF56l52lMYQGXTK5B/xcYbT+Uzn3wW
p7ReNgM04VC2P1cTGy3tgxV+cM2skcvETYv1EdOiuMWggnvMBtR0ovb+NOaSsTGd2U0iKyLRAKPz
pf2QPfRoD0mxO42s4fUDh9NbEcuWLmZX3d/z/yJLNumaoRuyYAjyZsAhh518hdFIQdxVWx/p4ASg
ww87WNuL47itACSRwV+TmG5Xe6RmsCp2IueUM489k80WroKePNF9u1plnyWtryj2hN4juC6il+Wi
vihHbFJkTJLorpZmTZKHqplIzcZa0NDFzOuNfesJYBJPOiSYb3o+DEXKoDyjkYK/+66PaeouqEo5
+mR8RNyIltFQ2Nnj1sJkCdUZOQcGKQNIOAlGPsed9BFO6eaVNMyQuTblAJMi9m0ziR7OnLeeebkr
uwhEG1of5jScpYgt3cxtN5IxWZ+M1oIc0HXsdFwvWLdjPdBmtPI3reveddvALELTeaL/BjWg8FSQ
BaiOU0ISs28m67wgrMAYl7yenVCLDeAMlz8D/HJE159ZkJat25+SRhwgSpdHwuaEiCaVYUfAe4uZ
qEIskec+3vhV3Cgur4Re4iwKOGq2bXq/gKaPxw7LTDNGTyrNM0JVfzaXHvhsJKhZJkGS4qyLeGxS
5p7owhN5nDQ90mVYK0KHPIC6ZOFF5AWwA39MhKf/RjN/AtA99VfGtHwzpKcca1JEfRLUZSUt5Nfl
Hc9UGEC1ZjGXcWmR8QwwF94b6WXPB6pfit2/dEj2J8rG5Qm041qBh+voQVYMhmp8lDgFyf5ahWIm
vum/4zpfhvmeWS0Vx5k5m0rWnLGKKUjSN5zwPmzixSy13naaYb8JksqZzGdk4Z/9BWv+zextTp38
GNdL/ciVxp7W+nqrsUaBkLaIJ2iSgHW3C+G8Ype+c1muHXSaF9CDKapyv9LTPU672oeV78yAxuhC
1fHTtvQzBXMv1+1JRPgiRn+uTGIiWnAa65XZ+UMRA72BUjW492oPyXNKNCLUc4YXrW6z70QkAzko
e46+AUf/2OvY7pncNq9eFRYOJfI2MotnSFZL2z5vbjYfZuh3RMkEtUUZCJANqy5FbAImYejX5oBR
HFqXetBH8c1eiMHRiiQmiEldtdCmjC7hAPsIcym2P6x3m7qZG+P1djynJDjfNLF/2JOjDQbBLF1G
JL3z4ijCfbCn+/ZW/xYy4qQRP1l8GtvTlZoMn/1WVlRfVPFxJvWL0vg+VsloUmdDJbhuthm2xoaa
bFb5uUgMiQRniQ16aD/T/l+8eA5vqFJ2C56cAqvAtLtDisZvMJ/Wik+Ng92itXer0kSJKwX7iuZ2
hvwvHRMPl0kUlT25ThaS5temoDeykFWsJNOQ698qExqbwI/+etLOq/FgBS7hp5rbZhg1lgPl8Obx
nT8WrlGpMGMUAH1//shzBnnECtjwPA6CHlqY4hZ5WfJOunD4ghR2QrIvurCWXqJTyZEYhWBpBglc
1Tf7Zv1QG1lXM28I1tKkpyeEKJqW+nZlWxvWkZh2MLZ5YgJ27BmJf6zIjQUGwTEQ9ivva/OCF7Uy
8bOwUqDt7ljR+9UOWCTm6lUlaotztYCADvwq27L9Qb4r0MjY+akgRjnMbFItBJbb4N91AIwIAuxc
rml+1lo6LSTKZcGKxs6EHD2CwjKgXlSEh1nRQUJqRcc7fV2OYxNrDhCZG7zV2i4dgVJSL9eTjbRN
e4dpMmvgwhmHtXdy5YU8mTWPiIdfGPGsd6zsWPGlorHVT96qFiYRbZdxXcW1lTtWWb0/iOnyPW3z
UZFTckSElEoIIxxZxCEyzAa9xTJ8EfHCfxPIuzZUk3XLaE6PiNXEf1HGIdiGW6plYhDArY7hf9Li
2ubNzstpHQb6zdgP4El9qCy8xM7+zmx3+x/dahC8+JmDqk+NrN5xDa4pqSXhtguUDeo2bYb9Ofb5
yikMdkep3iSKj4zwoJt8ueYv3tXL+NjBrcR7fpKJjG3B92gvrtyl1KI89oSYhxVeCKOWD8DQN5fL
sWcJwgkjD2nhoGnhh73MrvPtb0ogAoxS81UspiPSTjhUJODU6lOCcF0OAUiS6XD+8Meb4870EM0Y
P3ZQtnFVt03jlCq6PPT5a/OAq7QQiPyjSBrjXV4It3Hq8oKjI1a4raeck0kM2fbFGirFQBi+2LY1
HF2HX62YhIh2PvHmxJwai1quJWO09QkG+uFYUI6yTIIlw7TkvaEAhjw1vNnKfwFWsL6EVLoQZtUB
iXwf3K/9iZK4lkTsbGOC3wbUfJdvzIkFeaCskCGymivMXae23Wr6TCPuqb7yk9LH006BeJxWlICa
qlVyD6n28Xqe5wiKavTZgI2ApTC4AF98TS5J989RkzFE7or+oGly2aTBHl65h7E98QL6lFhMmtR/
gnHtnXqqNN6uPY6xVznl7nEqt5MkwAaaMG3Sm+bdJiyGGX/WrjkMZ9dFwfdqi2z74G5n/ErCvq3/
bHC0gmVEC0i46t8GReFZ6fqmY0bLwYdlk6EKWs9g7Ow0soA5Cs9Y1cupWtTsSUklEhcK/aW7JbR+
CpWudftEtfq29Rf6XJYvRcmyNOQIbI0xKnPp1D+Tpy2e7X4nFnu7uBF28W4FXdYHXkRQ7E1ejoyK
v/u3uKXEnBD15pUUHhOj0ilKT1bosc3OXuZ4Pi/qmgs0OetRkMK2XWEf+u7Ghk79rwMFujujSaRJ
1UhBb2k9mSzgOGbPS4ruFYsDAJezg85Ct8XW8oT+IsnC1htpIRKmu0Opp7yxt54hYMzExFRN3tqt
/FT7R6975lgNB5F0NFBpU5h0y3X82YCwNBoLPP1P3X/afRKCq+pkMgAkYQ9Ggn32ppuGsDO+8oVS
PlBqrQjzPiqvaGpn2/u4Snrr2ZbUSxZh3L2rqk/fBEEBUpTT9uzHBfZpcA8Caj6wq1XtKwT+3IHx
rXE3e1wONd/+4lqL1t86b4weYX/8a1ymTlow1YWtmzMEvSxPV6xDWMk7V9TSs6FyVBvCfvMESE2o
VI1oavGIBMf9LFMRQWpwOy2kb9/VJ9xDaB3KdInW//qqX25rNoWghKvB/W9llI3WriOB3Gig6cpK
XpZerUiCyx9SzO9mGyzvIDhJ7D4xj7WBL50ecuqQbP5LzHjNCJvF9Yoj1Tpr3abqN32p8YXZQBaZ
19qFGOuJqfFdOvI4NWYmT8Vr9spFIhxwmokGq8/oXyxqBcyUWxe7mD0tE8rp0EHrncQZqbqKXeV8
H7yhYYA6lrhvb1pomkt7nNpSQvwUILHHfKY42PdtgT/1Erdy3NctZ0rr2AZicT7765r/LQTUYFU5
6Ui1x+SlahUb2qBfOfPvuReGJJokLz+j7b0Ti4Qfzci5Zl/3pf2gPlLvs4rZ/ewuy3ZpsoRYQ/Ae
yMZMTFP0CIutLE8rCBSNmb2WVFjhjK4L+2Wr/uOyIai0SJT5VQgA0Qvzk1sdVlMzV9qSDXFztlAf
57nCavKl+7fxz410A2HodK+YzrUp9TxDYL7y/JJ/V3cq+ABR/VySnnpHVne0fHlWSaL/P3ZT6JhM
cW9O2VQMRB8ZiKtysd915n55+QjY1TS0yaLi/hYmuc6uwAFSLLz8h0QLz4bzybUWFaQwKouFUl2B
Od/LVlmxlVpkrAKxF6cFr0VC3DaEQjeiBOsyLnHHfh9KjqEBbLDUuKa98UfnIvHAbLJ0b+RM01UU
7A+RKBWh79JYQh5DJTNs+F/A84umVT2tfayOFEadyhbv12XN22C4cXxMNXeAZCTJpCXcxN3c0Tj0
KxrtTXyS3rzLHURITCRXXzZ0sKfAw2KU2YhhFyxioPz/9BbkYfdrvIwvvpQKIa9Ervv3PxLdhly9
/zSdNhO75B+qUW9DZfBI9LPhdZDzat8rIWLKPL9ctH9VPyqy9Dx6r5sNmEi+Feyd6Vz+3EekIttp
0cpGjEa4JBBTOhkeHXQlDvw0eNEWaqfRYEy+tyFJhmXifrTYVE8H85FFhfmrQ6oTJS2GzglTFu1g
gMZOXzGgGCjwTROouSM068Vb63Upgn+nZ5cbBLZsqlv0rm+9Bz9c87WvDUDdNLlP4NcYYTRl53A+
qt703W6cJ0MkgCUsFJ8LNAuL8+wxAbzsCed89rMIPkw67BoMV+oVmkKekCYso3rJ+t9D6st7TuVH
/0n1Ya/uYVKEsRxZ2piIeydF+3iZ52h8vbkd13/a3BEFI9cDSG0vTFlvSSAoFj2mih/w75W/HqRJ
pS78Q+4uQPyZZ6fGi0692PX/50KwR2E/rL/ljknDtT6h0rl5PD9wRR7j4g+TAq5Rtq2k4zE7Jf/A
SaP8u0oRZE4w8epokhtkdX157ei99uGMqy9sNOn3S62e3ZA3tnL2X5eDyakTxRs8CGOWkyQ773r/
dfr9uBwWPpSw/2PAGLCz8Ta9rWfQUUDsw1z/7xkaJlJwoaFMeqqTCkd4HeYLj2wbQRvLYG5HCOli
RROXgzL1EjAfgN6iBpfv1U/XTPZO/dil0T4fn+Qatwu3O8+DeBV8hK4ne2mKotHKT/k3TQMwE6E1
4eZad7tFxO2zrEfbym0a7/PSr/hI0Gd0mIKDxi9wCEYWF0Y1NCz5XcLzI82AhzBo3APe2+MfpPdT
WEYC/mhc0jrDM8A4++snkDQDfLNCfl2N7jiB/NIy0mETYyHweJqkbqmduFaRxoIBXk6mwQLMA0wd
87rbnBIzr9LurLUtR6hLtlwiaG7frNG0n0bELhEy2inmx0VFUcMVuYrhzmT2b41ivfzt72fumK6n
sMdR36DVACRZGjiS+EMSoSQJQj/qbTbhUdwCYj/2XKbuE7gkebcrJEOBuMm4eU49g6CROT859iV0
jzJcHXVzpPAV6YsbIWbNqsRR4wUonMv0AUyoxqOm6IV6IS7WjeMydIQLJKFh2K8xwXsC7BzNfdau
mzeZwM/QM7xoBVJLFvbikMl8g79xl7Io3xK01/tlWYdklRpT1itxcXvUKrwYz7Ce/J19EemUroeo
n6wsu2NvSGW0bObPdysBfCgMWc2g/f+H03VovzmA2oz4nWUgDzZC/VFBnB4oCNIiOYmG96wOGLdB
WjjQ4S1axJLiUgTJjgwngeL2qOzPkwwecK10sNp8rQHj1C9hsoMUQe5QHitzFleFnWvONjQ8X0C8
BwsWR/wk8I+JcDNv/+3Om4J7rKsZzC3tvOtYjkXrsiaV4RLJ5Yk7NxU30XPKmvGKbaQj52QT5ucy
RaRdeO43KXf6keOd0veYdsF2UknDxMZzD7dbjGEUOPPfAVz2xuiCxqrgrEqU8Jm88NSomwpwDZOD
MtOQA5EP+/Na5H6qYoZvUo7TC2Poc66WM0H4hRElQ/txJk5mGZai25uf5D8y8Mor1J6tcsZfBOaP
eTCbgZGwuTjP1XQXF3R2WmpfWMO68G/Dso5mtViWg//FhK2ic1QuDP0227TEc8fy9TuaamGS+3+t
rXZBrC2ZsIkr04KHKHctrlk/UycaOkTJs6LeAMaYeD+Elmini78zQSy7arXJVwT58qzQlT4CyPAR
rf5s8fUQdifTNrr4WcD8Gz6OHg/Dtca+0mal8+do5VZRB8JlGA3EEq+R44/mfDtp0i8NMzU5+plw
K2rqwP/2xGNY1J/dG2aeNcW+8ODrYsxrRrGpWQ3/JFycwEVl4k815BtEeaBLjVbhQ5E2iHGIFQYv
1qHjqUl/Yape3lHuogWE+vV3b5F9cc7rjhPoZOtnvIkMiaINPOS7muMeG2ZytP/3uRM6rELsXaEW
Smq1wbk/N3gpUeMCCHX9LlVul5tZR+SlUi/DasnSFy/PDPf1ZAw+4Kneg1EeKe762/hr0a6fPJai
biq1KvPrKXyVi0c8HDiF1h+6ykYNkq5VGU1MW1lCEWh2j4VdyjeZfGvsHOzPiKG9seMu8q4aLiP/
tlO4Aj+HvrY1YAU/8D7BvhmkljxPX0ORUqvy1Z5oggQamAd0v9sfRljYT/r/a+PtCqHiQg2S1CC5
aLuZMKD7oR5A1Jhe8SSfBji478v22QO9aOPMpCsjkn3tdjTE2nH5hsJ6jvE3w8otP04jfh+R9AhK
/GUTX1K9UEkfVimx8jSIbeDzKk7TiTwRKG8Cl+tbJ9X+GRDLngp4JeXXRDSgX0JhYKBnBXn5rBot
JeczTTdP5QKMCHHF5MPdHfjABb8VTsETR63a5QtqQNW4m/DdOxSdy0oWJDGnLA1maxLP1sXp3oy3
76s7Rwp7zzLeN+ouyOGaB9RIjxTDThNf1WSEexp6Rf/L3T7Bdf77uS30rhYgKUdg07+bPXHcbs/q
PcvCm9zrmcLv/khTMpdyXxyaBZ5w0bSW0Oi7cElXHYyci5dHKFvxwJJ6GbS1xlVhWcyYgSmuCK1Z
8y2pddkGHo5s2bI3V3zcGJyjj95U39WI6YOkNgQHhIEwdK16Mza4BNU3/bcL0w7BPKGf2Sqf0BBQ
QUpEf1a6pWxpX/5btE66HqU12WbVCc6/pqAYPrJhTSJYRpZ9+beJrQ633Xnryaq1Ptm3L3Hyt+LG
Hr74PIcEXPvv4SdmcUuVLmHlSViX3+uh+Z/ErY0YUx1s3B+7sMadLQHq+U1EH7bMjTvy1R3X5HGC
rOkObu8qNpJd7uPSkBfy3dSVznlUIvKF94dDpHt9BjsFEokPKCwHZOLpUDQT2D54rIEhC+IHokoo
eW7fjhMOUi9TtHOF+rDkEC9rnyzJNCMM4L+6h3ziAGvy3kwUFJoRV7Q8AJ9oitgormKqGuqsZ/vC
ZnUFpkI4lHh6sj+7qhGuHgUjz6y4FlnSerWyRpOWhAApSYWMiMtYMjeeztKRPIXbjZuV1U3xqCb1
fWDhYxc+4j31lCa5s6wT69Z0ry58iw9/y10DXi80FRBkPgvdZbKCOvHdqx9aWYZW4USYlKzPHtzq
iP185MIQOgY3Ij2ERsKYfOQ3uBv2dPFRL+3Lu1fKyHHGl5H1vONnqPzkpN1p42Y5Qm+fswpsnwBX
O26icx6T4sRd5BDSPRqVc/3JCjJwQskDjiQ+wQ+hLLor/sYCC5JyTjQ5Zs0Bvl63gftFZpv3Lsbw
QJwMb0wlrWfLAy5OyrZZHJOvEegCt0qfDOwOEZU4wpArNB54N6U313M+q5BQ0e4iPRJ2qkqT6ppQ
GX020sqf2+blX375z1QuanqTpCzqbIb33CSQTpWTwOR3CENDWkcdsIgcke3oDgjcKXOpjis+VDTD
rqL8MHRIFZPL+WLvnE0EtqmPAUnuiMuLKzSzgXzSXBBHsC4F/CfvDLW7kv/mYu9UEIKARQk599wa
iPqq15T64fxWMKPzSpGMV0NsvvOYTXKeH+FHE0OIvA0ldOqSgleB2ktsx8QjqvJTveFYl+wKbZYl
XXqJdBAMJREkdtsHYApWTTgFljwhzWHWclqtTYL66kXe4+H7P6uWBMFq7a+Ua7IkzVg7T6OQ5Fzo
Dl46mifySr53pLdXi5TGiQl72PUtLF6K7qyxNbsZeY6IamTXQX9/ZVDphoINLspEU/XfCqMdgNSX
PUYpDpWSaTV7HaG4wzSqMUts8hAv5M9z6lHt7bygCgcTlP8NqX4fTvo7Q2AYoMghDiEulZgq29T7
45hP1tZZ/la/5Zs/95EKnKwdX+bhFOqua/AdRrwZKgY7rLBeRE6DvY3jS78VdUsJGBmFvmCQ6o8j
2v5laaKSmx7w6YlFHMmTxRqrpvy/NnDZKQudcCw3c0Rh9qn8lddoboGDDHcWooct9+caBt0D5jja
G/4QUtXT+QmKyBuctXyaIKoMWp4aSp313l1O4btpGPnTpFyKkYdSy+6yv8tccHJi9wR9A5cgnL3l
ZnGyjHFL6q1cmxkNZxx43M4sxJ04q2IH2JjUKf4RflcI/xHEUa/T5eUfCyIHFFskbqe2Bu5v6PA7
Agw+RDjhLEZ49CHcw7tnVyFn0Q2hzGw/3mzlnwqCI0ptyq8WyF9Cw/CrB+bKhANj0go6we0YnV2t
fIkExuhIOjGXqefN2yBdTNnjhBczLr9+XA79Cx251iHkftUrCcZX+514Eoy+UFpw/E+yTxKk+sej
2j6Bbys8bKn1+tkelhxD/1qmvZzoaDLzQLTeL2aV2QBtA45QSFEx7JnU8S4kZgC5CE4AjAOYi7ic
cvqx5mHroDITjCVC8C+LkngAC7WKfhIK7djRMh0iU95NIl5Zqdg+7rb4mdqSMpck7t4XO9FBBSOc
zNw0RBEoLHRY37d3rzddSKgxNZqMsi8CIfl9EhkO14Rm34KSHqhAGem1w+mZNpL0d2WPDil6W5Rd
SpPvQeznhoq2hu61pXtC9d4J7I2zJn/2Y6RVbrkGje/hOn8MkVq14PrX+61hEf6U2xjYGyHAkP6E
vxpQG3mz07OHIXBhXWAGVixUlhbBkdnwsLORbd0M/SvQm45B/SrRDRiogQw5SwyhDRVM21bFdejq
MMFHQHFJW5Yc7WRly65TzgbwVAwiTnyUVigOK4DqwL/Idtp1BlUA0b16UXXYtCcEBasYYEqmoFzv
CxNKhQzF/Z090Cmc8eirSPgBmIJYHZCLHyTYtQhW2ad+SErucjMEVOYDyMjETFU4LJxLOqRaZkd3
evJ1n8I3xNUVjeShH5ZNIYPWNWj5tALVuFaesHFHFy8bLwkx79LRyHBZ9JdKDfGt05lJiJb5DXl/
exWex1OhMtQzT9dOM4KOjp4JxZAObQlKcECgVm5lwUq51rXBWznpo3Ewk1Hwns7X10RHBuJIkc94
mcjMKW3HmX0ef58oBbsiMsCptEdGtV5pf+PYHKPUkptFPt0VJKHbwLi59JISQv0WjTUfxTRfz8v/
CuqS8stjzkk17JGUZ9fzBbiCo51q7F5vA1bm2Kugo8NIMiLdzO+ItWqijTMU1yECDM0Sr/VtMFW1
DQMIcWtuMSgcteweNEJf/4fWrLKLkL1ld7rma6Hx5ZnXkYoBait2dbOBp7m/q09RAv0oO81zgnOh
KWSq/sPRTYPk23Yjsco2JUfq0fXWZBIzZWeDJMlNFxwzm8uc9q3tmozUmZrjvHezbcNJFgvrDaUN
YziefXmqChLVmFhUwJzQco4QITrv4BiaD1hMIxc5CCed5oLAO8tp5Q2An9G14mnvP1idmuBUQ4nh
+ivvRO5EQNCom6B+s87b1CNZgZtHZBBTHHm1CS//tNymvoNyzUqtRinb42UtnflRBPvBKrU1YfWx
/pBt+hdMe1juZ4ErJ75U2An3H1L1nzlYJj2M03ZmcAk6ztfp3kwsdcxkkhFYXP4JdMeQjWPW8x3J
nL/9lX4eTXTZRhMEECqnSu1LvAGOKP09FCAWk4bZVwF7mcdwU9fU77zRaStqlpC3+c8kPArHUom5
EI125P3PYMWsE7lABzVi1bP/6+1bVy3xoBiiZxy1USi5/7WdJuq+Q9GfS6HO502Bssr+GFytIVVm
5QTnk+7KAr/Zr1+4IDxWHuUBX0yiLAkJw+O8d8xdYtewgF9aWfIUlg88Q6sjc6W6hZO+yUebg+6Y
7CbbEoFOKn7qTanmQKc0bx90mAXxh0rhkaCwJnUZqPbMihHpeyQF8CK9jyy2RKFHh33E2AaTJbyp
RnQf5OAPw6I/jFyMp1RPb5ahJ96WI7sEWNaargf6jPnDruSuFBYNbwEY4RrXn+KLJy2rIsO3n9Jt
CwR5VtmSiwKeIAvjY929wSZmH+1i5CIuq4RGgPdLPxDQDQvupqGQsqlpMcUaKIfBwss0BPHyP8ab
9/aR1iTRWvW5kbXFe5OamkYE9qSQQ4LQ/fvJok0seiCXohNIjgcn5Ko06PVljVZtSwu9hWnnmwY9
XzV8ERZOTnvmLngVgWnEy1PRtZQmzD1xB1S8+itPZChWjheZ/Q6xHZFvKY8GVIWWb4i8FE3RNRGE
iZfHxWL1IZ5r5tIMEkH9AtKDjwZ3zVA/Z0kQ4pivB3PsdX5WsXJ3qMp1iTjZVwigDq/CMpp+Wjdz
80f7Nl9ipYDPwa3tO40MEw2T9K3jNZsMjl3HbKy/GrAr5jtg+X7ijWUB3XZ19H8kyukYMnHSdpSJ
MqZkJFKHE8pfM4IjRB6d3BgtBkPugD7OjnfiO+s8iu5cfIHJJDmkAkRNnEEQ+eZEERyHTUIGlVHL
Uo63zMiQr95ZONyvmOH98i4EI2zwIdHJLClFVkVoab4CCrC/T//p+BtdzrDHYufKN3ds0uT4yliV
HOaX8cn6IdNH4CiS1ecjHaSY6B2kZfIP+IwOI/BYD+LnDdRRTFLNWZ8BppSL8cxYv5l3ncNs2uIM
AVBz0HWTYgwxtFJgrMUFnBpPVXSfyWNQn8xeqdxhAYQK34LcROpGxAwC3v6Y3pJJciCJ+kYn5nwC
bbr6kVV1pGbPIfDHQaHHrGODs3sRlGFiYOnRjxhed564WDkyxz4p9FULBP/Zr2okV0XEdoRnwoP8
xImgMOjLd33WtAbuU1Ey8ljwJ+n23/26/992NgTKuoNCou5OPIkQIqDk0TT/ZxjoCi3xgzANxDq6
6u740X+bK8NwpBOk/h8VWnEvn+nwUI47EN0p/fGtaoqTo+fJXEX5VKrzJ+eF+Ho1uH5UmOYwMMZp
2h/q775IGjgDdFmC9555FIsXBNHxqqnGKuFobSZvhYHPDUxqXIGuloarK/VSzc0b0xIh6F+KIPH6
Aq4jAIkhRNB3V13y+PGrSuZMaO7da2Q5G12YO5y88+BxM0kkF5PbQ9YWp2bIs9m/dcpgC/OvJiqY
QCplL7ZPEzzqQ8oP40asu2D4oJTOkwx19A7L9tAt+uxp4QqpBqSJ1VSfNE9O+SDOz9sU0OpiKlYk
7HYEdsHz452KdEghiodGH7d4PHzK89hvf7X+rDva89SV1rG2Mvh0X54aTNNDCS+EPkG4tgxlSZKN
q3eUN51ebxADU7fIEY5Tg853kjXAVCKFhzdwBZ/10qyQewL1FKqTsYc/EPI+9fLl+9lF22S9aa42
tQOAT8tcYYkPaVAG+I03krmmAf9nnAvcftyTLSTQgRytO9Q+R5Icdz5VPR9yfTmxLLAexQjXbfdA
0qeW+L93OSQsQBT1XXUYdqF2CZKGtPMhh5/Y7GEmtDXStz0u8Lai8jcjJeVpGM6QOEehcRa+r+Pn
PbTx7HTO17HdkfgbVZwtIAXT4i4KcY/rOFYTD7+hwNLuPF0stNqGTRlSNiAfpBwEYk+ytrd5BFJr
N9DlC4AMUP3T+u6ZI0RNnOg2lw8Zd/T5aeUruPIhHK3jY0W5vc0sieFxlt8BUbX7gCprapE/LulH
0zjGsvqR3JbhPAw+pXXOrg3PBZZ3J7aR1tBqhusX1q4Iobw/e9uViZszmpkou+6tQqyGEXzvi6SH
zqw+n1AGDnRl3l5+i8YUpG4ZebIgbd5LuDcF8w28yMOOlJfi2XqRkuodyIOplvaDCZRlAilkdAby
8ee/bN98vZjfxpdjrvS0XnbEGHBCHiVJGzlgniKfVPrXFCWwHsmVEEw3HBr0Fazdd4lQ9+2ah9U8
R6tkK3nRxm8IcMv38eg5aduEOdsLkCSX2n+FXCm7fcn/wAuBKAqrQpCspLiK54Uiai9OATMzdf3K
+BEHyC9ajUGf1OsFwrQLxCF/K2xHO00n0MuR/Upj8DnbnK3t4U0UyKL1K/Grt9JGhdrTd4AIKFRf
O47LsanEw0XY0keGmsqFCLeLzGZgIqWYwTv1KtCHH+wSszdICWTgY5GPYIZKC1i0W7eVik0QdpKT
jqMwo4BJmH7b/IHvL5pNv9dUv7V+vXR2fOOIm8vs7PTl6yeDzjtTjSTKWOC2GJ/CAOPpvHXK780M
IWjY2fsfNTdC/uTx2QxFpiACC3pecAi3M7PduAuFvFWaSQOsRM63jm8scygQsk/8AhR2UjIENTdx
SnRNUzAWL3GKDqDdpGbG1R2zVyxq09VeN+tA41yb1XLr7C/tT7ntZbNiPBn8HvJmLD3X2cDv7stZ
ZYjMbUZMxldTvYDHPiZfYay7P2P5ABatZCIfSjq3Sd8OjfVPnYFDUBL9IFp0u0uYIv662EP1hAJC
QkKRTsUWa0b6jhthbQl5ebBAL9IO7U7qafCB3sDtwEj7iggpUTec6pYspsfPtMWjCHbZZ9cTUtIi
4N3/0os1+7kLymHiI8tO28a4/VMTnDojD3yz2cVP7X69maML8AfIdZvgq6Lr75ZzupHRjYeunYwU
OZeATy5vG6UbhAmHF7CK90ED6meMq2o0V9yLEMccpEDvPm7fVQCIFw1EzsCHRqtG2IkOMBzmW5oB
9lKRbkWWl3/YlMxUJ60C9HoNvk7BOkv/JVs6PBvpyz6FW4bQSp9vz+qhJCRkdlsxjh+TqKViEgiV
n7A/eEkX6oK8mFAYVa5FKvK/lLWpx7snO0COGr2nlV5RBfMmRv32hD3dWg1D2IgY1CwkZoZ3CBln
2PKEJzZ7rjJ4oR4zoSo7bpa7mrODlMWVboabJg1ze/ygC6lW55MzWih3Dx6bXZ72oHyWr0gLQybz
eeBE7XB9ykYFOviN83iahAvSCyc44dSMknyRJe0bEE5Pmsad6c/rHpT7jhYE5VwKSuH2TWJ8fNUN
+qR59dSarNgxnkZJeYpYCnrkA0KARp4P5LojJxbvcLXsf65ef6NowZLVuEBNQmeiWLav55cUeHSU
x92MTw944lvv4LVG8YgTXqg/010Mq0WgyPz7WIp5kMTNG0P8HK9ssEUDz9iMNKm2aqQjLyFBwfsB
O35jH6wsglQ3DCspLp0HWrl8mlcHpR2NpICxGSCvjYCNyqSDu1mIfjvH/BAbR8qV4yTdLJ87OmnJ
AMl+hUDWvc0ucNh2ZidefBUtRqYrchTVDf2c0Hq63CqJN1aRDH/Kh/d2FY+kb7kGgSYFDNl8cK4A
h7N8ifRoJ4d6fbGq4r/Nzagjk8UZ8LEFS9Pl7AGO3Tn7cHrzklBKRPzgeIzpay5jSjueTqbPBbPF
AZbgtV0bHBuwajPYU6Nm3LnrpJzrI4gNxubgor2QM3qiTrlierXIQJoVNY0PDSO6CMEldFhF7p+Q
4wqjXsTp6aLdEG1L6vdXJp6NDgl+kK0NvLcq6Pb3RiCmNp/jSx1bah9+3XcuuYKEWQmaPRERejhl
ikcfsp+lWpd7OSzZbB5wJy9GXq/+VGzeafF06EDdcA+V3PnCQVSe1jb5tKroIyt+mCVAQRVzSWsS
Rf3cEVbxWsl4ubBANEE4XjJ/Q6rCDdIPq4vVKw0Ny/QQ209E4kgHgGgOIMjMueSaRfjY7jDKguF2
FeKdLZDBVLv/13ySTVZ96Q6VsuwAgXj5L6cI7pbDgn+8SIJ6DAbbVtt2tcaztooAL0pTmpCmOwCf
VLpml/KG8WyPr+zdq9fD2/mBUIRKvHbzq4Xnn+oqRmpDMDTp5VA1ILyT34mjeNB6Ru2+WWZZh2Vt
aBq1EDId4kktr7lc9u0JpK9urp0bW15YHmh/j01Hh9mRd+oZRGbVob1/+TyRXgQvdMA348f4D0yz
9pqCsAZzxhKYEjtqLGtLEUUcSliW4oiVuNzjKLchDtW9ZxAxHwHAJpBSxe1oVhF80Oqmb8Gde96Z
Zx2S24RHNBosMKzoELJtpCNfIkkyYOqaaQXvBgA8+iI9HaERrjCs5QXjVoS7ZgFPTICDwXLsttPg
iEoIpiZvc1n3jiLl+EcUi6YNtK6rwbKvR5NIvBjDFv8XxFfnhlHbjQUIcyobcb6gHo+Z41txngdR
ek7FgFs1LXtQvokxVJcSS7bx5ewIBvhV9M3q5CdzntQ/NmW7oxhHvh8+fYPgWtYV66AfBwJZBIGj
8TNN7Y8wXOKgj6KF4gSPJ8MvEV5ax0zM25yxlKxvn2oVKgJDgv9jFVLxOB0vnbinV1sLmcPF4RB3
EKsO8emweh4Ay4NrBIY7XdjC5E2/gig7mk+hzJjhr2vN+rwR0Xo4SIWvtZePe3JuElzfM6NnWkcP
NLgzFwU2/38+83wXhV7hCOHdW6NBNM3I9Qw2mqYzx0o3Uvh/u0mOLOtXSi8p0iOuQ/SM3txGqSIQ
0UdXvcmE6A57vUhl5JymThxdM2XhQzJZ6pzSrh5n/FxAZtsQodO5ULPKn5plyedK/cbOm4Krbl6q
GE/ynMWuOnB81AXOKZy9CQHvJYyjEg+dR0LNMQxV+Df22Q+6wwdheMHMpsMKxHXsBIJJX5yXlg0j
3MxMlTdD/8ooyTK/f5gB7dP74xDA8KNshc6p50wekmpgPmTgbRyAF64MdqCRnQ5D8pfsXZoyZZfU
jkiybiOhM17bCvbHWltcApaKCg81+7b5vLND/gmAh6kQyNBJ7FTYT47ZK+1fhd/AGQZjaKqpDJpG
+MfQtJghYol3mi0p83I+DYgE8Q8rF7vn1SYqJIhldi+ItO1VMlx5TAqpx+Xx6SnA7UJROg9V64R6
dbZ/O8qzmdNM3dVi6DP72yJ62WCNXjVQzYdqJP8BvAYxBKYbro9M/YSlhH7pEnH3qmHPS7OK3EqI
tUR53GLAyrVwgh/71qRacKYk+B15XZjwwwFonRDV5NXRx8xnt19QoTl60790RM3lkSkOvhDnK4Br
a8eJetTssnOy55RPTIArKXJzzufJfBiuJZ0+bA6REHtHFXQ4NJTXlhE5MzbVo+1oYWHo020QCN9C
tgq82A5iMdvaSlCguPD9T/ngEufqh4mpI6PjGPNxPArElv1IXOZF38W9jQ+qxjLQgcAG0jKYUg35
s5iifPYq0GZAvirJj5beH4Utgrs6B67zrCj76beXy7Wzx/QLUObumA4SQQxpTrNbnXL4OzQvw049
LGMUsyX8hZZhrrE8BBzGIEou6bS3p2AFWONSPBR5t+q/JVtORpqQJTQq4cxK1wZDSCivvIuiCtra
q85fa0uaFSOlyhtm3G6cmD3vDAjfVgo6TZWl/CpZSnsP2t5stWIpQj8v0uDGt+WApNpWgO/aJCvm
Vuv6mLrw63oGsr5GWM7ZLVekVpgLX3bSuR5XaEHLgS39rxs5S7li5ymu+c8Frs4Fm0HMugiGRiiX
q8e6BihG/zdEISY2GadmneGV4Z41HJAWIqW2Zody/pc2k0BuxL3bePtp1u/D7h+iLnhM5mlgR3Zy
pWnXJtKGeMjLDC7t2nXfk0n7GemtklZpel7pstZOZw0b6iqLubz33yBKs01meSc7+zw/yPcuCef2
yTQ5b+jizlRUA5VofGpapzgopjNqXm+o349kVxZQnrC/daezX/huXMQ9oR/Kxa/QhMGo9pTG9/iJ
UerB22Fao7na8nPpwJyCHIJrACdl7Neq8hmLdTsmPrtrtSjYGoLjoibfiIa8gZytS1nS7R/bXOZS
O5++gGwguW4Ii/GdMnq8HE3eBtjcfP0AgD6T8U6BspzSGNS5Be278rtD7eDaiDGprjJ/K3+u8mpE
B0uStLy/gsqS8TWHaYzLNUfY/CePUevV5w6W8kdjvPF6aXnhxjuowUPl8es04d1raNuOYXNWfqML
qilRsJlGyn2Ukz/O3rfjSPAIQkdbbbTtiFLyNS6qcBUuPGpRwJBIUwrD1cVpL4+ny47oGG2ugmvg
aZND+XxMhQ7M9hBU0gRrrQr4ljLIDQyNcKAbOBAnbF9iUkMNaM2tambpelhAvqoXEbeVlDHyYGQW
2/5wAlQc5lr1qHF3bJmwetOItBEIM37MPXAkm9uE5ti7EvNWlM2iKB09sMkR7qx4vmLdr3oXgltz
aR2Ma/3/A6y0x0BWFt4X1rocenocIe0p2N0Sadd68bMbhnrt6yn1BzbHXYtKj5K29AcSxDkmxyp3
xhQVAddDZ2+y712YLs8DsZ8Yc8gIAjs55zY93hs8HJN9GWq9M83XNVs5/O4uyjbc2SQwwdydU8oL
GnCjczdlhRHaz1VCKH0gSSly3r7Pky7SihnyCknc/jqbOr5HYzNa6jswu4FqA129Z0MA+4BCG6bG
J2+cmVCRajRb8z3pAN3LrYJf21EDtgj7CwBD1E80rgdOF7vW0wUrw7rUOkB3vmA1Xn4fJq5Z166B
sFZD5RiwqI9JZE2wXkStZWP/MyaCVIS7rshV0nwXBBcG3WlhemAoGwsK7EjjqHG9Gnd+0PfheAom
V21Fa+x8zaWW21PEmwXR7myhKYMy/mYP1r0vLwSQT+vjoQ18agomIrjxF70ZMD7H5feNbyORdwSJ
IAuMEYeCT3MFt5pkXklH2+yLKcwnuPKolvuxUaitmZ8fXXigbkAiDoA2kNXQknJuT0UGIK8AT1Fh
WbYnzCPdYSI2J9r1fLWxoi9s/XehXhjrAmli+et44G9Tcp1pxzObZrAj3yppcSivOqChJNKPb6hr
U/HMQxZO5krg1RB6Fht/KmPA8GXK4PIZRt2ppoE7b/m0EtWg3Tkhcum3I9aHt5IoWTuXlto9+OqO
r/i55ozi8PTXZ8GDBa+FAb1Qbl8drqhXEztnQ4GsuQ5Ox6Q1f6oMLtmZJse04UbF+vZiXx7BmSfz
J+d7gQ50m3c5rbod/gDc5mTgwTNycACYQAiLjBjMO26SJFiLavW7ArLGTKBI7DLOJechdbiKK+N+
IuLvewflg/ySw3pfYAuTWEybWbaHXgsqneTdur0unxuEsTLfnlT67O7MKO5KFTKgs7lkAMkaBrGV
qvivRhn/DxIQXaMev1hV1LMt3WsbhGZQalG3+4deo3GmjwG7RAR5P/8xhRslnQzucERJbarkGo6v
e4DM/JzuKjoybHNHk4JX/98LL1O64JuftlOJMR3q/4FYB8laYC/2tTAkOeV6GGhhnCSMDpX5Eaii
KT+yPMOqiVdsy1T9RHLMfD3i+8l5i7wSmprKYLnSZ2HKcneaCyl2gv+4Po1LYTFZiZJ7zW4Hknir
pOjYmEBK17wE/yCGW6EETDXK1dkvK3nf3goz5O56CWu+yX802ZMbRio5QDcmlMeCyjHKvav1qVy5
FhLd4nLvDSUeBMuuvfERiMJtMXFviG1gbECYzdKvwgfC+TzaDWLMwj9D4i1VzyxFcFfcj/1lzh5p
lTXQiaHowjMDyhCFnjEA/Jm1IrZNFOx6GPGjQUm6jIb6KXEA96xFRXtudDHsxV8TzqpBO0BPgNwS
elnOy5hUgWgR1kK5uR+q70wWz7Ij1te9JeVme4c0MmieZbULbsFX2YmnA/xnaJxEIDjg9RMWgkOv
d4Y7QhcYShFyvWDb97Cy26MTbgVdkY5W6dYStLBddk5q+gZwpzRWljh2kY8V4qBNwltoW+M859Gc
NvhIxuvnk9wvR42rFKk+jgnqjSS4t1kZzSG881X0Zns2EMlV5gNCZ1pwRCgjDzdmWtyplL7M3Okl
smmmnVJ8WeVVgDYtp57btrMan72UE/KXau9N2qcNcRpJLIqj+oQKIqpwMwezURKRmw7z6q9Tk1qA
Cb65CoIaqKrtS5icXEbFgT8kNxri//nm4PyG6o/PtvQfOSvRv0o9WeWhMLGsqUZhM3Zn7ZvoGarS
YznOhjQJpvtm6HDhuv1RyiX5ow/knxqDRV6C0hJXlwbwRwBNPpCLxZ4+J6ZlTE2VE1tvCUzgSNYM
jkPqg1G1Jpudwvz2ovXIXMo0/BcmcdLHqMNc85e7kAVzjPsubbwSnGZTwfgF8AS9JAAJyVNGwFny
AuVRqFACpw5UJo3dM4ucoyiTtFEcAYlzDJINkJ6AoLOphQ8JGfhEK/2qWHwv+iA4fY2WNrwOnHMt
NHebG7RK4RIfuiHlKeVhAkyfiv4gcBrQ2ZDQO41oYp1IUjf1R6KLaFpntIv5M5LQN8RkGQwdku25
NuTbSH9jyBULE6+sZxsLmFwtlvf8vHdTXbWKmoKzIADHjE7xDxlYSTGfxZRB/zLVyj/bdLiLODNs
c0MNLqxtjMODYLYW4DYhNiSgUXP+CK+SEBnKcdnjykRqLy0mqaHS9jDXIyIztNJsv6UGpQ6JGiRu
eKvU1mZWu2Sb5k14l3WGTBIYOPpFefu56y05FdHjj/c7bDJIudPydv4MM/glXPkKnwCD1QMQpj8l
Y+/Q6Odij5RwL+I4YcJippiABfrI33TeAqCHZ3p7OYHeGOBjUMTSI1AwH+Qi3izVJTcwefQsyZjE
Up3aUC5VhL616t54CZvILTxjoxbpq+0KkYVTEmcyWD6+o8Bl/x5dlTr5ouv15kJcb9cgIwo+BWZy
RRm/xvX/ndRRCawyVigECLf0A7s/4gHWf7wybn4kw1c9jUu2e209/RRNckRJWopWS68Oew1zK3lJ
4QLTbxS7hop8Oj1VVSTJhDbXIgQM9Vd4ECP+B/dWcxOC705B55rbpeD3uE711vjDLv4iCWXy1820
HoPszJ6ymwkWeAxR4R6wJoUKGEsnmLoPjR1dn9EALdUFUUI3pq+HhXXy7y+wBygsccwtO02wxXZe
y9kxayHPc4kVwhYPhH+U84KiQ1SguNDSG1dBIkfoXH615bYNuv/6olyNcyeXttiMuF+rol28eAvj
Dh/ec/XIa+CbleUoNft4m2uwoU2qrJWGJs+Tk5/85dB9zyjkYA5NiNaKWwX/E2dxzPty+omqXdYn
pduc01crZkdENvENJmNFdjHAqOYCQKaOXiwLHMpx+d7D/xrJ1kz//vvBLo2QtqU7aYAd7aaXM5QT
GYPx6yNsWWvqrunWUZvIfVy9QVj5eFkU6uEK47R41dUkAoUoOgZc37kgqn8Lx6ScHZtz/tz7tidr
CFBdJb8COfnq+pB5tDRY4uDpBh3IEgEV/4IxK5BYOD49pRl2bJb/WzA+Ysnf+Q7FpPVmW6alsbg7
2UhKWfceOT+nWCpe9H5Sri7CFsWg3jRRlGC/1YII0igWk4QixdUiD33M2eD/wfZiCgto/mGkrUtu
cu+ncKf3JX5fDbJQEFBBl4bC2NUm/HBYdxLfumSw5h0nddDSElCGfshfQfd7llB9GfMcrxcvE5qR
x/falygvJP3F318oxwC1xlnSFfdHYt3odcrauV4nytiTp7ZH1OpUr6K9g91UAWDfjsTx3Rm2cbXm
lGFNi7f5HP2/iQaKJc07MZMfioKaSKiB14G9wQUU7Ix4MhgAbConZs61MERy4SWWe/Sj5nTJtOat
QuRyFuoOhI57VuCCyklGrsSdTtoTSNGY7s31L3w3aHMELRugZ/i81I/1ttLOo5BhlZTVMQvvL4xX
sPWRTVHe3AH50z7U1Lqy2Tla6bARIYAEXciiMCTovQi60FeQynWzA34kavqyr/dJnC5oZ/Vh9qFD
YLXYUGmeyScCCfqI279FszFoPmbdsjbNPLPUSck9srX78NoMKkqLgP7nuzl105G8FIFoxRCGQmDs
BKecz8JKLdjU2/Qx1HBu4VPOAxyvVL7XwvVwdsRz0YEcgSEMPXdS6JJnTo1oZZv0gT3YXMTRp6CD
68wEtkxuibedov77aOS6DAE//FIk6j1TxowAPnDc6Lg7a7HtoJZ6qB17r0ibOYPJO5raorWpRSAB
UpiIApUWBzlsBOpgMAv1T2OnBZrf9ImM2qtmmeYtcjakWgx6qd17gOG3pJ8NgdFFXvQj8I/V0qoV
kxnylcW61f2p94pPI/RigHag1RE2oUVndxlZuX/7oNOWEpRJ2vqNYK8vTTGOQGigai/tznPawOEy
VMFT5L9G83OiCMrhEFaFzi0gq+hCitD2eToQ6I6Nqme+f2ziDUE5dIOSWH9xmQihqEtnE6Lt8YuL
Nnn15Zm9+zMaf6vwUlJ7AJs1PZ/T0js7KCRen1Po2D0WB6FVU3x8vWHzfIV0JD6bt0LyPNzG8Dye
nR1nnQKAS+DS5f5G//b8B4fX4GKHWqqGTqFq4iAX154ASMGZLBGGWlKRCXyIOLcUN05N3n7k6NcD
GkUtCV+OvzPmUrxEAj5UjYxLE+X+AnYKJrWKmR2VxvoYGDXIOAjZajhcR2b7ZidEH09ZYlWoWXaT
bne5cxATAt9kCLzcZCEkEv6GebnhaN02tsGN3zOCTZCorENMIMax9X9uNwKZr3LF+6B7RI505UMz
XVmgmSGKr6Lsh0tcUbt5NCgRaBoWnFUbMVitSHMGYRA/hextXfTsTZ4OHH9A9gDvWyAkpLs0/kI1
e13qdij7HEoTlBcTkHsBveACmXmrKW1skfRpb6riqYiUwfeZ/iBrR+cj3Wkih3sGIKaQhgjjjzke
u2wsdEemwd7BoFgal8y6xKlwyLA7D3d3XUCqRk0pITOPopYNs2nsJ6eJwH65BYqZvnIJ6GHX7CuX
3bZfRNnBhg3Bp8nGzKyvMp5b/wrFu0VF26WXqEXduVS7YIpsAGckw1a6FChr+huVYPXM8IKczHmS
S4wNl0Db+lWVcviI+C4aPcUNTb9p3GioWrUaXOhKdRe9HBgBYbqm1h9/uE2V93OdOq6GItC9T2RK
jjcLArIYYpbmhUPhdfOrUISw4oXUhIwTrF9gxJDCD6yKgzIq1m55YBU2Y7sVOIqykjDo5C+bchJk
0TLIjfZRmihz9NjDVzmjDEJo/dUmrVCn8rgFft+z1kB469T7CV6fgZinyLxBrBUn8VRj14Gg5ugV
srkaHIXrTaQKzRV36OuXjIA19WKd/fOB+xZcEB0H/WRlBdb4cBxTOD+on7g2LUsU6zUwkiTsUP5w
DL95iXnM5nCHxjjdxmhWpe4mttKlV8vN8WpdYVrG+HdgcohqBV5soeZxs+4xPdMD3/xJqudMpiBl
EqEUMosMTi1fiC2STdTuLdb9dxbA650xa0tqIkSOs4yWWEfgCmzKx/h5IVmeYq+zYsaVzdLarPL9
Sk3CNraPv3zl2btj53G/A6G2owgPZvpAyvdCoLQy9mhsk+jW4bbsLEMQQapE1t22hsetXlBg+wI9
vqlwC7DyzZtTLA5zIapTiLtoJzMEAB1q2zw7ZKr8XBtGRKLulWd5BmThh2j6uvT/95YKYdlloMF4
JLSbW5YVJ6rZ/wXsAbPFBIPwWU/4q58FuARCTR87tGvU9OVMJidOAd4M7M5I4kLWnmc4s6R86kfx
HJC+aguvH2vgKCIuC8wLQCXcU/XsMumO7FpisDoOgoJyaza6bPwBiF6gNq+DFpnFpZJGKkEOQ88C
7VcFPYanXN5bDjQEdgDyCt8MR8SFcH4LVf/fhnkpAWIAvAW+hR28TewvcqWmler15a0//6DLzfeL
AtAUQxxD5O0YtHpk24+2GJE8Xnw8TtTtJexncq3qCBlWH6ApI+LSpxW0Y0USikmiqI/Wn7U/hZio
vO/fABaYXU2Ndh3Z2+dkChwyqX+X4zbKq9gQUt/sNKNXA70+7R4UdeVs12Scr9M/HrsxbBPPFbZB
b8TJF9sl/IQB8qzlqAWWo51649PTioOZEfBWxAOh1ux6ajrcSKgktl1K1ncXolAH7B6hkKbKGMFo
wt91NN6rj1bJSipi2PdXo7A8K+hYrsZk2y4xUJ2Q5wyIL5prAww4oIjgUEuy+0IFTiyFX2JQ5vT5
Mw+q0jIU591Iy2IvlPyrYyrOsWbCKax0bQ6mgsMXFqbLUAKk3ReqIqZ85CcoT0LAy+vOzaLtOAbB
SfNgJlr4JyslO62656gAx8YRbKpBMQl35VE+PCrmBa5xL91u/nWxQ2rcob+cW4pv+YO4uPzUMfa4
l0xZldcZhdWefs9bM2uZuu6oPLeQEkiz4EgdOKZzkM7REbqpzbBpp8VX8EUNRm9pXOxvtiwfmgVM
Qy7jhqg6CX/LL4ytB8V6WZNFRk2YXtJ86+IXLVYSQJIt+dB2cNFGmYhYb4NM5vUlzNjzoQwE3rxk
dm2E4OPWsKHUYp51op+6Jk8KW6bP8z5vZYDx56LqjNLuuapJMaJoaPA8Oc2py6d0blbDkB9/Pg6c
S2nl5xcaOeiDzqGp7rDyh7gRUWQBxKJH1uCRHMlkZVL/fHt9PlLcp/QHF4piZPvzuL+r2HjO8B4b
FdFvIzQWP4WBHdp0iQzVrwm+OZ4by4ro0YKxUxqlenRr8gjDdMLNpRng84ycJZikl2GQN4jW/ppa
cXzAlb3l9AAiICCciDiOA5OJlQz7EuJO3Us1m6UpJXwAGF0ah/TUVtaRy5HUbRcOiUhPRg4lkbU5
dSLwgUdlk0Lm2Jf9ogfdZD6dAIU5hp2nJ84i1NaCnhg0Cc1eUX1sK+fD7tIGVMYEHektaJNTOz1X
hMPsKdITyuAAZozaCX8DT37xTXdXKlzTfSEV/ikkvVRsGwVkQUv/EF5qxOtjyLcErMxAmYR1FMxb
SGsasAVKxv6mTRFvUiswspBErMnMXclvzq0Uc7anWqvjZ79EzV+BUF/H8CjfKDB/IgmcjQYfwasQ
BXsGrFlvp7HVPaSKHi+f4hj/bIepG3dz8lGp86PxGEI5+sxV4rJYVSZ1TmiGfgscG6ODg+H0Ab4a
mqBzywtONePCxyp03DfM/5QrXGRpGwI4AdCMQuHgZ0hnGYWcW6vTkgW/Q6PxmKLvEUXk9y3s3tYf
4y9gHFvjewDmLgUrhHf/lQArpaihtCytCxTBCOT5o8MIeC8p0g1IMlwa+PM8zJY/KbIlzhFPkDG9
uxjyaMtIrR1E7Zq4iNF/AJoM+Xan6l97ksbZXLN8PIsR4I281rWVeJ9WyE0DxwCFkqNEiwN/SCJu
s91gfr8jv+IXXTfa68ZrInFxzGwCQOA3ifi9vHZG4RE7ntXc+zaqqwQlHoXeypE0AaTUEZccnaL6
EOSHFHSXB5SmV7DPeZlb8yYFqX7vc391k2qj2cPERHMdFaaIySGMYGjYSawg5APuBrkdc6M4bJRF
k+68BY7nPg5GsIcE8DyMeskiAt7ZO6zZ+Bzi0HD0JKlLH8ilDMmo1FkA5mI2OyiQDq/nIpz3O/Pa
+xt2bpsEXZU2Yes1/9v/cB6Q8m/jF8wK19Y+akXpNqezJzFvbuV05X3hXaRHwZQc8EjpnDWqk9PL
967ZwI606Ritu+peCdDJuaMWUWyqJYngvIxIDVh3OUnz/L36vmERkFDAe/5tNY3ip9nr18sVfB6U
AUcJTdzKstzm6jJhItfMqI3kOChvOcxGKTPCvyYTkWkwsWbu9JsV2pLiEhoLzi49QheFMqeLf+W7
+n8/Gdk0iYbMyH/BKsEU8NLI7ZKzwctRm6EN8LgbP/OT/hIE3cw3iR7BnxShhQNXqld9sS3zdFsJ
UFBO9+pUjT/gsu54ogRQrSoIuyGrOPmWjVPbXLKKwf+KZ5yo7s9KwkXfLEhzicw+3B3I66IOHXM5
mqEpMIG9oyQT9jYgHb8iEBTAJm4ajCJ85jjYugocRx7wgQ5s4cXsu7+yOykFZP9knEDSlBPu/VQA
L14ZesmYVVd1m7WqcvJ41rI5hVoVWK603uXPkTjlA3ErnlE+P4pbYwZG1V/LNCkuiSujulqImL07
TS4qJCtaEMCk64aDF/UE42Dnad/IzaTZLpa372oXJx8HkcSoxvfuAJIHxPybjA6DdYvS/JkMH2tO
ISSzjO72oELx6Qy0MdHxwn398AG1lLRGmZaZVX6sijcfXJOY9J7HUqpRhqB2AhT7IO0zNwLCwlSu
qBbGJV6+az84AOQhJiPBb8AmV9TZBbKURVLe6BVsHeCijI9MY3g/+uHIVDSO7YCLXRnD1lhnpstJ
dw3/N+0O0GXDektzfH2e9lBjIblASd2UnovmROJ5jFfej7u6Opq6en0OQJ0wouuG6jtePURx5toH
cNN3H8GIJdAfeIT+EJms0LB2bJ7g2RDIkSacBUj55n8k8gSx3rC15PUJCN/umLyqBgIMRX6B++0W
PA8JuKos2QwKnJ3PVj8Uf+mpyQUd3RNvu/JFoF08IqSfngWnTf2wYv9xHZIENTru+e7izEM4Pcrc
tr9Gi1U9+Z5uwQI7KEcAxb1dA+iCC5eRWNuY4yHFX8A5L7WzJ605kYaJQBLAwSyFc45DXR1BnlOh
mciCZV8d/Yih0GqvJ3nSWL8i6uICnqQAaaBARCI2IlvI0smzMFoWkJF0qAEvEogRi58Zu36ei4MY
AeNsgKILT4JWEOnY/CZXejlZVsIj+CCfdHfK2HsEJ29Qin7hN4eGxl7bsEc4i9paTqRvXbUd6RjZ
4kzqJcoc9JsrTnPocTKysaLIzJdb1zbmm5CJ77txIMbqJOiEt/KE1AYYJCTdZZh46GLmD8mUp1yT
mH5vSCXz3Z9XXGBNv+N76WjdDFGKNrdyzVJjMrIBZEP6uX2E05UR2MPcSiEWlj3wWy75ue2YkKlf
zUESA+74T9iPMrQblE1zEWusIY3YYKHqVh/IedQABdfCG5SUbw0s9175GwUGOCAXfx/KuKGqqjhj
k/kTWbS32V+KLsPzn8/UMp5dgmUFke+7ufygeXHHChQMQZNyIUScuzLuNlGROyeHbps6eAFFtuy2
sd/ILMfQsjEk6KgpzXh81x5aakoOP1BH/eY6LTwsDcenACoH+2YIhuNENFfSNx9t3eKZmXbuuRAh
9OvHrjzCaN1IxEefFcJ57Pd4mOuh+XHkEAmW8gVHMCyPw8URXNJJnV73FLwwEaJuO9FfY0JQBJp0
mGcrrS7fvB0caAy5yERKGt+mCowokX3F0AhxtuU5GgDeIhzPYI9eaXWTIdKx6+O5qpuX/qpsuo4s
3w1tvOo9LUH9KLdCLh3Y3o9iKxucCMoKhjXS+9HySDELY52uscLtloHHQMA0WS0Oc+1zAXatS8Ny
j+DliENYBK3lyXwIbRho2WHIw8mWKA3u3CCMSp9y/M9Auf1D04Jr3nhEwijAIqbBlM2XlW3oixG1
a1Qtw7+bj0q9OwwuGlaJ5sKKESEYDqyz0w+9rSYnF9ztwHjKbtJWhqa8n57r5RrodzgTBsFr3dmx
ETUN50cNWaJqmABQIalGDXkT1zkgjhTcPDYh//hg4JnUP4R42vWpbjFKCE0uBrRXfzdO8Ii9h/dH
V+BOHfrKP/7azWWcCKhNweLGbJ76QkEgaT1Atq61tMXuMe5r5XPWEP+z0ZP0Z+68x0kNEVfsJmcs
JJBcTj9tytnVs6AGSuzvHNpX6o0gpps4Jc/GeBwRlEwfm/ll9tlrAsFCd80iACybBDyUjzYE1v2P
VlxlCkILut5aiN87bC9wjFBTPV9Uj2wxZcdZJ6F+6igRIVoulaciQtjLUsx8d7bydiJ5ciYFf7LU
P7jabWPedfHxt8ZViUBMy90l7VxSpxXVEnT5mk69NBumc42Ak6pBHFeCRisP1OCqIJcNwGfN60L5
6KNi5laVFhqBVt7R4N08xvTELPrb8Xa9JB2WNwIp0K0UPeADbt89rCO/IGSzjauUZ66HT2ESM9mT
JfnNGRkXoC1lMmIPn/xet2nICu3cUTv0VAzuGjdCgPOVakhyG8+La85E9nRIocDNmTuUCPHloUVb
ZVnN1ImrulP7QUE+9nXcuKUtF9v3CF+VnLne8ZT3DcbduTL/cHTg2UQ2ubLaij3NGj+cu3wO9FoU
zmrrf7EVmyBhdvAEMMbjdklleSndjCKOTTesVkp4UrWhGvhq5+3IsbUjyHwrjuqmY75zOoyC3GDP
u7vPWKgTJN4Byb6bqb6FedrWiIeVS/ug15EcdyAzxs/JYhY9Bq6nL8SqizvJKc5ofNypotPxhYNg
rfXRmdKAvl/Dni4eaKxrcw8ljRREGSfySikyICzrm7oVyPmcjN8bD3zJXG1liKZChFb40hrulMyn
U869j+umQ1NSmjGQnfFXoPxaphqNdzV3ZgieTL56AXOKDGJRyjwhBjF293Y2UbYWHuT8mu6FgeGX
N+N6k9NAn73Am8+lgzz/AL9weQjOQpzqPOcHDR16Yi+keSqtV/XrkkiNZe6id48YnsetRQSM3k5U
PeV2XZxaLqnZgwPsJpPCIV8hy1zXMIG5NcSZ4Mw0Igryu8LgeOkTGSpzEt8V9prN1k3j4NZVTTWa
0bacxvUZ08gAuezlsU7txqFMNvu6KWfADnm0s8uY/YOckHXMg7oDhndKhmkeZSlev5aXQTmUfNrF
+hpIT+AVpsXyJvpVyq7CeNfrpnEcndFWoLbv5Z1PZfACAbkhUrRxTaB84vzEtvOJECtDogMcfDuQ
OnuNa/LYXb6QJpMEw5zPLY8bB/0BvihTA0J2fp2nhGPKwXFutCDvzU7At7Va71kzutdak8i6unYJ
ivtEb6O5xu9toTzL9spekJqK168EJbFMP1+umkUS3KNER+GwcaoqLePadL4WeK6ihhnFusLoazcy
3+/RVnvjRos3RPJcpa0BsVO4t4t3g6ldkrfo3UFevNgCujsfOWWDBJuh8tLCwXzER+2bs4uHgmsG
2obaYSn4QVKYStoKxovY4IJF40qwnSOsNAFt+uFfUcS4ODeVbqMw2vgDoAXhCU1x/RRTMwurTHls
OfFxXa9kZCPrAWrXAMm7O881V7oRYgf9hi19QTLOhxywJ81uf7yZsqXE2/IX/RBRRoEq0Fg6m3D0
7aE3bEps5Jp7C4QgCWfIoMO9jjC+1GukMssGKeguqc0lYyyl39grkTb68l5ipodfGzn1PaYGqtWg
d4qzLoMzslSV6M+JDosQVWeFzjchakjKzs9c8x7dNyUk1wMo8BX9JsjSk4Y1lzqRo3Qql+7RT310
fBBmaZFu7S//tzbLeoBMvT8QqOesgI4Lo9SCigvlz3XWJVEle89pJ3Cj1xH7x1Xw1RdkCN5J4lQ/
50MHvy3LeAwR3Gs1gzl1jUKCI8aqlYZRbNbs+18U40ttcKdfHBsXHyUkbfoBP+oCCpNe5mI9OGtd
acz4ZmA/JsrionZ/ycGvnJoXShzGSxfYN0Q+dBGyAANMPqLR8Rqr1PQNYFG+M+CPxasLnk8JJrAu
7CGoX/qQkCPqjZkmmkJjWQI31cP01xl/TCbA52vWVaV6s3VCGm1qO9gBiNt6378O9KB0QMkCXM41
bULESTIo2Zn1/9iGyjOXEitnKIMY8poiRcklQz/tKyyMEK4BsXqNLp3bmEMWDnRgYCAP605nAajt
iY29B3O8aBz4m0VDyRQLFHdg63eiwj0k2gKgOux3jxTR34BVBqidro0GgIFcoqzLVRbwtNlGLZnt
nZo9Gjg0WiHNDhZJRDqxlt+k8ar3Z/MSonmrwPh7Rep1Bmywk1rBqVme+nIj1+JwAU4N3x8+qpgf
Je/4Xr7eufFRbv+OUYeNPbsM9UK9bHMYp1pOz7uj1ey28ZUVyF+WX47GQmUL/hNKAsux5C1C6lN/
Rio6W+uzD6Md3lT/E/PSpIP1Qv0mmIyBd+/njqnPNLaoo22Pl2jxvn4vsYJqgk+2YdPa5mvJEPwP
cJU5tHdiz2yb70cpiGPxevqpJPXCGzKt5DnMC3mMZbt3ZmRHVriJRT9pxfNFEeMsU+zFz51FFvbs
fq9DvZ2GMZlRxU7ssIZr2Kl+EejYtQkhqS7P/zl8rVoe9GVMb7VKBr88EAhfKku/7RHZTeBs04Q8
1QdnM2P68TuD8ddmdf48oi9yIjc9x4/Y96+lnu1aU8YutQ3Sd1SnFioZgJX1Z7qlQxWQoutBvW7s
COwVDQt2lviRfUD5mF8x7Yf+FzcHUn25W1gUfu56/+3oqhHGR44AtGyPrPbYi2U5ystLfkKmpLXu
Yi9sRkV7RbMWE74peR8CGFVVgvupg3/7xu57FETHxRo/XuizZBxMuVo3t7yLWEA1l6xBSFQpeJ4j
xnlSQUFplA5P3DKVkSBlMPG/xTcPmQfnC6tWMqIGhkHzYhCR8xVbuHAti4v0MIRcdwHwHuR4QLKV
3tRdr7UPNThjNeSrnQPsxYY8QMjLSKr5xi2lm1aE8XYeAEqSbYts1oQbkw3KIVMRB0X65UjjaySX
IUCje72QgozXvAStl9oDFEnXwOx57mCT2Pu4alZH5jRBS0wsdsQ+NsU46bh0uRTNakw//5nPnnaP
Kb9wni0VSrVPhKwvX1cIE43rZT/MMzBYHwHJCB40c0o3NjUQgPozPo+n2FAb782Q2HihlWVXrT/T
AdSJAM8pu2gRmQ4TjA37seB3zM8bk8dyzVu7uQU77DcVrs/jZlusKZHEjuu0zm4CplRA7lNSzKDs
vo/07bmzmDyW/0wpa0v16yyFAQjgK1H763fPiUbUd8uD3s3h8fltinCPEtNA9YeyqyfmYcaowWKI
TacjKALj1OLqd2AMYrdybA7S3gRkBnVmrM+N6ixpVJhk7/w8tctPOGcC1dHvbuYBlpA1oCsKg7l8
wijmuLvcSAMhei2FQW2KJQ6nk7vSOM6OGwkscbscKkOPthoLA7DTMNthecQnkzboF1XLhvn0QN4W
kgTS9h2APwpfatihn4OWyooPfpltaRwNimio8kfad9L6NlB1HblAOolCgeJfs8cMAB6vTNulPsw1
MobTstf+0qAYFPk+g55ohuPbdySAy7SJ3JDviH5gNh7+5O1a5LUWvG7qjkHFZ24HewdXLAOa7MDu
f18ruy5yriGVHlLjdIo5KY8gOLJQajOeLZ4Gdnkwz8glvZt1iny0N8p0lWcJFb/LhikICU5amSn6
T4vY5nNPFKVpERmLtoEBgdIQwYalS3eP37BaErKELIfo0yzoZrB/UIbQUbEkaObLYHyR/i21pkBc
3hzlAF9YD03Yu9ESdEkrwdN2jiLupKSrDRJMQ/jQ34EpvFbRl8t/i0k0gK9V0iZuf88Jjns//FXQ
anJoPl1WCMdnbisa3/h2S0KJxWgf2zG1iVheiZdLrmfEyNGUjkDo+zDj3RNqI6x2RdyUT0ITn0T9
42HLeF5MIqMXZT/QMEv9mHG0OxaO4PufDDReArb1cEepSDPn3xVuudHk94m+r0ubXADgNQomd9RL
2tbXpGeGOZ6qQwQVPc6eZnocJTQOvQgdkNbshC0AEGkypw0NiaeL7v7B93UGnDdgPssDKG7ZBUi7
gvw6RnSomBylK7HYfcVfX/6BJvz2EiK9AwyOvWzFvM/EWNQrBlMz2NlZfwWUwwuiVdnkA00wnIcU
/sQMGLf3llreCH/E/nQYftAuhIKQNTQdrGrgq9VqoFokOBZA8Lw1W71U1PfveHIJoTVaV8nT2xZ5
WyHbGB8qNxX8ST7uCTGIN1O2Ydae132PglmZWs3sWYP8u7+614SRQ5SKzzXcO49x09x9NJbQfB2P
HNtJjz26tbrbZUudEuNxWZmx6QukIrijMYe7eDJAdMUKfNxFbpkjFMXq+jpEYDbr/GabWN4+QDlX
dUYIX3IHmt5X+9K34dybhX3BXLpL9LDDv3HwUVBel39Cop4x7WrRnzr6eBOKVo2WOgA0m6KDRx4D
S+So5yCFLsmNiGHekmMJjRhZh7O6Y2vYu9w0ByB4X+nTMQJoMiAzcOhnTTRkVworDCO3tcgl4vZV
xFAJ3qCJMnunRWrOWIG+KYh2SFB+7EmLx1SirPgDJz/1PSgQkIvMwnphzbdjCKc8JzYFIj7gvly0
wPT4OmMHEFV+YmlrysMvV/Q4/3w4gSU3+AwriYwGMJ66DihYdx1ycnyI6ZBejNG7u6sddWGNT98d
4I8uOr1gTsmtIvMm14jT3JMshsgOXoOzxwxUKjXgxSfZCKDc0kCe9xJslM3l6LiGyg4VOfLWqiPz
Zf5eTuqRoW9rfm0hEsbyesqdH3h2ANDWJ/NkJXfQQ7BEpNrlTDq/zNsRSfevK4TN9nLKViY9kTel
J7+cHwN7B/jGQdMipjDkBWIpXnVWOV2LCDuyxEVPuf1NXupEz6gWDssLHem7PofVu9Ns6MdITAsK
D7ALac5dlgod+NGuRXorowkrcRFcP349dxR3USfBDsHQ4EA/Ay393HJm/j1e/bzv5F2D71xQrWTn
qBov4Rjq7YgbKmI1uIAJe/oTdAYTuto6n7pIQgKLaMwEpSFmw02gVz1zPDeB7N3zvUMOtwuK2vsp
uIoW4X4B64GwmVo65tzor4ldfbRA9YoeyBJ4mR4Fv5xayMLQoRKp75CPmZB7YiuYgw8a3XmC2u/E
nGrSPpnbEHu8OrKwmjpi+mLsWJA3JxBxBmV3GZM/D1wXm+AB3xM299lyNWIAiPShnAfAMUmUM3v6
61DrxDbU36rmAAhxYNi4q3V4gAw4JorUqTWH/lILsbLpdvXY1L9d0k5yiB4neoYMOFy3IuLvb15H
dH1Wr2TBirr3MhsFZhPz2e5kmLR1VuNQCgqGQD7K9Cu2GuuJmozfj4L/1BLbQKqk/wIRWxFzCpXQ
YVCkbacExB4SNdczygLJ4ULj2CkFV9V4LCY/dpJ8luASIvidjwkUgrrVM0GPq2WA99CayoleuAyu
OVgyDt7eIvGuUtF0RcmYLaI1FiIJB9IL2Y7DnfoRtnUaLadDWWrLtGUSGOOP6cHPlUaCnIiR3Gw3
+ccSUR0gh6/LYDD1nxhN+nHKEaAYlcoVRUoC1K5LaLrkMOZIlYGE6I6/AZYmulrmiq5RUDBlgWkD
f5l4domw31PhtP3cLBEtHD5r3Fl7V/gzq27XidwpSZypsKs2hjnBvJmKSW+NCllU8tyW9+CVBbv5
H5MaDTghMuJQGCjhLYmI2vzoPL4H01nmxX85JiL+tauPTDdWe/dftlmlJujqDcKokejrhhKRbYI8
VG/gWyR3sYHwqbN4xxj96cho3C60++5J2Nc7yHfj/j/T7ursAVksiMhBPrhH+OL0hQt2TqySz2N5
EMcrn860CrwteeE4nVqki5dkAuZlmzHnldyu+5aYRloZRAkgG1gi59ftG3cp1zHFMvQv0jDJ5GsH
jekCsbVfZhlfjOVhY1B5e5J3sWk1PbsQuijsFb9u1rKARSqyUGh/CDoferAS65i3zE689DMjBFoU
RzVDABgbYU+55o7dqMxKZqokGl3u8EJlZTce+p+4h1FTcLm4+5UgvvlT45cCXeawNuY2WxqxcV5N
9ouKcmYafl+u0mZ/X1xf46GNbdgfQDi4bPKEWJmkhJiYV5xHTcAuiwbdFKhMw7k6B3qKpwXjQNCo
w1YTxv6B6sDnPS7w9tggMyNcuWMQemaY7Jj5Lp3Asy8cxMj04CI977nWbOSh92zSXGJ2CTImbK4J
HbIzYQy7APN7iDqRUYHSGM5uIwjeGORBeK7IfSsTLkmiftGpH0sPeHbH0Jw+BGff9geGmnszfDIb
thSpyxLmjFv4KDfVxgEdlcVu75S/3A1ZANBSdWlF1pKsyLjgtt/04FLRVLlRxUBwkKy8XOGm/Gj2
PRmQFVWx2eSDKlaJKOJSVznS78y5E3KKXnu56y5QrS9wikl6IDv/mv0btZIKkjEc2Pjgqq7DWFuw
c2Ozhw2u05WHXyPhuDzB6ZCuPVgS/3VyI6nCbTs6Akd2QSyFuUSOwbWuQDojd1/QYxDB79bIBhOr
bk+9JvADQYkr7qdtflhbxVoDqK1BkpP9Rjoyewsr9WHFDlEmopGA4WK/CjmCuU/nnzRjioJTHe+U
JdFuzIrtFPEjzI+mYoxv7nOufImsaJ9QRT8zmyWrnfwe4aJ7G/RpVp8LBU7Rq72EuBZcOCZKq/2B
n/UeVvwXQuDHXaDfhkc6CjLipH/5KQzFJWc/QJwzfLtzP0lc8S5npFAWIc/AHs53MpXESGockLn1
YHe3+Jo2ZC1Zor7H1uqm5XOqF/V9h7v95pGH5+m2z2R6K+5ShHn4Ux0cnlS6HCwD/V0kpKqFCfsF
+6YR6K4MgH3X6xombGYH7MfFOEwcX1ek6RbpxBZlfzWb0ViFqsLukNIVaRd+ka7cz2EhFrbAKNkj
6h4+IcexYU6ujoXJOt8AXReNEu2FglE92MnvuozuO6JqXo5gPhz0RcO4mE6FnK8b70dWgSt8MQuc
b/7ohQsz70Wrudy8VJTLRykL5gHPKJYBKh/SQNEYRkxp4Wr4L9KiQQb+8QzDn+B5G9ajCWOhecpV
ZcfsqNQ66LHdA29YMDLL4sobuXoFk7N6se2zmJ1dt1OJ97jVVugqBXurzt79z+9gFLLGMNFEnExm
4FPYK/1Ci1U89UqiuJ4LHwvLi60mX/U6w9FtZHjY5fnlpeR2DKgDcKtYltjB7ljHCQKLKwqr/yrO
rmPwXZ8ANAwPjB9hSgDlDyGkWlE24mJEkQh3BhXcI1HFffkBlONzQ1j/C86bHQsc7OaJ3/CJBpn2
uFD5kWrY/XJsoOQGuQkKSahxCvyknsMR7H76paJV+wauwz8dTi7Pi3kB/zJHkU3Uhn5WYGVfmYxZ
9dk3iZuEu/tto3v1lM48gUJkZKe0GqUS6mpzijppn+wUfF6JjAsZnHjTx/mFZv8Td4/VT7ncj+LI
RHJYm3Z9+MkLqhQf8SvhrckOK/tAc+nrb6fZTPtTTQX6IHRK3PHLX3OQk+4EL8S1jEjVh4fHs51E
/mK1yz/LKRZg2KCYJBH2eR5E8Cqrk9g8QjOjb1TRa6pUX/LAVmLbgHhIIW98IEf8XzXEheZ1eBcW
YwbZ5ToW/rTSNS91y+M88BTnMrRixTcX18arpYnwTcDMGzxje8eIXq4Tf+27i76aktvyEHKDVD6p
YxmXJlJp8KZzk1mpHdrkh96CIWpPzZEWQDQmwOpnLg3rHIZ6a5FlMqJrYhLKkJyAciNjfJwEkZZe
OWZGMKi9eiXcatzFB6RZVE71FOqCJAEUIpQVoX3soRyAgvRl1gXvK109fGsM01w0h5Ro+pXbZ9Va
vpnUf+s2yjTXRBC5zgg0ljjVDJerp7s/s1AfdyspCHgjdUnMB2E+eTW8HlyNWRzttgyT9q+kjd07
Sc2NlqYjHmQaWb3KjFFrn9TmMO18s5oJ0zV+eVCs4pbfZzwBogxdt84u8gkqT3Aru0wBL0HnoG92
LMElTbA9EDZppG4IoGsEioGEVZxSQ3BUno22YRLEaL8nun6y5e0o8B1S2PRRSysBgjAQpZJqwe/o
BB5Rsz0ke3r26P5pjKZ/iIe3vsL3RgrvfxkYOb/hvV+KOGndRrQpp+N0ho6ysaaHqsW8/pt6QgBn
wI7BzPRblviM3c+q8szwrAyq+UVIT2r4J4WrPCGc1ahqCwCsy1liUmADXPHrgZrJZmW4drhhjS1I
aX4eASgzS+M0qTdIINsBPutEh9NnQlAxdm15QR6yAhXlzdQlWTaGeJm8lEn4OphbHhaHo2f/ZlvM
ZF4zZQG8YaLAIAfRNWKZsrXQCwrTnuUamz7zoxEYpSeyD3yXVMCNCIOeuD2j5+AKodiLXe4VjcGt
89goVyM9E6NWPTJNtW3ysklgdpTWjGQo4g0lp4F1N2nqYA3Hl6QvGDHCBsnB9IcHddTSmb8H59Bl
xnrWlqyEOzkmgdbWpYtyB7xRDMnFMZcnfT0Z+q9/D9SuRQUI4Fpy8UqOsKW3TZIZSWSZQMRFEYP9
P93bEZCWOzUDtbOWqQ59FE3mkiTJ8O8s17E+MK5PXOw+niYPuwpHA7sx5UXqRmjiFG4gVOKgj4Dt
3X4wXyl2tXUV1w/wMd9Rnq8qmM6H0wrAJl9zEr9/56Qx376xLz1+0tmVDkzkX2Fk2eOnKhiOH0hb
0H69vek91PIvCWYMqRBX/lww5d7H+9nWr/lK78SdEGWBbpdkpolY6bNWMh3f2pTFfpzUVpuOM9nP
ajSfb0H9biFmDFz9CuH8vtJI8e/iw7MZUGapum/zqUkXZVuwR4Q4ebylgm0WOGTKoRJqWFyYir+D
56+NleLX73ggP0PTk+Tfvk9srv3lgfQ4zIEGn1Rr3x+i/xjpBBjw1jiiURObBUxpjMKH7TeEyPHr
pk/0pGChyhz/Z7I+KTt2PYv7WEce5wxpJmors+gE3qotpBaaHrDVOmtqXhr6hInhQwU1hJXAOvmf
gVNYBy7c0LZG76i51ZkWPNnvsyaptDzMtvqAoIAVxnMk08Iq4YSjnqua9Z8hiWnO93wRs19cOdNX
NVmN2XMyVeXvltjaJHb/TCSfwAIGEbc817x51GI0QsyJp6fk5M2hhuIwivBkHs+jamCm9ZsWexHO
+Cs6Xz4VCa8derbBP/j8oEZ2f1Kx8xl9tCoNRFkEQOvCaJ+eb9Fy0kA4FqNN5aADqy6hX7MiMYVP
aFPQPTnXQv7jzq2H45DrjMeEKIdGs96Czom/WtjfW4NTgEfCY7Mqb+/QCOJpvRFnW+zC9yZswXBA
v6FlS/GyWua3wvSRNRQIJUlwN7oTkKpoyTE5Da4MWMUEOtU4mEz+wQ73koozMbNBKkBwBQN5dIDz
/3ESFUOjIM4aOhEiB2YnAzZHTfOlBwJMmLyYia0jK9ilPsjkxbeyBC8wYFEXdoIpTgpyMf/WMO2t
Vsj21JrZeXEY8xaTRxC09LzvBwHomS5UV8Tgd9tKsnHQChViDrN06q/gGPpUsortkhIZR4zOp9bS
1cggKfO8fyZnsS76ZCLlUQcoa6ARStnBFAHUuR2lG2FOgMRi/0mkv5qH57l8aarD5VLOOW2/8ouJ
t2ffW1TzjdvLBzIwMXOrV+6VT2mf9lNat2nj3VapT4lnVJojqQBEsYJzuZyNRLK3BT1FGGrXxPwA
nQyIphRQavhXSIvgtINxStd4y0D+3MBjqgHUf8Xds6HKbO7PDZYwhkTf0lOrUAwKA4Vu06AcBmvQ
ZICmxMDOIlg91rQdcZPPLvpMr1JAL2ZXD0oQM1blfl+QjIO3MAlfq/u3IUz7dQtk9BS8umiIU0pJ
4Irg4lbkEzcXkALNNOA9A1BPJF3KcTc2wvsURp1aHdkMY7ccZDX5B+YiJAqHPZqTJKt/gidYu0KF
0dh816Zye38ptsM2WFty7ogVrNDA50FHIz356Yp6BAyIs0h93EcvmZeKc8JsW0MmuqVWLb6HcYRH
OUQN8fwC1Wf4VH16KhRn0EjfikflPLBgfEZJD9YEb4SUXfykBU6uVjmxonDskQLXf+LY81B2++4e
t3gEzau643dKPTaVikr2NOSmnNct/GTIbMPWsgAHbkyeA24hjyOo+4jE+hbrDkXMqRl+aBqVKDIb
h0CoWlM2T+m0O2ySYjhIiESYZ6el+UNoSbP/pqB2jijaLzAORM8FHlXKD7HRtkPysf1tguUiMndm
3b1rQjoR0YvY0yA99KttzKY2Mal86qLKXryi7UtMBTM62iFTBC7tbDCiICyf+V41IGFBlAlOCzXu
swPzpLcsFYDYUw3Q7j4wJpv5731Z6gJjC1+OBHsGKhd/O56L94QvZORoi2Ci93kTcvB5TJyxQ/xV
87+InxXckO64rLHqefIhj/SzI/IRAWcLwwu+tBHjYVqAigx7upbDT9EimP9SZkU8Q4ew7dDXmJRY
++2Wuii+WfLrK7cD8U5Z2PdUqo6E1P0617EeldLRnF+5HIXvBu9czYy0b194oxSkAXo8eJtHxauQ
d5+DmHS9San8PVH+Ump4TVgOmnhdHf76QGkuSOU6J5Pixze+scLLAvjLJKB3iZ0tZfFOrV7DWF7x
xZnvp8IYaocyAuX0v04LwJMyc3FzrGgxWlQ+QRQpsvU73mc1Ah7B9v1VEVgcWzQNkY73FKFqCuVP
ubvrbtNcKA/CDbBzBKpUgkDUq8/Xm/k4fMfyBQTMBIqinTxNCcEy5RJsmYDv7PPGpiwuRiNFhbzV
zB1xTLNmHplRZdWTqcBrmTftNRqtoJ3T0GnPfRvyaCsC/Ux0SrSrTdDwAucJx7Nhe6iWHkYLwreU
XnWA040x0P706VbVKdtRtSj2RiXegCFcD1oBvq6T6eMDZ/qz016HKrGOouowQ6jgc8C6n4PjQj+G
5/rsHj16YMn46/1JflqcLp5OHj1Dm5aFMBV16q7a6Ke5GXiNj+rPMmUd10Hr4JQDbAn24tlmaWZR
VXUUaDneCsDjfHXtWcolWiI8UkclN2UA5Ckb2T+MjFNo+yVm8CjvYTAOojBz/NWEiL/7LC/C3sVI
x/WQ0VAAkt8WA1zypoD2saX6Wtgdbv5fK/tBFF872rg5pLMwC1MTrWXuKX/XydBkmnLh3wmjPMQs
0+UOyNoZv7BdjQjYz2RnpIv/I4ZAPuNlUCoJwQLp374jE9TregyNSwqEBjBSDmkBYYRg5gqnzuQS
hoGtQE8DFn6EyQEmfUc10Rm1Q7vT1MGenuLPwuWDg1N2lmdJybWWOYb0H7lDI9VemLAAEJmmoyCG
DS/NQjnSshE7UJN0+ztRI58uAd1hydww3l6m7w+0/WnZr5xS56mKiJxgDuKw+3C20bqAwqjdZ+tt
SUl3GZ8rtSCKuRWI0NddnT0XP502bUsERzaIw1JT8g4ABpWWiFCWEjPiJYqo1WGRLSFmiPS03ACU
plV9v5wdrk3QVtx9OVavVG6mzL28uAg8P1TrrZ9bDdxb8FBlNAJ3j2FsdA+Aa+KRAg4b3x5n8JbW
uV9OyhZVF/0zIH9HeboL5ks1jjKkbPiR3EQCaBVQiHNSVzAUVXSLOwOzY6Pm8qj3nhH269DN/zKd
XoazMapb/V208YgcyGQD4FkSSyGVyYwrAY9wu0d4JIlY/SJAnmbfi0/U+vb4AZaFKV2XWPrQKtGl
iYsbxuna6bTDGFfW9gUbwO6c2bvGQ0pqHji2fCJR/snvQmpkqXi53zWwX980fsmHYwH7FUxDK9D2
3853KTADWVIkh9Kc47xCCruMpigL3WNvKb5pC5RSn81WJw0IaGpMSfwTn9uXv7Sp4aFqZi/lWxKF
xaooJu0MRppQFScMYhbc36vmLBJRFBIJAfKNCuW3vY/yr1shDWijFLB83649wGPzD9N13z7tRG48
4xOIc9LSsp/HWGV67yYp7IBN8uitvCamIkheSUnKbjdAO5TeB9ENSuf2ZUkhr1smNvsaGSB8Ry1m
Ek+ibwX454RBDRHw30bse1K2A8qT/E/vIrUJBkSu9Rn1isMMRh1/D9+Sxt7naBZrUHfuraGlzRuB
wB5wYXBj401g0RthRyOlt0fi8WwAZtcdjo2VJkVxifCbw6nSwlyJjwMf8kYovw/Lct2UglLyTuFa
K6BPO5TWsJ+toZuIJYZgNYOoXuUUiJUjZsHLMVrYCjaOocIrqf8j3ovS0S2qO9Q6JfanU79E4uBe
zhKBG07APABRturaicmwFs8c8jJNDbIOd4jNEHiDC8QnRmszMmVsX5g8//HwdYBfCaeTivzzibDX
4qHFFsGYF0mTm2XW3J5VipqMbt9NiujOH/42WzXjG5vNgESx6PCA/jQsrB7y/LsR8M6Se0lcII8c
tw7m3lzMun1gvrSHGjawKcHMQ8kehRSUVv+zI82YUrpinP9d+e4ffotEYN6Zw5CbyciUTpr0retD
0Tqv68iC66zmaFRksqIttK+gBLOKyrfcSDhpCNO6qPoxQgjEnfE3mFGq9fNAWdi5SoIoR0sBL7GC
nucySNJsfjnEv/Ko32+ZybgTYW3Zh+E78S43GMA0s0cYlYDl0CEl8NJO+asoU6lQj5MVJsxZ217m
Te+M2nqhghae+o55q7y3sa2lB03++DKmK/6Dh6zgDGSVd+kDz9tCCRheOrmAG6Req/Jn+QMD22RN
A6GdUtbm83PGQHatHPU2NgQovqtE7WBrGMeBcYGfFohwRdwSnrf/DfqRC6f8Tsa/GQ5tpqLP32kH
2ihPkmF1D5vGRmprR+zqeh0vJDHV+kzdGxew5LmMwdkTtZsi3eogTICeCpA64QhWtpTMKnrMyCyX
eWJG2ndnlArKC1hjakeSc1GdOr2xBdlF6cVAuRknk+yvGz2o4Vb1G4B5qAo0v3PNw/3GT1DJ8Qx4
m7Co07O3Qvz4pQSf4Y095JI68O4QUpP0Ho+ZVd6d06aP+q5Qb+rjUxK38b/kkcyfjpMtN7aetzTp
sXAypnkztWF7/F5zlqLiE96NLChh9hpnLWHM66uamTPnu4a+ljgKYCsq31Y6NIjSrHD7VtCMkKv9
OgxGPItGYlSRw6xeiargJFil6YsitRdQz2bTWISTzRjiw4+Szs6EpdqVYtSwhcWUhMvtd39Z7xZO
IyMC2Mc+4OM74q/2zTAj4Y7kSDf1hKHgyKgrq0K+AhBv5G+mdcIlQwGJg9J79D+T6Qa3YWnukl1N
YLFF9Dx/XEIVxr9o6+JBwDrjfaf63vEss5mY4VsVRQlNRcNocaOcLxDeNgH+H9QWKOFA31lnRsvH
8Dw3HxCPXNvRmu+GojB/kzUdas5KdzPYsKJ+Jts+gORy7xGUK+B/eQMnmiTgSQkJ596q/LDscpKM
2s2K4S9Gu1yaiZsKY5mSzsK0Sy6TjRphMTOYbKiupKmDdweN7djEbX1rRIoyCXwSW217C1mkGgYp
aFL2uVwvjeRdGalA5tijAaRNPRvJ7AEYeRaFv3m1LrAPxCILqlVsdwu2iPNKjY/sOAI3UpqOl6iK
NpGc81NHwSMmD9nR2VbDu3XBY8p47uXC1FPzD6sc7GDNymUK+Dofn5XE6kASle1XuoDpA1o+7XjT
IJOYRrY1q/bNTlIc4lJMuDY/tJlV7VPAHwicmUe0FBlCF/P3UqKxyvwQqAh9IccjTNAlf+4Jkooo
5yNYkC7w9IAnIkmAkM2IL+DAp+vxIGPPpYIU7cp9hLxkOybOI8VS1mEOUXHK+4NAKWzYasfFqNfm
IsEwN1vnFI7MrEMFFj06LwTOengDFIIeg+rqbPb65CwGSxl5b3jQU/V57bLpeYrBoi9oXCTWVauZ
VbglLlHt1nbmVCwHhw5HvCsYfiW+HhDX7oNUnXs+Br5mowBsPK2KoXyZ7GNYl7GorPUynxKY1EDA
nLVjCDvuMp5xjmf569ziysbj9IN6+TSCUKw+SVqrsVFJslgeoIZmdJ7FRWSrQtsP9I1YL9Qjo1DK
YO8tmD0O0cowO7GrkqnFX2DZsB7phEIe0KtNTOPaQz+BUUWZnHVsy4LmxPSQ6Ct+U/JwCcsveQzj
rP4gqe5KVc1BHhSrc49Ywu/9GNUvvKAJ4EuiVEWiPkRXs8QOcPWjbPN+Z9a7QPmugGfelwHr0vgM
FtkWtikqLlaXPTjbCkVve6xjkBU8VPoIzACJrdcYe8l6RBs1yWIlN176/suAWsZfB0iPj4kabWtq
7nzYJ4R2/Wejjbc2xack2MDu2sMvv3l+agOY9732MwrqrL0cdLE3+hV4CFbppaE7wdRhp9K6hP0L
vA7+P1bcK2RHu35wRCP4ubiEsfFd0G1JPCXlTi8OOy1hFw+qNLDmb+/SZ45hn9e37pplpxt0sSwb
3KJkH5tkNPuDD++Q/KBUjYB2iM3rFPTi68PjzPLe3JqFGsWEVb7fO2aGqlKj8t7jQhmwCBtMv3IQ
M4RJOuZE4hf+mE1PDYPfTbqslh0PHZ9xPNnZC68LCy5L6EnFTYaZnGJCxwa/0j/cWjC/g8R3ORXH
J6rP/CjL7JQF2cltPOnDzGPIykcXw+7MHctll2euFRYuEw13tEdJlxGpLjLEdkYZHlJmCzALDOWR
P08gpHTbZr+sMoKVZHmtQpRw7RNuS9u1J1zhjaQmWeF7vY+uZQYp+wK+4NqAv0yOGljmKvnDHA3f
nRBbYDfERn9TPnwQAtBH6DqUAFa0kXPGDSbb1NPllL04kWGg047wowShcVQp8qKtxOgY2R2oToLo
qYxqnOOBBpkhBH9CqyuEqB5RDDc29mK2hcFeI9ugft9JWGOHbDK1Mt1lSYjF4ISXhcrnvmM9gYhZ
XslbqN2AuqoyxJ73zNN1rFdxFe9lR4ELTKIBYV1eoDAWjs0ZmBVpYU0gg3+xyeRFTOJ1NipNTt6R
K1Nc+0mFbArRV23qkjGNyMwDPITpcYK46+yZtyXS4zXmZJTTY3Baf4jrH0ZKPrPuwtrEW7SaYcN0
GuRhNIxc1wEgjlWO6O/QYtLKxg+xquT244CLiCsa3g0KwOe1WIfbu/lfszvdG+QLQB6pq/r5HH+y
Yxnkv56rY/ydmen7DXoBObIrPsB5iHMvoyvtpLaxIBJLUGkCDkzRkJNyGubA8g0WoCTbo6l10yeA
1SfyD7kK5Z3A3ycU6Jei/uCkOPmK33kyT7Iq4VBfazxk7vNZy7F7uQbfyBN3l840sm2zaLK5bRnE
Xy6CyC7m+e8N7e8TUbI/EduBqbr2RNlFfzd+l6hUIT7bgGsarafbH9mPvzJwqHUVlSuBDE/HbXKx
IEV7LOuGMrIJjc0pQT4AiJAaPoYkndsb3fXoSvP0XznxqZa6p+MFx3TVvRghr5zRHxXAoxgp8Fbn
MhaaVVuqQImzVrQ5utP+hAdmwDJzn15FyBEXCWrPmYVp7IvWqGrGeBFMnTBoKp31TtDfgMNnIkKi
B6NG+OAsW4kn0+JsJw8KFJwTbCVNjfxOnzIdsMtwRtql+fNHva0RptaNQyYty56YbJ++v7Fk5t7u
i/XouBwFBqZkjkwGzgP1HMjQB9lVdJhAcUaWJKyRsUDdXuPKyWaQb8iThy96scscUsHB/7zx8VNh
2/03V8zKfJ0h7KOAYC80GUa3Z9ImneTqmdC3PSXtjKD0s4K2J0jChhpzcmPZyHSQF3PNZ/euRxNc
bxdYFvWmyvm62QJ6QX30K06qTrkDnRmYsKh2F/j+hIeyjrEQ7b8n6w4s5lMf8EETjttXpTS+vNCy
yLPf5InJhi1ArxtFm/ijmqe1+01fyjGvWY4AZHfFCCgs30yDx5qTFf1rifdHHXrTQ7ftLacGEPY+
PY11IG+HZiNjO6nJf3KrRh7RIRXC5oWdwTnBqrof4cI/sjU4Ci4siulyiTF+tv9+LwCBWsuZR17x
Q1d2jzCRQpxZWsiU9hz0jCjRojkbnVfllt36xrGdv16o7yHcSi/EuuLh/TrVJSY0Sajvtkv80HP4
bz7xyCVhN60sXq66tpoCUnwLIoiQi/ZD9wfAxGBMh2tinaMX5/tCFhuNTGvCqe6qvSG2VzYQ2sRk
hNogLDLgozApg3BjR7WN9GE6tiHVgBe/t+vJKneYSQql0cKD3i+Oz9YXAavLAKdQz0wBdHIl/zQ1
kixofS7JDBDqmOh35PPGsXGWVWfBMJGXpT2twO8emIRMULeFbDqSkg1/Y4z7ICRH0ZPf6uP/XRtX
PCh/KELsRGitmk99jw//Ztk4YmuY+9eDvxKwP6ceqG9TL8pGXe6cDMG56ZlWTtRa8RKcjkZDaSu+
vMtwvDP34/ePj+qBf0T2hb3psYZid8oU7+PFj3ruINFX73t5rkfNSji35v3X17bduSKtj01f9Opq
yljenEfWkuZabYWeAXgS2gjByA8zhbl+HDVOxmHFGePJ72jp/8UX/kZWmOyenH1UlMt9OatUcEMp
ldYPW6aoQTZG/RBPWhTaKRkQ9g+4FcOIv9BtN3KC8F/aFj5dM+2pQl20+RomFmNs/5Jh/DF9vBo+
5HnHK8M/QMzTY0SkAirolawukbU7733UKXzODWWqCBlo0Nj5o3tvgfWz8ng0oQ1d9IpZoL3OkOA/
e0v8SgX6xgqg17E5pR4pLxfI8jQiEcHPDzii/vNV+3jjGiHqp4s6iZ2idaju+z+gtny45EwmrRq6
eO1pUEHenxFlGEd/sIYjj9zEs/PzHlpto+mOfbW9LRgahHhR27x7yBHUNbfN109DO5qcKAI0TfXo
TWfvn8kQyiqaOXoSTrJIcJaVC03hjrq57YPbU72gB8fCjmtE57Ea00thUeWqFivpv4UM3eagvmqQ
5DNZEdiBHrM+YZiqgPfJGEtSHbFgvHhJkkwfSl6E8V1hZqqQNVgPFGU+Crx0r2/5dElJ+CouCOFz
MXb/d7tMgV5Nm3F3/i0W/fR6fMdrPysO+3VL0LEwX0oDwNLU12ZZXNZ3l3XIiEu0IYEII+27awqF
h4ZO04QbS6yI08syjcD0JEcfS1UC3v3mIrNW70H35cl0p9HIfZpk5AqeuA7ovflcscHHRb+6BwCl
QmmrgPLAuMntrB306wsqYWHAeBOREHUB7vj4UlktRawxas40i0mE8c//ap3SmxkzQt4lWdWVBMkp
HBQAZ5oWiRMx+OLOF5d40qOyYvIlb9DcsdZ6skV2rWsrW3UXUX+SqT/9H/VGVCTwfDcXn652JcKB
if17XcQyssBPd3fpg8puXBJG/Cyt5AK8C1qWcTcSnIeD28sqCnsAfE+YHBMw8En5p0F/QRBPUsHy
Mn1SM50LsDFj6LCnYmBG65bDFK9HtN/S89dfYCRLcI2M4r6XMHSSqiWLCyHI8CE4X42rvcZo8D1D
cJAk7Bnx5cMhXR7vA9HTG6ryMTmkE2TLgqHe7qGjUQwzsf8glniNQWHI4kJlz09b7zpcghBSeZ3y
z3nUk2ZcrFkMAbbaoxFfKjuyMTSVfHEdbLczf7fOzz57QOKFnQBZL40HqFRhW9HDNlxv/KnM0zTS
BRQH8Ad9WAVxCuw6ss9di57niY0ag+MruZCn8ed5q6rXBO/tO871eiFKuDnUQeLK1IcxKxdTZ+mi
KuFfLQaZ04hKVBzFEEls+d3o/Q5o3J7D5F6xrPNoWw1iwNxaAXeF8C3cgSA86x0YCxK8KhLt9FCB
hl3cW0Qq+FNFjOecx+OvhKh3BsKBS5YNTLwUKylqAW7kCbHgkNZRk9KHzyu4ufVkB/3RYuifmy7/
BQtfxLjx8O1I7gecBQS3K25nqMr0O7qB8x8IlrL/HW45iSY1nLthTprQ8hg5n15BR5Mlc6K0k6pI
qQQj9hn4GfWqCaYEsK/MImJwKSLsXjLR5B8LMXMEsvddb43/c0IWJNu11Dq0SM59MblJq/dMIIkO
GlR+VaYMJhao8Cj4nVLcngG5VaLmh7uzNE/Bihzoa9MbRg/ybWnMCQOjoEsRLYBBenErbYZ7C3np
dvbN0dF4LjpHvBKPAVQiW5xjb7owNEKfOHWpV/87KjYBvsfiGos7K8l1X4rcpIzj+rxWOnfW+1vt
vcM5sa2ifnCxleLJqb4jWCkHgxo7t9EL77bdlWAIeGL0e4MjQ3sySEpQ758zES16RkkF5yh2aOmS
RPR18ZtBPRgLKRPX52QM0IV94YniRQwrQ2euez038NlKR1UP9R3bFdw5zKANU7rhbL9iX+PBDncC
DVaH8TV/Jkz7bffabxcyhYNYU+c8HXvQyb8IDAFUnfYFIRun1cJGWlH69P34waeps+423xXzg4lU
ausZbohce3Yl3hATu7iHu/WLKq7Btg0kfd9PUPvR4shE269hqk7BMPVQXwxZTVAeQyJSjb/4biTW
m3/dq/EAd3XTiWfQuwMNLWBzIukEyeLA6tEAvnmY0E+jwLy/vbbWXqDlL4tk+4LBTQmpKd5gQj7I
SiALS5QalNI+CH1t4T0Q5CiWrbF1Yful5Y3vHWFyUCcAQAzbADjfqpTaiwM4mo6EYzbIyQ/+7lmk
ab8pWlXPB7mhKZ5uzObJBd7qjvGPL9P1gIqnpZ+BT/O6e6MNzUpG49sAnmReX9Axl2eQWIlncdeo
hrUlby5RVFhBjC+RxI06BFpCmPYDMTIOY9iAI6n6ZQe3ZE6fF3tUcSnRV0+4a0hldoNED3yoQsWn
xnXslaC6EDHiADZxqGhVRqaMI2NO+YOMH8W0cswQP+rGs3mwXTkVUnuD6AHHcCxO5Nzs9e3PJPjv
MnTuDr+TzwGcdLpQPN/Wx+5DqIJODaYj1ixhdfs9iULu4EaAE/5F6Dr3fQQrtll6Kp0T0OqAhf07
cz3WgDScouBzh5EcoFw98QMoVnkwkDfai+ADfDt9ex45rjM8Ja8A/PZ7b9smjLGq+Masna8mh2jG
WMa2UiajO4eT+rhrxOf09pfjx79leiPzXvGRqxwj/FHpq0aMptCai9fvR1R4GPRUVjRAIwI51JaV
kp1f/7mgZ3HRw+eFj5JCqREOlLljhhVp0vh7yJJ8JGUp7LJ1/9Y+I7XU6/72Fyw+F0yGajW7+Vz3
sqWrDlT1YFB5tNBPGNCWD0VXTJiqYUIvWt3+n93NLagCWUftBx8Zu1lUJI6r23A4gEVVaytH0vCk
FDA3gxsUHLnWzFjdxGNwmZfjmiVcKJV5M5xeZynIFOkqGimyVeGDawzLrzG1NRDT0waBC9RjDRs4
kqP+7Ql0zk7YR9ySXeF9jgSCbQluQ8ic9YUZlxYYBSQWWHp1MtF3Al/zdhK0ugUpqprmZSMa+oJo
a16CGObDaupYrwW1v73xg7QOQKpfHv9G6MMoc+tK+783Zw9khmRaUer/D+3noZl9YvO4tBMGzq6T
ktf3LjN2IXbUVtZrT4Z3c2LlSwk5dLwzKo8Mi59IsEphkVyBpMTbFM3HSz5twK8Q6BDpFOoFnKzt
cesGZUbwpxCB9akTuAw4d3wrkq17D5YP0vQCDzbjxuK0G33A3u1765vBmLk7FRH/abJZUZovEnY+
Fsf8NbNHa+RZEMo7kobcmN/AWr975+5kcf26HWxtXs/yt3073JqmE7jF/E7nYR0OUbVoAc4awUm3
Exbi52bat7Jwky1A3FP4gYSJsc++0ypZ/DgeA9jMOsVnu8C4pPFoHKfsWmGRcI9jUXllSL5zKvo6
iDHyM4z8GINUxEg8N8x/eV8T4/hwFPIwSGUuDf9d8nGOxDXs4BRM70DtHM6SCTAqGSMQBbWQegHI
VtYmpwVL2J3qXNJ5Ml5g8JxLEkygZloBzovk/lu2DnDaqK/JB4hmIMt4IhXDGLOg3R5lNXETLwo+
OrhmtXc7MQaeg+35DAMS13/gnH9Hlvso7jIi3ASbXhXV3qudlVnPobYuJLniuv/wW58BblseJJAG
nLCGgw6+JZbtELfHfHSHs2+MTc3GRAEX79Rp2B9xsZVfJzwGz+YY7fR/I/2xWW9Jmq32wzM8nx09
WcSx/JZtw58NNqzB2MQN00hMKdgXjnrrUKuTIMKfMRIGjV/FsAFmpZSjfFqi6Ld6S7voyJDUo5Ej
iSze1ejhDouJ2auSLkiz2pv9m08nT97bEUX76kIATPef6gX+T1H15TdvyyN2Jt0PCQn2nQZ/EJ4a
hbsPgGB4CmV6tE1f0sDzxl//uw8joKE8DPQndQUoX/RJ80auztmXpuybY2N/cmbzFDWIS+Lf53cb
fbynEqvsLNFVYHgOIj3uniTxzpH/3m+7Kf0l5MQOVZVhw3cjZHEjT4fTEo10RbwmDsFmyOGAPngG
gX+rX5G5YAbgoJiClhGH+utu7Nm+2SIK3rAL/hkSrigN3yz6siOJmw7axpSEv5KITawg3Hexqtaq
7B21W1J6zx0qiiy7qUjBjZ1rREHlJYaKp7pnmNOWzROOa0uVYWBYRZT3ajC5ADvkpudKl9hF576W
+cnm4w1C3Lft0ng08l/RZ32jP0gaUKYrCLaw+iMSxvXuUVPM3+jzzCtpFJB1guGYjhdI1EpBKKIG
2RJaZ95gQL8DMWRHRJ6FrKr0OP9zNJzxDkS14matziFy0+fkUkW2PlEHqRRiKP9uqmBbTT2fU1vR
TxSnToiHXM9VjjDgVZuUO9pfcPUfLIGdO8RidCSMKUShEe2yXfBaFA2rioXj+QoyttZfONcbNVMq
AAQFT/RC2Zs3dS55v7uSDQ4LqN0InAGoovJqCC+DbnqpQyB8BGt+NwA1LqXly8Wa2TqfSrjW2rci
mBqv75mKtgvWWxJXU7Xms6AOLRdctLsc3H+MoQdRj0cj9b9SSPNF1zKf5bWE91MUr4B1X9xnetMP
Jt+sWn3ZK6qPMAmV8Uy0dSaF/pyPOwISD6K5aceZv4vf8t/KVVjZb+/BetWq+633TKC3TH0OJTFT
uZ5xNak+wbTXewfvJtrQi4IxLD2UhXg24d43r5OCFtEbShYf4fu+GHjMz0nyIlB3qDTnnT2kglGU
TYSW3G9xGlU3EuDAJQwVnP7tuyxhviI+mKv4reBAqzwgz/qyd7lsjb/QK7WkYCeAqo9OIMklN3lQ
ZRPch/7UCb1bfq7uZ3pmOhrawq6XFTL+eLwv5Zd5SUeI2QXodNE2KGmCB7EHKFckdyFPHnOwYOAR
sw0zDXyrWDafJzTEC60mIi6dvvL1bA8V7jQBflBmbeFggO6VVBX23+MSt5VN+AKViW3FoqeFY86P
6HLTkXAb4xpfBT8egq7y9fuP5uWfZ4eRLKLO9FlCUANxhR38it+VZgRe5jCqO71bXXhYzlYqBzUo
6rg5hDDzMcMfTMJzpM3YqdRJmajgvMbBjr7cc9hZ7CWGpHPuUWgUkV95r+1aVykDL6QyCx3g1zFg
UUln3GW+fim2T7wZ5NMHdvv4gfRSpMCBuuW/oB8EeTcwcuTIWX6wMg+RkbIsxAIAJ66mo/+WmWpG
aeQhqgrzPJnFvOHBlfrQLNPZDKnMuzIaJr5MW3EMCupVLbW+5PqcL6bKRr4s2ygtquCmNVqJxt8W
Yv1Zz4j0j/3xH43R1qI5o4MHAVAoDlzanWHkSKbT55P0I58WF0CUAtNIWm+kXaC9qXwTZTxY19SC
+O+ZaciHcMcPI3KJ91DrRvr88gb05YQ+tEnrMMlvoCQ2n/5D9zVvJbPHHXEzlP+W84cID/L4qng6
ncrXOYhD+uDPnwXGLqZwGvO49xb7nUzVcgySZhJcbt3USTyRij6zG+oRV2awl+KlcXFDwOLZCXBV
hwfUsAU4HRoEapDt9hT9BEVq1qV9FMEyvegBaeM2rfxbrJOTtVAXHbFAh2Yd2CHTMSyromLSrAZO
z7rFTIlPl/oD8zWfzB3vPXdoakFciqrEONp0HvME1gEuVVYCznb5FN/z6LL1bJF7jlcoX5TXkup5
mEthFhJwAs8o0/n0onBtybClr4ycRHo0s+SyMZi5noaXsezEk8yetwBzgI3A5/gIJ4FnrMGxQo6L
YvC/XBqafDGCeAzU07lz1TliTPc4kgzxs6VaSwr3kRmlNdTU1g+/cEkFKzJ/z/rExPwAY8qk6l4M
axqddXtlVACgRherSi0Ctd33xPeA3gcihAPbH6QtiyRiXY8lauP0cFoVKZtjneO9e7MyGEF8bLdo
42Lf7N8BPW7VGEHC/yC9GbcKiq6FHhVPbX8vObZe4UZTS9Ql8NUh/k7Y2ap2Lh0wExNpJ1X6NJ11
cr4zZwKxyGXj70PK1Mvr2kLCU+/Nzy21vacSfz6dJ+0JWmVXIsWtoYtEsSGaT7zl0SkAW+e8Wup6
i7VENRDXi60ayECn9Hb/bbOcLgm9r/1LCWkQL8iDqmw5L5zvWuIMB46mgqQuTeKcQQK14lJP4qhs
IQAYiDgnndd9pJrOV8LU6MyVTY64idIvejI53Na04J1m8JlZRjGEZzUhxkcaKvV6+czakGzlrZoo
YyoQHE7g9u27QHZvTQkhPIDHjHzMrHIJl8t1IKVpp/502v348eF3zPr08QHsJ8mE8VlLebZ7S79D
UDXXVqo4a3bPghPvXNrK+9bI3A2t/AjC3b8cz+Noayyai2JtB2XAEF2ZLezVaaxXrZ6HHKhSWWEG
vUyekLKAY+G5DHpwJR3KKCsZylajaxB2oG96o5Jf/B8HYBpA2bgaeJWCqmP0hNPnutycwoc6kXFx
19STO6GAd1nAS1YGAbOpF/6kuS01DmxgFpRKfMIFSCgGpzLdSONi0Cy0ZsNumULP+ab4eNXlc/YF
vaqfC5gUax2q8B6F1G3C7nXVHEnQYHy2+gr3CdW+GMKAdHos+JE8rrYmggSiQyUDYbdZx3vygau+
MrLaC4sggk5SAT9xb3iLFvzceOAQG99xpCfenEBuv+fdbgTefv+Krfggps9mlq83C0z2olwC0uUe
3gUQ2O2izkw/bnSjirJ7jM70EoAuIxUIDcdzoR9WnmidbmjYK3JkAtHYXMhO3eW78NQBaReTaW2V
2dfDrjWp5g+P1qRWsdZZ1UzHQEsot6h9IAtUMVaJHXOrLrL7fcpXnXp9MuupzEi0ezQozbgN7Nuw
dhfnthE5CZWQM+oibLCMID2muoJAuQuUH1MWsWrlUxbjnl4gjHhJGF88AT7G9srFfRjh/Xh1tfKH
Q69948aYpT7jO7U0HP78xupkwlYGTwNtHAsNYgqzJKBAaWySbDgH0fOFwQ0OyM1gzhUsm/sEOcym
FnCIX1Yi7oKJLHjQ+n/XussyODpadThubrFw0nFZ+F39uhzmxc+379zvKv4urMreF4AQCUuleBfX
zt0M10oL/aoBEiCX6wA5xIFZiC3KkJWhbHAFAd/muL/gslE6+Pq71IY2PO+m8Ja00lE4FxmsJR+f
uoOrq6otYYT5QBOFiDbhHrMHwD03OOr9JrJJo7mP+ONAsOPVqD9twz2bnpf6UE3/w4GVeP6NEzSf
Mi+9AKVQ7CYmmNT332xSsf0usS4RJb9tMppYFzPBtMlIB1AA4BypsZ6SsQyh/92Dw19NJDIiN42s
I8eXtHiCibb0ab1AvGtKunZw5GwzyR9TPhFaHj83j9tCmCZxfkY1HWcIpNIq0JDwqBYb3xqwOYzj
Er6c7NfxFSGNNTPOIkvpOkKp/eeScf3A9Excb1AgiDoeO6fWLpJUIftiaKNWMekXRrrW5STv9s5c
ZBNgBVy5NclrqmnziPZRbORzJ6yFRPMSEXDV+KNjuMWvu92eqb3ZqT+8h1hhVEwAC25DG3kcT6G5
NpkJIz31pc5SN1jzw+yOpm7qTPWRc0+F/BvPuGX4fGTLLfuylteQMlIZEClZMQ6UGC3s8XhR3wEy
3MecjUTZr1wsoOBfWyS6oCNH4NprvQZBxvuiD/eys8gaXnBsMFvLZ1E8d4XyjTG8vM+dz77+DCm1
pJzV7ZFEsE5VRJWfAGcNBForFi0UTvreVTcUgPhaYJT1gK664J72Om5DCcUh1ksC32Zu6eRqXp7o
4oSeTeo90dhgiHbqGRcctbgvUdtItcLYugKNmXPITos56dIGW6gj80mpIggST+p79RRfaRZ7LKZb
yJbCRKL+LmW9mheVSTy+nVkk3pz57+R+lOyPApht5iWozRCnUH8rt1aTVDsXj31PzkikaWBwHXQU
P3xNRV5MZtqSVIiN6qb91Ey4wURb8fYn34C6QHP5EZvjTH81oCSU44McqbYnjBWsDU7XUsO60gik
fA8tpyYYykB/uSKhHsOQHd3Q5jxkgjoFq9F5CIvqfnLJPnQZSpaEXucEzhJT1wr+ydc6Xu/jTw9G
B3TLlpw07fLSnKnXcZXcwzajhhVEk838GqQGaCmMBDOSQwEVJN+0QEePhAwTtuHpyXN2X0Z1BHCW
SY8o1TuJW0ZJT5/DctSL1YvSIZCYdulQXhS5jxdNeJxQyd3EFxwVGHUMvtbmddGjcyoJG/o3wsiQ
8MQWgnwYabO51BefEhJjck+nZxEfDLJFRqVvrcz5yAooEcjGhvB0DxF5asSuvwSJBniGMTaoYfdp
kLR3JBAMSg+7/Q4vqELB0XO4wkOLa4ecnJ+i0+WgpAKZJhCoY4RitCu8ZEyXQhG25PYnNodKZ1J0
A2nwJh0zhH/A5RbM1Dn3lQOsfGjUWYXTfLTtiGpmuUVd78tWbA7ixbjniy7Euha4c5S10jm+W+Cf
gxGG1c8SVfwld84kQs0QmtxwNtcCu9eFB6A3yWNJU9uBucLrF/fzqKSsILSNiElGfwzIWFl29hOM
c5H6Ykgj6r3KKyj89oJxPsHMhrjPID/6sgcEidubUUQyXntflGy5hJDyNRkPlncn6zFbg7iX+/Y0
bKxB1Rr1gK8G7ckhR54UyIq3z9rmBIcA2fCrohRbwUYLQ7ZZlRDtaAv9NopgeoOY8DGHJfO0KK3K
rMyjUjaAWG/kQo+5kWhj+iDY5NouKiAnG4noK/DMhBGiiSi1w/8LK9yBteCVj2WEXl3iJQ8gCHD4
JRFM219YrFj5czd+7VoI6CxGqkviW8m6/ptK9iRlVS003cL8KJWs5Koz60g5ouLpYiiqBJd6YaNU
vaT0luZZd1yICbX6ufrxFC0cgppOq5Ni9cw8BerVZ5u0ufnNvcoc1Tc5kGqwbZ12a6a6h8yG6pkC
+aJS6LTT8St62FG99HI8NtFFiUCQiSV1tJXimDc8fR+gaudVSPj2uw19mBQhFnFZvK0BMbpnObKp
vApEjqfgB0FxMqjWSsDFpG9tgYzVElhVJvL/M0vCE/E2XrWRWLarb5WMRKnNDjqm0kyFBHuEYfx+
C8keC19BkkE4e5iunYTgaFc4QMDV6sTbtrGo2VbV+ZOnJK5220DVyTuvQ0nXs8NBd5qHDEPvcwhd
9AmXSoPRUfDElhEH4HOUDrEF2jvQ/hPJFzaTp33ZyditADTU8l4KYT+ZxkBfgWfsrmurkQJdfo8N
C17nDeOjZIMskcODCvnoEvV39eaqEKeluJzTdFq2s4M/jw9No+jao+1P3dowuAguR5RlxzJ4rqO/
4ZVJs73RFhXoTj5Mc2plveQl2OOVLomOGEz7NWcEahKqYNdWqZBb9D1oc8GG2nzACfmLVU8RYEMy
bL+fkeCJ+sZseyxaHvF6WhBKyFY2ivrBOU2k6E1fk9RA+RN/nZTQH/yJX/xWh0HzZoz7GxU5XbOz
sZlvEllBLv00Ha9ZnYSaNhM/QkxzZAMrjiQ7kWC92M94x0PZySX26cx1m7aPurpPFcxF4Ng+SgKf
DB1lPfE5BETtmKqK49Okpm/KxLwXdhlcXWkQXoZ3x4eHY1uKuJQ61L4K5ALLl7Pkpj3a7MdoR/hR
TV+wJ5O6wrHwFbbTJwaVNn5r7ZpoDeRsyKgchoGq3ZR0uKOsLgZoo+i5tcUbfFrmN3hNuifnEaaa
3nM22Pzv2SJcU9Wt3aYSdaqP4OXKA1iUBkDnxrbl00Vnrd8q2M9U8dxbjDsZRRheh1MsyKFvHQ42
zbOQpyNfmJUfuaaA3g+eEQWhMEdTkb5ZsqtLTBsTOz/mzMf1dPipWwIOCmyFR1GlzcbK3pOq13bc
k5RCjsDmGIkdxiSk4GzIZtxSFNcerVAS6yw4LpcAnj8Ecg4RYCAtiSrgyN4wXePUrHEPMo6XtxK0
yFd/AAs7OhzroYj0e7FieGR+uXc4H6dInjARQ5icyKry5bOd0T85uMaGLplS+QooQmpO9mil1v4W
bu6HdXMhmR0Aorac7j/ddD/8B8qzQUCFrUBGozidibFuiOjiyr/k5NdAX5dw/MHBcSxiPfjQ+Lsh
0GZjzlP+aSBC5Hk1gifH7gFgonnYadhcJ1nHmb844HUpbWqONiU5nWjmmGRRK+0H4y2D3sS0I+dY
UIzp4T2Ftv6XpXWbF65uGGxIKG9siLSVs044vx0bZblfdJxuxxSyXsHBFgMUxpAaZ1HoMOo41tTy
Qv032R8DVD/uVz4tfSUPf2ZA2jPAxgpQsDdaeWIiiQnSEBHoSGFvmkyvB81MMXHKgSx8sCJs5F3Y
jVYGf2fHYlgssS5/pCd+QGc2UkEECDbLSj7U22EWhmeo6HuY381yz7RfWQ1Zs9fRujr1J1tNMQRU
IRfB/5PoTJVpOeejMiuEwEhex1sBbeA0j+8ZFSYgjhjeoQCnnBRd/+UYd4DT9mMVp9rWQIROJp76
ZvTZw3TGV7G5aBQcWla+Y8YMIzfMp9fsWUR6/MA4ojDDZgnG5lwN6PKjpAqqZqZh6z9BAo8wVMzQ
o5HQQQp2xcsaDZVfRmTiPSiUyuJmFvdf/idrCbujbSbZMFe8P2Fx6Vs7GTtrHttRhoMOUggkVNfh
SxIyf2IZRJxjCKTul497Yl5eJxBmBsHCT3ZAY0cSTqGLtsXPFSMAifdasvG+IJSXMPrAkmde4Jgp
fm9NtMAE86nF2xzRdtT3KRuwLv/GWvEHjl2WRgxO3331d/NBA7BlwUzll3fdVleKd84s8li3ZTvH
qp3aIvJ5QNXG+nDdLhe30Dy2mxSbG4kWylv+EdIsgcsZ5VY4uEjrFgKaVCJ59GhNFRlWMglukDzV
P0d+R1j2YqnOzVpFQkzYZL/V2D9bYBrM5UhVdhWGdFemiOqY19pE3ygfFc/WZcz90bPF6M1FNHLY
LfdSRAtAUiacOPp2fXRSxiqV01KEUU2Jg9tUjB/TjQDvCWvcDAQZpgw4Qi/PAn/FHsISKvpNaFZS
DrtO3MVvYDfQlKLWWvcmcf6yTceFpRvmg/TdN+0+mBgRkYoBdYafBSQ2vetCTnZHEJuRWaRLRpl7
IYsXSulGVXifX1jKJvMROaezt7E3J7vKdJuBAV0iuRztRaaoPiQzVkfaML2z4PONGIJdqIGBHD9V
A+WClammLOUs6qB/FJoqlIKqeiaqIeqnGDWSKwlOoTVUn3yyKKQotfVDWsIIWDm6+8LvHzYZxohD
RwfO9/bGatKWC/dgpnhYbcGX1yPpMMNhVt0ndyTsl7A8aoxUrFaA3GSRHl2DEZtJWl9TP2iV5pf5
JWbDdzwlW8v3cSNXTCg8nyHAUpXvO9EexC1dEWplvCSz3rptOuwx665zzuChADzBMAKfX+lL+BGh
76ZOJMj1DKo3k+fZ9WUniH1j4SL4TyXqdolEJah+61Ut1oXh4+tsF99u0EolMGG+s46SXefx0rzM
Sptc3AFE5GvfgU3mjOKbxNz18lIBnJJOKlss+9iFhE+Zg7YVioyPCrt68akYn58BkhXMbK6SlNAi
FzX3LwtHfv9nVMMPm9wSTSITHY93Xtq5w2OCkA4tIUQuO0sOs7lup35jevnuwiFqV8MimunuqYwZ
Wbs5ytCu+tvomg5ms4Cbrbg2GE6jrKKrBtkudbBSJiOyGRxBhAQ/vGPtb7l/535hFfDMQr2uou2O
r3OeBu/HtI75ybrkbO1MtqUA8z2URNaR2mSpr7xHj/x8bBHph0ZH0LdytNNXk+7JuH7yQYnXEBfu
al9/7YxD04yHzSDtXww2STuq6AO1H9KG9z2zKvjL0/vweoG9brtWnY16PN1S0qdC7rkrdfqizPlY
QcmCIK/RAo/xILKjf3KQsaDxw1UMM8H5s/cCvgY5c6HDGj0UM4YDKRUn/HXKCUyQCtLDPkPqVmt5
UQaXTHzaUHKD/U7nGrFcwqjEY0wwsq2mIgXggzqscexDD6WpwBx0/qo92YrznwbRJzHiLmYmeaea
oL2NR6/MGDpQSjYkg1C4K3MxSivREjFMKF6tPNQ7AmzerwyEPY3s6PGIzxquvCVRzoOvSD4hJx7E
g69lODxSu68rdpEj85VIksrTeMgELaWwjqkb8OOKXN2ss31Hd3zmImoaCJmTnDY/exD6BAKuOGnf
p7pBPx6Ada6hm6UAPFJC2P6DwGXEQadVf3K+WFkg5rUAHnvbpzQ8FsqaFvffNBvRInuok48+Y/eU
IL3ASAh+Zuy0XJRIzOfZmd0tqru806ZY25e1LZ6qN+i+7LKBa6SnWgFmXZlaLDVa4GHOZzRvX0Qv
RpHu+OO6OM6OO1IFehKWpRA04ONjUhwE0Gd7rV9qCwMzkF5f8xmh5syW0xY81um2IWLu24ehP5JK
eYZ6aAB0OiAnh+aKl5w0DGrubL0WD3Ptn/UxLIeC2AzhCY5/MnI+bLYdwvBUHj2Cq6YIxYlxn1th
Xoht4z317ityPYgXqljEV8VkVh6xV8RSTsmhWF8GJMcap0w40rZvkyPshP+TIWC8TuhUKEl69f6f
kgDOFikKefxleeIKs/d/GcBNNAb5douryrkS4OpLTrN0WKjCSD8IbRPdqlZYDQDvWbyqVKsoubWY
GdkTvPtQFHRyFr2t1i+RdrxnQ9msRgaFtk3QpjnIGWjrWFRptRuuICYDsuVQOyNfBteWXW13GIHX
WkKavkxmH35KRFHYnh+dEOpdYXwU1zlAYfme8tfOfSWv0E11xejnMbJTIiRvEvxgVy3aG6iuCR8J
dQcAoMk44vThdHVhOAgTM3kQGz8kMo7r6Y5X84Wj4fnyZwndZ1IotXJIpkoXymv+mIfs56F4qKAO
e/OGg/v6wzxmF4VFinI9i1XnDYrCc0r57pAeeEwBphIyAN3b6uf3BKQNh9I3gZRlOWtbQQipi8fQ
uSxpyVhRP45a3l8Cik197jwWRGPeezAYiHNKKdP3SSoIINHGNEc1+t4+mM5pzJG+f0QVYynvXGE6
9/l72tDAkTgMLfpINdMCKGuJFFwKRjTyU/28huu06vwuKDdjS5IMceRsVtSeHnmLul7phN8QsdC2
m0Rds2G+AwtuBI2NkGae0w11ERLlPFNu+UYiMxkQdE4yevXrgFfdUgtIMUYDdGKm7FyWRh5ESIUk
xEGn5YMdl4zajW8hyUaGBdZP8CaQ5B4pC9YsVvXKTcOMoonpOvQDO1lcR+R7Mo8Hi7q6fPqgb201
fQpM8gk79zA0uw5vgXWuAik7bIkxe4Lho4DJTV5RFE3PMtuYxn1b55d/IK/4A0mIG5kpBaiOBCFK
byZJyARATliUOEr8hGP04SJFv+Ne9NST4UvkXVtfQyBy4VNBnnHPuAqdKXzR/Zs7VzEm2STTiU40
1hrb+veeDQjm7C1W4vun1otWBhGx3RblsXtSliQ3WaWmsByRjSGOSHUsJrDhnR+AqxyBtzDRVpbY
OAimpNASVVeTMT1o+sHiH+nG1mhFv/wdQ6M3+MINU67Po3yi/0Uux7om5pUCAKhhBtJXnQBh+bx0
WbJVDZvriWoIKB/Geq7kN46ZaeUpC2MPrRq2ZrdbKpPjPvDBl9mFeIG6Epo8NpNq64rGDT7997wx
Gr/OPKVEVmIJuOs+NHKmYmevlkg6V6UVIaAfqcKYMqH+MR3zurSM4XEXHhWJMtO1sItLvea67HZv
bC/yvkbafYd5XV8OBg47D5u6tB7AQ7BabQRaWqar2kg789913xXK5Ga81w5R6Az3oDAfeBjl8hGY
Ou3cXtEqe8QphHUv4zL+Z4uBssbwE0WbubQ5GPoom1AtCVsBgV7uNmn1ttSmz/SoosGRGzBNnxx8
dpEm8OhxaZw/vfqwVh4yL9Yvwqh15SKsJw5eNqwISt5AuL/E8Ps36Z3ZLseesLddnsonHUruXK3l
if+hOApQ85wH12kSUuMH1ZmaxNhiFzZf2cPboEfm9xkJZdUC6QXIasZu+JHaSrgNs9tgLHr38vcm
zQiySV9dJQ+P5ZE+tRhAKqGIpzc85ge1VZW5N79Dcc53jq8dr9S9M+6n+mecfmRcGTjZcsXKXoxy
XUQvmo2u5mEZ8f3u2lDuV2M3AcrMN6RP/fb11boCqMdeF4sIMTZ6EY3rGzHE4/Eb8DFHRcTmu57N
l29akqQJ8iDH9oppO+mAQcU+9SjG2eZMgylRgrwr9XEkWnlXXr0QP5gM15kc+/KC4IccnjYcVMh3
68pz3YywOunZ/BiYNOeDtVAGn07nJGzEIV5q0g/4kgdpYarnkLquBTGSBnNU50llsfYXjRlz90kD
tCajgkV93GHyTQtVmCo1Y+d9R+uIB+Rcjvpx8ZgPbULiOil/3AT0FwPEIjEFpREjgUkqf0XhUeeb
UJrPFCDOw7Y0e3I0LS+kLyUlCM8TnmjF77a4Zz3KTWvE/YwYqXcJkjnMoulggxeyPhVIm2pI4UjY
r1Oh539KDNSI/CV+uEZtmtl0Mk9uWclVXpRK0yoAD1GiQrLMpShkNP9oCBhzTfzLFl/ZQWm5Q652
VorBROql6PG/78DfosFsXpzFWwTfIofnkid9ZVpgKrrtsAUhJYTB29JJBwRZGi9NQhAdpp+me/Hd
ECqWI1rC+AuGJru1sFJ/+8tDl7iusoMfd6su4Hvf1SX2UOiT7s/P/QgqrYodPeZrTzqy0e8ljoVs
F/vx2MM/7mp/lq1bNX92/J6mUcYEf3X/1IpnlQAyxBXlQujTCCdXbSbvWP2MFc5COSzWY+nIMED/
DoSsF7zvFicC7LU04qyt0MGs4iN0UMGeIdoVeKTyo6SyYgNsXudmjHXRHm6vWckfMbPvKh8/yc3m
IdBB2ke84FLXlJeb7y+6iQCa29ALL4xU4ULkeWrbfXjVf9ErlmUpzyDjm+uCzytxou5Y0YSiBmqy
ySz+7dZewucBpg4zn8EbOsQK7VSXO+XjIsOteyZ5e+6e2LJwAIJeGzwYWuBc5YfikIeBr0SJ18ca
cW+roDh/5WIc+l3ywiNG6AyeDSgZYrxpWnNNx7RVqDURv1UvJE5ybYiZlE084L96zMtqNc5OOxnT
qXu2Ni4lb1OBvZ9QLbLGd9etM4MzKMTYJteGYSCkUkR0NoVU/TgFtLWPOLaqb7JrWK+v340mLZWC
XHC5m0CDh3Gqq0VdXya1nml11iNZzmdlqasDdfNDJY31R8FZ6pIgX93jesk95BhBY4IdNsyTF5FX
jfBMg4h3YkHFkTcSROcLtE0KggIf2EefrBHJUfusnKnnSkbp+j7YTZK2JftNucxaX/pnP+NglrS4
nIl8+7fMHoIPw3e1OPbIHfkK/xHC5v5x4FRf3l6s7yrwWKzF+0zYd2fC7sEJHjLMQq5q4ahbHFu2
ksFLYMC68lTZfCpUCD6rpYcXkVap9geq6IaBWlaNeWzcPj5f0or0r9lT8nhk1kk5Oqv9qW5aoof5
hIp3l3wzC57tA9k86vOhqWCa2yN9OfmufAK0Au3jM0Y+hhRlKtG2TkWvsg/yp/V3JhURFnr1iEVp
QBpRmKqYOgF5Qr6iv0MuqpqoHSLj5L4c8e5E1+GEtNJCydlFx0UygTyhcFD628orroFy6HMAtAUt
bDi8XuSYI9/eYYExl5HPjD0WFKunMf8c4+emLCqjJOnwDY+cbmOcj63M23FWyOvROiRLDu3pm6BE
Qscu97qnkFifHmWNqwhI+qDtcHhHaF0zs47t1ke6A2kkzyzzvXkMKGfh1qrJoBfX/5CWnHRE9Qbd
2ZiKS20dHjtc5ipPEXuj5GfVhgRy69msHvQNgBJSIv7YQgAQLUmxPc5LknY8M4+CIuzTO2DudjXG
iOeArge2CiCkx6QcaU2dbttx4DIYl6fjLdSbMkAJSTn/lNwMtUErnfmQje+xqR4HqQD0fDGYiqlx
HTvbWgplp70HG2omDy5K5FXmpuaGBj5fiTAK2b/6AxuR2e8YMKX3oalYaCPY3B+JbSA5zOUDLmDP
op+DPBgM12y6KrxDTxe5v6BW001AgObiq1n9v1k+koxQllVaOv1Ua5djqlpEuUmDkLMB/Vw9ueOR
ClU9qSDkCHlLF8DuULI29Yn5fhdb9oXk5JjyV635aJ7PiF2muWNydgfhA7uPInUtftGkcI1XsJjd
sKzBB6mfNmiPZSeaKPEytNFcbSBUlDBpTbdg/uc7wH3GdWYXMlCW3ctuFFa1jA3jFA98wTtEEzIC
Bs8rHGYbI4U6vzEwmTMOcKf2VH/r2/doyUSK7xntYhp9KaqF8iXwcSSavzzl+yqILMfpga/mLUj0
xJ33/yjfZ2Fl6JsdweUhscQZboTC25jh0NjJCKCcRd7eO8fwkeNLGWQhw0baxxwhTaWInRESRnFM
seCsx/ix3FI5KnVr6fwbczpQPSzZjt29V/zkKjYzskH99Ddr+ULY3ByjbwURjW2xr5sAnh/p3iNo
nLZaxGuZ59S1B1VAsx4qKKimvP3sxCbbZXkjyBZi614LJTwOSSP+IxE06yu9R88gyPiVuPf5w+Tl
gmnIbBW4v4uaNLvL71H4CHBTnfLUW68F/2D8ogR89wWDeprsEYFlnJEAUSgTs+bvATCKw3VmIy5S
WbtA91tUs3bHbpp9FLmldlpNm0c2yj6wrm5CDDpwST5mbc2FGoo3Aw3D9EuiJU6mop4WNKtGeJes
Re61OK1jaOYLsCB8VcBdu8ohdHgR143ATVbuju9SQ3xX/w6wKNeZJMC1tds6/uXeuCgWgl/yziUe
MJlxUlSCnE418Rx3ilNKWoR+j/P+U/JKL0ABzu9OHELA4j4hLlh6ISg24KvygXqD3dDfERPiyNDx
VQmzoQJlHw6AvlliTcsB+lFKoxman3uOVUW8PKWx6cn9OMjtzGVz16gIZqfTxkkucpP0F5Ms8H2/
jTVNpolEJRUQLi3fENbhvivu0zjVWdtOSz1J41Qpwc5Z709Ot3QfJH5ZeWvvpOSf8Ku16x2KYx88
Dpu0CRfUArAnmIpvPOk3+5hGFeWkdfpWH5JHcmiJ4ITvPzWTSC/lbg+8kVN4iTOVyMh00cHA132f
EfCnrteq84WvKgAgq2kiFXKm0gfm/BtlxGH8OUfCANljRY++kkXEY5lMLleojdWXPlh8Zm0CBzkQ
Gjd3s9Wnhql2nx1SQKa6aAL/GXSXfoFpVdqkp1DqD9PKJTL/pjN90klw+VNvaqYt3AzuOiIwY8Kc
h85E7OP7NDITZ3DSfj70O6smKIzDTHVTsimSmwo8LiCCmAvfCW0v0edoFmM5x0768kf9TJpiqX3h
F7aLKiRA9SbbeC62hYA9U+Ui/xkmULt0+FIHWf71MmWw1GdhuqzX4NyUmtEkrFPf9aimnB4ixVJS
A9naJEj7D21yPicGE2es8qtKsPD/g6mGQz9upqndXZp1DYYs6K3C4aJUlUid8ui9zeFfrUGCIUUw
jXwnggCQIf+mmIvArtp4vxFICZWFbvTj/6F7vhy3jv1KFSn/zUuWrOZMEV9qV9f0Y0CdfMQweGaS
UvbU9sjM1lfN0ePJqRlrFXzaxAy32lnlx2UcO4Fh9ZBwXs3fpwUE37nmoLSaenuwRxsIJhp3hiBn
+8DVt9go3WaIuF7LS02agpMhGmOEKSa0mTbDWM/2RWSQtamCp3cTghcclowZtxLWWVb2lXU93L2+
5HDKm96JFMj5FvYVLyZsoVSpb/aOH/2IWyZx0KUy8aD6QxakfrPzuRYFfNhbgD7yJ5gTilUKHYCH
n3RZqqUrsi+0FyHfPr8Pfxe0oWEhoZ+i5zVmInOY8L0J+1vGnNhcDExYxcfWVBcqoR3ZCVqIzZek
nHYFCD28oM2xQ4eeqKFySUAfjX4WShr8Biqq8lTcjRi6cHkwR9nseOlMiUUimZ0lVnQXpPDlzNO0
wLZ0e+UT53qk15NGUYv+uT3ZIjXPmIetV0frTFVXVpoeMPJ6pID8S+qaBaIoHzC5SuP4EhRFnG5u
CQfPbxzwFZ771JoYU9ZAufWiNByiue0Xu0ERhsDw8EAc02MNss5uF7a8gNk+pyMATMZNa6vt4NTV
ghx1Pf28dQYi1K16YTy1j4qgzbyWiwTdxo8Mr/FaJ9qro8nAa92fUMTgYkA52ANl+pOR66nJAiBk
Cw/GmuRWFAQgF9mLt2QBunMps11D7BOwA1AaSw2Mb6uonGqaFPLVSV/q+9wGTWxQh32f+BVlA4xl
RJGCCvaBs5ku7XqhzRHQtj1ni3ayUnnalx0g+dwhlTVNxKSn81RGeSdqf1XdWvQ2K7iwL+/izAxF
SiRGVWiBrfgtnmxHIBFDkA3fe3qgl+rHlJRAeGyVDEZG/DayuUUASH1Cea1ylgX4mFxHSFPAesd9
ZDLQSqPyuLl4U49ZQG97iK1UeSCXsqKGU5YYfq1g5rpnsQe0ZpUci6DMnx0pyc4mCauZFNGnpnQu
ULu0wlzs9/IDrFIOOg4qxYWHiznSbWNAX1dL3e8NBp/MkIWXqjgrZVWmFpitf/Pmc09+Js9mJYXr
jGaypNKNFnD8ge+2QsFGlGkH4i4lMaK2D4mAZCNzBSYBcFtAa0rI+x9UVQVFr+r8PGYE55HcL7yA
lXssluFevz96a6Ny4n+7Vo8QrhNPDLitsgwphjTfDmcjTU4Us+H8OjVjGK4rgFxFJhri0DaozcZh
VAbn7JJoMpc0JJXyih9Yn2JstoyfeXUw1cfn08Lu87yfage3hK/7Qd+u4IHC59za8UTGgQY6Vm5g
O+YkDlyeO9qRHsyN2aWyZgZZGtCks7IZr1bSZhmDP4ed0tqijIgYNqisZeBIYsiBRAqogqz2Nl/4
W28I/aYhqDZJ/U/a2U8q2U920cbIZNn5oyIJbpECdo42zv3cqxHDE5tEfB0eMtt16xuphcMCG5xn
qaOzK84uhSCamN1DbXan27s83C2GaR1QTKv8Xxeo/F9COEvXTJDYviq0vFgDl5y4efQVBAjWuGpo
vJfoJbcXwkDlduuhPjkWa3L23p1yeJoY8kaMeYJ9/OzjEWhrJ1TYCgrkME+xfPLl5f2j/K8rXVkr
jHz6mIVt0NbqtDIZLupr0GlyOt27T7CPPbo0eB1EqgnLsJlRat2Lv/TXDK5YnlShlKadWGV0Bsns
fNbp0VinXlYVygSx0bSrzkZV1zMAJDs8ZSaO9BH4rgwgChQwZTGJWfdRsCiXc4oqvaENtH9t+8JQ
h23pcGO7W2gfsY/Rok7z/tvIEcAul8FxlYTdhxFaowQgGk2eAtoowpW98dOedMJgNP6lUBBTF2v1
NkfKTioqXQkrQ6O3rHv6V2kKQAZV3Ui+oCv8HpIUDiTHtloWhg/qEwv5o63q9SDjPO82+9fXwY8Q
bOUhVV+ZKDAuFBdFBxNvZqXO7EFDH7Dc+eSF5bwrh4mOo4z168aFplM7VFhVprVqzGkyQSInx4Cm
nhtOlGfH6CwVqpNN4DukOXQNNFdzSWGX1g2UFv8cIKUc+kY0I0qDAc/T/Dckr84g2VdUTbaj2Iz+
zHKORaOpkE73YtotYkcBCy+YMadtRjI0PCEkRfenc9str8FigtHbVTw0LGAnx+8hHIA+i96RjfKl
nr3MPqOw+n34Av0BBvoy2X8eiRBUkcQ6gPT3XdIxWHdnkqRxQaj0t8mhprSf5UOihxtoiI46uAM4
kSNCKCg7LnYqUGMhzwVF1OsqyXvnkHnqmhr2B/9tiQ6ssJ3vELtK/NGODrJw2O0ujIc5OzX5lgOZ
YdRPuRg0YHP2nJN7WtMwuw1yNbY8ukL1V+8/FGHXRwlgIcTTRiW9TGUTDSBJnWQP5MN1MIvu30tV
abeueffutKz/S2uvntZ0TnW9nuO7hL+p1Hr8ZHq4noTlBSe2OFqdvBG6fJc40yg2ampaFNjU/pTk
saor99L2pjho8ZH4BGTrxblrsJVnFzlSAX+zTbKXiTt4pNK/JIzMzQRfBKY1g5FVI4S4ZBQOEpqz
yAkfAzYa/zG262gDHBf4n3YKFRjd7PBTK1+X49tDJ9oxZvZDdZVvl3sTE4rppb4OdwUcpQMLzUTL
JM/tXcPqv8ESn+k0oxrWnR8XdHrblYGi52fug/C+vFo9CHkZuYh5LGW9NOHMqvytvhtoGdWFJJBT
yKQJBXEg+dWGB5/GZMiUHGpiK2xrJBk87Zcz4Fs8W/cjfg7Yf58LAEZ1AByfxwFfjTALgMV6VPIT
ThC+hqUePqOsNtTjUPxn3Cw4L9THWf+rnVa0yizENSM6zWmA1xh7a5FhtCwE9+CdThwCNxkjMCLq
ZyUFZsS4l4U9siwUphBFwVfgrmLbaFu1EQsGq1d/JneshHOAXgnkemabmE+Z4Yy4/EVQ6Nofd/Kc
p4pnNUHXu/cJgz/yPkIXuXeWMAxux8H2W14g6WIvFkwhgrDU2oZilC1+Umy2aiqFnJoWWsmrE4Ry
rjTMhOtcgSMDL4JFgyqcFZDdjXD7S2syMIE1NZRuLodsYIUUquQG21TSy+bCzrpMyqbN2XKv7aaS
6+WRArDnVUlQCdrQKLHM/RMD1iP1nVjXx0BVYyVRPAwNFBY0p3BC/cInF/QstRN2kL6T6lOIWljp
M0GzgCqE8O/G/7JlMOLt3EwaNXE3j/XSKPo5KmLn3NAQiWDXVZLtJ9iI1MBblz+IazDK74w54TKJ
AU1szxygBVTFNY3PsOHKSn2QfUmQ9zKmwYzjFjSe/bhJl1y0l7dOrsVSlq2FNNin48cergN63MEQ
bvdjjnX1pMNz8qlg2FRqteJyIUB8WqPTs+mgejr2RAOIe2OINzHUCxMgMn6ptCJP5MT37wrczAvb
y6bX+qsi8U2ajHMNlnS7z66+jIu4tZdiIsVF00/i5PaM18FO8JKk851y7ppbBuK54rMHaO/miaZv
adnmyrn/K3xXmxa8iUG/8TbXIGMH4VIXe9IZpH9zkR6ttovE4ZCiNkaFop4Dxi4P6lpOPUgi1XET
vKbAt9EewT2JpUefqxPAJ7YlA3bBFhiT3WrgAqWGqSoHe90XvNwLEln6rBNc6zu27qyuz5So+UGb
zAXjln7i+pnCieuqT0p9vY9JQ9f9rfUzDn6/SZJaTue/L2HvgnhmJVe0EexzfWvEnzX6qgUAc9NA
WYKs+Yp8MA6ouyPdUWOKYI8dkiM4KZJbvPuiOivggluCjetzAolRHPvOTALugUHzKvJNBE32gZDd
X7Hr0BwnVq/wo2GlyhlfYbDh0DdwB9ler7v5jibPgcG9dB0QZAN9IVUUAOtAdRgHxDJ0/XUUxnCi
MmkqcvA05K6UK4yRNqio/TBnVRADSSXHamELBa8v82M2dwUoSelu4jle+QM10ZD4vazWTvqICuEk
3CfYpD/Yhg2XyTTFKeLymiP0mBx7BJNzticuMlqFIApdT4TDNzlIgvMxbElAog7IOFuJB+EeraZy
iYayQQT1J/zn8K8mPjm2q3urYyuKzbvMvKLL2eMQ92g/F4GC8Jxf3DTlTlFidPFUicoIdFKPhJpB
3ffI4ov6L8H+jIJt8NVgbuuzD2Ho8RDlM+ZeFX247AxzKjTewuWcfkPSwDkMkwFgemMlZ6XuhpvB
Uzyx1TPbeiBxNawb5aXbET7mY2EE55ek/4cjdk8gbMoKthxcU6QoShCOO+It5ePWM/h53FU5F8HY
znjdMFAL8xhnC/32Cl/FARgI4RsiVrRGfY8S4edreZwX39HWgNQFs0YZmErv+GGkbFNFCrIvZeyA
N1VjIr6JG+BgpLEJmaBjl8gCoRLaeGJTff/7iplb1AYL26YYRYzN0A/6pxqOT4UNKmEb9zpDhGmF
egOosFmoS1RK71OVuWKyDXOYvXGscLh+Mfrq9aVFR8+YLuUFZsHiEAEv737RDevZx1WfGaC/ef4/
eMfAWHHxk8ynz06XSLYLPJnt5zTKFmh370bq99T9IGKSSiSlk5u2Nv9t/M75hVdJg/ReSAhB33Y9
i994TLTRXfW/pV2taWiPuB9haU8SO0yaovLQrxoqw9lYm0tzdWtL5W4yg69h2VgstP4yMmkDC/vv
S3PUU9GhfBKGRcBShFKfUE9HxYo/4RDS9VbyxiI9fX7cMcE6n2SEYXyNJanU6ueb5YBgpeqtOfBo
801/yVgoVQjn0VrrNUX6f4uRWWj8s+KeqWfAa/vY+0buncdr+QbCOR/9HCqvWqA6V21AX1kmC1lm
3819PMuhJkvNiqdTJr6EVaFGgpy6DKczQlgqQnyHQrdyX+nAKcosatWTUapImD0Cih/Gd3fcxZ8e
+PxqLeOphypLVWbPfzvu5pKxGO2ocRQSqb/0V8GJBso6Z6nMzWIY1Hc4u89WDqj/26NOMO/Q3SL6
DKvR2VrjD0aErl8QDN0C9qc4J8Hr3JonBGaYVn2FsOXOhOD2WyCRr6t83vzN4eDlSbY8vEiFV4lC
E9s1iaoLaaTD1zJnxggY/Z3TXfUQ5AMryi5XvRB8R9uRhVHSk7kocYc63WtixcAMIr9DdWXPFq1j
OGmhOzXb0XIL6yiLH9as6wFOylnXj4diZG9SdJTRNNGcTCFewX5vqQBLIhX/56w+xgBxKBEhYs13
4wkBRqJfXa2a5ZYxBX2SJ4v2p5PcmmgCYEOSNkrzmHmxMtZzqbD/Ngve4scxRAhZcCQS6+G0IwN4
NG2CAdgceg9nIEmbTTwNcXntos0amUmncU6kJ75f+w1Wlqw0myCRQeyCnFVgPAGPtAby38MWr9PL
/rVl39rWl8we8ZjHHREPQbVniz1wHPKGSWAMCCjDherf0w9aKki8ul1a5yhVMA244vMxY7lCufXP
oQCa1I9v86oEbz4oSRcSPuDFBHMoKhQClqAplduVjaFxRi2weAT5JNbt0eHwKxAlk5hMocQIC5W5
DNHxMnft3mql7BTW4bADMPPhGtsI+zWCoNe0jnDMj9SYtGf2ue2H3QmzxP6A+edjAmu8aPlpSmAC
sngc2a7AV8aNUhtbFDsxKOqzIudFg/MGL7JhQCdks2V6DboiSYaGCY0kWfzn2A1NAdN3nsrH2/Do
f8DFtflI07a9kdeZ8S/8T+p6E+VVKXdnwdqQCj+VYh315y4xTC3jp+p85V1TZc8qPRQ+ETpcapZy
C/C3oSW+71oP27/nP5sBsqjEpv+Y8zM9pqO+gjufvaXdfelmAW6j7+24XcoPoBhBmOG+BBOfxrR5
ytLC3xrwI9sOi64b9FvE8mRPztfrR2mAIBzK8kDl7lgFS3OesRwqgrJ6wGVqKgn5h1wLG2Lv+Wuz
RTSXSZCUSO8bPcTD7I4dDs1YM07pullNnYpdpn1TAt+rah7mbrEkayGwIpn3BZLC8/6OZsQ/Icnu
Hi3kT1K8Tg4W2jQdSyazc0qAZnBMO6HECSZKFGcws+VmTNhmQnczDxki6eHElutxr4iAevxTeDLO
7gPonfKKUpMTve4TYRB0cWTrH1+Pbi05oDbe1y4PcIGYg1DpXu1GDmu0wnQoNaklGwh3j2QJo+1o
+r3lN193BdZkpR0ggq/bhwaQrRBWZqrtE+lUAc3NxGbI+gFcOIGAsx5Ku0K6IELzCGF8vo5Jt4Af
+xAoJsP8W0Qmp+uHoIz5d7/2npsZt1WZMPp1sViFr022Jywf42gQoriEKHoACfOlv0J3kYpX7ff0
z9S8+ifCJrphXhrUG5DlHPv2OuYMhSqoBNfRqmPUQNKtOtFD5r531/AAYSVXRdntC+Uw0juJVJWu
II5mVGxROD9C9/FfTbMD5uPIQCZLhsXp28AUN6M3C7AqQzH3qot69wUa0p+Ib61P+OknI+OUTUGk
9zlUtD8xgIp3mE+QKGmM4w1Hau+X8X0Ft2HsXXA4hV+tF0eOqAPjv8PA/tmPIC2W1n0Yk6W2t2h1
DaXF4KI5TE0Yjs0K43fSn/gFFJ03PuiUx0Uop7Dekci5FcGX/c2W0XfM6ndDLUADGmRG3ch1vBhI
cbMf3BK2R/IHPnvmPOKvNga2Z9QhGNr5MPU7+JqhV4UBL6Pg9rx1HDXfnPLZodxNCmEyShN3YVIG
M+8Dva3I++l3A6+NONHL9y4+b341QsWSPCBERNGv5aZApO1I5xfEtKbu7cYhMhcfeXVDwvBbbnyL
vkNjNB/0RSpB0zaYffeNoypGwTS9TgYOUm1yL3OKpN1CCAsjuJSu0Yet3s5OVCGBp2EYCI+pQHx+
DuSlaWNnrR0rfzoyEZnPESTgCtl0vgN0+6hoCL7vFnjz08/9nK9zPvEGHbl0kCV/XKzHHQTDFUhj
WlvWVg37TZSGBqBenw7TebljYgfQkY7HCueQ0UtVZ5UXBTIHR9Sfm2lNj/D0R+TpY8IZvdr0W1vO
jdKoJbPMc7VHDjeF2UDe6cwPgbHINev3WdfWn58Vc6GqwxfczOINtQeirjXl+nkBwOE/4UemfXfL
RfAu976N6IkuTAYhwBiHkG41QlmZIQiuv6VpGKeg0F6QsYYPAg222hgIRV3JzLvgMMNAe4BNUzhC
Mp25/eHY61NjwnONVobjqadJPZqjx++f3R8NjwOFIT1EsoCGmOxbD0z7GYltDLCWJuAm5Z3+kMyj
z+wO95RVvkyR6c3ZnqhDiOKTGuR0hIMNZxq0il0xKMFJzfS69il3KDidCgHRwMtywvtHOuuWNDY3
Im9XfHDkpGMXLo7/14g3LfPIQulLImng21tSO28Rl8KleyVdJsFljLRdwiEJAyVtK+zxaGmmlgX1
ECWdxBax+ft03MmAZM2y0rs+fsr3oAqFbenAh/4RqcO7+4EbSuLvnZr+t/+CFZnHsV/xJU1iNuJ4
g3cIq9G1v5LySMk5XG3ZxDNUP9cnuM9e/OXNVtfkRQGr13bEOjG9Ts0lN1AfHjmbffvfmrWuSXj3
CJiRmaEpfx0SnxOMcCzkhdO2+17Lwr0cl4HVqxJ6pMVM+s92ojF3AWHyy2MBb1dFb3Y4PdaRe2gH
8Y/lhka8P46P5AHVE5Gt9RMcQMGgJEHBGsg1oUG6Dnpjw+/DcT7txSG8DhRUNtLGGie6FFeF+DkN
4FI8rObNrYmk2PiQNYHFiRDRZw3SykGKUzGy+YET0zbVZwwlto7BgjQjYeFK9zsOUHHnabmGYcfR
ooOirwwxmwmSzK0Pjon0BbMJlHMKBQVRBGyHj1UhXAB8Ln6HDfAh25e4oXpH/Yw4yQq6kOxQcScr
KGttpZdxThxh0l5svGoSbXBYnJqLgM+YHykB4u5H7+Rq5A083DvwViVdfZ9sjGM+BxCySg8/lU3T
eXwGeYmYyDZmCiBbV/SzyPCWj+U11TALp+o4Vgm2V0YxKBuCsZileUp/R3UMalew++j1QXUdPU0I
aeojWFGx5eGM7BwIfGMnBs6uVhq/5wAd49jjKIVxbVQorxQEFt45YpIocNYl8oDfR9Ap0geDLBSV
exDFJ2AYCQlazLNNByYiVO3zJDTQTakyEs60I6fMdlCxYprxo8Rm8aNvp1hmdi+CovTIQjLy6aaJ
mtxoRtBd8SSG6btTB2zFRyzXdya0CEAh9tvrfCE5jYSYJ1ZpznnyCSZLScHC0C6LSn6Wjd4ULcWr
+hlbyAH2q/ly9NZzhBZrDI4VZGI9yTlSYOYSue+eBehx/FdwZNWH2vXjw00LTgpbWdfMIq2nCoks
rzN42jU8gjI0H7P8R6JL4l6JXp+lWY2zp89AuPLe+yJp8wD+fdjc0aEaYRJ5NLqARWWMUX9CV+LU
R9QVlZ72oL13d+NDYEMl/ClsYR7QsRNcjuh50+fVzcu6ckOdTT/U2VBM15kR2yh4SzQInlbV2r/k
jQEJsA3RfrDFrihlf4T00/0jDVaUYgGB+uUrs+HP4rO4Ybv6aRNdQsgcu5MuTDr6iQxbpROvf1xq
ntFRR6Tc18Ie78l7ugP8nIXWLCfW5ZBH+Q2Z6cy1sCvsHqjSm5ApG6OuVBWD77VNINIykQ7RfGk2
kc2bcI9/8gjIE0P1za1tHYAaGYOp+W92L9hWcqL8VX/v9sSe69+flZAHzv2KtsPhuNcgqLn/LSIA
4TTLAYwuMZprFXeTbTIGfuYaS5VFSi0WFMq4TNZoFyy7dB4FYSLlPLx+qTXK5CRRBR5pkEqCaj/c
0qSKuGnGf8D9iXWnHcmfVdYL++DrTWFmxUaz8INJ1C4Gq6pbR/fJS534ZMfVLDsvl2YyaF9CGOKX
cpCTuwyZ+5bJFGA/p2LjyjIoeXtzKQbiTwUNlqA24xRpwhdJbXuXOK8Yb4DB6yFvvxJo46cSyJV/
yOkfbtlUsMjIJz7VfCtZ5TqmyvJiklwbsjAMMkVZyAefZDACI/KZs+HUa7uXbypw/U6D3UNPDBHL
B2L8mBdYx9EF11x6llMc8JJGAPxLTXBy4EduIuRRHIXO+ncMIZO89kGSglGxkizHphfl2evayCkh
fL+WcSQKC4aBQP3exnYxcLuFPnDxWIhBYSt6VW5/H3gRbtCxMWIqGlcg8vDMybpJPpBpYkvXhonM
aRSwoNAjEdAq57BxMT6TAoOpDnkc8Dy2nodJyaUdpRbAvlixOyT6u9ACFFMh+UUnInjcIGStPhWV
xRrzThPAvx0I7XLR0ewjSGGLNlSjprKodXBO16l9ecWSp6RBDkdrgxE0dxJsdg1dcChte5a6+U7v
IE1OdV8NItweWksd6qd5ai+qzhzYRISFKyNrgL/Q0+ULQKJFmx55vjZvYrkMrn5+9+6O+yaCr2T1
P0kK1Fr9xK4mFXnRb0Asvrmd8gLpTJ4KSdziV8rKRG06P5AiQ9PHyKO0gsyqiHMxtJb4D8+K776K
jQtMW2gfrq7ySUtQeohSuj2I+WqJtMl0m+FX3F3uMchnYrByxg4V0alq+aB54nqzQBan570Q7NYr
3Ll4jy7cIaCCGyDbvFf9qiIiUvioeu/YAVpmCIHK3o6Aem27r4RIbQpMeAEYH7ABvflNCtJSV9Z+
+doKO1JCbQo4wkjgVkn8cH4Ff9sFlnJYaiVXMtNvx7J4RlRJNiNMQHzxzxAkAvjfWJ0sDC2AmKCt
Ndpr3MCezeNASYEOUtPFO6cqI27q+kGasV1QVJkzqQAdKzxj6BLVNNHADr7ZeSP6XpEth3LX9+lO
V5/8NS1b0XBxujfIKyWCPCkFv0kNtZqZKPoWbzVViaKOvripcw42ax0gzPwDzht69Hp9zvaJkTUp
7zK/baejIlikOq+fVkJNLOx/UcpT+bOoQtbqFuhJkxqiMYVabWWfzpxfWCsDLJonIp/jGtVH6vpz
Ti9ZIuVDe1lSOLyXGjWQAYRX1ntzZ0XiqF/fbavvDKxpV8jJ7/pLhinVs1gb7WGE6+51JNnFzJ+m
EFG+mykIzWATBHjafHEqTybE5+NvnQ3nQHAPsbn2jDc04zOd1ObYtgk9CgpVuo+3TJIgUaDuoXSe
g2ZyR8P+FZfFNFDS8xDVnIq95zqBHw0/Zl/iAl3GlUorB29vgcxmegfbONUxMIx4H4udgBG1qJb4
Iryy8aoQ3LSYj10T6ZVTxwNQfQzRLICxjLcKj6NQs3HE1pAq5IL42bSujcGF10jUC7r5wpZg9K8G
UClfRpQ1o08DUC7NUWF45FSbiZYZVtIoS/JibbUMWXtlqQDviZnb4v2e+QfpyrzsbSf7tHMYcOc/
Ih4HTI6A3WKbqxJFjzCN5cuMR5IY48ZSKnsyIAHCuxM3GuJnYYquQX+D/ApX1P5zAYYFg0C4BOEF
/Sz232PQM+ACPivEXN3+h9zs849Ycq+X9KkiY7lNuhX8FgEKcK+8LD/Ilz20WwZg88Ir7m2pOdYO
i8PEekmj+uBEvlc3RFnGX187hRFpS57F/aQz/iWc1C4/GE5LM2yefPIe4vtCQP5G7dN9kUNQ7o7T
5KrU0Hg2kY1oxK2Rh0pswQ3dxiebDNpx92c3v4x5JBNd/+Xz2T2PRyjSO+Ykm9vFnPSA5bUG8Hbo
7abhTQVvQgKRX9u4LRA/LI3Dh02CnwY4kw2QJcaaMMAZEH0Xp2Wjac28oAzeejPR/6RM1G8f9oJY
fep7vH/DB1+JIIn3jZBkTscqNNUcrxGSfW418ss7dwEP6Qeh9Meyt2jN2u3+Gp/vLhqn1xFOnZEt
rWi/g9wgCQyMxvA26CVETFMdj9JEGbtaxrvfrw7eg86iwrrYE0WtXxVgY5sHggIVy4upbzjpXLiw
b3onAZuFTUVw92n8Og7k1WuEbfQkODWj1X4W+gn9XOVJoOZwpxvlX+RuUKoY73NCTM7xiS6ulKh/
d11/2zMc98x1OsxlUk1qhJdDXcWQs/+9NAAY0LlhYNFsYjaOmx2fNoErazSiDKM8R1xf/p+kXWVe
VoP/bOKWgXVBygebX6Iy/tfBAj44bO+Q8ewytLshmKPD/2UElEuMvdvmcm6+0FwHspPhvbMKhz9i
ap220fQXNiyoTnvuc8Nh+uSyGOzfJ0DK3DOwrUANlHAyoklb3X8wmiiGSI3PZD9PhGR0tDwgVl7Y
j5WoDWMkCM9taLk22Zcg1W1YA99uIc7Y/nB05pPSNeOSXAry/1SMSWKYqimSznwEJkt1igYOgQSQ
irKbu8lbE+O4WOygp0b35un+XsSoXeVLeScE/1jZ7fw3GgmE+VaoofIgoCDaHiYwqTn1NsIttlM6
6xmCtRohbvGcO91Z5Xzs/XwMqBJ0B5lJ6dxDOQP6aNQrCL+6XjT1Z2dKbe60EhNOMsmCuNX1WBnF
kiNsQJx4ghc6NifpyeyDe/ITl7oGpljPwhwI7MFmZP5DLLH6A95fH3V2W6FXPoG5fPuB8alb9wor
kfnMCU0m5mpy3mMz+Zs37KlZ6S1UG0YxJ4gZ9kRhR1TZMST0zbpGsRyA3NWLLyRkyPKfVRdv0y7V
3F9eXtidoV4nGiGCi71vE52op5WDxXgr1gL7WtcOjrNa+4VaoeMdSBGXTdIE2H1jalRc7EKMaCWr
vdnu9f7jx8/QESaiIjgvOeiLllbzspHfd33XGYNBbRfhgfy6cPozCG0jfMASEzQfPDxPy+7K7bEd
LfcP8kBCqasZtX6kGCM1LVGTQLntUo2Og+H2+Xc7dHleDFeD+wBwrHQ51BJsCxGxVegOLIoXAcKe
x2jRpcOrerxEDO6wun/JeJOQoi6XXCKQItCg/zs3tQmPYE+0RaXKU42mEmFx1J/j6S26stcwvoac
e9v1Owf3HFK21+tbcm2fO1BcZyq6yPQpHGcgQc4YtuqZR//ukFRhLdp02M5nJp83IkGtqoftxf/S
ij3Gs055sxQ0Kg5vb2nx5eoTbDspu59tpcf7jnylVEecIxlkGRpcOPylIdqKYurYCrjAen+IpAik
IEzG2FIaxhJ4HQi9+MPbinw6LHbGIdOdONjyZFqRRVFsEOYLWmWTjx5EW3Rv/Q0zy0FlA8lIK6z4
0hMsFl8c8LZ2l7QWHUMn1EW93C2SYfvmBe3qrwDnt3o/DzYPoktZs6vMsXyFF3tP5jp970jpvpUl
k7rYRoQKwZl+3K6qzijFQR938IFxCvglTrJg3AfHXHOwju3j1S9Bfz/Vvrrd6h01l6WyHAUDPjJy
KJNArUpQ1h9Q8XpVrWn5tYVZsfrJX/LGGhFEN4uOY42NtIFARy6A9JUbtFfyXAAyk8vDkKXk7POq
RyuTO3MTcrf+lxcXkdBTQWNnZ3yHFiKNPqh3PxrYA883mY7vAl4HZ6T8LBbSDOXbkMXHT0d8r92Q
ezp70X+rLaK5TdaDrDKNhtDyjoCe/1Bv3aKw2SxIMEGQjBF8uVDdPL4w0AMhPNUQJ8jQ8wrSWjJM
Th2LCNMAOYQK6q2CftRHrzdF4paHP2GZWE1H2ahxvu/jpvTwBVe4nNvNcEU8v6XOP7K9+whYy25H
yXRqwhBZLSlrviaa+MuC/Qbcz7v6/FtGVIZmw6zTQg+cvCHAZlcwY5Q+vSa6JVIOTZdBEVUbU8Ep
9ANfSzc/SerBN0VBSj5OUxFx7JJzKrDb5XnpVjAL7mjTsyCWKbYKbA/dfKghs+39xNFC7OECPAEA
tVvoqDxKtd+jOvGIWVgKXstf2qkZYFbAwuPr6IszdwTDJU+U9eSYptcUevmqaVC8CKUwwYn8RYms
6SZZQIz/VuxIrr0fVm969L+c/KaH//Ljh1crghtKWjABnTLnpuVcuIzBgcg9qt22JjkjLaYm515I
lghxzypSYe1fQB6q9mpSbvvUHpe7MBkYGdL8uOiCPvCioztPN1Hz+neg0gtPnuS5l1eLwnfj2TZ0
mC6GiQa0Rms7q9iAUxydgLQpNR7zgOgiASqmgcxtWZQuU7pob4EydeQemBxcnZ3vwtnEGbBuNWRZ
PsYMacqjPDxA55jxvSP3H09sOjvkas1C4dkv0EmBvlEZTxHjz4TxgfDQo03N6oSU0FVnMmmrNxbA
WjSwdn3xVx10GXWKe4yn6d+jJB8Nka92wWROZkfpW/L4cYhKK8l62dMQVN2IvbsVRe+/6l5ywPRV
4d0Xgad9/7xWCV8VVVMVIeUkBJ3M3Rs9uvw4T5m6jHS3TrRpODTyW7EKgNPN6qwhnF0jHg1MD+/d
1l5pDhzflud63IjfTAE6m6jTIrVfW7Sgcto7jYHbgatitRV3FJsQRFOsVeQ4hBP7IMAhETz19iUt
G+embMWmggFTaLaLl7/isb447kuPEyx75qOK2tDe2ZZgTqYOMLkwYc+yEndEmYZYpq/aLzolfVZc
7lH2ANvZbRZN8vHkBSQ7Xwks8tFKf0t10pb89+cpg8qEGFAf9UyzPvdUQZBtPmLO+jspdmEAn62x
4D2lKr0Y/WZrUv7sM/+H+NOhvZS0achDWXE6n6hMpp2GgHSxqhLHs7lMrFXs0wKb5hmGlEvx42Dy
oalNkbbupk2jCAAM1a991E20TVqgeszsS2/Vj80gwiSz8fcP3LJTJMDwiD/uwRFK9cueMMuFjATe
XxJ6NRwVIiu4/JDRgL0Wn6SMPapdjcN2zIj5M2ITR5SbrH3ljNcBWHJ3d8/7Xri0/DEBE+Vau/cy
rG9TmMzPKzorp5udtwBTTUm5CgcuCCMhhQV0/n9h29haJrPFTsEiroTdUcP/o6CoWDcChMAfJRAy
w/L/+LwUslGg2U7/mxmCYwHGhvZqr+DGri+4iaAIjeF38Y8m7gQUvdJxkLg8ZZrNZahwqyEbtkxo
OxNG62FKuSQNUgLeAn+LYBRARN+dJ/I2mtZTFvrqfC06veifJCNzGNxn8MqjSomuP+FTQRJt1lKv
rpXVCyqjFLuWn+SAritelHK2RjXSQoV3RG0BIqi/3DJQ3c/jrij0zerik/mTgK7o7ZjNdJTL94pM
wCMy2d205IWiHWSfgkOoC84uRvXXOaoMibdDu+XG78pls13wnIBwznHWjMCBamTDWSwjPz9L63Xm
uhiZ5Qawj+rUTyUx9Dn11O92mcFbcJxNpamOO/uVxbfCXf/2BoCaexbtF68guZXBog8U/aibQLNt
dULwF+7VuVifaBeLygDhHPqUMbbM3pmJ6nfFTplAqtv2fBUM6M6053no1ejJmaCMb4CJLoBVDOYc
jiRaYXf5F5Hhnc3Spd4/jk4RPJKfb7v9jtgLCq0DHkeBn9ilpgzEmmfqMg0dey2Qhv5fGN+zkGYW
tcv4d7uhStfmg5D63JpJy04CrN0rHC6ysRriZhzwz75lHjjsfiFyc9QMvND1/15PHNN31bupt7e0
FTGCHo0wBDPEbe7IY1qzhBpeUkmvYCuziAKPAr8uTajWKKeRIxz4ttykxWnyzLPMGONhcuqI8os/
H7zYd2upB9vrDq+kRyRxCQKm6Kv91Rb+muXR58gkDvihQPggQjFnZewfFPmZiyXThLW/jGC+eDHx
pa3f82wBOyl/c5BAlS0DRLgFQCJ5VIUQOhQWysZm3AfVHzfqMy9foYKN4h0Aw7FQlu9dd1L3XEwd
JXJ+9Qr4AfRpBsWks/m5fjEUveWG8mTDHMGMR7zGgcooEGavfh9c6rkTlGgCMX0VtfsiRgSVXWtw
rjVsipxxNe6JhZpXTZqi4huYktxOwXJGp0T+8ILFX6j2P8cGhvcGlNT0iE6V2JqIiet250wDihu/
Oi7jNLj33Mh731Fm2fTIK7775CCrpzV6sF0oaC36fBV9lsXgkKuMH7rHnwKiKYmizCzoLmz5yHbt
+UJJgkjmWJJenqXSsYzfdQKYUXHO2sQlbeW218+axuLMgxyAV0y9ChXRW6blBS6v7aXq+Wg/veBo
eeGZiJCCA9HdWOcIWXxP+g4qB1es6JgpMEtzTG+HQgJmFewe5wHMaPf5ctnx/Ko56dQ/8RiXbHfg
xA0w5Jbz09ig1sMEbDkJtiXVTHEsx+QYKejTjlZHM+GlFIAoOrqkAfzss/9QtUCOCGlAdqcYAGJ7
OW+O2iBBDOBubsZzt/oDt2uUNwVX7RnA6OHqxH2vGGDUsnbZsGqeiLMIkVQwt0zb7xw7gvio2iWy
9JuvuoY/ef8/0DRsqjrDo7h9truEkJaKv4sgUvttUvDMMLOMHc/CyDvk7GBnmu4RsM1qlKwhFl+v
s6kZ3vcTwaT/K/fPh9XRyMCxGp75fiJtjsir+tvSfCx6lsb1ljDB1pPj48AWzQv7fOno4vDNyXZe
oNHw78gQAP9n3nBE8gMmGFtDUfLCJRKD1EcUR51tIvlKkr90Psewk27mNJY6IBLLqRBRgtWYscl8
nk21OyzpP2HpO3FE7lEAYibHi3y9cjHzU7M1JF3c12jU9nSLM/K2F7SSXEuATukAfJVVRlLAJCQS
uOxh6aLEwPa91exOcju6Wj2YGK+qqtp/j4TuL2R3/KcKD4a/UgJKKtapRAgOLS1qHe9RmHvxbMtC
vA1SmY+hKy7gynbJ6ImeDeAZymE7ImZK2HGajNXqi4ZmI7tO+i5ePOKcKHYtK1J+32fmYE0kzat6
2jojhUYH6LuAIngf/uk9nDZ05SQsLOzd2qeeVXDojGcDZmfmyiaTRKG1z4gjp1alr+/zY6W8z/IV
e5qGr9zfmcRGjdfLhiizfjRRpT9BvT0j3/rRslRYj68e/V8FVxdwhnq86y5PBrbRqYSXDUNuKtVI
hPaIOQUP+YJLDwZ6LWH9hrsGoFhs7Z0/K6R45DDYyOo6i/ld+PF872T9X2N5aOljfKSTiUaLs2u0
RMG9M98wMbh/y27MwY7IPzSJ0au3ZZZHhD6uWyIerb/R1lKLFCH8OysfhYSTcHwfbVAoNPcVJYhl
RM6czPIf83AErUdBSiibGH5+7gxtnwGtoJgJxNV7vBOOko3/SfM2M+Uc2TWGnu5DpSOdGuMe1ypI
pQ2NcBIxUnNf/vmHyFPnyaVSDEuQ4eFLk/bCbaaoCG+SbiM9ui1/2SopWR5QjXL0u9pd438Pjnv8
4wW2Wwz5bNrrShYw/8UPYseHbPkFQjugeE7fJA8hJ7rFW/bHM50VBEJ5WLcomhTqZY/3tjYh6U63
ky3A+03CuvbnIxxVpR+GTtr7T8CubT7c+yYq0WqITPcBZgJI5c9vsRvOLICpisJkLow4b4tILcWD
7k/U/4htkgKmR/9PGp7NB4EOSM9t8rZOZ5S3L/zSb6iApsngSi+a2eoxfuFT85/AVuIpBXMqeHGe
ZQFc0wvgiw5TV7hHYjby23Wm3DsrJMliUvXKOG08T1yhvt9zUiqWFaoLfdZj5+X1E7H3ALMhzYO3
2Ados0Ozm9V4U03LlEanSrh62lC1ehqgRNrklyb0ox1ikuDmwu7LE4oxCdRGrWgK+TpLWuokPqD/
3Ck0rWSsPINTDTy+QwQc52i+pikSftWL6KiesPrE+5ab5ZNeN97Vi0cNIkzQkn8ETuXY3MArmAM3
BQe6S0FeVtFRd0vtwU7hlXYnK0hn+HRsFhwgMNepbOBRcnusWvXxzvHWUYFIR1nPpq0dcYsbMLAz
aRDnCe6BBohQEWd01MljW4IwAPG4PnEVfMk2f/IMlCVHOajACdrZF18RGIAjaeHrNoyVNIvMEuRw
XIPz7wMFS7aGIYW9MuYlufxulgy3agKThyr2n6zpLxuSLqwN5W8xod4Ko0tog4JkIqadEzreyW9w
IiknR57FcGjzC+BrwVOLgd4buY12y28zUobbHkK8RMvuLXY9z7uycPajRYlf6l/mAxpE9SmcAugV
l46rLG1D1nSYa/xt1yZWmASlfL28kbKfrpP1Xj80tn/rcFMevUYk11dTS2LfS1L+bADSZFL+b/0c
bmWfjeFiuGofta/zCAJ4Tu8kaHHDx608kDMVqbNDZs1fMy6bAivfN9HbtfHdWiXU9bQIb+hsh1+y
W4Rbhb6DLEeoYqHqMaoSLVtRdfuE7tfR78lRkk6+EZrj57V8/RldbDlEOv+RrycNPl41HEORAm3F
gaDnwf46Gt0XvxqayLqQI9c2tzCS4+++N/3Nhp2bssjz4SsnOYt+kkRZ4jy0sPweyMvpEPx/hyJT
bgN5ul1QAPkWtFB2/ZvZhm28NrsRGKikg53W32JaExZPEEyN95DzZKWpv7KeH5NCITWSIi4CkIfx
41AHSGc5Rx48707bLrp13oCJCqKHCPjTJRcRBCSOHz0nyWgSIBnGOvywGVMEWeT7npLMOfHRJRL/
MOrpOsAFtP2EP/xT1mY1jASW4nWGN3JAtIjQ6KehxJ8M7Dw8+R+EZcz1nJxC0KfSEFAFyEUmezRq
NiAV6kzL96wtylLdn7d2ZyGMKWPgnlWbV8ppiHeVNxV7a5gVBMmwNV1GcyOjHMBMT5YpxrMyIERX
NIAwz2ROsKVlr8Bd05WR2810lRAZzfa04rn+AaO8cQHABzevWalk/re/gLyy/OCb5UhR2CYNvLT9
7M7mHxm+pnCUEub4BOpN7xQgdxv9rBl1crULxDbhlqJJBvaVNi4CPP4KSF6BIY92ay8u6+Ellxxv
6d3UeL3gOccSXDvhXCUZkYa2woQ3XvjyT0oFqzk+iT7pKo1hnPT/6BXqm2lM4LAI9n2XaYsi8U1L
A6rLrMZW/LW2tzD0zHt3e/Ruk+n5VZ9aL8fYCLtcI4sPqcdSuRvJbLlCtPh0ybAg93qrjdFweQZp
7yh11iUr5FneFeK15JKEYn2xCmQpJ0GMAb3ec6TrTX7zSFRAh0KH3FnCij1Tyx4do+dJL+j5a4AQ
Ec9ochm/86O/GDmXOLZt9M6Sedidvu+m7rsUP2b7lQvKTuHHSV3RY/yZdaCWBj+lO3LmDGRTeGMj
a0BioJcsJHSOrb1Zxk3J9sFYDiymAnXhPPcXwnC4sr+k4JWCRStqXSyfXGSnlGXbDjbJuYUIr/Y/
48jqRCW1uytXMgi6XSeyWVYZvaAps+29ov2+kOBjFgWGmFjIPNiSJvP5CEPh1UWx9WHd5SBJjNOO
PlREL+c6Gar2QN9J5sDu0/LjYHUEeKHwDqtg6tYwxjcU6MmzaNuw6rATFEttoH4ZMUGN9A4MGEn9
fk+BYhcmIhwlocVElVy2y4Kf40csVeGJ2p2yIEteMWh7MZqb1MHJ6yD5ZjeBJk0np1ic/W8cd3R1
CeBEyFkQWqMPe4Kd8BA1eEVx3J4IAN5y90jhDYaFbkThHs3Eh+Xaarqx1h4FTu+gkJOszPwAy9cI
kXloTiNgKeIUlbopXX6mSm/dPrl/cokspWXMWLefYi99fKvEgedaje657pVh28D48h4hcauYdECh
tuw7rLfuWpu64XV4QKsXtJGb7HHSf5qLyxQlqU+G3sAt4AImsG+e6aY1xeA8Vukq3uz4+XGbfBH8
TfA30tzKMqOh0Ju/x0yFrTLDqnj7lxiTsgV6A2NbBxXwXxk5UVommG5QCTxg5pCkqsFKS8yJ5+mk
L4X0yt6LAunZb5OQPOSbZfe8D71Q7av1rigfj6FKP7OWDCl7BHl0+QjHRB9dj7gBZd770JHY7Ugv
eNVJ0R+YVTm5hqU6ZvEBA5h3UI9S8k+B2ti5pCLQCy5vmsfjkR00qfxTb/4YTuq35CmRXaF00581
jmo2ToeRop3o9tcf+BwRNg69zG7y0BmLfrHAjncAKMVO2VYaLtc3Vo7uUDkqM9UWfh22hEy7iuAS
7J90+7ufJijna9uT2CsvvQuQkCIPEm5nSH60A4ipvDiTtVjlWha4voeHfWtJpz4JkNxbJsYjTBSi
fSWl4/2oiLv27XLRKnPyJuAUl3IjiO0hic4M/XpvBFBtQp35mc5WCY+YDolS2ieXUs1Yq1p9q5Ga
X/QCVrDfsMymNGfuw3oH96ITtZTY7IXpKjqSqSsZfCcWQQK9UTUA4lPn2wB5zc8gPAMqAQJyHt5+
QCyK6P8lXzyq5rFMUKZHdbktX4DWXOydSk4yTkZyxUkdlDt4F3luQHFjRlmUeIgluE8oPmfr3Tqt
kHGSmPMKU0fhG0oVaTiQBzkXmkflpzm6OxBi6pGupVaZetE/SXRt0acBnNwOdVFP9SJcXKLiOMKy
JJ+iDSTMSkoWiUHaPkWm/6oV1113wPr6k52c50/A7NtKbqRy1xnGI9tgShCY47gMcr7n2ZhitJ9q
ux+LlhvN2/Ev5ZKXcQ+hzrKuB1FolWtb+KpJ+wsMmLFM70ul1CJB3//6BWT8eMObrtlOsNX4hkZW
zP0lF9BS9wjB1ikJ8FYTc7a2uZrrpWdcgxisOnPhWTqw+NqzSy+y6s4umnoetBW6qhZGVE5Rg8tA
j21R/usLP1HwXQHPXPTEey7Fsgfbmr1dFUvFJiuvPXV2dIlc2zxHI7bBHObfa3b1OQVIkjt8X7G5
enJKNqrGr7oU5JVTkEm7GnEs3+yoVDjOwb4UdMNKp0MRdWW/Ivv0UBR6Pgu/j8gOYgE7DKtuy7rP
bKc49NnrzZfFXeJ9x97SZXj9a062OdxqaWpWPJusihCY3/u41jiNm714AAQmNc3odVOr/pYxWAD+
dYcpz4LCxgJvcSrVl09n1ZUWvuUNAZJ6oTWmTK2Oxqxs+uTI82HPAycZ7SVzNEQfxvTq4ry9RMez
e9/2l+CgxgkfvMdjy51hhdbRkeAiFpED1UR5f5JeD3NGC5Xghpypc8Z38+WH0JkHIwG8/KuBVzw4
CHDkKIeS7I8yhQ1T7YS2wMYt9zlcPn4Gu5vwTC+jorqsjoSN2ieirn7pQt4sgK9QeQjQbeCcp5Ez
ANFe7xK0U70GNVkdvw7D2KGxYfDJ4oJjpk6zVm0K2xot9jJQhgPju8r53Z19v2JzM3K5l5Zo/5sp
9qaDy3mIZXP3y0WuUY4RvQ0c6TuZ+GfzYOsi2O60MdyO1EHh/SIsc/8UsNW2me3b2do6MMOXEcUx
z3nHqzMmw1O7av0GlwnpMGnFUU5vLFXdb+07MA2CEqUnQmGKHfwOc4iHfXNL2bghZdyrEArXJBtG
MDsYm70IG5la1w2m4n1+1Wx2HRTZncGE+m1yORGMI8FXm2HaPSsHpkBrmYmrKc78lHRAMRhgQZIt
4Lb5vJz9cIvWcadU0/ZGjRbQcP/zRpwfMiOW6ry+xkRJGAFUjfL0TTWhq+H2pfXTtfw/mCil9Uuj
QKdgChi3+5tBmOvdlU178vp4uvig9xoVQAOCVGIf7DTlv3dThKIPHEkvDqyufegADgwqu9annKqg
CeQ9lIiRURpRge4is/vjMSEjDYeZh/icMQz2JquoojosYny9WY9QMJmtIL0TqKE71fdN0NNQq/97
vRvgiLwZ960x6DiDsZr/GOWEJYe6zXP9TR55WysMz4VLTtKNGwclepVu5OEeUo9B/UKh5m6nxrXP
XQs/d5DbRcG3mV9ru0MlF6Bdp1jpI0nL6AcjzhhgUtWVY7LdeW7TS5ZnrurrjuUJuBcOjeAL3uou
Tp9PuR6pGyB1ndCUFOQEcRaJbRcXHUhJNz4A/74j+yr6z28K9diVd79FaEMHBDp7AZtS1pKNfEHr
+oaAg/OvMHu5wppIGTyPAcSR23QAWWLv9Ow6xlsuM3Tc0fyh7X3sioXIGOV38VZSjSOyDPZHgQNz
zU7EF+ZctcJz7B9txQ3cIwUeTrQh5PXkFT1tCeKLVXunbmmEB3EXLu6Qssrlq7WXd3u8Yku1ARIf
uogWZ68PYxKCIvGSjUvbayMflhXPRX+f/bMowCXgaFfyBq1J3no4J6vTyARW+/qnZC0G+vr9AFF7
b/QjGQ01i27GP4OivmD+JvUG45AJD4azJDRB9gTSLCT61fQleN4uVwSJwiB24fT8u0eEgsZT99qD
/ZM9vYs89wCzd3ikKReXRaoVUBPK7bruG7bW11NvKxWZkgS/v+lo2ub4SHBlNlZLVzBgDupySRT/
54djiRsC+EuFEY7jZ8tSo7AknneeuHdqFuHSCf3hI/gpKST8S9yBkdK4Jk4XLpHNVbM34iBNxDP+
0NmuMXd7tJpRx7zUdjodJsYPtmF97VBpLHeo2bik0vO3Mid1Um1f70rPU1OGAnk1Rr0bLOeQRaao
X813rfSIT/G07ErcjGIk9Xqa7xHH0v8JMLqun4tm5qt4BJ/+v/XsneuZmzPIxfz82YUdnyWDU37Q
w9zjUml7dJubbaWuQxK+98ZDkWZD675Y1BXixtt7Ilr2RBPVyXQMpnJLCT/ZJ0EeyEXPCQRWT7Fb
wTKGuSVelLTgZy2kIn2J7Xhr1cEjveAoIvM/Ad3UtwygfTCoLyUuadgLKoElDGPsSF627ZWUjHsi
YwnY9iFP9/bS702JV2+nMe2aX3oeu7/ergMyoQmBK1Zi2tHI2D9Fx6u6KZZBctQ0cxiKTmQT0MOZ
BaW5WCIM/SE1zZQ+mXPXTbY/FkiKUA3wFq6hMBZoHEhSgJoCMQ6XQ3VzRYXY5T/DF77fvA7lP9kV
DXROzphKxOn6VBSSaJzafFD2lIHo1plQpFgwF086O+4QCh6fjYa9Ko0AIUOXPSCpPlhXMdfOMSZK
ITdLa2rUv4RS4cI4OehTP4Hmerrolp94cTRF5jts0hrcLPLBBnjDbtjosk0m7G70Q1oRRt4aZ79T
jqhn1kKTtlf85Spg04zANY8xoS2olIW1UwjvGpkehGDT7fIR6ZWWapWw63sWRpLBGqgQlEtB7SwD
tGA6wEVSf+/zp+4yxuh3E3Y0HaUGIDWJdsZ8MGb49EZZ5Ap4c9KK9/S0s6bvsy86Bm3tgmQdUY8W
jsUlIp8DBZrPRigh7SPrc1KwcOZCSrOKBQoV9tFwHOs0qp7i3VA9pQVY0SxG5SUhXi7XTolzzGZ+
6JD5gcpAe0na6MbwPltvmrG9BSuBjk+FH0eDqVfMXw3qyaNQGKltlzj7si3CYrqBvEu3E91ZbCMu
zzi0vWkBtdmDQMnFvCK+vyovhSR42CXedWS8XWnVhTCQ5AhXfPtS5Sg8BAUhyasSt/1M+dcqyY9U
1MovPkMsYXhTDTTI0o/R4XDwBpdR8jet/GPVedBIaGAp3TGVHuACytAEGXgNZ13kKY6OwOIAno8n
DSVe0emw3ZziE8BDY4wsvG65pTnDmtqqtiou+DVl7Kzpqz5ByU9k4xX0+AdPB79BGhzLBgWwlEa0
Tn/3Z1ekwsnDZz05R/ZkDno9GIMsE0hOJFzhXnhZnsY5zew/vjMSouA+qqO8TEG3G0STHUuAMMiB
qdKeElH60QOpXvx2tGVptCMx95i05cfmSc1wCY6GlysZn83SZ+Rd5sz5+KFokfRO5SSOYTxOyH2c
iALnDuDWrVJYWz3mTtlOtYGo/YtknfEcR2cLcezFfQ0z0+uk668pD7W1om/uxCkTRCsdP1XYYDU6
U2fC49WUS47hN9U8X4rbpxVP3lL50zdUtwBiLIsiuC1WUks/T7JYtKkvd2Fy4VWy14PY9e/6MjDP
LjXaf7k/duTTiP77fGIP8OH1vVs8MVL8LVDyh+tpIBqfOy0ZoYKd2vp3jEIo3bcVBNlIXW9m94OS
iExyO/ydc6S1w9Y/8L5H91DcFljuec3eIhAWGbtrJQeDHj6kmRcR/lTiF38kxspQRYuCcxV5BdYR
QWi7+uR/qESUur4UXujn1n8bHmp8cWxe52IoWG/QspQpmT+bukP2vYtapFijDwpiBND7zkiFCOQr
hKxaB29av88sjWmQUSYKS6yVZxrRkQW3oGfyQJRAJcxF6gVzJfPQd+KaeIDhVuv85k7crLfFmWfl
cUgjd/7YIJeVnGcjxvpKUR118dHBKjVLNAgqgRvyGKcT6YPFXygIahzQup+KqZM/o2D68Kh7ZnYg
wY9wkHeT1j/Z55cqW33ERt19nPQAXpiqk/j1NupfJKitEc7Sh2o360UtK4ULIQkS9uv07y8e+0Eb
QKvwdUpF4ZNKd50D/LVeRdJQxihhj/EOgFdZeypmjAY6cCdj9yHZw9v020njyurw+kKjfPPf2g/a
ljgi8hHKhop7GKbYuNly0Anw6NaBH4yAZ/6Nft3GQGVQzKLdF74/xN5KZ1i2pUSkhGxbqB10jVM1
qyI/baLxYbtP35v6qaEBxIzfS2HHhUE3hNidD5D/eusSjr76A/afvq9RVgGkYXIhdBz4EJmCyyQq
Fx4IfRXpmNZOC+sN5vMumjwdNNjvhJZkmclkBtExv4sQMb9EpVFhtYG+ucOFTvJhmzF7soP/wJXE
EgsAy+6jjtXbjpXDcyfHt9zaVXXv4jLFaYpUVtTEquKfuarnNW4IW4+Wu2+4NKDWTlnPgi60/ygP
q/3x1VSCuTVIT1C8CzT5BB7GqQG6iXSg0XvorI9a6i61PPVOF/0CvxOdwaGEm8FeDEPuwQzTUpVA
3mfF8HE6BawpA9TeV0tRLgJ1PU7LWX6xFyCS4YquE3Zd2hqGMSMc8fCvudtAINSZ4GiUecxOvduT
BJaDi8SRU3R66Dnrt4mWq5i6umOC5Nc7DN8tLTSFTcJ2HpF0Hy42MOzosj+gH6sAB1vPD4ZVHCV/
OREnmCq8ESzYnOt5lLcdpQ0HNPjFR7VXXqLMK5iDnZW4MTvEPTLeYYnN63plmtRNtYwfD4fMXX0D
LydHyOtowtxCxOyGksySPzgLATfp9T2rpY9G9W+H8JCiNIJ4OUyNWQ3Y1PnU5YcR83u/kAU/PovQ
iuhF9IUWCKUvCKJ5STb4vTiDFO852KfUdGKh9XTRzZwe4B5Fp4iJfoBmoyyRTh4AjZJL0pEHxYNR
o9bjiUVZQsoEeCZJ3+dsmgfvUWMnJFSc9btTjta30THllQeIFddatUw6zZRlxDa8wAKZXZ3dWu/k
ZsQc+ohfsoqsb2yc505gwgZMFA+59WflyzNsf67ZGiNdsVk4IifcPeDuOLifLOwX3UAplo4prJYg
B2T8fBxHjGqWPAoEtr4tY7vJ30ugMZRDiajUpuqSmWeJhQf/yjhEQ8/PXxP4RW30pxOcz1eELgOM
dA6bj2ab+jWj5pMx2uHsrslM6rcGrx/KenEcO/bVtTxjJX9aODSzlh+zDe6KefnuAmVFqK7ZZtu6
B9Ut04YSyU5DzVhon4UXzEJThDgAeF/STMdcZPNKmswqkuE0Qc4dkvMBG5cqXwe01nwrXizJ2RXW
7BVJ5QvWYZr9dN8G4JIMjxKEs0YphkKJlUUX4HDrelx3xbU+h0r3w9+J95YbLZdxJwgDlfHHdxms
Z67+SKXLpoxtRarkIAoR6Khd7qvEITxDotdFGo26Pr8xV/ppCteqDsRfab1doZz4ucbDrnVl1sPl
qRnnTwDjeY1HKqck6Hy7XFqDyGkZVkDHHSuH9sMA4nV9CzusANp0w2joUo1TdEMW/hRF5bmPasrL
kqOf0e/o6YMp6+QdtRJ+EJY8y5jyj9CcZ/lIc2/jJcoRJpackF6NbiK31envvl9TFN6Z+JctDyfK
997vSvlEPGR7DCmrLwxzpb0yP6GGMI7BUzkl3WCcrF4c8ULAxmnuz3QPIk5tOmJ53CNfRCx+9oXN
d4hGybB6PPUKdym+Hf4m4Ydy7C/vD+YGhNU1Q3nISHZBByYvRmY+bgCB+fl8Aop9tsSaV9+QD/A/
3gkmd+t88lOyaAElNZwt8PyeIoTQnlqGisWWYxJBbG0z1s429J4qR8BlMXmY2uOutQ/r8JfIC8Jq
L2YS3IMeUMCAFY3sz08ykEXmrRKd63b5Gydi8nNTLo0Uh6qhkAsXxftpR0qxqtdtbmUPHeb+gVdM
2LOBs+0Mo4oz/YKDeaPYgjhELy2/H4ENp18QsRkeJDzNiG8k3eB2H6egAUqlY947IFXCSkz+5Lp+
qhCyZI4utmPoyf/fCzfsIMgLXwwZxDHnmdOMi30YeSlViSuwK8+TTSzDjdGCIfumhGy1EtSxhbSk
vXvC73KcL7EgpSn8kjLcdjgP++OOOv3fZ52OmfDsaFz/QTXllaBnhdr6EdXgLXO371Mm7Zou0BEt
8NfT8leQJPb5AZ3wtbuuonSgZmMbdCYBkwiFqDs5soVXnTlnf+Ec7v2aqj/bg/YYMJu0v5Iu6FoP
CmPhUSJKZ8zhIZAtlM/8cpVPVtJlAac+bGLLoDil7bF9DiP34DCsQQWTKIfycpxPc6x9KoU0CXy3
a9xV1JuJD+SpW8xP5dTFJKyIb3tQxQPDuynWKSBS3J195VC9N7iAkxPBTuQ+OxyZ6S5DPfkUddfC
QXfCZ+Nr+Y/h7EmBzIbWdurq5/HuKo1bBFlHAmIDsf35QTyr0L/cvDmI1Wm8ImxIuZW8MRBhZf1P
zuJ2nkZol0e7Co1zfrD+3Xkmb6VF19dNSE5EIIQJjhiBbdJ4lQKcrdVOlXCWEPqoODOxKdwBiBEK
aqpkdyX2NcNETnDY/X338gkhqJtQI44JpksYBdv8L3Pe/lYElftt+8BA+2rrc+MaByUBHsHBDEkU
VJ1Uo9w8zx1500vDv9o0uLB4RI4IjQmbn89EuonreWSU9s7IT25jwILnyLMHhiMjIW8Jx+4KMZcg
OTNwPo6TUudaqU65cGKn3MjYEBoPQ5+wy+rzsD12q/UVi0b0IupxcYH+pwHVEdGK5MZNi5oe2f5T
yvdw7FHltnWTFFPzplCcHL0A6vF7aijNAPwIpSe9ifDEpuRilZpZjT0Oi26T1dzV6tOvcY/VIYg4
K7mQ7ImWpsS2i+1ouLMpBrZ7uom3zNFx8KtaFZgiDg9aDwERpRzQ2sjb6eQlteaYBPZuik/Z6xJE
SFO/sSjexDjzZlv7EmsFAV+ukTECjCqMFpB2CF/vu1ozo5iR2nZPtbXSJsjznlCyl3ieNV+Ir8W6
173kP8Qo0q6lv6WeXrzaqCSLDtn21XqTo2sNxj6UDP7FGKOS3CafmPr0JACXP0rL1Lak+9/Dka4v
2CoOZni8XJLGRkQHgRKaKjXgQpMoAaRWqsgsDOZ+uBpq/0/V5GFZ5TAf+gm7TKgTgSmUKwvgoJb6
/DHvmO/vUoe2qXStndfM0wRwIMgks5dy06b/PbSNo2i1804E+Z9g9RCHMmtrgNsA6XzIyV0Umotp
J4WvFXQdfoHIL/kw7GzutZbefItP3NEYesPjvFPjEfP8KWBV1tIa5dn5a2/GCWmWFDDSHNZ+Oa+8
2pCsrmu2mMALP+7Rtp/0NBzHGoO7uzzGm0MmQuTl1JWFpDW9EU8Q3WltqIFoaoQvG6+nqZDDVUAr
ODpurRK/SU3SBkJk6hgfudgbK5tskk4A+OaA7JrYagsUs2rPRSqYqvI4p/u6HoYn+9EMI8/4gzFl
h/Z9qOtTyk8myeI2qC0mFJNLc39xVowgadtrvU1Gv8DeNA74Ngro5daKkCQRBa4TH3X8UaSB3g/F
DFSq6kuidMgAZWoE+7epxO4bExFgVG6VgMxG54Tv6dArTBL4+1yYb86JY++tGOkMq++dNJvqqpXS
lXyl1/Wngs8od0CeNv6CCbfONt/hGQ6yc0xKFDCfB0oFWMq2K7oDC2eL6UX7/F/uJdkpSGcE9DWB
OA1v+0H1qqbzTndgMYF5cgVC8UJfw74lMQwierH86JAlry+he91+pdQVTXq/0YD5IBxE64zm72em
J5L/UkMRrlCKQt3fzxOO/x3wfyiMr5Es/3C/doKDUiTVV+L7089hmKoErqxGs324QkSdk58bCnFd
L+13yDQvD5gOYx7A4DIN/Z3j7oQghWuDZNDDLPvIcDZeWqQT50/T/fcKBuI9aufuB2WpJvC7S8kP
Ti8WIRZ41Jd3ySCG4+PCw5ayikCzcrdPxRDMkKE4wN4JJ78VIp7dJYhqND0zNaLSqjb+tMzzIH/g
zQ5Dqga3/oQ03J7gEuqvMXK2szNnnruK7R9YrtGc1LiSdKXNnqnMlRaNQw9h07EPWicjocT8z/EG
aJFFXk2vAeeA1vV1hXxftlXl63lA2vkOHh7w+1AWfNOh3Ib3g9/w7Z0LAx+cggxQWuRSQ9VUk1xz
CSh5YphUMYHpI8nebwa25LoNAPnumNxu762kySeezBCj9ZyHfB6yIZgsHQY4pRgcoFVR9Y8xnegI
v3O+hgdgRuV9cBhq8LrLZeAmYR7UAaTOVG/RBYFrb2jn0PVmXprTmcxu0SmZ47sfUe8979To4pfq
NRN1Nj9U99DELjyeh23ODJbcw5tRwznXiwwRgXgflyjvClxBwkD2wlhflNYqTnaVoQivH6OEDXaq
SyeMiOroLOwJjEsnAi/2XDxHBMbK9k92lE0B+sYFP8QLINQasuOcZok0JOe/j+IzMGy/fHANoceC
lY7y9uIgrksK+HE96AO8H//kSBdWxUhERst7Clh57vcFosvBM6gqa7QaOmLdnAhd1GH/XFI/OGJR
BHZmFEX5VKTLOx/dfnD6aCfkCi69J4PZ64bV9OA5HaQ5P41o98xEnesyBr8gdaVA1QHOYGPal+fe
g+termelH3l9IeEXTUgtiW2Us9PG8/SUo2LxMqk//9McRKAUmiCoS5rl33uLMnYyjYr3AXkZsTBY
UOgHA2u1zaNdURsS3KDsmI1DUDVxz0pTyLj8SsN3smK1fczpGlnkqlB+XBtz2srpr5v50/A26+AA
MwNStTnPFcdcO9eMQspMLjg8REH4vmQrbYBiOQhSS7+QFV5FiF/WXE6Q7eKBjPi7d5AVwIz8YzMJ
rXFZ492icjKFEbnZtev6o1UYzO2fCnz4eDBh6znwYkjiOx05pzuHSCWjMzKHQGtn9amgRGcn1hxa
G6aYIuTzDLHRY9A7b+XE1hscA6VYVi/yAMpvrDAh7UN1bBva0Xk+RW1raK2PxVc0mgvvdGR3Q9D+
P/HYq6ClTrpcfwBbYJ4NJ5k0iuCVoy1B/4QldPxiK27Q+erPkZ1r2Ef8i0a9hvIFDw4s2il38HcF
S0NVDxQdAtdb30cSqPFvq8IPFlB37mp1a6KqSjwGZF/+Y3NUsX1v9ocCgNDfl6Wht7pc+6sewnHC
hGIYDHlfdzE/ciJVj88GJ6WAFJ+7yb9xCya4J0zgaTOC1JpjRcPWB0Ccj2uqbQAQbQE1d8g+Qwpm
tDOsjT9SsXqfW6SISrUlaaioPcX0TvltNvBDBClmIfmKYO2ApNnG5acDRB5dHUOhk8i1eQnP+b/o
gJNcXus4y/ZUHPfNGI+J4jfmq43cQ2H+QNsHdnR/XJLTB7QCeOyyHT1muBCD6UBG53x6Y7t61nll
NyJyzWvetCxJKXcV4QcnXIUUhpjJ5iYfei/AKu2JRUyxQwFWZnOTtIYjcG+VbsA6J/viuXu1HmGA
CgrFQtCh+zTmCTKAn7X9PWAAMPADtf+ymbMd4ibUGzFGWERcdauSqPN3cNJbEaUToQSPXbShQNzX
RJpnVlAlDMshLJnWgFyfGzWwfCaDWU0mSAoR07shb2o+uZfeFzeIfn3aBoSDU17aC/7dUVMlgaK2
i59ybmUAIsB9wLnU677foa39iFJ16Tp0cd8NPD0NTWYidl+MwyjDnyu+G7zNMp0cIZnybcY/SCad
3hoYZ7O0UsJBRgYUdWHwnH7i+DCgQQxDxdkA65si0kPOQbSj0OtJtAO9d4NsQKjVcAM56EmQOWRq
9IYNYPVh6OaimFwE5peU4Uk+WRlEH+D+IlfD8Tm3Z7Z+ewndDkfOb0HUh97DmNaXcj2WZXJRjFRr
IJK1sKL8FLafXcGuGHx9Blzqg888FRygT+ClZhZzvVuAnflI52kjRB8bG4QrstL5tx5g9TgXcUie
mgdV7fzAc7IAwPuPQWE1yeMw7w6mPEtWWzUThK/KuAmKSh0sGA9+KpgoQnY6eouV3jo47DVVX5ex
ehpg0RF9Xqv8s61W8zCByWAMvFAdV6UCs12bPLHS3FGsmIYO7aceUW1vEgAjezgCusRpDTmgnbh/
ZZ+NQ0PYJMSpFysn3t3IqjZqb3Tww1MC6y8IPcvujtDvBZ8yvEDEZkf3zMEoPVboChxwUW6NeVlf
SkddLoiYc+SntoXY/GVQURjy9Qb+DFK+11r6BZhXZlipC1mXUAzMyRx+rRmjXKd4PLq9M89hhHZ0
fc4TDXFNovP/2kzDgy+osvd7zc9jHJsZNcYiGeb1QqTcWTUKl+/U7wVgcYxQKEsQypTA7oiQwRIp
TJMRN7o2HZ7eBFQC7blfM6gXvHK0DiCMJLlR54ME/KbKG4dNqjeznqT5Lg66MX5wuhfxIrAQM1yZ
HLDUxo/qw+bjdeduLlM6//ZCqO9Tsd8Rj831gEPmypn1MnDo/J51/neV4pTM/pTU52fsjVCtR+Gd
0nYEIh3DL9nzWSz5ff46/kqCf8p5tTMzwIM0E/gtatEe+Kx1DCI6pXxuUHYB0E0kW0PcofHuMmpv
d7U6zPu6Wn5MMCuvn4Z2h05REoA9EFIFnvTyaAAaDWOmj1Ucf9SfX7qMVhfhOcmOpYZv97OyenIP
ysAXquCjpsdxz2ciHo7IQ5sE2VXOYeJPaCpml/YwqcD01kx9V+4vFqnP3Rrmtn5NmQoLv5FDMnN3
V1ygDVogrAvGU5ug9v2+nRjto2yeOY5NaUybjkP+benHX3ByF+rV3q/AqhGlV4JCmaBh5vtoiLzu
U7yN0Afdh9rscrF1evDbfUfK+dYf6BhGI7pdiiwzeykfJc+5lLfdzdyA5S/P5iCWBwdAFvIoKiQn
sm2Da7TPLNaPeJpDIoqIAHZRj3ZvOjZknmVOBEXcyjA4V9HGWrk+E8OQuYbbmEhmf+IsVuXqdsQN
ZOnF7RJrLExaT08oP9Qujd77UksH5he5TQgr1GHxMkhPgN+97k+QQ/X7KUXUpM2EKfiQTJI0xg31
MRN7rF1ZBXfEP92riW506EA3qugcn5U8zOkaPnY1Og2JVNPvwFhpxl/94aNkvb1UVunmm6naf4FK
rg6GgrWAbcdtmCElN4Mcu/0/m2/h8csTXOCp/L2adtQKG3WsCcs7xnpT92d9A3qzHu+XvdXRcLJj
0YMIRKpwslmW8uKDRu4EmxZ+RCCiIjEvOWXBgbZ0wQszQRRhu5FDsVdFuly6yrGUqg2tW6ji5QV4
sSn6bWp5hVv8bOrw6rKl+uJJaJh+hJKiJWtzgnAxg3kr4+x3hFY8N2YBg2pHgv78dCBIsBHV9Y9M
oCVjBpxuEmwDhIrqJTq45wFCnwejVPBZAOiXPbJJsAfEkqQbDtlO5C/9zsd8Zzo1nm/oJfX3wVbT
fe6ds4DnvXBHtv2RAcFFvQrnYR0pE6w9M9cYVAyyFsNrRm27cgW6hD+Q4+vMNly0Pqs0t/AKtpsb
1nkLjdrcBusqelqHN+roIdRDST6T3GQFBMuwkgb8FKa6JPPrlygFSHZT2a00WHJJPCGysyMXjtxq
Iej/P2PV+4Ce3fPNpp5dj/oBohBuuLYJGNrD9le+oAHF0e39s79JT6fvQv+INyUWv/CuU8JeL7vo
xXW4Pl7pM5NpwrdKZaJ5vwTW9kEy++S2GKL0ueuvlxmLZNaZQZl/sAflmtSXtyI4EbxqLxZnhPpK
JDs0L5MVoLg3lI3RIl7NxwkOIhK10rLCozW3if5eoQQBhElZFN9QVqWVwLlFeFA9eDuZM5N9ZQcw
fBmQabq6mPIxi4/+zrZCfbpbdSPvIbvH+5dfrdUWpvJTjt10ha8Cdldys7TVO3m2EL9kIg9aCaIY
rCML2rvwS44/ElS+r6Zdlsg0xBAP3fgBECbSqyHAy8BWylhTAyHVEPehuMj91c+5GD44zKuj95fa
inPg/txd9zSiO+3k2H7fJ6d6Z0/7FLGSih3XeNhx9+xeunB0JaHQYwEYKVkrKADR9JKC2lx4oxZM
TZLHswg7nwqHrq7ZN7XgcSRYgvDm4mcz+gS2QCgfaXOXkneA3cebq/+0NxjaAlSi04yjPfausuGV
Klg4AVmg+BoJblwbX41YYoUXLh79hGkrfctBGSuzDdl8ukOzN4H9jjyLBxNrHUiNY+DMM8p3klNr
jXZhX/lkLwazwZKeqQXyC0Sq3N7n2Zy2TOUGjQ+dRKLZ1R86Nd54v6wJPQCMP41BuG2H2E2G1bzw
2G5a10BC0qE7mvFdSjLKNXuQ9+yMnDOP1vKt6X/qN3azZbv99+jkICJOAXKvlBVtlSPzzl8qufzg
InqOV9YvMRhiNejVQNHQe4Arxa32PCEYl2sVmfr4taVJ3aUdm4L+DhIn3A9edq07XezdJQ+BsYql
UqKf5zvdODxPwa+jZMHw75wy+jYLyATypUdNIzKECHY/HwgBvjdW//zUaSSLFjrE8wlamjC5LQs1
234LJcD9PqQlbman/hU4AV2ti3m4Ex4fuEorks96OKdhB6RJ23g82WjI4hLFBiRJZtFVawODhmQO
MlrYBDcINEfiTV1Hk4K7xlVOaLKtrkkS0xyqaekcqERUfin/ad7jcrZQDjIcodjvrBmWgUAbTMJw
FZ89vj1yNmxlfp/L7wLGM6/zixSkzs2/3HG0LaAxBPZvSN70PLgpsBlQjjFIll47/md4frEI4f6g
PadX8WFaxbeglI+ZHtVSfZuuZUGFgirUyiQjAXMDZy928qekrzkt+6yTE7vmfiNKzSn1dZEIYqOn
lKMk6AZonpYaHzQBHTkn5PmTfFFMsH751GcPdH4H+jssxA3ayc2KQ/7dNNN+No0aGQMjf2RJiS3U
tj6IC6BDo2ioDU6JRKDGbYTSvMjoIIx2cGmrkyInuh38wz/Hu2n5sDB9AKu/8zP4gUXJ0PXuwgn3
dHw747WrJcYX7JxoSdXHWyzlp4CNFLlOqD6SDeHJzlhd+rYUO9+sOghWCb0LCDpE4nVX6qQC/LWT
CdTpRD/+Ck4vH7R5S+FrteZ08lLNf7iN+Ko7M/Vmq4D7qWtJrSXpzNGUSF2XXJN5nCm95/+6kiJH
EGoEh/+TTbVjHJcrQ51HV7GO0AsWhm2b6U56uvRn0NghHkRNFt957yIn5OoB9ojX0XtsPA4qKsWy
6FGA6X5zsJMWHQkwxZ6s+A2eGB1cbw43nLZT1arm5Tyt2HtLJHIc4ztHcPsNtVWB4pfAIcmWLFD6
klddGypDljpE6s2uXJLzbu+aNtYhTOKBp8O0pkj68hOgfM2UOaPrNlYFT2tBOacLldzvzgKBTXDa
VrIbba3ovGEdDrvzcJh41frDcl9oSCWtX2eezk1lDKexvnWd7Vob8SZNx8fuWbcnSB3aQMvgfn8J
y5T7HlF9dqffEkjoIASXeLaE0timc2MXhO9fTN84F7L3m2V3V99nG73SJsWYTXrnx8JzccY7J17K
vEpM2KwJouYEAM3NGn3IeYlZQMB4zJy1nNKfKAOwuyZ8AtJfyUl+/RkuLYzO91Gt749ySoTGvsOj
2oweEeAGKzOihNW5D6gj0UvufEp7GoQ8A5AO08d0WGI1V9O9FCwtNBgZ4WR82gbvATSXtzDkbNWp
rzPXO9Y+kb57OeifXcUWuDYqUoVEp0Z3zJjNFfzpqUygpIGLP+dnT4YSb4w7DmcHz5hozuNgywVa
f5FjXY9r0DbyME0u/WpECIWsJ0DiHhc5vl1vOx21tfF3uTcIEaN3xiDmF3/A3Ws3mJoANzcn+f/J
Lbgk93YwChglU4Eq86k9w+yC+rw1GBk6WRMa5ouoVXO6JjMdsOske92foW6EHXtvhUgaPgMrZ80p
LboN8DAzr59sMAO+nYbkZ+Olri/j4F9x4X52qKCMJuQz1MhiEHAxmVdVRjGdvFD3px8IvxUHO6jN
TBqX2quzcElFFMRO27vJA17MBPwO4ksMXWdQRVrAnoT+zjTepICiK14VrqW+q5ug2xEijUuwZUPV
dAI1a0ABMZ3EKDrPYa1tcVnpk7OqEhQjPPMTewcQ1IlX4PhcozIZWQZJofxhQXKyGAfD1cr0fpnj
0gj4IA8pzsnImV7ODSzB8jYFgb3avXRNF6z//U8mExIqHdHw3RymCiaAlHbpQs9j4dgRsB50aPYu
CHetuNbIiK0f27O8+n8kl6lCc/z5AdLCCWJZ4qs8gC3wDziMiRxHBdixm6/NdHk1I69w0s7vDTmp
MUjD7po4rGNMSuqcN3Vqvr6Ztgp3IzYq6g/2NltHQ5szj46HUEzMUZa6pkVyMl7QmYNYJunYlkOh
UaNBe1GGukhpzYpMS6q2ESII7cLMKXi9isMLOpYvzc6uIdIb77n5INYC6NSpZAoAREGTG2dB1dI6
vxJhAV1ztyAL0NRYcBcVDxqzci7amHZEKJbLpMQSnwg9FwR8ChoEqfVcsUUaeWU716mdOUbjDQKL
WfFEfP3WuEO6s0hgs7ZVJeVLBtbUXcb8Gdh60Xt0Dq2IM+K7FdSjCaUvM6GzWCjDvi7aQOYRz59P
wasaxrez/rui4FxpDeK9wddUZloJov2BmtopLipHlZPyS898j0nC3QAMCTEBuX6R/wCSjqG4Dp9F
nwteLpy85zNHRK6KFaeFmw08H9VZbWET6HYiqxMzjCq/xEl7ju9kziQn1O3hOhDrSDiibCVqm05D
EdyYQte4fQsVPLuWD3VgkSfDRmrL32swaye1pj8KNJ+m737UzAQxxkqu6t2QdiGzvhuVBxWGmSKb
VmFpMRB0UiGJgBaAsgKiKGHUhTJyc1RXJwZ//0VRN7/+O3lk7u8zwoqvM+ZU/jkFfr94ODGgscA7
wzqUEpGIFjWV0Xp2MgTGBAjJg8bvU9TLipJegLeOAFcnMclc58E82ebJ6h74wAklQKxVzmr93Hx3
LEi+lhcFNPLD3QZU6EHXRexWh0Lfi8jEtFnsVvTeSzc84Hw2M79eQedhVkgbFpZPlekq2I7+eEyo
hAfkkKwrMSrqr7tPAl+OjrUBjJpVjeHhgro3MeHI9g4e9oGEpoPQGGHAOxRzyERddNwIlA6ai2nW
8YtcHfWeyQ5sdG/bnQkJmR2Sb3k83b6TVebuN17UK1wL6M0JS4aFGxSVxcjgD9Ga7yaIMq9Ud0f4
9m45QFW44D4zpRjgk3KTJNRO5hee+m/X74o7CUvLnd7+Papphv4cEaYhh4vJS52pRuLXKFZVM3ef
UedsDKCfuzCSR0KBbpDq9IA2vBi5voNkzqEzfhHpDDZCzkQehbh1Woa+sSUbzSVS8ABye/QBlVMj
oE1n7ou3yJzOyRRPB5d5oe8S8vMgncnDyDn8cw2FR4WdibfeQqIyN7PztuD2Q0oNL93VDxF8/ttu
6Cc1UwJtWKR6FKXlmi852sgADbgIs+0692C2OPQjB4YfjfhPQAUBIzRUcd5I27NFwH8aCEc2HSoU
PF8ZEOjpdeL4JTLoiHrAp8KLMGEzSkSAZndW7gRVqSYu2ccfQgxUL7XW1+TAuI+bs+JEjXcJOxxR
+dtZjK6w7ijvOW2u8nEyszbN/Es9499g8t9TbrUQQ8/mskeXaB/06qUfFhijKWn/JPSrHRkgvc66
kWuBqunJCWhCj+1ejazwzMYNPN0oeHGkkgK6/YlKUeA0KGANeoJ9Vbkd2ogLqhAV+rfiXFb/8w7T
A0m5bpr9tK6O5zRqOwWf+DHRnGztNQCALVjBdeyleOVReiDFEIHqqPiGGrmfeDJ2f+LrjITSFGqJ
KZNVWk2kRJukSwKo6Vy+3EOnZqemp2GT3HiT3nBc5msvamPVxjke0JRyL5J7EBaZ7f9ZlKHvyGSA
02vmlOcqfCw/vwrpZsJ9WFTDU/Q95dKmWlZBB4cfOrmMJk/HfssdmpAfkmbaGKXvZkQIWRiwoz1j
OvFHFA5KZsaEfxZwa5x17FH282y+4seVnOpsQoOdMXLhRK+0ieO/LND3dUpmjYGUabTb6cO8CfcO
0raq3bsGymNahcLhcE7Sc1C9qFVXUR73ybomn9yIWLLdPCo/OEvBtoGSuQyTJXHbE0a8oxsxxM2a
uXaRBJWb5YBdTSJsyfkdiD8KSxfGz0u7M3xFGJTZsNzApotmID9XBVM7LTEWr2CcagOlI/vuAWxK
sKb6wQOEhtJ3LqF1UHs0MRYLkCeloscxtrUrdw/eOuuMFQnJmchTnUUPjK3M2tuBwJiRuJyHG5AO
AWz1fQEC973IvrJDuU2b32Do1fZpmaBlotJZ5y3nDUZIJa7GPsMx8JwE80GGy5zdbZmzupC/TlyJ
TumS0m+aUX91+joqAPy/E1TOYA7Vy7pnANQwXZfNashjFym0mFO8rCaSOEpLEqCMbCL+jkU9Ehw7
8Yy6O1/c/ZfXWmJXRMjXSY4sMtv0872kbQTLBEMEgyf+RUv6Kz08KnBe/lQIy1gNvRay/CJeoahc
hRIo59STEtijbxLUNyTDDxnXwXe/Xul5zP9dmGd1W19C2jY1HndOcWUTA9whbmJ6J6L1R5ErF7X8
8oGXHVhH/bSLK8nguURXdgW8ZqhK9DAIpGYqrsD7XpYNhxxRE2kSizTnI9yrPeNjYlESOHTLqM1l
pYinr8Qw9a95kx6VsrmQB5Eo0/+ReYd9bh/C1RJ/MbLrKv6YLrM7/hiFrnEPQ2aBdziYBTKqKbTA
mEZvfs87S2oywLRQQ3S3cWb5MDfS7Mg3MkoRv5Hf2bC0DDOxQiAJUqVCMgRF8ZaXFLSUQaWIvF/B
vw4po4fFQK/xR5UZ1U0SGZeL9Rapw0QbqCC3F7t7naRx6UPRI5/x/u1KcW13vX60rikNwbolBthf
2ZnvwefqlH/Ir8jS9M4RNm/N9qBD52nXFslYVUPchCs3ublUGE+CLOwKYivry2Of3pKCGr7hQhQ/
TG51rfNVRHfiyVx6rIuJ6CClEA6QFHO5Gze5qz4CKorwpR/0rpeEiJpC+9e1bAYb0mTYi1Vcu+zP
yoHgFQ9DxV65XvtuN4MxWgZ1amgph3RVGxA2hP42+y5bsYPtavMf+6NuybOvwvawS56J7HzwNUOt
b+gpywmVbL70J3ez7CPDWF79Ep0DDELeEud+yFIZw4odJN2F4NGfKOBqhx+NpfpOD2tvBi61cI0L
KCHmIQc8LFdDgAfWD2/aAR8/O3kAS3IlBnl0jnyLyPtJGAOOTOK+zZVvQP+aBFayTw1n5e2d1CIa
LblMhTzpn0ZwPOr3aOX5TqGyGTn1klB01cCf1AIpfaw+raOyWPIWbC1BslZX/5h5+VhRkfmIUOjy
ebO14/DV+i+URGn/lmjObv3NE3M4mbum4M6khvN2RKM3kJqBKMD7qCQS9RyZPyv8gpbL8ByzaeQw
rFERh7y/PO9K00eQVycDddX3Tr94xSDu/a0ditLgUsjPed3Mb9QjJ0WpCkzW5tKEIdN9Vd/adOW0
PBzZuixIh3KIdih8TaA+GC6cm/qNU40oFjVelWhsAooZhuaJOQo1Zilz39q1xc6PlxqEmiZhkx4n
CzkRAsH5GdbZPyL5aX5d7CPHrktInBmD1bahs0sA4NRGHkXdhFFsD6VKp0uJeetjc4my1LiD19In
D4sja4pqAJfuiK5+Zl7fKKsLbKsV390qqZvl/YyYGIqHW6Xbl/qxepa1n5TfH3Dhibe6dDiJozYr
wHa1wJCCnjijDkmwhmHApGSvCfgl+VHfboYTaicJ++y9k7MVmEHKyGtWxY5UdcsG80dGPRGuGlAE
fp/8lo9irN7w51+vMlLqIvhChfrOUrhdpCZkKc1T8RviWA418dfBAInKcDeVefhpQqJANbsqnBwe
WRj3/3tzMYCUSJDwtRisweMtx2OfEJuzEcA5bWQXLW7Xl8+MwYmr8ndkZ+zu7O/xWTgFsC9xLHg/
GtNDGGrIJjOhQnmeZsSL6mUD0etJ0P0+ka+VTL/0d596SKTpaRp7vMYqG4BCbTd+EmaZovYBTwP1
2/kwH8heT+H/8bQkK8MlES0SOfO0pj+JK+7h7p6nKzGrr+SzSN/51spb7aum7uoeYR3u37rDiMd8
ToK56qxQz3cvxcOKAg30LqGivhMlRQOVCwU5OUhKKuXIFGT81kcdPhMkJV1xlrwe0zkdVpOPO4FT
T/QybBwnyIcqsrf4g2q4CTHFPON9TmQUu3fXi99FopJvv/koXP33LLIXY29raYisRhEAdnMQv9ID
b4KbSH7XStXmjCNO/3ev3p5E56TAdNb/9dkXSIEQHRYGc/Zgb85YQs7EkeEV+Hg2h9SpHIkGYaAm
jHeBkzzDXlhPN0havJHfuNVtZdu3DPm8XiaYoIwUDRTKDMwwK+doXP8B7W3UanJaxOVfWA2zIM5o
P1wKxJyoAH7hGkSoH3XFi13f4GzUgqwdPTNMBKOA+Y+Viq9SmBU37/8qFuUumpVN+S54PA69gGZD
QlzEujmDqPX+Guy4sbCgRiw6szNBqu5s7N8JRgkjPaYJD8vHTIeGFbXY6q0LjtUZkuGwaJ9BohDo
AnnItsFYN84QiPvpNioC7D5DmH+d9RhbuNf96AbwNKyjD9WtlszS3NLpuSi8qZ4DXfR9i+ves+on
y4WWjnGGiCKxl+pwqGB6Au0ylFHea5chN4SugwywHLiMjQ3Cr4IrQ+pHzTF9iELLA6npbDhCP0wf
yOwmHFgc2XAq0UBNhvPK0cK4Pa6+IURggQdOwoQixlf7h/3IjLRiEyXRM+HPKDCRrJfXoE/EQHLt
/YqtDXeTVgnbRVewvW5EPQu2KRndxjPzazcS3meNG9dXcS/kUwslispvoIm+zdTR/LfJW5M130eX
nyqnqq/TWDFRrav9wDRtJoK6PzigToFmeD7f/Ruu/kfsS9/uaSu9Mb+3S1Gm3GvmnwQ7dQf73uNW
XWv/JgENapxmbdY4h3IJ7xl6DHfo9wEm1tmaD4VK021faOZuAtxQt21QB7fCEbA1Wm9bU+eQPtUE
8u/BVe0KClOCKb4tKd8W05vVOrX4kZAfJewpBVofBi1ky3kSv7U410ez07HjYCZ02Dy6F1WbtlR5
Smk4JdDu1mQ/hN/Bhm3e87pnPISNGz7z0G+VS65ZL6iUZtn5xvr2/nQvOd+cGZyZQzh3WkHROqw0
6X12w6UaHSZW6jpx6gLMTXb2l60wJFv//fIN5q6rblwlGXTQu6cS8rcZUCAiVCjtg0cZfG7oRh1M
Zlz1JJhCP+YscnCLQzmtD/DsKoVpEsn8ddAXnnYCm4f+dsITsye5FlFrbJ1aNmhX0nqXcFBBzwkG
iB6KWPCp6C1Qe9jJzoq/MAh7IKRfVqVTz8BZoQZR2fZpi574eW3aBjc28j9gF4sf0IqZGsILUcx9
fnOE7OfgOISNJ89kZFnCXPXkwgmcBwL7MYcjuRHWivasI5MvKv2xlj1mm29i/Ujo+HzJGwJ5DatU
6h55ek7U29+lTG8A67ZVoWQHRxX3ZF/mTi3vAwr6mlNlboyemkQpN483pjMoL5GGDmf3hNu+FLpI
qTvlgxreaAIEs1i8wGg/Ns3xy72O0a8spEWYizlAYi6KBdpWQvw0hMXrePT/EQGab5bctN4Ji6iK
UGhWX0VuWn/PxUYOuVv2g0XXCcXMrd6mBBGnoP3jbjGwI2h2UYxqWjLfzfepKy990qxu8JelKsx5
TPEM5KVwY+sSEQc2mPRmnwr61zu8EkQ8xe/zVBWwxtSHnplp1RHwF2D19bSc2K7a4TJSRmDVppS4
bqp/ELPJV2EjG+tZWUYK9jA9hrDg3GhfJDoHEm3Pgsi8k+ty0bcSWQUWgTKnv5FAw7e0+ZamSier
J1I1bLvtjPV7hf6OR/rzFO+OCTSeS57SqtHndLmbxK+QrshZ8DiBO+bWo4xqtpZKnRhVy56Yenrn
EGALB1oBuUf99j65ON5t3YL8JQBK4gnbICcYKEHQj6GP2NRJaq3SIzHQBEQ7/ubee5rUBlYxsZC7
5HQX0egjdW3H0cTskuMuBaezusTjWCc8Gz13+h97Gt6H13e+rofd/rm198Hsvu7dHQCvmpWezi3u
dQOlS5lfXIIp1aHnNsT+hkDIqXTWYuSWe+pRcZR5cnVMBMAGqttw0aHpuAsSbT3RFAlbs8ag9seG
qNjueC3pSUJWPj73ahhS0lT4ROpqSKNZyQiR3i5bI6JlA97LIzJfphd7XG77T9J6B8zfiHvPhiDn
FGTwDAo06iz5BRnybFskRQcJS7kShc59ojmI7V2nmBbloCpWspRKbFull8CvTal4C/leg49sk1hr
2gvvzTTFypKrgmLE75zBYxgWPgmM/DJfhMek+wSHSzL3+fsh2Vo84bi6B1REB3bH5N0ndPxCyk1T
6Fk1/Rq11l6bz6G+wT6CxnTKeFWiAfJgP8gM6/QLXbhiIgPy+bimFCGKGCkzENpCRh/oiCK1rF2r
1apK26ZmvhRlyfiuGrekS/e9axMbLdcWkO3D72wIshEnTSMPh+uT83wWCnVCf8+mG50NY9VYdQ0H
6d7ULu+40neJgw1NSbhEKF6Fw2EfmTvhYwsJiV5/47oJGNn2jxWb7Ia9mybzBPim5RlRDUSJB9u7
XO3HC6xo0djV55rILw291Xp+hbN7vk5/5RAwEhbjG+YWL1Wl8nrB49FpnrO5tqgaJ7lBq8pcUim2
sCO3x58XqbC478BZEExS9eyg55IKv3uscRMfvIhzx9FXe8muigHiEThg5AgykSSy5TIjFlpoEECx
DRx6GGwJULjKWEk69TCmfaPiEmfa6t7sWg1uvvk7kNNUvIfJopND9+UXMyg3XKihecw4GpxhkWNB
3p/EMXw1P+PE/HYHwRz7xBFNOiqlCEVs+sPc7cjb4jIY3kyG4oMqVN7u+UBwHTcq77uiaQObpmvH
eFk9nCH2ieEoTwIZcaByVgk3HUqc+xkIb9e+tUTj5MJ66QFX7HhVB+6rovZKBH04ZZ36cb7i4fUS
UocC/KsnMzrN4uyxGP3RDeXmqrTla/EP/gjO8W+vKp5DBxfX5w7x9gCHXjNFCEa1lzokO6ICj3SF
8ZZpFaGYZ3qHNT4y4rn6PG8QGq7g5gPDvSP65P/yloSok5PVZdsmoh7Gs+qiOoPV5oI2DN6By7B8
9jmOJ95XwzjnuukW9LzQZjyThMh9AKvUgeOSWopyUYg5ZSWyQlJUmkIi8gNYaIc1WxJvbqA5lL2D
KhHXjFt9XT9Y0tA/EWG8UJa7L6tG4ia+WF9tfuOrWqM/cVv2Vtosv486Rlwh7mHP7GpCAhix1Ish
UXdyqKneYfS0SdGV52yg3rm/XQKOJn7vow08pb45/hTT2gjxRdBUe8+JqeQupzaBhk9mWemrMoUy
J2wogBbvIfXbnJMYV2oCLrzbH5y4Q4e5kOGFzq13dDf6wVX6YowUC/17qpuBlnRANpSxSUPuxQ3o
VhQkMy9vsdWtIzOaZvaHvzctoB644tIsN9n0JlG45zqKWbld0KVADvO4D9sWcaaNT3XabdXZdJGs
x5G/AVljEo16LG6F9iB24VQqOYF6h6GDBUxO1chPnYEAvsQnbiEqTXgQubb7bfa2ROwRjigFWafD
JYAAjwdqvrUZvZZoto+QWyvNMOTguY61IxKF8tG0WEAjsxa50oApURudt5Of3Ue9nY2lBoL9jWlk
cJQfW+eJZBROFlk8mPrWTvUt7HjWy4bnWW4bZGOwwOBVVZJLb/I/ukqwXBo+rAobF6sNJmjVw5Gu
cUDGpp3vvjTS4buFdT48z0GgYmwf7BbElzMzU6bq0PIHM1eGX3VxPeOQHofAWUI7oq/oGf/bQVBA
1qeKhnEUb5KGWoG97G6mJftn9MqmwXrfWKfvoiJAY9bxmpslLlGE4V/e4VG8lONOxdP6b6dBP/Ru
cZ48j+BSl5CdGYtiPD/b/2VOk9gKYPCkC7pI2t0ue4/iHrsMMuCyeCoqpaA7y4VPeui0+oKg9U26
GM+33t4FTiV2gzg3y3V7H2HscbHjIEqDoGxPpbzowFBDe6fofea00gM6hqPGOru/j7G2Tyc4nr3l
blEzQ9TtCGsVkOUs8+K1zGJUNaU7VlQqCmvZtzw8kvCBcTF/TQrwy05W78NXTHjsgKLCgEk++9hY
Jon0b3ZbH/ywp3G8uQkafm0NVeGZHL56LBmuOKMrIKNpT34VL5KgLce8d6Vu7KOlYJVr0ahHjes8
knUUzi6Xcu+L/A97HTPjm1Eviyi2MEdvv+ybdlj59jzPqX2kYFSX9aDbHqhglyd2G2og32XHvmXT
uFFRrIYeQgs7472RXahjjqd2iEORfRAr4VIXpB+ZJULjGfOokWjpJkYjXZBA5n9oV6phToFd9UYB
kbdK+4WYTog79l73cK7bN2FlPlPQdI50XV1AQtp27OR/VP2LO1SE57kHCWkay5aa7v9Up56+FCAP
ZVFOI/Yhc+dpsoThGKPBgfpgqH6p8thsWKZKhNXLILE4nvmtSiHavjpoop3QuGWa8BgISiTuknW0
DxXcFK86YB3NWko4zORB/pTia6/AJO8W6ocLIsQr/a9UBgJe/g0rdhSuPiril//RKYBehNVsetWR
3T69z/XNRW/CRitPLjWA483STS9XYppt47Le83oIOhiSclw1HwmGBj/yAa9sP/ozuijoVdz3Dy81
g+gc79e0kY8dXTpTI4NhbTX89emgW7gmR6Tu+JdFcoIGypQkcMahLGc2iyRimuv81m1k46tVZ1ag
7AMOkyG7GfJaEtDvp4yR5JlG/jMVzahHiLKrlZSFOYs+w+1LP1vSRTXPCFbD5sS2GKfV4Fl06/t5
w+Qo7HG6XcllJIYx4Q9YtK91AUAA+ugiDZ3GCEEm4sPjCyc3EtXcXaaAg0rIs6/CBaBXGixvXPnc
C5n4AVGl+t/IF30L8byrQe7+/9tRKGuVmtQBjVe8JqICmFhgqeLiSZOe0pipTKxzdGvMfA0woMRb
5/S8fWlMIW1r2kx9KDzn+7VNa5rjfZ2QQkk4uBcJ6FJOqD/9nGXVUBdKcQy/0ylKQkQBZ1Oh2hUn
SCZ0vvvcR72M7YO5cFL8uPjsD7IoKp9PTu3l5trNr14IbeVNGNj8IaBe3Z/j4viq+zktE0RgABX+
w50Y4gaDitU7rnim3UX79j/QPUWDdWItMLi24OZviYwY26Y1tHsZpIrlincwbPOy561s9sVP9zhg
w+i/i8rsq+/hMffay5Ph1HEZLVGTkKSPU8msTvcMsQrRIF9w/DibmsDY5Z452/YDXvQuQwLKIbAD
ZdXUM/jVJAkL36GDT9GEr+0rZVuk0ReZdxLQHqMkbxqYk54QftHI/aB/uhLmEMsY/eTAv7F9W8Qm
8dfnfZzdItCsZy/rP20jQ6QKgkWHALSi2hkrF56YVmiNLsU3jGSK1KXnKT2Dz8+VqD1capoHV2Rd
M2rmPPQmpzovyk0tVzk+jUOY+d5ZxvgPgjLaiP8bC3vd1EYx5itCaMD+fmAetxeYde2RV/ih0pzS
sjvZ/iwV8yGuWay8RwOPvtyShXlYDbdBFv2vXQ2h8bza59KAcOxL8xymSGO24qu4uPOuKZ4hFzCr
v2qQLvw3txyAkUryIRQbcypn2Z47Fb1gLTUOAfrciboxwO8ojH5heLWj/XIP5GGXkHj6IXOLJDZl
PYLiP73aCJf8GqJ7i6ktnLhQBre+eWsITuyDv/ncAcDmrPg9XkU2KRgYuQZMDMwsJ4rV9aGVk629
HVmi1DGfIw8njryC8jgaZJAZLsX+IcC3gMGQndxOg7MpJVHb/yvAG86I5BP5cEmpE/k7EUerJZBP
FcB0fdECQ4Vn2RX//Zv9znUksQ3weYE1w3veHzJghVAta+P9b4zt2q+vYBZbIFfppF1F+/4qs/vy
w2RKE1qdzN4ZZbR6ZpYryY4F2qsj0DAWoERqcpSfWKNi57VBh0ragSQYq4Ex4a+gKuPF7/3eYzDL
jYv8dM/nXHPoOnL9IB5W9xnk4YkyLuZ7MFnDLCTlF/8slqw5hkpA3BH4sRgPHQWbUwORXwUXDuTX
ZYXX0xWGO57dOWZl/2PAn//4IQibwtbF0YZEj9thcITy+lQlL0LjIG/7tJiIR2g6Fy688KojyZJL
pnqZu7D5HIPM9pHk5MgSg3TTqRPm+Qlg86YN2PVcnm5tppKqgcYRBZrs2Gkqp4qm5NE9gutDo96+
6GKq8zDnGfhkRf4/FSnKqnRWPmhLHiQ2Dh9c+QLiGFVM9OgbO/uf95hcnv6lPqZxcGx0cxmfMaFg
F+a5Bh3VIGy03GkS02xKBWnU8L6nIz+YFLxuvFLyrk2dm3EVpxtphgH3gTMeXhBVrmxGstscj3ag
uA5nKhqzyDPhR5IwQR2u42rLaJSPSEL+gy/0UZjeRxAUTnum1xf8r+3EJnd9UtA8ztMwNlwFMQRp
kO69wWZXhdkQ8TOk6vEmmjSdG13Ml2YTMPdUF8TQgEYE/F7jL7bk4CKzIewGrHrh28vBMv/oy7kI
I/hYIegJ9gHdfCcIcuxEXBB5zlm99CSqumuBUdDQ9yytRABf5Y96tUHgrWfFirWHAEK1mM/A+h6p
0g0MDBPWEg7kcxlJ1nvLer8BT9b3txp218rXPucQsnVG5JXWWxqy9Yjv7HSkF7DAjj3f3SdPDYP8
5NXYBLFaWsIrGozk7V1xA4Pgjx7Z4jaGCw45ZxF12RnNO0YJXKGHdF0O/4nMn+kAMokwxbpcjEZT
JN2xFG3n2RzuX68sSHkpy1PN9FOWt4tdLrVLsovOv6OAqufE0YEg0YsbAvcEzsXOKxALmPFSBcqX
UgsNtWhcDntF0dyU6c91VdrvgrPlaMvXFqVgHgyLdhSKHpqIpA86lvh8PlsmLom6PhVgYsPFs13i
ODTwvdBR8N0wtPfJb44SLNzdw0Yslvsfq8Sd141xG5ROyEd+0pqKMKdUFRiNWmIPFgRxCFrPohGe
FSrOoxFArYm4nggm0rUMBLFxX2gaSsyTESuRu0x9jClnjgAibzhWE1UKrYsQ6G1DvON98tyXoOXO
+nIhcyIt88bE/KHseRLVAoHCORICEgl11j4PuUcV+7iyzOPhiym10cAPRjsmL/USjWDIiSNHFs6B
2QRNFgczOcQvm+ujZ+xVV65H/kJfzfVZ5HRph4djN715l9Lat24JLwKkDGVjVsMpNao/FdaIt7jB
aQtGzJpsm0FKVCBRWA5rr+0Urk7DXi2uxHwgJv63+FNZWJt5YKYqC9x7YQxuHU4VZeo8LbxRcQ6F
VlqFEty7ADIlrhMlpPe7KBEBiOrbU54501+vMJiAbkF9WUD/RT4s3VpONawu9LPerac6qiHIdq5U
j0b1+lzn2uoBhzTcoT+6IXNkrxr4oBB3Ko+Z2E3Gz7QYU5h/ad23xA0qbwQ+g+abP4UF2rSTWK3T
5kOQG3/mPf76+ai2S2CCoPyTE+dxHGLDEQJ+FxP169iAIKE3R9Zmjln2Qo/obEetEKuIXM12LHJN
3HULIiY8UCS9BAAz3FoAX4bI55V2c7TxZQ9KW7J5Tondb9XPM7m6hytRG03trjuAcBMYGcMeSuM0
WQICdoX0FEOcc8dUp5eVi3NXQeVg9QADhHRyHTNyAdwISeC57dNDfUcyzRP9G8j41WTcGiD8z7xQ
oU9xIJs1aHBUtXIR18DrQTkXKFlFwB4yrVGnXzL2CM3emngA4o/HrEBNTVK1iikzLRIhmromFURz
LP5pqCdRte7vY5CRFbnrTKGpSeA/zo0awG7SsTV/yHBlVc1qg4fJDxsxZE67Qxf2faAI9FkmoMPO
oWGHqQMRnRzoUByTmEybc16Tco04/971xCwsAxq+74MLse41gNYo2IrISEkzDJQ7qDd9KTeBkBP8
+C2DxrP6dShL8xFsLDxeZALsByq2bkyoTXiKa+586uSdRUg1FHQ10yIgqyl90mPNcsm/IheLbnEA
342U4Uh00wJDJA3K7Pc0kenZI9Rcm21j+qBEk1TR6XCkK4DbXmz0XL4GsK2WNM1xoHRsCRxV4ksA
z9T/pR7yAKK4qTWlURoFdsXt+x+RyGlGPqdlxmkYtCA4LXQvGJTNrKxnpSQnipp/Eo77ybFAZGLM
5OvVDV+ImFPSmwmR4LbZ3NS7otnZ98sQvBw5MmHcCMObK0qCnxFdj4CjMrqsCZ0mDyiIyqH189wx
sODyIagjAKaHI7ZYRc1ZP6+eN/8DdGV2gXk8OoxmIDuiuOZrC80nMTp7nXAq68qmRey8FMkGcxxs
XBLGTUV2XIgdBDpv+ttx9UWN7y7uR9p9VG3QnP1WTAVg9TFljt6kHU8Mc9Hcgn09SYMwS4FRJK8F
YUSpxtFgIluQUxWbbHjJFOckcMb6i9YIFA9EyM8lSIF2YA7eNXU26qzJaSjzI1nlq8y2s3KQL0yj
ZnnJEwInpzT1N/zu94zmDoBJ8BLySSQ973T+RfRfX3agdieOmEDkA9BhA7/nNTdE0cFqyj3BZJW9
gZdDt3YPjujJo8OMKcIdk7a+d4Kbw6AMnOUmJ1k4VbdTzO93QLEZ3iLvFZ5LptNnZI5KflG9Igwv
TYmx8VMb5Jas13IwFka01NdKuS47MI98C9MREZjReYNmu8r6++pqhIvGfl3iOZQ4bfqcl+401rID
F9pREcIsJTUoN+Ay6C7zPafZiEPcYx3YQH+eJ4NCjj8Lh2ad9Z333hnnMku5JJQKq4YeDORjoq6c
izHCdH4y0VjrxLt37/CIXBSYpjRhWH9MSsobAaoTCv+h51jBkxms6wt7evz0jAsTVPfRHEcReR1l
ajVYcS4mSpyeIw/J0P/2I50VrLHKvJbnTbmsDk6aRv0DRZCw8R3DvLil0EfhYMNu3RbUBBsEwCHh
pKoA2ou3+M9r88OOXXC9YZXw1VC4SL8KQVT3d6W8EASYxjy++ld485nPWgZq2kMjb2h8atbMON/p
Mx7aJE/kyOpRDxH2em3RQaHdxYz4TQS0nZaFHMLKkwNgWfe7ExrL8YJGqR82XgI/BPU7jQ+hJ07y
iUbjJKCkJCY7keQPCaoYvbj93bqMG4Jdd284nYrevbDifkz+XCdccESAWDegT44CvwmNeymoueSk
InES7hoxlAKU6THkINunVCDVEmgzqc/ZiVpT0UIu6rIQK+U7+a5CYP1sJ2U/ijVs0rXXf4NO6o66
a/aiB8g+c1VQb5gwxFGMDJ9esv4tXsHQtgHMH2LHMjiFEFtShtsDGnvJVUVlzrDIAid2TRSio0Cr
l9cbZivHat8++DhLmRn31gsao6vfVkz1NZh68U9WYrOwtxwGiOwMBM4JeFR4k+kegnjR/z5WhMBF
ouhRtwJMFYHtlG7MJffPab3jCqdo9AHKWxn+gJ1iiZL7IQ+TKHMXv43qA/XyksVUbTeFNx5RgjFl
UKc2UMbyoHIe84Ti3QKSzAVUzLnEZmup/i0yvv4vEhYjo1kXyVDOigyD8FW3semzURUEmZLUYVow
ENIOOonvf4XxQIQE7DI3d2oKh2X+KuYC3fD1HFmHuRUK9txwyB3sI4SRnfFXb8rNj/S0OsQbg+qE
RpL549rdGfAQDzdNgKdtdCuO9GbtAja+orJbFnVJxSuItxiQyStRDNbDmWxDhFeF1PeJbHyQpDwh
aKbSE1Nbq/gfyxrCI9HQTRf11QY0LZ9FYfzT197/9Z/lfdJ3Mr+nl1HsiJsXSchww+JjxBrQr9lc
LZ5pTfO2rvywxYEW3NnyUBCQCRcpw9MM19f0jLUXT87aWGKxrGBm9Ss+26SG1jmVP14cr+I9TJJR
ZnHOLy4YH4o8gCSSuPQoJ1kelcxW9rGZwy8blj6ff7eEb6T2jAJnGLVkG0W0AdgxRVXbdQ4pK8ux
+DCXCrHHVF6qK/I/O0XTYiXx/CXEp958Jy6bswHO6078K6ekH0QvcoAhsWPPZ2X09+wWHMsiXo2V
1pNKfn3/n+oBca9/WF9ofbieq3i+yiVWvRB4ZiSuGhovdHpvBAQ8rlJWXTXYoAgaGrTtZ45TTcPT
FPotBpv3zqvLg6XNmZt/IYE/fnhQWvr7dOZiHKkLAIrRTwd6ikgINvVr0+/zSPLbK+YwVe1DDWRJ
2N7nK6RxaVZ1Phcfp/4AgNWUu8uRkCy1eDPLWDgZKzQKHPr3lzsP3fuHDk+aX0q006oJ89SDXERQ
Jl3rrp1w49geRaDZRnulldDLx108EafqcxU5Q6AXUbO0kGgKATgy0qwTFpKo+yv3Ar/6VSqr9UrE
3sxcPPF+unGPzVPA/Qg+AIc8Lr1pxtHcDWd/+CI7eFCpDTScFyxq75FnpHxgct022tiHmWdQHuCz
g3gQxhgpoZ2ZwlWOJhWuoqhDUsZxhHDK3z5ehF4zivGAhmcZBIclc1kHeQNMHNW5Ywnqw+vg0rKd
z95bfWrL5ifVylQ4PNtTsPEXo4jkllsaFkVLP/+QWff4xnZNw8WJJoNnJssO7EazSyvP/5EYx6Ih
jRbxF2E6wBsh7AaZGl9DsMTghkdfbTBrhVZIyEc1VfHuJwQD5f24A+wmpFGQWXpNe6arbjxUS7e1
iIwu+DcBl+Xgyx/amoB8PKgK89GE2E3aNKbD/DOby6aHF4GEkreL/F56fWwMQKJpR5ZSMuR7GTpY
4pjXwaJmtvrPgHoyYlijTRgFG34xkFBc78moHqH1rmi8xl+r4Unatc0BTYx4OES3AWyxp/O3qHnp
LkPObYrSPN+sb7dGzhqn1/1E7SmiymYCKyNMcrjg1O+Y8zHjkYmGHWk1q0MFd1AjY3seH944aoAs
ExET2U+Hw4BqRfVeDwsDfQHP995i69Dz7PELj3vepVWIhBNn4n7z34iR9L8vAUL9Tsi9WHuFJkIs
V0bF1k3qoqh76jkVSs3Nbx+Ba5M2aFGHxf+ARW44diqajbThz/IrG6YbDL/Wyfb0ci287AqeXRsA
hNffmosAuRx0SX2zFz+YZmd3SLCrzPAzAiAkZu0dpga4NxwggI1DpOXIEvCCDiH4OjVJx73QizXp
PnpLWdXZMio0Awaew1yqnmDgU5M7MDWAJLk9LyAq2xpo61vCxmEaEFol0EEKH7yDdlkGGyZZHuPj
QrRqUSrendWcGgY/b27blyqd9SDloXBaly2h5Ow5dQgwP75x9o/SHSP7TmUWEHEokK5xdFBSPTOO
aTic2gr+BJEIX4DjFPZAuhjNFzf1ymDgb7Wy78BmX44ymj8BsX2F6HHJLiBYcNvL/6tjDN3Zs9l1
7xrJIHYno+Te5/+4rur6F7L/FqNJ5dMHVe5FxFn/f1aBRcmCb0vrGRH/SaTQH3MhKzG2QXYQ+LGz
pwuVnLgvyyCRUo1d7gK+3tCyMJNhXEl3QLz+4WPbOfNIlJpVXw3C+N1YXD9bodwsCfQOP/fi+NYE
/OrTcwMd4q05lKIsbxBNmy7oVZVajwYlkHJXZf2xLyWawM357O1MYvPnlDhk0DK8D/qnr6JezL72
YGeuHg5JCt+Ez0oTYbphrPqF6Q0nabGEAvmapFD6cbBwpOnPAVjW9r3wPo0Q/NY/ePSogZfVxObW
VDXpwrgm0cYK99nZ/DSNxJSIzMKJPYFavpeBMuItmyGLRnE43OGTbwYd/wnlEHmEc79dfc0MqeeI
dklNZHES02eIjpw6BcgQ8/uT+av8NgH0ZC6MUBLMQwqaJGFdgAGGPNk8GUs/TK/X88t9xbVyc7Ng
6ViJz+WOpqicj7NqzYRbhTBG9LPbRnYNQlq14KjcRkNYdu04vn283mKJyyp+qnCftdcdWj9YqSmz
YbUJyAlhjrXCHbKQ9OAhEhkH6W9GFk7DdS3BZXoAnIT15wG9K8T9+CUZ1WPgNKm7WLEwurt4NK3F
udLEozeX6Cy2tIBY5+lJ2ncu9WyoK1N2jF7KLPJRpEtT0naB5fqHsYPhOCZK/KI/4gL3eiwJawOR
d1+0U8khvFaIoCZV8A/CsEhF/MIIZzymaP9NePnMr7BWJi7P+ehEzove6W5383ceLKU1YVflfg0V
VXiWVADVvUVInkkr8Pe886jeORd2SqBR+PrvPl6Dz3CV03oD3D+4CC6HT81yWEblk3RceL8TrTk5
tZPa6T17YVDnTsW+CBN9sRw7x0sBfWv481QKO6D8Wc68C2NbOe4yMbR1tQR4NtviovN9zJs4afTn
tOxk7qNvygufei1UG8iBa2DTdiGRAqF5LhXM/WWU/XBWRJuQFqxbkK/ZXGEt42gvcR4EaH5wyj1R
qk+3Z2xxTMOBgwXi+2qQgzo93shstEBr6TSUY9chTh1tovnRvDFp6GgxfCxpDj8q44eKe28pf0M6
NoaTNjtjMTjG3lDoiqx1pFuvUZ8lDJhZGsDxu/j5h7wWyX02mobsSPpPrfBTNLIJ+60TxI+kfa9O
qxEyLU8rVg5gzADxq8Zr2JG4knqGM8H1kjpxdBkgi9r0BEWnauMEPkhE25zZwCAnZgSdCikheCNc
nnQJCjsxZS7So0qt8lcFJK1tD6CcyJcFoj56lLNMiGCN16gPixfHBWAFFE69nkTxHOGGQetscgUg
jaFI2/+y0BwN/a0ukH5PKwZ+nEM7YzZdfcuWBwDcdcaBbs5vE7qduaxnBAk5niwd9vgLWO/WxPyP
bS1J/D2c7/vEyCJHbqUmo8BWXl59dNH4BUVBNoToQKtm5IHfF9Qte0ybWwnllqZTYXowCYbOXDS+
jkXaBpW3tqZ18SPwGaSAoobd7zZEHi7w0yFYU+Qh/LxxtdVaEIPi+5sLw1vAaRswBs3Ec2ta5RBS
rQRuUsFFM2CpRw0vL9k5JLGPSRwujbTV4rhlSTBDcR5ygJH0it2pE9nzl85GdVUEG8KB+O846GwW
UgUkhu/WdzFF3TgX6uEjmqPEA7WsYcmDE3OigHm+EpLIOhCt7qvImmINLklzxnFavxAaAKr89foa
lrmIxg3nRQGdiCn8NojhUzB0DqHFa5mU/YfJpzUSWDdvqcs0JpGtCmF9BVTFmkBBnwuW/WQckck1
FsEEyaoXMRVREiNCn0w9V5adpC14cceRqPseZB42FsbmOAdzLaIw1LoylQxpoB7G7xrztu8Fo/58
fzyiy3IEZ3jpVzH0gm1pGpbcsTWTFdnm5M0yiAbOb9VVE7MiGuz/YhrFtpoG3m5e2uK3kfSfEDAK
1ziknOUHSFipb6kT9z/MEHcYVT1jlKVGpQ1mrIXCHc/0jUzESJ/u4+eLOgF9BkHKL0S09mWrlpqj
xbwpDSepxR7i4w1zOlBJgNrFWOBeAdXEUekmzPX57Rso0oF3JsZOjnEEeVKTS7DzuXYJfzIY6EP7
UjhuYwofo/xrUTWXPHfaAo62qzWZmqD9vqxz2yiRO9466gMpqi3xl1RGEDp2tUjVF9tA1bCa+FGW
zRmB4ynvYdCHqztdZRthKKLxmXlVqfC2pONPrRGAE9q++XTTmJ/eLpCEGp97UgU2YTYoe8FL8BBy
ZaT0b4/7lmhEsBQ5Ys44vMXiz8OuIja25Qh9b+9XCqbuS4PXPDBiRgZFFfifWODFZFGq3SJ4cUJf
tIJtWhFBshpMw+UhM1DfMP3e6XmpHz9IB+74nDFo+tGLTiWQhRNvbFKMMLhSqsmjxL4gRriDBfRg
sGOrmDyBUdfF0QDuSQHpMTDdXQ8izgqYNOLPklG4CVpXU1qK6Eo7c4ynPyyUiV8z4j075+d45kZK
5fJN2EGstBFo5jBrI4YJnorgNVhbu0XCD6JZQ6onWi1Fo/cFfXst7ag/GYMZWRQ2LrkxnLyb676h
Zhlt1+nPTTTO7285/lWI8YCeWYePJ710UXTBrDLph72gUxwgeTn4g9oP2PCLnmXOpS8t6/jbRsT5
iPy4hozwUxfYz6LIQLAoMsUDwrbn0hX7ZabtXZeZERAmum5n4Sjmcm8Z6LW2eUU/YswMbznN/Peq
KzAjnZ67vZB+MRP6uHkt17B2kXwejJkJsRip43BqRNwnDxbBV5g6gMXeZjrwNZpIng/o0rVZgBpj
BfGTGgZ0TS6r76BvJFXxJavde/cJEkwGEuA8dRLcitCGTqI0fc8q2sUcDYvf8/Oiabv/QSxdVXTy
WsVaKu0hmMZFzcxLSDb4WPBovuZIgsDMVvIwz/y6sSkAxE+mmyitKBhlHC4dKOaMAqmMvK+O1u34
P+Bq3wzxwLhPnxQ6q9yAs+xRq/mtNVnFvcCfShdfCpyvZoeyuXhLwMUQ8nqlmao4SpWhFDsvtsHx
ETkp16VkJ0M5m39btwvHUd/ErOT+4w3g5IgJ3dhgXA4mTvY+srJ0vvfFwxEwaLgXyNOP9VM9VMcm
bhZuGy5n9Z+NtasC2AGNR/1RPFAJ0jkt0koUhFzWNi+zDE6lEMXjV5uOfFteksZIHnE78f/PMSM9
3tcDgJawkw9nXIeJHAaxSDLnvyLq7knB/c+6f3//SAswkPl+i7+6uZWeJtSlLT3SNDzdcP55LzCS
JA4MMff/vJjElHPtqTQkTwZpEDKtZWPZLsPbdNBFBmE8Vxp5PaEer9WVjxI+S2zsdVRuna46cMT9
Ia085viRK9f0jCSXhIaNRxtD7K9dp7zML3ESAqwC4gU76Wj3t0/cQGAauyB2IKjzTjihePtZm31c
pU/hlRmTTwqHmOLkjJ8YpOVg7Mk88qdJV+HqJQ9xeIBzjEhYGnn6x1yXbOdkoqtYKr6WgxRIDbdk
Fe2aR08iVfAjpHGgiTFI3S+RX1LCnE/nLXzhMxfE34aYJefbN+LCPiHM+qLTY1Qqw2yyd+ih/ITD
5k4QJ5T48m1IPiTAIt7ZAykP+E42v0TCasO931DEOyNPrfIJnCgSsEAlBzLBZYQC/UtA1//gs3Jn
tHkfDH8BSOxzd2MYayPMkIinFQufqU7q6yTGyadVb9ZzxGH7R3SQBZJUZ8NVwQ1t2ye5X19Hc+H5
T21k8/DlDNX86z/f83lc5jZlIJmtG3tHBAA5B6yFbQr/fgbzrbsxQw0YHxN3wK02gQ0HF2eCwpjN
Ie3tjgxp4LwFc6Lt1PQrYhBTpN51axNNNEQthxC1fw3fVBsp3S9722wmUWOCy7Ca7pam0d6ITlmX
kqpOCAtVUa9+8bDlKRCcd7+XkWxneW5PU/wZ12I0NMgCkOr4MOdELpl2oFm4Czi3onF9uPImIwVk
ed6dLkRwVYJJS+VRWUXaChQg19Uk6UTxmxmNqavsdaJBztoLiDVXRMgGsrnsc1s3FmRM9C7c/1nN
npoN1R3JxMtFx6Sp0koB3X96rd52me82BMkiElDM+s5+yQ9phHm4MYBeKMeA5etltJYzGXC4YvB7
yXzWzgryQDSYfsRMUFy+m1xsNh4K7MZbBSnWao4rgqvhXm2WHuwTvZM/z+6kVGlNvsWMJmwdKloB
kjsGb9E9r/DGkSVJei6jP3/3flMZVUqhRiL/+tYTcrFVqoI+RPkqpsRdzZOgHVjI3OWHtr/az7jJ
iCcdZ8cc3Fr7VyTT1k8lyxreUcCn+RQ8R+gC2+qzYnZugj+Pkj8hYCsIejXqH8CXrBghXMLIANnl
r2Yep0FoCbZsO3o+brbFtMiKfkeqNjISdIKeLW0f2Isierqmc6cbYdGQh2p9X7CaLn4PnQSZkbsV
CjNhaiKveS2bgZnD3CgckqhC8WzYXKinpBp9+T2WO9JI092esnN32Cy9rvAr6+BVF5zdqDS0QiXM
oJ7Q4A6oTE3/gmhRLthOuw2rFvrNQrJI0+ul79vDeWXcVy8ROmw1UUvL9oPHqEdcuEFYlewcxRsT
/usbFsOHOEp2tOPEaoENGGW0C8MEPXs7c4EwJIpE4Rb0aOG2TaZept3WTHkrbenM202TD4fziSxx
XjMLbR3Q4vbrowTWGWxAMzMor4FJb1jHbeOsgp12oaA6H50UyB42g0B7xqMMVp8CwrQfh9ImFSy+
eVTG9PzcOz9mGNLd/cuFj4i/n25SqALQxYZPcyKaF1bYixOryeSw9P8RchebQxwT425zfkSxY4mL
C33p7dtCO+6hUFTgbmMXtGrD6CoXQ+tjl2ALF51grLNbZLd4GEiarGapTsRu/MWR2imfJvjR51SK
AmhfhDJze/v8N//jyTjUg2LnIuknqQEEa2xoR1YtFPsTgkHp54PYBRV4TU7mYCYkm1o1XhNAfZab
zEuFJ27xPn+pYBv9kCDfIItlbmPyRZ/CupFQobgyLKCuAQoQnh9JBrhwwmYD+Zxq0PpBxQCO/cxX
IjeKF7WfH8BNZcRTaMPM/ekvUKuiDLqQPxCq9lrf8GYyBKY7jkc033aTD0Qyvh+5/qfavH8GT/qT
3aA9fQNaRejSojCQsAA5IrrkOCgJkMnFObky0SbgC57l3uvqhp8jm9iFu/UZFR3VcoFNDqG0eVJk
9Fv3+ZxZLS0m7fhOAVud8+/T3i0NYDNsapBwz2YaM8zanzS0wcE7UcozkmR34iuKRmArjKQep24I
fP1kdd+1wVDson6TivTk8n/sXivXcPnPb/J+qwUv9arMvgbP99PgmimAxsgjEIJZrHgGNmEl8l99
oZaWNKC5R7PooZCLKFp/IyHAk4ROUv8tzYLl8Iayg5Z5i2WHqQ2POLyo0giygb5hDiNO8xhw/fGU
vIe26H77g7YThpDBSH5IWIgcBNQ9OdQUBaQSgTpXCcNlNXvKIyepDctW6e77RVFpe3ZKwrlPWtm7
NKbiks7MJUPsSlkHNEyG4aHo/Zuy4E/l/y854OBSSLwdxM3D7rKZCISFFNSQqS+ccKWsHHOdSTen
DQp3naEgFAlpIhmaG7qJ+MqpzZeui4r2N2MbuXRQrdYf0q6WPCcaSyJlh/aJQNMdcRy6YmoIKVt6
8kZsHrLS2lFG0Ihan6DKo0XRTTOJ1+5/YLEzfA4ukpKF4VrCCU6hBH+cZF0RCjO32+h6NBVq7TBt
GAVzujtQNkqunwWB48LoPo4L3nwPpFZwb5r49LMEKoPmqgVZLZNBL0+mNvu2QGMnH3RDiRI2LhEN
slY6yl70veN2mNBhz6IiiQu6qXtHrmplD7OHbN8ACeb9l0tnfdiq+XvlfjH00KmKC0VVwE3G4RFb
SefgoBMo9gVUVqQTCTkypXLaJTOWwbWGCI6GPUJgJe/SrDIA4KEaQp71/3mkp3VtmLOKJJPcxIgJ
hx0AvJQJ8Vuiz2BY+g8L7vUnQ8yY7sGrbDPF4M3s7Rh5PgpkemDMdYNQwa8deC6x8zbQAAUbKjqB
WjcWeWabJj6hsx7s33kBqzSgCE95KMkQKKnMXPdsvEPVACpO0jdxJdm/mf5axMzJHBdgorZIt/kS
PTV8hZBKrpPfRBVLK1qsTgHKsoskOGqe018kNPnpOpWnWzmsaUe9q/3AhB63qtJXTvNtDs9GZQrJ
R/Y5Err6O4xHGNkTd+nLjHhO0snfTLu1VXiL+2Ef4b4IDa2uojMjpGmVxH1evUMZloPVJVcSaKbW
LzvjraPHCBUagMY56k4XKXX+7FDa7sg8hB/TYDb1DqHrHbf/qbdwtjfCcXn8zAJxEjK5Ak+TR3LO
aq/TkoeDLG/6oP3UUoB/t59ksiqXNbrTjajUt4eGY95QfrHN3NtWivFoo+9j9weX0Q2rtI7MvsOL
ttUCMIBwkXai6BGfoWmwoYiT+KqrOXhDKrEOY/k8o+RCWqNAOodWZqg8aO3gfsGRH063f/vNpTjE
XQCvizZQZpn0RAz+ryACerGEfvE4Oyyn6+toiF195qxkLnxbhIu/QwQzBv0PKEjyN6p4019xKqwB
9CFEbcPNywPoXT1XmsBHGK3apuZNJ8Q55gBPnf9HVqVIh2Js/cMEs70Xl8a8t7O9Hso0XOqpdcZI
lVFIfkwMl5TC4mD+wUCYBBzUFUNavwC1YJFcOVo/Mzi55YZw0cxVY3OqvAZnO57i3lfsUuSr9ftv
z19M3+P7NgWnqcMH2OO/sYHkdPcz1VK+dxp8iHhG+cTpxgnAovailnSm7LTBXNaK+q7EHsQvR4Ji
ylFZrUBdXMWUxOLj60K0dRX64btwQHNCYlsfEOc4f+99nYI1mq6ZExV+LrsS0F5yK4j65y/99I3J
6T6fMd+BmYVmQycO3ENfKYj6LDdKyIxmq2yURB1atcxCq1VXOiifmWwZaeB5eVNOAQVQYdkyGH47
o+Ku85CWOCckmrPAG7SPbWhm/0L5qWDMKFxwRVOlygYYzigK9hH1HLRBBt8ZbAb1o2oRp60cxFg8
Rv4U1x624GqpUC1lVH4J0WFajtwB/QIHM9cLf8UwFuyfOz4sQ81L/CtdDtmDPDoxSNQ19z+3LRUB
M+eZaX8EGlLx6pAxiYkpCxSQtRszZgKCocjcj+AlfnpGbKFC7vQf3sBFFQbqTW/tArk3xJ13myej
Ulw2n+AGuZolnExJYOj6FoA8+2Z57uN1Q+v0HpM4CLe/HVcWrZ6+OQwosoJV3igs/Lq1TJ0bxKtb
iaFc8XDjc3xPPDE1nCxELjSHjEKriKc/Dvsf+XLTuuFvWwtp2yMJXuPtL38JbvVLmzhntE+3Z1W8
JNbnsGEDIN87n8POKokLkAIHfRpbMYcjYJojXxmWs4pCrnKRNLb+Qxpg3lp9Qm4Cf0Q5p22Q2crr
1KAYyA9gMQy7MhsO6XNI0119z2yq7mHQMu7txiLNRZDeV/QiezgC+8ZOHR17WW2OAdD3yE7eOZrt
sXCiX/BZoa9d6CT58xmz0YvE2tyiEZU0wT7iDHSkeLd3ZS6nyQU4Z6Yu3rxorZka5Ae2tzBgx4oD
wsGOQOKdXtwqiv2YE2AXQAiKZx9vsoffkCnWu87GCZssf2W2Lnke84clMZet4SnzhPfMhFmMkVg+
V43eym6pOFENGZ1qaquCkqSdOftAtooIT9bNhzDtvUCcMv7+prgCbrGBs5c8FVCAbnGVO9CwMGaq
GkKXc/ggrlxkfyj8cr/w/VcNnZSmDwhiDLTLqEl+eJ4BQT4RTDkvFVVoIvt1TyKo53XHEvXF9CEt
EqktNAyS3vlyEcReKAm8GBGJc1dEsZCJE50cLVh1tF/yrtHwJjcmtaposOKp6qR4HiUDpvqBrIAS
KyaTzVkU6b3vwDLI18SxVG35SopOjfFqQ2NKijNwlGCAJYpGk1m+rfSkL53DclU5/wqTaTIed/X5
aUyf8j0AlWFQ4wZyzdgklg4NRVUvtC+XRVjVrm5h2sGu69Eux8B17KCMPaJmurEivkxbygwUclqY
1pygRQVtwmz8qOm4OUz+QhGc9NBkde686CPKdzG7h8UfnzUg59qlVBS1DtFwoZu0W7kalnCUiSGb
PC/5rFcSRiRtcbPz0kWFOH33qZj+EI31ro2K9kzwsWTVNzy6DhePeYZYRqGqWVIXMfxGZtb4aAs5
n7VzEyPxAPLL11M9DhIB7+yb/h3i+1OSHmSTKZA04i+h+segoAVSRqzB93GE0aoSp5nCGwhEqFFi
jEZLELJwdLVxL/D9NpubXoQFzq33IFnZUEXfz2OGK66WF4mGhyXcBbe6FtfK+YXDGkxl265vcSfC
XkHXz8uf4JG1SYc1WzE6uzILdzNrqjevqjtXWDZIa0kukGK+CQaGBkRSFVPPKVY6MPje7dyPPAjC
O3Hpve72uH/orkMnmUKzSfx/yuJnecA0sxSSa7VTioonU19vXDGFff/hQrX2wQ6ITDxhptPD1lQz
GIyLxEZ39YNmJu68Co5r+g7WHpCh8yam7m8gyw0ElHpnOTU9EQ4zIMvZCkJjNtDrf7CxomLWnVO/
/BoANuCmsJrPR2l0Bgx/avWaVYsPDrDbgrtVdAxJzjfvNICyEXLBxbiJyRBbBlTTwhyMVNkXSyC8
LfdsdP2sMEr4ff9sGxcEfAD4PFctNHR0Tt1zxTefTk81INr8aw9oj5MV3QfjE6KRJeFf9TjyD42Z
WVPaZpkFccgGrO+NNqrER3Alf5dG5OTM/zfWlQblSjKJsFrc8bNL6nzL8XjZx03radCEMI/Px7PB
ijUW4BZYV9PnBpKc/kTQMAjJIxJU/NDS23Iz9yKQ5K5ZkiKK0n2QdF60VxffKREJa/+B1LRf6kYR
bA9G3vhZfwotBC6FnKFjCxmDzIC+Q10vhbACQowPLLDqQg6v5Co/goiYe/4gzPOa8qicpbHL+5n6
wCHVIT+I1BJLa4tKc6feTvLKeMYEqaPl7XeRtyyq2iOtMLZavKdYbnYfQPsladzBjJuCxaUXeO7h
+pcDgsOodYrwIDfJGLbQ1B1vKo3yVivMJ+BS85pgHLpjZc4LeGzp5C3NNIZEjPnfmuM2XFRg4g4A
Bc5V2izaByACvBvW7S0g0nelcw8BGyzr0XO4+kfzd6ZetV2U67VFMKeyxtvL1J8l30AIcQO2/W2u
OB2TQMflbE0u4k7a0LK34h027FQlgk64LJrqDpgNn1z4pQWpo7FrcAJ7685g915wnzpJkZ0O3mXE
OwpVLOGsKBtxCM0publhmOrTwfZzitFvi03EPaLgUqwjr+W0R6Xuf95/cbZZUNXVjTCZ9oE92W04
C/HcUZvKlMr6K6eAEew5Ig6qWeHRafrGvSl+76sNmQ0aHaNKUbL7qmIN04Izi2o7yAfQNXFiLnuR
j/ASSXcDTZoGSO6k3tGP2Hs0jWFzjFJUZR1kG2kLAESAsMkiM6Muv+wLej87/iNafdOa0POglbvM
OzzYrd5046vz29E18KK90HxLedlc14UmrwmNUvCWhzWZucW1z2TUQzW7fcrfzKempAjRTx7uasFQ
fjivclk2MOkmRk7H8NSwQcymTj3nXQ4qpaDJeXrhlwDm1DpMMCypOjggEvX3DYFuIQNoHhxcXw/T
XZY9bePVPiDPmhXwiTcrCYBSyUyPZhGhjx5TulIZy0nJh3CYhqV1ibqW3/2Dd2bQnK/vIW4zwJkk
O6n7+eMnXcqwlwuTc5jLQKkjU77MS/I2V6yJFy92tcXG7/eACySpkri8V51TzfV2WZ7OSgc7CzfV
vXq5uatXh2uI0GIcfZxp2QrMaVEJA8pDM3869JNK+uWqHf1+ujdi8ehfMdtVSYjVXx7JqyPOhSdR
9h70MsiMDWvuUIxw61vziQCq3FF4OOf4jzHGMa+W0cN5vGzX7N61BYg4cSYNcdiAgPN8/leDYTFr
UfcMPORwHRhVxz+fHVrYOTwqLOi82NkV+w7blncp6uKNdCTCb8DOL3ghvX10vPn8uOBOqJTwa3h5
7rAo+5KGX2Wmx2ApUuzbthdT1zHUUAftRjXpiglw5S5NBntNQ47K0ZPbVS7uocsmwl8eP9MndQ3F
BIRRs+4awqK/MgjTL3snGsfZAZH3V5LUw1Jz7x1FCCeRi3h86XxvqQCsIRSfaBm9gfNTDFLnqNUF
ah0TqhP0a9cSDqnLkLqdi3IYl+bXcI506imXiuwQ6dryeSo1kT464Wgp5xLaCDkjKLbrd4XRhQNU
0WFjLHY9D0s5NajRMcqNnY9B2/PZ5fFfc57L8L1VgZBYqRzfnHaQTHrZkNmF/KlHDRGeAhfys9Jp
LHJGgWglRpUfcmZ5r1OyYHvvXF6/9qOf7iHhCqFnMpDTnNWG0SUeXW3rT0E88VcrXkaONaIX5og4
kmg8E2fbfblSniA8PC2U980GTGnHA7dqqS+Evw0u8B5yjqzEqkFdi+8YlLQNRADl223+qsGPg2zt
f9eTlVOlvxL6YnatWP/cPwA4sjeyb1/wqCqEavGYbZgJVywHpjof089OTNNGJcVC1mIl3gj6nNcs
WGJQBkekZnrF2t2nNKVVb8fErJN1O5AqNGaP2yT3Iqd46y7FviDs0jxmU1KwUXTnImPAWX16f1qP
+pS0VDAUtONaYOFUvNBCQw6N39ia4afMIUZ80liMG9LmPhUcR48ylXtEUFiHPLwv4e60CtS1qZsi
rUb8RemGxWcp6Pc57jdWKM2onQWX4ZFU8DK5O93mrv4V4UsiTlvG9ehull9rZHwu3Lksl4z8GxWS
TzNDRfKGL0wnvNKASsjHqa2c4Qae/tnil/9HU6Aas+mGniCqmnvwrSJ3RD81vbWawG9lkV4mNXh8
+/DniOlJqngIXgbrZU7y3p5/4AUmNiLLLYoDI0oUyL37ZS9BNKsot24vZ6nso1n79t6+Jgl13v92
5MdLTNMb0w8L5hNABQbKVbzZm1mwccC2bOqEmEoFVeJzapy4lx4cPGQDJemWnGNumNUcwPGfZKyb
X5U1fztk/2IKU/URq9RCYVLKX6As1oEpCaOcNK4Ojr/+kDXB69zrviK0iLvSE9mjcAUclE+/X0DO
vZ7dY4DnqegmMIYrTabM6E163lsoKxE4LeSDQaUKD3oHY1g2L83UYoxpwuY+yMJV6DQ4aO3LZwBV
xCL9vzZYl77sEkowTurnqeUVrgeGSRDIHzzsAsKnvgFMCPNAtR1WFwqS0ZOyw39QRnNdf7BwDrv9
0+r3Xi9Rjqou1UREgnsWC3bTQ2mad0sqwfCrJFYTOHZUb3YAaVMV+96MlEbmjQBgX9gQD2VY6Wdr
A4ceG/hXtswLH82w4D3EY24Be5wKnyte2K9tA9gXmYLaMt+QW8tDVWK7t3I9q2+gB631Fp1b9HSw
0IkNpWVO10asuvrc3zGP/xKg/iM+hZMc/PoTTVmNlXP/kNw/BMr1wbTbTDIzE+tdttQ8y8abO+nL
EhcalBLc+tR51LmqZf5nhscUxAPpv3cW4pRJJS8avqu1gvH+n6rWmczAxQThGX5hM5/1NvOocIXw
knBJIH0jdFocGB8lWM4R/aW+j6l23R4DVGkvUPxr0FcYqdhdZK8f7dEFxKsV9ME2Lnt0ASeRI93w
YXC8H7UjOq4ad880oma0/TTgtKO369VInm2ubtAxRec22cBmf42/Bv7ukTxRgKTVVl/tqjwDvso5
b3Tn3eqX2Pu2sWOb64e80gl23cZ3XnRYib8aGxDiyN2WRHjVKUR8cI8mkwUA0lypqZpcm+lGa74X
G2q707irNCErAQpbQN21Q1XOQGiPJ4t1RNiCihUUa8jpZNg/wG5L8ThJOzK28QAmg6uuY6doHQZ+
wshsJGDgIlz8nnax+ph8CSJWTj/9OcdgGXW0QjECP0Lq8z4w/btNIY/L9jWiO1bh2VgGVpoKlkRS
rK4pSBBmkEQNYfUEZPp7vKaZpxU2lQo6g+CuSOakI2sY4kpBhPL4uW9uwlNpZ3FJHYpRa/0iu82b
oR8gMnSRtGtSPI6kTjJRdURTocIlV5O7yHMQFiR9qAKDi1tyalZwHpe7oqt8MiPBnk8w64pdH9Gw
2wbnzLSww4XOhaTVymIyFL6JRY4KP8WDlf9nECOvJODtlF/fwG8oXdYek6CNni/4zL+1pz6/wd1+
/3rdgu8aO7VHkssY7xzSwc/xdvuRxBk8qzVxk8unWR+UQy9dbNysmIstwl40woLP7SZodSbwwHLf
x0WRMJIXrKEt8nkodb7Ho3gxPvToiZP6jzu1HaE814ZTllr3OzTZE+viM8Y+lidk+OUyMiAj1Dwy
8AkufW7EFRgNV55nmTPoUNYuuTLnh1nibS1LdZ8suUssoGBB5Glvp3raPBJkwEGYMlymW3QesVeI
j0nO7Wg2GpX5rgR8eOwLNlIodOqZlyJb6rCbQ98TtidJ4Np4BfFfQWkI7QeHVESJRWFHP7DZr2p5
CE/HinfK9PnIZev48NsTHkSifvKEthsk9/JBMpWJ3q0l+p4r1MRo5yoeh7yiCHzJoiLTJToSAQjW
S7PSaP1Boxh4sL+6QTrSszA9whRUf1Hj/NRGMusMb8dOO9InCCVm7Oem7faGxizxihJOwdi8XUNK
FtNUqv/W+CoD6vZ5jSS818ufzrytYGt9vBaHG2B4qL6t1/RAR9H5tYJsgJZdrAxYUG9QvDxxUJrU
iWAfv7SjBSancePzhKprytBVgSxWNDdGP8expbZM5X+vU0Frhr0XJSAVGHhgpU1MVmWizQe2EDAH
Wa09G1pIb+hPzCyOSfRhpaYHUuBawLkbhb1hFzYifq8HPNwfQ4POM5Zj6ltbUyIjnYYLO9yC4+s8
i0Q6pCCvdOALgYU5gBmX6xbbrriNErTGye/k0gsl8B++rj6R8S2UBGcgsQCVwSVbGNLAH+p98LBl
OKzf0mjyf4n/tFO3p0KNv4mSUv/Rg3RBLNXHYbSkS3bFSvzWVkFblKWhv9NSiem1BoQbymfaTKwW
qsF91RdD1E29orxAZu+paAx87P7wqA8nukxVST5I2yPd0Kb4jYcZPfoUpdRI1v4zSdPZbYKGMkET
JfsVTCsygXIMetXO2KNJ4C8ZAdWearwUeosS8uxUKJvdupX/mNYdGDagrQislovz5HiuqmveuiDm
Tf72hQ1Z9k6wXoKaEkexAioWR+EjVgPXow7TSJvawm41CCPKOuteBJjqjrhJ/rHjrme5S5BVVaVi
CRXmsPEuXsReb6dFRi5pD8+dzuhtJVh8dRmMm33yHnsWHsiDJc5n+4Ecu2itMGiH+Arb11K/fctk
AENJSrjQBGm1sV8mu9OPpXCdQ0XNNnTN6KDLo+n5yBVcNmFqfWll6a2U1eOQDHOLlH5fchXs44OC
fz5Cp19SpSinWglyZctJdAmAvp9xYPis7WcMBT8qEeDI55yVmi+fW5NVMBtDm0qloPQ+w/CWlTMt
0NT0j/PvsXUAJZXgtRNyYW+SEg82E9o6M2hesYwC5kCJbGbLwL7sJUCtHBgsm3lJLyV+QGBwYj8Y
ssrVK4XWaW5IUU3aVhEPdAhDOnfaelj1Z9wDqRBYnil+ci8ZZgrSGW1plFBdeQhEgzDEgmaPmG7z
JeIgb2H9Lk0ZsLx0h5BAWVg0LMuCeUK6csTJBthY2XDz5igLPmvfmi7t/+OVPIfM94ZsPmoYV8RU
pCWaB613jYy500TSkW/H4dC3viCT0NepOBIIhYgXWKi6XJ4HAY5wQOSJyHI4gI3sbk4JWWN1ZcS7
gXA8/+RbDGAc5OgCSFeVCpnwpsxMX3ZBipPwvPPAioBl5BmGHhnUs/cWx8to8abk4Ngt1qpY6Yn+
cVTAQwWxPAmS+zFTBZu2y7BYcyHRzHXVaKI36ROCxvxSdcdoSyZYmMe0a5HYhSYpVhdR+1Hvl1z9
fxWr2Qz5qsxmXNzNBcLjdNTj0AOkcbbIklbiSXH5cGOxjuT09xSwh/BmhkWHtvxYvmGjKmy7Ch6H
TKBXwZnWlvtPRA26KJbRef0Xc9sX/q01ia9pLjjTUwmo3fSFGeDBuh4eT2QAU/pbAkyX3mnnFug7
Jfz51mH+qEawWi7VeTCw6ceUeT5h16eAK4vytqDwdFcYIWR/mxk6NrSD3389L5diUDCz4wIpfJHu
Puuj+4twVZNZZ4dETQLzr8CVQYikLDoaINilkrkR9K9DYt0Qe0CnJ9plRlu/nGhtwm7r3d+oLl7n
zaTFCFLvNF/IzbOkTutzyzTiCEwuIp6NdxD1cfuKdQt4Y/EOnO6MW+LE/ymEOkArJd2ns1nl1GVJ
Q+T5ViHQ5VTIg4OaFRKpK5An/hWGmzxS+HT4z192aPJVVN3wNrwhD/J6hSZyfcmuYQraPi9b/vSh
N8L+Fe9dYShcBBLLYDgWSnxil+wmw/lVue56KkzwG9V8Ckl/4QzlapLl+vr15s8QJRsWV1nYiCcq
HQKtcEDI/2vnS/liKKDuCwwhWyUyupUssUbDu8fPK7dLNTaZxPpdj20ylhNWhoAsgO6VwO+uM3/q
kDW0D02hsPNA/tzJbNsD9MWo0Dz5t9WLfnundmfgU7odj9MmlgKpk+E5qHzoYbtJ7cqqidGSGYFr
S3+lI3BAYvgE2OGmjRXLw1GmslEy4ypVMphJeA+k7oTyBag1pypUgkhxkVO+DzS/3MD9p0QEG+l1
+tu4tj+VW2CJn6lbpAfEv9T98qQ5MlLBc881DmLNILNxGZ5xkySNyf/CW3QfjndHo95w5G32bQJR
iiaccXtKLp878g4JloDZNhRvrqZ6bJlW7Q8d+iHdLYK60Twasp9e+zE9JlRHGLeBtgEmt+ICrtcY
AvGVu5y00bXP1ld5ZlUzTN3UIBZ2NLMfBEIsER8iWSzImyHdlYUdQVAL6VWnfca98QnDYugn9pnz
2vifhlPHcgGwerKznQqloPoZphvemt9I7ETTc1+0eSYC6SDdjhkIYO3Ft91lmAHHxQxgR+pnmRKz
m6zue1KKHhAhkOAgWXeGavS6ksBD01t4bZrBVD2GBy7wpiAUy2wlMLHioTKWuhAR6igg3XAdQ8bO
sx6IeL+mebo9ak3RBnZ5Ap0jFZlsS5UVd6guE/4EtM1EKXmH/i3OKbmBn40fj7rAVbakFuZtfKIt
2yjTka5SyadVCYmscXEVY12x+OvlSPt6DHHA8uZSB9iclAl4A2i/rXugrXCyd1ZUlBmDwFbx8Crk
5w+DJ+/PFzhKCbgjdm6Qgf0iXiXu6jsUHSRuwqQk5RjEoa8pFq8TPsE0kZAZpl96z+3jhHai7MDb
mMHTxrnNrwRXtGXACIYMWt0caI/SDYAed7JWzQeKfqPVfouGiv/VkvTLDMjJi4DebIOD7TaZGED0
LRzxmc2+kzdNzJQWncP1+XkBu8wxWjgvVCqi+7AgEXyJx6SvyB/8/WCCAKDXd6zuAx9UhfUK5Fk6
F0Fe96q5ipKrnXYh62SgN34b7ETVGdhS/IuGGZKSG7a2AT2jwquOE14xAHbq5ndWfI/qKGPZa/zk
rD1gjBoW/LZkAAIwxCiRTOOYt/R8xmm4iIfrJq1hVEgQXGb0hMlctPS8+gKGFJVlZ8gQY/gG1xqU
Rgx5g8FdE5fmyxhLAg/7JkLzriz5du+DZS0d9Ghlp7Mt4FB8ezLGFW+AgI2teDDIXv9QiAic/h1j
BAPVaQgoLkWlANVmKTWu93jisMBj/gb+tzyuZQNdJzFB9NpMtHscQmAfvaIeC66U4vkIX3rV304k
LLG4FP1D+U11K+gY76ptzMBYJKK92sKzMmT1siI1661qBpQHOsxLhElLeVMCjNxgTHA3pEr3iv0C
k7aJM03B0ipVbljM8zVAnlw1YdBsTExrPYiZoVS244RQXvaSD/3azEJpWY0x+up3JcNVtoLb21Mb
bKLlk16gUgq8RHVLZ+haGRLUwbln6WfEk5WBlqJd9rFID1heh94I+6/Xdk/fGiofIEtjMCWom9K3
5PFZ63hwGNcxsveinPQfMNf/Se8evbsWbD7jLFGnSLCbbuKVTNfhLok9xJtY2I9CyJGXtBOKmvhL
1JxfBTtux0n0xmx6cwzG9sjFPuGa36OfEiDncDYFwsHVqCXxBRyEOtFZ0uBOALrfPFD0S1v4KlqA
tU3xjMJ2H7WEO5QiyrhKzhEsLC4SG9xDezgk2v2s6OtvDLz0nEWLGIasFc5kJX/hLxusRPRcgs7v
ENuu3upjVnil+TPf5VTz/3LhePc8LKAkzQFGzh64hFUO9+82KnvRZ2z1vdsOCPkw1m6DUo/Wg1UY
vH3rLkWU8HxFA4g/m0BCSIULZVT1sg2nm74eISztSQqNtvl+zYDg7KBIMvyJjsbLoEP4oSm/jnos
4MB+hyCEKPhM7bFaXAD/1bVfNMuyKb6iLU8t61+bSXnXzbiBEfu7kCXLWBVVixm4u/K+ANXzdqLg
Jhgk5QRC35BKI6UA5NWLr09cHJfY+B1XXkQLbdcodGAl7ulLiJGGekSdkk5g5YE0pGI99aLP/m5O
b0hTWWQH5lj6GwVbNv/5Qcl7U9ZSXMRlXUX7bz1PwtCD8b24cuJ8jShBHt16CNs3KaC9Iy5my2nS
KS3Q0imJj/4GR7VlUuR2rs8UeseWufpKqhgDf/qEk+1B1ig1LDxxDk7VP2/dOHdUzWo+QmpY4W9N
IHrGnPZ9YZzcIDT5j5aNKuWauqv0O3DL937gnOlJqvdrYUZUMqVh7UmKHlRB00AqZswpP6HjXBJG
93RWi6p2uA33fpVMRWhbcG+lDv/orEy3UAB7PUSzc2/adHocZSyk6DDR84ixSuM3JKai+LJYTaqk
KRw593Gptfok4pP9rwhvpQVjgpwF4Q7R82KsMgNURyBDcZAF5plO2EJ2XPRSeMOOqk6zkU6BrD6X
nSXKNjsw6a8lkRVugSjAxVLdfk9xMPVUA8/KdIXJSSumeCTNYpcrQeQk2QgVg4lzSAgbQQPrVkHm
C6sf5ree98ITUl/vzZxXUKqht0QUaX671+Y5/CBIAcPm1idotR/Ngx+qPaSy7swfYX33kQnkTnm+
kuu+veI4mwMzjRTGDJ5ztSBERAm22WJVvCXuFBtOXCS7UfR6ymeHEV3dQtUHpQ3jxI5WFu9ka8lK
Jhn31DIQ/rmNrz9NdXX7PlwVFfJLkk8Rv1wYlMFv4kRQr8AJaV+4fRV9qk8V8Qn63TFz5rGJ0ULl
3WGa3INH/hR+ak2tM8UQbLYLl9NmR93wXZ5aDsBPsfgQv5/A36LS04Dx281wQDFIrUxdhCbIoI7P
r6hwwVc83P4xpt/IMVnIZJvDR3ZbmiwbH0OpdcdDKPvqe7+a1sn5t1MxODUf9uBhIAaek8kBzqSw
LxWCb1c96YM4Z2YSyQ5hDAi54Yt7U9bjd9BG57V6QktDFMkxyN0GzBLg709OSx0lWo3oz5czp49f
R2tKHlCA4DgW2r/guK+UdsMuwnJI1h3pEeb40NbYbx0FEJmHq8oaarzpPR/xyTY2g3JY9fbniG//
yAOqJmw/1SarUg6PQnlOJ8ejDEwSokmbUrZHCdXwJnB1NtEdFKIralFfos+QQinQ5BFSqvYI6FDP
yNeV8ePoFF8uDJ5HE9ALt1FEzL0JdaOWQy/inqqhnXGR88XAEjsEctQASlJiqFjXJOaDIvaagD2C
sA56+WMQuivgHeD3jlf1bRhxwCf+KFg0d9RzTD8f1frpW7SfHpv0cSCH78zz0Hf1P4vhrBWR5Sj+
QVA8QoveNwdlbBLseUJJ1PLvA2bCF9SOLC61wmBzE34eASR8RGXbBuByvshokp3ksbalNqBRCsGA
fNILFX7ib9+He8pRImAXXGZUwXHIQ9erdOXCj9PbHwcPLyPcYiDNdTZdoFmcrKm26UX6Z1IIjmXB
S40dvSxQQAJWzrpyfob2Vg3hJ6O1F9wTXkXB/sYykjtoUSwj3wdOXb8GPFDq+I1Mn/YIQGFtN0Rk
IZ7ZAmsLtEOtCnw5mK3eNX2VrvXa0sSxsqtT7IASWl/IEdVn3fbWYmPT3u/L3wAoZey+H9XtkexM
x7/6Dbw9+fXx6uA3+X/cAJGn08R+Wyqv4An3jgdJGyYfEg15RkvT7nqALEIbMBZhpBP6l6cRw3qR
i1tEIS/UFHfGRUPdyyzEk+fqgj48OnZkIWh6WryLlOW/7X+bEezRlxetJclkOAPkYV9+LC2H2lrK
MGWhKVCSnF0L1TVex8WKbzgEnlmYzn+PEB3cSnIx3P+OmgpGwnN0ySFdME6LnYWw4F6qTUmZo9nC
KVtnAdDbUeMp51VsxbnuM2cC42OX2VIoBr/tqLas3CIXujjjG8utzmhxzG3g07UpLUk2VTv9hETC
1P3K+WyUf/B09L9dgc8avQ9F6BmHW0k6rAq9JEefSl0QxZuLJwMpAryjt7jhG0ABCu5a4ccm7hd6
gGvbRMbXysk1VzsFrMQalYqTqYTj7wQUJUZZK30sCxmIzPwl/ZBdHJZM1K10g6/He2H5E1T0eWyP
q1K1d00t5UMah8D9PwjHuwlaQ2OZEEXslbQu/EdQn4FGCYvGeETEsO2N2FXXoqxiCPVpyqxA0GiM
03WC2cRCDIy4XPRAGZzuUzJhyLmEyx5NgJ2egyvcOx3lipdE5DGsN6cNKVmSy0WypxBywg+WbmRa
spRrBoE6Le5DAPvkRFWQIezZIilM8aIIpuErWoQGJcdAghADe5Re9pqGdJaHIkqPySOmSg2i+aPk
DD7fxmcLAs6+F2wjdbmNzsGYFJawm/TsJ445uvVjUx7ZEeMlisW46oMnhZxdbUfRH5lL7Fg0PtVj
R8droDXo3xZnc7sKE5LUcwyzDD7ySmAYFpL9fshZwSQd+Dl1gexIBPoGc+VS0zZbK9UnbM9805gp
MBf77sZDXwt/zLENsR/VCM8nqJFOgESsxJsvWAZCQWtzXxAmoKCsd4hANQvv79geU9eNpwBC1R+n
ZxN0mA9UjmiOmkRN4FvlG7mlSskY9tvW+uiZSttNWI9tIgIQ07Pn0v9JJ6jVWWxjVATQqSWhS4ey
ByLtwFdsFsPrx+dtZhNbDFmSK7p+90ESEcWfLIggU14Zru8W3+nLFxLW2L2yigNYE2/X8yzYLoG8
ReWUpxmyk032mmfmn29C7BzW/QDzoxZkkGpvk/Qbk+Sk70669hN4gDiANuGqFZ4YyJt1mnNFYKZg
fA+qg3PqNeJOgDUIHWR89ChNL5QkHTZBSAVvz30kKUDh2eYfwHFpd2/Fet2M8IrYqfN3wwWh/kNS
9m6RIDDbNqjPso6PZwXY2nD6xwIye5GYmY9R5zhn5v78Ie+4lwxKAr5H6E9bjipDmYoKq1bRDOpV
00uanlxzTnCSVBNdZ/9pXIdp2qzHm8u74rb9T6Ug8o4C3ayyAOgwlNwPHP6OrpnNX1xQm0WuE6O6
NC3MQsFBm1vpLNKiGzYemGeSabaP3encig9UhUn1VymOO12uMiD6zL/ZnCEcRR8/jG45qlwEC0MW
oRaqEnu0UJQoKlVL4QyNsJj1TTlbSpWjfxKw2Tk7jZUEBGA95ABwIRDDpgJ5Ul3icSI52uwvGjmp
5/XMgzcZPv+eqXPs9n8UEfLRMhVMuoCw4dCILd9u3Eq8r/x2I3buCJefLVhHeHoMzBmO7GgGkApM
pb7ZtwTjECDPYJuQe/O9P5QstDPsRiOQK9oHQOqyMKeVYVeXc/hmKJHnWJKk/sPzHPp7ymxxGyPn
aOPEmEKBJHMApHpFtL5SYLNn/BIeFZ8j5jaLSSCNLaOdgPnsUe9bB0BhYVyHQK/ntGwC2bdYsEhx
Er3gAY3y8UGWjz5qKzvRTJat0scTt7f3D7UPfNMFZY32blcweVcHk/hEU+4xFpkFNV6Kqm+GbQVM
Y4XJLr/JljNVjJ57AMyTs1wjl8ZTdc4XzltB0Kh4zhWdtx+UlPmJvhRmFtAfDlqcqbFHUzkCpyAe
i/QYHAjMpIb+pm84sUIJGzrfxXKgPL+ZQ11c8RCGOQ/UjDLOy+fmjhcIWUNBVKn+w0tmugSzDa8r
yjVhYi3cgjCtTKSeIDIbhS+GZ/kKfxmu24sOm+M4fV6HQSwMtrlv1nIamZA8mR6YjjpIAr9pVlY6
sx72LLuPfiRE8jXIAr/e3HkbEzQDWmMZd0NmTMVC7H3ysNX59b0Ajj3RLIofyvmb8gdllzMOtzu+
7m7nG5Ea7/GHtFMle4DnX8GLo/aGu5fnem9dnpuUpcynznJCsHGiuQrswiAxK2RRC/BP4fVVEfM/
A8H6xNZq+qPNaB42r8Drx9ugezDIb1hKtzTp+dflC7BoFyK1Eae/1wQvdQ4AQVs46DzSeAbp7Tha
PXJ+3AeIocT20c5e0lYYCCbFnMVdHPvlTlwEQBiEbP7JPSv6NdZmJZ6Q6zq+jzARURRgDveghqh/
gtShpwETYAakAXrUwFFlqBotO+hX2GL46l62AtwzRuE0UXpKbYMBsh6bYD2JKhHdS/esqd5JJHmT
XFad5HmP82RzRnnfOnVEPG85A+I+O6zZ9xQC1Dl7eLVMaoyhqyS2FahrOHBtoxynp5KX00oa0qPV
NXdMdbs2Y2GQewi+CUdwKLLwKhpvxpghOd4VvscxKJGKAmEMy8DXyTp8DNFz3Ff8KhYrXNBaAQzT
tH0dn3nluYT6De23ruv5mFvAR409UXraNcZZBwO1z5Y4mE1ltNQAjf1/qHkIQcsKZOI8KLA7GzL4
URJ7cpLqBe6DA05M457tVCM774mg1gngSas+KlaiFiBhZzOOsyv8jP758FhM0qTdhQZJwz3Yjifn
a9AqhwG2BJkW3dUSY+7w8W11v1PX7z4OaHJtriS/kPmL3wW0jFsC8EiAm2ABNgKcOMP4G1dm9NyH
0Hfn5m0QWA8pl/8M5cxIEG3g/Ej2XxxX/TOKSs4EHwnjqOaV+OMUBsDg9kp9KTVSoP2igGU9Yipt
ED0f6bgWU75Db+9BoOKkrUQfAxznE9a4KOVC1K2bO7DATXcvIcKdqqVXpxopVTnoh/dCLPznfyUj
xuBUPPX3QtqcxnV/3ZziEQ4eP/U3H+0TtaV4ko+dYBJjnJVy95u+YmcM6bNz++Ra6dnnXDY8mWXr
woBdWkz0pYup31h+deJhgrur+KmLnrmmX360M9gqMn4t2JdUFme+FrWqskP5vrgbGxdDHeOIpczH
pGsHrs2H2emgAy6j0vfyGs1vCUD3zmFlARfFOomrhMv0TlJ2eNQcXQKQpSCCa/XZzzexu52TY931
JY1g0VoqYnpHlRDXEVmzG5dABr7y1By8NAgnHKMUWPGHUTeR/Xl/Ep5q+IWAAYEqtwk4bvbKDkVN
Sd5Fl//uKUPllJQyh0RT3IXRk5JZhCvl/7M7YKCCf7zEIHLtFpAWulH12gLsHJdMu0vZecfy3rev
InESN6dZ1oIS6zBMAr3yDZDXfqXHcJH0AfwcS56misMxpkG7DiwH5eyN27f2VqMjBUCoQUcy95TT
MQWgXx7s8qWna0/g60vi2F9hiIuOqjNYDTuluttDbEPygX3Tl4LxBjfVmSIXdb5EoJ9BL/hl8jRJ
oZgBzFRxwlwKsNrfYE1q3j/LH41sbuSXLBJ4z1PyLiOZPzC85jJu8T8ObUE/8G1M0DTqZPpVgS8A
lnNM2wAwK0SOcNNhez0ZX6IK9iIpHIFCZ11Irb6z/SQytNIAJ3UkKnItqMamRmH80kLSLmNafqQ2
pDLkVX3zqYDMrbgT47tVafDuwq3VipKXbCvEqlMomESBfFbnovh1cMQScGes0Cl/nd8ICzEZecSs
EwFoxF95TcuO7EZgXMVCFjN52bIHEoOONsKHGx7yGX1EMJlIPCnloO6cipxCQKjzbUrglqXAvczW
S3uYwfgDS70195G/rvSufM19uHXPT6+vMe87D/IaWBYl+IhYjsB7ugybpEXByH9TNMaXJkbIYOYI
fqdcq1exwAe/rEgndoxCaVYtjtvAdUx4MPxZm2JOUPnPrDI7SezpqoyBgj53XLmDQAX2QT1VU9Na
AnL030he4E6lPxK37bj3m1EzUzPTQStRnIN82kl93NeMFAj0fvLYHLozaIZzxxC0CzucQZ25n5rv
Jg0iRuNZ6HDIRPXCM2NPTCY+PAej4Kj4ekbkIyD+WetYBkodOHb42ARC55pl5WG9r9wjY1tUicVM
o1HqgYoMG8l7vHnwIIufRn5zecSlol2ZS4lMWWRxAGrXHGfhOQiyagitW4ap/9PiDA4r+GMnkZ0b
wl3HhEAJM0ccfjsRYTd1HKENC/C1ToC11kKl4XMONxsWU1GmNVeOiOQpxDiLrmsy5GW5fHdcAlEJ
DWkB4+O9KCCMOmlCrsq/cBDyYtzubJd1+Y3RTOWP0JmLFG1GpktBwYHghdOxkHr/S0JRiJuIN3ng
+gRHqIPZx50B5dHiAldcAmbkhwBTobriHrgKRG4nkEg2UMMMROeKrBcfToIHF+5jw1p+e7XsPV9a
XilnI+ofFNP8StgQwCRv/kUaERluD5vcvwKX1cYveerkAAtRy3LkDo+DwUN21I09WcP2p3XDCfeh
qdy92RHW7uu5nWw/hQqsrApal8Z2V9T1h4Y0p+NkdLSsuI6+65X3lRQz+aa+REPmJE160CHxKUBZ
LzpSpCsdHeLQg/iH1ibybPaMNw8YSKQQ2laPvG7vskov0DeQIe41A/UBhz5Fyg+jhWqgrFusNjJl
a+HWtWe6vA2Okqted6TnjkaQE3DIRVqpPapvxVrEby9WifRSqYPnlUut/4cZhu/GCJYr9q3T44co
Gy1BgLf/pYMHBvjK1NLSHBxSOx6bomyMRsYdp8YKbfzJTeZqcasnimHNUPAMR2OB5G6uX/ezrTVS
chpJ6UX4mxDBJjC3vWnUDqJEM2QY7ib7NIpwUiAbG4KtM9HRI502up1wlhIIn2Pk3A9Z4G7vteJE
dRXbYGbE4nweiFn+Ey1eyOjFf7pqSC4RmTqTqGrV/i3NC3Wb5XbW8g8zU/lvFNjK49oc95Uc3HrW
yFoy1/G68QGyvFZ3p4ORMcQOakJLYOL6i/5mOFf5YMJjo1J9HMbsJvK5vBgoWjln4hz+ey1+i5FH
YOMbBGATMMk1efROQ10PyO4nPcUWSqv7fT6fjJSABX9Fwq1pWccyX1d0FXeiSn3AzoTYXkJrIlXT
tAFcr/mDuMpJRzDP7YkilA2PpfE/821XsePqBbQS5QPTDFJLDLUlS4PrjPQEnQ1Gn2YUA+4fF/6/
B+Pg5KluELhiLthl21rxr2NTFZ/p8X9OTk0iMofHX22TgpqvsnmERDU8IJ/ufFG2/Q4ajVd61foM
+4XeJf4AtWvJoOGL3BR/RNSoZwXEjcp5uunS+T4h0kJJJIPdERFtPT/+bMhjwFpLJnvP6ZqjN4u0
2J4j0Tqy7N6VoJlrWPsXRmWEGqq8ZuBDDEvXgr1il90vSsa93AoVa4MBbqSg60LRNNmtR77sZ2ak
CSY/+FyQYcIQzfOOq6TQluCS4+Owza8dO0W3B11BQkjpdaB8/V+7M3WvGwHYtUd6rKUFmyWZpdKw
njLMRPxuO6z6BxNeE7lIMhtlIf307NXf8ECx/pN7ZR+1opNWdARjnp2huXjaIDpTO3jIeyC98fhh
H1M+rHib6YeyoxloYj3SJyI9D4QFcW5/HYl6OzcJfV3hH8tvE+/BA0SkZHCqDbqGulQZ0gw14Qb+
6gH3EPWl7HsH3hpRWpq27NP8QRdjBz6Bv6XmauJveRNV/vqqSx3XJqwUGC7SQXrs+m8tBmuG+OkN
mLYvrwJ4gcUt18UxQ0DQMQX/ZYrXIOQavcbJn8mrs1e/D0mmNphcdR4ngEW7jHtyN49YIriuDJHk
sJlxYEenXD+Ej9/PjfgQRuApgLd2RuHnoGMPqN7cwCdLhEaY4q+hKdsGUSqVDO65k7acplaEo9WG
gMsZw1L+nDY8oGy4CCPO4RWlQ5kjqWKlPLxHPM02d+wQ6F41W+rOxxcZ6BiF0pwGK5wRR7WmVC20
zQXXiX3Pmp7q3JLBSbTEsci+Wb8QpkDkB9dns5l0N8bNkpNaxNDa7ROuVecGyzcIAd2kOhIJduMB
fi9aPyr3oJtPCMjIuK5/eAsFSgGZ9qhHX41J5p6iy0fYPi0EfcBse8mKMilynEjzBX/6vJ3JrCt1
viMryPGKO4X9lEhXeyyx7QjRUFZUsm51NPUz8kW6ifOH8WmdvHhe+HcUhs2+b9bmRmm0QxP2cb9x
HaKuvamQyiv8JPrsLRcC/7IVCuunfJ8/I+dlnW8iJz6MWMGKlNLAC0yvfXgSEiMmUAR7lvj2wqm5
btecjn9SIH0GhV2ThRvzmqPp1b8DaxuwMHSA+UCla7k+HgbyFRWa6ArQDz1VYAddWqJbQig9Bv39
rcmbuhDfAyxEX1P5Qrrikxhx/fBUjEODe6ScBykEcbOwhoHSt3NbPUvn8VdcGJgVD0MOgpz4wmed
w6xb2PZ/yrE8dqHet+F7wuHMxR/PgL+obxcWC/VLI8/F9/xkav/f15vCVRYvRHjuxVI7SItt2U/p
z7iwZlX9xXVJxlqcv5WcBnYie5WKZCWH4LgyRw2IzWA9+Fuccb64T1CKix2O4llAq7Ac1dIhLZ3W
+OQUkPFZfVXoFcClaSrxEKFFu/nNm6C/KKGW52WVu3/lRMYJ485vKqsTykMphdzGvjmel37obg+9
GA6ZvpJS3YDygnybZYxTbKCEWo3hsQFjzZxvjdVwdx144s+iv5aVT+T9AN26fsNq3HB5NSDyPQkf
0LbUt3vlx1wALAKQ996jK/ZkMJN/E7X5svza6L4EtALStFIReUrb2p8DrSbth1pFkRmPqxQXCwiM
e6TtKNvmFL17u+ZHwA2MtfStQaPJYnwWvZvCUBAzU3Q400w5t6bfRnLBLDcqDJBtwwrRdTyp2YOy
LDDyRSF18KL6HVDLiIkh4K0oQH2aMGtetuG/p3F/GDmWu0lzho2MEZH1MZG8T2rU46R7TuJiMlwK
A9jM3RRSIodNazGZxNET7DWl16dpE+07ea8UhAA0XmYggYD+YXnnpIwT1z3+d7bbK+PfjBhpBJIT
Tyd+c2QfKC+JOJUgs5/2gQTt08o1jL0sGiYI+WyyZ5M7a/Q240VvJzpkQQBxlV4iz1Xv9AyWrzsr
tr1YTKO7F+glN1ld/pEHAVExWIWS/DoxYx0ixhMS1w+pwjJpW+kTCWhIJtk4QJHRf7N3Xg7OGg8f
b6GJGrMF3vcq0J7qCjJOqWg7ERXoQbTWmrn3yVobWDO05df+0zWJXFzWRVWV+Bc7C/lZ8PtG9v3v
fAMjd3USfE2FNL6NqJm0JIvjGMQ9C/2KrDn6dBGcC3yN5ZSxkwgDdqkLFm+cJN1lvGcmijiCgRTM
50zpEpzdID5kGto5nz7BEW6HLg6wtMcfSnWcIC9ERoU8D/YcEKJAKgEZsjjQQSkYnBhWOIu9R143
nUK1rW9aaSVcce5blPcFOaKFGaXyUfFzde52PQc8VuMHjiCP7ET+/zpExprPzStRhBkDwnXJNZ6E
O09jPBIcCvlZdJ44h2Px0vtgURhcDPg2czstpxnQgJ+eevxTw1Ao0+y3/KTyS49ZDJ1zCiP888p4
LVW/xt6c66uXbodR/RJH/CFR7ZCpvuxBFrRP9ybchVTaYD9YcFvjcEJR7Em5D+36L7XXu4OyMsfx
6ogC+vzVdCJLXGznpouOnAdKhK4QWeC+Po2Oanq2Lxpir1xNH/04FJWxwcSFKv0KrFCxqz8cxMzm
NtBFHEpZGm8WDjFGbe75oyORo9+2yid/33YnbHPg3CTzQZgN7pn3V+jM+LHpI2SEhw68Up4cYJqJ
VG79NsnAm0ih9HOADBWuMl/l+brwFnd3Q0hw3Ux/i49yJPf7lE7C+Mh8ixPfHFIcYSaVU8JnrpGR
a32NaVCtxJ5GmGp67BRjJM+TBqdBXZxxJgCjvY1Tx6UNy/TIg7tblnPVAuu+ZFUDEme3Z574H3FG
80w6p7Iw8h8MpfVYozpg1sKg2YMSF22jicD9FQbon0qKXkgSySC1euVYr6SRku41db8Non2ubtcu
DiDUf6gUA2NZDAClFJ0GcwL9n9F/o7yky02oJRT9RtZPZ3cP2kiBiPIC+EJN7PZ37o8BiPwNG4jW
WxJvPp3BzpyWA3mU1BePiyyzNJZS80mfPRLBk+wAW8HC4yqFcPERVHJr4k4ZPwCpV7YdY7vPbjk6
LqylQSPL4viaQtSBzeD0UwvcipWpw+Tg/tEwGIYyZhI+H3UXKA5Ploxuud5Qu39d9QOrvFWJCQZD
vN2qL5kK9NKjc5c/LaGLshW0SU9B2VpzHeMc9ffDyicwBPsM6pXmG8S3lEDds68IKkuKHOxzpUNV
FAtGstLRl4IpY8UTGzoarM8t1shEUpShDpEGvskSzwIauDIzJ67maRH17Bcs/sGgUoLE+PCJudXM
GapeGnWIMchL1Z5HY8S0r349fHveN5qZX52WF7KcEWJJ0aar+LBsGKO1nhZ0lJ/WNOjI9/BQTVC4
VnWoD8pdzS/n9WfocE1VGrAGQizlNJ/QsgjgHtPJI3R89Wpx81BYFctDhwlx5+X0w8kHpaTqjAT0
zATZ6fGNFjZuS38nT+tCD4UwpC4p07YsuDTL/BGfKu+oj+27G3M2Adzv5smbemDFYnyeEGmRNg5l
IRr5WgxGyJlBzJ5g2Rpw+g53zQ2MHORFT65zaSLVkWIRDf3+eeRiqaU1UGzkQmoFvYQZ++LSMjmt
C+K0HqESlXFoY0K1PSnjql0hAymarAtcX97BynUxndWuvE3gdGmN36L0CbUhoRpl8DNBpFa8MmCz
UnY3ZyeLOdNkMbZhNIjDELbrElrgIM3mAL0PaTZyNQ3oUcptQ6u8aFK8MVM+fL3b8gzhLVzFsW8c
YXLJtT23mHb/5A83O5lv3FnRY7g1nRVJYEPkfj6z3pl3SpPL0ZYQgBUvd4bjZsVzgmN0NwH2ISch
wwEodR+zQ8p4pgJKXJ1x6+x/YJXe9605LoYSgeHz65pYds+xVVwqo8Sgy6uzi6BIBNdJWcBBHErS
LtZr10UWVSLjMTiu/gahHQVNThr0sx5b0707ZzYHWQd8yCg55uc/BYOWuOk1DB7Bsuv2/f5iGGQ/
8/27gQWXOXm/w/hbTzcepOXoYKOD0yWVA7Q44E4r4oU7lY1nQ8Ig8j/E3pfTZ8Pbx9QbdHXhOyqR
bl0GhTyRsA75iY9QJCHX1wqGUtvzQ3A5OiOChBklaGJNnn1wRHaGJzPOKtFYQ3YHpDFnoNM9qnKV
soiIqWTOenUDhpehcqt8qmUCDaY3wuSf33HjK7Jdx5F+LtxSsq+wcJuFKwgKeUFLKs/aPPqUGd8A
inP4zsLIPzMiBAXrSP4kcu+8HR75tdKA1fY6H6Zf/E6w+iNc+UIsjhiSdA4LGyYKUwxxYJ6iw7p+
4nZET/YnQbpr51lq09I7X9e0yClGKNVYbOPWxAoFhUtdSD56NC3Mi4MFxydTkfw7Jx8AeY5JIzy0
WKCXWbddTJ6I8eYrTO/9bPyUZ51AaN6bumN+/BL5rmAWpzcitWv5Q06MYFsaRkUDic3/PV0m/IYk
oLaQB+t7RyKNXxk3+ib6qgOhOii1k/EuvuMG2Hd4O3xk5d6KE0itgxja5qp+syew84ugSsHK4zFq
XutfujfykPvgllKXp0l/f56+J1dk4W+iDxZ90VuRfrXCy/pR6ryElBPn3Pxn5smOehHtDJm7uSl8
vWWEWqwrFow+GGIU15CAfTrAJBGyMy3eOqwutQOEbsXWkXMgeqr3Df1X+JzXqAx85F9YVEBPPhMt
Tc2xcVQA72EFJOStuMJorHs1fkH7KXRZpbiTZQuJOSt7T4zeLRqO4wSeFn4A5omZtGxX6aPheYWA
48Zw4OiqVLKnIQod7ojjGPNCe0iHF5bpbnDHTS0bueSBbqC4hOELUo6Yl28jjuR4Ygc8b7tlFB5X
f1ShAHvgbRM1U/3l8YQUTZeM+/G4OJIhYOBiJr4ZQrTEJ+4WKxdwfWcFtGK+stAGzveDDPJvVe8L
z59YnvJd9ZeREzmTkz+FGtN3Ar/PKNS/STrR77Bv0egi8/S3qP9/p1Flg5pb68Jmm6r8hkkqcRTs
GSl4ze7h+rbkfQsKRVQ8QWwZ54I4l6x01JwgwQuz0tlbnG8x+D9mcn1ejUxKATAsR5Ct12ZAqb2y
XgUSjeICK93DZGL8WEqKnAf0AtGKmBipE8jXGtc0iD/7UYFDNYJKjrSGBXNBCy5OKWf+9puT/kUE
VGWDDhEeZoyJe6biNItK1YUy3FbvhlzW1hopDbzVp+GwOPhxsBJY7Cj0pBgQSjawUYHZigN237pw
RVp/Kr1AcJzZVDMmhJXuwxvuIWyeAGa+aJ74ye8wcU5MccQsiPXw+LEKJRSLz9hWcvCrQ+eGLFsX
7ax9ff2BWyceKoC186FxrpH1HShPFpT4oM20i5Zabg0Vmx3wgri4znmz/SctfjDvOKMsaXbcz0Fm
skZ3NgWsO20VXMIBd5LGNKVMhybJQsqAAddc4z0tE9g58BEoUkNkaY+Ybc4kSSWjhhptTEfecwCB
RF7bmeXXO+pW+QpjJRKfYGwr4dAOuiT/LLqOl7bHMTKcJv6cO336Va0J9qCPQOQcpxFI7UAG5lQI
9WNniwufM6zfq1V/3X7PpG1bjRPBeNlDnzq2PZ3Y+3YImUqJwdRNvIMoZnE4ldkkwvB9vL9ZgR7Z
yw+wx8B/srdKJi2YFeOfZ1WPv7eqw6kdtogUUEf1bgDiUKr1QQKb/afStLU59L9zrg5jo24WpZH1
I9UAfPoD+sbRM8+PXX0uuJTA7IlpY4YCpUZeTm76EzN9ReBFhXNj0GKFSdANK5K4L0WNyGWr3q4x
5kgXa9EQirwJn6VgcC8lhSYaEE7sg4glDIdtboDgSpxoRZnNvRz492U8Ms6zQtOvheCAA6tZJMQR
D0sIV7Qdo7+zDzBIgB6y3sbavAYdkSBvG++Iyv2hv4os2jAeFbhh0MyO6rrI9+NnlMoHU/hJzpVi
8dqpRl11P5eJzG0IuCVY9ubsTuWgeM70XMTiHf6O7ossiBy2HhQnEBBo7iIDAFxvoWACjlJu2f2F
v2B0tyb3TEdAM5ypcZeyfydn7HaPJnhJlZWaZCJgyY8gEpRrLI3VghMl6guyFa+Z06z5X1QU7tVu
1n947CxB7YToQuc3N3vYzS1L0uGEussasACteXYptdSnQ+QDrXDw/+uymmBGqpXeHY9BNuU5qpC/
sZYxZeFmh6OdJvX1KHJTv3ieuTFy2DSAeTm3xka0EA1XtbHJnGF1TC3V4HHUX/7WHzs3tvqoHzPc
s8dtR8oomRNrVP8y4lnvsLNP5u6JSuUXS0bav3q8qJs3EIcpsokk8WBAvB/LP2kqc6Ymhh3/6YuJ
luokMsNGkeLVQ7J7AEcsKWCalqfs8AIAXWDz0sGH5d44NFbGa9L3n6YkEI+WewXN2OebE+EkwvEj
O9S7S7emgxLs2eNqOCadGDkRCV9GkNK+fotDVD7P6GHNVwjEuSwFxw7nU21OqfxtQO82F/F+aIj4
/3V0AnXTr45uLhNe3iijYJ1D/BHbesYhzcTEU/ZhCty5uj1XMbGUSJ3TBIa4NPPThSyxnaR22lSe
gJ7FJJhaA8P8iPHYxd+4zOZopGKKk7pJFPsL5YBNxTBEqSYBeGmcLygS+KedxuVo51P53HEsHJ+O
b58F09AMirsEPmMvyQ6mPeh/Xvhl/Y1xoNSnrDD3vFr8h5KPUVGxzRC8IC7bKZXgCdenX+Sonlyi
sC2DaQVje0sEFIQTGaD3QiXNsdL148hA97zSar5vRAff15n0JbcspD8XNZ5nK8yFjNmcSMg11Wxx
ionAJVe9sxt6oRz6MdO1fxdCn0fgEY8TyfbrLFao0K7e2IERA1wRp4HNjLR7WYl0Mf+QPBpSvdkd
nyEgcHr5XKo+9qYOWKn/T1nbhX64K4LnRYkt74y5P5unbgPddyCgiiUYl7K9s9OXIvqrn5DI2h/3
uaGtwiSLu5DNDHefP+13wV++N///4BmoYoenYblZ93iuEgh1MtHjyxu7ejvpVlhyWDhwjcqz+yPh
9X9frjLAQEGvrhx0835m9eLeMyrNooSqCVXA/NhCeXm5+7Hb/vyyGWLkwkaW6fT7SZlUOpbFPJFO
/B37NzHCPopjaAHnJn4pTJRgOVC5fCNRbaRVT4bHGwaojkH6pXKIJKFJY18rGafyrKjLE8lAsPYv
gD/siaooGfXaBw3IT9FdR/HB/yWITFGRLQlXunImAlRMhsLIw1pBYNIkKNyi4Y3IOL35sZI/OUhG
kn8wLgnz4DC+0APu3qh6y4V3dPBHoD7Mghiwn/+Ym6BshGxusuRhpzhP2miLzo/Dby+/jylhP7gV
cf1pyzSikIq7O37P2CLUNwOKsuUVoQHu8ygJDGVu3fB+W7XgeYWKarVgUhBuAesjSHntDMB4yX8/
UkFI27Gcp6tzxV3zXWYzu2nMYrBoJxIPg2TjYaVo7yltrXcWWSldCNm9mj2Ds+Qq/3pghSNFE9nh
nOgwFHN//e1m0KC7LiwqSRY1+qhquIvgCwSRQrb7nZWT5IzgTpdn8eGGNvUVV37vaVI2zXIBU7nM
QjTtYbKmyDlJ3FQssF4AtXwv+6IYTHZjWeK/yAVCJHyCn1z/fx0nAtiM1FgJ+1KgRA/E07h9uTIE
bCjGj70VXJd2vIbRD58p/RvYcBDeritlT/5iYP2ZloWE2HM/8M70l8BgavUF1Q1dEIBzysZ5jAoG
96aGyGPMrkboMsSJmg+yIm0JndZ6XLwAtbRz7Kmlobd4WRfQva4nSSN3xFLggb5xhBEQbbHTCabU
mjPIBWbT/ODFo+8t/N0nOdANT3rH8o2FDq364hIe4OTEoNT11e6f14V5jvAgzMmSFHct+lDyM6v0
E8/88WOxNIHY0KBru0XQ3hdpcQKvQrcyq93ZhKGcqfgq7utENFO1cL+/UQAPrBjSqfx8rlZduk12
XLNHMXUDdY2tIW5aurhZBy+nERZIhIa2i95k5xgg5O27OUfNKXnkfOiVY2bqXU4GkXcuYM7RHJIC
cexnGRSuUMWyu+Qn0oJklUyjxsGamtLDH9ZJX3RA4ls7PEGq2BQm5zFRWaI7dGpj5IQpVKZ9Q504
Sr+dZHOugVO1Ulm+x3lHi/0ZQTv1OxkxQNCXwk3jrGMmeY8j2p8cQnbX7GNw5afGJDmm1nzbvP7U
219M/YdYP2LsEYU2l3Aw6JRkyUi1h8xjLB6IEQ8r42xoDh8NbiHPaQf9yuFTf295PJe4gZj63WBL
01B4LxE9jBmBVx70YOd181DCC0hKsOXS8eMsXuMX6B2NinR9IY+J2TRnpNkCT+9SlGHuN5flIuF9
FUOLgfcaOHGu9MTz6Kx/48RTEO9uxbPLyGbiaE2azDRjhcjfT3vy8/DJ4mhkphRSgB92JYbirfd3
ML6X8D9Q+chbC0maUfLQo3y1RmLv33JNOhRqPIK4lGcSFH0R/yeyZN9O6u6qIebcpo8O+PfCkGL/
z2HLwgV02nf8vKCP7PMQbCgj+3lS8zEQNFxB77Utj9owk9loLTkBhXLvnJ+oeyxjuFhxftxmXuC8
C8g8AGRw93uG0ZVkSRr+mF8i8JJUa1akWIBpB9jvuPMr61wjAA5+mfqx2J1gavMgg9g8ZzYZWGfy
pvRr/L9Y6MW0thjvUMIhCpKDM1CyQCsQw+rUrTuARYjmptBzzJGd9ZIzgY5g2vNqJKwQKCgbSdBR
/6hY4iKOIQ8tonZy4ln373cxtlpxWQmamoWJQbNX1EU7AgofcKRMVmCJpOysmnUeEFqBZ9Kj25b5
eDVBtUX/mWoexQc2dSl+sRteCXuwdsiwfigyCd5S0XjPF0Ui/dq/Bpjt01VPc59Lz79vb24/gNrl
QhTwe69wItu+6gmtsU/UBrFWwjPkLOU9lqY1dS3vTxf86J6XVuFMnrr8sWdoy2HrLgYIamG1C66z
22l4S/fsHAIoVEBTSTcYaIot/4eUoagleed6eKM3k7vt5nhH+GNT7qLm/BkdFfsbkchpgesbtZ5h
1v8wI60yPiTLPpei24HkrJIVeWq3BaG/vCSprMe1K5teoCmDl/C00sVimxImK2amC+RjQsEAAmRZ
SsWq7QHazjz5+2VQysanSDACqLE8IE78kxNcSmKYGmbeBJSABbTReq8DOiyOd5srNNLRRYuZZPPU
/jTUzM1zV/F5T6/ZXXLQMjQMJ75Sb7jSePRzsMfdolZqEta2j5ZUsnV0c+PUswZgeU8olehCBieK
h219UirP7zDHUZPaenNwahY1FqNbhtkxETDUGj251tbXxFNeqgBjTOR/wgvli/iJ53IH+by7FU/n
HbLT3NmMhvbmhi4o9ebOOKg/XzNGqWlSTk5bn3bmoIiHUV8rErshzqLkCZ0zz4WYe3HmtgYDNcOX
rhhi3AfqlFDZbljD5d1zI6nqvMgoQ81bWrpC8MFphH56jzWDHJrUcK2xiwfQts7Wa1aNufOGmHay
29B2j8vReDARBNFJ6BBq7mO1v3fcR1Qt54RNjDaBSwsNJpBwDu13dcAUT8VZw88J6GMv5ulEyebV
yxJj7jw9lCkiS/nO+hTAJjraCR339iwK3yLu4Zv4nOIBwaNn1lMkHZ3BQblCpm9XokCWeX0DWa54
3a+6u6xTDi2g7vwYsP6oB3F3VQzTvUIB76zw1SK8qo5IHpt3ONdz7v+EeCbJVaonXko+ErVBQfx3
ELbbwTdlzjt1Nl9mvFLfjSMemO+/oI35od2JsVVcdJBqa7ES6DUAP/TvYNancFlX+3llXDQJps3a
HYUkcIemJ3KFQqeZLEvUMqrDI7N8WoPONgqtQKLejOsvCnMB56APq+XrCoJZGFmd+F0DH3Lw/mk1
pAe6Zfw0iRdn7KxdJqKJyRMzvH87TLlu4d7eluNmyBrcWJpFG4tqM2sDIk6x4oATC7aYFIdGjwAY
B5dHafQZQiG47gzAHrP/fxvvzlGrvEk/zRqxKicdMr5E7yKdRNCRd3sljg6rMlCM339N6wjvOQGd
5796ZNX08z8eGEuyLfliibbZgTv5TpxBHyfWf1lHYZsHTnud1pSRNYo2MaUfnMpAujqlPNOUCW78
0WhnsfC5Ud1i+D492WC/nE+GIFvOrVBJ1ulVbNmn6Iw7+1E/9NyT+kqqFvmOjs50vu79WeXhV1X4
tMa7Rmhhy1ev2sTQMYvXX5UKUmq1CF81PzE/pRdSSOM5HK8L2VLVeDcTifMZSgJ6h2zRuweBIvhH
McxsIbMUfCOTP0Zt0j1hxmBqDekB/GbKUsBMUCmMkhX6TWIB0nBAxIrE0s7ExNAo48juyjTFnQfe
xD7tc9V+cDBIZrBq2n1/SluAKnQE8ZqkCtgZmBtYu0VnSLCNc2lTAjl5Zg5Oyn5tDYd1VNUUU6/z
Pt5dQdGNitWRnxWJyRrh691fwetUSNG/CCFVxMvztbCAc89wJbdtzb3KBhPrZwayMpnpF6eWmxCr
21k0CxnjdPF2G/Pte2ZK/++iMrnCUZM5Tx21k7LWOGrrBzxWurr7ZpeEvQs1WL4N9loXMkWVQ1cs
qn+GWwqcknYnnD9t26ZNlpd2MR5O2miXpQGeTPRSveRDLVhGV3Jp1r21/9dmSRSiJ48kPTGSAspj
v2w3qeolfFz6ccb/sNXTAkHkC0n+CrUMJiKEbUEWWVB1YkZS6E6OTGMOxYPWmROAZ282e3R0Cl6Y
r+xVyMvbJkqE1AbfEIaOTUrKANUVFWd0zrjdaeYWz7CEJrVvoDpy0ri++LGvo4E6Is16O/ifTAeq
LxD/mK40ZqbxiPI7J+Tc9rKi/1GZG6N2AiYgHQHL0xY3H8FM2avXKOY+ALlynUxb+m3Hr/zUG3Ia
mQM0AH8glr7M1Gx3BQgpLXANwwcoJ+2SOUe9IGf3EhEoEd+RUnSxkeCx23IW4t8AIkMxE4ao2akG
Puf9ZK4kSqBa9O/ewV8iXCqL2bscijLslqq0TNLyXpXJFsbZWv01yZknLJMOdNP4EfF4CQnP6PyE
pDsgukJMuiP8Ono+/GqDHohjO23C9uB2HUowXv6R+BNxv7DakJc4887s7VSwCX113QfjPLx6mq+m
llaDAqJQXcKorraMo+3DDrhqSzzBSOYaoH2WZ100MfphODBJcuKRj+sD/bWMVd2n3ei69LWXI7YI
o1qLZpqzCBlOv+g90sbiEfJaPuPjB+0mcsv6Z2hZnhWDawSdmifodd3IZ28s51FhxxzcF9sDdi+e
3c0E1/RKxxz+aivVpeQFISMGOO0t7yfWB4tIqWGh+P2qBoa7LtkUO09vXRJyPUu5ZASzAK5maM/g
Xkab+sgcqk1nLOCxREYM4IEGG5olAORzRPHIHWKKb3BZ9m5GYeuK/PVvi8wuKAmT11KhQfcHfEww
qa9K4UnjSYJbDbhPuOruz51JQSl8u9iQFQvpu6FKqY3W2BvQ1dopBSWn6u0LdNEz9jd5olx4lGtU
Lmmn9Rj0ux7fsRmzKCA7ALFMgy+vY81LicCYAqbKaICT5fmP+JSLRrhaFCCOny0fz60YuPDS0XZS
xrfS3qpkhoXBoxWwWEyCDiN9Lf2eMk5JosDMntObNz4C94esz+B58t1C2nsLW9vZ8jS1AtEXkwda
vOg+HXTErbNK1k111x2Q6MwvhzkKmQlxIAeSJDsy3AxUwn1iO3F0iTWFFojiOfuWBl9AIUr8vByX
gRUP8De72GeCeaUbuMqYQCdiVTyDiyEda4PCUtrYJcuMdlS1zHMPRRBPd8nxlovylDNH1DaGuK1u
SBM8VNwveg0NSFM/vGCUuZeAWf1bMStw8hXxQVfQK2jKGGe340Ee6+fvFKnHZGoIBDwz1i7wlfST
IJJEemlsR0hai7kc24Qd+swP0Gjix7fCENiHCaVknxBozQoCc2NeMtJnALN87cdlq+JGj4ir6PT+
MU3+OY+oVR7DerKH6gKfpuPiHjWYEfuURYMLCYt6brmuCOqJmcxMa0PkWjkZlcHL5/vMIKCwjXxt
4tewtwg0gBfR+5xVgJBSVnb7B3ZLBUrK8XzdhaT4cBAaUoeIbgTRgxQoHPIyepehOkS4N+BT+Umb
+JI1KZXAc+PBjKb1HtvEMfNujGloQ9J8xtY6a7QQNk3HCt2hvIDwFrledmVvSxJY8HIfZ/J2O4SD
8/hragA4bHoN78EW6oxS2DS+FAN3Sto60e8r68P410PEIUpi7SjBrIfVaworRs8VtHlx/87VkjFd
oG695WfIqXi5CfUaAhC1zWvPBMbrTygziBjYPBmEuO7RWRdzDh/NyqwbxNiWT0FbbTWY67W7/Pze
qoZr6b+kVPF8beaPt1//B6NGec9iN9b1Tew4rKEJZoTYUQu5SeJ34WD551uE/oiiFYS1mkj4Z2uC
C0RQv5Xk4luXOVWtqWRw4oGmy/sc6skaxzFdaicU0jVYyGIbYyB4F6xSX3Ro/p7IGy2Cre4Az5FB
kKMyaTnHW3wuV5Kb92Bb2gq2Stj2XndYK1Vc1m5GgrJTKVC/R/DFSeG7ucvG7hqQiqGR9KJTo+dh
Plj5FCjdiIszItzgBOZz9kAuxRzBA+7L3ScuI6+Sn4tZCviUbrShKMm6axsqOyDsjFdW55KelB5i
cTnT28OWG77bj9fFIGitgjuREieuFCgG8lVE/Eh057Plsb9cRGHHqKU75Ve4ZlxV7S5X/A2TJDpl
A0IFyvjooJc0jo9tZLng/hfJ7fQX0EQRUmyPArsr9HvdMOfgDDTlZzydCf7jpFicI8GX9dIv9ptX
WvTzUiMzvVaq4NR0EJH8hHlEdQJolrGBBxbyAm3SfkCzo4ene3cHJ4MvXF/8Cv9g7Io0e+Ppkvud
wXIfn/u6s0LtGBY3y1iP/uczzUC0VTdN71Bml1m9utpggiNd3MuJqrTuuC2dod3IdYejY63Jpc6T
MLRx+Aezobur34Bu5kxANBRgUDy6C2ieGNHZnpvkKlpLG+LOm1Q78H/rx8avlfFXBYjGK0wIgApQ
I2kFrgEs8djRM9/hHdPwMVFY408GYenCKg0Ox9ScuhW1DYtpT5M7yqpnDQSBNhgnLVHp/YyJOQSW
XA4/ITD63c0GkV27N3et+zCxjtWBrWmxWQAH0Ad5Yau5pgWLlv6I6aeHhvORZOmn/1PFd1ph+8UZ
k1Pm5EbNXEKrcXXRNsKrGBRK/Ee+035528uT2AcgeH5pAigKiKuhaKs+NW+s6tH8ZKVZMI4yV+cz
zLDAwJgrwRCj1BHWyXp/OK9zTSDnLi1sUFNnL1GKU0sdgmgXXG7f20A51/wNzgPDcoySwIL/3kON
Mk0fQ6Mz7l+U+vCManiHMtmZq6EooERf0h3ZaIYCVQRF781rM0QQ1um2+HIiAp/B4x1FwajvydAp
O3w2pZ2FK7C37/gx+xIrIWtqQS0Zk2Ch2fi/efzWH8+hIDqiF5oa4aIsak9n1mz2l9z/RIGfGIn1
vDucGYUOe2rhaT2iGXT4uakxA7bRG8AsrEw+p24likcSfX3ym2xv8pK41Ng+i3X/VhdA1bOekN3d
0X2nXNoUYP3P/qqCFndu5zkE5mwX5xsnhW5b39JhryGVH/dKiYIM6uz0f/3N3XfffcHJkUu6azsz
gNUEpvHoxygYkvso9aKFhbO1ll3gHlYaFWSLPGH0H95/NSG8ZB0503yI34ns/J7JwJ18W+V509LW
RarTkZEzDIfqPG6ZgLlVemoHHVO2D8+qS+riR+f5Va2o8b2EsTCySTMGg/TMKirMi3nwk/0sqBjW
RIZMleG+7xm/iBBt91+qaBaXJ4FbHShj3SvhRHmqX1vMnqfd3MloT+GFFe0kZlncatzeUbkgFwis
zzqKclXPSI+Oz2LIaw7YrALGRi9X+ooVp1hHYwdFFzMGjq+h9kDGwGz+WeHeBEaN/2sngWfO90qH
7+NvGQYUe/vo4814TCC0xDegw36UsEg++N2wx0Sc3ZOoQ4S5Xt0NDdtKbT5XAX/VRmCIbgmEK/N7
5GglN8rd2mlqXyGBvF/fk5kPk1Oeyf79XACGBomJL2vyE1CvJ3BEPWKtAm58q7ZdyYtiiaMQ/MRh
TcA681UuNTpWiXRte+vNZY9xWuk7LcLmrWTaxh1ig/OOhuzJ8bXfB5jin33Mk/EqonogtQDlURM8
lERyFFQ8QoAKU4pE88IggIcjgMCENd5dd9pvpT2Ciml8Lac80Y5PvNmsYN6fzLrTcNwWnZeGDZ0U
7WVG+SKXB7tL8oMFKnfuxt3BAUxHurTbawEipXEhBaNpFW6ELuMWjFlEe9SgkfxEtBJMzB/JmgkL
i3GqIgxVdwFrkhRKJZn3arIXb51/uvzF1i+75aqRn1r/T7QyTiPQBVBw65uPRG0leH7jKO+E0+hl
rUexTrbZpKNGmT6Kxu7+C8pE/EHLvhQl6tF6KXwWnjYtbQnEFY5M6caBWKnrRcfAv/bR1HUTyRhD
TMffZ/9fS2f1P9FZjT5Sj3M8KKITKzSBDL7Ius4TzCDWA/F9EuaG+8ZSQrpeaXOsJt6wK5uJU+Dp
IvXPaCqub0VMknqOW8lhziEouVFses05sOeWuybNcYtdUv3KABqjRRB3of4TRXvMdObYnxOxiL/a
I/ohL2D2U0iuAFZPYc2006Dh6MV04Y+Ppz3MK75uYOKmrlwZUGltJOOa9liW9xw7PXLx9gsKjOsu
mgiLc189ScBDXgEZbn6HTKVHniaDlbjMDjfulri3DuPSta2U6BpDg2D8xSwPlCwyUJdIIzxJwb8s
ctng4L1BcjM8KddmUp8/Wj5jUqDN1IenUIqka5+o3ERwxDg8K/lymmlqVYK6EKzV3sjKFfN4BSK1
686+CQRPGbp8WTstBJUwY+7Wbx2sI5S3rDyA0NoISFVTeVOHPt5iwx1WngFbWi6bonOhg/lsFGXB
+kZaMeXDaV4JQpZ6YnzfhaulLEKR/DAAF3Gq78guOp/UqS+31vBJ0LZztgzolgCtv2xpF8+8qrKQ
aWENYx/uxTRv1Mwe3Q8RKJta/1T3jdvE6cO5EWZT8l/qN+QsyUwSkDzGhHzqCp/HjIeIbEnB0DQc
5Zl9HauDwLCy40zPf3S+ye8Sd86PA+XWJ3CHylXK8TOMPR2sBMlWR9g1hONlkBQd7f0hfLVujL0D
CPjh4x4YLr3Q7uW2/cUXv0pAtAQASBGdCBSoy2ZFi8lCxmPLO58A5mXCrNDzh0Cj0HszoHwiuhPy
zTNx1YnMcxlHLkQlcLDji4vCOfxsn50lBsgGNXZG0A17i4HyiI7FMesK4CB4V1btshUB8T9qbpmB
49ufFKzQp+TeYTayGUOmOJ7ZCHi4CSeHMV9Vz86HwmXVT2HsYuErQrV55gw57GouNKfPUGDHDAPW
6ojhhXa9zOUXeQ7qygrmzddb+lNRg/bH2ekExLx8U0nb7mCTJHbGLJpTo2+6/8bXim2Q/Pe0Vxxq
fLr8+t9RfFmSVF6VkVMsGYc0gvc6A7+O9fZiUZs/I+sQ7hyC+Oz9cq74ncQ+KzXYQmbDvx5JTnzr
Hhk2PwV7xYtN4lQkrUk7HTpY0curAZ5IG2zfgkleJHHGWU+fDiZT/TJSEscDzGenX0ip4q9JYT7r
1ACmqsXHET6gZ1pxT97L7Gf77uKiNRFpxCQetmykAvTS/VkRYpPH9ix0MGOkY6Zi+8zLrDiSJ2Mo
qC2BRA4fX+qHqyhrMQg67sOU81/l4/g6xxMDOB6WLBJUr9X4jFZ+jLroIB7cK+9/D0whKTPQfgjp
JbjXcCYEqWloxnaJotWbQM7soot3KqW0ibFwvw4ptLzgOOcFhW2vYK+97oB5O5taSsPtkmqyEUca
+OkjJpQNw1CwBS3uf6lx3Ar/gtLQQhbs1K0hdgjL9JSTSXj7BO5w9TPGbmMjxgirevV7NoZ+6jka
BUCR20+xCZM+NznQtnvMpnzkMU38Sh1dGgioIjXdPkaX1FJAYpFdnTw9C82qdrYw7ii0xZSHtXvj
kdazxUgF8/UlZdcHqXOykHE0uhwkIkXIyrQVl+Gpa9j7MciGB9fSRZ2v2v10QQxh/w+IqORHmVvi
eqeFFFr460j4UGX+gbf8Ir//OjsnWCHfDRdBWa5kbMF5ll4HGH71/R7jBf38muUcj46B6ITIESda
lZM3OtwOa217Vl4A7oj7gENaaZ8BgnxcT8PAa45mUrXoQMJ21sagzXwPP13zAx9gq1uW/DSkId47
iJlll0ffAnmhpX4xXi3sFV3Q7x05pGu8WEeXjrdCIXHsplmGdQSBG8N/Qsei7tulxVVEdXUFdNYL
Ujxq+VhM46U1CySoUCi+cgJfCML3b2g0Eoz2WqCS29QOmNAgOacND3hl/VaGOQMqosO0uOpKu79c
1pMqZGCZ0L+e5HOUmJzTeI1mePgiXkqO8d3ATV5fCrMt5sf3CQLq81ikYWEZx76gdJFZmPxgUEmS
KjXWiwCDwlYY2hbEzQ0GuXepbCn8cM8985IRzC6XEyM5MHB+EMmH+bYwdnBDRptI+1y1eLiXDVac
OuG3hcfeMnthJg1FyvRww/O5WARxuqpG9RjWGDANaykRhZ7Jx8gE80IIFE9THnfxkLsX7Cm1rC2h
LP20KYyMdOiLPxJ918rIfkvQ8Gmsv7qHHN38n0y3DsuhAwB3KW5OhISkpxFuDSNWYbmhsnJKOhG1
Z7yMJ9CW/idRfgSdW9KROAgFLfqFl26oabJwupYzBfSqOI3IE7vAefww9cQaXSRcSeynxWphke2s
ZNXCxvFrcpW4HW11FkuE81+1Lxo9LzULZK17gfzw7GdS4vVJ3uSWydd8ZtQHbL6N7Y0gTjrjoia5
6zvr+2aHOnh8TFKKgUzaOMyrvTyDnbyQaD0yc6ptqFIRnk4vdbDlXrY73XL/Nn6AoeFlGiR66BW+
RJGd3K3iJwYC8Npm4f84uMp5dETVRPKgI+H+0tMpBM51dzwhyCCZjwl30B3rP6SHsuYxyFPp8Qay
bZaJFKw7LzApsF3wCjvy+mxPgHMNDVia3Ji46tQP0tuzRJVN0wwGQcQprxvFoOj0aAvKT1iR0AdH
0X768JIAhs+O/a2A435y3Lcztf5BZbWBDQylKPQ0L1UOXr5YmKWdx4naMV3fzfG+bwgCAytPDX8M
peqtleGEPIWXCtvw3AVcgaq6f8aHYuFBN8pkSf0IQ7cbtnDA6gSKTKMAE7PfH61IzjYPIGlb2YpA
2vHxlRD0iFOP9pYSOCFR1/MVUGx/Zfs1NdjLW6WTX31yP1NiNHxZYs3axBh1szneaH8MzxyrOYbo
5V4SygAXdlAmhpEELHu+j5rLsLHZ7eo3rCGq4fQHmgn26hBIKR2i+K/Gx4jo/tEZ2dHSpbtwts6W
rN5M/hfVXj1fFIPFEGHPP6TmGZ4ajoAAwUk2ExOAnoljYoETBRQI8zeVmJDNKwjJAmbIxMp/rKmP
Lw1viOH3madpylCNhOS2bBQh3qy9BMGeXIlR2gWmlbM2DEW7MqNHmh5w4yz4sf30qiOzZ4Us+h+o
UYxqcR9wfZ6IzMnMr9F3Q+Z7H9kCYjYFD91VVNq26oUz7Q6Ts0Se0DGZHOjUTHmur4SXVIss4heh
vszV5RCqBh122XptwscAZ32VB1PH9y12IvmotyryX5RhPvgBYbkGY0lL1Icq81gGjtI34Eq4UKLk
ciTE90nvR4P3LXGFuMkYBqEy7lj772Ksf+2jvoJPlVzI7pJVpilQmE5Rrcj6+UuG84rWvTB2U1/2
BK8Yp5WI8rWnkNjZh3OvQi2BXH0i1IqJLceUeZy5p/heudMRqpl6s1m/sAtX8wG4PlWUrvVH044B
VaWv5taVVZRYjSM3dKVZ23yaK1XMEz3ULEogbhdccohyOeUy2CH1MZ6MCe/Opi9BMfklrUB8jRfk
L9xyXRUIvdNboCbzWMytZSeFLaoujiOZ8Xp6k/Q11TeE2pZTc47uXwdmyxsZtq2bK89U3U2wBWBd
SC8nhWWy17idSzz1FGloyCscaM90FOuonwgxx+xSq+T0YeMtoY6hTyFKhzqo9EkL2DaJ2y9eAvk1
99Vfjc7VXCN0bvEN90cAimv/ELlkx679aOZmW7AClo9xdAQZr9YJBksUauPrDgaOI6/mB1qsnX70
Kc6hbsVBX+PFKMvgWSX/M/TBSEDObV2rP/2EP6CqxmKjHXr2G6XBXBbCZgSP3N1SyKdRiBPUXSEO
5q2ypTWuq+tC0JQHbHHteP5yWFXPLhThT55kWjDgj0RMKidcJ87lTjcbBCegv8CcxIE75Dk46zmM
bzUserJJlommRjSLRiBEo/4Du2Ce7uqiJAX/Zo0RdOiJUTFm/g/V8M5c61Wf7SlYFkukyo0ca2PL
3iIw35/I3qdp3hlN3yLaRjbkncsUhDDeHiya7V8bAtk1CfZdLJdVezujDkfK0PdVhmeYyxtUiuUS
wnrL1QYFHZQ0jDDi2Ttb3xh1BWLGm5PU3g5/yd6Pre2Q2JKAJ+G+ZyWB3Lzkzk/R6yiuBi0zNIkN
dhYsr/qZdySSo+Hv41r+qs5qhr3HLXGf6muQNQx9lbciaygmcl6K4dRgPX+48dvORhFWoInFi0gF
TW5rQqZT22ChccmUs5KeIKbg/Wh3G7aS3IGIZ/fH+gI/ATSAczFNEB7t1Z9as8Ai7YJEdMtdiE0Q
/nLL1n8K8VhQ3wWbzqEJh7tdJAWcoA5DA92/DJhCTva4XyPg0nb0L+0yiwfZy/FWgWeDTfgVtreh
WzLjE2Qq3C4nz+qfw06d5MmS7OQUYHkbJNTjiJq6hZbS9nvmcL2o8t+9x9qhe01EG3fOaaHMzWSq
NulsqBGHQxfmA7BuVLIsefwI05D4JOEeV7Fvanrn5oWO/Eoox5wWQ4z7A/8Y/PxWydnbauBJpp7l
PRDa+YtD1aKcP7VQbbFE507b6ZP+cKOR3SP0w0S5sy6lQ3dXyT9Y8dYAlqgZ1Pc7XiSPKSjqdhjn
KdaqezRpE1CkdtfOALRAIMeRL/LTIMKDnySDWlVBma9Z2ow/0dh/XRbc1gVGFA25Y8xpqsZQrvy0
NUiOMgj3HZvrc/N73eQ69qiJwNE0+V7ACtcCaXQprFyev2x5XRX8PRBCWnB352Ev00y2GyN2uBdY
k+mBdHJeetIvUHoA/mvZk4uoaliT2x8eRRLgt7MWCn5TQ1P1r6zd4sA6VNkFQedeVdO2DpkXaIV0
97OtOTWys6cDZ+EIHW6PolkskD4pYZOfzJaDPpX5pa5mxd2tOKagJUjZYzGaXto6oHQX9JP57FU0
xVh9rrC55pSoqFk5r4DAxGwu356agie6c047QEN+OF+h+f5vieXs8dJnYMWWQWtehjsK8jqJ+Qmc
tztMeiJtbiwSjrw1NkLoTUAVnE+xmjl0dQHzK8vYUS7m0X3a4kc4uQypZ0O7/JE9vQ9EJluWDJJo
aXC8f8o8ZaDZbezqwIHrh8NN79c02c43wiixx88cCB9uq91913IWeMp5dEnHSOvOTkmhCCuBn/WP
hTQYLhJh6+mr6ZU8C/yqC/y7l6nWxY/hG1RP482LcQP2rscTT1M56OASP6UNroXNURG6IDd7cT+4
Ei7CBsEltz+q2SQv5ZsivUfa2vo15MNt8hk9YmH1Bpu78VJu87oSOljRugh74tsjOOeKpeu65PxK
TE6FET25miITGEiAM0EdTUxMI+/fJx/Bx3AGG5cMpqf3C97wn7a//jDSy6TjtVF0EMUAuby/ZcOG
Hi6FJ4/dbPhDID3opSDV7MndbYzRZvDupzTQ/ld9IDOAlnvIBr6uv2v4WUgoTMpFPkT6+zGhd/p8
kOGLplOGMFL8PrZT/PFnuEjqq9AgsgUryksZWoy0Jo/p9wP2nHFcqOF+PHvZDPTNt9xe+8rROejj
uzqJn2Y9AnDy1p6QNdWH3PQkV4NQ/Yrx3bPcaUOVM48HGHZDdmR3Yf2M2tWxPcbHBJfgz08m+xeZ
QySpj8h1kHXuDKstaP59SGaYrf8doqz5EuRyiGiqoNLnzQgXQtontj+vj63suNYwKesWafvdpewV
uzDb4WPxfBWhrU8rjXydlELXnbhjKZ3UVDjkBf12Su1Tf/Qytlgv+9UFXciNynbhBc9gyqu1TJbB
xQd0WnvUT2PIIlxqLByzngI639Z28lIrdkGhVzcSGoIRVHjSyAhZEseoPf+41rl3KlSPptSlHmXj
aAL7FTrzXgh5nOY+R90sQ6/M6kDvslIBdWxHiX5OslnTX1rjdtZQysUikl9d9GwMJbp6hfAdODcn
5K4pts4SwsmdxAw1+cra4vT7IkMRkeGZHH97P1f+O6xqYHDq9rkf9oGA6WUSIlcnqU1fXmFguEA1
cfPiRZNiOEjnFF1TiU5T5eqvzkNnunvMJjAj7RWgVCYCFf37XhnoTU5+xx9oiz+pmdsGu76Hn18v
/ccowW4M6Vv1W62ov0H2gaVf2v2w3H2tC1+kf81Ebfyb8N7RR5kQoQ1cG0sgURLGhx3NVpuJH8mq
oGtjN+Polp9W/wsynIB6y2cn7LGGgN9Jb7Xv4a+soI/v8wT4/1BXniZZ3BHSJdZSsMgc+bu1rDIO
h39/GaskRH8mP7UDugEG133J55X+o7z5Q4a7e9bFsXdijoG4bXk79aft2UrTvJjcnxtBqOkhdLWr
JDnHUBHrHiv8RavT2VPEWjetRRvHEvgWLGieHQUWaPTsqDiSL6vodLGx3hdxk0IiwFhyQcvAmm6q
yx7bugJnHjDtcHUJ7Ux6+JGctSP5bDDWi6Kd4iakQWs+Xb9UZ88hw6qX2y4mLwSXVqFLx5T/AUcF
Pd7AhkHVHArXn5REknidpxEqYzi9QGFqrXJyfceAP9GJVohG1DTsVmGSy3pP5kKS17ArIpsgbAwW
JkUNGpqb9HBMeG7Dtoee+6yo+DIMwy318VST/N99Ku1S4ReXd2APtnOwYFc2JFF37Gn9Db+ivxfg
UBVMR+zXqvCNRe6Rkbo9GGZJQT6ttGKVFaHWa61KOc8qPKwUKPvQaw9hfBjYYXmzzi9mkvVn4798
cVtIOpIIvLeMPfYLCqdDttB1ssYF7cb1sLj8YY/GEXweEhX9MXLvz70BfEx6LJdWnsAMM7HcvzzY
6D4Axxb1hTFZRESkdZSiK71kqv+vMBqYeRAetQvkkXqTepkKV9DO0tMtuYseNOiNQBWDXbKfqgA6
pCK4CHWDfnxlidzPDnFZse7i96rnHozSiJlAVB8uonzxhjIUHA8V7XKM8WTwi3whXLe1jBfpTRrd
9j9VlUtmKsmvLHFwN7SRdLky66CI14zYv5M/Xd/yTHSXlULNqim1l4+7v3dR/vZir9JWSQXl5ppO
EHxrg1jd6gIiEhiUkxefV3wF2as0d23aQDQoJSmruHTQjvdFVqDBNYN/BcUnYujtmacEtZS9eEad
vNCvLo00IkJEVhRrm5kE4o+0/F6Ud3FAMNTW4z39Qjki8B6ORSSILI1f5OmLDKpcjMDhoPx6N5XI
iHHl3cM3lkeJLz5FcvVOQSiRbTK2f6+q0+Enl9bJGAajzVZMb8KLGqAh7F7BsjAnf69IJFxi1bA5
ZfPejK8vMz2O6BbBetyA/WydzPJOYDsWa9+0jzqD//Nxs0aW1MqDeBx8/nVFZD6GE2L0068brRHJ
oRyBEWKocmTAGu3DieR7xjIYBsBFOKm/oyALk4b2a7ecArLaOIwOtCmzsr3CAbL065rPC9Jz2Xl4
BuTvY0SfS0NR1WD94XCDt7b8c6Xe018EZ1d5/VrnQgcx/yrz3Nas2rccQh0Cl8zj1RX5PWbk9jzC
YW4MWCj6QWzW9H9FZFvkgr7ClgXagd36boF2f+RgiqobBmqqJU2WjwjltvcpVCeVHmI/6OyKn+5M
vj6nWxsiwJvhrQd+YjunP/M96gkETlS7wFkXjQtJ3N5wB8dSdVy+ADhE3nkQP0iYP+tNIuKPdzp5
72YuEsNac86Vh+6Vkz5CPqeX7vdQmHxeCBTn4okRw8hfJiCIe9cTYg2Zi/FQFdALgYz5f/iWO8qL
JoGY7mz41J455tyqXvtcR9EoBAl8rXzJCRxO5oC4B++hOOOYoV5rzmfW/SiACTwuGWAyY/KhLDu4
FtFVughEvOidKsUy7g4VZm897mteqHzJwCKh4YL2IfFmtqeRktgwgJGkBvw6OAClR9Y2HhKS9goU
yoFCpd0/ChZAKJcqsxwoTuI54Bltm+beLlUvIg55Xu7BVNTKECflh68769CgCTNpfpTrZfE+jseE
TqPRfjQP0k5pQ/xhorPWgkaLUbmK76pWTk6B/2coz+Cdg/0BBa2naylDxho9SLfUPYPGulHG30HP
n05zpYYVPTP5YI8cXV+X+Qy+JG3Uy9NpOFiINq7mWdtiBSdlt4Nix4Hkx8IIPTxLcX7umtOLf6r5
q9dM74h0tpjPtM0cVW8UBA5VGghFdIocCn1RLWhrajhVtgL3fZeG/X2vn9Owc7kjpMLEjJj8OOAj
25Oq8DKWk3/K7rCLsFW+5/k2m8xAw6OEXobFHNCqIar8Qe02HBBSzmgsUmX4+bEaBwVKb1OMz/CT
KUSrv+wjI8hiIPDWPKVaOl6SU5qmzLdm1RB0vJ7nMBMWi+iE7qKovRscav/Y6WqaB5EvINcxLy8O
JXUbqE1T50mdNaeVAgqMgzWuD84xFRNpUkz1Sncu/m59k6JIx/Fin+cQ63x+FG4YC3yxCoh6aVds
w2h4IjH4zHlSPuXRPFztFaDlb9ZbPaCnppJiF7tkQ9A11vNt0/7QMDrS4ZCZvaBsg3MAuh5YwEyV
083lGHVi/eNTlrsNxeOWdxcOBGWdISzENI5RVwNOwSMsUcfNh4sirqkzinmOiQNu8xE9aCfP3DoW
Z3VkSn081htSlo6t+1RZ4hCB9eNXIHxDUNNKZRrwjzHno7PhxOcf7oNvHVq/iz/WFAiK+tHeeMp1
rP9VcBgIQsjnmxlUC6yip6rDGxP3bvjDtlZerRCOn4vv+kdDcytB1FmsC2nq6QRxoUAmGMCOvh3C
eN5cmXTzPu5rmQeho33gJrkjAfIUvqgvfKKyKpb+6ebG97KVMjV5JhSk1S8sEsw1jGM4EXh9yq4P
tOgL2wrcYaOqEzYZKJ36OgGeVI7xSvNCKRtc8aZ69YyUHyI8sp/oMSq5uU2ixcQomb5WabQzMrst
KVIyGlrE6RXJZJA2o8/Rld2Ztg8/gUgAx5PIGwATjHl30H6bT/EeckNx/0ENRNxftIMGv0OGvBfA
lS/Oet1Q5/e7tVFaPospF3w+7JjctUCM+w1jVgvRr3IkNoCB7UoZNhruLYWcAdnApbkn06B1efUj
66pNR5xl8Zf8RMR+ITFsJJfUxu9V2DIckOU7PjgFBtWmX2/3Tskmd+L0Jptyt2PJjoj7EoOdvIgJ
igYGFjXniWQRxVF1ehYnMAocmCnsMLZPwAhIOjx0KvZsazRyoJjlTFmKX9jf6gqXy+Gsw7plffDx
SGyOkiNMsF+IG/lKdELW65Fudc2Tezo6mUeyTP8EC704x16+2aU4pX+BJWYS9WUpsHQ2Fsyr0Z+0
JdGQN4ekxjJbW/oYbB0Kg4vUES//KojBpUszhHLY7Nn1BwrmNGkrzWQ8F7mH6YYij6flxwytFytM
GEZgiFVZ2tZ+6zcSXT9SgwsYo34kK1DZgX8ytHF7cWlR1mM+PaqBL9sFXkZMZKKwWxFdIM0uG7HS
9cV0GJ8GB0Ujpn+rPHdWcphvOJzaPo9kq1MoB2tQqaE27NDTwznICrajFc3G+pXy2suQmWxvK5G7
pKc2RJ99IEISz3KLFYlaO75Qyzrtf56o25zBvwp157NsyaVpqe4ycxcn0uJi13HR3TTbMsVvOVR/
VvvQl+rHsln81L0kahKix0H1g+ZCutCLBzisXeB4hCCQZlam1SzkqNDx66A4tK0WGPMf5akfT/Mc
X4zR/YA1FYpd4So4p5T65vEuZf1CW2jOzEsiOFOEop3rRLaOjs6ndfcPje79l4f2geJDhi1imzIM
vDgJ9/cjY4X/NS5lVQT6JbiaDHMWSr1RkM5MrXFAQOvKIYGBSI1wPdwJR7jtd0JRL3A2gAwMfdtb
Gt0LQpx7Mg3u8xZXSXhQWYYeDYfvJEAEe6M+SJcr2zBrRXMmgHw5C2zChXBop951zKSR9/HyCp1+
cUeBf0wScCSDWqYBg2wrUbTRZJgu7JJMN27tvAr76lkoilat0NgP66VEhgPnXQHCa1DZ8wu3i2eN
8ttQwJ6b4RbePsrnqlOLYtrL1IDkXiPs1QLhq91yF3RDIrf2o4pMh8rPm7gXiFzn4V7i1d4SyeR0
bUy3/D+KURbTxqYPTxvMomdQ10DVSJoFutgtxzma6m5QLFQFOWpzrdXglNe8o0EB+CxjWw5bW+dM
VYmTV0NN4jiMhuYZjnArhwlLmvyXzLcfZa/b2Ioq9FUtO8lO12wQp4I95eM57kSwH0oFFuGetutj
Gjp6+mCfcE7Dqsfkb+PFeAvTXTVEquEkz8FRE5VPf9wZgTTDwr4s8jfZC1YjTjc+HEvwO/KlxIb5
ns/BPK/GVhXpMrTxcoYCCqlJfp1GnCo5zgWOz+lOthmK6kfc7kW9iEN/e7QN5dMfoVRws/CeslND
NtIXBMUFI4hff3WNOiAtLf8LnrYQkB4IgFiQT1g3F/ujCEGX8GcSuZObP3iWxtpO5r+mvFK/MFU2
Tyv13uzRaTlLnGTM5aRSaCZxZMbroD7j1rjffIWXiUXKDcDK05EwBjXDHECJh9TdDAtJP1MDHYpv
4yzvhSwAidecWGEMkUzjZs3kkWs8+4GOAIbXgIzUFDZ8JyqMjEdroOqGRn41SdOQP0AdabLlt7DD
ovE9MpOAf3QOzTmU/ZM9PZh+Ez8obyfDKjG035Ys8IphwujTSYBG5t1tIcv4kDBXCqpwOti19WG4
juGRnGBzH8ZIta/I9KeMRvaTyt8JMJEBcuqauFsCvHt4wRqUgvp6Rc2sgNDQiVdIkw2I83FlKiEJ
xu5tpJgj++4N0nj5JrH2RTDwAqRImQJTHAZissy5XwoOiqPOFuXt4zoPrqBT16Kw4g3rAid/gAYC
fbaFKEUYHg3JJxHYUwNuPXnz0DOVUbFkQyN/9YB/9UTpzOKLxAZ1tGKQanSylzIJ8lqckktqAjQr
jsUuc87Hgc1/bfr5PV09NZvDcSWpOHjfnZLRJ/mBOy635cVVmA5VmiRVVgDkaAfJjRgEWRFrKuln
FvWY8pNvhlxaK9ZjlhUL89pVAHP70nXAfzLS36HyEXApB5acOnWPskCZf+8d0ycj8OoFKcyp3tzk
S2Dd4JI/sKcUzLoxX8eL8e4vBmeuG7Nh7oHLVKijPUI/pbMjkZTNU9wsJTKdK6DUlLXyfqg66Pn5
eSUgVPMMIkj/1h49GHKQzlEEbiHbMFAkWF3Ax5bYKcmMATU8mFW1s2097tEzFYF5oeINVbXgal2k
P8qAR7ewhqPQhX3fULx6C0e9OaeCAmj6W1zY7SctHS/FQluwaPo2t1p6BXgwRIiekWhuSavbeaWh
i0nF6Kqv3vSizPd/EgnQ6fNPWYXGV2J961TGPf/AnXdxJE4JBpj0kkQ2fv86GdoMi58W/Ny1UTWm
cMnhZwy0qcwg03jLLme5pOHiEXgCcFEmbEkOoic0ctIdxqvrHHOPdrMzkFaxHRaxIJPtTn/nKBtT
/9Hd8NPWCou2hcRCoYatXp4LR6NBP4EHSfirzBsNQ6vGci1dNYQWW1NWo5L9MNoQy7db6eZU5CiY
RaN08XIy9UIOU6WPWmYK8iIJ7ixWje7IT3aI7kPkxo3byEZ8DLX15D7IBPbmiuvbyj4tGTJHS3gu
kK/xO+9LAA4AHFytQtqZWtYc/bUFB6rddzLEy6RrNNjPsiH9C0zZOVbUPs/VpIvsWSo+tVuPdrqN
lUFyJ7N2gtYuXdUrxldb/6GWaXnhLPbqUWoCOizdemwp5uZ3RqtqaVM5k2rskDn09I/RF3mAalDh
9zwk+U0lFUkLmdNYVQxSuTwWAWUbaZG37gX2GmYDKWu1SRe815tApHQ/Kl1uN+vviwEVMRpo+2DH
M90Y5tvHdPazag+zixaXICRD1Fx271s+Fxjj0BlbOPfYtZPXLYwaqSY+3weKWDXOD1Ud/I2nuC8b
2nLhfizl0bZFwyRSu0FK8xeujGCJhdMJNTUOpeqfdCyy3uxNLCr6Ujt4DfYZZuvN7GT9Rh8GomPS
aH7vmztz1QfeeNnTy5LLsrawX8CvWx0KwZmRrSQ2w5w4HpxBL5nP+PAfj91g22Zhg8d5G4k863Af
QJBoe69ZAuZXi5HIosop+ac86xXkRlrxXD+G/NF71wxiZsh73ntIGGgESlPNiIpcoQEcFSSHfTpC
pPSohVj7TGLSpXCvTyh8rXkYYFjrypnkXLX2m1FxrTbEs89CR5YkqIVtMKV61EtkgBVOVH6DsQCO
sCm4IgCQhoFy4slibQbgh3fNBdmtBUbwn4Zpvb67yy99Snj2ZP1MVRpsEp0KrdeNlTmqB7f8mkdq
FVJzjBG2HGVtnA6yWTmgaSn6JqckmUFko4hClKZO5MliwaZ+1ULZZPEhSPHvAIxR4KuD5H9MOo+h
cRQhKNsvRUID8W7GLpqmDVElMdhdzplb5sRjKvYGTb/yXJR1EbaL9s8o5T+eejhYyEP5KltVMzEI
ZP22GK0VRCg7w4wK1xp5RO1N0TflGsnDJhHiGiNWIb7gsnktxYM+uwmmLcLq7WWaf59K52tYnU/w
Fb4fvq2j/bsyzNUlQ56MkHzQF6ZH2Zu+8lGwQmdSwklqZVD27qbv8wNeJiyRoMrYwX1XEb1AnS2G
lsBdeNxh5hArst5+tfZrqv8kSOlHNWHv3rx2dU7ghLo1pucxlSU6fKxMF5bZY0K5oJWECKfWc7W7
+Osp019DF4lG1p0Nk0rlul/a+eHGS+BWxGDUF30SREe92xUNJUQgw8cFFUMkNtYDW0UI58SyVq6R
9fc3LQXvLIdXyB6/9M+vjzIMUYJh8kcmF5GYORubBbeX+LVhaBrl/kfKNrj+ixr9/YyQLDlZCZao
mpzJlqKirkk725VMjAhiv0ymRsAIc3vAnwG8wIP6oPJlCaCl1YZ8KyUL6WOC8EzRRdRbOzqleFqt
xR/pjHl3Poz/ZH77ib/7oIUv8qpXpaP7Va8NhHeflPK/KevjQ2g+NVn7c5Nhn+VKxhAHLATvhtz+
i9Dhd7uwDLEqautmoIecU3dYZE0KySGE/X+jTS02MSEM7GsoNJi9+plmtWOtSI+31/XwO/KiSEfw
faGHyG8XQsq6rpNdU4+zNWSyw9dl4Ysi0ca3TdcGwy0+0lkhgz+8Qi+2JL6U59Zjm6M4ycDJfBwU
0YkYoRyvbQUIb5HNFkCuqZNriXn9Bn4PbbL/LLMYTOxSUyZHh6Qor2DNcGfiSLZhGGAhdPdYp89d
BD6UWyg+rzI/2f31LEYemtw8HuMROLNoQc9xTMnYaySxc5YCksECTdWv9iSnQEicw3VXQ6v6HiHP
m8g6XXy+3c2G7Bivi4UGTF36PsUUCzuZfmEXLCXqGfzjeQSiFnQ6pAIcJP5q+g/it32vL2FYFjqQ
4S9jGU9/6t10JFpN8dAk40nBIBZc8HLIxnyYr78MiViYBM1jDQBeUK7I0R4pe3D7o/yLrqpgGUeN
jtNXdIeYy5LIwupgC0bLifB2bKf7sKBPp5mbCvlgwmy41bI5DH81aqIeG1wrpiDeqiPxO2aPPS6o
G7fYGkWbwQ0r5a4Fp5FxqIUCosyp7bCfbnepuaziE38TgzzGWBKAyRLy4T3yIkXO91W+p6KtMx8B
qlA85RKfI0KjHlQoDJ6ItThOyBSu+kf9982DbvHD5eRalnlp5fANmgdVd/iaJHzhvNaNuiiAOsKn
sBYXME0MQZb4wLI/7K9NMDdpH62Hi0i88ZW2P19VWK51aaBBcPJUJLhg63swFxV5+OnSxUkWB1Vr
yJjueA/Srwem9rC4yp/ohuYxb5edk04j3hdE2rfESIEJPwSk0BzW5Nz/oL7JOmmhMCypZlUDTlWX
/Vsij9pLOC27P0scLxdWGhKFHlKvj+TqL8vmCZAnyO5UGHMxNviFhG2DEgjhqCi/qH5TzygC5iZC
1p94sqrtxBavU6GUQJtqvXBs1rME3QjVg/gXaLRAYsyjMP18gp2UTtFfiPSH3qvUx8fmIoPkl7Qw
51rrJ0xMVL/YcVPE31HstmQqTtj4KB6uNSb3Rh+GsBRMj5xj3WlhIMSznesgwbyiGmrFVRKOUteT
7HF4WOSVXmbDUuxC1R4mt0EQR/vkJALQYam/gUtjDdoBEdMGgyD5ebN2ow+vbp4oKZUAG5wk0xg3
vBG+Btymr8Pi8zELlW38i/EC9TqYez3+LAIJyXbrWsYvz4AGOpMdtjDMqUlrJJQowENSATKujJQ1
Ff8930YryXNHj089OiyUr49fXEqfgHtsieF6hrFQiUAWAOm1TF5OpwgN1RXdiw/XsrZm+6c0IEbc
MXC742JNZNMEh3Xlfg5aW89jMEAJntZ8I+j8LhaJDa4v0VxKQ3Zk+3k7gEsdelJT6orKiPI141KI
vpUI7meEiP7jc5OvghSw4IX92MvCVo/0VyvlfoVA7yW5PbdUjlsIn6ZWYmTDx/glJ23dWBsFCzew
jwqy7lpGePitrooxAB9lI+5wv7eTQY3QZl/kn/hHt9RE7JPuAxg7qMrIgYirgRay2TKYXN0LByGj
wpPTjHP6GTFiAouJUG4TF/fA22rspP9fbvzJIBb8SmtSML2gGClpZ77yomx3eEBh5aMhBurU91/0
q7ywX0s3EuiXfL9jKO+K+3Rm245GkHsW+kjgLHSA7TTkBkg6ly0LXWkx3ZydNgI5wX2fN/OAoGC6
VOVOMuUQ7so9SFCsk+Szrw7NQbGMDsoNa9VDeSsMgn6eBQrHvWxrUWEdcP1sjKMYG1EX//9uiVhM
/+kSmieTCi21csSzOpQKPWwpZe7biL1jzRAw8BcaN0wSewRbg6XCqOVJ7vy4WykZ81H7qk1qbQVv
3EvAsOzafE619geevEg661zjzPnmIr611Ae5n77WdbY+YQF20NgHFzVQQRpo2qnsCtp4Mr7va4Wf
Tl8HUr+u6m9JgGPGQa67E2ILv/M3oyeiEdmxVVKThFl3o/L4g5v3ptji/DFX27nwjAhybjpBUVwh
SLEjdZJ8fb6/bIi+hs8vD+f/temqQM78rEpC6MPYEfZM2KqArbHOVgz8ny8bQYz1eYPnarF7cuMh
FGIp9VD4RoEylpmgYZvIzEsgtwuzmk7BeCCMjFMJz+FIOH1Gcr/XuGLufhIrYVpT7Nz2QLWCmbVk
T5d3ywFEseUVSMhChF+IOvJR1yzhW+KCaS2Na5ehSCGIiLdAqe8sggJdbIZk+pkXl0r0S/hKZh+K
S0A8siWBA9fSDQLl8SVFBdtMcK7O5DwTMXdKrgF/LrOlzPLkCFLKO4DVE86b2Eej/dKVE88GlmKH
Rhdi6dOyKJj4Biu2WtSP17PplCQGlfrB5D3GhAiXWCNwgPvEuhrPkrNMMB/X8EIIigMdaZDSNqVq
eSi/5RvVTOmc1hXkIwwJtiXh8P1KDkH5+T3/0AOEQU3DFwjG0hcwxY/EJ6A5ZIbdqVnWznzENAMV
zPLxkmAJZk0N/uM6yj1Q0BTqIenVnhSc9ubDbrtbMq+1ufcB8GPaKj3CnOecZdnLuT5UayHkGWdZ
Fh8+KoTCqOexyDLDAFYNqrlVTfEk/R+3KbAhro4Uu/4SeFNoH6//lZaMBDpf9YhwWlvA2ciNOF7O
vfyVpHPqfll7cMT9E4ufdZNTC5mypR2TfqatLx5Wx7LHwvA5hkeSOT4YaA9qQ8VE+Kwpg/CgetnD
A/+Fh3KQe3lCJKIFlkWgxoEaW0Q09MLjUH1ubJyPN+MScLc68YpV65wcvDiTaUCkj1e0FmQ97V1I
ApS0sqiLUKY7Q462Wa5khSyaoRlGxP68uWeFZphW2Oi/qUaUTN4DJhAVp8o5NLgmNSZzziO801of
ZguCiC0WzJbOab0XOnnaWBNwjBWexiVzn30ZYWKQb3HtpW8mZXiNW14sbvO44cqRbKwjQnPBlESY
dzXwacGAdIDlk0n9IgizF0ywjLy8go+EcWC2ylK0sK4oNKqQYf9TwGnTh9WN98bfkSF/dY7kcrG+
O5DRrQhn4vYFx4UHF+WtF00xhhPN+P69qFa3XZAgWu43aIDGg7AuD2yMf3HdQomb7J78rivElxaG
IkdGSoiQic0U3Mqx5WPLqVJox/kQpx9l0/zkCUafh08Z/mDxVD1SEI708F7/VGoQNNR9qCx2tTC9
o5i/7WNEH/JtwsP+ZsgIsxHqPrPLrTCm67ryjK1VgeKcwh6wRbOTARhCRKaQs9SAlQjWH1pxIINN
LEC5cgZ9pnn9cQZk5+gkjKUPBcFzuzpb+NnA7NpTTUYym9qr7xyVheN/BnK5DCSEmNeJUuaVfv8h
CrDMq5LWYsKUB113WJjwMyAYpU43krGWLyknupHdwzNwuXBvlV3wJmSuE6ePXiwG4oKXMV+yPq30
FNJJBRbSMYaXGJ8uSGvemPUjO3isuhw46br5mBkSJmVa9xbAeg6fyjkmuZ+lED94iZANZE/mRKhY
5bB29NJoe3rCqXXn4YvfnESAKbffldW9WD85Ve59reoHfwKDUpM2hE3OPEwwcKMud8gCDD4j7GWN
G8uF+pC2nxfuQgx4B35PjcD18LfmjW9N2BLW8x0JJzEngJBOQENi/fu7ugrmIfi1pgURzZC16d4A
oVNGU6Smp1MutAx2/fva9lhYpeKPFBuRpRH1TwiPnZC/tC5uf0rpHRQgLiWhuEhYAAYh2g3l79IL
eXvfsMik4Gok6yd7dVIztCdWVNLp9vSvB56+ThDvGyKhJJHZLcMyKGLSVdMpBtxEt3LiWYn+WB5g
EC2pX0K+7Agi9n48Qxp8xVlR2mP/N6kKT27IqycL0SmCBdsUNdeyPYAijcbH+H8VO1m/++l14Pkf
gbtc7u0CxUJvAnIZM5x9rh3vTnpoMmed6qH4Z5F96AHP0UPqSoZlUMlXzuBezr6MJrJr9zuVc1Qy
sn5jL5OkeWaFu2uy0x+iOV7g2fDbJ80oX2KvTbdcVr5v2lF7a+hbWq+RPNRyhF/gCONtEeFmltvU
rXoeoN5CqbxDXsDegpDeRx8hFs7OlqTw3tGAMF2yiBk9vE4tkxi4KnS4BEX+DGTB5gQLSZUHdWWr
fs0S+csgZczceTEtiipqlhRwrDcmGqrC7vxm6/f9xbFX50d3KQkqEURcXAysvFM94yCz9QiSrtgn
XNdCe+eKNjqFtzOru1XVLXnKAPcZsq3N/J/sOfEDbCoUY+lXrod7cFAXyjeB6gIh457LA1VFK9so
ohf8FFI7+/GBirZfGRuy7khxIeUOwTUB3+40OD6Lbou39MrhgWCPoNEeC7QMWGf87MGk4GDVLxXP
s9hW3Ver0aGm3+1gEPvFioz87YStcKe1JUbr9z3P/dtP3l/2ulYklRXAZ/hgiO5d+tmqR8N6V6C0
cYKAfrf7TIpUJFDlYFrWsGlf8+5K2cNMC4laERB9wvHqo0RmR1FehMtNEuwmD5n7KgyuaOxkGseo
5w8vtXDyWVxDcOqPUMDnWWuCMx6M0kfLMycQ5FFCK7kw4wedXgY8kj/IAsfwOBMuGjZX2yx3xux3
V11XAYFimzfIMVyphM4dobP7+A1V7gkElbpW6kDpoggy/eXtU6PSOcMDb4f7MjiDNgo3/wTY8nYJ
7afcoJs1U8pfRHNz0MNGprqU+kslO73Na+NFw6KWGnUAUMj0UPKjABb/nYVtTquxdksTEyTTM4MH
Nic5182nOtwLsHo8QF1u5a9mBbdYU6zG0YgoPsjlovX3r8fhqOiXSOny0kY//SXj6nqrepG8nfVL
TCO/c07UekYw/L8W+UMUvEH+8hyLAlkYVIJZF+m8q9xVvIWJFBJArfXxLXjYdkS/sHiI+bFi+AhY
YQGh/WOfFjiULBywnYS5a//DR1gwrFLj1qgBgvsHKN7EVNivKpABgAGu+x0ahibpWoXetmI7OpYA
1qScla508qcJoITsT9Ou4fJBNk+At71hlXBoUVu1lUVM49JkpcYYnRis4IpkbyvnnBx9ohNaIboQ
kwnDPxypSc0dvsHcdD2JPLxh2NHPFP3P5MwHQ8SK6DF7V1jtIEHsSXxwV4/VZoc39AT01D3YQnqx
zKjhpRP6jLAC6DgV2Mck/+sOYrzIhng9PD3hXm+OjBYRiQgrV2qOCxGjKm83yfBGSwVLiFDuI0t2
Tisby2kiVbtqnVdwtHEMzIFHQC3nLZTagfC2k/v/oCqDst9ICq42fMWNmmd/aVKQde5oRqnB9RrI
VSLuGwtQ5tmuxKsdEXYVSY+kduzw+SZIlwBJ3Npwiv7Hs47AGQcEQtD2eFi5kQpnHTEKo6G/DE0B
scAsDDbWN48+j2e42VXTUW/pSKm2kVkln9SA6LJDjomhsP0LeiDxXqjpkKRXvQwrkue6nq4I/8+w
SN+u/ilFUskyuzhfm151NV/W9uDVHPwrH+wlakIZvJZpya2Ml1f4kt/B2jiJJKItJO3N1UL8EPe3
aWe0vcnrzW2/zPRWQSoKSe3k/oXrmI51BrnyxMiqERP35IdfiPqA+9fzL1jphKIr6RgQA/MhUqv+
lbSPtBZvLy7yLh/jgplgr80vholcjr0LdLWBEANNZbnJ7ergP2U96mIOSmXa+JKQDQSOFAxk+6nH
0Tl+7rmFncHm2MmcJyXf6scVsOinh46oDc/fyV7aJ25DebA0gTbkLae9Jd85O5cs9d0zvpvLaQMC
/YxfNMLMQX2yA5Kc5rOW/kO3ceXznVIGbX/8tFwWY89hwUyafQBYI11G1UnY1722KOlNNNy4tBOo
8bcvuvaZ0lyrbx/35zSi2vJg3s9PfKOibyhC9UX6Imjk5WWMCx7rXvj9KZPypBzpEFt0JoieWkTo
0M+LGaf2uMIx+RJyvtTzkqDrEGNUBqOC+NmBVrNCd0DfpIumZcbZu/mbb1If8itQLStIwLLuhdJT
QtqRSfSwGN/7bq4uWFuYKamo74Cg0jW0oOzekuvboj8bnd0SG1iIr/hCY6DlPJB3A6DgcuXq7uQS
t6pOJ961Fh+9pcgAXTeVXtzYzK5oAlRNEq9ZRfEZtm9hAZ3ZYW3fKQY8wUberEDoFUudZR9r7I4E
SB7Qi8xrNajRxklcVtdCN4qHA1N25GAhwEf125FNUyv7e9CWuyZIcai5GlbC4Xstby2wvK6BwdVj
fL04amRNl/ZLjW7QTAjuMLEuwhTVMoD2Gz7X9hsS3gLjp/R44DjHN43dCn+etfo5UEkwhV/GYBJ8
0ti9yZTnr5gJMLFJ7jpz8ZlTcB4zr2yKAnEZJ7s+VI9K2VyhFJzLfLHxvGyQ3cbUhCJaPFH7Adx0
eiinnYGe0LaO+W+xp7soMOY0930/EmmnYeSMtoA/5hKHONExTQbzq380GPVlxE+KyOOAL6AeNKWr
ehfmYNFIUhQNutfBO23klJVXeF/Ckg9b5HoFFiz6Dy2asgbc2FA4bQCrefEOS6fFcs7xItwePGIE
JgytYqX90NzpMsQemAZROS/EcN9/qwYkZI7kaKVBDxkpncFta1llyupN6iDq92xuSFrkOcl5SKsR
ovPNAo9W5WX4M+xTYRTwNWOqYq093s6grenxQP8USBrE6cuP5qVQq3rOPfJa/c3Ej++WlM9QDjWi
Mq2PvnTuQl3CTR5mGj7L2LXZhVWp5ugOKavKS5+6ut+ooB0RQKXDgxVMfnQgbZQFG/6iiDeAbD7F
4pHrJkABXjQz96ET/MOxfyuxTAohmF+iVqq2nAeOjfShvAjLYzJogadxbNSnW0uEP56fsFlGsxtC
xfDhAVB8U4MXONqdcL+0TmlZ/juDUovCpXGf/ilntBZiWd8+/I/vyFr/AlY8Lj4rFWn6rL4b6bxC
WTgEnzXA+8p0xnRu6DgGMPVIfpJVjzjptpWHz+Zatx7id8I3XkT9+BaTU2dLaRhSsu8oaNT5sT9C
igUHGQc2afJJMTksDPnGhpdOfRibW+Vd6yqx9RtLXrbb4Js0sycYskm3GB3Sspxjqdf2l2ByZBCV
yYMzD4xZC8ZungFWCFfPxrJZLZBskIUNaxsVoCIxWsMxEHr6esf8ki7j4fkjukMK/QlndxWBufWz
UL8cDrmIw2+6Auw+V86euQj6ezQGILr6AAMeOP5w+flOun1m8ceHou0zyyNSh154Jd8rjFgTE4Wy
oKI8NhjS9WWxb1CObOUMcwGTzVzdzhBxpPTwMEugpUNz6Q81t64EGmN54DfYQ96rHjKcvCH5PhU1
gWw8/KyPPiFl53Sqs5U8Z8z5sUcKePRbGRDKMwWcBclRZlZ/pXi5u09ZYAab8pGd6Ba0cVX3HVv4
AFm/erluumtvhu0uh1ng3KXMrc4wIg6Qmtpa1NHeo/cyYIrpKV6rtD9IWDRMfOtEe2B8YQjuNKVp
CT+/LDMglJ9GfeoOdvqVyRKZaSk3wqfT8ewD0L4jec0z6CTsE3oEwnF2hgOE/+4yRVB4NGKBTlwI
hH5QYVU6cLtpldX3WblRJdI89ugZbfwvIN1KKz/xJQTiKJXiKZpUr4Z1VXoLFafQjr2gQOziFT+P
LXnoaelDCKj6XJkzVyAPYAtr2ryauxheSklJEOJPOGRpgqE6seE6QNpbewhRqybnOZ6gAB4uvOkZ
n/RMXhqCCeuQSMiUOWc1g1e5zy0NfUFOt6AtrPJdGytd/od1qeyb/HHWCY4r9xFNoBVFvc4QcqyY
JHxYuTr2JnFghjg0mobUz3xHvinbPmVP64G8XTg8PqjewpYzkgx0W77RSjvRd8OsqBg1e/Kanl6l
NB9UamiSbttIqAXNrOEK4muK1Ych1jT7GGr0g/g1GU0sAh7C/Bsup1ayY7byGDbEXWxif74/0pNP
EqVcdbDjQZg9CAdCvgKbzbR+1qPzLQbP1qfw5pKkurG6yqzwdTq9KsDDiPEo2vfv8U68YnMjVLil
T0d3Vi6yd689zDO3SEXmWC0pTHrUJIVWnX89kOMvERs5mOynTBDYD6iFLCLQLdA+7z5OPLKs/SyO
LXsTcQStbWnm/WCCON8jqX4aQjPcJFJ3Mx/xgEIIpblYJNgbXABLoY7ofkpeQ9sasHKmEpfOhQMV
z78wX2p/hnOTm9FVNRIpxUagAQS3GkowhdestSXaZ3nui3zUtLhSR1hH2oTzyhgDCY9ts/tqsi+q
sndwuRfYTFLGc65Zq0UWnwBAUPmYxxSgRKRGcLUYmJifm/azpHGEVTdEBVA8FgHkQovTiHiXJ4oJ
T7C44hW+MSNoqfKZXYMwckQzOypa1zSphLaj5zt1JjGFMHQO7L5lLeD4YRzayAjL3P4AjOf1N6N1
gE5J96Ilhh/2HLFXQQPjOfaUt7rVbQ2NtF2xN8bCrtIqaUxmNx8EbreaDFy7mbjXY4b5k7Zqn03G
8FJ95a/in8+Rqb9+hvWGKdCg9F/K0la/kgUhdb7y8sBZhK+vb2w4u4c9cM9BpImOR6D+dDnBkwlV
R9Hk1tsLAsl6RbNY0hZlGXo72lrHevGprGzkz4lhe4KO6QfAcb4u2dBSp1fjE9ZeRsO2elw9Tmcb
E3tBa8iwUUzNSx0ZonoCv8iHWGctgIsKWl9BHGYQsuWtuWhTbkh75EKFNMcI52yfUEQ0iCzjBExZ
yYx15/ELu3fAWLpspTEJzns5ElDejaSWjR5Yxmza68fOSI6VXsa39kAp/3OdlZSieRSRdiOR7ceS
1Z6B5TeH3rLbp72D0eIkD+Gd2rbIC6Ha8A5llARJAstcTUEwOFkrqEnmLdXEpwTf2S36gsY4cKVZ
U61SGJ+YgNBM6kaRv276vUizhmRkGg/Y1La7C5AVT/66Esfj0gh1ZzR3Sc1UrBU6QyNpSScHkc/g
PNspF6rx+a47ypikPV8126Rk8zt/CD/KlCAhscvS6DAW9T8NsjWqYGfU5k8lOz9PJ9KumMe8HMft
yXi7bBgjYSNbIkkwII3kZ5Npyn8ubzrVJYxmM+ksC8BrFcReeqCH+K4peFw64ykwiXCroFPG67ks
g/3lDEXr+4BGH5/YSUw+nOIouu7pbaN538OqZaGhc+2ly8XTWur6CU/EAAdkkKVnFKubI1rZ55h3
sc7Mi2CQkDZWrT4RqEQqOgjOVD9fz8YIcY+y8nSwXFjU6FAmeWob0via6qK4E/6/HBFG8vO43aWI
LVjkI0A3NppDG8B9GjNx/ItPJK9M8njesy2i5SEGd472+dPkj898Es1PHwtRQ1Vvb2eKTWAA/wzd
i67zZQgkYsH7vIfoHIwXiDnXsVftGAqWn5iJgA024Hhv7qq1s3Sk74i74s+HfR6dZmZeETKJzCV9
fny37x33s6LG2+IlhnUx2axUV4qdguKm7TKAKHedCICDogZnWJoVwuhI+IauqlsTkZhbA+LShcDx
k0jaR9LTogfD+P1YEUu/fAxNOyTdUfhcDV8KOXDW0LdiTFirC5kh3VUhb+ex06d3ipGBgAP+CUBa
jJZrLVq0562HukjfAP/Zc8A0kcPca2hFioNxzhVR5w2/K1VwACWIWAGSdExUiUt1GQMfG10Jyv+l
26CgwsfTfh6lSkBvwMpQhZ+q5hW0/KF9UJl7vRHu5MKR3lEZzB1idg9KEOrBVVk/D5B4QLT8pAn8
wLlWkg0k/ulz9unIzTohs0id+BG3qL9LNxTr3z40Kr6lyq4nHsF66yxbjoXYaQAOXFHZSj+8ADuC
8luy5K1xNXu6aKYsT2lrrtuBk4QkQ6FZUxO3t7R61tzIcGhOc7p3iJbWQERF8v+jLJiQYpwUjWFE
JKsoQqgdXhdgcIWHNrF7fUCqT0S7p8k3hwwL+PAVLB+JT63khDJpZ+0+xqo8+nu74sdjteqOd++V
8jnXJT2ZyP9KYL4W8zNil9wjVOE4zTSKVz6RnnEx4LHdrzNrgxjo6LNT5iYJ3dXvrQf7S0//Gnwv
ThuTxrd5C6RYiNmD8pKqRSOS7ab99OghiSe/CDrKlLWxR7BlhHbbhWak7zHR7TWEnzy+BUh5PLEo
ly/0jTH47Wd/qDO6TIw6QtmRKmFtib4N8nf9ZCZXf15ihbkTGNcqlrGGP1RxQ2ne0uKy1ig/G6+W
b63GL0m6BN+ZG/YpRCcVKs4MVt0sp8NAosgAhNVvepQ9ATgf6EUFi+/d0zhwkP3esGMVuXm8u7XG
wGjJf4DOOtXI4Fb9Y8FpWgBNHP7+S9IT2MaKP42C9IrXiXvNZgTwzzLExG1F3NpisIAa6k2MaDGM
fdA3UvQ/GoZioSebbvbqG0OZ+ysXNoEjjKQfLsf9BPMzu3lOv3x//KvtAowOweHWDe76jCwhiDe0
1o3QKOtsaMyHA38e6PA3tW6ybfIJyP7qlf11U31iozVCTQ4iXfwPGh0h7XuVfgy5lGL2zesYcd/k
G4iii1jY0Gf6rspxeepleJMpMDQxvIOu29x3v1KuBtRXpDiVbkQsM37lmoUCn0ACDr8AezqztJvE
c7i4wqmXd6f7ySHcA6pLf/5EmG0scgkmfR91lFnWc8J7edSaAb3uVAppAPQyCiRe9k/h6GE2f4mY
qMeFkGwp/50VWrq/oIWjV79e6MUC242aDlKJq+brir/fWS9gl2HBZ4eTXY2S7AD/Uaz+vwWMq1XV
SipudIo3BJpe4pkgQIkVB07Z+1XmhMzG3beQzTNEVkoa96XRJ39xsKW1nFHBgLP6gZ/fJZrpAPVQ
z/FWWE/Uuso7csp1RUvu9JqY2yJdj4tYhdTUJhLOmEwlFRJ11UM35LT9Cy4pvUxTdZZ28IeX1a1Y
9bdWwnS74Y6qxxaZNbi5hypf2kDFjmlcCKLxYxrOyI8hY0qCcBDx40x6ehboaPDmllWykZGNTAVY
mzRoDsOz7iS/Yny9tPbLDVwv0+N2nQH+eiipsF7oI0YJTVdZAx8Yhq16WBOyVO/RFCvFFXzeW7sI
oEOee8TluOLF1xP2oStPkH3zd1dHA6CpcSjrWOy/vma37jvjvMiurDLf60lL2FIzyX2jM5AUyYrL
63NXQGiVuLSAnnpy/HD8pf36ApxGdXWlQuQRL09unjpToB+59ckgsQW5/z89GKWLjEK455Wm5gnv
5+VkGv49PGPx+khrQ/bj7kRaIzvfc+jJsyKPweIVBK7eH+ify6NJdkWlhSTQ00Gz3CfLOuAkXiks
rwoS0n33f6ABnFkNOidSroVLyBkSxqSiPg75/ldqdYmJLq11JRjn8PLceJBfNI8ukiXj627ptuxp
3kFv2mHhB2xTe+83zXl79wNMR+IX3BCCDF5YJAve1BsL2tZCesydYLYNYRJMA1bnuJtsTpc5hgiS
kOPGeVFWXdaqzoQcBikkN0E/L8m6TLmxCciwGbnqMHTzgdOeyHmOQK4XVyKdQcCumNH+zpdV88UA
yig1EDYSOwOVKNQjNVmyvS30apXnmlElu/aq2/GPeWRNH+ZxIw197tA83pBLZpVzHzvurB56TX4X
a206sVGUeMVUEBHM4Hn1WESGdYncjYeSH3huVCYwToGPzDwKVVT7WeO8+S2oy0WGXMs9Gc77AjTv
Yo1k/wp3zK9DoQ8fF2H1OmS37KzRuEHGmYeXCnd1aq4Tdl8lY+aCrw5k+xlXMKOXVVH8YfzADKgr
pyculGkxSVPt9vIQ2qqSOBIQnJvYnUyRmE6uESGOtP3MPtNBOGyN90gZVjx7Aw/qY0rm4elnPPCJ
kcVAH/OwHHDh1NN3u/2y7RARjPvVOzKzGxGnpO01ys24w3rkxZFAKEx+iyFZqGfXxAeKrcVRs0qT
mhxinR6bqkQN8p1DdFRSIb6lDNBodkzIsRiSkxOYYPJ9wLX9Xs/MBzk+S+IciMTbdhq1BRrMT3aP
nY+4z6dKhnECLyQjn1dKzgjVtcUhtdQUZmCorfNVbLp2T7FDWqWVsBnuxcBOjnsmJWl3GN3IIDAG
U0b+FBmXWtkKWuBT9v4Zgw65BVs3woz4nSIhUAem+GTpFOyswfJ6pQuaEjx4pw94Ut0zBJNp7tnG
oaL262GYFC4nA3qfHivIbXeDyobp/E8M6mUZQEQ9MRQg+SK/HIZvOd3O7c70y5sXyna60w4yur1C
1JyKNUtGZMlWqxtlmRyUJXzniRVWAt2v22fRdH0NUhA4lrpK4nfzb6lTvZzscsByJ0xkNCxOkGy9
8gS7Z+NvnsIfnuRRtcssZSnPvP7OBGU/2MiLKNgvFqAFKrhfGCG6gxa+wTY2pjIsBreagqfFDxzf
O9tUk0oA2qIMgJ5hU5nkSZ2Za5HyNwMZOkSXXng/7zL5vOkJlc6Vzph2oPIVeQ7VmjhBe7f/n9xz
cf3Lfco+lzTBGlCSAr7VSEK2VsN3DgezPvIRVqO2axNdS2f5yvwOb96aIixi2nDNRPbjTSL45Wjw
ftERMppWyP/gBkD3MRoh7nrjHqaVqM7jzpj1eSjuWYGX8V1jg1qK5p9BmI8rX2GGeXZ7pGkRON1T
ASCaPzcf++huzN1mpqmqbEh3CGbox39nTsbC9cFOLORLi+segYEqimLskKmuNXn1Py8T9Msxc1um
Ajyk+M12dNc00lpWgDH5XqDHcVJokw/dAoH2VRqGYfxtNhiuT1tCXE5VwRLu0Gm/gnRQiEkjknCm
rBbEOfL/RiF4ISO4dDdQn2rM8D9geStginQb47HaC4kgjRTBLNXhlgN4gCsAmrhOMcWb9+8T013I
rbD3wSiuud4z2jrg/jbEfDuu+oCkZodcdljMKhFa+VYtdcq9A5QmFQ2291Y3rSYOfpOzMjBJBqko
q6FE8PzqXtw628jydcsjCGVWpOe/eOPeewgZhCCOVSbozzBVsKmTP33wDSYUXSKuieec5Uac+9GC
qqwHQYRMuU+mcjnESRqf9cYw6D8UJqMD8cDtuDxTIJDHM4rBs8yOerLrHJ7NH3wUjzvtPC/4pwxE
okRtY/4dM3bmT22aYRUWp5QhEMCYIpaNzRyCmH+/xg3hNQQmOLp9OEiAm79An++Lv13GveZXLgqt
TPD6L/cqZ4IK6YMCz2x24whM3pDQoGnMLY75/JWipLGgzwhR4nlQ2uftNU3Z7KUj+uSR0EdUbGe4
/wWvR7pDTqsjc9wno/zRBB4SAd6nkhcvqqpmBsvNctajSx9irSkZ2jOf893HI24AyrYyHFqftgsR
M1C5SZHRgOjB010mSSck/Usdzl/dKu1YBU0dcQ/QP9l1KyR/ajax5G7p7c703Jj8wrL7PcEhOC6K
dqlno+Rt7XmRrfpeRIXcye0SqWz/vDlagQWyO6qNYPYjGXk6Ii0WI4lb7c6Bt7hkWipr7TjvuIWI
cj0bpfs4sTaSx2afAh/RYH/vKCCLqLO2KKca1vt/mv8lFzh+l4y3RHm6swcBwU/PMbvkZmyxNtbD
vb3VW1A8dq2aJoMvL72HiGShJcT8307sGbBv8s3oqg/RAltJ8hqdt18Ac15n6I1YP6ZbLhT0D4TJ
Dw31JCVHLHmMQZd36Rzbv6wCFtp1k+lUqiRwTSW4C6kbGG6gU4mbmGDFm8i9EvBTDyuVkLuRdJa9
XUBaxGHOaOxuSgWAgnEHu1gdCx4L+MFiIYVuavw97mHKRCWNZFvNhLhtWSnFYO5SAEBk/weFsoiu
yNa0WyFFl7fP5F6ofnQ4cOMx4OhKaJi49mp8voYCBNmHDpqj5pVHW6DTm5N0kBSg0nY/qJrOwRJh
QQz9nhMVaKXMpjMCx2C68FrfO/bu6c9tIwpgNmx/JZYJoIi9U1S3WMBTo/1GOVqlUZ5D1mWIxzYK
tNfIMyMmLad6ju7DGwOzR6CsJmjnBkP0D0PHwj0R5U/IxKFXPSnS6y/uI9MsGfbpv7W5ueVlhcMe
+opbYRqcT6iMl1BWnghEuwUIGOWL51l0xShg4VT+elbJhv19BT/ruoA5fwvVtZlUABbfTfzZfE+Y
76v3rPbiQQfLbQDSo73TpQq8EAOyBk5PI/TgyCrSGTpjOV67SNpcXqTR0xLvsKYNpvhScpUuGSZC
9eQcw01CRwoVqOlT+QvK1wGj1DN535vfpogHV/JCyzeZ5J01gMW6Y1ErVW4bBUr+iLQHiRbK2saI
ocd065ZjWPY2fsWR7rnEPtojjc1BHgXMeDNAcXBLXt9iBU0boKwyJ1fXgdE2c7U0dxQc+ejDG8y7
w+JxpEOJiBJXCT0NvFNDso9KGKjk3YvWnqlZ+8vM02S4A0DS2nOrKCR2Ad0gLAxfWcZRylQXCHBZ
ePpeAibQRssI1Q3YlRbtIRBBVXE0pfwrhEzNKpmVT9dbt/CdvCtE9fq1AURi7v/f1UKIVvx2Kjwo
fONS2Tp7W6ePzDCyDOs3uqlSMXUR01RQohor/a6XrTYKmf7Ua3Yb8xJMZHxGXLEmmctBwErUb3lc
9YNRA3XjgiBVQe+qxBp48Dp0FfbOkHigu9MCgt1QX6Mginb+lfid1qc6kM+grXOmj9Wv8e8zAKnx
ncjkgxigFaV5env7XvIAQyz8G7rEaifGNN/0CZv8iVbaZ8Uae2UhqzMJwAb0MgiEGeHf4fnI9l1d
RQjmOsPnlGnshP8DjBPk65fMimbUXyGbOPpuHYAvvA5fziqArcFtn+NszBEWnsbI6PFPDUHwtExk
zT0+t4t5fwvujqYVutQFYL4KEI7mwbg/dfxIY9E9FHASXXjMyI8RUXMNYCjozvRGCjUbjAgSt0qX
Qc/+6amASokYWLVz4RbTAQ+JLwvKQEj0axhCfDfguljTFCZI6A+UBVh7U6VgqLPiDi7A3smx4y7P
g00Qpz01kHagQXiPBxxGHN3jDPm9znKQSH7hiEosuWzrWEIIvbn4CwFEUrtHQso33UVg+KnN5MHJ
Te7jNiq2rUDmPIYCw/cRaXIufwRk43SgVfJaqVG89XSktlV7Z4SmPbCRX6/rO7D16ggsZqQBRPCX
Aca1SLGlO5KX21kfTBz9MWYo4zAfRh3xqN8xJzuEqYBSpQHpVHw6IOm4SGq6CR3F4Gqr4Zy1JYpk
eDIgyLjidZPCN8rXt+7KpPb/MLM5yaACFr8yVCjXUD1R9aRCM0hbvAqaNqIB1GRd92oDRpHfcwJh
X3RxSb8KdX1I8AW+miOfFsVJFx12jmGqCzALNIm2lsBD8DTshvRPPI5e1RbcU57lbFesILEdiUYo
lh1j6GfgLRAtN1keDT/a4oISmWTwtoT9OjO7qld7FPY3oC1ioGqaS0TSxvZB3IaRx+vykzZqbYkv
TBM2rxQjGm92X6Gyf5YXzOMO72xFtTShlHOgdiwLc7P6j6d5PMcS+KBFd39nElQBw/08cInQsUAy
7TWxzyeqQrBHuriET/Z5TwsU3oBUuhkYGKRTYJ04gsdyBL2O8vDb16Jdl33RDtpMrikWZIulK1JA
UxWV7P3pGNOkLGvXYf8lA14BZK/0kZPCLmSVK7KJqLwbfHWa3PnZcwvejwk6O3xV4uhCbwlIyMdZ
YHoqcPuuz0UYTMooCewX9SQf5UOmMkISUe18DovR9H7yXhJ8omIBsIjoA/xknWAxryMnFDOs75cI
NbaGcvK6S5SIcV26hNHtyM31YFj1Nqw1a2O0PfqPPLjSp9jfJ0W6rvATiTK11GB8g8jqr3YT4eat
36VH7m4eaBAT5E/3ivSQoZPJN02yLkd1L90JAaUsoIz0buih7rPXHIro8Z+sRE4KmUfwjBjbJC52
e5eBbr249jWorasH3h9qCfyq+oV4RSjBmM6bbDvn2XJgBdc/hWDLwciV6/pXIuQiwMro19LEl06I
3j3AdMBexLDx5VBtZupR42m3icJODygmi2URWmvIP81ZkBUGEL57kMCZ2PhLhFfPbnWbNZVLcsfQ
fab+R25B980QHjpXeGLJ80cOKnhuXeI1JV1qhn72kNgv7TUe9mX0evUQOV90lUWbXv7WwR67/1y/
T3O2WYkLQCH7slMoVBIn2dqVWJcLaayGR6+DuSp0XztkaYe4smLhCEzfXWpmz04tf8ER0sEV+g/h
/SZbpePcyXsIW/dApSX8BGiS0URaYv+yMvRhiKKu+XGrnzy0IFFM91hLVdXSTdMVM+ks9wd1R9FI
5Z5Ol9CwinukH15EOWjgGw3zWpbrVSMrTf35nsdNLXgK62X+1ftoeRROmeoGEbGmjawRYs0L7F8U
DTmckFouVEty483KlNBN+dVK7OPsEsuQ1O0kxJR8Du/jMPZS4evsUohHrvgEo9XOzWMVHWkYO/0V
nFvvCJ08JOKbLcDSgIa4fQ0/RvkkTMHtsyk56QKgdwqgAcz6srIeUHf+hnKoiA0vO6qX8OWvFEDa
ZrRn42IqCXbt9449m6H9woNV9NlVOlzLsvJYltxFe/BM2hrlNlV/jgIlpWMce5lpI8kx1zRERGUB
GTm3M/C3y0koCXw6KNZHGgOIH8r+NLIInaE2X+Su5f3FC6eRGTVqkyt6IdCGqF6bsTmpa43FkLJK
NBRpxpbHMRj9uARvAnV1OftWPm4BhMK8J94Gfn/814lYfIHvi1LAl33gecEC+mm99K89+A52e1Fs
uvrmCTl0RiB5t8JZqlijNLbzpyJ0j8r/cC5H6GTJTz4zBmdyCaVAuFLP+07vYW8VCJ4QrUxK0IIp
SrHPDxIZwNh7orNv9Q5kOSUaU6uFJ2fp77Dq0Jjr5hUl+mMrm8TTDqa1js+wSl7ZZd/m5IehzeeY
5x7Qw5aMKI9pxdE+mnN0A9BFWAWtIucsRAuPU6EhRtJtA/I/ZW1GrY4lQsf31ZqI6pA+OMTt3mc9
ngqFZsCt3C4TKh7LvZEMlxEtA6nA+lNoMjQgFURk1pjlVaFO8YZJiEc4v60W27DViZ6m6WMzEB9o
ZvxQ3zQa91SFMIm/v/T9Wljhn7NCjCbgiGfmN5CxL5t2u8PpFaGQQKwGGPfSs81LbqZGpMD4lSHq
8mTYNq82q3DFNuXcC/RiSWNxCt26e8+QZoE1hHanC3pKptR/cuFDcUYjQ+A8L26lEJ8Vx+T7tQO4
E2OT/HgjPrmxxcjvVbKGrdjC3AH1kGLsMi3yxBNhW+n07As1PkSS8K96lGmxlFw2EhiwPMvv+NjV
qj/QXlK6COaX6lUhg/FkqUapur+X6B+Ksfsgn1PUg8c7KnKaI+ND7MaCqHRocoMp8UwgyCcUIycJ
/Tpk1GTXN1N/auRQFQkWOlTUBEnZChoHy+yT36QmZVb5cjDtU8RhnFYtjH07eHdeunjLsy4qY5KE
pUvJvU1l2d2uKVM1Xpu2e+4vnPGfIgp0QTAomSG3yj7ovRWD9mP5dDA9cGWJdfaJXUhNknEjtNqb
kksDI0jCqhZkUmu1vxkm+Eumco5zNfIqyLAC9f9E6HI709klJnA+uYdJkFXJtRe+eseDVQcWQcpr
VpI52dtwsBPQnp2b8tL5OzqE57rDJDt+1+V42OKe+WILYBqZ58xUfGWgBUb9aWE7JhI9HaHpcrHj
jcJAzEs+05jt6bFzTxAvzB34JNkeQvLKgGLKZZC1yrmeSrf/4CngBXeFQQ7w6Y4luLa7qzsedWmd
FJnirgUMT0mQ4spQUZn+lg+y4k0xW0kj56D57R/te8YQ/M2eoQ67t35I1VSafAW2RlK9pIGHz2ZO
cDOrYowMVVfwmMlc4szfWe6sK1JnemZ/lG0jc5VZOJde1eZcPDGOrFAcDyYEMocUubnbLAeSuc/R
Y15mdsp9R623XciUjpYazEupjK5BaMQKYg3yhDtFccLe/YU0ZIUffJ7MeW5b4ulSLHyBHdCnhUKr
Uh4W5bomL//UvaICcVlt0YzR+XP0g6Q3o3M6Amy9/MBEVCr8JiLjzVqyba3Hf09xwWSagZSh2YNE
MtCsg4zEKe1nnXdksq92/frpQZqA34B2nzpDvheZ4WOfnWeTEZmqHXNpetZO2a5EIMAvs/KC9G+0
DE37rvDSGEl8Iks8BdeHyDrffj59dtAjZPzk7McjngXarQLwoQxS/bNlds5ljZVUt/kpG7fhcSFZ
dYDra+ZugdfLq51NCVv5aRXRTuoV92j8xy1t9ON0xsUYoD6cIckTSf8Tqc4Qr6wuIb6nv7kfTbYs
zpP7RnH4ji5LGRQp/HpxBZ/aaxtHNk5vRoPVrepfZa9n1wIlUzkj69+rYfcyo4Fczq3lJ9isORog
2I9byZFJrHFiKGsucUoR4OuJyArpM05Ls+QPslsH0xsGaDvikOrfZEwBh1D9SdXWf3sSP/CBxqB8
w9/R5TnWPkSsoEQ4RNT6WdtQgPUGd/Mm2Gxelkc20M9shxtvQMqDTzLmw7NqMr1CwYnJhIx9q5ei
5wzqbI2O+TS/H6MPBgWP6eMMM3xmrlrjETdovPF8i7VGGAddldgy3N2svcUILdesSzQHQo2BLnG9
2uiM93YgifQX2yx7ksw7Aco6qUhcFZcLLq/RR1oxauboedYE6vkXM2BcPOUjC1ekACsu1ST1sbF/
kGXqEJPUcVzK5f+ajGlKNKwkGg+B1MZK5k6VTwaIRjSqogT/Mf4UxKPkc/s/DGLMTnOoITLg914n
JEhWEeEEhkl9W/YxZ8Qw+hgk/50QiGsC/VIxgDCZ+H2yfpsXjowYUOFVYBg0bcijXnzv6LBhthz5
qXjfTSgJ6chhjg8W9wdVIwKX4RkPrlKXo6tD4wV1vFYBL7pl/pobcc1HYePqcyCs9bMMTzvBM1XC
OsKTe5Q1Fxe7pvGcRtFVmR/OUVPC0deezrZgxZ2eKx4K5+FETpOCNLgk88JRVdqXfpmCaK0qZqBZ
TnCtoqkKNgdO14Ds0VrGuw3Fzep10Jk2HwcJVASN6ieL6RP2lYDjl1LYC9xxGuoIfXJ3tGSM9Wlb
e0DvXFhQZGYvpGJj/V5X7xn0ydh2PSahusiWwJtErpz6XRQ8dHnCRPm1u4hnrS6PCmhBlFRgcgOO
gVXiKh5Zqg4MamRZyfi6fXQ0fjU7+2NsnSQziIa7D3eMk9jpnGKx50PqbSsILdlILmzuJWT2yllK
OC/gEavJItase1+skF+K05ZSUzjnslc27SEozVQZCIOW9KbdMn+DeHCjA4Srna4kA1Bgyd9Thplp
d0cQFI8Rd3HVI/v9/7r35iZq1hhmLcfEP8u+Amqfb12FcidpEhVrJvVRVWWLhxuHK7IFACkWPOHN
qcva7GnRe0p0IED+o2/S6sbMJaZF869rZCK4aaQ/MB6jyl9KVDlaj6qCGrPXH6f4OYUPxjG0igE+
jkk/f23UBt/IRQTU7YCtOenVIppQGBdbYrz20bKmZ/aFm6QQjytmTeqSJV9q+aSZ29rJktCDEbwE
jQeY6evi0cmD4iichyJ4nuVDZFRx93WmVnYyPIUAyGsBEJ5aHuMfQCXkBZd/i55v2i1usCl1Oy+d
zCR+3O6uqfpq5hp6SKpLXjSAoYm/pemYxcQ8DtL/TshOWWTt0EVitLWGPWTQwvteMo6j6OWhvA8z
Zwxi3dikODFCag3ptNDmxBgI4pRBJFFiYkF8Vy19lPTQrb+qniK2yZ2n6GEDRKl9O9YtXiBE+DJ8
ROALf5SKkx6zVhamhmIUvppvglWfkeNvbVwidb+HnMB+Jfn1PBRydD/j9eDRMocNQKLB4IHX+uOt
S54VTJA7iv2vcQ7cAfxlgEAQYoKjnWBPlyuK2Ol25kSBBw4GyRrlF/p3Yz1dkfqTFtjAuL7amvKc
q7s2US8CGrGWmgVusilS2T1QM7ONVxHlWvO7eHN9K4Gtg4QIVVDWGi5OHa96BljuQYU1NWSG7hra
ItI4RpTknxIke2v4YVt3d6fusNv6h20OLxtHtjuiPSvcnsLP0W5GCuYiLcrUyq7dokkXRu0BjnCm
difu/ogBi0p9btTqFmYWyVcITdcacqZKonoAq1PrctLp3dIftALv/Aqg+hXtac2UxpdtpTFOKXU/
Qe0xZh0JK1oEVM/0SGpl/08xCx7BlEGjGs1PssRL8PlJLC3zHtuTtp4iRDc/e5mTrZ00TvNpG+Xu
l4K2Y/td5BuIDjKkOyr+mVm0pR2j9xHGZ8aB8mTVcE8B9QJF1VjRoRmxnXyNC605WsQNiRBmoWuc
ftOaDyGOAc/owCJwLalumHFxdv3cCksOo/SB+7Gv7nQO4AZ/PE3pesnBFdC9gh9LdyLGruUBtubv
XCbBCptjxU2K5d+V2fg6p4QDnNSIMZR94wyAaPX7QwmaxZMDhO9ILzmG/sDL+cB3Iyy+7m6IsEGC
7Uh1Vo10HODiqS1BGOCb/GSjyHUgEdXdt8stgZToEnuzsD3UXY1albPS1aQTwrrwI4zEHMBOOU81
EXePtqN1IdkNDluppOqLX7xLFT7HO36JmUZj4ih6j/JeVTOslRJa/0v/hL5hH90prfvsSZVWRf7U
UuoW/qCpIELlMb0y8rCim0hvlqrYK5cQq+kUCilcj2O9sTrSDV71gyEGXoQjwJksvrfIRXbD2kX8
VYt0UjOZK3IZOy0/axshAIQIUI9Q5O7bcGgClgYqojS0MqvSHlJq/qrSkrRAWI4h81BMwmyt9Be6
m1R6ojIzWu5wroBe/iFC9nckWc5f7nbbBqOpTXj8EOGRI9fGIAZcS5efBDDS6o0DaWdUHmRsgLCn
iKh5hgv6Sz/Tbzs9voeWLLRzlgKPPLrJNvdQiuNLg8xBY8FXe30mmNwUhaqVIxMLxxap6sFe3zAp
SYuotSAOp9ckbjQ9fft6ZWiU6KftC0Apu3Po/QbTdSAPJANVhJKe+qjT5uAVHp73lMkgP00Hfnns
qcnmySURGmms8FVy5jWGEYyJEfzDe8Rv5RmaFKZXvQ1h5V0OZYlvNiUuZ98k2irYrNXp2jN4i6sE
/vwqS9BppjHrxV4JLfUPaqX4mckJNsuMbKRXDAIERpp0Tif4VbhNoXerZxe6ki28GGRqx4F5erzx
mnRDmz7BTfhjn5YykjiWwH+NRbJ3ZYH9JqqR0W/G3lIQ2JFvctFc55Ny103Cr2o/17zn0qccwr31
NaofvwSmcZKkjZnwSPALPOAjtVlvfKu8EVDKtfk0KP4K0g8kVqDMpwyDNZSPRgmJl11oJ2bkajcy
pYUhjbYpakb8/WC42tBY/Ydt2c63J07VTxcl62ikdjgXnwyVGgfT0EzSRmPpMNKDxLu5QTspWqL/
ZzzzchIHRSmK+CFoANMT4O8ZEMinUCM8E+sMUDKMzIhFBYzNsI1fzYE8f6mhBxx43t+jKlluhlZ0
yJWj3t9u6aEfudn21KiR2TYe311LfcXzwNH10APQTIhU5TrHRIWlmW4vpi8LPk/2XxGE+9N1LQ+H
SKiLdhG3I2cq7duyXXcmI221hxHdeDMLqQBjJcVi3HGukDHt1di0rBdQv7JpsKUw/P37Pi5v/rgY
xVRa/6YwUnw/iBuJl0RBCl9d4Si1dKWwdFlR9TQske2XcqA0Hke7rtc3zv8vbFE5naqReSuLLZXM
HBGuDgH/0lfzdaFJ2lbv5gqqZbVVQxMCWRSBHCEebuxLOz6GN+Jxh4DNb/3OrD29OlETONRfUT6K
PoQAfYi8LYs+lneXlv3dSX6+Ky0MTs41ZBwk5x1vC/VIQ1LgqtfKjKJKzv/QYk/Pv64TuiHiKwAt
LQbxBbcW1IS9jNtMLDHBLbyhDKPR8XkF1D6771rtE+jcxefXHdSoYGDfKCFzmO2iKdKvBMYznbJO
ok10ZJpRV/EHWRZIo87RE1HJlphNcf8pEohVfWT3rMfyJG0WMJMXy+Sp4sAlnxTSrZ9J/g2ys8VF
YLux+DdWcec9aR0IM2JBt6Hcqbyl8dKX5qAHkslaB0VIvZ8zZMLC/arWE9awpmeobZoF4f9kT0AR
LbxA6lddCetIKwfbHGVtAW/3ze+PJ+XxfBMGZeqfI5SYJnVLZtJBfLe6z+EakofdUxxW0eaCpzQ4
SfLE/iZlhg4GfGKDsNsA+ZP/xmuEa9+Z8jd1Q96JsCg4mGevsCMUvYcU17OgN7MoX4U7sIXngGZT
m2b7JJwQ6RM6I2+D0j2Mn74vjdzXQce23y8jozqkFXGFzvl2uA0JB1YvdX8MygvRjK4a71mJK77L
Z9pdIEvTKNa24M2bJ7ful8uvqBVhPuo7q0lzVNARXeIexU92w2PFbh2hTNEQjaL1BMfB4W0HClgP
4Ttm3jTAzptrKqANRstp0+rT9Bbgg1rsVm9SiFw4KyPNyXmO96mpcLPYnQAgcOlrlVQBFm3YPpq/
JS5JsBnpmvvE3MK3AHeUvTSIXecoWb1xljeDBBNcmtBvw5r3hB+rk7Spoqbuycr7G8ji5lKy89Oe
UsCKPog2rrXhHNbav/LNy0KXDUTYcNCnytb69VBGIAJnJUk3lRwP0v8Yp8rdQ55LSuiIMPZAe2Sp
ttkaLSDaJsPQCrYYkPFcK3SrWdQjKujlvomVuBOXTVEixHD80VgVWgMJewMaO/SVNCyoqdZ0JMfH
LhJuYeZh6kQ5jw6L1q5YllHyUK5Z0WlUh4D7JXEqW4ApWnzyT8WYZnnmYV9Im4PNAU1SKw5k9Fj+
MYLKpdJ78NePvURzE1LMVT0d+r3uh4v96vpBUGZ58qyyx2t7Kkj2bbTAUCUhzvn2G0qkHW4tphHL
iqdEeZSqlDwxFYPwG0lZsCXTEwQGc7r+G8mXPJcSuSY7PR2CgY3A9VcDTn8FeqYrm/4uy1d5mIQN
5uYTbXmIaeogmNXrr3q1t8z2GjDZuuOZzYyeOM0rz3yQuqBlGSHR4SerIffs8IkyPpm0gx0uKWkt
Qs4tjQ+pVoj5NycAa7fbyxRVPD3pJfSxZ6KwGLlpyA+VfNy2a/GNP3L5joSsFERWwEYbGurrI/fn
RTCWy4YerjubGJqW7CxKW2TNam3MvJzN+bIVR5QtoWcMExpzyXOjdIogDFcEnaceTccvI12CC7Ff
gVghhxae5cZSV+0MzVIVWnk3nBZSoV2ZvBr0wPG3u8ZVnrmNgH4f3B2JTs2Bcc2EzuZYWQtHKBy9
2E5oudYWib/Pc09aseW89nYcVzhnyU+5u5KKkhNPko8sxAR2D9AhFSWAffX+sENT0Rj71lOIas9w
u6kAYzcizARXSgIzxbSSZjhK5GARvbiH8PE/60kgm96wKZoVgjzAuRfojQVRdFYRsBpx/R21JgkJ
lxGMO2MSx9/fd5RcKSvSAVxvMW4m1uMDUwVUafn3SY8bgj7FI0xxdJK/AMwbxMzWjlf1b3isyKAp
GXcCSycUIcmVt9DkeEa0h6YmKtFCObcYAYJzcMEIA5MuYzDb/E1Urp9XCvI8smgoibf5n6JqhVC8
bCrokKRGpNfDX/Xy4nW2pfP7ePgVK4Sh8ztkdPrTJlXt+dd9pbSR2SXcoYTgEwnw/trKdKH8wp0g
CvyTRab9p9tq6ejQkk9m0eVFdLutF6wB6ybCuh3D/WjOsgRIH4rNdyXohYpLv+nb89zMgfQfUkfC
ZO5fpUDTDUSOB/3ZnvgJ4VzsfcBK8/ufwuc6lSoPwau/Rp2wRyIXbieIxPuuU9/JT617WKbQli3z
KwNXt0IRRAToGRn0rpbuDN5mrZxle8uurtU3aSEdQY4RBaaf+u7ufmKYSnbK1t6KH+k2XxRqtvwL
+eWjI86cMjQpDtUtksbK4g0LG6qPGgATCdhd8yXYoZSDabjzBL0kgG86OucY/MGY2s+79sw0eoF6
WtQr3ly5UOPkY+3hw3ax24XyEn9cadV+l/RwBGeoVfWDdRy/ui7h/Ua5YwhPumIH6fb5QLgYQJmY
dbphl+dnaAlTDnXegVWI6BTu8goXvAXG6xGRQKofqRu9Whi+5OvTy12vr/AhfQqwcV7x5C8OhfLw
4SzEE55gq1GPTGSnkEAcCHfsV2slbX/47pneU3E7KknwUWz1mkjzVqrmT915iHovTNRyDL65Xfb0
767IA6HDqlBPFkmaKvjKhHKU+TvVKEGjwAv03ssVYscJCACKZXlvj3PaOu9vM6YFVqF/BPEcfLGO
Tpgh7LYS0x+tuUFTnCxUhlJruJoac8hY2d0IIuq2Mrus+eo6rqLdMCMlyPAY6q5x6Ajr43aY+waR
PhFVRBG9jaTiiqTQ6fNHPjuVHpdmnwjD6/IORQW4KjcDp5DX5mCFekxH3zXuTn47ml1xJpu1g1I0
oChq9P4x06Ajr8nIKztWUC/o8ZNK99amIAZkobIvobW6AYw5hUXvbEL8ukY2E3Kjtb6rJZM180F5
FniZlnTi3sul2XoNt7C9YRIOtcqZU1Z166XTbZ5/+eIf1wsjPdjPYJAtiJ47Twg9mAR1lJ2Bme0E
MsrW+odrQuVFrWVwvPWU1DTmfgbbvYEzK2mfMitYzSyCLJEfj70S9AtsvUlyvyAVWISp740YbrQm
CdUM6YYcMMm4VjEn3MqeQc/QUcNkCWXfSc3DIyvbWWqZ+hIQFNuRV/7EiEx8BDc3MbckI+lljqFj
PibVZvZsVKx9WBtesHK6BDBNQ0X25phsG7+3YTGpk7oE3XN40wVS9LwF1sPm/9cN21y8lX/rCfor
9AgwMlqX0YblyU2ePC7InlcGOhrD/rOz337YTTVZY2atCY+nAwSBPkZqxMMvMQJW1lJ/th0BD1a+
GXdatc7KdgVdiuoO11FbEmIBDdoR8mfdbvNnP1pEp0miDlSHuukv2LOJpDAZ35cEwDw2FNPKlYZG
POSQxrMwnTcv5727DXvwnbhWHhaKbFDEOseJXK9Gm7W6xlFaQtqzQN7VyjLKUepRaq9/Rft9VMz+
w5a8h7x8+O75O9H2hHbhZyz2AfCfW+1qk5LgcOfakSQDT7bTzEnNMCGzYeOABNg2koKPrLutqzMA
Qof8jpAtwHyYFqm8tRRM3ZBt0iFduSj5fOrIgRqInPUcYqxbrkm3D9FheLcLOunwRV3plyMc+pBx
DkZHAWbipcy0vmcE24F9rbT4/0HsrpvTlcxy9A7MNeynTMuGdURu/NE+M1/ZWqby7ex+d5I01S06
EFy0ZaP8fZuygvlGIH5F+Y9dPVey77vCuK6MXDslmwZ7/w3KaQ5lch4f/gUvIqOzpxgivyM79kgH
BpXDmG9cOrwP8A/upstefU6E9FGOa56Y9eEDfaj2TSg6va4RzrCGDqKutYqBAUdhWh52A5NOFdh0
XyxciX9ucNksYfVXOaLX0lNwl9bJ/rDtVSFHUL7rFsUokI0ZcHSzlEYL8o4L6PyN2PkNCL08qwHT
QwlQevl2wpYd3MBcB8QvB773rDpuX1YAXz4rJb4h3hEmMW9QapDV97bbobE4XcPTS+LcQoJ3ITCT
IqATRx2RXKAgITVpIWXUu6qZ3jgv3xkvig3ySmpGU+jFEXyHZ7/7CnxTYJ4FQCuTgwBcdOq4p5vN
gUSjp2uKItXpbTwcjez9xr+xgH29RNTlpsUY/Kk6mWRuR/BLU1WauiXzJ5xfc+jBp7N6QA5I5QeU
+WttHUcgdwkvbmP1xtyxq9ukLijeVN5o05duRS9KwRrQfn/ZeSqqp187UDSNCwkSPrxUoG+3AOJg
LGJWWsQmDnTQQkc5Xer03jzOtXZ0Fzf7xm1U+YEVM0lh1Fq/eeax56492j5/duJlUEoZ6o08bCKt
GqRtyQ6otyN7fjeuKbTFTmjshTP8uWefFEY2SIBL3ZsBuQnoaO4UXtuDDOBEPwLzvEOdg8TKlncN
chdpCH/Ip3EhrkFEY1WnvWsJPQgOLrwAORH+QnFYG+6VzAssZwelyCjTF4X0NeRYMJhXYC8x1i7r
eQGdb2NjFRTp+KfgTqrBl4pYOBosrGaLOsJpmzX95nVKpx8V7dmLZ4I7C6J7v6MQhYsSvA2lGXZU
dt91rj5ElWBODedxcLgBRV1ah1R942cK+lHdA1hiqgWUtiEUNxHheQtykf9HHDyc46XQWu1zZWyI
tKKYsEQGrm2UMuENrb37oXsNCEBkH5R+H6NLXijjIYVG7oa/i5Wo7PjR8nXxv/wK39eTrC+qZ3XQ
zZ5snPjL7T4qF5MeFFNn1kaiCwvcCqYbxRBZ4LVnx8lcUjY7jchzeumcTvhCD/9w0vRzim9eJjRD
mI7EQC7J1Tif7/xn6KTWal10YwMO/l+ip/W8QrnPnEvVK06pIBt5BM21MpQYh1SO4BMmMsjCz3UT
+6Dt5EnPiR4xOoVA1kyn1co0oGk5/eLbj3kV7tT6mcywFnE4bz/x7Gfk+6tSIVYpxXLJ5BvrH+pE
qU/OyZGENdKhcTWC//8USIfXUN8RQYMhP4Vfw6JAsOWWHGBedHara3PjdLbO8+sshaoHo3YbO/dR
ByMk38kItBOZc3Ts2+2XiA2tOtF4BCrcpX/qtN4h5EomrzD/YYz0J/sX6exSov1Bzj2hQ6QDbKZ6
WlJUcR/cLp4/ZsFDGA2xe9EMMtxcN6MbsZsEJvv0kbfAMsn9GZT1ztffeEfZ5Ek7gCcjo5qfDSwd
kbrf/u8jpZ/Umuc8Zhw/Xbl6mf4HLpj0mWAoAPPWvqMSEW1Ng6UDFOJFOvkR+To7s+TjsGhDRXoT
Z7D53JLMO150XBAyuDn+gTFd0d7XRy2PqSZBjqVx7iJ8whm8ld9IowtXXwrcrmFiwEvD6JSpk9L3
wXFuvqvlnPd3m9MiFqFl/uyt3gEJT+mFD9jUB+TUuISQAThdvz/gJLfteEW99kif+aDwhTwpi6cI
LZKR33LwLFgfOAPP4NCWD+fwSoTTuYmW8KT4dkXJAZQiT2e5mneZtPe8icawm8mXenbddWGYH4ns
XEvgbAg9lP83pHW/MdhrK45T1lMN2HuPHB1SV0PbcBWa8NvTNJe84J3bS+Xca3UTB0TvFocokUAy
7Cr15qjrGT90HcaIySMCPbDdxsOwNqoGc3ek2uw+O7RpzUw9NFh8NkQ3kNUDkcXf8+LMTxOeRWU1
QZAW9SPkPsR8NVnoPLfpJGBF85mPbRb+mi4YgQTEuqpHYqUGj5PJ/kUgbLZEtBlv/7VZVPlK8dYt
EhGwdsoadbTAZScCsnv/XOd+0O8vd/0R89L2sVsYgEn3ZNF9D2LGT41PqO7+qv+xX0OkX8X2Tcl1
01T4CrPVIEgFRYbLnFQdTz1oe69dG7Ls/+5f2hUkqUDI8uyZAsN4BOVDjSYhqySmuaPxaJogoXpB
ua9r5sjgsdG6kw3hZUHycPRmP1bNrqUC8/1OZH+RJQTLG2PUWL1ds9oHmdwkcKT9HakSzn+tL35v
9aYjMkUEzMxVdG90DFQG/W+af9FqudVRwl2FdP/NGYsUResvNQan5/IpRBio5kfj7ed8208fFAdW
oxS/3dzRDnL2PtZ16947hlioG67MqepzP/2VLaU9ZvwHYod4y4u0VMnLS5b4/bVPvUdXjBK+3Ck1
JqyPUKFBrMhjjoXPCic/bvR+/DpN7WXq25GIFh5XKoVpqhvpR18PWTg1QcnVwlGwJQEcJ0jTidp3
2cqW+Sd6qnW0u6SNx4xMdOptA6ZLndM4agL5pAq0CTCMFR3ejiU5O4+6T5islugaJhyFshajBneV
O0Ah1rFNV1+rCJxyd4jp26j1dF3w17D7P/7Yj4f7gYznPc1Hm+owLn6JhkinITBVF6gf3glAFw/Z
qp7bE13UEKc0EbUDvFVKLvzf4z2ZZ1U1TrLwAJeum2988EYOEjByxD4j57WHFR9A/USCn2EanOUK
tpdZtmHkVyk0ocbY0D8xalzpNz8MZbg8HblQ2GMKVykU8dJUoU2LkPhVZKh9urucS39sVQ9HJ1L4
r7GWWBfJ4iUQ8/0We3IrXEeerSy/sRQpIWdqVYFxAekXL15lA4vXmKE9jcMz+K+XxlmlY08cHl2I
q67M5FIwhVPLzsClO+djogtgCjognE8IOlztCU4Yb6fSf8gWrE7eC0rG6KF1vmUJfGbvjIRVOlVZ
I5a4Ot3AFXDrjOYBwVdwpZtXJqiB6yd6CaenXc9vT+XTtdLXj/h6WAmJSj8LbnvBW7f2JScA+FSU
dtq6aWO9GB+izdrRv09ACLl3c4Cu89HH0CQ27kcSJVl1/j+9nyr6bNi6gcTeDddqMrZmCmlZHaOn
uSHnRXbYImZzC94u52LMj03Cl6GJUnlcP7Kra+C9isOie+S0dnMAwif8MPHnJLM898duudTnYnkS
Yrw449ShBbJNu7Nc612ww4DfrfehYzY/KqPRo2gM3I4BOwBve7/EWGY8+iUk8wHnxEbod7RkrC5a
+FpXnWctkDL5FiCwgrcNtzMRCj5FnNwP+g4JzjgWZgHAd9B4Eq80sZzSnQ2E7ftJ0TM5zb4BqOe/
ZIAm+5HVujQQ+GNE9lg+IeORqq4/mBpTU7gTUkxdRNvA8XHXvZXTxs4EhTE7a6XFZtgl38iYqn9+
qqgwVXyYP94VbDT0+rU5A9bxRFlpduqPdEDqA3Y/N1UhBeXsD/AS99yBwtNwMVbD6B8VbWuaUGW8
AujxnadorST0eKGeeRkJElnMiEE9xFzuoFD3R1Ky7P/ZnX3Wz004XwP+SRAMNGv1nO+YeCe4tpcN
r+o4R9SFpL0kU3nAyh6UM/1IuoOlCOk3Krng3457M1JNCVY1B4icqSXwqNUSDa3RHiIor6oH+eDI
DBd8T0HTaclHkioT1pdpSvFC8az8UYhkS6IIiJOJ3zK4Yml7pQ3ctX9YzfbG1+OdAIQ4grRNzqVs
e03DUdgQItuj936goRUxz61ysCp+OPZNFZRhlS+xs6EpVU52rSx34l2+d48aHsDCJdt0FQwEZw1Y
tcRGegskZXPcqe9+N8XTV4JhRP6mk8k/kmtctrx3/JgUCTSl/j86olLKw/ffVOHFhAAMCS+2FZ4b
6gtjSOBqL7ufi0IajHn4M56qC5J5+szH/jeA2WifHa1Epf9bTLxvVAIPPDRzeZrF1oeurcazdwj7
cQuvDW81tanMSaZiz+/5b/nSxwfzkIuDPnJsebdo5nxQ38DaRqOUv+o/pMFq/s6u6la09XvbEYcR
WgoDX+HFB2RLv0YA2QqXXkk0G2bY3NIfrr+hEu8d15kEP2dvQyCD5te4xqwyKqZsg694E0YxiCEK
fpGfe+XsPSIQVA4iPjqQ/Yo4/P/59hEg25QIELcJdE6rsN7jErF8DuBpnpHcbDDv6HysMGK1h0iT
7Dq4V1aARwko6Dz65qQL7YZXJP1atgQVtxq4uSHkmNrC8sZMJHKiwm3Li70/GvSBWENgFSGfxoP9
DPQV4/yNyxJ5a1x3qKA8E+qMw1Fq/erBTkdmJ/wOcksNDivLsjV3rqmoHA5pusQQ1f4xNWvYHYYJ
44bRwFn36eVi/I3Lmd9kcIqgTBU1FrSWmE/KsUZpEtCqQcvjFomHn6dwqJQdMjWrlm+/9QicLki4
tHE/2wM2rz3AImhtXz8ZNkIS6ni7E7OU/bE04aK1DUstudJRg/PRIgFYcjXH5UUhx7LZK5QdP3KN
j/N0VQRtKMkSy9+9M32Sb0aSJXWZNlDoWUFeyENrS4DP5Y4VZquHwmqOdhS8WFMiwIem739r3P7r
O0WvsQmIX+iz/azm+iSNROyx0JNxKTx7WUrW0vmcMFK1bzpu7oEgZ8Ll2K6Cz4+lQBQpwGoFTLT7
+OeShBelV99UnOTz2mwQyeE6FsxbrolLw6kEQYjCznw7O7n+nSdFm9sALsXUdH3tSPAnWW4xGntK
WmT4S/Lnl8NhbOqfoyvauFVlhiccrpaTX9cGGNTlf0cnJYi6oZjJDaiKo4XrKIM/iCYY8UGJGAnm
EErOhiMW1qlctarOztkhv3hyDAjy33FG9aoXcRECIHCY1uB1csweo9Mpd81tXTXtIeweGIWJtHeI
gqP3uN9I9OfiLEhsBr/wRdDVB8ptMQc3wjijG52VJvrTgTogsNGU/3YJrwWrmx/fXQNilSB2KNTr
I12PRPhxzCQLj0SPrRmQvPHUZUxrLSJG6ggACkTngTYC7jVOYnuJwXaBy5+3bNKn76rs+O0pPbng
Svc0SECdcSX1aJ9PncPk3a5po0at8ZtRRfYrPKticuQmyFaimFRWBBPS5EqM2J5o5eRNUFMGTP9R
6Ntr8wdP5WlZAf9FLp2wGh+KZ0OjNdcwf2bzQGqzmg/gdGbvQKf+iOujVP/6EBmMhlt146di2QGU
RTJGfX/IG0hpn13+ipX4/9eicwZ9tcx9RqrEdFzNyPWkfcxyYMZr/Xlxhu+LewtspM87e3Dkx1oZ
8YreScV3ZQYp+Lb1KnCO2KQME0uOtlgWy8RKXOurnJerz23jpPKsmtMqW1V89SWyUMYdmwbL8KGY
MWY7utBg9g3D6ELWBY5Nk5Fv8tRDPztbuJ3+n3aNu17GvAmVVn3tz/PSZ3GWldvZh/d3S0krvAlK
wcSrNztzgD+yac15/xbDU6pMk0633laxYXG60F26ytMr8o+xBll1mRwZzCCiviFwtWjDEazRYySi
vOIe1Z+mMJAdAaTpzKj8pRgEMBrUXK+wHOOMYAoTccwsbqT5CLkmVcsnqOdZpu0Mb6Lc4/MfqrYw
/TfnRKWBvcVn9dugeYZoKIotgrtPMPe1eBvIKXvKyEVyv8gN48E956954Qa9zbyX+xjkqNF5KJiD
infws2/1NnEu9Lz3A3nntgGSPOYdNnjAahbjnJ0t9ByF+loSwHCqWg4bkauPfeu6hYZa9ZjHgq6S
6j4FdygfoLSa3PMf4HcrV00groos2IRjqYliH3+ylhVH1Jy/RrRq5mt3hcIhVzWaGmBjZjGy9Ofj
6tjeBTKMFN8wv+ZMCYUqXObqqj5Q4+jhTs7FHtXVuEvoS86gdS3rQrvmJvfJTe7Vdyc37x5qw79y
2nDAcZsrdho6odLfafIRpKBv04ppf+7Lo8my5O3W7rG5TrC9JKuP11PvyARMv88AQRqlO/r8A2rS
ACvc77Q1h9KkjUqSLx2HMNmEibMdDfIHkJBKHLI8mmK7LMUlKYcE64BeLT0X+7UfHUyPGipMXJ2d
4B5AglbQQh9hmSGTJcqtAV9LYukFXK7yXJs194ejhiShOzJUi17T/qzG/i4FBp4TKf/mBgBg4Wd7
su9aCTOQHHcBsdeJe7pUXBwBdaG7Vk+iWGlpA+lPaSFM3XdXuYK6FotBNHNE9vu6/fCoW04M7uvN
AjuaCdUvcuxx1iD9ziJZT58CYS8FW+MKKBOqeK6JjwV2eXxNSah60Xa/2LnkBpUgDLKmrj8GHcA5
quWmow8zhQ2YsGCahd7gXy32Aa4xqQ/ia2QiWjNuDDkQHcn6hY73HwTSjx67bbx3ESjivo8kVNZ6
rSXEtpFnQ5GOiJ8rtoE2ShvcKSlNAuyGL79l2imEFM6eGioFl/Q71iovugFLydkQgHi+evFKpKQv
7dPC+J+pdW8/5IW+nI1wFn4QImHptYc7xZHi428lFyTjaYlKgJ9434LtbTtIqr2J5hq2nUcAlUbO
3+UtUAbZ2aiYexQNCT5fN3sN9KtrjLui2bB4XDBYe8oEp1l1VOv0L8WJRDuS79J4VeT48taMYxkC
L0C8eQcPbQZS9/mjfsNRMEw9XW6jofPnLdQbK5cD+PmJEG/cq9Hy7fMObqPvEGKG6LNcLK34oGwn
uiEsEM0HWL9kNYMIlsN5HjiRxNWkzhhLtJ2LJ40WTJUF4t918cpT9ZiqmD88PrmsUVkxHghESR5V
AQzEAVhLaffNpaK/771IDJWR31dBfc7wRvq/otb9T4TE3tyHsKUI7WQwylXjJmzrIVh4UE3WkMqA
fezIcETJ3nELCYWasHCzpWULLtXVNCkIWPb+BDO+bdrmchhSE2dTejRU9sxIknmYCC2YXBxvo4b+
LTByGbQwRsMeO24tg0b4s5JXOqiPRB0owdKy76smTUm3DX7KssDSon2zC0C+0CK1JA/FI5WTAbcS
xwgZbAxldztIEwzWyu3nku+7+9+EBI9eRn1w/8iLofkjyrNGWvCUGZ6H85VzH5o9tPCrgaG18dOs
umXi9tQmPMznSkKm7b1naeSyo9mju3umGj3jO+llPhRXl5nt3RS3FtO6vzPRuLHpYOtAKynTbkDk
aBvrobSO7lUwKNsj4qpg/Mk64Ci3b49P6BAPnOrMW5SLjsgsWzZQEfAOfgVlQQqUBneMmoc66ZgZ
vpKsklnuBvLDs0NoehaMKRJdbzebYtG5WxA6boonerw72GshRMb2snmxaVr0BMyRMIswxamCcY2X
fuYLS+i819/nOZt6/7RjflDrPhctNALdDaYmfR14/eCzVLY2h0zkZcEqyfio2tMziqfBgRABeLiW
vAIgdUx12H/KiZOHQuoaoqrI1r8/XxsPn9lykDzRbMUUEFCmDnLcHSTWz2BFW1AvIUZeFqXnhVvL
B+FXxzzcaq0Ft4FNZTEA0fx80dnf/BV+SdnjJ5g/ZduOj9dLp5c8XaCHRAxuyIRSADwJfFY27eqb
IgmzOjJPpPojmVnW8k7bueVR4UbOB62v6zkcrcf/7Qf0VnzlQ0EfoVtgl/nFqEZU68FYohYXLwAL
ktVc5kOLRChdPrnCwi9B5U2lvUDAtN/K0pE4NCGV7zXkfzy9o3KOxB1CYbA55Dfa3b8Ge5Q5Cbv2
WsLRVTfZBlPV3sxqcNJcbHnsWtDZBU6vR8NA+1PfZ7BmXIstqhWe9wvboOcTBMtwlQPnyvAkwUSU
WLR7QYRu6d5eqt0loDzbkvNRW/9wESaLn7tfyieYZTYnVQHgpo32pah4KqLS2vUWfzHzx8q9i3uG
yYZTd1XORDpJULK8eOXQIsuZJBdWF1+PCfb0Br9Qw96ZejeJc9mU6Xx+x+FH8bToI5JIFIFhyfq6
h4hvPwshdRexs9Ut3MSKJH2yrxjMh12MYO0Nte3ueOeZtyV9hMjpdKJU+qvs/6J6c4Dx2ncXcVyz
AFmW5Xq+7ogRR3/tHgvsApZ1r382V9CC2laRyg/+lPTUNR7SLRj6q9nSs/C53oPNrBWcBkL6MW4V
EJe7RQq1AHkgbaS3v+niCLOvoOV3qLRvRwuLkuMNLu8PowpkoH23IWkIH37zfQhrjd0PjhrmXP/g
mf+/oJsyTs4MmPg2Q9/yUsf0Zntt8ZDSWaA+eGTpcewEIY1pvW61lXcPqGK3BwwS+e5RJ6u0d80/
/P7MVyHq4jJk+HCX8YUj85BJX7aFv8HZa8MlN7aZ0qAjKUD1Z5ZEG1Ac3/eb7Nig+92FZuswZwRA
NVa1c6ZtBlK+ppE4jQNoFgxPCHznsQqWYQRD0cbhvPzUjt9yxyHOg1u2vaB6SrBx6/GKrpp4eY4j
qR7bvoRbnvbQ36m0uVg197UOPcYSCS6SlFDIZ6IoIoDCftue6uRod1P0fUc8kpPjZiY8I80pZYGH
+5YYsyUJ9epkAsocOXKqckVO7rFW3fThMyLUazubEBsvIi0WsOyK7ODA+5lYqrI7RduKtJe1RbRo
YizshbM2B3TAxbbLx+BMWANFvcYRgfH3vo2R+xbpUJ0JCn6pkBEKkBGv5x9mNa/gfv9adfjKT1eP
PO7+d7eRlSXqGc02sB8kNh6DVvOPKRXR0f8Vr8a3WpNgOSBYp1femHzGM1oRnYiEb5smIduPxVZu
o2uzo5zofPDQ1kdpv8Gbs45YXLVWUcr2KEPf84BdPoMhlblBfBhSIgACaXmsb+8aVSvLjcauadLj
QvfPCfr5uOHMtYEGhK9XKfiPh7UmA0K4pzrpjkgYjOaixzb8x9oHehE0Y9y2C9R3s+IGo/Tl2+FT
ejXSYAYuNZD+vPbvaHF4jYTqTz2jIKkD5MNwgnwWG53x6NpxOCWnrZ4W081uZcc6MFCnxp02jpyZ
MfsVrePgfdlLLEwdGISU5T6q0aqa1/hw4ectKTCr3jnGu2kUOp0GjzjEbmkIEVU1/jS0gYtt1UCV
WbcHw27T3OBc04Cfv6jll4vMla9hmguSXl1cBmyX5AJE6h7mi8br3mIk1wYdvtWuGyUSBFXb0nAh
kgpSXIa2NDDljz/SlUS9wgirVpa95fVdHezUEtt9AC0krxaQWvzYjAzkW+QLaBRssKnLG5wYOmws
+GpfGLk49dhzFqZHHgjP6a2K9qybY+gErEVcqy2g2RqHFYDK5cl2GjhAlyhxwaQvpF7/HdBW0IU3
+cBTaU0FnHPeUXcVbEbvz1AlxT/7oC+PdywH8bBEyBl6zPKlxAN0yZL0Nu+79wOkCue8EPvKqgr3
tJofp1O8AWU8+DEjAeuNvEFpeHJJ7VMVZOCvKYQqrb7wGk4qdCRCm8vvtL/0/if6Ll3cgpO7jLuw
7lSjy5Yjh/sLsvdVRVF7Ip9SqceuNAmrJ/X9ykektKto1h/WrfRS7J01vwdrf4OG557JsFhTBUMF
iUfAGlzwXeY8Z7Ay4wKwUwIXcTqtPb7H5pro6dfnu85KqkKCw8injPHqVK9InmbVefWmqR+r0++n
ssZX9Hwj+vEGoAgJznMjhlW+yRHMhIAEJ6Mp4i8fhuKpSICE7WtK0POdps5IxsCZopwcvoDOsv2A
L9oGNF3m5U0S2zBTw5qWcM/sIUh7Fy+f2SxfJSdLjDPSKbfnIimqXaVbP9vf4r9/ZSHtojFXtztl
0CZKR1jyynz8xzWOfmxC0CHitO8natb6ynONgUTIEzYAmMdYcnCXKRBxo9rwNeN6mP5EvsF0DigA
CRJElSMPgh99Vg+DgBVMLrAGDnVptBArxpDJ6Y4js+X6y0NFLGAorC4q4sxFyYCmz6GPz/tFOaif
faq7WwI3wt6qJmat9ZAfvy3ta6zQ/E8eX6fhSbZPN313wrlmBJWEsXFbQs8aKAI45d4c3P0Bmjnc
R/YOx2ggLFuyN8tREpOWpruTFh3DuIdEds3Kyqhpn0Z42rgsSRaSwNZlXHebzvl682++Ox2uBR6x
+YXsO4w5OmqtxFhBFUm46XfTU5/9RLcmzSemwC6yi/qHwAnpH2hO9oJHFoSQ4WRVxJ57xZ5Gdct/
dQhXuRSXe9f+SsikVaTiErWWS3RjCBCDJgc/l4BqXYj7aWc3ebgN0rIW9xqIEZw0Dykqx7ZAKN9R
S7utUjvlHS42CrJb2GDBovE9HS4DX+0QHOvCo9Nhq2kir/ZLlkggYfk9HbdiSBGA/ml6buuMIeYe
IczZDJtLmqlJXODB/jPSSegKaeX1LzAa3MRpp6L9bdrg9zOrP5Rt+vfXHupg+5JoWoJFY+VHZb/b
c+TvLWHQHQKzmXtM2betutp+BrKLnFjd0H4tmidYCgec8617BJdb7DorTvzkjNzKJpEXb7x1Shht
V5gUsGAE+yvyyfq5L6gYHo7NAgxpX880VLonsKb/5ZKbMDUGrY9pQ44ouIO2keQ3iQkzYRNn8i8Q
r4HWVGNUSoRB+QqpMLd7oDZGswZMU6be2JaUqHZ+sO303W852HnKovWcwGnjz7dhrH34wyLIwfi5
MN1MP4yHe7gJLAq3LDhOvDWmknihdR0veEB81WJdvU2W8JP2IT3w6kJE93YzrZLfrxDK5oiVeQsl
9agz8lL8LTOpCY4jtQan4cwY3MiBZjXK+LimgsdsqgRHEQLNDUgTywN+64f0HON1edSFcBvHIKka
IDbiNNwxt2UOzpYQoffZmGn3VUK+1ilgCGZ+hTidBc2HRqNWzAv09+fVtRGLhORFpmCGrYmST9ju
WdA3J/V2mR6Q0UsKAHCujVJzfZaZpgmlDaEbUSAxXwJEll3nkrLxZTQH6He/T8N1yQB0v/L7BZH8
XhgXezzB2RCGfkFsTf5OPfLOFoh0BUj7xu4+S9T2sRB+MvnQkc43lQJUjt2IW2DaYF0XHPbWhswn
Ed4YsEIn0abTWTnhPsMrpL3NzKEz/7dBWCyjf7F8yLFrHPKPkr+lM/XIvGCOLt143DcfP1A2iMTr
jXfpzFMCw429aaOTMeY6gAawAyR7298PfUWTgvC9s4sPqxYfQpYdu+O2jqv4aY8atL07cxKAFkhZ
5MvveTITd610m5ghK4gerhDQxLvXDn5FmRpNZS5ST6YPe+BYK9KuJ+IEDtJId6O334i45kljaHg2
cOiGa5cHuSIQZ1F8t9lIQGv8BVfjCp5TxwZlvt92fzZqbtjsSDmYIh8UzQWLWpyJitaLcYEkmQxm
7k0Sst8zowTysP8hoebWEdIoKv02Umi7MAgKiCl2XkN8udTjr0S+QeitAGhuhVsB87QomOLmJxmY
/ZuuA0NWnOS04Ie5iZuUBxubJd53wVYimrbaUPAfBw9Wj073tsmmV3gxEDREnw9XZL1kI99Y3+7q
ga87TmAwGj5jGlFomLQwmmQ0pGSHJrzQzU6HlPrhn3tc/O28/TUA355rSyAQJcBYCYS50674Hah5
6jvv4NnVzpoHK4XsjKEWIYC/p7Oo0+fuVZSc3Jc3jt8FVVL2KXPn1+UyhwUXmeRfEuNQpn/jAqv0
a5VZvhTAP1ee+fTSLuCQaxdgAmNFR8Yn/zWkDTJEONkrJfQTw7qTxnTfXbzPScwZdKqDMrbt5opi
dnsfmm+uZixUbGT5+bmzDAPXNuEXKTo6EpGHhgvS5RguPNVWyq38qFCyscZfeCE+XyZyAoW74mKH
l3JRNi10qWrEErL4B1JO2mOjsz4eyhHe7icwcC8l79TwrNbpZmS7+PYmySNQXC2lMheyZ0tV2zRS
GNV5KGTFD21uClW3rm9Gu+vz6ZGg8uBpRf5nD1WKuPmsdOJqiGfbwuMU40Ih35MlXX0AE+xa1Hws
Narknbgw8u6/YTSQOUSbObYz9Of4ZRfaGs5s/wJs+xvbxB8/WNBCmKqdja4U62KD1rD6u313DV6p
eIS5fwrFqOJvSa+VLbw1/Zsj2NgGSrL+eeIYvvMA37c3M/X5RephrLsAUlKejTBCxhhxCSyHOmEl
3/AQWyaaYsunHAJfeUjK2MW7tciECbG4zmeknTv+ymrPrgnB8DbFexaQYA20jAehVGK8PWa9QUTC
jKojVffy2Gus4FRIRa2Z5og5FDURsxTMyT8ThSBE+1Qr2Xs+HEgcgaD9J8szQmCgT8plDI7gq0bK
vy1p35J0vZ9AmQ48JhQpni25ffDZsojTyUa2KfBJT3cx9KHwo1jpy5SU8DsZer5URu+bhFoRm1cN
wRJp+o7hECJmq1gmoWOSI7jJdWtJYy+UGodA02t2xBzP0a4tsp3qlrIfozAgOaJXYl3O5GrtW5M/
uKTnujnuJzsUiKCSSCB2lw56PHiP9DujmlqEe9If2uu9m9iHxxSjfouTtGI4XvvFXcpM1BS1lPgs
lY5w/o8+ne+ENnuDcPKiUnxuYCZjuI/TomYJNwb86MKYbADCZfHzv8Y/sVZ1h+CjyX7zcBnuMtlZ
RYKjvIEApT/4aZb1Lw84uYQg+RY6m2AMarev2VMiNf41L6eIy6zKb1fBc1IOIpri7zPtSj78GTY9
OdL3zu5ZeIJsfn3g9omVZHd+0KMFhfPeRt9EI3iYm89/qwOBb5famoKE+T1ZiX3/j34ZN/TrmRN/
Ktoh+J1NKmmjLqdbMUsc3QyG+gVXR4PhBpi1hwiuvPnFGfEdLSPxasKyT2yFk5HopOodB5hgpA6w
NLSjR0cOkxAXOlLzNUYyDIprp/St1XKMzjiAMIad7IXTAfpbTKkFP2W06BpGE7xkt1nDuDzfoNa1
WKKLVafq5w6nKAlXoT4DviGIYpgAPgtNXbxxJYrXEcKVZZTMsovFElXcGIHjlC2nYtyK+gCa91rV
TvOFlqRZ9H2j4H6lPKTLbrmVTPP7jES60TMoCdfTUweB7+9a0CAzlTG93HcfGbjSj0X3K49gUxMN
2IxknzaNTSg+r6ARk24hY+Qk6mFWiBRD/y3kZZligMJLjZoJfyTKnR1e1T8fYiuLFsFzEiSFx21n
XOs5Zz4iwBooO8hvfjAgxnVCcUGTwYkOj2goI3eoLdiv5UbIFabVyAVTESZsiFH9X/IQw5iWG1cc
rQtQbB4M/kKZyDrpYRuZZRY7ROjFJ9sB2A08t+YIX62GcQzCu+pZ1hPRtPCRU0dLfl1eoaNEpHO8
cItYFZrh7Pq5llwXzAsA/b3fXd+fRdTBw5pdCKtsOOdOiaBJawlW7iQ7ivkGaurpZHNPLPsqe+sK
gj00BvrJLQSFDwJBLjMzePeJX8giK8lDvCHNZQ7GIWHzRXDaxJqCqNPSTLEQ0CaVGP0SSwAxAb5B
Z91OBNjfzFMp4JNo5sUrJYXqlB1y71wN1bQvmqU9LoVjfrwYr/CR1wRYp8xp771EqAnsSoi4tJgQ
xhg9rohgu2kfXHxdj406T2rh/EAkl+0DkOCeXvvRO0fF9s0gM/JxW7BVngGNGFg1NKC1RYxfdwnx
syBxjaQs34oK6i1UXS97kl7PY8GS5ZwQLGzlFY94qD+GxxOy9E2Vv2xK/NS4C969omIDo6bCPF/m
b/mPe6n7y9o2SaH9jnaH/MANHHuityRti1UvOfd5fMl3Kc61UkPCtbL1WfTPjLlb9kQxZQ2dKH42
JgeZMmE/zBBLBu8xhnH+YC6kuuwB4yWaB/d32rpyuHEw9zj25Uwbuh2MoiAr8OvWhXu7nc4q1hjv
5jjyBxpIddv1zM/8ek9jPbjOw0zojTt5qGgyVXFx5hmnWkR3tKvOvz+FmjoNaVR0AmgwrlSz60wS
FT9uY0uG5/vh2iWL4R5eC4hP4a6XHUl4WmmD8x0mXQvcF+Hnxih9SUsH9Wkqhxgqgt87dlfD3+xe
zL8yWuCqPyWWDvTYS9GTha9F2Xdo5CkHcGBRydhvW8C24hlUPko/jU/HDvxoYencn7ae9nrjs+hB
55mLDpdI/X0luvS+U7M5Eg9pDL7rSp4JikrCgYVFMNYdENpKlQHMviuOCsd0KjGBZ49kfryzB0IE
e8+n4tHrA/a71vvXjhNajG1vrEzZY/GL7apmwdYqF8thOo5+7EoH1HVWmR9KY1ho4jruoCs4FG8R
thWFp3VReLo7BuATXFNlt1X91My88Bj8WLShQ1YzFwTa7O/E9B4lemouDbVx4vpJvcL91D2AqMST
ELAwCuTK7O3I7dSQMQZFIZCi5/P8BDL4vNwR59YRdK8WjlH1xBqmpUZCjuKtIU9tyBvNUp5Whi8k
8+M3q9PZAr+DxOOrDmWQrUeKpe+ij96BVYt5uw3BfRmWq78Y4YJs2CpFB197SJmCANp2jMvCXsN3
x6ZkdbJpmQfu7mbz+INwDKF461Wt/aE0/6zPVzkDHOjqvpomEafKj8hjBc3/hkHNaMVDQ687lOmd
yA26xybfkITlD75Z5JO3r1T/FriS8Q8fa4Ohz8uXUfYzWGExPzE1BRsatRglEd7VFEg9O1xPzbjR
jVQWTZcp6r7BMAZ5g62vM0bVYTMI+XLOcEKNuTFkjXZxP4A1NbJdlmRcIk9QkGvLg/ELNweNSfiT
szNA1bCSQ+3waFvIrUGir68hiPl7zfiX/+T2ieu7Et7wSvLuK9SjEtXsz7+1QjANa+KnEsbqmRmZ
Q6F+KR7I5hgzNCm9IQb1rVIxn3Unc3h9eUeINQK+jNL1MOnR/c/oHKGw7QYrMtZ1lW9LBhAnwDpo
wtRLbSOuABnvF/ER81xJQ2Pgpn1Rd1iQq3arKu7qfzE2uT/rP+KEM7uarSHR20VWklzQtWEbsQHC
ojikwTNFmRtUXTQ5LTgauUSEwIyPCUr237EzVhBS4YG+jn5Td/nC9VEauHxY6UkZ6cr9ryEVMyRl
Mtpf0qDc+yQduMkBXJjqq4AwFlCiZYVs/BQVHpe435Z31pexKvhopPRngWdpwSolQUbFtASKUhmQ
TmIIrS1iWiLDtdz6OTJzuUgq1VyiBihf/IWADwF+JHImJssctUe0QsK+VWxxwFdg0FUatkzO8xO5
uu6DoELuRqWgeIB6qgm+SiqJ1lygG4unxquMGMXhftx/r/LvgCC6hdr9vTMwq640uSaiVvsn5JUE
yjY1eZAXs0+65O9dVQIh1z+boSc70pNtPOfDzRHvGsRoqrVC7zzPet693ZxcKN8qh0Nhe+M4C4Vt
kMFV0sZSPffBKBTOu6Igcu9XWQeu74KvKY1AqkqpQUJXXfePDIT6jHmKkqYTfEnHJTRr4QJTZ6k3
tWTazO8O4NwpzLmFaQg1tFN3cPeejzK2/8Qzi6hM9T3v3V5/oikbce1C+Bkh+an1SGa5GgRtVO3x
P0MkIJg68RBsMDe0szol+fHWRMniNVkp4JFyBmqetsjOc8rDEuCHMR8sm98CQPOqBiL/oMBpqf63
Rcuz33ztTYZ0DG6Ftim5cYw3ScrOwBytvjiOmz3RG9qfKZDHnPxEVeWvbeaVHiS/sh0tIeb4N2n5
Njn80Meh6acXBhBsL7/JQnfiRzMEJ0dzAgowBJIS5anhiz6oUGn7IaDkHEPvKH6fcgFl9zAj0pKT
Z1rp+qHoYXHeUBNUSNfyL0RRNCwrsOZHrKaILcyxz80YuqFuw+L2TnviMPC+YrriamC3kOZ22MNo
lJnnrH2scLyA3opUh6n+3uHJgxzHcuaaBXt2IkNZr5tA4Pq09S4mGRp2MZlO4RlDwylbeFrF9unz
UwEJqFLw6C2l7OV+kgrBHFosyyoKRNBj3jDGjJC0KY7sAi6usDFvuYzjqO9kK4aRV5qIkMVkVINq
S9NEJ2hKdMoHUE3p+2bqc2W92tP6p1UHFGb5MSscKjPUIDFajs2/NOzBt7IKGoqT2a3II86y97W2
kdHx5G0A1sSgigyu9KxefgfKUzLzjPUa9gEwco4NHQK9D6WVQo5chAMvC5lVMOigJ462FB30C3FI
vbJfbqPYT8Br7Ct3U7ivFw+TqYmbt4LykN9uev89HGYsdsRAUoIzUG7DaC49hRp+qSLnosV/8yeW
bGh3Qsz5ebX5T3apFZDXwNVfxkfEgY59UGhVOukW+G45n/80SzRGqnrEC5jftEhsGWXGhXWijBVt
gnSZCR6VXwJ7EhCHLVIBR32q/VNhjow+MdESDZf4+Wht+WFh2aLDfS+CJITNPgI+YEG9qynxmQxl
CufroSesXfxabvAvo0wR6MxPwJ8iHQy/xttJsJclvGa28+utNOxe4BeYIR+71GyZ72HLRT9buttw
awY7jkA7/vM0fZgLAsp7IOMVmIoYAbbOi5teN/RgmU6slyCQIlML8w6owejLFfTN0f8PXiHORbBn
h7G3c9c3QSXyuwZAxQTqViFY/p+mWUcVdsFucQuHI+ss0CxSX0HRXIe6iswV7VIJY9ZkEyqgTCw+
Rtm3ZauzBbs+jZbJsuxj/fR2kr4KZ2SlxtclgLVdumLOpcnp6jXRM3YJ7co4R4KMClWZu6yJCuma
fWOgY1lMhKsPQz2Dqp5V/IuDxED0LeImcO8Vd645OXXwUP9rhVaifScUe4tHFD3UrhWS6nxsDLjl
6GBedBNR6zBoLim7SlqcQRhSrFTIJE8tg9qzXzlsuDvTH3LqCocb3rjNzuxlGlzP/ZQs4a6i1e81
LMcwteXJhW4a4uuT0WPBQt8S0CACUuxXcq0ayMynTxY4t5Fthrk/yTeyYDjcWtaprRcuBWX7/SW2
RVUefCsbahoM/lpn1o1qknC7Pd5/y70RaSdu9CBUJmuqYXKbd/tjypQe7dgLrqcWfIFFh/RX+e3L
81ID+GJJR2iw7mCoJh8ltkDfzfPhXxBH18UWI+TKdFwXOAlqCCASggKMAYZzrkbFLHE88UD/v6Pm
MhggUTr4qFsIKTfWZ7Zlv7wrirtvqQL8RQPv0OCkUWCqhgn6jbsgJcUdt2aCdU5/BhvJBsUOBe7f
NZ32rQ54bLKjFxgJC9IrgrkTuk/QQ8AF2ifY1JnMULFjIyq3sCQUprTZ9Y3tL9aZFXefw8qNC81o
V67KIWMocbOS+csQaJvzs7B21Rf/MWpBkrFwQhw/DRr+C9IylzBStvkAhJlsrUQyhwTb7QO/aJ97
wRHqegg8PmsmcbdjLUbu+jRKOyk5Fs0Yu9f2gY6jBjigh5qPp/+EMhK8JiMUPnd4ksI9VEs/AZN2
a96Z1iFprRkl7gnXIITXcL7lPaqIFvY9rNc+pVOfDTs/EAiq5hsO0AsF/kCKUh/V8OHNg8Z8JG31
p/o6lF0+kn2+oywA5U6PmvR96jva3Hxe3ci8aeCr4GBk7SjuYMYuPGrq4LyWSg5HVfCZxeTlsK+y
f2KIXvC2ML8NIhvl8G+IxSIrxE0sOjtJBhEnvztGh+f5YIiDwfWqEhAosqR/ofDugvVrDL6VcpbH
rg2XUvVv+PWo6w548unJauxuTjZ/5xw47xDeeHG3apGK1weUaD0ZfH5iDpYg/yknTTeyd250+UVr
/SUVjyarwNeiOtstHEL3ONnS5puibcHdqNugAnJNIm1BdKgmqyiAqywkyXUk+gP2CvM/e6ow26zj
ijdtww9kYTAMP8taSZ5hB+kSpvw4qck2GHSEawA9MXJCLqffRfQkOhalC8uAMnznJnNguQ16Hc0V
v4ynnConH5kAFRjUzwfRAnJw/X/zt9b76Zn22lhZoUK68xeNZkC1yQQKn97BRu9BRaADzvIRHofv
m+ksp/hVF5926xw2cN5SAd68qlz5QRa1GWOHtv53gOETI5wkdK+W+34KcEEcZmGp6JomKRbksJCP
DNwfXoMp1D5GQ1YTexOVgC2hTCav01nne6Ld/nAoXcdvrGWfzHJhNAdsOZDDL992nDkKUsqj7TXY
t/D60C9zfuNEJtgTA6KzlNx9gd7Cq0AD08CTpPwvwtv+kSTV1DqEGmt+LVYrAUQ/SfB9fN2GtiD8
nmNvdBGuIwxoFeVT13PghePPqYI0PjkBJ/16/2SQywCqt8N1m/7C2hkzJSZ6F01P8C4DBfYr/ML1
U8lYU6YdbqmFbetejcyqCSdzFdqGwKugf8t+XCENN6vKrvchO3GQOfI/WtN8Xp7pvwK/qq+YdVGn
Zy70G83YLQ3Zx4529I/iMIolfv72GzUzasP0FkhVqvqre2ekgcf0V1ddzN63fJhXjPhCooS7NVdo
ccEhYSZw2alUi99IBhWmmqIif0tyazJpOpXKgT066xn0ebxez/iUlFIwIVE0pnEgY4Wfzyf+05HO
DVnqKeluH6zCHATL0E6UHW+a8WblKJylnQktiBM2gDlsnP3wpu11aB5FEd+ZD6cYWGjITC4W1MDo
gnv07UtPv5qpOIa2vK1HXDbe8TGPJT/4W9YVRVAIz8PdE7hubEFJbswBExweS/RFs8xUbtPPSwRq
nsusf+XgzzjOtuYmOLY3qbKt7LqxKIKMStO55AfdpEYaL/Ce2y51sYcpJpDcbj/1tZDtpSucTT2w
XTmuxhM41sEY3QddqL3BBYXjZW3R4ah1Mo6Yqn8dKZDFXSooDJuxv+c+Ls78nnJUl2mAfsPq6cVO
8SHIjBiejNsmkDBxMOc1hK4xbcpeLkSHbugzYIsmST7K8x9tOwICfrioyr24EInx+P7ft/uQ2ZeO
7FXLGOZlqP7InMa4X9DteUKw7CCXQMUlYqsoeP7ZIcfpN2IzDDbkacTFb0S2Y9RugMFasmVSCpDS
P8XNdtzKJVizQ3BzOS3GB6NWCb6YeoD+9Fl24OyOVofK7m4zeTgTjLkaPaBLvDxe/22sY6Yt/B36
HiQAZJH8ntveWtAVCpYmcSH/Ahka7QYW8t2nKG4AMyiIQF/NAFkQA49/GSKcrcLlh1xzIGXMXr3d
3DnZrdAjZsbbWaAf7MNr+szsZxAkK4w8pm8VOg1wubUTqYizTgaDzdDllGVp9hRQ9uAfpCssZPka
yjyud5ES9MnTRqfsxYpkMc+xUCdJXE0TPo4ZONwlQ9XlPw6NYyQs3UVBBCott7tY7d5TtUtZA9sK
YLwyLBNzXpdtqtyMB1aOzSqx3DkLOT+d4WC691zXL3hAMTJxQcrcCDiT0U8o/2TFGz/FwbAe1tNE
atnirupzms81zyZPJpk8jyrKcJmpk7Ls61ic1NY3WSkCKp8oik+OGm4vUW406kpb0nrd5jI2wu/P
V1l+ARnNso5UI+QSkRz82Si4lugphmGlpt+DtWvbkxUNTu200DSlu6yArzvcZ3/xAfN01tlHtdm8
ofMCo2luTthkm72iNFb5C9keRcqFemk/aNyf/fsSTqpUdxO+ej2suztFE81oLVHLL7pERndSIFKI
W7DGaSo365v0uSPvZ2LJypAI3nuRMm/m2prnQng4a1rxJvE+3QvLp0OV1F41Sjra25vncM4zxV1C
BybU3JgHlmG55F8ZjC8ceR3/fBZSf9RL4Zyz2DOgSkYuk0R7oWGXZc8vhTmN/44CoDMG/R24yHst
IzkBrUq1JjkS4d309Tq3KzrTJv36q00qWWkMnHyvE+9tBQhCnyOjZ9dEREWJXLjJBSc8JY+GvqZa
hofYW7Kr7Y6s1cTx+G1nw7e8GO24FyDxUj1tGsNiMHOM1VluMGkDAMejCJXzTUiKnBL89h6VeBAw
cK50YmpCjK7b/utsYr9xN0j72LD/8XvCQCKEKXeFoAgeo0dIPJuxO0O4KdDuCqLMho99mcEwnWyD
NzCMqk1AUCffm+tKNBIcW3RyhmUgWr53TrbCPrZJGZlXfZRtrhKLxs1YbhXDZqv7ht8+6jmTVhI6
IA3fu/zflCtMXHaiCuJvb8irbqtSa/4kPyxjMyDAz51+BjUtM0CipKX3fLv9FJGcevNvunPyHZPR
EnCOTHs5GT3rOt8C9813gpNtDADGAt3+VvzTBi9Kn53O6FnR1WrmLd+0n6vInR3svSlipylVr6ez
Bi0mVJK30YBwN8ftqJQ7hy6zZwzI0GfRiwoKWsaUxQhBc8Nj6x4/OLMYYD7pwzLUN8wC8eGrCRSK
RGFnIdWCesJW82CEX6+6BxAqVoTHPipTujxHlmfqzH2ChxP27M4b0hu3I2AJdg/eSETAD5zpg6KP
585ioNIhWhqHL3Ld/dO0UYm8M/XsxkZfP9C1iCDAhJndRFHnsbwqhaiQ1vYTax0KRB0VJJkMgAVM
bcwCSWQgRrSShpfebY/nUfqhXsfBoDvknxZiFIVJC5FhUkVDj74wj7NKzDxM/qvkRWDtjUjy6qQu
+qfMKmTdYY0euWfWJ15cnYkLjTpt+QsR2LJonFYm1YOyno/u1LEIE/xOYfOUttFwJhuNst74+gdc
kgDL6e1fjEI2+Y/n0U+KPkBWo6gqlvttbDnDKBdRjo0fWE59vwRPtZXKXDIslaJ5C5JRXwOoLFFo
KtRg8mTkpWMr3D5CmJfWo/ONub8TfboVTHI1WTKqv5MMjcTxOKKjTQafT1eW/i2P0mqZDOSp23ZQ
V1zoKUz8UiDXaVeKO73xDanJDsr0DvqQFNLUIfbyYtg+VOWi283gXgca2nsm4Kp+hosV2AKrmK5a
XAEVlKmjvch+Mhkg3mTaiHtyotx6YPXgtj4ivqJU+Lw9iS9EE0/lmvhi27OIEzag1Mk8Mj1F/pCx
wgcr8oMtHJH5fRXvcDM/9cZFIuop8+Pv2jIJEDctRQHQQYBREyvNHBzEWoZugiMtN6vsclDWsQPS
IPRzuLrzs3ajyX88z/ccLZfTGLV/Met9jlQiyVv7FQbhzaQfQSdA7sZBN+Ar7zgtjE8nwrNTQ1wo
QjSKQLAMIdIMfrQeh3rjJ4bhCENKARnnQXYCO20RY35sltJwYtNlmDMGN/fd6zT7JsLMSwUTtXLg
oLJTDJP1ZBsoDyYAh0TuSpjhUEBvN1/rBx0G5VMjYRv6t6o7lLkXdrxn3X0LyEACJLBKGDTrjeGl
7a7VQEMM5TL3q0fwynKyftN4FrPMY6wgwqNrM1f8JoehCZlOMzbzB5DNKwLgCK7AwExzovJukA/g
/xNxE6LHNqpFL0jqmNwsdBZdQiEEklJKpA+qG/2NIwwUJ5xggXp1VmpG8xEvOb6V8Eano0HStP11
mRV0PjUKHG/Nmf9iwEOOgM6GT6TBLk2++gLJyHOrmmrmrVdZPeMCSMVfW5XuwKX8V15eFPsaMmZm
Yj3cW1seL1N11C7GYSUOsw894ZheMu5T5qtxUauXhrxQ1V2Z5ucBCjWR6zdDhlovtd4ENVzKd/Y5
WE8bvaayXe1c9cxTGxVWqhkaosmQFErgUtnFP8zrBZkWJhr60KsXWxD0wWgREKiEBhyPp/Axqbt9
yOQh521L1InAh0TVyqjEUO5a7DuamUhSR3B6ibhXFiU3nUuqMDwHO43WblrQMLnlvmeOUUvt907I
yMl+R/gQKf/MtcMEp7Cp7OkXIo1XjfCeh1FRhqXfBaX9wKIhaKrimppRZ7VBalIPvlNxqLzVNCgm
8ljqCMt3TRbVIvI54pHpbou3YtobYNNJRCc5dWpG4TsAY7QLvHZhJd5APSxzEZWQUJxNSbT73xlj
tUDktQajHWFjQ9M0NKRDoqqJ1FLuw37Ol1YTEIOSueyFfsNbSuP0V9ZnwiHA/G1JZLo4Orz70oBl
irnXseEDYKrZigBVnjWusXfDXmgRqS1memKIhwLts2JvH6l8B4Y55BUS5TBO8mL6W2yXkJZl+bNw
S/p2ofISCuh1jxWwWTywbbcXCJHvJjjpwFiG3ETWdvg4GC3bVRvRNYGEdvzdD7GaQeFDQYL2yIEa
gpCBn3vjzFWNbWaUvc/G6xlIsJa+3KWM/dxE9z/QhnublNUtQalVOptHVeFatlStr3fBttAR2+ek
NyMzSW5MSKP/UfsMjLg+s4wrgOJNVfNwpeeT73zyoeEM1p1I/UiFk5eONZdEUWkf30+7E4VSL41t
HkT6TGAFBfBbsTAGhZK9xCoigCJHJBC9MlcxYcxXWI8xmbr95qgCQxWlnSj+cpdCZ6jfBQ7xXK9e
/PzTLtPqkiOyYDyVMgMAGXGn9VBSFC1g3+HnqVaNBvBx2oaN6Jtjjg2ppUzZ5RR2R5E4mh4JxDgZ
V7klj8Oq+3ZL2/kR66T0IvZk89FiXygdwFPq2/hvNMvg8IrwOECreN0+jsnHv/VHaAS+esUp/PqN
hPPEFMmpllXIYnpjpb+r2vZwh0eRuWTbCQ32OsuWDlpagciw1XQjIaaLFzYR/9AeldcyZ4yIxWxz
kt1f5SntJY9MoIaN8P5y9Ixk65itZ270664pMU0PiQ3Ap/APKK+sc263fLjTohnzyz9CIRM5TOFS
qZ0wfuTesgERFs+aFewJ4IOT9VLKgkwaCTRBX8vPAK1XrXjfyFr2no73AaRMxB449gVL1X43p/Rf
/aJ8VhhXqxzhlPXEY8e8CJ79DHwNzLh0oDfAaX85rRWa5skUF3xQz+h7Cpd3A0Se2ywcL93gOZcg
sjZdThl5/PClTmlcfwvjp1GsTSMDrCxd0xiLkdEvno/xX+xc5z8FyjGThCr6fG2Wedu8HuZL6aWn
wF4z+V3YPQOnFIf29PNMwM+bfBdvGBGgNP0r2iHxUffcMSfo5uxHq8qWKmdMcJuBUGW5l1Ar/Z/n
F9bW+nvx0a7yedBO84ymAJFXzvSEawzk0qBZkQg6WICtDppErMTr1qDd0cVc3vJOpufQTrm5i0IC
8gT0klray24Ws92doFSXryw33cuLuzQ9zPFUH7uo1xJe/8unsMaWLphGXGgs4YuRgkfTldhfqTHC
iU0vJunSTIwMgY7tZYAcII5GKo5SXovVC+MwR52DvKClYwgjynjS3uhjrij8/g3ciwzqUCq4DhCR
CA4GnEuQDjTmXyuDWL0EKuJsvjNzB/jBtDSutFqpqW1xHj/Dz+heuL5tlp52NCNHvc9/H6I+N1Dy
6ee5gE0B9P1YzbpLB2qKcBykRMlS4BUiV9fJos1IRSVZghOtX80bJ5QxdBhLlT8lSK4n3ea3bykM
kXP+tQyueuRzhz7NcQrwewT/mJRaFB5tsY1D816R800Mz5XZOXHAoKgGR5FHsuZ5V3zekzzdUdTD
j2ehTb8X0S4e/b73RP33/UZ4bLf68g+qZHgMyPtahQ4EXsqvWUr7kBTv1ZQ9NhpyJEFXlRx79r/l
9YesIzmauVsq1DeIvLem3TbmknbpeKfx1U+uC/NV80xVCGtjJtlkisQrc67GrkLQJwl7cy6hreda
kA3yA8aXhHlKALrCGLY+gj92RTYmj7sti3ahBe1aRfK2WV5lr3ZrBHYNrcqvp1VaXWLTA27PaGoA
xT+hjFdtI5dfwSV6Mja4gglAnnDa7AkZeGjz5W6+eiSVR2xofyWRFjIBX2cbULnRqsbuPoTtXMpt
/taclxT5gF67pyJBCn3nka67F6LQG8iDAvHP5+ul/Recw9XOX6QQkCSGICxLjcymsPuXKzk5JlNl
PXaBdyIgoMxLKILefZftRfnT78+aUbLV86A1nj8xwcTZVIxFmVSfPeff9I+e7ynaNpgfTgO9ScLl
LtcIhxKv4JtIbduGC3a8shGV8ddRFX0+pMzGo0RTzOopdiKDVBTFlMxEao6PLi4xnem313XuYEmX
iWLO7MafMjprou5e9JcIY3LkHBYr4a/kRY2Qaw4HsJi5qw6UfzLuNc8aVtfYUYrg9Ec6l/ORw7fJ
hcJJFXpL5xnH9qz9bK3vI8qQslk1pS1atfmt4MgtJcFwQbPoIYZnlKB3qKv3KX8pny/WPqEU+PBh
z+ihitpqe70TP4S7UhW9FN2yTgr8Ck2Xst4Ef46Fz+5gm1Y2M3ccSLOTUoSGJkeLqIclJmuKGW41
7JFfof6JRo0e23XMdR7rkWVY+2ds4Cs39AYGrNYZRH/nWlmhQ0BcV45lsMomzhQ6clMQNLSIIIIE
utzwtiindKse/n3z+yY30CfHxywU/XvnobtKl7eJPFbvyO8GNfT7aXwUixrAh+8wgxYQHrfUqpev
AUfZJAL1ZfKfW4gqdeNNZpGW+Ov27obmsG4HRuGVMQ8qb789NQ0dhKM7Y/+Ksu1b2JqbaWlVpmCF
XJon7M5NnNOrdAmY6y4U0L/a/5AmlUqmZQqQsfQZrRiYItJj+CF7s8CU/QNetLHl4kOSeGqGVb7P
gtmMHT/iVJP7QRG1xgl1rQ8nj+PO+jidgfnL8FRh1gmc9B8tzJuqMl2rk9LL+OBAoJkqW299f81b
VNrBpjgbgSkqSyUfnEL2Sml2RxM9OoQAU9PBh6tXfD87u2GVFgkEH0hvE9Zm7NCM7CsX6hvMP+o5
9p+7u9QD29nLW1JCQGiHMsYktpk+ZlwKLrCHqCrmERVCDpBy4RnPYXpooHyDfcODsb8IL5ExBzMv
GHLiiDv2V/zPQ4ceRFaj3vx2eB8uMJnT5ige3SjAz2rkontsX4bBmN/HAvxkV0g9VrNzMJDphl+e
KINVRfo4BUb++gn934qUn9GdSeJANUmvxQ48rWT+YGoyq1hOmDYm8/qtdS+tzqt7Rqq2udbytJJP
KoXm1qSXefyNHLs10LVwyH+95iQQysVNXj4rq9H0veJcod4Nkx9azXsENeuutCfqKw5jscmXPb5a
zZPTMANxZD5JiscCWznt/+/1Em4xV2tP2eJGtyCSbVoaQ3dXATYS3r+SynChsWUGKDrS/ym6YUqD
xIu0p7d/8vbc5e5Fx4P+3AQCC/MfEc6jsjF9cye6wW1NKfnAsug542pZw1hIQI/UGg+Z1zuq0jS+
mFHzr9Od2Cl5ww7fK9sAQn4X07msovLEuJj9ocE4yZggnX3iPDNTws58HazopDl08ctIkil8JfUa
pS6s91P6zeGHg981oCdBuAE2dCY8go4NFiBknVruGzbk5AIUCBJ6d2IDQTXchY19B6SriySvs32R
KgtLVtglmvEyV8xGCFFaeqC6qeTYZdOz2mMIvjWaqqSwmbFz60TRsssrmAspomG7qq7G2k9oosSW
vE/f3lDbGUzLQQAXGctOs2QUBz56f+NAUQaFqhzAE4kxS32HFjzNrErPjF0icKRSfNmZUd3rgNRV
NUKtEk85EYzrz8M4/qXeyXzv4uLsr8/ha8C5NAeuB03H62MeaXXI7fAWSMPW9ZTD+o+VlmS4ePCo
FKSOiS9OkABQEa0GtpT+DVmGjVMPmh/Sx0+OhaweIOonkLwMWxXsHbescmmOZ1/2vWrfH+vQaOI/
f3EouXbT4Qa72yMkue0LZDCg3aM5W3SmRPqz2s2LvNaURwenmAihYKgQTm7NLzC7ARKxsY2YuVrD
7O2wV9D5nyrmeYqQVLPEJkyqzbXOZLoQ1RCBbkWzrzwPEwTGo/XVvY0hXqcpGteonSv37cOjsnsa
8XQPVh2P1mS2fhJt/CiPZUQ0FgwrAhOWlDD0c4StyLgVFZPVOp2P4JpTRgxMdHJGyAyfhq5ZEwAy
4AN0jhBHMpkfvEms2AmukRNcuHUBfOOZbwh2IVS9tCBqHGEw37rRqGNXmsgPd4bUKv/6YQSEI8sH
iGIsztaXKIsByHokxG4m+WWezWBrm/rPCsEzoiLylbJIcYXK9owXYiK3Wngz4mC3p1ZvkBPTq1oi
/YxfifwXOq/CeAVNwNvcjTtYhH39ul7epRS3/OoD12Vnk70sYSY1NObArOX75n/ZlUFq48RwAVKC
0YKUzFnr8K3VmUED7Kofys/6IjKnRGQu/Ub9OlKMwRDJnysAFoFd7NuPizeJSaaDkC1UmXi4Dkte
6WR8SvwYy2cVGM0ajWkxOKbd/SVMbNqCOIlwZaByKqq9efFjW6JYzxODo5yU46ZzNSjIEusICn6y
7uwayyHrqZEdq5MzqFDoUqny+kFnFeoxxSMU+QHQCvuxrkyje7tgcOBRs/6ae/oVT4Gr2FySrAlq
wP6TitMotBnGPP0SrlhBjoAko5bUInXgBp17MjJv55p8+1g0k+eq6GpUSnwlluD5SeVQddwXvgjr
C+2BuFoYUy9q5WnxLmqP+Q6HvO5ivsJ8Yj+lN3Xqz21EsFNWnDXKhpfk03++TkxC35KUfoCa4Vef
iZ01MS+B14Qi/5nZUzG8CZ555/Mlz4ZWP4Lxno44Q/eooEERWQlRPNh79k885vanIwV+hTZIZrkK
VD2hy0cQdp9Of9N0FhJPQItaR381emgMrOf3eVWHL7jnO4LSQ0lfthoJ+IaN8Vl4BZSuSLPKyFeZ
RXbQVCnVrDGNlDY6I1dryVldF1NVWlFZAASrR0kvXJvdLnzUTR5a4Aov7c8g8kx34I2fRi2tyOPo
kEZNMOENmmolRMbC0SQUOvQfSGJR7Sfxpe2YlsLQL2QEL7nu0D7GpxZGV97f3H56AldcsUB03pHH
++y+riKo+f1KjZFzFA1FD2KaiakCSKhBIWF4aQl0i1uPzgIEezK2QAT1HR49TeAzemt7W6p8vbEa
Ww0SGuTx+HzjMqKqAFQuIDoiBjiBQ9kljYDIBA9QCYvJTTMK94VW8cJE6a2EEIC9wbpgmOVvs6s5
Hnny1EwZDsQLEWG9LoY/KFajqI4LNLJseQwn/acn9LWoQYzf3MlyZZ8CtoE9sPtIEYzP9as280l/
sIwb78gFCD+FUXzaGVG84msr/7EPAjGAV+keGCviPTEXwH7tGq7bgcEdopxBqpsPc/4iWUPNc4QZ
n3iUhAKDd9PC5SF4BMuUepDyLedYi7cxq96MJjvtG3OXdodXxJ9XwDUNRykOMDhJuEBVV+yHGkaK
C/nbTFJpnCSI8P3zJVE3MtPGfKFCbgVOgDdp20u0OMVZAirMLcgpmK8xJ66EVIPgFN+yC7G9STjE
0dxKfjbjO39Go1qujs4hw9zXCFtAototY2pTJyCuiBFDf4y34X4fwqHEouM0mDIZOQJxzA8FX2qr
b5quLvzfLR7ttYmOjsy4MFw8YqpyZt+9c1FFG+0oel1ZmpSe4x8BklsWxotNSBUmXpgr+UmQfw5I
fzO7wLoRnCUr4W2/WzNBk8f7vs7M7dzTvPttmQE36b9P8+J7/9I2VcuhYMnsYlBimfyZfuGZlTBJ
0Zhy41/dZlhdV39tMQ4/albSVRgUMp02GNrJEh90nY8HrgZuwsZfMnUHXxqT6bLi2UIjEHO8HEFZ
ajMsxCTAlq9F+jTAhAI+TQ22LX2vzxsJkV1p3BVAVdNyLCLg3VX1sOfOykRij0O9oFue5/0Oslly
ofVjzbI+klvnelrw3WnyuVK8z9207A9wU6jF3GVZx5Uw0VDgN066cddPiDXzGi9WKzknLmv8Mitd
waXyl8wtkdkU7O6njfG8LNhI0gmzCTe+ibvpAH+HsctoKB2nQ0EUK3pyRvz1NAwuVV+u8HYk3yfW
A1NgNp1jMSK85/ZQqH7g3r2mFcfayjK6zViFaSXsmNPgY0ap/cqQRR7jT1FxQa+vUVom+4ojcsiA
rcqamtWBKZI67zLOaDRxKFrVjKHRTHznRA2yhaF9WJj2I1YEKG4MsupiZvKaQ1W4AmO62v/59U3H
H32hc2PfwK1pFLwoGVdmpZXuwcyCgNqyg5x1n/fbOfMUlV5eGgvFiCYxbG8sUQhqC8kEvPyirYOe
0ngtrytAIeQbDzwwrYX2rqTSd0RggOn+xYoLPYkbWqlm8a9kG2O34hFkhl+Oq16S3R5yWID03yNv
6jcETPk6tD+axEWkvhsOj9HPmxl796sb3BZ4IgdUCwZVZNoqlcrEwKOc+328LH8ac9ORUxiuQciY
GlSTq2yLe0V0rb4cjvWqUjmE7uBN2Jdej66FwbwUkx+WdjEy4LuylOWT3f13kvX8A91RTMd9tBn9
X13fzMsATQqf9mcj1B/1Nw92p0wu9PjqxiddSwPivuscmd+/awxNTIJUiKFP8r4LOwa0uNbklLxt
xSbiO8/tI62nE/i1w1Oux13eptLn/HOxyZiE5Xub6XFryGKGboh56YCfNEalWh+lC/p3NyUMBjc/
MhyDi25n1vR2kSjSjkNujjJjWX/AgLWenVgLOYo30+mU6WFxDOxrAaXKsfZOHLKAcJVob9Dwt2Vn
Lgj/j9jZYY/9AebGw+DZ3yOk9kqEzNsrfFkE/NZ771PhEExa0PpZ0stYIku3cAqvrYVr5mmlYhxC
LH1Ihnd7bER3pVRg9h+bkubFIAT1gsMeB0qDvbMR5kesRsg1sGElEvoUcL3OcGWbe9omozwegMfg
hvN1TcDd1hXzjvkk/aH0oB+/+lv1mF9fFzQZ4ivu/MtyJ9gvWBldmbVcS5iB+qk6eU4xwcpT2Hc9
MaWE2NM3iJLLXmI0Usg3esxjt5Saf51pCfdgWv95QbtUCWTtCyyXtRa0u05qRVm1kvjmIUf/5ZmC
6WjiPdk86v+YqMt7xz52vgBjQOI37OW9icHzKxFsV4FL5GF2xTjWXfWmxeDl7KhOrnQ7YwXyX4Iz
Sg2LlxezJ65RQQXKIYdPqRtSrG8yBKW3BaNLS+ZoCQxP8LVNQhobEfQ4+0GyVihh/XEqkgWs5uux
Dkfj5i/BGY4crQSQoe80Yaoc9vzSwBfkCxV3Qh+L4EnEib3/lxASeDTMycMC/vprPovHVu6NY6jw
6fo7noG9xLgAJZJYxRq/Objp/wAz2X7errV3LKvlHrXm82/hMJPukJpwSNnarktm1sxV/fmXYnMs
yA5OVA6f/VGrk5rznLwOrxwo91gmdeiQCItJw8Mc8Ivt1P3xioALQK/lLLf/NCBo3H5g9IGFYyVA
v2/UywCxfemDumxofOH3AOqKfcjC8GuqYQRKgOF1bf9cmoXpEaXOelGQ30vfCyohhzSEb3UfvNUf
G5QxdnWCbGdMPu6S0u9Pi2JL8xSZqhEAofl25lOJuXGE2iZ9r7hVCKnVS5tk3ZjATaUd5ZDLSwfM
O9N/y4ZMbG/tNxyds+p2LQQfHmYBLwUwhg1fAciTBC222I3UvVQMr4qUMVFqryZwAQ+lH9KhPsq2
4XX7t89/ZHNeDcqUn/GKPC+JFm47lLQgUs0V8td8kBPv1KnwC21yyWdzaG9HIRxnnIofwdQthNo/
S+tAVkkJFLLTe0x7DxxPVbBTrb3josNgbV9O0Qx4pWTMANEMl7NKPYNL2t29Mpcys79jceMrsgfx
jgjvJ5wrw550HCT4uiGDp1BxNAeglLMWoGj6T5Mc68CtFWE7uZz86IBPCEEwypIRlsgwLg4cTdYw
dtzTjAxJ3jAuVUvoJy6xzy/mcAAxnznj12xyE4zv17B9XyMUqmxIAtxb5OabgSxDm+b8HFPBW24t
pbtw6Ll+O5w0t04gyXyh0EGcyY16DqaYgovMGanY5OG2DnVt/EARG88w1nwuhxOXKyi0g8mxcZp/
tRJx14ytofwFz56iqb3OsbV8kXKdwUOnlGY6vO2dm4bsG09dGEm5UWIF/q59e1qUI+0baYS/PbxS
6LV2yMgHbYtR6lN0VHtEqJv2BBhmpJbDSqGV1z2IsDvv4I9emhjTQI2aGgRr5Hd5B0bm9jlimZW2
E+iRuV3x6RVf1kCT3ep8BURSslb02XR9eO4O51mA0OlJOhM0ItfL5cQ74Bl7bSexHbTfe2uhaabg
O6i7xRvmI3N4lVbq9fu1hHjZ37qvzdTmRehYah3pGDkwpw6wqyG8T2+CXpJ1DRr2svnFP70UjPcy
m02hRLsomLxXEnYUjjgdkl2fz5ggP/9+u8NvCINY3ca/BWX49liLdoKOYCrMBRbk/GO5URXp/WR7
ZATospyf0dMLyiDoOffm0tAOUR48YBLLxwM5GJ+wby+EKhrtd+Jpep9je0xw9MfR0lz31Rf3wt+E
lwiRBOBP+Nk7ZVBuKik4mNeOMzkML3+DwFPs1HtFuSyTOEqc67VNvovg1vSUaZoNjYwxvDxMcvRL
4OYLSUa1dgrK47T8xvslkBAzXMIlcySLq5F99F1VxRSIbzKN/VRNNzLQkZ2as8tboNbnXbrH6f9q
cFhu5txLlGS9kmWVhEnHj2XZrIEbtZkGpgjgDvkU34qFG3MviBYzsLi/GuCqs71jXwJw4C1+TkLy
LMmU4HZCsF1pFnq3FksccLc8yAqqT0MCLWKMdFBoI3wGEKvbm531Dx5teeTEolF4pCMfxWLu6NPT
xRvqqRYjfLJdGp4HA8/vAn6B8alvbbfiqrwh9eJObB3McNfw4cq3NjIJ1m/7jTgbYdQvnn8ENbup
eX9Hrg1m8zK26aQ8W1IRG4vuj24oyBh3z+mR3yhG1Ie3Yduy2EPgai7Cvv6DCzUDRxcjc7xeXVb/
2bxdvkxbpvpak4m7qSqLt9uZpv9owh7WQAvmqqc/wDEQjrvuLCBzZvpvOZcjf92Pcmwh8gQHPYsz
owaeqgApjR4u9Bm3p/2OMDQWvvMHfKhkwXkVtFjvIx3RcIwsRaiom+gWwRvRDKpmk/5gERiw+qiZ
rBOp2q6x3cdE69aeR2yeqNH7PegcN3EQzY6jEgmHKFdTZ0V1joYENTEqJ99WWkkMJGHkde6ySi7e
+1XPiKKjltgZVT3VrE17fQi8Hw2fqFRF8YE995el2e/4P4RatV2kMdsWyPf0KN7ncAooHQZO6hOL
tXiH5Vvct1P9cdjAglGrTALGrFUXsbDHfv9Fx4wEl5CgeHUud0eLiLZ+0xeJ7/bVbIx+vdhUOb5B
d+et8gydStywv2SSNZlq2YIVoezlQGeaIpzTGc4LirAOQRezNIgLkA8fwa3cw7kwdJ15yufV7/UE
oFKBvYkbQqO1ELL/YNgsg30FIex/FP+9rez0VADeMJrf3E2T13gr/JnpWad1s3ZAZ7AA5sgPIbGP
dumInjkI7r+yhmbGkLMrbiex8MQ5450zR1baZ7yJWv9ZRgLO689whXKTI6HiKT+uHBGYjzh1JR7w
gGc1jiaa8xmK6vNaj0DMdOlZsefcUep7bEzxMvClSkPRS82qeFEopYAn30gn6HmNa/4hFpekmuNs
nas25LEzZN1ulJ3+DPj+JJisxXujbKpLsiIXELvfYq1pMoyXOB10fLlPGO6UYPjRwbHLACBK5iR6
8+OBBSPUWVylaJwKuI+WSfndKG3KxwPlQh8OTbETt5zqaNlRfdgHsLuLfuw/ewnJR1HYov/CoiqG
MwIk/DXEbsK7FfLViaz2LMpbnAwGD9Egrtw4kgBSvK9LW9HB1P0KuxW9HjIIbKWMbRu5D3qgP34h
NeKogKjvMfuoZ2Xmi722ivBDbP5SYSzvS5PUpSuLQ1vP2S32gGPzhanQgbK1q0tP1NZIPIW5rIEf
nAGWbyDKEID6cf7DURQviB8my5FbBTcHcQNdZlon15/GitUF9jpMkCC/+cgxNzaAvFMQzAHGTgRI
qrc6Dba+C3d1PTV7C1xnnlHqtiD78RX1l9KhvPiEQHdAyBmbWIBLyvFejXgbWC8daFBpTSKU62Od
0MeMluZMxSfX3Kz88yvjD5o5aQOKS7/222FK5i1UhHuIigY6BCKVd26yR7Rs0sCzd6OwNPqb7Cp2
pq36TVfvLiKDq27EOG7HCjeONiAslW2w5qKtKvrccoCvN9xSE3qV+2vOLs+vTv/Rn6oIcz+d/2/c
8WuOqxvmQOrEyyQBhkAY7SqCU1QCJqHg4S8d/SZidJJF+hNysbrrFG+knHnDsp9NQgkqJ2asFJz8
ax7ve2l0DU0NqGEuz+Ouh+k0xd5oEdjU9enSq0daM6vJslHHo4wQSGHIcTg7TbdmTV7NoEO6rrr2
6czj54fAy2LwUGq6NXGDvsf0QgKHIdypLJOnLbqxenUSZZYks/YuQnkA+JnR7DG3MASuIMaH+deH
GPymgGWzOyOvih3taFkxJPZOP04Dc4GxuGJBLdoZ7VSi1O3fryIIuyauwVluqDSuONI5qX8vib7X
Q5S2b5nf7RJVPnJp54wX2KG83gygao24IF0XRb4m1EGHiNt8wgYGZZ9X7uL5tWxYCtRELoNABqMA
Avqr6t+mbnSioHh4ogNhiymq97FY4QiJQw0uVPCyexS4QeSus+ueNE5cKYNfHVtFQzzY8RWueKfy
J3h+/b55NTERFfooEl4xNYP7OCj5bdCnCirMtAKh09LKrR82Slc5EtQ7/8vNswIMiGQbLRPTtVK3
B3Fs8qRViokq3fTZ9DHZmRqu2hbbyd35fViJvKEWJp8BwH0dSK+6bW1av84sSaNKmfk564aO59ZH
1QH+lHT0Pw+uukLbS4DsqcN9jvfZ1iVAGnS+AX/amyEKpOlT+SVGfXGc11W+qyuM6Q8lFXkttd3R
4FzkRfz32viCp464XSBAuOlkZq1SIETgGE+2OqYWUaHTmNLMdDmzYrzuf5OuiqBjsPtiXXscrNly
dPiOiCFm+Xc+DhhhBfSyQR8BGQ9Ia5c0KkSVizDnyw7TBe+7t7iDpEh1Aj1kszU75u6vtIeo8uaX
rwfaYoxT+SMVSs+dFuuEoSQ1BOk888f2O/0MywALop2D90t0hERVAuTx38MO2FkaxPrqSNQV2zdy
zH08/d5Zqpn+l2wypnue6Se2In90TeHpoqy4GX6oWd2VzJIG6f76BXaER6XPCjZnxvQp4YiPiAee
jI/a9xbYywe/2wED8t5arY2ipEaub5m8yzBmKnZrFuGqdfr9rRKSb8p76Nutj4JwhxAsmSPRA6D+
6jCqRq4BM7xV7vJvfb5OpqQ5S+XAqAZJOBXUO3NwNiqxYQpIeAtEgkUNzvgZ1ydoawaxKEhJsEoC
TN/tiIMQao4f2/+C712fBdkU1qIt5eKaEmq0VgkSKGHqPZrP6cDpKf02GmGTBM8vuBpS75XtdEbh
nxTIIW8wffx/N/ZrK+wCIRXLtKOOVt/crAHp5A+7oyJR2cvetB6MD4cq03WK0EEr5/G6xBwjpuje
STysaGc+9cjf//GJ1oeIdWvtsJCeTpKIXBoByY2gIW1chQCLBiay/N+LqdWTU+Vhc4lQdNldhrX2
xnbab1tHjAN1iGUYabIRwUQ36AZsoXs/elt5FgJvOZ3W1xJ6DmvlOeyD5GoGQac4NYoNJNX/PjXA
M3uxVoIPzNCvMxDSi7Zmn9tcy5wBacYECwpADtHnirTJav3VDC6y1zqihh7akkU9xlBJR3U1hliK
7g+4lfvF7H4M7wNQmXgHbyIGC45d/I40N/2Ac1TdnVT3lM3jQBvbDGNMN6my2697P82dLVcQf96Z
F8YT4Ys8/9S5fdA9AN1yiI4kSfbM5wk57Nzroo3Elcnt04V/YxljoO3VT49xcz/oRasziXuLFZzv
i8jMQU+sAmjU6UcrHF3ToXCzzlVh7nDvhFFRkuAr5I70sJhp3fxtXBH1MTGHQrD0wdUbNLdhlLeT
i+K5eiqBKXiWWQvSb496k45uD5/FYa6pJTlZ7jMxg4mJ9VAV5fsF76ISMcljWuBV2ZC/G+KdH35b
g0UtoshZOUdYPm5zaXaZLEanXboW5sFdUanF/ECa2uQRHqEDZ2xWS3kGuDjuBrDmxbegP3S7otuJ
k6mew1kvxDiePPlOj1x/jIe018wnly0vLK+XIpFhOVzb9TFGom4FdG7IhmMvRXT8atGrF5d11bK4
x49T9M7sQs0EHGAYSaUdaSjowqRCwb7hWs+0HsgBubS9Q4aHxuX7O2JzF8ssAk6n8sqIrN3NAh2a
J7h2TF3KJjZn7w/0Y6IvOpJdj1XOsElWyUTpjN1+e8/ggWjPIYqprqv0SFDiNxi4lkyWQgTXWpD3
6UIOk6Uo2db403HYbTMN/N6+9I8GSPJ3xFvm67U/A9Q27sEiCvU3j6SOxsW88sz/q1wVDesIEAs3
OVBcZ8iZZemei31bH6K5qqVd1YI+BDTqeXQtbtTgQxG/lyoDbfDUX0AI+xYX5sOgAF3B81R8GstP
u3Vf2JLcJ4wn69/8SPa68WLfQzdEyPwkS6PMZ+7TP4LzeRUyOwxXiJCErb5X7zsYR+0wXUYFNRFi
ARaYnkgda26m4KEcoqG3zi+9oBUYPGRL/1+DXyMILvYqM0K2ZksiA1AzVHnk6FWLQt3i+/9xvb+q
Q6OWYApCvZxcT58rnGRbPeo29naKdeCW+Ix0KhFKV8UukKALGfupDd7e2dNuEnMXZO97QGOBPV/1
5DDcGnoQ/9JpIngxBHV2PlB+fqfislTj3jFW0+WmsK87rJ9clbQAIhjqvzxfLzyiJ9z07Dp15nkN
7UYwrw1TrwCH6Ozij/YRGv/LBgg8HHCiaIEQ11l/NmYyeS64teYCQ/sBBNC2vEJ8uOZYxPeIAFHR
/87wn+HLCI4B1TSrMBzhHopdy7fqyHAtmpcnVjy/QM1I1PJYpj3OXCezOsrjTsk9bmHauAtdpQrd
gObBolx+7jdxz/1uXtgS9JVNp3eVG5bD747kSA96/XcdqrwdJSTp15/h/+1ichayW9/SMH7XcNmB
EUeCXvxVwAd/CArxJm/HGKmER9J4IJyxvrmfeyg504xCgouDGC+Q9+ArK21NIOiXvzh1OmxKuUHd
IwndwqbrR8uqQCqxM/HaqYy8d64Judyf8U6LFn8/qKPsTQxY54uWLWGDwRAMevbyUELJF5skzdDN
jDS5aQFqKOAK224Ih0PePFfNfELHyesLNAg+ttl1Bi8EfSn1OBrKB4w7c53YJknUHd9jTlAeokE3
PFvN3+kpkMsD43D8WXPVLMOHPS6+7Y39eeFMOon7quVA5fGzI+mGkgxQRqewBC+NKvGRE+TZ0Gdu
PrgFqlGZd+s6Lg13hhij+6784OXo649p2FsxOhp9Ix0I5go916n4c0P41iK7/4kEIm2/3V5llKfH
QSqPS6u1uDekLYUlGyznxS+6o2SwCCfghX2K+mt0mcvbFWzWD/0NzUR0+X4wtyuQcVn1b6WsmUgW
4v8/wkhOQ18AhEe2XtEXstygqVOjYotaD8D6DeTUiT1bs1IIKBjifakGu+a+yyJ9fkNLDXOP7Q4X
wLZMg0BijQ5DQ6I25V2xt7Nxr5sYSOAI7DJc7kdi1+K0PrF4I+hCvv1VHZ5YrpwjxcC/UNemyeR6
VcOkGlrGfr/urVjW9+/vKSrMbRS9ISoW3i80rwVP3wfUz1DzX2QCDeWTd6dwlQh7K7PNeLyr9vts
4vPb3d7MS2q/ak4FGCzrjHWuagq+RmWWRy00Wbmgj+KhyhCZU24O2efIPZy1+/q4zz+MMT198UEt
/DGwqHDrHSB9UapVVcTzEv8FUJ25K+uzrb4BiknnXH1OU7EGrYc7Sby8HYWMnY+C/Pdoq29Isb6Y
wDgcAcQJIDZAFiriF4hoOYN0AwcPt0/16ycpZN715nlLSuVGyu7tTV+HHuxPCfKDdJPyh8FqVS66
C+E9tw0S4lNjsm3PQcu9UdvvZq21SizUn/g36Dy78Rh+FiysGaK3WUeAuBCWQA/CyjNUG41+PeZ2
TxNpibA0yJB4bcC+qxtSJR/8QZbMgCQjCRD50R+e632g5BwTrjev6DW2cGrcZ12rNLWOk/DlVlJd
Q9eFtty0LL6r5Jyd3LNTXT1CX+Q0qNs8wNhuvE1Dx8/hY8LH/mkNRoEKhAlVKwSt3DTvS9MlKdz8
M143UKIb+rhZ+F12HX4vOo5GBX/lTgawwcS1I3ZXBEy/g31LKfz+hNzSAwc804yuyb4IIYAQwIFa
2jpDjZ6nPK87iILAtssl9tuzRvNIROnqZXdL/bo0p7Cu+uDdqhP0mQ6fTMlCpLN4wwGO004bPB5I
DwwA5/gCqPIq2Or/+MMUgTbOtK+xS2Gk6e6ZVG7Kzk+vQI9IevGwTvZ0GYS1qD6BhgOd62iuMRhq
y6XCxSwlHxLIEsSapSBOQXkAuJXl+hbmV1/0fLTHhMWHv3cQK4Lrsae/68b1jr2sFbVLehtbQoY5
p8BDYAyDqRVrRn6PctbbxMsNvAnH8oYV1IKdh5gNlzts5b/6KYKXzYPd91+EwnLp6liEVTfhiR/p
CP/ijKPHDa7Ff1bEUHiD+hYCBhui/xJQ4/FAtbyvLM71taTb9tmkgDsRVwOq04PrIiyFVefaeBuC
5zcZU92m6nFYB93DoAUL2HNKHUoqtFdRiShIsOKDC94a7U1X/YTPgnw81a9qbhUZHBtTBognNTtG
m0jfWvio1GEHTG2IEmuHRwwgYioNKUYsJenAE53V/qSENnKP75kJn9wCubeq0U159wdaSh9uXgV4
hAmlpQM2+acN65D3jOm4xHuXALI5q1HO2YgiO0AGDrHFK8oB4VG01C9hBcivMx0IV9T0315+5Kug
GPe6gRZC8s5cclU8A5xi7xX1zI3/fGlbWLmhQ5vXb5qddPMXHFc227mS0BC4FDjrVAojKx35Il/r
EgUyqO4bk+2AyNFDog8z9Mzd+Z8e4yoJPQgWUuAQMjFgY6BQV5E362S02x8CWFqdWVz8i6qlgwYo
T/QLFdnitIXNhK6vbJc7KF6znGjQKnjhP6879onVIa0G3rwE4Ux3Pp2nh+SAp7tE8ofClmn08ksy
qYctrLOUrUQyh1Kw6i0wIQEB3msFWY0TetmTOo2o+h9PDeA8BX63FGrb35aWTxyj2NP5ZoZ5F5pn
EbYfx0CnrGd7va9MfD/SFMF4qA7v0eJHzv1HQKh2Nfd6de7VXFwn2qtHF9luAC1GKIv0921jMPXx
9jh5OVNk9x7YYiU7FZn2JA/jlqyEIIRLUjOoCvBqfeng9+Yorc5lrr9si1SL037V4r7BEu6JKiq+
tf7yfI8w8Sc5mMca9pepxYgxFjPYr8ZQFUULtKYCxWXzP4ZDaXGFN88ywUEeKuGKotufzTZoVQ5y
EDwHoAgU0Bab7JMfBEabhu4TNYEJ/SPV4ffR7+8yPE/JDDkxVqsjOcyJX2F4C93xxAJRdoQNxoDT
HxjYrTucpejbnmHfZetkLSFFvJS5QqjJek/sPiIoekoQTdrFZWOS7kmP6b9McKi6/7B1qWort2xK
dp+DZ475dSEvh6dEqUvEGbMiOBxiuxRWKwKLoYZ0j8mvQ+x0Q67r83mOGAuGFF2vbj3uQ6GSzdWF
dlMlHmed+EsQSHce2i56mhH/1KZ4Fj5oZ0N5n4WKOiO61rGJSN5L7kvZmOoIxUHHLdCkjC0OOrdE
EK7afjf8OFfvN95MQCRN6iwu0Uq+kfs+ZWf1Jejmzy0NnqCMTY8dI82/v8H5crFdLgzYR4lSPio3
ZvKIO3fi+k7kMWirsaZMmDc/3aoAdUFkXUlu9vApMuufXM586812+Af/S+oWEuS1LOh24bDEjgpQ
3krx8tJ5gjm/15fwS/RaU8mHhL0UOV5jqI1b5YiCepmNNZ+GBgOLJ4+B/xfBJ1I9HMaBrIILDtZ4
w2TcJhA3L54TGOf6lLqomdhSEx3SUEBvPCxC9atn5brcYzZ94wZuKTWf2HAbMXUwKuJDVUWNtnNa
pqfaYuU31EKQ3cK+M7E7SsWteCgbHhFYUorwGj2sbtBE0c0lh7OxU939aWvDImjFTKjrPnnFgSol
CdJihRAcd8sGWHkKQZOF6yT6O3glAx+fSvtIy4VMopYiaRGncA1hOVMWHqaD3TGxYmJSpZM4F/NN
k2h7Nid/19ICMK2QdqdHYCePrBPaeVh9bKD2Yukak7YXjjlulTENK1OKs0w+xaagpsGQNgt+nG0B
tE3MWdJG/wKUEAI2FX+b6nYhVIQjtipjKp3cRkyMPB62m4LrL1HQFHl2FvejC2JZWLhWAnqkKeqd
CopXyLsEmhAK+shdUe5J37otdFY8xOm3YQKkvskoaHRSSTpEsu1iTOlFYdHrqzQ56VRWNShErzcd
SNF/ixO0t0YtWjdtS7MkbE03Swjmi0C5gUqzpZeNI6b6EvtBFqtftn7jzdSV6kSbNpGz8E05U8H+
YqlluCE26UFdnuuPbOccdzjJ8d7wA88WUlXPnMVp3+fhehzfWkpGE5JJce+iQvGb1RJ3HebrN0K7
uuD/pQ0MMe2kHwA7GJkDTarcDaNl+Z8yHRmv6xPrN0R+AIa3q/o4rYvrRBtqF494Cu93HzFWZYel
88Nvaw+j9+HiaswO9FM1D5Pt9n8hiLvwycOpy08vV95/G/IIsiE0u1VPk2ADgAzUYBDSs2+enMXZ
B8mea7B5L6JSfu/aBKsZ13m/fH2FL+SItOWv7h8B1fpJBdrfTWUuuCkGoQUblDemc1nkAtF4QAKp
MxBLaQqptdMVHyFZztg8BRnz8yMkFdErXgKoOSKWXjUJGdmpXyG2YTjHglIe1t70T4XecQakuYvj
SLS/LtBunye/ht8l4m07+f7+SorKzpKEoK1dM8Vdlm1A11ciH0say2cpyitEL06tDFvp37arqTTt
WZnJvSbeWVOdYkiBdUw6czpuDWsotSjbONaP/OlQw/i6OjKV+s74FyVHBgkv8RIigDIFoo3jnCOx
UqjrE7g8uXwu/9sisi+d3U7h5DdaxxtyQpqTMskXMuQQWbDdtruCk2G3qKFVL82yfVOLCgZu6cA/
7t3mstLqlGS7VkdHrxDNXIr6/WygHRHRmP22KCrFl3MuBilSPEbCn2VcA4/P4/yt0IbAPcQz+N1u
JkIOPt0bFYmcooJzhme6tW+IV4XLuoTvKm2jeT3ukeCr0RgpcqOJZqoyqKGwSXJph7NGLiAZ0qRg
yzhZUE1L47Yxedgec0YNUwVYIrgCo/j1BVN7XqmUVA16cJxszisvAc5+bPe1zFCHbkBuZAuTqHnF
FSKMZHtnhroKYNpOv0Yw/LKe3OI66p5VF03mu9iSIvD3FJVo9ZFXeIO4Gv9AhasF/Sx1RgHpWXjz
4BbPjVeten+knjt9Vgs1i1fcvl8/sVLuZu/vHjZzNSowUDbF9XCkjU3umGmD3h5j+Fm6IEcnwt/G
WT2WSVlVI+kJ0d8/0G8oxygYau8/KMVjK02DI4lkvzPZwWN6aF8z7yZBvSqWntinuEMYUhUgcL20
cq6yD0oPnt2yD2Br3Q47r54uymwOwVD+CeCbmaIch2TCCwJCpBCHh8UKphmhTxcmw5Z3o87vPnLb
ogkkPQxPVuO2upCrzmtTwDkJ5B0DR3o3+7za+J9d+CKUuofGtQt2H9VGegqm07xY3aJnV2p9sNCJ
jR0gIFr5yVAQ3tE7DNF5koP/fOUQw0qUWU1RnRr0QCPuAQMq66tFOYIxbaFZwET7Wpa5C+8j3xxO
HA5a3PgQqw7KDDmP6Q8t4jFnece2PhrqRk1ZayG8HuLgsFdoPMMx7oZGLIN02jjp72ZKVEBAeLxw
qutv0ElV51U0bxmLL2n7KRToG4YVz/mBcV5dtgeHRnd3bdiyhq79UD0JZ19cnO3K458fMpHbxw+Q
uQm9PjFsXk2liSOUdQqy9AtZiWI5y3/F2ib/ea5geFpUzQDLmGBrLifBqIo8Dq3VKd7pznfTO0IQ
RRXqKbjpv8SJsJRllZslOuHMucNew22Anu5X/62QPD1VFEAPZCgfdZxKfJLwPbCmQ4E7WgBHGpyu
s0ZiUz1Rv0m1oyu0KqC4GyYSj+SiaaFVVP+rMpRDqQmye+j0W8fwsiO0668d8AABYUFj7iXOdtwt
PuS63UevSJ4BHWgrSXDSXkWjANV1A2xZ3i7RVrAN4jhoOVqzE8mZvL4X1qugCiLoA8RTub3RfAHj
ITQpusBFWQROyCKBiSPSV80m4wsmygQ4NwNdCEA+wjgICmmj6A8vSvm0OBRc07ii6Hto7IUVEqqp
8sQOWCbxbOykX6h/OSNHEqpk33DYYkD2WUPj3Os5ry0Wey+IAyo5pzpNIWOSSrlfTz8U4Qtng0Zs
uUzQn2CAYqGIWnFAzU0N7VtGucHYAZy54CjGqty2VPg6p8LUvtsdpfCB93RQSVY1TZcR3u4uNfLO
xwFvBERvZqEgO9b140/B5hL40SlAWiNMHi28iTeeZ5BjyMqOt/3VvCQkF20HqS14s1SUQ8kvg/gS
b/Q4CIiPvFJwtJ3OLYEosRM4Gdl4yH9TnBtTrYGq5iblpHZSNYGB5jwHHtfLDCDz+WDL/phJdJQe
l+507PB2qVN6Or9YopnrgXTCtleYgMMxucXRMNARaLcJeUAyXuZUGoQCUR4nCM87ohFZePFqHnZ+
QJzvnubbhciX1eyG39PKnlwRDlcouDx/REu3+usa5abo51KDWc42oAaHAwTIiL90M9Pcqy5HIweq
UTUbNRirTIh1WRukAHLyMScmSojpj5rIGfp7Q1E+FORjem0OxDfDsIIHbG31iNblhbCnPecj5AtS
2lWC+tL4PrMb1isKg6F3C4CK/7jeDzS5Zz25Ig8OjBGbn/WZi1ROzgOvpgZ/HfJsr5QEfdm7xyvH
YL94kxglSagGG6xuO7kdFfwYaBtAB67mMCNMKTfG7xmVxubsnjFT6VS1F3J/aLhPvUf9nZNca6zT
CdITzle1NkXgCT7Wjrz4LODKwu9JiOHEVZeXr06+cMF839PT80f+Nx1iMraBF2bjJPsFDNpqVn0w
ix+87+YrezrR228AraVsxGHh45UVBfN8pFtFzFbwrdOZ2urrwvxVXoMQ6VZEGf8Z5HHKPYUzeFRZ
e584o5xxNpXd7tLrOr45s6K6Ywtq/w3ghGJxWOvoGoQ7TFHWMAqiqDrrYOGv44t6eRyVsIAr3zpH
wEJSb5JIUmfTD8Qid7JwyqY/0spc9ax63rd/IRtaEsFiw1ma4jCdiskEHJBb9DF9zmwLbAZp6/sy
fMD/SC93YSG363uLYx4ZG52UDyx6pheQTOrR6dx4pvVSGyV/1FcQ7kHwE/mN54LN8y+VHMLuZicQ
i1nSiDCGB1EeJ4ooLUCl+5e7MD3SRFUtS2ACLXBBynqgtWYKSufMD8FjEUe/aJdwTLzlRbNWhXYx
Ox5KFwBEZYC4vGC5+6iR2PTsOFsytqOoFuX6/Ht15DrCKh5cAfBEkMVRo99jCATzhlY0m4P+ResH
u8X2mbXHDSj8q8M5HmrnfLxlyKH15qP2sFyNrWCa2B6+TAg95EsbjaSVGdKnWRc6TtfTm/QF5GPm
cV9EezB1z6GHz+RVx/02yZ1+G114ORY7Rq4GMp6O+DAa9/iTfzNYeHvCp/LDU1xoeR7MIETC2n9D
2WVE77yPrzbNZIaxBguIUSiKKSJtkmFDtzHkfJA2RhBssD+X0PQOO+XXd/oxbkzySKZ7J258B8CV
jE/lTPtYcSyF7YiEpJ/ROk9O3T8B8/8lDBEWbD1khaKFbXr/lkBeRyX0kGppWly5tOf84wRUcR+p
OuYoggbWyZ20CAPlqNp8HePMBWie54NX0Q1DsFZsoJ8ZfC4r7Yn1KHomU6X6tT6evQhiak5JWj+Y
iXmQ9dt5IQB6fHqeJik6klpY5L4CAtBGejFBbcsgWG5MB7Dt0AOhuwTb+UmLljVK617KhHnuRKIk
n8/Frrubj61m2SBWpbRydf+q/U3pRsmEihoODnN+nQohQqpv5LCJzYo88vnZx4S6pVBj8zoAR1z1
yP5rmvAmSZc9Mg9qbXsQ5r9uBndkz9RAhoJ46lVuidacY5BKQJ/gUvypjjSjvnSRiCeIIsDAbRZR
ORFNA3g9WtBN6XmG8Vi7KRdw8O17hhRfaITGzJt4fxhhnXTNMenrka2qerU4XZsaS7B0w4in5NjR
ZkUZiBEXaVuJMrT6dGO6ViGHvf/5Q83KXQvLHV10oOF0q7D+tCFMYdhpZeSoAZIKKhQi71VFW1zM
vAVVt2gDqk/LWzJrFQBDQIz9YrL73XL73xRRlzko3FZPgXCbwKB58BjfbPSNKmfgHA99x6eOXBvD
j32dwpVOTt1hAkHGwJsxbtLybd+ncaGqS+0FDRss8aaqIi7K7i9uoHePGV5Zmk0kBkhNo5MYZ17W
GsM8bCufu0KxF74ApNF281ERQlMunAG2wCatOfB+XSclyQYOL/8YcfbU0oFRKiSC5A+513vMbz9m
+2qGDYOKB1Fxtqdu6/KNFOvgwk6XXITacbNWacczpd8Ewwz2Jmal+8/xicWbdBU4X+1zM/zQjC76
SpcQ3ae1/3Mx3wHSFKh+yXSgeox53wk8N0fthGv55lpPj+1Vu1GYabmWLUl7Xzk3mhOI3Xhtsvn8
mlAZYtGO86JE9/GnVycJzT5I6YpV/ikBCUTJnMxCsknanV+LbOqU/TN5Yj/uqUymlte4rmYEd8bu
dHWQY4j6CvnO+sjh5PcrMxvAoqsfISLOcF77YdPNTy8e9oogDsKp1Ps6x5WV5G1j+Pm2MWWXZWe3
VH9dsYLHvz9ssWTNuX8j8NJKFneeKta8saUpKFfb37rPqn0f5wPXboQ6+xMgrNT6Su1Q2OxmjQ7J
R7vng/O9Sf4/Y2eNdVSGZBwfvJ24VrS9xUMTfb8UmdoAVyf3FDTm7Bvs4r8MZ+iWsV+ie84ouP/C
PF/3PCMCuwMJPBN4to4EzsAZxVYXaeOWhQvnodTHJCvAl9wwd98Sh8Wnx2lenCAx85LftkBeiK7W
TMUNX1cji+qHzl0lK1s13t1gRo6eAczZe4dsFJyA32AzLNRWLfX+WY73VL97ZyRAT9HeU6Gb/UdG
sgHSPtWcWODEigXWt65cppZY7A7wMP5OCs0dLywnnzico/2LMIfFqwxnfkiufkKyDON3QHvn4XVw
njbL8LEFiKQ1YOw1Gpa+AcOQ6H4TX4VMQMiaebSLa8sZLIeU2bZMGqtx3eDpjDN3hEj5jKxIhdf3
DplnnUfe9JDAgWvBOi7CjDl9neMIswunScP5l3UZhSMDdtEdG/JK4P28ptKGauTvNKyQzsklO+KL
Mb/R4qYWjnGM8phhWhTI6E62p3WJH0x/bRzjyXv8wBpK+mG8EPNQMJMvL4ubmh3rjY6+TzIHysGI
miesf9zVXmyMWBtPFSvHpNM/U5/r2AnZEkIl3H6qCAwvcGhyd2NQ9ZBtwCdSq5hlw0U+b34GQ4aM
FwFaGMZQ6yurx2d0S/qZc2RkUpT9B3/v6QBo5BSbB5pkQBcvbFsT1/TNTvMxLdoHszc6Vm9Y0cDU
M4O+gDMxrdLOreYpXkb9JnjKfpwXxwbZHGK/GJzgrOpMfyxiRGCOHWVGhAGg7B8KaKR/4d0PZJx6
fsoxIEqlDFwLmFwbKVQnNugve0GGLczvZZU8xnX74d0RKn6ZoLmgGf+waffWCQNe7VHBSXo4QT8A
mj/n6xAvfCKcNKFKMLsRSRpvRlpV12f6icpqRDgm2DlQR7vEnyZ1TZ5/SWnRPmcBz/X87ZHqvvEi
GpIFKsHquM0MK7D2AN4sRpw/fpv9XhhAYIL1UqH+M3WJS8LalEjoqlqyqbCzFkGaIu4RE1koEv9F
hhvnJz4/+JeHOg1tzX8rjtWxxJanYFpJRbRhvGShD34ql2La0gY8O+sdaB4vUWwZFm/NUkkXSgOf
ssWArHGZ+QKp0OkM9RIEkfejrE7rarrXt5Geu6s7ayqYAdEzgOptR5opIDH3qtmWHJ4PsIivJJjm
7wHtxnBylsoMxMZlnSXVddAvIenMpiclAcm6xJJG903LXRGmytxK7xqS5o0//tCrB7CaTHXsT4H5
roL3Ufmnv0nCYj1JkXpQmC7TpajV0b8vGNNB0e9gZPyuCgkVHFTOH3HoadUFRIb2xKaHi3ynJHuX
zetvOBEFv8JqCazJnrXpFn/pr0v8X2djEUiRDwpu0uieeWvA9Ar0psJFz4e3UnM58PRIOlffZ8K+
ZK1oE55u4RDOBsH6V8xnzClv8e7qH0DxRGmkOFGiZHDLY3Dsgu2IzYnNCUTETH6fs1KClicyMyy/
cjz05wzz2GW1rvRrjmEwa6BS0jlCqqzvYYa1qk48p4RizD6EEovZz/HzVHkR3LhWgmqdfBuvBWxc
Qw2h4bD+Ldbh7yYsnzk90vaG+ST7/bFcjuWEbRzLwZ4UdQvJA3rXhtUY9gYYZyzYNJ43mObuH+rx
7DtxHmI/Hh3HjNT7eB2jYOQDoJ9BE0UEMV2A0HYxVI1DYuGsLe5ropzmHAYmCZl79EHUZUOnuVFa
j9Uu91PEP8AVqbtSnpQNJAmN0sH/rqXzE1JuyRW5X7shTmznZfBcU9OFFu6d21JVo662mPUC+QjO
5fMttGZLMQ2HoKRT5YIBNZPSBYDmXDCmhsqVRmIEWwDsyyeyG+6ErfpFJWyNYa06Jc1jBJ1COX4l
+cCLKiwHYZ1+/7Ud7nCP4lFjp90ezAWuum3dKhMRUhouxWE35uE3x4Pbzse+KaIx5Oe+msjVVM+t
gpGaP9MkhSCGC+zMSf+FKdpDq9NIkpkZsKTUJ3tAmua9MDut3IsnjPzc/O0ReKeZsqKilv6kVjpA
LaaplJJ2p3iaG4O/5pGf2dETlpfctcAhI66A2W9XrjMBFkSqLbnMDilkf8zzWBlN1mm18q0shQIP
tKTcd4lUPo6QFXW8jF8HZISJ+fmMcjO89KtGC7fuN0sl7qHIqSZ5V1UzJYN8jeueYpW0727HQe4d
l0l7HwLhS3LOw/VHFGzB+MgRGU4Lk9FRpFMqSfzBW6BVorLmeVvP91ov2ESENRq6JSv82eCZcpAt
L4A/QReEy6EipXO1xhw9p5TgC9BeLpOhX5c4mLxw4FLnWbyQ1XomtJmwfHrydTMvBQtI7YT4Gd/c
Wn75iF0tq7yXpJ0vblGadd87T3UE9mGObCdAjUr7vWG1XehdFx1OGrV2MYEKG2wAJuOjT56+ez4f
j5k9H4TDF5TWC9TG9BYs/hmgw8h4+0/pA80r54CeIRLxo96271h8LVGDx+kmPqf74siH0/fhv7/C
7nzYwLzPY9GmrCmbFZVGFTCUn9A7bSWzz0SRW6AxMsc/vhpEzmbixPbCkHGBsSsz/jEyzynGKhtm
84q/5qGe9riCwxDnXbXn81S05nc8hXb3d59DekfeVZHtPwTYDS6HcTwH2utyXOp1Wl4onNnyiQfv
ThqHAgUTNaKZmMCHlI8OlHWCji+04X/jz6Bv4xRx50rSgLtrdx0vC0kqJ5o+Ax1TE8OupkuFcL+h
y/PrZGtLi7lJwRxhjqoUBwn4nn95JRXMdvnAFt5xK+JLhWBfqvFQwWIN4W1Wg6hBcwW9AKgyGQ3S
hWuKQvAF032S8ilq0kk9NHgZYAmfglZ6M8UUItOd0iZ9lavYKXZrqKyeleQZg9WCalbEPhIxvdvs
PJyvcfM4VPZydmKZYNVQjUdqjVVHfXiX1udSFfXcTn60VX1RJPFEXrP9Dc11996vii+R9Ghg6vAE
+m4X5/NnKxNoiLW4ACfTeb1QISy7Tgp5nmV0FjL4pj2skdT1QzWWLKgSkwQHxXsMPN4Fw7wa/UUd
h+fkFbSNQnjGtPyce53qNPWIM003mRJTC2T8iiVO2xhDoBuPdAOUeBrhrjjmsldkzFWVM1/kNdMz
ZZowSja6xyXqtCc/Q7CQbCqASEP8PAe2LvkHawq0fqE0xYjRjCguBDVfhnw/Dwq+AW5W7Q/rQTtT
kNRSacH53zXpS21VITtf7YHTSPe0hLISqlmJ7iutO1s6nRChbIadusnEFYIiGyeCbCVVtxBHduyz
1ovQGihMED40UaPGAh8VE4JFELxHG8jWgK4eH2fBmcDYZCsz7Dnyf49Vtkc33yuinju66TfbsySW
8SDQQ3rJItWc79YlmjuHUn08CJ6DfrvqocoB2qVLvMzad5/ofiY4qwK7nsJuSI6ykP3wXc5pPOBb
+VBhBUr7xEb0dLyz48eDxUA7aeklxSUfHfhPmVDKpM/AeoMLApPrlsDRQDWZ6KzXv0GjV6NeXHHs
N3nxzikqeqBn5OQLESguWfMYD2sEP+1fIElsR2HlaGF3dOUwzR9PWSn9QXZ7XWIa9RXVxEpyZjb0
eeyi7TQ6eUBsjQARauYxejpwq15/3VMh9VR/Go/8lewDWtH8DBquuDdo6Dwnsnn6NnbYAYioKfUH
m0WDRLjell0u6rHSdHR4AqwVKzimQtqj6nGf+/+mqXpRp2sY7pWaIBvJvoyXdYcA09BGKwaY+kop
17+a/b7elTZKaGce5DWhwzP4dGSScW6eHAtdtlldcwcWrtIagyqpv+FfKXtVB79YNghBYEoeT1RS
B/+9+ddE/Umq3ezLWQYbW5oNKTEOAzDbEaVokiZkAlgMznNeD6CUoxd0Sc6wP+qpDXzNPbtjf8zF
zKqLk2DPEEO6jlbUM8Y/jdDHgj2DS30kBnbUxrHDl4gWJrtnzh6oNmPWVECGYnBOhKpYXd5WY2V+
Q6oVvHa8hHU9fgeOGm16+bb7eF0uIBiTzA9rgJosB92hVoDT+xwSfbCZ6OuJ/gwHVY8UKCqVTo/l
v3CrszNnERMQlQo1eS1DKrfuTPr7r5yaHCdQ/jGqkLRvM3UmAPK3JqIaRuDQtEBFYNPW3Pkp3AzE
PYtQV6NcZrOCViczKMsDLWA4zaQBHMWaclio5hjbHws5NZmV6zIxQuZsdp9Lv7l0/MWjA1IiV7mu
tQezUyTQRowpGARN9P/alx8FHWZX7ybrCLYHa/oWx6nYL/eky7W1pYF6ZGChtGB3iOajHoy8awuK
jYWZhHUIIi4QMcLrPZBGFDfXtKOr/3fwCw625abC8mx+ZWVtCGztKxeUvEeM4dBDcejUSAnlvaxa
khNTIeMJ+MzmIcS34m9ulAcMPDwkE5G6ueWfg5yz0GVp1XREKSOMIG2zlCOQyXwzCSCxH+y5Db80
Ghs8qd6ILzFW1k0ja03vNmiqO5MVcYz/233d+ynTN2nMPQi3KoLIqRIeH0yKZf6s+TOo6mghoxY0
tWG4w69KYgrsRq61iLC1y/yGMg5aEWhrpTcRw33pakOfB4QGcB/hny+16bh9cjBa/g/jX/GzGwh8
BVTE6xOuX3IB+NAqin4r2ZILiZHSwNL7N9sz+kfhf2NwKquyYM9lHiAWcOPBmqBQNOkPGizFA+RC
90dh6+vqOZtqoVVImXO4NaGugzInnXBiH+CnkM9OS7aZLOcBlAq/zI0tQsei96YHx2b3woD0R0pS
7IlnvSZlfensBAEWmRbuPuE3r9oPmPKVvAtsUSvQuoyiqTIFReo5TFdhq8tRov1j1Ibz90wWMv1j
PledNOTtYXQHRENz8JhkIGxZhHgda1NYm9xVvkzFj4Lb+zKIO779Jzi0FszHjSx0r3RNE3BRDZbk
yJL/V6KF2mG8pRNt44IJxjjyaympdq8uMK6B/VoW4zGh3aZX7PlxjHk63LBqf2YLacB3JZb4rafN
gehL5HpmUMlbJrhr6DcSWZmzon0P2bxW5SC0UQom32nk8CCcKOPoqptLGImX4grI52T198ENYp+I
WvTHl+9jGUf4xZKvSauQwkzyZufpLsZdG+LhW6li/X+L8I2K+lwZtpY2/HzwfZTdoCSWMGjQ2ni/
SEGtxs56GWeK3KLZfr6mYz2XbOlawV49ArEfRmfMSUGXJDmQkVLFiCyyRGFQy+0Xlgq4x7yeb20I
s8lKNVD6bTQdqfDA9YTAoOLnSReVwZdEWRx+wdvibcVGjGmo1wFpe7/8ppvdMh0AR1E1wm/Rg3cT
YzHVgzCmgSzp5ysxq93ezrT1To0DY4SIYJgO5IpLaI70qU764nOQDRjFYI/mjdMit1G8KcYoyDbi
vlIcnNyn1uODlWzamxHMT7w7+qOKLWBwA1yhq7TdM9UlajITVmwDYp6uFK/oMK7RJR/9t/1OiFwc
DG3KkSjPUDZO8tL6gjfwpuFpH1b8Xwcc/Hj/Z09fsB/+4klBNOY5xjNFE33VvbHiRO+b+g9E9IO7
S64SfG3ZiN9E6pgb/Fs8wswjSjZRxyGxqQ9DYOf7a+DlxgciaKt3iVGDm7n3+GB7EKGqxC/yCHDJ
DXhfNRdoBo48szxFYGesdVjZ+TyOLV9Aie0Qh7wZ5iGDNWCB/qCD9OdQN82usEMfSut70P7E0Tpn
9hW/i3bC7s/HCy10UeZsa7eX8ELW7nkVJaNgoFp4l7fxXwN64Z+5oNlPb7ZtCxIqR5sxmjCsfGcT
+jbbgreniwVWTbu0Umi8OammhdwHru5AuzzXqvZTi1SSi/WR/V+ARILRAglRGsMR8bheRosN7Suf
VARhHpkx/4OQ7QGKzpuApEuudHhYrifWH9jfcpyj1Fjus1jrKzpbCgkp52pKWp1ftzmB1joaCbPv
vTgql6UoKS+ZmqO04KDJ7faSgZkUqCa2WmOWmG8zWECCv3rRGfpLq3MEa2RBt0Q9mf3vQtSpzLlF
xsOpDDZhDy7T0ZaztdmjG40V44yIoM4ckCF8s3pepsQo3wzLX8iEE0SvbETyU/0k7JX+i9vcgzLy
DTGfpk4LzlYsXTAESFSq2c1A45UtirT4gojAb7FwmjaZhoRQAL4lLgNBXkLFm64oTBpnZTpREVoY
8pNW0HeiaBVGpUXJdLQk3yHEWIRU5vkFLQB9vEj5QIzH472fNiNnrC3n+2dRubX+GQ7ETflxz0GD
LNmrVn/zdw0b7S6AHoItoXxbIwtiL5o/ro4bLMvc84fMt1P4dIyyiySUkpWsCzkc67/SoHJPwxE8
jw9lvqAHCo7Pbsz40/z6B0JBLSqn/lOwVFF1JAP3TBY25MbZM13t1EuJSGj2aYSi7861bu5zrBiR
vZrCPqEPfJcVzOOiC5Qy92/P1F/Z58oa39RhKNW1L1ryN/mOsSJNbUA0Lh6vzu/VLbr/dwgt1Y6f
DY8vjvTAOo2I1t3DOrr3nTejIqjrgaCB/0A/Vj5giBKG65axP8asfou5A+L4IavkI+b/fRZOi7Ek
VMeudRJhKkv2V04lcEZvUt7svarqzWMNPAwjK+w+LISC+4LLMZix4ejfHLLuWCukzxTktItFxzhq
I+SxXIfON1pVUUUb+L4tLejWDRvx2wXTXD5AuE8D3YzEIgHFdaDdQQbXobuDdg1BLW/lgH8E65yX
OtflkFYjknpDwgmrBMZC5TQoOQEjmif56GjZACCif65vlNiKFALLVQgVqp8u6ZVWGg1nzTg1zw9o
UPd0lQJNUhL2ah41oXxkPZ543mhiz+PWX/pKeBSoGyYfdmKTz/6V6G33QbfAcuGTJ5KRyhXPKjA7
j9eFbdIQvF1OrppRkBYCQSpe3TkDSmNqLVyG7/znw4z4cacj95V8y0GfB+cQqOQ4NDLUEO9Huwhi
4hwLYN8KOX4cnsOZTtakh5yj39JQQeiVaVKxh3ldaERuuEbMEoztxPDaxyzp0g/kJ1K+tt11KeG2
UB1leiQcwFbB717Tva64jQyxqtldm02yf2LjliHZdQKNehYazwbE7A/04TEcp56PP/DLL5dPZGYZ
YyEIk8GTkJ652tFgv33pdHAKS1zO5FJoKGzukf+79MPf7n4dNNMGBOJoWjBa7sSAhMmI9q+TYYWG
goL/14VANNhv5J2typCiyawwIXnuEQdRP5jl4z1zSUXeP8DlvRg0HmiDj/GgzU8MsjjPAPIcRa/8
wR2M1I+lA8+4MDw5JRCpun+wbxl9yD8vJz1C2pxR0ppZjr4DwnAhOtt9IVzuGtD1Hq8jVwIskASd
V4qTIZ6KOyX9fXtiMHRnR2Qp/RkJclvN+m+G1xYzKK/FBJhFqQn+wujcmVji2PI/ESuP1sm7A5L3
RMv2RIlLisx5eWSxyvRCHIfNVFGvDBxNXZ/9gwHrkKgSjNTPHupLH0XMebTmpFLawzfXBwcv0O4K
sSVs58A0laz9w6NMf+mqu0O7gaA58IrndDGyBpzSuWnxVIg51tEhG7K3Egi7QAa1NLcRKtY5LnBy
0ZVAqPpsFW19Zwbmux4ayrQwP5UVHUFDyO8xGfJrzepL8aQgCKsnahwdJcN3utKsCgEj7WzJgRDk
sm18Jj19zoZf/rx4z456DkSaxoyFsWebOi7WfI+dw9L4MYlp28n4Q5NdrgsspozM81/sH2E/phUC
KUrCqiae9wsHpkeZL7oJL+DWXKaMaM9bJIYSCPCdeAqkxu69TXYEdXbGKLYJ6kSN4/0HxZn/tR9l
8Y9c3hGfVA5VVjMRn3uM2+2XKggiY+4dV1ZQKJw+o3ke6AXHkkbwhV1nG270gSPefmLK2+LgVokE
Ia6yPFTfDl21MOi45CtujGa5zrvXi5lo1ifrY08k6wyVtLL9SJAlKJ03Man+BUvstMfgjNwptHzf
VcAI2PqmHG7Mp1O/CPy+QtLARNml1HnStPCh1LPiry2VCQ/7vSF3zHudINESEW9EZrH/dEgGtw5Z
z144y8HXoGoWxXItvxaRKJom1R3S3c329cIlRahvY0SY4Nr7qdhpe5Oi8qupeowIM4t4DGIeif3H
sXPFhsn5SZSUjWi1psbovzAGD4CvUXw3ohACHlFDL6dZxY4xIiv/Kg66OawhobBFnTBjbIyBXihN
oCO29Oyh5ykcy1PsIBUv4Z9VjdspbU8TyJd9d+EcV2MKOWDxZwWC681llxZUt2EtxDSRcl1cTA2U
zpC2oGRgdJJoDpoIjy8/HhIsT1Ot1LNvHaeyi4wK8PIq+KGpCNkPuEUVNqvOXu9W7dpPAFJcP+C5
pd61Idv0BrTH7QCf+MM28BaK7hmeFndoLZMzsClGJTpJ3ddYgPMkEHN5mJUjThCjX3BDLDVr0V3c
jnwbOmH0uRt3T+boviED5Oyz+SkQxKiCK+iUUaOC1cq/EbjmQzMOW5cdGDOXZzPl1jzhs5bQ6SYJ
ja8O259uDnYCd7Gy9yxg8aO5nXAJEIpypGLiOaN+tlG8GgHzvWv7CsTeL0iGZY+a+eEcjMguPuSD
HeI1R7d+YpiFwHqh4JONag+xePmCK5Z8U0Y5Qa6XOfDMOwuLOGSJ9iwAY4lc2CKtLfIJY9R6yr5t
uWNvSkvecvH1lFjpI1QPvAf9NASXmgDaGRE9H1yPsUSkuctEj4HVaeHlSXo8M10iYsUXt4WqbDgy
yu6iwd+Xe14UW8+Tj9GUjkBnQk9YOnN+6owCciPySyreKhAbDuq9rwvh0DtA5ac/EgGPNK/35OAW
cBWXdfBFG2FbPhrwyE75XGhf87jbl403agcS+XtHAGDcp6d89fGfibCpi3ka0CpWfdBtNtAS/twn
YQGxgxxBq1UW3ZFOEVX63FJEfizQyJ7h/euHbTQQhk0tEpEJdeDMyQu57glEck6fPegsepYu919A
oNk/NaA/YcQH7w3YSnyTTn29WDRcV8uyk1KKH6Zxbp9s7tfoAOJ0aor030X7EfTmQHYZ9Nq6AHDa
KtQROPzf5WrJunuOgxY9wvFNlk+Er1MbAxByl9uHEyJ0MZfun0DoLzA5okDHfvLXdotYS5YYdXmS
3aVJ0KoClvq+5GZYPFiT9YnfKs97/X1Rwjbec+pfC2pjrHOLI74pKp2TUf+rXQthiK4HuRjrbJU2
WbtJXGYCi/D92G4DqtB2qGJ3NOmnhdA6OK+4rSikztSaL/1W+CzREArg4RuFyZ2M2Tv5P8j3Hfgd
OX1tbGtCJ85QPK1Hm7YxZetosbyZyTnpGuRMM50h3pjT6nmo0oaMMDOkipnUxttj5rix+6x6iNq9
iPwibpOqvbtSE0MsxMsOaZeHsHNzqw6yW2vvJRmairNt2Djbha0pTL+v+35dsqJMScwMa7iOr9BU
GXpqIoMNRABb4aAir/5mFZjNHDb8FhEPdYC9Iq3gL4wVHq42iNnSnBN8vvZIO3m1TBB9s0VB3ZN8
dLQyfxFwuD9ha8MhRCMUwGz1faFevpm/k3We+zWL5yW9Hk+lT9Di53t/e3d3sixD54AejNBy3Fs0
vWJd4tcJNtIxwI2Xk/qHJQ3uEVkcsVZ7Ab9hHplxAzCMe3SOjsJZaGG4P7TGi211x5IfwGW+2jpH
SwSoHVdNadH3Un77RhNlAzCZbEbw9imZIZw0WGZ3lXiDjnr1E9RKwZJK529OUShVo+nCi7kf3s1+
jb6ITiOdVFJwSCp83ylXNoKgZB1xs/AcIox3yQm0NfkoGP3lrMs+JVu7wXg6oTFAp9TdwUKAOaqY
4jTh4wmfTXyOfAAjeemKYO6TwAw4/X0GirqCAhacpX3NLTskOFExp+r81dqHgJ21IM2K+PlA8egj
coimjlJKFUZLVc9StMIak2kB5KNzqql+nRVWOsAmFspXlNZSlQqMovk1G1ypsp1z3/hX9hlC8p1h
HfyvVOZQx8l86tJSeOg4LnD56/LFTQ6TksRWeelkTMY3HPm+ix+epfa7dzFuxHQR0Dy4lMTRzgfa
f9Rw9C35HoWBjsM/8jCJnt4F3ZmONCwS4SgqitSnIZXJjOEsWZpBNfVsOUbR1BQT4bAVvDaVDKeN
OshlQF3JMG8CbSmHOnGBWKl3oPvDtDduTad2h1Cq6+JsqAKArLotvw7v32/CA2kpMj6am+T44Jsq
4OEpjUbmZ+UHXV8ZDYNWpxL7k2j7inE71l/FP3xZ5YNcJipbky4Gr0dhJ4xgRyVjYrOmvqHvfAFU
fFMWf7+N1I55uoZWK0I+lXgR6UwpWXGUxpNiJy+c3lDXrEKtHOnFEwBs/bJXrD9/kHRteI1ROBCC
fVzuhTvKcKzl/tLqwZxfYkFUtFsbp4lSBZ8DTS9ULlgu1kzFeEaYfT/BI/i90GqLzw0gSnAxgMlJ
rklVlUOjbe8q5FIynCHsfesYFsBElKxUyPmPw14ZO4deO5925NkHi0EfCTEJRJMoAwnyiYT31icR
sJu/Sm1F+9b24X7dHlWQwFxuJq18fuEFNWsJAbfGKhEEQoELHjAZNRxjVGL6x2jQh3+2zVmaPXfz
u9RpbIF4hKPhb0w7DoXHABSJuty08Bwq89U7m8+K/O2v0e6s3wFLrcrX3oC3ctLuw6NRISZOeADR
KTms9431Z4zc05pmWNk9OXMp2ujbZw1BOxE0Dy6LWTgzM6RYyWZnO7dK1HHgyPIi7QO16W++dlMU
+J/nVV5ROO6CSQZQyJlvudBDDKVrJHF2UVucwpswStf9qge6eOUPR521Ytskfnw3rmfxslQnYbdl
zjBtbgkSh/lEUksgLLAICSrAkWz9mf/3VaF39NR6Ml9NQDQPxNzrqvZ0EQIJKfVJ0ljz5N/mucsZ
CnmcoesuLboMCfogt1blezJ7Dm7QMDkVw3vhYV1RCR9m1aHXGwlcUevTOwwrMFAg0bkCIS14/iLl
ED7UkMgLlbv8+M7/TUZikshNtaU2Mp8VUr+y7HHD7wtfW8wwTywv00juVjeDXrXeMuSj9atVy6bS
z7HnOxXkwZeyHL9wmmULFAx7nxaWHKZ1wIv1Rk/wVhRDrf2Vy002ITvqEYuRHMMXBugllcrhEE2h
azJV/VKKVN8jIkh6epAcPXMyEgcegTiPwZFf7dF4/PhXx+haCRJhhr+h9rDUY7XnugnH+kLXQqt/
i4AbPyQfiPzIAj+iGgJfHK/Vr1IIAdCorCAywCBtvOx+0ctDBtlVh0jmnKAM9RAAM71SsFDzYQrt
I4XhJ3lts26JP+aqOZt+8HMrSKBPkHMQ69Mx12RzpXzzyBz0CYr6DEJdrvQ6yIRYHmU0jlD/MjGO
WQa56vKHuT4jAZZGT4P3SfpnVQBVsT0PFZ04UG0kv2UJUuFs6DW+rul1bLqRpnIWFn6bfjd6o9Yb
ireU/Ut0W50CP9G7GPlaRVASbd5woAthS2pGBlOYJpgnuE+dEPxoPGUkTWlwVEZkACiFe5MGg04m
URlErYNiWZRn2GK1PR+zqkD+Pv3M9NZFaGfqC5gT2UgyPO4947Kpv4pJjq2K3PxUQQL8I72+V5mf
5K50ZKUHRwuzvxW/EKGPIxgF7VkAGmsr750l1AjCJBUNEo0ZC4S6t12QoL/ZJj6hMYco22iL1RHU
uQvRuVIFTfkzMC6wP0GZ6XncWyq5FAUs0+nBmEv70W2tdbpCqpBE7jZqKW6hpZPyD22RPxYww7nG
sWWzeLBO1eL6GpM82ehU3XFZojmxxHDeZulKdbvdyFJt/HeVHTP8x0S+neQBr/4bTJz+Pkh8ftW9
BzQAm7bbH/+2oxkevbg0fgoZ3FGyGd/QNcPRnSuVh4d4VmnUEItZbavm/HFR04X0GlXnQEsZmNlS
Ahsxw/S9gtE0Px+7M2vvJWMQEXRggbH30DClZ2IlAc6Yw0+XmYpXKLRENCkQJEZopHuhAVNwbS5m
pZsV/Z7YEKAZqWjvbW9Na61fMbmm1YPwqogfZcjMyvntxIh0TtKa0GNlOcrKhuOnh283A42b/Fnh
OXOn061ogbzOymya7YMUQwLNeQAxnEbhhYa3szjWQe/wFiYAQM4IrK2omOsY6t/qdeOwvK/sm+YD
1EvaDp06dOeBdZ0TOlzwvvMVS9Bm+e4sIMceKyydSYXg1nlGU8KNCEWl077dbIPWn4W//xN5o07/
ffw1HwVsip2wVAyNdic9zJfIjViHZUHdlPwYpQkvKf5T106xMPKAMcTMlrxWqf4wYo3trNTdz3+L
HLJDMJJfKKBVWPJFiEuwZcmIeJLE5CtKfG3iIOZr4dkxUdvVph+1ZL5/OVhtiY69h65lGsIMhKnM
XlcOb1wdytpbFY3qJ3WC7e8AsTM8Ttwm8LouEcGY4Kzn641e0WfI0bmHnWAt66kRDYINKRXNTR9G
GsdHbynl7VhTrd42MaJNBx5URArDzAMUV8CHu76JZTm2dI2SGUmSuZLTm7PIVJxAEdqN0u+qluKD
Vvst/l7geMX/1OmpPszETZZOP+PlHoomYI4otAs6lBIc+FnpM1FA7RO5c5iitk43rzt8xsCOYnvV
HU3lY8X7+iqK7faUqdkFKo6f8m4jMBFEmGptkY03d61Oy/fnWEp24klwm8EL1wDeoqp6ZS7V8hy6
JkTvSswLpe66HZd4J3ddO6sPenpmu1VQUeaBFu717va//XidS67PrIzDISfnTLwpbAfBsdFUTRDQ
pWhjYC8J6hHQCGTtVh+CMAn3QCqywh25DuvAD+NvEE04u9FRdkw6cWoKA7Pa8L8JSS1VWZTlPHaZ
JkltN+I9DlB0K5XMqWyIWcuRsKGNJXvFA35X0injV7rpywng7QITENUAVlvm0obcxPgbVqWyAgti
5lyOPpSYQEcnw0Em5e5F3CE7/UCpcIhdCTx1Mk9faGdzFxIrsYfQaMW+1WprIFosexMT6LhIPW84
HTxCh2PKHJqXgN8+oaAGGf4jsqzfDmm25PgrMQCh6gtrQdsEGNcIkfaBsvYLFtWsCb6Ft2qQIomZ
UqTd6g5iPJeow7Gf5eH6aXrDdF+AOgC85YB+/E6o6N3+8anj+IA5HJIWW09fVrMUGVL5tLS4ewpl
THYcH0+kuClUpFKfjh0lB83SLmEByw+UGB1L4zPywojiA8MRa8NCuVlVp+vgyhxEPC5ycIHWa76a
er1skAVtZ7e94ab9LKkL5O9Rb3006J0Fdf559zoa1LF+ECXRlieabbU2J5LSenk08lYCgy9+ssp3
26aTl/awOo/Kau8bCihKhMOJ1al668Ctxe2XUqHJAQYKsFJGll3GoCJSCl7Xe9HARKHKWtJuG07q
BMQDRrOnv+JQCtn/gYPkoJ3+zAOjHHkLROLw/uZ6iOwd5wvbNoiSUVhvsojyO4BkSabnq3FtzwbT
LJweAIHmVzSMmkOg/OeaEq2FJHbSr6tvZZzJ/kp2nA4+evhSk7eouezplwuyfwlowselk+z5Aba5
P+rkTvzIOTkEgKq7hyQeK9p2Gij1l5vc3R2W5pzMv1ZiQZpTsgjP4RAmY3IqnDhwaA3P8R8cjgGG
G5yR6MUBQupFHilVoEFLigghEGoIxzhcH9MAwJ6DtC6UF8JE6P0ZaENfV1WERwJUAv+/QJl6+a+H
nEp/g++ZzTMKEmmt6EyP8Up2n/im1CjVkYYHeZh+szNULmRFW6lTIxOyiDQMA7aM05Px1bcust9a
YUbm4bX2DJ49uRUvWooXfUg63h6ecJejNJx0uMreyhet6nTJLHCoUqEeKwSybOw6hBT6bEJbB2rX
6MBN/V6av6t8Q7R/LDyZfDq53l63ODg8mZnRU1jAyc+hnAq4uiOD2veeEoP5K8RMcZxlR6THVrIe
KZgNtmeQhMGHwFzLglxjWmcZSN1PRR8mbWioj5Q4+FKOyTy+Vb7gwcqS0H/RPkxb7w7UhuDbrV5w
vczv6f+jYKE/KeJgx/+9KEJvNKoIwJtq98mFka8IrTO1yI/7CuxTHZOJrwqlbPzDc5SVCkY6Jzd9
Q8kXswU4HOIXW8YbfvQsnIojCwHV64pxrmQsaRX/v2novrpIkVdIAp8ZZKQqe452pG4o4pkrXT3N
K6uhD9YbN7Zi00zUCP1Ow6/x9QSHCwYJjRx6fW+oJ5EkSipMUcCjUrU4jLMhcwBeftJ1dGE0ddJ2
zthsH+vZ03H9tXpJ7Oztz3GdRZqyhx0aivDn45CVtkWmSYGDqNUngyB119uz+6o/M4p6tm56Hk2L
+hApSSOGVttQ2h3OWxri7q2KgOkv0GliLN+U6w/8h/Srcw6g2vlwBCxlu/pR/U+Bve7tlDzQ/QoJ
L5U416F+gpc1RByElTk5RzMhnNzr5+/+PyWi6h9kW0xm1MiCuolnqU7TF/AeIwnGbbfEoJPPpHRU
8TXK9xd9hhOwUEIE79A1XI8nteVuR/Z2QgzaIiXF/T5G5h68+pX1PZ3kBVGGTKmrVrWkcoa15Ts0
DUOz4B1OaK7v127AWDvqCpYvlFdD3yg9+KBMqJdeloLacxNX++o2FsKo3It1tzdnNJ/NIdhtCRpg
QIwlwCrMpEq9wAXwXBhZGWnbGRdGU0u2CcU5UwXpott+AO9Dj74PnMSFnATYxs3g5a3eHyoJCf08
kHGaev0p9XT66EDSLntzIaApCD69MzPrLh/L/ORW/uGP0KMI3Jtywk2frmocFP8GhzJFKr1nEmYY
9yei2LxA8ZRAXDRreUfwUe5TZaKfbQCxQtLKW49ns2YiQkOsrRMMgKGj2FHsD2DqcWGiiLKh4hcA
3XbprOzwYV0uigd2ynzJT1KZ7trHYUEgmxyOWcdnQ6BBNnmbvIaSEil046nGY2O80BgPSwriYx83
RwuH/loOoQRXcJM6RH4KH05oiBRHTbD/pCA7bbaIIHr3cAYtLTx0sXkE+PKWv/BtzA0N/UGfCtFi
jLG++r/06ZrHxpHVygQWoIUaxslorQsNL7g1tJUbjlygONNhdNn1VslA3MtFHDfKcFlquQxX/JLy
4Ny+VfRYrszwLF1D7rpM+7tvgHGANdYVeCLnml/MBZ4CjVo2quQ1XO+3NIF1m2PB9Sw2+q8DyH2j
hkEDY1rBTSGJtlXnx84roKJ7lNv/Kqr/hTzmJuqTmXgQxfGH48/LXUKKa+I+tLscHRCpisqPcB+t
yNWqnOSwnD48XWwIU0/0hmPe7CKht/uaEPXw7t2NvT21qEQVzPvFt8G78AxXBhiWf195sOLVralJ
ALNPNmJmtUOsTHUpML4jkXWQmkS1udhFuV4XiMpP8h5A1ilTAcYBTwSn/YX0V2gxmnRn+qOY6kWc
NjWm2SgLApQYfY7S3ADynWAkKOui6jIpHOS0OSn8UqSGuwX8tskiySGY75KdV9eN8YXIRykCa/XE
D8po1kBftti5M9Evlpu7Qh4ZIJVaXulspxIWmZwM179DxyiRYr6hLwxTAzI03nWfgsvn+uVWD0Dv
02W8pBjKQlDvShKE+q02gP1rXDn79tlgcAbH300PmOvEs9dN7v4bFGZjWQsjd3PtYlO3W/up8fpS
0Mjia5EPLQlfPyAriKk1E0/edgT/WSOgHQgjjSbVr05fgA5XwzuYq3U2bsGst10/DNWyLqNYYOJ+
7KctrfsgkFfz1ii9f09kpASUJaKYwR4sJIxWL7+ceulFwnQ1iwY3m15JqVyzFzcLKOFiNYuDl2+P
7tFTQPVV269PTJsHVOSQnXOcICwUY5MDHE+SYxi8FAuZY4NnAMdqrAu9MZqeQkgtBhtYh0ntzZMD
CPUvuwl60kUOYKU7fqs9n/vb7sw1qM3MYx64SeUOlGHgEAHQ7pfeJC4HSeiZ0I5XNlbijpIXNMbX
ScHSx/CGbpnU4iKEzU5pxaZoNR471ek2S68ZqoI19B5cCiVCIpUaWn3kBOkahU6//AGd9NxzeObY
Towes6jXMNosFSYu9EG4glw1wmYD0+e0xxOCmf/SmUKwjg0s8DdNQctiQYumEqeRpoD883/IEOUr
ibmCpLoquRYvNeIJRqW2fKGSRp3qg7D193w7i3mjKvPnya0zEuDQETMD4j0ox91NiYo1TTnS3Keg
8bt/oLOz2Ife1PlNZp26a6hwg9hegv7AGA467XeXStFarnpo0AAO0cxrw9fPt4Irj4KakZFi7RVK
aYTsmiwkuclNeu+WEoNFbXYJ2MkWmXXQ54NiEbxrY08b3fyYx03t6vUHQtwIyJA+xPdNbDo6e/Tn
/YXn7H+BqQpragB5xw6tYgqRk0hLgosXfxPavesVhywKUQecLjjlxralD0V8R+5pEiSin5KckOYu
B8x7Zr2HSjPQkjfT3EN5/1lsIRr1B2Q6ySG9mMCfkdw3zIOez0HLh5VP2S+fTQdXwdJGjNxukcga
N9euvCRJuCjyl65in3N5ej9pVUr95XAEyn3d61G3xkZIPkm1/iX/Fqkbi1HyS2UAqlqDMHUk/Se5
xaXzwpkNoAh33k3jF9m4vOIEtRSznWUar6prhY3RzJiYtduRAigzmsCJz7NdUcgOdQdX+6JtkVSX
rfh4FuFFWE34+5IfYwnNqWLcrYuWZMJJbVDys1KmU8m867v7OZK4rBbtg5TNwufklEI0AE4M7xGM
a5wcQr8+3ChNlHbcKpmE3PpaXrHIC/XEAfwuHFbGnGyP0THlQ53JHtpoJk2liruDTWdcHsLL0mka
CpOH2ias5W3otMnTzSjQNTZSPayN6LQ3ihWXfk15TNcyzGgw7LSAXfhqtep8cFBxsxOVOqZayy98
p454RkhSg5ymCnkzG57lHvul4nHOts2gRVQGZwzsHm6Kf5ihoByinZpfLPLH9hf7nc/wLBjpFGV1
TwSiN1wUaPtz61CUvh+C54Rg2is3m0zCZhE0UPL0K2mfEybqp4u8IiJziNTIq/xk9eGVo3GX9NeE
8mjRenkZ04rVLQCZvLa7FRDgc4kPnLLG7oAmVEWAkeLfHzryTTRhMd3wtAra/4yIhQj7RvUeN5RT
Ck4rgBxpHYbRQhNIzL3KXmZQwnqCN7qmPK7FVfdfkdrEntE+N0QxHbwyxkzvaBv6eplBzXIHIQiJ
MeZZRCcy1HfH4Da/waSR2/8o/sGSByVnaUddHAUmK25vCzaimBiim0mrrYmSyS5w4hz7TmxR4+4g
Ya51WPPU1rnIlToSkcpgD2ruHWQUJSO6QS+xUlKELEU3utahN+UGXKFXXKUHxmddsQq7PJ7ycMFH
OuVTtf+K1TQVkUko2nThl7VJZQTP+tUt3xl9c8CIksqUoaxYOh1h7egsBblTvFfnKohCtP7d3BBs
LGrVVXTaBfli4EQ+RosJWr2IUxAaZ1ROrlDUzl4fvpK2tkQ9ElZWohAdycn9o7K9e8g/8uBcwqKa
ei8XgtQzt65pV5Q/hoV1yOUO/smywC75NsfTSafWyBxs+IPLq3U+frkiDkkd8vDx6kMp2mgmjkgC
BHsEv8Ws2tQpCqswHS2lxjWjdydTYhh7Moc+cbgKJyLSYj7ZYjXCewdJ+Rx6eOkYRs3wEWj7fz/S
nPq9wADnzxwYqD7Jre2ojA8U0/cqDFUpfI+yl+9Q07bgk+QxwFiKGsX6eFxY/6HsBMraf7vYT4ml
lVAZnwH3l7kfUlj9siehgk0IKmnQUyfDBwCWu5mpCZv7P6As3/XvMQHI82b+ZN68v1YliMkKeBoS
EV1HTj6hf6hcMqYUUahLfpPnlrD6mu2FmVvHNVHBZy56btq3dqpjqzV4I3UP5E0iY56hfgV27HYI
PuYGnYMJzrdCXEwrMMhQX4Wfu5ouJ8aA75ito2OTEpVn6s3ogTRJD+YXdJcG5onpglqiOI5XVnTX
n2cQmzMtDXnBd5DhoErsQWWPahYhloFapJydWF9i9TtVwgpFLU4ihabPAPLM+dvKJOeKFByIN81l
o6x9x0ljB0OtCiIocIrkSSGJF/RYA4bnv0RiyK+PzxjrF1D/7DcYyJYzXUCGOAsx6SkybKnmOkT3
mVxRxVpZjxUYm5dV8MyZ/oS5E6yhtAmOgBcMeUiTAOZ2ghFEmrT0uZqa3wsZKsekKLLDA/d56164
vbYpU/rAScazEGQJprRqrKC0vZLriPVbcu5+oQs6lc/ffaR8puazuADRzZJpGSQsZ+7lK+2UxR+m
CFSEM7Pi9AUGgHAKHAN2XoBqix0+lBAGc7wOdfMbfruYpvydg9jwca6kKBLIHWWURpKVAZl53m5b
rjhTPgxpjTSyx0wMv3FWr6ZBCDJlukrnwOfFOgWWxSMxV7qpkscw9+zcdVHM+DXkdI+zf0HnppZ2
ao7m//2BfBqnescIz1KX40VjqYIMVGO6/Or73A/o2gFGodG3TCwaNE2FnxyaLYTBibWKIn8Ym3uj
2kok+L9IxyWGT/baWzvjRLEMICrFOmYIv7+ddsmdPIw9Ct2eKoek/n1QgahC5TkpN/cwXbaesb+r
UBj6S/cCcdsC04RSQ17jw7y1z4pVbMpTOv1dHWCc0U6j0OhrzUBDHqZO8z3avIgypS29M6cPySnN
JVOmUkWmYokglA8MGo6oURcTSgxP8wyGd7d6tnT/v5h3qmARV9+Wcdwys/R2HRXKgb5Q5Yvs1q94
zgLKWEAkWuOmuq0hke2SNB6f1byRmKXIwr/GVqgIWSp587zc5Bd8jj5mHK+x6TP1hwWP0UDunSNx
kRZxJUmbIYz5cBu2fi/wxq4PQnrEMhrptJi6pgZ86x4Vx/6Vy3sZILqzfS9iwd/CgHlEdOZ1zzCE
G0uayoGm/sNDW9fSb9RCPQDZenbcJs4A+bO2Nu2+SV6VoVjoG3BfLo2SGSiq0tzY00pvyjIyprjj
2XE1KAShiBdHp2SfKsq1km3IxkShANB0HNc+yCbj6wDojOp+BiaD/y26CNLXiSGZkSeDcYDTinhA
e+IjZf9hMsvmlOPQ6iUhlwGJE+HwWmVcwubWFhGoplNBW770L5LlY0XNDhbEPJK/h2m/HmPsOokT
9CP9nNe+NbzDbBvBubHrf+iKIGJ8ga+/GblTWATwrobqyJZ3EOjTVx5O9j6gqXzJL5GiAODyJ6xe
lG+1CvS7cp5WVxzDhVq6tTXlK4zIPEC2t6cKO061Dx4BpvJkMzPsEnPHJP8BjPpC8g0qgoHDNbaZ
yCzkr8ujHsPKB74P3WMMJ1xhvULPwIqdFERgp9wxE/5MgPz5E6EJ0B+WrIgRsVZ3+jW0X+krE1R4
kLZRbptM9jkqQ3L4HJU1oorbeoeX0c3r31GXv2/ski2GWTR7Z8gQdIFhKyXQFK/7xDWac4CRvJN2
/yz4PwOFTtlsNC8q/pNp++uvj9LjDujtYwRK3JsAi5QCHtrTqOXRVjdQrVp3m3f7YomwDvDg5MSq
iIAkDL6WBMvqr5z6ipueCZykSTUnz8/Be6MiUYZbDdQFScCeqkqOE/0WG0w1L9wqX7s/rKbEA+2l
BH5fVIYycxrdTMcKGWoYTu2AOaWvaoR2xNwljodU1/ccDyyb99lyAJjo9GkbKM9yxpnuMfmVateD
EDAQkXwtWWrZK7LsbiwDlOwrQgdD2v5BuRjSdz+Inoc9Ulz0vhM+0XU+gZ9CcJOZpZQMARQB3ptH
wTY4dLcxQOzO6fD6+OKcRMqA+WNtgXK8sPG79ba87ewTdueh9ffs5ypoE6fxL4jyVCIuS3/XObpY
ztu8ky8J/RVSk6Qpt+rwVekCHwvqQVuPd3ChQICOqLSD46x25s2jthNZK9WXb7SJlsaX4JFZb9aW
f3NWvC07Ld56Qpnfh2MbDuwOtWZrBP7OddEuvXkswKTgHGvuU/Uu7LXmFSwommQU94NOnCcg+X1L
yMwXqXWL3cHkz34jhJT7YL2i3q2lwOIQrWkRAQmTlxyuw/2/TKLZl+d6PGPrpizV+S+WqG65z6W/
SJK/a9o3GnNsKCsGlqva0H0njujyDCPCZshojOtT1nZtapmXAhWPz2pPuWefv/TicPPLl2kSVvJN
rxXz9G34Dj9TOLn6ap5jxcxQ6ygmgvGqRctJ7fCqjtvpl9+L3W1K1pK+DaOkwgWp3/YvNFTbQil3
QwJZMgxGtHxskF2XMvUxVFDp+CJB/gizMsLSzXukoh7+4Za/kv/Q9O5wDvsCJ8a44XlxCbJWT8Vo
jOpzKA3iO65NUE1UqDSMs4aVzokDyIL8OTtoyzVT70+VmMdWPSRz5RkXOw7M65p1CqeusCq+qVm/
abZE1c1IrTEw9pimSgq87vzrrRED24EheMQdVdel5nYV69sUqx30qiiagb87s1U/9IIiWI/xRqc6
6suk0kvFj7ssR/+YNxnY4ImaPb93+x39SeUz6CF1El2sv8yLanA8YeKVPP0UZ0EsIH1vDAhMfTn3
xT1mNg3BkP74hDoBZ9QfNth6f0rDDDJQlp6ZVK5+1sQvvkotYasA6GtCCGOJ8NFM5pDmRVglRl3G
2LeKvLtxs5e/uh9M7L7Ir9Ud0xMa+bqHB7Rt4y8aT/yANvfCaRCtCjGE8M6tU/9hLRBhUzXVym/q
G4UmRL8NCpRSuZREmaNl59QiiwuUVr8LIP7t0ekOwe+Zt3M6mCl+oxL76VAGUAQ+I0UqAAGufxQm
BGYA1C6HNMD6AgqF2LPfeNa3kz817hhM70hojsmY3tGuBRYkbYF3EVv/upTTQxFYz5LasUxY1ScE
e0GbBVqDnVmauiVEvZTg0uZYBLkAMO1sFoNDZm6MjfUiiktBc0ms44nenFbqu0pEzfgl83Y+pmwK
/lFbupwBos2IGuys3Kz036lvAAvoM2MZ+4V5gFYyTRIgiTrPSFpZHAjejborD0wMlyM+5MmA+vbV
A0Txt8F4y3kyWa34gHmem4jfnypfSJQdcqZaSr3QLbCwyHX+RnyTPEngfGKWEZX1zXGDGfsoA+02
U8nsxggRNqb6IweYnwmJAPepJffUA1OosTPVBOItixIbFN3TJbu3Uc8TjEQ/WgxBlObguEzjMX2m
BTV69GX+TRkQKOhF/mxb+JSvJzhkVnVOVmeTeSeE3+qT8wspaQFz7i7Cq7fnEq1vuig21vIoNmce
depTqiYjlJ3jz6Ojizox8eTnIonmDSVPS95msTj9r6ZFECgCFuzniE4TpqvCu6CxIMDSX1mrCsjc
UpQaiN71nVRT85mjNDB/6QeZe3EhZRXqbssGPm0QiNVn39KNgDY/Qnb9k/0SuUe+eZJ7tysTkEiA
VJLujC7+ttEYo7HZ/KMJmDZJssACKoDaef2WxCD6a/JYGqTrQG/8KXSb2EPrIMkFjZUwV1h6VvLJ
ADqHHIsxtYUNWcezbmnXLnuyPmLU17nkSdL1dnnfduPY9wy6MlQrryjIi1oV4I3UZKUQz8lYMs+z
LgXLtLoVYKldz3AZjvTjyfdkk3A31s1a6czuwK6LFwSMw57MDxcHAcXXtk4U8nXm28yWSZrnNIFt
yVdiRYGGRJ5xP3RtE/EGCwUojoHUEhiP/PN89FQHUGqfra0mndP+pAXwxUSG4bf43goRdFM8uPrZ
4Xj90pbkpsge1Rv9zUUAWhkOjveNnUYg1hjyK+PSp+q9hn5uHqU/dhGp5P8A3CAP5obNS3e1ifE8
WuiWgJKgoWkMugKem2DVVwrPTuh2aXnw4WZoJU9Eqc5mfKSYmDCyf9C2+CZxLV2CmEz3K2/KdCei
8JHp6R7EXd0m6JzmTrKa/3m9vD146OjZ/Axoor9ZwLXNQTlCoy5zyTxpbQ0UVawnr2GDrol9xnva
K9/yef5UdqEqSiMiAgfk4a3VeXEQ21xUSMje27jUkxLX1X+6AzZW3tqFSPfxaMbx61oGg7hmRYvR
v+1uGGx3c/g3a2fGFHZkZH7PLMFLAD/UGNsM4zj79QmI01SsOz88DnOFShI6beycDUN7bV4LLBZW
tIdYhkpJkc36TyTEHKfF11Vh/TJyWy0BTkWmFlSAx1cKdcGNE4yVVXdxel/+e7FghtXcwwAAvwy6
JXoCcSXDj/QLcHk9Uwr30sknMW27fToRvHnLm1Ni8YJfLR7pia4Cjq/Pv1vlMH8QAc2ArgN/0AEh
vUvsKU5P0pNrCl26ppukyiN65HoaBLfRx6q9K5ZxyuBDZg3nYveQn3ZiPp6ioBw5lQBnBhgO2ug4
JqTXOeVfU/Uf5rRPeWKTH/uW0PeLCpNGoNleC4BVgUkzjoqB3LLPygkux6ZPcA2ib5L5miCQpX4J
82UGepZlnUHsnKX3Btg9fKvsSq3b6rWKmIKSYGsyfzPnI9ZjHTf9BgMDIzQhmlzdumbaF0kInH4y
JWFqvJnkvMlso8miWayXC2vT0Zyato7Yt8YpA3yia+unWwdKDNT1nm+xvRuMgtgeOCQVcTM18giH
4uhYKBXplJjSfjUA0TsEBSAlF4wUXLGkLScO8Xn21exVZJ7WgfKljTr8sCFU6av/l5DtktmQOwwu
ICXDmryYl15emLgp64IL3rGn1BRU4vB4A/33Eevurs6IwGuY+ny9anHdbiFC6Luj8RdFBT34AXDX
qJczxwLQt/joJIqkxGTazd/XS47N/ODHItD0bndW8dO//PPfF7azb+o0CyBZHtURxLVYu/B1U6Q0
oWKXQhdcZ8ZuMnHF/MoZt6BrGKyAN1XbUwes6a9xBUiZeXRuHUWt8LQ77BqoP9tyeHzYMb8DJe7Q
ualUuhJ8l10wxcEaRUoFNZYFkY+0ba5G8IYkVKTX3Oz604lU+Tn9lZ16YzG+fH95G9SRhG/Eb77n
i4Rro9k5bHtYbQjc222uBOr9Cd32of94IA0rpOEJdIEF+qRvixX9gCfIaCUDowL5ypdDGM8JLsJU
gN5gzEfos9sBGbMkn6s8a+kKNzSihuD3lQ2/v7YKrjY/iidqqnDObM0Zw4Hm1JiZrsLSCf3rNvUG
sqVIPVQLCjwMOSf9y4ewVnbR+vUCjSx1aul7bzLrFbTiDqAEPIw1187gzNhx8wXA5qMlX5U7O+q5
GUayWWGqKXx8Ib0+LKAUi75T9fukAfc3syGqmDVtGm1wdneZOBUQGDHE3MrgH2j2EXKj1Vat85tc
OX9Ibmgh/DQkR8vNr6OWvaY4bEfdahhYAv7vOnH9pThEOiXs1oJbXGs2E0qkWCnGfk4/EHVm0wSj
2095SVOwFsBi2vb5+KjilIQQ9D7hfHDbEo0mtx3tkuYlwDjAWXS+PE2z5eaXggPWEs6McLOSzWeb
nzdiDufhH6gM5bptAWgU/LqLF6M3O4oo9XaWlEhe4a9KKFVCyR6iuKN4IjTwWUS/LDzdLRnVdRJU
XyL0RjHYvEX0m6UKf979Bc81/hO/4yrOQ8HQ0J7Ivx/j971BEFFKqj131b0n1wVCgVsr+G1/JZgF
Rrr8xmLXxF5y+X8VhkBItEE/XMUdHZHg3dOozq6BKje5fpAyJInWvISwN4Ool7rVfNTAePR9aFln
9v441nCD/e8jjGYncOQ1ssNSXoYw7NMARDJx8cctwq5J+dNJklAfMpAdjAiBPyRFARCCv0lIhk6A
KGgNWkwvYqQzsym5l3u7+JyLeAxXcUah8lJZJ00XtQcC32wfxsRaVjktD5Ugkb16G48zKMk13aLk
n0aa9n8NKEszgqH9jyIWyK5IItKkyr203arIaXuW3flUz+d9A9pwIR6EG0eKpf+2SG0qplhTESNc
/oQ9B3mR4+duS90yk+cOIAe3H80de9LyceKRRJj4WwlqVv8f//EBGaUMe8ylvLjF4eZ+3gx01H33
o/mOgrT+nMYiQVVLnJ9i68D4RM+bzL9S2EKQ6sNwKzUIkiXt04nd2Zb5N3U/7Sab31sNQRLiJXV2
nDemUaPtOdUwSc3FIaAPp2JS9H3RA0HESflAIV8DIKUKnkSswf3PDWMU91rIC743cs76G1GMLPx6
/3B9zNgZlRhtzX8CmiE26HPsvcO+KEBGxGOqZVqCgDXA+mH0kpEHYkFfZzEdeHf1k5sobEu5ZdhI
d181OHLXFVYtQxzk1NELCvSqxJmfVWHbmMtXdkM1p7y4wu8UU+upnbRy+CsEcXsdrkj8SmZ3TLxX
u3GzN9oBldYuqJrqQvbFx0QgSIutXNG/kqeex6guSNcVeQuNlETeLdCLLW2JMdopug+NhGgrNORB
UZ644zaPYdadC4VxYMHPIgDwAYzsm+LPq+n0ZfD+aVUXZA59ddh5J+2ys589V8kTFcAXNg0B7rbJ
GqKOBB784vpGQiTbT/z2FMWVrCsSFRtfkEYtQLLMt/bnn+wukZ7tAOjC6dsDUI3gWK0jvMxozdne
h0ewwPchRS4lcH+NP72dnRNAELUIfUTSfKgBYis86f+ydu2zh2PWSMlPJ7w6cLWz+/i9zNtQotZJ
rmK2bRFuFP03aMJLtDT/az14oFRmYc5TC6Q3jG8ahP98+2FQmWdbjQaIvTzVljyTv9gOMnLQQIQe
yDkbK2S2Gc8e9dws4OB8kIu+yb5tZYAiVcCJUpk5CCFT8cfGXmkYGRfmqvfgVfonYieOVxbuZlv8
pKJLdPtbbdDop2hCA3AaSgnXdloQZHdWkxfcF0SQ2IptJL/f5aIvS5BS1v3qltZUsLlu8xzJYUoi
hvrQPW+DMjRxSRHTsvdUuxxyu1fngltpDWsO43zdFapRk1NzSO2Dhii2BO6FIYJVVxsyRO+yBiK0
IZeIKqPQ7Bit5s/limbkwcO+rT1Wl/ERakFwfMO+OFWMAbuze4r/xl93AhBKoqT+eU6DbX4o4RJ2
1608kdUJPbUsPBJMPf5e066CAN4t+r5jT9W8c2c0QlaRACbTFMKljqUHcwP8NOMGM6TNW9zOKpOn
OfeXGoxUw+bgGOYoCHrDEumI6UWfObXHbogNPAWx5cOO+s+KRER1uBDFDIi4QVPAzBqxvez3nkXe
nsw/EfJHzWdV97QxGyfs88O6QeydzXS91Xn7yRgJNu4iET5Se+i8JhRCRvFYygmjqt4OkNjdjpJo
2CAx37ss5RZDNy0zEB6bHNbnlelcPTZ75smyApFVBx/2rd694eM2VBixtMsuuOaHQijjcSwCKZh4
C3/ulTXT4zdaSoVp8bX7ILKP8ehclkR5f85jhccmn18vt13XibtAMQoXFHgSl6GzOhC/uQc/Tq/u
nXmmVG2xQQ2fV2qmsT7aVVfMhXU4gbB4ss/zlJzEbWWibqm6hsx14MXcVDpfllDnvIT3PnitPKu8
vtoanM3r0VbiGZVJG+clSGAwPu2zSNsT+25Hrpz0Y0mHkc4TR5f1/30Bz5rzWQwEYJ3CD2uGv7PF
XRFezMK8mVtuOUcP9RpxdQ1tloHdRFay3GlCAf2HTNIn5KITqj1SQOZBjgy9sFuCV8kpnqw62UsM
Q9iGO08hR+P6aoNrVs7qk/abgpEGylBqQ2Z4yH8XFpKGIJisjVafDhOCkrCeiRUOXfaeG1jinbAE
oYdD7zzJ490LxJu0tii97BNyFRIUYST7+MlAZwWU6LHWbnwUubeTEMmrq6tep25L9jh3w3J0Udvw
WX4IVFceQfNR0fZQ23Aefvvti4kYxti2r+Ya/qQCQaX4iDpqjbDatkdc696kLYc2GIyQaTU0NwYR
70310MIeNpRuMwHa5vSCBfqAOCk2NcaiQqZChokbYj6kJyOAtY0dRioPoSlG0fQ0+00DEvKMp7Ue
ioqIAYtLZR5CwGWltLxqp4+tQCgPQAhWJnlgMy0L3Sw6JVbSRFQYHuIyIFg2FS+W04DWmXskemkc
enHhLz7gQ3CQHryZli7JhH0nrhQItsyg0Xs90z1xJ3LNrjjpycbjxbnX6TT1aioNqrlCWeww6nyf
oQdG3PDEENQmWFzjG+CAeZr0L31DFOUFUfAzkU8MZmITHvniMAjNkT5x2p42ksGx7lsaLE4BSbWp
ouYlXmwuqS/lJVir4Fzo3TSCYQbi8voQHTJFdfJAOFhqpyqspUZLk4LpscA6bVEMRT8uS/3dVsQf
aa2008Mmwz37b4lRcUqcG+cOm6zzPAJLCIWrRSP+88C2qWLEdEcdg7Be6D8QPSLcmsE+gJlLzLcO
KbucLiYbgF9C7A5CTd7AO2kd+yrTgfszFE33DFyk1U049KPhL57Swp/X0cnDCeJVk2wk0Y4Lh8+m
g6VeCwitpKzBHODVMTUbNa1wkbVdHLsmIWISMgnSR6JLNiZagpLsWf2vsAGKyq23rsur6vNAEBDU
nWqayW0kjOQCNZ9tA4erfOfGeuQ1qfa0frcncbQauHAiIxelyidhJMmx9+xRVM9fN4VxEaSLY6ah
PPqxRMmhkblS+1uuJFWyiNxRcgVag5A+F+9oHudlil5VzY2RRXZfaMUVAmpo2N8kKilqGmtcOr8j
a4Ag6Y48u6NxZD37/aIAxcCIOvI+XZVMEDvHXhG1GV0nRzvvIXLI6dE6zlxz4/2pLrlVTOp2Abxj
sAvB0bbzuwIzenW7IMO2c4TrmXtcFqM0lifQpwUgSj3EOozBo1lvf/qCt3sFSRTSg7OBjKZBsq3G
wrY+6+KjaZfMScyiTL4V+6nqZDbARFi3c0r/McwZKFCct9MsWbq5qR2D8zpqGquHvaQGVkrDOwwd
ZmEC/YRgslRI1fXN3D0xY/MBKWlzAui+Is3Qs8k2VaYoRReGn6Yagt9OMa2IBDQB6hOlibyqryFf
195wQDN5rlUcGvEfZlesq/fnuVCODqwK6+MyhPj5s/JFuFXAw5c3ftx5oRf3r+kCw9cTpMEhDdCr
MGGq+xxAgspVr4iZdXy9jm3knWYxF+2YmHd8TNSNczUuPYTSbwXce7ZQjPv6rSxnKUB8wedcsFRl
xFbojEo0VYP5PZnBFcTi7pqA8Xa0gZIQpM4yYVmu0UHQhQUdn+xso73fxnpYaMjDA57McwbDamML
MOjeQDaz5An7ZYWebp2prl6dJYz1idVKqqRqQZnm3O9la2dV4yGmopeL8vGTdEZZTwrvhbVPHKf0
J/64NBt1jjSXLqwPFGQFBGhiplsjUmBMpyplaoKpo3Ey58muOpp6YaqEV3wiAT/Zli6s6KWPATRV
t/8HfazrjGU4ivR491UWhr6oiYzeBzK0Dhknv48iO8DK3sByPyaEcWF8F7mBcmbnp3GYB780hUuz
V7nn4WTekT0jriQln8VQBdD7F5ufTvs/+mcIVwqk+NtIH1VKL+y3AtC10ekY1w0Fq51DIwIX4KGl
9vNoueXa8kPco6OmBqnqoi4OG8dak611dCtdWhOcXOmyz/lUiZr9eYcXhI6kGlJfQL1eJy3tYy/c
7Sg1K8ca9HyvBrpIbyV85Stvt+Xn32rdfcU0d4uudrH2BjHcN/IWBB5IVFWAYDIKujFGZMsAJpbZ
QWzk7iMk/DSfX9xfjxGgbr/IzDecVTxl+fqOtaKMpPhIjWk1Y1MmhGyYYH/GeVuYhD1EeiyTL8Ls
WHMmnbl6Vuq5Bc3AReEsUKdK8RGkZM2uk1Yg58lzw3dS9pnY6TZW/js1yY/y+rt5Xia/8YMyACNh
rgxcn+oi4KnP1cxkMn63/Dn3paBeg0v9sMihj67xydSdVV06Aeos4fZZ75ixxycR+ijXK4rFGKvm
kjcDQ2uDn+SPjlBx4l/2aclFAvqL1nRirzf3hw+w/WhaeklKNcESG6V0BU5sxsrpbM6g4qYjC6/7
Fi05D31dd2UWNKFZRZa8Dnpfw76ecNEnI4G+r/wcT7Uu8XU/QZG0R6X2vuue9C5KwHtrIyyI70bW
uB01YWNU17mmLJ46BpmO1KQYKpExIXid6TCGTXF8q1xcGOlGv5QQY+cC8nFKOrH0/0G+vltlxLKJ
mH0/Y0HyofZ2Wn70bMPiUFIOEsjij/Cw2Z/DgBc2fphUwqtvFrhtttDnCmsZlDBjBg97ICtgBHm9
K8zesyRmElartBCj7S+bDVOWw3+EOIq8XaSVr1qhBptA7WX7Tol5G60N2CMcbSWjxaOyKY1wLEuX
M043tgIzR9QU49X0VYweRn93kKbKbHPRWsDX1ambJhRYI6+2meg2wZt+fzPG2ghOZKwF+oauHQl2
0auKq0av2M7Jc5dcM2gkb2daX961YlC27T6k1lM+6g+RaRu1E2y1aSpUrU6p9Oaa2mrTpiS+KrnK
gdhSH6M0lNJTvo+qIbTGhVtEo4kj5X7R+fYYddwh1Y/PtjzET2X/I0BBtiFGVergfLEcxJQPrK1z
w/zkBMnQShFeYkb6IqVx29K+pk5qAwcfO2Uk8iHlTTY4bHqCGHMqAXKi1yFHHob852Qbhk7Tu3nG
3uFgPyGQLJY4E1iVc2mbIEfpvLqYvw7QPkv9DgN7ec4mnNYUMpEJVFgxhwXIjEN9A89tafAsxG71
hhGHSzwmyb4upGlzpaNAOdEtOxZEVcax+C4PysHCiyWc62aT6yzRlYtTo+nzyknrwF8djRS7xOhn
bUANZtfIokSF2OxfLlJhgpCvdTWTwU3j7ckLK0WVIqBxocf7yPKDH8iC4APvyZE3EeoG0rtl01JI
CjrfnXr4BIll581SUfXheH1SVxdH7wej01tCKqpL8MYZi9qInBYEfizjuwg+oU3k1dFIzYmf73jT
TmK0tDbHC1EbzM9DYCbFoDfVaoCW/U0+Mj4Bj/jxe9uBIkWWCESeNSt4S4u4B2o0zSzrxzDayIQB
tUtVbgq1zre7J0pz+3HX/pWR128zFbgSKz/csidQ+Zbor4jcMC7YW1FeQQYFz4e/yv9MpWqs7Hiw
C8pVBknLFBSL0zCxu+Kjrv0NqwyVfMbOa+ZCH5QtlWks47zluEnbP3SrVMtlLMHAmfQc4GtsJ9oh
CHb9kKXsCB8O8c1bO/EtJymVzZUQ8NyKwfDOASvb6V6YvJE+M6/4CXrNJBmLh7PsKAI3G4gDX1hg
obNkTFbOqjGd1yx29O9eAhDZbnEbv35sYgSMc0XnQHf17GPzubaXSvHOQ1G9UcslMDgd8aX+E141
VVNUYuyqCGceCE0Mt46huF2EEJnaRGmtu1CImSJUH2bQ5ZbbpYB6QB6ZC4V9c3cazUbA338hskjw
7LE7uxvwvzzUtBnRY0kNyq3lIdPBGM6q3FxWGWdMZ3TpEZs91zqQgkwQJ/Wa++XnkScUzFV5FrsT
AKmFfm7rDGq8WT72rrU7CUULO1pJteR9JzelLXUpoH21AOHue24lgQCh5Bj9nhSi9YHNWf7Q+Zyy
CUaXCf7ZEw1uhqQZ++KlV2N2UudXuiovGGYv31gff0hY2EZcwy3yFAxCSG7oyZUMAJofj0gYphQJ
35XRziICDcbJLE50RxFAcP9MaegfILyhqAg0vYpiNuH3/dNkcSk99a9ueP+qiROXRDwxH1aedfdJ
BtESfRTaV3YBumoyhScP4yZQ2BF5ccQkK+T5SSnQGXjtcZ/+rhrv7wF+mt+PjK/AnguID1pV/eLG
Vs6LF36ZHXAzHWOIj+Nuu/FeRDZfwqMYmO8EwJ8a+9DyB2EgMvfUyeYUy6g0e3ChkAw1p4Evbad4
kw73pdXD3YkceN109yaYVoeFqsEaIZgV+8Q/sZ76lxhGtX29qhqtibcxo/Er5AwUtShUgKJoVDLT
0Bd3eVaRdurBki1jpLAThlsX/Czej0x3ed7rbJ5C9p6SkJVzA+zKPrcUqZftUxO82hr3+DVQiB1x
uR5/Xqf98cJUJTnZCgnJc4CBWkN1tOhPKAhyOuse9f6F9PND9RuosSlYeWvU2Ixc+8+QAF0LmGFX
tgxZtGob8KzybLkJ6xeLaacyyJsOls4VTt6kZL/RS7hsna6g+/BoSUN7ctS/Ld2pWFy+jqN5W+Y5
ifF0IFmyoZSoCaHXA7m03FhFVAfyPvBG9EI/Cj6f81e2Bh5FJs1r6STAPffuEBWMYxDnamITX3sD
MGDIjKWxIlaPGVljFJtLF6HZ1upcKReLK8AMkTzDjx2otyI6SfuQpk1qq/JemFAdA1Ssl/7VJxcn
Z48/OKrsQQUd6LNRXF5fhke4r7wv52smdTQoJa4hDrjqFmuopzYI9wkzFaBi59qwzWcDpegVxrnk
GDpi9rdhlVdGM1Ki6e4oPiwzV/uR1J2A787KLH5z1xJL3jBMM7IumiDRg9i0Y/oGHaRxuP4c3Vck
430hvutbf0Xbqb3aeF6b7WNQ5eQdXv1DHDjqb/qjQEpl+E5Ong2W4CjcbcUs2TWHbmdv3SWwW07e
8Rx3a+9DBbOdPgsDxp6yql67lmAl5Se6p2axdp/oK6UdDMBujbMzwSaOTxvC3nvDmiZm2C3mYIy9
APVZKjVzM0RJTeh50fNEbDosGU+lWCZyKezc6g/O2aSAUwFChm9jkt0c3BNNEjF/XSvEa9ZWlmoL
NLPag/RqADn39KsNroKKxasEddGAf0R9rIA696veJqcYXyQku29h5a8QKhxx3qF2aIFBBQ2Fojiv
QZvVO9Ru96TpYQFC3b1uLqXgHLdP6N4s8S80YZj72f5jYhqz0U0fMibqElh8FAwESatVdFLE0W4c
U/4clAu526Inw0yF6XTK78g1OUPMA9KkOB6DYGwcbKpOqfWRx13A/lB4NBTSK+2GDPu1mLbnsHW7
iaDrMY6NC0LJOTXzS06zqUVK9D18A431ldySxvAW6v8ET7bCn9h9brVzxe4eUKekp5bVBlBG2qUr
i6NRWsMfHgbulO9ZuXHdd8SkDBdgf2yQXU8l+TgRxP3CvhG2WfmpmXuBtuDbzelVR5z32RUaQ2OD
XRBPm87v6ZXer8LDYB/V1CAsqgeO3Wfl36n/zk+8xkEnwoSxxmAgFiKSh6nrHYsYccvr6/wPXgqN
SHUdneOUaD+6H0At+hrNO3H7Jv0Kj6OjPTm3sf/qDBBsG4WzeaWRMqukZK2ZcBnkHcdwgRzXu9rh
r3Hd9L+XQ1JlZSEl82U8Pl8xI0wBhhSIlsjy/3zbE1T+ZmJFjGj+7xA5utzzQaKwkRgi3nr94eCF
620ShMM9loa20XD3wVvgquZiEh9CwI68UOSMva4hw9sC4gVOUBvpUK+lFDzPGavc+FVoRESlgPVE
RpFHHiiwismy+d8+zaKLsLL7Oqn2yxEmPBTSECaiS6aiBpTgoWVZdhTvPkVc8/C7JOCGCX23yLR9
cZQhbONiIpRAy/uCwi3nle/5Ygtg4kjyJoq7W24jG+J76D/P6rrSXD5TtJ2aaB9GO7Da6uLBma6n
ewJhcPzc/MbDe2fR3jKiREfTkdTCWV4ZQqwSBOT8e+qwTpCKD3ld1B8NbnGiXKmQbfEh9CoZrtM1
AD7TCiyxAzkzYXzbWaHQvY2H/le09rqN/5aaQcOteIv+Io0D+veygqLHkeyh6c6Bv8PMeRp4LSC6
Nc7fi7xWY+r1l+KpLF4WpIizmz79e3n4RULzcLFpnYvByrCXkIzD/DeFhkFodWGGF65TOPQkaSca
jUU/FPjeOuZZGqy1hsQC7ccyHwAiuZHlbuC+/KGDNsp5H6oWh97OVBMGJlXlltcNZbHo7WlyLjpo
2CII3EAZ0E942MJzfnwKVYR9lj+ajB2EUbBJuj7k9us2rVfjGcLiWoXm68rKf2UrkqmzaExQwwNk
54ZgKl/VJ3uauJ3imik1whE3NByJCvVhcwTUQjHg35crKV4kTAOWU57H2nj7Hgf/RQD3IomdHcHX
Omxg65JJkwOjsTsDxQ8bvpjjfEdayuUiU1t1Od0QXmPmytU2Y4OZqFHinvnOihGdyCmD04h12OxR
YAPmwZFph1SX/fTEKxJt/1R3vaOgnWES+747yQBIGMdBX69aZoR9N+66LW6qA5H+Zz6UIL72/3Y4
pZdA2AxEbb58JtCFsBz9ooONZG1pyC/ORn2gTDxRam7M47qrUgbdDN59HVR0jwdE8uiRhFTPzkHV
eMxalggGKJ//4Czm2nDy344YXFw6bJ3dUBjHvSQmlsl095ovQNK1AawuzRMAIwvv6svLizIwDJOF
5qYezdaSHsRh4KH8Pw1dl0OMvHlRuoDr6rZGOCqtBJ1yqMnM9JP7B898otQleHeARnoILYpJNhCT
6CgDzmZXA3kKICWZhnPert021bE7ZY3RZ/hozsvYO/eIY9UGUKq+omVXSCp4W+TPONzZIldru/74
dDdtxTVbgTX4cJns/BTJoD+BtyzFcvmoSWjsLfxtNgiSkGf81jkx9HDXjTrG1sb5woQ79mzGGqdj
vesWHYrKjUbNbbSPNRuVkfURHbmVgsSgoGfYMOLbBZk3j+C3u1U1dQ0f65DZlPo+tzgIXJPpY2QO
lVFO6A1cETB5bkQtSCeuExoGr5pnPjUH16RdQyN6mGMatyKNd5OHL+wE+DZGZpqQTlukaDcS/5by
jtWBHxkGFtPFsvWBMTAK8sv+DTH4AAKVW580LSVg+5BvXkE8EafTjh91rhVbH0eK51z2gUrdoI1G
3PKsttnqpOTj0S/mCVSWnqkn2bwaY53go2dMdGTc2VZ6e7HWr8/GpWZtD/CEzJwjC9cgEtazL0Eb
xh9Wm4IV4DaUcXFm0u1i3ha9A5tIvAofZRMgP0zkZ/DNanq89LbQViUy9j91hOCGLj8T+rXxkwBt
3tb0ldMI33POnkHPskj4QzhVch844p/AypK4oZEdRQLSeuGzSDxovmavHXBbDt2L6vi2LXiBbzyV
4U9q+jV/dhrH7oxiLGFsk39A57EoQ+95RWydWTFyUeNEYDadmtmiV97jEPsPft7QZHEgYBLODDK/
KW9ym0TehJG5k7Aa1ugeYBzgn3edLPXgcmtSRE/76TT0gVqOkecM4dFnt7egWQtTc0YxcTvR6z2R
wIShsstIVsUS3rIZYbBxLjJgLJm1kGzje+UGuKFtbZFpngVC7urOd8/NsApot/Tsc0DkYehJ+l6S
mauJGP9INyDaSn8gkMo65tu7WV/TdYgaCM9nv5dcAVIXe1kgftUWs7mvnOLSh+rJk1kJ+uEb3xU1
coXKftm5QqA9jUFq0rSmW/PhR67KeRRhMKxL7RkiHaa/m2WB2tbMGSD70InutFJLrTPjssabw6MR
7js65HODoAzIyEL9F3hlQjG4rsZfwARSvXUTzP61jfNn/LbNzRG2of4KfyZr0VjEJnf+eM7upfxB
SqiM4YGs4/q2VFRBgyRgor05wbhn4yu0FtCZ2MxdCgGP09jDwGrCGq6zsl17tTkSsxO9xThZCR1U
tAbP1BFqKhYvnu6AGqwOtQVT/GxidOtB6clmoUqAEenDEAnmyaojVAaHpO1/gmh1pws7s6GpJzaZ
QKVC+xBkb051/kHtW3vkPgX8m13SYEcxgSHw8NlSgAaVu1IAYm7LNyK6X4dKRoJqgvyfuu/bak41
VUVEvb0BGDrnqaDkAiqL8K+N4zvdGnQoxFIpz7nm7HBGihwVzixDJ7o3iU7BYKo3GtvujFhomyh3
XaPVj6UDMMSYr2yEzKmWwrhwM5sbhgX1BXDvnL5oY7KB6Lk35QOrW3Ul17nZQUbgDtBkBGv+Xx2i
VaOgjbi+TBcuy962R0vykf2MHgSTh66sXgL1FMZRgGVkiVPcfpxIqkco6J5ncQqlHaB2HLme5wdy
js6mEL1q0f4b0VV5vD1YSJJLQrvr5OpT92mYZ18gR8cSm/aU5yAsAaq/2WTBkXTJZK85ks7SaH5N
cvHHAJrOPPfLT2d8ZX/vUbYVmj+orVp8TRCPQTuZ43JVeTLQike49t3wZFWmhJlRoCJw4qOA++GB
8LKqsAXjqwxMdpqOPEkSvULubF07T6IZN4cjqqG4pC3g8c9OPF6KPtkmJj975Oi/xhHSRbT4GfVI
YsbNM7DpOaQdXooCxxUGVoqsmG+CTtQNaaBmWCo7JEKsWnLOVGw9T/y5xggIx9p+6eBgbGgehdYY
RePI6u/GhhISm8UbLRUgq6v6LSJicnFaq+9QQje2KpN2u+UFLkaDzM4H/mAiJ5w+nZKQF3Zc2ipr
vPqQWO7DXCT2KbMR5zC74LcPwT+PEHdivoTckw/uR/yZ0oM6lhZiH39gPgX3LPCYc7lXQlJxf3j0
JK/prbJNXfaLtJFGaHbX0CyBOpDeTgi30tEdMH98H+G+cmjXNu3OqqOglfdO9rhTO9tyJIQtVeK8
KtJqwyvFdOTZDHpK0wa/LS7ktYedWiLuUc6GRdm+tu211XOXWPK+Hsd1EJXHmlVZ6zSMRv0wjeMg
JDT2K662F8yc5wO4E54n/57aYpRiO+pjlf8xn4CfmeEjiZKij8gbhexPjcz9R7v7HVHg85ItJ60S
N427zDZ5REgnYmPC0LHi9drZGREhJo/kZW5RmTbmmqyzVNQLCnzC2So1XAtqlQkm7welEVMSoaAh
tR69NL9p0kFs2T7Z0odlvl1gXWCyngS1YPlmDsvlaZO2urvLSVuG4KOOMTCGPLMhonqSFQldyV7R
rw3PaBiiV50t44vS15KFv0Tgh5nqB9lsurI0xdn3IrukpSeTbSBIs6Dfjccc6bngAgsxp128mcxR
bV69PAPt1pb86OkPPv1wxgGTipZk1h2AWl3DkkbKi83Jd4JUh+Lva4T7Z7hgRzWgRvCb0FPB+GOd
J3HJavEWA29yaxF5DtmTPK3ObsaibU3QYJVJA+kPyyVfbcCHI3X8RKCFUdMzHeOKnOby4n11SP+x
h8rx1kfvKJVAFGls1OFWBeFZ9JQgYEbuduVzurudGY5BL31x+n45EhKIgZied3XhTO4uvZZcFqGM
5OgB9flVqB2S1RMBEEzg9Ur9vBAO5BD6Xy8W7NynhOJYB4DM189fzpanAIJR+I1S+Q0VaFvz9x4j
jYlnKVG4cuOqJ8GyLRaIyMqkFQiBMUewUIDrb3zbYL8g6edNF8aH+LIeHMzBw2jifEIiI+mgpEYf
IFj/911yN5U83gGzAkdXe37szNp5HM865TsxeaPflnnPNn2VMC7hLEe4Wp7bd7bDhSf+9SADjAtc
q7BVm7l6L/bgH37XDfhlJZOUkSkfOin0ZiaO/htXYu5M7j1y+lCktyJb1yzuRAC3CSfE/szblMpR
ZPQoacIeLRsabq2msYnJKPo5Q8NvXBnDOaXYp7r9AWxfSrAEY5ELaXqWY4N4r9Nieq3c6rsSqbpN
t/F2EyOHePw83pluEzzhTqEv0LFpBoxRv4myEqW30yFiUS9ebsxIwiACcm6mlFxVJc+w5dfJ64rN
b1yzTQR126tlKQsiWLbnPNv4ZXZUqY6ACFioapr6GK9jYMr99x6XAHzSkKXytLJQpNJ44McZkHXq
uE5AP2xQ6dqD06lSyatt5gZXqx1wqwehxeoeArrh2b98sQJFtrf85wNO7kGBSQps9c08laZATOo6
3XpYLzARg7c0OcuNy/KD54x4VOCyMf7Tw58FBbNF6cIUkIojhgI8vLs70zhjQF/lNHhEu7vYRs1i
AUoHEq5rx0EFuE63+hii1M+aosNgpy+EMMbehWN2UMeu9UqCvOeE+4weU3ysC5P4LcERTPDHxqkl
NHeHPJILLNtotGI6v2Cg9d4FJY5Jh0iUNWffGM/ISAIXjbSHTd4SxOOFVGFSPuNleqRgRwj8pXjR
soC+Zd3EwCeMKLUcHgtgr8yCbgaXcG/QKErKQOPXrFZKtbaKHu4ex/2bVy4b9vr/i2qb2gDDMXGj
laklF3SPjVRQ7aiOnArSS0fjHjZLd/n1U2/3yL58xfbU44jUIZbK5GSilhUbDAy1Gmb5gBtybla7
OI1nT1goA8qoAbhJxAderPJrqP5MAtCvKzI/qhhU5LuxWwIlhUdZXOI3Ts7ABQI0OVpBk/yqvDpq
dHS3IG4PHeTNpfEa9P0AZrHJBQmhBKKzEWEPMoq+WdTVSJxPFExExFrbu/OjPTWdn9pkvpl7TJwP
QWhB9C2D7pykju8lI1KSNIKK4UG0F0Mm1oMMRg6tKLmqXHL7cjAKvqqb2kbcBr37dSJ3ZItmtd5w
0Z8FARY1iwJzdsaVXy9mWDeFKe7142Hknleovmc2pjC+jqUcovFtxFrjUNz9hpNgTJUEP4EHsLBK
HQevUL8W1/GN9yayXNlt+zT0XwKMpFz7qp/yZJmU2etUhwvpIvVA3z+zMkh+M6jWElSCzjZZklHU
BhiPrt3S4reLlFiFS0C744rrBYyQNLkm83d+Y9th3Cb1MxK3GfAogrG4OoC0WJfN2X9o02mP+paD
RJF7xKuIt2VqO3nTO7V34BSXTOAejTu4MYxwx4ougJfluYWNSlnQzXDc8dV71EpwUH0K2k/R2Lma
KYcC7iM9eE+wO9rAGzxrJN6NiRUKSABIaHQ20k2mV/eMXHEwuJCw1V8b9XSjGpSZO/yUdxx9qILs
+Z0oxjLVJrSHYHjnePGWBiqX3ELiEprfk9YO0QldAq9GZv3xRtEdj2JOPvk/Zn9vY7XKbKOESOEL
zStid0rg+3pPdnRJCM78VuNIjnC3pcCJAtCVELYfGjzwgIMJGUROiFidXzgjkh/TD1rS/1z9nTLZ
bqwjjuyYUGYkli4GPqkmEe9h2MgNhwxPDzlUMsTqQBw5ozFjIH6ywgyX4xyyrccP1Y1E3LEIybNX
H8Aj9n7ohBB+FqKNEebtQ2WWmpfQwMRdqDlrzR01sYGPmbheHX8J6VU86Ok1TxtlFiL0Rqn12CaX
z+jgul34RyDx6AfpdZA1l01ILXOrKlmqQ4q5aS4oX/UaPFJFVaU3iuxmfDZ58IZwKSelrOQ5z5pi
uMKLbvyiVlO31y7lG77M/1g6yGEMQWvbjvKnLblS+KBuOwwrbCc4XFFY9OY4Y6B3tQAPh1v2R4a7
jHwwXDxbDbAqp9FmNrNQhnY6oemz2DaWX2Xy0Gs0+TDnMB7HlQUz71XmDM+mzXZqEpZnLeGtN2ek
uB4TzC6PwvzvHpD5DLdTkFNAfTPK/PITfYD1wSAFs4ay1fXMiPqmfN+0HPgDtoWJuYPjqRU6zlGN
L1R9Ax1lDkgRLPX8KXfVNF+WcfCvF49DcyDIXRfMpJLUPTUqp023bXkXfECoAf080y16DXPhRYqs
jF0f1jPmmI5n9T3I/Tw1sE0w142pgnzLO1A00oFrWlxtO11NabkSLHpveE8yS8EGiKOxnuMcEQoD
VMojghoSkDJzfuo1z5brjL8y42ZTDF92u1aC5oQXLnoO1J7BvLcDZcSwwtgLkcXfVsx1D7FgbSGH
29xtJI8E9oeNGfO+xA0URgk/sYDuYz3Pt75flXVqFNU7U0Adfre1XYFpywIHy0ZH6M3bFYwHEWZq
sPLIf9WxbsTARUiVwKcYhRQNhDwX6+m+vKlXVv7O/pvTfMsHrXsDvPSorOXpvronTkH4ZZXxQ3Ev
SfMOymaaHFHORSzSunCktY/pzlbq5VPV7S1dKJ3+PlagnmGqBTV1WU3yroDUnbk3SYkT3gvtWKD1
rG+b/tLfS0k4x7zo5pQ2xptDLmJCDpMo43PLwlmabXklExx2Hte2cwXhtahJiyUexME70OieQg6S
rtvb51xNhUWuNLqsGoE6no+KXx/hCUfylKkKiQD/o+jxPPOYEPm/cfXhKnxJb0nm37zu5PjlRGwx
lcitmhKKweZ1gfDmKVYiLgbm9169wpBHuWqMcBunWDH9TbfJXTy8E1t8pESAALL1kqdgpcCea9VL
OG9x1ms8JS0SWuqwePFs8qdAHVoH94mfSjGbOsoT4RkINLPhmr2PmzSuzN/exEUjiIRGo1Ejr7an
c9joObrW/AQUowMt73+7SZGtqTqUuOne3zw8pzB/cKGZUHqSNDU6HqFezD38nKBcO83gpjtRjQOG
fe/sIE9WKOLpS6qNcLVkBgRn3j8u/wCi2xjzYiSGAPUU7/MOjp/B3baIBa8GFf9I+lk66+9l33wI
2gAPADkpzIO03BUcXqVSN+lg8Yd8YAAEDOFNzHIAFpC903ow9XEjy07VGBvo4wG2DkcN07JLUQnQ
nugrWsrTzPMe2Ze33w/hodG4ZhHvjgfHoxxUQH3FyCLv3K1YveJHjAPvykWPsXTrXiZksJ7YUFd6
1QiS0kvWpmvYMI3i3ITUu8sODizvd+0wjed7Kv93uUXasZgAN13jBhxZ9gGkKJstiqzrq6P/QygP
917sRklkNmetTEl7RsbQPa7tfWURaL7O9gJYyEWG/DfWtuMdQXFr7Gr27ffCHOQVrzUqwU/5vO82
0sAFyW8vYZTeK0cEpOB7ethdtZr+KK1H95cOj4Dg4ziPEB8kst5WUqSyH00U76MV+a5UQqH8F64i
m6asXPFkw/bSHUtUBfQVfkGUo+zRGCAdqn+sET6Ik7815yfQry6eDFV51dYNIN4O90p1g+3NJBuF
luPPu2Vrd0mkcExvdugLcfV9SVl4KnVEyvsHyfuZ77GphD5zkWAmnnsY/ctvAs7UMWaREJzOkjcu
yEQH0o8ufWY8TL7IowPS5YZosDDLDYrQOQ/Nmd0qsm7uf2uxJOZS7pquhL2HV13fGnQLGvpBYIyf
srARhVJ8gudgh7RPZYkRRNv6m4xAEDDR1Nlv9TB4kEy+1MDYtJ2g7dLNV8W0Tu+LrILNEE7lXSwa
wAbOm+IXmdYFsnXbVaJGEIO7U2d2pu39408l8wTDDfwJ3h7/5dPWSX1mvxvHgFX5Uc30pzVP13/N
BhtEANa5Wyj/0D+3ci2h8aodS8NqASa7PkrDY6GdupTCBDA9CtrQ4AU6Cj2M2N4IeHr6keaS/laJ
ciN/tv/WboH/4XfgaxyWttpuZDpkibVaptbsv2DFXG/jG6mJ0xE0N6VqUZuFO67a5tT+PDumEMBc
t/ykxyeg7vSHxG0xqmj22J5SJR9DbufkjpFhnDHYBUb99ldgWMX/dFUnDRGTeMQ2cYcL3aq1LRY5
395aaaihSEzfg9xalPDuXXCQBnvgvB853kl/b2hHpVADrbP9VYtH63TusHIEiWiQLPc1T8d9o/DZ
8b7xaj7LPaWFrbeEgJRbjuQNUo3DWIlVb4jKI3OmLYG3toSvZjWnW3C/xWWtNEm2HtonAhJJGHXX
eKdQL5P4ttNIff+oHn0gwaRQyAmfT1IY/EM7+dMT2qTy8GU9FWs3fMbKAcr6Ww7bA7PzzA6NYzgI
QFQ3N31kRjhmoMqj8ufXh5Mj86hBH8Ich56SYYlgFYTFLxerQdNyUPd+EqLvQAGXUPr26vPBZ2Nj
JGoh91gFqZvB2dqnW5WPO3gP0a2f4uB7JbyTMRW9PHBa2fVWc8BvCXLtHupFoP8d+AZ09JsfLZEx
R9H6e9PW7uVy3mX07yVb5nt0ByHsLCau4AVSXGRdUBiEViZ7wA8SYLYFPJ0K5Lyn1+6DPmXcx1MP
Eebh5iSJRCt00hHPSCF4XzvbgU83ONQUdGrzHMOM7ikEow39r7lzLop/KowlehMKVnWDU5bnuN9q
WerrwveShFtG9cesTKfj6EAaIqjQpdhwJp04OgQSymL4mq3/MdmYEra4iphe1Clp6UQDd6az5NA5
sUAKIVOl5nuSh1Ax5VnxVc8XJBJ4kI8NnivvFLuM9UuqLTSLZU2uvfCs9dHSG8dBomNuz4ONvM1e
tVR1d1EANMkgdan0G8nbZAdSEbSHmuklB+E4JUheGywteyRzLqupzeb3yT1TjVDH541Rl2X579XF
NREgtvB469pvTG2xlyyE5cVN2eyGKWLtrrkChj85OOLNQXvmJXpSCHPTVNu77fZoQtTUdo6S4b9g
hKVg+Yg4VT/w+W0e4ZRJzP1qF2I6jtCBEBYOz44Mokh5JEyAbMfh9Whmxy0DVlX0WUVL5CJH53Ch
K8kmI6ou/w+rhYYsCzVIiUq6Sh6ijb+D3ELZKiWdCLJDNK90ylNosRJ9g1lQmsCXO+yuHZ7eGS8x
443xlgkY+sSrwHQJjFuS/Hpx0b1/hevZN6sD9DrqN9vltwfyCuWTjhWV2hPEKDMW+unVDxKFXqqT
1xfXIly+mFcybMAQw9J77G/92zV2X/UEtTrAYVnLOQRUf5daHx+7TI6f2xOJUDNWfC0bGAouAOd1
tz+fKhrfQRPPKulWErKMSQ9BXlldZF7GOTlGyozU5eiFb97Yt3eb7RGcqMlYLpTwOXXjgklU4ukO
hzkHl3kVSauRrhE1BFpaSN+D0jdUkerG++6ZBIvJBVnEIB5eGn5i7CuPQs1e/66DvUcG8VVZSi68
jSNyRBjhyi3rI5HDWzLR5htJ3REsVWXB71ItdYMmnxNSGYZg48o9SiAAUX4ViZTf3baUjPLiBtBf
WH8zsaB7TQj5HmtgMkimFSSHdxXsV6ukFiy34Gsm2yEaaG5uThA+jbhkDJtOjaScS4RKw0zuoQiT
doISVVBlhbf87pNoZ7L0NPoBxioAo2Jyr6jmAJ1JabFPFG/Uysz5fPS5EwabHj1e39Btt+jn+KOU
vorHmLbkzIpVLKCk3dBifnQ+9fhOtevekfrbkvA35h3K3Rbc59y55SoakDqTVETJH81NKa4ISVv6
VPz31iRs3/cbuuW4wKkfVSPToIyD93DMWCC/7TF27H21W1Usaa6tvqkFKd8gTiKR4m+JWQTttHxb
LC9DhFO8DDJZ1jigYIiOjsCxJQvRMh+tdYyXFPJwnsYFP+O9RKRTCqU/pu2SQ+rpyze242IlQZoI
QIANhj/oN8SrwkAZ/lbi7KfdoDQ0LzwW3lec3j7PzlbkUbDDFO/u2zA+pEtTnetr6dj9aPY0TPNP
WwaUDXJLIVvTVRTeAU+OkaivSkNhA0SD/A12rs4Zbk9ANlzFWkTcsNhV5WGY3FqtryGkav1tgF/Q
c7m4f2jgrndqYMvBz4JxSfm7fk4lzX5fNz2w4xXnvfRzsen07fJGsJ72tZI7ISY7qGmAe3oEqP/G
6WVJSbhf2a1aTgWvX5QdAzJRHwTkHdvRlC8vU2nV0MWHKr2y841CMNkagwwciwzqa7k+dDu9L6oD
/osQiZA7RB+OXuhA0nzkO6FMDWIbEU27Wr5YABfJF+AjYjg/kCgNW4wU5muilfolYEop3yHwWdwV
8C89SfZB1SzBElWEHvjzcQhpuzCLzY/bCvZPLXiQ55sppq0/dNwxxjG5x7ZefrwbxIjl/yaNDv7M
TJSVlgZQ9RzEXgdo6GWHO5tCfQFAmRr9xPwXugbVb0EfwY/KNVRmBjrnTpt5/76grNNh3a3XYTo7
ZlSArg9JbGwwv+Jc/j7WghZu9bug/60La3V330yf+bxgAmanWO1Dld3ijybv5QQ3x9Nbd0qyj77n
HQGmkenP7d0YMTpXPmUrXed9kEgo9GVE5h2oJtFAa5NyKy+tDT6V0xxUq88QLeTviHMGwj3Ua7gN
Hc0u3TLxPcAV/MQ0qI3J2Ee5+Tv4RJyws8kzPxH7S2qY46XEAjno4WwcE0xY6SE3h4/AAyR5jC90
hDu9Ks9yzLWF+hdHnhVYOmW8hnsr9a23tqUtoZ4B3zwV4AIG40+zaDyYA7nR9mwE8kHwy5Pf8yXA
DGOEjv4eCFzOqWxb1kM1UGbZO8c0oD+ewoabgsmKuk6HqwIWxmMX5zPWKXKa0G8lX348pqOcSGwQ
AnmuI/72Pqpg75sNseUbBZzCOsUp0oSs2hCbwqdN3KTa7322F9VUnDiOgtk9PVv6YGu183teWaCy
yGB8NkPEna/I8qepwFvbaIM77uPo6IrfLy4/rlqZQXleL18sNetgJQ0Mohl/hDwPSUW3mElhHIra
EcT3DT95GwPDrpyK0ntd9oiMtz+OjUzgfm4UTxaVMO80TmoaRu8jMDbeupnf5KvGJLmabBMb5BjR
ZM1OWY3GMS0BWr3uvDdYquCjleLB+/IpIgAGUYc7G0BKlu2sFnnDMi3YN8xXb1pr0UX5L8pT3ibc
RR1sNwSft8+t+6TdnRGZlkNHynXuoEWPz2TZCgb1WgG9Tddjrtl8ZCPl/Ojdc1jinAkvGgrvxoQv
5KaBPcRIoj31E//ZnOscPknjkaaxxQxBRVj9W2lZlubgOr5aB9T3dFI6shIAyZm4jQvtwHp0JZeA
fGAS60GoVo35sZmz5NJFK6H7E3+ry5RD8STCWXe3jVoq4QTLAmrcwDdPd86V84qAjKuCYoiRozx5
a7uCH/uOVfLJfaBWprIfOiS3Bums2Qz+VtgotRqlo+yV5sZULdjaqrlybwJzjUn/5T63QKgvDRfc
0Xa5I9tgV42ZQ2AP2M7G8bZmFH+riyMXNKhRVjia0wtBSFNujEeM1vG4U96fXGy53MXI6WwGwgpK
Bg4eytUv3zhdRGPze7tG76ykR/X2P4JoSz/f3hShwy4CINkAM5WED8hgkTT3d7qOLDZ3R+YAjg9i
+/T545lpvU+9vPJgjGnniit1ZmMg98N40WnAR0xT7ZJlOBu1XJtOsttBKYzfAV0yKywdUi9bM9un
w4ACbcpxlH+WBMYZW9WvuyqSa+0EVDFE0lCEB3rUKV1sJuUQ/5yTkeRLenT1QB12Cw5JAIANnnHv
Bk7CptwC3/pxi0BfdWFQ5rkEHjHI1EgsoNlW0dC1xOpfseINJTF+CfkOVxcVDk4nqR1W0HKuQ4GB
afOBvklZEmFBY8CQcF2bP41w5dRIR8qh9M86JC7SIYxgWb2SEuHbwdIC5wCX5ZpWJvnIn94lzsdd
G38cwwiyIYJrW09fLojGA76dRD1MfJJZ2MAagsBeh2vnkg77a34NdPcvdGn4HZ4L/6KWvRlBbw2v
A5s7O15uNNbsgPimnBYTSwk2nrwU1kWvXciZvu9U33vS6QVpXxIOUEtSdYR6zAjwXQR+N1e1tJQX
2jnvnA/DybG7p2Mmst/2Pgu+QfnV2jBv1F3XPA3UajdaWI1xcxDG8qWB7sW7V3O384e/gU5gU0n+
ztVU3ggP7G+zwwYOMN0uIZdNkmiEN+rBc5AbMYC0CT8j3TcXKXDEBqqaGWoexW3hdzeTRJ1FNPw4
BRH0UdYqayeFhdyfm004eiFwx4fctK7n7yqOkzDZtArIAOfOKgBnR4TCkPNFv28QbIsQrDxOJitW
CupK0t2uB8Fjc2A3fiHPT8ZMgcDFo3cMQ9KDT7D2DmyqfR6gT8YRP69cmerQwAdaBp8mu3MtHCto
hmZW+9+eTqCDIlAAR/QUwU51R3QkVWROFb9dJm1mSbEQb+Zx+5VlYufRL1Z1VKX84TaEp0pV/UFn
KlM3TmZ6l+uYgv3VEbDc7MD7BeHVso6j7TMOz+SLRhYQGIYEeNHjzOLtUdL14gklh/NiBGkNnHah
oNSF9NrJGGZTYtod1vcyEVoiybtJR4oaaq5zreFBU/arJJYUDsUqzrZC0jVG3/KemOZ3rr88sFSi
xMB/EuWymqqNgrLYfgiv7iQ3kwvYPTjdLX9uXmuFnKDiwliOYMxEgG0onBQAMFVVD3+EXNQCO7kE
EtnbkmDLiASez0O8G1Y0ySSYm7L3mdvAzv6lhevQ7AXRiCn50St9WNOBW7ZS4U0ygQNlgnw1qjj/
qUxjj+Vf3f8Hb6g3zli/qRtj6enFfKNTPHB0bj8p4gWic+LxusnvBXZpegnih0VZXujCpb3j1XOZ
wWFIjTIVL7XCsS46Gy2UlxEPcJgDZZJ9g21p9V4v0895l+8J++wMxL1yoKZx+ZC51dVBXDCUEMB6
OUVA+xm7qn4DfmRazDTr37DqxxyftpYy1kZ3EMTpMGMK8lRyyoLLBoJ2i0xZSrfbUDO9m5ONjMbW
KOlPhm9ttEW9aHQ6+qin09ojtlCtmrwQKo5NqzjV64sC0qVPHzJfs/oirMYaDbLt1CEDRUJJFxoL
j5At5hFqJsfx5VA72/DrIbmVRnZoRvh+MIBwVd6PCLW38Mvu+/l1gI0LmlnZVUA07sjA07T5PYW/
lh6kxygXWcB7N1kr/WE83fGkQAnGBcp2AEmMgKdQLmccACjC/QpueXdmxATbykktZ01PdKe/DGke
V4SyVzgqo+M4jOUlgxk5q2mdMuCwo0a3VA8d0PhpzDz3plhFqTm4UA+tiAsAhUzFyUrN6dMYf4Dy
F8xlB+b9E80p7+RDgoZqtt/rk8m1p+thtSOX8flkRy4K0s2xF0nkvtcgbkcTllxZkDKNIP0IBNmn
MPZODF5WFNIOCNIbZ5SyehIxwfO6okHvMQw/rxAcDfdWWn1g1oUhkjEfizkmruGozAZ/0G3TMmFD
8/+oHDisZiE7Eoc/22zr9f72PxtPVu8Xnd3MNmvDg/BR0Qp5/64PksOsl6o1IcL46fUTFoXnV4DW
TVD3ucxwr9t4zlEjDn7hM2SIBTq2qwWyfUKyqUAPesUsp0U9icB8C4GXwI+8Qn7OkdQ8yHRIoLLP
FHyZhHe4UWCOnEda+iYUR8QR5BIIIFYZuIxgxTC6BUThUDKGuIfd5tHrJoR/xVNM6ni4CZ1wDxAb
X+46omL9PbxLTF41IVxMONodImVP/awvDSccrWtvoRYRtJt8uMD5PPCkiluZJ/q7hC1YG3/Vebjn
Pr+fgXHYS0XgG99IsAvrrwVgW24coteWZeeyzCDniXDMBbPY20TbH95uV3GG4xq1gBfI40fn2Wdc
SG2pW4STbIkYTMNQID5J8yFKlSceKLd/CNQl1L9EHUDS5MMcn3n2N7vSs39Mhx+s+yupyd/4mLB0
dWop4daPLTz3xOj4FYu7B3Oe9leqdcdxaQGb839KSJSojsk0acBQqHgdmYhIEKnnLotnBqFQTY3i
4burDF9fy3c+F4fbSC94FA95+lfjiMTTa0g6W/6JRpjqpgTnB2+xkIJ5RHnVGUtNfpnJxRb1lGVX
Z5r4C4a1pSxxYrpKhIGx4f6sVVIzhsArUahmpdscqyonhETkyN3M0zEgUlilMoF22LaEkh5kcKhD
vGeaReWt3o6Be/YiKqxAmqdM0nuxDUJaKGU2CLD2HyZ013VRYTwHCimOJcR8CK0m9AlDy0fT9h/0
LK6dbAunsRPFcQAg/tUTaQfDaFi2uZPQbNcL6goRTDUSc6qNBQ7CzcmJtCGxbIvNh4OvZZZ08uqi
8spDl16SBFu6LcXk6hJV9IYWu6gNn+lSd2ihSnJJGcf8TO2aBPChO1OwHRVbeq6vvuU5xzXEn4Tl
L6hhsLADSYNjcOkapP3/lmwYxR2Fq8oPPoikZsJzRWzA8KpTcDxUT10gV0fUvpZONSviCf87LWq3
bhpNa3WphZ0lnA5qUEUwJ5MBIFKXfQbrea9JtZJnCQlhZF1W6GtytxzTbFkWVji2RwpbwrXoxk3f
mXaouWwKd5H/wthQOdIjkMGVKOJwoqj7zohpUuNIhqYWsHaAiLnJwLhuT5vEk5L0QmXAF7G09KwA
uXb+JsRwnPd5jauQLHwNsC0JUe28z4dgcQGZIpnoNxPqpxL/NeSHtyOw0VeaB09F5iB5G9lSBzma
xHrcObQ4zeiJaCcQ52GFNVQJQ3eKIVAi6ivM1vP3wkQE0WIVWHBsZO4sgJDYsib0P6N8doGey/KG
ECCo3e7yq8RJD2Zt2Jq2XxxU66SOdVyH6T3aAMTdQqgyOsJCN0hanHpfwzlJe4n9ekaTBb8erJEY
UGjBgaAi59Zm4S2SvqTJVK8CJLdxzcGD9luv/HLDQ2nOrEvDUWEIVrg60o/8xsjz/qBvyg/kGYsq
/YR8snmmj8fTOaAJ7TzGuyg7xmkm3MPM638493lwwhWDe7m6USBgZRUDAfEcvOF1+G43PUwf3m3O
YztcZ6w80ZkwQfUCfJT5gbcecyY/Pv0nYkkIHjxANs76i8kM49GgcQO4iI5VHH2neqKg+8IhYy/A
tmlqTux2UcT4sKlLDryETw1lDjH5GV3fqTDbtvioCGMUhZ7QrTSE8RvaXoO7bqzswG5Wnf7zYGGd
aiPtclM1AFRQcOxIrPJlbwOhv+HQPCc2EixUkyH3QUKVeVRHGlXvDElh7Bscx/P1hR9EF8tZvdJj
QaPcbYQD4eZhvr00be20Y/gKZElNKLsjOfVd+BHkxm5eakNSry2FBZCGcOobdqaQwqiY5gYDFXy2
hjWJhf6OQvzeB3pQPQv/smjCQG65FKHAPmavSSWBeK4Nr1HrMv7WkhAhmj82KXctuy7Sygs7Uzlo
Mcjgyujkr7RP4eFAwpc451hhjW+rmPF9QE1uitUh0tXIl4nzxnXuoqDHCLE4RgwueEyl/p+eMXNx
1bkYLI4lRoh6URGS7rSLh/vPggDUgoBtFQ/GaylrWGzbdvNYjDk3uBYgFwSx40oqoaFtC2/mRzdb
r1ADfXbVUiOyhrwZAhuQPyJpZP4eTQexd8eaIUsFpQ6PZJQY0OUlk8lXe2v0crB6mzEH7I1cHbt8
/wq9AnjtBDQMSrqMfeDFBe0q1q/2N82CYrwrO/elkyAT5V+0qm7kiNqdT4CuMHhUreQs9wEmS2eX
zqHX3i8LDekv/xyVTjVHXIieNhHV5KYsY6HSj3ZYKSP3N5HmtAPkQ3T3CTzqy3MNZGn9I6kpcc1O
eXP/KeXDBZnf0Q9Y2dpLEGP68BYnLPffZRGkxTAD0gLZYVZELOlxuU6MJtoUU1lMNt+JfXUgZuku
AmWrGsTfNjPrM8IbK/7TOZlCWr17y2yZ1QQmzyzZSWtYzreBSCdSYANRtjIl67KX+73T21yrL8uD
eDnyLoXmTqv/zNJELU/Wdz9zc3e3Yj7heYPeCpUEVyPqje+VVOFkGovAAkXtNySPZPADZlEgdDUo
j62X8Ofkn0yl7C4lMDPrLX88SGMc+WVDmFp+IVH8uHjoqocRMrS6TFCjcBWjVWU9sj0cuzMZ6BuN
AEVelY5gFQBP0U3mb6dBI7joqiYucolH6n6doOKEgOLGRWJjPieOK0lZTBlmiwLaENmNH6IqRw8b
2P7VSsH3doyG1mCKj1LlbxZPShIc6R3TPWqXcMhNTtoCELxLQkwGlUUM2DsFuZk0U9GMtlrBmJ6X
Qh/QJNMcbUbe9sNgMPKkjk8Tu9JLXHYQq+TFejhUAT41UVjSIZ+hEYAesCbJvYdPSDGWQKJ/TpaC
xySTecmGrfC8HZcLde+UO8niSx272ug18LUMfL2eI7/pW6cU1cHjhZSTf58Ewsm4tLEYlZ1qmrL/
Svkv06nRedmQfMQhp2wacRfgbUYrfPWXMgGbclcRBhHLvxxHu9HcLgjNJBKmwLAFzmudwyB7pir5
YOF5Y0iuFABPsjUA4/mTTUAw70byojuZSUWfGQC/Faw8A4lKS96vVPFASU2DijSpP+BhqMhtx6/j
KAJ4JuoZy2muZMRuvjc4dx/j6f/cHZIk417GFcLS/1bQPxbvaxC7AjTLSsFYUzMP1fAFihZaPzaA
V4R/2EC7yuywoWvJdyJaiDBMgY5ZefCtetuBWkHqR24QD81YKfVYrLffhBCGFomgR5Feqq0+CupJ
DTtdB4yVawVI8d1noZXoLuPHripPVETzYo+LeKbx3N4P+td9FbtL5cCWQFOIHFA3PD/4x0LRHygK
Y9ByFuAlBEp8+RU8TdgNbP9JsCrZ0X3mwgADxDMchBI5OjypN6s5DdbbewMHjZUpISPFXVCfeMut
ByftOD+phFhhrXoGIFReqA5JB1StlWP3SuF0aE7y4UuBGDmHk8uM07DKNpiyRmxqFPPAzUHt4r2Q
+ddRkay0l7CTl900cphZjUSP2G4svGahpe+oQi7S4yB7eXdxRAFHsqWdnAl8+ShkZQQsdGhx2hrI
iJ0WUk44/B0tHoOFtIuzNsIOj+98iMK0Ajj2LlVmlkzNTkNSo/M8at6AYRIUA8mySORwYKJaiGEr
njX7XL2ERNpdE5onz++/gbC6nwx+pcFTHu3TDPBAdusSlEQl9FwlFIuY4Dw9QmeYNaZArvncd7eC
FHVI6frxVeuVW7HN/YUTZoLRVk0HtgaCgyh60o0Duicbc9rIQl1HTu2bQIuTC9AmRUThXXuPcyV2
XyZ6lDFhrhx9WF/554vMNkxAbw5Si0Bb+n2NYdzQ4pn9ZW/P0ompiV+wcGQGlvvrZT9hE6Otzpd5
/NDlBR4JaZADU071sDECPNPpuLyh7N04aiDPBHqr+59MhOYPit/onHS23xphW4dp/8OUBknrYO9v
wMUxGmGy0eFauF0wtFNMgjsYNagDL2lV9OARQHJpHpuOqXV/99nZPU9hSOSEpgx+SpF4loO+gjem
YdpQnZd+ievnZHGD+qqMCDaLaghLOMYV87epZESZfNdxOOGvmdHOUDz7T1bjWiOk+dLoz7hx2mUj
+tcJ0ri/69PkepvLDuYo+bvFGM+UE7vsYkaePQ2B66hk6WJK0Wtyo8rTppOoeiDgHSfOZYLlCsmq
4UfyCy2LNhWyDIT8B/KnDcxmGgpxqZdAy9oPLHlu99aTNs1jFBupZPPr4lR1umn7p2kKzBaNeHXN
paOrn0TY6fv4wUCex72Gb8I3PZJYFn/oxppJvmbuz84c2mtbKnFSwN6Dy9mAAA2RQlXk6Et67m+Y
dMljzCMA7P3J6t4xTEFGWpCX26UPH2/jOIxSzndSD0jGrYS1V67Foh9oIgmwB4QDzozA7oFW28hn
0NMzbJjp9jGmL2u1Ix2qPeVEu+IE4SB97GjcCcO/Bu3+nIwsoC7VRdVDYmDIKFLwf2DvitU7lmv+
kBhs1ATeB+Tf4jRd6ReW73929nO5eU79G9ypD4V4+nXLl3PfJWSJi4dQ120u96sbIS3cBWiJovdq
abc1Z3jSrObd5EiB6GHuKS9lhUXvfpFRAfJ7yHZtOnzwM/lkjkMtF7/ZzILO0fXkkPSXUtUpMvde
utPAmZoq9YkcY3YFBPpfbOGmp/89rzrnaeRFEbzKW5sexoO7ycFbRJpHCTEwn+rxMsn8uQzGjP+J
i/Gt+ucL44+3NQToNaVG6Px/hhqmInSFYLiSloI3TfT5x3lhPO0naEePi0QkbCEuo0Husa9XVwmZ
BSf+RQagKeyM2SVAXKK4SZitdlZnSqM8bJwk9TG/dE639kYUkhp8aS/qIXC8iLzCY8bbDo/BrSCO
Uh3toxn/MlmGOV5pmP8U4d9g4jRF3ClkzI/hiH7OZ9MbbMPKRsAJaQfNTWc28zgM+l3IWprkbB94
VAz8ynbj9iJYJwEF31h0IpsSvhzJX6hT81eT+fYItHUNOXJ20DTI/OqMkzBUYUIJkAoOTXMwJSTz
M7R1svdLeJu/JWxg5VEjgfL7/jeo5I3JENuHah8LzM74tEKeT5z4wM5IBVXzd7ISaUd/FQ2NpT3K
2z7SWP7UcnBUWMj/V1pfMLqdaoTzT39CfqJps+sRwofloZawUBm26lNpB6qChSp1XQPusrFBeZMo
mpMPdZESfAMz6P4+SlS24377E7bYXTXunze/Pssdvtf9un3pI8d6CjMK+JxQFl7CHDL92P0NfGP+
XJQ3uwFpuUcAXYERdA8XOqieALzlzqd8rLJXKqiqpT7wIbBiXPJWUiLZS1FqXBcAT8Dk8SyVTdpb
6Zh2pjDIx7lEtdvzMCy/X7+9NeEvAfHCryrktxPO6GDVQoo3bYEQrKiB1BpCfZO2q58MjCbI3gbq
W4zeNBa/5QQamiHcJOaOCMM6lUvChyMZqt4+oNZhAZYNi3IadgHo+soPOK/Ri/ytccexKytQ5J8V
+KSIFnyCmu5b6WugDJjV/Vp/5ChJQCT1pWBVDdfguY8yb8peyxp8+BdcTyaQRfVZhhCJvLDULn1h
QiA2Q3IKaPBFhGRWCoLARFFqq2WWz4+nY/Q5u+wSYbt6f1t4gvdagk2HG2aZqODJtjvJt2pwAvIx
0n0KSGENlSjbeBmj4BynypP1FJyKboqnyQSCAStr2XC1u4yvFB/d/JHsIcomQe3UVV/fxPXNp08B
wMcZAjhquejP0wDyeMlj98Gzzh7fgalqwxNm7LaTBKnHPxtDIPzUmTgeIhVqZXEeTUdiXqpjvTDm
EvYEl7QDTGiei44srwTfnHSYIRTADq3WU4fdUpb18sxzqUJVOjtf7SyaXbzeV9y+WfF0gCfw5vyJ
I7B9AusUfnNpIvqI36FQmw1BCVDH+iFajhXrDWeGOiMToeD0g2JBPMuFQaDanpmzw9nj/y5dpRJs
J395z1v7xiU/3wH3BAr2vjbIyAO4sHBXNd3p4sAZsQRT0cyrgBUdXs+nvyCdVJhcCZxWZ4pmnnyr
Vqy9TIgRpJGUEo2EdzF4GjtvwA/vAv1MigaP5ubN/nWtRLlPDHFGiW7rHXIHk/eQBBwsXfDzcYKl
g2lIKqvSLewdoPUuzkhSsMWLS4sjC18sm5kKxQutDYYIQdQ8QuK4/yjj0g0+BmLLQMM7hYRKsYpJ
xiSF11mvY0ukqmIN0pQ5lImitz0Z8qDajykIwQdIlkjlg1TcUVHCZGK6T6Vtt4BfOHgMuQKRkT2W
90wNlzF0J2pp3WTsXGhsSfqTGNVylxoDtfzpTivNmdkeNfpAoPJSvz019lRQyn6X5zvuVUk9Uxpr
+6KhRLCP0xtpSERuxAXT+WMmhJN0qmaa4AIHkKTdhPNbmHuk3eXsuafeAw9nI5GRpfc2MKMKMrOd
xJfH6ss4EiLPV9YgM6qTym5IxwppLIV2RsQ3YWT1vtn+8/U/GwPKm18NYhJqFrTvJjqrMY7e+Yc2
546W9tRDvRLmghQjyFVoDXHPc0x5H67e6WvyahhBuHHwWx7aIrrLvNo7SalRFgfkCdzG+jgPJotk
gS+FTN2n3wT4mvDMw5fMKbLbxP9AmE05OIq+kQZ7+eclFAAxDFI6/mo+749y/Dt7G5EZLkGrdyl9
OrT9XaYY6V95pmnhQrouQ2FZuOmKrJcC/1eZsRJkmKveLxNNlKyPL1/pN6VbogzaVArURVc8MMkb
jQGVV6i1VcRZXsT0Sunn/wrEXu5zJ86zySHLD9ObEJ/1bp0qVuih+zQDxaju/soSQdmCJu8qd8a8
ceXC0zk20JWjeMaJ9tjewKgP0yZ25dVqIbG2rKyWZsE8VTqX8RSejd+YPYI6CbMmfXjw9vdjtKfp
UqxNai5BVPNeGYKHVaB+kd4wOiSpOi/6Kbb/RkzXwPmhtagcvgeXdIvQjtPZDJmy6xJIitG5/KJI
yLBJ4eF36h3Steq/l9j7Q8zKqpvQxwirCxLxQlyEo7VcMr/1WEQxq0tgvjEc1QwlgL0PHWfuY1Ul
FhpWBQF04HV9DAzmKtnq/XemMbKHxtVf4pLReBn9dfGykjJ5Lr1+MD9rbI4FRgdSRDdIOdn1x+/1
CWo0rBNlMFgtCWElrOompiMz5kkLIyc1YkZ9w2xXRKaCZPaOYPdq1kniWBpD/dY92386FTMIEKse
5/6cMVWvw9Xq6uZVHvHQ1EuY5cPfonG0hghmySOLTbr1WK8N+jikQsMty0GkwpLZW7Nks98bVY9b
C1vOx1JFCfs1y76wZtjyKXZJAK4ytTkUXfu4kfIK63raO9J+BeLMhFJKMGIs99rpgp2EedJalaMe
mi9YEzYI8p4oCwuVzq+hmtluPBqfaVzgN0Oatm7Z2m4OGpEI6akGn+l0/hl0ZkzEcAIIzLMeSASG
29M5mZ8QzqpAEbq1q5J5xnRHy+sUShJN7Nq4tznUCaj8DhGvS1/EvxWzuT0qT01yDd8/r0pN16cD
DqvQbfFeF9fQ2IHI2NmGxM9D/TfaKH7SfVNt/1Awd/cvFCUcg/MHATD/PCRwoSYpXCavrZCXiKtx
4aKmQjpypAUJSbTsw9lXhJ9C6Vqv134BKOe6xRzCfiPyMYl6C6hx8juVftuLCde55cJJZzR09vR8
6nmlkRUSOaIpDQBiptm9bToMrp3aXb12c5lIGHr2P9GVE9m+/dauvZ8/jHROZEprarlXXd63/hna
5FvZkwY0OM2XPjYsjXWPFVHMTSk8kOeF2Uah/0GdJ8Zys9sihXbtH5YePCGQ5IULIgBABr1IBWP2
4DfkOiohbfobL6tThSTwUK6U8tfPmV1IJDlzWIvDOTB7leMJeRPsG+++xC69tK4ZgwTvetkxulS4
ptfOQvOV12Z+A6vyQbsWbD4RsKkrsqSKGYD3K07YPFq7z3GhRK1Fh0gvh+lpWeu5+UVt46iCKdTH
eYbT3tWn/qOF9PFilpgicBS1Szn+9LSThHA6Ar4RbrW6hXl8TVWDRoex9Fpq+ksN2qua6bDRM4P2
ZrUGTo14LBxbQ0BmW/KZwbDnAlx9LgLNuNFrPoFpqAJEjoIic3jvi7fSyXfben8+09lctmx6YtIr
epspQS2qZVLrdUz/o6pV6M+dHM2qj7qju8tRp1lZ9/tfzG+hI1o3pTsJa/5fbzElJdVqzWr1Wejf
5ONds0wAjicdrag/BuXLZO/8S3ipH6T0LhGxq9Z6Zsf1J2oNyPoxrbIPEuPFe9e5Lgr4mNTu5rzy
TnwrWP58Ex8oE3tQDA0/2VQ/egB1ka/cEgzsdKmUjYx445Q/EOAVVuK+hUeZoFP7qQjJQvnY+gqt
VZNnAkbaneA7oVlwtZ1Vz2gthfVEP/9INnfGB5bzE3uZdDHjgkARIi+MFywrs2GQwALSaVv/nxI8
hn2FwS7r0F1H3FsttfYuI8iPMd3SokV8yezV7gWYnAJkbm09d+H8SEEvea3rzzG5wC6eN5GWnZKo
RdmoOe3f5oGyUs+jlRrxt8PApGro02mIxlcbqTnqyv0UMCdbcyv1pPJOH/4uYuGaQ1AXzFne3zl7
vIn0+uPyL0t9j2xm7FhvEI6viY7ZbKu2aDwcKGoM1xompKYjHxvHQd3tDHL5iNzaadRI3qEZlBqf
GcQu3fqWgOw68IuegX6tlvy0PCwdeOzDNblgNAqmRLyVQamMgKvJ/ubB43XD1f+Fo5nghven8iGr
57vFdfUzf87bHgf3Y2EzNIkYWyDeHtUvPGzX7q2YKdEqsgx9tNNwjmPm2I6DAqqf+CVk5MvNctgX
IjkDWnDqOq0rIDS7SqSf2EYyNEsX4dj/9oXMQERuermkaj9S58AHg4RZHAAW2OhE3kIwVIlAweTb
DpEQEP60NhkT+pCHDt1yI29Qaa7mJkCF/4yE2sEs+w1hqRPk20s+NUinKrfIpqIFdlW7zspNmU4v
jpLGtACH08lkrgnqN0Yk9YmYLHwDTMdsZcWg6uLtbDjL1j+kO1L8fcB98jVdtZ3g/sT4vlKBeZTT
w1BzPBWs8QN8ffL4yAU3njB+FqV6jE6xIXAxlB53pIvjs2hDZ29iXfF53bLRj7pKcgR1nSGJ8ipv
DO5tTIKiNL2l+KoMrE8/tquIswG/7EEdQMBLsplcHTaMwA4J0ChLNpBKZ7xZ4TFb//qJRq39FSgJ
nXvYCAa4nVH+M8F8/dedtXy+cxE7rTMqjgi2fj44jQ+ca2XuSvO3xQwuL2q9CfLauvVhBLIAyPw8
5wtoRRIxxajqm+Wg+W2VO1jU6yfNth3I8solpNb9jekB5DcI2d7vyETMqtYEnpzzeGWt1G7+m9XR
NTpBfknuDXGxmc1fFei1wpTLXc2PIDEFONiD38J7VPTXJAml0s0OL4HVw+zWNghcMg7PqG0vpLrd
t4+Mdoq7VDgnsNaVYq5klJBrcU0ketYTP7fpPE2kguzbfDqV7n/DtR98tH5asH8gL7G3DgP/vdBO
IrCuhbxF3DcCud1FOBNTKGm6D0Mma1AeNBQ9kPBwGBRYe+CBM3UaVr3xApK2oN0yI9gXzjwtewBF
CGsq+7lfNxcM9MoR9sVI3ORA265ujczdkaHLFKWR+Zbu99fsS6ai3QOEazeqd6U0WEZgh869WBOZ
pSmI8IUiINY3l8k9Ehbydhr3mzFUwHN9ul/dkUXeFlSkZaxRW93fEYD90S6v2FgnhtaqBKKB1V/K
M+AXh02faxhNhfPVWWYA35p8vTi1BOYCYmxCdJe2UB8pLEWjFZP3bOondYhT4Z6XFv8umYd3di6h
6Y4ZzEmRnRvCR1mOiyxKJzfLr8v0zec8tbDeEgFawRz9yv3KcpRU/WtXH+v4bIRtfctv42oeyQV/
stfwFB9g7S2Vb2Xnruts1h1yzGwSPMFu/R6a767wCJGQ5410dixUDmhdRdfozT18IKUId9EXHoRP
0TbHMVlb7yjGpW1kAO/NS708yY6c554PRkl/YU1Ondlznp8yxvvscsendLoEK/WqVMazjX0VFCLS
1lL0VZ4QSAtVVxY54f6XMYZaeyjXacZDS4k4dx0P5e3T2/48sJvBRtRSlptcApMtgftg2NO9uH3I
QiKt33Wm+Mk7KEh5IMz3DyjYbHz+duy1si316CAUSPLiAmMAXhuJl2D1dlkkiMRdzRBBnm91qvN5
brK/AHPwAeQSGGx3RV9W+8/5+elohAv9NTFYW4rfdXCSJFnkhn1+zHRZ+uwx+xBVfv8wwOMCyJMG
NteEhCBDd6cjU2BrQE3XvlZas4YnY2qSMofHBE8rsIMivlH4w0MBBqFd7mjAyKPkkTFJOyqyCPPU
KsfpzafTJy6cSujGybPiDgqjhXF8crIpP/fxGF6PnMtv96fIdk5x0ExQVWuDNyCRgcBvwQxoytgP
/VGL5rOFmLhPe1n9s8VszXMrc8gRM+DbZtlMebc/ijiwDVcUjZMAzmtYznYTOa68GlhQPeL4ugtg
YPEjTP17TLI6gpvqyE2Nei5T2DMiMdsezFZc3F9R3Gb0Z3SozIGXAXWQIRtx934o6I8Y8GuJt/ig
SoG9Q50kiXl0dsz9olesGqXVimPh4ZLtfvx0KDA41lJT9ZYubcxCtqOtam6cjBvLNpt3ipi6fp6Q
QRVkDZC7y5mBg0c5ZknkcDTHmc8N0Lc0PDxczprqXdzeD0wag2RGeVZcYC9BsUzuLmCE9KOhtLAO
fzxWDZ0cHJs3J3I3CEktBLoLvuUmXVK5ZC2r3RScaa1SBfId8ZkaBX3pA0EN5istb0B4du7WtnFd
ezUl7EsBh46QEslWj1GbMzhM3H6qfuw/wogga6hBInVtfVHMq+ribDLV0JxzOF1AF1bVWNCKMKwC
YUw/7sk6iueHXXOIZ2EF5+Zbe9MQQoBfrEEDIPBF4OWWcso4NJYD1Q8+fMngu/HTOBFxhPgOAg1a
kerm7y+bgr/2MQrF0OxMetLuQ3wx26/tqHTLPoPsNCivhMBBS488ypjyRSSuZ/1qQSRfeZKh5MQr
jv+/Ug/tdYiLlzxbv8+LFyXvbAsub5BRbnk0wFQ8+KiwLu1frnK5G5YAXqLhObxQu2gy3nDNzKd2
eUOM77Bc14RZkW95K+lO3KWNKq/dZ/amPrdHkhqG9Zyik9yTUfMVHGDQlhOVMJrLcvb3zUPiAYIL
ULHCf8JDp+AfClOBSYryRMcwd4GTjwudM8dAu2fQcOBbS5gdgn/QekgfsIAmjOtbT60DfrJR3e/Q
crKcGt4U8gZm2g0odDYdZFFIl29U/OM+YsFtzHDGnpOt/fHPBB9WAm4oHlJihlXpZIAQ+0lXiNFx
CAP7SBNFxhCeYzBgILzzyyroSxqGBOYxF7ypv6uJ0zDWobar/qsf1ZnwR808Nehk7HH/uRiQu1BE
ib/JdEIzZiH6uCRxWxlflTiRRQ2Bnx+/book+XPFVVeIWGVf7jWd25OqdfRHGXqDhbpp/LZToepx
azjOPQ4g1QDQiOa3TaCxaC+8JwyH4a+cz0wZz941zuoGA28g6ECe+5KiK3uMVsSlexOq95IWST8g
XhrJE0VeujwlcfuTWFWetDQSB++nIYIWmO9V6q4TPVUWrTHMTWXx+JOfLj7+yozcYqfgEY1jOP7Y
BtbeeIwjF541zFupBQQnZo5rqwB5oAhnokB9gDJ7HFmfW7CcrM6NLlCjqiUh4I765KxdsQ/8qITe
koJc7F5Q4jDDY7O600N/Hr2la+Gwmzhj1+yTCd0BnmVfM92u9ZKV5IOT4TuUvL/wVzlifnRrltiR
TBslv6Qkm+yQ2SEatz4rT15O1yfZnrW5MQzhfNqzq6EdycdKEJU6JVSNnN+N1LkQGkFYrTOGX0xw
Vm2MUE8kw4BMVoY1rlkQRyXJD86CLvUMA6tXjsKw16mryl2cpQqdq3z36gmR5UJWClBP8qFNmepH
9A8JAKmQBiIKVdPbF7HEXY8RaVBQMfq2QZ4BIdKLVeaarH7l473pynIQi7EleuLX4wcFrLC3DxS5
D0pMnTLC1FyqfRWCnEM5MhC5pgwuVAti2TLuYekkD6Tji0qPUOGKY1eQNuWuXwziQGfa7h3WbTXJ
PaFZ0hW1MgCr0BxGQa5eRu5g/9yHl+TG+lNgCVxT0S4kp0Cd/BYkYex3WzlmgKOyEc2CAuM8qyps
O0w592sWlOzwU8Wq9WS63lked5RaGtO88UpX0wOG94WFxYa0PoSzCWz+eRxI2aDBFS9uJYmVJt0I
x+wyoC9123SZ67zEmWeEmmMQSIugvdbxBIJh3Z8r/wni8EyLFgjRgJGunT7iNyD52TP1cNskcyO4
QnNWMJlk5kH2SICbVZhX01mn4Z3cyPhMxH0V44nfe2hIeuN6JBmLII3xpcLJelOpEhIx6lM3m+ec
HEoHCBw2+lfmpUpgyyDMxDHsAemHqEv2vZKbIyw3VBzwrKiMLcHX6OpIWlywrbcFyBuhdnSqszsR
JkEIqqUHx9+oSMX/06bEUyZkTcg3ll8AWRQWaOVFLSec4/J7/YW6KoRNIaAG6WQb9v3snsUlobdB
U2Sa6yaPcKu4b3YAi1W2r7TVR0E1F1CQpfsah08eN8qC4zn4tRsVH925BwBFN3LMcSsdV3pUIr8P
fkDFUuWK/x/GD6cQDtJJigghqZgsKmGbmSJJfygAWcD38Po8qoKF32ZLGWs/L3iD9jxRyM3mO8kA
y8prdW6fyHMfyZKRxH4Ulgff4ZVZ6hyxB3EkVUC3Sd/I6dOnBFH0Q1bMC+OYrAJiV5gNNVRYqmku
jGrsV7LxHkhRCFDijlH70VnxqXQQDtUWU7G8OIeQ4z9l2cpTcboFoefyzCRC//CH25ZcmICkWQFh
5dq/bUHsFN6aE1LB9qkgcds1rwdp4e8FUM843kp6SpTNdDdZ9rzwkKonV0azf9y7SEGbOz+8n7x6
EaXqkVIN2onHgsnRtfawm0jOiIWCM3ezkcA2CFv+eaR9g3c4zN0J6bips19hUYmNjkHyy0rVJCzF
dFOdjjrW0YfVnyoIWtq6Jfck6W46ReM994hWEkhaO7ApYwhE8ZVxj8yZkHSbY4uCdougXqmctSZK
t0R5cvOxsgMcaVmIYAt74Zqf9+cKJqCTI4pxCsGcPMwZBlLEDpnDi7+21YuW/A+QhrrOySJXJNB8
xFKmlq0UCUbp4gGMYEHl+TB06f7qUfaLfxoOkGI4lnz3AVPqfwfI+oUzaOpbXxJlqY0pDKZ+yvVs
7PvzYRLv4jLdvn+TWpHUQbpHW5vH+M5X/MlgzCRG1GWd/W/c++2Bgkyf3717+Um6FLMlDU/lixao
EWJoCp4ggrw38WckRB4V/izA7xmV76JzzOpmEgRSb0n6Hn6noVqIQ92txn97gDy0WMofFmZixdgz
byiuZEYxiuBcmRaQM3tvplfe9h8e5ibbhmSLw0BONk5GtZty0y5aw/+xkIpl0eqp37cSZww6Na0H
zuK6abyZptke0GlEZSJNdBrydmXHJOMWsdlm0WkqYfH2SHu0yr+KsHkZvpBJHlT/USUzksEFzyDY
NO8bV59a9V1B/mL2jmJM++TtcX4EyKzxsLT4wkdy589j23BdatAuGpbEnRecQTA9yj98zhwpmly1
boq/87cugXT84Xoac77GCqqQqrxnDAtjmt8sOY45VuncRCFdgL4OgNXJeCCqDltCZNu6TdFwBQVo
SiKJwF1yUEYOaoXdnsy464PEK6GP9g5sIOC5XqYtDdFRdHVIQnFk/4MHFuA5VUjui+QTZhatPCbs
TRKjRiVSSGIpmgZvWJg2bklTuUrsMQ304Vo6+TPGvW78+RIdrBAXWRCcBLtGudj1b/s10eeIDEc3
I0diIRNIS+CyEak8Obvm8nODfqmNJkEWsLAAE9Xbznah0/PY9DpgVLN33C1ud4yGUloEmGFA4cOp
pITv9j3+T2G7b8OvZw/7OEEyQX8QiZ0unjWVA/VK0H7Izecf+LzQBxLJWg/4bUg8UpLHVmP+y/td
rsULzToctXW+05/OSVxzNxE8TE+ML1nfY88HTwJ8h9ZhRDWFDXCGWT9D4Wg4LSR8NiHYz/xEWCg5
tUA56nM774GDOow5/LXjoE/U3fajwxsZ/CmD9X3r5rhaOOjU0iEYz56+ovTgjsdEcZ15GyB/ifR3
V6edndSf6n/3zouzRm47JvIzXG36GZRvcvBdcjNYxdsnz3Cco/zpK9UVy65Aw7yLUFSO30M2owW6
cKBzrVkiyyazyZcFbqm2twjdO4Z0fbCPdNGluKsuYQfL8IyMLhxPB2bwNbuNkGEki10wEfI1Dsk/
PcJoAlSbUCaAR+F8DUguszu6GTSNkyBdaOYoncCC9vOYhu0voUgsx72OO7YhyHkFjfEy9jhPIn96
0D3SPXh38qTd36IE2h+mQlge+pMF/dZAFfltjxkQMekxf6KLF7Rk61yHb5YpZEWZXgb6TObjjdek
x6F5xbzXBCoBcKxyJ4nQBnuX+oa6dUGZEJhx9rT0s9QZLHF5KWYY9Xf/Y5W4y333/8q1Lc/nkkTR
xS5RycLM0zMLSbxkuIxS6RmmsNW0o1rjbnmOwPNx9Z4aJgAfGMCOHvEQPc1nPjvUYX6ZGgqy4q25
1gg3y+7YuzSoTwPoNIbZokwjqhF6lJsBUmzoCDoRiXG4ieunjRWlT7NFGzj0OdZ8C4kAnO14mhav
sKp0hL0GFRFc+JyUelB48m7LAIQA+8n1SI1zaV+Y1GUfxD6SywJAbmK5iU/mqCZAJOKcdc3d4Ijd
ESda+xgMUdYzLohpLYANNr58mmpRP/+Osvxo5FOFlU46/nK2uyvo+NwJKxsiu/QyqnER7reuvbDv
gnuqwzfHsUPERoWlPhGTpD0C/z0WhzcFVFQB/D+drZTLRlyBHJRpIZJIKZ6vpN92KF7B9kY2j8Q8
tj5BkOFiGovA0p2oyRSGikdihLYETaFkQlf9BJrJtAol0T6nCUQdSHHmvBL4rRi7Q4D2+Li7SyX4
rXUxNW7IuRlwayj4cWwPkpSUlzmUMD6rFdlj9cbf7tWVDhnz/CRblouRBn/UaV5lhDOREdOGbnFy
Ml2NUCs1li54/pDkkCMmKPfZmmPIiwcPNtrKGT1adWzhyzsegomcW74TP5WtxYrLxSTvFiNdFj6p
h76ZnpCT7dFKuDjbTd2ZABDM0Lv0lbMkW594zcnrX4OGZB2RkySYfFcRp3jwFuK5JnMH57/Cf8g/
+BjvACsI0FfLRZS+QitDzHK3GrF8agSSt1eapDHXB35aCkTCQUatvZNvC0ZCUVcznDHsA11k2wEt
PzQYDt+YPloxripwHlIq5sc8jRufgm7YOM4jHttPCOsucxt0qp+LlxJTuRiJPZ04+9zleRvw7Qv9
NRzpljmuHGKGSiF5K1Gz5ySDRSNlY5zpdQiEvMnvSubtB7C72L0/qO7G99FS+b7ZSmt3+oRApHGM
9HxPqNDziCxhg+Igur0SbCiygMgtAyatvKBJ1aC2SvzuAxTREyrPHaQezWlrvcHAqVWdDUdokR5s
1CJ14ZxknFiGNnnMS/XD3QW7goU7OAVuq2OaPsf8TSF5NtNTiGa3mo/RC2A0QFpIYw2MOg4zCU3P
SF27E6YvoD4f8AM7zYAIxlR4Sd4j/wz4nwnshjMJFIbXcaUYmf6wcE74+uxgGIYcWCnZ8S5YnAsY
hYeulR8jFWcwaoW79yVtrhInuJdNrzlEZz8mjkc6phOsQtFQPaWaCoY0ElnPChzPXh6KZ9Dkgl2V
6XrQMkzrQtEiqyDxpbdpFn0Lh+yiz2w272xp/h6HXtW5h5rjgBqHiKT1S2DxE/X5sKvBCOFdGabC
iIBAmbDmO+4VoipK8Xg/1Oe5SDmCryo2rv6AIvOxujHUU0kIMlnRSk6Jv9734R7PBhp6HOhkFtpD
i3MB+ZaoVH6EiM1qpqOvA9sjfVeOPJ2mPlWTPhArq8IlVyiFIbJ8HMlDcFJ2uc3nPgCYJLNVcUFg
KGvewV1tFr89+gV7B2BkF40wZQnsak5WAFGgf0t6g/3pXfXHpJDUui/x9Y0Ovy0UM/U68rV8pBLz
0ZnmZo2f3b4AewQMkBsZPBz8ppfZaB60Zs6M5JbE8fbjybiOS+TRrf3msOuoMZA97gE9FN9PauII
BGJKHJn5auOkAa5trmmNSBx6Br3ooJCUJA14lk1/9nCcOnl5B/itDifUx9uhfU6xBJtDYCVzkD0a
K0P0Dkz6BpCCOG6+EzdBhw8vPd+7mJweDASDmQFS+seHtJtgQ8DATd8qalkSIQ2tHByoHUbKg9aP
slCaij/msiDEEV/pJ/TLieIGsf2Rw/ntfPGAJ0//pUiFWL9LElAlFsk8yYXmwN/44khryqQJ/Vr6
D/QM91bFBxt+eI/oCZKkVNA+Rk0QHTdBtwRhHQBV1No2w0CnvZmyFdI1Kvs/yDRM6AGLgNTCN21J
+GvQdeI3HGqMzhEo4D3reQRNMXQKauytek9ZfolD4dPv2H//tquckc1wgzkPCc7Tu0gnkfOR+Gs4
eGkl8gyF/VXLxNdoWTQjICmNPkyzqXIgddkmhQNzSuoOHoGfVzZlGYI+fSkGo1ps1nLEx1Zaf2XX
fVWSghFxBHpt+jd0GseCMwDyg1hdBK2toT2weL/ohRczv0WVOCEC89FX4XKzeW7ySABOIQPHZcZC
ax/kPF0AyXwjOmgIz/hYz/9GKGFLqwvtmAcj1iZvL2B3/nqBKxhOvDyWb7ECB4Vb0LvKIgdfhmVF
ITN/I3lPH7t9QT3NfrirjysX77ckGfgNg50iUWKAlbv9E1nRJ2sL1n8PcA70pH/PcQZhb7iuCaLc
x8nd+4VO5+bqoL/ayt63WmZ1nyctudJIfipWhhAhGlWXXR5mt8h9q5rqN3dcL6o1Xz/dC5s1yGLI
Q68UmxjalepINafujZIojA2JcbzZzkgRifUHqw0HKHBbmYls7WI01QjysG+YMLTAzxGEiP0QFhHf
Ok6xOSgMzlnW1jAh94Fm/JOa0Zr4oinf0huWJTwOv3yeUdBobg4MAlvZ9EPbaE2YLemGu+U1wnHj
frUvZHXMfcqUBwBIeKXUQ57ID2+p9ttiipyaRmXEoasNYfBwtdOBeYQQ4PowPkh2FGrMz0vl17Xa
AkZ2BVpoW/q8HUI4SxNrNSrWM8g8xnHb2geVySNUqHj+eTDWLzdgII7SKYIDRvj6lXtsLpTvKg7J
9BKadHb7kXrqQmEdzWDYrI8REG+Fl78g44w1i0Ukkf5hXW0x9Z74jb0yl9Ug0GiL+WF4Jds3x/1a
5ytMMlZAWlaVyYybIDeYnWAuBsBl+G/ufkXUe+Bhk1ZCsFxLXpGc36ryFsNZ0kb0Ya9i1d3ZLEmJ
nm/aSRRjWzwoH01NMYaKlX5Vo2+8npOf5o6ZWX4kZgyW96ekCeiWYLr3O/3iQCIZ2Nu/W8Doq0nN
Is6ajRFFhgH9q4nLuMXu3eMFjSQOkKlHynffMsCEaGgh8PBaFwT8pIBayNxntsCBdXbDd0KzCr/Z
iyPoMTrZ9ziN+Puv+2H3zj+gEiFvBukD9IxS7jdFppI8Vr4o1sCb1ByMRaT2efbqVR8qIIM4KTsI
vsYQFPTA6KgM1ANuZCuOouuW14YtOwwgFwkjdTUt0XwrWjoaaslYsBAXHNaTOZfSqY0vG2ysvBWs
gutMI1D0jts2hh7cjblXaFaaGPw9VLGkwnTCWxMQSGyabXeT7vtriKAtCG5uoE22Ybfb8PX7lSta
k0d0iU1xHubi5VsnAZG2M4HXd0N3UDo9ToPHRb7Tl3io7pvriR+bZWLNvEJcYAYvqXFxwK+1AO+m
va0W8Yj5jgNZhMKAsU0frk9eSguL81xSpmIu0N6PAqxGwtZqTMPJFdrZDFertw6iRkvMKVOZCdt/
WLiM/kFk9GUWLB29fwcm0J42sFqkYU2u1fPhJ4MbELJp75M1ceE/83V3X0PNDYHYyNmp38nmiHHr
2DIKMwVbH76U/xI4UFBHVStn2gFURj7OpB4UU4iCjugLDyN8q17L5krA3aLHu3hevVJbz7pHHwvz
HSImMkrPN3dKAooTBDDXOUNmSCGbfapBFo6eEGCkzy0gr9x3PZ2aGrRtWTG+I3m9YtM5Lo7g3IoE
tAFM4EWo62gCxo8SXr920YJ6PSbsbzsmgUbXtMjwJGSmM9LSeWHqqHUnHMpZafKRmhiY39u+S5ya
O07SkbOWoKimeTEYLKvSdmnamCczQW1nT6SRYryPRQof5cTC0JmWhblt+TjFONhvHffNEc/n77UD
u7VyCZshma1pfdF0JglQfD6ixwh+JGFUXkQnpWoWYlwNAlxRSXD0/Fy6XcOGkWB+UA7TwGT9S7U0
wVCzPSEfaItzw/wSU9lgdoJ9mWl/ygMJxcJ75x9chIjU5/Ws9Fx4bLvIOjk5pB1Ix9umw6V7FcTr
nTL/i8EKgZUEVi+v0n4dvmCQXG8PNd+1bYdYRnzYYA+V9xxlRqDXIx4M+cGrbXXhS8OhIDOOkKUO
wpWrMjDH5ZHCfvAoTn3BM0mQns7r+wnuNTQErc5uF1C1WNEzfxFjI6izGm4PxG3PDnP3+9OeQsO8
0bg5RM30lPP/7UKgzyY/Dfm8FbtDMjS3c8L3NcneWjVYh88lQWTq9YWAqZnZAbYBuD+9ZJqSu5ZI
HKg2b3mPXEeD9uQDndQLLjgoGyxtyeaVJ8StJ1OkLOor9o7pl6r/NtZiXk0k5BGCApfCLUoCITWN
sBv9wKTJTqB3Uau2qi2JKUk0wLF65CgUZM65393ImethtuZH+JCDigbYptJ47iOcT/reW8LK8f2e
ztIig6dzPa3RvkpadecNVyeAKuswNAAYqI0/NgLmrSkorsvF6ZWmASySHZq65owXdH5cRidkD9O+
I2RuZAzD1S6u1aPvhzuWw8pYfnnCwBjNwnZjQLxF+4ASLJCypVLLt7IF3sPEfOm3cGw3OqPzkf0X
hF0DBddHYqvqg5+eMjmqvcU/aMerI6n1+HPuL4nIzCor/nfm/PZ6gZr6ZgWQGmR8ctb+KvIO4DIy
/uWcHC3GNfj1ZMb+YzO+kJN3fuF0Dw5Jmt8h++1v0gz44l12ZfEeUjXZSTDFhqwvSKn9T5MC8Y44
KTyUabNDaNLsAqcYJYV8tc7Qhd8Mmvz8fNitVD+jOP+NtL3Q4WQ8g8LnttEieOxLlafTBq+VPZ+f
odlmI2gYKYrAms7LCGy2aCiqLRC3eCLUHACdVil6HSELvyPKYPfcIsZgc7nvNUJztwhmQA7IdCzI
fwI34WZRgyXvRBJ49la3RC059LrzL+XpQqmcjPowzDWhOx9Dp4lKiXfOKHy7QzEDd2IgfWd77dEQ
VQgB9/0zTLhJxcWpIlidnWiytM5EI3Se+LLn7dWsK+dQw0KBmO6EHE8zijwkcH2rK4KMw9iyI/nW
oVS6duSj/y+ZkkzXCbGOmdfh166vDizydXnYpiflqKqIEzEu4Lp/Tzl1b8yLbgUaVGBXkCNAPtKN
0KwIZBPlDFqO2SjSMD4lJ4UIRD7UrJ0ilH7v/B187kQTehdaTlJVQlhLurs8NaiUGGwkQ0nLoMPp
Frx833d2P0p0OgPF4elrkc3KKNTN86rnlc+p5O90EPB1U2OCaGJMFZNgTqWORlFfrhFW62Zt3cL8
hdg+eJ6gyKA3uCkejUIOP18ssn9KqNcXxCPqLb0KsIVxrmzy64iiT0qgTUfL5xsZRiR6iN3BPloz
Hi7NU34tMBTBKhpzL7PK1Nxud4ZPd5S7RWmdR/Oe4MP5ObBF+Wi7kGwtsNYpKAP1vDLaqJ2FBnDE
sm8R8jmSSzLS88aqODD3E0Eje1YJUavqeOsaFDroCM/HYAr01ZDHs8VU04dpl2gysJxA8QeXM0cW
uW6SODRZ4rHd0KXvIIKkwki+PiBq5eE2U504aGANtfli2+WBJwuilmNwjDZPFenlIjix1reENEt8
ERkZopkhKcREPkw6P8W85XOj/UZyKZm8v7xiX7uPBCNRCWq1a5y0PhaLCNM4NARK4a2NeL1CFL+M
mJUcJsQuAnSfa0NRwJySfsieFPRJkx01agqvIv3Ln4SP7ESDTSROWNEEEE5VpqjrOEmWECI9pQg4
x4nGsxFgEnko1KODXFzS3cBSoUVQv6qTPtRCSInH6rAzG0T/urs+mKrmpr/eRPPqvjzG7GENvBZB
L5dW60QCg54wH2gnO+GR+grc1gZxMCuEg6s25sFYTd5pQ67WC9G3x95VITHR7BJDKrbQrFTj0f3F
2GMFYXBniaEzjII5xqTeyt2qVJYrWb0Etflpf3FbVUnfSYnET/ml1RKGtk9aym6GtIwfzCAD7wNA
PBmSshX3eFGbegQNH8t12PSe/wG8c7bk+NN1dRoSH7etsT/oTrfE8fa5hmCoX43+3voxMnyvgsdn
VDz6ur/x4DwCwG5LEX0vXqrYNR7FWni0RvgUoXU/V/0KgT5p1xvj88pOy0pIXKRSuW6/OzGVCdmG
e62Hfe3aLYKYpgSAgKA0qaBkhpVb9f1MeoMUvC356GKvKqmrgRIn0BRyIZfdJbS4YUr0B74967Cg
20EH8izNyzzWN2f/rSOhNUAVBPmy8LV0PN4BeJA6tznkjFRkjWAwxg3XVy4WNxbs5VFBaXfPMJmx
aMn/ozMemA9WV9ciXFdlbiFYusKp1WOXwmvXvuPIRcLEnlHN94Fe6DcvHaSA8oJ48BgQC2bY3JVS
qDnBT8osEFnM1qQwajtyZdV5sqOMzGwV0WTJSZ6PBQJvcZDR4+dh/RqcJJlC5wLQ4h1/YauUWItX
ESO3Q7rMXSlV8gLxA+mb3Lg1ve6UlUAD82WZlw1hHX8oh1ydE4K8g1L8Dqxdi7lQOKB++HCQ4LbZ
RCuVvVXcS2bScrbMHVsVrArX8NH3dYcwd2q1+K7KGqJHKJpQ/p4aYxVT/6NEoKMyRfehk8xHeWyn
KyXv9wiXicFCbYBFpmu5pv1swrJKDYZe6PhUYHMmNis0kqCoV6Hvs4v1fc8JFo3AtATkbxucJjDT
63cIaN3c7FX10mlDhVOcKajMj8NnqSalZ8+vpTqvko56sPYWtBodIAa3IPIkrNvdMphYj5iIt7RS
reLkaBkoTPbPe7fGhNptKUWAxP24kbWNbo3GNs4wWqghxwQK5a8kwlKWF8BVJJdoepCgaDak6lp7
ST5RoDDxUiSpVeGnsD1VUITquKCtIUHup+TrAv2NzTq0duTITDIDCp09CcZs/GBXqE3t4EHACLhL
Y1PaT4Nw07fFzvm3uE9VChQiY0Qa860Y8xB7VfL+ICdNSDN7MYPFeXncnuyxIxzPhj6BtsFV4ZWY
mwpD8ZWz+KKVV/pelNQfYtJwKBsxnaU6mabwevdUnGn00V6BWBp+kyixOqaVmRdMu60NHPzN3k+H
BxJ1r0tQSGNBpU1J3imx0h5imZLABezMu8YGQMw8LLdcBzNVwOxArRcWb/BEq79srcBJoUsGC2WY
TiQ4C4IZQ1ISLaEdY29ehqaw3b9grqsxixgydPIy2jPoULHLi+0gSZVLmoeZQIMBVJjDsQM2ouZR
x55e16BPyq8vHnZOnDTRzUKPVO7+ox0i82RNfcoB39410X1sbXTZ+ztg6Tq7+ztcnNjFs8Ko7siA
uecAOSIheLyuGdL8pSHs/+u9zIdL0brOdVpOCLTWrqrIpHVviUvr4JGs/5ckVTtyPaAESR5ftzVz
aAWDns0nrouq8+JBLJWfW6hxSHh053hj2cN9HHVd7gQfZ9QJi7fXjw66H6pOhE8+14eCj/erV2/O
8Vpb8vmyn9vBSO4I59Uud7qSK/sYmsF2LlwoibiwarKsfVtoDinYqEq0AWT005D9l5SwX0EMS7+W
2ZmHU3DHBrDiPgOyyBL5gYUJihXieI6aTuSINF6N+BBjhcYxIEs37cNqWGlOr5jjcpJxIwJYzHkW
jdd8ozkPpZKMgoyw+D3GV/MZkrnDQMFLLdV2iz9J3MYJEaiZRfZBipW0TgeG3qrxD2lpEsWrcTpY
Ct/b/pXPXnukUflj9ZK9FPvst1KGWcOoCctqRJTPnwO8bangP+x18IP3nguloM2xQKWFSfyVw9+B
E5LpWIzSTfwgJZzqyeWYyCwg/a6Bh/v/4m+dV9hnd8utMMyc/HVWWGE9Kp0YwOCq9r2kLtL9cTmD
TosWY2sxZeL2MTgQPaFeB6dveP4nn/i5ZuHjGI9vBH+o6T9Y/HlmLGbKQlH7XErtylSqIJ5HhVvK
Ekff7RYEbYTHobyvcxPiJHjvVQX5AaGupwyb6qGJbGSwBrk8zivxl233W//yO11vFnl2jIY5aU51
GH2VN4I1dgV0ToYtrONtg3aIna1+ihPmtiyjVrwagRW2NJOTLW26azNVYNEaWlptppqS+ffZeZ50
MsOQYSo8ZUex9SWY/vUj5IYmfNE/KE5N942Ku/ym5W7f+6DIXVA/5CrEaOIwa+pGVKKIn8yieOh+
OdwW5fCTWgN46Ise5k2oOplC0e9yVa+OR8lFWriesE2i3n5V4N7ISmmt+siZ8C8f50/gqYzKodqE
PMVzBw6zeBCf3N7DNp0SekMjj9h6AiHZ9ruQnzfH41TY+434N5DH9oWDAdoTQBwP8sBW8bOKBXG5
HHWQnKINvVaqCCyFQSEu588/8uN9T+cGxoozKClcFGbUg3LzcO5GyViwO/31q/NBZ7ls5oqwyblD
bYcY58OeeKmDVpdM39eYhkpg3eTgPkq8wzbEHh/JANVGL7m7i1eockUhsEITuSnsAEYxgGj55XYe
zSQH16WdVInj65vColnZZzDugwcQKbNl0BD6ZpJ+SOKrTv+uQisW+wWAEPCJXqr+wHaxW+hvJDcZ
KzkjKRpoYoYHaH7HDUPHERCftPGIETnI6v3R5VwX+/WBzXb3nelIw9bQMzk+EboxZ9OwF03G+rZR
MgHEO3BDHz9RxE58NxIjOaki0XQyNoDwqlbv2mx2DqV86q/6hDUT6EVUvVKsAC1WWz2/ed1mOAl8
D7xVs3Nbv4oFjsWHRKOjUPY+Mikh+/+3zB9yNqfvOi8b59QUh4SHCQxeAua7Qc8buREjIwyGeSpZ
fcXOrvPTBmCDy7dQimErfeS3gkMpia6CAAiRVHADhX62mR+FIURgR6NuloYfRLly6v/4LiZoVLOd
SffAJ0pU8eDEZbhcFL10BAtFY02BhYLvQ9oLdJg+8VerIChJz9ez3EAxhNZx6qusx5PBpic6pzVm
A1WrwI89xncsP5OntlY2Gx0eIGe0/MsZJ6SlnLqGU9awLgN9GymPYYOVFTeMk0YIjsuwd+Zv2zTc
l+5ZczKvjHvW71e1vGQl5zjk2jFAUqf8sLoiNphf/ZehWt4VOm1RG5osJ+UtwZT8LJEOnLsGd7hY
oIQ4cPm2PXMRe/U5uMOyh/121dzdsTC6o2S9uJ4Jw0PHsyjYFaLN/PGBor5djXUlIwXZUA26MXUL
Gsng7P1vi5+rOpTvikexA7ZofaqoxuSj7x6qDumGIigj8g/QT7S26f2tn7jcLssG2RlEVmaYznPG
E2siMEPO8jN/iau2cBY0EfaWkmMOs2dSM0CbxdzG5Yg4EkDX8+QDepCbl/drIu3vMB6txPF1kAUS
CSuEJKklLclfh+EyNJ/tT6CMMTkmpZZQWG2Tb2iylg5hP8qqqN21yzBfuyg71E9zkm6h23Cuy8WY
kK1GV7aV0RCdCi+ZIw0jMhZzueH1rwGLwQksEOu5k35f/gO8y4Pt5YZ7TYTPH4bfYfxpAG3jlM7v
BRYdxsUnItFQL9CH4nisTfRmmlqfjpCedXxAa9EUc1zm0J/jSpQs6h9I3VUBwpEHvY6Q/7Uzibns
EYU14lwFh/9wHeyPEdS6bsxGNGZncd31ylsA1tFFk16leLQNIfZ3OcsjxMcm8ZuRBKZ61v1NbbQ0
uEF59E6K4nfEtxCIkDCwlE5TQpgEC1jR+FYX57LAmqcett68SVMigl6aj07xLl8+xmtNThMvrkJC
xNZgqZ+jgvaXjqR7lOkfVMz2ZWeRHjJZHxceKMJSTt7u8wKbIydUHi7Fo6XQkW5ddm+tl28i3iP8
x88YaCDCkqdSE9TgzYYyH+cYXpUKbVspD3NfLK55IQpYpoHjg3L4bo4hJ+K57+OeZkuko2UW4q4a
KiW+MePxxXVIlvebkoGxyUoSejm8aQ+R0+OFIcU+XlZssExFFPDealBSPvTfJazolyOpRajyCf7N
RZfT9INfSjy9NgozAq5FKQJw27KtbvempzY7ywgsW667NROK6XHE+fzsaJrZCoNLZoYXj9QZSZmY
K4Mxlt+jVPxjNrUNZvLJ+5ufA0TYvCCZXfrL+C5pY4tUBwtZmRfMJ4LwbJAc2tnHTqz4OH0Z78iE
r6rRv/AVCcw/mae3zdVz41gmb+PU64DkyJS5MLpLsbaiOBneu/uFQ+SuupBTaJpHATMnXAphdmsm
InOAWMynLr/fXtcXCzWDQ82oTepB48yjuCssQDBMTsaWV4ogPHzRMKJxCk0LLO7JPW7kblrcayG2
UMdy7KQjpTVLrdT2euf2rM1C66CmDHMa/w9gDsaI9/+yVrdqfKqdoy7y+wvF7+qltVwN1po08105
1B3GetFoRxKVEOM8vXK0/C6gVt1epTY6zwUQjm1uNX8xQE/0A2mqwd6zaHov+DiIHcEv4CASEt7d
VOg3b2b86IiNJJxh3+jlJwbBdd1SLLkIF+u59ipiNVVPXDb3c24MMcD4mTvyoJdsV1sqx7Ah/BnR
TLCqxletvkJV7zuh1cnTFWWtERfJm5NidR8ugKSnuxZpJHnH3JjlJ5tOM1mgDtx+EM9Zw6kvKkwR
HAntMPaZm9r0+/asY7BNuVKbuPXprhadOGgJLaqSCe0Gv58ZdVDwOQNbX/x6djeC6RgiUvPjuOn1
1KLGFFO2Euh7ylbuU/CrcRx+9yGIfesY8oz8LpGxHMlGNPbAiFsO5gjtd9AxjinuQLz7s9nBTJDl
enQqFbTBBNmSVtSYu4vXrLDyyLXu8BezbkpKd6aQiGiC1F5QhZeF6Ede9pKTy0ackxCBGvgETXjW
yfJ4Pc/mlpOMUUVbR8OhQmXGdAuiiCX8EwNmxgCGiXvPwEzbHwWN9e99idbpgHLPf5tzTaK0VfS6
TBY8HNqSzWH1YKPK1BXDR/1saQfEHnYFNEhQqAiWecwsLGH5WMp6DMa3PdJ9O7+Pzx5YJ+PJEIk8
Y8zuK87J9JzwKI9vgrks2v3GLX5JfmG3/oXhvXZ0T6RUi94G4tsKeBHdKDKTd85RQuRWUlZVwgOf
TJCBISFUB+gOqh0ay/1CjiL/sZtTGOtg0W62nUSvPapCWlYcrYAaL2cRZRzoQlw6bYo7SEKRkkyD
HMaZtnemo4qNxJuHXRIujYoAztwrA8c7kY1HFq0Hdne5YNKtF4ZQg5s5MhK6Le8xrlljEfGagdV7
S7d0RfzPvFLskWWmd4fodB8LEkU2fahNFckgB2aXx86pG9OyJ024wTSYIf4RbpMothtS87RXvoRa
RvQvdpyUA5AbgQRGtqUt0Adf+jJZz6i4JfPwS4OY4p5ErI8Mot99ujt1TLs0NNveH34bNh8X3hSO
Qtu4xkjzN0D29Q/VR/Mvi2AeSeBnmYTBvdHDTvglizuuG+nnlW30LXyLPXcKHLIenaEPH5BjNHPI
kAjifqoo1UmvZvnWr5aa2wHaLT0W6kagGml4Ku3ihZFs/avkkTtcCIxfvkIjNy9FMiOW6a/O7hJy
6MbPcLRLvh9TWVMObQKL4LsJEMb+pOUAIAMcMFPnGgL9YvDQvXKu2MzKJeelwLbzQiMFg9O5fq1q
JkB+CrGcz9/kI382fUZxfUbdt5um8or5teCqqHifLtCISsr3psYHwLpH/iwQTMr9gpknnJAz7woM
mW1MaULeq++jV+MxU8lTvOyDIr0F1vbqdJcGr8tWukBWTIaxqo13HUR+i9YZ173JLeASmheeK8IP
64z4QQJnpFcK9+pKliwY3TxT2bTfkOwXgIDFzkrKtoAc6j5FFbWC1bYtLoScIARNbNntbdeh4Uum
vMk1U66BzPFAWx2vVjU03lSmNmhrjrvFEvKwm/irsEkdIAqvSYZNmiI/JRrVreayqpd716JWay41
wz71Y/DNx108/WPngPqCP+FNXNReube0RLTIIgKlUMXWvY687A1UuqCVZA+t4XTQltwrNTBmc1m8
VkNE5sRvyrp+lf5H33Pl7HScfAf+aQxceNY0uQ5B7PE+gNKK/rZGmILS3aHU/v+kcFDWgvpq5Uky
T1sYmTQsc2OBN4AY5NaVk/aDGW+JR6pNtUg5d0GTaZY0c+gVCeHa1fe7bmvNw/tgATiOZ1i1AOOp
ItlRnc3QBANEs+wLUfpal7eJUNRSG1zy37Y+GjvSBLH46i22eQjlnJGus1333NDPllIRKNq6Kon8
97r2wS7nAPGF9vuOjDHOVagr5MX+H5X/44gDWf2BLCzfeFuqfSPfil2GtxaxzpBQUFrN0Ni+E8e+
IMj53YpUCjLtDemZg0NFmEHCh3oWpxpDVUVzJA4/RZuoVymFBvehCnWs5xlQe5aBYmh70orrHmdt
PeEl8QD6AJZUtaWsOqJsFSUMUjQc+2Ha/uQOK3M/aCjgdKIuMGaQmgBibcNexcBEViPe089juLQr
ZTowqYL/COYkT5XbAP1NDWRkgpI/MvHHyrP/t1et+/08FyPtxybOBs9d77W4Ja9heGOx3Q2Pd457
jHpzM3hxVdzTEGzrvkGY/kSQOx3vqOzvqjA7b5JevD4QGy1ANr6Fw62ybgjz+qljpIdISmUzVqcv
z5AnO9FXnuZI3UwNfgCWNjxJiO/KA8gG/stkPcTqkWaBZ055YZ9HfQbSurHtrzWG8HHYv5zyqsGn
y+CkL1MdLHWtVCU1TDYop5mmnobSpOGYW6kiEq69V294ekqg0QUhaUNezm972Vz8wWmIRXdckNA4
N7i1hA3BdDybL0RVjknDTLn1cFBBbYveFnR6efjXHcfeSPPmOQEedS+q149Uu5TxZpFFowaP7U4w
hQqXq3S80eX/3iboZN1os1YPruyI7a7yg2TMJmpEjJGquxpxh+AM7tPC3saBB30DmsHlfueEtlrz
1LMf7c1+kmL7Z1yvBvTKHd8wrkMvlGuoocHspQ4l1tnylxIiTFjqzM3rcwSRR6FRwbEMx7A7/cl6
qOEjxLtw7Xwvs6dETFKrZuLQ8BfBbyAAEX3biIqIvGEW8Wv0rPjCYsjsLr+YxchF9F2foJmzE+M7
NPZJxVCy52zH8HMlNrBIkZ5Sg/RHZ4CqdaplTcKFxoL9sbF+MUf6zdjjA4i9j7DX3MWWoIs+bglr
wqk+7ie5Y9U2C6jBodrLLbPGDx7Fb/Sg3GtebnRtxNUP7BpVBOEcu044BbgRVS6A+6DbBceTrVep
KWu6ZSVrjWVVpiMMH1rxQ4RTyrKo5KSgJFZzJC1ESuMC9ViBTG66dvKziFsmrUhNPcH1cU07CiW/
xcBLb0/8ZxmkXK+WlnEZkxahPy2xU2UoNzyC23zb6bhs14yI+PJsRJr6fTTKn7Wdh5toh6w1Ev2A
UxCJqukS4ClLB2AR3Ng0YqmopEWyvpQft2mh0RPYeIc936Tn7ZZu+EBA3LhMnSqP/SOgxbLwDzkR
gll/YVtHqsUNTnaOVmP51M80YZzyy2ev9yBTeuqGHgJfjmNmtuj+UkzcVDGjKQ3eTpVCkb3xE5bD
kcVaT0xa6px7UQ4+SMhIDmkOpyU635lTQW65cXknju/JZppO09ZRpNE2hewk8gD4s5s4SCVc5UZE
ZZ+42oNCgVAt4TfRIxKx6jP/gpUr13KLTu4ZV7rPNtvgwta3MfTPy1PDwsqwE+649H4YtN+feGkF
7tx4Rjs7yCnybbqz4IYlaIfDELmqh2F0qwWf0ne1S3U2Qx1UH3rECk8+HxD05s9AKZM11xtZJzCe
OKLYbm38+FRw8JnN+Z04iL1fmqRbzA4z9g4GNyLPVIX8JgYU87pT8FIBgn6CpuICMcxyVmNr+s67
XyEXuUIH4ex9xHxRTjtCczzAIeIL5lHTtIAdH8SPVKQpAarLDNaFFoI9ZZsJ0dKELKFZWQbX2Y9l
VpckJh6j63qi1o/YEDDLpRUcH6nOrTVP9CgeWGS8opCG45zNsCj3xgzil4G5NZs2k52qI3hQh2B7
5YZcffphyZ35P2AfQVlviW5xkAcbGAlJomrwW8XhrFF2hmKB7m6p1iec6CxeXuYFa502PoiPJuBu
dGau/pjo8uEjAPPfcTOPj/7UvaP482Yisldnk0+R1VD4vf3ByaLzQFkSWbKaRLQxyC2y6LA+/vX+
3Ycb1PGQYWZGBk/DW5xPpR+OagYN5VoKaXW0s1mVw4UPNUlYzgUxAwqSKUmz+Rir8VPZTAZi9PMI
XUji6WUp54xAECqzIAS5e6/gf4GlctrVOc07OL+D3990SuJ0jkxZDm5RtzIa/o9wc9n8Am57trH5
gqeL1/AjAfJ3whIZ2jSq217T88e2VA3u0UkaQKwj0WhvIR//wqZJWQN8/lMzLl8KKBs21PNLv5Yy
GospC7JCNo5oVAj8zolaDVdXNJJEnJRjgSGotvdgBZs35xoQMWO8PisIQKQIs4BZZ9/XBrlf8szA
rSXGyRCkc7Wdx1SPeXbiXWQ8LHsi6rrRv3gmS5gEugJlcqbRBcSYjtkon7VnWC+a/TuyZQVQyKiR
AeS0uLiJxQ8S7VrMKvLLTQjAbGZ40vMmzYdqFjaNBUY1XFLGgtw3j55awTd+L7DgczLoyxBBXToy
II7KEiBlb9Ho/J34aIaUzChCoVLPagXnpzCle0JcfL+Wurp7q2sEVuxWve0rWRlWOpDkNJeZ0h1v
aEQ+/cQMKAEdjR+HnWwIw0RUu4yo8TqpmHCB0lhX0C1hiBi64mPOctxBYu+dSZNs40Zvmoq6k5Fc
bk32/sr46W1tjraJw6NIlN0OHT4zDbZDhqMD7ZiPy1QIZ32AyZ45kofAAIMPzuqFrUuF31DJWZ4n
lTP8/rolc5vUZArWBZZkxyOcgr+bkO5osaU5wJAB4V/JgtuycPlMd9XniTXlnSyEfs7JlbgJ7Dh6
JsgLmogq4McexNRMnkgUjhxugupcNdZhkf4FXJwHTTVD9JrMptWs5UbS2qhWUYsrho5Rj4ExufTT
P4cEK689hGxBquUFMq/hHkaJQDYBKn/BpSKtOOrhR7AuENXnhpkm7dFdj/0AhFloNU9eu7frcqIC
P8OD9V+OnJG0KRdU/uF4AJeAPosSPLAwSjo9GeXV5DHGhn6vin5Qlz3dZV3CsdjIUI3MFVcSNd6F
+3cTlZ1SEgIharMATOo+asiU2TraE8BI8/t4k7wFQpyA4uMHo7axEkg7/as9D4OQfN2M9O1DI8z4
oR5Sew3Ql57fH89hrP3WP0l76CVBPBmnK/FizTNXvjPcLpC+7EWqXBoeLJnTKKX7+XgR+s91XY4g
CZjSstVEem5/8vjpVXKXEOje7FISTXcCINXPCxYZF8/cCkA4n0I+nXzLKCEpprYcu4gtNzpIFVeB
qFb3g3wROEAvknNeRmufivQVYrL/nNwqBVDRfctfvzhYxJjfv03j3HF2LJG3dJ49wG1MbGkA6QuP
s6hW8m1YKr3sKWi/4a8bzhizlsEuihASryX1yBQsL0xPBbG/BOcHMB50+5MuQviO5N7y7tuDiVrS
4NtJipSMbVllcbo/MOJ4k2OvVm+1e+sulHMtbaJjpMZd9dVvhCRlSDTfYxymglTmgsSzVwdu4gqs
AqnVG3bt2nYGJ8EzbsWUezl1RK5AWeM8apYvyJslLgX7Y1SzHuEf4fQKZ3p9FSJHFNyOgzntSpXJ
ylALCs7odAImQCCPFHWMFTDzXBVWus26v5ymt1plB87NIrjLBRefUr6GyfZ3mwdYDyp3f6iNqO4m
ewUHvZbaBX4BsTXhMgzp/x+F014YQDZ8NydKg89mO4m87C1IhlLVU8a1xO9bbJj51lHe1mf2sp34
5oQTjMd+x5D4GO2f97kc/mgHfTwMFrwlnLPECiXNkjIgKXaLkD4MTZQzdS0LOW7oXbXJe+gFjJhp
2xWeu+JRLnSpDf3W6Hk0S4Jd2YudGV2FntjDWUbgnRLQc/cl3g+DpsJWgCPFLk2Hmfk4rOuCGu+1
u5d89nqyjtODfmxs4XUrLJFmL+hUXUHOVGkxwE2MAYVfVwuIpDNdRnlL9Ca6Im1hmf25Y29Wqu8x
JHcf/Pr9SEzbUslUXL3QqDg4p/6Iky+F5dqs+tmfM9m39Xnow9/z48hQFZxltRGpq7VNANvu4Lxl
2pCyPqYKI8qEn4mNXJbpCMgkevdKUIz3DW/tEC0d/g8Hz4R5sodTAhrltKMCg2e51QKroNPxa248
n4C4jDGYsfHKM+4U7LxPe9GbaAwRHF0Goyzcnk6LMO8emR9/inFfdEVN+UR/86kE9ixG3rjV/HS3
YgluIFAL94SmWelqeArXdE8GcsoAiK2cVSfkk3UV25MnLD2iDWDR22PxD82Xg+3loH+CoGyWCXVb
KRT2TmAFF7yCeyqXAPUQBv52OWvtAjBjQwKsiYxBYnRA/mE67L6GUFjVHIenuwZxnn95ezHMDGEm
24B0K6W4f7GLPH2Qm3uocXBG9m4Ux8TYMYWzD2rH0d8om7qySu26g/0WsJSQucHQgY3gl7s3XE5Q
TtTqbkYvZA+gstKyBQfLvD5QhrcvQspXas4eNflX211ZR7H1vVM+tPAkYLzFthb42InOkX11Pega
5APR3bGXvl+2AKWwvnv39VP65xppRluJFKUh55Y2xfmetKDKoQxRBip43GwWB3wijQhIZpg5XrLZ
LRs57B8thMG6ffHi+vSbS8O72HFF0sz+biP7/CRRk7nGDCpDYvoDxicye0JQ5kQcoZoMGtNYFe/w
EqCEq3WNqQsXEGctv6lJYGc9hUWMekvTxcGikyHoOVyFnYyMl435SOMKgkKi2es40S1ckv0SXsDF
txYwKTOigZc4LEI7iyEAoPBShHXYgT3OGjceH4qMrzUBVfEq5ULiE+4s4W9Wgcd5uCpQsJcvUZO3
HWZculhYaUhZJ98//HFZsWs4w8uHn+i78fEk3+JtI0dBLZpNSTaiZghPVs15xUu0hE35xaQeDBr0
XXskmKyTfvH+PPM1W1RG/rqBUoWBPCu3I2MkW8m4cRIEDTZr2jHebfkrNuXCcBamWJVRpcjlJu+K
MNuOlvqj273HwiDze5ErOHEV+8roJpIEXkh64lMgNYKMjbMHrrrWc6/D/5hggw07BzSdBbqfhJZ3
C9+HaUljPDlNo8Po9Weui1VZN99lm0o4K369m2k6kRg6j4hbMHC55mCUFQyu3Bw+lCIzVRaQVFwM
eBAkV/8cYIopYQ5mxe7d3upHPNA2dXy3vjsadST154mY7gWbtnoR7opvvcxVjDn9BXQG0NzL2WF/
mZQ3RaSbryEoVATOqRIlg0FRbHEV6NLn3lQvQScaxDUPn9UfDM1UhE6cgRrHV+fA/LT5vPT3cwqM
m0NfsKsmW2z03Alp2hf6Ilk2pfW7mXiJilmr/hZvZYQjzarz1jukL2XitLKCto6W2RzD6PfWhnVS
VBHdghzPDuzDzYnHailhGEFLFHu/xbOgBc1TrP2dyNPaOL8pvO82cwDTv+ZJzbhVSXzWbWQTRRMY
Ed0tEKVvjrdTRqYkFN94vavQ/tdBZe36BCS5I5/7mgOiO/+jWCGfkTMDA6J9ZlDvccovbbLpLN+w
Gb+mGOAUPjEb7yaWAS+qjJprmMmMO6SSnzRA+eq0LmVnUHvZXh7XTsy9f4/e8xEK12yIboA+im6j
iXC8UaN72JUql4e6zdUaFTyuRHNHhm6UYRlPNEuZoGFXJZn260ewlPCi8JOJ11u5y8rHv3oZJEgM
HVliTtaweB/5RruscOMfJcSMhAnQiFoGpcRW7c592FC4162q5wEGp0ELNesNZYITtyOkV2/3Bw3J
p/ym3wBQ9fO4CDn6MFYJT5sOHSN8H1YLTp3Bz6gpTsKPnTm8WnDLbG7AiadrEk1AZ/a/ajQ2SOIo
ZLgtzLvWQQbGVWoaLeBjKtepzhzTVP5oh37vhHC/0sU2d4d3NOr5CecdqbM8iC8EFpsqEN+e165h
mrsjKNxnPNxG7QKlBVp9d95u1n6H80VkjRLLsim2gWVnencMAhGrBOToiGq2XtP5k2EiWQVWDX1L
XDnIUyooCYN4q0/xPYPNmGMBmumj2nJHD2zu/dIu8vV32VOlx4iBO500brGA2nIhVFvUU0gDXu1W
OYxUlwvyvXFSTYmX++Pmpx6aos7VFWBUJVuHSfwssBQjuFlxKMQuaAb6yau58/Fv/jsertLoN1DD
KZzP91mT0vcszkEvX1V/AuMHiQD0Pt+8FQaTSotr07JSFIwLwzQPx4AzxoQ4jXMUTyPglc84hBSL
D6ZOU6ByEmVHoT89qEfUnA1K1H1v6BvDaSWoZDw4MJZoAWMi1UF8cRPhdiMOoSM6HU7c5pnZL612
hN7fpybR6dusSAlo8Ps11SFQ1y+qW+74vGleMhrv4LiQQgp1eqlnda7bhDOrw/Lh+Ar739Cmo0at
W7NUzN3OTKEujq0hG6A5dCDQO9KvYlYae1po3XJD59qD8V4KaE2JkxjlbHy3Y1F4QcPcu2AMoF87
9cLQMC2uNeurw/eitQMY2jATcgkXEWCDZPXtBoIfWXUtNdgOWPv4/dfVWmYkCk+V1eW2LVp/V0tB
R7RKyRGcoVaRVWDRmTGrCJW9lOYFrHhXwrL47li0oWLemjCVtejmVdU3ottdkgIBRlPwGhacsC2p
FNtb8lYCDbUsgXeiZXgHTxxOBGA5DhmeQ6D5SLCIL090EdKTmL2+vvByK+iwbw1eIAdBQgQ+DQG9
RrF5MofVyUWNHK5GYX5qrWzAxpuPwPXfJ/76XJFQAsElzOW1s0JJQgdTAnHfGBPW5/NaHaqSv9RC
KVzPzWRCPS23J63aVXi1Pta2qLmAgym1R2MYfhcm7bvqtcnHaPe82ckaqgTf1KfglYGjfxBYAv6A
P2dRSMIJs7ERjRmmxUy/EhRL0Q9sxKw1k8MoAex7Od/NFYqAEWjpY8jsVngbBekB3MvmbLuA8bIW
6LoCGZicpuYUev7MOBfkCSMK5KdKd1IG9gnoqEnB877rm3VpiXQuS+YsE5aFNDZ86uUyj2HFJQe9
ORNELRiAsfbWq9ArQE7r+dthPumhDaJS5AOIquI2Z7blFRKxKLMKGTpnsidri/Up9yn3MvZRq3Rk
HK/rO2eP4AN1f5jSlJjgdedfK06Rk4tZnxyz5d6mRG+FeW9avDY3AvMp80kmRVPmpbV9+Ps51lgO
lsuF/WrTZrlSeCF9X0qmQsM8lsLDk1AvIYTD3pmr68owFyz1NuZhpFk1PE4oAgw8i/t4snKAgrbw
thPjxtd7EoVttwoWijBKclhITMWVPl7EQnfvlpjTXOHJTFz+WEPZy389nwixNFcbtStX4wqQHoXU
77dzPt4/lHWWj9um0YXjCmui6nsRBd9cQp39XqsLiHZcelIBpywkT1GIgUpctvGuPDrPEMSXvjJu
ynhpDrGVe3GARhjEkYRnNFgkdFsQksaLSUSKTJAG2mTTUzIz8ypNB+xDsMnlC0ZReZCJErFFS4ku
rx5bdwltiFrwLSgrNVAZz1wz+/tdoO37m/bDT7x1wvzimh9eXMNBch+vBgXcTkBQZV9YeReSNhvh
kNt8YKKa0Smy7IWmeSeyIhH8fM2uBufIXYQ8welcDBH4oJW8dukdtsNLgYSSyM/7KI9sWEAMbO1S
e4aKgPEbXe1KXTA2Ds7lD4se9UN602yCdnOmgEYtEauDQGB7fsJ8G38+N4KLgsr7kZ1gcdezCpTL
OjCNqsaGPt39OqwyqLvwQAYsemKhGWWk7BLEnkvTR5vcT12dO65bZ2xFCQzF/qCGkfJZAJB7t+zc
B0jqSyxSjSYlc+yjmEavpZTO7MewpQY+Jblp3jE28GS7A/GLkC9bfKn9+1bFGdmQ5bM8mdrelhUh
EQqd3N+Ha1hWmlP+4g2oJRUf/53Ax6Ni/9xMpiAq2KBvuqSKsl3bgcKXm2VfGh8tC/XtjFf8DpMW
f6WiPirOtyIiRF5edAcopVTuh4vXdrrzGzR1j7qIILGGAsB3HftNMwBXlOAWWcj7OxP+gfP0Xyf6
tKEA04Ljsz6yoG+lpy+oqAu3RnprpW3uH0UHRI/kfiSKfnRzLVShWZXRZUwzfRAusmA3wfMlXsmS
XuW8X24NVJLKQcYWisS16lzZTOIU9q0bUjacj58JlOqWuUN+Uy2h91OMxbPf27HX09Gn1hWRbmtO
gjdRPFB08zL+PSz701y7zfAqk5eNXt2uTIWHDUnXkPha3dLXjnapQIRvSrANpaxJvED+tXqUYsxJ
xEoO3ZsR5pw21HWwc8h5yzFgM7qwuUiubPgfkwKyuC0NEfN+8ikDDaAY0Ktc5RTqtTKtraq1xz70
H8c5EEfV2ij20XOdrKaDZUShCMXlK8AN4JHPYaCoUL8qoo1xA10faqw+CB6qNvWcSF8ZUR7kOJoQ
JrUTTQU2VwVhQhsY3TcAJmS92irydRrWaqaPgrirdrDFzyk83sx6FQGbSbm7mFxXcgh31hL77OeX
W1Mj0JJppflVaAObLHejJCb90QfcJDFkE26R7PR6m00vQFHldT7wtV2gStM5Ss/Ye1eoXTOQFyXf
NFhjmb0x8AiROZMyp5XyQn7F6trG4KTsYoRixcZWwUkwKcAp4QXxcOLZfdrHh0bDzYetGA141O2J
HmoOAvEO41YnKRhERMRsC7EcmkjqLxCM9j2kk5o0uHKyl7jSVnrBfdLv10OxEaiBAY/u6rtTUc92
R210x+AGZQ6Rlicp9JTUL7DOkbvyeFJ7gRp389EXoT405la0pnNc1SLqAcvfRR0chkVkKTaRqzdY
pvOXN8H+fwKU3nxA6MxuCplSEQEN0ANk4UJ0A9zfW8Zv8oNOwKqsaUyq+BweS/ztKWnZ8lLd3H0H
+9u3/NXr8qrAk2HdR1iQtnGKspD2sza+5gIVu+nBRSsy2LZXrjGgab6BY9UqcwcFJrCCDcoz1Unp
aJ3AICbwPYygnSjEocBNpUsu/o+mK6WxohTIzYKFgddQLPNwOHDnPtP4FRxaVyesKZa5E9OR49NF
smPlsV4SEiGZn8Zs52sgJhjPrHnDA+ak3+LUyP4nf60+PMRT24n/JCnp8HKzD4dxZ3+a0s82vO6B
+OXqLoTKgo3l65NvzriGQOieHe4DwVBIJJ4cNfqj1ky1fBuwoRBhGwzoJbNY3x07Pbdfx4YMP9vd
pDnX4fq0dG9PwaWJm3UaghO2DuqGAWFEHfGLd72+iS7NiM+DMbjgsCffqhuN+fB6k1ZaUQQ0bAY9
EIugB7JOnflCpWXzK+Nq4LE1KERx4xQ1i54AydXCR/SpRLtDN6HIdadKMZxr4rZmd5bxqK8U6O1+
J3mW6I5CPaOVMl6WuenXkvuAswQMl+MGM3tEBghgDdH9Si5dAeqlpxfaw5pqvlYmn/YXve6wM76W
Y2+DTNDQ5/HbJMqUHxaaBpBwfrKLxG2lr+7+2Q2cfN4ohomEVuFRMROAhp4S4N76oTeSxi+IEVQJ
L8Mc8r3Ps+TTCwfstotD4aO0hXUNwtteeVwvkWQfTBlZXn1RH8PeMbxGFLnEeREV41KRvKT0nzaS
aro0gGVcvQ5a4aOGxuwGEdiAVB5FHi91wy/5QGj2DD7zN0klWXyCr+yDaxiasrC5K52rGnkOrgd4
LnF9JHTgd+2Y01WnUW+kz+4Ud29cE75rW5TrWZOXSStJav0XjIg8KYzb+9xQ08vl2cPSLpqhbbwb
3Iy0BRzjISyns6y+x/ef0jkPdza7wi0h4y22ibdf8oxtukJ6aQivkgPS+XyLyvx7SsCZVN4U6mSB
V+KHSTJOmGgUoggB0frrcALVQwdc7zvuK+xnLyUsIa8TYOz1zqZ74VREcVGLhfwqvlh5kkUz+944
RjYbXzjd5biA3Eo+lVgcvq4BZNAXWDhHh1awbH9OC4FrKVLCUXCN0QtUpGqD38r7eZNuVzicMVS2
H6MzmPadoxISIdr+v9Q4ihTglbMTw7PaAOGRDaDZ90nPttOiKyuEkmlNblvBxYsKAXHWZyPyFzEl
OFkuz7PBAM6TcV76N6N/rMGEHvv9SGX8woq2AEdbrw4ac3Yq6whmRfL5AsVEgbgbHA827sA3NHUi
DZK6Gvf+ILYPoEEV1QukAKXrqZs6rxV7hPiHRknER+wWh8OcX/+j1uuSwq60Nvrc64hsBjKRSP2+
5294XxetHxt0EAE+U167Y6H/s2MsX3O8m5ez2rvJdFmNENkSLEof54wPx61Svh6WcnXMQAJwSqRE
Q6YOEM+zGCzp/HgTakgh7u2Vu5bzQ6oHFY/QMztGMzOfScY/Z+G8HpPB4CTJV317ghLxcmBhkNv7
B2TKHlFothYMVIAs7jwJQUD8lpMlb8/qx4cDikMgv0pTsnHyHRIUpyRMf8yGhsADZi+5TlnstTZx
ZAn0WkgL0uCQpsSgHcod9Zy4WFJ071+Y9ORZIgHJVeWr4yoUE3bISsHH1zA7H/FLjmv86kK0lGsO
PTl5CkkIxygMSv149qvum5oaEdAxuVMRHw+VGszP4T2rPHVTgebTnLSiMg0ngn2uL2vI9K9vYezp
DUDI8nIYzUVxykwoxHjS/1yLWpGhRrGM8gos8e3p3s2lLBWl/JofASuSQzNEuLUlmHH/kHsohtbo
HHwb/dn5N9MQCpnj5dqxuWXtGKRlrchNz849CN/Uu6FXRiHk8S5qsg3+k8U8m6BjjTdmd9NhhxGL
YFVMSKN0M9fE6iviA8WGfiDYrX88E8oj59ihlaXc4W3dSHhHPn0OXkGBe2URXV0TCvOj5lCYNLnw
uwiteoesJ2lxGTa+hQSZQ2dcLzDszzcfqmqYWyPjgOPMNpdM2z1qLpoMdKNP0p3yOhXYin/fV+RY
KYZwUFGCMrw4PK9mH2omkTVqFIKMtyDzXshhu/TIdZNwgi1x+427J/FdZvte8kLQbPn16Y/R16+j
oyE+mWIxkx5gHyIsI2wjXvO/5gDX+OHIRoA0/WYp3bA5C6Oigg0mChRPo189f3r0E0ePfQsY8DxZ
1M1nUzUowIT5LC2ukoutPHepc+L4Pj3IZyXErUGaSD7dJj+GiM0qJJRdDSz57lAx0fEG6oa3bB7V
oQsKqV1Ivini0TsX0rRaHiNR/LqJmvmQqNH2x+Y6NVlIc59XPPFbHRvC9GSUc+Q4MtGcn68zUNB2
3IZCnnuXQX+lFnGUs2NKaqF2j7ISq3mIUlqBPv211OyBx1PmtA3mHgW2j9OxkFmcSEEjPde87Zg6
fr9tph45BjE7fpKETHzqAFI8P5HiGkhWCDrCJAp6+AbifxYMulYGGTK74EoOg5zOny6IObKYQExy
H9UPpXYtuoeKhWvNe45AttCf8biOsLp0muwuMK+xnsW+LdqRZ16+eqNXyzv91zYYVZTwhb29E9Rx
GNNrXX+VtTyOywi6A6WpTiwPrkKfTHBYX/i5dErrN9/tvQcuJaz2+HYMuix6Dq2k7RP3L5ak3r3z
8ofxTXb9RykYV4zGFIlHDri0sn263Z5gX7C1Y9ToLth+GNdTDY8sLCwPwxDVNMoBKgRKbJ2k43dy
+LFSwQdjXfACruZBz7l4/48uWfYhp+i5MAxlV8VINqk5zyWzp4OPpm+aAg3/khSrWzT/aLKN9Ebu
I/p8GNceQVZjn1tn2fFtt4cpGC4sBVvMNaAjSGSaY0UjP2ixXO8yeOsUnUF6wcUZoC0jYJMs+yt7
G1P/kP0Ql+UFHz5V5uFe7198/QeRpsEfg/wT4e9N59Nerge1m8n9Zs4qxajTWlXSuB3khxaBlXtE
+0Kl1pOnv3nJgKkCP7s1de0Y2rTaxaANRc2XZwkad5j8BUetPfb8m3w8jIgwmlZ/LGH2M3jk5gct
72bRgovWEGiQLPOIpV7C1+vtstq6IOBj6dWRkxtW/SHBS0r96M7ZdxIZ+sbYCUXi03A2B+kApYbZ
XP0VylG8NpZy+xh79RPdtDibwG4PmJv/SOyihDFg7E27oRUuBtYB5xKlnybQY+aKdizwCe0+zCiz
Q5NpW9fkgxaqheuEvKKUX6LdmKRuEquu4YDB5ONhT14Hek6mwvp2Z3LvKLLTIzAyVJN1eipMOnfq
AGA8svnxJLI+l26dMF4d9e16yLCkjJI9HGbGSixERmnLh8Bk2NHqg5PGaRbtCBYn0DUh8tj1O7Bs
7jlpMPe+ltaUnam1hNyDgZcP+3/SKOylAltBwIskDOw7ApCX1YkH54iXUQX8tbFjtWE5N3g3D6Hu
S1zNZVgxJzSnZFDPut5P9arKfiNh0tapttVnsbSftdnvDGqyb0GHFUiISZ9CqGJm8BS11ucZCSz7
JJk+Sopqo1DmhXFb+F6+IRmaYJfyQqId6c/jIHlc+6NJ66sNwQlY9Sd9vOq9ymRCpBgdftZ4Vwp1
miJ7pvGYttlGtgnIR7Ck3fmqQ/ssW5Hoxytkyyj9uLLn2xBodhiYUWA2vuRq1eptQ/ohdSdKIshX
g2BvLGvYu5Xo9lVbYgODduOg080cpciGe3+8aPPTXEiTrN8yRrBlPtUsRiAcFKy4QM/TIHFpFJuP
FuZ35jiYIj1pi63tKQS9IAVSlgaZdreNEF90cLSFYd9HF5/KuT/ia7xp1QZ8WidHmq3ywKxYOQu0
iWaAHlGDGBjOEBVlY/qoCFPbNLrtUTDup5zT7Bf7Z3VYRHRbBnYYzPpGRM4UrUf2kpyRKAe5bQv7
LIgazuubR3Bz+DJVFfPyA3f/+MA8Zixa/lE6rbYYwRfN80yb9ozsgvjt7LGj8PxDB0banLv4B6zA
8qdRZTrqexTRlAeRJp1KvaP7FegV5wdychyHn0wbaK1IlI9OYXEKcIKARwoXK4SxcGcH/BHUQp1Y
fHna5nZtcxlEJvnnFZg+ChrGDljla2E+KziMtzmbMrDL5yvr+FLLGogrh7xOfryFkYE4yKPUHxCe
Lk6xkES2bZmQ4bV6rI2QgFwMEDQOOvt5rNmFjwgd0dNjmq3W+Cv1eueoCmDDimsHPBi9LCvxdwT3
/4fXuarFn348S7lf9JN9tQG426XFvg0g3kYd4JPOj7GbLZbdp/i9yTwFRTluji1XVqdmgiQCvcm0
qd8y1y/2CqaYX+RGwpuSA2CFwSK63qsmTzUvTKngCOkpjNlCFNfDPceFpfgQTaBx2j+S4MN0oM2p
8jwr1zOEPt3pjzBNKilcNPji4fLne4sWiHduvxW9/z5HH9xjHonw0JM+5axS0+Bvg2bum9jDYwJG
wRZtcDO/+CZRtDy2HAdhnZFpeCW1kXQ2kmgrDGR8gT4FmBcSwTe93bj69BprozbBsjpoyIUfx7qa
9UQ5X8aOl+e61jcPmMZ1tvn7WOKsE4/A1nM+2k9dH+SEybQd0gekpfoXbOY4Uo1UYg63K82UvrEP
IwSYiI5n77DaYLBIb4SlE+zTPC9JFS6eH83qhefcoqtkzdOlZb9bC2AKZIjq5MtyJeYgdFbr7l5R
z1GRtI2Noi7/LkTzNhZeMkGGLKx0hU+a+eY96dCh7XnY1iKwaA278s2YZ+hMfMmi4Z6sWhamE10b
3/GtpZADumQDlOwff+rLLcKfd2u8Efp7rRQh7ky8RpS+89k9ZI+XY/jDX8D+/1DK471ESfPuVifu
NA4sleB7+10XnZ7vSmytqRH9IHmMTYTL1Ta1/x14qsEam+uhFrsFZ8sBJW9Fee18suFIhMVyMuUO
RwNNX6a3t0tfu4UG5bDh3CYi8xuVNAgPJW3TFXvfmc3katiMoZByepEuVCwEUm4WDd041Tr7U7LX
LO9EMWcgiWiu8YR4G7tezOHxGW/2bzNOhKJIMFfPj1LV55V4V1KGTq4Cyio3LcExaksiCYhvvZAD
NZAcUuIc8oonre3hfiZbogz0cnCwTLn2vstf7p5ov57RyReKtRC8j78kWEqBPuc4+ZFUmYh7PbAi
CVj0xWvjLq/LpR9LKxCxYa8vBWPi5WckbmFmFE+7EerdwBHlz3yc1MrDM2LUcfY76KK9NcIsZwdM
F+prPi+RGdmReFUgXThJx2iQwDL/3J3Z9NKoLD5uQIP5g/2hLZO4x9ILUzHkI8xLHgk/w7wGVZGL
HnaLiJ2RiWbUfN+604h4SASBuMhsS/548rc5H86ucEX8T02RcTQHGEuECmFJ4zlyuTm1TRYQjyaL
hjPaNXQkDIod0g+WHXvQx61rRHZVD8xUwtdvi1vtvn6E/ErfvmXEemfW4OCytZyB7a1yvE3Q5k6M
FA/Gnlw6M43mfIanT2/60UzYghVRKbVJ9k6XNoXZ1aV/AhpRPQQFuEXYaojoXBTXvxp2BLel4hIo
PK1hm83F5YJJNChaS3UsGPkgWCGDaympHVtJigsdGWgEwEsV6QB9UIHJna+iIVDwg8/oiyN1u0IS
0IMFl79ej+ARlS4Bo+LJyi1keeCLj2RqlY0PNpFuWDJR4qcwr4RhOK5cE27Z2VQ+1TUGXXKmHCAh
2aUHnBRVM+3nldFi8ZSLSPDr1UPI55lpU/84rk1PVlH4FpmsA9/zEBfcd++lNqnJ/DPFv59JvY1c
vdNHwpywxQLg35q/ZD/QaOqkiUfwXytOtIa9xg3simG7TdtgCQ5Rgn9MMRiZFCnfAHFRX/Vz9NMb
egFmj4ry/a79TaThmoHJ2x2aaf8E//7m6rLLFbbYZWgJHeU5yILcZfpdDdSXo0rqCrjb9DQm1gZx
sYYu3FZGSpipO1Po1sCdh+Nb7Ap6XLQQGq6wpF77klhZ4VqDu/HbWN2W79YGp97sDQ++GZsHBuhu
W+NIPHfQcz0RmMsjfruf3NmeQLaFIZYqr6e7i7j2w2+JO/7+rNhlfolJDXfQBlmh/0dfRl4UegkU
gz7Xmb0CuHaRERT8YZ1HuOR6+h8psEJbF35MS+FmH4PAfHRUPDtqFi9u7EROIVQ9goCpZEIccXn1
xJVdo/t+mjW8ew+lOq5vw4uq9stQ24vKfgV7LlQqU+Vl4TQJgbY+bqa04txTwu6hXjm5sUm58gt2
13L5U3Mbjd+mJLy9fLrUR0DrAa3sOZvzSKJ++jFKlHrUBItdf3AmzTyoYmc4JEw5apvFTktqtL4O
U0ibFxVOIZ+lACDI+PPffb7a63cyg/r/1ALsu8U6UkquEOSKTpjQ40kZ5aCbXoRREuQP2Zz+SQwc
JrpqNZYzQUFAEBQXY0hN06Tvna2qAkyZH7tHrZRJqOnBUfinmY55XWnT8xVVk1gtRj5xJAPY+6wJ
4pGGFt5Fuj4HVg632+RDCBMYi3oz/dlTwRWGtWzNunPLfzxZYxmhKy92Lj5NoXfDSU2Tdf/0W9E+
AjznxkwWHi2ucS3bc46sTWM7YAKHfzhu1iwexvIBcPxapc3lWyJqXfA2U8T3XTPjKimpjgzKymXd
cXfrUCGC4fOWKfphlYU+LRVdG7cvE8p0cJTrcVluKvQz4BNO+vkhkwwWzVm/EC6nSZ07wXPEttL5
JDq0EKSpSLKKX/ylhuJwOC+Qt6W72Mg+918AfVfD6MM4MANYrLctCN5KnaARDwJyowxx5TOLcV7w
ssnTqzp1IRJRU1l1ZHDGpzaCSs3dkyEvG9sSGaP+VV5DORmdlSQJsqZw46Ag4Eol+XSgVri+M+OU
IgMuw2nuHIBsOgw+0+8hUFZqk2SOJj9XRXLsMMnwyZHjuFt8fEvTAxQAwrzI/pUDE8Rn56N3Vjq9
NT8wNsJO8YgLahN4XyFfuvhRVf8iNVfhbYPUBVu8u92i2sFsjLuIzQJHZqQrI+V0O51oK0/F69bq
TZRNoKdJqi4WxflLppPjaxrow8LZ2eDwoXxAa+ikoYshuv3On7P3XYi/8gpkbM7mfntU1sjm7OVv
pfwbWouCRLiWVXX4yQozUk7Mx1Yppo4psMv8A8tbXGKbB90TxaCS9dHfkFwSQIntzlEqQF/2HEcF
iLaKt2w6EyygKCcuIUkdQCJlBE/+025mSeusc8qI6N9/UkOxhdRMqCHyMeC1xBGE4n56YP7wxDyD
4JcVpR50En2aVYW/gc+jTSS8nNUnCDJNVHy4GKfGe25CLDUr5aYQ1KBOJIes3IcHjoA9Fy1Q61LL
CUXYlphH9vmJneeu1w06AbgM7YU4Sjtf3qtVywJF2Zf18YenlA7n9zD51pFTXMWIbvNS85b4M1XC
EaVPOM4hLwkT1nYxy4Ok5+Aau+AWxdkrmg1ShAyDFWR2Iw+86WL6aZMIUDM0Stn6iakaRG/6MIIe
Z2mvIfF62az/QtXUCASWl/Mc9iV7CLKEjeKFfL2OvByNDF/yLoBwxGCk35wW5P5tMHFKfGAuyaUw
zGU3q+5vEi1laTRO/RW7fqzKVMZFBcML2ADiOT2sThvY2nvWHzQpjb1LyVnFRgNkg6OKKA6Nxah2
KjCAmSZROmrnbz2pgQfY5trweo7hEsFyh4Oe1hrEZIAf0L3FkHHqXx+h7CkDasyZuGDTZg4ymyav
0a7dtsxUU1az5JYHinyGRjpXLWwIWNkEayMsu4ncFOMcdqTGd0PiZZ7mxJ/i1VOwnjoopwkL7Wv6
mS7J4KkpRNUga0g6/OdWx/kHIplUjzIZnQfNPC71uNSjepxreTPkPcXmA169YIoPzViEdiewS0VX
pL2LlfsjqIQYydpGLCiBibhJV0ttCsJ9iLEwmP7viA9I4pKameUwiLCyW98mWLOwT0W1WGy/kGhV
1iuFj6WzWZwzxqwIW//nkkwlTIsYsN1AoKRMDtED/9qsLFPAxeO0/XfYURLWOSs/yvSnd/UcAU5/
fgHhTrgxzrqXtJniFvcHxMi8djCckNd4ahf+jtYRlxDu73SM1++NaUYaOO6QePsOdDHQG1VmacNn
yVI6ro1FDDSvBXNGb3UFQ155Urc94WTlfhULbmbXeImFUuJxt+EUuIvnJ54Gz8oJFjHT67Rti8G0
SPnqdkjvO3HAHIjr7FL50pDyoCZ12Z+pYr2NROK+TTBvnYkJpmzlP1mQb1fQGDIoKaaTL9Zags9v
ndPMAJO5UUndAzSLMlGuEsba5akO7RlTauKGLwbvsy11II9JOi9vZtp2ff3d6sr7T1UY8Xc5/xyW
TpdQUKs51Da57tZOxLrjRexyIIzH5oNOaOzb3Xw/tsaZy1+Doc8sApEMdjCn98RiCAxOnuqSc/mR
QYUGbtVAwXOqeprLBmyYxdVlryeUVzWrCs7R5rofahvWQqcV55Sz+l53SEYoNOKYmpK1VqE+nPcf
vJmEolryXemGlEEXBgvnFWavs9E2HICazkNIyqbbn+aWKM397a5rPUAUG1RAvOo0QeswGGhzTyEC
RYJPpGo3vmAD7Kqcn/PBHsA9AprdLQ6H8kOVXpqX7N3xbnFDWuKdpT/qjWlWdPAKJmtNk/eaIDVB
45QBxmmSEk/U8lXaDBjvAtyBT5TrrWtEzZEt3y4lT/KlyleHpvv8w5/IdNcYJv8vPrZ6gi80Z4gJ
ieg5S62O3Q2fPBSh9ifoIcNUq+W+Rxt3gvY++1cCZeA1aWzUOOMvi1GYJHaRfXOWXCzHRuklikU6
XvmKBxyoeOtXRzloN5X0kWpBtiFpoLesH83STn0BIssSO2PuD0/4ieWFEPVekwzPfLijvc+dYsv/
Zz8pelMX/AAb9cgKMK6kAuBLPLN7Dh18muWTxp5+DLVKejWFrHTEARjjzOi9yS+oNmAQuleTgQJv
XIMXK4hjIKhssouOJULQo7uLdqIPTD7KXkUN1oCZS7+OqgD2ZhyB2mjIQxhU301Q5ePL8Qj2nlIG
DuAdUTC1+rH1nRSRHun9iUf0V2U3wAXIXMGjunvl0LDh9Q6MD0r4eGGsgI9zHPvy1aN5Qj9Ko1lG
Z/AjdC5FrZu2OeBVoHiSqfkeJuEAAiamiPEePZkch++YpBghFaBndACZ/o6hSK0e0cOrGU/VTz4g
63CamMr/MXkUbqW4F0j3VFbnhOEmVdcwj8LfAfhGtrtAOuwaD6cs8WQrNnzi46I+N+nmbKI3mx+X
v0MpY6nfeqdgC6lYISD9RcmGlg22RsyK5+bUpeSp7+7vHzndsV1J/g66E9Wxok3Zw3JYjep7V9mp
WjAYVfqU51vOT9icJcnlExvBb2fCqEVrwpwVFO26NMgBMdmYrMZ+S1saP/J+Htf59pqWSbSGQnHu
cNB11w0h8LAE7MhX5z4FO9LZnCLbWZjuOcJMVVKr+pHO5YUFMbC95C+mI53X5Nl1D00bWeu6GRMJ
UHrM0CIIQ80Oj2f4HlqSzjXjfZ4+l2Wj35+zNQEApsoBHNB6g1a7CfBqHJpeV9lGnU447WNnv+Rr
+QCLQpz2mHJkOqnNju6+g/THxxYB999Wfe9jy4cxd98HiG3Uz1whaEBbJHfuwfeBYg5G+jtnSEGo
2qyElYqq5yArcW8U60juNTDHFnTt6zWIjMgnzo8OVv8rYkygD+WoHE7ooKtyEoeZIx23hZFIjUML
me7JSMRS0d9DL9SFY48UAvNpK7w5VHYv3faO9sdXhppS7egcw2Vcm/V8MniBF9DzE9r1a/D2OGSN
dWKQqgDzZaqEMGQg2ooabh+hJM7qzhAbiuieKfVmr1j2bQZwtqYonPe9/AJcs2wILG8uX/JGt1AN
4EZDkxPQ2B3lMZBntqp4V+1JzZhjR3lnunGY5N8hQX06WfQFTExkjqZRzxI9UfpjIqOiipHm36OW
e+gH4ektNws8a2KmLZH/Hi2ynde/aoxgFRAIhWNjGhbrdzF16OanRGLXrr8H166hXmdSkllEa4lV
XX7cnepVy1a1gm6xx6dApn844NYq7qtBnUe63m2KAbB68rJv81l3NX2b7gs2DGBafOtNMyjGFLn2
uCeVuyXniJHtjs9x7v7YmKADAO4T4PRQ0mel1dZ2NIhUFfzPtZs1FKAnPPohhxymYlpb68j4/Ojl
KYoCMc0htOpex7r1UnRl2WocrQjT6SRu1hwMx+M5p1zDyOr79qNWANK2IAApDYQ79EcWBmPz7uCA
47EYBadSS7O+uP7kWqg9pfl2LG5AFrnajsllcvPkrZtCgj86WnrgSzxRucA721nBHj7/GqCKzaSW
foXpjaX2sNksSTQi0adlHnRTJbEaB1SXXzRHxUt4hh8ll9kQ2cs05iaTBbvcDuainEch+36N/Cqc
wEn3i7keTwXrkT8W3cQFXxhtngd/vnaPpbsiiN/K1S15gdZ+ISb5BX0uxXXT0uv9EQ7GtZ3Sbkre
W7E5zMd9YWRnp8etcMfAzdcRoWrlkaWzI9f0aMj+HwA7KcgL6sAplID+ouQlQ+ZifzSmJc6PbNok
czkCCHCuJ+Wo1Qv1vDgHRUm9G3976O1EJ/Na86EVRd08NgPlIYZS4e6SJRj7jIaGxTRka8zTguv0
5ivLq9JjPtY0IMIfJhvdRSbfTcHojnMj5II2T4y0JkuikCr57gOjuiioJvOKAyx4PjO+MMa7OuAX
3S7jrr31FPRGLarY6DXOtA5zN84delNCF5xA6yBUKUQLt05Lucy9tzYn/v+FNxEJJxM875Er8rpF
GDo/ExUV/v6+piTceXoZAHZ3EDY0FZ5XWZDzMlPSxamu7nsCxMfzEkTsI4bi4Q3RfMOg/dhaTG8x
h/DVyGDbWJzuUZeZC70YstahFNTkxxudvrfsTX0UuzHlXOhYwmh0oRMgxC7Bw1VoTpHhMAWXdW4H
8hxS8tu6xL6r3aw1twfiP/blo02urtb8x8/QPFgXOMDX7RbYXAZyhre4EvIvI+ME4dmH43BsHn1G
puJH9woe8dQ/AfN/rwEg/oQC2dTZ8j4MkHucbWLUTIxL0V7ylFBLXB5NZ5qf3QaTFJO4y9i5af40
R343zuVVdCqAkxWfhpL6pnmsncMv89p2DHs3xQAsjeQJnHfI46v287hIloDRb5HP5yacqPVWb1Si
BfUvfrPofRkFRAeFYeRog1wfks6ezh6HO6tgusUor2Ff6qCCKLhYQPaoKsEhA5oOrJ4KNk9ZC9/a
BCXN47cE9A3sAh4VVn8Q1Y1vONffQEJLawO+Lf3iYsgEGHL5QASEhFO3Jhow1VSN/UFhuO2YRns8
vckzIi2nFNOmXiNRW3DmGeg1TU1jwqaaZMmZ+DuRooODtdX1jHyRbfBhIOpBhUqeKhcS75XWF6qV
/UmmhtYw70vCyfsEp6dnBEIIVn8Zm5/tQmYMje5lKK6eszRylG3XHuoaj7k2sxpN0rzAKDj6ItgY
PlGgfiVuMgjKMkG2QTiMwRjxdU9gplXkluzw6+Dp1odmTEUcu1P6EPzrUkzIVaUuU55asTyQhOip
3w2vdd0OPOhhxbVZb+Ojc2gJpw6+WQWb8uwhILNhgDBOnA+vElpjvExPlXgliSI4LDCh9qzXpSdO
arzmI+7H2sb9QboSS3AUjaMcW5qe8+8GStXR88W92QbCZ9ejBB2tz3pwTsLdSOqwZPlV0m2SSYal
UMeZof423dcjBZGq9WVgR7ghPtESS7+9KQgeJeh680K0UVZuWBSPjH7fvlMfdok8lhAKZUCbDAW0
JLFiv9u9M0NFFht/YJkTMjvoIfUlsuHTvWjJZFzo1LnQSOEdZAhycsmnQmO4GEshFvxML4NmJJ7I
o1qsKgMGlgfUptUAP7j7cHknXa9bDhONE+bDkfEz1dQSwkUOKC4LIIEtoTI4z0SJwC4w5P2lGk+s
gCqClnqWfI1HQIoMaJD4ptBhjv216lwZj8HK3rLNNmOsOIiGUoim8INk+84ieRPNXd502CCiWU33
iUnfhbnYVEQxp647zD9Mb5jonUHeOQQ3n3Cp13I+d5q6J9p9GHc+YSvFfyTjreT6/dsea6Uetkz2
KPZGMdOiMeKzW9Pr3GgsPNXMhLEaxc3jgL99sSdzBJ/zVZ2v2o9sMxIVtNy7AU6lrzcVvXy0qbpn
WlX2GY3IFO1cST9SqWCGSYeucryefMeNr9ubWTnen4eSdisK/TEOMKNNXv7wtwpbwURZGhlwjE9U
nv0UFOwv9XXGZZ+D6qNTRItPhhwUgfp7P77LUNNFKFV/wkQIl3SsIB3WGJhKnzf8lHeaj047ia9Y
zMnoTlZ+4g3z7EpPWfiX+GdH0dgv5AYIx2TkK6smlFucwuHNF+/viMaXYRTo+CTjYg6gbpE9mHxe
sTU9U4BszRUtsKUQidjRCj2a45F536+uzZ2CXDQba/FHNjtbXSgcRjozQibwdSCvPOQBxFR+GdVK
B+y07RtQen+YXiPNrU73lZzCvwTsSAxkvTZJe6NdcnKlYDxDbJKyJdF9UWEtN/sSiLjj9F92mCPJ
jYBTR3Oc+DgoisGNHO4dA5dO8vAJbuB78Pub8iCMM6d8GjXZjTkM2J9AvGY6LN32VAR/WSsXTv9w
20jxqg/8iV5Vhdyp4/ToZDAhKrcB0mzQbYGA0YEmbiuDZeygl/V0+mShwKeiQkxvszlPqWS6eR+X
JkPeQhi31ahQMgfxtwi1eWFmkt1De1nsbp4yH49+lYXI1K573XdDxcDp8qjOLeifAiHoeuwEtTtn
KF4/EHHYlGKoJtvlIszluhIkPG4WpTip8d2eW/U+PVIIZm4hUpAIz374w9K+gHCgExler80fRfYF
u1ZCNOfayIxQRBN32J6sfFlpTUJ9vcDk31PwLCpAB/q4C0fQCTksNoQFauV5H5Slk0XVqddwlUve
9DU3AD0MvTffszNwbAUk9NjuPj8Yu8qG4rTmdH/9ZmPnmjJSUjAOoI44OTzURrJRtAjBXGSTYXFJ
o1Q2RQYS0Dts80gFW6yoZWogfB4WrLarGZ633FoTlMQFRnjN0cM/gjGo5E2TdF35sK7D5a2pwoIw
CWyZfjkbo3nkcGLF4IRt3bO9PEh2ds88IEdIptccRTe6bKVFOWjuEFG9pLxVcqTnKGurpejzlzsn
UMpNLZFpf8je95Rj90UhRNXy5XCzJPf4oUXnjoXEqf1zpAr1lcz5p+/hLVz5tUiJBxXmbz9fy0Zu
vKI0FRf1OcJi87APCDzIzMY1z8VnvgTYorTxESgo4N1K2h5ivvYHHUQVSy/sBZU6b4fFmrVVXaGt
ouyihK55K+Jcxc0AWlMkUJYSSyMZrqfnr6T9WmWebTrRnfqcH9e84WWxVjbTHwXcOR3Zf5gFpXEj
kX0lV2OhD25wxzLRU9207u5ZIwaztBGpLxF6w80vW/K69xtLblmpYru/QN/QFETGpyMKRZ/ZTEQP
o5j+aO2oCQno40v2Kvie9HCvWjO57jFsloCIACWlj0TeLJUND2LXUKWjczR/KmwpjjNkbrszcOTa
GBdWwnVvzBWXh7stt2LI0V8iiZ/6/aaBFZRofIXnwvBSg8ke8iBiN1fHFT+ukk3KJPVIFdacsiTE
fd80fiT/ZJZgwjhYFpwI0ZRdoovbyThg7tma3cDXWRHczhtORqwkEnxsJUw+3YlBlrQ8TdDA/yXI
7H8wGKrp7VHyelC7PFIA3vMuGfpSy6OIaKcJY097cOcTFPoXo7WDQ49ulpdJuMcGmfz9CH7u9ZRX
BcDbipu+RbjEC3yGnDrOM0/IwdNXM/4M4Fkl5KKSIYEpdtgFuzhQ+DtqQmZlk9vT80WoRtIWQF5P
WwN3hDiU/AC7MyknOm2Lnkl7xo+iGOGZXJMH4GDEACh0Ai0FmRALyvoPlVTtvTgKwM4NjGS1acY8
BZjZbo+lTB88OIr6d4B9+asa7XkosTGoplajopeNJDMe9ugtYQ1EGjukA/vpNCpYHMuGEvu1+wWk
cgaWzsT1faB7h4Y5sMyFydmOVHalvqPSjuiq/oZp6IJW9KwcfEeYBg9LiFEcOYgZKtJcze3OqDFH
i1HUvJURfNDJ+a7ZdjbgHZCncfHBBs1GEyft82pS16fuhySBtX+qUnibtzCyGNxkofltY8cEVkWN
M5Uy+mumMIsxooumZEvY/czmtS9MOHnwvwCDYz1Cc9T7v5D4Z2i3K9qbhNszafpesNg8RVYNi8TY
fMWN7gcBd5cpYL62wZhgfjsaqzc0d9UApgvAjSGqrZwhrakaN/9KyCiSQBJJUpJF/TZPdj+DxRMP
TAwdo+GMxphRmMHwfonuZcNRMuaWFEV2GSNV3YHbxDJAi9ydHUcYIhTB8WIz7jVIdVGCthUBGzvh
rB/HEGNJfJGyKmzo+0zHtPyeNEtVWoDiB43yaukiXlL6euzGblmaooXrmdMBWzVsmpFr0IlWQJKb
DQx+vzD+oYtY+uVpQGdHjFPG/+ZFrKfoajohLjOA6d17/D8oXsPucDZVtQGF48I9EmUlDvKRFsQ0
7N4BE5J+tUssCwhEHtdJdwWZtw/lXMPpHAMn8jgqfT9tXg1XOSz9/jHRj+xH9neS3HNSkcXklfAy
ZoCdKK/3crPu6GqIPdhr5bX+Ok/+acHREVrZguOrtDbkiHDnQPTsBOjr+ub16sXUZ8CtSIzAO2Vk
HkiHx3px9otmROmEcFHdOaLcc6gzQVcSSl19EUaSke7/mWgsITsGus4+uBst08hhimu3Z8J6kZKD
LcivUwKO3G+fpvDEvDp31MZBWv//r8NKLzNjl7j2eNJm6cVn/1TSIuRdGUSNRibE2PWrN8tcoUk9
enaRIvcst93kR5Q1yqnGTLt5CYoedjBf0YFSuIfQpqatK/9v/rBwGp+sQQqZqC0nihLDMpzMQ+m/
tgYaCUeo/AaMk5T0thjRfYhLVb9foFQtu5ErZjhlWePkF4DSfyujOZKDFARRc3eE4alvV/beOLyw
ThlSl1FTJ1vpIzV/+rBjHYD/7xlvJUMG1pIq4JDB1v8pSG0FTmoooqBcvniGA0tVJW7kTWw610kJ
9096TJt3v6OdZ8xm7m3FdWyee135gZQQucm44Q588JtbCoCO8vbfQPjHnhSLUhhllNZgoJvtWyQP
QYiLP2O4HMt2xAxtORvavNiG3xf+B4HVz8gbYPZqMzgVYLVhZNVTzlElpS6xaGa17lLFlnstbQvy
c/AC9V3S8Itgbr0URVYAQxU/Ou2+qEUwpMcGfxnt8HUtvgmPFarshfyFJBpcDu0PhfM6euGKB8Sa
ygHdT2GCjCAcMf3KMwciZi3CvqgRPHqy03WR/k25EWxajrvqfEfgm8TknXwLmMj/tvhl565QNpyO
/LXJyE6/1TaXQwuplqkHFs4kkUL+EVta5vAuBGNPOp9kfOhNjUv/rQhE6AG/AI9/SoRKVuvzGt3n
ZLeEIgxObaUSEEdAt9ELF9XtyJYtdpNuBOpukUkaEDYdknJmJ/ZcpVvs7MSYLBKT+vhASeb9hayo
pX8NFYDp8F/4LDBlZjBNiyg47WHWVtgleQY3g7CpF5Vfxdh5EQ4Ube84Y7qB5x0VhcCgAlDzI7yE
66zFoXyx8o/M6OXh5fs6ftxK0MtUAyuCmYlFRr1QYwt5R+OoLooc6rTov8FPjsW4X0/ClIYgjLSq
5cZxzCfPkkUWPsTbFI1Abv/6MqWS1kIIX3OhFQI9GTCzNdCQPfBuPNHUqYHUXt20i+HjiDjdN+L0
ULLBfh3icF4x1ZOCRtlnFW+sDfVRRfWLi6VQGEw12hPr1Yq2YJIafdooe7WwteSySy5I2CoUNUHa
HaeRTUOYMz59BQuWacOOdQaFtj6cfevmI80zEGCUSBT1GZJZJ94GhDPwbASAkmgMu7eSsF5ghQIx
8BYMzG7xAeaKdqILOAvYtYImKQrHg1RUJvpv6e0dHhU/Ns6XUJL5Mv0VBF220F1bi19eN5tbUTmJ
OBcw09E9zPWrt8d+Qc6hrNV8ElTCFz8L4Hm+NQ10Zx+FNFuRwtXOY5CoLOj6Si8hKxPL4ySD+6q+
AKIBlbLnrLXGhREH0cDXCca/UM6kajzfBuq9rd2E+HokWuGqbiutVMO5aZDvDoYAqdX8ZnNJzXbT
e+4Ojxi16zekVbdeegP+qH8bPPcFJtQ+wjuRiB6WTfM7A3yb9CsX+eoU7FBh/39bIH2A0h7nwnOz
ONmqdyKcDnaSTWj0d8PK5ysnf3G7kuBqQ9zfZyQ40bVbZKlUxpkak2kgog8e3mTitKSocifoN8YH
+uP+W1ySk1Rm8XrpOXgBw6HrLMzncV1YDveuBtBgTpyoCvBkUZgqYUQlrKj8ghnyjXYWb/Jv+V8s
yO2ahAFOUZAs8E742OQgpq3cYhUwdhFs7BuJGgVAAHTTbi6B1O/QYliTCL7j6TTGNRP9/Gxqd13I
VgeV7QuU63l/uQe6W/SQcNIU6K/8rXxJNhtGN5YgbXS0UhifTYbA8VmMgIIg1LahXcHkMh/aRb3f
IhAxDMf4hA7nzQk0W4DWgcTUBwJY3wcvRoHBlxpqQM1NpiixXxS+d5Mx1yLoUe6ALqTXeEqc2zak
Tasa7yAOvYKM4F0wOvIs2NeLWV7Z47yBt4zSugUHOlXQARoNjuM1TSoTMGrMfBHODi/LqHQPFvP1
96P4WayZWzBANZ2X250SxvQZMQJbcJ+DpNxQ/NhEwWcgT+XfvVWSi+du8u+DwHKF8mpuGBkk6eRT
rlKZ09UFz7lldTr6+serWejV8Ynz4/tcqPd8MZn9de+sEhrt/kRj0ze2E3lV9wa+xxh8gbLJ8VAm
KmksmcNd1VXn8a7zYOlWfrThlZiR1cPs/tfcQ1Kqmh5dlOGPdOsTYkEJDaXB8FP69nzQPLy2w2nE
96poiDhLSnxVe2RFQx5rISsVwHfuQ4N9ep5kGWkStiFb15xuJ/VR82doXkazYsTrPVkT2ubUvrzM
bLKyogmIyB0EHUgHjMqGIc/EPzx2IOBNbnefCen/VhTRohg0v583wWW4ryKIrTHHP2mwlzPWj9Qr
AwAOe2iukyy+99rvWBPqMOvAoSX0CBwkge2lfU7S1jLeN2av8PmkvFL4GeVeiUz3CM5r4MuSazBU
aZ7nhT6SiWy6r9wwntKSqLBIzuXtVx1kjyBe48+P2tlqcn/khw0orCMD2nn2qLbhFKVCUjUMaOCx
0S9tUgsW2Dakmb5Mxbfro8HzJz+cIywEk/BY/n0WtyAmve6HGd0CI/4goEQNf8vyuaYx32nE58F5
9cBDc0aEVW9BlfzkJixmhexrEsuj83Kvtu8vglHu0pubpmZA7dbJAnb+tjCDUIhE+YaqzI/g38wO
OMAw8z/7fs9vQpdAcT6ySd46tCPnKFAvDotskIafhXOXQxiFFFMi7oq4nOOeXD5xeFx1xm/jwdkt
Ko+B+6hYh0E7vubpX3IY8A/nRH6XjMx9jJ5ETH4RFWZeQzjoeHA0Q61NFpalbC0CUtu3SWNyWCcg
7pLvhV62RVdFoEuUPLp+UILY8PT7Oro0jLQR2yB8ioSTTNif+kLY3xRTVapqmtW9r3iCPk2IHgjo
TLDMJI2bxIUacURFhW1vIF8BcNiCHx8/+a9vsMRPo6Ro4AJPLkOVbJw+OXel8HPznZKfzOJIyhjY
SdAFPwgoVSq4P9w5xVFv6MCiXVsDKBxWnyZPI18g9bLmvrNZ385rkSj8vHeaO7vEsDEo1IQjMzw/
PNOBsoRSvhgrY2Fjx6YjiBz133OfyB1avpPJfhE3VTGZytncq+ZXAW0TvZMJGyujiYQdQq4Qj1op
VtY+ReS5uzstkFfqoTa43Ai4RlhET4yeegihDMqTZmeYC3mcIXklo28RQuvkmDnGvXETJ4aqhVUc
lBx8dbBjMN8sp8O36APCOGLn4LsrsYAVKHTPlipNecm2HPHGuoISiJMa0jWcYmJjMR2J9aZhrGk5
bBMOviC3h9b6fnFkYlxlTY7DFObbejKZqMWpWXIiwt1FgWW11GMjsCemZDEBclGBZ060hXb6v7qX
7lCbNT4LLrs3BXSVZlsC5wIlRMx0lFCrfbxJOCZ8P38PuBtlGAkOZfj5oFImeGLcfMnvdWD03J8D
8Te6dG4OfVVG74Jc85xHnCVfWvUZ6P9DEISnQjdgLS2Fw90rR2N1ga/anopy0EBbFuWzBRyTntzw
V05t73Zdoqpp1Dkl/HqhoPTR3GSHpUFnHgsMlaPmHGbQrMI6Xf7faw9Ywl4MQaWbnnbmZhwqXIi1
4ZtTohMcvCphzKNtHPCDuSHm+n1A7UvTZTQQz+2EIQqljDXPHuenuOwLq48fLSXEq2Mv3QpUpdGe
v+8LSXLcQOeXJkNV/7mY/IhWHOpAdn9UZ4tXf+t+IL7OoAFqu5loDlnFRfaHCJl3mSEq3lFn3+Gl
a5lcrF2qln8hUcnv6K2baId9jne6tc/IQ5V+1dNmZ9waIfeO0K0UfbkklrEru+WR/RiuLaYeDkD7
ga2XuwbPNIpJ8cxLjyhSUqzst1ak7Wg4qSHalJ9+2BzbkL22hlPvbCvYqsq0O9F8oHFG0lgkFsEz
VWzQ7SDsarN/yfaUQQclzAJwAbyVjkBubz8O+CIqjvcJLbED5+l91fF8BXSHZf64gBcEE39W2lwx
OMDgjjMVG2zIJP1zTczRBGDA6qI62VsniR5Oc8HXnY9KpHE+T387NkqiToxqDL5s2/oETUsRTx1B
lEdQD/QPZpTgGCUVQZ2maErRuC++bp7Ui8qIhKeEljMY4eE3veZqsXJS+NeEewNwVkpVeIzLiMYZ
HwYAc6NF1RhSV86v8EkoB7ugnx5XzU+tulBrufxUs7cO7P83ZhMqWyrc3LGIceoiYu273qzwGiQK
WnoOKskuyGDDfUiXu4WOmgN5xSe8uw0UCRFl2RHwGOZixM7BBpJ9a/oOaoEiinm6v47EFlIpDPCa
Ian45pYg/nlNjzCzpzR7E4eKKmiLjyCmxl+IqQWxSu9pgiOjMWN23fbzSGgCeaYhvm+bVNy0T6RM
rnLyZyDHY7lJlEB9rnivU4bL53FHuLcraJkE4rOxG3SVTlA0oOToGA4Qx+hIytTqoJC1GfJ9ytjq
bjdCvv8IsWRxelcce9SY9NgyR1EJCEJIiWiOOBiiXKKDETOsA4wZSPerbpGTu43zD85u//b6ONQt
4nOJpv1yUGxVAKWhxeHrB44DeNStAESbr4AF4rrYBmxj108L+lNK/TDML8o7AA3nq25kxutlMQGc
0NyJtNkIvY+BL8EeY0yygATMnJguNXhq/sSBuccnij3Yk6ZSJ37e+FAXb2MfocfkbCzHZTkTtaU/
JWglERjIUfFGpmWn9uYKQlKjV9rLG3NEM8qH4kViZIImVGGkFhuvd65bALp8tnoo2sgAqb4yIVLR
BS7DjIDRO9/iM0ehWt2RVW6Cpk6uX/MQvQyFWlb1p0LxGGiok1fvdIjILXmjUKctXbqO++Eoiqxb
dMSVS4zm3xQac0k+JJwcW2FkdBKRe+e4UfRKREEtg0711FXZpmsaGzBQuv9blv8r++yuhh4IpAgP
f41bMfdMS7z6v6BUng5hqMOkhMvrHIACv4gRIyUKrhTXw8XhqCEGUIr2f2LXQVhnOMmgaSyooI6w
xDfOdEChmBQ2AkRNafgDk4w/TvyeQBi2DsYdDJDGrBVm9Qnr6eq18WtJ8eNTIvcTnJnzvlfJQx9r
FMRtXMu5eHB0Ct0K9IKpdlXpHy/WuVX41NI3hk2ZdC69DEszgtiCnlXCsPyPchOkVt47eUMSoof7
NI0DVt/eVeX6+zeQbRcKzMv5HTfMMIh1h2fUepyYok/7cWulFdAf/7rfthWEjpUp9YSzm5oMB3xj
fexPoxc1MTfQaAQrMdsTw5uHW5wWzlp80TrCCC5hbzhbU45qYlbcpfceslrKKTjaddrnGmYzihte
/EBt2PIPzIJ78U5IALCq71kfGHLaMJS961YWGPMfaZ28X1qyo1g77a2R13ncEECMICL2pT39eYpB
gQPab9Xl1XqCcmkUHDAKDfV3aailkZSHxvocOOLl7ndq1d6i3wtrnKEmXADQZDzuzMYs5A6Z1aPj
2m7dLkrSFkE0WzwADfT0SX77wTB3RZgt4sODgwL5JkthWiJfBqyS1L9bbIkGXOeM1SuBwjDZpmgO
77+gUmWbjTz8pInSXXNN5dCiJSw80g1eUxMWXPUv2awcyQC3g/nyakWEXgTfUyDHx258JjCSer8s
eZe/WjEuLVdmodK+VlETtV4vfVMaY1nCC6cvC4RN22pLrUX1QwwajFONUaBCJfkZXM5X1fNeH8if
eWWYIz1j756C+bTuXowHc/LVBlTJPY3VnP4OGvo3MIyRC1kBSgi5UFKkOzORVIJyS3TRSq4jv+sg
iiaEdchpUkdHXIgoT4qDg6VZCV6QYmpug5/pxRSpKrB7jKVrOj/xlr1iiocsb8U7EfzAKHBiEv7s
wiKomPgmxz02cpwzD0ENNcbxQdFCWul3cKv2mTFUdEFYd59fZjQJ05ZhtJX66qzHovNto5gv2vXJ
OWxL3Z1ETE4cZBksmliU9q4X2msyzqh+2Vh2ISZs8nBpWUxUkh1oKwytjVFHPyW2eRq9Fto2PbPV
WjMOlYVpcPHO1YwDTVgWGK8GBJo/3dNAM5zJeCrcNCj9CGUMqvV5DwubbhYOUu1e7edrcsSq2x/+
jTBEax0tF/hXiZ12zaTbChehg/kV6Iqhm0QsHDag+IQ845bWyw6530JDT073gRSn52MCBohkpZ82
v9KxlgmgGln9bQkvsUjnesIj6Efw9adY2EUlr71eg57nXKU1p/PTYvW1xn1CzOmqEQum5Qawg+hx
hkELPK1ZSuEsaKql+FwnSVIN4QLPBWlK1G2vSiTMGmIW3s/EUR6G2z6K272Rx8O/gJFu8Rz/x13z
u9POxNWmapH26re0EYxNXp9h+ZvgMTHZIvhF5N0SHZVz+ikEwXipJV+oBF9j59oUnJO4WL+KuEeQ
vqZdXNapv99k2S94KfqkGSi+s8ucTvzuyJlEpSd60Peht/bO3rTaA0at3yrvbtAnNqftsXapldXd
sBzHFFU7URERER/TVE9sPUu6AoO/VcYoH4yvrJ2vSmKPsoIGleoPNbpUgwQXCdWoCtUaannv1mJ7
fC64uaFxWvOgRtNiNNTmL/hKHr9eYESZT3Na0fa2DhTBbbB9oPxoqjprnKOSQ7lzzME9+GJYRtoj
85+L4S2Rnb0afQzKftOAIsYL7QWekmo05ju/1BPEFGOXxpVyFOGXUaNQrrFCx1CIF/y+hf3VPR7R
5RuRfQEs6pj/9zuylCov1NWzX+D2p2QUt6ZvDmGmnNfBoC/UDE/9rTXiVrquG9jKW5WFJz128Z6l
wm7hvEMmiy7JLGUb9820ZaQmiePBvYfn32WzMp2zvMczHbq1cnq5PktreVspcVpF/yuIg6oMYH6Q
uZkw33M7bu2SLOIRT1LFkQlw6i8fSTi4OMIyicgOhRWUpMnTUZ8nu2MZm2RgL8DhKe40+pt1yrtm
3AkCYDZfxA7G/PeHv6YMLyoSCvU4j05t4QaeUd35mW5O14lmRpg2/jTIgLn+txLhCxsa3wS6b5YV
auuHs5arCBBITvmE7uKnQynhvsPMDpcVJhlpW6dydTftYHs2kjAQOf0MD5Ta5y+TqznX9G+Gn6ns
ozeZnkGEjoS8BIvVQUHnqbSXwqem1NywKGQT6KSYqRKVDgfL5z6CXr9A0aahdPIXHjcn4N8iJGpx
p4fAp051yFZGmZXbsE5W7AoaW6DOB1F5civHCdhNSM4sdC2IsOHOzTT7oZ8cPJcd/qiWtT2RvP8B
r0AxryYq3oNVLWCv2PKGsGGGGjFXPHSGaUe/2kSYR6Y6todja0FJkYUbEZkKNwV12KLwvIpC3Cuy
7mzOH7S8QBalbtm5C8g8ixqQRuRUFtBd1HA6y9Zmfdl/1bSpG1B6p44rrvE+p9NTdZaOrR51JZej
XruTOL+HA+1E7w89PEoAEvT5oGy3KGFKMP7LQbNts4oS8caNiZKub6/eHsxWafYB2/D0R1G6hK08
cWg5sjaTP6FV4IF6DyYU0+uRv+gxcnctxsiBPNHIhBVFIRt6LZjwiXNGNrbtWp0F8XKMilT9PmHI
1trhqFkp605+mkjmysE+UBjRXZavrLEtI0JlxM6bWvB9uH26yllSjlHphOfyid205wVP7PJMxP7h
UEpbsjTJz1yLH7AZHZ2Ri3jEr0hVypYnAgc3NwSSFDTWrKVGwiEC1R3vJcUWeiMx7/mQI1p/S+v4
AfrK473g0tHXch6miEfyU5+xxD1lA1RGZ2nrFIUxa7w4XUTCn+WrygEIg5FO/5WCwZPDIBVbvSZN
mJRwI7UGnpukft7tqUeXNYSsmgZGsuAHGs5Jd5sxQwbVT02IAJFMeHI2p583ZjKPq8QEv1sW6WQN
aPwy8dyq4gUWe0oV4p/kKOgKrwDGQtiVE52aUBkyZ0ggPP9RM5q2T4cw8cE9M4oIHz9sbb1eTo7h
V3qLad2VpsntpRVBxbivO6c81T51Ekj/nmDkps/jY8htJdKhnU1HQU2xMDUeHy9fL7mhWXZD+JWw
ySiHd7zr6bcLlE6jLTtusc/aCkr9D/vagKZfhIR8j1rtFGfzFSGRiH36JY0a+M+XhbJsgzpeEgYF
KbC8QnvrazFAJW1zJG/7UYEwJbRafwVqDJuCcrhqPCYApMNG8rIiWhEDK/0PpgmJbJX9gNPK+xL0
+3IVbxa8ut9Yp3JPdhoPAYAUydWGoHLl8OeX2wUKLM1K5GhF8xFECgcxTfL4P7acHSkI7MU1/KOt
QpeDrU9oMRNOoju0GhBnUs632rqxoSyQ6QsRjUQTA6pyU6tZx2/XAsc1sBcQaTwk8W8SKQVu1Sy/
Q+kFPAOryhF1/N1BRQ7JOuTQPfX1+q07/WD5EMXlStdJQolI15eM/j7p16kT71r412wNMw/E4foO
hfvWloKsdaM49XR3DB7ifSO2Guht5FA5vlArzvaZ7XWusmoPn7gomITm1emfTYdpuxGjrVtjHubT
RZBWqHN3D+JafNq1KC/gq1EDi8/K119Zc3yaMYHjQWvE50ZHkq50Av+9h5zt+XaHz3s6Ay3aWioM
oEiaCrYVTnGnMmiiTrDWYXbPZCR+ORp/0wYbleKtG0sGtP0E5mBLGb3r33q+Cpzl9CGX2mPRE+AO
4QYpK0pFOg9Zlj3bDQxko4oBVB8ydli7iO/bZlCVXTYdKxn2CKPkHlqR2UPZH1XO8mBOHwQXntSm
Y+vd+OK/7dzTzJb68f0QL9FRb0Oqbx6x/Eq2c+8vSLL3aHSFKf2FZdrSKaOOVMLmrM6IMskUI8/f
dPto/Q2irV8mdcKUUc75M6UDwimWGaR1s8PIuuhNzEMgAhIbfPQfmy1l2gGL0DoGzEdfTsCbhEMs
Iq4tLCySLQPGCnKjCpUjKLy8jmACKTtVVHx5U5VbJaSXA+NF+r/O5okN8NwHCDPISCSy/B3pehmo
WuuTTEXSkuLs346cJK4GHwZVl29nQY9J9SFgTiMyoJBjJzB2HqMe69SNfEPB6gICgKRuIysLrRi4
rzo3c3EWk4ckHFvrIuB6JaSNy858V/W7GglniUDftkBUmZr8Wol5HyDZOythmgIbsvx0J7syKiYD
KtKYSVYoW42+4sTXCp6S87omZZhjfgQ0Q5IvMSuSWaiZFjwQj+hQNoB37SGM7iDsJavZhJ2SiCKr
7Vb8ZRIz3ThDSw8/330Ga6zN+4LPKB04hM2PJg9y4oPYteYXg+mUdMcx1dwZLDs//M2WWgTLePqK
+w7qB5X4Gk48zfW9vq+FQUlkGM0gk6zK7PU5zj64DnCg/p0psovHuOftMcRUp4tnSBFdFvPSEVUJ
CdnW/XASqSBXqKiVlHEBwVo8qtOnxa93KlpnhaYzFtF1VwIzm7xL+qriIGnKb+PmTBQNnA3lqL6R
a4imsPeyvXzfh5+Bws9dYCwPO/yOBWVE2ZCh3GXuX9gW4Dn9vflqS3zrP78mbIFsL5WB/LN87WOn
jAkeTkp6OAM6vRfq+VpDOkA3nsgAbYpfAJna5lLt92GAMBd8lNJxPAnRjBY704GDp2gb98x7eRZ9
7voc7BgFbfgruVWNuf2lSjGMmAu7vnF/GPzJVrG7qGXABzxVtvn8CZVeL0Dbg2QGHu1EumbLpp8B
jGpCfkl6aQ6dNxH0voZsrvCG+D33dg2FYiRgLzaVUQdIxaoj2WTQbRsazHstRROgiAOkst2+1EC1
4jB9TcC6g/qa0dkg8jZZYoseL7I2SUJsqenH444JIA+sqeriu9y1LNK/GlKXBixim9R4c59hVPtA
g6HhCfbCtyrXBvf6CeDnxIqg4WEtY3bMOSh87bEZkq7JcDbIif0Q36jS0nD1UQDr2Ii9GPoR9O/+
FCyq/8wzKrORLiFM/LrP1iAZZRkw+1c0BPLrbO4HgSbGDdHISNoLyyvaxLwNOolZWInQs6O6KZhk
MrwSsaz19kM4JUA03cXoBMeRRCY4zFtvImue/CTdXgMAy9LUsRqY2Xdn/e+mbZ0oIrm7PHkdfzLe
Yt3cSk3u7EPF1JCo/Cx8AmW6B0qGOOFysGVZg7IiiBa1KC1KR3hz+UOQPXYIl7vO7E32eMSD4ot1
E74uGDCZRX+bW9+rdzgCo96pUyMiV0CRhiykVdATsYZHjcp3b9JUAcq7eV3qWgU/jNm56VXqyW77
RGcFBDntO/9DwFZ2qeti6XF/fIqDGG82O9ttxOZwV+DC5ho0Rc/VMi2qIbxeCs8QmZqrodPjYHar
AWrvA/XVAo7XGCsuWR8hVMkYRd2LHZWpPlycUsIAwO6q+TY+3MH0oJTfRh0UvQc0skAUDGiP+WuM
cCYhnG3GXKz5XbbaThbZfVIkW8S87gndQzJHKLaZmMWy2n8l5wUU8I4nXvZd9nRoRqNg6lV4VrOX
JECOuOXhwBBDy0GBhNwM7jsRNbIiLLqB0ZI9ZQZr4hLmS2TOAt+YMIRLvFnAhMovNrdSsFOKGKPf
xwjPIakq5DflFvNIpDJB67FpUPrmwLloROatdKxlu0UHqVbi43z0JRBIP6DLBlmSpCp7qiX4e+Xr
Sk5w+TjKg4+Qgued9VWY+bh/mS+u0XgNm7HRXBji6zy62WxsWIadJG3UCWUUYd5CbtFZlxmIjDen
/yWgULuwcymZoEw6DCuU8gMsBMzTPQlV7+7atlTo+aiK94Rqo2R7Lku+yKqGESClf6vRMFdJqQs2
C59Bu0smM4ZoSdnhN2qyeCEN4ENVsmt2VFStI+nlPKH3wrjmp5Ibe8d1bcS8fS2XVjznajtDccRQ
tGsRQICNELYHKiGqBi1IF7BuT8y8AQv6iOHraAtl9k6ct677SECsupnaLwKwX6//RG5hTIzWfi5T
eMDdtw4TKYN65YzaTCDq6qAYck6m8i9UiNVvzeLhzwBpcDIQSfOjs0N57marlvSfEcOv/vVs8YXo
RZWw0AP0mKtj0dBasX22pKpREzXHtbjZ06tc45hseKl5/uLFD64+7Bma4t5i+PUgQJAi3DWlvVjw
JBWtOwASaIb0llbXzIS1alQWgFwkdgm2fQ6yS25Ejb4ObRgxSHUBWW8T1OVt0lorkOZR8+lbt/Hk
hBXv7VywRLv3LjA2ilM/diTXnxyNj9zvlV3fDNOs7+H0m4uDMUdGKI5uTyObP16oJUGbEOiDRJ9O
rVCENOTk2zdAzzlkAnNtsAoM3z9r6C/1uxwMD9JCx2BRyBvIFjzXb6orPCjgyY90mAx+CyLYqKsg
qe9LE3S3Hd4PM0icmLR0LcX5TYyKZYiyj7DBfAWj8awOUeVrlYj+SyhvKNBXqX1/dqO9ZgumdOVP
p1bDqEY+hFLP8m+Xk94ldnQOSI8mSc3Lg6/GCP+qN9lJ5igrDuwQZBTE5cwyfZJ9dyz/Y7WgBhkt
5AIXEBnjw8C4jyrMQNAy1rP45gcTDwhJl/nChKSiOLzr097m26MkIWIMcwGCBH4szL9dOx9FJwUG
g5kaW8CRhK8kny/+6gm8vz2qvsSsfz/ONHx0ZHGeJTZimW/Y1xR5Dmrsbai1shwBSI5znqPJNDNV
u5hqh3Jnm1ubRSW4m3FBsIUQe5jEkHQecMV0zDqtsy498RY+tdIM8eFQRbIUV7NMvkVkw2vnK5pQ
WaJDiXr2z0cC9FZCSSk04OXe+HXkZf0V10W2wwQox9lcW82qgatEIRRXdU8QE8wcTic+0SiOPDoc
6jsdgcTEy8HcBJtJM74AVqM1yHjeFRrFNPyBfhly+BN6gvzW31NS0/TD2/DDocOG1AjbO60J4cdO
dJZ5yTAPyUg02mrHhdyGCYKLR3UQTaX6c7pBBt58pzoBXPQPpDscxd2CGnxk7povBRWvk2EDkxYC
0O88Tki8JhjBqW5Dv/b/nMK9vbuif050+ob/Ivksaj9yTB+dQDkBXCgYdABzIvpWworJSVFyF+re
pG8kr/1r5h11O4zBGa0iorBIWMg8KZqlPuhkdoYCbRle6AgM2jfTxaX3lSsJyY1rj8iLeK6BjwJC
taMG5xHQ7/ITVvnEGhVNDv+RnoZNH1TallwHWTHEJ6TsIs/S/FhL4ZK+Hq7hDZLnAYXNSBhoCjfZ
ibWzpZ/3UAVtthkJ8f+vky7nzpJnR8mkiAL5L4PWMOebeZXOlPeSBa5FsgQNcP9effQa7+lhpHOB
OmTAN915ejwYAgsLWnD96fN5QfoQj/2Cl/IKTdfkHwD1TqfeWLrsML6WloFLdOxeM9oUyiSkmfCd
LaiKBPc4+xWoBkwUKIMjbAKs/GBFfQplKFF3FMrzvCjae6jffbdu6h4CN7J2OjkY2c7tfMVfcbrs
WQbRq59DtNANJIuzdY4fv6i1RIyHF1Eu27d2uBSGTGY+eurCdrlS2TP14FCqrtbRTxqcbb5iBFwG
WI9TQGFy0AGxnD5wIaGYjq1+zkIwmgpD3iGPsFxqABTbdSsT9/RO2Bk8fvh3JXmOM8iY01Pkuvpw
gzHIvbUEWUw7I2pFwX50bfquxcOpg203uGwzGoDSOttHRF6X9j0Mo5jdYKOP0FPwHri+hndbfXpp
F1GAAgXcGpj5sS/oKE/oW0IXfsDiwXPd4dafagZuFA4rZeEDgsVZjq2ZPWK5MmzvUaR9pqB3s0Ib
flCG7x441kCAhbXMkL0/Pfr8CsVLc/fOuHdcFgayvmaZEqEeoAV8LFdAPgPhAsB9CfK4C+V88r6i
nwuT3U9wU9H92Z2pExwxQTpfBp2XcmnSPRQ4MkgmkTJot5YUM9yfMtY4Lqj5HniyNxCwHeaT8Z8g
72vipUcZMpQS5XU7p+1kABo8l9pi1Fls73UvplpgaawQ4YuG1ysrcHvSusCKv03pFe/s+4kyooAz
fWfQS5RBYc2ySKSwvn6l0uLfdKFGZWkaP2WTgksxA6utOu45XBldkKC8TFM/NnLixh798z+dMPQJ
IdLvRVAQ8Nb39k/Fw4pYWD44Aa1RlE/1pQNUq+5UhobHWRm7ZvQNqJ5XN5CXBQOubY/pBLbUIASS
EcV0N/1eJ8e7hpAJTfuB7GYvNZcAPzKi7iW2ym1dat2PtF90mEX6nCzLoFQl2gobEoDH7aWRAiel
1kR22kZ0GWQXyZ7KsYiFRvTpAg/rGztNJAN2rmnWFJ2Mqir4jvGaK1swCpOwebQ6EJzcuG91LxwQ
eHVOl3qajw3MACK57/5/CtePVpvvi0rdg2cee9cmlWudWX455xKLP4ZGmD6fJsq1TjukA8BHswes
Ry5rH510TBeHBnKj6A1a4O61sv/nk29RdRZI03NJfVkIlwrdgpVbm9uopzJoFoClsYzTnPFYjurK
UKz9qEDWIWl5IlxC9AldhO/zOpx4Fn4sh71httbgBdCsD7tsqwZjXM2RW5LVkTYcb1djkR1Af86U
/b37XnwshiRplTHAisaIxL6ud2P+8WIiYlOusj2CxgkOP6ulGvxVaTKI09PTNJDJB+emd0EiDDay
WoeC9+L80+YtGS2fvZalz4hO67MajqaPY5ytJKGVoqMgqafGaXOt250H5czg9dsAIqqfQaIyVph+
COb9sSntk0fuUQKbmEFpxkYe0MgMVfWY4wQlF2IgG92gjVZfk5T5hWq+yzhlz1DoNVHXOJxSNuch
BoIGQkbuAIZ2x9dY8ZBT7j+qiVnPUZdxyE9GRLEDFhBtNJhpGfx99bUoXYwTZJkAfOWUdG1iP+L7
8ul3vzAa2qWMYLGoycaNe4rIfEB7VyoJ4dG21vvz5uOkF9LNfmyk+NL4BI0Woqry4OyozOpLP5yd
L43LNa9q87fJkAUMp/N4WO/vtmom2ymHAZaNWKj4iymV6Xrw1UWeuWo3aGHnnzNawnnj6MEnWiGN
AtRFwIl41jMgo5iflFM4/6chLNiMxRy3iGKjmcG8hoqtW5lwYc6Xg42k4O+rr7JYdCvQih/VgRIN
6kBW2+ue5PcmKZhxJChg8dv2P8uChBoCXppdyJuXXbGDZ/VPgujip4j+KywaijUIcAe1PlZk8myI
iWmFmj2DUnXHmrkXlgsAHaOueZazAPT7AIQRGgQUFCE0omGj/cTrevnSEZQkxWZ39jNt4PDfKMHv
6AEzlvj/ERxptiblVXw0QYK3lNizOh3eYnWDsByOy0iWFDwM/Lvb0ylWZBMRjlC0U+Kv9Qda7QtQ
iy4UVXtsDjn6sykYjWwPS0TJrCdg2AFRQUEX46mBGyfKvte5+MRc8a9SfwrqS33z3zmnCUWxOxbQ
k7lh2qlAM64hH3sdGogYZz24Al2HnCyJy4aE5+wJU3UBKeZhY3oT/eSYYXZ3JNhHFzxt+9r+pBcI
la6mNWSIiI2nrY4MANQOI/+zj8IFHMt+nFhaYgSgoHZOgNBt18spwu2rU7VZDzosS9q1wuUTiR0p
aNGOlkqL+T3kLhjjV/CJ/XFaJazAOF+aFhnRcDfEoidwDi4bK2i6S3EmR/9mE9lDX35UFmx9UZJE
I9MND902raYdtvj72Le+BMiUGj8llgi98RYNZ2ad8ybWGh/6uXkgDqiMOBvpLjR6cK33RMGLNkVn
WCLZV6wX49MHTgzS+rdcLERBVvWL40Uv9vfZ+BEq2IxD9EiG5nCcWDUvm7P16jLuoSZKVjk2JB+C
77B2xO9WJEFMrmipRO3SA3LHSw0oK2iexnd4o8OWtt+2d1qBIwOtfCTWcTK7txyfxcUETbo7+t7e
PdGiU4cWl21Dar6UPQtKwDwoCILaH0joLzeE6MzFDpMUzy7JqHu3ypXbD3CjpvM3fo9xrdaMkuNr
Lrbvs0XOIYQlfJiUx75lRlXPXlTgA0j9Eg2rNyZo/Qn2uAUHfzZMnKoReh4lhAAnQ1ddg4Ay6YSS
H6dLMRFgaQOw+a5UHrugAzouBPbxwLVSOjsITcfxE1eh3USnuiZ/+Gj7HuvlhUcqu/8gfTlyr14w
brC+PSbCMIfjH6jrNk90wIHEt4atRMmCLP7YkBYOi5OjBe0R/9EQQ0teHylxdRop2NIadFMG+hVa
WhY0LREQawcA6gELIuwwTgIwTf6qCT0MYxW/0vxczz2aEJIrp4/7Q2DjI+ClmVN7vGr7OgvafN9H
36Vlwpn7Hk+M6cW0rtbFVflbTMRyU0qTeQFliOIbd0q8tKno7YzjmmKGzRH18twPCIA3OosIk58t
qsmtVGAprhVuHSI+kQeN/Xz7vAkgQsGKsEjcTId2L3MshzQ7FgFGz2Dhk6O3Eyh1JEXu2ldodg9U
vwUYaxB8Wuqb3TsN1F+xMxBNs4Lf0K/7Tkhf9sjmyMo7xNfaHBgbHluk/T1/BFSGLoNnVnyNLl7X
M4CbBtdtFBCDJn9M/Y/N9HO2Pin5M5vC/rWnmKmMCUf9G9vvfW5kv32T9XKL+xrEC7JF3N5jNRca
MEKUGk512VGHO+aMeA4DTmz8Z1tBAEekIyXdDj1xlme+cQza8LK/T9imrAI77QDptm7pJifaj0VU
XzvuUq+bPpQKtfI3U/AtXWzxKfWoNtFBv84WKpTkcmBadSK8roe8Ide4+76E2PfTIuPft2EUXDKD
blPYAlUW7lQkaAAMi+7R8wfkGvgDajQMBma3HZ0zqM4T0gULovHvczBmu34mtlmeddL9Wlxflyao
rO5nUBEs/K01dgK272sB7LMTfY7hCAUm8mo0579MCTV7MqBdqy8+aveP+tdbuNIJwFcphCCDs/OZ
PIIeR93pmTMxKOw60B4M+5od/7KCoZzy5oaMKQ4C+rV3uiW/OXrDTCyPBwgjbeAwIy+hs37fxEpH
55TmFnrlG47YVeRtT+wuwWvzVVKrLba+OeHdlMvCl3kW4s+SQBver8WaDFVeRx5VlY7P+bppRoYK
5Oc0Oui1ykiGEOqIf1S4NW81m5JUMFIgfDV0B9dr9J/4nMeVpyNBi+ZEAkhkPl5NmWEfTEIOdOUt
9KIDaWIgw09jAyKd2RRmHvevWbuHZWtvC/95DZcJXBZt52iiBqQHmRxqqtWPbKaCTvBoDf5hr4/W
lJXz4k4jvkcEaVYxzFwTcwJqApmwaGG3t98m7xQ0UbvkewYyoKkuFNupc06+fr7k/F6UG9qAS2UZ
0XLUOqovl5k0oZeJH+pcUh1jVa9T2wK54gbAfiqqySnlMt4eq6prsIK45bsthWYhjr5wCHjVU3yX
8U6Oc7kxLOP4XZfRtZpYehF2xVbRRIxTT9pP7Wy6msbMXcdGDC2pbt/zkJ6fhusF2wlNs5BYeuOK
wkhy9/BK7b9JkxO8H0MNIqf0n41Zm0M6NK4k2tHJj1AgiKMhBlIBXkjBKWs9/iXHasAM7U02Az4v
xlNOlhtKn1QW5l7plAZ+nSLSB+qPdv/EPtKBYlF6v0azt9WiwzBTGsE2OO09PYLK8mQ1x1ZbWnn7
rhqxS0kdECDTAM3lnT4EV2NxFdKYfkdrcZ9fRpwOHE7DwZ6rv94bn9BytfTRdIXtKH/K4PDsczhg
qKmiqBNFv50Dyecw3J4fzm56+ANX8UYo2FyNyurBhiwL7ZvUozlCrvpWxWDclszfiUIQZTzLvXmj
HnBgL1YBZC5GTLtJNrFjVWp0XDluF2CD2bSNrLNRYWe3TCuyKuE1C3+TjV+B05Y/TJHjeINujsz3
OMvjb6cGgs0yqantUEbfEKBPykrYWRRWGsGm6PdPLuI4U/61JZ0NNgy3IZ36miM3eoDp0pn0TatU
qe0c8LbYzcMbxy6fHokGK8WaSoMrgRms+uWCbqeKWRSW8RZv+/Y7ArkVYiW/EryYcKrF2UOPKfzx
PPhKYFGa3Huu+s9qjU4BPxVBUwIe/1pcYNzgp3oGPq+oIh4RKCa5qCVRx1d3m+yzDaCJckBRWdsW
X4D0EzzIRtzYRmiPipGHc3nzmfXtSRsdfTDqeAIGqc2gYHgfPwsQumlV/2uBz4Vt1rimkSHu9q4f
rLMhSMfqsCeTZuKH45F5SZGmcvVFa2KGlbscNtTjgwI38wboKDvNJ0D4PE/qFRtVgtXYOl5JQAIr
XWD1CCg7IID7aeUWrwhbcSJGSNYNMBXsfZlWNCm5b0LcDMZ1t4UB8XaDTTIqXi0rQ7pz+d5Z1g4B
yvgiesSvLbcMG907gEVxV7VnN8BFM5QbrpNkrNMBCDoqjeIp9hM824rO+5PR3j+ijyhORjUf4gt4
xzu7IxQKHJfBb1b+fEJgHWzJ6BHvopyawZoAcxSduGyBNlr2oKO7QNQq8aFdK3IMEeeWbYrUP1OV
DsKz4LsjKe+rMqYjIKvAszuw7ozPfRIMfPdWFlzxo3vzBkD9n1zEDqqxlzAPPI9kNzIuGHyJOvB4
IzOY2IPEbamXlhURXi3H6t2pNeUGAzwQLHoawogG2juEcLf3Wy64HGrdFxyr9KxUNNYJ0mRH2rbr
Q52k+9dr6otNcC2hwk6v6uC/BxUfkOqZiM4EUfMV1h6X+Nj6zVhyLSDLPmE0ogcxtnM6Wq569KpU
NneLqSEkqlySGIJ+pU32CsZn4NAWJiqYacbLCIY7qa+uf39/gX6dJHuyMzTQwZ6sw5I3Or0qhewM
tkqBIvdvHokSaB1xlKW3rUgPMVckRdYFmuO70j7zRzcc370DryZAwftrKhZrkmjIiz+PQRcrT/me
6GXOR5Vpz8bNBm9+uffUZbiyu+ZreID10+OlTzPdFyOBohJzHWSn56wQvqzThmmeJUeI9OA5371e
KaCOhUXDCm8YYl3Xn8RMOMDjcT4gH3yByhRTVLpboPXA+NbFIyb3jOQ89KTgoJjNR2AxaxrINmT4
uMz5FbJctL9uLeoTo4Z11i9wU/6ESa1pA1NwwR/2KqW1IKxmmTJpiJM3aL5XuJbbwO5maOVj8G3I
ruyzoAyGi/+Y+vLdBAlvFv25xXT6Djodi6dRd65FB47lVxadX6D7EB+u+/FoD+jH5m0uJWKBmPaE
QtO9rRMnASyi31dzlWsWpUXBJC0hPk1vZhsNZa4UDS25IYCnv+Vr1+oCO5AIMbWN6z/TjfdThMUb
S1QL4LTIhMBL5TkTStdTayGgvWXJEzbJgwy4VQIL6m3bIQ09u8mx3kbrY5gfzs0JCAgT4gtnVkwu
8y92lrIXfHUfn7MbQXS2HRBuWey88kXpHB3a4zmCtImAK20Hv/LAT5++p42FZjH4/mM+Ft1NX0tl
96lyJ6rTQqDqqQgH6pCLRI+kzfko0yQQ3H2PfpB7ExarI+M43QjfgNygraDqeKhbrhuRZLa7/R3Z
F0yG107tPQTZLBtTO4CV8laNfkHmighifFpEbqCmdTO46mBc6mcWTrC1JKkxjpENBHvYjKCyM0dT
8mVdUnRDGDVXieDtRrXk4IqHwqlot5/W6Wo3BdguNesqP8v7M2Mvbce8WP+7wLqIyFecNRZrN9Mk
1NdArYQtJfZ5GqTS2Vh86buArsozzBoq+IlymKtLO5mChK6J197vklBB1FEjomoOwc/MLpRnSXme
n5LZf+8O/lwTthNwmg1ONCeyyA9b6bX7ZHn4VodFcskSzJGAIZftrURVJPF276SvV8LOSfztKFUt
UfLl5+o7IXTFVbhy5luGdqwWncb0lvc/2HLfBB8PJnFrQoWfHaoR14bNgT9+Bz6uRWirVTqhzvkr
B8OEZo0VURZSRkxyPcfk8U+36myoAlhW1aEanagckFynO2zfL50GUFmtPwIrr2OAy/h4pWEDv++B
7jH8llFLwEOKpWrG+5X/63/TIslXVn6rxF15ZFJ9NuGSYETtQ2iKDDvaqGxt/cZc3UixLe96Y+AT
ZpYTVJqK2+lvdorqQ85htP31J43M2GenuTF4Id3FJXhUJIPX44ELxaAvPTJUtIbOnhNHD7gKT83l
hSdFWd03Z/D0nC1XJPbysXKIvIEGGdttVdCQt3bdN6tm7fu2VXhXmnGyx3knwqeQKRXSuz06018L
V/8juHIaANB0OIIW6S49ylP1X5TRF27CapK//tjFg22e5+c8n3Zn+ghd6ggppB95oHQbnb2w+fVL
xCY5iy62zzlN/MQDB8ONNUkFataJr2jObCf6EDiX1mXIVsU4WKdTdQ/N19ySOgmrVAP6gdCk8OlT
mzNk1iCZqRtKc10MG2XYtk+KV0sYX61z+HQMOXYige3Fu7o8mAvl9THuGbAohHtoHdO18QV+Sz7d
s2eKxWKVSyeSRQaBaVG4DS7K8gyVwZgW0W3d4O1/wrYHr91bJj5KUxGoNtb6GernTMXXNyVH1YHa
Us+3PQ8MjjodT+be9D+7KBHFzM9eEvbozkdO9tg3Q8Hsb7fSa7RvrVV+OPdYMT37Me7JXV3sgPrT
ActO7B+lOOPx9dqlDBVNF2tNOHd8EZ+/oFK79z03cPXDrJsrx1MRZGgLMBnSpFidPvxipSYlneel
TBZyd0oJHghFttxunEAxsDFVAGq0L1aajP1I0FFhUgvoRsFSGLzcFpQzMQCGsbGYSJp09QNoTzZ3
nclf0mFwv1XGPxQrKhPB5WqnQGpckZcmNQ5BS5QPUWK38KRO0K0brqAsYTzzo/nTNA6lMQwVoOHt
wDRn+fZMOXAYVLA2fzpKwsgsLuLHgXoFvDzSZr5SOiPpt/R7UvD3I/h/wrI65CQlWqWjFj+7TKP6
Ia1xIGybJAuO80rf8U5KTse/DUZJ9KAZbj7B7loOuq6w/KjycGO82dJLHruMVGePZJBx9gC0sjLe
33CB97Esc1fOoVg4cGbiAL6QxNQReITMkKEvqoXEx3d0MYM6kZ6iv3P7wdVYSIZW7tBudt3Ooo9r
P+JAK04KGFk4TbIFT6qp9eOAObhbAkarL1sW134MzsBdGetYqk7e7PdmF6IzcEsaHUpsrpJVVUGM
GBYOZUGWQdXiucAl0bdzNQz7DeydRnpSITuSkHTlhMGExS99HZWEmKPNuWwVLPErJ/RR8GVgZrjH
OL3EiBd8gTvqhHLYvZkOWmvCqe8X16SNfmNN0WIvkTAqiC0gxfRvIAn3RskJGryCLQX0kw9htqXN
yBuE6B/8JibxfhchbCofv3GCeN32WtWwB5FLZxDxT8xG8iYLfj+L6bg4i2Ae+VLCiJgfwb1WQTku
4y6tGH42Iq/NZqNCM/NRyKuqTPEw+qvcr2toRxjH1RQ2Ub8TD5d0GM9fjbo+L85V4iPHyYssGMQy
KclkAK4md+itO8xo8GlANhKxKo8H6jq5xZJKXqEZuTjzPsKk4VslwGTJg83lC7LhSLfun0UzcfWO
YPwXXDSZZ+4DI0VaOI5dlMJYmu0vPITGkS4iuLpA3CQdD05LfL3cjVJmaVLDUV2f0KHlo6ufRbRh
ISLRcaAzXrQbqrmYJPzyzISTN2aRRWxgcLztixOP0nautsUSoqbcu1CEjbHv9NnbpkEm3jIHdFTJ
cZxSa0dKqV7U5JkOzhw8klbeS6f0cfDOFgEBsDu9EKCRLz12XNkIp9QgNw2+obKy8EFX3QSdNsOy
UfaZ8+rbpDR32XADkT+wfXHDt61z2DU88fYJM/B/XfOzI6OMoYf4neT3Ws51QBSsHGsrDrvAEzTz
KP6XjGPYEto4XMqca0HkJUktcmPUHvfRU1duR60F2GP6MuK4njlTEhjSMRNLSmv3W3ohFMfNG0M8
0k9h21aNQnDs1X95qcjcQzjO2IC6+/WukWk5KBC+/evATB2Onv5HsUpfIZ7go7zVo97dgaEj+k31
6bU0M1h53nbAYkzqMS1OmYwYX8/Z7LwZ0TZLNSkEGsk9eXSURRPfzUaCvC30R9p7ocqu1HEEwWRl
6fySZyWWMcHpO4SmGrJ27Kc3x6RKzE+3plu/Vz4UUnrhtmgT8uPmGqcgSafOWkvo3/AiCqqgHjSq
bF/090O+D7nHueqI+LLWqyjzGP8znrrXQQYtF8IDXgEvKMHrjN8bc0BA5pBwGjPs1UkfQymwTwxB
djkJMYrgrI/pQdvXjWFeOA4OG+8P779gyVg+6VGF3TfrQI8Q2BLo+vDTcTQReEz2vSe1biMP3IR/
dvSWNaz/h8n3uKUvvHxBRs5ARkqlXA/wOj/RNZnUbc91ofXsbqsdrqV98Ckk4xeaqYzEtQOgcFw7
DvGNjM+O6c/PwvyXYvdGc4iP3CTesRQ6WV8Xh9MVZm4tsU/h/dInB8XI+LqwkxinrN+6A+9Q4Xut
BDU71J305FRlTy5AzWmXkFL14KuVx5Px+oDa7GqeYEXBn4ivX0X2a2lytrQwKmBmCEb4rGWgrEH7
Dvjo3ouZdHZ2aVC7jUGsmmilcF9lq/Ig9/mXVsQPtXAL/udydQKOMQ502drKHpWELZURGj0Ucf6R
S+Jy6O+5o11YhdIxOs5EXNgNLliZ3vHhhotoPQhUnkTiDC3Kpqtxoglge4vm0x+Vu9Bf4mraCs0E
jQXVZ4Pl+g8sNTs6g3DAhgCyaBluGFlc4a7jcTVZi6LQOY/WujuNxGuzI0GnnmzmeFHAmjrzyNB6
ikhn7zz1rhgAnVWiBzARWHvC9XXsOAqC7WYLP7MUqlc1lfQ+EaAS7DIUEwN1QHoZMmj9093eSOvc
7AI0hlYVr4KBhgkPkYISvNm+DRALtngXP42bcjhZHQfAVuHsPcoE9vb3yEC2YNJ4aNxnm+PtlMlN
z6byMw7l9UjFuYMY1Hwki2qQvmMzvhpbKacwKa/fvNGL4AMHIS06L/y8Q7I9HM0/eE6W8kojquBV
iZbH6JuyWX6rtdELlka+iRodnM2WWV+u382v1mfOHg5InVzTNpDwQMpsVLBeGbwzZTyVW+Ze+p1p
luKBn3zntMPd6Oim43zK+abFMi7B7bsw+pDM/rgemLlbpApJjNIQJyAqmd1I/mzU0Umiv38OGGlH
LyRrr4jsBFtexNZywXY2N5PLCDDtVJYdYH+pTY9lOr20x1Sc+8b6CzQR2gK+OTqzsCiMm3mGp7EE
XpmdPLbQbKm6s1zgqjwdYhYWFe3fvFcz+LBgA7lCZHSAodhfIgRbPNWeTiFENPVuoQpyUFOQpW5J
Kg8w4MDmuPDg5mbrgAC4zZjK1mPT6OQdz7d+LW1o5lcBq2Y3WU+BXXs0/duoCtiO+7u+53XfGMYK
dhufhYxAedDk8bwXx51z9goDqwccWsub2LnW867uqa4KB8TljpquaScxhG+Yp83nqkVUcu89Reql
LfnFlZPYkO6hI6x9Fwpk9sSv+BtvpGBMejCHU0sACXulzrxHx1RTeKbLAqrrMA07zf84x12gPzAf
PJcsfLCS0uGqUmrToKQiUe49cXlGIJIfvcFLU9bSyrC4r4W3yqLtvieAstU9/uC14ofMihlzAWMj
xvPPkSsIq0fp6qpBnI7YfKAtN4kwQynM8y2LY8ukHmwmJaq1QDqDBRwhEmsnyrhHxMtl9RojOaTY
rWL/umEBwgJaOMFGxVG8qOOuu2KOX2KefNfDhG0N5NIF9tmrJpT6QcfYArOnubs5ZH64AAuuIKqw
xJ4UCBt85Tw0bl4MgGjyvQ0dshqslEkZYrsQIzoZ3RKp/oZRZ0/oGPSVdXRAFFuKyt5YIdo1P3nk
3nll6EpthPuF74SfyvBK+wHVQy+3WqvKsHMFRGJ6nXrJHw0KsWXdM7u2deQQ4Ml2Mzv6jgzJvEhO
gIovbz6tEVZLW7gnAEzdFvrOMgitAfh/gjvVEq9tB5FyVsDnthLiqha2Nnbk9uP+JkSc8jnnBXLB
B5uXgEw46Mf+VyfdOq5PRl6b1Q5Z4OY2H4Cu/NzPpxas+1RYSSHvtayxAtdHz/0D3h5St17WG/4q
jyM+6VtC/tkh7wozzHtY6WjAPIcew/lI/cZFXrSPoVM6TDLqMGUPoOVdO61zfuJrlmHReYWoIWvz
8dXVcNOohwZzb4JR6csORCBz3AdLyr3g0daPp8yURqM/JzNDqNLans0MYqAH01tIsEoxECgk9Py+
scDabKlJb4MbnNsYFnBnQbxrcMVY3QImZHkr2se6tGLONysn35shO2l2vtm8bDwQfuf0dTN6qx0p
o+sJvIUeym3wc/PS/frDMFt1F6zeecDVj5U+iS01Nzx/sEeFaWc1qgFyiw0GdUy8djUzkrt7aHBH
NlTA+ikg4bip6eabENouzjyzP2CmD+HRL9vT3W2ZEKbKwKxk+cwcU3+Zqlb7kcHsKLw7fuYhee0V
fC/EXjSiDxod+OKhjT41Y+PUIr+bt6Kg8RNRh5VZJryMMMOTAlgIzYyqVx0MRZMOscvPqtHo8ccP
awYuM5mZJZwUtiBkADCQn3D1xWgr3L6nCgTd3mOS+JhLfF6YgdHsgcy1HKUS4pENhbaUUXrkb46D
fa7Cah3KTeHGWPxGBk0ngY0+y1Jl1AciXQgMyPCC+gy3O8PoRSwFhEYkNoubUBV3L+1JCI4oRpMr
LGBzbbfDhz8O5i4WcuBQilmc6IEy8trlFkOiVbKMP3Z1nYsAidtv1+1Op1azhoFnf3/7y5FXxEC9
mzu+0Z48IsmXS8LhVfM/DcfPJD853BoUzbN+TQXmHDRKFXODjUMqFNglHfwMCWjlwrsZOPQrql04
+0I2jQvhG6ve/BTd/J6VDkx9TrmrmC2Mt7TrSLGieJoa8OX+kIpxrOhzgst903ONotk09vLm773X
nFDSdmLAh1d6AzTVkt2mA0zoXcUnX7Xbt7M84HgYKCOyvrOmJQ5pjz6n+Z3+vuT/vCnMh/nhvkV7
0+hf60dKYlson0EbkLoLF/9CrgBeSzc4lz6biLNtG+uzPpfAIok/ivlceONQNB63WtiH77uvAWdn
QneufqLhpQFN/0t/wF1FXxvIxVFuMFw9o8yQaXThQPE/arI62g8ONxaU1b8JEJdpAqJgeJQqasoJ
IEryTtePpQDfEpLqH2w6KOuQwdmnOnK/n5yCT7WfWawXUeNGKcODnE4zBnSDJm4MXfRX1DHHjiLp
xMLQLqzJ1jeQrcPUIILHUFALbVtA/1Fc9+gza5aMBvFMnmCwoZyATTd+ZJlo6+4kOXXoeSfbPwbC
ICsBtyiekrljQygW4GTKbrHv0LvsfyI3NR/bt0tfhT+tAhlDdgJEjxjM6MJmCVEcQZGk3mdAmvaN
W8KrrSEUTG9FJ6/ptRjoeM3XwmuMzIjC4boV2VGk4XIsIORU8MVp/wHpBZ8KDtiL68s/goazwOJw
a/0+PEeBMndkA6ifV6Rngf1pmxPzmKq0agiVCrjVFgRJ6FX8epxVWVdYa897w4exlLuIHkG4MqBB
kmfVtzPIRJA8a+Nsdx2P3CRnVOzUJiUpwtjkbmBgN4DWpTlGZEpaxWhzELcsEMpMoIbp3wBF6xn6
Fux+Ov1nyU2HdKkwTNmnUvbqWdOvB7oNIZkIhUxO9FtsdOiwyCRZtA90C6poSpVQ75rtdaJbglxB
2hSc2TAdfVclaywvKhJlUML1N3Z72PJygrrJDyFprYgWVVSLgB3klC0Id6+vTDOi/kaXmvlEmlVa
eFLANaAaC9locFF5dQ6h0WetlAmcimoZFyjxIHtOW/nv++FP3Clr4OX1RIh0vVKU3j5+J88CV9OK
S77Vp6B2u9cEBEn9HNEnUQ92p+RcZQrb/zNwWouJg3s7xae/iYnKxOk6NhQqnbi/yKXaG0kn4yOQ
uoFDvSYElYG8Ru2ep8OkpeqcJ07DQgrz2j9MAqq+v4NdbYD2g/M9iE3ZvCLBLvBX07GeuCaLPptP
eesYMPddQJfMeSVOVLksu8w1d0+370Y4Fsof0s0+iH2q5zNDclbuX1cmVW68ZuuVxXG48apNgnuW
nWVvdvLu2zeuVtG+mcHnGcfA5pOZNZPjGjjnoRLq1kuxHwkaQQPER3x1rSdoaQiTR+TyIryy0N57
osVeiwJKmettZaArpMfWflG6hX4ApxeNzuCFIONvNoTjGlu8/KTvlzYuQcQASlT4VH+PCr9SzE55
rhUZjayPtRmDPvTC9EmlVhlB5Atn3nGHOZKnAMdPL36IKppeRK51/5xIu4CYvPyql1G4g8cv1MrF
3k20Cghp9UOFRitptq0rahrQWUAHdYmvr9ejnpCuX8QsuR8n6MANPRBGI/EiJCmy/keKwlHoeRXg
Cm7cv4DV2F/CxETD2oxypwlmvZne8OrvmgmZUw+HCnRxqvUVpHuhxsv+9mR7eydZhpntNy+gbj54
87ZXCIUrtMRbm86EBN0WmiwXlK53Hi9IL/+36OUvzaLHGbLJOfMJigdWQ1P7u284OhnuJPC7cr3Y
lAIb6gOWJplhP0VyEIL2rFjPJWNElRKmTYQM/UWo4UHQefJEC2b0pjfpx2ktYh/JeyJd/kcEyJXa
NT+e6kZLNosSM7p+UxAdIcNzbH4DiwQP8iZDWzdoYdpeRqga+vbcpkyDEFdSmkoMWEom3BsYE5uW
g/lXP44aGixyQ3PYypz2jIMxjST5zlyNHL/RNuIlqLgdFtjTwXeCYIzkEnoqiDV+e98WCDc7Ij7D
NTnLEm0WP6Ux0lBXukGh5VlsIfE78VBo2lLflhpa4yKNo2eXLBs8fJcMJjqRj0dPO5m624aGYUEu
Qj+prNr26XoyKJchVyZtXdgqBodE7yGxCCQsSLKKvgDhqv3d7bDiPGo8aKZxwu/944re5DLHVFDX
j13CZ30LqUXlybRzPP/Silx5RHo1iG0CotmU847UTAB1ljWrdAqQQaWaoz7p42jnxuSv+soeitRd
hxZG+8KwMzYNl27iZi7rwZOvJ9FwarKkk6BTZPTxlpmDa7loyTBQjyVvgrAJpHY013ORJVzLrjN2
wvdXD0qJwwKpkybOt6M29Q1BmI1MPiCBFEPpAeyjOBYD4u35Ruf7E8L3irQbqlZgTQ60hq8IgRrg
sPX6Y0JS3Ax14MXklVYWoyEwKGGv23xcqT2D1q5ISvIwF3ixGHTmqXEl2CAne7dQTf/SUr8pk82J
NhfH7J8ld7qT0zYu4Gmq25Y4JDurzX2HH678bXUytcEznrH8b5NJqPV+RtJeyuHVREV7DIhCup3m
e8boyP9P5x6bwtnfHzoAFsl4xSbVGA1ZmdyaEG1YJtxXQi/NfmDPzH17OFNuWNREGv+mEvlEHiLG
r6bmd+WjaNGxLfM+x522yQnWXd8Pzj+1w+AsYmDKVHexMn4KjuSqbLud5+Oz8XgtMHV5RWVvpdvD
pl39RppUSCexjtb5QB32uggKQMpPJ8RnczgXYsOsL11e64gwHgttpy5vTgkHYQacDMJ6biP8ULJZ
Yd2WK/zGiQ/jKPq3fp5EcnnIndyGETauJn8ra5a0K7dtkEAM9DIxa6mJxpx0LkErh679K2JnfaIQ
QgHBdN8+9+QXu8efu6vXO9368WjnCw9WJS/3y4ErWfvV8hoAiiuqy5/wvkxP5Di5MIRvKV7UwceU
+5vLpFPHzwdj6duODWG+ZZXoUSJpk4tsjE5p3mAp97UYszPYc54hqvpEmXhtx0sTDwsca4R0dYWV
K+zDmLJE9Rxcf8qn5TRNG0lkJsrDCUV+EXkXOjPVhK6ENgwRxs3oM0biJiPOJE0zxzNmZDbq76zk
szTjgWmPnwdohtO4o7UEfv5foR5/6He8A/DJFHnfQ1wmdm4uPzMYij/FiydmgnroYBpA036m2syR
diJXOIA9I3jTY9V0rTe023aDjhY6AoXt6CXI7hxhUjIbq+1croZuytPTjmKJevyHjX+CCxHTzw/a
euoDsaKw656UR9gAPsL9nCJBwjIfPcqBc0pdBNsRDdWr9GM1tzrOLZ/WD7z01hF9J9boGU3CKspJ
5um74DM+nrKQakM/NSaAo9lZ1hH0/NanP+FAS8yr5hcEg2oO50vchAmLP2hogmZf8n9SsiG08ENz
t3fA/LgEOSI7UVFJmLP4LZangAQ3QwYEKtJbXOTew8M85rrkeCZP9uRh9HVoHP7bLl6ntINhLmSF
xdZPwqkF8M8kgqGb6Wpvttjz+H2neSfrLODwLCw+hwUYqfL71a0eag+QDfZeG0cl5o2HpI2TCeKV
f7dB7lls4PKlZw+90gKQ2wrHkbBRoOwYsIgJ9Yc++dC1cRFqItobA9iQYDv7Svy6OgvZZvUu8W95
OxkfbYdWYGM+RX8bD4oWPcqFV0Hf8stZGoJvSdrd63C+d+pO2roNJOLCW6TmhKlr8paTIX8bYc1j
pQWzpxDOcn8+FbDgkJWd2hVIqmPCRNHcC/rw/yF1amA05Hx92eGSPF6BkCrgh1ZBANjXI9ysp5s8
ejxhvmqoZ9RL0vfMLF5nLjCMTZ3ZQu89O7khgbvTic+1Yok8fPgbjXD8v+2tcNIWJ7Y9k2AKRUHK
wsjkscwzJHRjSR8me2jw1sLL3cO28tNuFWAYRcCm/RYwS9bVywMPe3DyI+FIbqrl5cutvnBWT5Y5
1fxWiH4YvxS0A8v4XO54OBC91s0sEMHEsWgdHDKbtttGRCFkg2OiOiOCBsOnda0ewxYIAzKZY4D+
iQsiNi7dZBG/1iw0ooazgnqq7/JSfEu+pzkCoMg/Vi6rVxh+ffiSaPxsp5e9KPCTqPGz9A12Pm9s
5BfNyzUWty+oXGz1zN/BkNnXXJa0huj7zBKcmw/Hg4chwXChzZvLxen7wAxj0jQhIYUxKtP6rvxb
5NwltWufcK56KZ/sl9XHpY/WFHzNFI+ZBF2zLbKW03nog1I4qvrbLHy0Btd4Qgn8vsvWJyqS5KGr
VB1xOTvRZMPuVIi428nb5rbNSvvlvO+o+4oLkuPGMgqxJjX5usmcG9unhL57gMRcK4up+Xv7HpPy
FM5btdddQQRWNE666vEHITz8Ft+QbAQDx9vLR7VpyyyUjst+SPBBe0y0cutFWnAnItabnGQ36J1K
wqy76YZP6jYKCIAUppIN/OEo1f9k4bHsEfCoAnxAmYuzqqtOZYlX9UmDrjhskXSgwkWJM1+WuGH9
ubq5P5MoP/hIw+uNipTNbLo9uOFRxBhWy5OEkwImmlG8dLOysaNsCb8E1pildNYiBLGyQEHmVDgy
i2qDr1l+uLKirGPLdxnt5QmO9zpnig0pvBXw8EtQhqmibC14L2KAI4oyAaVFHNkpuAKFBEOCY2gV
7HhY9QPdBvuiFmw/CerfJIOtfWqrpawJ3ZAUgd69D7x9dCVNZA+cdGLmElk+khcGeV4E5gccFs07
FYHv7PeiKKRuWOD9mac+1nDKoO/1w3r8S5a6UTrFYlTi2+VG03qoI5mJA7zcAmB7nqXUWc+aRtuO
oXlIyVfQGhm/dHirJujUqdmZq4qEt4YyRSi+0IVQbS5SmHM5bchIXrBuRSAaO/XX2L/O3R131tO5
rVruhQxe3dFVKZbimRR6tr0jSmxHYybHVZ0oPq1rmrIvNqUF05KMhfVstUHMZYWU+UYnqFzAKEXW
5XCR80rLe7e1owxEhLTX+4/DeqGUaUOWTc0xNSy1UJngyF32aohN1HpFs1nJ8uvvKQijws7ZVqmG
RTIVtikC12cnIi3JaO8A97bWkemDYEvMow+wTo1NT7QQMc+YOqn6Xz/GhaL44PBKnM/Wlxs6i6xX
1ECqItfSe4Zr7jAMFfexFo3ozk6ns4U/lgv5pTtV9P02vn4cLmmLFMFTK8Uezf88/dBJ01EP+75h
KVU2NsOT4T3s9TxArozn9ZY/H42RQfNFf+5+S1WEgkD+84gfqPZt7zayAK4EaCJ38blVla2L6fek
nxWh2ZbCN1HfZnbKwi3U7Po6AucKLfne+LW/46sf1X9jUGJQRRgPNeshaBMdXqaHtxA6BvXbnM6z
2tMgLqCaByw0UirFEA9et6DfvEghVom8ZgQQImBT4rxpnqlSj0EAioNRKE3j52sHQTOgve53talx
BM7My0ZsuudhWeNYWhWgbr0pQsScJ2LCxS4vSXWrTZyN8fOTaTZWFMM/AHq+JNSXsu6ygtVvWFaP
/F0t//IdtChAoEeY0ZkZi6gyHGji9Q+OBVqcHs+LCXHnA4mssd2bLiwbQEX5AbX1br0HjmhRN/0Y
k0cRoxhsibE1rXAvk6APk/kQtV7fguIkiYUZAm0SBRImaRIRYUXJzwFiETGErZzXyojF22t1U6er
VWsERzEk0A4HNmcLZlBS8+r/1/DWzJCzdOPOrpnngn3X6b0TE9SrnGiBHjK5Vt4f5X7NyJYUciKJ
R/V6HE7WaUMEMBM3HBZWktmC9uKjiXAEhRScYPM1TL3bD9cUzm4bG2sQN5fic4omZeDBopCnUM4t
UeH3kk0XnXsSw5C6i0ZjPMy9Nx450JUfwXn9Y057ewgCHxCDtX5tDymgBhUCQPjB74yPqrJWe2Qk
+98KkDZXPjQnNV8fT+0hwUU/zlU/WE9GSf7fIrStpy2mg79/7/Heq7la2zHiwKRNn8ijVxaAJgPL
zdwMuTmlLL2Q6yoNmAR8v9nllqZnePcNa/O0kn0Xay+S3+z407GqyZhsJ4n41TBN0sDLTy+4lMFM
bgpaBEm3u+VD7ri3kJpQUXqHYRfw7shxmpRfI8cc1cDaHSM2W42ZBwCiDokxzElKaRcr/acd4dR6
aa3mfGy2QLOP2Q00erVGNZkaiVKLBfhAOg6D3loQYLbLelxO4hhpQT4fLY4Bs+70G5GRiAJHA6x3
1Nvxt9Sh/IfKVuMRFkFXvai7RStbMxFm2aq3FiiyB1NUtbXDced94Oz5vCKuzSZWJsZBow3Kvr1b
ypjh7jg15LMSpmZ1H6PKBpHJe8fPsUjO7jOl3JscHdnG7/EZuzki4X7qLKlK5hKdtn21yVjKww2w
Ba8Vocl0/1ABGfiMZFMvJiWVF9oqCFjMDA7unxVdVm17fwv18CQpGPjDMEVwuieaIj7yEwnELlwa
9LOMercygh0THKsnijAiK0yGAyYRaa05DfNx2IXv9prWgS2MjHYSAcqgVFZ9BvssuC0RNxl491UL
yBEQ65L2khH/G1JbAoXsO3yhiOopj1w1aUSKxgbWMghSUl2dnS1xycVQSeXW8Qj0bM2E4TL79oIX
kienJrfqwQV5toYsTh0x7HPyz5YNJIK2JJAsoq9lVsqgtuXiMeKss8kWQBMgUu2QFQzEmZRLRX0T
3rgaRaAmdz1EEYt3ktYNgB7HG88O6J3hwKekG5ZfEMvJEWwoyaoH4ehP3xvrJz7Eyz1lFI4A0126
44Ec7ByRo9QfGRrGuKLC466VvfvK1GVosKWnntnFmnposukyA00OgQv69uTQWxOgyiDsV2afRVLB
BfuahK+7/lL9ADoOFbdZaK/KPT2twe2dkY8gEv5dumP6uX7V/uXOTt+8BN6YsO7TEFOBmQROQYio
PKjCARIqluEuClMMoju3BOuhQUnpqEcPv+03nWLp441TTBhhgJp8BUtU1TvrUDd55A89N1AIFM6p
ge2hFUJehEFwvYjHrpc7Bz79cruFmx0O3g/m9ak8ulFvDpn2oTmsCg5TTbBqMeoR9iN+i6eUjKLB
iNkQUg8gn+moRV5dBpt/VPcfFR8Thdkh4FrLexBGIO6r6KMEFPU+i1CKkW7PFDkW0mWgGV6bRY/m
5+E7iW7iRvQq+dIUZvvseLMb9lw19jH2vt/BP4+b2C9dyUu1HS36ULI3byjhHVbXGN2UKcr5K6z8
JUMmnwM7XhfC15wRXiHACC0mSxvj4Ob710uMpEXmiHnOYITiHzYSAuLVCn7FFSdkDLtBAupvB7g2
vKfg9uBPBlIYbSVyivONf2JcdoW+o1ELUqtn2Nc86QfQp/4WZG4RySbv78TvRwllO8bSYW6/twHB
WfGz2q2kC4B0G0LABUpxqokzP+zE5PywhVPeq54wnViQKWAIQpNhKOsgosBlWC3Fd+fzqgTIme07
SeQZHKLtPiK/DJ6PyngK9veDSBBHq8OPVczaBeC+zDIqBEiCHtlIiJNt2nRZ9iquuOeFiSh01xrq
qp+Uwd9UIaQ16LvoBCLoE0kSo/OHfjnQmEn/DpUuu4Wgs1SArujKf7inGLsJdybf8ZmYDnrGxXDp
mt1bC5INWb/6zXnC+sy0FE4Kkc8go6hhAQZLoqRFz2JYb2to2DfZa/oOz32guxTIcpN0xSXnPfB5
XsAGfLSlu1F/Kx+KIpCz65fLfZa9EzppOmP9uJet8/NeB+yBLgZHS/ohRjZsAbpemBtF8QhwhkXO
UkI78qx4fud0uoXKt8ZYsEUwvv6nrZVXps5pY8vrqllyokqIoeFAGgZ6wYJ3rDcjk+pfzkTSlqgB
6okwYeth5JP7uter0+BRJwWKzRdVq1to99A4DUnynCa35Tj9DZjOm9aNaOEm4ijJL/hDqcRhbIUC
NTCNq/cSZnSpF/AWWGeKWNKqR4SwHoHWs6plpHpkA8CJsYsKA5hmuoQ87pJcsy4FgmqSR1ou2OGI
IdwuMPBOxKqTejpaXdWvJq7boGxHnmRS+IITYdrttScnDedNl+u80Xgffn+OuihZ1dZX001+0T6O
F1Htb8CI/JKNudHHEt3mNmWW0Bw8Nqw0ZKJHZMAabUwxAtSsqhKBZ+qntAYHqM24uMUK9btBaE+Q
gibzfnh+lLesjwnCsml3dEdOOVtjw4sb3dsO5AAQnEZMxUqQULtblyjqZCuVY2cNPDiG22I/by1D
XQuPlV0u7KSHnKBscO+qgKHWjJwSgcwnXwbpCyR+JNTnJPeYDO7wXyjOmgGyC1iw0lS+aWgs03L4
54QcXnbw4zVAJ2gvEAsvhDcE33cVtKZiyW/Ke6p9X5AOMb3af16YPaok76soJbDK1JBTL6uGaEwv
4GS1C5OIW+hf6hjHsfdyB6YE+YNT6kNCEwLbfbl834Ayzqo0hoArcBzKfEz0fRczOi/DAi8PqH41
dwI2MvCq6fdDo94TXbdJ6tiLgvq0Ze4xMwqxkPARubvNY181lrD1RYD1+EHcDXLKAfkv5BcefNX9
M/XiYYsXa1LsaC46Afan7Nf9HE6WQt0+063PArnLBxa8/qT+SYo7Q71Qrbn7t5D85v+kgHibWNiX
LoO3Nlv8A+OKvCSLGhH05LiG+Yk8IWdTQAUDokNtE7eEN6oI7GUHbUzPg3zKbiDlhN5PhfDUpDsp
hureSn9bLDOFCdMPrlXi707z4cqx4nicBHfv4qBCbTCwLyXGJJCUzSPW2PBPB5CVf74iFDK74Les
r/phQZp5fGevy44SpwZSS/JZHGZiYmoe6QaZsPt4YMNwCbZUXzX7vb2T8cr+YyojFJ6b97WU/5bj
5DoIeniQRcYtcpYSXu33NXoKVRUxaFK+2X+JktfrmqAfNHUql1Qkh+40OuuX2RQK0kgp707Tlwtx
ohBuXMwPmevAJY2He1rsv8YfaEdBNNp7QEQeH6sQJZUQs3pLT8vVEHc16STgIKobIoqH+cwZ5ZlJ
qZIte5+nJO46RfpFe45jKeRIJ209VcYpJxyy+6OEaxnrun36q74LBUwjqZzLnItd5V2LKVaGPwWK
NuorFZMGy3xFBL6afeyhe93w+pHLUr3nQ0Oui88FQZxIpB91DL7mEB7Rb47wIUcU7IwroBHtDg5k
0Rhq9i6LmmHWE6jkV/SbvqRRqS5IYGd2bCALT9tYOpvU5KsB07tm3/9p20FF3N2bbpArmxdqlyOw
prCpslVY1qEr0WkLk9oVUE57Wg9OxxcQ79I4/GAMnOKw8nvuVaTwU8DIjU9ZvbIjA2LO+FyMpQgO
Fsv6tRnR6FsO0xYvccOnmTSzHLhZ9ytLIpLG5q+vmi9M+CQmUSzct269mwWDjU91fbXUF6CXAzfo
a00gBzR7NS5zmbCQsy7h95tcJQpUW5ucsAfMeLtDGL6i7SmfHOsLJlLCeJa2Z+c26gs7WlLyGuV8
8MuGdKyKKm13E8dLvobBKa03VBEXl/O33YZkeX/qn24yKlRMVup15FFOubN1Bro/KwFRNIJWM8jE
mbcRBL6gz2AC/AW6upLhtt7f1ENtZhMLXPK8lNISmEc1nhSpskoFYg/6VSh+RNUJeVoQIZvx5zUE
P8HPaHLVbyp+WB8Nlgjn0WJBwW3y7t7AETYCICtcBwFNZss47XwbB1UXcVqtdOb+pf/ACco5Lg0l
pEnDRRPPkK6nBAhPy4vEiJJ9p+mHRkgnLspwNA9rtni9FKELyTUmOIXTOXDNzO36ZTaGnK1wizL4
cBySGGDjBtjBOv9e1r3mWA6VoMcO/aoAGhIst2Un4tSGwcraziuYWCH+vDlADZTKewIWqC7wsZ92
PHpe9KWA7qjKDdipWEyLE/GjJpMwIRNYgl+0wQlXOJsfJYCV9pNPVgYmU78kdrK3gWXXxGZtZJxn
bSw97IjfWasdrSaTE5E2+fKMm7tbMqUw4EmR5dbppHMr8A+6WrEFI8apX4WfvKK3i6ukTAIawIze
hhPdHT9d3cgTNNOJUTi9S5G8tCksngTL6tiY9sOlr1GzHb+Jo7PoXmTQCCQkquTzjL8G1dQOEugs
MRPVWiw1Hx1tzvgS6gnzyrZCXyKMhtOncDDw020ziYAfTp4jLDATgQWc/65l4lqiHovDmK5ehXCL
kEdnzY7D+sUqME2ZVRxuDZHq4RC/j/eNCiDnlESjVBWN+mrnolEoUfM2kaR1voZIpmtmJwgY0mU1
DQExsXoFDpdeQh/tfgz3e2rrJu3DQXa0YUIdhilKLpy3+FVr5GCrLU4q1OXnBkiFSDLuNF+q1H/v
Op0p6ErDgv3/p3PSk7hnjap90Ug2nl9ZYEVR9tK6PhDH+6X2tD/MCdkxHeZEeGMMwVHlhQdPitjQ
9uCzvG/IcWAeXArRMLiLYTlsY9M0P+NpChfEn1N/Kj4YUOVomdbgs2qJaBHO1c4u+BntatE9gQzz
dbRIhh0mGXkcpmCmVGA7yDcCtQSD4Yz+nC9G2M1bceoaSHLrjanvgpvG2pDRBj7OeBioASIr8kWk
w66bCwBFTHZL940tdEoQxlN/M/Q5UDYKRZGSZSNDXuaHbbqbWOTS4fPHnQgPK/YZXlquUoUfOEJR
iWjg7X/fFF16vtwE63KdZvXVQMTq39EKcFyxalJLlFE2OXZGc8IskRGPwMquku8O0YAuorKU+s0d
4gnS2kl3ZPHhcG+k7BNcJgssvTM8kqDMqi4EJq180WtofWiyoVJZjVW5QkUM8cKzPt6R5CJz6zbp
SSARCGFzBGdCNeS+nGNH4Sivz8m6eIDmh+K8Knz7gHIqoAGQ15jckgeu37IntQZoLZzxC6eRKW7B
CSAuk8e6OmErSxphLBuKJ+U1ewxtFyxjlPwDzNWG/a706w/ETtnyEdyjwOrh6pKST7yq9TSNdzxv
vSyn1lH+jbnkJ+MAlt5/XFNn/uMsh8a/7U+dvaAR9qklO+UAA/QGYcA4HXtPrvYAVMeMULjOpF1b
nM/uoigenV+NJqE/cja0M0UIet4H29nMe6wBUVOcwxIS3LRi3KOp55HYvr5YhNg3D7OrOuwG7vCl
I3dj+b9SVk4FZUePjuZlXE9p5Cz096MaMyScPwaaHEQHNSE0BgANsxDyGpV51Ic8I3leb+uPmJPY
QJojITRfia2M+td8osCvsWvHcOPbwATP+gADilYwaCCW5SuJduXrcUmFdTtFFcUoEG7XRzdBSTgB
uyxUHwSwfQ6Qtlrejdo5r8FMPMst7SxjyKCETOgns/SK7pYTWkD6ckVhAPT8iKJhoLizUVDi3RWr
2cSjwwFgHoo/fxGGeT/FVS++fX3XXImFZdxkBWcNnt/TtcOqJY2KJy6ZkqdJk9WVSc7kk+THSwtT
cPH9GQHJ2JH1NG/LFJ9RVwnPhaT0K716ZMTH8B4mM8TokAoGiaTq5SwOH+TD2RIXf1xUGOfff03r
Ww7filcAjy6gIB+zPXAjkfDWaMOhDe/hr+bnaOI3JUt0mfJGrFJS8x0kbyBbs1OJbPdDUItxAHHc
iavTC5B0ddNwRJxR4QTrCnLm77/Ezgdbndf/mW8BOwthOpdEZf4A0L00+hLgT1the+hOrfe1mxpN
2VeBrcxyqgBmqOYn26YWIkeP58cbLPEAlknpN78gdYb6HfR42uivlcdaIlCWvgp7gbtGqBxNeZPS
tg1Cf4/u5FNj+hH37ufCrVujcqi5HU5AWH7Z6E33CScKcPMCEuNHQyb1BaZbTUVs7oKlp+mp2m/9
t6TAMkfbOrLuMSD5GRV/E7xudJqiIeS6ECGev6IWRFYPcEqXIcHwRCXcPGx4qp/yFoea8KUiV/hz
zV+8UYV7/OIQMwOucLWqsfmgKCiIq03ARtu8i6FPOOsW7Woyu1iZWBJksvCDR+o6uDWjRE3uTccL
CfrrRdRbQv/Ma72KE11oGJit9VimOoIkK1NpE6iG6Jxh/QuKKgDt/lovkHwvCyRNVMTA81i5HD8K
SRTr+bE3DBT7MDB+sOT9wwELAvXWO11XepCcJnkddeuI2cIzoITqNBAOSAdGvpU/MN4RxlI61SOF
z1mNvjFcK60XUE7mUg5cWP422BMGNhdbDP5y7yzncnFmX+EyFAXWfV0g4up9O+M1rjTPCPn4qW+S
OZx0zYXh54uEMhMSztUORejjM1U4FqX1mUgK+e00tuiZ1PiTD1XC21pukFMVkKswKvmzgzTwziN8
MvnnSJTKK6TKS96aqmmo+XPfqELwbSTy1RSzDGCQM50IUu0iLluNWjvy9VA2RUpcMDhFblm+VUgI
BNrcsEO1N9yb23JWLe8QRhhGeS8h2xrbigt7Xdpvu+Vd5ISW2AD8/9RLEE1J0Vij9lOTeiP2wrU/
imDr4Pdx5ktGIQJ6xIsLEb6l/BbU8TmehINl1tGrg76m3H3Vuth9l4nqPmakdmaqNwqteKqVTMXS
RdVfuizYAw2DPH56Le599jw0R3Tm391IwtarR7+HIC9jO2ivVXhtivO+iOY5R1RDj92StloSfIhW
8lzxoXMUrmLkAI+5UAWL30rN4devannZQTAGT5S1Dhzc2HNUZnXUwmKTbZjQXysAwIi40pZdaErV
lUyVvZgHlVcQY4LVm9p1pKSBUqXaXaIvjUPRP0F0mnNLzZnIppEw06anNhl5NabzwpBGshPc0UIf
TJnmBHoseO9xj7FiHfiYFoGY8f1foLg1Yc8aRDsqAnbwTL95q7sQKyovDsmlYuI52Zj95LMWtBCY
U/TNG2TrtsIMFFo2NriqTWevOalSlLGydcXmz9MB6wYXd3dQvZplyS5tBKJsZ5ZZHKkFEMZAQ3iL
r3DFPMut1kr414YsmmwJ5qWEA4ZoCR5fBG1AFb9LGiKWxBKvJL1f/jwIThCJeRoa6kv+2wlR2p0u
GVwddLbAMBeR9as5qdN0glODRcQQUwH0pxFGsiiZWFKKxuUV17NJidNZ4iAVmnQ7UY5UsswkQkp2
+tsZR6eFshHUnboVzcC4T6tbtUGL6JK7/0J72C29h/mkybAheHEttlblHi7rk7TPMDzYZ1Mxfto7
v956lEOlfsnLa2a4FpgAtNdVDGNolRONPFhTqeZINqxO5IFeZPgPsBKI2g9iD6h8kfD3K5Q/HdVN
7+iOpl870wjCd3b2WaVh5t0qQT8MTkcA9xh+g+NkZMQngFTRo0AVMuWsItj8FD1YCyn7CLU2Kyrp
xEZquUZiFJMQLhlVmIFip8Hted6BntZpLlV/V1l7IVwYXvYrMidzhO4VpZ/JZnzSE79Html7pBjJ
hNVPDqAxtIP72gQNsMHxDZp3/ia3bQCLPVUAB0Z0JgvBb6e7Wz8I5jy9QsUHNglj+ZVRbCNBvfAF
yP+G7+zgq+H7a162sj58/0XkiopbLfFkC8+k55SDfc4GLfD63O+o4Y6ogHewwk1JLCLmKJbXVQkY
J8MxzMnlSJoY2AJoWkH4ko4YbzTbzq6gY/uRwVdqLImP5NT552JGFgU1QomCHG133XhqViGDE0SJ
voGg+8tLmeEqFYT6xmbxHmnjt+Lgn+ririYXB0ahrjRqFyDRHuxgf6RtbnHeZ/gS3uf/59xmbsQ0
S6V/UwErn4LpGRa9LX87CMgc6ACRXcnzMAlIMxsWZXzma6Y5TA6z/KDdk4S4yEIm9ZA21kTL6uTa
i6czikFISpWwnJ0SqTg/I2tWOVDOqagKKUKZW3Fk1XVob6vsCOZvJ9PBeXSNMSa09xkkS+HNhkD+
LTI1Z+gnZgXCQwJlMI3/piOOjmjxPW1PxSRgNqUGNLYUpm9cEKaawyZdJwjsKysO2sASvOmTh849
0vGh+uTltYjtCPdjNaKy6vkc2jcUryc7e9tzZoTMPxt8mtznwfciXx2YIVRn0fPK7mjadMZgjRnk
fLV4KNnIVomwrXO2bA412bhs5G9JHFSuZZ5OmRS9xF0fIeF2y5n5fX1mmcKLBxEvn8NHK/hta1BT
g/pP3n6v4/lucvIiS3LF8sMWoQgk268utt1hNfaTNmPNNEBJwv2j93ZprdiHXfXiyH0rmbd6V+MT
W3/Seec3GFSVhw1DGd11A+Fk2YIkSBqbNRAZONYSKbdvSXM60r03kGhBha06ZytJ0BNX7f4RSwTa
Bq1LLo5FuTLisYyXenv96WDOzkkLu8jlpdZpE2Y/t8wlX5PcoQ5YAewH4XQCzegoEgDvy0erHT0d
KanYmO0/KlnJ2YzFdUraV5G3OwjkU7zxEaZLMhSo2HriYscEynzaSXDuHzHe0AHTynS0DohsJ+39
qQjnfGczKlpFs/SQo81QRRyxdrcQtJsqi7FTkUg1t2DzK5d1IhkXZ8p5RcYQnLjiml5SXM/8a3O4
h8sI6PtDcJsjQbrDlzOaNIneakuLWvLGCrXZLKUuTKRaOsapIaULChuNVDx3hIwqoP3tDYy1oZbv
asm+YI3YDUlrCF5Yo9piYgTkR4uaknxNiWfJkDlyFdTkRDSXaNK6hK6Q3mCdYxJvRmM2C1D9MmDq
HQ+NRIPfgI+QbyHX7Jup6yve7Rl7Pv5HgbxgDUofurE5U+nm18s81Z+zyophO/3xwIIksVcG6cLB
IcLSZHoRcdyVK6J4K520mhHaUXqn8zLdL5pv73rFLMhlxi9FwRKED6JbXMjJU3c6NxhzBD/us4TB
s3/ChWUaoFYlmk0wbeBkpZXmweTcEcLGN11IKmdOZ8xubOANclUuEOU7x99ZTL9z3xw+th77Exnw
NSKBpLymUsEXdvqRO/CC2DttFczNv4C9cmDUy/SU6HIscHiHRuVRFqsObUsi+HKrSkpY1KujACJB
2FUajj9du7BKnDw7KAKcpiRPy65kH6t2YDx/MUICFgnfH8B3rHzkr0qf9/JTgma1q454OtzkW+Wz
Du4bSllFhQMj9FIR0DMNMZK69webjAFuBs06Au+cdhpBYZ0++EkvKk1pAJwPjNQ5BAN7gyEK0Nd/
QgTkIGArrjNQS3wt+OfreeciFw5Ffa0x7f/mYtUbdaxvI5O/5PRaPaRSB8yS0z+DQiuL2VFd8trn
L6DD4yMeDiOuSc+9jabufpz48LTqLkpGdTtLOdhvnMa1ohfD6frl5kR8isK8ojHu4K8bZliBOpKu
BLfBvfd7vDhEhHUrbLa3YDxm0EnxiCQFD7Q2zZvLNiOcDrsndepv3o6db2vyPJ9cDBUG534eSAg1
CobkMF26ulEDA+V7iN17p3H5DFO6hcr1lMDHSwETOPoVimAlTyqJ/mXJ0GZP/wb/b6pGH5eV+H/g
jaHyzL5tMw6s4yz3DevhfbyaavivCjWz1TxLVrvhbo0mBuZ14/MHKft+hyJxAvYOtEdV1nFBoTIc
XaLze2sgBeFjZVGvZ87h3dAGjwxgL5YS6SeT+nUqfEev+kcOj5vIUXaE+32y1d6xZ/PaZjxZn+2t
d9Y7f/e9ZlEeCFMFuEM6WkYwWA5XhmyKMqmKTQVE8+Ro0Ndc27osGVA4onbBlkWpZX3l2X3SjaHJ
n4WqylTqr+VBgndrWoOObrhMbbSa9Dl79TbkTCT02FgymZuk7Mqezk8YyDqpHaDXPQgoZ+Nsjc+T
5zflhg60pm0t2IK6yBKV/8hNkikdgjN0J6DcWMxpaPCUIoZt+0tHxEtjzzK74imOJxOpgfNyyfcA
AzSJh4eBrgLL0ev4X2MMHQFzUcMc4ktQPmwG0wQqsBxq3m00kDsymdybJDp+6e7qqaZxXMFGHnhD
5lrNnQs3JHVQELkQpuhuR6LkUJu1290vv9zhymdQdNmSD1+kvqXUR7TVfWewyFYELDhG3WmjCO09
7wov0RwAiEatQ+v6UH27xSf3qTHDUg5squ/fNM8wLjexp9ClcxojwM4cNTQbcp/ojLklZYRQP6tQ
9DXIY9+AspOjOqJd5QBRsMGLea2m/SqDlJv8PjEL6RHMeyyCIbAiyD/5klkt65rIYVTux8aYLMWo
H+XW0W81xu6iEUimoC+gDLjVa1+pIFerKAuq5UROy2+WHturYHBLJFb+TDyQOPAVDuhwM/eF+hzq
n+kDVycmTUqm5PSRWmIJIpVMeX3grAnYPCvaVCi0Um8WTP8Qdo4bKSXN8MaaHzbfIL054F3eY/Kz
VpQIasxa5MzaT6hqrGwnjDqo2+eVCTLX9HqZ+Id6ECkYOFq4J0K04InYm7638qcRHgnCvLhDPBg0
sG6KaYGW5C4bNFNpaBhCoiyMgtiFFCJkljV0iL65r1iKiRNEf9R9pVr8QMu9fdblyqqg1THeyfXS
3GJVwPTT+JJq/tdBYodzk2hq2xX8XL19A8mE4EIkJ42I6LY7yvtMSuOYWCjLOXNghXJZP7AODiTA
Y9Ja4fkGWkegJKN4e9E0tsNGF7rudOTIBKS7PcpD8NZHqZ2Msb9DtfcoLKFh3AbZAZ63auRnmhXw
gY9lU1XGWsT0IIQ0224/yny/TQQRKgupB8JM/mhxFW21osZiFh/4rOkVQJgvOgy6NBhmFqsmcdRl
hMi499eGR+DoB1vZn1bII7QxwIamJuRFIsvM1+1N3gKOLxNc1e5ZmdEJOzEz69j0Eu8890itA8iZ
uFfcrq+VjSuMbQpMHrhU+uzwHuNbuuZ9E4kEDib2Rh9mziS7iFNuZKpfyD1U57sks9HmnK1DMDLG
rwjgUGjLyIEkhs79qeZV9/h2A7c6b6+Zgz5pqO+7Ef1G+gsWn2q35eK78hJptcfsi2VoOjaA4937
izkcezh59FAHBAsDn+qkVoxJoWogxxxA7+gunPvnLAHvXSSjl16hpRqnJwOHjHb08cWHXLM7fNMM
HKhS0K6j4rS8vY/DbLV33/NnNDACaUpeBq7o8F5EkGlbSTnedh2Lfg7SWWFr2KUixJYEPwgRelln
Ywe+Xb8MXI21iEn+oNpCCUzcW374zNIAl1mUzSBlGvJ3nJfV/kObA/PQjjnfhTMUkQ5t0IwVdo++
BVioRQQIEOk141i0NbK85kbq7jQq7uHaca6q1IyHebGDq8ids8u7yX0YqcR7VSqjc7smRp4mfkCV
WXEjjHNI6PWKaR0xcQiG2uGjfLDmorDLFFKpsAWmLRBAGtNpfCcw+FTEb1KbOo1rx1XUoGvRkXxY
Y9ITHRambCSaMELPND4DQsApfJPSLcZIoDuWVpRolq690oOL6YMFU6fAcL6Qzvpuz9OBVGmLhtH6
5Y1KKBG0D/Qc5w1vhBNh0zii8kH1BO6305fnVfqGkddU++4YT1JuUZjXR+cNlCRoogFWSnzeeVc5
SEK2ZycFRNIWFsT3VF9SD4ZRduJ6gpzrQlL6N95LsAohyn5uGN7FJFlNC9lyDvCoBiZfG1Tit9KJ
BHDy6kiRruyxo0OPtmz4C33ZN8d0iZmT34IG6XqCMmV+I0UM1/Kf6zQETgfdrA4uUshgB3UMiAP/
pMq6y63meyWT81hM4Uzckb+FwSFduP96/7x7ZcOKmyaOtijmoxNr6/jwEUEvIWZYWjhIsD+ge4iY
KAdoswuILPkAJiFcT02yqD4HVdW5uxd4zXsILZfxtsYflrWK4gKrkCx1XR+FabHyQ81+Jjgk+rrl
2vLWKz5Bkax1mtPOkHZadWzhlhG7/PSjn5N4CpTPi6lOvBmcGp/rlbvP3ddP6Jn/uH7joEnu2STT
1DAjkOn9flLwXf8yH3RHl27QocE2wq0gpLXD2DAExya9ADxy8Y4UKSinqwEtBdeqRmbVWRZ4+e1M
2386EyNp0KoKQhnsqXM/UIFRuZpkl3EP+T5/CnWoLFAj5Lj2oOlqokzEDvhNOP2hlox5m65eDula
14Wxzm34LdLPvyDrWllJ2JNEUIUmajCUbNCe7uv7xeaPu5COUio46H3iouf1RZI3pwH2rqzVGYrN
Kl95IICbETi8bogWPxb/19XEQOvj6uj9BDvsPHsZLG0t0eIFVbv1BgfFbaUf4qjJ9G+zM4k+zaxO
JaUbXYviqkZLTE3BmFmASJ9UXK6zRIOEpT/eDemNWzJL8vH37yeUeYRFFfDwgT2gWgyFufOkZGLa
q/0NrDh4eUjjUb0hLh8gIr/WqwlZFfPFqLoduqZSURZsBRye4/91y+yL6SLhDPZV9vzK9ufZUbg+
Yctt+WL/GpeIWxZ0cvHN4yDJjGPTn0S3HPPQT6+A9zbQo+FEGFdIKpT3/GkLvSU6cw1BMWMnAifJ
aAzfE0lAYbHBZp6D5Lv6+qZ437SihS9FQWv6TLZ4jk5XdfMnZ7zFIjf9LA11AiZPxF9xB+AardGu
skdV6idylK4B0onsy0/WwpP8dbmQf4y6mtn91XXtyfMguqibraXcmme2WZ6kr5abLx//a+KNBbvK
qmLbU8jjfEL7iKNB4urfYMUjm+9uV0rrp3hPMh20h7mb+d21T9TiuCE/c7IsK5OctqbY+UWGuJKq
XKL90NlM9b5wbyXq9w3EQXm8/Bb47USYeyYzWnCtHyHuuMjUGN+7DwA/g7HItB5ohtKf0761UVTO
52TjCUI49YVvmjb9T/cM3Mb7KwihpDDR3uP3dfKfAHf5CtmbxpLImLeLTcVYgDuidlBl+kg8jnwH
LKZiEfAsypQMqtX1Klb7KI4tNkzlai/8LK13jGS7Bh4nPGLzBIgpl7tOcJb+eIxLxPxyQS4vferP
rkvR4AdAqwFpUzs0S58o7YGixU/v82ATnhrI4rbAS3aquCR1mjYiwku6og6UX0x9Rgd4FsbOcLYo
/JsbLP+UAuhsbvWbsAcf4sAskcRghIYMGlmSvq89rmUNVd9kv18maXW/wEnmf2hBFGfnzOxRFqcD
SxlggiiYLP3q0cMimGG3TKcEe4CCzECvXAj2nVM0eOHt33sK/yANdshAAa8V0CvpgDG2XbXvxcqa
O9S2uoVIYsVedmN8+09PVyKQURXvNBdRBhIi7cUTeoqg4O7MGMoPkjX1Arr7E1zoYoEgHVHOZESj
IEaxJrRacAKrTUcVPrris0J+vGfHJVuAkHyURyzKbM//ztNuzlSfdEyUxcNs0LBoomwySGh76fJJ
aUk9Xc+ayYr3izL6hvCt50FfwBsDnQ9gywUpfVD0pE8umH5qAGv7QthmQT13XxgkhehUjEHG7Yzy
DI6SnLG7qs2Je7OfCD9mI7kZJlGzaVSd7uRfvcg7k4mIY8Ps2gyD30QU1x9tK8hEPa6m+BNDfvXZ
opWEMj23MfSnEDUHDVdLcewjzxhpNFZXu1IIZyxc1IIU9hzNW/8LlyVfxxriRncR/eFYpMsrUL7p
Ad/Kg2Cbkin6VrSAaPpmr27rYvZPljLpJKlPykvj3KZMQMqyFyaC9FoeO5YIVJoSPKzmMHuS3Ruw
XVdXWPsL0zE8pnnrd8TgW2S773WpKxjGeaa2FQd37IwoatB69q/zAAq8SLCaKhh74wQsEZfqznsX
PFg6pwS+D03teIjsIY0v2BCjRJ6fHmT9ui6E8qccXz1t+/xmUjpp7obvO/MplnO1lnJlHODTvujz
yq0j8MRHB1xmiUTXJ64oQnHHWrDl8v1rF+bhMRgtAlBo6zQ7U0NF88H4g8fV3Vakb4R6MJGHsXLO
0SaPpImej9qoneQI+G6T55DrUyV6Obi4nwNNS0r52sT2G9pBkQjrKmzF25S03sO7+gLmRVI2BYXz
S0zDU+A+t3MTmmwbJ9wy+yARmcE2CHvb2VXh3TcRsV/A22QvEYxitypPPdq61UeuMjr7ckkTJ+eK
F3i+D65C+X3PhTOktBnPCiH3fU2JR2u4/0MYCG+8B6bERT3fBn4kDYGet0UGT78Bj1cS1kTz3S2r
DDlrm4sMVv5+/y2370nOTbpRVQivnI1Te7iiG9ktsBAkj9CJ/NY9wVLsBAHefHYoylzRuhkw1bS4
8uSGqxECsoGW+QsjFGz5Xm5l7txwdu5XQ8FOh/8ZKN80COoOz5zqWub6m0XamHlfq2KK2RXnVTw9
gMsc8Wlduq+LQvdBi0zwDke8EnT4SuFZKZ8jkKH3q3AAR1baGF5o1okayC93m3Ci0bHBqVSWWYNl
oeYH/olO2uUJmIAJWE68lP86oVPf5XgB2NzMKcfNA0RuHnmidRTS7d4oJ338Sqp3TQ8zW9lCTH/0
nVfAwyZqrX93E6uZARMyv71L/ONWfvE74oLunZFy+3DjuyzSpf1ETFxt6seh8hGNoE4c9w7gQPrZ
C/h0AH6NI2jGaXEr3KqEZzKviWCOkUC0hhiIlBbaJjZPgNwvSwJaoWdhrGt0F++LRSRJuT4RoixB
f1CejCSEsee2jsppBJ7n2sVMXf/fvC5Zek1G2RiZkm6uZNnMvPTFIcn/tDrGo0pUS2RsObFyGr8V
MJVdwe4kmDlqc8dCcFZpw0aZXP4fFzQ1YCrzym588mXzOzPmrAN94K3MDpRPi3XB1yYL332BPIvz
vGEEYnW2ZjlUf/SrgBofZIHeZ7I27ynDAxMix6iLYhUNlZJO1SiaBYMa793j3h5dFy947iWhslIO
FK7eayKRZPqT3/kzQJCeRYwCXJPqu28VhPwD4kw6k2B98JwpOmtd+tTXBKfo9N/fjGqTE5erDETO
Jz189DhdhlGizcpQF/eIRTtHAwewm+LCgaOZn90A98JHP9xeFNnz8qLoCx9L5gAvtUZY0Klx0SpJ
1x4l/bgAAc4a7R4rWp2nmY9eL5yRmESTrZTu/KgeO54W8g6EBdaZcLSke9bHOhb6g3G+domxkym0
no+v5QF03zgerN9uaUNszBBnRSkTUxiPTwiknbdQUJsCYmF8eNdgAetHGeWOJ9/kIVVbKyZ3zB7k
Ay8sj4KPI7rcncS0HB7qJ4nFYemZO6zqNR4JueUCfMm91sSBoV3ZOUSmkrkbaCJC8e7gOK0SXEem
NTZJmvA/uR5TdrI9C8O0A35M/9f1uVE0M2hAJ1KkC7ZOJ8xcthpD0nxAj74y7ejy3L8n95F5Hwdz
JggnQ4urWMLq8b8cbECse2DJIw4GNcZH3bGjFvzj0atW0KYfWZP/F++cOQjaY2FTRKxmcdaQIqrF
1uyiTCm0UmExL56KZAg20l4w4F/i1RpGJXSe5kfQ3IJ1ECmmr8PnkSYIlPdNtyt6OLuBhXSHFlZD
7EI8cbhMU/gujl5dl1bWaKtF9nhW2LgzuKAjisFY11mtssDQ90Gpotq94tJkawoaEyfgI7zrIfcy
yTmdXQ/8xkQWtDpOSO1RqMIcSzvfqx9Rh/yrVAELbOpxruXz8YUf8LIWzzC94QXc2ZVvilB7Qzk+
/OHBroagLylomoDkG6LSzX6iJzXY0Py7exgNUFq0qLpLu7UbzLMqIfrtSDDchnwGkZHcq4zEYD9j
DyiugQqgXZCnuslbrft1sHgK47dXapXTd0uQLcICoIv/97KWGYfMWsrQM5XOegsDK0+CN26H7kEn
hJ056HTnCBmWzom3+4PYtzh5F4+ElZrOy28Be90XovnKHcG9sqGtXNWFI6dz2pPwSZFo2a2Qpzsl
UN/HObFAvfvEljTZO/Z4bO3/tTFcBx1lIcKUwyx+bJ6nxy+s8REYYXWQgnSY5loTnqo03xRdYPNm
5bIr02wTrjyIK8dq5haHaY2EA0m5BHdl294c5qxlhAyvG3ggrBex2Job2DjV9GOhTiDiTx4eoZ7K
fctw51AQtEQUB9kepSWgIV/72/gcduJtO7zUcEBbJmy8I+RbwQ7Q65p6jEK8NdFkxU50sFHsCCll
9IpQchrLnj7K8vzq6xiaipghFHu+Yhzr/r/z3tVOqY7WGDYcM8hQSfOEr9FtMX7RWJWafnvkLPO4
PDT7N7L3dzeUcJhBETCkysQ5kvSxMLvi977thGjzuVKyxwsg+OJh7u62GIGGxp6+eOh/Ext59EVJ
bK0zCGnx4YBUVTR1la8MeedvFrMEgng8vN5rlsD7hE4BJxmjAvv9/oJyA3Ez1UzYGnvjbCoGZ/W2
Bq7bVQWzeFu+09lwNRh4QYm9j/8xnBv2K8IqPGnvqq9D2S5HmKNW+rXZwR9aLC+RLKhpemWhZHnJ
e/Yp+t5cwmacDGynfknHrzxUhYEELaKgJ26xTaIIvlqziMpipo1HDoQyCZT29KRlDbMVa7tTiB9r
DfVA22QJ8IOfGd9Rc2howRml3beF5XngQCmK8Hr+Y7mT4dW/LNYt9mtHWUuWpOgbXbesoZspLhjt
d7NaGmsYoeSZiD97SbmEuU9ZzczbR7pdrVsL59Wknu4M9CFakIObVRmPIJIWWt7LrFbVm3rxO16T
H9k6sHgG4HHpAo5m1kiqOIAWGS3yU5B1o5Lz7JrHy4TypVgOBknWCthoT+5P8tGI/jjFmsmq0Y2+
I7u3ibYykWGByRx0Qabxt5MO7w1S9/yMOA2CgDLq8vZM5eaUV02A8cij8zxTlm1nm5jALyrFBn+2
SCpEH/6wDk7V7oYPqD94rxV6C8PzEe7lySAibJNhL5oRBerrDtrmDWmG/aj/vrKv20sYalp5A1Gv
5qLyaNPezmEJs+5z6enq990CL5z4UI0MMQ5Z5JTBks+eJN3dxSiJRRxfO9zIT8WYQHaGNqCAIdyD
Dlv0a+rbQ/T2uMPtcynRmiYzpwK8YnkBB/FdsQkDc6zC5aB1im3wautEx8ixI+K+UaPwB0mzMHv2
PlFai/3cOiBMTxi7HXF6rzyI6Iin0s0TN6BFg6DcH+5EHGsIWQe0hQiEnPfpJ2TlzdeMmIZMU85B
OQlGvmlVFPTVOF1IA3xX27ZWUw8L9ZAwqEOd7Yhv9bzIVG9KIVdrgP8N5JtB2ovNZjpiPwE9tTca
1MoXvVcg/ZEbbmqV9qoKL9Pno00XEejBiR3x8r9/H+YceQWb+jmRLK7D86eQ4vX+DBTWPHR93SUe
IvM/NkyMWC0QLGLwvV9ltGkSBXiQ6Pzj+DKeREtq3KhiVlSRfTqAUl+8q76sW86lk3Q2dSS4yUdo
SjORkwhUwizIr3jp1ig3vPU1Q9PbGGxxdeX/0hpVpvZTCeDoSIRMS6YbbRfTTbXU3ZoGRa0oaGzA
wDi2Rbe5bciRJymo/eEuiGehlOLDOZxknYSUoXFTZNNrYu8MqMV+NzQGTuu5nrdKT2YC7xnfMCwm
yZlgmKxI+7065gRxqrd6lGrLdiltozdrnppzVcAjPYKOJkJnni8NhRCJBXIv+Yz7dmtG/lZmJTk3
02CRFvweI8PLWGoSOcTw62R5tY/P4dk7iGQV+SJyK1FRU1WsnEKUit99Nhn+1tn2Hlqgo4odnMDz
Q1SKtuksik52oP0dFuscSr9skxDR+wyIxr0kliSGa3uZUbTj3xksaJyI3s7Zl9zNrWp0S7O1aUUp
ao0Q7JmgsB+IakzASWA7sQfV3iNGoImb6/fF2yV5C6q+w+4qDYzQOuvQyYHNeUE80+vEPk01FBQc
eRM5eppIoX7aTYWXg6YfBAwCFMzt+gWrWigNPlGXn1u2ftKVTELJj7QCsxsWJCXHEQSCR+IFSvmL
K7Btp4MgH01twxNwNg/TB6VLB8ENYfsKoY/ZLtZZ0v09TZjqbie9vDcxTyi8wAMiKE0mbtzZWAg9
zRxeVlq4Bd6tZTtc7EXTER9zdu6dxqEr1fmWUJt53tAl0HUregVzkn/2BuVH5hImP+VLGPbf3Pwf
f/ITPPqLd7vE8gONQoChnRSTw9u6M5wDiyN7fXZPyoT26Ke3LJv59ajNMs0YLq89/TSmyxWyf83k
HgBrmBefbOGCqu0PWBB1L1DAJekpDxJ3WzYkxsHIuO0VslfhEeU9hihfj+Dcn5CztWLJBnPqJtef
XUikJGWtKN/IhSUREG4I6CkxcQoUQ022oEcxDtahYlZawb6xV+2irTx+Saotb+V/L7ToXvOBtbJD
8W5UjjU8KIQzhqWiQ1ZYr03e1ZnZLeHukaUKg4j5vNLRgiS1mzlahH6pHg8mAToFBKeYQE4hBY0A
FnhDvZqxWwuTSHcTw6HnZdctDmLT5MawQLSTZXPlZm2pZZAFbsZXermcuXuV3L1XhdQx8bsIjA2n
IV3gE656npqWUGrVdCHpKl8pxNyUmAyUEgHNqnzHBgsMleUhEFVNYI3RNGGqASMLJQgyEMzZ41Np
d8GzXVVWN93yYupN9vItfZMjBXj0hKwlnFM91tqVKYFEn9wGTHo5Ogdy37OkAzsmCA1jZZ1UROae
nScJZQMGqfKDdguxOgldt04jxEIeG6rVBcS6Nu4sw+p8J7KnsZ0yTUTIA/WHYWhUUawCWILOk+vN
LP4OVFSv0QiTGNVoR2zjcw0Fc/E6wVZpoofyPS6bUbAI3ME48sH/zbz7ud8aYFi2fRIxsBzZ8i0u
vo7HrnQifa6VigXfkvqw8Six3P6xCIY69RfFiLDA2C2OvVnLsvZBB7WmC3uyqwI9LuAp6nxjGsqr
jCzf4KnABluH/KIYDF83+2ee8RG30ZbUvxU6RJI6cHWBPpcE6nWU772ihN04+jhezcctp35Jj5FE
lYw9390JHDeLtZneLpupJ1q6bgNqdtgkypYNXm0biBro8+kV0qgWQpxLqyvyrG1oDJNT1jTxu+w/
ca7mNK9d19KLaTdk0d4WDBO3of4BFEcXsjoEM9LG1Ix6X34UXKQ960V1k3IApb6SBzWkA2j1V57M
WbvbUe/iL5uQ35XOa3EbfrDzSIIfB1n3b9j2cMGG7l51fYcVhyFS27CaOjxEWK4MimsTK4EqWC+x
oKoKy8m8fJB0QEsS9DcpmjT1g0/aA9cc+c7x6n+XngN50DwrQhkh+PWsGZabvsXXNbCv5L0X1oMW
eU/a0uvLTj8zDRkmuWorQ1i3WkLznC6yDDbxkQN/UR+PZUX/Hqet2O4XNc6rfUqH5hBZHn7BDPBn
9m8wGlxQ6llfY9yqojxxbqH5yyC2rMWWZFLJZVavB13oOS8Y6CaZ5VXXZLzG0fJgzFwd37ECUNJq
hTU5kUIlrJCiX9uuTbCuQ6z4UrqXK0hEF31aEAVz3wtSKpmGnZ0YLaPi75E6oLUsvcAE3S5QwUn5
o76WslFah+QfFDFkmjRY2t1yVWDIHwIGk59/NaY8sQTwwof8SjGlqogvDN7N6oP/ZU2oYhRFR6M0
AokSywZmq3ItJL6iUCPDGaIwk2+Any2Buhljm/CpfPQ5eyAwcrXYRLv2dLqYXhyFmQp5JbrFgPbK
etEvEKEAtWgPxlLuj+GHlWm3pqS579pjGkqfOrHf18bJDOzKJV/OLbjJCWbJxlI7cSDpPLDYCJ7N
H0bcgsu0Hd0I3NoWPPemQc9yxZ9co/oncCTknyxu0U/we8RGC5a1tnvYAww4wq0YGIeSbxiNr3oO
q7jiXme8YqA/sdoD/pcxAkXwmEZxFluvMFkSYrgWBqXsNEvHpFEIlSB/VSkBlymEnARhKBvCMvnz
SgFHDM2FuUSUGqadww6m5+CN9AICVXxVyTYM5c42CrPS/9r0vepbxHJBzV7XayRfY8ExtxRtpMnI
zhv0WFsPvbh0ZWBX99awwV/pMVQkuRnnvZvunyL+D8YPS2CIc5AwKbRJeSkcJiniXtG/ud5gpuXm
T+nTIv4N8ukuQUQxeNNpJRuCoKrWbLxDGeFcGK/M2yp2Z1MLf+TmT8MTEn7Wp+ROnq9Fo+c1hyoc
NPu4n6oqNQGv4Pf+9ToXzWYd1+ucSAjTyUdBbqDn8p9+n3vbwlExDWCJ+UvNg0Z7MJKCdVUepiQJ
XpRSKgrkWqKJdeSfSZm4OBL/Xs1MNUGA2sPGSCek3Q0sYOP9IOb5wTmp0Sju4pWpeix2OJKfidBx
bzEQ2rUk9/5ka0dcyoo+gh0Ghwl7MXHBmW57Xz/JPcuZAUCFkwCOv/f87WKmqMVPXTC3KUfaNi0j
dEyRslRZX1I2J+JasHNQRqu61dmvh3PdmhSa8Sz5FslKQ1m5NwH1GMwZw1YDr6TtbfzVnnlnpTph
NTwAmnV5yydXYE8dFmCE9h1qALoG9KLFkPSGWhHQ+4LKXOl/5RyWJVZYfbTZccnDxH5YhrVlTJwF
1ZPALVUHO3Pkp/g3oe/7fLQ03UTO8myO9TfjypuAZGpsSkQqfFlu6iYEA8UQPecO7M9t5jdp79mD
rqHCCgRbSBCuqC8HWFp9PXtOAFyZ84WHG6FINOzMNpaVTq/8+agLyZcZtbt4Ut1OeYp61gAVvDd9
sSsaVUwmoLkyZ5fHW54Al65D7JzcDBWxPZ6EIgvFpf+xuJcraF0tB0hDkb1tQtfRA7jNSaGhFsMH
VANF8OUefBajQYFxOcqoV1QyfVwCmSh888tpf1ka1ylxEbJxaHlJVsloNwruZM71OEtBBXW4JFUM
QojclIzhlc7REMFbMOZ4fIu12pP90vJA3RbjmJ7uCEF6sJkA/E5V6ZNMl99qfGumqSnWF0ckoBx2
atJCcI/H8JdjvfVB8Cs++ywUjT3HPRJlo2zU/P+p2KTE4+iKKnDbRuCyLW/+llt1x+8AA5nTlzOs
GF7/g8R1hEbcEc34qKDuW0IcEopG8qVHULdquBZxjvITY5dmyZpE4aktmk4DmOGSr3+gPAQ+LS8k
7xV7hRt9AaNuL7gjuq8+CdYDsQi8hr/U8kElfhreZKrDR2u4Qj7VI20NkXpkdtBkoh+d1WsN+UnP
00Gcj2cyhsBVFAxKkyqYxgfuXjiJ5SJ+wtBtsCVibgA46NAOyLb1VH0hMepp7ZBLA1XL1BNwfiNE
f+yA3f4owuNGA0cj6Dmbzx6K9AEUacROh25KSHXE/+jwkBSTiXFx6ysTJKbXAyxDw5iiy5JH1gV5
I9kjUrro3sIOfk5Ffk5PGRIlH1KqrvkBdeU7VaIcTJgf3LH15Ap3qsM2/Ss9mMRWKqDE9/3ObHua
gfzUl94sOqpBo5p4EZHZ8EdOSItnIEJi4qv+PQLrCbJeRBZK27aOEYI4drI0NKFsa5q01Z4Uk5jy
fE3cMJR2XMyHRCmgdWkOVIDYF/a2Nq2mBuziFQv9glm/l2TmEDcX6zjz6ApNmbM/2cpPzzbYSh65
mEnyZe0E72nMovZMlM0NYdZkOq47+SdbXdLSQ6lo+FFNPtqoT326nF/r/KybZhYkGUAuCU3P53fz
bKf4j/u9xWIfHN29s+TRP74tS8Kpk+wtCfMtXcCL/3uSMOlKVvhg5xezprB59DtzlBTxqCtm2jpe
Nz+lrztTc+RVHOXHPfs0g9maVESihEXdo5Lx7J7+U8yaZDv5BvglsQM2KlCn0MPzku9JtUfNp/+M
0YYTKoXc9Kt6Rlpp2FL2gGHtMAKmkuSFiGCfodUJDM2EOGLDa79PVQLp8c0nikst/eKC0FjnZtqH
goQ/bLTFP64VNQSzE4J57OYgcBxiNVJjJPzFlckFRB0v4+l4yy3Jo65LqzrZG29nQqqkzEtBIjtI
UbMFnKCDkEIplP+KbZgDzFVWJHyHNyo23QWgPbxvNPBidWH7QjwDEkvi+o6FnFBwn1CyD1AsJmRa
5qDfBCY1kvziyh6KzQMfWDJfknN+2OkDtWJJTOVbdVu0QyOsgc/xqQ7BRbSrtR9lBoe1PeQ5yF9y
2sarXCaCq1WSoLSwYPOVo5h2D47lYB88w+d9Dto2jtsupWAKZDT0lk0BIbIaeH5emuJN8qvPX5vd
wPN5zQOjx2M4WrGCZ+Aa3dqYPilM92wHfHhdbUymn5QAHgUa4P3W+UY7+gIMaWpl9eRCS9LOgzKq
kpuumNbT31/tnYGKC/kaXZxQ4pmwzREjzqaQOH/Sz+2R3IKDhURaMm34uRd6JKMD+yXPHEhGfrYZ
MtDB5jvAFpz+WkiOGcj88jPBwE0re21wKHitbfrm1DQ+dVPLSlChtJyJrPD5+Ofb/nEdaSxHlkEy
J99Q4LAz7qJzQVqX4n7Lvg7l5xnfdtX5PT3nxmPhpvnrpsq5F5bJ1LhzRrpG5k4bAYdcYNVrKz5j
SSYpHwjmygoFYHu4WU5dzTSmTq/0m6G8qR8GImFnsQ19z4eGXYLLqo1jBsnNU5g4GUcgc/GwLeft
kWFuTjzRilfvWCkk4rvvWR/Ij7c7RZSEZgEfDxu6fgrODnaZaBNl/Kb+6eIC1bGiwB8OApq2RlMO
+ijZWKvAuDqiqg7BzNON3wLYqro0kSiK4NWr/HjTJsLMD8kGE2EuvolP7G9QLaixqUNjGHAs/3SA
ZFCgX8WFPDynCwGcBUZyxbMfBFOjAH6d5uEzZv8OxBKTDgLUcheVx01KDIqrPGiT/VaDilddpYNg
a3H70jvhW3xSEv7fgapZ4RtI2oL2HYksYgQsjsq0ZgUk7pfdo0iMYl6fq8IlfbYuATJbAge+DefV
eWFxBUjYmvI6PBx08tcUZ4+eg+ePHLBr0Ohrwp0UfEP22vANL3qLIAHma8rhbS/98iDB6rgI6fOW
qyxo+KtkWhPyAZuT/Bod+QfxJ0mFMYY856/GlA9RfKH1Lyy2VftUNLUYVtF5+UPlKKMiA6W5KVBs
M9fmzrnw+DvcpSkXO3s3y0x2/WYSrnByo+K0EHySMP3MkVaWpTVyJ4L7uXxQqDoJXwV5nPHGPTHs
jJSGz0E2/RaxZfn/vpHDVsdIIiTA57XlaS3Mkv/EqyPo142agCvnow7TX3/fmNjVIWeMwv6fPBfH
8qSSZRnA+7LpkzsEOucK35zSD3KPEkgaGAAmVMR8qjF36WXUM8o4zpIsg7amWLEilXYgKR6+L+yj
mJH7kn6AVP9qGBWEYml4pnjsl79WQH1gj9P3Mwp48FEGZmpV/znxGZSOSWtB3rtf4LSfSwld0F6M
WkU8AyNj+g178S8o+EQT0I/kHbuAZMjAGAdUGJRy31R1JQvi2IVPZUYCWEnqsuC+pJK0fYkcD+be
ogtbTFTHfo3eg3U2I5aZwRW91AK6jZAdx/VuLJeZDctnUtFzgcN3N5wQUEE5LrvGDOITilUR/jXd
oZmrsE8bCEqBbfeMK+LB4O9DPlvB4SbC7E+b7FmE2YVbRmnce6U+0UFSh3qvhMwrrSqYID8w99B2
uvB12d1Ety+idxax5VygtyIm/oAR/rb44IH4OZM/bbQkZmnTTiDDxbU1r1aptRBqyfGA47gdBPTt
7Ou8SKBUh1uepAhF0DCj7NkU2LqcNbcClaquJC6r/AazjzGlFDVOtIVY2p15ph8Ae9PlQ8kys6Kt
K9IrHxBM7G5yEl838l99ETnfomCiWsKcQPu0VdpaI0FAI0QRgZyyuHGb5G8dU9YH0n2raHcmfxrS
MY3209/ClCa1zgVIoWYV2mkg1lYvUvjlPMPHT6WaMWlQpnz6dTOmNdp+jd/9Byk3hjKXKg9guBve
qJ2Bt/mSbA0mtGqWf62wu7Gqj5tnwUvDYVOkqPPt8e+4DILhTQ7p0OZzQic3jHAIhgmUxRRXXvrn
yO5+89ZkIiMHCdFJ6OuLw3IXveRczr8VmltoomNAp/dB1Hsohol2X0iwQqTPJozxoXre+D5SC7ZX
VTnMu3OR5ZGRkg6Yew8Tgw4W6pev8Agylpgd3XiItyH3oy4gJfFXirxncnf97rKv3sd/Mjr0AxeI
e7/pFw572e4x0hS9F19V3WjBQopLR7ScauT9hAFrj+CFN9ewFVNRbz2l0Pbi6qUTQvNIBxA4DnXi
aC0t6qhj+SFynlFh6VN3YDwBbcbS5JPcHA19OrcQzj96B+RW1jiQI+Zb/AbogGdCzaTl0QPW2ufo
hM1fRmie1Pn5nJoaT3Hfir4f+YbIS3qpazJFQRGdCqZUT/Ve6Vt91+BW+8YVwXkpXGtdHiCdrUVn
wVhOcNCI1riKIiNOxyuGlIjqr5U6+s8seyIKXDXUgLdeXtsPV2JJRBMhu/C44tjst/A49U4oFHqh
DUIfDoFswaN+zPaeg658XoqjcH75hCGvpiK6mfQe5faD29Lq6Wxam0V6fTRT21j4M4TsbQ0mQVgE
v+PO/Eo32YA5Js2OZnssNX/tEftuOWeBdefc6QakFCaR4oF1wI32Ivb0/j8oZ8RVxBivkOqsX3sB
X+3fSTIbnYYQOV6NdPYqImh2QrM7tn4fgY/CuK0aJHFBtpDHMZgBaAu8nUdiqc9V2tI7dQReJcn2
f/NlwDpFBXXKhMao2DDItHnxcF+rpHVVPYtuH0/iu4/E9gYJe6K/6tQXenCxH/fee2Piziftu2Ni
fHY9NWtvTmNSRGy5DfF8W8MaQG5wS76f2ZCkUKVCUvNeyZw2T6AGZAV1olWuZ1OQcBuJUFpRxsX+
oc5uI8mwLdGpgc6uQrB8dkUiCA6490f6dvZBMSHXOvFEptAVlXocdnyDPkXBugEkelqNUXlkhh/q
N8+LNGz6+0bASJaSVsaRA/739h43jEmJu14L3nLjHSxQllQfaBBXJTSbnAZH08buT4eckQFwV7vw
ebO+PixjpWB2hK7Cyk88eqBDLAYGGkpwEeL8bLIgGdp2BieQMW61PAF09Nas/5z/eAeHmFixSyjj
D9yEzFVm5BgstwBnSe/m0t8Oing6JpfPeGLyIJWN6GD+PstmT10rMyirAfCumjGfXHn2suTtXswV
IeLrSFwYi2sbxtlIxo4GYm6XZuKa24EXr8mQrMlxeuQzVnBwVn9EFHI5Ds8sW3sAjDLvvewY2geB
xyfkhpSGqamAiXKYnnKPrRo/R4sjGGUbs4djDFi5cpCfb4qx1oPxhFJjWztCvJ8tR+BwrtiTFjc7
yZJzHVHqTBmqStMYqCK/rTeP+4p16U+duM/7uVEQsh1dPRZO2LMWbjborCUOmbWpYYL7VZkKjFdZ
uCXDijPO38mINCNz8LXZ+a8Z6mk3jgbzGN2I0lFZcGcB6I5lNNIHu11xcW1QqpT8muAOecV69gBv
vz5bAiT9LTFU2ttuFDLsgqc/bUNOtq4dTmRzX0MwD45k5rDv8Ek7DewBXF85R2Uz+WYFBT/PkRRX
Xcb2ZXocBoPviyTLrdOAl5mff3BVIGRmRyubm7Q/wL0FvZGVetOh48Sk/GPjiQRe/jKAMQ5MdJBf
L/iNtdDObdVu0oMvrtUwKIS/5ZvgEAhcG2EfrW2st5PgAlTQ7nZ/45WhM07AjB9Qd/0aKxGQxsIT
BKujHwU4OSSLKdAWoXMxOdX7numdeUYaZE8lQucxYNWWmRu4cXe7r0Lg6wUhfGnTSoU3vrZI1QjY
xcvTEXXDbJKOIm4FSt1tFDYEXZdpZ3tOUx2WTEqZmxunaLB6o0qqZxGCXSkDpkukt/Zip0xoAxI2
rru5gKsjwJPBo7Jv14OI2lTnj3b44btsIO9V3DepmHmZ+ArJhanmGvZkaPHMZRHbppI5KeLo2YEp
QBEZXItIZEyYGj1sEM0WFuJAq2NphjCMxFRvPrqjmiUNhfwg5ytxp53vS0B7d4YvQ/BdNmPTEntn
DBUW3HMnlCbeboStMvqDBVuGrCu89AipaaLMPDTE6G4n7R39/0Z5akRyvv8bfj1rcxR+fjlq5r7Z
llRq1xLJ+xtiMOOfTW2pEWpd7yZzXeEuPszJd/nV7gLSWV2YI0NgPwjIxV6F2hkLuYm1jz+UuT9Q
UkIuEWbyeZu3qMYvt+StcJ6qWTUUTDfZgLtjEOSln+iwiQnghuIUckP4TrfLxP1D6ikZtvMAeylF
p4WNE9fFHr+Axjk31Fmk5E4Te3UJSO7HPunpiu8/AN8bDjaWStT+LMdwvvDvDSV2vEPaRKDM6okV
jckovAiTyd5ZH3fCgzWIv3GXDMoG9bWrtxzTW0xL2ntqiNu6mJ8Zn00q+5iQ6t++/HFHhuCF+get
QrFB9nMbJnVSVQWGHXvMYAAk+VXotcFInUetL6ggV7O0MzjDmeJQWhsB6ebBV7E5U16SUMaGyJw2
85MFCKMsa/NUuiWDPvqCiP70+UCRwDolA8XRU8oWPQhf7ufKN4IBm0TiAVVamYztoqksYobtyjxo
gi8UkDpT44jLmgFHRnwQVFe8+B8eY4hKRNGHPnU0vsDNovP16o/Mse7ARhIulahH4dTf+2FOwr5y
eGad1hLK9B4V4Y76j2CV/POXaAguZYx8+W5DIOBVMy/TRBryAGAWnjUvxG90GODezJijwpVl0/Ov
4w63tz5wbG/bodm1CuIZ3rWs7Iszh/q5slvskw6sSlMgZ+l+IQGR52WC01DGEq/tENeU1Cd9bcqb
Bu5+phLVCMCHdubmvIOqqWOUeJ3KQrI2f5uibdU/rm/xMk4Xp3QNx17yK/BCm67GyCJXaHUw5mSr
p6KdxhW5AkunCnua3JvCz2fb4FrbUXNmFZgC109Bv/pav4foVk0pYynTR46XNGsBvs/00bHgyI71
/m+M5yCbfjP9W+pLKGQbDyCDdC+EvbysLrycfHBY8dc4ejvtRNOJc25Y1ljQD2LDER8Gg+xW8dz6
SHEa5ZM2LNQXP2ZO76t82EiuhtyKFZHNnegWqnOtEyttOJbsQzjdwcAWhNR0F7uiV9gZX0HR9+w0
ef/i9WHtEdrJ5hrhAjtl+GCQeCsDXmrMbXyh2oV3wNabjSPuhPexfET1mCdol8KMtygXMdFYC28/
fLQ15+cznygNlTP29pdRUKNU84LZT4ybBXv5yyJx+xEDj5pRKiLK5WH/owoywo+TgsGEX16ehG6H
Qv74fNqsIuKVmVwOW4o61LVbnvTHq7oFk8z2Ks52lVP/ASbMXEu1IZx1HSB9DoB6JGzTjwlE0ilJ
1Q098r/s2nLmSz6Yb92cRItwiULZlkmDKVpygrCnAFxQa8M1W1VbBHcM1E+DQ0yaIY9osFSpVvnB
3Yws/lf5/AKX9cM2erJ0zSqRXuXxWWDR6emIW2bhfRviCMlYR45CFxZmC4Ub5ilfVZWB9/mESZUD
CeaZK911k0Dlr0lomuDrdExzulPQ/eTtv0CgwhtMmDxDpZHR1WpnyINLKdD2RyofTKtvP1xNroEr
GqkNEfD6vgGWBLrqRh+zeNYFkjarWHXXr7FGQ3XxHYFuk5Xm/NRY7lK8eLOTYL/chsnkcVrOxlLu
GuYqzP7oeV6XYOaSl+uv6kE83d9YVYPKyQQM4hE0YsMrTFOOli8TtJCCTFOVCbiVrMLZpZOxD87v
AbKPdZDTkQ+Dz8ODmhaHGQOczydQBw5APulMrqp+iqSIj7/2MGCIfYwXgDRCOLXWRAvgHiIGBbpu
frjdliAqV6uQKtz2lywLzno7vr4RuyBDE7yWlk3RsLhCGgqlffx534dZhDqHtnehXDkyYb77nnrg
vpEafKGXWMdUf3/pHGq3p0mS4BFUl1l33kbvFA4/zfUH5QYnsmjWtr8xZwaq8gWaj6Xlmsh7/qr5
TJgUODU24QPpRE/ACznAO8K+YzBVOyKwB4aW3k/hqUGLjcAasFCAs/pzu8IBOkVu0WAx7wJiXRH4
Qg6DLm2mnlSKBHZsBZXCVm6NYbBt8UJzkQbySeFQXt6GySlEAAM+juDtMVMsRxZkLyWoe6qYtrah
Bx5H2B+WhqxYru3w25/XjRcDe4YlqI8a1okr5g/Gvyq7EdRVlGQu87bfEGsdvVjobi+jWDJaGcVT
sKh3fACZKjB32bcPcV7GAJeOAkN91Lq4lpdnVlE7is3qcQfsCLS7zGXGkutfRLg6/A8DaiiPh8nf
rMai8CcWnYkyA02/KgYXnvgmVCJf8QGP+dMZzEoYdLgodlF5rZ8WpqZRw3kHd7xgvOceZSee73UH
S95jxDzXwUnXkdXtYPKM38P4HrXoFM3E4+xsS0cm+on60PHhKzTbGuZQaFHtdMkLtJi3DW4luE0b
u/t5qtskInklsrm7OvKtDEhBeVhONg85O89Sohf5qUo6cXeq7fZzg2cnWrrLcddyCgIHBxwmj9/Y
A74bbkfMCjY4Sc5lnO2s2a1bl97g38WaFJi4KO2M+TjGhaNHMvVEJUO84L9eFRW+Nr0APE1zb5gJ
exdUGca2Gro+GSrhHqf3XNDXeCgYdg2Fm9EudY0tRouJCb5pQZMiVVEqEU6yPp34wC38ZYn36Zyw
i9iPPmR9PntSDMcg02pk2bmbNy6kOyc6e35h8nLjnL+hZqEoIAChzzqrgizasbTuAJXJhxVg/tOE
/9W6c4qjAH2RovYQ+hrciqjRd9Cb12Iby1iH0COrQDGVW7vmvqfPl5AytTqmJUVW41cXhMUFd9ia
9RsqIWzmq/dFfhjgLFuBShVSbcofKqau/fF94W7zEL9UmDO9x8KnWr9Et3HF0XwBSza7p0s4FZ6t
/66EU6uB8QLzLrVWacuA1/NjOv7oMYjN/684c2EirkWJW0YqqofezitD748/gPKwmjnD5gND0DSw
T/e0JDDxFV93L/JyfRzMxjNOEvblHFHu4bWEODC4oR1hn1A0phmw8iDJGNaHvm+z+qxXn83PyZns
w1cDrhCXrCpxYD/PxbhdVX8vOxWTJgX3R+2TP/RIMy094GJyvw8tBs+8Ja+qYNQukpzCAHPxVN2q
Uo7IMlSP01LSb1Elw93og+PrleWYsV2/Wsky30upx2ouWMBGeQMRKfHP4uf4J0R5OD8bChHNG1jK
u+d5nLuZmaXHOIoO78t21F35nf34A1KSyG6nyGFpwo6G0qCe4n5E3/BteFE8YuChkduuWcWPsh2u
+EAGcMkXDUsRYXpK6fEs2nRDe/hWwrH8N+U7xi99RH/F3I3rsxwKGbx03K61Ma0Py9B/IfppL4IF
mQyza95ZQelUFoTSmBnsyeS+ln2FSYOKF1NXI32qFSixD8dUWpmGAJOSc9k5y4+mPjiKxTP3OJH0
Ol9FVlmouzJIhEcKilBwNlbCHEJNQONRVFvChTl6mzofGnha3MeMLw8CZ1K2lXmqum7KCb4oexml
s7tocHGInQFq6a0ugAhhEWGkQyml3VVlGJLRs59YT4uOxYQvZSDtqm1qp8Nixd5XQxlIUKJle7vZ
dut64DXQRWN7Lrga28NK0ZA254oCVJHNn37VGe9/E6mJxJEKBWe/Szxpcq7lB/0Ok9K87VtpSz7s
q2ptQ0wzgzwuRH5D+qLewUFs/txr8hcWn0rHMQVfHppwjeWWEZBNokjAGBOV1kOj0Utlc2Rl7xVq
GYJxELghdu0rbqRoEefIdfo7W6yF7lk82VINRdrhU6M1Sl29NxXOttB+rkIZTPGo4ypfn3qN2D8d
AaP1LvDftyKxjGqK4iE19VNtfd3Vbud+OMf2zUAtB5UK5e8TLedtXaLByZGpqmKzxkIZ67IBQP88
0WQgrfuvrpAa1LxxJ9dHCGdIacxbUbCaNaskEZRQWk0sFvdQ6uZKafMT7yQ/Y80ZCxrPbes+fFcR
n0eXPs8m09W0kkpoD6ymRWJJYV9R/wS1VhdUEbcknlHoCs5cVQsFVhXjdXymZwCRpH6XNv68utsI
Ogrbx9gLZI8CZrGFSL4RrIcUX5PtJO7XVZZ7oRQx3+92pXm2DYxCj7997hSobe24LkSTg4wAQFKu
0Lg6t1OgY+cKjun5cou+IPTAmDEI2NxYDVbkCpnT3Gs/7GO9Qbh5+RSuzSx2G17/vgZnzwiqAAhI
FrkYWXFbQDdYLDMTSPaRBdPUyDXsucG9r+jMkF62qamcoR/IYwKxQbxY0d+Q89QPUA3ZheTKdXgG
oHOcWaew8+yEZ4tYxFdI1UjGNz4py4Dl/t38PfcbwxlyCkNa7vunLiTlal68pw0+oBctVnzV9USE
HVWYYsxT6JAiCTeLp2slUSCvmuac5O7XYInpSlsYNI43/RIs7t//QrMMGe0bv2kI2FXp52992RPk
6SLS3gP6qhyEtZJfQ2wbSmwmp2lBRw8ZKTR9VSdhM4GSgGQqz54gEE72cY7X58ROp0eRRRRtWb6s
vXw+M1zN939pf6iDHXP+yHTVlhB+lkDVBFZxC9v0VAFaX8mq6yqQsZQx1Dsv+RYiu2EbascHbS81
HjCbFCP+4dvOgOyS0VIrFkLjhVOlrJimrHYeZMsDNrtY0eAXtCBVgoJ4hYoK9e47Ym2kUiAF7I6d
XuKY29iYdlpFOOFr1OA/xsCLo7121YjklCA3Y6r4vQ3KhVCozava07YFtlU7wQF8KgNcLr6yiKc6
aggMbjuCCMiPGJ7c1jc7fn7oSiRruOOPLWgSTVAGkA07Oxg5C0VqpPvgDxyYbQG6UdTr8rozOi7H
3IixHSi7ny0nYd1DU5KG7rFkzXYT8oKnm2/rsfALv7Q3wpDTVCd8RCOso7tVPTIp4O7YrP+HDD9S
18A8yTDRaLS7uCogjDNLM0FpuOs45LOE3dNQhir9btkAaMCl2nerS16rrTD1DbLhn/hFrCFp7vgH
sDDIqfcrkjeVaWcHh2t+f/JCTL9apUlPBWYw0kFYpc4dl9rCHoaMGXiaEKbW3TjvIW8rYCulLkFg
TDD64xa3YOn/Yn0SuoMXxgtTVEIQB85B/HgG9wa/WLRMAh3MmSDuhIqriNHt3OXDifKEgdcN/e//
Yhv+s1umqOCHbeGWJLNmJkCFNXE1S407TED3QcL9aL5p2RaioXpuqLHScheAACO4cgsyS67v3IDK
7I6mEKIfLM3cRU6rrL4ned9BH5hlXAqwU/PIZ75Y6uip+rRc7xns02Dqasvc8LU0VkPRIKtod68W
I1iPC18AAMRwY/aGEcCiLv1LEq7QvPU8JOGdM40MdOr9JdvK7SswojobVIPkgMDi7d1qIsTu5DBH
KoChf1XJVA3NYzoUZB+G1dAgtE1hfwljqmt6WEXaKpTPr2GwHiwnDHeWhy73CNM5VqR9S45R0a/W
A+IbIHNtoUpMqQkseHN3w2Hsp0yAUeVTeXF9gdWCUQa6ybPNI2Fn11qGkJsC2T/2d9Qn1f9IX4sn
1+EfvKl1AMt+QxgZ/mQyISDgV9K7nDF/V/QXNiVf+fxvJme2NeTOFaufEX6Je8WIqJMWHv7k5lWq
4LYew9MfE8kocHWeIGX6fos0rIkq+rskqehUhHo2tX/hXRLmNJzFGmDKbZRSW4puz6MgnXwgCZ26
wa9m+1TjJz5XoXoN3QOVobQ+Ml32cNHqiT5RqqSHj1hwLtEDAvdZYr9ETVjp3McfFcoOpOgyco+H
F6XlCeND+KU4qvWZqJuT9g8szXppD8ykGfr6jylYfBvva+PKsctbJTvbIjgbBmCYVrOxfx3SwJ8S
g8rBX/NcsViIosWo1Agd77CfyyysTe4rHzZ4phYXynnMev90Wf8G8JpVKNOl3Q2B2IKS71wrdTLr
Rfq+BMlB2fEZGMI4ADB4W9dA43Up3OAYBb1w+Gr87QDyQQtNkXQ24GYrXOjlG8UBP+maIXQuJ938
Q+R3US14RzTzO2DIXtpG0wZCteoE9U/W3V2uumhYbY60/UtbC0qkHWa/QMT3KadK4MrPV+iT07f7
VtIEbXjWKgj5kAG37ovRHspVklxnxp6w2y+lBsAkymHF+e8Yevv3KCiiD+Y6StlBAv+eTaGYySV6
7qRD18nsphZWoksyXK8/H4n/Kwh96ZSwaEdyoyv9dkuzarF+j2WDLLpETEfpKMmRDWcmZ1e/7XMW
5sd4p+qQYCciWln4Kb8IVpacdsmOaFyInpKxHAblkPqPfowwS4S/N5qovuxBR714KTlLi2uQJWvf
dBWoUwMpTbQxGmDW0lpki1ag74zkxR5Qd2zQYkO0bWooBvNBz9gKMffZ+738N7N2lnbqD1/PhyrK
X052VWBUu8bKGJNfl7CIKuUa60+Ljebfzc7XjGYKQVpWNuyWy11y6tVEHdyJVmoWP98F000R8s8C
UsnaFxOfQd99PDEwu51bK7ZEAKTweDbTP56oSk2Qj1FqHwKa57hWJmHfCruUwGy5h5yoZg7r/D+O
Ti6EcfK/w7Uwl6DL6s+4V6V4bgGFTHSh7A045VE/JO+MwaN6s4YONYkC4D9CNY6KYuiWdnfwOctb
LMKGkvQ+M04ib+OhQn9Wh+p3oVwEsbCcyV89J5ExT6S24o34RQuY7ToRd/p9dhc8Ezv6/hFLhlVR
tr6gXe76kPVjSyR3M07tYcp4AUtolSo1Ko5DgIjs+qiYzSn+1G8SQzj1URqub3Skq0Ezqbw20Zg4
voYeP6GRmpKuymcN0REhgvhLfHtj1BGEuu0h/EnFWfl6qugeqw3jwDVSGfTeTcOdqI61UEwaxpDn
aINKVmOHcBdTg2e0s3Sv8ZW7PPdLCv+YHjSyeqRRVbvUc5hW+iJSdsJI76xn86f9gToZ62LUTEfY
lrd4N7N6c2wi4yaiQ0CwanNv8APPjh54d54gUaWdQ3VFst0jHVpCi+32VYjciGQLBDKxUS/hU0GS
XxASVglI1Ehbw1woYIdSxcgeVQ0pvWWzIRbU6LwuIqIJ9d+HEo5rC1gV38BS6zdrT7iRHnRCHjVe
84+Z/3KEMuaoy9LDm3FNd23MS8YvZge6H37yd4KbQBEIlzLVHhNYcS7J5QUEsryUWn9ZI+tVCv/i
UEPIeRASmSEGrYqh0fS+TsJPsBR7OvjKNcUzaaotDPJqugnqU2BZUo/vRPrGPimNG7C2V6P8yeom
hTQTao8cZX/qYF1pgAr1ACQI071w3z7sc3TauHAhN35PpWemVY8xWW8N8uvx2YNBX/BNkr/AwL8I
/25vxyfa5+QTEMt15YjtlQ5QFejV83QdPXIxOus6HDvEtC7hjM2e8ef9j2ql/7a+cCY3T/+uumar
iL5EmRrpyggcu/ufVqySBmYpa8ohxtHPXIaZsnhkc62hR62OEr1BsXVtaFDujToT1hXUNMom6SrZ
+KHoou4ByBelVquLtlCLRjn8W94EXmpLMg5IrEXjclH60r7W+h2xpJcSz0RUbVHac1XvgK9YL7Xp
RN+lO4XMu9K5sC2vS6NDTcD2r1d3/bcMe0Ok7PwGhzsJ0BYLRTSU3JP0/8y0blLoryEN2LjUs6M1
lcBU2TuoX1/GXEayXqA8ZFWwgUXHWBUEWKM2UAcslyUmd+uuDZBbyUF3vKl4hSn0YFS7rE01CXYZ
XMwMB4lwtJbLhDVVXg8RSvZTzGHytNW32hVgRwAJYLe45nHHqu2OIaW+dYtBEz+HL2l0jaXPEUJZ
Sdnbrv+bIp0YvuBjxFPGhUEdkBqLW9EdL4jAPpctrQk04QDpUlInigYDysd8c65Lx/IJsRw0V/fG
q3ZJlRJ4m+vUCjWSYs4ATuSC955nTsSD2YfFa5c6Xh4GPEYcAb7xAGHQcwuWQ4tBGv/mAxmaELIY
r9TmNelPti0Qt12/u5pa+mQPSgLNulyX9ClvsIQa9MiOV5upPTX8/+gYUvJrMptSyYbb7wncbfN2
2ngRo3euKGHi7D06jQhKBKbI7sPXnBiTtom5O0AACNJUOUAS9/4ZAxCjLiIErBWHB01nIjiz+nxM
xJZWy0eGmXU3qVTg6pXACf/DYOZvI5v/XBPPFuhih2O6S+A+ovE0kGK9TM9avlBZZUK8Y4tyQXGQ
U99Cto3H55+U//j/jQ1SUvLhScApl3DUwh3+7OOglFdGu6YolQLlXYX1OwsyWbGrUTXDyubyYe8T
eEgoMHKP1fHwBHv3aWhIqKaAwP4tPH+3XexffTMnVIPGaGKnTHniLAewCIVXNVP/E4cKwdLeRdWY
x7eyUfqsEmp/ElMr8Jkai9LXyWhpZlzWXzQK5Ad1bmQduUIt8AC8uym5lGioWE1m1HoqcIFJgTqi
8ddg35CT//Huouv8/YoqxRPtYVJAGTy3hgzjh8lbcqV98lKEx4sYeTxltsnYxp5So3FfsABfpeJQ
uhEdRw+RkmPhMIM5wp7e3otky8ziM+/P3GF+ADGPBr/UM+vcsY+i99Yy1vQ0l1aAdacS8oxuytji
jUyZCkhZxDRuXI9bT4fXG4V/YzDXYjbxUvWmx3V04a5ww/dtuiG5UlcwFOk71VvE0l6k18krEczR
lolegXawBwWfJ0PG9rHZvKJC+qXmPF/4ATr/XS9vnateyT2Z/38sn0LssViZMxd7Ni3kr1B3a6wE
tiAZN54Hxo++xD/sebs6jaVUMWWUKOY9gkhBW47JZwIOJ3LNoPn3VvGadZnLS9HrcafmzxSDJzp5
l+w4dRd8p5C68JYMIi6Se9UaHslxt3uc0nJ7B1kZYsOCTFu+3r4XfOuGvBICbM/CT4+oB0QwkKdq
FDNVFDbqzApj2dKWivKMww3g5SEKLBagWEAsBcI97mOI+Teknof7JTCtHnWLkujCgS94LZsWGrGA
Z/PDPZdgh53xfuh5ahKcag6tWNleZpaZn8CX1cjh58cI/PJoCu7Gybx32kObzAS3N+gHlBD1jglQ
kwIyX4ed0hDJE9yombLyIa9bcleYkAA/XkF2EfwANzMccPTq1xda3YPSNjE9WFv7UahhT//f5m0R
I6bU0r+8/JsaXk8ztdxb5uhz5iJBnATMFnjYOhtbbt1WD228AkAUDN1PtzTyXYgAve888D8iYpZi
q78eVK5J2UPjw6tE12+45ktiIjQaobYy6eguOJGJljY6BGNgr44V807aVJE+SBDwGiFrbCNwqEyR
27pHeT/8UhYmpezIGgTGGwOyI05MalCbWKCAPJ02BLgUULHNdUPcjtM8ppOfVHKWsV48dnP8pXl4
+5Hj8lzr5IFFuPOXtVH58mo6OvCuNLCwbWlGOpJ+mgSiYCTSODlP7sfeTFDkYKDj5Vi5ijX31Sd+
h1zLLCFsX7Xwx3sTb8L6e3NZzwVsD7RH+t8UU8UoJpwmQ4El15ZossOLZgehESwpyHavinQVS932
4oe9mLX4K44d3/cYo1w4zxgu++g1HPnHiBQsptZAJw4W+GDRZClvJcCLpAjqTSzxKYtmJgsQl0lO
CI8cpt3HxbFtOVPUXe19uzBwn85Fh3lxrCE2r0noelJ+lZkFdVq/O6zBD3WvuNPeOxoY+qPespre
2TjQGv8mH+vbVJQEap99QkRlX+SflKGsTkSz2KxmD1L9VrnhrpCj6vzshuAVGDWp07sdn8lu9awj
qv0gfFGpUUE6IiGyKOzyjwi8rhqubfixS1uaWKPcS5/rs0RU5raV54bmjXzPlhLN3NyoHbWSneCU
A/vjl231LIn2eVVPR8ccnpvt7wS+d2TRfocnF1Vnwg92INPIyKeUndJH07arYJ8VEBB4SBUj7aBT
Oyf2DDdcMlfnJ+JQTcrzh2Cbe6i2jwcUdJ9GKVuo/HDML29sIQ68D+69raGVouoG+RSdE543AttD
7LEuhv21pcXe2OkV/Xpdq2ERITRRRIEp7hYpB2QOfY6D1RQ8SMeOa+SmyeMM7To9ltC0Iuj+8TIG
P37Mf0hz8p6F+CNpXbHZ8fuNz4RtYpumbmdEpRpg/OkYavL/MsxYxX1WccFVt8mqj+gm4t6y6hfn
vq+XHWKzdSlFhdk2QHzYXmOgfr4uE8UMSZSwlBRtgYL7hXV5eydH6P/usYsjEbr94JXHpsNf0zLr
51PM3Lg4KaZJH/uuoayzt0B8Dm9nMP7WPpqyrgx5pn/DbC0/clCCiiY7jByFs/ik+RyRDhEu/lCA
FnCzJ2qdotpyrQwfud248Bxb8kLsqhrmq0y9QOQ+g+Vv7FfPe7xV1tKVEDQaStBwGNII7aWYESsv
F7xaqBOTiz4r8mCKBaK8VT5ddk7MP1RZWFyLUmmtMIToDrMjgFKu1bJ9lgwR6rdkCi7nXd5nPUnd
e4wRJ8I+OJ+AR85lZ7wzWfkX1uDUGAkoimVom65ABPmTfLPh5aUwOTYwgZv2RRv5xRWo9yvDMgTt
cuDZ2FBzhjIjmmAmwEmd5LPepUTjHb7FoEsas6efXdts5RHt+p1qH1O2SwGn4Mkqre7cNl2bZsJc
xXIsViVNf0ZShSV3P889MHvRqad2X2dxf8jmuO0AGKntDiZ8FA+wsDJzyPcBvGkpb5a2VQabjlxd
Wm8XbZyyJ0MOMelp1hwEHKXF+ph9eFIccjafJHiPXj0PONEkwq8ojAvrTyo4mV3xX6oq4sHwsZv2
zix6h828H4ObY9/mOIfSuXZFfaWAy/Fs0W6u3EaSs/5HyIzIksIycK9hJSgoUKzRNM2Ewl9MjBL5
0ogtc0eqe0p1mN3TM8f0zEWRc3M2W3x3S4skJ7C07zE0g3HHgrQWGz9+l69HEB2aU4BRfYiGB78w
YtpAZLaP9AgC8Jf0wxV832kcRn95+cs93fdH+yvyltBHlcL4DbgBDpEkdkR0AYjHJFLMQxTGg+IX
aMMjt/snKP2JXzkz6dIM8/JW19D+eDn8wnHVqpVEi7U2gdxCQAAg4PryULu1DWyla/rVM/t28R/2
KN4Hf2WF7PLZbmahtLXNrAaYaJOIHxD96QcY335BYLF9j2x9F4jaYYn5wGPN+y/4ZqeRGF0j0tvU
ttPQ8j04qZhZ+750MT5qBQB6AXjhkt4log26T+XfEdltaLt+XxQTjAXdP5+jJw+0WP9VpAMNkbBo
fXEG3teQpKYg71GJhiuNY9diTR+CjiLR+r3Gi0SKAVRHbb7XvxoRzYWyjvYfk2V+WiLvDHwXoI6E
QufyzYyO3ABMO7H9MymJlQza12xjRY2ZA0aczNu7QhaIkrkQp35ueh6KGOCysM0WxjY5VfwgQJ6j
pePOH4xIAiCzUlp8zGWJS9tnPlnRxmKYar/P7/5xqmQ9zcnLgwqwe3c5cDZZgkRRCnpUNqFEVrOe
IYbKp4yam1JShq0tsbv7Wllsesp64k1z2tbfyzxGzhpdZE94rqXtXE2pgWwISe8kSwx6RvAmF1s9
AoJm3g2PJd/C9L24+7TmyXg4TWUq5Vd25VYaZVfFR2c0CwhYFt5It4hZpo4JjAdYbnXry8DYHdOh
IYd9zAkRdFoQu9ZtQInFb3ePKBaStiu0X+riinU9i+dpCGgoxlFzjrHdVx29WZGqB2FH7LlKkRIg
jqzjdP9yeqCKw6UIhdFUUXtT5QlYYNlVeau6nVdKHyu1ph/TfBB7Yu71U34LdoEcnnTug3nanH4W
ayI/tTSK+VJaiebTN21qog78Syl6z+k33Ra3cHZQ30ha9ln5vkii6T4BQYC1zihLOnvOAWPfJj8/
nFvnmkgqNruuydbsCYoMOcAnmh59RyRL3CiN8TGKoj5K3pQ4TaKPBxJaWqb4OgC+hSDwV7dDWxX7
DsRk5tko0zhzNwPV0Z1Ov7M3eSFKqBoO87ujkSWdiSZFfz1p5azlt88h20p5OIUlqWpoanE82NKq
JWMp8wuOxlDx1q/BkbQdIaSAytyrmapfpJ7Hd6KpkOZZyQVgyRCRQzf75Q4MomdKqUTUa0dAdCEX
3MWOss2lCaXPwKQtHX9sqYmrlOxei4n0fQPHRRu8DxqI47Qt2ieCbmllV2tBeMft9WWUhT/EpIED
ZnUYjn9WcCJrnhyQ07Jaooh6pUigyZgyPEYVV8GZ+qm8BAq0t0sE4sH7V2mfkLzfyWwnaS7RxEgL
i3C+Gfq2sWsWJU7PzwoOzdcc1/7N5NdmZrOJ1WR8oQYTDT1LvDWn5F6TgvOADCtZ52ahAG0rhmmF
35lqdSKygjQqsCp3rL4ff01FR5cW1k7CAtIxhjpdWWmDJI/X+j+uQHdbZ7iU5TR5yzkWQCCwvS1P
QRb5obBi6Ptbek5XPBKdwYqfg/eVjYr7hNnuIVERVAcYDw6NXD457K0m3QY34ZjxnRzftNPbYQ6D
dIhcYPZRXxKY3RtI500gFvdS7IAWsOKEdQvbJU7Q4NqiQZLNwJMcyuSfo4Do3v4aTfyzpnY17P+N
YpR7r5n1kMY6krcQQnrNsZ5v7HDAMCoAoC/zVGo2PaCp687a7LyZByYedARNWDduG4U9Lqjmj8Xc
2zX8luH23xPDv4xkp+PswZuYYcyQoQUaTrhiF5hQVunC7bx/WDTRlzQduXDs570cB2ov/MxsUJVa
MmB74fXjisd/YP8d5T1ubPf4teX0Tx1aVqGiBufAbIvcVp2SdYoptYjDA9aBUB0QeBGtJsG3fHzn
lzwZ66w6D+o13bwsepw4c6ePYSRIz6iWLzawnIVscFvzQD3GtZZS5YeOow5TmgbiynikTKyklQA/
/NkoIutrDYayTidZqK7mUARZp87XvK6QSRnFUfZis9ka1QQP7SYqFZhaWfZjGu2fdLHHi8FWXOwS
liBpBMhJRWjAUu8ubKZV62YR3fTJ9EiSWIQ5Y0DQrcl1i60ondgGEv0O1K6hwvfBvBVNp07eumut
Jdl271Msayu0NcfRTDyV1W70RWhlUK57HEiQry8UyOghgxeg2nz/cY5E8BjTAAPFlZxh9pkX6Mia
AbWvU6WKbrrnQutWEfzhmaYInKaGGVqDX1RIZK71YEUmvUD+MF/JFIYouBpCKlp1rgb8yXTBQBY9
ln/yq7nuawDClEUWXMl0vW94m9A+sj1SDvYIiHIEhjQMtvUinAZGtH+w0VMhWLToTFtrvvsbawkb
JtKEX3nTxoK0hVLy9YvN5pVJUNJwsXh0Ic8RjLzCc47kBlC0zTLyL3IpDxniRxnNvjBeO+BMw5hV
z1VMp1wxO7cwgbJTbVHtazq/cKJIL04QCemZEliGdCGosZ/2IORmo+76/PgEi/GiwaFgCv5hWoIy
2PpUjRr41U4ENadLLbgsf8vYV8B1T8gMRAqiFtwIbjtADdhkPYkg8bk551kHCPfXwyuAH3EmW4qh
UC7/octj1xgmfYC50uPhYcPCL0vYCEJ1ypLGx/955giUyLfTDXGeoUkVwJTKEpNj7VlzWUZ+nAeB
kEEquqWgf7pvY/UkFU/uwBoF8TsfxKTzyfxZbvdS3u+Z6NS/F9a8k7YJjUNsirsPyOow+sJZI5du
CdUtXDQ7JbNAz9eiM2lE7DfumdvMdySTnZynLXDczilg5MW5owpmY14SOGOnRndTOazygsQNnXir
p+SaTaTiLlvWfQJdKN7g6n15BtP+td9sMxN7WxxyavGnk+Hd8Itr54xVY9zDZG5iBlm5u6ARrduj
kgiXhXXnS7aiI6Z8tfcZKNUOdneOaYtWFoLxWQgddHGR6VfA5G6UAc/ZP3AZUPvsEaLDbUEweDby
C346X+i3xcFWBy3Tf6Zs2z5k2VInu/sRLqdpCnrVBiUekyofBn0SxOFRMQGjhourjwiPXXKl5hXY
tkch3cCmQeMZT3ISzGUR4JL/NKicNp8d/M1bNz2dXUXYD4bW/+EDl3vLLJoDcEHX/JOvleYkiRU1
cRCvUv9BZvO6ZgDujAdH4FroasQZG4UucHnrMjvZC0eMrcthPVwJhfVCuYRjviLgZflWU0jfnq0V
1l9uwG9PDmQEANCdmqhoP3J/rxX4PYUF1M3cWcRYJIfloERyytKTkh50bTGj0PTU7y8P7Kr1p6WM
DqPpINElA9vwBJHSFehVvcZHr7QhpS3172OG88ZlBENIhh/fkSGmuvO05Jf1ReUf4JxkZseqH2nm
x0y3i7X+aCLscWKQSTAli5q4CS+osS2MpK/Gam6h1GuEHKyyehyuQnVqKV2K8NyvoArcE3AMT/uZ
ZA6CY6bL3m9pwD5iA3hagrHXVejAsR84HK4cm+ua1K4IkTcB8PV8yUwK/BA9yZbdaBcwm9wNF0+h
xHw8gl1x/9TNMM/mwRIbJvm/GuaJx+pNdye9FGUYr8JedZTe3zbhMxnTE1V0BFeT9AiFQ/Xkp8Ju
2HGwwT+KJXGiqbKrb58NufaL1v0l2EmKX7iymvqsmLDrmEnUlRrvpPfPBtAhPGq5mEsx2BtaUu9F
R9jCIHIDxfo30/uBZH35nNga001mNdVnUmmrEP6Xi2opnHEvp99oGtS2jpcBBEFO2AN/SQK4aKbE
kjOFgqNbfpQVKEBQexrbrF2rHnOhho+HAp+4XhOemHUeEGHNSpXFBKbjTw9z2k43DmV43L9vR2+5
VJkUzSP9jWncMs6HDV0tFESeol5PYsA0ftcHEdPW7g1i9oQHCqbcS2WwKG+OPC6KirJVTXl4ayEc
ivaN+3tjwwX2qfO0o0XR2S71Z2ezWMPNgAycSemJIvHzUM3PBPRyd6anE63LlAU1TONK08oVv3k4
ESPWRyLoyXedZpDiakdbnAvBJJI8HxTK5HoGT10E0gyX+JcezGQDQJYGfLR+OAKrx0i6LlMGQPMK
6yON0h2g1akk4yfrU1CHIyBlo2bgcxQyy/VrLlend2hncUeBucjWluJN+av973EENa1sVIFAoD+S
IVBcMp0hAWHN/3k13fyBixmlpS1MVv4ck65SzWswrNz185CGKF2aHqiQYc0Q9YD8D2RGWFTZ0C0X
+sdWCl/NysB4g420i9TOK5uy/ZGH+WS1T5Ce4lQXZkFGdlBJO5t3JdxdPjxXG+NX+6e07Ns8KjXj
n8U9n8T60yhnI61ITYVAb20vqMP/iwtaorHgyMQvgwBG8CqIOMDxo3aiSiK2rb3/zSmKaPWcsifN
sp/JzG1p9mNehSt/UXNaC9xXaPABrht7WeKN9coqp5xy6imFVPQ6sATl5j3WKSQpeX9PW/MNqK5V
n9+WshUxlSpC6X4QTiYkhy3CAScHXvbQu6/cG9LVvhTnLTcf8ksv1p2l90IYA9L6wuErwgT/iMzx
j3BCFYvi9vkA0ZeTyFNF9ceFmV0gRH1lmKIx5PPBYjpIffd0+u8ognhjsP6EoBGOmjuMO4xM4J1/
qFh6awrqwFfL4gcUFRkpbXS8E1KzAQ/43YUsc3yceJn7izGSWVBvPhyryb/T7KjIeO02mpYiFfgh
dzwjluhMYCBYqRwf3qOG3AiHxp4nIG31Q7O9RFGB6k2ocw0J9FtsKeYvPaIP7j9kgDpvVhHWlbXC
BeoVbAzUnarbACY3WnjiibwdHaZCWsi/d3TUS9gJelHBjBzImt/zJdNGm2IsHVAtJvGCtul9GO1i
+4F3oWOc/QAlUSHF9uOgRj/xuAAIpCVOH3l6IYIbpUHvp8ML1l8BxmvcjuNAefMadqFviuH/Tw0m
QJ5BJPf8/bbTJiqpLVCO+NXV0m19pEm2Zyh3HCmWK3HMSyRrAVmkHbP3K0lHcT/8pdXSG8W6CPkK
iyRaW2PKzUnGETVwHPDbtTdA/9l0qK+Tjodx20ddOOcMAh1zpAc1Eb0ByGLprWLivUixxNRjxIF7
UCLZayWBYZtjk0vgdsIgI1jqx5tvXNG0H/LANFsGvNczJTeSbJymcfFPMSEl7O2F8VMO5j3xVJqB
fuiQoYzaov988Mtj4A2EzK+BbAerSnJcyCRCrvuh76KXyW6tfzglsazcXmG8YGuHaglYz7uMB1Dn
SxCP6e8qWjqNz9teVv+PeNCJSMioIXWlhFgWia6CUy3lv3Arfd78o5mVVqc3NPH9lMaGTqsGonAy
Kq12xo+jM4r0s1/DYMnncj9D+3a8l4sIGnOkE5zVTn5KaoDG6IBbi7eBO7DItQ11K5kNxZaEftZk
xAvrhYYvta1qbjzX/PO2qL0A9BeqDMWwkJYqh86QaaJiKBv2cMR5IuONaKDhqlwUcwtTIzvJm5tO
jBhjF4FKaRZtkT6+q/YmGEkHNX6pOWE936/jkMt8CBvvo2yYppDsbj3vejhqOno6oip0Y3dOC9oT
MTYlapX9J4WvV2LnG9u0fRPwlUu8ooA598ed/MyCiu1tobtwsCO/i4NYzBpZNKgb+lM6EIcCQ5RB
San96EgYiF0Kazf2CEPSsf9iiykw/XLRVudKVAw2lkxhYAJp8A/usaR6Z2mDxjRM4yQTizvfNFfC
w7FxGA2eY4OABSTyrHT60K7vKxTsyH2lQMmdXMOBrVty7PG+hTYy5rzAyAk8BTk2zl8URN0foxsQ
stSdIP0MCg9skmbf+7+DihyvGKo6Ac0Ciq8RT3odnGutZ2ORCEHEEnjVJafZTopsca/TkRTJUYFi
lG9IQwZD9+Vq3mLHd3a4E6TaDl71CvsRtGMWX+CjAwfqLhb8/WvIEDhkDLSBwhpvAoYTFM+OAo4p
yleHZdVWubuwnTD8ANV3TyMWJHWjU4lmSfQfkd1ddy7/G6LMI4+xa+3k+L51yK4ZRqNCsCi0Ba4/
6Owg/deHau/0T+AqWAE0s7Aim1JvBJyhqftj/U4mkrmmqY7nlZ19U+K4kfLOA2Ucy3fvvbBSmcZy
ncwzo9yKjKMqotsaPibKZKRzsWDgLhBXb8CRa/sWFhovVHHOAyZkYws7Gbms90IGtd+zm0wsxDMr
qwu4EhSlX7zN+/z5/aYIo9Qb7a/Ygl91N4y5hjNynwWmBBKjZxO0bZ9ddsV8hGtnt4u7FDoeJtXp
+BX0mHUlxofsG6rr1TNvnUki4qxH7o/IGLF1A06A8BUZs9Xcv4to9n4+nzRFslAovXu449NiUbC/
AFs4GrWSXy0hA3XoXG9iIv8TsrRpzySoIQW/mnnY2fwP1AeoB5qxdP6LdmysvkNTn7pphbkyN1P/
YTlKyR2wHYSKXHhWpo2OQD2YIRLVwAnrH6ZXr/4Zz8C84nSEOUBZJWa1xnrFECh7ySYnUiE+6HMx
Asb+KLGziTs7fkn9jBo9zFZxl6QL3nUJ9z3AhhqKWW+041XYnrArg5kDumW8UDJY4xVljdPD+xu2
PPQ1B9kN7lT0SzvgiqLukvyHzh1fyrcbcpNh7Bvsp1NDx99A4MUTcUFkifmkGDnoj08+7P3ULwSv
bR9HhhNKoHNINHm5Xq8UBuVNNXzC5mjgShiNg55xptT9gqz5MBkuivyx9RcLrbDrdEmSB7Hrw0wb
iM5VJvBl9kHWk5lQkU+T+dyli4ar8BkZTopi6NK2HU7tYq2R6UE1XHnSpbyyXSQYQUS+ANM9vkc9
OK6/+nlDq1E42FZGKeMk0fZMlUxY1oNqDn9IVyIwUtbY50T9FAch/HX6FUArbQ9+pobQS5NThHr/
UQ16X9cCDLRv0fwvnk1dlYznobVIoQBh1aW1iFckirub5889jjNV6hr5kDhVxO0KM4ghH3CNDyLk
WXEX00g3RlIpRC1Ge8KaNw73gNp5INkbZoFEHEvW1dcbvH7ql5mseu21hwDQAnK3vHRxp/Gnhglm
Iib0t+07GlkyoR5XC30lN5OiVgWDNn9YoqwEUV9EhkAZ7i0dMQwMYf/qHTMYHVpQdh0eUb2CqVI4
2aGgSCevluIWOVU0pdcl0xhnW5oyXDhNkzDxdgHW183YXokn0Bau6CxrAtUuEFAEHjCIywObzmOL
rTQ8GbqfZUKngqEMBCBGQn63l5sS/PleX2fOIlVKj0hGBPLrFhm5cbqbA2W3FYOaIxW8qq7EAIp1
Yws2DHvg6R8bc06jMAevhupNDOmMm+T7FG6TppmWSa0WDkteKTetue/XZo/o7KVxZt99yO9LRvg8
SRGK71V2+UlXpm40F4VE5fnAElhS7gMbDir9wcS6UMHtxexMVF1I+p6LbyJeUfUAVUWc4eoQ57Xu
O6sAenx/QKK6GzTG3dttKfYKVCGCT4arNqf6FAmphoklq0grU/0bhmziatxTV8D5CJxHMeXvZ7Vq
7Qmr5yt+bXvPHQUIZOS14i6+1L+2Iz/UEsAOZwmmor8MU3IB0mk2h7fZWfxuCR/AukcyXt9mtv0S
aqiQsqgZwY0P7cH2yvfZujtDKJk5GR/1+maG9UTQpCKGtsP+jwfrbOsN2TulpxnLOdF28LOpuIb5
DayOK/biXh4OqUH/0Eg+UMhHT9M3oM9KzdBdOnQCgG3Z/PhU98OuRFSOBpTQ99poi53E/uVoZsgR
Z2dlqAoYJqwpJUDhiFFBcCLIxtO+L0VaX8ZzH1xfA6fRPwRStQ9AElqHq+N1bKDSK2aelWgFj8d7
GjvnzfmSHf4WAesB4UkPc5obTVQbrtiWWDObb5bj4w3iM3a4MDaZiWLD5Cvm0Lc0YJ/K2NOame+n
uu4w6RWegwvNcct/lEpDx7Wt8e+dTUgBjGC+sJEG7M5SRdxIk7OLYfA6HIVGWtKkAMzONxJaUXS9
yPVsSsrc6hJ5mtLhUDUF+m02TdOdrnqQPQcLX8ix1ph2A1VZTVWmstCV7zHloZfvM99TLfDRdj31
BP1O0+uGL4fZeTMRmAJYcN/qydBspKCdcWHIPzLEIp6OOiY6bLjX/AdRCzyL+cAXJrQ8iBCmZDog
4GU085enc+bKN7Aa0ZIEvGX05Y5ylrCDZzWZsjhp6kQzBjqTMN6cQ/Uz9qCxVndVaWJOCvn2/e7h
ijBvf8OBWSLg2nV/KkTvlkG3zikIV/QPvbLHbkyLuqIrSIESWJqBwASJmNwDmD57TE716lUWzUP8
p4Ab9ZGvDDojD/4pTxQ4qj08R7cphoL4htLVjmvjI0PaENJtYEul/uNJeed09D0UmvXPLTqV+yDW
Xm03kDYD7xEH7amwyrQQwpf5/HnofWlQv7ceTff1vDceBYOo5/+XQ6OiRLACHx04s3FZN+bgnhOn
fbQCvd6kO5XtCm5CXkY7T0BHJdpU+Z8lRfHlwiRMt5GFNRLHv3mYLwGgV8wOMc+1ucAv4WgHzu3L
wwjrvlTmw51RvWbWOpfN88FhKJPeh87r9DH5E1UsRIuPpjfPT7lp8c1otuwbNB2le+UAjKNi90BC
IAOLKTms74hrBtGXVUwxxflFi+TBJzEvZ4W+FjPEnUH35l1/6jLDyETH3gPu7SYmJxZrOHvhsOTW
IOHQz5Zcdi5SNpgswE7daceS/ZfqwFYkFmOKqorv/BdUI0rnuGQpZ0wLVNB+TSUVz92/kOJFX91s
H8inx2HadlplCGyUBL53sOSQ2YH3wj/rjqlztJPnKJZ4s5CG7+YcHPG4fzfqEjT8TdsEU/Nem5vG
pIKLAiTWxsjP05GTcv5LYrvDEUfoRsw7Tf2XpZy79psi1ND8pBvoL+JXRgZq4DCiICvMzcRwlMON
XzjFLTfXXDOik9OXbxNUmH5JNoagBd02JmERXGcQ3wuZiKBxoo+tucJkCFUppj/pgt8lyI55edVT
s+psYqYlTH/JEcUSBFiqv2G2AjVScOfLobKxqO1uejadn6HGP4MS20chJlJMYHIjXzUEhVJPcwGT
QuoOzC9Vs5e5qkWc4ohZ3P/ey4IS9EjhsR9ZyFqWUMqEK4OgEd5LOdbK4nSzh0+imk1kmcMw/M8j
DgbRUn3xDs6CCtyoflEymjKg1ZVy56wbvoqRYi1npX+23g8Q3MSOvM9A11kjth1+kl355YFUsiGl
iDHjtWv2nprEHpOkXpTux+YIAMFosb62YYTB1EBDUBRey2R8YgVeSBXtr9U52axuUMi8dgrpqhiH
kRVtKQ6sd3C70zzEd7PekAFHNfE1cIKU1ZvS4EecrWi3E7QctKuuZkUTvHttjB4wEytgbOmE1gzk
wmRl2mfitBfuMHggjPENWjVPKegWumHwDzXvqLG836dNcC1+9t2cOuXkd/XMYBfErtycImKl7wiP
nHTor2Qx9+14RdB32qCi/k9D8WKjfHKG6AGlAqWAhdiR/vG1KO7nbERzawzT3v0EMVPkd9J4wVUE
uf74UIy8zPHYrn+GNgp67V2oSnOtLyrvaLZZEYW1ao/PL6pbaPQD/fH9ovUkNKSm0wn92olVuQvg
679wdAasODfOM3tFGX6rshEmgZ67rmnBBVIk3HKgfDhIRNS3TuY4IDNw58i7twgBci4QSSmdPsfl
KcIJbev335b2oppDR5uXahHImsv456PXMyS/Uh8+0Rvo23Pwm1Wj/rTfXEUVsgxVnX0YRVlO3K06
9NrP5/1QkYAEGuJeaCHOcVhlSzZOZhJPoQNFAFqSGFx2pqie4zmmmfRZ00nykWjrF370P111MpZO
B2h+H+3HwA/dQ7iwe/8aYjhhayvsHAchLbYD9mmFpq0btlSmLNCqXP3XyGG0xrmgfjwSF9tZEmfT
n+6N5VK6YgKeuQSHie3KaRJ6DH80A//nqsEuOL+wuse5CiSUebj2/M/942/94Mywv/ZlWHi8qzvY
yzT2hFr4HGX97KGAz4gADD7AlD61eDNypEgVJX8d8MxyRG1WkBcjV6xrn/EbK+yQBKxaDP7yFl4K
dHPCKX1hS6KYYXV+M95LKuHz9K5uB4XO1M8RLCDU0J6FM8Ay7b9EGgJlxVupCGt1F4xyzCvtYsqY
5UdHRDDcTxcZ2dsQHhCfg//UUXNS5td12eBvixnekxNRtCL1juy77jwXUMpioTboMXIgeD1RKv3K
YZPNwDF1RIKQ1mEwXfsNyXVEVIg140A1QKPuLk8AgHIlgfnIn35G1F1irTc87i2RTANSIcypxY5s
DtkR/mlyGQJe6hffzEkc4VUOx38Kifsdgr3YFRo0xO6Mbr+/lRp00wcALkdpeYr0oK1yM4bLrOnL
SK6GBc6KKMnC+cPLXb9HNnLLVpYzX6j9zlkzgDvhePKN59qAX8yThYSCnsx/f3mQMi/MeQ7aYOkz
skne9n74Y5RZqIX67TdtGu5G98bIKrUIa9sBxbr/d5mjlEzQk7TaeRzjgwxmfkc/Npf3J/tWj/Lx
SNK/DsXJ3QiFI/jrcOdstp7pcAj509MkQKOXHFoVBr2OHvpDsDiHMHoE6d2bcx/w/skAf4DebZ7u
pjOmVkx+D+XlYkEmvVR0anhnHnMvNVypMTR5ab7Yy83fZy67CqEHB4VopGzGSJ9XMn0ppE0Oin+c
O2BspZ0VLzUfCDHOovteVvJFuKK/7/o4QrbEXWvUk5Jj8ZLAkvVyagbHQVLiZH/T1J8i03oUiXD8
W+9M8Ap+jTQtvO0/gemsTmhV/LeApoXZhWPJY/+S568clFzQVEbv13APUnLsMRNWwmaCRyM4TbP/
lug3RgggsQvHG2WAjIzDsazd4AUh4j0IzCQ7Uvadhb7bhyjsXjxzp6R2zpx8SmjqCjS9MnJdyH9a
AWQaamQ1+s7TL8yJgKEpzw6eNmrf/2ynR0Ydyuonhajc4s+L8AzYTze2kq+LAPC3EHfj01I7Jx55
2A==
`protect end_protected

