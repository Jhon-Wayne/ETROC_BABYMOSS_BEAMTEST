

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EsXeRsPajYX/YxoQaWaSSiCwfBR719VMFy+WbPGh2UU7Kp1+dfK2zv2NuQUxEGnYh2IsgOHOYx/7
4D14E6T+Iw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fwNmTuDBeFQhprdSkaRvfqp+4JN2uTi2veIKP9lTdMi6V3vFfJL2e26ZwNopnqXVxORqcIxB7j4G
1obXJPT2WSCL/0R7vCUMg/xfDg6ZfHRQ4HvE6Q1qt2f3x2eHE9gwy6LqEJ8d1O5yddIUz0vAxT3E
MCeNfnm0nCRZRRRR1XE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kL9kQOh4E6UtbQ/npzD9A5qvkaHmW4Q5TOqEPVqfbEiuDvKyIkPxWrP2j08vuQIG/7EyOqE/kj5s
ywoJMmW22K+cqgqvRYX4CWXFmZSBkvNI1XANVHol7+tm1Q6zcn4x8jo3f8GnUuBouEp969uv5TVb
C6W8kRmH5VAQXDtD7qgbVeYKswRn/GOr03sH8N9Ixf3ujy/rBmCmzDHZAfpgrSzHpSBDLuEk/POo
Xr9RNXhKMiY0o/UKBWTOczhocmLcg0NMSjuIOOn231vhyhTbXXcQqDAcqV0PuqZO7OgMM9AUBcta
f5wQBZ3NAv31WeWX668oqKgjV5YgAh+FAy4XhA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RtCEHK8hoBVXzxMIwgNIEMWUxUkR5Pqab6pK2iAMH+eKzf39R1Vn3oDa1Ljhrvx1X7iUngAsgX/3
LcmaDU9gqDte6ddNPkmbNLHvLhT9m5FvOkIIYEvIwBd4IBifYnydM1owSggUGKGtS8XQry6CERrW
2IwC+w9nzwdB76vItXdw1s4IymWgY5uwNq4//tpnCTkR/OMjCa2f6M9qEfWJYNlBJ+GXDAJmYmUS
wk9As7MfL7ue/D71kahi5ZCHlR1I+tDM5txkG5hGeVCdvwQTXth7HwqgDY5sYW26p5uvO2ZqvlfD
UgWjG10wynX2xKhSh6d+19vsIic1nRD2zh5zJw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
R3wbUw2LtZKD3E3fbP2KygA45tQjKS5V6VfkBIYGo7BlcceQkKo0rH9dIS4uarIFJdlyweFapK4J
ePxAwMW5ynwhut3dqSMsEu3D/QC2USMsVE09S32y+GwiJIOKc4yR4T3A+F+DpWiAENZtryn6RnBV
jZ6etPI/ggwkkZm9cLyFuFK1/x6BNvCtmDYBz+NvlP64/yJ4zISqL2xL7EkNUjtPoWrn0H6hwsMN
LWmwS1HAvRjP69CtcKcn/ZrOsenLSCoE2qMOpIL4p9JrIN+PO8HJDrOUWtQU8AFS+CmCXdRF4XvA
aw3d/kbIocHUShnTob8znWjsVn39/MpEWEx/5Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NPgqApUBvoFW73rFSKf04YnhBIrA8CIHSiW0X2nssipI98eewlp5fI3AW8Y627oAGytBSN0EzSw6
6mWHpipQLQVJA6VeUIO+8/hOLRzTb+XgsgFpVaE2fLeCPOj0g3idUo0VTbgU5/uqesDE0Vbbrta7
T5odN3Lm9NJkl26/v5c=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ejAJ2cG07D83mzglv1+hg2mXZeeRNlGMZpMWRYKoOLgMgbw7dHfDf5ZV1yQve7ZbrKv4ydzeaMEx
8KfLuTCue4KY6+jlpd+KL0RPlmYfM6m/B1rwwR5ILj4xN3GdnDEXXsiMW/kLFu6ZLoD4Gg0fG+Vt
XWxnZfKM0dgbJWSRVoxq2KanJ2PlZ7qdlRIn3DOrtTjcJYuKzzGfxtNYdsTieTfk3SVn5bI2qSkC
3ck6p3do36oxO4wtfit92yihFVrV0gxzgLHMK4c2SX5FGVkm5jB2zgUjTl0KTI72iktv+yeDkEkh
cO+wtpTtK7QSUkTWzCgR8DX8WFsIX5CNO6bleg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
z5d7FpSJK+rLMCshZ/iDhwX4O52NXk0tJCOUOfHVwd38PR/4BX/ThQQ7LwziwtDAa5Af9dUoWjlf
wqAgOcW/fMwSc3z3jNhu13J0fXP2ZgRc8XCefU8NXQrtGmHq2POa1RPg8LW2jeYMf7P5noKPQifM
B9RvAyETjSmJPW6ktrre94fR7ktcDLgwgDDlYSxx8Wyi5Gzh+3EqCU1KSfWUD3z7kO5Pp5xvjFsp
BLkKMVcn4UTwBds4EUCkEdMbAmUziXnuwBLvb0t/vTGZ+MLbF/z6Rauw619SvWcEKOC6uXZIUm7E
wdJdo+nnXTS2RiyAt5gyZXa/6Vz70Lgbfo3aJKrKSQi2Y80hdRVRhrC1ge6HD9+Wg54/p7yMxZpY
I3tfhKDckC3Arn3f8sfi4W+mkE2mEqeG0dvMS9TVWKWoIUyDd2nCcV3mZL6JlGTYBIpSLlN9dNYF
kXZQx+3lGljieNIcoqJnu/k4mTukVPYzwX3WFqHD2Yop48Oyb9S76Jdd0dK7q5iC1+CsticGG7zi
2q8+SGZfIEMzyI+Cm7fxkvA1MZ5fU7Vfrn5u8ReaavxJ8RsOcbcJMUtHmbwu6xY6ZU3XnGw/NmuE
r9WXXieq1qoTRMYow40Q4YAIf6gn/MrJ4sgLlp/9Fv4arxxLFBGFsmfqFtQFawFUmy2ROZdqRnGg
YiD6e1fwiWEewNdrFO4gyj9i8StrM7JRsNFYAXt8m1+Waaxv5a63W1wCGkWxgoXcMY4wna66HXIQ
qGudutjIonqfM0bwPLqoxgZ9vWhVrzMXwP5vjhwyp1XFgZhQ58jf3Esacs+a3BDpKgQ5hwAIE09J
XxdeLig2DZ1sNBDOxYbhKZptWQbLzjZBU87YgKKqGDsAynBTzWk601b/fMYaZl0G1qAVAPjscIFq
/GxHykBwlcrYLqLRrcd8vs1jbZM4ZLVGRZ2NDFIbOiKakg/UfFbyxIvoGN6lqzT24sFokm0aCPLO
yefHZiOS2X49VUlNk8A78CyJWeLjw4hrVZEx2eALlgYm+EFb9lwjm8ci8SOmtzZ9KYYRpkCPTP8r
pMScoAB3PUFixpeqNFbDFnHtKrp8lORptjg2KX2bJBJfH9qL5LObPcBayTLPVJ8RmQCkpYKk4ugl
tFKgGCQ781w0li/zIzfVklVjx+rwd2a9UjL4VRlPGlkPbbYlO+0tSddkCgoZ8z0U2YEAx2P6CKHd
ssq1HXct3JaoZ/VRIHdG8JJePXyuaUOTg42cJduu9tnC+3Kmw6KemKteQSOTLNjU7RAKt3HctRe/
CQ0ycAEXTxnNtR1WrA+nzJQUK9UYR4Vfq4MzRPvFmQZ+V0601IVxr7rMIUwc3MKFZo98kHH5olEG
jw31CvNV7Yzp/5ml+/92AwxgKH6QLJ8drQpQ7R6iE67aPcS8zfCtNfZHHi5fvjJUu4YwrP3DWqJ4
kebdNZQ5xaMJi4gbxNyS+cffmzScYWC8fg5o9zZnIjtYkNcb1FkZPhv5lDjsuQX0KupuvFs83BLs
upJptTwZf1JLZE4C83/dQmZ2WrrMpz0DlZQND6DybYW506qogKIiGv0R65RngrX/nz0QjD8oln/I
OZkdZFtFBi4Ut1ox7CqhtPepOdjhaR3H1hkynHM1CBN96lmzcxDlXFeInQTRENAcvmlLngj5PHRK
VkB7krGBfU0jWRKNVOL38+zCxsgFocDDBDT0WDtv+OXFPf2kYgiVk0arE1v6K4bCbvigslrd2fAD
+EI4BFCPQp1HERUE28zzR423iFj0anb3ufCdhmu+8MFhqoC+wkaSmmCxlP/mN81syfl6+8pXDfzB
NwzNOA2HqmZWFhJFRVYEVJ9Ssk0bQr2En1547FIkFtlRnb2aaXhbKH95mZwZsebgmoQFce9RRQ+O
8OLG2naXzCZfjPDYVx2zV8e5AFCIU/DUZiQdNSEU2JEu9M8CToMqFbkG7cqcRRLsz9+TC1mSFrJt
m7Xeg4NoJQvOixaoW9e1UiLwnkW/4Vzl5Yqbg06sYs3vsf1s5UjFvBwk2wS3pRtCYL8C/XSnLNqQ
aYyk8xx8vVlx5uJJ0U5cGCWHKhekbdv3yrVOLcC6GJTj1oX46vICw7xzJFwLYZPNhSfaN7185r77
zEYMxexUjP+zIrfW0opa66FJ1sSv3i+oKoCU34oFoAWBLxYDnr4UkDTlBeZBTzueleeGBOFm3ZWV
MuDG6bf0Ul/EpygMsPlDAMyS60G9iQRUeyn15HAmsUyq9sKV/rvT28FErQTVe85c3L2ytS2vSw9A
BUJi+FY9SsHloZ/6lrDIKmudDW4NCa85NEcLIpL498sdI7oSHi7rfLFkEupy8nDRr/Vl4Nl96KeO
VqSn8uJ0iK2apN2uxBTHpTjrZROYQzw9mBL5frFWE+lW2xx8SLXpwi+uDzS8CanDt/SkKs8WFpqA
oxoQk0yrJ/DSPZVOYdke+xDaDN/qKOtQGqvhMj38pRrLjMMaiMlYMAxbropmF7kuBEM+AidlTcUh
3ttyoZG+lxAdQVZMhVLHG/Cw/DJLtaTV4JjyI5LPLUKuash0wfBmkOhzAWuNI9le+/4UMtdEzPFW
3yYUWXTLv3/uBERScg+kQ0ILn3GyYlqUMWFrn6690IN8kchxP+j5UlM6Ra07hHutm1RF7Sjk1qhF
vJhqIu+JvlbvQqGi6uoz29Lx9aSHc9C+7JUC85CbIhFDWbrBqdZvLwTSjwGwllqGA13aM6S7Vzot
wBoBqq9xMrqJ2B54hqNDcYJBQL2xzQpOG/+RUo/SDdCrcsQEuWVdMrVPMccC38z7LtS3gcCXkKhr
clp6Uaa1nZRrQAYnh8QGyyKZ4zTeODFyQ/ZwOhhRF/rgHez3tolPRoSPaJjrIlAA+PHKGlmxV0be
AM6I2MFT35e94NuyHh+NXSafUxzBgZnfxHDEYcQ65aXxElhKIYoLY9/TGFR8hErQHWvcbgZKMOb2
5i4uoKLNzmeVT0KxE9qbim4P+tYwUAS8piRbY/264WYo+CNnuQp3OXVYAfAhkwWvvfASPn9Y52wj
70mSCrGnpuXAuEDQykYYmvvXl+xIIGzL8wu8bMyGJ++xiTFLnNpG8r4AGBsjN8Bh1Ozeb2uvI0uL
CuLcP1ywFFkuFjS71kK3DZt7eYEh//ACUh/gRYMtb5KoMDr/x9BZH2tYPNrkWOYivbC4QRYNW94c
Vmx1y92rCdgW/Ja2lJI/riqnM8cExjyEI3x6BSlJ4TzYSBQ9tmDnMW5bDOS7IlM8GQFgXsAXbV5B
O9VhKVKO4b3jvw4J5iS0z6mnKgSob7+JaTjbDHHq/avVLtmwckEKqYMbfUh4rKGC3wB3NkRjeQtk
kNVx4OeIBy7iml7h6OWSeF4cOoBdMyJsTXQYoHmNJrgQ3Sjh4Qb1f2YQFDO6SlLm/nFbS/v7kic8
whIBiK5aCwifeDH0lRRsAKu8EF5ZdPlnWSr3HJ5jt2MY9kVphFXy15UpqXvI/aEQGdWs3xftclmw
vyN1cKvMUkJHXZt1x+XuoxaIVAFQg6nlImfff0gxK9+dtp1n0NU1jN8b5HR3rqZy/XzJYhhDk62z
kO7lQqq5AQGHmL3n9o7PMiRxJn68scJcHFgXmWb5zcWTP/BCjTaVS4+gLxbtPsEmXv1zXjd+Z8PC
byHzWIx3I66Ost22HRpI4Fo+gW2z87XrPNC/0umOdnvoP5ikQ7bENwhcQU57OQ8LdFCchKqzk+LD
8UIDVnuHEd9TsocNsz4Cq0Pf59OP5dacvvr+BfHLsEVV1mAzv3TaSoxMcFD+QqiQWLONX5EaSq77
efFO8ZfsTX/Iyu1mY9R1q8/NUjd0WLLt36euhnfp/RSHy9Ddg7oIUFVloEQk6H1l6PpInJJyNb0R
QQJopEpsEPL0LClzOCbA88LdTS0LTEudFl9VwPbFgjLsNv2TJ/TIjUgR/kWCFsu8sIVeiRkhPlcT
U7A0kSxWmABaNrkq8Ge91qj9Qy+2gqmSJnmECsAY3KK+2PDpTD/Qhps91MKIv7Iu+futZiQJz9WN
y713Y6frPLYPDzz7CHSvSPuiK3Z5njHpZXGrk2DuLDPC1Jr/gw5zCr8e0ZOHctj3p7F8SEQimJe3
uOkrRFZUM4h8LlbYUizjcHV36Vsyvw1r7eEl7LBrEak1HHX5xnn4Au/bCoQCcZpR7orZEIwLOz+T
qOiXF4CVzFYyWjGJmYIFYMOx5yQ/PGRarhBtaFpUTbR3Jm/rQzUVSGR3oGLa0T1MzhYEKgwDGHXH
maSWMNiQyHhv+D2v6EX3YVWcMLXrZeniS4lWnKIXYWk5lLXhQJq6PZeI9ODH7td8r5not2srxleg
fPPwKelBnmQDEaQqK6CnUf6adhDc42JOdn63pPctPjObRbY4WdCZ7k0xlzEZS83q4xNOAeyvrzSG
RSAO+aNs5JjxHSq/zeaxCquWuQQUulPpl64HpYvR+cWcP8fLfK6vi+G39Rbi0kq9P+xBMBp2Uhv7
vRb8ylsvsCfaSo50pfBX1EtpjBWlljgr/gEBr3FadMhhvhtweVCGL2n1iXvsDAyUNMn4/TvRa/m4
106ejvJq1vKJf3Xv96Ezg3lOy9NjpmqJ97ddFTRNdXAiGQKNL5Qa4M3CAAkMIbjmMhJrigE1eG0y
6AjPOGUd3i5sp3SmOBHjkrJUK7CSxQLqRqXZxg0fK1FUKiB2QT3IUEJLK+EhXtzOHk92BbkgM3hQ
oKRNDjFZ2fWhZ5YulxQsEGR29j1mkBTCP0Lx9DstP0BQW1CUhMWGZ49QTZuafcHSzPR4/YAOrX3k
0DuSOSwlH8Aencq8rmekFzuS9Vqt+nfODWnx1RFGRlZReWboE6ohNk+dmacXO5pr2Up9lLeXXK0k
ajmO0HPuo+xj2NadGYTq9ZvLJ4Ahp72QrVphMF+9uXDtEGXcRTpkCgjAo0dk1lBMCl+jMc1x8Kk9
BIAfhgpEwmfHVkJGm3lUP0NpKfdQWelYraO9DnC08CJXrNYYGjN3UBbe2CaIpAvIbBfUUybjUPp7
qB9mFLE21LdmDK7aux20sZlZQaxWXpbUq0D1PPtCo+NlVdX3j14iXZMLOpgyuorjc/oT8QZ5lOo4
p8TYtU6uxW9LO645Q+4lPa5xZS+EZnHEBRMIRafC7oLvaX/Nwq5SWFXToC8MjRcJGO61CMveCVGr
j22aofU1NmSK1E7CaxU60g2g83MbivmVDnAZr8wCxxhYukogi+jDvC4X+xAQI6+mhDYEOqiTq+wp
077lBF+btsJj95GA56D0afqNWkG9lrreaU+0heq5f+V3GFjIkukr0JE97r/E00zDkDFk5XAIeV4W
UaeJJtidc7O7U0U9DXKzl07gERG8qWjlq1xqKCWBP8KmkC0a5dIp1VP70MtyL3ecD1KeYT9B+9yF
EeiEHj9PSgx/MXj5h0GG+QgUmVmqWdcRUt+dipBzCmA+nECJflx2WmlOfsuO45cQ87nEwfTX8gSi
48QF1NT4bpd5XLF6USXQiH/HUQGqf4R3oIdJVIPSMgSlbM0iaPJDQV/32l5qeI8BMXKzO6TTumFx
R2m15mmnDayzOKBPH5aU+YNhFOt80THOxVQPu1AvXzNqX6CaqUJYoEhbVY6aPKbl28vOkGC0L86Q
mO2DlmCpNxU435Y0/HmSa/7WeW8a1zFRFwB8HXGZu6EjSDzRTzBEphCh1BfBaQ8Bmd4+AaxzzYB2
UAnwFvbo9geFdlPFo75zZJuohE0FpsfYCBs2IOgu0ipdrYtHNY6RSazvJib9XUC27CignVb8aA6Z
xXWQA6AfV8uGC9C+SfvX4MwZtROh7zNEO8eySsw5k9AVMHv8zVmZJMk+Krui+CUBXwOZ6rXbTDGT
Zn5ENR+TgbHsPCKijcCfcSl/b8LfZwFLI3OH4lwyXqrvow/zizdS+lG1Hu/GCYLI6BcNuxvWPNiZ
+MU4TpXziolTPSsloV4oY/T5w6qZjaV6+zlZn2wxjgbPOqsZtxiPOh4UjeafRwLos22CPIJZZZkH
EwM9T3N7QqMY0bNyNf2k9X6irmZUW9srsHq+UIBoN4gNbp3RyoKl4tCVKLfYsVcjHc0j2IoGnXA8
yXMgT73inKYsG0c5ll8dcw6l8EyPSgRkh0IJoVKNtvu5lA47A2YdXPVTd/doQrp+/c+vhVC5NWY1
E3Dqbv4vn/HcCO+/RyaL9rBXte/sqV2M0TDrt+967/mZA3Wx99Fc8vglSCEkhoQBJO2pXG++rMRE
1nBmOW/81lPefqkkXQM9yQ/sbTwmjmBmeXwyg0mkZgphZcWj4I1V+ANrK0n6N7ERyIPv0udefrmC
AQzzyA8vZ/8i9Wd/Ecnhf4zXA/If3FQsvqLzl4/ZdLEpJD0KqhCNgbOFM6/X6q/svd2DNOZgoRRx
JBHVvOXaKp37x8Q0JCbjVEdu0100dLHgejZvafy6EtryYgzIKgNTzA3aCxD7QzEWRmrTr1BTshdN
+h1Iiubm9DdFkM+Z4L+1GWZo2K/rNgh/TTbKEJWLJmwlQWQUT19ajx0JYDl+G3uxTIUXdDUPBHCK
u33X/02AyVaqTkmPt+b5idnzw5UUPbfYlwDgzAL6PbIF7tz4CQeYESCytiyP5CdgUfldBzB6TlKd
NrAVD4XXhLFicbpgDN30RGXz8/HaagLil/kDjySBZdWrqaaacY7Iwe170U8XvUnCb1inJ0dpd4RS
riJzvh5yLGk7fC2iPcRJlU1MwY5wLSvGlALFOvinbbP8LaeP3aWrhtjKKCYYk85byJVOEG6dlFGb
t/VMCmQQ8tnpftI9RzdmvShws4Y31+dDQOkPE+m79UVPppLkYIK9sdms+c7T+JY7vzOP6mI8SUhn
P7x+5sjm93lch8IB5QPnVm/ClWb4OGYksrBxn2lVEhRwA/iXsA6ux7si8Aip8S9KF1HIkoleavu9
RQJGfzDZm5qSuGVpsdQpyDPUWxkN+hIa1I/t5zIGuqwmo66Ob0uR7lrAoHm8e1D+MEvFWr+jWpcK
JghPjnVWSPNQs0bEK2B7OPYP2e9WnKnGk6Xe7L/7HsEV1jDrnwyBRuOv+vGUrEDci5atGrZgSHFB
UGp5jURpHIPekd11SqIbo1nkSlexfier+mZBr4kt16s6k4i35kcoitk23UglhUBKEefBC0rcGvMt
lcrSGXOEe3sF92CSQpDKiPWeSL0DzLWue3MltXXXbjSKBpAcPf+8U19QIbuLj+YF8OdFxzCfP+fo
K/qh9nQ1JG75wYXCV/+zLjtuA5vej8ZGlfPLRH6Weq4CUUP4HzZhbzqP35VV4FXEGQMeP8/z0Zh/
fGhF52LJ+2bnE/lUT9eCV+PQKElxPrkV+Gr36dHj8PiT65TF4ntKB7QtI52oBVE/miy1UvTg/vAv
0TorQU3jp9uQliPHzdiyo9lgiH2ylxKwgGXLGn/emcxgjO+7lMV29WTKUzlCM7/wzIABbRFBKbEh
910QWZPLl3QhtqciIDKEYZzMngJjGoq+4bE+eV9MX4bkdzZ3KwlelboJIBFsOkNBFhtPLq2GVtFx
bcCuQzhxFo4orn2F+Ey1MM3fgajHBcAeP+EWxhH15k0VXxL218JNusekMCkNQzX2LRwHB0TIzjn0
bEdiRZmjY3GkobW0RsD5se+7lLEnAOP8gYxhZ5vdNBAuvN/1nEnemRy5XvFo2vx8B6KNNCfcIrgN
wekmzQA81voKSYvCKkKCK7n9WyVoXWWSNAXQKGqFFEgU3sccDowPKhGuIDAk0464StWSrkipNf8d
+e0hNDJquzOQbd9R3pnDBX0XLeKo2XjpdGO0+LofnzTnuRliLKHfAtLYZAUa0HB8XE5KPiL9OJza
VK/Fg07VRTXszbIGogJGDI5FDKSUThyUi8pw0NEV30Qad4sSThG0PzoL4OQg2rn6JtMDJhg1Lm9Z
8cM/1dAORLBCMQN77NiTdj7iMZLeUVbJsAMv7meLd2anS7zLTUhWgjlxkNqKkMLT7mGFhbh2vfab
rdBsNT9778CT+LFcaZl+LWp4fGqqW+9pe/vyw8vP7StJmFAAvkGjFTNEFElxqmkkiEdSe1MpD4Bw
xEE1CmVRwQDvOTXWQubZzYEn8DImoMygVthqsK7Gq4Fh8lT3vHLKEbUCIy0aukDkMMf+BXB63f+O
yZWHD7m0A9KMMe5nb9KcZz1VcqP3BbIfSTM3KA9tfdVEwaiplrYyqocsf+EKQ8O380x1WqK1+JA5
jWrFsEPaLwnDFioQCg9g60PV5w+JxU8FgcNDvziIlWHrwjY8pk6V3RCCxyBWkvRfMiFIfjW5NEzj
RXuV4jHMZcqEAoq5OJGfUPh96cIp5F6clEL223p5wCNozGpeVwzKvTqY2H/b4SUyk91/sL6c4Trf
v08upw8cyPWZGebetvj72cvAljFBoaPvjk7YcwcBapzIEkjTUsQxBAolL1Y5YfFY/VpKFCljLpwo
nJtKR+sLb9aM1wM1qGJS5C2VclLCOcEXJ29iQgzUc+kWk6O7n06cF/HSmASqJtC6viXW34F8EwyC
RyCxZl7J0keXEtrtmT2255eajb797pUBVXmU8AgUp0hBNgwxhHA1AYlPfMKKYCCnojkbfrTfbJzw
7yk7mcMI/kuwkz0NOUPMZx5soij53vJpaGHmbceQ51a61rcVkA6wyIMCCXy0yW7jbpqyAxiWhP9j
Xv77kbXbwVfHNWmtBSIv2T/myvL9aREpy7/asraa4vsHnH7rdgVDpv+QNWy6hbp72hnCUUTSdD5O
hP/JeQZ1J6mR1d2JWEljJa0CGmdwkObSSbU14am4qiko5ZUVG6MVDPStC/7XInsmxL1Y2ow9oC2E
+EEzNWCoPtYBTh8Fo1MTvYMDaA3mRibf+25T+CeWqLiR/sWssrBaX/9Tj1SCdy7SyUewav/RWN0g
MGOqFnrqnXSjkGHPVadInnOhL9sUsNbbnjccMnyxzKL8Zd0A9d9ZLygVcVkrKqfqYhos6foiOULu
+5LHJGRUItQ3VrO4CXJgSZX7gnFd+LgNoz0ia7OVTjb/emZ/35foztxsW+79RSLvxeHL9jhryN6m
ODGZjs5NWkLW9wWkQEIJFl15l3lASOkvA1BuylVMI9Ne3fvqYdd63K0q05uruspEWAyZ8QHa2S+L
3VEVsc2uH8ECSWR22Dvnc1NVKrEf+wCFzUoK5ckB2m/UTvg1ZDVdw3eOYuBPf3GdW9QVvKDK/Y4/
vSUqMkQmYIH6+yR0gv5rzYOsHP/45Ofxs9pXJAzwINhx3btp7g0LW43uutZaxAbWxg6khs+6aS5x
b9M/GrBq5KBayB+MMXM9K+/3bCKhKYzO/w2rLQ2rLnYwo1Z2HJndLCTrIFYUA50LVbJ9R0YYWwGR
HMh5v3UHDTTLmIL79trPXN8Dp5pj0+lE/oZXgrgw4PmxwDI+qXBfISC6X4ygD1itfSaTs5MmJd9d
Sk8JCiHKyxXjqjM/7J5KyMn7EH1w/3bdOYODIbQ6jEwYU+f34vL9mGMJYPxFjPUGlZ6KYM/qYG53
7eTiEAwNgqzwKQpMDWS4AL0B4+7RVC0R8FIrHj8IktsbbHmUQfvx7GqoWaavXQiLZyB5pl6YaDHz
LhGyy0bavju1tOY1pgdD9Ybkmc+Cg6uUg6oJarVmvLVDYxngEqY4uTBBJIQi33lMli7iPswV5gGG
+TigMhge4UaSMkCDb7ImFc4N+gLESywiMhfO7dLY6zQr3PGN9MCndsqENGDgYMeSNFDbkN0/ZTeQ
vUCtglCYzNjuXpEEo0H7L3ltY/gVBP+689W0KN+3Bqv1bLtH3xM23rZwLMdSK8yuSHJVDw5zzHco
KA4CzXzm1uxg7bvNM/dYdJLS63ZwwpwGcnvlcg8M9WgjPhj02PYMEEKt/JYTOKHTo7d1XysVr08O
HScU5WJbKBYGbhFGNeCTZLiiFk+zj+Ng/hg836VNt6I6sFF8yT9FWChUVW6lyD6FiG81riq+1Ms2
aY2iNHg+yH9H+yGjqk665G6RNI2gVYaWVzBwtv+iYX1D20FqKl1hM9vwRAbycRFHcEanPBrV/S1O
97psGpx/0up/lMmM5f4MvaahDT7bu/mpawuTcYOHc0GXt96Jwt8ZqMMV39LP6mr03ZRUEK/ZVi3C
L+docNKV03VXfeivjRtSvhDMp0zYS/Uqb8+/sd8O1M47+NvVJI3qFWvPiOW+hHAiOC9hcnEoeq4D
Slo4WkrByM2OMesLlxl+jjjB3S5ycWHN2Fs0WYZXml3ZmdwB9ClzKIfnKA17gNNHQupHQvqCM/rO
Fr5F0By9P3GyzJ3HnLxuTw7fXrcGrf3igEyG9cUDYKterLfO4K4/ezPe9TKcHM69ozf78xNi+74d
IukX9mvu/B7LY7ac7QAaocFrllPK5mDCVEOfU8xKWLCPlXvSuPnJ1gjjms0ESRuGtGFDSYcSoRFY
rTyiZRdQISP3x+8+SArQENWqOXAI10bDrDVBMk4KNLX62HRaU48OGvvpgxptNKyISJs5AYhgxsGR
bIGoQVgksp3YoTmMOsnq85lAEqicwAzeI6XzbLlENkKOJPtSlNPvD6jIjyQuaqaSC2K5jklvJC7w
shPzUOYdHGYaj6cX3a/4ZbA5tgB9Ecy5alPES96EMEQmAdmKKWUizDGLgYIvJs5pIf0IbkUjISvu
0udzNt2vjETy8wInB0kSzRXNBompIn1bECjmjsrfji9MwxFVjxGnK1JfHq3ugMcqeD1iwTk08eCM
naMgm7vVFKav/MaxxNxoVycyUgfvJswDvmj5+JeROT0kMR6tXg+bdXUeU6DSHQyqHA12mwDNOvV4
K4beYOxSIIV8xV0cEavwENziUaZG7FMWHxaNmjhSTfyvqdy57PaewiFdnfEY2TgGEZEvJAbwPgmO
3/n0ueq9Ulqt3bQ1tjkrnHDkDu0ncUziPDg3HEWZhqyv4y+savLRZo1nqQJp7ASlY6cyvl8SPoun
HZq+8+GHXbnPEDGSdSOaFRt4MlcJ9pBLRXraiA6H0Vz6IfYoel/JqmqNssrx879ejjoEoNFaY8ix
HShqVTF0snLUCxCavVjU7mbMSc9Uy3lgwT8DjkdhJj4bWk2esHPegK9Vnp1bDIrGe9QLq+55B9r2
e4D6exSoCJEMuvI6WRr4V3bfy6e2ewrx4ElLTrKBpowUWaW76hNkhXMGqUKGc3UzPW/+zLBC5Gdp
0+VaH4Se9Sc8nmdGfF3qPLE7pK7YqYjA5T5wDIOJ1+vDJ120sWTLqDzZ6fRsv5P4yW86W6bznuzG
WhdutGv70WwIxPgjZ8roT8XA74KcJrW7QHBl2VSNh137S5DUuspz2cH1M0d4izpTiKBbp2wXxm+9
7GO0eGd/6i3/WKdzfGYuKjSoZuGs14xN5TULoWDx+xPq4hkxa6BBkk16SFGmKFGLGA9FfiRMPl9F
F0dRrvIfDAvPm8Win5c1KpRy8r1Pt/yKlej5H4xGkoW3zMRr7lgRI6UNGDpwZVyzW//YUh0J9eZb
1Frk/aq5miPpe8kdipNtUWZ5FucDW4mJL+ndv87vFrOSY0E9qijVA6vPaluy695pqnBo3ReWQ4+7
BISqfL0fGGc7vHZIDYsvpkxBAZ6mTY/pyjQQrdnRVUpe7Vo0cEyppLl5Qo7UN8Q0GlIz+9VbCIw4
HlQBxRR2ZFJMQ6U5cgjv96VtfoPy71SYHbNBKiEju91eVT8ut0riPFtPHjPbznGPJpLGnnmDdm73
i/iopQB9oA9X/XP0D9s4zaoqstzx7y0TSnNRf5QDT5FZR+QRkwNXAD3v4KSC31c1I47M7OvR5bEH
Ca+iOdTRWuoyTZM0vZlcIi/l/Pt/4uU6Ynpo0wWfhvWRKS4DurFDzq959L8j/N820iO4cSazLs4S
LqM36eBPs6BYI71d8qvh8Fil9T6fVxA6ZVXJNjcKrWwal8n8GPT4Sz8OfNNVULLw6+ELn9h6KGTk
Wr5j7+evDk4AfCuX9avpQ7JU2/Xgjk4lvnHAIuM96ErP1rTcxtZrj56HiZDCNvJYa071DyRdfDvm
hVpqXjMwR2UdKDQtPKbBIYro7w6Z6LbZx5mZPq8yV5WMj759WG7BWxUGFa+TDc3miG4hDj2zdX2r
okXRLkoVKP46suPzK/m+c9Zoi0UhiHsi4M8e9Jfpssgm26+uToVORpJ+63GW5BchUOI4N/bJlXEK
twglAQc8s7AjSxwNOAl3QhxESYX2FrKkwAx0cpzDaQ8x4jVgqmeo1bQ+U0jBa2DXB1HGz15FBJXJ
fi0rOStEWpRh/ymwyHpKsmroOdpyZBIKi18br5UMISYGTy1ga08QI7Ds7O1tFqshjtsEYfHyUNbP
9UX6caMCI1O0wT+F952ep8nIIskSkq42ZFvfG6PRgmA1+KUsBGjdzrriXvzC8Bs2DgA/XHG62ncL
Tlck8m62gd+qttKfco7ZydRfaesXWKBx1vYY8D08uH+5VIjnZVQETLLZv3JKDw3a47PCykhcFs2W
v0FxSsvjaq780TKP+yq5bX/6gtw5i9D+UrkTu/ntEXXDY1WN/TCXR/r6hdWZllqpZrZEZ2hiJJ4A
iJuNc6fd5ljC1XV85Chis4IzZKWusSU/hY8XNXLCisyj0x9y1jTJt6RriDbi/zlRzxp8OJT46TLL
97PyRejf4yVuK6DmwbU6W/xivbWkWwvmFzGxcjn5uitwWvLB2KjJqKT2XjcvGLIMa/pTe2+/KuRJ
E32pD6C5/tRPIfQeztMesLPClGZlvTY2LoayxYYhMPUALqLmP1sYI4wSdS7hsxpTU+2cCXf3PHOi
n8pxn3FKlv2N+6aNDNDVHkcSmIKT5xbPUS6nwifCUtt2mRmbPOuF7skMbTeI9splmPDDhsFaLGxG
+SjUGQDmmZTLs9yHZVnmXCFHPB+jp0z2nwr5paTRT5P5T17CDqChs1uojqVjKz8epjrlI5iSKv5C
FIsNoEZVSjCd1r6lQJ1ESXvhcLMVQgliv04ImiEubzHXStJfLp9pCcq6hZ1zulVfAg5QEhbob21M
CTmTnjlnrX94xiX8mNV5v6r2W4yVoDKBoRziq60mIlKqM9CyQ1839z4jR9Hg0b/7Bj3fe3I1Xh/T
ETFeTRV5SYthf+TXYnonKzHNJ7mubNlPgSHeY+ZU6KCZpL5olhPAtkUmhbvBkr9Ho9IuomM+n7zS
DqTC26vtHW1mYsKd/6f3Xt/Dd71zm15sCMxjKYK0oOlnPydsf8Z+TOANbZPIWjJBauNrlXj6cKqH
9NVvLXrJowE1nTI+n37Qq7mMpWOyCDuYvbukBrsSykoFRrazNsdto/+7REgDearGhpA0BO62obc/
7O8mLYiLB3aGYXOGPMzr13cAzAIEyjyvpZ41mpcadkM1Q5ezQ77jsjrp2wqkjC+J5hy0uhgjrbvT
OiKqESDecdZNENodKi1C/DDQJLpLPyPyXNtkp2WOaxiChQ4K8PcuUT9ngqshYD9ZHYpsV5NBzjso
Pqq+Q03hrnVDMvix9xI14zCCO5Ql+VRQe98wAkeIxeyjpnju0JTnWJ0rmvbQK8nvfm9m+Swr2g24
1dtsRfEjktbw5ItiTKav1WPfeMOMNw/WEWpoXV/RQMkzCg2GCqcR1TSvUyEH0WPg1FvxRPcVc00P
APEVRjBACtdt3eJ/1pr0CUfzMBeWfgL1lW6Z5M6jAmP0ysmehgQaN/CurMsoHRgQHgBLxT4fbGGh
UGotoNEsumTXLrQ1KcncKGgLjKZv2SdMhJ5HSXGtE67cR7K/AVsx1i90pMdj8lJpVtOJzgGoifIh
1F4bx9MuAgPQ9K2Oi6xLceLKYbK0UKco5+8OJS0QIkOzPlIGNtlEcMmfrEuo+fMiJUt+Y57gnao3
uyx627KLHJSKeeOb/DgQcTztec3gjZWqbpxVNW2uBWtua6irusZs3ewLmBqDFRHEXueLdmudvKmW
/s1rhGm6kqIwt+pyB7jb+iGxMdJMxcALeoj5MaczXVKOa2SgufHTeZser/nJ7QJgwlMMgfrhLAGJ
5KYVr9LQSSuyQiGbwFFsQDFYGN2gKuGpXGdAg1nJrr4xvQIO255CTibX7rPrsyz2oRha0zk8LNjG
e2PbK1OUIa/dVX1DuEGM+d6HVwno1V7EfrGOjwSVvdxvpVluOTRGcs3beP8KfAWLur6HcI7uH1O1
wTSMxSQlW0NWyoqx4XdR7mC4EswuIrzn/8JlqlRUKmutj524jay47pX4ZPLdIq+/ZOZNq3IXv7Yy
+rs4ElFwiFr0t4guHSFz1GDHSeZ/9G2hxLXnopNDlbvV6Kg7pqbdCzYGOjXXMJ8L8+SecN2P15oP
x0G7m964RSTE0jYjUbaEMhdjI99+0TPETG1Vv5TybmR5qwGkESjsH8MiiEDchCy1X8uRJuaIKQSY
eoomT5x4SS6AoqP+ArhUFmPURqCM1QJKqdsNj38uBrKuPeRmsMETy8+ex5KpvMTSQ7ixt1OGnQcB
pJyA4Jay0uLjlbHVlOEXjt5KvUKXcAbkvUJE9BFsHdH0TXvltOwae2II1Z3JXALtdCDxWclQORSE
FNnl3yFYxMCOh+x4wCh/1D+cKh9M1uxS1ECCEIscJIWW8Wy+mZ8I1JBRuxLXpd8DetqhM1XxkSSa
ykyvb33R+j/OK0vFeG9KPohsSVqbnMXjDKNbmQAe+0wDdz98Zl8iI0ZR8BZ/Ckw+OIKT044Cm3hg
OYw/WDpw4zCH5mb3gQx9PhtOm2cqTzKO5WGMQoHJR0R8bqYW6wadQ66qksXcjJcNM+1iBfIGVwCR
+9Mo8IVm+2uwbGC8uf2ZY+tqpAL3aZEhpr72Np/GRbc/B5uiP4A157uelesy1kmVhVt1HGrWBN4R
mc/O29Jq0cMc2MqM3Z9NQ3dO/bV8U6amudk88/bLLRyLIppoe0xdfUoIRwJMUm/9UHDeP4Al/ntL
he7W65g9A5W4oFxgcAz9VqHSGbw2kheyj2DjBObyxXOSe3V82slXTH5iwDWY2YceVOVsoV7Tm5/Z
JsZDPkaWep6zHG1LWICYDvhqFkMnvXl25sMwbIQdjk1S80vvCtFekr+UkwFb56q36Rk9CGFi8qKp
50ZRVsk8U4Zb59T8nWOa9koh3hoL8sftSenpYQOh9BljwwMGZZkNWSrJCp/tGkSN4/hMrEN+MvhG
3DmDACqPvuz2aGjxUsd3iS82H6KgW9yJk17MyJloo9M6pXeGofNSvZalgADvG5lq/A9O2RE+d7a5
f4buPROCJS4pDBtkOH1s8e7tVlCl+ATJtCaEt8GG1CbMtKMI+Jt3d28/psGmV+3ACJnxC9aoV3s9
KMGm3iGQFb9Ey89QcbtTThYXGJcaNaXfg9gOR7l/s9+qSMBKvHILQBjBEl6xoBcbkLPy2V3oUX53
pXBBCnitjPhXCsQQ8H+OwuClm+EkOsMDTowDS+pNUOUP0xT8wZuG2G7GrFPEk/W5e3BqBlGIu7YV
i51qjiJsLXkS2hxjb1ov7G5+D49lJMMTOSwH+2z/S4kAGMRGeJgEVd/Yv+hVoW3ZALVgml7QMzxR
DHBPLgX/3CCxlBqjmNiOeiKk085EEsNyZkAinI0gN5GZzR60/IHwT2MqESbAipKv3TrFQl6gZcG1
DYz+s7BJdew/IVWrUreWRSts5XMwMujZltiuzTaIgz0L4hziVACQ2tdbRy/ftn/jdubFtrzmQaoR
tNeMyNbnnKvU20ozRXcs9MygXkM41JIxkGFGhYDLyD5T3ok0I3l8ytvC+XO/rehok/33ZeBNbxq6
VY4Y3wlS/FBNBnrq4r4wLdPFWsjOHv11/jwAyOpa6YHmozCRGnc0ywjmkJsjG5KXu9BIA4uRTi1B
nXEh0pKnHJvar5ZGoSkMHioeI0XKnoDmMUyLHJEFp/wYuEWvWDvkyJwMe7PxZoD8q+bqhteXhDD5
mAJ8NyW4bmhMYOo/MQ5+HR1CGpFO/q+SwAmGQR0KhvnTNXYRgjCVP2zoOedgenIRpw186gyGE5JT
VOCeMIUhp4X+1SvLTo7m96M7vzvw606lSMvbcFacDXI9KY3aFBXxzz47XbRWVe4I5ywQ6YkPTdCM
cex6qDsvhtHTNaxsh0oGc4mMUfFBXuKVovYMFCVagRdTTypnZJqh5hzRZpKkkL8NsOAT33ATjUHP
8PVi9/FM7VDcmY7CDH1A32bSdpHbk9kWWtuwNkmO+qmBTrbdo42NYl928RlLShMcnbweD/SBCN1P
spHJx1B08Lt/uWeAqXCdS6BYPU6twxW7d8AOUW4cN+uV/GvwH0S01L8NgiCgxJynobhXyvQLwDXI
xYHsrPINhueOkzOZO/h289kaKR6wZZUm8xl1WZwbu+8AJkOpqDFKQAJJgLU2dNikk6CoD9Cyi6hT
nd8m2R1y+jezYJ20iVcsWgamaCQcEG3GIE4Tbj796yLFTSs9xOOy4k2guYa1J/IIChw/MT3GkQ1C
WAGeLQOhZ2AQyhVzt/G+AbXfdU+fAdbCywdtUlUFuRksbAFtcyVBpKIBo5Tc+rEr+vz1v3/OrjIq
rO0B6y6u2ecVHMz7vYYxl9fUt5jpt3O8H+cJfvsU907Ei+eoFoXSCq71z8/GZNnj1mEiG0IkZ86R
O8qnEVqbuZ5Aq4F6ii8gtiznj109Oz73fHchgTr2KMxuXMaEuOfdmmZy8pUeKi7VNtKi6v3YAoc0
RT+0nrzvA2rGj8yqGQ3QTKuat3t2DCs8AcZ8x/kRBSNNYKrW/7keoDD/pzDb6wXPjTDx2NYfP7Et
Wp9U/pv3Byb7oYW3hhuygKmVTbDVeU2Xpi/lTQ/VczXj1ACVjhwFTlDQ7EeWjwF4m65hTUSuNrtA
oH2jGB5fZ6AlpUKvOu9m5n8QyH/DoM+eKYotOJ+0MLvbSm132YA9RGIWZ5hwIiSI2RDNcdHyunJm
HRtVh6r5oYgfLlo3tdvA72TfGzQn4aXsy9U4EArVZXCU5QFrkRiQ2FdOLSGFTDnGLyzqlIL34QNm
Bl9WmgGXXcAPgwMZaccqqvyTB6pd6giyZZ6FSySnR76GCDSH1KQ3TPXwDprDsC77h98cQpItiDLc
jQh0R202G7uPo/9STiq+CJsYcri3m8U28PI7NE2r+nBuGi2cHKrN2C9rBIDUAfEgo8h+uvAoGabu
bSmzBGSJFchlPcbsHwDG533BubtDMM3yJF0TUKzSz66Ohz73aHzWXz8Pubgcc221ZfhejFYaWCB3
P25NFReIuNeGwullde8Y1KYiJ5WngRgDVctxnhfFElgnsE9q1Il0xxMP1iHQTwOPYuDkgjFjwkZz
pGBXQ5NmjXFW3v91WScO84/mA7sM6hpVOkutN4yszrGjtLwi6snS7cqeHE9CFCZrvgTO0Kqxh/CP
VbisFZMeUCflmKMTU69n3QgxvBlZO0RK31CCO6I9C9ipH5Fv0vsRAY/pnVf2XBnTIEDnFUmv0K/s
FksIQs7FTB2iyfwv1swCtgDgDY4Z4XZJY3i0plMqbFlphsPx3YrIioavdAcEogtLBzxVsfzHN2UG
1jLSwjUBC9jPm1D5IuzgYoqFASKq130lCfwyC7ua0lVhVvW/T+qnttmvgexutjyw+TqHR+gZBgsx
bB2f1UeKjcVO6ifJo/zKu/0YRpi71crCdkWeokoH6JfZOEmyr8JVzrDTgdlRfGWIpV9KQX1WnJ9w
h4dxcV/foMX0YEMR0aH3uu0Ab8q+WesRJ6ATG6q8cL/cIKpba7vK2bzrw9SEIIogTASM1sTGiiXa
yU4IZMXp3jbIZd/WFH28H133/TFDwzFN1UesKWrJwZd8V1W19/c+HVzOBrj1gUOPTeKZx87Pk35a
If3RlGkDbahM7UzFnPb5xCsOdue4RSvFr82ntHWOXQRKSJq4q8vm6chugT8y1FHWraFXXIsyzGcz
topL+ei2qkVX2MQEN8QmYuQemwXC0tghQhBX60TXKa96SCImEQ5wPkylVXYpJjhgwLJ3CpzKyyiC
eTKUj7rIBzCOjX5Kk0uFVDlDuZ1BpdZVjWabyoEL8mPtfHQaaEvvJmm+hXtQUb2yTDhFjAdbNJMT
YVKH68EYZRatPnwZF06xpq4NjWj5n1ghstEItqut1JXh/jH3h0HPSvImCDq4YZPt/+vIjXbccJPY
kqyxKP6bkJow3KxKcaSCWTMaOhMeQBo2QcquL9HDIMimBifL1OmYThNIHTSrYVboS6ysY+X3kGq+
PeP3AS3TzmrrGC+NAzfXCz47VHrEhDsnJ2NIgcrGcCkEqCBQH6Opq5WaiE+P5DuXSvocAwoZprsY
DvxXVqm2vsCt+n+2eZk8iruyzvedlP/rUPPHbO7SLPG0nYgczM81YizRZafQHlkcS19FwVexN3G2
ZeeVNndH9p9v5JQMcihrlAm9EPcSrTnIn/iOOjgRcK4ajII5/rh4QtrLdz+BjGOKMUMpJlTA7Z7s
tKxCpAx1FHfKVtwM0aeHKa13KqOtHuviVW3nJ7fJPiA3A3apQvrfVzDLPIlNFSIh/GtNhKlrbHpr
bC6LNw0NqIIEayS2YLxL3rJ6L/+NaFTXMgvdja1ALcfpUmUlJx9aimzJueZshwzlfEYGwFNACaHu
1cL6DtlsUObRZ9RuaU5Z+9eNkVSbkJjubHz0p/U62VFZ7lSuLmTWl7KMEiasqpEkwHeNCbZKJQBz
rIHDFQKN47U8ruHrLU8ADNxESCDffyBZNedWsXu5qSwC8CLYV6JCrUuf1gbTRIK3vC1YC1/3Z/80
884f0KaeFilAq9ONlXwHJlvDoV8X0C+jy4v0VhTcNaZmjim4YjHDP+BO12/KcwMXsoaJ+DMWaWVs
0rhARxkO2Dal9bw+jV1pusrdI12NRH4ULEgFcdL1sg7HfUwecZESxM4uSDMqDheEZUpD85jBm3ka
oXQ6gZmaNsztvzxzPpwhrQvYtKMOce1Gq84bLtMyrG2v0vKY5xkZepQ3LBqwc1SEKBJ+/pR/Trku
86iWGEJXoBBIHJSqX8YdhVOv5iQg+J0bvNiK4ht4jdmDGBgzmI7hj4OjqsrRFpvbs7FMCZar+TXk
6GWg49QXcmIrs5HpntAnmxMki37+NP8bZig3EErCEM+C2+bfUxHXjitskDnwTNKD7OdlB5fshG+U
60cvuUx9VHu6/ec92WUsl8Tg6ZJuccE2j1iTP0q/I1v1lZRfG/oCOjMzAkUa0ub9A0q71LNjueIa
bV4rcdDzv2OFJSmCXRpsujDJXur6jL9OhfEdpyOHipS8uytHUT4Nci1rK7b6Vqof0w9Wlf1EGBKV
ACf1HSu8J5tp6FPf1aBkVwwaMFDy+U1Q2Ep3eMsgohnPC6f3VtZ7Sz20X6j3SYy5QrWzcsmPWKLU
a5SIWP8F0Mj34+JIH11whPhvVbyjExchspYGl7HR1j6HpD0KjCZ3RE2thvNXxBIJIDS3ntIaJPia
Z3fYj0o+hr2iBjt/TxRk9WINNLsDiXcYzYuHctIojH4nJh1kPbh2xxeACyZQVo0mqX4kSdqvPCZI
Xz6ncvY6CF0t/x2xWQEbe2NNoFQSjtlzQFdZChPiOgmfr47UdYcgaXIw7CaKa9PaxBF0IkHuwQy4
b09ya0cOspS0Y26hZhgZgSYeSAt21whrieHn5e5TUj3AIK4vBlbGThyqnR8uXGueE7fIRaufilZ6
Y7WBAjZ7QmRADEZlDO0+L4pDrhIQzokdISTel5b84bmimY+bFzS+hwnxt2jzfuVaQcjWOYmbPz6m
sZygRHjvQT19uOSflxaXaEGSeHmy7yWaEclTm+1gw0Hddg7gJt4Z/2ZO0VUt7JiPkVr9M6uo4nji
md9FkPI236xUD/mYjrOLaSjqaevKLaJQk25trmu7GiuGo2yLskfloLY3OUcGYJrNoVFRwrq3YJVb
IJuXRjdliaUPSMCFgi1wNNzyjgSC8Z6KjasUOryzkEUeFcewoSVzFBQhrsdaIIPDQVHxcHUx344X
iGzxzfFfGfgwYOCkEaEkilpuefZz2D3oXaTflPw8ent5o+Bo773JLxomgcJtwqvoVXKfULHgPszj
6oHKw1dTkG6/ZnuEs1EeiJTNNHmbiWyGVZkQHhnzcDHl8mdOosqOs4DvXIuTwVAoPDSJ5+jOLoEd
Mck6s+fO2Z1wYpq52X+sWMaP+a+hB0s2cR733fuKXmR+p5PrmtcIuoAcQHTkUYGJEvt5tVFr8vc/
Tb2mLpbotINO2voAM+0PGEXIq8xDvI9Hl2K/App8jeebyQimebA94YkywOY4zO5tZQWe8YbPuP/4
7iLZptbW7O6CufVA+7QNNnbyUzI3+nFdeJioTeS8HVr1CD+sWy2rqXqS78TGDHhvLq033bCnXx3n
lqeHJqGvlboTcvzVsoRw8L541NgRnbWBWI51LnBwTYdwsVM2pxjttT5BpKUXWLiA5DIbiLRWGy7r
zVd7EOxw0/MRnEMMeG56ZF0Mbdz6aQsoJBcgwxlWz4BpnXAyolaQbKEEuh4hVL/iQePh6IYbwIIx
b3jjRChQgcg9t+fem9umqj5DQ7H5BVVqP4gKFQ+dDCzxCI0jFLIdSoMpAADdKVcgLQ0L4curolg4
bG77QpStgVKcMV8Jf/mlnTP+8WrIhIPO9EsGJYkF5BJ/7NfQFm9/9Gm0gQTxIJeb8PzYs4YLCJD2
FdGL3u04RipB0QBEcJx/dZ8DiLXsPfgp0WXiXMDJKTw7lYuruMzOyHZdZt71peqdEOO/bej/AnNz
BK9GEdMsf67v5V/vvI1b5B7vDF1l2KjcbZ/hWtZvCjMYgl799BQ6pdzFraXcNR+mVnq5WGpGv0Ps
oge9Ahq80f5Surz6sTjD3i0yP/hW3uLuuzIIMinMUPulF+8BnMUZN2kq9nu6Nini1lO2wWJzld1E
MmsPYIKA1vE/3lpEaEamaTRtSHp3UAQ9/xOu5GkZYvfLqb/0IUJ7QzV7esdnjG/cUV98hs0CYvlV
Yg8L7i7/61U7uImv/EvCwKJHyZBxMmyuQih/ML1V7yaa8BJA6NtZzYpYOFX0AcdXyNb5MGwqNt+3
rJMCmAxV+Ukljji5G9xQ30vCX/941teqRN8ID9G2LvUSKMMpFrgJIpdxL8GEQwhwEx1cqgqcWeVO
+LvuQ0DdtVtecOw3zgECoHaOmpjBs8TnbBhKZZK3TrOg242mRWVlr3oJ5FcaWzSHuL8fCLaKNBSb
POL7/P51h6MV6znJCAPQtGemJ1RAhH4fhfmJ6cuzcPheTgsgXCEMUbJ93vTQt01m3Svj51/OQfn6
mwRkxOop9XW/ok90RwpjKcaZWjmZ7IZJYySfxVYU9h3vidnOPZZbnZ1QQQ5CHKl2C1Awv4MNB8CX
MfhTxkE7c2ifnuI20fylMDEYX4NrvaISi56aF9sQ5FR/n4aKyi5oxvqTNCsY4VK2TfZLv5VpyWnk
3wCeo+SgZahnelVrzb+Z4QNW7x5lgHvZ1MByxm0oWkpeqPGUYOQ3fwyhmZBXRPgXifLQHkzvUjIL
RikEx2GzXXw2kIeepRAEI1x6Rwqsx6dzfQkV2G4gWPuV5ar7eTm6voyLLt+X1ixMp8bhZOdWF5X8
OOw9G59MXTNgxy0/OnU3CzBii/6tzXwuDlKA8x9NVX6P0hlarGjGauR+k6PScaYY/K7FHhPVSX3p
jcS8cnejT98ReTMDiuWM3MBMrKc6gE9K21VN3tX+lQGoI799EbHEveouFVizlPKPObb0NMG3JBBi
vonI1wfvzWWxAZSpIcWBven4xZPtsRSvPZTmXnueMMvKUDoE7OW11xEooJelPKv2PE66U2rsrHod
mFMTZ/a/h097xmyF13+zt6KBWH3gyQ/9AK/XBs36qQKoB3UgSV1fluuoOose7JNs3DvlMcCOQp9W
jIoiVJn2BS5MyFjNnN0pbUhKfSone5uPL0gI/WWuO3ZzDD8SFum/GcrNIJfVWYSfofzw+KGkbsP+
iUa6nE89PDr6z9SUZu7WD7HHWhI5Osg4GSOB4x1IqU+RTHqka9VH3ob9LCmYyDMNN2ZbOgW0oCyG
q6Iqjk8bIWeIL/T08r8GiQWhFccfsIhUcgPKe3YCD5GkvVeDlzYkXtMGnUK0FpCVW7bb81ljkW31
enKLMaQTLXiXRpV6Fk8sA3FXyRv/DYO4kgVSNEgnd2D+RldEsK92E0yI7sYqpNrxUpR8RH1YyGYt
B/0IpndTkm6xQdpv/bIbv4t13GJ7E1jQhk6n6WPhXnO1QY2fWj4cFf9BaiSxA+3AUA/9mcHXktFc
tQ2wdO6jcrIa7LvNtWSI1A2tAGL90MzeVTj/gYJ9igrlCoY7xDmFFvkeF3FHQiTI3iyWnT6obHa3
+J90qyKa+YdonVDBVX3A0C5aH8uQ8neB+31UfF9V5FXypVVyRHMwXSpnRGU8/CoBNrxfxGJME/Yn
TNXuPpq8KW5uBrjiZTANMAAQOa4DIfGMcwtciNWAgwzclMdtHsOyW1LY3VcsDeAIrbkdssFRWjpJ
wT/DSca3/2YeXrT4JFI9Fy2txOicq6cWtgDxbyPZLg0zb0wfQY3pQgfnRLuhcHBvhLYYWSY55o+Y
BrTbo0Gm23HXlVlh2p6bjVPY48uslF2IsGAJ+gZF4pavqxaS3cQqkjxN+4fkEW7lTeuf0B2whFke
q/+6++GXH5n61ILLkS+vql/SvErkh2FzV0+qzK/IRgHp7nBdx3FvVtJKXpdMvUjbmk1EhsPqJvz8
lH8UF7gHjWzeyvzWH1YeGCO39o7aGRlmzOJsy/PF3zggfAhls2D8dGIIb+qhyX6nzpGUiKPM4u9L
SI3skoZ2Zo8qGvss2Wt+zb/K0ZrBToAEcF7p952KZvJ/HPAil3GPcRrlNFM5zjEuR63TxSWi+kER
yplxLMz+tgUjHaxG769a6gX1wrez2yXYBh3b2O3ugFyIjVn8HMFDYQfks7PYLTHHVV82z1zR9OAV
Q4oH7GvWusO8DNgG1QyPRufuF60nSxwrDlyTTcL/rJ9eAxkYykGJCmjmqE8FQjtiroH00aO5Blfd
JXKYt+FR2OdK4fQ5e3zjAdGOVd5y/lmyXvn6hDAaviiwB0h6tbs4gdnlkEkcK5+LsnjeMdrVK42w
bPs3MNEdq32nMsxAhKswMwmJoEKlxtWbgP+14jftFqaKKKGxyKP4z3MJGJo4JQVhinXpg7+cQB3s
XnBe8vUNly3vJCkYBpEIvjWKneaitlbdMv6Khv3L2T9+7kq8VK2l3bufkb6AF52BxGHIIphEkhkZ
Ke0XhHbU9iTMLsstUxY2ZRmLz7UpvI6HJLBgOFWjVKI4V7/L2W5y0aBbnjeCcpTNPOPFOrAHJWVn
4V5CcKJ3sjm65FMklj70YF/EqqnFhOTJZotcsKXLN7JMjSdzWDabnJ3z+IHOPvlb02Silx6Vzwr5
HBljSoMR9pJP4pRpEKjbmAi1eAhwlQsC2fMRu/+BiKqyFl8Bor372v0dGutGq6Fvy0dHOeGArqvR
hgtV1HSAB48tFYsjH4BYL/NPQUbAJHmsS6ZDU0CSbd5YK1hWHd1B+akVNv6GasUuGh0xB3DyAzI7
Dy36N6eBVpXaI1VA8kLu4fuRP1exYOj/oiP+DmWB2cyxL0386RQLqXYB7yKGA1LRzaYpTFwmn+AA
6lA19L+SHGyuXpgx0EzZzDIM+Sj5+fAUY5pjox13VtGf+L+Th4cx4ygpvR1l0vGVYN6hgxLsiSy7
7cTDCG9Rsw/DYhVtr0/VcZeai0jsCuk9Am1B5rfwf23klTuD6FLlLYiACvDNNfAO9DkAoLg1bwzY
gqkVsdLl8JCIsiM+e9YBQE0becMg1gCqVqxw1vwU6cyA2LdA8iSD9lLID9qOgvMB3vfXQvRc6tmW
VzyRYdiqWGUC9OLpAKYFHGxUGhl52sAB7GyUIlauevTHV+ARBck065fsOA7eqarmH93P/5pMCBCk
37PczWLToGiNF1mlKvUTadMCslysa7zlk/CrbSXgT+rt5HEUrwlxSFiffu1eGQjyuv8YnwEtX9ow
Y06l12Wd3iyYaNy2ZrFmu26uAtXvedKUy9xXuG00BLqUB3m2FyNt691rUSAiWUssXokEMKft1aUy
6jaPaJgLZWYaqMbb9cuncHPDfJt4CgfhPQqY70nr1kORV+p60M+GCiWZqSn4WdEp17eZHSUXKs7P
6gZHOu+YqfD1gKtAhzC44MkjPc4NJuCJqARs6OB79l7+xGYBERpfexXO4UtSUcsXrRhdXnrXxE38
I8Avk16A/ucAlzDV9Cofjvlh7OIsuOL74GlhIiGzzCl+1ohteZJ7P4hZpG9IoBj84+ziR5d+F1CU
lKi1RWEoNzxy6BTQGFcf4aDZhMa7Wr5UaBM1ASl8i8begPn4oKmKvK5hgiq+OnGi1PMu4AcAPr2c
HJ6bQ9U6iU8BwsxvEV91F474IwTi/vnamPmgNZvx+brGj1gQVk/TOjq0nr+AnyvNG5LPs9f8vyif
A1HT3Z09Usp8+hcWUEdQCTMVs2e1MR0ZyDE2Mfu90rFEFMFQnScVdMWH5Xt/t/pROdUmS1vycKMO
GTkz6C94ZL2q1WJDOqpxmJ3cdAro3T1v34dHy8b/E5PYQCt92dfcTVEC1Av31xrCs079wmDvi89w
7vjfnKHriDHuvBL+qrXoewuYDrrGUb/cr0bytBcoPr+twkEnLenfHuuOYvFToF38C/fwFGvOOG/e
iic20kgi4uGFp7y2gK0cf5m6Sx93o/Gulda5YVsH7l5dE5OcwM2hMBinc7t/7PAGsgOkp1+YEQ2Q
b2o3qGuPBUF7wB/496gH9VJxn8+PUphH2B2s4LGxtbS7auxe1V5CpPUN3dWlZoghfOwJiGKObsf+
BzpF2MYMUexhhBBw7sPvaZ0DmmLIwbqZHonDGMh0pi3a2F7ivqmA2hjOeEDT6FYr2v53/Ffi2HA5
GPMbTjqG4urpTJPjcTu/IqP99utXjY0/bDlnSokAGNNLIlLZACEnfmLml0MWc2Guyq6PgKwxQx4i
a7MDuDr0nsDOshzy7nWxVCf/QxcPkxrwzEWicWFZdTdB+aDpjQCAqzGVdpwfHVQXWD51WmOYgALD
JuFZ+AxxYysszryBqOPUDGd6GUINstRYqlArR4q09/1QVgY6NdQZgcS31l+646eaj5KHt7JSFF4u
VdKZJRm7ttN4tC9MXjxOzxWEzueqxe3ytYGpwYNazLVND2sBI7zTcYDJKWAtPeX1S2fAfc9uVYkA
In2PKHyqK62liIu8rKxr0KFZtPTUaXsGElWbA2Ce0Faeeo/JtwK3S/6lkOdIS7OPM/TSfBLkgxtn
RhoaOxHVkai58A86e1r0/0r+cAHqQ+ic/oB2b0uLK3K9L8bHir+ANnFt0DyvXxtf64kInO/CowtZ
oZCuhkvFizfYUZJqmfNwslZVo2w2f2P5qFHg9ssqHhGT1mvSjLjF9liLqqQx1WEXjIfiYQB7JrYE
b+ZriQk72IpOPfGMftk5hVXzkeH48mj6+UIhYxY9TLxWtssMxCfsLXCMs9ksCnFUFtBy9tsyx/Za
W5ZNO2FqH6+BWGtEHlWZH2U9NnJAfGraYKMenWJTvSs8T1yFchuRQar+IeYFTi9fhhHY2m3sxPtx
j4hi0O24uVLTxRX89teI7VGmFg1R3qz2wDLQmXDpzFeidp84yIQL52gYyTSxsHB4/RsuE67yGavA
mJxQwZsjpzJMcxB0EZlGTQuOMMtyfcLBUEP0+PwT7lOAcFJw0w2seYrBGqeT2aT8GXmGA5JOBJ+6
xDeBb8/q+oFssOjGVl7bt+xlTYPD/zJOUHMA7f0zNFxsAAVUbYkbhpQWJcQpEnfe02F2GfbVew7b
da9gyXaBO6jJs46KnHNHLQXmZBt3uceK7wnEy8218pX107WceLgPw2e/PcRSezrnoGMfpgjzNkom
lY6waF/p0UPEauFbrvAIfkO4hRMjCFFv8TtAEAc32ULziHT74cOt58EHQlMC+QAGuencdne1wZPP
6OEZT1enOolNxhX3/TZ1BoOZZclsU+bulnNOgj89kGWB6nUv5LpmdfjMd3b2UAdhS6tmWB0YFKy6
d/Z5Mk44SDdMIr080F2tw2Y2VuXLUi1u71vKchx+VgViKi9U3aO29We4ChqYMu2XzXA6/h12hOBY
Hl+lwi26whHo1lZVrD8nYgDWrGDzDnpVCWDpgeaP/1xhJKzurbln7AC3sl/fkvI7z2GcBWknCakw
5uwsY2JpKTtX+k8Q/t7yNjzRYOyJCqf+16KhlDTtt/N4PiVnvGF2m4z4cU35VLp2VdyxvGHhAhkJ
sMJePoSfdoShBRkU4pn63CxIKyYuuLodvS2CX/65J0/zi9FCtjhi5MuCnq3BV6wlcPOMr18QvLHu
OUtOvLA/TpzcS1hquT+DixWYARvPRKqd9hpi2YSDhFRgImbqfZ37RmLX1Fl4u6excddbh0QFARY3
iw/i7bAdOj22hhY0azoM+wjpHJkpHnO7Yq83dWhawfBTY9Xga/IkODkRDRje8owyDnqfGUk8dJUS
fGNXGdudcPWC773CaPjpxQ5vyHGsRiJtn8TL4hKh4UTZ3D30japXtExwCLAHTZbkEcajTKe8z9R/
lE82PjmCOUXBDlhRp75e55KebIvX6uhzNk13rZZ3+cYXiEm8ydwFN4g9IQuFC4pUbRQWtI6jsis3
l5b8HegeX5K3KfhgPK97tAuBS/ZWV9ikIpuAJG3ZLFMSBvcoUnjOrHtvYxq8qKhEa0CXnZiGxHDf
tuO7Sptf8Lod8+FEmVRH1xwLfZfwV3ST7USuF7Yy+mVoyXcq3hAWP1a0mfl1q0Rc+tKgs++7fNuT
NTAWmRySx1o/BcsO7A3HEL5OTfttV0Lce7VZkTurvcOxBqXQMGGs3FgRo8TeV+q5E8n96TmoCBL4
t/2dYnAOO+xUsEiZe02VY5vzASQYSHeO2vWEcCqykHFpFbbZWhc0uig0l0Mo+1IacO9GNwhOHtkx
8Ogys7NRrypdDb8PcgdMLs7OdSockUB6m1FBerQW6KnsHVrpL4oyT0C3gHcGOLgAG9xgf9McGRx7
7/k5sv+YbqJg9K933etAoVcpARz+HGC52s40Um7bmICXQ5QLrzvAmWudRkE8an3lfxfwEJF9cAZc
M09CntUBEtNS079WdqjAUhZQjf1O20KQUj2JxbPH5QrUu+r+KFS+Kd/CBOdZ5Sog4OK75ufRXvif
LwFUd+sQaQhLFKcDxJLCqS86y4pIflC+XD1/MW5G3qhdkakFe9mE6RnCK6XFuyEA5kJeXa+Q217F
8ovAYnyKjmomdR3hYE2MZ5K+gqdmuIJZlf1ka+MAStAPX0hOSTMoA8qzz+85cd0FazrRWP/B2R/7
3pJhwLHxo3AKVlXR0NF/G9M6g0rSlAtEnHx5jD2SDz6bIwdNygWtjQ24Ly68OVGjh78Rtyh1dnfv
2Iv5HEMPOqSgHujnx1o8+m0McNsuhesdkzf9fMypCUG88ekkNeXpCcOuYws522pP1i86oHWeiSBD
Tf77mVjq7Lue2WUKo23zBFainlSHTPKIJhOm51mEcc/yqVTIqW8TaZLfdziufCjsyQxim9fVYLOZ
H857L+VPIjtllElsZL4GE4aAyG3PH7mZeISoII36kEmUlEvoYKgygcuWMkpGBCi0gTFc5jRCoN83
Y7zew7JkGXggu1mlAtjgQiLs9yXgnimrp/uNby91yWPGaznjZt3SboIV0RmPIayVqO/TITnKCClk
blU3LiaoreuV3HDvVyK3cf2ruWgT1qjD6tLPjB/IiHrdMmitxJxVbNb5fW7j9OdaWxPTBbsOdivo
FPaGydzU8c5+Mx62qfl+t61goOs+9hdjY5U/exXbUsm14OxM/rw0I9KAW3N5VOHxvaWYxJ29PtG9
dhelt17yoLVIXsbZtLE2ciou6xOui7Nx248OOwPwBnmO/QL3rDZ50BwtcZp/azqrw51ZS823Sj+6
faKoCNfliixlKrfUx+0ANPX9RUhejiIoPSxHJp683PnikqgAkixDNFU3v72RhPHDvYEB5Ibr/BhK
KaRauuXs1u6tW07358WS2TW2fI8w5wBHOpTMtCsyX8N9TB/eu6Undqk1s+r7wG25KioBaSVQ61jS
11n9aEox9PbGI+xWjiR5dKl3X+fDjGm8DhVU72Z0lXHSJMEBAy9xGQ/K12IukZZXvkPywbBqIT/9
2pVvHtD23sA6awGC2mMBDgRdTp9a0/Di9H2OngO+3zjj1R2Gd2fN2W784aOZ2ger+YgB++gq4rlx
nfwrSkoJRlS5uPnYRmdEwlw8mRolgVOgOKc1UPYZhwwj2Ihubipre8/CqHwRGex1X3ZZ4baIUznh
BeD5NYc5g0ZMdY7Y2tWz7ueHZds5iNoRNSvyl/vHl3Hz8YcpbBlbOSNVawViwu9fJCIo1Ketbwhs
u5BiMIsOqTGay3XFFqHc5LeCkYPUPZXNwTRGnAPNcUVwzJZ5iZAIeJhfM6qKgohCaQOTSwGI5EIV
zoCq5OVu5C5jPj3Z3p21rypAZmebWG+MxkXAz+T70zVoVMNFLKwcYESC37IJd7IF5pWXINdhER6t
54yDwjjJJhUVL28Kr05DngPQ+SWXWCBO7Etfq3r4dtvwZdllGi1GnQTDMv95SBSaeC45nprXPFGx
5W3TGLnfVxjkiTFhO/2Myf7dLl92u3FgS8ebIa6HijBkCYTKscGazCiC8YHnu5+wqmif2H7FFA5g
O7m0H8NuStXITEFn0+pJx+p9QQ8Xb6v8URaakJdDKWb/JPwN4PR91U7xcOa/sTGHgbfLMBORmbNd
WatVDyCI4g8IZ646R9IsU0qdKva3xzOV0R++dVlzasbrBYMOaI9Ga5inl+sj+Jgec99IxJ+afoAB
utIGuRYfJ+xJLJPQ4cfNc40+bUTl6M/bQrmK6a6nPGU4eQvesK9LI5/WSs6anKeIZBgfHYpDmPRa
45sQM3voU0UqgIVi1d2WrJT9itjkmbtKFISFoVsR/H8ebRJ12K6MNKZzO4b9e5tOalaoa7tyx985
bLedsPq8V2uXDgNoJTJZ+wn1mI7aXF0H+Jq5i9gk0WuoMWizjPhq+iOeLGNp8u74cydcf2lXCSdZ
hVM+WAd5GTexZTyhs0zAxSfKN32Lfd5bXGlnD7G4tJ2bSYKt0ofjuMCyU7Bwe/wSyoyuVAXydWt0
Q/iD3z6jNNBi2vej7Fx5P2FMmjg/WKixZ5LKCRlDC31VTw4IXOqNfPFqIT10r4M8lMFlcpKwhzsF
mCbY0hwXrL0vlMvOq2winQrYP9efFk71gCziCarmtAWv6MXEyBVoW/cMxOLVzu3h0LTOUkWhTSF2
32lutpMAyUdEsAwoSsdL+uwcbrF9BTa5oKiDulhu3YHYIFo646p7M0H03eqcL4dY5PHexI092llY
jklJ3qxdWP0hW0dqYr8dTZz3CtKZSnutsseY683YGfR0r6aw2MqiinsAqXJIs/EXpGM2hDIj2LlQ
E3S4izJIAWJzNcJpe5PHdWacisEsWnlQozy+W3UFoWS2Y6bq1IT3Nwhx8Crac92HhWmsbL3AZ1IN
LBBZ1ar6fKpCa5JXMGfO3qCgx9g77o2p3MtRQAO/kSROI9DVvG8ebX2b6a+9AsGaObfmnabAvTwl
yZYL0wcySJdXwlzPC0PrgKkC+py4+tYzEm0tIPNdZyZ/wwHgMhHMfwNRvv3pZG3o/JVe5HBpPjGI
YtfwAoH9CV3dd25pnr5dkVYEy3MqrmbIMoQyUR5e37A/bEGCW7d0IoezXAKqv1omgTLAZI4H40eE
sIpHCa1kyg4tn1KCII2LE1G2pIuP9uoSzl3FdZc+kLMVI0urUewqe8UsUSjrMTSCqY8HVqy3xi/T
D7IWqRvh4kDODoqymiIwjNeVvDyLi+28mCJ/gS9KfbcY/GJx1WKfwY7Y/lwn1YCGP0hsg9d8Q5av
thI1ZZ40fbLwqEJgEzZYICy0f9qQb1Fvb6NwqywucsHdAlCA054vwg0mYwKoS3IbvlysA19srhD9
X3QuKHQJADqvVpxirUlpX1oZoDpPLQBtJLqyHUzzlshtFRJzQbRicQjv7FxJOln7U0LIb2KXny3i
S+n6al1RGgC+cydzANJweFQP0/need99AHeY3jxS9rl8LP9q6GqT7ksO7lXejY5xFGtblGTB5Qgn
dVRgnmnnVmsK6Xcw/NQbOfArWW5UVGfXPg1DspPoiFf8Wvov+Oj+/KDmZ2ZXNROxmK2UFY9UdLEk
YeyYRnz23fAS7WURBCmtvTaDyQuiVi0G9ba6jHSXnn00N3nASvUJy94mUIeEIEpuqpO9+nO1n1WW
r65AgY/BMFqYKA/OdCZgEzWGZmN45dMrmtUE6FWVzGsdvI3JLYtVqcxbKPaRcai5sNzMWpMWAR9+
gr5zV+0Xbw4bejQz1uoiNti4IIrGx8LS0CUH1MeKPC3txVZYBnbEfu4J1VMkRzn5RO1TeVF28Xa+
rL8xhIVJH/YOgdvTf2uN8gAI8kXdXjrKTbhC69o2xKPwg/lzw5TPRGQ4kIOE9Pyti0QR3TmawjeG
xzMmyiP1B7vL6ip55s1JLh9XSKFplW0hz5XWgGC3ST4IEeRMDy9Uk6FYY7noTpdIA4RAo2OzOAlg
XpWHUmeVZZRJ8o5b9P9N/hzPhk1n/MWNvLx2oIPF7teson1a4aepy6jMVLCQEwWchoBT6H71epwJ
ovZvlsmHgRHr8set6rULp3w2MfKADWOTEreZ/uD0z1PIdYrV0SfJ105bLRYipKYugMbXcSR7uzD0
CPKKNN/amWrHdI4f2C++r//fcLdbpS11wp8+wQfkWUZxy50XnY0tUGbLEo179slGYWlcSnfJBIF+
TeQcr9uGMwTgwK6KcYpiOI3ZdiATzuHp8FJDQCAdzrVr9192Um30BH9RL+vGzVm89ajWDc84xDca
kfZKRp4I0LuGOiVva/GTL5OPBcp0VHbcDwBUeu1oBlTZu3g1Vu4W3xy4Gwd+XCdqCkyLppDxbGgu
b5RvcRLnRAcKmO11RfY9VFXrQi/AeZ6Wes4stEszns8tc53TwjmAIQcBJEZv8xbOyCbw1Em9mBsV
/MbOTzxFu7S0QDvv1yOH+gKy6VDTWAqRIyurBIRXf+oOc7Vm5OfDTHCgC46u76ND3zA7WZjcJdO+
2i2vxlp3jo7Z5mA6MHbACeTQKNM563vQ34B3yxkpyKmNhwkYcSlYva+nuXrAfHX6VfVVnMnYpBiT
8y77W04A+hN+WSp9BIcUwecY3GujuXx+eBRWwl8XQ8cRlyp1wq9moKulnFqHWIxL+r7692VY8SrS
NtW2FuZd1kCBw4nzRlvrKDLak+hfFaetN+CXjre6TpO+rhgDbb1x5iCki0m+xSoQDiH4b5hQDgdi
JDeCS/xZUUIuHiQZsKUxQxLPUEBGJiuWQ7ib028kgI3euqAdyDDfuxJDuzW63dB/xHx8uyGHPpkD
HnQ7NBtBiNZHo7GgZ00xCp7hEnObpNHG+DzgwTn22eqQu92xgpSXONr4squ02BZ1aip3a/54bA9M
ED4SsXdBGM57V3ZSBtvuRY2KWuUSeDDE3hKA8gAQzzYYqCfe4+uQmQUzLFy/kiu2fVlnFemL8DsS
/x3UtTFkoz8sDdL1do6fs2yWqUbF8r95FgmNRvAIBEha/iT7v8RJTy1Q2z4UHHzdQCrvz9OI00O7
7Q7PeuqQyJVOC5tDePsrcQkrpfnGSi8Mu9IUlTLqh3O1TojRn+P4FZrYJ9fkNtMxXx3njlzpPfKc
Ig/881sR8M5yx7jNtL4MFotXLWSrf+6uZd4oPWHO5jmziIjuO7mPDDSpNeB6sqLtzII+r4+5DWe0
XLlyyVKynDcjoRHm6jG++amUFPX4AUb3uAEN+oQXgLfgmHCKYB4BaCDGyFrzGO3WH73shC9PmL9k
nvaIzWi9kTgdmHo5tMbelZ1FeLIhOXC3tus4oo8szmC+hCnJA7ebNpLHiVdrZp6bvYSvd/NJ1Wh9
K1p4s5jJksSdDMswPPjI1ilc3oU7YM/StVS0cIzRiwGbHBLYT1h/TOt0wlm3201Cbdytk50ybrPX
W8bU/NDeImoHGMSHdEL5O5JEpgjh3d4reU/mUKdh55ZeamVoJ2Y+q/Fkcs19arGg/TTQ2xFleILp
CLyQEpLiHcz8DAB14eSUkXd1BQcLFKq0KISWDCH7H3CVhcPLRDB7etVzmZCso3Tc199hHWspJ4MH
w5b2w71IwIPV8jWwpj53EOnnyNi2M6UhPmTiZ+K76NpEQ13LIbzukqq79rVeqf5bNfvpP9+CBtRW
SyeQ+GZ0/yWIfqsYyOVI5yxEgb9vV8FpfaIbJ8lZ7DeZukXhpb42tMO+sTjz2skzg6w7D0aWQxck
HflrkRlBqM6YhrkpYz0pQl+Y9ebxy9w0TcpmJY9iDFMKwWKnBazR4FRH4EiTheSwwl1V+EBNTv5P
BHTgTP4HoZP/4rVbQOjr82jTYHx06gj+BCUKO9so88fc9WF8zOIWubhavj7mIiATWWZl9+NZ8foZ
uQNQCATXej6YpKqJNRkwDElzub9NNQ2nl1NCiB5LAEmLTx6ibTRZKiDB8gv2a7A53CAHfkduTlmn
TkRB7DJCE5I1DwVsDspPuZe+t5hmf7ozFSRA6ouUIt8754AZHeRwAKjxjznsUI3/iS5DxNrAQXv0
p0fQbWiKTgLPFDrc4FEhb5UKqg0tWYcs+6i0Ftosvwor52MAWdgpy3sknN17wHfJym3QM+Q2kmwA
tG5CX+moEO1PWWXr8ZCl5q1nJcEbINOhzAkxVaj/lngC1oW6i2WIjtSEQymZmGVykHqTLWuVK7qr
kRgMUS3Z2ZyBlUra+fiz0m7Hkbm+0Z1Wjy53FwIfwTxH2OYG41ywA0SaHFsxEkxOyH22ivJZEFmA
2qnGlHPORfr7lDD6KBhgJ6fXHqzvsVF6VTZFZjPpiuVyEaaP4IdNU/4kuJL9sZF3q/9Lk7nKyTDQ
Lik9w2poB/uYoIhknGg+mT6ltvjQRCwBUqAwoThZljMZI3Fw7sd597AZaf6/A+Uqsex0JpfZfxO5
sW639gM07q8gPo7wckvJHZt0LIIA47YB69Qx03p5xDhbXwuQWiaG3OX+E6duLQZ3swzJJuHmmYIU
a/5JYU4eOCoIO7X1dYCpNN7W5eho6h1nKoCO/a9S/W8qRVpf4+qrJdVrtGOkFYOSFrISDnkhV01s
+VLg0Jf4D45cFRNiJG3a4j/e0TeedZItHwIVQ7a6JtOpP9VK8xZGY+AUv78loolnPeyGyR+UZN3h
zrd8JROtxCOaXdfPD4uEC+UtyaegTwkbZzxx5VwIUPNsrtehL+agZY2kH3g4fpU2m3HOlPAh5u3v
j4rdf1+z0JKyH1/zqyQs9eWDpRabcuiGbW2prKBmUKFhaOeZrzsKmF8fNEk16hAPVOQXjU4y9tMz
tivbfbS/DDUet23fZHXTTx6XYzsJ+1DjjGMQJcY05xH318tShl9q+Kuqw0e61P6ah5IDpOsYg6Mv
GxEPBaHqm1NaZ9xOn4rocSMORjdSGDRP156qYVY97W1vl/RAE2FkIoIqbzzwVfB2EFv/K9Mb5R7M
IuefAomUS4ytcLXQirK5OwfyD+IlGCmrSnrAkKIKXK1LJVRHm7MyGDHm7um2h90eQzmiihH7/mt+
uNMT+J8wpt+lYAvL9c3QKNYs7mCH6Wjqo6i52xz7+K9rDS6N9FLp8wXdgkUIGPwu2zmvRGx5ZmUA
66Sj2Ry5j0IaRydFDthut2Oqm86I8rwylov7dPZelIc+uLzlK/gGTYZAPWwkBbHoKDo+6+O4wjc6
J/a9h+2VMxPO6s5naRCeS3SODKoYhMLZWqQicF8e9WujhCcDR/YElHihffQE254SgJ3RS/Jx3+9O
e0qwD9nDHkAnNHPnWT9oFCkJy0oD7Uq1t6vmRXHb3jn9WLpBhS+UhCiuLRTMnYqROXUUk8RUSo1Y
m6WPO6hjwRxQFB+lBXR/bsy7Gr09nVw43vyTrLvxofqH90bhRgXII0IdwSZo1YHHKBBxK2JPSeB6
7DocuoLGvcK54kfW1eWWOQV947oJeb+dY3BKF98s4iLltIIE91VVz3gMD0rng6gReWyRn21eyUrv
v1xd5i13eliD4OmwGaRSTlMcxgvuLwlsi7bFVe8gJ4ytwOS1CF9yNSi9FjfK6THMjKZFiFauxPxv
vCMrV/gxmJh1s/zBHM8Aw4QPUxP/X3dXa5RXupQfQ4BSRa7V4mklDx7UWMYud0524Qm6BfBMBfPY
AJ5IXeL9kV75E77jnrHPMYH3Vv5Wky3olwkhVa02KwLHCXrpBpj2uSJ5x1tPAMXy3AutBrqe4sSJ
TLH+qQtYqqrBPkSWJe1wCMXpr41ZhTWdp9wTuTMVnVHWvKgj+c5fETX9LYLWvZiAy5PBZvp9b15Q
NMhBSqquHkhfiOTj+L/k5EgxrXlQRMb6d3aWdBnJeN6bzkIVYiCOu4uuCtF0R0NQLmTFlibiXfCc
/1E0J9b5SjImiXPDfeswdXVBo1K3J0VFnXm4LIs7o9Qll5ePcLYRpwDAGjpUxsfiQ8Ff/pRaSU6w
FIpq3va+/SVv5KsuFYKeEehT9MrzJ7NPGxXRlpFWg2I7JcgiADCIHG4TH8titTKlui+gqgmxKSQX
LuyThrNNai48E5SPdpu8pDz4PUp89cET7pAuHYUV7fsqFZa2s/IbRvSk12ysTaG5v6pMHQKEAkqf
gjLYjSmAJPPDhOw0d+qoxr/6Nx+DPNZDotltavHgQS6dWbApTXRrHwFYqsjbZGWs+cbG+7jLBWwM
Ab5gRFL354C+4T9H6BXb7bJ9k87csc8vWmVDSuLK3MF3FPCX6Bhk9W7tIJDBB8iF5DMG3SE/CSMx
x1bhK1MXRkNEVldpqNJyMSVJjn5dZAVv571gH93SAZNl/worwTYyStE/RIcEufvxvKzDU4BAFw00
FejeFYyny6iBvlNYKg502VoT4qG5c+ThnxxpCZiHomDCr0EEol9q2nwlKqxEbWaRrxR83FoeOcGZ
truwIGFyGznTPGLnI4tVHMzHBlTXMN+YCXSOvBuuQCG0sMjCPi+sdiy1PoMGbqwtgzlk7weAFhgy
FAcrP8qBq/LseS6X/XMUdf8aoSgIQfveQqsduGdXbqXofdrLkYFCr2OcEhuRRV/zM+YdDOhnk1Lo
y/4Hkb5LK/FWRtF0wGl3GLMxz4chirEJhQp9xTO1g61x0ruu3LtuxElpOItMZq1G9VdmG7p1Q+lj
tbWNIh+Pk7w96+MjkMdcu0Pr6z+FwYM4LvgcYIsfLTloUgsSEdMpKD9RMwt6WPlzAOHStPewhHjS
RxSjFpUrvlC8WqWeXcWH9torg8oBw5kJDz7Af8OxJCMbxeeas3fZHRkCtMBZR8ae/PpiX54mnxHE
3AUNZDlOPTxpT5H+9+hrXvfMH5+sZ+yer5p2LzCx9E2C9CnAbO0pvNndXzJb8aIJg/MkzjV2YgRe
8EBxH0AIjLM4VXmexn5M8hs8Vc4eqx66CTNmsR61WVMzlKkJs68QZARvVAeBAchnW83AK/AEpaIS
Ye76MubhvdX+WqEs9SoyE4sbR+gnDLDaY5FQ+D9O/obRSlfsuqfdaPoNDqKm/9H60MTMI404Pw8b
wktk4C0VMgqBI/jhJfak56aVnGWxAw36G+leUYjj6ErE9lNIAvyMoumm1qFu/JSjUgcUBRbB9qOE
A47+VskmVwaeNr3Ie89sGuJb9xcLsLaIMFCdoDAG7QiZ4d8FQTPvJRQuE0wZhXjkBgpzxfq8MCa9
qhXGaNv9w0mwRQQTM9DG6/V/QhzPSZzCIbZJvr0eVFFsKD240st2i0GAp9VoP6KKCmugcolvqQKy
yH7CqkRug4VCZPUi4RrR6mDQWtpxgvKfaFZVf4H0UPhEN8r4UsHQru+iaXdZetgqyaunulkBQOrL
j5JvSVa6yCv2ghRXnoOiBYqK1jx3vHBoh1XKgxmNy3l/ORWjvv8QJBsZhkVWsswMBR88V9NYWT9V
pCGt9OwC+MJaJ+2VeMbbkR+/SA7pV/N/sJcmGONsrxsdVBCu/pnk+/feCvtE1SxHBcDV8HI7C7GV
BkH8BgrfG1wUS7qHawycjPrwdgyfvZmXokqmOuBctLur9PRuxnVWZ4d0bWOQ6cYdjnN06LipO2uA
OcDB00NsLmyUdePV8Awgb4mV+UnaLPgKqfJ9QWsR3CeEY15FOz40aMNwkUgg/bBbo5Nu4druts+Y
4wLgX1lqHEG0+El4C5MMeE/T25ltJzoob+TWrF8KRTTrjs5EM0wiYzSPy5aN10NlVt56WyMF47EW
VELWZSmIBlFI+ZiAw0L5jkoraLH2fve/Exy1eZVRbmJVlaIlPWnHbkaRfyqHQn8llonH5EgR3BNQ
RRBF69xv9fK9156/rDfQ57R92Uv5mmPa4jBru4mxuprb8M+cCAQjaE9aybi1qGyTOGe9kH4qMc40
S2wkPPrQsp0Vfae3TXG4TC8uuxf9otlNUyfq/hWsbnwUM6beA1eqh83Y5Fr6iq7QRA6REZOY5HS1
qWkQj27ge46sFrbo5GIzlAY1oNZBUhDoWyge5OGii3jiQ7KyminYL/S9Nl+ru2u0CodRgoAf1A9R
UjsK1ohjuzwRuGxI/6S0asFn2ULtsxecv9wlpfqnyk2DS91I2CowhAiQeuv4Z2LPZbvcb3OcmnkM
PcKrAjkYpHIkm4ll8Yy1IeEI+a4lSbckCa+ChUvPo4tHe+7D/uw52/ZJE5zUUsPTSu7UgVCsSKvT
3ox/matFK9IH3FzhJRoHU7DdpCp7tjIWgfoOFO1bW+M22HVfJDjEXzqKXOfIarOqNF7pGJDfMQIK
NOs5Pn1LlVgkND4ASQehhFuStrr+OaRACIhPYVbXo6OrEm+g1syPWr6bPr7kPk5gjxey+tBVf+NK
HOJ012SZ+DrBuuDXYnqz/gO8THcdhGR/JZnqHZjtCw+5LJhTyKObUExZULcLE3oT80g3Flxk5/IM
8QBVFvJWrox1zHxwY7NW1nVqCcwUy4GZRJXQIE0IuVcYlS9YWlZaH4xlSjJmjBCSULnygdvaXmtV
s+t7n5R9kgJ8RDqk/LDaL0hS1dzvWEIxpvV0TK+oNWD7btOCK8VM6C4nv3eHQdIgh5Sj/m68FNI4
uVKKsTHfrgh2gFIffb63WThdz3vLPnRFhgEr5WBQdn2do3bXfVjjEY6aMnAwBeprbspYXRC9dcYE
NxSFJlek6xV+0yhrn26182GtpxizIyHFdXlVc5+0wZSiWp3/ZBLbwgt0hb5lJIGCVQBRjYD3VPho
2XJdAs1zGZlr+zVvIr5foeBIDkVmgK6307WA6pCHWmRt0pwD5TbXpwgONIEpppa1Hg766xxwwqIz
eTAWyZb0PjDZLzpErTKyFN3HHLZFHk1IulW6mbFz4QEfX8Y04M+1gvemdGMDtArj4CydjKv/vviN
tmFFthBNqV7eKEPfJI44rNhXfK9HoGnLT5w1KhzIw2xPEsuuiKxUfuRO8eeXVJ4d+35F/MeNEj5W
Vg2Nztt9eL52FsE9JEgXAwxowsMp398j9Ws16EFocYZd6yvKu9E3xRnFl1j+JEJnd8zp2x6+J0aI
s+I6wCvvhmkVz0KBqPxnyk7YlLMiaG30MirARUc0w9s4h5sUHRVwo35BeCzzwfschRxHDMWFzEJG
N65fHadXVh/ayeJuuwa59HExMmtTOA4voE9+WOquiaO3PEtmW8X7tNAdmWCZpIJdrdcmb1lO0flH
itTIzK4g5gjYF5+dYnOX3amz4I/xwH5clhrSO1r0LHA0taJFMydHVhF1f2U+EIZ7GwdaUHOR4ySe
FBvGjtescdlvoq/NlhpNIe1bG5zTgmCyz4epgfX3d+OIxNgb9LRRjDjlVuM+aluKyffQ48+4jQdq
vqdoya/hUVFEQsjb/IbwLdn8FVKsWIh/rh4pHBdC1X/iR/pEzMAWCHOMq5FiPrCwbt39uglNr5bZ
Gme6u0VLT86V3OD+dIGByNnV2wrgwKa5+H638wtEJ4CSenMKC+622fY5NSPVYXfFQo3TDp+A8y1p
ql4r9GMDCQtG2jJeOWOsGq0Xu64PPkarXZ9fSHHHw5WloSOutyIShErZV6+mgfUKDYu9oC5pq0Jd
nmnynHkri5xi3ewXheafGBnceurEi9Bkfr/ufBbCe63/ijytT+gsc5cIlEfyI8awQDpNHU9F3aWM
YW6f9YxVeptqjTZKAQFoXQasplA0PiZNE5UpXBjC/WBCaEaW7c8/k9rBT+GosylyM+X6f6DVOplj
Ra3Ytz0wFyLwOXdf+xTUYkLOHM76zZKbB4rAwYIu8Kv1o99DgEsuqjTWlTrwXeObjgDEJlCvdfsg
kpAsGPk44Cn6vA9ct6dmLyp0hK8vc23Iin8eqeWtA7udprM0KPNAz4G76YAcCDqfZ6Xn7ctcSQ4K
1ph/OF9oQ9bb5XTEsGDmZ4/yD41To73fqtO6CA9uyq7kamTIehUbHJnCTpwRTRthMMWyiv8lnPH4
bGuevYr2QBa818Sg5DjrcKk0d3zo1mAJcqd8sAAI3fWQWwEyf6Z6aadPieAfVYa32QpcJWxwHtak
Rd0qTZyobE6FaFrDQVzg0pY7YQeRDpshYMYkBxvpu5X9s1WunndmodTVlwtFTnmeX1oDb4qXwrDX
H+yKhRJ1uN7hsMfNlDdXXNCiaGF0b96ovzKx7OJiApf/1ox5GUfyydn80UQqWaEyQUPlr9Uu3rpc
avkXUb8vM+/NHnL63zrGPgVsAyCgawueEHBKvUvYrC5vyW5fcpklXQzMzZwhqnNfV8kwMb/LYWJL
9gLvb9G0ZZlIT3jxGu1BzorEj31U/B+/4vZlEjP8NoqfK/XH+Md+b/9E790/tssjPfGA+ROdTJOd
OuO+EdTwvy8247Xz9Ze0kiORWY3xRE+6jtjSW1TK3LuE42dfWtoTpIRPZK0ouiHw3aQmQIKtMo38
UMawxMJrmVh4HCR/CyF4pVBlaYvpty0N057gAwteZKhnhEmLhPast7QVe+DaZbP4nf3B/olxToau
SkYz2522UWwU7rC7+ZPGbrQ8DDc+GiJjwZXcyXWFr5tjk5jSfE0JoTLCHfVvEUnrn8XwoI9+Odxk
kmaLJi2Fk5VFNeodMtNZNRiwJDeZRCSKHsgosq6q26yxJbwDopB0XxQBgZvdqDvfHc3QLoa+XGIL
z4jq8FVWbrtUnlwDWuWzcDEvNSZMp9s8qDjeYPR1udE1t5p0fsQLWhsLmcFD8WtkQYFy/IIHCYfC
njrTan09WvQy8LCQPOcohWeNptl2i+d8y2p+ZjQ+20cH27kOMh85eY9AntyXSi9PmDbZG+ZnB8A/
zPdqWHHmqCOoz3wOG3mao3Udx04X6bM5qVDvShiX9Pd+S+guJ9WnZyXcl/voK8nd/4/bMysMJo3n
ArCh2qv/7wHyv0f3WrnAIL4S422ZjvJCM0/bGbDkfqIKLbP9+rmAS9ONYdoE1182CHIREQPn2t84
1y7XjNNBeSMbj7xSE2JlXA5fTdHZoFaRlW1QdrQJQmLXJ0bqHd0yJHihxwVQwG1/kcsFvhLn/hIL
KB8rLD7Ung+wgJ/ihGTTrIBUPcwwBcBdY9C/7BWcwPvVH7pHIdS+N9oXqJg4qV5Ir9f5Q7g54DrB
iQNGnZ0c0+QkcSv2JOAn9vnpI1YOYOW9D23XG6B/GamPcMif/ZspWqscSc3lVwfBsmylhsJXT+a8
DXBDtrL2WjbK9/Zb+2vf/Ux6HrvDXnzm2im66pygJNJoZxDpJtGZK70Db+t+uFgdJ24Cp/a3KUJB
/ZlYBA1dbbMfJY/FBMjeSycnpVY5bXKamCVH73yFSkqlCKV8GMl9n51rsRhO8sah+UQ5rhZpD9fu
XKD/a5nePRYYyGNsRUlxgbwlJ223n8MsfU90RirbPMnKbxyGFCRrpXnhIyeRVoNg9BmDDfhjoNWM
rVCn5vQOn6bTHL/yNiGwmxgj1ygC0j0w44YXM17fUp36SWERq5/fufjXdyMmx1Tzxwqe2wwJkq9p
QEMoNeAzKjzL1PjiNxKpsHjl/VqHKKPDDFKM/Jj9nvT3cGNCwqA5uY7vLYjdnCQ3q2KK1/PVR6Dw
wNKZkQ3WfqYOxiSjSvQO0rxN9CrKG6d4GH0u8fPLcZDZ2UUxPf4vPhzO7Wm4ZPPEB+930ADxNj+A
s+LLxyahxni7TutBHtl2jUx8+v7qvIVEO9H6EEktcVegieyXzEtUhqyFpzPajIq5ZFjgQTgjVIKJ
S+/2Q/y3xOMNeYdvpR/WtlEvV88DUp6OUkAxneXnNsL7LE+9G0vZVpIgGoxMH9IkwIHUu4wB4vFF
OzkaHkIR3Zr5kv6yu3tT4XU864VUZVx30jx7XvmTVRt54cZYOuYBD3L+scbSpku/PymV28TxlQCv
S7iGu/NZV6Mkz4X0Vkqe+L9HwqqotWLBBY5g0+Sac/Wev9FfM9OPm+mx0feccYu4SS+dcvO2/UI6
MA6OycJzc919FRsGPdRYB+xonJOCQV7UM4UzJO5ed+bviTB58CAOL+bmPGGV5PEK6xL3uE6JXp82
3fBn8CLF/jT5MZlnLU/n9kJDlHvmRI72dAMtHhXi4fuLpybduPKR8mY7u2qb/O0ZiWN6nqjNnxyD
LMxUM0kdUN4ua+QCKWfmp7P6g+ceHSkmxBV035RyNjlFg97fOytRCSBfsBQ+9r7pHmtzoSr0PnkV
Qs7aXxCAWM4XLfwPGMhGmUFSfgJNL9z+1D1DWU6noWCSASK27+CsbUR8XCJs892TSHrONKARXomb
xZB+/7XLq0EGHJ3jXTCkb5ash9bMpmv6vGzS9jWBS6JAWF5BtjHg4M/1D1UglRY/zNdewpkaMlQJ
koQBxqBVWyafbJGsg22Bc5jwltP5jDqbhZBHXfBmvIH+NAk3yhVZC03qp2gBk4QEdXZZWnRq3Q0Z
hrB9LPLjuwsHSdskw6g7zTmte1+eLVw1DyuBumCnm8JhBFXsrT0QL/WAx6pPojThCPjTDyYEKefB
Yn9gNbP1wo+1jHQdmlhquaopLsK1TREnOCxUcPAxLsy8o0SnlLA7qysBh234587mITtdzxRlRGCt
uMGhRB6/jPfFFGskVpdyE6LiYjodG6wLW68grdrSdPMyd+sgsCxT/1faqtUwMbEOgG9qvstG6Cs+
hht6ysb+5cydFh1v8Hak9v5LN9mRNxsJ9X/yfDJpBQ6S99yjMvxFhJoOczfBwZohokOWLSpUPH/u
bQTYG95crUK3O+xaM7Kg++vfQXNYyGKIpfuMwJD6U7hmK3Cf7wu2O+R4bbT813djGlhhk5MvZqe7
+SYlj+LfdzdgaIsUtIYVp3EAZItJH2INT8QXt7HOfUKKAaJeNQaCv761CdLTlckC+In00wvt0hCL
9MIEzMPH9yinrquqqjHKR6NK5K+HLpAiV383uWYB36lhmHepJ18as83e6IBswlreKuNCQov7BehL
yhh/gCsN0jgxwAxkA8nTNOEJ4q873/PjI+pr2P4/sInFj4zZ9745ekrWntftaIj2VNgROXy79h2F
LQWRsN45dV/e1tNDT6L96/bm2VLWJdFHw77R5DWB+9TM/1QUBb5+vuosiui+72ok0j0AMYGeXw60
lhOX783ivHyS4dFQ6bqSRdtz5TpsQY8Q3pMtDOeOrRbOy+04OZ4KMs9Kk4KUhKiYKTBA0If7lEEp
re8OuhhpkvZR2wlZ5tZD7kPGlPHewXB66TuxQqsVODJ0GK7/7JY6wSkJ4JTPnQgt+zPQAkN+YCeH
tH+o0tnDfu3av6hONzmkpZrJfHXdN77b78X0SF+K9SXJV59Q9vSj1BE7OPEhT8QFHjubiYI8FbsR
jGAjoBEgRHZOAYKwcauGsh+3NMW8OOMoJH1ZKqXa/r6PYMafqa2tPnKHY7W4DhSlWR6SCEmIrwc/
o6+af5YNSG2rzu8Wjqv87p/o35y/KvXmenYUzsAJFbGQ6N1mX2QlaGdivWkjP6P5/t/8UqzoaVIp
UzQ1jYkKqRmm7zw+diQt1ZpCotcbWRTeVceH+egto9ZhDVgN1j0fkmjcB+cbLBLmx35uPidFEGa6
2fXi+6/fK4aSMIRz8/dN3FVVSUEZTE51XPI5yY9xPPorNtGzdceGGDGYnVvXJwtWg3ubWQjfIDWP
7aivMvgtfEm+ye2OHlB4biWjwiI+P4u2bl+zie+NhIcbcQ+175ZzrQ2SfQiukJ0pN2d/iiT3GbVT
PzWptf8bq4L5g05KrvsppnLIGswi0qRZnl0RAI1Y1cRHnS1g+bEW0mnQ7YTKxLrA3VwkyuvZCQ1N
hDx3QmBj1ZhZdJZ1Q/Ma+uAhd13gxRVd6b4OcL2LEk0dEOEvFRVELOzvmNQ9IAt7c4PiNetJo9jd
6OJW+nQ5DV7LlpMZrIRAMVktSuhkHhKRQhwym9PUVzFc0dgDSurbPXd0shfetrTC5h83OKM1IhsQ
F08tdslPc3oWp/t8VLWZn3cwjcSKFD8JJ4nhjfJQRFBeuagYpQMZzvbsDn8P46kopyrARgYvypvC
QgI8fRDUpL0GhGkRRmtiKLTo/FCM8wtR4K4FTij52aKht3/xGYjjqkPe6VOd229RbsbaC7NxN4ko
ztTnvXOyA7wry9RIw3sUOoTsT5W2B+f1jH6jmz1PpE6vv49APiZuocjyYroTHafTmX5bxhmEUBUa
KpiK4dEPVO+BdIQonEVe44JAj1A+9IzJGSXOEwIYPOhuz9rp8UtpoZjKMPwNhf1GcrX0ac5JrRZy
BrpuzW0T+nbdEKJrNMgz0FnyM2541qQQpaLXePaofQScD60fReMJZ+t69mKDfXD7K+WFYg60S5Yw
8aCA7kgSdNfCqyT8G7xM7bDh1PM4THd7dzQrIqg8r/23BpPh53gNlrOZGo0NpMdK61nOo/yBZxFX
a0EfF9LSnb8IgqkYcFgQ5IZL8kriWtHTpRWEEufTdJJGruyoEAglMYlsTEeRWPMqpC3laSAn/IkY
IOCwnRuAcafZ/dxqZ9TzPgl1pJf983zET3AklEGQvvD7dFSK1N2o3u86afm/NgBgmE61OqLJA+cW
wXvgeC5/KWkQs+5SjbHIDC/7EsqwKbSURko2CKXa7ebP7IARb8D0nxxLjzEX82Q+kQTQ504oyK3J
aJbMkDkQURS53tXCjfEvP2Brox0LGJtlH62O/4riNazy16ZhhBfPb4SM8c/nEDKIyHDqy+8mQ2dI
1tznzLCggbg4rob+fnN7ZTOZHDwRiJ0TwS/Jysw0R3viMyaug2wXgNDAFmEkEKrvB6JKvqp4z8RG
vGDzpIbq2fgJUXGnXP83LP34g9r2IkaK4XjxFSXLGn58Ol3E8xXWa8IpYphsO1cHZVPW3Xxf2vwN
3+WdEUS7B3ujZRWWj5ZdYPW8Skt3po3eR16UGRBfLwCbv5FoZXXI3nYtQ1bQC5lifiCigyDthxLd
dqGGmltlTtg8Vzk2dnEDpZIthVSsCQeisnnOkuW/ozICYG8Mr3dAfofCntu/J2LKkOQvg+ygbU+k
993SekYMjA1q52fPbYwhr7kyr/TDgnJVe/cyxO5b6zeFQZ4EolOW9VEDsI9eMMagaElkCFROjuZ1
IQTMeknmTr6IkB1xnlkq3eZYjhVCI8j4qqyjh5pvS+epcDkLwFXbEyycplDlox8juw4y5Rrx4+Eo
s36MYxN1Fgs4u8azexGugUyTFQ2s9QbpRE7CaaR+P3PikJU+zEGzIAPWEw4wQC6x75lN4CPppeQz
cxishSyTjfKkP4ygM5w0u92ck+W+i+GK9K0nJxHuFVu/fpTGAML1BWwxjezypWd12ZnrDMJcC31p
hXoFhf/VUHJVHHAAZWx/ZWRG/K9ZwPvRFnpbFUhKLhNLAqiVgOnW0V5cg6ZgXpZ+3Vjo9AZcadqv
QZF3rVo3gjegTXTowdGTxpk38dPCI3VGDs1GMbT+nFiASIr1KttLZSlkUqKQ600LxFx+ZdWuLj+0
ld5XqvZwEIssza+M9ybUhzy//3FpAjeKw2/HnfZ8QGjAoVbDiMQzxURYHm/GTzd7t1XfmTEvTZcY
6JzmHaqX6nhVjoDJ+tSZP/K+udHmG8TmriONXpH5JNSxb+8yflBhLAbNxoknSd4KkOxH4e1Oht+M
046zno7tvNGVnN+pZ/5k2HvMpBERfgHNyPWqA4PTE2dfMvXMaNoK+YPEuFmkgPmJjr1C7/CT7fqP
fksKMDdi0ZkwzDbaY9+ySlCKO2pvYK3cVBuyNqkTXMOeXYanaJuWrJfemfmiB/OYbFp93ZjGLsza
5P6KgBT05l4GYeAQ/d9MAX0gFfhgmQ6nmLcm3Q0xmH3ld9QwMs18dINs7BvQsQSgA195v2HmFDv2
P4ChIYqTyRmwbv0YE7qFJjWFGfN+yiYiWzW6YVwcnX1Zkxacs/wHj5gi8AxyB9FFbeeYAWSvSfz1
x7CVnnNFcdfG3BksZ0zhCeZ+CubPDZPsFJ+aQM3aQjF3JoZJN01DGdyLWfza++aapJDz1mTTN37I
195MDrYDucjyFWKuVpngk9ukZQfWx/kZ1p7dF0eLd6cOTtfBsE32/uR16mmN4C1jGWfTqPTXYTVo
sN+/k4CBRmG0aTYD/Iq2Y07GBmxpyIRLe490iTCWbThwXs7btOpLS724iJsZPId8dP7myhv3EIka
ISv915BjxocFkXWhoVJqLtKAStPlks71HChvnPbT881VKOR2TstwI1FdF/QH6YXzPQlpfjL8fogd
qZkV8iJabkb5mNCNxgk31YCnhaBlg+3q2Je338gh2GOIVncbd7eO6mFLjTUaNDUTBYXfoC/fJfOV
DGx6GLEkyeOVy0N4EY2Xbj4vxYIKO9Fub7G3DwTkdUWzVFtI/O17px34u8FdhFvDZUR89bYgR63T
ZUQKHhA6RZXHAuaVv47PDqcnpbb9nIODR9nqKcdD04+jboxBxOLTuVVymYsgWntiJbQyUQ0wQsSQ
Kv5D8Tg3UXljCJvaanLAww8kEmAdfQIHE4hxRjmxZms6R1VZqyxkNuYsW+YvSpG6O5HOgGZJPm8m
qVWOF3m7P8UXresJbEu6rDYWKYldUtGkOgjH9K+5d/KMRQ6g7noT9XNw6sSvKPijdBKBcw9IY7E3
SXDSkwzIZdYkjERgiVcC0HHvfnTbR3h8mhB+xNkpfTu4skOSB24rWYHHHM2ShGfZ3pu9PBgDXZSu
la88wtWfpDmFMNZsw92gt+pFpBZAmECAPQexJtrt89vuD7oNy8h0umhvRG7Yu4R5iWv5ACvbeYbK
Enp2EbAtOyNSxAd01AvC963axJJFEGifhBH19XOqiikm23+/e57ASAyjyrL34+Wv8grxbSM1SGY0
jmJSAuwOKAw61i1hihytfC3GngmtD8EMDchWenEWQPShI/nKJFknpez85jl8tSNq9AE4zesy+JBi
7JOS477ZuTot8VfW5kARrmicQf725FBURI9aL3K/OwdHhV9xu11+rYkq1l4pdT7tYAa7tQACSFuJ
kn5qmINyV9nKXkl9Wl3AFPQXKz95YUmYNnEYLFEG1cjS8/up1mytkao4Ujr07r2mVy5ipptkXRsC
BCls8+tkL4OwCMw4mSsJy/0TfQ/XmWnpYGPNZ35BCL+bPxeYMRT76aSkMXtabY2ydZ0Cm9bigWIf
i4UkFOaTqewLSb82H+VRG2g6JBI5xGFUo+fKCg70xeqrXzXUDaMybLBICViGNmAStBY1QCU16TEs
nb0O2bqgxxsjD+rHK6hDwFjq/DDsP3IxVz9ReztEHqRpV9MMiJR7PyduWhKSnN5RtvsAtM9+82C9
milgIUGUfgusrKfOaS6vkEysihtzVdIF6QnBnE+U/SxFEdUIMPhP5XvV0o3PZi26KPhLnXYWp9sG
8PzrJO+riKeGVMcDm8zr3+w8xCS2xDdlbYMZTG5Reid8DZNm9NhUexRg/46YmF3iRSppHw2a9pcy
Y0dwsmeBvqHdV7gh/J0TsGyF2HKETdeeeNzLZ8ed3hGm5I0pIu9hVVedg6+ruqOiU/3arIunqnuh
XrEzGIn09pn2KWejnyYi0rFYp5ZbVyQxfi83R43zIU5XpPYT9w2hlSos362oDfBf98v9uTW5emXT
hzauDtk5422Qfx3sacp7TMLRDZr4j7sCia9O2pJkMpKNh4B6/finWBUvK5ZsNkteWZdWIDS5XKoz
xaUOfRr0PvmlSLykQrAJCSRsTeqZxYmg3bwZj00DweC3/JEFn/A4NEzt9Gps8wfeBeM/vocMxQna
IVaf55lgUPf99W4fIjdLGroJjRo5axWE9kigDNKHBMoCyvYz4GTh6+U+1porUZ0nPJPJ2llmKnz5
xuQDd4hT/8ftJocZeP9+KqYricAz7LjMDiiEtecbv97LVFvvU0cp7oU//6oNQ/Uv6FiyqQbjGmll
UvnR+0rGdoEGY5jQRTxPsJy1fECORqv8602trZNL2oHsKrPkp5c4wf3LN0LRGpC6FKA5Dck05CD0
/Poaf3HF3q4fyaXA9A68iDa5hLBWHW4Lw0j2jkckQk7FcE0i+AghluCQS6wTjvsOu/LmbW7sqsu2
Y02zQkfJakYD+0kZwIjDa6qB7g0Gxk9rN+WkJL2kEdTGg+0LbLgek/xTSFbWC2wCTYhbUUToxZFA
btqevAfoI+U2Es8o7JTFHPSr0K/hXJkb7MKuK1Czg81iPV1WF2+/28CuU1NS73IX3TMaAMGH+nT0
enlZN5/Bh6ZwSl9x87dy2mvmA/DjXIVDstLjaiQeb4n/sLpEYgrrKoPhNiXK90DkJAnrZ/X4/LAw
8/CFsZFHi5B+s9x2xhQfuq1X68qojlVNRObZXPDyTVGsal1Na+SDwAUyi1i8WF1yuV0TmVsx1jNY
Zm8PgAdJ2IHhifiSmNtQUEUoW0UEvNV4L728PyQtZkuTuRdQjxpVo0gweSf/CGaPCHQsymcpyCny
AQv0HnRWmL9FguP3yaD0Tw0+W6anH85j8W7F5IzxTtyEBz7T/841a+I28p+PbbM23bmSb3l7oYpi
iy8CN8Lq/oh9mww1Yh+pstILiH57+9Kh0/Y+fdrzqM2asH4webDOXjyKZWn0jLUPfUBfn2mInopO
2HEhp7mE4wNgCzzy0nc4iXBy/oodhZtK1X7tCRSml2QsV0yTPIVk3Jd1IXhhjBdpfjSA21sz35uU
+KD9dyBzdreIZOGmKhnNMRVisXSTPMR1ZvpNPLmX3Pqkta/9eX+PYP3C6nI0amJ9Pg9yj9e/nZn1
RHRLYi7hDNxW7gclKu0vr6eu2euu1Wyq1MPoq65UUSThZ78mii+zXMukgOa6HJLw070KQin0xrGg
fN5RFr7cxuNLkXHGFprmTcxeJTs3rFv8XcyKEKhe8CBHrT74IG4ZiEtr4m78kWQP9JNEdU+H8kh/
n0HKEr9n9urfGjDKeHFgnPjWyt4N0233tWOxv4UAnfTgAA0jbAcFWGtK5Holg91mgTP6Ju65x/Bj
k2/BKiCACcuTSwAPto5MESwo/QHgchIT9f4w2z0P6F/IlyJ3VSvGaLrv9AMakI+iSq5e2DHVpjwd
i79ATgcqmVuRqEBl+0gH7h+9Lvufq4XRPs571sK2R6k+A9X/rKhpMLl4BF2o0lCzSKMHdl2lH0W5
WV4NQRYtz9dchirh4Uci8Itki3JVgpmX4hC0nBpwoM6l5oYx2QOFAT3PDmk3mCkp3ZiIDcPSJ89Z
LdcyohNA+8NgPE9hg3yq57i/CVpk2RusTHt2cMYhclJV8GQYeaxhU8eLoFziUZCHOk5yT39LrKL7
zT14uFKPT+UTVOsTu50gil9xyDtWWGCkoaKRDorlH4w2cpaYKtAWQ+0FajkQe9EiIIvq5Y7w/tWh
JLH+ROxlajeqrl1cXs49r22+HJi5DglZwRfGaZnpDNWyqX1ojpi+72d0+vo/PgM0cSjgKkHDJbX9
JBtGiVBH5xrom8GxZtKHab41MbGCKVCou9/5yIAgy9/CmqNmFQY1w6Y7xUZFjp+9DoTn6t5ieE7v
mHflHcnP/PYvh5zK7uHyZPn14L/kcNL8IHP6QEhBTxNCtpmLlVTaYHRX4nH0I/RsizyXMj7ddnmV
8Ci3eXLh9t7qkHj3pQhvSCSPkW5vYD0gmUWuldmd4tgZHSazK8o4ynm7t/i8q9GL00kkMOjBiWgw
5f4KjfwDvhdFW42Kph8X2irVdpXIeaXhCBdCYPuS39nLQ544eP4mCc6K/poommOvtjHwNPFjnoBm
M5FOqAvDmsc8CMPGqnomIGDtVQRuJw1mPzm+UpfCLfE9kCHm0+MvnFfCaPX2tfLSRC4oA4+9BuKx
2NK1IQ028b2xjXlwsBtOvvLHRemxpdiUSPuTaISX0ChWOS4eCpgSABZFoSnK0vEq9GvMxgrhY9Yl
J2mGJspDCT5x08aEYSsD7FJyGq7agMtwFtttRyND8Tb2/bGQjVn0l2rZ+rTeW0ekzSmkbkNO375T
U0NN7aN9UmKYMNldpHeQzch8sQfjYotGwUqyIBAD2H57ztLuYv5ESRSZufWOuebaBw5d5UZvIDhD
KcRMsXy2TdY/omX+kxBWX9oZWaPD1LRCw2uuxKN/Ul9M4sH/megq6mFkyzRi7ZTunqzg19B3Z/4s
QmSXG4f9DZXf+t0LzHBCP5KqhhPALArBC2sFg7rP7qWGGaEI45ayV793Tv0BzqmPdgTApyBJ9vVS
e+qnG1QWvfEgUcO1y1arK4qsCoBl5NAtZWkzp+448WWzwSXBwNAiPMzydSN/XR7J0Sr85Th9vkAT
TRM5wYLlPwzFiZR1iYc+qhJROXvlmxs+SIWmi4MmuTsFZnFwIIYFheLebry5DirPpzazjuhSb9EV
JWRxeVk8yHvvsRwosX74mCs6P+NVsvMFTlA2oafirx9d/scwKU0niWkkibQUvd+DiLUxnKuPl0tJ
C2IXafJL3gJwFUVDx+NPGAE2pcO0tEFugMKdxBY7IvmfBZLfLIk6LQcdV4c51BWRQLPhoOmn3oyS
MHjaFlAb/Wd9oiHZ6ImcR6mVOA/Y628HQf+eUZ3cedykVS6sNhJqD2bktu5KGf/xgCn/SjcoY53l
dGeuYjKsLHvapRQg3t/srfDQoOOtpQwUcUdH9qYTb9LVuneUgXK2iU0IxFuAuNijlK7ccOZ/Nd7e
Dx+CWqtFTkuzD//XDtnKASMHLk/tauntKuSbFtJRD1LEFpXIidPDtrdGduayeojNul9EkgRr6Dtl
3/kuK/WJdNb8V5XVSFQjqB17C63n44JJo/6NUNU8X9S4oof5DH7lv6EEOQVQO3Q9662KZLgQkkHb
Z0/oA1A+ZG7lX6CvL+AtLK/SKRI1OdscDpeY8AAyOJw+fGkbJkL1St6ns8JM6esq3eUDWDmv2Dxb
i/t9Ml9P8xWy+xj2D/yRFrIDYSDvpDfvxT7dBdv+cWpbofMfrDPJeFQcAPRlPeRA+3cAxhxO+5XR
z5wpqtnB3WttWD6/bSQHSDW8DwKjBFBuuJ2lBR8dP3KIBq63Ab2p+U5NDhY0kNR1LINFN2k/rIqp
6bWS3bxMV5vxYjUeJn26sp/jnez7Qli0eyi48LfvD0/bFVmrpr3gLHrwPn/pQEltojZxNYzqykdT
g1a8xsWf5mIPJeHVAu2NbF8ckmKD8YGj9e9ocIcqanEazB1RVn98pxHH4hCoQTs5OIDs39g71gQi
+nJmWIRLcHICBUza9ywGVb+ZrELIpW6113tu8OiqMxknemtmVukQ+EysDDwd3inIcNLmmzllYw1/
OKyoY/LFJwE5tSulTPOIjzi+tdgE8ock+HcL3vE+oMJZO/q+Vp4kSe2xMiZSGe3a/dOxf1U62SUG
MZtohnNKsql3dME11x0hgyHE0XDJTV2+L4xlLdCxvowKuHzq4HUkMvit7bn9NF9Um1OictUD5n9a
bf6vfx5M05P1XSpleFqFy5F8Ni5Z9fyiZqz20yzAZQ5YcSzLF8ZagoLCUX+yaY/jW1Z6aPHx6BGg
lbq49SB1ATq1LSy5dMQMVmA+SaEQmP0t3ucwm0PnJd0mJfQjzpF4JhFxDO5WPaVPQLmlhcg2xGrf
H79P+6dnjuGTyYE247hmbBkDF6FRcUyWKTA1V/HxT2Ba2MC+9zuEPWOSn0Gzf/9p+KXp81LGv0yU
DFPMMC8rw+/Cx9Iwzqk+DvJDxU06293qT1zDQeORxS9pqM0FA+X1z+uWqjT9yzMKYzTNFIZE0iBF
7okxgTzPthvuStJ8WpEiESCLcA3LlmLLbKd3P4xX3oT04j35qGlZX+iU99faP8QqG1Inhb6YutQa
73CiAVihxr8dl2s/xatPgQDrQMzXEjwKQ2PuAo1xX9MJ5Q2pdz9zQ2E+AZgl7IkF5E02GBXrRVr1
8HggV9fK04+aLyjfyvkSjQhD/Wh2/buYPKLj/IE5CcLROuP0pzKELrIk1w+sJpdfH5Sp74GL/GNe
IM4aFLRLVhI3Gz+qVmKogq3mX1Nu0sgI9OeqR+0LwIf+vK5XGCnWtNLPSps3Leddi9r8NGnqoNwh
YjaLDOMYbmH8n52lknfo1KLc0F/przgKyHb2+1yVNUM39RoDZjE6ERZN5tf7VOK35TjWifXAerje
fWtip1RFsRMXVvT2nJX6aNE8VqhAvSj6UQuq5TArGC5yA/8+zvPyLkPVNi4F40RYAYALZCVqtDcT
zVzoobMBj1AclzHwNbngoG8Di4Erwbn2ZF4H9DHJfOvrH3xMC2zcx+zCPJxst05yPVukf/OCpQM+
sXXvAS2GGETTFj4aJJ1hatCqFQL39vzoab7ArxDSJ36WVovfe/sPAfnFOvW/XwSUpNpnfOGiY5R9
zXApBZOs8T6AH04z21lQYST52vz2tTgl63oRYHBPESSpl1L/WnmtNofxz1yqSAztjbpZFwWI6R/1
dCgHc1ebz9noTjnKVdT4XuZzGRdeo8vTbnZ5y9H5TAp6XipXARKwl8FYTttzO1fX+m+CA0saJchM
RX/rhUitr2+39cYo0+JcyRba90zWClH+tPYyOthfy45MZ7xJgAOy7mNrhIe/K6peRnCRT5yAoWSb
PgapBUBwuRx7ODASUyHewTRmCxWM3/9vRPVFJnVkM0ew+mUWaM00hCWzxwz+y+BiYanCBZCXzAy6
aRQhODG4cO19RwHOTXhbXTLuYAyW7dwb/ihoK3jTSAVFKHLEjzcU7v//Q6zGpZKTmUy8BVsVTJIO
PwQpAzeVPi234DXhOJxL9+4DeNK+rzmofbIulCx5JrcF0ST/JBl26PDpo63yZsO/sTBe3lQriwTg
/K8TgzpaOE0/9FEdpP+LXw2YwSaCbx4LkU2nhZBmBvgzRtjKymn8q+ggHu2z3ugtXbiHHDEO6THx
vrwssUESkcOJ8Z4xvIi7jH4YgkekZXVrYM/s6bcPqOqiWuHobZuKzB7cjoXyRkbJJ7jt+oo4Vns7
bBiG1h7fojVLNQZl1/9+O1vYPHww1LW4FYKw5nedB3R/tSicOATrq54r8ZfUyZbPdcT0SxQaxN0n
OneEvltcgIy/kXPtCTc43JLhepMwkDdWQbItdFhk+pROEgzlIBFdKUjp9wlv4m1mNnISQWDr28w6
cyWrwQtDu4rEsrdvD+HjtoP1R77BcHgxrAE1+rs8cHNAZizOeCOOu3i9KXOkQFjg1ilFZizY5BY3
ppluwbuu3zK95Hp3wvoEaLWj3wazvXht8g/6GYgRhmve6LaYQ7NrLpbjwmdTsvggROe4RGP5ifqm
/0zYouWBTy339gWKdaMZeoXJ3SZHstRk1jrjjpEwZ785PD8D86ksFwWZj9su7MqJb5eblhjXGKMs
NrgIqXNau3Qj5SJbWOv6ndT3YUnRbisd/aDeyMZzbhCKEhfICQjbNl8s2HqtgUpfmXhwBfaRU9by
mJ2p/EygHVkN+xPi0UNZdLi2mRALvkYWXZGVJvo2Dwb0pXDcAL7e7LICY5MlOowz3TqBcCJLOxzb
nigtDAOPTr6cMom55i56t/XjROcdiad8s+MIl7XMlQ+/m+auTlLtrFN/g6px97nLdAJ/t2sQp/u9
x9VW+aOZbLXhTI633Rla7RN57ojkaodYwYLLwQlhUYjM7cwlZ+89G9A21SbD1QA3/KCkAjSTMfS8
SlhBlMCL5BgxRyjMS5QzsjW8Ckjl74NVL2rFYpvEdzBcQjfZLWaBDHtONLIp8JMd67mUv9zvqYtT
85o4DtdK0lsatA79vjhGHyRw/43TbWdgmsHF+pEfyUci/Ahsq1nEYStoyexSoBLEtMOuRBuS5L+g
PnIUe6h6phGIAKzJMWtam4IroRLuurAPQPo5e+0A1noTI9CqBWFvz8dlAO1kWv+WcRMY3bKvn/pK
E97H38MXA2/c5GNbFn0cY9BTS3gTGDuoQmCdMRrqbhtfFsW1cHWsJryorx+mmotyemOcQ5G6MYXm
FjkkaMkE/QuiHx4927yVXvV5hQB6Ym0AdiXrlKOi4v85QSHq7wC51se4WVTDyvVPqNOItzXKQw4m
05CXzC4+5kr92jxfowXM6ePzU+rJPhLaKhtGKYMhj6dCDBVrW8b2B6c/jbrSIf5hyVneZXDHzUFO
qVnBipdCRVHjV7Ko9UY2KMKzwQBztGipcsBWQW7welYiNamWj/83UGDwCgtiRyZfkn15vxP8lZEP
1TpzzWn4RoFICiI0hg/jnoIGrbaAcNs+MKUy2E/fT/mEDkKGRcPalmkuJ75DZU0fPnWI2Eu1hcKD
9haJwzZj7TpD6rMzbRHNIsd02WU0ut3dyofwOGXLm3UOGadX7fO/ioXfh5c87wGSMuYzUjNJ5T75
Uxxn0+Nzaa3TmSU8GRVQjvygQiLjg6a06yzL9mGkCi+/eUwtYQQG/DlX6ElF0ucrY/1awzILe5VI
hVVELIPd0OVSvRsrbp4FRh7NT+IElcl/YAR/Lm4lqPEjCZiB2b3PgaCsQNMIoOHr0kPNpRrbXx05
3bLaK+S0400RCSN14kzT0145odYRK127oiyQ/Q60qAwFSTUtXi6amLPW5pk2cHQeSaele0qOgXJz
ap0MmHNkW0cTPB3G81c99T6Hi8NJHyv5H2mjLgkisP5djrSmx6KGF6kwPRyBUWU/PqDvOcAlZexP
Q6Qz0nBteAS1P/Sua7FTY9VvH3zBkhnZiobuJECtyZkZW0O3If6z00HS6YqLQEzHECv1i6/xqWul
WYuR9AuOI01WVVh3E4jvwpo1X8jVNuE/De2w9halBTzYdg4kQm5hXGdFlGIMYuy8R8xn6Wi7LblE
c8tUqsqGlgwNfbk073deYyA7WYLls73W6pHVCSOqiskEo2cSfeUlZJYdik1QmzhCbRh3Bw4FTGu6
5RoNPnn6ztd+d2D2FmLQyoCN8hafknNEobUDk/biNWG26SFujySMsnY/Ua183EL/Bwa6VV6qimVe
BOE/hYw9ld6Ek3+JuI7yjO5lCiONvyacULB6owKHydFbcPRiwmRe2cYn+ync8aGn0b+2OBl0rRb/
aq4DZ6FUu/DcISw2IYx9L52+vyCzn+zFgwKCItzYQyABR6k7NL4bct7fZyp++2ZWfvqgQVJeSZ3O
IXUavAlKMhKjcKL04PQIJ4z+TjWc9O1K7CEwpJnq0Jl51+D15tJL8RrXULCtfqUem2++g2qVUzeD
fgWtUsMjGgxscdUsVDNnjen89C6rAmO60a1Ae868NMsq8rcCqdKEStiJQEvRS5SgnyFIJgm5aeac
5uHpXBbyU5V3hjHxRZa2018Mnqh5YK1OCqacuDjjmHJu5P07dF2ja5sM17NU2NA5BzEH6HhQbNRg
aDdwcMwNx66M1A5QivRZ/21YXbEqoq/Q6HNb2swHjiW0jzIfl3dRf2kdPLiMGhEJNEDXWwOrG1d6
5z+RPgtHgZFSp/JXQJXuAWQxuklzPzETLyzolDRwenYPg1aHI2p4t8mrtMx9m6Zuc7KogSeXqT60
FDxAlFVzNVBHbnioXbfL0KY/vVLxCr44GFdE1Y/zUx4MoaUUMKPi4ltHliAe4rLqADw4Bu4MWF8Z
FUQsdZ0eT4am2iJpBtM6ozV3+oqB3a8Ejl2JCtaAdcZGjdvC4q6vkN42mvhQqu/BJqPrPayPzAJH
RWQn5lSlRh9ugEoNaujfauLSF0BRsVyFLCBNEY4Rmg0L4VrzI3NhO7xzLYVtJ649A/XGK2oH7rQP
6HXw6xMM/zIdK0UXnxiWlfqVy2yoAIVecqnQVgAssWRTehm5Seku9mk7BBdNHI95l4iun3TUWnBW
Y5ez56W0i3cB5ErW93nx6vDDZvxA8886Tsmmh48YnjmoW3IW554lpQen5y2vlJVgVoL6lYsQaZ+0
jScXEhjNBzdGOXmnUNu4FQ/3REoyHTTGLGrYHE5+/jsjVA5+SNBWvFWBZhovmGU9Cix/ngshffZM
5anY+9kHoY6DW4zYu+IG4kVE16DGat7wT1oqdo2oGdID9ygaXvb1qvYKMxQk4cfORtfpoa2RmKrm
QxmOm26p4M12ohT2N4P5pQ0bYzDwN0BF/NnyetHzLVlBXqmbm0+0tChGIWPX+hL8AVYFcm7E5bRA
t46V8jYBQlx75NN2i4cR1OhzM75pEev8v/kGw5MB07sQBz9jz0tjgUvkF2qwUp0M6trvnUIocsvi
G/yvMqWgaDHWRhTb5jyjCZiNiBvaWP6SafQcyRgUFlkIorgvlU+MdhjQ7J9Yvdx31UG6IdpqgPJ8
MRpDVP9mov9xIlKMmsAUP0TuOH2pvcl/JogiqOrDcMxXgOcyckyO0gVVYv38Z7CYt3gKOWZbAawD
t97p0QJmKNE/7amDUGYl7LSGm6h1fmxtlIKnJwhwNbZ43xgVhQjdTOook7flqx3qVdukW1AEBsF+
ZLquPek/dCPHtRUcpad+AZhmeFfeOo8H2DLaPxRdGegv/iV7TDHfdXbfCEU+jp4BlStb8wHtlwVu
jL/6tD5ldwzRGL/xdahxuWTmVXIQWwkZFDSv+fU6k3JfEwH1MkYpz8z/7UYY4+adDvIC1fKPXHJY
pVyOz38arjLDEnjiSRakOUMIroKXyubUq9fEKdbnTftdPVI1jQKXYUEbLrNsbaPzCnaKiVmofuHw
UBjtSnr8jcUacuqNd48ROxqCXWr/MmGQQoPC4bhzZij1N3TRK1LgP6CJTdIos9T+CZRYY6uz3Dox
dNGtsTboLM8JN66cecu/mFVyOd1erIQcTgA8xcjADlS5bmoi6zXSYVoMCnrcf7+4yKctdZazANEq
mjzwzLhka2ekID3ACDWWzGhw/dY/xAnBhleBjsw/IQ1CZ18RAJLiRBcYjLyKKHxkl5PZgYDwuTtm
QBD8Y+C63oH+EQ8Acy6AdXCWgSO/f9FBCPmmvzLPOwBJSXvDqjLRUZHvRqEirwoWz5mRdoK9KmT9
abSKZikjWOwscaYBbR4gYibMNQQZsN5UkLTMG4MwNsJ+wnn6HBJUtX7974i/Jn13k5/dmg7xYMXf
Xtqjm2O+m2niC5DpHksGBX5/uYaAJ2oZ9qcVKEXTY39RXI6GKiyFBYel9O+jmhIVEWsDSQWud3et
D1/lDK9mqozaA4X3GE//tV/U6vfnYdN1x0x77URQiXWAJpMGAfvYwBY6o5+vRtPWC73NJCQawa/h
hr+hI5byzcIWP9I1qHIpwJt9amDX6qeVS/dKm14v57TJ+w1dW7EPDCFRWUD9gAgoW7iz5wn/g/bB
2OHyB/EONhHD6XNb+0D8uUc+lINVy98AuON/TMF87L8b2knIZ1mxwwqfRD7C4sdvJ0uSoOOMuvuE
4Ug+oNvGdCE5YHn4rm00L7ALSGPFOUwGhnHp4JrC5KCb2hZQjmocw1HhvfAFIHznUCs0BMOSltI7
N3bbaaw794mYjvon3AjJ18FhmOStK0CiyD8MDeZW9pEH9AI3PQs5wNK1GKIWnfQ0A8cZn8sB9YI1
F/nRmS5c3zRt5W8+Hi31H2x0xok+gdpECHIW1UZs8dAbsEM6z9KL/RDW+dqd4vzVUj33ZidURkET
TUqJu1hI/t9RXG3xSCI5oiV1Bm6xaqOOu+5Kk/mkqJsnh2i9+WCP335xPS0yKI2vAiMPRXlB/JUu
QF2bX4QbEAGYOhJgga3yyr6MaehlCkZkmJ2JVO/h52cB8rcJKGLtta13Hw+Jb16fqpdKWaekidI1
ZJnFjcp2ron/Y5m/oRac+6W2RalTXgi83RdFhdm0EVyhRmluFGB0C6JuXrXXddTZvGPVZy2Hh80P
WczqbRtjrmkfSF3/cM2I3m2hrJ7tJdcu4Eh4aoQaDfnPdErvtfgCQUXGVDNmBSxnSvTVAA5C3hmA
HAGOS6jvF7lFW1L4Q0st7sf3FjV+KGBw/dkbXty3npKNDxeY9VThTo5QCZSnpAINCZLx4lvpLA9W
plWUtc7/S05iXpvYwqnG3XjueIsW5+Ai+KB2adDtSb32Sc2YQRz+q9+ckENqsrO7CMasX/4Wmjd+
G5/eu4ZhDZI3jy42lvflfxfWTqMGBBEoV5N9EnMlgaEFJ0I8+SJHdba5F13jAs/H/ki5NnZXd+rX
bWfXKvdGPRCqKjiRZhy8/hP0Bg5NWuR2Gbw8ca107Y+kMKCSob0O/AzWN8cBJuMELQv+iU1gaEQE
kbrYCTn0oFMuemxsce3hD6HSM/4i83486yLhlILpoJ/RtdqAEI1CNq0FC6y4VUInbOthk3ogQoZm
pAtvkKWWmTQDENnvS08tJtwKRH+QGo8gHBvWURkiEbq3LgqixXNmn9AtodytvB6R/sb2kAKxkoa/
Q6s+ZMhCz3soqI6L0R6gwwpp3kE6M7GlhY4LJzr0x2Zr0KYSpjXPJMcV4YEdQaJKB12a8vXgmVru
PtPWfpRJPqetXP1HnVcaBeIGgzd2nv++n8VBN6lmrKaMW+rKE4jvxny8RpBkP2iGOynDtbJoto3f
sqQsfxKY9y3fkjRTMKGQ6xnwZhv7ETs8fp1+ug61qq3pyUNFqwlZA7x8zJlC67dwfjWVup1Nl1YP
495aVwP0GrDjyU/d3wK+2R0WPNXdKSVgv669zfG+Nw3zT+BXmIj3uPeku7kqyhamqPWaZoFLqSlr
kXWRbMyzmQzpcsgjUKFJsskBnx8Nt+snMzEaepJAV9OIHmmHIfxeLAomhWFNJe5tj3tbALKVEky6
nXeC3fCJrj/cOTCUwwTrwN2S3ZGPfrt7BALLr79VPiyo5pUSOREcPx+ZF7MyqGl9AJlZkQN2kftn
GPZGnIC9sCBd4Da9CdcUa+gv6o/VoRpG9a8Xzb02ZMlGRH+iAnPWAYtNQRjgbNr3As/UhgL8ZT7H
30KGXkCu5fWTIG+9Mll0oNTB9OAC6GgVrrjNTMbQIpklVbJntJaGLeYKNb08cK6qD/LuXDqSXejw
AhsPYTQpNrfbpLWinCoo2k/MrtOsoV2TwJlQRWOQdyHB317ORw4E2Jvr6OOfcYx54bi1owssVr3k
f1Gof3dG5UgWe3gxNO75qZsq4FOw/NfNSipY3L1MpUGQW5JJqFjnSe8qyIW3j4/HnDqIvyIRnSgV
VT/HhfkEIERebluEOtiE6JFOABFuzL6H0P8mJ2UBR5uTXZf/nwzn4eoMbFh0++/loTC8XNHRYv5l
ufW8ruzdUOZtrQFblxqJx9ebQqUo29VETpyavpWONzwcHhlsFjrHou5JDPNQw/CDYgLX3CpGa4z3
gSoj3Xp0/OmoqClmesR5anFYma1o5AQOiKzcz6CJgf6TyZCc3QuFK21hK/bjeXoKJi4E71Hcp31p
LMhWnJ9+VcCi9s8wd6Q4tS3WqUu/GY/UFCVkoKVh9D4R9C6+fCUthtwH3s/E/HDLRxNtsfTGjJff
NKevl58CTyLeqhXrUnpl9cIZvk6K3a6cfrZtvX09vYMqgxzYM8SfPxHoG6kO+Z9xlQiKLQzsusK7
c4wpYY3pTUOSVTCjA1AK1QRDCj1dEFnjBCv0GgmocOBdh/kH1RxTx3WCTizv/33r9EVJzCPbrR5z
AQJGMhjjE13F6KoLUxhB/tvCYbA7HPwOHhas9tmi88LzZugDbiNk641mzwibZC2FDfhKd7A1C2SJ
/axOYgPxJsKmxb/S0vNFB4vpr+Dyd6SqXKhftHeNxPAiCV1yP9boiqWHNZJZbj0PJxqNXMw4CuNp
xC4GwoFpLd1DnUiUfBG5dJMDuK6Z5T+krxs/cwyg9ZUrNSxYSn9b/0rCRhQhOraluUTtMx1qSDCO
dYbCJtc4bKkZrCH8fHZ0LUqhgdHJkGiITRMclp5vIZSSbPVGmZmVivScPFZnwF+/vNuvc7jDwwi+
Re038WioFVidxWurUGmRSjXp8LiIcCOnQ9S0SpY+sOOPRIKKVAOWj8lWbsHtEaiVHFlopE4oe6JA
tzMb+AjaesnpCtWotPaGfibVcPItHpRp/sF4/dotg3iSV7NUxi8tIW5LBSf6CkX+VIb9P768G1bI
pcjw4OKU7yjhVMQPGDKxpXmMfSsioSTy6JEaOIU64r6LaYkIDpIqoFUNM3N3wmena2L1cQ3/D4pS
je8yEkVunBH311zZLFs3pYAP9MZEY1M18+8UVwM2VaE84hzvq2YYJKfGFEkosNWc8T4BulrfQNsQ
KzrFR8i+rkJrSplE49/pVnPub5LebWr8gpJ+Xp8uCTUBghpl1MZMXVtkg9pGDlr/LN3TXm7D4CUB
qbQ2cCsUGP+OHTg8fWCzK8adqwCleg4fGUm/V94x1VHOncjkGvqF2djX7Tmp5GXmiEdZmcxNnYSX
7phgEfbiQBhrKzWlYN9pLXxlvKKx5MRaQnyMYT906LZaARO7nD/VLWndNWv0XkFKFSIha3Inu40z
LKLCArVtYVDL9PsaUhL1gQaczIOnoC6Yy0svSsbEsTjB71io8LZ6p7okDvSdP2doYVWd+2NUfYOg
nlRArQczJfnMjBOuTPUWh5+PTeIr6/fYmQMGpuz2a6PkamrzPIsKTlLVui+3lgV4Ujqf/1Q7/a3M
x8rQR9woc3BBQYzHwrkTUPPzfQPW1R0A53ZQT6LXrrKMVZ9EGYYuWX66dccsGyVEZrUnNVLD1dCc
pJiugMA3xDmeyjl2GVb1k+cjGU+31LMX4KycFZZfnsP7GZ4yYNKih17e1HAofKFo/Hls0vq3Ge0r
KDpl/o4fe/e+uECV0I/VByhzZv5y0hFswezDFhKhOVBPjGc+4UDyzr39YIPX/1En0kAMzW70er8+
UCsDfv05GV/N1z5rl1if8Jnl1C5tStQiE8YaxGOiJyjJPeLPJ+OZXyyXtB44jxBaJLSAdYi0kXH9
6qDCGzYhukFnzf90IxsUoj2pm+1Fu+jRL3Dvn1oiq5lqN1uHcRwX2T36zW+S5Qvx/65jVNKzghfH
QEOpXaIP07MEQbaR7GR15f4YXt/R+TA80xBQEegm+wXiZ8+fBK5dEiU4mYlPqDwFI3ABC0fAsmWV
EeSLiRNmmB+Vd447EW+L4mhcG3UruR0XxVknRUcvLPkmKwUvbEWVupqRbG30hY84rId9jJS9p6ox
aZbpTAiZU446waLbI1L129qV2t44gcsdyet16BpdTF4H6TOXp4Zr88ZDzgTT9ior1KL6o1YH8rO6
zKRJ/aUW9NNHiLTKWJ0KjSf4gk9x8N7wIa1A3x+sY0NqNXRwvhna30Dvi9Z61gabKLopWRe68tDt
msxpZS90XjMMcBSjDNXvjn+R6MxXvwgZTPWr5TEyDaHPpdqgjnQvQq+plSUdUWfuL8+lC+dR/ve9
dFmw20i0KP4YAqYucDJeQ5kjYdMKyongcSQuvWYpJd64QuWq2zpDzmtiF4gnio0ZX5Ei5yph9tnH
uc9UnlBuiNywYi/+zDij9d09mSpCnXoVpsDwvGueigbX8duWeQ5Tve4GHkSHBppIyO1ewY6fHdLj
AoNsX669ZXi2ky9GZLnFQ1E+DUpe+d6zXHslIYFUf8vXiBzWcySu9IumbWhvQ2GFbg0VLVhMHIjy
NRmk6/0t9+rH9fHjE0xNW6znq1LylV/Rq+2Q2UVl2AmHDaxv6gozIZKZ1KbSja1FS8KfaPo+Q2rb
sivKHamrKA43Auz9zuT9G5OXgmRy/E66Xlx70l4tCJu36E34gkEkXMrY0Vqa/flpxYg9C2bKpMbf
cvhYWzKFrhSKAFdDxduABnKKW0rjsVkk74SA+wQJsK8CbAsOnnVL2HKHfQeWOFMi9h1aBbg/LSMt
9wSRapzEm74euIDF2I85mmRfXFIE5XkthAd4aSgQ3HfCvN8LSJdWoLUa0Q1ht9ERgS0wOf44id+g
AOrUbxSU/KtUBPKfUhdsglOg/IcE8nsiDdJe5A03LJEnqO8wUmrSuVBN4mh9g9vD+fo/nswrn69Y
6dnU4uS+TsKerERBpn6r7vXpv+3vZDQK5fk3gzQlwkuu+/cL1ODq9qZaPVXblnbdT3cbzd0XvJA8
+DcSXfutxk+bpMoXP73pLmguZJhIJpITlU6dmLXLhOa1rKhdUnSW3Ev2p0ml5ATZH9nzqWKyl5tZ
y7EVY8XnJLz9gfM0Ic42Xewa4X/7RCleRfxratflz/4lcBkPoC8WsIaLRlRYMZb/TQqcHATlW0sN
oOCcZ4VgXdVTwVQuEWIDKaUuZkZNJymT5W0xvLsAwTPiQccpOvBPpXyppy2K+TTh/p2XBuF0H7G+
mkc+4I2DiBsCzD3+l3nePGqnQGpBB9UtlEw3fJDBsbrXp1z17g2GFTBFXvjxP/8CUl3e8v5QtlDs
HtWyK+fiNwA5hGcyEal2spKvAjCXOi+h122e3shzgRx9xhi7WDWAjtqERuTtiSUCC4voPenat3MB
u36XczKJuZz3T24Cqk3TXDV8pd0VAxooDNjCEHuuqE/z627CCQk61UGmHBX/niammQzH3PAczYnw
e3mdDHd5X1zqtALMi4UdivN+bOta/azjybvDBVoikkD1iCn24JaEX/bcq2YMVNc0apVmYaxGm71T
8s2Cie5mShIWA00v+EbsX2P+zglKhkyzXwVvYRxZxqi10hTHX4QlmftLRpmW+o0yA1NtPPtxVEtf
n/fakP47mj/p3bps7Ep92yeN24Agkd6mzHqPKu+4j6ytVD8Lg4AD8nvZdfetzDEl7GWL6U78JJiy
mnukMoJPzk4YARPiiUiT9F0y+gNFV3VP4KlEkCL3f/4sJi7/LSFauAwhrs3BO2nEG48/8ECJ28eS
Ob/20fEbLqgJ9tIr6NxxrHzDQCmQvHOoBSj5/uoaA0ChsckFATeahwUWL91BbHE0B9lhGECmLqPX
8IhaUoNR1JIuOD6IhdSicFd6CHoD+E/WbIUeK/Snoh45Rq+e4r4Lawjs1b4L0hZ9DjShx03yXDP1
IGvr2L5M0uKREY8tgwmDGM/TBxS8r0m3WTy/mjkhNL863Odcky/fp/zBBvVqr+yJInYCovvnl62K
TYg3o6CSMfhm+lHishSF9HaOEevGuzhZfJLWOBugcJ2mD8mJVMLErLESw/ZR98xyN5bOBUKMVmU7
aoCCj5lAJFKLeDJHUNGGJh+2jnBHF8NsqTp1kvG+qTmCB/7zgY3kUp5zl+WDye2ZvU1vRauye01Z
Z8Yrp00i2v8L1NVQ8ARlmPn0q9/JCyZ1UcViaB4EWff9GytM3z4l6aBM1UDls674TE6pmxWPZwEL
y+4GdSMKx1WTls7oYv8ltpxEGx2YD5jDn/jNld/+ECNkIAzTOuBzFX89lyQO12xAqriRLm940YWu
QtF8JIF3c1GmVUzi7jiNRjbGwG81UsGP5mPA5zBTnVKQQ0YRrOeaXHyR2vBwzsyEKGQEF//Txqd1
tI0P7Nu8GEaPDxGi439ARjTFosB5k0eHh/tsGvdAaqonEKlxQsJDwHLjBlLRgfB6JkCQspFWig6T
H1yB08lDC5ePATaS534bLjUZpsjyIuMi573Sg0pM9NuNWJ1d5w14xuB5aySDjao8nqH1JTWHAiT5
VGewph+cR1uPIPVrWgxcKqKIMQdtAw9oAu8FSZQS5W0zSjkCP7UzdEloT3a7pfaDOcqbIbmqGGrD
KjBD0AgIP7kc3GywmjtyyZ1TKtQhXwuaxaT9OP4Szlr314bD6eW1BhvdCipB7TOu+YzKUpDrtSqi
a2Fgd1HUXbdQYLZilTaZg6W2oB+drJk86dyIISbZL9q285puCDyrj1+9RGBowpxCMZVfBs//5O8b
Tor8Iba6rGyNHQXyApoWK6goeAhDWVqC5r3t4fK7JqnNrDDyK4uLUBKzbys5qXYYEEVZawMj8aaa
ZAV1/5MiGz0NrjeiJgKS2SIzBqqpFs85NftYmOBoEb+IWSXC1O38XvDNXMtM6wVzhTO5ishT16FE
ZP4k+H4kDDmlgpKOIfTwD1jIWcNmkp2X6IfpvJ4K6/hB7OjRGL/n/wTGonriIOuHlYXvLsQNN37y
c1w6lS6dPTKuJfcaIRKrYSo1j21BhzPZgqEuCUj9nh7YsHnB8B8r/LU5LNK1DOKwLZab5k/UGIuH
yJgF1c0qMuajS9M3oWvs+OCBbRvHk+2caFtXegYgy/hmaU48ykI0any8616cEkImAWEu50zcABh8
oCz8D/PVr7FIaQztWafbanZ1NkMCGaFkl0j5FeQT06a9QzrtA5OBnYeLE4E5o0lB7JA6qQ6AF14v
EJx21jr786vrm6fksqR83NCf8Qt8076wW5FPYq6wK8E2ddzP2qUcKz5vsz9H+eAL274zFUOPwg2u
xhzP5rOqBcYAyVe3KqrzouD7MgYz278hMhVcl/fn4AjSsxjz5k42wVrhnK2nNNgAiVGC8WwMsbcM
3im6Kd29+4AnqXjv/EKX2Bg+702pPK4DZb89NJZq13ZtAiseE7M49qAzX10V4wHdbEvTYZwqnWo6
HUVOeCo45vPK2Pp98NcYw/kM+Ik/XO7rpAseXYYvL+ngyHrZB725VR2hfXWcLiXkkSeqCWdk+HKI
fZ6N7cUz6LvYSGeRuqJSr9xaPfLX+SbhiXoGrpcHriP2Vu3rfIkYS+qnA+eN3/K9vHDW5xNEDS+T
O1nSv242yO8W1AVWMy/PmSee+BrryHSxvM+qbXlC468YFngPLohKB3uNRWdV8fvHc5FIhJo8mLx6
Cs4FD232f+EhS+8DR5v+3EKtyKO1Y8w4z5oIWO/7dY4kwnG4uHdjr7K4xHFZKH3QY9PYlNkqJSZd
FE+9eOc6jkgv0rX8Xo/vSIGVPDFxnBvHCyyYEMh5Lb/p4shPozguu/j02KIIC5ayh0Q0VLltzeHB
1k/XbYsoEj1oEO4F4j6FXMsfn6bQ2sEHpa7HB/WEptxgmkZfTWz0ibNmQo8ElfWjUbhYl1G++Z7X
RJsVVl1oiyiwWX8qlqvnk7So+y6OMKoumAwywTesbyFyz/HW8qniGvdOPZ35U/sfyl9OD5X/TLO/
dGNm7So3/R5IFqRR327Rn2fl52wb3blPJCn8Sp4MKB3xL+8FHnd7xr2vOz/nzGBhlsBpbPoRs3QI
F+K9uGwdfe2aK+GoYdVmBBeWgpX8H+zUN4BK+RXrux9/WFPxgjgHWXlf3VstzxeJ0IHplHoshHAL
7RnFus1R1BUu+8VrVloYw+vjJ2NdvMAmBswSRzuwQ7sNiPqWxf86VpMl1lFQlxeISnEgEDQMO/PZ
SgiGzsbcBf+jO5G9IPasyCf+JQfYc8Mn6i04A//gNCMO7V2V4zXrk8Zo0yPODYDulQZwXvnUyyzc
LD3tl+3HENTbUX4NXDsXohHf30Wc+rDalQp0CHRoe/Izta7q+cvDdTizxfYfCMCQPj12UMc2XidR
xfDFwuqO4Dmzx6GoF+1e7aSXtqJrsjc9iU4eYybQu4PDGXYyTvbAvUqEzt24Tst0HITCQfhto6xc
gkVCvQI0hekvj4cCo5C9idOISze7KD+nhiIVjJpwGQc6IDZ3EpHReHGIYXFmM/w3q1fUZaKGuKjI
t1l709qYEpWbpBvXHajiEiqwE5lrqFYQ6votNGrChckEOlrzMa/SDDCj+Cy2YdpAyeietobZlnVD
rTAgaW02S+15nsc8BMvbw386nzd8SUdjfOd5ZZKLCIYpvn86UoQe8jjYXI4ojyPve8mt8jgcP74v
wao822Sa9C5PVxcpkXl7O4P3I+HcUaKrW4eeLNypSjhip8ofdVmjRq9QtTmnfa/ZoZAKcCbTaKcq
suSK30ZYf3XqYLk5mbpYXBDVRl5n1xe5Hd7ZcZlLf38HXfrSPyi4utUCudJHWQc7QyCFQYxLQXo7
x+dJuFoyuk/p8kBYW0RFVGZCfJUv1KYLd+u0pRx0xG/c80BdHHZMQ2dhFAevSxGWixZ8XYaZtLKI
UxLzAgeZHwJIkI+NwOIIyS/R9ubT0iqALBmzGfj+IIxel/ojBVakm9/kwA1+2AQadOzuN8PmRbO8
4hHNe1mg5ikN/8f2DcNGRPoldPa5yjxCoaxToPJydcx/8ChiO3jN1ZBn9J0lsGl9csj3v529xPpe
HsZs7PtWoGGdhFSmHuUt5np4vnIZn8Nud2qc3BFwTdHITr6gXugvlAZy3mVrDDSIqq2UddW+VYef
B9pA0GP2qa8bB32T1ln+KzTz1aG4ANDyqLbowBNIUM0MsURXxhkt6gsbj5G8th3VZFqGjlyjbtsA
T9glxadO2bQnIu8b9yzxkbCfK1TAXzP/3klTcASzaQVDyLXmmIddz2N8pCyeQEivU/tl8WMgljB4
E4Cc2VsCYaqHLYA6bvDVkRgXtDJcWs9HebW+FO3ONp6x5HaGMX7Dc6zQPqddsMzp8CJhL5D9A/TT
/nhXlGd5bcWTJk7rhLmLiKeGCpGjE8VXyYL3kymnQmUMwscQw/IzL/7mMoCK4DTNS4DZkiDet7W9
iasz+aiAyBt6Ciw18yH09KKDWIgTBVEfTDjNVzhXRVm9TtZKtU8MHysESsX7wXamfZC224njSmOW
zQvEVzxKOXQ7rgjsfS7NCXWykGhlbRmsnq+MZeJDAM+hgGLSAPWwcWyf8uA1nE42JWeX+dvfVfVo
4Ti25FeGIwBBnVYcgetuN77/dLQYzaOhVsdIkQLnWT7ww1WG5RlGSYmYwo+/7vL7fEEmV9QuzDne
aOoRDLcZVcmEnoApghNWkw2YjoiDF8EJEN+TOSiByZc0Ew2SCWmq3L83EnGB2GNgD11BvSlOhCBY
CfMVcOu1N+IJbcWweCI2n5HEaRlA2dMD7NzsBQJVaRtHGR5yuaxiv543ZBXhNG630CNirHiW2dQU
A7R5G0Z+kE2jkNcv5NJ429ZI1W6bgIXzk7ni596RxWiKtnlTlFLf8sGNum8y/PmdTLkLUKR16UJg
y9oe8U0t9PoCoXEwYpZF3qj3oijqjwuyOZvrrzmmuOOJRqsqK9U3vZPYiJerafDJNtj9IQ+u9ewH
+6WICV5qvvMf5h7v1BTWj7rXpx1PdxP70szGI3kGVUbcKCMaXIEJXg//iGklxjSoJ92Tocgx1Lxy
9W0l9XKw/Gy1utnW5IQkosreY5+e55LWZt4Z8M+3W2ueRqR19MftdAuz9qUpfXuOaCtD4Rik8iQd
+SeJvlzZeq4GoTMAcXm+RRl0g6b2kaFYWkIPIG1oqLHcpErr/SUS36XKDg7oQ39tF/jtxQ5Gk6rC
mwThAZLe+16a6pmFOOCjm+Ad8AF5gurfneDHo/AApnfQluVrMXJRt+bpYfsfyZT54nI/Deowuj/s
kOswQ7jyCzp8eNKgmkhMpImbvAoetXkGXluOKeNzuqSRRoE+y0OLvtmiw1AYqGR3WpLvgSBOygiO
OIv8MdGT6n2xu37Ux5IXRgjwHs81qToWmgg74l90IDmjOvwwx7gQgrgkCbr80qm/mii1TbYnxZHt
+L0/GQ/rW0Q2EcoP0cdUH9PJRelBSdLrrh8KF4zNiE93AJtD0ZNhDGpyTou/h2YnF7nMb3zO+tNg
ERybrNVCsx1SeULzm9J/C+F4AKD7hDl33RGOzAjY4uuQFrYKQVEVcUwE5/YtarAMsFBJyZOlpDnw
5jcxryO6WXBUj+5bi3f3mV48otchqh6iW20N3sPD6KQTNUVuYJc18xxFoXcm2oW6ZUof+mC50xzr
mDvz95u33MZ37+FgLa/xMkxJp96LbUxNdGA5ktRgk42RR//12XRec5GnBIbwWwjpaP9NST6+mvGI
J9tMdDtBMHFuPXPpCue3rRCgx7pKpvh2V5TBYpA6b5XFZdf9zbMr3FSk12QxVCohhtKk3EnpFpVz
OhbaWhT86XU1t8iipMkwZzXVgodwx53oIsyc+1a5UQ9Bb5Cm1Mh1DzBDX/y9l4jNOr6q/670XrDc
YMPiPOo8BuJtBRl8G26DRW319w5C7DzafU+8D1yE+yYyH2OuekRBLa12eGJH0FDN1yvp909g7wCJ
ZDb4kK26BxWvl0yks+2FiiYVvp7ZvXglVjUYiDdTJ86mAvOm1qDAhP1lALvBAi7QBJXwEEHQ6tbC
m5r00JDA6TX0vLjCzAUtWJuGHHo/iwdWOxpBgchzViadlnLJIolyw8YRWnUxnUo/4xaRi7soHMdY
Q599ZQbRYOdqRDq+F0vKHAQQS9vlMh8ELYc6PCX14qTxOteVXhFKYgTrNq69/bOp/tvmwFizGFgP
e2EYxDtDLDFHayNkfa/KJA0x9GDpZCJRteUvLn+mp6dmHSqHQriac+79KHHnZgi2hktbrXUcO469
ydU5ipzOgE3ZwoVnnJncxQsWc+anZ6qfGSzLaE2+9K1rgEFBFg37HLvMUB2F4FV98TSRpxvP/pCW
20cwp+0JSAx5veY/NOwYMJN42AugqoV1rCJu0Co826A52bZZuqTtcMHzDOtw2P47mab+TOudtItm
TRRwLnTkugg0B0Jxezk3mUtJmvsVkytz8HCDHmrsYrJIsdfoS68vAIGrs7JJne99QqXSYAHaOOL5
SZL6ZDQXlPFLsifYCfLUD+arG/cP7/SkNDNgU3DlGNUkHWXCxgZAXKTiwpxTQNIexVatrRiayg08
BqAoONxeBI/KYrMiGGD9tnQ3GIP+Fy05Abrd7XdVz/GL++ke20SnINyG6HrekiYegJth69Oh62X+
qTzPtFATCHVXN+ivc+EZgEX5xB8Cx2+JC77JM7HgQP4cEUuauN/3iCs0RMo/ngBhASCaC+YWX08j
tpDwMZbDC3LCZpRkgP1CsOFuvD5erBU2ncS3RFu9SU+TZsRvwENMH21YRVPBGJBANMx3UjTtXCq8
ciIVy4SnTrjLY4/mkMQhVpOu2z3uBgaZoKqjUnQ7cCj2wcvo+/+LksosS1+2IRRw35zcOmzv13VH
STQwR+FvJVi4x3s/J0mjM1PZ8kafBF62jEBsSMWCEjA6zpL764WX54i6nfdXA4ntTJuFYvP4ZBRn
lmkAcMw0Kv4Aj0mgIYFn9WlqofF1A4bVgNdsjNEqmgYsQYpnZEUy3nfN5DyUDN8luuQ8v3uduIBU
T4Vz9YHMMq1JnVIZR793LUTyIv1S3LeGWvKCny4v+Q/Ha1NrLDb2dWV4iBTtbF4KD+UAEBjxlq+9
Lv5e2dNmXdmKv8rr970wCDqTIGPGOq/XjUIH1YPqKqc6OyKtOQIs4JSyoFTCFr2Ir1L7rjRBW9ck
UtnMDvWB3zF0zNmiGnVU3+DQ0qeVu6njdx17teeI6fXJ6PYqQbUDyrsRCricPmhxjvE2pBbY1QHm
JMceRkVhAMQemYCcPS3GyjwjmoqYyz0QmpLLW6JrW7DIDn0PyL+7dkpIym5Mlor1drJd4sQQ8TGk
ACAw4yNpghCjXFVtBscEM/OE6PvpNxrwg/nH0/vPOqu4Mrz3KyVRC7e5Wy1zbiCXFA1FPHK4XSWn
kOJkthRcxnrUFxwA2AGq9xNfoapCdsodU3xyFqHogLruxhiJblRV7i5ZnRvhaOeeaA485MkM/iP8
zLCjK6AlJ9VuUoA6KOvvkKT0fpVqHUDUO4ViEKFtScvytxlPi11EhUh5m1/QEtixt9AzdxJkH81U
mBsodpybr/V0mBRVxbTo7nwt1QQZT1D1kD64cak7Fqp/zyfWxwIRvqJGZ433wdp31Q5jyfxwzQC3
tLBflWe52of9mW86Qw/6sl3Ls4Zhm/rDKQiCDntK2aG4o/z9B6qj085cjW5DqWvVBtrMcO+4D2kb
LlcZBvOxTUcoZMmH6f8vxJKia2xvqd+liPAvUXSf/FrMD6Pam5CCyWctNSl0OB8ChNVrLyxw3E/Z
rv21K8rTJVmNCfO7+YfJpGuikZ4ZY10KDKJiMFAr+D58UGj9uWJXjfRA7EpIACe03e5N7LY5stbb
947TZH8bWKED1edaOy6BfAwhuMqFItYtcp8zStTa7AKcNcxf+h6xPHbKbx6KJsglOt7t1QnPDptc
dgn55xk/I8Fihl+2T/89gKUdFHYAJGQHYA3xtyLH6k3+GI5JjhaEMfTe2iDVFiJ6Px7qkFeR3uQ/
YSZQewXH6/wV0dMkXPfB0mENEx4MEDR4K/aMu/4X3NH0BFaIQkc7Y3UodfWj6ID2bFGW5BHAaiMg
/1eAWH3qQglp6tDbLaAt9I2Uj+Iq6Blv9bxP3wFtE+k2sdvAWh/Ps+wv8yiYh+gfKpwF+ofIsGRY
Rx1y9kQfjZl0qiwFIKeJT0NDFh5jK65JW1QLTOWnTphsVHeue4fUBw8nsYiKpR0lG0jX3YXDE5N2
PhaV4udvbZ3GfPBmbDAz9Sx7LQpopfYSboufmEKIx47ZPcrY4GZ4GT3ECStxo56j0HpzPuMm4lGk
gWS8muAGJED88nhuPMi1A8HuCSHrBtCQeyu1eskJe7JEJL1qt0YG+HcM4ZOZmp/PncCJGD9lvKBQ
bFXQv6agMCcuMomqMUQrIM5DSSJMRc5mydzEwIZwznkH7i8CrcoH12OkIJyRfTycErV3D6WyJ0TB
pjasoGeN4R9X56ffcQj2mp4RATq2nEDRHWG1GE32uBe7rCHmGPzwcNJeZHcqu3L5onMp5mQzrzgV
E09SNGZ+3GGOqt8k/7ZIuGBrB3UDMLpNNaOwc6CUVMZUxG40HRtr3AfpknrcaHQ9Ayr1DWX9yW3J
QZdPH+gjGEQ3fmEHBr8hZHMPNs5pWA9rZCEsIsUtjuQQTq21HzGzrQY+ipVVFZd33xMobUwHSFX/
qt/32/sN12r72fqhe+LknkkggjJ6JhZQQfbC3gXDPPJQ/bCvbxo1lg47DJwCWZijD8Y23cDlVH8C
Df6ACsnroTMNpfGOjmdDXkDkkH1168Hs8ZjHbqpGICMskPnnz0aJip/02amrH8hnw4kf0Sx2DV1b
w16quj8vVvglqVrX/pDVIh23pHeZdkWOXGufnbNx/WjMG8J1hgShPocLIrTpFEdjFHaH47PD86t4
yWsr/H/cpoDdJ+rDrqoaQJJ8XYBHu35yD8xO/ZBngN4Elk2mX2Xp79kT/8ozPpIDwxN4yvZLtXYO
B0aShPDiYc7dkuxzTzSSea0+p+04RYBxV4SiHSfaSVdT5VJ5SMvtt7kc5AQDHt8ksxq4iIrTAl3L
c6ZczZJbBGGSMmnXkI1LR4ev3BLfHPwxYQP89MANomdHgNJU/R+1LSRAE5McYd9e0djYKLc8dTR8
NkXH3/ra8LBluhRJ+n0mxAzvxC2TtkCE5MMHoyI6U+pQrroiI6udijTtBb5KiZkCZOS2oDA8obDd
MGg4uuSBVIziahU0k24ZUIfRgzv90nZfwOMn6IO8UZEMWZ+NKHuBje/nxWUU9FoGO3p/Hknh2CJr
tYIp9xMuemtmLUoNEWYozolCztfO2c27Pw7cOYISsNodhzuezSbE7rX6EJawz3HHiK/8LrAIDvj/
GE2vp+5tNySLGbeu/Gz+JJO0kxp3HuPd4K095ZoaGsMnsmvNgCfcnQ5r/Tkp0t71JEs3Bj0qLV13
SK8ElYweb0YsUPgVprBdDNg5NOZupfvbZhemL0l2NwChK5RF7E3y3mY9nb/qWf2HLFT8saZVS6WH
32Ix/26z0f7/ruJsijpGyHfi5xJyyR843jaOJp4AvAoREqLC4gBGCmcs8mkCQC1QLB5WfaoQLo9h
mSTXW6gnFzsmN4aZRNzyPxSK6V5r6NOHVNgqIQlg0muPkuws6qeVEUGVV/gu+7viQziMCdaW7edV
GKgXZQvc7fpajPUeJSn/tBpRoo94ijxeqFkWWV+Loil05is7hqUPrlcs4MstoW2AMZ6vBY4g5Kiq
h8//7fEAc/2jlvQbWl0+HBCR0BW/iW5gpBKB0+m6ZADlnPm6+THNElK9FRbrjYRd2rL+FjWhTn1v
QMEhuBPF6ItAfw7UszWP3pubL4lbzG9f82/KVVHWDTnN+/16jETeLFE6H7X/Iw4jPKbMiD6/ncfQ
N4UxJ+OA2uyVl4Aj7eJ9yEpQPnlvGRBX5m+2g/drUuM8+al15ujcAs0H6Q/skmchXejgGM2xjVnq
9pJG4Q+m0DDHMWGl6XqMkt/ZyI+Nr4i0aKtU5oP3dZRtGwvtfDcO/43L6RczKDQ3AKXMfC4ebV/o
vtI6qTTzsz5exKLNuCkhypnnn8fjNrrdjleQsTjg4b3aPCHzWTt9wVpl+7uMAsQtVRPxVIbKJDXM
n9RzLsp9U7x75HazaZJJleEqSaLiE9yzsO/1MvgBnEZNOZ6+aQBsfCpKF7U0oHM5lTXwzwIFnJUN
ROY7iqkhy6zCCouJ17mrap8HOuLsELYwgMYAINlNRCCMZsLVeyHj0jUtzu3lfunnWecUDMAN72mW
J1nL3TTsbg6BrbPQ2wiG4AbqqoVa2AuqvoVaRn2omfVM49+TiOlnKXzQrxQ7xIY7zHtGo2rNrP4E
XODN+Zsp5K+BaNnbykn/pwduFD/rhl8ryJ3pDfZk7np3BUHk0rcU4I8a+1wBM52bJZv1l7zvv6Q1
mZiXudheUS0SbDIoHaFzR0uHaPWaayJ+L2Ge3ijZl3MpF/bVjqEpgzv+E6uO5lZ8dlnpuDMuiXzi
MntkAhMPyYOJsDHrhFo0rEivauLEr8o63H9fqRaGu9pvGrwpBGM7C4TBmaxzYxHlGoFHEuGQjROG
E+GK4Wos7hfF+dVuFw2SCmwA9eHa2BtHzQ0roJGSGqRpGy7kVe9uUpknH2DTIovjzvgkB1fYJc0Y
b8y/qDRPpLM1nRWQaeEeg1ReEip2ANfvXzlpS/kD6/psgUVLRoKZjYgmuQqmTuZ7xaNw+JsHPVoE
aVmMEzPxJ69NI6JPeeGpeTPaPxncij0/XNpov1zi4/HVPqu1plGLf85A7iUMCLE2cuNoNZHKTsKK
0CimeeaaZOfJyDf+BKYi6IcfQHHlyNKkqEnrk7SnMIB/rRet3nfAJCwRIPshCUcuyHrUEf8eueXN
uvGe7NN9HhzIho+jCldejrfUIqVJcZdI8Bw2H/EU3Zh5m+mjqSjdiyimxxUPIYUI37Fbv4zfHeqf
lfWmTThnrfnCDXP+tYns2B2q+DQSJ77oFcyGtbxWO+BBKwVoRqGz08tLzX2fBx/E3WXKSMD2SWrq
R3ImRgmnh4ALjF/k/pf7Y7W7mls81s8b4U0/Zt5aBfTR7NuqHMrvvmueARzvXmRHDDR8VjUVetV5
PvzuMVPwhaponcSllUmNT1e+XVBWL0bxBgzRzi4Qul+QTs207DaCGd3k+Co7MigyXU1XIkhjxR78
Nye8xRnN6xj4V9dCx+aBeYDOOyvJfN8AWsRgtgIPVy4c4Bqi745+JVCBm5cOHxlighsAiLwTE+hk
Vk4XAUaGS7kf1fGA7p2V0BdarhTsHyThYnn8UbZHlv5PaQeyPBZm/R8wl93PgEiiMYZ5w0+3AiId
UdXpaT1ZvJK2ffivN7Wb1wq+WMaAcnNhHH7u9Z1M7GNMPa9USjMc1TouXm8d2ETYltxUbQ1AFBiT
zB+km9Hp0I6/3S5dXrIg6LENdJ78FSe5xQW611dalJXCBNxtnfN9z5Kcablonp/zAfWBZWQCbl4R
uFH1Da4TkqpWVYJ/7D1GoLIOFRZAV+YzAvnqPWY/CAvklxrt+BOZKCxv3R+rKCIL/V/Ewg0dxSQT
J0J5WXyepF4wYJ1G5DQbgX2MdF7aYhq1cNMHHUfGTGjTUQaG6TKjkcKiDkNytSHmqNZk5/XFRJ9d
N9JAStWQUMSm9Da7GyP/z4b9GSIm+UliD2rlD0Xg65m9OqKfx5Sd2czsxHoAqFsBsNWG9pL8zpHV
qadXDMRHAIzJPCIOoBNik8pNa4h6smztkgw+3FLrUz6vIXARCPkBQyzKTWSm52oSa1Nm4VxsFibV
O9E2jpGZza2CGxjEwL+D5m3nP1VijOzME8X0m3w9mF2SiUgBlER9Faqkof3dcYo95kfrvt3an+3G
EP8hjmpkt4T2pGX6JK+dRdFv9L1U4BJbaNdb1L582m0pGiGk53kc7QunndNjEyViDK2HtoNihCgI
KneWSR9LFYiajwL/KELtHW9JTZfRWLCAKuxDsaiZTFa3CgEJu3ZpAZgyQwsfC/CinufOkRVpNU+C
lyR77JSpFbhmtaPmX7Kdz+C7P/zIYuHaDBemYYeVeBN2hz24/tMe2XHdQ8AhmJ47oNa0I4AElGEt
3mc5NNbSu3hIOabAoeukKMmsnGUtylBwVctIHWrPNaq7j3xfAVuv0eQnUtIpVskbscwRTbc15bWO
ajWohOiOWtoGs+4mRzh1LpiFwiwiEL8OC9y1tkDRm5jMGyQvG26YC6bBCg8E8evLjk1ctK5CBdNw
nHLU9o8SNpuAIdlApXJSfmDTc9yjd/fp67fLwCFusRGAT3c03nMT1z6Cgo62Jr4rMDpxeG0Mg98J
T5Agb8lnKP0kREcjRMn+YOV3/kFSnS3+zTPFnn5ZrJuTb12KooGkaF2yfP5LA3euFz+ZV4tiD3X8
5r5zi5zs0RAq69dASuTe38Ttzakh6PJJt73Wb1vDZaOoEjPAWxDOyVqYJpCfXCFruPaPRFXbvUkw
iUTIsjlTWMzgzshzytiRoKH1TeqOt5ZTIyxsikF7F+9MTkNTPwMXUCIRGWhMn8Hy6K+2ccGMXR8l
edjg+lfqs4msKMoPj75S6kpnjO0Zj8AkLlRzujiwRJu27NLYb7fXJRs+zaE6LRc7FEG9ez7yimIK
Y3/LQMgaJheiDNYheNJKz5WATPOj8pEAW5KC0CjnKBelEw2sPgpMUU7OciImw46i0VQssSm8WNkw
TYqYA9KvXF/z74wVpPYLgCBarnXM33kDlkuUTZI/otz325yl+7dKPK29AjTDxQcAEhdr3Rwp4cnc
sQACbsM/BWr06dAjRGuK+1PKaxSnl7Xy8lq19YSI8eCKVAuzEZalobAh4P60zBsvvaOKak+jfDR3
2oV98Dvs3w6tZTSBJ3M9TS6P9Cv8HtpoBxJlYitbWuGLKOpS+T1lY9zgoRAzHV/9FJH06ejsMiFl
ut1uit+x/e2nmyG92GkFxW8/xrUIWDXk7IaPEGJwIUL1tp/K4PVaKSkse4kgX0PKus72L8l00sQw
efXCXkl3lyV2PP6Fddb5nHw79ru6+KJ10vCQIPms5rIeFAPT4pIFOnzvMmKI8JI/7EWbgM/3n/9d
xVHnjckjVNkSF1qQvTyrCStwdNzNjZLDUFLNfxqDN/VpWnSMhC9/dGT2zTFYupx9tGxJnKpIVYDU
sgXoTcK030nhoDMidHca59lYzM3S6z7AwmkjkzMoegUgBSnY0hRKkWJ131cMmAQJILNerl54DV6w
JRCiiuMHIQ2Il6ycTyTG0FRoYTxblSiTXZoAX9Eo1pYej7OuR4r44hrP2UckhhhGf6rKWvxW7C7X
PNb18ahBZ+J0DCxdPGtVf0cG4SwWX/N8TDdU2qNncdxAAWYLkcKjKybkhwwEoYSk1ujMj3uoJAi1
2xeLav/34L1VT/1MwKGO42BIELvNJnm948caeke7Td50kFrUJuTof/EIkhKD8PyB5w+78f9+n8+z
wwsdWgx6YUAFJ/Sxa0+kSgVUpXYqNXIRM4Fxq3Dp8eojSMGK0yo0uxPnf1HDnqyRCB7F//On263t
OFhFFYN+acn6bDNHcodaiWUUBUuJg470DhJ4va+XNUtNkd21ElJoZDNVR42wYb8oLNpN6HlvASJv
piV6lPVE6Ge29UsBhU7FHyE3WCO266Zgwuyxj9Fiqa+8zbFCLtmPzXYySuILOFGgxwr8VUEga6su
TE3Hu4unUguBLhhx+2bgTbNC9WYagGz93AianM9G0SEDGfdrWi/3I+RQE708gnHOBLT0ZJL48xL+
pnHQ4Um+XRU7dQ3xIg329+cwfNzhkcdQp+oSKmZurYBw/rdcB1TIQXenk3X4yOK2Rvezd+U7n+nE
Vrnyuugz/ukqlEDoTrfnqgg1Yv2BAn4odxyat0MUaUcv2eLHBOTvB42Cd3deTPxsPWLDuMkXhe8b
sx08nnAUo6ofu9rjlxLc3kcl2TSltyBDNOQOHGH094NlElwHFNZQsoRg6PT+Tm2DH9taKfI/eBFL
W6oDmFcPrFCuFbhJl9/e3uREGebagFfSpPJYwRhJuHvQ5KTYtrZ5Ek78wFoYyDRzzHr0xoAOmR43
JDSLK75qyYB83zlnPlJ0mEfICKcw/z+3ZFZcCxLwSQ1qqZWkX9j8blG/mVS7+3zUeqdYs/OeGRCu
qMjHn/LFEEkO2t/9FYCGJSD778LbOCYYdBtxNYQfDuUT34MzF0J8d2rzX3LYfMplmRpv0zl9E/fY
Qdpwq0gwKr3JOZgnKL1hc7VjejCw1CB0eefULkF30/PikXl21NxMPT7qhb/1CnpQTzUlGJFUAUjj
WKqS0ds2m/3LzsiF4wDEMowsuB0mFZBQVL9whRNe8IBHfq34DX3bf48FzdDaHTpOu+YxLsadi2eW
CyIsaYTS/GryHKix8udVnHVANqEUqa6VYY2iDpBcBIaYVxwesPfuS05Sh9wObpQCviUie9+DVyVZ
ivsWIe6T0JT0TEiDPrM3xBuvvK+S8pgyFaPwRymnyzpnLG2r/jXL9GJs+EY3xkQxbR0UrV+ryUWU
KU4dX66c+5DnIEVgFKoByLDm+lUIFkvUE2z9BAnSuaIfKG8Os9Rly50AQgX9cxgR9Pq2dNAUOmzH
DIv7XtrYjdszRHsB08N7EBXv/BsxGSsvk/0CVLxgkDva8PnyW9bhulIyhKGwPHM/nBLaEV+pzyNt
fwapqiaVdEvL/ftgxNFDByy/V6DB056EqQ6ABTDhTfkCGIh6NbnB6U86HdZnOiO3El9qhng/dkbk
qv5gYQECLKeJjSKVrOlRNDEQvNG7yejyPAEGcpnzOB6m1aDPvPokeQswcn6SVXTi2B1okAkm8gxf
9n5VbkZqS20lRf/AxAzmoleWjVAKNlqWPHCqro5PXiCPGoDj+lGX+36tRuFXhvN62WD+ru+k6A/X
hOEMiaM3+rQJIAYrL0f+JBlrtgNoc6IcBLxtxT3IvOSZTarWT8wPXHRAyFNlo6CKnW9F5SFWjsbh
oPXiDK2lAh4MnR++Rk7IXv8NP/6THzXlaEZ7D/wI4MJd09fHfbZkIs4lOfOPU2P3xAtWHXncEsKC
yGUWVCx6d0LLYyt4KxPajqAm/lTCnZo09zytLXtjt8gGZLnKlZXuO5lYph8/nPewwh0oKyywANZZ
ZwI1yT4NA575Rh8Zzm/GER1nrbj3IBQm3EFN62ZK5Hz5KBEhEERDT7/2yu6kdRkM5rL81GaVS7AE
KIZTtxxeembJ+eYGuC5KdSh9FncQxRcnhpPvWI5OrW/raEk5fIxHohM/RPNfFGWIIJQOsLHhhh57
EVJMsQcAEPDXsOIWUWtU4sfXhx6pD0aqV9o13JcahJwjhx5rGD3tconfwwUGVwP3hVax1K4wgV58
jnxK5jZt8xQtAmuRv8HQATbvJjcCELqFZWXSTM5PPDpQ33ENpGE4MCDGySi/PTw7eqARstjR/N9M
tTId3Vc+V3hVdYC86p3mcoDFc/rbIeQ9NvJq8UfxJlPlIckUPTgjpe4+nlacW60p/fcIM9SJHM/t
EN3bT6AN2aNf4HzuIoVY5tZM+pzyjrMMFyARP0SjhNSY9noZdzWn9p4G8fr7sNaci0XYqL8s6OMo
xBOB00Ms6prRgg6qBzlZrXbdiGLPsUsF4oZNdhDnpupIfcmQ8hhov/q/H9eNx7zr42F2nS8Eoedo
cUlBuAIHWAAdnN6vXoQcV6j79MqThmL7mXEfD2bXdqex0TmKYAARXPCdBLbmw9K9Ib5uqxgdw7U3
jOkoozR9fJARuCmBmJXfC7AWA/5rHQnf8/AniOL13QenqwyZ6oY2t89aJcV+ZT1CXlrbnSLMdQf8
+unYEnukrG0Pkf54VFGLo6Z+cV9IyxCJN1HtnrPWw89xevn0lMtSVsWL36ExXF/NCNdDLk9jOxPJ
pDb3a1reigSk/aksvw7hpIrLfQueMe2D5L5g5u7UJfnIH9fgIJWLApd1SaM5yg6rilhW1Ql4HWsJ
S2tBCFVSD8wN8fQBGiwyscc1/4Dh77UXB1ZV+4wLuTXxEZl3zsH8/qmzWQju3dvehuY7foRpK3gF
LS+WKRC2TuAks5oSVSkCXwmR64h+drPLbYuqji9srYANc7ZYAeN0PISa1j9Y1YQMdhee3Nd6MhIk
82BNuM31B34tzub4yQvVBy7c2Y5G0TMfCXaRe6+KsyIUFSJZOqaTkP/SnXcbkQjlefcxtHg2n3pU
f4jLr46KXrnazj6YRYMkMiHcKb3kwaSoV4vO4vL8WcrkzKKhZY5BVOGRrzKfx03M5XoyUqbekb90
EeoaZ3T316DeCFOMf+OrqEpk6pawE1CKgVb4a8uvV7uGJZOkVf9oCoCPOVA2vCJhAiDPBGRR77YQ
RIU1mHl0S1SK/RaHSlJqfsk9wn7yczaQPHhFFGYP/1YeSvTak3SviQZBxsmBNYhT+BMT7j4e5j+7
q1RxEvNAq+I5UVWeTr5YYlNIOVdAnc7JkitMha5FsN3Fj1bK6/91N7/t4F4tl48GKaV+UD/tASec
M/2RoZVs8UgubLhX7CBJNfVJDNOQCwmiTdnJKewCcwIbc7xMkkcLMM1cZC/LbCwKqP/zCym1Q3U4
fpN/ZATMlgE0DveW3usVhb8lLD+RSo1U0OR2UUVDZW/bqXoLNUwd107rjVlGQ9pt0NgBktDlBDrW
yCuhs6IA2fCnuyvkmXzeXU2AmHHW7xYkvmf+dWrby650OZ4VhJDN2GqW418e7L/nVZ40H+qDxhdd
70asgWZmYo3dstvHLvwp1XBrmbPmo8WaCLkWd36iNaT+3R7xTEqTPdYYmmzZFjEe8R7OzxMAqrM9
hPtp1rjHX7QrwBbRxBsZKHaJiL1afJti3bF7sI4VQjThXo0dp+ys50K9+f4S44OKp81TuL8xR/wR
45I9iCi2sUKRSeFMCCl2TBDSKkDZYWDTBtThseT3zxFae2v2oaiNSmzJRrpEBmrHw+jT1ghxwS2t
sKqufohKo1hILyuTWyssXah6PLTwlf9VbZU1G/MQ63YRdlnbqD8i/Qq3iHNxXb683PYWRXXflQj/
M23JC4C2mQbmhi3HLCCWs8byw9V3g8LEiddQMU2v0Vian3M7oQ5R3cSL0UPChquZbcRqicm+Ou9T
CujKyWX+PkphccNnZ8OxDAHx/wKHLLLLBuVQxDx3By6TgyuiAyLFg41mRxfXRDjS6bM/B/M6JqMq
WUuTayJWBzqf5QTCNZ+msV4kNBZjSClE1ofH9Kl76AEKqRUSsRyR09MycAKo+jMRkbcwnB23STMm
eHzdT/uBolyd0pcK1PlmC6pGAhNMEZn7aR31v9zlowNnkOfGHDsIXzEbJ2Jx9iq7LZ/HU1FCcixs
zRwE87Ai0LVBeAb3pveHbGU/kOoFSWra5iov97oRkmHKOm1VMV6gEk05NDjJR4ggieM+DBOIwnAB
QU0+HdTdTym2Bq997Mc1NhqNEPjTVCBqkZQhLWH/w07F7EcRHK1c8fsmHSp5ocJsyjZ6A1Z2EY20
pc/Vvvsah6da9UEpVmfPFIwMoBBijj7Fn2AFzB+KH8bLqZimJoDdGjB7GaiVbbyySfZD8AmA5ZO7
bAGlHOYZwM3dEfrUYZfvn+aCEeS1asEzZkb0hwHCmWmNUFNm/IEhFGwm7eJubpettyfhMK4xyZIl
504nSMTK+E+i0aIfiT0/KE4/m3WJQOZUq100ZHjo+7XOLfA0aIL/UC9fWAPA+R0hhejQnz2vwkGd
nlFeTWGRjKpzRDDyNnsQxJQH9oQ6hbVCmIVqU3hktpcJ0GIlUXCLIVSGSjonxLs2jG/eG0YeJgvG
EeSZi1e2p5OLR7FbmjFTsxYK50R12/sUzSpUMWEx4USqNu7xvOqWATq9s3nFLQomrSyUFnEawLvE
o9kzuIaIqtNmgOd/Gp23PPASYSm2+dZhIXFe0dRp81M0AaP3FIUGpgHaZyeS9fR3FD5/7yo1fLrl
b44pVnmgFaiiFMzxU99XXWra6jYi68GD3KD+SoJTv1dV/07NlnumyMBfg8X6OFc8IfP11BQLj/mZ
ZWF5IauvjM7BJWtcFFDD8aquOuvG8Pnou8vHL5wRVBjcv0fVbG+SzWKliyovzkNEVOybWgaPNHoz
TMba3trwXe8HNYeNgXWWzHsG9iSaNXh3lJhlpzWRAHw2PXtp3VXOD/RmZV0z51KA8XdLkTYGy/iT
KxNA497ohWei98GlUqfx0wR/+DyyN4++Dc9wfgK0bnoBJaDFqWLIHQSR6skTzoK956AEQRK10303
QYk6j5ju+OixQyVIABKCfPppkQ9ciwHAsbKaOO/izib4pheKZjgACDPO/ZSZsdDqfYSSAezgK0hx
j8to8n3s5LIUDhCuzoCpMnFyDUAMYtHW1K7T9RUmLx/k7AR6ymgrauVUnPpEAnCZnjHUOJ+zhYOh
aNsS6SyCfZZrQ2yCkCteGm/LAetIVThRfj88cXSxhBugzQJdL9fYWQg5WeeIpQC226Ug+eL67eHE
klXvdrJpDJMoPwBByoc9kik8tg10VgplctfPdtSiR5SSj64HR1Hc69r/v7vXtfsdhzbxtk2/LoAu
UqJNmtOZcO+LDztIXAxNegnwzeMDueJg+C6kVqlhM21hI8bOXOuNzyoevwc8dP/lt+L015CKagIP
JtnaKmI1P4upugh3mLUcN0rlmkslURP2r9+o7J728UZlDiJmwobyXZ31iigEKECQ6lPGr4m82HIS
DDtu95PPZdvKR96Ie/a8PspY+ebdX3dRwYLWCpnUg+4o4dn/tM3ctDCzb681B/ynCpJGud++4AOA
0POcMCjzzy2dJNZ255aF8xHGG3tKHejRhXHrjugEVBrYQDUQxzPXfF+yF9Mv8Gy0P0+cXvcG5H1c
wVTriTiPt0ZafPpYC1PzJF13vvEbK17vqILLAZJUqoTjAS1A3t+6ncQ2HrAaddmrth8kiIV9GBdE
DPV3AnAhtqFbHarCt1woUu6g5xzArHjXrGxgrvo4F5Fr3s5ZQ/x8jFOihCiYY3kPVqUIcT1br3zU
uwTOb9f4plaGDLzhF4qmPAaVJ6oV2VbIounD/qfdMLXPs989pndGe8RrZ1Mcc8GDqpuY4jeh2gr/
KMODN0gfiJZeQboLwDz7m7l3djmJ7zKUnZRyibViXj/HBxxCB2nxlTuqwbVZsvHRAD4aP/JGMRdr
W+cBXn72fJtV5+nx08VLM6qNsN35hkln08SfiOd1eqJVoX7GdV9+ZXfPiNRw9aouvQlTSru29Kwg
XCnwcX8hKRiOCZM1Lrte2NzJjDIwDQ2QjNGa1Y/q826qUAqsiHNFRF2R8czowEezloQOSoKrmTjr
DkYnPFqQcn67+SQb2GC/jgfsuU5FPjSLdxW+i6uMYxuheIbwJl70NqU3SpTGIo5XdrbqqEkKU2TS
pr87xE+OzLxrIoeRaTTnpX8CTjwLHDQyGJ2F1J67y8MpUxV6PokmLfVOsa59q8JAUR40BZtSVWKi
axRmxDD5RDVgFUQdJgjz26Y3whhRcwh7SaKGW3I/4cTnAwgdh+TXoqaP7yKE9TyY3CUGgHlpnbAb
b26mFl9WTmeWXFTKCFxAwkDlWVx1/qG8S4ft9A5Buj8f84hrgBregc2hoQ2VhMvgOlMRqnHivm+i
D7rQPC9C0qR+MHxZSKxXdGeo7RbsHuWU5lRtwwzhc2a4e2VfPs20mFCyCDi/y9Ts+se6xtMTR7bf
7LMSG3emczyXDJN1e3sJFkVMcztD7ycrg4iyXSd+Bj4FTRJwbxtfrFA9j//VovTCKltBYxIMH5xM
ZtNqwZY38WLB/6xS+b6t7siN1M0AL7tD4QDwKWOs737fs5bh7sRwFhwCpWOAhLh5wk6ia9vyC2xa
jtPbJEQVvRApu1KfzX/nFI9zOA9fxdMLDZO79wpcZwqE4ygB17lzh/K6ynvl/7O4jyYEP0ld4wzn
15W547EI3mLpQBaLZYrVR+unFbmf9YtQ1jw51MeihObiKvah8mnqrLdhu+Os/yrv3nBZ9RFlUSTD
00S9zktJJyHCmDH8u7YrGrctdpSA8ZnK+n2UYtgHfCOvg3ehjmOwoiRAr+6DwelGbEuuP6SDMriL
a3T8AvPer44H9BaW9s2fuJyuCJu9lBKMpL1ExZ0sM2HSlmFrCKy1w48AF66ZowlnbZfqJ3+Q+hh5
1LAA655EPhIFI56mquCgAriDDBsmdmnUugD7iY9PYEJThm8xO+lWew+2qvKIzA6H5JNdMtQwgNJj
lsiOn6Am8xdDo9+GvhSEliaV/xvy/y3KuEjlD9oCgg7xk51r9FnJ+jWPfXwDdFPqxeqB8LrxpRdP
m1hD8b6TmxqAyOdqmw0Qkxr3TujUEvntaPGosrFykz1ZPQkv6oIEWFQrI8IcLAQbtLRfXxrSTbg4
YCEJU8YPYrYUl/QEtV6MCTgGC8SUP2bFD7lEuH5Rr8uIJ0eAXPQ7ccXWxR4bZwWvQn3sf+v/e2uN
VHIdQQH99JJ5wRtu83AVSt1B8jzQuEjrBw/Yn+l4jLSIwimWgC82XkTlRk+4ZY7W+7ovuJYHGAyy
F6fwD/yT6oqdzmcpo5clvoAYGeVuj35QDHeLDLRRmZSxvgDee2Hjp6GxzJDhn/n2PL0z4zBZex3m
nIwW16UwExrQNmIuUjzPZHDIrGgBbgCX7OqAdZzWfDh+aFQmb1rG/zFYyPcfBJX8VMIeQxO3IZXt
JOfIe+gIkjqggWh4vB6U9f+gLWH6/YcxeBTTyUeXY2aMD3BV00TXO0+5dTVMS+tV5G9AGPFyoHq/
q9U51n2SXR6GiPPpXP1rtwl1Q1XFlYOpjQ8ALEnsL1mGAIozUvpxvDvg9Zip7YZAibprb0T1Ksi3
fm8n89b2P0huXYi+KFDJQNW3tjuCRrwTM0GMNDEtWg+faYR4VSeMf3mcded9ClAz5GDw711kvKRq
yhF/xsv2BRyRk/f7porxZtkJRaYVcBxW9IMHemxCQ7i2yLb/6dJB+QO+7nk87RsSD3rK6zrcjdRX
dkmfkgVrJo/gGcX8d0K87AHqU0LFsY4SIlLKDv96cp/1tAtnAi1Caa7T5dWm0sIl7nZO1xPu/trY
KLDFbWtAoD7+5xX04NgGCVKqYD23T+G124Q9pe8TTN3m33M32lEwnppf8A0Qm1+W184W3H14W/Wd
p+1Clgq4K5OxQAiWkA9pOGGKPix3/fNg4Rnr/R72VfDqVn5OY0WlGc8ss1KE/52FEUU+P7nwXhdl
06OyNcdQMyUkHh2gXJiMvL3psVz7vV94Fg6rnGy6F70yftDHnvDNFseLx1ssHbfqG8ZpQ57yqk7F
EHxcnSCIb31s4Fj/JhvKZecznjBlMZCqtm1vKLhnwWl8MGDDGmcC/GDRtXd/sJD3MMvmXCdhHUZ5
AS8/glyIr+0ZhYNgEYO4K4rsMbE4RFvrGVBAcCwsBJgOHPR7RMIxShBM4WTU7w3rpTKNcXK5vL0q
VwgamXE3lUBRewhqq2EKEOC8hO4nEFPEpZ2bRwemMkUIc7LN2kaXhcRnxi6+vQZb9xFfJ72zLRdW
cgmrZA+r/JwVvRcLqqsVoWXntiIiQ6crfCX9NR0kzbsm456PRl13z65udvExuYJRemMb32pWHnvc
6waoGjfIPJYvcX1XcA79L0NekDCOoI1KYFuA+YjvyAk9l1ZHSYNXAnbSNH1gzodD7ud1Rzdc9F1w
1XbIZMVSSg3IGUtVcWx+jEQGtguWQ8jO25r4tHV+U2pcJBmEWxPdFinh1ftS+ZYPH585j4aY/wV3
xDxOxe/OChp2bnSyZ5T/T5i7kIIoKRQNPgNU0z3otorljRYnW/VRuAp+W+QzeOkb1sQoRIgSmgZU
JdWGzyGFv8GEDVQ8XVgRZKoG1HiRco9aKG3QMUeIN+Kko09/ADjHfM+5OIrSTlyjz2jN7c+NVuPu
UnWQiro3Ea9Kw734MS11oeuAENY4zdTZhDYGsFxFkqR5my2xB8BKM7YgC3NqoalDXySLI9gYmcSI
nmlxH0W6shTCoCm4YMn91Ec5sUwk1ERZLTHS4x/heMTfcsZmGTS/2NzuelEhMSdxHRVl7cOAwDr6
bwcpcoLTvjvuZLuOWZbxymHrQLxvyA/OUd1OfIxB+XurB2Yzc1qiis7sz3MF3raAfm+16XMxGwT2
V44dmFtS5R+1JBVoAkKEtootuY67SRu6l6IwA56Fa+nn86HVpBXyYU5gvDtt9gT5zWwlxrBXwC1W
pWQJl/rX1m4OkSYrPRp2P04YuwRBvcu3lKo/Awd4DejH+1mS4MiA4Y257fF3mwUb822X19h8mvbP
gQjyJVqlAqym0cjOsdwDbm4hIKlPIBmBR9Q36WBdGPwkF585PgyUfBWxegmdIizYtRLevc3PBj2A
Euboh6y0mZTkYj6vlt+MengbjZL1IiyuxVWWrCLUKVrR8ZBUOHpJza8RaC78ncXu77Ev2Ehua930
H0j/j8SU76JRs3pZq3RVNb0fAGCNEVlCkhvP1kEbJZGtWampSb9LH/xeh5S3yY6eHff3G+omK/GP
1BogKc2Glwp8g5Tno/vgk5M9v7cuZHrs1qF2Z4oozKl/p2gZc/nT5hGVO8NyxBvQyYGkiCQsvy62
e1cV2TcTv7N3r5pFBowHIXF70wTTMaYyZjLHIS3HpCw4p4MjcW+4AFqErGlO76cCKNJjJMZ8r7ta
KxXK9aP2bcdpsqku6qqV4356rB42/a6msZjoizmnCDOT406CqMPsfmZx/2fBpz2/IVqt7kHV6zK/
VKZUPKbbplYtn3Wa/ESIDkmPPj4yIRD5gdBYvjbe8uA2dh1FTQeiDLHVABuhJ4iuRWWqVIraas8D
RbhK7lNw1rhJAXotUGmXRxfv63o+7V4tZ6dlv2ukBMsE6mvX89hlZsA8X6TxvngIm3XCHiSi7Ln9
1hzQDp05otK+sc78WkhsLed7BAn1hT45SJmG8LAn3WpLXMWCdiM1JJbs+quHBAF8rVmauv1Dscdo
UwB4Ms5BCV7kX6rss7oLWnyuvMIOnky1UcrsEVTpoNcnRx1ghAYntFPdPhQjiInXk+pYpRTggovw
VeIzD6LSWvuVGIS3e1TBOsWK6h3qyIJaStndKmYEWGIbPRCU85pvEjk69o47SfD8VphPdh1qadbF
9ErsrihOf7Q2iMkgz1tIpTHAg8TQJ+ep0rDHHw4HKRzN/Y0TxW7WFxV3cq+jRRnlFQaFZ8rdBeRQ
YTf9jvcIk6DvdIUpjonlncIpSWBYGRm0v+13iZ233zc9WhN1dWBfel65M0APpmOUobjKEPATjsJk
dH3UQYZaIKDwWHPcpQkZTZr8KWKI390/NdqLwN6ckNf6kMR7RUCi79AXhKXiAMQh4IPzla39wZJM
ppUzYhzfITOEAg1HeMpZq+ByeOrOSlLMyw/wNHT9LEbQiPH+Dj8yPz/NozK2Lp5O1f7HHhwoM1TD
VxhhTgWmouG9pMZUXHzx2SErbzfdChBGgAumwn1UZ56WSclqVrsNdhrVjuFhdGzu+Q/hgo1JOxeK
zrpwmBemUEX8T4jWEE5dE4D9wcErIfWvPiS9M2GYUA/aNl9sVkFWoBjbHkLSuhwMwmqjuEOuybeP
oxdAKxpRRdAmboRAff3z87drXq+zKW41B8uQU7JBZvqHuwlmtz2GdzPbx3VQ4LeU/i9//1owMHif
INXep6iinNyIr1Cm70RJXFff7vNiBhRBmmUplQb+LMxHEPHUgPpwtxtc3Wu4H3R/bqPjfRgkEgpA
7vYGjkUigtmig+aB2P2zuU9+7vEOwx8cGycxoUEVnnA0IRbzN+cPLZw2GgxCbuKvspNbOxniDwBt
Y8RvwFYQI55Tva6aVtpe5PxsSsupMboxpWuIZEA8HPFqaZTHY4U9gBIKOlC0KtEm2i5xfYcP4+6a
r1Q7THufz2s/rjWLni6J1luE9w6kyu/t2XkmgvH4yZViTJT1tYOVcDEwdYiDUe402Ek/ZZRrj/re
xuKngKK9262Y8sAG9Ihj3XaYwWpS/wVyVXjwySMed1+JF2FkgUxXy1+a8GsQeSUWheegB3oYgnl9
qAUGgx1iUqVEqv2nf24Jng0C2br8YIeBdIHo66AOOy8nbBYtr7O3nI10otAvx6ouCG6xKNPD6wX2
XVgViy4Fvc/wpB4qZTRYCoWovBbK4Ah23usLXJB4g3rCBkcXqSeuIdNkozmSz1g9CM2v9XqgaLqs
vl6m7Oj83acvPHquMK5+IGVhKiUv22ToZ0U2AZlXMD+p6j7iiitR8R/t8XBlJKStewNS7AWDAF8o
W2viwCl5LBPgWQ9i6xgOKYOtUvMda+L8QdEBI6owVi6wAJ9mhfAu8y6NANBKQjp/H0hgI3YCYnjy
HQPwyeYAAGAEtO+y48GIvpHf+2eWYvjAU1p0TrYky+5v5IcWndDMM1nJsAnYnHDphhSjW64Y4Trr
SwANl1Gmmm1WKE4RkLjSGX3BBrXRC7mpk0YwtYwLgROSKC0YoUt+Jn9hbgzZYiA+VMQHX541ix3Y
rn+AABfUYaYvyrv2HIu9tYGpu3IaDDSr6AI2p+xVr5cj6ZNbw3hz3j1vlWT09+kDHomLZL7C4yiT
KJad4p93c9Bb4NUbBFW6YVA8kUdJARK/CHuOygMEA1TKzfDYqALK2AcU0D6M+c2g5NYC9vFg1/qa
5ptqlZuccSc2nMXj2XiyasBhMsLwbKmKKU5WrUJaQWQ0mmhStrtZhqlzuQya8vSHoTZEcvYoG2iq
gmOKeRDA11XGS3EnvjDm34b1uyKqROEn1Fqr6a6SViI0WElfKB0XwWSnFpcJ/ws4ICU8ljrY0TW4
q6+T5FU27FSIBFupSd0ktVTrYZCbO/T6EnakxiG1yGMxactBvWYxVGAkKQ1F8GFbKdeQ2GuwrgMQ
LZgPMghs8ZtVP1M9+r4iD+lgem0xAF6+d8M0lQ93FaVAlB8X7POIU4oZ6OaZHsUwNKez6DZ22NSg
1v5q8HzZ9PlNrVwTYltwenpJIFwKKod/VelviTxys5Vb7jPs8XNNFBG0nFaz75RDpkUQgOrvORov
oDnf6rZ7/tSAgMOTWb1Z0kseW6b//5ks7fwDxv3HiM6iBIh75TZj281kCLCyldXcZ5dQYJMp52lE
9QrB+C2hc4va+c7tRofCX81CYA4iMf+rpQIYrGbGpeM3HBagKg396v3hnehwWd6uAtNTfyn0kRZ3
3YQson3Esz9Om2uvfoj9/Fg8AU0340SYuaP4uS7PkYZ19yWBAYIMVyOZl8b/5rcyvg4NneKWvp4p
m2zAgVoDTn04amyABpTm0vbDaeazAh+3GidLzaAwGXItoi+cctWqEa2H0ppphp5jUt0KSDKOQxAK
UDtjLikFm4Z/GMlN9A+gLLFJZAlUNAykyzhHpYgUIU1VYdMEk2Jzg1MXFohXsUHVZVl3a2jOMfi6
RwIba07oXCCRNuxUvcaAj0qQ19HEUkjSgo3fKlpVs5yMpSafDxF807BkJsuorcG+ruN9MEQuhrnh
F+MdFSJoWUzrEK9hZPqxMnxeZfPCkzgLJpqyUosPlRedh0y9ommfzYyRxGBao8t8+6l8mRWTYyPL
5BWlzMuRRP+lqz37xfi0BT1UXT1i+7MoifAXPUl7VJfnhOLw0O84T9/faQV07y8Oi1WFJ/yJIgrd
eUMmAyrL/sSUtW4M4MrjCZ7IP9CzqPoc+jiQAsTxy6i2cmLKMtqYP+nKfz4g4Kna1l0nk9c1WjS4
dPLK4q4lIiJXk356qXg7OQB3VYSr2aB9tXgR3z47zVxA/3vzvjBgMeqjXuoUssf1BXB9Onwc/9Uu
8n38OHv3IydnnvbFDMmNUhIo1ej+EbjhrdyWfeo/tr+gOVtpb7WRyCaovYrCNPWo3GImGYvppIDO
jeg707OqfsmiFXBWSmrjQ8Co16xS8ge0Te+3j8KulzwEXzO2SeOl1u4fnSnZg278YMEJFh43mm3U
yhr8w2kymog0VZ52c46MHEXwTCszLmDJdshIMBx0M2ZUJs+5RTxJmeyTc3voOjoB2SBb6I0+EHr1
ShbcTvfJfNNZCztEeo8qSrZXHrMsM+UZIsjGrBWlvjuCws/pYsm6wTS9cicS88HyPNIj2z4HQujZ
UspLLYQ4fnNSv17yOhCZdFVZ6wpoxFY1WK0iUbO/ACBmz5jy4Mxai6u6bIbuaZFI5EnCLqQ/WSew
8r+ik+3j+GZgnUs+ZdOZ2FG8JprrLTxT2M9xpY4+LSlD9lRcx86RgPdoSIc0rpYW0RXGn4hyZo0x
5kHHo7Gby3EywLpbKTd12e/aKitxLbQaV7lsnhWrAkZZgc3e8rV+9dOB3gFXsxSDIAEM+22doVGY
Ea3ikqIWcxB6eLQVOE3OeN4VRwjRUCCQIlVFbrM5cWsBAM1DXu51ZnPHMmAxFP66UM/uQ6XW783x
ox7SOuG4P223MO9+oTmTtTJKut+9KDqR4vOteE7qNEwFJf/6d3/rO5SdNSLXnjVPQwniMdsGTzP5
hkfk7m08UhO2wUEYbpXJ/l1bofbr5A1jhmauba6OCmZF4JAg4hlElLy9z3a0TGaDxr9Ef3GXmU96
GZPVW71Fv8Y8C2MtMjAHWEThStnG33sULNb0r0erb3+FvC3BLVGQNFR7GWgHXlDngCyEHQajErBk
B8KZAsQNUUctm3L8V5PBB8ag2kahKT0FjlIJ4P4Be3egMMKYS9r5LOHwEg676xGYeD/8Caw31+11
Flc2pu1MqFqJfCa3nMLDRgEc/FtiKDNCCND5QHtnG/63zUmG0yZexxm48GVKR5cJFc/IMRON/cXO
fa2sA5+1Tb1H8hqvOQ+dG36hvZ+PhfRpjFrmI+4j1bGuFwlwEUgPdix2V5/Zel4GgDwn5RboD65t
DruzKXOvBTaVCxpd6Ce2GAZ3ImpPVz+uQtC4VYUddY2Lg7pSmXFDMltWGMpLblyX7vwvnKUeCrRx
b5is8v9ZN3l0EsHg628/Qaop1YNuGcAHDIgdZfaONrSWAVNn8G8j/bUuhIgUo1TYMs5OktLFn/UT
XwmDD9TN38kZ3q0U5OiY4l0dSRrI+ldxmWhQ4GKDGMFjyXQnRtbzNtjwZG7pF+jdKFPxxj1myqsU
nQNt078z/ZC4HXk62xE8QeEmZoeMmHqFmFTDqx/GDHDrD4cTOuPBtosf3JHGXKUDbhvCZFLtLgM2
Efw3ab+aKMv/NzjzwOZnjouUNtFPlEMx/uP69xlJAoHnVhWP8apJKG+HTXJTGka51Jla/FE6OXFe
CIpVqM9hOMmWSHVurrvOL5ZvsLsq6gGl7Jiw3XcU89RWhIJBT8kWFU+7IT1dFnR4vwGaE5UIqag9
2ynAKtQgRvmVmfJo1442jmIIIIi3G/XQzTJkbJz7/4ZZTkO/SnpLzXAn0lABxh0qbFW6blY8go/l
ZkTrIIpcYZvaNC2d0ZgKntvbtWoGHAfswfeLRzgzKukykl/qyCTUIPiPLX7SzOaj4w/pbhRH8oFT
OWhuEfT3A7Zt0GMZ/AcaW3aTUrd0FMl1OXod1IBHUbpJf5BCFtkYqSTi/TfWYU5tkyTzo6nSRfob
aSl2lBVeAiN+kGEIws1rz6/RnGvnAO2YefvsXTWYshQVn43BYmchZspdyLsZXv/9rT/wbGQf94ke
Ye+NBnW7tbhMDvB4fNsEhkFHT1CL4nGtLm4D3kEfuLgCWrOaEwbdCa2vr/8uvLfi8kmqRerpyAiU
FCmXv8lNF/sOwXBaniqeTsow2FdS2fdpunnlQuDuYCKqrEmII/hnX2v40bFpDOAvT7IzMm5/omgD
7gy/Hudj3Fhmu2xrp04ACfSsPQDdyPJO/4pXsqn4O5vPaEjIBr+v1W9qgNH7wokDbNRuvXtwvPvr
JeLG8lEs0mpnlR/L6v3NzoeelNAfMjzFHxl2X99YvMcf1WrL23WQTN8nnwOr+Ih3aozmZjIVkUlK
vB6I6u35Xqt1iee5oWEp3RGN86C2syQRO1peRMGT1gGOlRF2nAzLyCkWgJq/hNEv+u65t9w87Cud
TGlQtxBTYJv32aD8i3jpUv0nkOt8CU5zp0U8zjcm5sZlftRD4q2Q90EYb+G9RzMpqXK6lBCbYKDT
QksKfKHx6MooRNXVpcpIrzfpsI2bNPRRDF3HZNpRFkRGUxzFLWicumUdF0CczA2tOBYfrmY7bZ52
9WTIzmHXkgROyrPfr/UkTs0w70P5MAcejYR3JokPAouSg7j1vyZoPeaeLOwoiYZDgsKj8Fsit1Jq
w7ZpIqsa5mj025+jxQTH1Ko+4Z8MJOuoFb/0kdVLp6wkQ5jqbeXHp/xnzyJPKLT490PThnqO8A6J
GtVSEIbq3iNkhrgPohcefevksdRD6m/eo6doUIquZ22rfa2ivJipdPy/rgCg2oJ9UdaY94WX9yXc
uIdPpCmKePDdIlqKCZM756MHSXYAB7actgHkzNKW1ByRG+POCf195VBsQJvOA83W9FnpfLXtgKKX
+YpS9ud93JYVUKNPkrLt3pBcTesvf4x/oCEi2hItP3m7n22aNHW59Y+FrQ6D6cxnvHLwcYCTAwk0
mgzpcwREqAKdlz1KKOxW/XqJWkqeog4GN3Xc8V+JvoJCswX9UKHujHjixLHsjV/4FkHv7DpfpC15
GC3iKbxRC0RUmJ/E01Codz+Ugents4kiZip5wQDHQn4NIjmffuTBMJWQsBMkRgNe2c0dp+s9ofFK
ZM7ji5KQDBzlqN1wRoNzih/QmC/tkzqTbvl4s8hoZdporsT8kQN4t0xTpaiIW0gH89qMT1okdBIK
GNx4Ae9zdjFAFGY+Sfim7WXjUcUG361rX6YBQtnu+qK7sPJI6MHCY0wUWjwVZe6DPN71VnQW2fls
rbXQS1UTP5KzZiUlUqcjCCtJlIFx8VPa/REDm4V2+XP6BTc6wydfS9OX0riGeleGAHHcrCzAAUW0
4OTDuGcI09ZwfYQ6IZ+pXdCcvKYK2MeEwPCjCjJG9w9/GubCbRT91+hKbTFFEADbkaQ0IYsj4h9T
c+BoV7TGrvb+jsmalgMNYj6lYKqpAIbznLlpieYRza42EGDPmxuiUpGnW01x9SCsPoEpL137QvHl
Q5eY7E4TtCGDzVM27MDBANHkz1jyoGnR81k2Qp5Z3p6cSSwgfeH7VmxYsrtX77u8Coz7NTlVihOY
rBDKeKiTsjujRncKBYr6iUKolzjW0a4JGLRixF5xzIxapSr02xOqoqG76q1cKMqtUJDZftt920wi
S2t0U9v+u3YVYHDoczHGyA7yS+jhfYaMPsrrAxeLrnVVFDVZ3KofAmbg+iJyPUB0kmXSpgKiAuTv
Ml3YsRnLXV5i/DHBekIcLMpqE6W2vqIg/QIAn2N62FDew1s8LIFyB0BqKxTpap1q5ySMbJd9+35S
RZYGjsGIPv6HF8qseWgW1L9FrKdfUWDMUdjts61a0TVgbgy8zyDkQRW+Y4Jz73pZQua7QcqfZcrt
e0YMPzVEBjesLzqF9wkWg6W4NHZG6AaWjBn5oCGYkXVoapnRUOdiRugZtwVaap2aX6dqJbEs/bpR
u87fX4t666PDJhXqAn+RNckJdHJHg5TLuBiPiQ29E8pDJlsRLEyz9Ybbl/3vTG/A6uDJywy/Exf4
DI/mCjdY63Gjyj6Z+QVTfu7torf2aH2aTBfqJdbRV8CfAC0e8n/GU9G07W43Wfx+KZnkwfvw7V6c
7gusSYQ0FXWaMSE3MMi2TJBvmqKcbnavKpv+brUi9yEPOUH9pCZ5WGD/sTLMV0srOspxyT0Aba3q
xagdXLYGsaBtmgQR1hTKtzrCEnh4D8JL9B1p1k2WPpgDoDs0Rl6/thkVsK8zn+7PWoX4rZN4TfUA
99zjW1+wt7Qgyil7KC5vILsmUt8MvQtmC3uAQXTX9z17mckxZUJEPvU1vGwBEJflEIts+dBoO0so
0celTBQfKRQ+5zstJU3/i3sTB2y/hGLTwqEnJr2FBEoaJAa0JsEFQkbah97QNjdQwBOptM+dz3RD
QHEvrnGHbgOGQoknc2LyB2gPFcXAyNQMXzPTTdO1lkl10gQEhQInN61sXUEoqhK6KBDmewHK8vLy
WzBM1jvFihH/wf3v2fjsdO8wA9QuQUxV/B5dBm088hPROd3xlZfjFUlaUxF0ogspZwh0fKO93mTD
bnsOwVy7KQEpHe1oGR9iIJgOIqUcYYMb/xVMYxQ0vyU1pVykCXT5+pjJdAI3H5MMoihTCHWIyr4b
/1NuGDkmpK5w8UqhCPA8xDfKiljDAerkNDHLIj5sHo9iX0K+xI7DemsClzbuT6nocdQYyrd0Q9mE
/Bg+pV11jpVc19cHLdI3e0O4HZRoku89DNE07vOpRHtZwis2BXvaFYYcj60OVL8puVfPwaQZrYjP
+h0oFKCwKfjtJLFHruJjXC06Yak9Rfs1VctMaMt7D4ktG8s885dHuCH1FHmLaGYbkfwn9zipAoCH
l5GcHbtlsEWT2v3ppGDOJpCZBpCLzDI/9iXIOt27FPf8P7G/+oAHcrHfo6KhX05aVx+PRXBBNz+w
WN6RhVwr56dXT6pFPsSqBl1SW6ynkEwbZi+Hnuqbsj9vqavwhs18iOA0uzs/6aiuTtdYnLvLy1Eh
3iRLHjucviLGJMawHJdTp0kjjPQKraMQQvD8g1iqFfUeLWEKOS9rKLQ3MuOWlh/9XB+AGtdm2W/O
OYg8ZL+fLSplnlQN9h3qpyiZsNGA0lqYm6xIjcJVJuxsU/Faeb9wCxdF57zKwcmRau0KCyRd0ccX
6RsXwXtd6J0tBtQwgbhSVV3ARQDf2HS0FJ5tLJY1emy7AfuWvR7nmPsKnny8s1dbBBYco1KFatgW
1OsClbFUlE/2CyMUe5flm/BdR1XLx6nVqWLgnesz8aMoYnbEopFJHZZYkOgCOV6Lm1yebS3WXZup
zF6Eq20ICLrW+aXZ+C4jvFtKRU8OTOhkQ3XjtyliIu8sWWJTRgnBN8465STYOWL5ms6mm6auJepo
RaKWrRC0cz1UrLslkg/ox99TSDboaEeW6NyfJb1JmCOxGaZ+M3UWAURW5PUNRYbxk/w0wUfRjS89
tqESqsbktHQhurHxonmS8ViFwPSyhxqJZ62TGazKEKh+T2rxW6sAsdXTikm/J2IvQHKWXdLoVBwh
0ZXVGyghz3yGj+HyHAlG0nESgLJM3GtIa5Qj6RNkPz9FkyghL9KxKQSaPOAV2INEh3QEP61l317h
rGQTF9FPDBkfJnBv5pKUurUXG1Rmq9QOCT3n+tbfAtnZFn/rIuU6j8m8pH1EQmPdHevMooWSeFal
P2P0aKKO2R3ILMJnFA2dYGAwSUYZhT6PkRbmN0yxrNy7GEWhP3bdRWvgwG9CmxS56MolbUkUAkvP
1SVE6ZWO1+YMHQB0SJn8wtfa9aMk3wBLUzNQyH5rf02wzR/RQbMlPZy8zar2uVZ0Llx9Nt/1szq0
xfuEYA+z00L50By2lAlX3kXrAX8WzLgtNDyEizOE1JXpvtUZXz9nquQcegAbuIKZJKQtDPLCwDGo
Es3zdm6fQyETwI1TZiTgwfR4b3Mh++/oy1ms/Dp1UAIBoS7Q7YuvBYU4wrzba4/iBqrTC5KLG88h
FrtzzHqRpsQgQIjTCNkPSS7kxM0t2Q7aYaL3PqxurcWM0dHtNd7ebWDwA6Yh3UmuBOZcbDD/5jpk
zc8ccH2vOW2RbR7UmNgvxqG4gVFJEWocNyvo+hTCtV6Hj2yDsjLK77OGW73iGAdLie2UqTi7qojB
+igvDnbqEDTh8QCC4kDuo3qFlY+lgMT5fq6fDvkVvVy+Y/Nx89sqa3ASxYcp1vVBfZJ0OnmyHsRG
UxL0y3TlzsfRoLcMuvQH1SG+nv7V9BnSYhCPv+Cq3ePr+cTnLyQlgi/8kBNmrXEmqq22Wt7NJTUF
P/OGoZeZDJYJkL1C6JvDHDbPMS9pxLPB3+KYoVNkYCMk8l10u5xf1W3y03jkjxdLtXVixL4xoqHd
bkmOciNOCiho0fMa49UImSTZVEsZedi1ILGM/rns8b4ODQjqP2csV3fWgMIx0QrdLcwSQvCGcqs4
AQKKf4o+kBxA3lhC0qWFAK8OJC1P7odakupNjelQpvCaUZRcGBYviZ0pBdRb+WnrztaL/rbbkPEK
9kSmezveEl25gw7NqKbMAAlBbp/lWMGs2OMvk7DpOAetSjMEpqNo01H6mVP5Jwegt0PyJN1MHNi1
D4wucsCNAvZAVeVlTKNoOxBlHzonj7ZMY9Ks1ZpwOHnL+V4IIk0tOpbd2Xe7j0+WAAq7yMh9L690
ZnZ1Is5ExjrQHHIl37jWRItmHWzv/lHw/SGjeeeydn13WlHPdzr78nts34WRbMhpgm7os+4GBBJa
k2UHrooagvvYvml16n2kgj8aYLYGxNCPI9nP8khF420/NiDsCD64VnHvtHEejIu8xm4d8owhIZru
Oo0BVhnAlE5qvOVDfNwawO7SFIIdCBWWDnUrtdFxVatgTg2i7Ib4lkuEbGZCI/WjHxoMZuGIjSvQ
FMCrP+6vHz7E1aPt2Y1r6eOBGRQ+mNFqnFeyhEfIUMavkA6tYNt3aUvBmprtRXzCfiAkrbpZVjAr
TIx96FtPQ1ozoqitM224x7OplC9lUpsueXo7EGyPwS9sAukyoIDbQvrzYVVLSj2wLHFXIsY8D2us
Ddq6s5UHCCNPZrIVb1A+S7FHKqWBt9WUHrBw0hP1dQosfXEiaF+4MP87C8LmfPzFOIfYm5YwMeze
QnYnQL9lvqxcdsa7usfEzpnrs6KcN3NPGQdrLN/XobAEwQzgyCv6HEihir5p9cG+R+5wMaJvuYOa
vfMxH78oxTAyILEHnvq3dkzhQQJAslPK6kR+Emee7HsVW3TOcv2DLsyfUIvY5kFSDabpm6sbpGz9
A9zduK1VohmQNBPprAW+SgDC8BUJA7icb1dYSJt46eOqK49VC3YcbTEBMBj6i5dUaANZ3dp2VPH5
DL2P+zvDY6omfdcgLsYy1cTD4vn2u+pN1aep9rerMBamnrjwHQ/QeCHNWlTAZ3G3hZiW54ibjZGG
pcZjHmuuC7VFizTgawf5zscYBZINHDgRutwiur7x3lb4UyQKovcJFw4NbQhnNP0zFbvE9VJPFE7D
+6olL5HzPmxeYvfgpaEBjlhUPIxTmnuZBBr0yJGE1lYehsKcq4AzTit7OKmboiJk8+zVFU0hHaid
N4UgMp6lIKVVJOKs7fB6bEOysLliNi6opFtI7VFQVxuU2B3moFAO8qi4XE6WwPmE//HV0TieQ9LH
QoCTc4A8SV2rt2AhQEq5UWZVFNidfBZ3+6JLaRurj08C/wZJnGKBJBzRQuk7cyUbJ/yG9qMmk59t
zSeHWIvT49SEb5SrTs89R864jjRlbGZhwHvYjzLW7q85Swd6oPy5D020+BFEzk8rhzEc1+HWtPkU
gepR/xmSGsJYwTCprPMd+6fyEcDSYQRunTX9ydKtALdZGbcLjh8V7FczY1FQ8fAXkfEg+mE/p6JN
5f/DKkHl1IzNtvYVou+KUgAxwJs25V/aB9hUrLV67uC/aDJ13WOsuP/RFnRcfJZrvPqpnSeapzgW
9rTHdTz7YK+bTQrt1Lxq7zg5HYJeXHW1makA2AlFU7a9dPS9EEshEzYYcJVQ+E9CzCOTa8S1je8/
OJpYhNdJ8+aaS/7supWbdlXjGJ2L7u03NzCfBhAgJHmxjfJGv9gYA6rv08p+RW9iNTF3giqDe/Tq
6Og5+z94IXLQfS4LSqVualiffTKu4Au0++klLT3inAW9mms7i+oFz379wI0BL9XmKpn0U3Ph19/S
3DtWj7mf4dmHZuaU1zG5ixX8nbPVYtaEzYZJFZT7OfMSe4v+AFXXjEzRXWrt8XBtXNl73BiV9iAI
oz2saQAQyGumLrnHGT7HkIrFBNAJf2v++t/7ZxLvQFDEi3qbyXap6fkVMC3Ui0ktMOvNUMjFDkJk
TRhrG3UL+85EX6n9XEZJTAmaFCz4C7Pp6KimBu3ccwWFrKpW6dWLNyRs8wGfsPhtoqIWyJHXwAPC
ZGmkdGNianll7+SHiyMRwmLtwd0pjP53r3dsE/NVQfzOE6oQPec5trv9nwlI07x4AV8feJH0oLsA
up8TtMqOOTrgj4sbqDDYdd5DnsUPBVUpJmbQTx3zvngzbWY59QM6GCWHbslochIPZaXmPJptXeIF
wyQ3umE7yrpTKor4vh6/G2DaoHEY6BW85GzPlSgHnRWtBz1g6cbZOPE7CDF5z55AOCA3uYaLyJ7Z
/E/YlALwHRKeEpTvu+n3ktBU0vRT7kSMXxysWlYyf74zMf2DryKPmJ8QH+i92ebAk1IUZWTeisb5
jbjzlGZfkq/IBRGjd6ECrhg5UNaH9AzrVqesTnGlvNMMnGEiYIe6QEqDQ+WGLLqCziFRdSVAEnoJ
BnH7x3WWt9zWgVynBwUGYu9UfSLECRldz6M4yyMycNdOa63ympqK87ywRiI7kxlLzxva6vrXrKQQ
FITiJwVAu3iZwLJKZOTkOo1MqyMMVG6GsBVszsJAotikb2Dwh/6Gg4rWTSFEVPw713ouQKdKmMgk
OSn5maL9lXGYEZN4sMABNzYA0LXvGSHQ3sTEaqlGsHIfq9ucYJ/6WoLHJ0wer5WdUV4NSqsv62/o
yLc+9wTlDGKcurUqzwTVGSGSGSDnDeh4DcVc3KY6Q7eKL/JgBkJy2LnLtG98C1dBjmQnPsbksYwT
BjkLWhgrqPdWptxdJuSeVi1wGqFt0rG5xURPUX7HiqBM1yJAM1gVE0w8GRZvH+9ySEVuudnH1mrJ
wBjv90VDCOgJhxs8lsFiX/RKgV2m2wBc68Aiz+68apa7uAp5F6plBDE/cj/PWEI9YBni0ykxuoUO
pZWbSmxj5vXTe3CRbKO7iBW6TELoGBJeaZKOtPExbj8VRyNxPoS2qvik6eOU5sBCDOn/lCLEjhzJ
9X3CFSY48utTxLXY1b8l+Tcec8/AS/Llzh+ntRrJtC+o2AiLeB5NCkLNjh33BaQAAATNoHA97Non
uezBz2wZxCA9jv5edTC5hlOTNiLAR0/CIwVXzn1dZmyAMVQd7i0dVhu2aDmiQBFZI1IyDJ8RzHbT
IVECMOzpwrP4D2ZZWL5lneUzUBaYQ6ibPPgdMjx7Nfodg5Lde5oIOzIOHa+b15Gg2TBOjv9tMJzu
hPNjIXXI4yPyMrNuTgXwJfX9VZrON8L4u/yrB/OWYTMaxOs8XmEDKRS6wVUqETWDz+t2chk8bycC
tiriy6VTw3Fdtf7/dM800EySNoYuqc2B8vY5IM7SUxV2lVfak8oSzLmJ6pK3zP+PUS6MZvM/Vh0V
CyWUwK4nkbEjIvzqwIr5PK/pmaL1Mbuq7gxq48qIqE1sSezQVCf6weOaJON0SKz/KMq9rsTtqOv2
jVbORHn9pN9gzBVOXn0p9zh7hKcyEwSEJ9A6bPWgcrnnGE0s8/UJBTZEG2c3MYUnQNTHg58FhIRy
CH/gqwqkXqhGf0x614azADnK8MNItA8vDQwtES2VBkCQ899vwcZUpQTM6dhGb0/Sw5J1+l+SaVWV
IvuH2ythOn7vsZH238Kd+vzF+93seAzHx8S3Ro6DZbSn458KkwEuqOMY4czW7xv+2mh6OSzjuSIg
n2NWwVVpDVIQEmpy3ndpeF/+W+U9PM2mM/KsTiMRqmwPU6yeHU+2PYG8p1MsnhJ7hfvABrXVs9LG
FLEoUP/ptSBR64EiKT1pUwqEROCwgYcIC02BtRkSPTJ05bKZfDeN0FAIDJExbfZjH75TJKDAwUuT
1rgk/uhl6pebDp0JaO2nufTylMmG9cc/kVrZDa6ytAdCIg3j8omTsS4o1rGaIJPNk3iUh8L8l4q/
omyD3+M6IIDpbYB3N5F76jNdcKojnRQbcf50w+S1iMfSYrWiqbdPE+Z4bIkPogctBKeZHGC2ZFqt
nM70eYPpGzk4hkHpTir+8J2bb0g7N4Lv2NGVcygcB1tVLTpLkRrcRvA9cZeszz1QgMqZwDaQLjaS
zF8jbc/pS1U+30UYLnLK4vfVP8WyKOvb3ORq9X/NY6rqHA0pCaP27fnoK5oYJcVhktx4FWJxfsdy
FBQMBZz6dw90545R/BNVHzq4FEoCMPuYQ6PcQp2gA9oBIhf84CVpOPtraMApPRy4zhidrJQrx6yT
1gJJhDlR8Fev7sz5xnXjeg0vNSO/gfw/AZH5Ztt5l1Kw9GXwk6Zd6YxhQFj/lav9z34w9BUB0hx7
g6C0Icem/M7I7G+YtA3M+5lY8hrLCNfqCr04GKLPbrIYLvGeXMhtIh5+Wk5kHoFNE4oS2O/HHLsT
lSyp+PYOq2A1uyQDLa6nnUpy9EoBCzegkZOwj2ybCB3HExoW4y2L66e2rofhGHSzYCs2uo6sNO1d
TwNFzaUDbhVxFaVWn3eRHKAvzkkAMcfzoDiwpqRbmcmV9JJuELD0STMigpsdC9DP8WlZ9g2Jkd16
G4anMaELCtqElF5RcO/Gc1WBR6jx9TY5frSnEmsLb8XafxmfDm1005WhqhIpi9q68V924FRfAXfG
SXcDlhPjeYeq4xqHZdPFYnxw8tV0+BX3B3tX72ksvbBVXXe7TxRVCpIT7UE6gCjJTNvJOazH2ANo
OQCv7pMmKKbUGw57uWrEg8OKKcuGW2AEdOHAn2TvIyCO7XCsbShaxu6GDEoynlsX4Mvah2nzOIGO
qKYRQ0s5Z1hx3yLkgl//TNSrSbVYF7qksb23+RlqDwKC8rvoXPrPZOxQ0Ynt0cVTCmLVEqVBBOq+
Xxyc+j42ztochbj5/mnYENRnqSfl2OHCGGfZ3dZyMU4bfGFOD2oqnfdtVyPC84Pu94ylBNU/dDDY
7Os4++z9f7sR9Td+RRaFiUyvJqG732PKDSNcb3csrYxxj85vhIJGzRzsqC7L2COPQGLzXvZBfCUS
fWBOSAHKrzEN+BU4AvMnvGMPiOInnKpBu1pzSOlMQSWwYC4jyGU6ASvmlJXOerhYmDcu1U8Z2MSX
KKnIYzBA6hm2g0sXLveI5xBiMb+KRjOVQVyeYCFBXnK6pMVhGUUYYf8b8ZLHgL23vE4iokY6hI52
pMVi5V4q0+3tJb4OgFtSNn5AwLWni34bTlWRxnjX4HN2FoMrN9x3qkR7dgaH+kaoWqP/TzUgfvf4
uVT9kl6B9noNWVp333voQlcrUvMQwmX+rU89GH16NW9IgpBBt+XTdN8VvlL3I7uuzgMgghC9jHgI
9f0b471qZts8CfpjVqTXjpuHC0+hOltBm2+8aPJnuIZppK+1EZ1VJ6iI7FWYiNzU9GI/ayqq1Tau
1uuUAv2gnFvIqo+ysfTfiUq0fP4h3fxNzoxE9ZyaMuK7fLHditVao0FcOgCNKUKVx1Q4NwXKYgPh
5angridjg1DPZ3YL4MomRtEvXQoBY8oQDiuFfPlmadVIjQ7//V48VZLcXifBpg4PnlxYD/pojJA6
HqJG/Z+saZ8FbVDk6a1ajRCCM3JC7kNaIL0h9nqtEmqcR1t3NjbGNSr84FV+csaZktP12qnGmfzy
80SQSE/S4Lw6TOv3aHR9frJG3AwjkGr9FPBlDkMdqMi4y3bK2v0WjcSCjXlwHKmpFC4zLyRkIJrI
0Lky61ajAl8PyTpQcpM1V9Jj0t54Q6m6Tnof5RKT9t/vLwMqceD/3TmzzwCTgJYujuiB7b2YjZEl
mJnyK3ONcB9m5Un6/hnxWnjA/03cBi3+dV0sx8WzgyB63LUeLsDWSVvmUlV6FdCQ1Q3rR2FqAm3h
QfB2bKAHL8DMuZGHJJtWzlyWF2dKwG/7MAVDpOI5jtZ6iTKiYLGfAkSaunLk3kwFhIbgoLQTKVQm
P+NsjDBc2OaW7mgxtSzoxu5uLC0sHWPDgOxhzyP/oMEnYHKwa6ywPkyGO0eIZlsSagIEyF3vxDZt
2D/u6BSgkFUpdRtW8AfIkt+wYyyyoBv4R1/t4wKaPkIDf50moK8a7vXibfph5kMuQQe9hybpXukp
IKQQskig/3Cxnra4IHqnG313ogkCpkBzlMXYEDk19Ayh1dubMWzxleSf17BZ5JUjSHqJUyWeOIwk
4yA5txU3i9T2WQqX59wco7Evo1iB3i1qkVLD1hNcyiPuefi4gpCrFDnTyFUN9bvXt9AEK/y46NCf
qkHw3PLYiu8sYUHYgVfJpduEgq17Huy5TAkog6AOOzg1sHcgmhBXGUpW/Y4GUPZW3Du4dcOZO/hJ
SmHO3RzQOhNMUSibxFdf5MKHJqx+e43a67ox2g3e4UpX9gbFrgbIwlQe+r7CZipwauHGQ+fUcDV4
gxyGuH/JT0YPeMYfDC4ZyohSxbVYGrR5OqBpvBEvQCRUBxsU8G49iisGuSiBzit44RGkRWa2ej5W
ggQLNEbc2dZxv7ahnnbssFDvTcNIomycD74+DmWS/r3tJUsnLDz0+p/w5iLctW6u4gfB/fo/8/wy
6osZtbGVgJfkwk9xB65iBgA9pY20i6gup35BXJmexPHfwOWhstuxKu868CQYhr70bLw3Uc+9vBW0
K1xAOMFhefxOK1p+VroIogB+zIpWTSvZBLb8x2LWyOCjtxfhXXmcelspy5vy71Pnn0bBeW9vVgUk
KplNDZmKbwpeln2lCC8MfVWZZuPuXyg5r2pdzY83ZTT6wkcgCTIHYC5NVMdUwocDsNoBYPBe86Lg
8BhmNCb9fugE7w==
`protect end_protected

