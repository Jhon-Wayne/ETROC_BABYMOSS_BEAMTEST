

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cn+MKgScMmuOXqDja4nBGV7WBeIF/ysF292lfgaKjpujK0iaFYzIB0eXWu1mkHfQiveaObVLOLk8
mrHpA4NCow==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lyXUbl1fNyCoynCsgKvsnxh4xSVW7h/6+WXSvHl9VdQRm1K5kCFQ2kx6cA9GQA5tjQws4LhzjH4C
jiN86wKYjDRH3aO0ipukeid3+Cl3Hf42WJLldVcK13r9M8WvFiA8f+TpNioyqUM09aStqFjdSjjo
csyM4N1L6gYZVbIwZOI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ocYp5Q+x2567q86I1MGJbRTpHjo6XgxppbNT9mGuUHy62i1N8b9FapDfB/As1HxRsllExonP6L4i
nOrPFX5dqrfhgwJzsoiJa+kQoi2nYY4KOnCB/Pv3Scs3TRpf2vM9w+ucmXI+o3jD4h7K+rgsIuZr
FCyudD/onJvsmis4CLUUX001F3EFidOEU1Q030HzWCJJNPr3CSJCNNoHPiRhh83y8YSpsqXjqNTb
qItJOecjL9k1mrcywbi+GE7p8H60wh9osKYdQVQMrETxJObRc2pckA7TWFtDMJerirE3KnEZvIsf
rkobt3565did5AenTYngu53T6wdatItFn3vIuA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vOCsY/SF8gPSqD/ldVKm/v7jmfpM33R1VJXD0UiCtFFOs1P7Tf2U4nhuNP3HANg0qD2YjaGQ6myv
dlR6lzeuHoYmZN/DUwZJGSaiuM1h6qmcn8qFSCISMqaoZHDjixJ9JrSXtSwMaPXqwy3RINyRZxZZ
n+tFIFvhOGXInTnHa+V/8xfZhzHNthwln8CBoCm3vnx5oPwRDkJfP3YwEDF4x4X447JPTEXORFnC
I+t/Qm3ldihxuP2e3EP3csValIaPqAY2BoE1dXhtaXAVGywLawKNeUCq9IIPVqj+KxyFneku6GTO
rnMbpLS30BN7Hk0gd76CeIpd158Kv0d8sEsmpA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dhHD5W3lGGtC4CZjL3T8nBhCONi7O+vACUFgJCKoGDg4NGC33+yxWhu78fODvPCS2DpLrPJfk3bA
djnpMpnwkBjzsk3CeFcPREHpRWWK8maEH4z7l4cbfw7kGO1b7+ekrWpBI7kV7eYckr9C0k8Ompl7
lKzWRDsnDke7Jkm2xJPdMkOOACVdIUAXKGvSGFbWAwk5E8Rp1UFWwqjmBhVrZ9mRxRT8Yg3dtQPF
q0TNwwUnijSFIcDGKDKuZ7CNTFcQuy/Tc8KslLW8lYYLxncygRHOjdaP0ohBUBQua3Io4qpRdfaV
InvJO9Dh+lNQuqdcaJvi0JXgF5GixjCSKmKlqA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Pz0913pmzb82uZOhWjEa23X64ev5vHsic1WjUUDytBBbAx/E1XSrB4wbUFgywP/okDl6EBGDGRvX
hoS0WBJe40mrnz7XPUgtp2OmS/NgcqGE7AhEty25v+Jxpgtk9CS4If7npTe95nuyFzYHVToQP4KB
6/HKuWIfxwjB8zuKPC4=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I2mjOeLUUoNbFKbqo1sWmTLCRf6eOvt7iqKURENUw3Qh1TB1B+bnN/F2rG994bfIQZsB5fvWkgKN
FG6KCYNjKLRpH6Z5OVJR6fOANjgDmnm49QXLpsNS4efTdEf+OXCcVzbqTKCiqtvuRScAI/nsT87x
y3rpJipze8j6Nlb8T4cSSjZaNmboEH9yPf7AxUPuY/HaH+yXbGP7PNWIOYU9iBJ+xgANh+c8Rbay
KHHeEYhxcnp20ptitbVw1sh77xQpfQIoY0Bv7zFymqzyeXKX7gS+ski/Y7A9b9aGTleTt87NJDz4
ncJx8n/LI8MaThS/7y2WYyDJ5UJrv2MXzJNvJw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
NArW6DLgUTVMfz9J0RNKQjF3uOF3jlAtbqr/JeNuIjDk12/bNt5GhyuaeKPAWWF8nFaIswJzvCSL
kpluCruNEMaJM1QFzTH/uG4D6OTlJtZGYTNP/eL1YyWFI8ID9cJ2XC0XO8jJY6iOTkHg0PE79y2z
sUa0jx8a1lYowtwoTgnCvryAkokGWPrqW+rSrdTJnr/Tkf0Y+/4AJLyiVbsbe1goMTa5R3twQWCn
QPnyrSwgxFkWt/IzZ7lVUtGKyhbAYfcriWRh3Sa9bbfgw2IBwqQ2hapWpM/rWgsOqriI4F7hwWAj
+2EyNGKkymLzMaiSwjEk7z/rkB4YTNUJdza3NGhmeL25nrWKYT2zkghUe1kKVybDWj7ubZ/vwlof
Gbs4bx4fz2ejjA+vlH/2UklUPm+DmhIy+jcwWuzDtjgHDiRGdeDgxquISfmyuaiwI7k76XEECyHg
w+EaexA7LYan2caKcegIARMdADSFgdOzSWr2T1Mg2MN4erCN2YwY9J5aaKAgMAf3dveHOZq+6Zj+
7oaZDlW7RX+zJYQDBtC/P9SGlrJb8z4z1dLpGbz7vFxglplExNh/uwnptWb4CpffDtuyslq/dpVc
sFUCvIy37WQ1/DX3qIJ8TvBtw/p1f4mZvSMGfTnxhvpgkq0eJxhTsdWIklV24qT1vNHe1DEflPYQ
O2X6P3pigjQ6ZRwK7BMkocrNLx1Q67P/105F8nw8YO4JCsDPZn+hF6nCUsl1gS44AW6NT6jQuKSX
MEglfj2u2tAE+5FKmqwxdP0sE1KBF89zLEtQvXKuMpjIjUCi/JM6PtDIKR/KYKIsgCjGculvbz+y
+y+7TnRuuAf3qFO3ajphvUJaL7dzgaSQryMqAgKZ8oiknHbq//ISGvRkTWeE51aw6XmZvIxvXUSM
0BMsSMDPgwpm4/oYE928tTNWOVaIYDKeNsieSsUQvH4N51PWwSLHBJtRZn/c0ZUnfk/JQmZinz58
vnTAjJIEGMQv+dfgNAfBELV1ZppHyniJqm/z9g9jLNqBlI0IiIseSZ4g4xR/b4RETk4oi3Hy74Qf
SlKVqnSVvscVMl7HMA7ogF5WEPidVOiqd8IsnFHUW6jgAmUQhrBrtiT8c2DfoD/CT6KRmQiLqzN3
zjW0Hfr45KdY6avG++OZHcnRx5aXPIz9IO0vFhXUDiSpOU6Qfkv4ASpKancsgfEOehMIQQc/kWBv
JEQklNeh89A/OnIs4r/3WLvZdE87BZwmasVstpThT6JPhIHPEGfjsn/1g7vu9QJD70URLydthhQ7
3/+jDIKxiXDpaTyCXrPh53Xy4+WC+MDV5mbCdd/Aqo/QLbZaCfweNIaWS4U6EiQ+/L8PVIb3I697
9HqjLRNnEgM4HDHZXT1tv2WQgEpadZfBTXROGIhCDUUfr9vwOJJm7RL5wMVcCtH3rkVf5WhN2LJ6
AMZ5VBQmuwCX9IOr2ICpnfiQXb5C01zdXaENHrCHZQxqYTojWzooboQjtlTW3m1rp9kWu9lewlL+
Pss0Sl8diTv22U0Sidonn9gcNBJ08Ym/W2czgFsnhmcR8+199HC0+mR0DTCDKHygkMHfb/H5huNg
wAuGDpUMtKtdgQmuG/GAPGM2RiRZ4CpbUUpI7Z50oNxQwxNQwVJ0qLvlyB9wvQVJtXoAu0tQBNp+
r+/VsnWLciZoUFeArYuTTX/YywdcamDQYhWTK8YOXGQQnBG3ctpfY8p38M2KrjTUL3oQKvn+Rg/5
Ij4NGN/BPKTy22cAO3Xr+H4QGQOZzc/FtUbeZEXysybzH6J0xemiJ6jBGSCcD6lrCntuUWxRyZhd
kFpM2ez/7rl354TYzE+/MVevx6YPSR54CdEXo121ZeDc3UXD0fYI7X9h8CuEPmzcBCxop4gHBfEl
v2FosB613IN5ZPkuUHp9vFAT89VidAoX5ZOzBZR8jDONuNjH3/RNlZSZROVpgAvWQKlyoS65ziiZ
6NMp/VipcGI+JqjnhX/mw3qeoxvUIKutVXuegPdVL008Bxwja4918EhaE/6t0WX1aKd0b9S3a4ZB
B+VA5Vjf3DHjqRFlv+HjwWG8e3XLmQj5wz1CKRrEswWp8kdlmhG12EcN21s1k+SikubpxLKnKeaC
q8sFCQYS7wsBrXmgS9FRu1N8gwHUccBMhqUf2m5tDuZHgRmH22L3ASZv5Lef9gVNjX6cpuC+DY56
ThBAX36pkYxPcNvtN1Ku207MnuuLrpohe/TYPnon8zgOi81H9vTrplAIExZzriP7pxC04gqBk0QS
1uoNPniHy4RNQgRuFPM6bFaXasTjR+ql25+Y7ZnD5Th9uYL2Nj5kS1Zo+KmwZN2SJ9wy2f5NWqTX
ctMZDphYvgxlzVgizBte78CQ66dkEHRQYxv8o8oPBDxVKQ5ZOO88+SM2zHdlEiiCbdJTz1vSz/j/
gYq5sWa30511QoP6jg1770ZcFD1wiQHLkfLYdog/9sWZBcq4b1pS/0dH36EAqx4GA2mYFHmCVG7w
V+NffQymu1kAcUyXevt2J1LYeqCtvJ0I8HPKWhzbvyqb7A8tb7a0hNqxr7Vp+BzREiNVmw52Q21G
gL182eRXUrNBvUYLqGCVOlnq0ehEFyqng4GYOIUv/p/C6CsOcFzNyZQpg+ViUnF+du9o7APgBmTz
HlRO8tib5s7swPIJh5iO8V0mvtwWcxa2HTP7eZ65oPkq5d8T99C95FCkvo1eEXorq1KwPJ8xNMtD
EP9o8PPnqHPwhqW6oSqVDkoXxGox8O0WuE8amg57zSGUbpX69XNvXSOowjFkL3zC2Sqn6NxydPA8
KDDwSKAosZgeW+z/2OB4hJeR32GVeXsuj9i3ieQ4Wgr75ypCruQSFAPTg7LjFwtCfIzZBPt/+uyG
LKmcXqKW1k+o6CeQdYo3uucTBC9WBb71Nxgs7/LS/6d1YMId5muBA/abmeLVUcfeWJVUKckYf4uo
Mbi7a8YcYX9rmkCWP0+UMdBy8IqaL9r+mHYHEUFBSnd+fBxk24KJ1tEQZ/3l3o2zDS3w4aAd1Ro6
rD2/nVP7n/wi3iUaJ+/KTnSWipcIs3mSKaJUACWiBvsbwUORzapRLG8sdN5xRVojDGRzg0itxuqg
tbsE7vBEiYNSxarqAPI6qLB1fwDLVQZuZJYbeAglrT2wdQKBZaTd+1Zgukq8fsU6sNdTxLXTjceb
W28TTdzruUKilL45XAaPnoC90ieX5TjaZ3AJxAOWzYYpTh0b2VvTg+poj4kFY1vu2JmnnqWnRtxw
s827AYIVB7rPP93Kus2rVRSafWlgMCoG1FNpw8XA4K5UTJq29Zo3V8z/16tKH/TJI9pDjoABf3RQ
6lWx2d/Vw94Ux5VLHiilEbOZmVcDk5VbLhuaNNrlcsWm9Z5XHtg6RxAJG/kKKU9I4xC86ArsES0G
uSFTSY+2ADopq9F0JmqnNfndiSY+WPzFLupfQUPKqOTS5rwqKl0DZJtgjxCMIIcfmrIBHozatU8J
cOAYHY9EwxmixRXsLPlH02DsCD/D9f2b/6gMaUtGcoxGVuCj7ZL+c3K37dXRqAY/FDh9tF09bOCh
B2U2T5VEoqWF919CM78YGw5BcNuL7ECa/+9/nqk0nl9qxi0py1jduqYCkA1mO0r2uP63GnKDuZYJ
zoTyJfTxkxDbRCD0+g3WKMHQFGFdC16nnF2iZlKOv2S5Obg/cEqmPZys4GObzMMIoXeM3dEKgB4x
RneObsjxbM7GqaP9pDNRO0J3hCEbtd4cjPhQuZukofuHrpMNGrFC7o0ojftUPtJj3r/7dRyTffsN
VEB0UrGyW2IvpfqJZ/1Ywclx9+MqSPUaR5F1kb61IjklSr3belM97M14ei9OjluuQfAMGt3qhzrm
yHqkBMnUKwMVkpoSi2LUdibSELrFlEFBtp51PYX37xjjGlyh8u8yHJrZ/nCUYIAslLKZ3HzuBib/
2n0qh+orgdzPLurJ7AhBYyWheJDgDmNm9TBAVn+QFq8ryLcbyrlOw+zkmPDcw6CbwUU6earkFPlw
QglWo7jngkzvqFjvaQjeKztoWm3sQba91sfu3BVqny0UxjBbb+blo8mDpZFP1VnEjtgWje4xzIsb
Mms6rwDyTdLHUNTUuFgAlYImYBS1wqsAis4JxuQa7USaxX5vpcNA0QV3nEkiRnjBqmFKOGhPvHQw
X5+EjJYEVs2NMKsGCGNDTq20RweQL7nzo0l6FWaJNWPpQQKJmgsNZzihBs+hPsPxFHEaUsmMu1tn
zCVc9lzmIGTBk6wGjEKYZ4/lZ7Y1IQEx9oyqPTRDo+89sw+LeyscQQgOBHAWEDUtqzxh2kJa3sOR
EhDMJf06KBo5SePtVBAdLCkDX1h5lcyNgPTNw6thlAjuzYO44C0UISLVXa5X8LJirR5RpGcjiMUg
cgR4JIx1TJBEAYpFbYKtlYJy+2XoSyv5HhkRKlpWcKf+vbdFDpPG79CI1uu2VnMd9gBNZ9eWit8x
wQkkklwkAbpxwnhznXYuE9kw5Upvognoza22Y7NMq7J9bQNIkvCHTTkImjbxRkSn+Jlhto9kuES7
7Ljc7NYgBZ8W6n22cyeEWHCSuXDyYy/8AvsthXoNlPsEurpytp7sl6CfK34GJ4M3ZvshQWn7gi2A
UTaeUf6T8tpkvtXGayynsgEl6SYoSLBPmDvWLtQFvDOz6LhvpteHOm/0Ntthtsby8DgAjrIeQDw+
77uNkn8YzSBPK5BRkmgHazjJ/3kyXZis+U00Y4CBWS/aat4gkXwCkkWct5/3hiZA65YXkIgUBxOV
ciASZjBkH5aMFIMJlVs2qOhTR5JWl19gf1OjVxFqBWvv7FTkEmWDIK74PdH9YOADAJ+3Sh7ujKf2
ulfkANTobwXRNxE3tX5m6VXt5QIh7o46uS5ZAYxRFaYD5K3ctGaEa0rPIt0eCZq9P7msoa6bC7e2
bnynY9UWm1nqXOMdZvsICX/u7kpVRrwQxE7mUSbH2NPF3444bdAddswPViDMi9ECd+c22SiD1CI1
ryggUDRKFpFBGPWhTKNnw/C2/R44vMmJPx2UMmASpm1mm1JOsfmQrnTVIezV++py7AP4UndXhQdn
t7lXPD/e/JJxH5/zMlOP8gDVZtQy49qoJdxledZqTGi3BrFjW5ntIg+v4g+lCFdYjFama7pl3KWi
paofC6TO+NhRuyL6J+kq3sq/XzkiwE9lkWigxr+BqWyQNJiiIaurqtAuOYhnP3tjBPUTW8V9taQg
n5h0BzrBbQbiyUJeYjVuNB9TgCPSwdI/+md3EUA3109bL1ORQtZTOCaMMUtGCaUdF6JlUefLkaBr
3CLUDqy3m2V7JuOP7mxZ+raUgAAJtWZpZLTBJQHj3+Gn6pbXCkBGTO/JW4lCSI/D4yYt0DrtyQTs
BHFBrUV/0++1ymCy4bR2EeGzZJLQMP2m6iY8coq/jB+aMoxyKmn5njsz+vBaaT+943W6f0FVma4o
pD0F3STjXao502F/A2lyulcM1oXVefZMgpGjc1xQunm8ZSfolkZsv8y3GzwVfBPSEYgWLayA+GOM
jMl88AH0NyRmY3L7tn2kewP0ekdxAesagUbzPRGhLHd9lA24I/wBRUHd7uDDBX7LWHH4BYXt5H2+
elju9vRvC6m4ZiiSkxc6kQS5IesJjFyMfxDNiaOpAs9ZXYpk26vU3nXS8fb0xWGzEQB2Icflv3R6
VZpGeRckz/+emq1NJK/WB5WwQYcE9zzV//u0iACLPRr8a7fpMRCknpMLn1UPW51ejl8r2HNoYVu5
cPVzPxsknuc2eenZ0ixHHjCuh4P69MwQm3sioiHyZL5VTg4ue84oWVjNgkyySc04TmWpUAkc8F8U
LunWKickf4JK8rbxycvgUSBSULTuzZ3w+bFYJImLy76AYvfaCpRtMNsBxnhiNw6n1XXbc35DFY/F
mf1Ez7CTbe5V3tf0ONLXpmGJaPn+RFpV73sEqImIEXgzxC8ToZ0LBCfiPJtum5shOJoGCfr8g6Im
Kh506BLk5UY55pmDLNQmi3vjZTbMvQ9sgvSGI0Ryslx2wqxrB1QfOBIEsCZ3etXxelUj6gPz/TGp
FzzV2zrVZc3aqWHgAKBlslnH5E+5jKwTnOHVr3HJYFEXNRNZo8UzJJxXrTgHOgp+eCOvoRB9WVlI
ZehWV/kDgqGK2YveBi3rSpqJnQiEYLXUBZqLDKC3s2cZFPIHOTWVIbdfi8s7HvwPYJdDJ3zv4CFx
WuC5Asz2fa+GxEs24rOZARN/E7an1BCXgtnzOqfttQGtjNuFEG1hp/d5UZPhxS38Y/P+0trgCDuy
XRxko89vG4651bg6BPAucl98DDMjV0SMXGzPivb2Mfik6cu465FNjV7/xQkAPD05zmRbmBb8WeUj
LUf/e63MpcMz9N5GrBlV6CtemUkHCERcroYuiODgknBwe9rFO+ydzRbsaN90e2PXfFrGAmFRZhlL
EE7B57uK2XCORsPOepD4qJhPbLu8JgZ5qz9RVjGtbOYl7YsM9jY74rszl3TE8Vw1ahez+LxknlF4
qyccr6OR4XYx9n7JyNi4gsu5V3slVyV+VFt41VR74Lo02EqudfxpIbaT97M+bLU0TAJ12vYprL24
zn2ZkIPIrmFmXqdWx+9iIflHb7kfTKaslKh0MKN62tUkmAcWh/0tpVpv/zhPEns9JEii/dxukKwf
ad/NV8d8kOJqQRfoHnXIju9nV+9oWRii0Z/+UfLJz8lasfaFFiqBSYyXWFFBt42Ka9D63OBf6V3U
Xn+7q5gd9LFz8vVHm6TT0RbdVRDo+na0UtVdI2zkyRpem+2urGGB4pJXCYsUyUR0Jt2q5AoT38hH
lk9F7UTpmhnHIq28O5PDb/iGeUTc9WEAKRHzm4i+qWB+o7nwnAqs4hH0T63jryvMrfktIqtbJDQH
HBY8QD751DZzFNxeEPggKSI6F9YOINibfhHRky+QThg9iSH5qNGC5QlLLAJCy8bGir1BQ73poqzz
LSvqJk8HsdFVa9Dkh2XD+EXErTUk+QVT7CYX31dIObh/VjahaS3C+mES77yIJkk6YxdviaQn9Sfl
k/4TN1TI2dEt+TlCFSS1X5v75zaI5WaDJGZLiMJe6PEjnkvuLoDfadOHkhPjQQU22Oc0cQlSHzRR
W24Ev3+jaucMeL5sPp0PbQVxScGaU18sh4TcCuX1l9Vp+Rj/dKVfY5snICiuihjqlogfDTO5+AIa
6Y+G0Fe9fYHpHW5crdOqqpoQD8C3or0wy3DXlL2Lru1mtoZobI1bSV1FVO23qitMcpYY5OL9psuO
BgijaqoQvbCNQ/hC3dTY5zM9uufWkZ801iIgNUXnH/iod92h0cYgOm4ugHLe9E7K9toO3MXN/PnX
yq/fvldnzbgU5Spdg5PWII3KGucZT1vAJKY2lFhvpN4T78VpgZRyyV2BeVxGpHACJvV7jLCa7VlV
ggugfllSTHr9E9v0FVRxE01bmSvI1k1Ta0Jal79fR5zC/HtGZR7LKs1Zvqn32G7k+LKc2yn1qBAe
9P5x4x272uB0Tk5GcomelsSlB62aPNSD6QkBcsXBMZZ7fFfnjz8hYUtQVBFoQq1aw2hhLaQuWLpt
5ZzpQifhHo2BPpIDu9yOA8NALnVjCsayoyCKTy8r8LPTnZ7Ecw/gmph3xNazI7E1kmlto/Lizuon
QMGsU+EKpRm+NAnPBrIBdzioovcyZ6YWR7F0/kfhReQjhWxMEhZPPtqkHkJlL0iUxX2S4ju+fHOf
vlhidH+sodMAqXkOpQcYVs7NLh0KJKTEb/7gdf2hafmbzD7xIzgdy8g+TjnNY3J6eClJB0YrZ4hG
zGeW+eLM86UZ9jdZ0j8OiYzKIxx2e520CEZOsvD/yfaRXpLksUF/6HR+n7uZDP3U9gSEo+R9GN1T
Tgq1Su79KTNzmgwcb6j7EYR5C64EXvMkvMoj0/vNF1cSbVprjqp46PKyx+0wvb1jJy/0r1gBkQVA
KRfiiqjJuaPEEh/kOfICoD6tbOHPNBNKZ6oepPRdvAl/xPZqcfmHe4y0AX7Kizq2u6AbcaW00Kda
X/1kAs8i9JR7XG7gHebpmB6iGGly7LHLP0aXeNwRz4WJXLwOGjgrnO/HesOzUWurIB2PcGqXUM5V
kdFhVInX9NIAi8mNte/E+sM4izRKmcY64eqDv0sxLVAg65iFhq4k65tDmKNO9q6sekUXOyh3mJ2O
6rIDivRJxyQhYUTApaWns/Ha7axeus1uZDZpc0nPJipqyuKk5WeifdyQqAXk/dH8aNHNwSSD6MAI
vWHKf5D5py+YCfp0ymxxIYb3ZQph7fDq92ZY+BOqKSwuo0tR9OZ5htd6eZEIiESUsOu2DMsCQwO5
7k6ZNwSWdhxDQawntkCFrqSTB2/0DYin8zuY8pAEglIE9lrie9NoBufHvxq81bAw9FpT1uwqeJEU
9rzLbBfmtAV6Bv3D9vvzfJZNL35tF4NPQ5/PMpst4rNfVrr3FCfC5dRb2Oysj0Mqw8wXZh7JCqHL
YKTKa/glRw/UpCpiiCUuf2jzB3VQft7iXDqRDhwm2qJMQEQKLs9k7WvQ352TabrY/Yo37WziaNQl
1rjCDgJ+jypEO6NPKLYOM+RYfcWm3REdLcvm4ySC/vBMUGsd6gQsBQ0c9lXQu9dPHnAjRYymJNVP
Zq7g4m5xDxteSvCh0MU7NAWPObIRTfvvD62BahyWlfMl8Nrr2QyergLs3VkpcGkflAspI+payPwJ
kM7h+iagRXmJPv89j1Hv5y8pnTBZtJFGkIIPmfZRQBPFYihxvFyHuoQ1p9hfzH2A90b0nPKK9ooC
NTMlbQb3FE7sCo5Vu5yGp7sLr0Kcuf3msOL/D3Q68qB3rrl0ODof8GrQIm0YatQcjJdWP7jqbH6m
Y2+z7ex1N1c95j67d1QIlAtu0AYK53J63WoOP05pwbihOpez3fl7BQS6M74D1rupzlYaVO3Ab+wG
wPFkx7cKj7MQZ248zFCBW0RCm9Eg5OPKqZpVYPwb0wsN1WrWDFAjvWy0A+71KL2C04PRzxliE9qQ
gzaopeC8nRhc2Gk//SeFBU/+s9PTFxF9dj9X8ythSAzPs+8iiQGk4jWx901MDVkk7czfH4ZMEBx1
jEII6cLdyJ4h8vQtubnDgEgaTR24/H8T5BQbcuHBVF1NI5uv1O/RtwxIpfmlVrVpVZjduTcznuVp
oqFk/Ig8v7t4zLsJWQevNU20KhZ9VseOfL0hm7t8rSJkntv0V7rP4ENwgu5HGXwEF+pUvZSDO8Rw
efohIxlOyxAoKkjz4vhzBcJG3CL6fTaeolyYYqi39KQ60p/I4B2I/vig2MnaTC0IDvCuNa71jQYI
Lxep1mQFOHiBrS+KR6uV5UlMPOx162+qtNURRtg/bdMseuxR5v+Xbv0yJyrDhj8PFinll+AGw7Ex
b9S5KRLezfOi55YJSTWQ4lSvHPh5tG4NhpWm9Wv5OatDsBYV7Cu325Vp7co3PxBsvB5+qmfQqQFX
PzP4jCDgkiIV1u5a/WVBByjsUiKQUM1YTcyA8usO3KIFQDK0z/oE/B/1KXwdGj1gQWzEj6x6jVy8
n5LHngG6n7nTRern/rCtPlMiA+G34jfqyLXuigMcMRpuRew3TYfTUKVEEJ7gDk70g4kMg8a8qlnQ
T5uNdT8efXDmYs8JQSrKpB5XGlc/6UQzmjypLQJAh0TAT4sLu9UU3C4gsl+A/6E2gdVtFdhlgaT8
nIwERV/mHaontEtkC4epsZHqaC2tsgTUrTl9frkbMo4HE5GUM2NAeTvrWRdpncRjgW2avquHl/9h
DO4/BazW+ZBNW4jyxbcZ5T2gkq3lSWwOl7Nvp57BCreJl/6KZ5g2fP7Ofq9lCdDzsVtNhPEVEBP0
TuEJNpFes39imSixliqqO7N/oaIAce6SuZkzn0GmKne2TVdGjlyOX+JEOXDwnkCi19PaqirgEkRM
SNLcpFraKgtoqrsvaMMQjvvc2eoj9t52cf1sDj/hz86y4kJ08NdPf51jM5qyUVu//Ncd9IHaE3+K
Av5f4Fj46Ze3jh+FQrXKZjPYpi6bfMTzhwF3BHuc0UeiV9+2GN0901u8Il4jVgyNjY8w44ezbS/I
/Rjkt+urJnHquYyP9UzlQpkwnJ+5C4x/vhVXGCoQVT2pNUDPGcejtR9+K7NTfknhu1JGrYwhmC/N
Aa1ynhyqa4QuTuORHW+aFt/EARjf3TaV4TUD2v0jBs80b2rv/FAGIDDea63HQ8v+0+ruDkGWAXXS
33aecX3WeSdpMIHfAjH+ygKc3eZdsutk1PWy949gwdCFC+AHjP2EEM2ojqS2Bdv0UoiGjYYPL2nm
z9DTVHwxF93mb19igJgDr5W9D5RlppkGdRk6CPHvfWNcSf4sV3oCNjo1oWlC77YYifykrUlqdYge
kNvmr4pL9IjA9TXTrgf5UAufGZrAS9V4xIcCb6sp8PU7m/PcxlWivgrG4FPoo7rWEbQ5vaMnDiRW
X0DyvrxnCL5NF1ouCTBMlKNN2EDtdrIFGJq9qFhFQY94c6KikjIf5tyFpHtxpj9fb5Vs7HCPaj0v
dW3viKDwnJz7eGXLTPA7ulE0o0Dgax5CB6QHhqRTUNKctr/BoepMyh9UmJ/8bRiq8C5vVhUrkAF3
Q9zh4sOOtvEZkf9gO+fEwLtvENwFkOLMdQ8S5R1NHvzxmA5ns8HsMkp6QC3qH5yKjJjDrXbjYkl1
0MXPiPlI4kpO46nMrik/52JL/z5kl6i7I5kJKcxrKrHFGZ9QriHP0vTLfY38aHVkn7b7iuGzbeJ+
x1LDg8ga4pmWlkagme9Hi1GkxBps9D6PNuusVGmy5jnE3yiwkILcY0mLAxci3Rsx2IN7+PPuBWs1
NBlC1TVHIbCEddywSfqswqLAJVwMFl6xyzMI5OU9OmLTju02Yse83Z2rFJXSfQ8g8Z9pvaW8gLOG
usCgZesHJF2MI2FVKaT5Ix/OV7yF1Oys/7heESGyOOfwR2UcrxnQGWVU7cdRaS3gdffOXFDgTCLu
/0v4ccPxqdO2E53vIQTc1hF0Mw/Pm7MMAsaKmshv3d4BVHa65l1lQOH/ARzrq0N1lIQ75bDn3JdT
l+DvJYqRySgll3Rz+imQ9NXwMCb9ERYrrQe/O8zhtb82DDtA2+4bjCzzO6dtgT3EaII/e106sa30
zt+pwI3woZDE6hePYE5H95rzDEkPj5pY3EKBEGflp13IJGFp7LB54XffqeCXxitrVccmakqQIBk2
Y8n02ZMe38tY2sZmXEW5YCJ9HYtiBmuvgUBLKlF+W1mRpJ9mLrWWC44AN15Em2OX3ZOkYaDIBQIY
o9ff+v8tDcz/zj2DS3nc/83s4gQRco7J7v2GSKYuej5DzUYRLEJlGZW6X2CH9Rv5JiUtTUOK3+wh
lNvkuwXoKBVSRQIr5VdlCkN036iIdA38ZefVIONhon1kLQasP9fkVmvlSlwiNUvuUUFv+b3MnFDV
VPXA0iU8dg/8aGSayMUl2BfZ5A1LABo7LbtzrpNPw2Sq+o2wVZomz87MNGURbxoAShVviJwPSyLx
hIK1eFzfvZV1HjprD8HLhJnaneH213HiEKE+oqRiwD3lCwxV6hyHbqKZ2Iso9QND2uSLT06yfKD/
oosadgNEELxbRz2EDGPn0gO42TOzPFeIsjerZKrTgezwt84QjXDmkLHNyOW9w29hYk45t0MYOgd8
rKu93dOs4YhcwMqokQWMKxAuMR8/WDr3lktAowas3AJf88BU9q9T3jN+ZRjYIOmDm/iCdkzpEaJN
ZBY/YJstknGO2ysdumbd5AaXXtASW4yGiCqYlj98M28+USlNZAuONz1hTUoCvORNS4D9OLj8PPIu
xw+7Sv1WCcH8b34oOG2/kD3gJJ4ZE0MhvrlqFXNXejTiM0Qgiom2rbMCURu+VqyX3tLowlTF2kN1
fRgmKnv+AEscWS3KtP+AqJbbe99vC8aL41rIRhNREdrRSNlCDc4+EC61rGGdQOfBPdy3GjvFP1yC
ULP+EFj8EGO8vzjvszY8fbeTnHiDOWcM7qXtJqJmV6nD/UOi4rgWQJ9uvPWajRxpOyHELNZd8fom
lDYTGY4m3knM3h1oOFnbv36OtMNCtgGc6gE5ofRU4zrf0YuiQNdPsNwTAiMgGdxNLtor5J+Avu7k
GvvXCGfGAoxEpWTGdCdaCFCw1kaWGpGBMDzExFGfZZpWKZvp/yGwmNsApBOfCwCWGNYDczydwCE3
Qd8Gr6o1Fzi4/LZridhs944fryFD5NmfUySThXIvDpoVJgkOfOFs16Dm8/cgoo4sZ7jScEyQgsfd
EUwAor14dSS+hTiSx4jxIKW9ztMUOd04pCEdALo1i7VnSQoDwNNBpVfNFsC+rdW3g7oTOkveUZNm
qrKJ8ccXDoVRtUh5byMdM0+PV0+6IuxmgoSptTOUI76g+TytH3UzXnOw+vryP83Pt4UY9YmbWD8l
mYqQHfTQFdj+UVXBcObt/vtbFxW3AsCz82paz8Zs67KGx0nTjCZLA7Z7iKQLtAqF6WieY70vUARI
4nO71BJ+gPog9AD7C26jyGMv26Rc737zj6al4vA91bra3lPRHRf3KiTHGtMsQt4ZaxNn+7aF1Waf
Ac+dxTHDhPzqQedBDqawYvWdAsbe1P3YBdNSQGuO7kwKQrD87TnSqSoJ+zNujZF5SnArMGDC+nF5
APugbMUV7Y43FXj+Ehu+qQJeVAfRUhH9V/KQphn5vJr886oFBd2XAMOV/wFIhL9LrNf00dJ3GdAR
UedjdimoavkgHROn8zAaDNyDvJUdTbeptUScbwYRVK2OcqwgtsRXg4YeZUFqddPXz98CbwJvVOma
DZOxnRXl8w++/tys8as5/L/uvrThVr4I0+aRID4Gru5znYd7G7fG11d3T6nmTCKQD80q16Ma+EVo
ZYilkcBhX8EPcv5vQOdLAdewJ2xMVgzRpq5vYlGIOIahAUGZZwbRR5QsitY4A3kg5Pn+rPcUlFd1
zPGdXN3Jg4VvVffPuTvK7gEPAurMQi538qcsCtjuotsnY3XzirdHTvgIn69QWvSDqyHkKViQSZfS
K7iWmCNV37d259Y5K7D2zA+hBypvNHSVedgO+EZtLCsn6LVkgS77LVTt2tK+hVJAxh2ESmW5lcaR
fQQf3V7dQcDtEsg5YY+ipeX3WpcgzL4dJCV9B8cOvH9+sEVTuNacnJGY4vNE3JcfjpapEG5tSynQ
AWjBnk+y9K3M1Qcqq9z+iSVy6hS86EUhhcbh3w/gpQJuKimQfb1SPYCd0GYI4n88+Eei/XR/LsLa
M65djtntss16xsk2gPiAf+JVBy7bF1qWBxAKas+ttem5zdEA2ucaT31VYnyQ0zfF98kbQZ5krZQ1
jKnU7tT5M654j9L9zoQ/K/5PcMsK4sCIUc/MqhdCNuQWRSXHdbye/N/OJMRG2PBeqcEWzW6Nd4dP
H7z0ysBSIXJiVJ/33RCyGposF4ba3TNsEVOdTz+SRcGtOFuySvtXOkql0SMxGAi1xu1+umuXhFd4
6RHOS4AJ4uwXMRSpeYT/AdqdiE0sJuTz5MBUz4jWVDAJ8SwiaGJzYCHleCnZ/I490NAIyZkgO5MZ
twYagBmq9KmqSqE7h2jkzAZoTbq8+sBopMqlxMrvsieusTbt2c5c/KzVXmIW+fVSEomV5TlLvfWc
xXI8juoBcyUmHxqA6aSljhzNeynX5tdmqFgtnrR3KrPjyjVJ56u5gzecC4jBOyivh2RZmSiQb4Xh
JloLugVWrU8u2G6c/NhDiL0IPaOH15TB8Ya9p/5bNSZJ7/xOxcAfOOp8jSpUvKGMPGjXqGjBckJk
2Bepqbt3FWIU+hHDNbkMnnfJ8OE2scLeo25VnxMdMeZAjtsyMThrUfYSK7nscGw89UFely5rxPlr
4gV6nvLYxorxt5WkgJsocl5AEwzuvRilltp9iMVxOfq3ypvgMrTUWkvi5VbkoeHK23Dx7Y0KZ8Ps
64A02rXaBgP9LhYgek9B7Ye0UWatwV9wquI6IG6bNct1aE9Gq6sNJ6kUzPQNoHK4oATvwbhLN7lo
w1mS6o/vYrLyLUmYO1qch+V6N5Te3N2K21GDAT75Sx/MJHNQR1rSAaZveEwPfJGi5SNmhrLJY/HQ
1RqVnWU/sCi05ODIJAnj3FxktGNtY/MJh58bZUzBAZuhGkG1jjoTGqZLu1wTOixcGiduhrMKH/Dy
PKPYRid/MZ+yOBmMRVqyavZ6gmwh4zsQFyGCllAUWiHUVcmIX9YeLoWaFx8IpCfjUVGlX4ONJ2NT
6ccH4GuI+EUtYwaj4QcqFmP1D3WMEI6oHsinqga9f/VL7ehfKhaP1sjFWlTeIOf0wHCvPw44jugK
U3v0DhGlsChkWDbJlmkhbMny8jySgt1HxEUkcLGAmNhkpRzCiV3aqiQ7FOpsCPbUsQwKRgb7rkqz
rGSe39vxAdcuE2GJsxk45b+J0HBarl1BvA+VHoAZjG5CeRmNdTaoVqRLImI89NLpGe9BkAL7zu/f
TXwkXtgBv9Jtvsiok95C1mjfMFUomMWm2iHiQTyMFjb5y9lJtJ/SPBbvUaoT01T63GluKXHwsZQy
HBFYdEe41CQtHzxtEL0ehaDe4ZqC+KdIh0Ar7raJoVW9IRt7HAANSj5LPZTOkTiwSzd4aG3b39oA
aswrul/87u02NOuTLA2pQlukS6/AAQzstV2kUimvtL743YayXDAk79qphJfmll0qS5iNGC3nQrJm
BGCzorA+YwmQSm6qtBlUffQ2I37+BC+Gg+jyiuUnSWytNvRjHqHvxirSa2wFU5mZhchwHxePRgrT
yV8ZZrrb2rTaG6O4vO2pZm8zX19syCNuTB66CrzdMW1oRhC9Jebwdfgd7HFw+qGLHpbJTWXubqMa
fKaRGgY27xCC8cGSTM+DhZTw6u5G7NnJOKP2qhYR/KP6BZzwa2y7eoSI4Ynwgz7/seVwk31kVO+2
T/RJbduVqCqA0KY1y63WtfDH+xP1B4y8d3pBNq+tWUBshZZFsIA7Q1A6PWXya9FqVCpvtebIhQT7
oYUVW78OeqxFD7BRLfJ7B59Fff6YrdhMkbezOZdDIFHpXutREjyuowJO2j/8OI4Us9GRlT1QApBQ
fh+f455VfIMcFPGqQu6/Inz4zAdOtHySkZXh5dZZ1zfhm5ZOC7km5lO3RqZUA3BJrEINYs5RDaBu
e0MRBnqgvQ7DQQ7TuTMq9wZ5metFrG79t+EVQupAX2vwhRy05EsBpdYu8DwqHZIcIIMveOsyIVeP
xLk4HlwSeEXEnvlEcymEIK11pP0eqdpmUsaqj3TPLUJvKbYx4Xt4+7NhMnjP+asgUiNyzQ/oWzdT
mgmuqc/Z38X+/apmxKxK8PmJ8njMHsLpU5s60CcOId3i79sDaC+Dak7FFYNX0SUNYpWs4yg+I7a7
ocZww7MvbVwK5LiL93FvMfxKosB4q9LgQi4Ir9le/Xzb/yzM28SL4QE6C7Sl5doi84vc44i9cQdK
wErvG+5W63/DF87bDt9TOXiweiVdWyaKLaDd+uV6Wo5px7BoSY1vgMeUt6IjxAWAa5IYKSewFiXq
6wYwsJkIzasg1eCFu2r3wLaOKQsTy76FYPCFGKgz0WIZQnt7hymVGmfIOSj6z6L5SznNIKG7nOA5
eu3csD15y0G0xHFYC6B6IfEvKWdEvTueh7ttkMqbmrgERgL8Z4FDmyxbHqy/5oU1zx5qaJzunSXS
C6qK+0NJ4S+mOXQtR7KK/nVL5HZ/GrPTlgccytkEIXKRTmtwlnqpJ05jvlqg1LfHtOpotEEQocbW
NF9VgOcdmDO2/5j3jTs7vYS9cn7DxoHYbR9HiOBNuOqWrl9Lxa001n1SVyTKfFeey1cQSMg93jQJ
NhP9cJcxpEQrRm13tQce36dngZ1eeQn+IwCn1CXfGwWceeQjhP5sgg+syxZQ1BhDgjHSbgE4ZL6u
eqE+ZhQ4xPruqClpCIiEVbajIcU181R+hNY0O5Vu1ReN95uRpUW2auszmLKs5dIZ/q0u7rnx3i5A
DRJsdzXKXcwKvIv7iV8k659vWtRz4DTy8KgDtngH8JiakbYm7VSMYXKCzfQ3cvU2pWoVenl/dIs3
s3kBaA/FtIiKmvIYfEmaRHm9F5ZT8iCeAu1Zvbr0AzLCo5u06hUF9ff5XlCRcK7bY9IFWbmfxDdh
7YpxpSJuSobUYBtXRsZvk5fsqnjYNBduTvqQiiL1iH627UFuR6sARI2MgtRblWjr3O4epQMToBUz
UBxJW+QmyKWQBqNlf6ejylrMQsBdjw4zAwYmO+KxAm4Uan53puqcyfjo96H94cOSQuAf63qFU3Lz
4LGibGOPknMOVuJixg1WrZetgpLyYAgE7D0upsL/550t3w5DmI1a3QHSeUecO2PxsEOXtbOnDDmK
ghLws4SCE9ALoQTwlsbi7xIGW4ROyFz2/jRL+Pp1ruVgimNmtBExt8oAInMMAMEl8eYFIC25MjR0
cnvH4CvVXSgReee53/XkxxvBYohhFget9azmvqe55a/u7U7YRdk4PIYB0h+A/QxHgXHoozS7sIPo
dsNr25f/LvpVXgm2+JT/bEHUX9noHl7kaYYJjTzerHUm418ARPmhXxIFWrvOWb5Vd4BMdDMDkixY
ixZiv3cdcWvQrCPTIacHFZXACYt62WLqLJQMOtCKoqo8QIjJFymvYjHBsYo1zgzP6xPott8CeUTI
eE4Z8kZfWsWQPAhDDj+zwpo5VG85Pf9iZMkSqHRLh+J+KYLUjWFwzTmYVydJ8IUhYnvsG1JCo4WI
CjGmIyaP4PTgYI9O+otmCjiAv7b6B9PxIA+kR0qWlXu8fjz9zlcxKEeVrWHDhAUE4z/Rjgbp6Txl
3omb2Ubr6ERp3dq1W+hln46hDiMsdW4QJCq7sXyKo15gD1oX2mSllPNJBlgq+lrQAwskgfzRDnh/
JzxYPG5j7OGDtZqFkH/LTVcrkT8lcFERFTJ3dKllzGpTeCu4KSW6VA7PiIw/9h3j3Bp9mNaLVjjl
itYAXvhg0AfNy+NKhdq40josKQhTMEWtmQH/Qo/bgDKOCpt4xQ6hIf91w9165W58uJ5Sy3d9M8Zi
M+Ffqi6bfiiWdfbP2V2I5cGMZtSgDM6bKzdkAew81hhxVi+m0U5zgrm/zGD9Ar88yIq90ZHqxQ/R
pM1JKQ3nS+U9YJXRJGMjejZ7TTPzFPf49uMu8MB2cNMcsCMDGJikTf7pmwvM9TP1MFZXh2DhHFtO
wLRQwHD4PGPaxR3o+8rkP0MwyUGMkomIjIWPLnlhbbxXzJaXTswNZg8qghoYAfbvsmFvRe/4CaBW
EE0Sje/Ug+TL7oCjQo8XKJO02R+fmotGUpRThFbX4f+7n8maqGnjdMobxfqtJT3ZWSpsCzph0o3s
zPrfASiARd2vOEO4Ewch4JdJBA4jnXuQ350zp4WvlbZikR1JRKWCL4453uCUXr8TCevq7mVgyljw
/U9aaakNWhVrptApbjIYCOpVCDW6bqr+RnzlEThYIsgIptIAIHMu7oCBiOEZI2kxzIvgyzMk8CfK
zZnYvWkYlT7wBWq6putu305gpQEX/2gG9hsXNatoA6eXKP3EmWBbFUuhF7e72sWLJukwO/DwNTID
MwV2N6XCtQljlCCHaIpM6BLBIL7cbtMYuNIt2xLS78HfctMC4vUPmqwgHIcbcDoKdilwrx0hAh8v
O61VuKZLQWSblum+O53a/R9JtCZLRFvfUS8sfeQcCEj/0T+DZLI0mTF9gcgF8Tl9jwnUnPF7B8Uv
ft0qFbLDgcBMQj7rcIWcErmBl3bsw3iXv/6QKYzueiBLLG1tJ+JhR9lrDubSAHCFajFlmsNsGzem
uEi8nHr+//fmORe4tgf5fgBMC4mdRC2WO3f2goNtQA4q3Aod1L8EH3t/4wOSgVC4dlOzA5wm7hOU
Vw/QRUszbuxTDhDPw2lhLoOWHiQlmh0ZOxZ+66cj3vaWwgYf3BbVN537YAySEipWuMlDDgTzf1Ys
caMvyC+ossnAq0hrArbMERuBKI+qvNSq/cvOXinxww5YsxfvGApRMBrpkkGTDUNEKBwT8RObfavm
l8vnsoYiX5YFpc5rYUlkS7fup7bySL1Oljmy7lK8tGFPsgrbwdmVK7T+AUaBge6be9KHvFyTig6h
0gK/JNQkwC7AAoQDaEzPOqd8MDy8ORNjwOuYdTSUGuyhwOyxYlzRTTrd97miZpgD6+YZkeDvs7XY
CsfVSqhexwmp2LZDJOscRA+jex5GWOw6anvL7l6aPe7UdOO0agTiHozBsoSH2/hPHm+eJtJe9zzM
M3H6yWY4Udf0sdktnkCJHvyRsBifjArq2pKXyIu9yhUdzayLPuZQXO6n27oSCFrGWMIxOglTP0an
ls0y/iWSELD3nCE8qbHhFi0qkJvaMPR0E+LH4/viqQT7TQoImybvrlxmpY0Ka534LX7qCiiDzJ/Z
OtndF/D0aQ3gUczbjo3LuJh08L2wWwSlAeiLMMpaMBcHkxoJxb/YwSJvDwOj0gQOzgtbq8Xy37QU
Db40MSB024+lr/3dV3w0ZTg6kOMCLuJoxyB7Zlp/sZMzI/tMy79m9cxMMekAkxRyzCjZAClF43Ke
nTZ1bSGDdR9f25W16GLMxqmkd0VWtuURdImE2QChCEsbsV929APikMX5p+sTKqmFQIUsvjMcSD1y
lFlntSm4Ubg5Pzh39V2ejUeZIv3fvBYbEiO+xLkHGruTvDzs9RZK3aaljAtpAXYfaooajM0k3sqp
qsTxYo3IzLbApWZL/e9hblPjfQ2/mR7GgaXB07Yqnsv25o9tTj6N8x1Baku1occ3If0M6bGYDh3t
5Bbg+0gKaww6shfDnf7Zei4U/3WY5s4Hg1oezivn1IZzZuH2w5dd4Fch/+Kmw7QHK8KE0SW/9a23
6dwQIJUVprpeXWSoRsBYTR/v5X7Ln0FUft5yp9QisWhlNetJoOKs9+TG5uW0+t0/guqhLMOx8qZZ
GZqgtN5IIXYVW15XQRKhFVYBBhCaecR7KaG+WzbtpFEoLVvULtdUnrJsSpgogys+4fC8kM7WatSv
Ly/DOV9P4sgHw6yKCk5fvJpmMBuaKm+vrp54XwvILZhlgczVc4lcw+pciFjO5sruTCcQv59ZpcT3
qjpFRPqYZzZLWMyZAvS4zi+mmBTM2EIE7xnVjqsw8Hsu8newcuod/DdM97AnX6y+THA9sunprqxu
DqNfMX7jqDD/tvB3Q/hGKJPlHjmcEQZwG0Kgtitex8NU18+k5pF7sTMpFoDrf/zQiPXEI3b7MtZU
zF4F7my7787vLoadv8NQolTVAq2/ZPl9kNr2gmnPbLG+pHR+harJz55SrIpn6hpZsCbH/2IUpNKn
0J1fXf+tMGKXEqhe/zO0ih7PV8S5Sq1drtTVLor5xQslSo0oKt9RcgTY5qwSrY8XyKFWGvK7ebim
8Izmsxx8Gq+NLFkb5h9BXSx3S3RYI+zDcak3NzT8vHCSF4DCARcJT+/CH5Eh4gYfxwWdrLXKj26o
mikZv9+wSlGNtczBm8hLN9AzbrhjtN4L1m8DtTOhyryap1jvvQCGE69ewkcx6RVoFkrvnwW0OPd0
97hmqk82qbfNr6BMmBb06q6lWFMa+vyfS67xwCIvzQ5GA6poH6l2SkGK9Mojw1IPq5RtxK2q+1Kc
2NYvqCtDrVZCADL1xSKc+RzE+HxWM+TgDwzsYHh2hgI0VgT5DWj4gz/EP4k6oxbY13zUco6v2tRg
B+iXE+TWJRNbGO1bHyOYepNmzTHEf/72rHKf3K/JHJxSdkqfhHNy0WpkDvSBV/LSpj5G8DIUD+96
X/9G58LuBAvl+uXhOUNjfGGTSHRISCX71rqQE6ytYyywK4aPU5CiE7OqwSxaqiqPn5XsU1VDuq1J
Y4Wuq0vPUo5uY8L2ywD3Tzaz9Di9piw0qFpF9DIGMWpueLg/PTR7fkuFRUqPT9d7ogD35WO+8NKq
LhbR4iApFWa1BnoCJjWSbc8dZur0LfjKnH0dJZ1I6XsddtFr2gEv9IPWDAZveWAsj6nU3kJJBF1K
QQz7Tnq4Jo0xwvbYrA/EQ3DtnSB4U2KwqEbQU1d8TogQXRL+fhMjtHafnQvSKNUh3DWuRt6JYQX1
PpKy0WA+tQ9koHI/bSm4WLoH6a5kyByIqx+tkvFQg3qmXJyf5CHpCzhhDx48yIRAnEGaogOxe1B0
tp42bGHMudrv2nKeR0MYgtzcRTOzbUgdt1IzYG90O5c33+TZUAENmyk5ib89MyPlTFv2kgLbRnOv
qxU044Rof83mKn68QTqrylsKmhWC06FCPx0PhDgykrlZk7ZpLPBGNTbZ7v81bg6U9aeVgIGlCIQC
13KKPmilcLjT8cI9+Km0qsQKNZ45NIJJiW0NnP8RyPGMP/NPg+93qw2mdnfTBA2g3qDCyBEhYmM5
mRek+AW5r7viBTShvGzQMjjVNkbmmqG7VPFoI68/+upz8aYUpxQaKNKX6krsP7jHvlIKANAcokfm
G/ScmC/tBmV5Ie/U443W2j/9CJlFxGAr0cA6W72irqvK4NnDnyzYB4PIajWBUdMDA8zwx7853emo
TachRaCmlkwRmt5MX55zEHNaiRtfw+pRl7LqiS5cgBNYo+gs9b4/yJ90c+lfhYWccI/QJBIz7Qci
CbrcrkwDuqjiohO4SGGyNi88sz8L57F/djXj3ZQm4bhcCf7WepfcYSmr78+ZRsZt7R+Z92xB0AmZ
GwFWcrdLKXVgs0/V4jQSOi29vVEYmT45TZpdT3WkuggyjwhtxgN9WHYRsZQgfXnHdoxo87jzc5Xe
S2n2sN1hJdDk95mOD4GTLSK99Q7k4hMyqJnutjb3QGzhJ2wfONL994vgL+YfD64BZoz3Z82mH+mL
CVgqwr100DiUbxpdggZ//u4dv1Ff59lrLOn7An1L6KcmwazEpcb01JbTOVAJQNin3gRCyXwjXA9B
cIubKIlkZAo3s46UAIAHXmsu88I7/n7NQONi9mMkEilNdZno4MulW/JEZ83zpmLN2uqfxpP/RyEG
Zfs/0h4HWqfP0Yq9cIBo8MFCcV0PBCQdKgQMFdTXxLLJ0FWlh+t7z5dkulqM3jib8qdoayS4WzH/
53XCGbxEJ6Twb4jlMP0JrAOk287/JQ0PpsW9He6xc/zdsJzja7K5IEYFNiLxV6Rn4Y+ilMSt2iaO
EJobX8WpERF5KV572DtUUYkctrsi10wzymzrX6v0GR6agmFGZrFVLzKmHK7lC4+uksbAPECuEkTz
TM1ClKq16pYUIdxZ8U5uzhZLLyuaeY2V/C+0K44+rV4d+1Ev2WZXeVdaxjocTSA7QF1ZsmOz4ocM
kWiF6CJc23IOIt5dU3dqL6T+Z02oRUdfwOTm7N5+V1TGV089g2yjNswohmx0voJxcSZQwSI44oAc
ffMea1MucXVhRCxTCA/ZuIms0MD+laNfBuyZ+8BSakcGF5t1zWhCRpo9AXLGs2H5X+Opvat/mzdO
5I6YPGGgRl8efu2jvmZEzN/MtKHJaLxrrcqDELtGDNYN9kKg1i9MsQyBFzMyLv3KO0VSbeE7jx7Q
/RvQqPen/5XOVoKP7tp3vtWznNilg3ZA/0NSfWAtAeqmsUikzyRhrFbNcGaQ66d0PnpRWMtqrQt4
x9e9Wd31nJtfFmOo9oGP5mWC0ycEIH7BKMVc+kd/VXHsSqoxskFoGqv+l//Uq0eLkxtY+ey6MnB6
dmtKr4rmkF66d/V1AToHNo3GKiE0AvBFVKtnAGspdIHgEVapcvZHxT5fOP6e+OM8WmNGz7FYmLq9
zwETYcIpV/SBbZKjgO4p6hpDUfWD8eT5sx+52PKVeiIMx2C9AWrL3naMDhVnxiWZc9FPJkc3ndST
uzJpZbZiu7nuItnSHtjlBxItX6lprpqGsQzYU7VAFrl4Kz/6XA5l0FBI4bu0/wqwB9QhvHPJtsDY
GY9gQDsHZmnS0sYb88JXTlwWqcrz5BAocgu82Y5H1bd/N/iZET6DaDglLaRnfhB3NhEFhrrH7tI6
xDuGhmGcIKGFFSgbG2FKxxkipBju8Y5oxILCJvItCNQbm65oIgG5JJ4Ic0doo/H/Vetn9QImVXbs
3QxuiDPuHRuSSNN3wFt3AZvZg1WIi22wlr2xH+dYzO2/QID566c20PGu/PFcRedWbmrwHi/p+7ud
DC4ya6WtNRp37T5pI3GUpeZ9ubFzmmPSd7cg9QThTEVuw116c569K4r2EU7N+9+8S/PWpnf03R1f
G2cP7dRqcKXF4pgif9XYIfbgtu3rLgYbHKTpJbW4YqZ3yv8qAfdvUTU6sZouWOD6TbZr0DSpAyqH
TtNXhKfochAT475Ws8M7y5N01fMRJTLnqOs3YLJzHEtBFz8bFpS67jpT0IIsuqPG6r1Sla0XBVLQ
m/V9ZGhrLHOrag+BP4NiOWoIWvKtSduUmwitQLinH7ZVzSxxfpHzBkBzyIO8Cx2Zn9EvTY3n9B3E
mPsde/dkyI5bUbkapePflq01K9sMuebu90O4DACYexu8v7V8JJW2NsPEJQyNCfvIGOu4/nXAoBcE
W3q5IdnTv5b6wVSRF1Gqz7JFbxbJKYJGyRJ3u/jOyUrTHTLiwj+hfLiCoXI7kkJYGlWraXVIOKHz
z+2dqibB218O4qV7UbafPXDF2OVrdv44qR4NqG3BIYF2St7OGtMC3E4mTMh3MoulUvGHClPg7ips
tt/LZaNbl0yJqlg1U26w4DhXk8WRcQvHLzFChz81uYHXCbYwiqYiyCcj/oL5az3V5/cwx/Z3HMAj
L8L5YULGSrVsFyg0gbnhbi2oCVW2ZgctLVgfEU3ouTOIGsdohYYNX1Ek2Eb5aju5Y6og4Vu0bIBN
yMzT79fPAjJq2apYBSxeSbhUMNXjDwNkbKg88GJB1YKdY+jmCiqZyJsAprYn5FpouR4zv+Ms0uOM
GXKqw6D15vSQ4W6v/OLq+ci0FSM+fgJl/P9fN23xlYqYcC8eY1wslBPQoqaMHSAxo5d5FrkYVWcS
IOFDiJtqZxzxekC9azLTE/uRvXXm+Tt4gE10qz5igB8zQ43tfw7wheCmcdGgoKHgH1/ki4HF6nSE
j8JYl4vdFI9+ZHv7dtP5TRVsNLE5oKte3rVTDeU0PkOIRT5rungdbQm6lwKjjlAcG1W2797y5YfU
py3mHJ7DKyw1AJ+7pEp7GbOEiKc2CXjZvMePUlnltQgzv31/LfPSDBQ3FQIyxM2ImnATj3bDTNlB
69cm2O/4D4wrPf1um89deqt7nDzlvTH/RaYyPd2syw+x3NAxgdczlyUjtSYPa3DQzJ3bf114NiCE
QvLGK/V7CJbYXDpV1iacmIG+IBn2zT7g+8knYDztTRExmy32oCQ4DGXS0xoPAXAzGB9K1RGsbkBy
CP4+KE4HHyTMlWRImDeD2LWb3h2tnHgzHjlE6S2RyLf02Huaw36VZrh3ARKHN77xZJUWhleW84YG
Lqi+pj/b3q3gApf1L/mT6b4i5exoZjDDquncZUaeKIhzgzBuBQgYp+DpHdT3KWxTYwfRE4Ww6qyA
IQXw6wXvWztAri5zjHqHQPjgA8+VrwO3b6PpZpBcWpvsmijunUItcUGk1/16GNwh94yi38p5hRxL
YO0fM2I61BVwWavyhmmaicAPM4SGrQDtgnXCN/CgnvXTBSua+Cc8FAI+PiHkDArr5BprAs4pGQKz
bi/DbkHfXxxzi8l4xdKZIU7l/ks0nOLLZAY1tMfI/3/sxlDAVFJmg+ZNyb6MF+hNPyBCxKoetzst
EOGqhLUPSsG5hvWp3oS6JfDYt/UE++dEvxUqP4xqJ9rTv0/YI8rBui5L+dVdQGd5o7jo9K4FEU80
4iuqOqBx4OuczbhpfqYL9J+ySWuAekToz4SH2L+bPeV3XM0PCfxR1YQwP9fZbbSe5BLJPbhVfer4
RqDLcgZi4pwSMX/FOq+HTthBbIXAepw1LoJiUVj38uCd2iHkQ+r0U10zjbhYoChGwGvCl9na2ySa
eUhhZylk3YoTEb4eLgB1M7qHDZr2+YMPahqOaoZZDRKGcrYVG2QWIg8QYr327piHep9k4uHwuWS9
ME6kfSHiR3qUTL/pS5yiXcomLGhJCRIuOz8eqw4ejhYlVg1U2XvOfZPVh2Z3vdO1IkmYcjJh3MwS
KQz3KUmtQFdR2+8EJ5N2RI9AKZCKJTlxwbL08bnVFU7y3IjjeX8CIIOfaGevnpC/x9eXUM7G7wEO
zfcJFyCdha/ctKKySdzeeaAjlJXjj4RzhztxNH+xMpoXypZY5q5uwvxASU2MNhvCjcpSvWVUSTCK
pmvAz3ceX1IaOJCuKzAxNYBduWBySq+GRBl2axcMU9QfP9IHsn3dw5+C43iSfTD/YJYJu91uYv8p
tfrR1vbrOZbUk3Rm2/cQaNLD7yR6Tv2E/Cn4w7vxv32EiofoOpnEFbsOrwRC1FRpaZY1QEKdgo1g
D4WKnSe7jBQScTBxku4bOACvypMMNRI1Et7DK9V06KTfSV28o0FjWUOzSUb5X6tWql5KAkmlmCh/
UbQMISo/V47af1x5AfNhn+6YQPe7gPg+vJKcWZdE2IvEmOX01+P7OD0WDQO5nwPyOwylK0LrLwkm
62xwI9KUI0m74iYY+9Y4jbjCj+7NVoLmakJKaLkoLx0DZUi1Ke1qAiB/JA6RVg1GV3wmJC3LfaVQ
OBCjs1grX0P4wIsFFFY0veFbM+FF6pFDxTVcbSEi2PkQi5lBuarJ5T320XZU3D7kI8bnGkb+a0k/
Uk8g6GnDiFJXBxvxdykHQNNO7/6tvyN79CAhQ80S5Q2ZSsdzel/6keQvrczNy6TnQSjjAPlBKKA0
4iYYQq3J+vv0zfa7dTH6QzDvPPVee9kK05FbbQulWX2E/BPOhDtJPeajmsBUYDvK0Z74XJe1xM9v
TVl6hvZwEliF6J1haLCDryNUCGnVEiUPTdB/c5TwU46/WMFD7ObqxM61Kmolh+LwQSWfABadynT2
IsaGlrPRuOTwPbPvZbksVRwntqsP/jrFyRWAT51MvkOl5nD1iHbYpzfxUooI6ozh2/FvyAX4ppLS
kDSl4Yy3/kt0hUlGB+fNWaZqnzIsIcvCnxQLIwtkLbVd5xKFvm/GnF4hu9V+IHtjIlnxkFuH3I01
KsTjiqf4btFauYsgNq6P381J7bpyE15j0efD6dgLJH/D5FshocvpLBUnH24oEuSGKYr2AKwhM6zL
pTC0xfEPzwXkRJMf35vbsN5pz7L7gLY30ILe4zIDa990mdwtG6oHE1yEv1Xod0kj7rOgyutHFg+7
Rdt4S3WMiIqNZg4gYAooNLkKlim9b5jzBuOa2Q9dK5/9M7kld0QoRtH8QQYX9XliRjGUrdaKgQYU
6aKGBtK5JAp9K598ATsMphcVPhDdf9f1aK3N885Wn0eepipwUmZ2zDtR4snVLlGN3zbLKjqlrDfW
cu0QPX/0mCxwOcrRiuseWuUTmT9X7BdueNw+dPl4gyVwqGAlKf/41YekUrfXxLVGJfTPb2nmezdT
sPYkFqHXQQGirXECro86r4SW4eaFuXyBQyQXWJ9JWSV1kni0SCHAc+mRuINaV2QpeDNQen3h3SZt
8mfzt448HYNRUTyevFvEeFcK/bS/B+6WVNhSJm0TDxiSYI0vzUeNz1A3qCr92QBIlgMp6GgW8cuE
rfp2JOzCTmrJz4QB7G8hpIctmAGwnaw6fS69iyYP5HGC+rgyjfB9+N6kv5wQJvZ+T41tl0zso3Cp
MiDIKJdOFutw6MBZMPI0Q6qAyirW0wJ87YowziLTQh0F5MAVTL0PCPTpw1ctIQ55UXan5zmR3juH
9z6mM7QsntSSZb9peQ09SeThQOEgrQX0auh1cBmmgvy3jud1A893ESgRQ9JvW5Z9pv6ksra/uiPV
v+PdGasiE1e/93Ehjt//OVSlVnb9GZ6W+2ZI1byeyuhfjWddQoI7P6ecqEA/R3na4zFZBZkxI5fv
Dd1beiIyfYIHjxHZV2xy/KAFn7QZYrOCVg2S/bk90uf0DVIFyVCKh0FgtqBgNj2VuXm80q3DTy+L
mVKnAzU8X+d39pNGqwjAG3kSDrAKtljhlrDkxJC3k+Yw0i1hTcyn3bOh4i4gG/bjGL9JV6QGrJ2u
PIi+GcmR6UPq36RVkVanr7pIVNJ2q6PlqZOb1KxDkxF3PuO6x82Ts0xt0/MJo2Zdl4BLbyfhpKJU
FoRfmSttHU3rkFHzTTQ36oPsI7Oxq31mdw3yuJSXxlaL2QTLT8FKYEp+2lqwnHD8E1qzkM0K8N5j
j1NWVAyFrAxhEqJWEje+plPXvPeKc4xCLI1LgiJ41HwgukTTETT8wk9Xc580L64F4ZFg9OzYLQQO
zdbRA7FIs9B5a8Ar6Z40WjUpTT3T2GHdJmFgtf/bdY8+Kt3ea+RJBj8pgjaeMzxfzSkCuz+AfBtD
RE4Zc+v4TeWUbi3cjlC21O6Tx9D6xTCCvvjF0Hhq6HQPUn4BebLMyQpPoReB0Rjxe5MbMKWk/zb9
i6c3jEPjklRfjvKYTGazRVKGOEFR7n3UKdOtSuRTXjp+bCsWAsra3K/65WfbkbxSkfoNACAEpAWI
kjQSswGddDrrSXdyy2fKuHccpRsLPjLh4fMXa0J0jclk/pHHiDZ3N+Qe4z6Ks/av6adRTvJxW8LD
VZXsb/YfoJwP8N50LTNqxljZy1JGJEfC19z7Bt9soGHpvmOVyYWrXB/AOeqYRNdMuTwUxlNs8TfL
hkGHN9zoCxcSpUeTxeSW1+OJ5I4Y5AkRiFPDnxhojyKMAtbqjsB2iWfycZ/Dd7GyaPok6K8utW+E
+hJbNWnATw==
`protect end_protected

