

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DIIXDeJza+sKqBrj4qf+gSpQ5HFYwUFgPgXoi9a/661p1fOh7GC1Yxr4QhwzfxxbI2esRkgX+RWV
O70wuqmd6g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tc3vvZL4Z4/k9lIOYWoeVvOilMT9DFpT/2Qg9j3BlHsCcWm3A3qs8Rzy60Chth5nEU3HV6KUki6A
hRQKZNb1v/6vjwTmXalrXjELjcws7f/IYaWgZmjVdYjpJE/aoPqNISqRAxye6F73bRYmttkSLsKA
mpZhym45OoX2lTi2dYU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qQBOLNsTpDaTilOll0jbdzN9+CFe+2YuHpSZBsocYQBx4tFyydxFP4QWzsgkpKMVj+vgHsshU0FN
Wu3IvX6zwtMbic8Oj5a78zbLuCwQAJkzJHVEC33oza9R+KKTeRuoZulmj32txP8npOqkH//3iN6m
rbkJ5ZuVWuWTahdk1WIS1WH0JMwmkoMmZOzkIvY3OwyRzQ7J4JWsuGgUCQP2UiR1wTcS23zdZ4if
K5dX89DOQ5XLDZRfGBzqloRoc2KLKrNKj69bM6afBdivLgfZpIq8pSaRYrb4D4nQ/NQLMqKVQM7g
UtRkTmmMOH9irg/EZkbw+ma+qT3UysisXvIRjQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FnYKQSPwFxsA2Tic0BZESWi6Be2FIedgCX7009o+DpIyXr2I2/Jxc6RNA88ViWghN3LxaxRvHMEk
pR+MRZPIxTWv8WVlO2x5IF03WAJs9GAB6d9KbRe6Gs/fOQS8fMMkXpyEq4+6dsQ1yT9ckah4Cdmr
T2dV46kU3DtfOZwlWxk0OFzQSvWXEIETRCvrsGEf/mlDvxo3c99T8p2n/HDBiBrHIY+98bbLLHvl
mVYYFNZpsys4uRT/TVeQxVr2Ro29URGWoe0peT9xCIdU44Br4X8OPNWGJlsWrkooLMv9dYIUEfQK
VsblVGzcgvRtwlSZRK4G7ikWOKojLVBxgIsuhw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
k/CEKtjJXdiEV2H3DdiRA6UDxaoZt303yi4S31RTSRFiDtNKXEWX7hAbczUxcDYrAZq9Pa18y/Iv
ju3h9ViJ/yaF+1n8xAYTxusQZdevYvn8leKkc+XbCxi8/TAYj4SQ2bTf4RMijly6zLqqO004hHo9
AbWF/Tq5CZLrvf24Df0yyJWZTL2km1BM5nTE6v8B0iMxEncPNncJ1g0VKySbcBDCh6+IdZeFDvjk
siaQTjWx1gj+MKrM5hxCdh1gK5aVhC9As2wDY0avEH+1IxuO6QhBjnWFKX5v8fUQvgp5zjSufCpK
Ff3Ce0pbO40TcP98XMg/XiCNI+dX7w8S194wMw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B0pRxV4llSbxSsgbT9dwcuzImsNM7Ywl/K0BGEC/Mw/vBjKJqOpZbs/20GVssjsAwFuJAwsuRvU2
DcscqGBWo/UUVxZ1dW+/mhv8EMGY/gglmOl/jSYwQ7g7m4z3an+lZM1T9/p423pPW8FVM8MYisbM
+tyxyBR/MgTmoxWxnA0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EHRObHCL8AfvkiomPbt7c3iNsMF4eZGxQ33JWJrsuaoV9trVmGm8vEcVPWLNhGAeekB73BJR+LiZ
zi9a08JnSoTsgO+46uuuGrEM1IK8husQ9MqNyNGRTbups69htwaKPx1YLtc1M/60smF/b6euaSYM
JSASlMnD29rew98IbsycQiGsHKlati+Itr7j9mPAlgM09poau5yONp8Qnq4dT11PG2FAMF9RKNCl
UCdKh8nmXtEmrpJH+V95f0ogErBgKxxAVi55Yvtg8bgVdXD9OE1BJxHTIDLs/OWMstM7CzQdhFwf
ujlmDvylJDwTSbP429MwLLobIYUiMwfATB7Cqg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506800)
`protect data_block
TJ9aEWUN0Gl+GXys+91LM7Cj8b2StXrCqAZA7YqTq0igFESH5cKz5Xdg8gFK61+kZg2HEGW3QS3D
1yfuHEjS7i0/oPq0rCRU9wQyt8umkubCSKwStphagVVy0MEwn7nomIv1SJGRzFglViLrrTKneFGO
bFVK1zXLq2ujCcLdkPbPpuSEp7QSY2YMhQPL8alf1Is3LEE7+cZ5HlTmaSvsOIqfG5MpvktHs45K
eh0GO1/r82XMX9hKnGbz6+UijWMshYRPXbce1Hru34pyKs7Kn1/ELx6/IpMoXfY9aU1we/3Q96iN
S1KMsEJkqQfZqByLQO8/eUddjdwQBO8xF/asAnJf967czdg4ZaVbZKms6V9+AlLLQ5k1wo8LPR1B
zwkqYVSnFA5RKdUhXR3W+0kOc2d37zSYHGQHA5hgHehm9+PxlBcT4ehtu9MhWhNoJH9PjyVta2UW
K/EnPI2tBIj6QqR1sZ7k2VNRX3IM/P65SulGfsdvWLKvv5yZYYhpo1D9bzqgt0CGwCUg6Rr5p9jr
wcLr+HLFDHT4ZQecJpGS3Tos2cGycAAV37/EaHvma92IYjNbC7FR2Amsgspj072phEdZ4Nt5vCSp
FE4Rb7cqNjxSQtrUbmGQAHmnU2rjqGMDL26pbQFFHPbK5gM5IfjUpR7TyXchwlBEJ/zyMzdtlrs/
Aezyvl+57INmuFJuHuCZKtSSkiRTqQ4w6fKzkqxQjo9PRCEXbZGQpDrIfHsIbgzA48RWK5wB63M6
beKPl37uL0b8XZbLx1fVLhGQPDkaAaLRH0eiK3wySlLT3iyB5VeXLBeDFAD6AFCD8ZgPu6Wt+54s
VdU7sulBRC71g2rC/aWKlQXrXNGI8mYdx4Q3cAUsnFaFqgmk6BRYdxHG0jae54NI37BVoTvgUtQ+
tt1vf/OI3w9YhG96Q78cFqrtWQbjrXW7qKxoQQU+pBjtCPubENJc3V/oe4Fdtdfye6xTvCjrBjIa
yRb9np22fv7iWaZQtWqnXZbjmgWPP2+ygfZjqS+fWS4ciTmdeoAthQB4ITW1WRa5tmfbRKJDGnfN
o0/Mn25yzcs2rtB0aBQjCK2XFa9+BKJl6x6nC9D8EihvlRewPDtBdl4wiD/KHmAXMHp+FT/cnNbN
qbWTlfV/NK3UNlUykmHP1p6ccGkLoH9xUbtJnVnFGvxCkJxOC348jXZXe+q2YDw2T9bSS9miJY+J
fckNiGuNhhkyD9fXFUG2DesnLSRAHc+m2GRK4pV9W0Vu8z1yhzhgR+WMCbGM4Eamq9JLL6LgcVrX
iIn5t5z1FweiXIJMVr+W96KLpsevuWKl+lyvIz0AHHAle23YFjacNAHA7y0eq47dZbM7lfqVpw5/
wz0Q/4U6gGpF/kTEPjjZ2cxVKKJr5C30mcQkwDRGk/dPqj8d+W5oTIgsJX2YhTMCm0QWGiff5u8R
M/n3C8PDVpc/dOck4qVbQzKTfB5x6rcU7MOAOc6orAn8Do2bzn7tystZC/V7jC3e0IjW5VevcmsR
4X2y1KHWco7Tp0tVpMHK43E7v80kvU5LzYOvl598H57x/xdw7B+/fzhLjiZexmmEuYoePJpFJ8oY
9DEAiTMK5MRyivtY55VjRBBUPLjkb0DnMDacgS9KX4RXM+6wBreHXuQDEK5rcPfsUBXIuHvWtiPR
VQp5lTwnL370u/V6O6k36xLgBrMjh85/Sv0RaPmd8+jwJ08GjO8Lna7RsH4apdnb5/4vfH6pbUS0
7t0ffi/KLUH7mzlZYhRAGgWDYFwE6WBdm6Exc7OW0xHl20fzwtC8ZP8PRfkhEVUEAA4SkOJpNcXE
d/77ljgUxkV7yk2GNmr/L7tcEs+r7QD5sQ4QEBt0MJDRO1h68vARCHSZcIywrwx6c2jv5VKB28nh
Hb5yB4It72LW5h6qleo7iIOJd1O2X5Q9ogEmjwnpeIf+Wi5KgzA07XzftfCzdxs26UaMnqsrH/H1
jI0aGNU8tgNCQD1o1o2Kqo+fXJfiohOocukEZlPe/iMdvhjHu8VkwGm1FrYFvNXnJmy2KDvt3yb9
/R9esabl/Nr+Qwf3vIxJVw/yKaIwiM5cG8qUFOFmZBi3ABanq9FBM4fsZIvvnobNFII8n44WW2j+
XPvbn5dYhAZBHiZvBNtlNECthiLexArnHXmTkTqu7OD2/p9nnvYnqdlGVY3QyMgoaFgakPpPdXIi
Sb6jY+s2O+Q4YtAOfP5F8PHyO2+NuJ/EYZ6eMla5AXd9Pp5xUTCi1uKkYcXlX7+f8USdEEJsOsrj
Z9VkIk5QUN5xJNtHa2WxgfQ4/GhcwnxD4NGOpVcrrxqSSBvLx7yojLE+huuBXcEjaspJUKsU5ddQ
eXB+WbvzErtQxXMxI+2mpcqPinqSk026ENTn/vcEJ+Km4vEDqM3paAKVVs1tLbJMuGU8Bf/qN1/O
qYV8HO+ScXymwzEYXQZqB8ijUjOV6qeL6Sgilknzd8Dp7+irjFmK1I7ig9Nq0PeaLxAUgoAwvGCQ
2vT0nu5ZvHK5r98yi36o3EuK8oKaskqk91D83TUuaDDnqpOTtTgg1zg4xH4Aw7Tp5a453quuev8O
SdAuKdG/w+sn4dEIeQGHMQwYRu4wyuVeyJ8gmgxY2CDW93qIvykmoDE7EZ+hipMJMqS6eNkGArgp
acGATx7YYMOc33hmNiNkmYcXWH7aZvkfi+rzCwRBXboU1qegjpD3DP58Bs76g5LxjeQbDWlDMd/l
tplclNv8nOOqDwLYbJ3D7mYR+cbpTP9i0Vj6OXblanmneJo133lI1I1B/X5cqATmTbZkbJTC3U+B
T10i97ea03EmoxL6HtJ9Xt/d8wdt/mvDK+DgQhcPVovhpce8iPx51jktjZLngvE97s4YDm+Z/89Q
Oxj3w1i8N/Zvbv4QIgTWVk3ipg0DAxf7clYBLpeBom5Psvfz5Io+Hktc3f5CvuP5GOqjeM+Zqj+n
OmsX3loCyb4nv3GGWl4moW8Sq0EPl5ZQzI+9x/6F2ZAdSm1X4NwILjf9/tsU40NngNTFH0A+ksKV
OQ23kJSyzvkhUFlTOy77ejvOYNT3FSxmLdmLZ1NULzDZj+EGnaimby+wTHfyg1vMdqHVn2bfPbqt
LOLnwVwBL7g5pmhwLnqZGmk8w066S4c9OTPmQM8fMegbVHilsUio7nglkN9ylKm+k95rUtYs33yF
4iVy28iHiFCkPN3XYQsKSHa594C85suQhHTv+g584iwW7COZb01nLODas35tqsmLQxPIbmtkzOOE
pvATg3gFy7VesJNknbIVM1R4mOwCslN7KCIUYxiWLpC1hiIRmZ5mo6tazEjNaukmvsGuC5DCdFQA
4ht9a9lvP4hxDkASMj3dIJU6P1+gemLMyHhK9zX1VJqFUuy1JNknAvNnG4+n4Q/QXiKSSsKc7gTu
160Ps69NlG0wZYOGMxagPNVTDz6MuENkeixuYvcRzd/szbZTa+bNh3RI9tg5+utTf9pFf9S4E3c2
uh1gRk4qnCH6o/KVL+bVgpcLAikYjo0/TtFUVgKdCkgDgOKfzUyWg+Kqw+NVsrSgGOschy3XhNiS
Ae9WphrJfhYAIZGL9TZHgVEUefuLrmXqeejzNX6PuEfBv5Lu+SFyaJo1hfkHPNwyKHeDOA0d7UDB
noJSHPswTvp+g4zUVZ4cgrbQSraPujC9fdYnFcBrkr66/js5m0Fio+Mr69JvFR3necEcgrXdgyHY
qi+wkw7jPbs+wsdA6/66NYxVLKhd07KNedQCv0NCRZHiwNwQrqJ2RtqFQGsRLNEwPYpM3oxFjIq/
RLCXM32mV5Cr5HwdC8qBnY4Y2hgRAcMXm63NSL0Ryp6JmwLOnxse+XSvZDHfd1d/Ao0IdPy8oB+Q
KZTGYYQ+tRuY97+5oyyEALtGSi2SrNph/qztevQ+NjYw9uyUesaCBvjre4C2kKDdK/cDXFFL37+U
I3Zp2t2x/unzxoy47aoGvKqTssBo8eykGiu5s6MFX8pmuRppAeZW1QPztmTyK22Lr4r6R4rfH0n/
Mb6MROLdVyJES6gzP1zxQkrz3fuDJXx+22JCc8J97imqVOoyoKgABrhuooMDJWzpWzp7DHCH5JNm
CefEsP6IA1dZqHDajHB6Lg0nwwGThBEmCguZPQy37lmqvx/U33g66L2BVBC9EG4aOLzuHZikAlGP
5BmWOl0aO5t+f6463U4qSs37054Q9qBqXv/k4jlTJdNXx28GHsCFDjGzilXs/wiSssrZhvbVlzNr
zaD1YlGVcbD2XGFjT3iF1HX1IZWoUQ1/22DNvy3eXzVckbDQ2wuRlWNxlYlHIa/qIeL/g2DCJc/A
i+zwGlYrp8eFaKrdFgUCEE72ykXoi8iAbvT+RoxFQmpRMDh0Owz07IBa7TQtFutBrwIluSMSTF9v
Mfeptx0gqq7w7haTiHnx81SRW1hKhDFlSHlHKWTHDi1eRmZcyZT/X4cG45N7f4jVegHWAdlcdz+u
9on/bIqL3QsoOpED5Us06G0c3tlvjlT1LXAiNgGlLL8OCdCovbt+vW1STvJCM00wvla1V+yzLymI
ovlbVRmGsimOofcG+XCA0CU5vNBnSN2i/z+0tJe7VDIK3qiQR/KKI4B1cgjULGwXb00BIWutSBIT
gzfaoExY5revLfY+WfkaSj+6mlNrFtOpE6neO7jqfZljEfvIm+aAtj6OWrvHc4ayALlqr3h0ct0B
g/pqYrRPFpUNcn4WegB4g3gFpqE56rl8g1Ps1OGFdxMImHUHUQd2PeYAnXRP12+6HY70ZDxOUjql
9pjSnqasZHk1aSv1PfG/YTrATCmpNfZrUxYfTzI04cFOyUXMAgOZzgGw9JPL8mrZX0G1k4QtORsW
UI38HWq1EDTrae7C/FLADKyDcGoROWRQIvJDdN2Nn8jsZzc6u2LGBGsNzQTy64Er4kPimURUSc7u
246y0Iw1ZKgpk+kfzma6nUVcZ7QhWRF0jI08d22Nayw2DkCbxm99wzF12KSewCGdemoMTzpDy0a/
LkB4g1WvPdAbezM+Dx7ISCGc1dArCxXWEea8YKcU3BpSg10/nkY8UaTCtl0I5/9RfPKUHSfNupRU
iEWG09u9cyZGx59DcUn6y+aD7Ne+Ki5gcVkaFCJOfS/z5dz9eMcpY36uh9VdzuAvzWKdrd/NRVzk
g3UV4NQws38cHEY1Drc9QAPEunwFk2m0JNBXGfZVb9DHtFopD+lxbrXgUapJfpZN9mZBcEHbzB8o
DAeeqaUewHXedEYTAqXVGNIANzGUuA196Cv08VUX/euuIX73oqRFlx8JWbdy3LD9lne0Uz3DNRH8
i2V/DQhWSbrvDNqOoNXe2QzOWr+s3zROo5UrJTWGI/83vYxz2wlbKj/hvLKpewjhwjyAFIntAvlI
z1UPDoejWn9v95Ab3+zxFgfzByTKXUZ0pmyA2EMdanr2CHoxy18Z6hyx4b5XNGW01WZP4NO4j3ro
Rv7/6JVQ5X0yi+4vAFgrbywnNYuJvrWBHAdWWx3ofUzYCVQFDdGeWssdpqoZDAt0/ao1tNfntfyj
RzTnQ2h1yoQaVMZEl+S0oAF1wOS+NfvbfpmkI2bb6v05zmuaLRMnh39XsqoGTc/QVxk7Yx/q2Mlh
KRJYYbOl5aLx31gJBjmifUNC8kHSP9ChmZ92cH96B7sa/2AeRO4Bg1Z9XBL+xrUI//i7C6AGevTK
FwmWFh6mbXnrdouRMJvC01E6cRR3r0harUHCuVGb8jAc7kBBVJaI+ukWCCVB7EzIWv7KIGXH/1/y
XgtJGO4MmDwW8pBGqlobIVfbnxOelgj+wG80pIHf1ECrGkj6iT8jTYTCNUm75AcdGJENQnTQaMHm
yd1CI3Jly8u3B+8/5hXNHeQoiDoWAma8PUqZMVxuxx2B5RyROT6i6RRO90lnqijon+Fj77rshpxJ
6ICb8UMbMEMqjoYB+K/3y6x62IUeCWchKf6jSDlYVrkBEvg+ngyQEETiNRb5scYqfYyYq82McGHc
HWzVw45CZTeaqhdFzstLapGKX6TeKn1v4LS+RBo89QRyx3uo4X2Cr3Lf8hEZb0oCBj34SGch0Bnc
56hxT9T8/nFWNAGAwfwUUnlbeGV3ANXDLCsYRsW0ZXv6VIg+X4LqxKvtSQWT2nr6mzW5BzRfvY9U
S6wqe55yrqovxm4YJrNR59j+z31wDQ7BSOe9J8kEJZyNJAqNSTaIBR7MVQyru5AANCxzHytejEVN
0vm/EEN7XUFNd+8e2tftmvH8jPT0owd9zLq6NjVQEAYdkdhdH7P/TTVUydNt/VyDWShdzWnRPS2N
Kp9QII3SE2zWjVijfb53//qhihkEkiIY8QFsSw3h9w5otMgUpnH2LBaxahupXVfJFomLYiYwPf9Y
a5MZTTMruR2Idk50FC0HkZ63VBGJdHnUAjPGkJvaNjbj7oXT1nMKi8OClhpjLt54vnEkJklSKmrZ
TK7x2Vp7thIh+PqIRE0UoSjVfE31J7RgDx9cWLGClhGrjGMIPEfTDlVTZDDLzg9H4ns67eqToQ4k
6GceF1hVy1N/TRo3E7xJ4yiHDA4s6Tm06AL2pv7EdsyHR2FrJKf5hi4Zmk68ZUHK5ICHnho+AYXW
KNplGGL8dVTz6+EC4TTPWq9KAJ+xbxA/eNDnCIVlBY1v8AOooIXmP+rXWiI/Zj+XthA6ghqSd1UD
CPZEX2fp93dpRQKmRlbbM0D4RGANh9SSYQmPBn8CeAl0fMQDeZvy2pEVUKQVSCClNakBsg42nf66
ZUap8PacosgxagGdnQhZbNlwEWgbKWv6C43v72ePEde4wmTuQ94dRfzTlxu9gbUlpuSS7HRO95ii
E8C7WioLwftH4wWaJ/wNJuDs/6zwi4/RJJSAGDXwpp47wYbAoyEJqE2k0MrxEmDeaqy2jO9Lrn7Q
zkg/a6GLQki3KOkHCR+NIqXMlki1OoFHjAaEGixac+zV3bevmX5DpiSTqQ5Rj8A16gk/XdS1xvyV
tdC6f+lglrSGqg/yccn5UOhn1cWzj7ARWPJENfADZ7zIT5FIVRPQcF7eX5vxilruGu2KNe1iaX2a
mHQDq/eopl6P1UaWzelwSPz95K4JHv1SbxCNTRVZGghp5O0QNCsMv7twsjAl7j9oHjJvlwa2OWaW
WVVqzNXG58RagG6AC0NR4K7KSDg5BJRvjmPeJLzmRbCdtlVp0ipOttnwAnzafrkh/QztWqT01q3+
SHyLQ/NVXuK0cD4jWtrP6V/g8+ofkRRhmZoTllXNojw6L3XL42xzp7h/qV6xf49bmf4vTHIglvrA
/UEPjidp7ASzuVx2x43OncT6d7RF9HZ6egJXOI7/GZTwx9ARuTupQ0aXg6w3cmmkAX2Jr5wxQPll
3ftsTE0w1tfiTpBIsCRPVWYuqDbJdNFVUNOg6Ecs8XdoRLq86uGTX66pLxTU45eooo/eH99jteNP
QOWUq+S4/B31p+UCCmXTvzn00ypSitj9S//IrROfq6ofl/GzPYS9lsAQSjvmK/8HlsrQvNuJ2MUw
OCCOsckOZd3RoidqAxDxpiTNEBdS6rmMrd4QINL+IB20MphSbU6nfWkQ4nkggbX/0rSB5Qj26RBt
5cQN03sAsDAcNv0zNAAO0yCrgo8xqpmlJuNnCqP1luLyC8/2V8ollu5+G6HIeOfGTwDxM8eqrbsg
exumN9oDAckr0lqUAdB7ACAW4qNOy/pEnSXPkz7+6PBQYftbzKshRvQAdQjKONFpIEoksORd8T2V
fUrCybPElmIiBb/a3MYyni1cGkkmACynIXY3jGmTsZSOdO70RwM0lxCGpJPX9CpKF9dBnQOOHtas
RFMYImbGlr5Q9Gk5gsGbupBt9lOsL95dn95F+yDLC9xldHhuWLbPIBwx1pg2aUJNki2JSuPGHqTn
Jji7gY8WoDxMjUhjU338pVHc7kGVQsMgVKzOOIoUTOLbSpNJ58kQ4bZgLHHOFNj1Ylda+lQk+E+3
T2RMSgQkYfjHxFw5v6MOAXfdKyO+lFPrvhMkXXeAi0rNB0b/cVhhkitnBpPrtwtiZ6qR0jvFrsBH
GzQMKuysbxv9hpm1FxWAzRZt4WlaDvAqG0gXG7P1eEMSRY67qTFHjcJE2I7dnYXnfJv4jen+D6Qn
7r2ivTX8zxaLZU8sGZgNqG2wYcoWHPGWhkagipc45u6fVOYIj2+S5TSNSwqRV5fvIEwsgc201WPk
9G69WKiWggnpYXDj5+w37xoDcsvZMJqKANhrD6LPFqkg/XmQvSmUJ0QrAhadJZBZvtEC5Qmn2I9R
uptkjwh3YzSdoExkesPVqIJE74ZEI92Ue22LilhaMI6bfkHQKUkM2zin79AI3eSDwgFp2BZ3N9rd
/q+Pq0pB2n3j8sl8nGCL/02cc0mBDYYJK2OG3A5D7hLyNA0IBpLC711wcg5gvjncbOJWdGNzZmbV
xwmy7kxJ1qBrq5une6s+z2Vqzh6X/zOQzr5ek/BxY2Q35jv6XGwbF4xyo2Ws5CxeyJgDykXYvNty
o9l4pJS+fEZHevrUORk8LGDq2MGRCByhWDEAj0rSMdPGmPxXWi6PJRjhFGRMhEfQ6EnSvln+Fu/X
lnHPvuwPir/5wTVn65SjQWmF9gaXMBHsVwJ0kawUU1UeGc3G8Mz/+pMtNiMKSNDsLoch+4xFeIhf
6svnZ+zL+iHGuORr4YLluncrP1ap3PyQ43XujB32iODRtcvJlzJvaIx6GG9EYWomT4KnFWm4WY2G
AZW53EqIEn9A8eFQwSvCAq+LZUdtnpU5dcoNdzFL6gwhRqtKpjiJi+2iklCTecomPrlrFERAteM2
kTtFIgujtAkMSncnAAJR6HEO0Cr34fD10k/xZoB0eDkiitEyWcLhjm90h8fJNnhwmFQLRuBvZLQi
PwNVR7AS/0GgO0Q3TgUlE5LMey6Nbd8aiLv9Zwo4wd3Qabk41E0p6JmY1C5TM+g/7Pa4zyCqjvr5
/tnNp/Rtn3JaljfAujC9VvTLT8GsvH+ZEVNyptcZUElzRWANlDTJ7e7Sv4YDr8iSBhQ/9CnjMbT7
H2PVjPhsPcn+jhQWQTXCumwKNdz0cHIYfGqfBJrUgLlS/SqfV5p8L2vWnvL/THQ6OvGqy+xxyKND
0xMNyjEGjau/ecmGXiu+yJCrKUmBbVMhf3n9GVFNvrRbd2OCup4TVLOC8rE5znQN0hxIPGezokFU
a/QADlzqoTLptL1qtqRU9fFw7DpkdZ+F0zQCWNSCUUtBkKqDuc7ji9LrIMGvo2IlTJRyYz1+TH0Y
+TDuPa9ooESboDBtxPzFTTPr5ltWNVPC66DoVFWj/4LTwPLjlNl7Bph4ibewc6eypDCBlPcEFOFp
IgsXoli85wtHrSyqx+JTop0pveq3a+mmPAUzvQLSqETdzVw2dc3CIAxHBm5+9XF+rpoBRLjEle64
XoMg6LLBM7cPKOEwVkKinxZiUos9iqf+yCY9uiGFKujiJZqCBHxotTY5N6hhP5T7v+KIkgB3Sqv1
GgRhgWVT1bXz4hvk7dmn690EHSHrJNngfnbsQr4miP1sd6x6eEHSnEL5lYcYOzg50u16EhPFxtps
G5eQ4t1a2B6qzxonzb11U/M2Sh6epn2tL5S5AnEidwcbJ+fFVMQ86lIRhynRV62HSv1tPZm3Wgva
+mw0Yu+cIFw7L4zP6an7Ovw42Z0ZSEJDqPVQsy2oJXgq2lZ8fsUc5WCLPOvruIKLsJfetvpmM72i
z6nwZppHZnfFVdKg9lzaIpzs7vtuVDb6eTlue7uA17XwFFuPfI0s8jN8JpIKJW9HHqNTlsRK1Dll
ot1j49zZxU/DlYFe+8Nh17x0ONoYjKUtj7RWEJeD2BDdRfPuOwkVXQDZk4KiHIXmB4AgzmljSYfY
I49Bnh0cOT3A9C6xjRxVZDWYQasR4t5yWj4I8c/Fgf1szHVTG+EKnE5w8+6KU3jdVHapm2uvFtrJ
dKecYpDjARbN8djgyG6ZTPbqzJd7HFa8zJ1ERVhq5irudWCFmCpsZxr6JgEm3wR+dkHu7rTtCIbR
TTgJgUeiOhmQtvsVNpPcMBdWsqtncODk3sVp/95mO+7NWBPN4IHRBTlYFa9VdrkuEqKxbOT5FlPK
/APja4m5l+W5vM0pPMjyomKBA8GgUh+sPYeUpEjRZfhtJguoAtpZqmDDDUbJaD0+IqLTErxrRJZ0
ahwgcmjDAh1YkCW+WAcw0TZAFpjIgzv3o3COnShJBAYT+l44WoahO9xx5HqVKZHDtyhKG6GV6rwL
6mpGQuTvd5wBTahsGR7HSWUcYTh+mPKgU58ARXQSsU7DqtJj0Vg7D4oIXf8USAlshLY9/qw+SxLf
HCwQaKnGwNhNssJpf5M00OtsRlVdoj4f8pB5ZWCAvIFxYHSLMQUjn8VaNzSHWO9iv31qcobeJF0v
cuMkDN5Tm1vSvSWLdVvfDa0g5nJjA2LAwbN8M/dDYM1VcN+XbaypuD/ubWL3V9wvHBkg07QvRjBj
CFPvXk0FOWG+dUbuaZT5LU7CKcu2EDLlRMXz2j+HjQy55Ts2BdN/lT2B9/Rbie6rRlC0VTPPaMM0
s8iZvzFIGPsCJuvF3AO0DkaOiwqeIzz6YEeFR73JEN+47VGMsNXB3tPIgPuGTP7/pDq3O08jN9Yv
RSVkovatzorVDjSfs23Ak56IJfaaGfBEKadPXHXiW8TAC6eeFELdfZ8+LarRyrY5NCGlscPDdw4u
s7nTaljsSbnMbwUjEQM235GnUqv1GhWCktVf8cHXzwsPfDHhQ3uRU20OUFm6A1rR1g+4boaFggbL
7/R8rJMqJLMb/GW9tTvvJTBzu4I6DLuqBs1GFLIr9WlBZyRvcuvpCcewrBnoAKfixDScznzkb6R1
eV4JdwgA0pxXSGipBWU17fci68ITXmonSB1jVbRfvPLJ4V9Kj/CdKTMiFI4+08ZxlD5b/NqGHcu0
hc6Atqk8ZuPK5v3zg0Kdce6kHVm5onwWXlHnUhijcfAwti3leGqFMGuOWrVCa+F0yTh7eA0QxNyB
OuC4imL+zaJSHgf/s3v/kNug9QRKyhv79/J6E30Ma2MZph93mKn1DjQR9KYAxSTHwWwNNcM8GgLP
MNhVFORyG26Xur9vbr/una6CcidWj/MLcQajapGMPBCc3d9CZbcvDtzWFAVH+QHeIDLmnEaTaZoC
jKEuaAJROwZRg5U68qToIvJac0RO0peyV1jTTcoLdN3bUlv0lZM/O4ypmBn4DkyWdI12AkjRmeYH
gOaxtXgi7Mzy4BSjgD1rtGDkMXnneK9M6ov40lJcf9E8x8zKguWgJGvqs7jVXLBlJN/ZQ6LoWtbD
T6VCXC3t3pC20yN3SV403fwIXwl8aA+W9VIO/ql652PiVVaX6zfNteTzzUBhUHXYTst3BfX1JGKd
dFOr/VVlECfo04r+RAX5HwT97X4UcW2NRgLiPPyBsc4XfAaB+3xbXY5FB7SYr7/m64gHmmK+7ab1
/xIBYfirNWaWczhRCahBlJzjrYEiZkLwtLIoKhCjRW3KZgnfh1fYild29GQp8QaZkyC9vmbcZ+LO
YrL6XSGG2ppw2wxhe2YRvkXCk3EdO+uZn+JgWoHtCxLAIwwqfOleeQ0seMb5lXZCn312u+TjT0bY
7W9tMzt7wkZokdfKDR5h2mASLXYO+c+tlQrVWsWVU4UTpsTJbapHKM+8LH8g2agNn+fWIHND6TpD
uimsUA/XV9fz3ZV+4RnxIBCMv5pcX9jjWnh++ujtzoJAsV14wyfqTiAg/URU1WPf1GaXSziss1yi
4CQE6TLDNwR/2fnLuUJUmC8L93WveMtAZKaB0xxEcxHHWaJj7juJpm7ajMl3uGzHQywgE+Eko6Km
+CzrJ7fpU+RJQRUIQsU4FUpngOBZ1gsKstUYSoU5cACo2iTc/zdR2q1ONwW4PzwaeStJfHWvnIDI
ldq3tfeLkvxwewDqZn8cvujUPZ9o03JraPz7ZFQuf/oRGpXEF5G/VTqvtLXRfrOrMitQNx22PMsV
wIMakQ7AGnN/rSLbr7kC6/h7EAc5LDt2HUdDh8JhYs6VRdyD6u/+8bTR7SOcvnvGJfM6UbVzX2Qm
mvs14x+WWCF66T7Xa/c939oYc6SFn3YEK82DrYraVBEngaxLMvfphQVnAZTZFL5U40nA3Z61ue2h
rjKJ22eCeugkjNh49F8UiQjcVpr7cE+YFliyh5b1gjhQvr7FjHo/QBLmrRL/bjp3t37ObXwWO9Ep
EIq5hSCs0wjniXAU3QO9P1DUXKLpQcwBYz8K67o3E4GL4mw9GrdPxS86+LIjx9urNqb+v6nz12MN
RMDeexE+c/1zP5klpI7Hv1hEIVXBkaqibB+xdEp44PKqzWGmnC93jscc9SyW7BY+cqlxVtzSzSb3
7rDIwxaCg8NC1l8Hhp9g/Ush3ol3EPzePVT/YineNMrykhQlJkEnS8foLmckYS4+byn5lgmQUA8t
NRt59y48XsE1Yu5lc/KGT/bVwiVfudKPSvI7XLiICmRy1wNKrgIx2/zrHZTVFl9VWt/JiE3ZYPh6
NyiOntlNB20sFkvyKJCxC3kybb1tBoGoNSD61fNf46rUiNRMvYAIXiCcgeoxZJAxULKtd320py+J
0HvG3omIplryVrm3zDGoNViaK6dWTN+IFIYp6AZXfYwin46dqCXPsS07d11Eh8udVqXG56D9gvTI
3w01RjxOEDZOTomKRaQyY8pQ3Q+ChTbjCcN0MpJO0dx5/JTYgoJ2jC7RlAWHh3+KLIbKYh+T3Fu+
8HJzoo3fXMxlNTiGMK2andSWEsHYwyHWRkcNTD0IBzkheVs5EDmDrr7u2x9fwlOIPXAwo+rqZlRb
fOsxyqUgqEuntsyVkl0xGJ964TyCBfDfXb6bez2zpvdH0FJaVBR6Xo5mn0Gl7w/2yE1L9Z3M0Tko
G+xwqU+Pjvtey3TrlZJY4sjW0XxRIf+IUKetTUASnn+eK9qUBjFg8TkiV2Yyyd9xC+OO14KrLWo9
iX4juDPtzhE5xqpLt3rt86tPLNRp1UTUgYoc7hHSqfGuw+OS3d3E8zDDGpBAAfku2rv9zuFcRYAt
9vGwyT0CBDOaKizF2xszrr+9NDDTaAbacr+AHyD2bY6BKqh/ck2mxrGRApN3y/IPLTUw46VeLMNU
jkYMao7hKiUT9es36+wGKFQpEJco8NQL9t3a4Io62co85Q3SvP/Ge2hWHyRvpSn9CrHtmxP4SJGG
VQVZo6SoYhL5yIMEcd61x3UJWQowNz+PSy7b0mo2U3IUnm9/OimMf3XAZ2lV0cNVOyqSB9kcZezC
4dmkEFyKLf6Tlfqgrtwf83CrpdDFccz0sbfA1wOToERCy+WMdTZCLaUlvahWE56/wOMEtPq8MHn2
t6ZRXRDclpBbnBlaE05beiEc8N4O/ca4vp8MMCpRXcVrcuLOgVk57l2HFqobSHKezOSU60CTCc82
naRNf9iMZtVrWr+nx6s1C0VobM+QGxc6OBDh1MePPP6xFDZZbu620ZoZ0vndE2iAmJLgtaQ45Ma9
aZywokgEIdtYrU6tQDjMVOrFppeWLqnWvLeGWvqnYVuLZx9xBZc4X5bIwCtz7avahDaMq4K2BvDI
EUaw5/kgC07FBRg5sByJUWQSPu2JVbr2Bkv5ysHho+HikHxE0HYBPJPMKx8AXtKjka0vriKkVCjE
EeiQ+xE4S2phjLbLDowXrlGuKeIN4KkXFWefJrUqfso3eIKAttfP3Dv+n8yPU4oow3R5kKPtmjQX
LMd4WtfZ9XkPLPqQgg2mA2hV7l/old7lG6oyo6VlD2JOXq80amQEd/eSFiyuaDg/x0SoQH4C/EdO
WkKm6SLU1ac2wohukmGwNKTU+6NJhTCzEEpyjr9ZC/ZBuF9kEM5N5cZINLx/hZCBlKyiB2vbvSyN
bDUpTUViZlcUGqVkQByyUsLNHsoAi7ef+Jc3j+qWH/YL9kaMTvb+rRxQ8wzy9EX0tC3E3tFMnKUB
vkPnyreHuMwZR3NSw6T0jawdK0DXpTLXruhhDfMWg4+LHxa88xFenX0UzRKrm9t26JsMFKBFiXJS
PK0XZjD4u/7WfbJwPGMgVfTED1jP9RyjVx1jiwfTiXA0Uj1o8tngA+AJKJz91CF5qMaOsj5S990a
bypWUS5rCUTA1p7AE1qzFihnU/2qymLufJhaZ7rpEB+J0DmuXYjV8X2X1rUPsJoQW7L1QL06tdvk
Gg+PmPsfCQZQjbRisrTZyFvAAP2axnDqgHgXLQFVJT4TRUqK4kPRMYYAEEv1z5PLB6XFvtlejwDF
8+CP1GBJr+YVrPMfjC5WNdat+uZBGw5xLBo+QzGVpd3VSzEDMKxa5m7EtFcUbzd0sPPrj+LFRTTw
/rtIRvhOFIp9XWucEUxDmmRTmjpQmO9lZhwxk7q+9z6ZtcVoeFwzfDG7Wjn9e7KSfyIwQpvSrhDn
PlnnF/96l4paf7Wtl14Ets1r3/JzPs1K4pFnUVCMyAFFtNo8XywPVa2r5x0fWeNM/qHuCsJBW+c6
KHhqqPyuBHxF4xFLtWsJUnCYuz+Z1wda0Gll0lI3dbM9tlUcSs2vkVCny2ZZ5uC9Huq3bXU0XqVK
2NlKR2e2Ciyapi4YAY3RrjyAyisT0TfLQ1IOL7MJsOVY8JkQ+BTUofK5npuWWBoN8hA46U2rYrC5
aPso+QWnT8LT+ERy7FqzZasNM0Pa/2LwemefBQXI6qWXhAnoEXiXgJvoC8SEIFMbb/LItG7Qq0En
go9S0rBCMMaRWbcsUyzgwDC62qSchMMwt+e9opygoi6MOWzc7YTU/VEtAU4WFCaoFhdGro1zmvQ/
iGlWgaP3kbpT693D8vRBh0yWDhXwRWkYALSmmHJlpdk4ymMcBgJZaj/i7Eo5BynoWQZtCv4aUUXB
81MOnKVTSRC8rkT/QjKOg9hUCyYfbMNqxhVEsfUm4KT4GURKK+P5wu37TRH3HsVG3P6kM8TH3S4g
uLGBHiSHaYZDcSGBD4M/p1Rn11DBoAmWUZWs/TJ5byNFOQ1Wt3aL+XR+v4iFVhvE+9Jw6ftkLQT9
g+YAdmasGtfhwPj9PZiM4tFaqOGOS3OoIOihhxTOkEzIJLSISog2Tc5cLkiqpfxKxBXTW6qWz3lo
YB1EGUiKgEJ3sK4wABopthEBCouCOGHV6IlD63c3VXRyV/5OGLfL2KlBo+BQawbn0a9FlEjKDix6
FdBcP4UffMu2/htAc4RhJXYDl7NaH/0rfwMHU5g82+DW3CyaQYxYiPb6SI61lbu0tBiugcmRqUdi
mebjHZYfd+WWBQQH8TKXPkKZvKoyIPXyTuzt0IzOcyAXsQKk2xQQeoIw8fqSHjb1pFjs6PkZOV0J
9G4w2oNncB0TxrCkmoGuWWrOFqomVjqcGRq1g9wqGP/VyX7ggSSqmrZKO81vp6AJ4ch5PAgFeAV/
W9qiyju6ps4R0lvNCAdtc56CTZlqzKg1sGNyf5US+y0TRxCuWGBlzXZ9r6nWfu3ULdlTxpvO78m7
wzTvWKp7ZU77ZN47q6kiUSz/oNKpDozSdiM5tZXWwFl1iooPzUO3JvaGf+vlxwPr70/tvxagX7Pe
ZN7EW2dkt0SyXH+eghG+kb3aeLTqn3abch2wmtYtM8SCHwTcBXAQMUby5GUNADRGpsqdmAvxWLjT
u4Jgdw1TaPIEpyMU6OkIis46b6iElLhHWHS/fRI7bShCSeODMLa7VobGTjsZGjkTwFRfVmgeq3kH
iyBud75AIY0g743epgA/c/57o0V1nXCTY+Ouie9jxyzGxo7vnXzvmXats6WBkO8234y+IsuemwSg
sjiP40MaH6emGGIRkSd6d1QXMZAoVUeSW/e7oSQDEAhreBzBd35/QBlhA0sE7unQ19ltJZzy6jdz
anfHX64d9+L00m8PbYS5YM0BJaqGIbljTOT7Gl37XOA78gtpVYbezFRY4CpmzhYjNNVXVVbJPeki
oLDGQD8Rm2oL8eCcDMtTcGwoBUS64Pdo9fDMTZKYzsTMUBUu+2avLYX+ApDjqHLxOyheKgmkuFqx
TjGxFn9Uif1ufhyOsOjyLT2rKYusJI4ahWUE0sewWRgFYAeCLcmHAlW89dK2K3BqeZ+/ljf5ENHf
rOs/EP/PvY5Nd4IeHnUotRn3J8pGGw6JOoXhaQEgwhRgodWa2sD1HPE+7VSLNnsptyHoorx9NVUf
QP0hsqyqoNSNKuvctiUJ4kU1TA5Z76DKKr48ztbvHz10l58CtaJLybfqn/GAlbOKOxhPR664mfxp
YnGwS1yIc41PPA4LT0ivhrNSpZLqc3dF/n+pUzJcjh/HIX0F8Wz00p6rb1z+GlHPtK42x3OYZ2jo
v1avWHPv0ChdreBdfxAbxPj6zzxXr6iQTKERVtEo5ys3UirQdfsfWGlf5PtFBg+LRy2g6XT86oQO
87FnTqd9dC4l6QnNQY/7NaH6uMeNuSKRGk7CjJedVGNaZSs8y1nCWxU5OTizsRRH5RZxYgKV2F8t
EUhkIX29H61AFPR9bMPTbulzx+30qc3WMR1B8KtUM2DUwwbT1bkTvcnL2kCX/grnkalsCwx34DHe
/pb9R1/WnJsnNyr6Jl0/ltmBnyrQXALYn3KrqLkLeDBhrqAZsIjWdltMW0Qlz2Y7+cL6HCND/jxw
Opw/Df20K2kDeUdj8ATEN7Ho7qTt4dYh3B1RoVzKBPiAACHs39YKLivDTqtR3pTNzyuAfa7gCYV6
zEatqDpzJx53XPpxnNabpGDWTtMgt/1z0CPB97sTEgVIzeJZU+LTN4j5gM7yVr/ICFjXGyLJ7L0q
WzgB+0eTevf19qWI3LxkybnIWDKFnUON2kLGDJvlV2PDLvl4uNWmzyS4Nf6Ck8nnhf4eqkPmbVbZ
qw6pxTv3oXEJ+uoW9nKh0u6a2fDI/MuX3tR2AgEaj5O4NVGGFXRMe1zNdkFQ0T0G6mpJNOKIleG9
6Zwz07IrojBnmN8QRo1joCqqyhF1cbHCQiGcvlv0tSrKV33ND4viBQJSUuoaEy01kXeOz2FldETe
xQXqidkiAkyZzhpo2xEuVA5j4iL9PY65zZdgavToyaW8VQ95XZBAqbFr2OujJ6aJpmyBtaEQ7nUK
p4fABVXDohAGiVW92qD2ejfuzHTGpPlbomIuCcK3AavKNIbS8mik7QNwCozZXLRoiW1xU+JKQK41
Im7CSFA34WNoUlVAI34AB028l41wXB7J/dxm+LaPENsnLAGhynIFeWqkxapNGR4kmsz8jaIdXzQV
rdW2MHeZBTLJMr2q5p0TRlotgfv50O7NhMzAOwAHzQMjDc/haGWfJ+yYaNAhw0oJAlbS1ny60R6h
HD6dGStlXxBzDHbRNkIdxfqDSXu5UTaXB7OZrTVRGX8/yyACWyMJpLnIcDIRRue8CTybxeBzYQm3
6rqMIit9MX0OOEZpUacPLG/YgueT2ZLEotSl2nALJ2W+hqDw+SRc6/uClfb2NN6X0hsQJxZX8dVC
yR8UgAyVxcNd2T3/GUlwQd4T1LGJ/itrZ+b1ZbyPLK90nQ0IIf8YxgeEVH5zHt+DTothtVpOIlXd
2lrP4PPYHQQImWtTFl89Htbcx45F37OyVUGCksQ/KlT621rF8WO4nwbSKz+chCv6yo6WtwvRuicl
zOnl2nCLRl0C7HSswQNU4D/YZ1B+COiB+o555x/cCSXxHrgq0jeeXyXu6T76naUSq/zTQ0A4+x7K
wv0GfC5B4GlS+nz1A1+LAMHyn6VXHNrLTeiCGxUtXHlpEBHkd3BhhAMejuPhmPDOaL/FYjolkJI/
UgRUsQuXG7ZffU0w+/ZOMvxPXeIDs/F+8TUjQjbOsp5HdrpcS1UitH+ZmrtyWEDqXMtit7/wnaKO
MTIL9p/ldoPoq5s1S0DiF1trvgqgxf6Y5Wz+SNPA7Hd6qjDc9G6SwXwGueEGwShjX2ysPJq3obJf
ozDoJY3I0N0po0Z4hNbrID8lAOBNLswAmx+6Ba0DDBQXfS2KLmKdB/E3pncdQS42dlUPu7GXh0in
7uFsDosApNjNks56t82/pxlLrgQNTjxQV+d6YnsZhTcqkGR2VhEO/4v7axUtBpm2gpHYVD77EZMv
XVSra2XRuPlc+w5bl2WpDC/FfPChHBd3aCgzUvYBS4AWTE7rXXs1T88dt2GUg25XkneKIOs0xXus
EX3RUeu7Q5s8IGSC373LgI3Dwuwb4UlrHuX9jjvsXmnF5syt54mV3jctzMa+pln/uvXOIWnYFGL0
SN5tZrX8SQlbkBjDIHQIeJCJ2GCPafgikZhtobuSiqZDiJ0xQJ08FjZQ/mADWgRVvZap78uHMp1w
UKyyMZn6X+PDhzVYU6IhOCbgqZ8/GyJ4MGgL+xcR8QxIHPzznRslnpMEJWeiOIT3/Odw5N+LUmKq
4JRXII9CnHjiNbi7We0QtrZxeKWu7G7xb+XLdZCX+TcoGqwMlJ6UEYqt553ecwVk5omw9rUmQKwB
9r3zEDephAgsx3gxlQ4Sn4VvsCGlkYrifO9e+iZMGBuu/0j5vzWJLSMnQ7RuaIyx88g0aQeMiTgL
BysgFdyhF4AsmTn2Jnh8+Oh87bdMAC/2AgzevhC1xc0ZDudHgGstcwEWsLJmA7v7di3TClkD2juj
B88l/5ZntZ/DZNMLeiRGvxWj/AHb4aaGSKl/bwDVFCbJwHVZ2VjmXW4BDJa+CG0a8qnEajleygCe
cUdhcBMfhD1mFVQPIFSf2K+gow55fLXyg/RxbZ0EEzVjXzJAUSIP4ic3/qz/P5/CY7H4jR/2sbkf
BoBy4fcTTNojtNurwcmX091xzPBAM5VjxS3eKO8qpbpZU8QwL+RaAkhTlIihjYUyCuyF5TYenYB7
HMOUNoXZ3tW4NbvnvU4XPHWSCTMmaRhUwPnxWVv+xCgjD5HNUaKXYb1NZjlKQOoNLOUz+TDOPkDV
L6Guw7mOKDTh0KRCBDr6DOwqbiHX9CDbvR+E6+ZImmBdE31c5c1gQbNzApaTo0J5PurwqYXSkZyi
L+mKzx9zZflofkhB2tVmukCe/4KsDMWMrgRZ0DUJADOt6lfkMlqAAPBRol2Or5IDl2PuDHd2wegH
hbyl0nDxZ4UpXiA0wWV+lZ+R8VmTgTE2modbqBZrzoC5hI213cBQ4nIL6VkPzo4cqzhpyXuIPmAW
w4FTKX8eLqHcUzTvmaCVkjvuihxj2nfCtXvwJmOaGjgKJaKcT7XlTDAGzS1deNAT7+K18SzjKrDr
Khze/lvZxvCpYbhXhiRL45TXSduT3F0GK7UApFXVjGgIuIdu85VC2W095zbJfmwnNNzi8m84tUty
/7/E7kpLiAtJa/9hVwR0HbEPK/GtrtA5a5j2cVgUPRLf00Yti2G7c3W+6yG3ZESBfi8zHn7ZSR0N
TIeCu6yNNNgfNxChehkt1Nyd7KPW3SWpyLM+Ry5+mDtxiEhZiXXFqDz2eAuOSWsZ3u5As7wkHHHd
KHCANUkZbBRQd/1W3TxfKNoJVHJXEXJ9HTR0C0H5Ffnj+wqwhPT/YLNy5m1xjpk/rZFRI5BiojHL
+X2Qm0gl+/oHXNZfZKa+AeGQ6EMzYD8bc2W/hRmEZnJ+V+5yfe7N14allYqkC7ux0UbO5MNtSyf1
mEIt39zcdK4wwQra0JzoPdYCj++Rfxl8jehUmvLnsUVRim4YnwUxey/jGoySvCLIfsV1nCMwBweM
VTpgOP+EOixpF2ARl8gzVPrHONvRBYws5q8EZu5GObauElgwRzaQ7PKlh46IdNit2lalyAQ1fW8p
IlW7KgkpNSkaNQpYvjTr6flWEtdkRwf2QiJdq04uyatkVH52KQEpST0LabidAzU6wkQ/F770oJNG
JdmUlfEa4UVXt3mrhWKMC8yvVz2roP4Kz9Qguq7VgX+ZAR0rRy2OV7IVic4Ni43OAvr3+3bdgvnX
wsr73N0b9GLdIdkEm/OtufFoM7YijxtowzY/50xeULjQTd5EgJv9pfVQoKwgs0QO18z/i/SKZzzg
3oefGaMk4ytwArAHWQErpwNGqeIr0hIZ0EzTMRPYE6L3JFwyOLyYfMSBZWNKch//DmSSEY9zbyeg
+scnzVqn8SXw3aSyagbWGYsTlUMUq/Z1SjKBtXoPwii+2zUPPCNJyMW8A7YA4y9wQLyAlD7Gijzh
cEUyUS0vcHqpILFS/jfYsKJO6Nlrg2AvMh/86i93zUcLddB/Pu6DKMmrfJRo0jKoz7pil8bRwZ9K
bXDQd5regdPIaPfg1d7x8jSjofWyeA5ULp/0d8kUK0V2xTzd9dL+GaOnTo49zZP+TdF9ipc1HQGf
8goOvA3S4N9Ct2HWO/VTm9nEdZmmVtcz26idUBKFhahPQwuAQ31ug+oDH8JI6k5M4Ct3pQ4d31cm
3i63P0497eC1mKNB3FhcboOt9PAHgrcF1/LCQz6PJfF2OTTEXhSNZcyYcWKdU5Gf11Rvb4BUt2De
WTHrtQNnMyxSaiDs6I9MfNEAcEi4AblVPsg/XT/0ZuqM/5Njx2x9HCLk4wBdenZySJ6ZYAEJOexZ
xAtlnw7oT3mdI+MB19HkH4pW0oXlIC2oo1I6zGZ1lAvt1AWaBIet6qGMobPpNQrGd9UoqbW93iAF
r68z3D13s66LglkChTsKL6XIqP3fJDXyhYcqireZlkGbV5n/fwJTk43p3kem5gVb37MJb9AhCqy0
Pz0dl6OmPl71uoW/otDFngpBO5dQhTtFVRhEtquVM41bIRYyUqafRoQ+7iN1D8Yl7X10r2TI9qZt
ea7VDqvep5WWJI686NdwXcOgn2UMF/QNP6bRv52hP4eecqImZqyVJyVFNNG4/rBzf1bj1ClwFz4P
vM76mqAUMjKnAA6RHF/CmpJm+jAsxy9VcoVp/RPvEl55YyP/wiOWarrL24D+VZc3IicD6A9aNAss
jvDS4g8A/UkQgjtDaEPEJL+OtHXVzE5bs/34ERy5kL0ARnwY8ZjhzO2EaE+Ggg0AaOwO1Hx4CNmb
O6bM6albkNPQ5Sh9zz45DDVVNd3On/nSWAnj+9F290rYKbgi5986whEVEUVTjqZt3bkAf3MgR2i5
SGlrj3t8Ys5eRuwnf9UAljLVC1y/2rjeuyQ4fZiBtzNOp/V84VF0uuCL+mlmIxz/ysH46sPMp2gs
V3rTRZqBDcomX3nl3L+0Cxn8MA5QXPhIuA9ZiVubl0OYE9pBGHkiSVoAbWkmeQEiVAsdfhtN2vUU
SXOGA1OyoUNmxoQhyzzORYWWcAYNaNGWc23AJu4j7R3BmgfGhYK5BwOoMGfXLWjKpu1Xe5dlOFGU
03cY7p4t2VkR6uOgn66el8z/4pUUYkAeasUOYvRq92kS29alPCP5kcR9pM98IUESFcbDWSZHovYA
kY9DUSMPqYi3/ltJ39x/nY8o5MrITZFMyFtiPqYPSZQGTFObzje1z1oJ3uiBcYzL6cklyF4yatb3
rbgD+3eVXGwvOZmTPGNLBjo/tueDbpFDXDsuJ+s42qQ+QnqNmi5VzhiBJxpDiypRByzwxEV6ULfo
DC8g8hWPfJUjn6P2IBCPMv3zsNZNVn5kLVoprnP+1toe7rnwciGNCs2AXGsM2Dz9+eOzXrEfm6d1
0P4ZL/rymS9++pcv2D88+EbUxrctACoiJl/VPfEtlI26qr6RExB3hU8QpyNg4ZN25sXQeV8IDx0n
w+A73FVG5GcdUbXyBNdZoG214ddBFClR1vNZZrZmJJQvRbJxBrhltw3LQDziVtggMgTbDB/K97iM
48CygOlDzdlVPGeZi4f1BuHReJ6X7gup7f74dfTrS4NCbErgXKgZakQPBR0O3XjpJG9Mge43Dw2e
yGuhMlEJ6tFP2DIlSQ033U0O4DDwV4rqy6VCEl2JKzjsxxc8PPJaK0iBvez+QAXX64xB7bJlyujH
6hXwA21fy256uT6ALzeodT55owSD6TR75IwwW9/MJTnYjHsjPJ+ouldxDQio8H8zxxP3qrJIId0l
WClSnI3AnBm/YjT8172gUxZhZj0TLV8sreTPWgBjULuZDA7dAb/fDaIr0DohFCjK+JWYX5FVyUA3
1uZy/JTwNhgJgeKcvdbF9RSX4hFHd6yt+gVGSy9+ItiHW/BvxEAcPviP9z0wGDaedKbv7r85VNmS
PSEnOf28XyEQ/izoxtMEOyZ9xCXzSbekF9myo1MuiuTE52IfrDdm4PPMQUjr6YGmAI5DAQu8W2z3
dExidvrSufcYA7F2MQneOA36I/EcxlZ87U2P4NMSSkNyaNzg3UsJGjsy+BZhUGHCOdLr/8B9Zr0/
KB01H1dNt0McI8Bk2QwISjXYphnqkVxkn77zqo2ojIE3UrPOfLqrTjp1bWaZNvfeVGsfTGqJcvaP
nNHFFuk88bBvhd6WzNs6zVvveYwtSNo71TSKQdEDEHKS3gArtRWn9zXqBTV0t8E6NP7qOjqbS7N8
FUMABInL19kGQFMRXDFd8hd3qQkrNmoeaKbLfqt3qNxLuumUbI/psGe5qyOCL0K/oeFwOqLpV83L
U4NBkKHmvEpoG2U7sJ0yiy+r+fTWzYouWQ8zEqoOd7q8zjIKpemB2TW0UseQ+vY63931hy2NhBrZ
vxOPCAdsF+bVVAYko5rPsnOqzCqAQl+8U9cncUgTNerJsk1UcBUu9WYqr2PWeBB+gcRT5tOalPw2
V1SumAwJJ4kB4OjucewefHYXCtSEGSEuM1fqzYqxm4uAkXWVXqUS036s9i4nYSsK8BNgawuM8r6n
biFrJSEiS3mzpdhwAkg+5A136TT4miVI6ZaqtoDmFprB5a27Dn+DvDcNSWgBu/oYE4oJpalGPQUl
LFrSh2zL0K83FW3uCo+eurB9TUk6D9Gjbj1SL+XI9+rJSsY4Qf73VsybOCMFPz4g3HUDiawgEjwe
MBIE1jfKILSfIMcx3YOvc3u0iy4ccVpLI47W37UF2nB5Lyky0UR0t3LRyaBrxUsQuWnKBhXkdN93
CryJpoiQdMwmGrxVQUkZaH0RY9GpgFN2EAEn3MTllGyvGDxu/Zk5G3vuXkEImIFuWItj5aDHZM5f
ADssBp+xdM8Ua0bazb6YoUZVbCDganySPVDVc3S+56phbDX+NWx936sMOzjGlD7RkvbU7sj4Irpn
4Irrs0WqVwOeMC1a01FxFNQFJr1qJX0Fgr0AgnN4RqpUikdwMf3VgdtOXGV2Kv7m52GJXFZLYWfB
EKQuG0WaW1FSa7pboUfxsOIXGwoQ6ol/QKNMzfbPtDDNlPm2LcrqI8Rd5uMPJhoYX89tyjrQ6OZo
21qKdVQMjGvGZFPnAwz2PkKPe5/YFdXhy++Dj+AvaoqODHtdZtcZZEG0BDe0owKa2wvFEoSoytLp
ZUlp+FolIiWCGj8H7BJ+vrtHQSsSpBd4cAg8cYiPnkd+0eFZdYnIY3rv4eGsx1d0+qbpsHtAasS6
ynj4Ke0rcMBIvpPaIUrUAMTtWvBBmMShJkP0nhJkpwl5tWyDgrVbKPa9eafsF0Nss4sA++l//Kx3
cHDXG+vXvgWLC11BjMEsO2sqNzG3a8AadUnUdpLFOLDsyxhD7dwDHwr3ykRT9Rs+S51HC7gAsWsQ
pa06K37U60CD9umlrKuhJWSJk1tof2b9Gu1PVcxIYuwuVKQNVFjfwF3ZSNUm3/raJxTZmrm56DRQ
tbQpllCrX3UCgZDHKPmZdGr4lRGt5KmtGkll6Yzz9MoQuSkpTA/82FRGWRG5P7lNFsIDSR5wea1k
iTmPBqnm8GC/J52+4wQM4kFv3zCssde54WPDR9exPt/f5QuVruI544nZIuuQG2DeCWrOZCaweHeG
Prwq5hKbvCOmQ+mi6C5FfO9dea9kenXwGQsWAu+mNMnWYxmIpatmAZ4X1QSvKFODNZDNPUhtwuJL
vx46IHhZogkpU5SgNwjoWXrYVZDLdk7o8ul6Nr7Qe+QyJhobTso5mA0HRdk8stXZCaAJLp0Bu7+v
PelMcvhJFA9b4fummGDIlOTqSu6uDzJAp7+oxUhogtkxp87Lv2i/TTDI5xWNtC3fnbt0cSLW0YuL
biHdoEsnCqjI5AGAN6as7+z8IOwT6/VJMSEWq04NqEGSZY76bCHQjlLcIdnVLtHMKuuy55CB0bk6
4aFdQvJvDCyc0bvRwcdm7OHjcxNDQeq+M4mtQABNlNmHiKS/zN6yQDWv1BorvnPsgVZUtBd+dzW+
MutNUV75o+ZzCAZB16atcIVpHl9jc4HYnU1rRlJ0dZ8YNB8kKwqSCF0AWbSHOLrcs6tFOqQcjWhq
08SSIpT3nLqz1UPog+ld7lIYVQBwYaXmIQBDiRgHU8ogQ7QUE2KR0Vwq3FRq+oY3zgb6MWtvmnWQ
ui96jnvs5oz9E+txVD6f2Ascb7hFfnQfCOwCF6uDyWxju6HBzl5+b5G+6s4J51ycmn1CySTgiKxX
Wwzuut1YZUWnP+RUlNq9etIMNSFf11R7fh9iTFgKuzASdH34yWqgzFKAeyzruOtnfRU5Ue8Q6ckX
ClfT86Hm1JTL8eJkdLaYBh1uvnVOZC1IGiQu03nZ7ycONecmaM3NEnttD3m04jaIvUi//vrry0yq
Os+wmmEtrlsXj+90OohPBKFT1XlSiQRjy1dAof2hwICOAX+sIJ8RS33SVSPpPipINw9Sjulqmtkb
oNNSKOt3i5QrJB7SfWzW7AN4O6QZHHgplatqb+atRBFGs8SOJHiWN8Osl9Kh/LRZIzu7W2vYXIIr
M8KtJlN+CmWYWuyrJDGA01UsNWPw4f8uidrQjpYoq3Wa/7KDb96oxcKuIQnn77ZG+CL7SMx6PHNL
7GWV140wB/HfsHCjqqB0s4H4tSQ+6Fb0lMuP6nSlUFqYEa8cQLmbEplIf4exbaKji3KpEYnRG1Nf
8QmYEjZhAf7v1DeRT7hQ/ulSh+DucSM0zishQhp5S8V5IyY6+9bbVbaHWQgh/o8Z5fnmAdH+t0+C
V/J2wMPp/SSe6SBzkUGlPzQ8H8hx5OMjUi59dvcDj0gG37/k54D1Z623lDEFpulvuyMSkzOuNrFX
Xd/aVPlPgROmTtnEf/ohuClwrgmhRlXH3GFxNsyLAZ6hzR4qYvRHtQjPrpzAeZfZdKRR/pDo2kMX
2YVw8rf1LU92Sjp1eKI9zvPOOeXc4eyDlekiCgE3K+NtvhalkwsTdrt7edvtvShmF0sf8ZivWTgp
MjUd3Nuw44hXmkX9Ej7gAWS2nrLcsyiiUXJ3HR5kHpeqj76DHQ2daFWd5yicR/1ciaf+hNNVWBMq
HO2zu1XLMxf3Mszkzf5LrzDg+p5nbqXZubfe9DxSDCTXkyTerrxbsQz8upVF7BJfcObWJ+kJkbj9
a4VE5S4hm85K4Bf9zxuD6uaPzjnazKMTL1fkzjc4hxkQwwMLA/mEaI9DWdsBGTH4XwegsNktm9Yd
oQSYrYqzF6IYwpxrLzPy7tpXRnqMrkzAdp/K3QHYZEBbbJ0cfx0V4EE2PlcYxygQeEwnWsIUo9CE
73FFrEw8yEjynmJbbwEexk2tmzqjP19dabttM9t+O07CylDBnCkgmiaB5Ax+mzRNsS722QS8APfD
jWOnU1NfC/6Qs1KsWRPScXGi+cQBU4PoWlUOpOQfn8pSVB2o/kX1Y7onq8JiaqvRHmoLWv1Cu0pY
laG8Ezecn8UAhjyevInb8EyoUjmKgcNtJByO0DT7snnqkLt2NaihvtUYCf28nT8VZU0EHfifgR3A
U2jm60k97ZawJ9el6y8vluvljG6oI+QUXGl8uiojOb7OGCI0nTxy37r4CNsTEgTyWoGLtSGMfmst
DWwGTzTZuVgvg+m3S/kg0aCRKepv0UCCUoCQ6mhcGuUUa2U+TR8GEoUlaqvug0yK+85agRzGOdwI
9JvhgK/Qt4mnB/Ckf+ET9h3tv39xCww21c/Yt//3wcRd47jr5QrSxgAZ97YgU+salI7HGGGUC8ff
wehVEZUBRLnVV56cV5JrskAA8pWjVC4A788UZMC76LbQ4cqZV/k4r+0Op8tLKYtuW6ZgZrwlcBT2
wVk6uVDlrFiuHlQtvIcowwh+KSkcJ+XVIu4yu0yfKQV6bwR3kdv7J1/Fm9yjVOlrdLwayhEjQ6Rt
4hR2OkydXuZX22/QRC0/TEzX9RG6T6scv4eSkVbdymXqDl+W1hc2VlBYigdYaHJg6QdWAufPnjRr
mjcNe1t2GRWVkfKlbIXdw48yNdnABGdA26LpQAjHFPLm2rttP5NdusnXGJlcR4tqb9pxGB/klQwW
THfrL0e+H8f4rtvGL70Jsb39hjXWfZiIMTN1O5Lv2FGc+cZJBWLe6soaPxHv8qhy2pikQYWkV8kZ
L1vFxhMCGOrdv4oomG+lDRHLo4q2ozUUdaCDPq2WpeOTy43ZtDSRXWI+et0lRwdrX8mh913LWo3D
9nsFp2VCPwjzFkeISpP7y4ItbKTpcEKa83zsaaZeI0Kilbb8xUKWp+Eg5kFYdJohUTuQhJfw4/UL
zH+dpIPzE/mqS7EevljuLC0OFybaoqQui1C1S8yDR11yCl8SMdoKfNpgJh54AQvOspIwCDSsaXL7
it6lwR7SVf1xas/CQ8+orHWZZpIRfuokYA5Bd+yY2aMgxbfvZXDoERNesmFBTPhYRcZlw15W4CDC
FmlFqPBQ1A221Aw8AiEDk7ceJD9DNxpTZHTeMprYEpt3A98d30g2yuSLQxmug+O8hWsETc07qhuo
qs4tsdIZzC1GfuHKqHCg2SaZsIvF2han5Cb/EWAiMdhp+/dUUuVOxRhzWLlPnOH2V0Nd3aBMzZF4
cFd6lNrkgXhStI1kjukzsWrFHkSWYaJNvTaBlPkMi6XK34VI5NRaJClmnCp/zXFIc9pIBbJ1aiKf
Vq773bOmnDlpsKaH62R9Ru24aqso2lSNd9nxoePTcWMbnv5V8ON607eftElYJbvaP0weLxhTf5eF
MPniia0g/PPoftS4kQAzGvGnnv9vbr7RjzzQ+H2FOgi6yqBLT8Noabsv4ivIcEiAfSjBamO0rbqj
ZboRZ7A9f9Lgr9/mTjCRg6DvS4hBnVOluavDexTPhq8wnOykUfXYR8Q2tGMV7QRnVk8zAI/yKWbq
u80MqlCcxdkGlNM/KunGcfkQMPp+IRLrJbJ8/J74/I9nZp/vpcRLPMRH7oqVRRv054QKYQGqKiT3
uy0b4bMUiyWEbv1uDTpvQ0nW0u1k7WH8zW7CWsZJF+t92aQNjTXbuF8I8hbcOnYPj3oRFrrF6Dav
Ks5SeJdzzkyP1iUebKkMOKIQA2Wi9+bclbRfh8JTg2fkdR5cR5hZxx0QJPYuvrVxOFGc9ZXp0sVl
0wruiXQwmiEc3JoPsbb20SJgDGyEEtcpem4OzbgYsJxvOyyI7RTkP2tMoyn+mkUEFQGSVskb7Qwx
yRvB1C0+j6CW/j1k8fmwGkOiz79IL0EXtWY7LQXpAzpzWg2G86njUj6ncwuF/vGB05vgx2/iHhQU
JFM7PGQAR9G1QjRCTZ/adK6VO8j+zH0Q4MRFbPcW4wtxnDkYn3c0M2PCIyKeGc21FJ0XKzCBDe6A
J3gGYH4eZYAt4rw3C3wcClwe+0DMt5UvAjKX4jm7wYPLOgus2Tre+lRoa+iEZp7QxKQ/OmhMrA7V
c3TKHFSZJXdQEoQGGgLmTaxgwp4rNawHAJRr8mJlkJ1ufWvpAt1RzKV/y6Bg5MwNaVaSUASJs1bl
rcrEowCoCCToyqLG15qKQSe1YZ+7/Rwb9dRCs5dNr6vMlPTBXLX5XGCPJEKK6aB5jz6uEK0kTQQk
FaLzZqrfgQsR1PguYq8uXSBc6FGlbDpLyPuDxZ197bTRD452I1LRNGkGqg6MoYl24IWbWJVLSLz4
tEiaL5+zWWzEmNh+XlBCxtVILpxFCHRxk4CmiLl+z+iyKKVz3jqBDcGH4qn2mCsFGhzwooQ4zP9b
bLGH5uusu5t1T/wvK/1uRkAfv84C5k2FGlc0h3mf44o98rV1P077aC98GTP/QxjT3Rfd7RT5i0c9
ISzPNT07PH9RX21HZ6ZR1QiM7qjE3iFZdpHJi30nNy8XrkRFd0uflkRe+rVAzeYtV69PtfIEJjdm
4SuXxbcbNM1CwlMDlvN9hG4pJunLmAIhIp8+kSaFuILXIVTlMLDsbSGIqB+NEQ+RDca2JsVD2YoG
lnsx6KOOdyDOh2C42qMnARKsDv13Ta9ne6za6YzmJgQ97iUN0tJiC0m54aB3XpdiUPrhAVXFVVso
c4yOCG5cma9XdfV0lvtTzeAllVZIybRqspzUOcjC0gawNV2aJjHMZM1G0ushO9GgAkHd815nQVV2
bFRVia0QLGgMt/8bJqro9aSeZleo2eEaQTC/K80JXeXjy1qR2XC27irMW2Ki7FN64u9DsTf6y94e
SRZa5YerEKD3icskA1INf93Bv9ANsHbRRz8YrplGFX4sWMfUGQiNserxIlJYVGLaHuPPgo8sBSdH
C7UOuPnM/FCNr/nqU4lJGNpNtFUY3Rze8RfFljAnTrdfRv8NZxLyGuMEgJrfSbuxHjWcBFUxMn+G
RSEvQTijhXkgZLYSJmpGXRIlbcueEHinSROa6fNRA6vHfAYcSXgGkjSMMA1Y1Orr5sObIXDVgfC6
/AL0WLyY88rGGLZ3an+z0tKohrFCz4Nx45j/v0m/+MN5Mv4tUla0rXOVWCHA5hc7tDk0pVL9QJGi
QyBnTazSJYTvdLcDUVcsDvKVtt+Tx1tH0yrfiJU6JIs7+F9SIMyYtjTlmnc0l/11GTZB+q6aGQ2u
aEnjWB+AaMcXfuve3aduEKeqT7GqH3IftEPftmacSFsW0GpXLqKNJuk7DnzquJrMU8rXT43I8c3J
8QDDdxR7IxC0Fx+lZZ1/zAQBy0b5kKlKQ0OoIo1h3Rer6CcHQo3dOofQScLqvcO2feXWL0QddQju
cjtPluW0GI37KDFFmBP0htDNwLbhHRBUfverIh5vBJUXD/Z0OEI7R2gcJUQa7MBsL1UpAU3zOLZx
DVR9w6PyfL10pB981TJ6U9Vob8Z5oQElYMPCXzvzwCO/v6dzbe89SlcxqXUgFfc5JNnloAr+IRL3
T/sY/+QkwKxqbrrtcAX7ZGomAcBfaCSivAvlsBPZHLpfG3LYYhQk5yR3me44TzsKmtI4qgQsIpOf
cjtiXBcfi3xuqKpKnlchgHU7gCZIq5U1KUWUoRl6D4wR+V8JwxjL8iaEn7UxNTaSCKgB8rE8GYxo
s3pkmZzldcMxRpqTynhM5fuNODjG/fFUM9hP5GsQ+5DAPWGX9YT7knluxKq5DNFjrYoWa6Y7PFg/
RXV6v0V0NIGALiM39TsOzDZIcmuape6IfxTlblLNEJNHTwAhr3w3dx/uDXzE8Yelto0hmjfJjmQX
Hvgm0lVSMCrBMHq8m9NZxzR87qocf0ZwLIHnK4PlJbDo8XGJCNJiBhwgbQt1PbDd6D2TWVaUANMk
5p9KLQXG971KHdPBGRWd3gOGd0Fj1BRXUZU6gwyEmNL1L/kHayVL8MouGYrsP0eHdqCtNJ1VBpZj
dNLka6YxQokT9EjxBPIZMLsoPNKsyE33tx7EjzN2cAqecw+7bamtFtfD+ig9Wl8Shz+MVZ85Hr8T
Olef1AvQJEQ5o2295I6xA6vB8n2w6ll8r3f1cVUPNGv9Pups9ij1mvlWwLFGzO9MwOUkVFjYVAQf
df62lSfCg2Ufb8NbC868ng5f0SUIwIZmT5+FzZRC9aKGaZDvuiOiGzbY+I0jxHJfBL1Sq4RM/RVN
kZ81zI1O6cFOgNX5xSdGsjuxzzrucID9/7pBQ1zyPPWO/4QrHxkeOX9g6miDuxCbcYjJGXo5v2CH
M86aoYogDdeJzVDEp4K/9jHB43FqDjhQP0yF5963nOVBKQMiBBySIswdwHzBsEa0I9P4oN2YhvDW
QDhuw6x1O3a8Tj/zirloEYNKdK/CUFS5mCeyWGVi/MXX32qB4vnuBtQlyF4MhK3TRkFMO7qwnhAd
wgCE+vOmqXB9RvmEXFaqUBs4PEj1t04PKxnyyBsTyI8W46HR9Zr7frZYe2ySNs6lJQr54xXdTcIA
FUi5b9X0KcgnQGEmQpN6rbw05ItfCb7+zl4mntoZldYCHsiceNFXVR4eP34bDAE7WsTUs0MoHvTE
Z0nvsHhk75uRDuVcJjHgFX87EwWGIIOh5qMCb8KsXiuhe7t2vtAv71H1lMlWLzteAY+5BsnRjY40
HHJXHkM5FAy/vHA/3kA/Um+s2HyRpratK6jRZqMz8K84AbpfnadFivwb2FsvZEkmyqxAq/5LVHVa
SBVxV+nv7A11IZgz7DvA1A7pJT+GeVQ7eDheTsmrb4762cTBJbvfWpy48GKvNsiXVVF55b9DH7Ly
OenLwxJfvf2YAchAG2YbMv+Ee8LhEJNtCoNkAn+/VQdT5J5MxZkhf0pJppNaV84jph1ezGEl4Bi9
cDCZmNHDRzwH+xjT0GESlGu+b9juBr1I7LU+LYSEG1wJRRBAmpUrUsBpb2P2Xk7kiij8j308SaTk
ZnxfsRDUiVvC0eIwpuA9gNty8pYQSs0S5mjND5A5uFSKpFnVLf9gIA0N3iFzmKnOAtWMvVoSSAii
zEQzuTagqKKVulAJM5FtxpuGh9uIDGW3k7bb79RwJxKTNjWPXcOMlHw9Gl/cBIAazFVkVEIA1kMm
FxoDzgHtFBAcd4uGElwRxo6GacAx2AzvKc2yVjAf1/SUbH38Ry0pY1f4JEPEKJhqRij1b9PodBmB
ml4iTuxO6UERNtDVJ7IUE5UpMEDOgdEIWxCTlY7SBorrsc1ujE4QWuXnKP45uXdvzEW1xJ3S5cHL
soYWvwVAYpljwmIw3aQP1dOgF8fmHOfPexQ7LvPxbmLGaAZFvL9da64CQFdnp590fxnkSfgPuRhD
sWTI2Al/vJFp+HYWne3w1vcJOyo+P+TKneLs73P2d3cWIRKsSWZYiWyecDHBUj2HyqJi4AGKEIlT
ORLPXqdEJhtTk4N5GBe07EM9m1Km+IojODiX7pwN6NBm3Ycpyam/uAknViUZO8a6Gox/a0j6eWeS
XgzzorZLQHr3DhsggPZQE7YJ/ciWC72ZSZRPWWe8BnnXIC2j6sjFgsueNRJqhgUfVqNzvu8FADRx
PoIU5YFdvBJ9CA+JjToJcqDqJhE3Af7pRlZEEOWUq2Oy71A9etmphfio1PjrR/fhXcGGw3nlqsJP
7w/QjvooEhJrSldNHULc8GfBmBylDogRzEX/I/uhgUTqgs5pr3XahPd0J74bW5/m4WsvxS6C7pkb
ZIjl0iuva3abC2raFDqSAsjlz/LdkYoy2/9vYAqPnOZGzorJswdR+gpjQ+Yno739Yaw2Soob0Tz1
d5Gkn7NWMDph6cZAV2KdTFQ3IJgCatiKrj2WUsLIFV7TKIHIyZ5lNChtYG670odreFbMSasME7Ra
ZQrJQUPPxU5at4uDKzLGkhJKIgsuEBylSpSHJJ5CKjVLFBnrZZj54wXW8jZsjG3r74yAMzZI4poG
RM2+JGnYrzgpqrxJxmqVByo/b8qG/nIR+GcpOtwB3JzZGJTKN+EPtdQGs5It31gq2Yv7u18Tpbof
lkZiZO5HjTG1G1OLlBx2Ve3CHlJbQIe4mFJ/bbP9PZ/hlHAIfOfBw4tbJo/V0bjrmfFS5G/w1N1j
Uu8yCj2A85RqFF2b9GWKk+EBjD1oHdhIA2/xeuzqY1LAZr8h8uo2qe/4oANyVjcmdetw9MuxEfxA
aQwN12gDolnk9KNKaPVJ4q5xUYVGobjBRJDoUTiUfyTxgL5oNSz/bkjxcKZxLt3wxaKHxHVTjLI9
ozG+o1bX5D8VxLMIBlCYMt4pPoHYVNvVE0bbUAFi1pHqaFGwr84ZudclCveW8XDQTqBV3uMn472h
TP0faXxg9cOZmhMcC7FPZAXalkuxPvK+B8TyBaA2CqDgGlgP1modEUyDnRWK1aQ8v/xElRylIXxM
EbLpWH78L0DXRmYcN9BjtrDAsDHGCmy1q8x9ns1J6f6K4vJJamfYM9jeDPZur1iqgX5l76aJ5zPk
LcNlQTnEIa7M/dTjPkdEkoIF2qBPt+NZEnCqtQK/NmfsjNdu1R7KT713ZixuiQh9xrMzdV5dB82m
csSkIyeiDZ7GfFX+baUeFtZTVG67bXhhuXp1p1MuM83kvsVRlTrylU41lWcRoyZOg3e1EgLvCgm7
yj6Bge63RtgED3nNhFHjH1Tq/KL+EkcTMMyvl845DYi5QJt/vcQxp750nUs/0DGK3hcbQFHCjS/D
Di/bQqAVeW/YVWxhlLrthEsJZHeODotLh5SPq1HcYFOoBikRn4xKT0C+doRSj3SCmrNfk30CvvJ4
FNuVA2dkwQCpvywOpIe12QvexTBrEtXs7g5X0n9HYFj5KZyN7XrHTjn29EjRXhs4p9+EZsnnGP9t
zBrEg8WVM7XMzKSrf+y9LQADifyDOngLczNIFl6EFTbElPygtpH+vkgDsQg8Z1qIsNGVDg2iM1YO
C66wpP1NzPKJGmQA8zWiiHbble9noiqlystobeE3wSccKKZ1AhfZQg8YpHXBe27nxbyvSZQ+G7Tl
vPgPoYUlaNHc40I5dnbBg+a/s0QPZUqQIdpG6Cl7lXnfK25kjfOv8v0zFLNNEtTuwnS1scVvL66c
C6oeTgAXCD9Pllk5uFnNFacVewrRkfhzOAENWt6mzM+O7DwZUAi5/vc1FUY+emNT3Xu4P8ZglJas
4rGGlPNh5HX6043/H6qnOpj8ieRdnRcBJeHGd+VZxLq7kLrh9BtXq4mFxQAgCr+CdWXDqwHicBlI
sGL5X9iwkUyfLMy4QOLtdKqyZPFMCS4rGpNu/c0dGBG1z60vuuiDH3uzkLZ3TF2HZaqrjFpD5FKH
b26RO+NSRPfLLU2gDTPBc+KTdkOGJmu2yKY87DAmRYikT9NV+y0VgH/uxwuxj7HbbwYdKp+mCi3y
xGjmjrkV6qRtHfFyotJqvvYj3JO9EovGr7022pvO5uySLGegVttLAi/WkjylLrhfjKQmoqD3RRIG
YcCMrQGnRobNg497hMLEdtjhuxZEyK8ZXAOF/RDwFdcKyrjCczPDR0MFsFNbaVWKOBIehkzjrt0z
MRkwA08sTZFN6cpGOXhYvZ6KfwNmggdH6b3xPZJT0OXjee6i63NHV67w3VgS8Oq54JLXq9m3S4J8
kKNSedz617uI/othkmwWC4D9HPpfxXwdaeoFiOeyqYEi+iF4Uh9V/NLh5OpU1snrKSMFnlWRVE8z
I8mbUloMezTTBjIwTIpdZr7F3ttrdBaJEWzfyYiQDdxmQmDz8V3/KCVJ5KukHMwseSK3+ObwgGA0
MLmTa3rn0ajdla+rBJh5wqQ49bcVyWR0iFHwWtPPaGFblywFnmnHpb6dhJ3+tu6f9KPtZhokohHG
TtiG86lX8cTzMouxLbxediCFbEkAhcGlq9sckspggmugCioA93VFiXg7n8t8pUHT7G1f25TzQnqr
wuNb+Sx5Srjm8Xml9/H7OFvjCKUnW5ZnHjyNae8HDU8t06OWjVOqZtqMnHCjCAecmr8zcn99n2Vn
azbLp7MI5CYVldjXwCWzrazZid70XtQaCnQUV+XLvv0uTIIiEuVC+MeiIMMvkvN6D1jTkY7BZqWq
gx8uo+vBXu6tmwo1WaT37Co+98FwCtClxDWl3b1fHtP0qN7YXF5V917URYtYAHjd8rgX0/RUfLhN
+Z2gTraQY9YHpF8BCPuABX8RAH1wr9TplomuH1XN907yGQLkoxz40LaNvJdUG2ZQjU55s4xrtBV2
u4+nuIPtEHsvAry4VG4pIahH+eMZva7Y5z4qspNUlJ5pu/a9wFvqhpiZR/6mfcnOxGAF3pnzD+FC
ijLjH1dcdfd+Acrgo4INk0aAcstCKnEe9uSmpriv4/HyLoseZ7N+bAAYrSUOUQGnvfew2TdO8xxY
wL4zVOWc9jytloGfM9j4JsOyR4PFvwtC7RnH7HXRJJCcqweGa5XIPa1mzelkWABXMoL3dKpoRNy/
r+SwE8fCc2P8t299kFZ/RKCVWvhn24xjAP51NDViyMBTZIVLpvCD/1sum/bx396uQlW9TLOEaFKB
YaGZ2CkW19zAu7aE+Liy+FxOK4NDoPGk5JYwRrdOzOam05pk+0+mwClu+6AntBww8uFeX4sY2HVz
UNRwuKC/pFGP9JQrsXAyWHbF4J1iNZdJ4309hCAxdyIgbQC4EQJSY9dr0v/Sd46b0Gh6w0dy5jYb
kOOggFRFN8KozTFEfdIdPoRtEcg+MylJJwLWBFBsqd0/0qokZi5HP/xBglClsDODbHn30Q+kIDul
VKrzPR+VD7PmZu2JQ7sY3RMlByWNbi2LdwdqamVSgkZYuOU9wlGbvoMF4c1U49qNpGDkE4UFft0D
rbYXYEBd9gV3F4GXwr2BBh/pqjJEuOhoWWV6itO7Vg9UsTdXN2vCz1ijybIPdcBPBxCSvciIUWJ9
wgYr/NTJbQauFAMm+AJ5Vs3PnDi7zz3EtFzm7Mc9YIErf1QXNTUt+ElwM0zNDODo1AL8gGR239hp
8LdfrPUIxOAFgbFzUGg8p4OBhz7KXy6sR5fdmz53xa3wMLmwjw0yfzBraZWaSMZYT5xE/lm5hBqo
7aq7ElrTsVXT4d0S/ToSS32b6PkBLNZE4mk/SNTXbXHXB7JGg7tTEHpZz/sB7QpxNCctxTX8UImK
nZoMcobVitlPqcrLNhiLw9jyekst5jgLn+sacINvA9AAWVc053yEdgsAbdN86YEnVGJVArzNyjz9
Ap6l0A2SS03lBh9lBnYgqH01wbFz5YBK86pVV+rzDiFoebM+aw8PZLzC6nqKipHXg9G+DZAR/9r+
gPk5odD/F6qgGZ8TPenJTDxfJ2y/Mn8/u0gat/p1xFrNDu7X/Vc1mEoxsqiBnptmBQBQbvPe4zIc
1QIY6OnyvKjjh6y+N4RELdf1v4wTINxdQ767Z1N2RByuz9CpxRHU8QgkQ8MqDUjGUSvzOsXm3Jaf
wUyXnoa2eukvic0tf2uKszK1U5UX6d6bn5ZMLjI/A1y3C9GMYMzL9CsxjgsbbgA1F7hfUDI+UiVg
Iwbd0f2W/yGwOvHP9CT6PhZWKbnqD5MgJ0lEF0dihJ4bOZkiEj3RrBIwAsr2Ww34BqLLQ9yQDdoY
M8OT49UIb1Db6tykgn+2RhBNP8Xvau/8Asz+TSVQIob+T3nvTvXu/cjK9Ni0wi9ZTddlyb+BPnMT
RrNCXl47hWNan9Q1HaJGaJYBGf2O4k7njZbfTB3WK7OSg95LxxViB1IsP08yyc6RzjnD7/6l1dBj
0eymeWPnMkisAd8C/qI2Jjp7dC1fE9+lpRloqZy90BrjOHX4uFj+WdS4lpcSH2/B3U2LCLbYMuXc
4mnqukD8dmDUbjHOnjoB4kb/SbfSdo9pRYz1CSXQqLt2/wZIxJscUIWeLD/Y895vfzB5wFlksts8
wnyVJW7sr3zEClqVhYrR9KsrhJ8merGDzpfsEcbBU0smiaRZS7oNyIHxlA9n9bOpbyqDshGLHM0R
L5KkbF+tF0q9LNO7JLRBifQcYr2fRg+jGXq+z+LqFIl5Ifa9Djyl/ir885J+Vg55Su9N2KNkZEXS
tgne6AylPfOhTOcNuHSbrMBoi+vVRG/mPoGRAugutg/Q/uLMvm6XDALBTlLgUaGM3G54SLGXheWl
g9ZS9CjClat7qtwhBDQv1oAu1kVTyB1YsuorH3/IdAQdy7FtpuU82sDBxRlZno0Vr0us+gn5Nj/V
oaqYyAzQaRJsYXb5CglCpCKwSli3Z2z1ItGO0nBoi8pCouVq0AruqJh4yHzT9chtz/2uRWkYENBS
fof4EW2nJexgQXXQmiS0k1OcpkPMwNkV9xttFVvcB55usTWaf51+L38GTmC8Tbod+yMsD9BM9gwW
n3tx1POnOk1urhp4hlK4kes8Vh2wpbLKuuSAJej8C3r1wCB73vrs2+P585GtRk2/n8x0/4Ru8LZX
1cLTIy6NGAq58tQCR6qajfUKSbIDrhkH8Pe6r7RCnQ1Dy38y4wLpPLOKAvZ5wHY9GJyv/ef9seF8
NxKuBgu1PthrCoUqw4E+WZ6nAKNba5ws2RztbnO7IyCwM3z0EnlgnLGcThkyOYwkhvAj/YkRwtcD
p9ogOtGDVXHoSG/OH4gR7aybORX6wjNr8LKIPYw9XTFoXRC3jEd5fVqRupo6Pj1kTO6+apZmgza6
VxJyp/CBfcbeRRxNTvLNgMVdUIfttQQA2MXvXQI1zrHKjPXbMb/8u9KUIoDI7RSjtWgthVlFQj0t
rdd4NRlN1O9N0hHrcTAP6C0Rx4DC/N6IolwvMooBBRJgZ+vJ5F7WHEnfmzlZSFOoCMMZV0VJzlJZ
VFo/ziXx0RWr2lOIaWnuAcDRtlR2WhH8J6iEal+DcUr18xQSuRCE4ZjnTMQFa7vugYYqfYAnGZTs
bGlIXGpK66ORLQTWbY14+qdM9wid8mMw3ZQl39GYkitLI1UCrLFhTdIoQQW9oZU/Si3jKVSKFR6E
Om5yXNEB3iJPRVks3sksb+/jWZRHkeapzZq4CxK/eeSgapAtriI9Sanpk70VaDPG2d2BXCZRrDhT
pK91S9fTWXghAf2P87X3jc3i/PiOG/Ltho9ZbC+Y5RoKSlo47ee9giB/ZijLO0KgK+UGHXW/oU55
rgPWlzk+Mjdj5FooucCjav+3GCNm7UsN7gIl2vcTiQHq7aXKXLyuWz1SwAQCKJ2t/l69jZvESp7V
sfwj/ItQYdV29CAOR3SjKW18c9b8B03J4yWAIRl276FJara4LzNPRt+yFh08kvhyv5f1UdNQN+vU
sAqrkQwIGr1d544qm6iLpQahHIHtoD3bNaXC3ovwJL9pA4t8+dm8j6R90EkRJ636nMUdWTUvuK4R
92x3ddkzYuH+CgXJo9/vB/zV6BTQQVFHHxsR1Im1DwJu7pZyioQzCBAVbhPUi9T0oBEv29zndJNt
NEmqpjBQw01tRaIusarI4lbCv+USYvYOjlr42RXs0Ovrmponlb9gVUsnnTP4NIrkVKuOOUn0AQ2Y
M477MEG/rXxAVvIa4fMwVc+TzuZnucuCFKtp7pV836Brz4AXDmd3Q2xeCEUOwqASk4hxM8vOMlzT
mDd65V8k8QreBdQpXdRTmRHxVDsmV0Ly+T1jvSl+NY3nVtgAXbAjzvQjdrYYeVo68H37GCahcoj/
SaM2Qij72kss6YReL7WC1c/s6PilN1WjU73TxarqjNpFG29zpUaoS/r1ebhTa5hsdH3GdNI1zwtm
Ox4CAz8h5+p3E6Bd7J3k4pLyyzCjZYP2HHpI3xsVjGNqCnRSuyPy70ueP1f0chURHTaZ5Sa8N73o
NmOP03ggqmBzuStM79tCbzJdXausmxW7TH1rtHQFTOApoG4iL9AnFImKMdzvdluUTI27j4oj+saN
+89MdN0s9GkFZS8K8qo/T2kUu5ek9wdeH5rfkCOIW/QRkyyktkV/HVCQy/APrYngxykxn4UO+/bE
M730Ru4FaqQsgwSR5npVm51EklxkQqs2eQj9/bFrnXaVrQxvPTUnq6O3098BJ+NQvfqC08LNNdDt
DvvW8m7gpAzn924QSox1FZoxGuALwH6XtrbfyqQl21R1n8WjzXX2JgvvJF/nE9uHIAyZ53wEXkVO
lue8MEl+Hls6ObEMgefq71unDC8pH6+4VqZ1nJiINYs1VfX1BQe1rDJSvtVMtsM/UUkprtaTSP12
a21rekPgAkWqU8/jR6XU1YSZJnkjNc6IEYGYmzb5AZKTx/fcBe9Avt3TwBeJI+YoDz8pJt4wLggx
HY2+QDCcsyaTd/FMy0F6hTLEIrem555+fe8gojO63+yWnUj7TV3pe23wfukVi4r9tAcIdJDI7fh/
nMi3mDT/gEohY9rM2WtJlnpXwmbfYU6czJB8Gkm/nhP8YClCG1IKKkgu/BA7HqXa/+Ui75VXr2Ud
DboB6Fb6zxYAbGmHrG2ukffRHoQBXMrBFySZMg+PUgaj++XGrdZpL91I5Z2R5SDRzbnKOlTW5yGv
gyMoihkD0u5Ag21yFiTiG1mWJn92qO2lDAIeAJSrYNF0vI3cqmnxwISpZ1cWr/RfRe4g0rc4Efmk
LtCMnPBF3/A2UJnDyih7iXNLG0W8CRMQRIkb8PqyXwnGKH+fbcpDZrmfjTFrmEjeHNmYkIjMERm8
PwZy65VCPVfFSMWUiwtotXkksVyrcdr9qqBFiHwHPbaMhHYn+OlAzZTq7P1o65RcC47bfdvmMYpe
l1QVcKSkzkBrufbBZdW8UQbsdh91gdWZ0gQiK3fp/Hosis5YGKEiwfnHxGWM83OxX10bgL4ogNRe
tmZoWLgfgkaHfDrnKSYOeUSUXlXG3GDdvQHwxzzP5K3pt+RSm2iqeq1ueCsum7F2eyTXaKpmjuWf
3c5LserQLJsOy1y1bPi4JLoKxFEwHwhoOzn+aYhs+ir02qC4lEdlHxHVaIw7LvJTuCNBSm8QBUzH
nJa/RzZMPpQl5uSvTpTKFky2/+3bBy1m65EF+N5f0+YXKd3eYj+BQDJNt+DWpvvwRrjP2oNUb/TU
Op32CVVkKQjvYohXe003crCGIlCqv2XBpQD2SvpnNtAi+qigSeC1CmYT+DR2SINSf0bdiPLkg5ZJ
maxN1YAwcEcztz7Tz3iGMmfoQf/IEfYOnmtu/3zexlyH7OGckShrcnlu04Hj2D4KyUm2Nq6je4xf
CWU7TWpFQEsRgt/zJRpGmrLRWg12cEfQEzw6qoWAjfdikPnZS+pNhnSJiMHMHpMDA4KcxRWEjbwa
IxLw/hrcExHjxyRRXlhoyWbucfUvhjGhaltyGs6a4LrXZ1c7AQuf/xdMs3+E5Tui27FI9YTmXiFA
7SMX06VPMeneKl4P0Td2LeWxrIgnrn0DrK+33J3dAfaWD34y7RVyBc35FQtMrFzL7h+d2AjlguJ+
2lUlDcDf+nXvRWAhb3p9ujNGRA3naPD2Q5o2AjvSzGI7N3wbcRa0AuJXFxATov9Faw5v3sHmZsYT
8umrcmvKqF+mRwnIghMkLcjYiTJ507mkiMXgRd77Tde+R8vzgsHFVz08Nn66cz9gKHUkMZabDLPz
JaAdVebiH7Uv9N7dYTI9SEAL591PtouD6HR98ofXSIv9umjZnMG54Fv7uNRa/CDZyBTHo3T6Ww55
eMY7v8Xy6M9GYCybrkhsPjIB5RpA5JmuLsomMj13Fqgn9YvkFpD4kL3oM55Cgu2l2gfw1WbZsElD
u7E3b0pK0+6OprmTpun1QClgZ8MOu2oKHhn+KvQImd2e6xNmcY1z8Mc1am4pIdVKhQKIRi1qqy8t
prXl1V6yqe4m0CEjwMTvWOlKPvjS/jJT+an2y2rZtZjzKuX7fpRvdaPOXrCkanWlJnveLNNItVRZ
Ka57jfD5ABC7NN7KKdlPlzk+/padwvD04sGnhFWPe0U/9deiYupf9gelraR9npw7mXBlJ4DRfZoD
C+GPZxdAV98Q0qBi4xAdLeFeAA/mXFaA/XHlt0bKcISGyQwoXDrw3GHFyH4FEH05e1GbprPM9wy3
vS7Aso5PfKDQYwDwU1OuaT4LbF+Wf8v2GOmgnzN8e+xgoHr4lCq3UNSvzjjBAqTVSezmdAHNhndi
i3uTvCVB4J9+f8x3i+ElQlWbw2Qci3nfblqzM+x/CuYU3aViw+9WSx7iSTfqrN7U5ykK/0UNSIcy
Ow+2gBIT9wuPmUMEXrNVh3qVS4XEfoH9wpHCgg3fWYGyaejxkjurej+nEuR8MXQzR0u4CI4SDidx
+gJ2Mj83Bqh59GjJqLO4MoYu5WgV7iXO+uoCYSF3gCxypQGTltzBtaoTHLo5qhJoVSwBSB/pSw3K
Zw2a54ePGk2/pYfLFXIPi6xS/EvKpzpsiEbLvPjW4jnYFmCoxOiLhkeeEuNvSQCJeO5A6hijPO4B
yLDR+fbTJibLNxYf3B4j0VI70gm7KLC4ApI9E7q4GUMm+bf5zG3yCRNivED05uNAAodtX8I0UGct
+Ky2qwnvlWLDrf7+C0gueCVT8cTHFTZybmwmOjy1K9fsN9MoBoMLZhTS4YGlk4OvtwTdasFFSd8x
bsuCAa5omdn4JkkEdQmAhy9YTsp6BwUOJoYGsr7Hj40TccTQL9d97LqR18P7l7QRd5B4dIvt2cg1
ayKBEavd6ig7EJbxUMh1N+yfvFmV/rDww+04DE59vK/64kNK2wqK7EXej+VoffbTqPlVm+2LJ57l
uKrFOIzxii2FW6EiPEeLB/VuX8AjIyJFY9GfwgcuOLfh21de3eL8W1mFoAJWjZXh4KG52cox4Wdw
9onZMyIwZuQfumVkW6L4mXK3fVCQRyMxcCofOsOqZ9lGUe+fXLC7XZhg9mivFVGPDjWAZzOSl+De
LDjoQH2yDHlZH0taXkEtfimT33M6D/Egps8tGhOvCgsbttoTiAhW7WYZjTTUFZZZpCF+wArbA2Fc
ufGO5LElIqQM3g7iVbY/TFrtHMPJdcRIBbFGwGHLcJCmfgxJ2zgk1/D5KtfVEMxQhUYkaxPYVk3I
+/xMzkkbtAqCzIyK46lSOaZyMjuGuGylfl8wCg4GUkN7HtSd8l1TIkE1KlPEFoiwRh4mXvpUr4Wz
yiHzuAiE1HXG+HCGSlT0KxNMUG1+VrleIgJNZI9xUy59FKvXjUTMdn11S93+yNVkxX5xYnHqS6gS
EtA0OeS+0gXNpNtMIgt1Qk6M+UJ+KlmV7jvENjvJkRWFZdUhA8udeC9/TkSEdQZHe7l03aslZfxp
xjpHfhV861HrcT3TGQ9t5qtIg2YiquwoSNfd96Gq7GUIuza4kA/x4SIr4BSetmFdFCmp36svwtE0
Eb95EdHjBsgA6/jZIiQfmc8Oma38HS/VaNnQfOCkOmmIsPbqh/ot7h+6Mpr6u0FAsxXqDi9gVIs+
G4ZwG9rfN1GXiu31KjaM6q5BM4ssZzPo4g2bLT+CxgdbUUJIw1iCNjckixFtXK/utKaJfUbDbhlg
IGEUS+JTNKczjBmLiI+rtCt9AtP2Ko49YhX0l9b6Z4mqMrpZN2LxKw2QUeEP30KH3S5zVZy4SybX
gweC0Sc5WQ91GsdwvxTqCQCWbvXaZ0jwk1dgX2hMcQEOUXmHykLmLK8gEA0vm7V59ZJ8Sm5gcRbH
s1T4u2Lc6EpBBM/W9CwcfqE8uJWXUeeuKzLOJ643c4gzjdPhVgF7qT+I6XS6O1iqiVnY6nQ7r7jm
mB86F3P8MF1qkPp5NuJLx+77eCENeaLPzIQs+CKtVQFegjLP//UcTawPCJH87Z0vxPnNLF6+Sx5a
dGbPAlKSiQu5HGsWlK0eU6dpEyuhomVUs0J1TqO7AIb9raz1bZswGY418H1Kpb7s4tYFKiddzc6w
2+CX2zddzNle9c4W8Keuji577tfYsJb9KHQiKc7HVvEtFxaIjpf3/dnxHuOz+2t8REabKL9nQKPo
cPHUl5WWKx1k31wUXS9vqwGQwcJJqDffTnKj9MBUte5CvLt3CSwJKiiPY3woUX5mINzP3IWowkB/
WeMOrWk6ThROmgwmv40GO23JrL8MJuZDAcIvzp6scpvRI+9r1uBZAYPVKEtIDtnmsGmQZcvOd07H
54VGRnKl2heLCEpqMxU6OyjSVS4XMg4E/ywsXYwxTLWeZhpGRSJNQumxSiE/DW9SyioOHYYZoch3
7XsOtcrowcIkW/9Rz+jd0HG551uaD2iwKUhrSquyf/sHMs4xcsRw4a9kya/YBSIQMnf411yj70vm
Hqb1FSDGyNqgCGE505Sxz3H258D4PmT/UkX/2BdH8JH0JFDRGetmSEguV5mxKaqv5BoAVLxvPG+z
rf9Swpx1dpbD+rLS/3r901d4uLBiWtonVyAXJcldh0WV6hMxH/uLz+FMlSJPXTO+TlyGQql4RxU8
AO8HHTLHH9XeKNFVugvrwmpDM/IguXwjlCVYI9XII3DR4Hvc6xcfkoYXSmvzxg9C3PMR4a9Uz8lf
rv9lemPo2srMqI/BTgtStnCVGgKFgB4tyDWG20P6VV3+RccOPoSHIwKFt4Ozyp/QQ8LhW5SblRGc
OrWBaglp7JPRCeUihgMn0Vw6unXbzolXPDCDnQEfEo3Ss2VM3RsVGgOU249JsSrNdW9fve4++yeI
o4Wa4dYl4QZs9KOiSEdCYFP1G1F+fTDQIVZCOzeyJ6nu9nt/ucm+ZLUtIZdRKR0NhQkTay4qpELy
YyzG/zdF6Zp4Quqt6DyXMViXsZ7wFa7E7dsJgdcOiJioBZCvi33MOyhBxEdoqK8iiHhtm3ytAoOT
kkMPfZqw8KAlHHlUtPOy8jjmfaF53TSV9nerKgng8OpdBJPVCNQFo5jwHTOG6ujyhSb1UIWXzgIO
l9VthlE591UhMoVkOB0IVEzGKcmqYH3Qq0op87yM5eED8vVxHbhQ8ltGtPyjoxpC/e7BkbXdSMke
QkXyAimzJepKzvBqcajCoA7uznL2JDxjzUB/rWpQ+IAWy+jFA2Eu/k7OcIoUBZNqjqN/wxWWMVCC
OKlJCEWTsVh1uYKDhBOCsd1VybvwhdF3EZS3dUzMLUF2m6VRleIXfD42mP8qdHIbAFQtpwBvAvI5
gMpdwR8KNLaTiaMUuutpSuAZ5i8O0b/0IGY9GPgKntq8hjqX5IwB9M41c0IxtWgi3XRrjlT0uyX8
/tFpw6c0IR93eSD8YVlRBvL6F2NFhNXOyOW4MgZCjsfPZJdoWt1ijkHfdPefAQhW0eNwKJFchSWT
JyxKMX+SnHNxiDYe5xE8y7ClxwXfsYK4tn3kek3W4C4NOPcg6pXkUkjXJaPXq6SfsOh2azQ49Z/4
urYPdMzi9BywWoTOe/am4vTrnPITGYCPrA7hocALdkZXriapb8Tb9+MM+hlpF9xko8IjO2QculUO
Z9oHjVsrteHkutnRw42hSJ1JiKMSC8uiQ9+qecXM2TyjcjjsTDnzWF6a4MrDy2gMFhpoL0of2hcD
vTIWQeSb57saS09oi4a6tWzpWkiY6lJwgY1rEyUtn9+RqZhnQrG2wPYDqit24V2xkxzo4adKykkS
10n6fgqzPmiLnKnaW/qMm3keWTzsOG3GJuFwe44LrRX9BjDIOt9TxSXpANyU0f+sPbqkNNK1Iec1
M+hMPA1AweQ+x7hg9lb5L3vOadh4x91/5yQCXQlBHBhBNRy1hOXpRgqt+vdL7Ld9m1yvpx1rKdkl
B3b7gHE3EYKLLXtWDmgxCyOOJsHdxeSPJwm86ZHlGYkSAjQUX2xOruGMggfUW1PFOxQt6fvQSImg
+MxtTc3sclvH7WdC/3NeILltwcUt7QFsdQJAKVO4byCR5WgRZBWq/jQG7C0HXlUXM8jsrfn5tQ+K
kJNlpZ6XZJUSCRj+ZOI9zUZiALC09tYOSQMe1xw0cDk6Y9e23/utCB7UuqbxbNUmTgBa2QG77nbJ
zg94kfcx7xsLUV4ipjC6f4ROEe7wFGzkzyuBEtDaM5ba8+sAjvHuQZXht4Otiv5sx1O/ufrWUy7Y
rDZ7xBPRf43B3ww/KJv+obgpByk0G2RauUJ2rz3b/pX4jDhBXW7kc/uOmI6zM54PN3vnJQLW9bI0
w5afzfJiZT7Kr9uUc74ERmllbS4laGVa0dc1xjaV5qmkoj8ando+ho0OTSPNEwEx9JONDdYfGyug
yuiD2abaxmbKRONDkFF0m6QUXXIoWSy+f8MHaQngu9XvexPJ8s4pI9quy2oQV37qkB5qs8IKx9qT
aNAatgbdT9NDlIOn+hqoCkrhMQTvsLhpwanIUBmndWtT5IjiqXGU53Xdpd9lu5ERed2N0JAKLGzl
LSX2E8xUc7stwdhhOpbW+4N/6mfyoh0lgMafj95DFr9Pr0yWwdv1XLW2m8ODIc7g5XXkd3lsg2oO
GARLzXuvDoX2zrKcakamzFERARbiVZljhVpvypfAKy6hhIx7EsbrDVFvgYKKXdWy0mbM2LDG1qzW
KoOEIzFPEXMumV1DZ7pvDOstJPZu7PhxW4IlyEEBF5dA7l5wAZrGhVTUDfW7PfJWzJwrCW2rLP5S
vfM8U3y7sclmLoZUhmcfODPyc4eX5OvkIuSKbNCYfzZ9saz0HzT0TFbDnXUN5+F4XFVc8n1Od6F3
SPqvX5LGXhzT0m+fp8yhekxEig6RxoMK1YQacGq7Hj7BWRMguIRlS6u4cLRwmpz+9E04ERpoqjVu
FTIDcVdMiIkjmv9KmDrOCDCQHaUXl6k72v2UCxFaNWXo5R/ti0T1nfSUtqn+FtnnHNOkQ1TSaIhU
080uPenk6gVrHx0M7WmLRCmsnpd4+oeYv431pooknGhE+SNBO3EcM+M8S8rtwmy5e3zl4Lqs0yo8
ASNqGOhTeTF+0GblIPBO0dTBU1GoRaR4snZWrRonC4YT5JdrkEPwBXrII3JmyhwoNxov+RIU4bvA
h0CO9Xhd+XYufH8thNH2bczoQO2w2qzYcwBQMEM7GCdXRE6S4GFkX7PiiqqkcTYHgHVFe5i5+82Y
YYBs9lH9J6n2Uk007z9f1oYdKwd3eFUiQyeQtQMzhJ0Z0Co4rFSF3gdrvJQDnkRimLR289DKjhkV
OcxMo4zdxZVOMB06pMLNBB6b8Wwlw4b+l7H4i9dBjiFMR+/E1kWQO9ImZqLyRV97c6rFjTuKYgEq
8ey6us0HFK0PXS4BmWURPrFwrqhXXv4AQFTroQqoDX/+3qb7e8gCzec0ys/HFzgcbWGBE6IWjI1V
l4IUwrrd6DQwl7iJyTVj04Pwk9EsxcWNnf+5xVu68wg4LQrFHFlMw9QYzFGQQYuqC8OiHT2n3fr/
3L4kudYZIPg+JJA7labB2/WQw7rpsm2kkcVnoDaXL8zyPGXwJBmcjbNl+tYe0Uu2zVjZLuT7HZC7
O3IDe8W9iYyvLOHR8dZTAKVIuYvE4ZbfF6rHgJ/nWsH36e21CzjvU3TnqfNxxMaaY/r+hpWdix63
T+6ZxMLXQohB+K0Wa0auLDK8J3NXbPobxMYe59cVoxBlB53D3WgyX7MBUAOl0s3EJRV/+jFO8kzL
0TsESoohUc/sFJpBwjO0Vu4YKmNFfvae9zpQMqDmg22RbBBfNCYkKHmMzBOX9ihxmmhpoDJBkP+u
xGNuMvAInv6/Sk1OvZBKVZkyAnZf69iMXQhzoSLfcIFnyp56POIq65tICfoKwOI9zLJ4N3l+BwBm
FP0sdAEHEPfVfsRVrqDuMBWX6Ytv1UlE3Is7WB/6WfzIWM6hVbqwCS/MpzMnOE6a/S1jAiWDnvXM
ib9Z6o8+Jk1Wea/CwTuzb5fuouMnlWcC8hJ9ShcEszTJ7FxuoXWKOZT0easIypP9gYFfrefBJ2kF
+d9g8VmgItdFSmeUVSrLOPg/VLHIreFaMwUxyDhh5VsyuP8JyWj4cPEn8+4B6TW0weCRsdiLtsT6
3jY7sY23AI9rfUdEhpkAiRfwdyUXNBpsA1n5APepEJsptQJ4bPcEyjTNRXUc5oOA47xejys8Hbd/
/ycEt2Nm9RcWEUL6ZcPOcBTK416bI9ExpCb9aOxbmaFnZgQvuodPKfVGsSCUmKDix3OYCc1wmU+G
ZM2euj4kJd3TdLQ+PXrdoljiSu6e5jwAYlS8+tMVyYYnDnirKuY9t5OFmCVkf9rR1ldgPYbcPYst
9C/HSxttiWqZN6weVfBJV9b/n8YFurMTMMu2Dan1GWv7IG41LjPuSN9ETt0/AsP/sAtvHKg9MRti
D/cdApareqFYfrKGya/2gDQe55QV+eNOSBRNcV0aRGoaCj13sC49dgQjQD+MjmmF5mAMS7FSKkCR
JNT0Q6K1XtBNiSkgmyzj8MY3CwVQ/NrRHXjMA7mb96UZVp7bFJIxAVX1uxWDu8tX5sqoSvmIGWtJ
iQ71MNr05UPLwNBd8/gvxcPtFMP7Yn6/wNgsTI/OefCvamNvjTRfw6Dvj6sbwsT8M/5PXAHsVhOT
/B+CoFUpV+YtOP9xdgEVpnxMAA+JKp9DVNxvBU2sBngKaf4ETaYRpczGLyK1verj+9srOjkE89hw
O5nXyG5UfIDXiF+nFVTu5pHj0jnFaPG38xHPpJGu1f5VEhKwPekGCbdMtsfqYO8gOYcRxqQK5FEv
C+9Zu25rggbHo03p/GXRrWYSk14RaqDm+5TsFNJwzqR48Iw0Pa4xc7gl/ne90lSu7p99Krn7KnLM
mqfnvSshRP/3daiXAYElLSSl5D+HmQp/BsYqe1rlZyNsCjvtM0o+ck1bfmNvGxnCM34dIl9a1QB5
HDYjwb0x3do8P3bEtUYiNbuA2beHXFMeLPZG2atcN2MBFYlRGdRTnypZIxob/fyotqnADHG0COpc
xhjsIHqexubJMIdyllQTpFcGVBiEJ7OmwV8eJ1ZJVEuV76kMGz+KWfJDETHTzjomaKcQkbcrYb21
VJFb3WwlpbZaLYO4pyuCyA0z0OIYR4q2rjPJhDH49hItvCxZ4mU6S5gLjgu/vjxkaiw3VzexVGgu
EuUVDnAS9TFKj5oD53evBJZhgQa1X9g01qayu0L02GVLuKyusphos/7320METsrIwz6lVtLMfEtd
R+M9yepM6ETws4qwoj5gcOPV65w25Usid0YkaWQruJig6zm7a475fS5mZmo7vWNsplJOGelrQ4mR
w88lOHQnM2OtVnGRxgMtg0U8Bm/1BJgK+0CLgVSp2kJCa5HeXI/QJqS78yf/2YT8jy90uPB2C5Nh
jyieOqCU/kLIQeEfeOPkwvTF3Z0K5+9gyx3NHP2oVz3FoqOzM8fggRJcf0I/bb8Uno+mnhSx97Qp
b5OSn6CgNhuxn9GOG++57j5mYzYGp1GqJ7QNeA8Dy0t8NzLDUbh3HPT3k+8ppNODqV43sdAw9N8A
HD9oBaXz11HG8hHN9wfPcsWZ8+04Fe3aSowwq3aU4FnnDnFAs5etxnzPeRxKgRwE+L37dXepty9L
yjePzJ2IjAmCgILd3u0OpxuLiMZXkksQ32N55/ywx08LE3eZR9Vj7457DjFAf2OSiy7Ycbpnizxj
CI2Fmo/kLa2i1iP8dPAIz4gSLi0hfFC0DcbrxjYPwSvVtfNmgta8rGvF86MvT1fexFhMacpEW32f
PgHUXRc3bz9DPLUuJQGset0w95oFEr1QhXCdB0doOn5al+vhNP8N6H20Ui1URDiItg9r9Shb+y7/
TMuozqctiET6Ehg6YyOLbYsOXxfENoMSyGvQBzoyuSkDqaoIaGoeeWVf1N/CzsViPPYUjSR3uGE/
AYtIwZQ2vGF6bQ+2fQoNrXlszWMF2C61uHiKZizmoX4diQF8ClMsXdv2WVj8IhEvhZ4MPfo0gcbt
M0QikdxzEOrUVeWmDBtNjS5uHc2JjL4rePaYhejLLRcMSX87YSqHYxBB9gHvFabAvqvR4XSB2PzS
VLalCTAyo5iUEbYxjMawPACYtcri05JOdVuteRwQIcfuP0HUQO7qqE/w+o4c6Dj5PJl3jGrOTc0w
2tnyBs3SfJjW8u8ceWHuwhpRu/QyTxAYko8CxfeF6uDfScRNh8k4UhDGOFpfa3PlYCrarII6YDMY
7D0hfg+rpJo8VDXSDYc769Tvr2aE34eor4KKo426W+8uqllaerX92nNqR6DfNvoWulZDAPbzDBPO
lsdJRoshJXiGjUYb4f9M95OZ5SBJawuz0Ul6stQccbeZvWDBK1q1KaqZvIMkZbG2T4liRsthkrOF
FOjIpZY/c+brUc9VTV4P/hqPilowCiuazqhgjKWKYkU6Jp6mWUql7W2Ak1SVIGYRTZ2sUStoy2qV
07Qt+7KdVhgrraEfDISsLjhM0b6CMkeWG80gRoU0yDrkY4Hyo92g3GKC4m2jFKK87OTSe1KsDEKo
YhNuDUCeWpQ+oNn6tQGErlZqwPfLJRunZitYYbeFOdmbNUsVATdiA4HbJYPpLsQ5hykwxYxIysGR
7K6CxnU42vX3aUI58JEHmzVH61YlrPWAybkep+LVOmT2Lk90XrNwYW8YkiKi5EYFFeVty1/btbJK
NJNUagUvM/1z2U3i95N23L/ip+2zVR3q2DnpfVWe2ta+aQVjjXmeWT1TPHinJsQ/G4+hTtxa17nL
rClU7UUZYetycOuCLLuYFDxTtcRIn2Xk2ECDYziqDhhcw7ijLxM97RkcfohB3I08BXU1d4IHnpop
+3lQYJYeGAiCi7bUUw23PrSGjO0IOVn5dAaEBVXEGjPF0CQM5GI/znEssT7LKI6mDvIcDaE+JoTh
o1bRgArpxt9imIZSuVSfmDRS8JF03t9yU7n7lk0PWARpBojOdddc+Pv9tca8QfElBPgAImkb4Af7
Zn502PSHR/Fb7fhS0O7rzLSDjy7cnnboX425zJuznNnKFrD6YVVGnw8e5a4jENc00KLtnryPtP/A
qXb9yexXCQeCQFqnXlpCqUKHljmhsGq3pfq4mVK4StqRnDtZaGQI5Gc8YUObncJ0M8GW8FBwHKuA
WsGeyYymkQTmtVyptRI8DHNb1yzPaXvwlHTV8CFeBbEYI8fnV3WtQrHFscQ7KROfgHdPAI2a5Oiz
0OI5YjSV+YQEC46rsVBWF633Zti16p+bJUvpXHjnZxz5d576IoNISLuXLFpHRv5obsqgX+TxWBem
WNqgEMU/RR0fXOsBZe/CY7fgCHbZDLkuvCGpg5aeYNyv7ibLt3n0SkcQ/9f+W2CGAMDRyrpoSv0C
5BIEhRpaUgdB0GdY91TLF80XDNAOgP/tAdnR5X1qjnn9uwE9vP9XsMuy/oORWzToa/BrfEutu+Vn
swqjVEXL/3FIqwo/pDKEdVEcgw080cBNu3sK60TWV5Wc50ptAlB/6wF/zNr4TfkxGwsY/4W4KkuW
9+r+lEJEsTNoRdwvCE6myBqBO/CTROlhWyuvOU7YLM4NswRuCKxpfGF2BAIY9z0ApP6VJhFH5rKd
94UpzQGvQFruuIumJgU5Lw5vgeZHD+3SaSeNe5qT8AIhv3sdh3KfnKN2f9g+kPJowZqDGB7CVeoW
F610B9lMVOKSVcrN83i4snHtIzDzegb41APC1idLi7VoXVwz+rgFdIc586Hte+QcTFJdJZ9MhrOh
XGzTJ5KCG+/3Ch/CoCMvgq4pPSHeS+5ttQqLlS7xYvkYTmtdGqyDExJqDlY6K2c58kAKJkiFkMvf
7wISb/KNF0vB4yZg7ltOaddzhgiwc57K+yhQBBJGKppR64EJYQUUInQXk1WHIn5m+Nlek1J9kWrI
nAbE2fiHB8aW7OKkApgQhxMvslEYmG7gsrlWdufhSF3H8uUGr9zk+tB7yujRbkBuVG/1Lzwbyeto
DLZMQsCgpMWYhZ/xICi6sFKRODCeL4k7MAzc6+2aIwkUD+ZuWUoBjF4iFGoTd9v4f9XsbLOz/7Kb
GzMNboU0041pyVSlY9RAGSa+7fvJJ56CUUZ9PTwABUEw8AMj+y/k1aIMmar4AYkGP2QMxT0PJIbm
l0BgFcOHPr23gB15XVgyHETO8lsu/iKa5nSOPCVfRb7hn+0Njped+XA2UBr9q7GExC/jSxHA8tiF
HICB/OYGRUcwX0sQ9VV7TGuTwGORs9BXsm8/x8v/TxwwIeTSauqNv63LCauTW/e2hce759pBAd+9
n5rKxYvntdJr/K4Ag5pOUXT7TmGJphNlGffentCkAzT1llJESKqWLJBuGkPzXwQzX8x5VKxZO+Zo
K5EJw0gZZRF8z4TasqbPpbaHvcWhcTwU/AiYtMJaE90lVd707A3812o10BSZY/kUyYKA0eObMzLz
nZ2H/xYKmo5kxz7oh0sk5UsKl9TpidVNO5rt6iP+/jsE5K7Q70SBvr8Damd84OMsjYNlnfLHIu6N
sghHmmud0IIQpSO32VybrVNhj8GeTRaI6HXWajaxAbufCr1/LdPn5nhusqzps7zlBy8OO2FSS7PN
zgS8uTYzT4DE1YFNrLCzd45YLYtg+4YxIvdasHImGkvv4SAXq5EN6kaQic0Ya2iSUpH65iQjA0Kw
B73MW5U/68+oam7DmM8ZuzZtzZScdBL/gu9uuAqRYlYCfFE2v17Y6kUMbR2lc6Ftpi4yfeLDM2gj
WDygbKj1oQ2bmXc7zVSC3RO0CDD/eqMMiFYCq3vnxKY2novqn8/JqEqSPJhlv+5Q1reghW5lMQdx
jpU5alGVmHdLG31mDjIfDnfni4MCv05LWSUPvzVyJS4zYEHbi0Y+N95uvw8uxs7hkIOPbUwHjt64
UQgJq0pSPy88Oq6dTmu6+zwUAG6jyY6jOwmiFh0lcGKCZYO1MLu/TpwvsvP4bFw98ru5sIXCKtDG
cjuaVBeJDRz9lXv4rrZrx/iw0dow0w5Pj8z0byYWKTGyWx5AVSKMmLRP3g5wsZbdwwiLPSLy+60c
Ypn3nopJXs9pcEfwfsz0PFCYPNxuQDrBuXsFMMkmKYJ14+OVNo8WxdkbQocV7BBbwqjlIbkGEEBE
wi73NFORqHF/FlWWh8efuFTaHjy1JP0jO8NKUqHgRKcCzsFcY5nXIMChnYKxLTEQhFJ31OWI3Yz1
MV14wFG03QXxv9yENu6pIx+AvyNpv/sTHiJDLNmP1zb4ooiUCkcSH72j88W+9uxBeH8YpR9Y13jt
m30tn1wfJGBoJhQKvLrcQXOiVyMQIngJIDJrlBMQuDWgiIZf08yBqjAE1iz3Q1ZKgfWTfoZiTJtO
0xGbVZR6EMBLYWk2t3cSwePSvvZoZbJFCVR6EB/2riEUlJsWOvM7aaxSRxMGBiMV6uRcNC5wUs36
q1snMf4qKmEKG3btyHhDmDmWYY1pB8r+duRp5WDHDbHg3w5137Of5THfO6aE9gQ9Veu1s+Z63nsO
fpLnZ7wJXu6EEG+LAG4ljePVEtV0fciWEcR94swDkPHSD97sa6/ewQU6SUfR0vXlYw1OUfdbuVtD
efSuEFQE7vcXQJnR+YrgM2OTSWFtjOQGjAYya0JOrxZdPZ/+DGwaoTcUkM3HMsrDdoVR1vXXiGyu
pqIt4BieVOIp/BXASj+gopwLbmHMQ1bv8c0fuTgJ10Kp9uIyVC8meqFPlI5mOZdI5XHB4yLbtBn5
P1Uhid097ugujT9PCxTycjicv47W15enDO6Kn9dhBTTjAgqQnVSRgCEDZ8ipo3M1OvOMb5uYzVHC
qj5rp1P9ZRSfVIDBpGxgnYBLVxJgSb0InhcnbITdQXUvNiWTXOQAVMQehDYNvM4OMolUW6RjStaw
KO93OFp/PI4DdDnUkb/1M6Vhg/FgpQm11Eai1t6PSUoM5jEpoBLR2YD7H7pFV1VeIvHL35x8E5IS
GhAwebOFSHo0w9j6Cwm4e11+nDK8qaxWi93jxeNAnnhqFgRqfF84WiLdFIkL1MArtQPlY7oAO9Xc
rYFfyFbSAIeQZ3bSozeuContlgHETFUmwYkQsBRdqGlcPRCfcU5UyiUQSifxLYbDaE/Km7cJsUhF
0w3DQ+SeUn0oF2pmtw9las/TtqmnaH+ViG4B2LxOFrk8Gwo7OpdHsOVzxlsXz2c2j1iKJPLX05+Y
sQa3TR+EhSWwjKES71YFGnA1cQmXKmUJA9xw/OMH6y41szf/B19Q3w6Be4GRNL5K4CIxNINe9NMw
6WJzRZ8PFRCGWJHiDlag6pods9IUBPUsXihSMC0lgg3oKSpEtTgsZzaUzg/xE+pMISEcjv2EvCz8
nBQnkB0eolYBalPv7HZmEoBAsfnKOIxaCzW0ymhSgxyP7yFo+lMCbY1H4BRPP8FFRXmuDyrv3UkD
dc1tn9LHP5pLSyFc8LYLY8kjBI0vudSb+5Vt8AHbJsuBAxYfcVQWhu1bPT2SLqpzid6tvzRjoBuC
GR4k5/iJkyEiC9wusU1O95nW7Uk/cC33Ap8VMEtkhar5V9E1JD+0XtvQInvJpeagMqHZVnpzc+Gx
jnluqI0lvcTnPkFSnFG34D5iOPbV9c52gpNwJWzUIv7EUcbG/663AvEvk9Wr4wkXQv+9MNbUnj7P
b0CO3WE39nAaV6h5USVwxMO5w2MTqzyK+YzPR0+Gz8DtxuzzDyMIwiwP043EgqItsMGrmrjHOOr7
iLOcSopKuXOAS5sTZkf+NAAORC9LKHP7WeRiNRz5KZe/hIE+JL2ACDhHjC0tAAhjdtXTol6JvD1Z
Wr8eBqRGO39lGHEvQnZ6VVVI+12/0jKWKU4BoQPY3xDK6Zi4428pj7++hWYmIGkenYzRQ/NAlyaC
9TqicGFuIVm66RT2N6PwvKWdLlRwAyydcjV+yPJuuXQkHAKHjpWqFu1ahVgRwEO9yKhg7SUm6/sF
CjhNjCSd5DSIjuqiT9EVgQcVZnSsz74mKPNq0uzNDcxVseS9n2/sq7FZFg9dYzZ2jocefNUB+nmF
Ds2knmswQhBho5GknxVge7Mbcf1JY5jXYVCJveCD66PesFol1+u/VDYClhOhkbdcrLTzF6yw2O9H
zYvNFGbnnx+9kZR4UFIwqLbUzPGMgYZKNuNj1sR3Qn2i2zxtkDGaP1im02cnfXjpAGpqs+YkC3Fa
/tHYgv1ruwkORrvQzBvEJy/DPBJlUNJsx0c+aBcrBcGRPF+DjoaH2Xom4eCrK/bIU7jZ1lXfmw8o
AM7gNR9kAMi85F/sWKTHCZMaI5YtOz0qHIhhUeVPI8xBCNNt9E7acGJD0JrLTlSIY538a6518g2F
N1GwPxcJnaNazSV8Ww2P6ReX2r1G5xrkd3AyCb+x0kHspbL31CnLhYwWmfy9b8uX/Q0i5LRdYLZg
Gt80rVHirWespp5D9q9I5BZQ+Qw2CUbdNUNRHSL+L3VlPJ2Qw53mFAihROblPt0trN56rcIEZZyU
kiPRyiL4eLsvZMSBlTBFQPifxuzCXQAtfjVMo8xn2Qb33xfsspqAETRJCCt8nj4J3pgdPUqjpCiN
1TMyt+QUvC26sFvsbE3iOG7QjLvctNKDvN30/MU+FYDzq2oP8vn83NsIaRyiImT6+xwOLsR283mu
ZoYNW218EdsqCM8uzA9NeTos+MJ/07qrvvhuYtFAZA2WxLUdadjVoXP9YrLb4cLVibBpB31vk2oz
T+7CyKtnjSbBw94/KKXUYOWHEQzM2SLk9UPoC+SCDhOy/pMdQTk/IXo/10kPcyIUF5gDAbPnGow0
eVz6XbSZKESOwlXdqkmpp+QKihr8nMPcnZoNeHQQJCxzRjRLqtsDxjfc/1LYkukBw60jbOe7vR/+
WhInTLx9fdHv3TVcf/ljLikOaggUTbxDtAnDq5UCd2/FYdQ5VB1Vg+qjdsP9fxp+7xQr26rjNZL1
w651UKJUDjxrcVIpPe3KuIsNQq27nxXDl2dolMI/ng9B/zYftcUxECkFy7uV9m6TBTNRVC7nA4+o
RKT1BLzyPaMj3pS6bH8oEp06TORMQN8Jsq2/Ha/A9KheHRewjn3NRDKki7eHGBIkAQDdJP3YYIip
xBcLeMvlsgj+1c86NHYz5cJg+Js5Mub32iLhb44yb4djyb/7aopPU/wCR9MnCJdBChTbraBzuhHK
bA95Uy4CUDfEkvb6HIg218Lit5LvfzqhLK4OidM7oP9slXbhT1/PD8MDZueiE2svRiroMLuVljXp
LTnYjDigMrgBKFOPTwsiwJDu6s5dQu23gEwIVc7rBsOq80zuSh2mJHwurbsFib1IXLoZiOysKSuR
XeE0mG2K9APMQaV+zoTuRKEurFTOcKHqcC9UtqDnNtfw6XlbShglKExzwjcEvIgpICMt649evgpZ
PrJ4PVYnhUXqyzyVd8R2/ZK6g84l64arTu7Uz54AOfBdOV1jHGVe0Ifit7Git3aTgYq4GsS83LI3
z2mIzQnSB/jK4wKqsMfnnVgYfrDBXAMsQWCpXABqPwWEz6Zn0jotLEu2MAQIAITLsUk6Vg+wbSZP
JuQCF19i9+XapQhuLdo0dqxz3YYIwTVAdPYy34ZmZ8ORUdHvgsy6o8d7fCoAhBy0WdmbHv+t0/No
hoB9h803me3KX+HL/tgcXBcDar6lUWI0Y+Zv+UPHWmxCDXSk8wOlIwE2ZaPRU8jc2vjk4bUO0p9g
ElXMiuXfSR6R0d9g0YxEn/ouinfxIHNiQRBmQB1KPGcRaq9ax1h1smkLgYtc2T5QWIlojGF2vb+Q
+XlYySwgjl5Pse38eiVZoCB6tH5+/TY6Euu/8nPDad98iCdYSLe97rtr+w63wUTrZGc8HyQ4gH91
NEtlpadH4clxftBYPb5AiO9W4Vi8vX9KqArkiDU89m8hw3TNu/h6Khef61r5LXqnyLgE3CIkS26T
gwzSRs4CctOksgLlO0tQ9dmyngDRMvzKMN6hgB7LZ1vkMkIdShyR6kU1GBHvJyVFOPtPN/9R8T0s
MaZtOWjkfSFK7EmHL3ecSsRMPyRBW6sCoLGPnWqyIxzxhjRkIQWEnoZ4MHT/iMcE//lpWzhYyqsD
gdW0n7qMA9Y/xBDdtMeGJ8XJ8WI3+bmhlxNPm0eJRUejuanchvyNQIqXMlwKuj8wGZqXOmWNuAZv
mcs66BPNB/m03apH3Zs2n8FHnkBG7/twaynQZAk9BnZv/sQr2em4n1qpYfhzcLKYltcAsuyvn+7o
3+FMduw8mpUQKV2wUgyU6rh3zylVuPtSODeO2UWSQ7VsrFORFWRxhghRiW8BoOg6wDvGbJcXfIBS
eRB2Vz2/4jP/LtHqWxAcihUCTGqt38AG+9pJ3FxE+v1zhekYb3laYxq8efQHeCsToMlOwE87j+5S
R5luCllv5ozNcXfT9i+FZt29/A1QL/W3YDn8DdkOTBhAICLuuqiTvAu3B1kVBzVZaQOTwBjtcmnB
3XxU6EWlwvj8crDbZGhapr6XA/dXIiO8NP4Yx2MIHelxST/msyraj839kSNqaAhrN5R9+fO0pdSv
4zzIK1GSkz3CI4Azf/sJy3mMyuxU1nNqwkhze0MoUjAlpv9rVOSywdH0A54bAhDf5hTintey8OKw
ugBgUFFZSM0CezAoroJqaWBQpToJIvc9uhdXJuRJie3ahUNDt6mBvyrc9Su0wchDqJ9e1g8ftpqk
NNOEtoJl8zlarpvF8SwMcX4MQGo71J7IkSfAFLXsbY9AvLrpyKMLrs1SjCXEvTR+EUC/DDiZvz7a
nnWnEIIUH5WNOFXCBNqrUDFAypbF9cZnekmDVq/BHCG5WMZBAW4L5KQS9o/TtXXcW2FCr2bcRjS/
Pe8gePQbnUfjv7riudF10XWSM77xckvjzBdI85RwfDlKFFQgmzUzgxiyGZBOz+UM/ib/OZ9P3KEy
gIRZuOvx7VwSzFqiYBwH+n4OyP1ng9h809roGAgU06Gq14K+We5bQNGtruCNdNqNhJKsGpHYoS+T
aneU63NsvpesZUH01Kiw54tUISqkPZfRVCUiOW6XN13jRg1uVfIoOICRBPwzaR3Ty5p7G4l8ibhc
OSqqwjXF2NTgWMlrVdwNjX0qNG4iinC2GjrXRl2sPcTZXVVdOCkjUGoOHkMvJaW15/u8mCq/rAb6
Ia4a754Hk9TzE4pIRx1ojxXX1PbkWmmw2340SA2o+3bzilYmwHiMpcR/tsZFBzv2aBqI0PeUHHCF
gNUq/Kbz9ZrdPLi35JABk1npn4/1YBFHzkSxb0R1mx9rtxO+RCSt1XDzlsipC1iyVi1aAg8w9u3B
9eJjEXaK2pY/H2aa+3Q9qWkC+iUjuqF9Enn7NAa+UcSWBFth1YgM+bsw+ZHEAWo9wRkyj3YILuFV
MFghu+CiXbjlDjh7t14y0VcIYsKcT6WrG3j/p3il0rX8FN+seEmcvQ4JiGkbzeVcigD5A6AApewh
Iq2uMoIINk3I7Ahs2LEBRf4aJhuChCTwNocSGIhCO6OcdPZQ/N/9ToVqT8dUwStGCR0rjpGbVt2Q
KkITs31wmXGXBeh02WF19VPyHQEAJNChm5TLsr8eKQzn+DR0ntQYI/07g/BdD44lH/K3TfLSnoqp
wH0sYbeM1KBbqWJYdye8J1gzr05ak1/5WM7RdSrGUs3ZQEGJpmKKLEauLsb7Md4vkgn9Qff3LlSF
XTAKNnbOK+3dKlv+3MkBBRo1XIS5lC7VuYDSl+CivG5LzxsM+C9GoGwxl1+GCD1hUSbK30VIVfsy
NrGKR6OlOqxF3k0nvLMHg6Vr/tI2gRE9zmN/JG+snExPNqCu0rrjR3vXAybjdGpWotj3+V/i8oEF
zxWOEO7sMmYMhT1zTEXzhQw7jlm7XsGotXmxuOrAEEnYHfhAHJMFOEkcYU0/hwbS5Q3TYIVm6yng
7JX77g/TohxpgtllD6JV47ay2XXF/wm1KTdFn3TAcSEIpwqHHqbI9JdeKSWC8kqgJk3+JG7EYxxo
mU5eYYvDGY9ZYf/Wms56YuC0EPe86NF2fRHq7QZcWb2Oy4hc+69sTXckoosVi689D1q+nMO5lla1
4hgqqKVCoQEvxQrVOOkP5FQvkiWlaWjscSkpJjoN0LmMJEDwlqT/aggcOyzUCpdVDhJl/atcR7T+
Psvw5AkiSbJTbadnYUDLtDL8BtQfJEMHgb0x/8qQRVkx6PBSdXgIhG+5TnCE4xjwXpK2vk87/BuC
S+oomq1l9xf9WqDMQvePdGilPS0XO3XPe/+7+3U0ZPJYg+biwgaek/ChTuZ/nRu5NAPuIrocHzKM
EoDJIeXY9pPSGqfRTHyWKlXo8QeyMgzNH77Ln5tjumbJUcBVRpZQgz/nXsLCSuMg7p4GG8ODvpVP
HUPUE3voPc5yLbIIdX7BQwO4CkINXZOxDXNDyxi5efSpU9vToy8pYVgw3vdmp91dF4kJjMRwL3Fy
ikkvlKUYwMxwk5G3uaa0gTwrldg69oM6oz/F9+71B8380d/8CbCv0YNf+IcuJBhBBCLn5lHmEr+d
EVwtCFor2HJ4n946kPmJlqPuRR40JC2eSBnwpKH+jq/KUlXPXoBMpcaoCG5AcfTUWdEgfO9Jz70l
4cX7uQ1LsZUzDp3vpyIEeF22nZ7aGAda6RF8l/L109oopTGtr+7HDgzXiTUZLgnWaNNnA76lx4TE
SjM/EiUjpLpcAJ8esy2rtuOde/EWg8iIPIlywzS6+73u4Cz2BjlnjRtKhjYqkcmZpYUFXLqsfS0u
t8Saqpza5AyW+kBBqftfA+WW9L7+N4inRlLdieG0dnhOncXa5+X6t34SJqxjc1L3vbvhvt9ef7yy
0Fy9dBW+6nENUpPizV9shShj4o1FN4dzxd5KUgcQr/CAvPEJ6Tb3Tw+6uzQM+ff/TQdw6AIBhGnf
xcuuOf2xNSqosJYgbiOlnWRcm45FQLFSQ0knkgCkBxwIpIph1os17O97e+fFsj/n+D4R/fGPzcSi
JANGZsMhXSNA170gpJNCTj00FGXlpg9pJ9aY5CyZrULjGZYOUjs7xWRQTGwJeM2+nRsNlsi6skcN
KwGetk95JTWAWfBrJ57Za1XVZizZSlpsCTzdkTdSzQ3RL6x8wDQvnvbyGLlJRlCa4w6oQZpLxdMf
nlCQj5+IKmMdDUPgq0YiFG1Iw5N/OwMK/Q+ukcBi1hW1BGhxSvZlWuxP/c4lbT3AfMfSdidUnvTu
8GgRUVjEV4pSCtqCfMLP+dGJMqcdMHFHHEs+tbjXD+vPs1LxoXoMnXB4dhbZXDmcnS4D6nou+sIM
SB3snHEhqPVgl1uMDTSj5QAg+jkjP3qiB3gcrT7UyPSdgBJ5cLLebXoFvhxAZmdIo/aKjAmv6WlM
VRyQ8JmXMbjTBBeN0bvznyXBp4qG0F/Rr61h5HUiIfhaMWtTG/pClghFicNHAaT7QTq5VHYzNq/a
48miSTjouTPLUh0QejJfNOStGRk9Qv0dI2QqOIhF/+5VEd2KCe53gmj1jY9jnvlcg0S0rOQ7k3e/
IOcNWLJKBTKACnih8ukkbel4+Dioe6yvclPdbzEhc3SQ8AohmUvjnfgOsGxFAO4KPvE59TVO2Ym1
Vc11ucJolaDJDvd3kTZ2QvL5JWcjr6/zrZRiNX91ITGYv8D6D0WXWwdcaEMroMJnoguLbKy/jsCT
nFSxm9xh3sKsFIbhPIkjTDhWEijfDqa26Kpc0THCd3v0MpIvEHuC7PhpFnv6jExg2TyhPLWyI7B8
fahtJ7DA57Ur5pqS3JkbsdfykseI6TjyuSi2ESAk2oymYQ/0tvktSWhDX4w2Panbm34ZIwqnN1MC
3qHCgMpPibZ/zWoRdYDE/Qus2ExFA5iFXb/s/axpQNLNUCa+hayGyZZ78S4nuZleTZJ4iU5AhaKo
a6ffapSUmW+pTJ+yyDlBjXfN/H3ru039reTZ3d/Zue4lhg1Nl+tRB09XvNWqi6ObaUn6h3PHeS37
Ub5ORZHMuqo5IhuhOFZ6cbTaR3gXNF30t0ssy9X3+pTFqvZEiNxSRZcjh+MtpnbeIYRx25goWfhW
5yeCTYNC7PY4pQ5RV4INIMbpW/lVPnb6uC+g+FY/ASvzVumOfI6/3+5AQmAdN7u7ngN/MihN+iz+
LpUfwVijiE+6anVyYiP7W5idGHmUMLj+rWmpoBUO5Ruy092fkB4UfVnJxpxNrxepXxGo9iaNfC2i
lz93QY3MGdRkLcTm959TjYtYSlFBjEfiVx/tm6FoUf4U9IGs2bcwg48bdp6rR4g4JQh8XH7LWV6j
7BDxuvxu0MDTYXVTaqtVBS39ceDb44hBPLcLiecTU4O8OvmhC5TaXuHbNZ0b8a6L5ExS+TCP86RG
/u6WOcs2dIXe7ZX5a9SrbGUIGQNQlTxurGsJFjrZTT/aGQCV/Uu8QczmACiT75aVNs5Euf0D2+qp
hPs8GS2pAyUAcYtfXhD2DvsZ1/MXN4ZC/GoohG3rKKdL/Vn4yikpA+wAUoEpA7tl7zGnFh3i6QBN
ZQ7P56pvAFmDdpu9/0R7v0OxSNWzSAVRdxjSHV1dW/d4k031VWSCsdpJgFIbcWIUYVVijNraEEpW
t4VFb0SPXn6150KY7X7siQ0q0sTNT0Ra60D4WDbl1830XHhGXy8mYSUwsSPpxAwQz9ej2KlAjw/J
uGoas9EQdZJZU4feh4qyx/smHsDrLksDsWUChZDLmaJO1GTXZ6mfOXY8C7kAsVMuK1DmNt0wBwY9
StK2i4l6vAqi7YBujBwDDL80okSW67EEZFAS8nk+60Mm59Rb+fXrYLNXJUHyJ1HrHOucTFMYRdOX
jChZlr9zHjmedgkAVysCn+dWuIxlFnWJgzNyQva7T9afhdsb91q4JG/eu79TdTEkucqNN2DjkMki
DzLMEQVIUcpoplH3BtpaMIyECq8UUBg88UdQWjMs5wegME33J25tzRAWbWbZ9ExawEkjIa7PCnEd
e5J9WMnN1eqeSaqYUvKzkvIv7Sx1MozjjTQWlZMHD+/SULjPBU+h1agskITEWnUh+eQrlXsF1dut
jw9gcaWBHdjna/jjzRrAYwyvvhn/vNE+7OdUqd7Ywps7OFMTgFiEnOrO7Cdrgvmbzvl5Mp+digYT
8BgqVpCyzXwgm9tlfX4b8tfJY4n3DFsarh0JqLBvCZmSUkJNHvgFWzl1tSVj/pbnjUejL+7IY846
pjiVi5EmPU5wij+uMaKpqYkIRmeTmdV8IQ2rriOSUp6pD8IPqgA5m5f/MPftVP48G4J3CowqZJAI
VhrFOUP6FA/1WlTxWb5b6TgxGh8zsikFFdaoDDsRAEhnKqln9xanxkgBm9cHAQDNhTzgXTeMb+by
BnxBUCtxFmAY84lg7arPeuBHxTyLUx+cmDFu3cRNT1PFFwGgz1KiDVZ9iLMIBIfJCAprAgr9BtZ4
SD6n/uDChZ96tSVWtLpVFUb4URx1dpoTKXeKtvw4mS1RhRjFWQ2F6Ir7HBUcyq+R/ZcdQtUwzfqg
8ff0MSrKf28tnGezVsiFlLXVhuj2KzIqd9GE5XFNDgIVREA1FPNWZpw+zbHhQBRfns3UfB81VE1K
3s3Bt18fVNd9LYtIFyJH6UlZnXozq1SNGog0/sWGi8ilDTxQLN+cHn1zat9B+bZ3qwOga0Z0qdp4
AQ489fIw739MBaw04V4Hzh15qKBMbvtDCSJ2vhmlVNip1gnbYRaE5omXk9w7JfCf2tgM4zDnHPjE
H/tNxhx7HMkxCLzpT5wYLp4XePP/Uo4iuYDviodLZkOiL0uJW806hjBEzXopQQRKK4Z5WuSgj6qD
fn8Zo2Lh2wTEIDZ7AnTRde4xc93R+bbvIOPuOD68qYA53tCH7OWoj3zz4cbHsUmUfjpPkSBw/ubz
B0IwvasgV4y9rQXLktlXUSrworPU0NnE9BWBmXAI41ZjTtwlSuB1pN8yJKw9kzQniPN+9aO0MCy0
3abBZ0zyeoUD7LwudifJOYbK/9KXuRQQOvR1g1qVK+bNMm7qVhmX6cmd3QokzCdaKz+8xA5d9sTm
eY0KyqDMYTm5UHiX/fqbxxkMC7ZMgf3YXmZLT7xJdbWdRnBDVsTZwUz/Bxva2E4sJ+u9mcc+D1ob
5nT7y6LNJ+LItqmCIb3tdBq/qNZtM6JMVZKZMgyS1uTfDMX6ks5HeHUU1wkNhmAK8tmdwgMyrB91
lgoG6QiYP4y6rNR7iBjEJzFFvxlZqZxmFHHBMaKXnN1JDirU5rpjDI3FEIWOTbBamEAUXs6GMpHc
Vu+TSB1nmvqnNPeIt8cMP0G0R2HX0FLlfbtexbx0Tlv+rNDOWMh3BIvdLwtF7PakqBoMrBrAWXE5
GtTxNkUaTAIv6kG14YD7nej2qXyOiNK4sSax3sXZO32RvC1PuDmB5wEzlkMe6mq17M77gvphjm0B
4C7SeQknGktviNPA9SszkthKc/wIGi1JSbLtQOWBGi0XOul0nQiGHTJvGkeCeKZHEousu4CkDXkQ
zs68MIH7MXwnLbT7nvYC6BL1YJSb6rdMrgvoSbnzu4rtb1MdXUE0VUQGfd7JN4ynnjY+kkoPKN//
64wI/Glq2TGDrIwWj+6Mt5h1QxKZiI2HaqNqpSpfg4BHqNLiFBVG82T60NaDHNFspWtNwnRXD6qV
t2n7wq+hLAhu3yX2794hF0ak0eKg05JLDPF0O7fa2qdncveLo2yXQ4t+Q69G2hUjkLG3uX5q1mFU
9cXpgOZYG9qiFkhpWbTBVf4FtXZvQRZaUVyZZbjLsen5gHEbY7L72iQawMUB4qDqtEBtaO85NA3G
MR3saRGuYbZ0gDhEWtOSa6+TY9gr18ro1E66E9cAn8HQOXjDlnmY13wp9f2dILEb8+Ja8I4xgsd+
nBLlwws/2WokKDcHlUNrUYOTJTSVparg716iCqQIrJPjRKfqFpyuWXzkWgCDYSigylHkYPRN5E9v
N+b+LsGb2uOy0Up60WZhuj6FYu1pTQHTdX958h8yy/eGS2xl+8ptOsoPPHqp81qTFrBCwrLh4pzl
hqs6dsl5X/ut9Ag1TxMZUT45pxz4//pKs7in2DqGJz6yi9RWXBjqBsIwpkqJeau3dcspdIJEVeW9
jGQOMxW1pbVQ+BL8ILuRVCwg/K9+dgCPptNOuCE2IhdfGTnFPTVYMnkxPoRzeehjANJGXx86468J
iBCCk/SuhnIA7KvMcVac7xGUnTQyJYLJvxd3bH+ZFDyiGjSacrdqd0GlNjakZ1A3GgiAVrGhEqCk
NK0fN5VS0ZT9+ohmwvO2vZvwLLBwMQE1WXa6dCbncxVSoPnxdWqr6Diimzv3ZOMWFkvVSPskLvV4
hXmESsX/xvO+hCJp17xz8cOixNxfs+41+LmjlhxZVpakJoeGF7O8k5jrUwYd6gchGp1w05uz44/0
Nh9AYK1PtYjtgQ5F9bEf9plFyNn6nMEO6dfZj+8dsB+8/L/+x6/ZuLALdOEK9Ov5SO2lJw1fytI5
fOa05PcuzP6XuHsWh8kD0DLa+NJaNS2Ycq4jyadO4oJthW26VeA26J0PzksxURawY/MEeaY2AUiY
b8z2+2Jhv/mOSOszx4eAHSDasmuKHpBwtlSk0we2PyfcElWgcQyO++UE8wvH+/Y81dlumNUbjBSo
VoUB5F8bwU7mNYYw7ekn6qUnnQq6Qvb2RuSWZUe4m6JvNIKhhpz/L2+bErmM9Mp4+gxAye0KXcrl
SsPpm7U6CIWVb3wVfMKS8cHfvXRF7mczqGfFramb593Yx3N2UWlZYDxYyfAwofZAjryTflegKfxU
c292IB6IhNl6SH5zV8ov5SUOXr+HSE8HDuTPLiYQhSygW7fQxWcVE1qdvy5oFdcK6YpEvbrPzdha
BJ4vdQCTyFvRH50uwYaol0RiZktpSGzqxb1AuHo0pa82Seyu2xrpNyXp4sWCIPzx4PZ9Uc+BW/gk
NIVZn0Zynd6ebDycoHsuYfG9JKrGbesikuuIbMtkfQRctkO2swY2CUPnIjTueQA3WZRaKAoUKGVO
jwckzaJw25oOLE9fvZhxeo5nZmapEKnrfHSjo9dAFIRLpy+8O78VByFuLRxNBEH2QFiVUBr2/+dY
GbcFVJq2EBgs9Yb7lAbiwAwS9vreRV4gDe22HZ404UjO3fdRwf0AAzqwOdFZd2aurMpMSikM2xBG
dXO8QbyGnQtBYia7Y4CikTIBvBuuvzdEyZr4HJhi1dVAIyLhsBNfSxguqWB3yrb5B49b/gC/ubzM
1742lsCYiiJxWRynXM5/zTtLaOyLegjluGiraCbXZtIqoMEtTAJH2F1KL4++SJvDWZlEjhvknZdm
2QZazCqGFZ0W0wVdkZ8MCI9ff0OzaWysZYvY5pk6r9SLSDoG+5mZZ21OqdFsTDYkTIFkOOXl2OGE
8gUcIDhbMn1FZ6kXdfTddGpDH2qU+yTccLINk9Zu5Q5xFz1hUv7zIkHU75KIboRj3WLgKIDQQf/k
e8Df7VqR/Y1TLBG4uTdVMQySBPO9N1JwYnBsEYQOjY19tn4tCjUQMvaTLZktObUXXUhw+aRiZQ0i
xEzntXJbFA7wWErqk7zmxyWuTiM5KrChweV7pvkudF9U1jbfb8SVyHPRyJO/REuBbkVouunbglAI
teDpCFD/JeFB3UQ4sr5+Rxs6ZRTV8EPGOd7g6zx4z/N2LttyixOi9lloezD0M3LX25fLKJBrDefl
BvT6ChNt3NY6HjKQ76XSPJoPgZYZNUIGMNhZ1RjkEmEiFtSqZR+NbHHjeowXtFiO9K2bu0jKephq
jxHicau4FZveupS677Edv5SeIyiVX2CQurWKI0nNPFJ7k+btZpsEbP8Iq81Ip978PZNPdF9A81zH
W2/JfUlV2j58zEawJqB6qBaO4buq1OB8ZDYqWtxx+5OKhe/z5zRpXlH8SQaZ63u/5gerBQL21Zyb
fouskG+/0MnP6BsNlL9Pdb0prdhXGf3Z+pp4W87KQ9F0eP5S5nGQwYP6K3ksfQELXj58FbPlI0xQ
oMNSroZiZBRnb6Tzvx42ES0SIHKn0T3eIaWXeYv9GLCCgjcty8CcELve2jQg5XmxpTkmEXtpibV/
be0Nq/VEdGbAcRol7Fhr+jr4V/zyY4A6seSHa7UzyzON1YggP3S4GUwqBEXE/P2SuMnS1PFS9OCG
YLLD/di7GQnJSZzdrwbyCnQNNb0yg5t60G4PK3g1tW77CdRVa0sGB0CS5MhPzQP3Fn9Ypq45Qhkv
k7It/WnU9cot8aCegNE40Mfxfj01XePGAZAYBpUiLdcKgGzo29yf4WQAM6AVm041QVxqvNAKwYO5
YkDl+teFWIix8SAV6YQ8KvFu33fSPeoUI73RfKt0BASPGkrWGvzDrwqhgoQdK7TvjrXURYLs+mjo
fNRrCEsu+cV9NLWOFoPnDzloRwlzXn+mEXfmeigkyCKgdjviIdZeyieJlYRhY9tHPplYiaXmibvd
/BkWN6rICEw9A36/Ty3QgEq5YddkHpkxPyXoQw6eXcO0pKmVhByPTRDHDWRp2gyIZGfWObPG/nWW
/RL8Bz0jiQaSzm95SyU/UGegGUfhuFpP6hFGD+hkx7pMgEs6qak1SQt7bbEX0UHBdckLAzCiprIj
/nwlYTxTSXeZLQxehMcqrG8yIDdyHZ/FrqXWr343hFd96NBA/NyK5XxtIo3Fc6E7aqv0rATvOb5b
dWpIwyZik4yOSa881NpOROOkah3VrNzlOkf8iMHAAglbSthxgrmaazh4rJc+V+Z1u5hCSaixV3i5
hASreq72Uub7lH/Nt6XihOTDuVauy7fd8snj2E7/Flwy2JmtUvx81dLPSA7MutBpy77xoW/gLdQE
1HaA/HTianqik6RBAJpjDFtXgvRC1tOU1vifo7nlQrzGhMj/24DHD253JrTSoqkl1H1o5NgPGWaL
BQn+zTNfghoujZZT+5pZKVU4FyAGTMGQJevRHFe40X0sjZujCwtNwm0aLqA7CksC/M425AdqHtik
r1j8TK9+aOBmtPeqvVwpcamcL+fkwrlCn5Xyf5wfmk1s3BjvDPl/WBuzibimbTmDrs276l2gtuwM
W5yevMIn8NkPUbjDLUwr0lf89kqvLlIgdTTKTplU3BtN3VRrTZx0GT0FTwHDVukq7LV4RfcPdPF9
8TyfnrF/ht9DvAKQPWKOROgxoXgN7ZV7FqaIEKtAvUuwB02lUNznTjuqHuWQMW85VMtdrO2JBeIQ
r8p5iDmr3saxqEpXGfT9/dBS1k243cMh8pjOI/EXyBuBY+MxYLX/i379FUXNnhkZju+Yl67U8QKx
wFUCl3isoXewOmm3/1yo+EF3/D1FRczsy5GjSHB8GpAoSWAcOfNg9Mn9wh8EwoenTutAJ3uTwhrj
kADSp9XhPfiW6T4DLTjLCjSwmXC2WN73ru6SbdHqJKA/7kXq5j3C71/1GGQV5BTi/ExKXL+GFWfA
yaZIvzWbF27ha6CGwiHPTI6s5mtkTLRNoiSOCtbvPnfjOfO4HbFbVphk1O5P1dfCWXw+6gLABJT6
DWRUNQnGUHfy+IINq+N0oTHxXTTAvGpjPp602qSzcdirbITfE0TNYmKpG4cM/Nj+yuVcHIvXfK/B
m+oVW2WJo0HEvlPDqFzSE9FLexs9rr2ZqhacSDkGWRm8fBIVJAeQJ0F6XRkhf9AfxlnTOkGWbMvr
6nrpjVGMOf9l2gPT3f2I2MHtZb9IJWwrqIoW/ANZGj85A0pI0DPtgYTHPLmChaV/lWKZN1Wwlcem
8CdDuq0zLhFX4sT4efazUItjjNWjlYbpTANnfwebZHJh7CgyQbBwXZlR+A+RYEmXNvGjLGPer5xG
rIrEOxNl1rgskXHtGR8thBzOQCtR3cRzehD909k5THhHpB6+XxSd3PiJNA1RntyFNsR/XDV1WdJ1
eLjnDLMDafmFoBpICBhJNmwWdYtOJRJFJpxKGQnIxEKY+kHGUZ9HNo4/3XMjsmqJchmTJm7zLsT6
LrRnLynAzEQi7S7ZlhdsJrABSvqxUsIeRiyrwHTl4F0OpghbRmEQj6InXDe7fpX/2qq2sPENfY4H
9G8lJpOAf2sYz5PVHh2VZBdh1yJffDGit4IMhvHq9qD/gEYnERSt30casHq7XFptSIwFHN+An5Fm
KBTlmp8K9KMTVK8ok6iQxL22d6niJwMsS6Vviuxx6v4To4L56PDmtns2jBuHjsICz7GBBDV32bbd
0fJT6wWLC3+X0ci5lQFjBlPBdzX8O379GIhrkIrrIuU5MUJsIMy/rXfQuWF6fcgu+bKqN2ZmQos6
jFYK3wfi2PCz/9F/f4A29uo2ZrI/LdSBTKJs3aOP41FZzTMmlGF8G0rekuwpH8u1337kG4Nkff/t
1IX6LsZRwutwocQ7FAza0tBlw692l5AJ9tXSNA6ZpP0xP3xLSXW0FdPwvuzXA/W0qeRwCGkLCr/z
BiM+j+gBGNzLgeFGXdfatbZej5KikVWEKC0HeNbTmYDeO21NFvmfK97SXSQ3vxfxlom9RWDW0bG1
oeQVJ+t41iv1yZ8moRCRMgfvWYdylOVpoA8xGsNbnxBkBYnTvjJdQor8KMlBR5FrnKtOK6artFuQ
oxmqrYVQwQGoqJL3rC6mTO+7U/od9+LjkWMIzB4amLWhcg1f9kGwntlZU0nHXGufSaCbHAD7ykPy
hi6prLGnaiEZ3bVyz5o2yH5ofKt2H7vKqZJ7x/v9UZt+HTrJZCCnzLPUeYb9V7cod46PHvMXsHld
168j68ELIWr9b4MRGxQh3nEvpRpfTbqD4j4Ft17BKnlssNWokmRtNffYZ2XhR9bqxu9YOQJ19VUE
7McBx3b/3kPvF17evGr8TOV3O1lHNtohT/YciLpLP2eZSsEsdb14jPgMvhaIyMvZFLGSwkyGbPwG
IGYmTeQqVGuY2+y8kxhX+9OCmQ41BhNFylWsL2xB3hdFB2lvsD54+M21Yip2LOWw8AfENqN5oIYL
GkMLiYFauhvpedrxg+AO1/8JtjCg9+E+cdwufQ55MLB5vuOCUhtUcT343He3QV0a5i5C1rYtPZ/b
cjpdYZj66jmIgSOcuMi3fIjmEqRUZVUCAQp3Vx7xZIeiUBHf5qYXiC5iAveQ8Cv58yVF4ku3+rp5
B4r3ImxRaDfIkf0gTaCP8WED6nNqFvyjPfEIMUqvnNVD+PxetFzD8UtbCzRPsMpitPgZOaf7pQSx
ub7vyyUD7XvG/QH4F/p30mD0b8sQD2TvDTt3ShWCFTGHV7wKaVelhZLT4v6S3jDxbpYHOPK+L9sK
exhSAnWT15FD5QfDNhJtGAVMBXoVVaM2eDTvbTfofdln0nIEfEt75KrrX49auMKpf02cL0RINClj
80Ip8EDMEgr4/lg/hKR8yKAl58hDoNerEtb4hSk9EUUoQS64It364N0bf7DgoBGbpMGJG7hY9UgG
IPHMCv3B9WM5AXYNeCBEGJSIa005UiFEbUFo3XEt8ZuuU4BXwbr7LWViS6/Q4yYU7fifCoHCY6E6
JRwGOa+TGSDGaIYnba9L+deLwFqigorhwI0llAbTsJF3I8FhED2Q4w+/eGsvCqlr1XDMNBv4blpi
FArsQzQ1l21276bqjKieMpUaMkfZftN1tl/oEiZ0HdV5J61Sq9nCg5mwjNiH1/902nQp1E5qA1wP
abtZpJ6yoQYpUSJS2NKXNvCKaQQjdUmgIGh6CVxcWRvKhPTuzl3iWqC8/Bx2LwTiM/87dd7ZLTj+
8wdqBNRKlcBbeWCQTfLTbYcXnkeVZZvJnevT+gAInQdISuU6gfyvftEiELmrKBPve3xp3KBGGsG5
S+8KFwr0t3+yo4w8l1I2SOBlaYZ5KSZTrVmUxBRiKq5kj6WbSvvcjy5RF7fbQPyzEflXdf8a81rT
hCdL4ci5pePua3qHt1FQr1Aq3iiQ9GqV1O390CxIpYePm9b3XJky5HDiYkEPiJaqhbfJi16VAseJ
wZ5dbWB5GctVzcTNS7DRV7ZWW2yqZJ5/qDzSuqbstlMWuVfaiBvPPNI4jbSzQekb6aRP2zEzExvk
6Tv/ec/5f9XUpyDnuscy4FxKu3Zsk87FBJMt4+F1x5mQcJiZzyFj3uC5E3uz5NLfLpNNx600dvmV
wY1GIOFghCoPJSf1STinECiRnKLFoQBZaYTcSMjIQqcHv5ny/vknPCbHzEovJPkKkNav7SIbuJ9d
1yPkNYKpMVVNnMudE9y6X3LvgLH1zinoLx0t2hPgptH2eKVMYTvKFsNvbKYt9v+VEW28+HuCvcRy
lUxHuG6daRMEQUAOq+x41ZnyswxM2EiFT8wFMzDVK3DVi0mO9uQIJnEG242sGACDpVRHrP1rpV3B
jdkg5cxytg/xFBpV9lKzUffHMUIc+ICyVGXJCjwyNocQLNkZwRthqGEvTqPu73+szSjffp3D754A
qN36z8XW36BTDO/P3ft5DtalqeCU4j71KpyalusiTak8bGVOvNd0UmZRPssoOVyClj9uhbiV781f
zGMlppB/WSj7SZ8+41MvzM/McB1R3cqVs7GlY2XVZ4CF++dAHsxrjqtM9D460GC22NIAwMGat/GM
X2+JSnvXBihVn8j9vDgYruzY7kREgcN5ZyEY/OyK3UTuQoIWAHVYeq2dL5jVrADhqppcmN/YfWdh
ApTYpCsfvWutyCxKs2WH30iv8iZbTgBMuQHWu2HRzcDY96riQyU9Nx15m4/VT0w952WQOPAz1LsE
MFIvJkPaer1h3Y1kLpGSiufPe7AkeUaM4b7sr/fAE0S7Ass9LOknTFBBD+ypyUKmQDjgQUUu8FTM
hVQHrQYPtlWp5ouaMLVlUVSW7KZZ/eFZ0hE2+OBDeRBqOJzGupfxdi2UxTgq7Zm3e+/FiBPQAMXn
OlnCQvVHb9wZmVhQD0Ju/4BNtBftXEfr8YTNgVL3lV/7yfLq38jHJ80eR9j6GxHZjGyDXJXadf2H
YaR4vi8IrM7WBqaRDuzSXUQk1XW8aR2FopxE5fM0CJ9rcWvscJElWZofDUZC8qMPfxzFK+umtXky
qSJZtcmCI6Y8Gf8Bl922mFz2xlhL03T4ZFnC3hsMsc+qwTA10ijbjo+Xjcm43RBEb+7DW769hQkY
lJZa8OyEKTkxvavVG61a0C3xCa3nlHVtMma2RpEv0cYBa70/vEFTfUtrSNkfM6ztYCME3g9z3eAO
HHejs6Q0JaIOZ17RGjUi24DfBDj84O8tKEVgq49p6kWZYljtFD5PkFW/QbAxwem/140qLe6adktu
NTyPb8GxK7j3QSzrhKtjxBwXRfJQdo9yd8/tVnnRBueJOBAvH3JBrNLLLziYVpy0mY0r3t54KsLC
4b+WxJzrBBqrt5KIbwsrt75Qbf2gRLxiXq/DSKQWnZSwa4h/SQvL2tIJ4NXzLVSXnGN5Vq1VTao7
FNc+yQhavEbr+rUoU9bMeq6myZxNl260fGAxyOcHXNubnHB6oa7PalgyohjPEBQ8ZmnFLzoAhxXB
k+lplJsyEPqI0esvN1SHF1diqu2qyqlSS+WLTj3tdvR9MTyi7PjoI8eH3vO76x3pSz4i/d/wvnHv
eQ+0nZx2mFFgrTN/6tPApmNwNSrnM+xmxKEAdUAe0cJSWaY7f4XtcrOEBU5uhrMlCSTIFLgQNjQL
iqxOTkwR94QKqTjSzbCa1WmTzCdaPfHTogIOHsMH4yNV+yIIgq5051FOmYR3Ta2RQKmKJZ4fgerB
a3WvxVnUH4OtHrI6pT5xcpJQU8pBMIglmZ8XS36kn7OpotxHjXTbpTg5tAdiLSOIj2pMXd+xLxlQ
ZAogjGWt19mjVWgQpat6kf7opZ7nwimn0K+Ya7qtt+yTZMXxEMzOPdzSzymH7La7ZtKKG7auCJo8
Q7F2DVGxu9bQg146kIeGGwJ1iSf7gHVpB9kwYu3vtA29PGvekALoTHm9+KV/mlmoUkw8n5WkKiPf
iDhqAwwJgsaxKtiu/qa1mGV2yfowLS7CptKFpuerGQmZDgygPokz2dm6ruSiTfTmWvrXgOcMQ/qr
qeoOTaIhT2MhsrwthKJ/JHJw2jcDFPsNC/mOGm7v9tk1CivozvIgn+5o4//1+xxZlrm5dr5NO7aG
cDH7m57QoBHnZSDQ6N3YQG1zVeqLv6Mgrans5ZmiBuBmHHXdheqtbD5twIObSOGSKDA3dGZSW4md
hfMzgVrN1ff4SQqnBWzWBicJDjuRRvT7W1zhx4T7uNwG3Yvg5mqqSOvBPSTf0S95A07o6rqVAZVS
MVkx6dSQvx1IuNlY2U8X0FuwpLyvRxq+dLXem1/laQMOAvGvcJ23SwZEysf1fF6Asm0l29AlGT2X
0RJKGHuaeuC7wbh3n5YckFm6ytJlFMPUkctbBTiaboI51lTvfmBthVbY6lYPhLS8fpztLtzkj4AJ
FVC94+TvxmlCbORdkEb82V2PmqbNEzuyarU+QfGzIcO7HbkvX2AqTGcrB2070kNZYxIV43PIsDre
ugKnayXJB/PEEJ/as3hTwZKlkac0Z/HdQqhViL3Gh5fzQQpAYEHb2eOPpVNIc0TIGIySzaommhMt
QqQf/kS28uOGh2b2eVRLtUykZtT/5rUutc+NQJZYRB6kwATd0ajP4zoQKMYVVXfVJWIwsIi2pHWa
8o2kZNPMzGGUj/KCkMrtTF/USTQgsLBXEtDMGrfWQMW+D2wl6jqfVpWDdy0syiSyNXcEyKV0XLf2
PuNEQvEiVlNFEOUP5yxAJ1j0FGKe7cdU5dCjURdNKQp4oF7Pq0JgLpP7O3CUHUYBiCMLkteDKRQ5
UOzsKbhWvZN3v9qD2BKBflqd9N/kJRiZqP8Z9X3GP9cOFfH/OTpMzIFg5HhvDlZLvAFY+UEgoKtR
cXxk72CA3nFQTfwmPlYvrdvwEsJc1WI6AGPqrwTWS+KYoji54Ji45/BwNFIQlXSMhWXHRKRM9ZUz
BtkdbAL8YJ54teZhsD1lMEzMMr0yimj03Ekh5doFISp5bQ+6XnPGV6tHVUZOuM0W8HdpWISZMqjX
CzVTsJHFhF4IPqk+2Pr/K5wPM+zxWZJ6IU6w/UP7pIF3rp8OyZO/jmrF1iNK4BQ+KA/Hbj7bb7AU
WATTWv5ZzL0gvyaCPU3C5j68xUNIljn9OgeWzu9gCBc7ca08QZf16xMf7nSuQ3232SzMAX75xI4g
zjj+4cOcl12w4RZy/pL7FyvNh3yD9vR55XUwAm/UnG+oWmLRJYWwygb/Oq00rgdEAVQzsNw/BP+e
bLSyWU0eYvvjsEPajvcK2eOo7G6D3yn6NrfZ5ROEDQuEQRBDwHaNS/N0zQVKb8IZ2BSw0umtPQHm
BKyyQHykdVaU0lw8suwlm2+9YjaIozByixNKgh5gAAHgr7VFqvZq6FJL7aAhoLXDcd9g2cUiJEM0
r0xj0pixFslxLwtO4pWH3Hfns3fQdfCIMPnvjcveHdT4zdSaRjM+ITYNuwomWXkEM7mOWGhLR2Iv
3bWqpZBd4zRVkgh+iJ1p9IwO8jpHbOqTHKj+CUm6lCxWmJFjCAuYdU0fho2idlIE7ntasyzy6YaN
kdmwN+HVIQxmwIWggVYY7KXf8OrpNYeeIr/iAgkKJkXBrmk4N5QU4/bu8mS8OEuvVf1REDEPnDMB
BvRXmkxhdUaPLyb0HXfyW6+O5AMGwH3Od/+o3Vydwn1K+Af9aIBHo5uo3MJhyF1OLQSQCQjdJFuT
Kr8GJPweHilENhDdYCI/tMPzLct91DaGHlgyqWoOI3g0t48oNgBNKad002wc4+stKadM3ih6KjOS
xXXgtD2pGeUEMEA2XatNgZuBTsO7UfHBOCvclx8tfmrSiYFAXncXDLirjEPX1S/8HyZSUZfM+bNd
N2Ggempko9m5OZz/FiV69wkV90A9h628xIet0d+aF1w/9x7N4taPh8eCy2WUnTJsSJaWBVLSh1J0
zP52wAJCmeLthDeSCqCfYuny7O/jkHVxz2gRQPuDUZlmaJLQvHlx4gDjg1t0MtiHIQvhfdM4e+zb
MOdai56IDMiaaut8uZ5qRaGqsD/Y2CQhDUScfDmeQL00nhoKUHd4hKTPkpFk6rCW1PJGvItmjvwO
ymEwthiFYF6MjXfozHNFHs3Fsz8Tk2Tt+ZcQE8XP6WgjscarlWx5cZCa1PJ7ti3NSkutKeR0f7Vo
BcRFbCS4UIWmL3Kb8xGY/qmcpLUPQVI4/vMTiCmqP0sA0UDByfFotWS0Y35pZrEvMgwhG8ZmOtrs
0Np3Tj3eS3g+drx59tIcCRP252ZMlYkwdqqNoe9wDYmwj3ELuW7XL2oFGN3pgstcvP2Py0gBwxOL
zlqFocGcaK4OZtYRgbnD9PM9PQUjBe5iTuvq6o+j+NY88PEcQuOMY8o1LzhX6O6TPDirI3oP0oZV
/GBOjipuPcH6PRADAHWBNgZGLa8PkkXOWX6olvyfaXiM9SW+IUM6dmJ49tFCHt5+wZko+GANN6V6
qUWOSbjha8Fl6W5CpEYHBjNc28hO/YMeN+d29qR6OfhMoTQsThSHj1oTo4TPa4Exajo3v1Wdk8Cu
fd/xSwDUP/weq+yM9t0PjZART4R4ko4RUrUcaqGWpLYybaCGZ0SvhORJh8j/JnpBvqhdQEqsWUrm
oPgkDNDLdsNRCc8NFv/UKrqoffNoCO/wX1OHcyUPn2ktmUTijvDQl0/wJNbG5nzJ9AKkaGCBZuEK
AqA5A2crvRrd+KLvsMYVL44VjntsDDBVYiY7f869c3kXIv0y/wRi0SI+QRtzLbWicUfhYS/933vc
Yftai4tSrpWfWiqJes1M1/Tc/P/Nhz/VewD6GHonUAxaGDtDd902HkE5oalsjQc4fM7XBIFcaMPW
2hqhi3qNLjx2FpPRs79Oa8W35zsSSxHp0eyxLf6lUw+2eZdFQloD+Lx4DcBaol5s9hQ6MTZJtzUI
uNCFhxic5rEML8JDdJJc6w2YVHijft+7pDPL1POjMr+XKT0FgrEsqlYY/9F9wW9Cba0IKtXpbTGt
ulpYSZqBEzeuV1uXKPLs9J9qb9VftsKmk4e04FA5vFHJkO5GeUI4lUPVgUfP7poUnn2he4w5etmI
DbkHOjQhXozSxWy1pzhL1YrgZ+R2rh+qANqrTQ4WpXHCPVSeOvPIy3SekVAnEUHopJIY63aOqyn+
KmX859dgRfobCVncf9M460jnbehAcsz0/qMJVjoCbyPZQcZfZZDv8ux3tXcgUyl3t5rU/F7gzAgs
mhTyNr/1xE5O6evcuiq2dbwRJhgEpu6mFdBHUr+a3lVmNWcVP/b3+ymA9dwmLrLHsnzGjfwRccB0
jLoAp9XCJi45Z7Cil0mu9Hx5JZJcq3tft5EA7iYAGJBPO6oJJr/WaoB1OU80E+8jo3D1dxVi1b4X
JsogwjX+5gNsMLXCeT/1b8D/Lp6ymYq5Ak1gXYX2VDQ1xmD2gsIy1lepkjTgruhfHVGroWDIXw44
Mbqn1PUJei6nAt/Y2afc0Qn3DCkbXEpC2wIEcNm1Ew3FCSTLkULi9vz4QfRkAb9FAanGrCcGcLfS
BM3nBY5FRWUdFlOqj5sMuhL39OkgisbBj3rOZs4w3/mo96aiEo2yI9uOtiR/k29uEP+7y0se8PKb
1U9nb6ys8u61LLU5lWi0rdeV9Sgwk6+n/b8ydubYT2yIK6xCliEYVvUFArKx29VeK9NHpT9Nf8Q0
DPa7hhIowop+6tmUpDZdY0KvLEqmPPfbzYk0l7rzxcgDbXkkzwYrOesaqILdr9bkXkDwAF9hsOoV
HGQN7+fdKjxva3155W5djXtDIMtnRc9dqfG1r8hB7TtRCb2Z+X4UDgwLuKA907St7OKGoP+M5hAi
Fl2IKWv8vheX+7rs4ZtvgdwfWPktF5L2busaJmZ6ohnm74SY5A8ceqSehAyIJVR/fsrTR7qbBTDc
HL5RqnBON5arEgOyXiP4FiPLsoOnWIvqB1y3B2ad2t9ptF2KK//xyiiXW7h4Kqt4Y6MvQIvIyIDD
utSOX0PcihvnKSzPWKI7TniVlmxVsj1yjRDnq70sp1gaG5Jm1rdf4/E4wx+2pYVNPhEJ+pYxCgc4
w5epsa9ni8OMmBbdHHcKMpmzcgbrwWtgVBMpo1+6EqUXWMkr4k3ZglDeacBXmLe7AC1mbCi+i7td
GAf6lspUdzW33sD3xoOkfoWML75sH7gW/wRZdTI8cK8uXr78DXEeDIkQROgE/TaY4jZI1DSe/akF
qr/rjzm57m6gQjVAWoa78qB/DXKmZRO4cJqh9osiAnc3C0OFKfIm6jTDVIUWTijEOMUTMqQhVoyL
WMBwNYuYZQ9FVgWkHK6UtU68LD1vUwbQ4IDm9QwrHC5O8DD17nJjqJl5AnQWsYJZFEzf0w+YyT9C
1Coq0uoDLUUecNJ58q4ispNaCwNeNbnF0HmIDwJkivDpC0aqazYArKvhq93HhxtdvYCbjtgs++kR
Bb1I9g+NeFkFv1Z1lgQ4MFITDEmP0oXGMh10kmdr2JMrFX7uHLa4/dGFFV/WTgQJqEl8C3epG8ot
pQuHeu6AJX8GFu1k7HggnerTDrH+Ej2oiMkkjtFxk636rTBLOi+bMayq4mtAMz2Q29N3/BwgCTEk
umzI8IMos/AjaIEqdkcSctgaZHSsxwx40hZAusAyqt3r2tJ62BZbw1INodPsVlprJCgeijA4MpA9
uXPjr8GC25ZUAewlxx8CJgkpy1KKQjfLpVGdIcFCtG9YuQ6d3aQ//EnfEdq2RQn78HVWtLiFbBmy
TQJzT1JSMLrLLj6oI5/bAou/+5DnKWEcjhzJ9x1ogabf1fh/aD3LWu2P1BEYDTYVJJ0RREAZ3HMe
gh6HS8bLXplPcSlc5X5LCu1LbXTOmAV6J72TL/rzxHemAuA+RMV8fKzsn6hiN+N0XeQko+SKKDzR
YDG2NUNT7Tk7Gp+VOLnqky4G58KpqKtJDArsQZbFO7L36HJtfsQe1AkVx4WaxYVot47fTBEGOqO/
fuJTUhW4pBcBvQL1k7e2ooiaA7xqLvYKql3prqpW9TERMDCX7U8YJLoZ/plHcmWyWyLH+11Pi5cH
TQlcEH5yWU0JqtTJwGicrZz+CkmSLEm5GkOndzJa+pbCePmsPMAQkysoiFOtpJwisSvdNZIneeM6
4tFQ9EPWCq8EriS8i8I2AgiKnfm1RZSROknLSF5JTQrVxIE7sHrijHNux21xpNZEJ/vy+pR7gvPw
LoChbc5P7pNlchp6xUlyMwO/B6jPArioRLpfQk6Gl4P5N1s9EzkErD+L4jhKAhaJ6GkbC3nI26Ti
MmkQkMaH7s4LuWAk7pwA8Ej2iZ07B4Z7aAlpGLcgHfiaxuYotcOcL6kXZUcItkupWd/GQ5Oh3eeV
7TJiNXp3odgumROjyxtqCYE0+NCHow2Lxbf0eoWYVdPyOPQTQ5G1UGTZqly4Hc5AywImtYomImNI
jRu0dD811UMuKGY8xVfzAVBfJbEE4j8aYZw2UZ1uwDDhuffBd/5tk3talSCdzacLyS869abGIpze
OnaT0XtP4oM1EIt7dQzavoD+he6ncX5jTT5RHvMTQugtQQA9b7qOKZsuS1r8ng223iGJ9+qcF8C4
u10Oe0SH9e58nQhDIxEGbcgUISGChOZQrigYk8deLJZsbSTcaWsmuOgwzBOqC3gHn1JvSCRTXrLC
57RlAeaXWMPTbtvms6a2krcoG/3EASLHE8WQhT5TslTREsP2BURbf6hF3YcYgb4qFh9pI/+tVO5N
fzOXbtzp+bNXAiY/84CkY9qqucJo/v767tniJ0Lbm8S1rmm8ZclIL2f6Zokp00FPbJtLNFU7pMIl
O688rdQ7OmA305nCUn2m8s0tGzF7sQbSk4e11/GlLRDiq3pfbdS2fvKv2Gi2JGJ6NDcmKgxfiI0l
XJpaf4PIwoCYMsNUk2BtIQWDYH/obxWFIhI0qiiZB1HgXBTkThNPfWVI/czl2Z5U83/pmJgb4gx0
0uPNyIhss/MeWS2oHafVk+J8VeTCce7YT62JSbv5qIvtTRb6gJoSLYsFDIPZq3TgKarx50lJiQJm
9zBkP4Ho+GnoiteCjUggnI4PF1OTzdx9yb+tkwtFYXJumQdg3PG8+q4s+wLFIu1rZ1fTfVFGSDoL
w2zg87hc7LOg2xXdeW9YI/uo6Vv8pAePljiqvS26sCpYKgx+XJrlXNgPswgTkXGQXEyKRkmNmoi2
+HxSmVXAM+UbDTMEp80v4AZTyRjL+gyrjcQLl6/rcaTsaxTpGvYA6e2Bi4MudXJAc+NSZ0EgwMoA
NpCQDavrsoxkrK0fRVu2wAOuU5quijDSHQdhMZlrn708/zEqJoh8Z5ewBNWRIR3kJwF0MezEmdm2
KM5hkdCCPOsmzZM72BQr65DyAzpZI+Xk3R+aNnI1lH3ETAe8hnozNxehuO4iJwICht/s3e3y6UhO
Ovgf5M5X3P8CfM5KPlxJlUX5QJy22YuJGW39YhjG9gjQL85uet3b/ckuYSWhhxmDR1eeETwNgH8M
yvzjRVPEx7xNDvtT8eCiiv0S7UzXHsPiHCfWVath+yLICXGcKt5xgOo4h8L8uXaIs92g7I70I677
x5gs1d1o8+FuBwFr+eFk8yTAhPRwCBsi4cx1YrDehWrLMv0z5XVeXfuZ6i/ZvAi0atEp1ZfYIBka
ZlSSeKKSk+wAgJnAwvcXHkXPHkrqCEDx85yogFfEJYdCeqgWIcr23oGuCsdX/A4J43+a0li12Vyp
ZBinCw3FtbDLQbFZ1kHBLEjHphSSHAB7rwcVTa02Cfzg7WRRi37im5mXcMxPG4HWyKaDm2EozOJq
yz9x5JQ25zsbSrWCJaUeIPVDdF14hiXZ+LRB71/3xVVaVPmxuSqo9bOIiLx/XDFgeeWqxBxLWcQz
rCGtct2c5Y2DTlLtjCqLv5mHiYMbvfyUx7N9u9tqpjK5vH4pPzpzz9E/pdOCRHVp3LeylY4r+AGF
ggagi3asibFO9sIsbxWL/Cx/d8aTKMkRDWFRINnS0EllRESYHKUnrwFdtL1X7D5VqePdoBiqEpiA
TZz4YNHw4fyvJjgv7OqxCFSRW00gdGmFh7sgAD+1ZpDRdRiQm7bcKgibsDBV9AfjtV/0xT+NyVU5
EUS/Rwh03P4vpqkC/cx21ho0PU4OY2s4Jb+2SBzyttur4Pwv2D9vnkvLFNyS2u/h7pLtMmdHSRH6
t5DF/DiGwneRQeXjW1xNl1FPGz4o3mwZrk4SbFXJb/StQmC3CxqsF0hwvamAgGeMBzrO5GRz1xUM
fYgVJw+QBG+phj4hYa1NUrLQ11f/xlq0XW/WxBNNxozqSvIyK7cTuTEun34jonz6XwmHCulqRzwt
IBq6iOsIGqw17h6yuW5hZ/mv+XP/Sq4iIJfVZX2feBTVgSO1RiRIrAtgaHlp9ZdrTbk0+S5d32EP
dYP04ZfPOPmicYBqFf3OrFZ8gnAXqyQCH9cvHQdiPQVJZLH7bV16BMWGTAdBD0A6aSIxGTffaxwf
ks6fu8istu0tlrLNXWSRQowQXZvZAGQUN9O+dX4tueeL6J/9mgIXEsYOXEEo+dy5NdmVBw255FBu
+eOWZHapdSBJlM7thStUDgSJKoz7BVofXds7yCkX2WZIUus6dmOm/h5Wki2hq91Sc0mQbEHuR4fl
AJAdKR5uN9Gijdc0y0mxuTfSG16+aWN4Q86zDWsmZrep33xEMqQqikzupvDbGnt7PMBUHepKfrmZ
ruB2cAJKPIQQvCgydRXGKfBo2510aIK9PM2l3LVdHOJj/jQ9EGhcY+CzXvikeCi1d/zQyE1FghSF
Qq4GK1UGv1CkHlFXSueak/D0vQMVvP/kOXA5Z8Bq3DzyYLnl46nY6IOEIU/z7bkCfJ6UCU/zCetO
CTmA2SMZaft3zBeyNrVWGrckpiT39W7TxZW5D+T39Gx+Zx2rXVpYMAZCVJKMZ1eDPJlIxv1Y5MXR
nv00irEfgdmppLsTQqCJsfsePNOYaNFCBHveiol0L8+0RbrmsF2RCMTZIb6Pb2gnIxnJYO8igoZh
s8uudlQgSRuC7zrp5CX5jj8SutZKQ5QmZRQWeoGiq8Oq3i90auYop3CIv6Nzemu8a7cxn9j7bH1O
dcI5QKm75MXHE0VcFw/bt9+5ZjXmv/+TwL169Y2KEiNKG4zHMKgaBBcaDuiB+CI5lZgwamR4qLml
EmA+Eg41quaqXw4E3mAabgPlrp4jRnYgn/SB75QELTj+kWmMffvX3Qj+eUwQRBgol6Uue/17MLJl
HKCVXdUPv6i8G8h9Mrh0XivHwGmfeSKaFQ4HeyY5vnZixChXhiEcFTKXua23hL5uQA9aoRPVQgDb
3ZY3wH5KjlOwng7C9uPABFSS0KPklGTHsQQvWlid3HD7af1/SnGv+MDYO/u/iePkyC9NQKzJ9z3h
lhiweF0ffQpxsP1SwiHnf/IWlLG2w5vfyTkiYF8rsAxUoTcBTR4NWTQtYY7McV60CsseKusnTD/U
80iLJbsndZK7DGYiX25V9C6qliDQRCZ6VgcNxvIvXyEgfllXtP3Wk8bb/b4/3GFWOGKNnQby+7a9
mFpSqPiKQrHwpQpS78d57tHElvJ9ZSScEJu9zpLqX2uOc9TjQePOFXuAsINk7jpZgbzPyCB8P0rD
y0E+shMFj+zY+4PQrS2528FnZlGvxZv0gpqBTYbG2tNn0fvSIL4x7ubjwk1N03ODCMTnR1wtgkNM
tbKCcdxbNIWjzt6fz0c7WsBYbABF9tjnMarq+3Q0U9uZOZ5+O/Mu0spxoO9khO3xYhK4d8SKWAL8
kYkE4aqoHLrxX6ErpzqOP03Qbo6BamRcSZXfdua7d3sFOfVHw4Ksruj5Q1PleTezy6Lk+w+0lxpL
f2tuYp2QIJdTWAG1RT1M9Og3Op3dxexva9Jkoiif4u6w+Ddh54PJRJBfZMaxyU4zCFfJk9b9M7vx
bA3AagyOPDUwxjio+hmbE8bmEyQqU4QIPdcV0/s7Z/ELjO0x4fNw6U3gObHWaVAONsfG8TQfEL7A
b8rl7ha23ecqGANLj8wpgHLYkSrFBjIC6hQKcE4cpe54boxr7VdAOXJu4XCdPznLLliz+oOCKlzJ
ReB+reyATtM0/+rYr3BFEP2L8HY0S3txfFMty3ZXfp3HjHPEox+Rl0R264cIIQrP02MS0xgYMVJT
ocX72Bde3ty3EeuX7CZNOw2IICOnxR3469Mb8B5ywQ3ladJDg+n6+Ev5g3ZaVGV6HA5oOA1e5KNy
8dv01ohzfu//aNXrhqin+NAPx7mNOWHo8Fl24FvBnUomOlw3CcofuB4H+XXsHpuoq5FqsWGrvRLJ
1fD+4EgcvL79fVeTEQxkHbhQbw1ZHnr/HWxcXN8NGEHuTNhdKCj85p/4IqwiGmqbPFE8zIV76w08
x4i1Wkg254uqiw+YJY7lVSwMsWrPZS2ID6OqK6oWx7r2TA8iYzAm8Ts8O346IoHu5MuJ1pwiFrbu
+U8P8NbX/QBxm1G+FwFKXJz3buuCvJooxIQXAA1TVvu0NNRDmL4N6SqGEYtEopR2kpcmTSLDybvz
KyEMh9Np1krDELsAL8zq+Ox3gKOU/eUOgx+z19DcNiqFQJGeZVR/8T9bjKVAM0V/cX32ZAElwPlD
/VIvb5A+scBvMdGpxdlMu0gxnd7sXQGJML8a8jXPd0PNgoGKyD+eWLN4sBhh8jSUZ4IaBi4kOPdp
qt0DsCCCAzVi/ZtckuWN5awTfi7XZvZ+0W8u8wHLcbR2K163hHKjdSRdEs+T7+G97phbx1iXjG/K
ubldzF1MoxyIi2tQdwBpJff10IE6uQLu/7XEDTflJlErQQxwwRqEYZLBJpToRD7hwwYKRDQmuADB
v1KBtLMmnkA70DL87A5nxsQdsWbs8MMz82B4wv+BDgZOoHw1smJAEoXIQd8uTIxcosOX6DPN0wsR
n74bRhS1Z5xciaUfzTGKdGWZ6Xg152zI4IIvfnTpGOnO7VBa978nALcEZdYfziUY4Ve1hjmYTc83
sot/l2IX0MDoONvY7aJ4jASmyyUfMDISPosc5JO39TuY2eh+48lwoqiLpgVaefRf+VjLBfFolLFJ
huutobHGa/bfX/AQZkNGEd3s6R7mwOTDbi++/88Ox3bDTlMjbMcbxzZ7/upnTFfNPVxqQym1SZ6N
d+aSX4gIxIq7iJzSQswgIlTjC2wrorAiJ+LfYRrsYbn3oC6LDoBxnYyuT3thTIFcf63cvLtz9SUU
HQFORmIhql0OLazMiAtpJK9RCAjz1UNy5EjkRpcmXhui5+lFllOa3toEKqEs/vJPrLYAjTQdvetK
qkBXGr7GNA3BGT6Wsk6wdlaPuhAPUBbaZ+S8WgNIjA9JjlkC+CO6LF0Vka12XY0Hox8zePJpg49b
5gwj3CrcTVawd24fI4BNE4HUZ4bAPaSA2tXHw4ZNH57neMyZL8YnhZOPbNS0LRP9MeUUG4pvERzK
VImSzVUPhsAa9iV2JoUNNFmiM8RuFwXR41wv3eESxbQur4kM0X6DLqhIiyxS3EvbC/wwovSzAB2R
a6MknPlNe72nOfNHzinvVVZ+oZmXw+F+zPXGH9d/T3t2d94nzseOP5M0ZhceGYLzBy0m8bp0tzs+
it/sZ3t51t9oO2M3TvJNLqEpGWT4xNdvuKE4eef49nEdefm24ni4Y4W1RLgk6xrqVfGRVsmTSEqL
Az0dJLt1AEmWbDXOlhaq5yIyasAogppzD3ImD1O5tAZZTsfe13p/8YCa5Tco3cYP0Q/Z0EjuEDm1
z2v0jWReoekwWdKdo67e+g33dCqW/rHT3MzdUE+iqOyv0CNt9aDgqlXayDbQwxXKnV0dkDVqiaP3
InvHgwinfC0Fh4RztnWS6SsYf2iVf86tLBmXKXY60h+Uq02n9ZTi0tOFVIhg9osMcKUgJrwowdd7
JNhAxFNxVuy6v2ZcpDQWD28j6kTGrKP6rZgHYmoAA4jfvKyL8kLYI4z2ucIxVjVKumZ7ZBKxRPas
qgVxsSyrKMmydMStEfzBFrF3rUHOfVR8ysUyFqocyu2KkSGNKKOr3xtQvxTlRe7LcRumkgXx873C
0Wa6z4Tt0eT9rkrNVe4a8tSwSgA8O+az8gquIbSjXNp4w8riE9BuLZJsAPloSfMjUXrizbvs3kRv
OkJK7lXwop40LYrUtZNR25LFm5xMVBWXdGzsGAVstZMTJSW3UOJZMZ9SbzPMSEDrUId6lfpMQPTC
T7B3RcE8LKqRwR/FDPgmCs0MFbnHdFs35QMW2L1DtdFcqicQKQn9hT4SQN5LuJi4nGLW8jRAHaNN
4tKrQSY69cljRGiiI2hYtJCxNKDDTless/N80YEf0CV6Y5Lq+0qK5jEiTPTkUrlpztpF8maVjV/f
bNSvAwQTIATO73Ef0CyAFpyfmg0j6GrLB5Lp5heGupHRq0XNnU+H8xESBY8KY0ma+huKJnSCz/Jg
5y0M3f6qXyI1a6gM5yJzSY4lTKszv2QcHUjmxZ+d0EacjPJRFCzXHVlMtwK1JgNI07Lc4AG3fKgR
4Nh7lfNTJCKh7Uf1YSLaxk1DffdHolVChYo3NIE8kAklPlw/gNe00YS0LopYLxWLcd2CTnZFsLdP
5LtT3qoF9Nu80wo8KZihFt62rJbNwthQHDR9LHnIAAzjW6RcdbL4l1p/UOHNty05Vn5aMlsEu+yZ
rxThaWYM+Z4gDouwv1O4ApvXx8QoBd8JZkrwB+xn0NXsnp+Nf3Vj1ckcFbU0N7OUC9FHxtWjcZXf
5OKOd+qklpqT22wcdshVv5mkTPO9HpolTfUhYkdk35v674tv0l/2MxP4z69gdOlGv5yWQB0WLEKT
ROnhNCcWeU9OyplgXrPlhBhUFTPGf9WzNTcUbcevgNKKAx57OKTbL0Ab4noIRwzWKIajGTB3zYLU
T4k5Sh4ctQ/4ZEQVY/emzbQFpBdrcOinztkyqtyaXv4yyzwWamAHLuSshTljWvKviFosyqyWI34i
v9ZFFce+I9ykByGQ9X8ibcNDayMPML6VdU5njCAf1VnuOyKoXB+mkSWGLGy2r+PvKmqW+20Z3WiB
0Hwf1q0F1Ih6bwGPDtXV1vew0LKCIuXwCgmtEwcT0+QeMM7hHA0YrsExUjYY+OPeVh9w5pT66u76
c2FURJrc+ylUf0I3fJNTqN7HndC77FHgBxou4fzceDhhumwtqp1t/J4cEjbAYhrImDgZlOSlP/4q
MC/JxgfqYrzhjUA0aSxeDoo+QFISOLdZJAfi3Hab/drHFdZSom7tyYcO4LplXZ9t3908lgIbuJ8O
xNPvzghB+VeMLtwj2Pl06dA+toHc3rS5yIlcrjASYvDDDmcXIrmCpO7QUWwnZ0T46AeHDQZGN5R9
rt9Bop3d3moB05Ly7V6J4Fx99GVBAWLZvjGctdu9m6FG6kx5EVry0uY5EPEaAgHD67UB6uvPlO+2
bSuU4i+RqUKiiorp4cZq43duoPG71fcmEFqhxHLSwOXnU6DCFqRe2lwk2cxDNAybo9BSVihO4z25
cLkgmv7Z1xh7EI1rlj1ofaQvn3oAWYENfEUrLLCgVqBTlWws/z6npflDVqehyi8mI8TmEcCivohT
ZjBhs3URPIUYcJdDOM58EzzU5nIHEWus3FZYUgh8XayNGW/RijDzj5PDx3m6Pp+8+7UR53Kk86dJ
sDn0y6pSXGuN+w++22SCXcnJLmO1cf2uDxZvRt6tYH5V9X2U0/VqIsnOQV9ubjT8PP3rPR7EQXQF
SdYRHK2pv/9JHC2DVfDlQxW3H/qOlbAFn0Ra1z5jLAWV8d1obHyqgD45jHzjfhZCrqstm9smroqp
qjtCybIMfPqx0zp030KxMkVh1AdYH5IQVPqcxtQc7dJV5zwqs7khJwy8bprK0UmsJ7EhpyEvN6Hj
LXyilpp+Tv7WUa5gFGn9SJGPo8jV041GTnjPZCXM5aCk1DUymnzV54lBSM+AL/4WK0L/m2cWyujR
uV1WJVwLfbY9lWSbMN4iU4P5QAWM46FmqSIbx9Fyn9O3cKQ2ON1UTIFwQOG6ntCQs1ukBmVxM1PM
yaHxQnw57NOCpov4HZr/OjDrfqegQOSHTcObG2JfSc1GA9JEYeAVK9I5HJUHX4KZu9vqvEF2eM9w
TPriyTAgnPb/gNlvCNNufeVTDjKWl+mki9iolOYFm5gGo/iAAr2j3JxoNBfnIVcsmvkUFxqN5FlF
TQbwPKnOYcbDmMlrZhpyZjyKE4lIypnb03y5lYF6pmJu0Jzn1ACJEak8elGpabCWeCN4uky09LzX
MIcilgKk7QDBBaiJTV4spy9r8xgEeZrfruFdRm8Z+u4dAxwBV9stSV+IJGqBobMS+ycxDDNJq/Lv
v+vo2ri9LwXBkSBV/kEUzXKWmuaBKUbmxZ39w0Z+DnL+yOZ2PET9394KncnVEvJc0iukge3+iLV2
8+m0e9B6vvotCeisk0lp6Pafzwm9NNdjJS9IfIdfudzZl2iMl1zeKGYLz+BxbDESrfzPkdbo9Y/o
TwctVJ5tvnsEY8bJ4XSAaozc2f/MK09wkASzfK6+uAUstSY86FB7JNIaq2bKXOZzbllrsyWXCPTG
Nh4b+ckyt61HltgYp12nhrB841bGZvLDp1eOHC2hNBPRsEZ1ayfgg4UygzQgxqM0gSTnMkrpc09a
iysCJj1qyyxpAklCnCU+Cqwqw9UkqQrgyCs8MnJZrJCVsIQmRh7R9m0IvYjBqNJV73S61ChXavLW
VYLnuc9ptdmBGN9AI8thj294YR8XDRBa28Y/xdBN/vlTOEx/hpQXTDl5Gw4SSqeDbvVcNgKiom7p
5ebYdMYw4Ek+ciha3a4F0uqhj4dLVcs/Fy6CqoKpDXrotugrV6nO17tDpcLsZ8wFUbS3kYvEhOrb
wOs+2VvjU9VvyECfEZceNu0HFlDa1FZjzIDmG1ro2Knj0KIc1N0tj37I1YEugvvh3eB5/TESgt5Q
tewCcxhBCYd0IVsissOHyr/Ql4SbXTR3ZHW34xA/sgITNMGHcBKCa5PK6qpeaBIHroUdd9AwqXf7
GtNj5GRM9OvU38qckGs7qeHkfXgyCl/Moi7gVmMG3GOBeM8XOcIGcPsNXEA5AGScl50dxkNQ1l+8
J+0U82lGF5QvnV8/bMTWJL+xTh4fPRZw9Y8NL/+5d3sDYjJufHgefCK1SbmIWEjfU1rB+1bS7Jub
8DmBPZQa1FDjjtdfpG9Wjct2BTqHxmCogq9avseoCRQ3+jjOWEDe6/hXuKIZB31yON74E5MSSqQO
6Uf1UsFL1/s2+zjlUpANsDI67Tg+tJJa8s/YkToAbJwyq4SqrMoMziLdY93bqIbKCcJyVc1K9eYj
dzlnrA0F4HxfJ1OmZtDal3yO6duhNUiBb1HM0FhNyiyRMPYL0e8Fg6Y8u1GEHNoWBoRDY4CL1FgN
PEYVwsCuFBcCoUZjiZMnVxmerGRNH3DNY6Fzd3/DHQYJlnI3OsjGnZP4cXeV0cJuJYbRzQ9BNLIt
0GLssK3qnzIJwFABpVR4juG8RyRtqCfb0AhVS41jHG74ISr1S0wh0dc+S8JwIbIn7Fa6xn+hdIvV
dl2dhzKPqGzVrDzqjdd4IL563xT2sjtDSpIar+MsErTZ8aOc4yltwJgsQkiRGh00EOHmEHt50NFD
MuXBk/mDWmvnZ7FyROLkBRXzYH7twkPeqCOJGs6tI+gnQ+nu9dAHT01D6qsaDFxw81NRq2KNEtA7
VN+IRZGlKDZVzFZcz+JiuCShLm+r0GVZfYUQZ5i7Rxu4fD5V20rCXjfvPj/6ocf6B0Vj8KonhBlL
q3ExgwJt+I09gUz/1je+HXi5FT0nLa2FQ+2IwTALHLxUQCYJFmldjgcXjYFeDzj/EeRJnyeeKAiw
Cp94TXmkxXXyhmAQ14oeTAPAvqk8U48pWS2CtLq1SWuyVm8EY957Ko50WJFte2lUdLwZOkk2XPim
gOQqBw/Rk86O+yqpO7dHiosSEHlL+BlT5Bc4C5g4EymWQG/bvzT35GxywF6MmVSioYaQ0xqxBYmI
QgeetzzRuCdVKr+M38VNEx/KhaOaseAps8atwKbfR5Zf7/g2S6pOKKZ5rSdGXKxgvhUhxgDHpYi1
pqg+sb5HiH2ZnGcPDC1me198sjRA1i2kt1ZOnUyup25PRnlUhUKK5btxlNgWfb44PiSbjqoCO5SQ
eHNbHXYniAz49tu2FFMboeXvjH9o7Ja/1KPvkAfCibSNDRGEN6CBySWY0alSTp3nUIKFOAR9HXCs
Uh8nDU9AOxPoI19R/2uUqqKaczkHE8wcKmsVUe0GGP7FkLlM9Ow1pvkwIbsRciQvdCkJhQMehOwV
EYZRT+2b9rKw/Ql+qrrLYxTzYLGjOQgNV8vY6xScVhiZNZXAkB3cgySY6/an+CtH95t+xBqxN9q6
fB4fd5NkJJIavPIH3SePIKw7geFxR+9SmMkKJiYHQrti2WGP15pM5l8jO8j27Xc8N0uTCZVietnM
oRqM2kkGOSESBQaQ6KQdLHCRJmJSecLpaAqRJ23bMMX+bRhWfbUa2T11qvVEenOneB962wqnKHg6
8dcuNUIr4BglXsS+phehoSC2hP3U3lJAnjfIsR8hwHq1dVwadkKIUBRUG0VkJ9FQw2CyErP0/6dE
4AxhcXiVYfPKUItjb3JSiyBY5FcoSu/u0vhALdSNhRgIDAKpX6/J48r5Z0VF1pljjp4hF6UaFCVy
v/BuabgrMna5ascS0dmpkaPssmrA6LaCl5waKURyROfObhPbT7WDi/KmrP/Mtk0qyDsAjFDiQQHU
pw9WkmCTpjLZPxXsSbkHJiP1123DUSTkNfDdgplE0SQVDv98KUtH7g8yNVOKtCK/UFkgvY5fp6oe
wD8Ge0yaqZ4NzBQ2SPPPERNuEi5xWDDLdCNovIV5R/lFEEObsnnIRzPITCY7w4quJialyhFbAnM/
g9QfnLKtnCHpnoHFD65Xgc8XJIKJko7O3Ld5m1pQpvtihr6x0qGl0/oELAmqG5nQYnf/pMigIjuz
NVtIbLn8mouvEfwBxxmTf2xZI4a87+IbuazradWS5xSNIlEa3h7spg+M6/woFVHYRnvIM++ULQAM
kF5RvlAWMFPhYHCbtrTCJ6ixDWFXfRkeISG/ucQvWpp+Q6OL3/a9TkAcKwk6zSVTCLGoyuDs/yPF
kZOf60Q7m/S/qAh6zHex1MoOYRDU6S5cd7Lp3yMTK12PTsMJk1LhAHWT8uAZXRzz0KuvP7N51F10
iVvFurYzFU3Mg60u7dK0Vuig7LAre5cXDeMi8j8X/bvLaaJrl53BriSetuifqNniqWBztZredVxH
SlklrmreeyprAhjeUeYCFbYBZwGJsAfT0CesappRQ/4iaI5AzPx7ZKDxt9N00i/iprI/tZ1Usj25
YCVngJDSMoN8lbuo3W9aoyQlklqKt0jRj6acB1U1bULG4sF/WhlY9NO2ti2KCnKrh4/Rm3F9+Crp
Lv2HMT8k1aHP8RZp3bv85OongTnXKy5iaTAOjLLFPT+O5pnROhjoZtHVdkrez7l8IjdWNA+wY1J4
dNXXSDski6MZv5fxFHfef5R/8AaV4zIn6CwhamOQC6OFjpugDt0TqYa+BjQfU48ZWkuLRYdoV4OC
TqQpACSZ1qtHhrTmBHHxc5NN0GXiLCgw2j5kpk7CiaV+qOb7pp0UY9ex+KXvDgDH0fKLplNZDmnn
9FjwLXByFk6bNXWknRmCEgb1agHfVa5kEN75f+hb94qpim4hg7b4ExyFpoLVC5zwdhuQgzc91PPS
Fyy6zxuoOhWAGmRKBe1dcVr+dRNcMbGorPFzl4/d0g2UbvbIfTk8XuylGMCjNuKd/RwEnCavOCQH
zz9733fYWOJ+bnmBICGnn4GdiMyYoMzY+RGuZ+CYWWPyNWGzFACq2DQIod6Qw0VGZnzXzkJK9JsR
OmWgJu6fTxj6MAml+uMIaf/pOhEd00rgGK1AwZ0ttz5YrzDs+OBn7LS4IZ3lwR2M39+28UIl1mOC
zuAfRZJHaqg8mouA4KU5kbJ2/U3/jaU4Le5WHFJb8Qw7Gakw8AVWt03r5P6QeeWBrvMfacZg5pt+
E19mbYex5lf4oCHNlvI7q8BnkFyG7UjVHARJN3SUNHvbSBpbwE+WHtvqHZ3bFfpVtwW0Bi/2MFa7
f81CNTA5s4w2rIxDy/BwW54SBq49PUAAE0clZrLREFJxt7qNnkiITd3FzdOsROTaaXOo7EKht0rz
2kEvrV0x09WMfCdRb65GAPiuspL5yNeJvAyfisfba1U9jbbk3a/xwaE5xjoybFPj/W2AEX/SQJ9E
h589R+zJJCKY4yAe0j4ArVOEFUxsUvUnETbWESTq+43kpsmlHkY4gsGvKJaLuFovZSJxLhkRMXYr
zTOACSRlGHnEgcAn/suKHaJpZkxWVLcge6A6/TmS+fuh9YFxP8H1HsYXY76nGV9E1CJLQFddRuMr
P1xNndOzWQCdkR+erF5eJUYxRyBHcuWec9hgz1icH3mFr1KVV3q4pvSnNZXngjYanrvJeZVpWTvD
O7KfJZ/aFw1zrAyxK8/RIErn9Y36R2QpDRvlbvESvBWWANSlpYrvA8TT+3EJUnI3eC3odxS5imOs
rj89J3W7dyso47jBARwL3fNzxKs+/MUmbx6NKvkxJgiJc9f9Os2gSBqQS9hfPmNrFiAr61jT1qWt
3Ky5DN8BVJV0V+Z6K//xmlStr8nWIfMBMztTUPs8PU4YkhhNQ+qVDEqtS/lqVzGBfnCUKUTA+2D6
nI7d7kUYo7o5I8Lrg3uDHAdLde49+R4khTjtThSBStfizyFpw8tCEePcFhRQNDQnDFPDlx9LK/OZ
CCZC7gS/t4Fta69JZgWgafKw9cavq3OCv6S2cXGphYUwUS3H78zwOHFYCgvMcoUQ+6rdD4uKmTCW
Opj5JBkMb4s6UlgGPe07eiVZNIk00We7oBbuDS0ml1zq1o0zBGpEd1DghvkW1wJYo4l59tLe2RC2
KmmejFltgbeEFO5NyJLr+gpcVJ/t4N7Mp6tx/W0Z+5yJu7g/aekMNDKzTWpIAGiOzbo6OrUhbjQA
bTOEQM9KyOUgmJMvkwV6bMTNzV6W1wz5SjlEgETIq7t6mFLsQK5xNwECBYm8sNH+Ss6vBjCaJXyY
rHe0+dDPNrNLVMB37J/aybusuXzI4FmppaaSll8n9RQHSfhGOlUcJtKLzk1aiOoZ9Rn2BlNT8YBE
3w9STWvmy6jvfCd1Ci1iohSjZubaN6w/nDSHg/gPa2eWp2mHanSFDlTBow4u0M8RZn9wK10hX8B8
kSWhL8Tv3KZbcdoaMMGzQG3Mk099q2ilAEPUUt6HxWUQouXo0xc5VZdqubciyJ44mG7y2RdCbsBO
sOR2zVy+QJlIPHnJXQ2+IxvWvjBmPJ4b7Q474CVQGx1uVwHvjv1UTjICa66jS87jx9z+uWoIfsxs
J76zMQkhOrtbXZf8rngHjwrd9312W53DRlmYX3QbufzB5ujBRv8wHYEv+xbK1iKjXmD8ZKAE77aZ
xS0r3JAuSzegzbUPXK4H9w5SZXDzMEYQcMRCIbcSMhYp6v+C+UW1ak4WsckRN/9t26YNnn3EHExo
WAoDTd7caXT8A37nTQRMaKDbXA5jNwyF59nQWht7aHHrgzA5ac88t6fffMCVXqHDr0O0c+5VyhHq
Qwm/5zbgRcw2ShgVN6Dql3GpCfwqffKZdlABf5P1QBn4qF+aTiXDeZ3S2FU5glKBTHhRMu5dhYTt
G1rUlLwZjnpeRhwkjAU6lZNN57xa/XkJayW8kcWpRNnn8NF3TQbUWE9bTd9TUJgNcmssraugKmEQ
RvIL32MHVD2AetUWW1tcnrvzA97TjCiWW7fHJybiyegjM1PwulmDzpT8bmDm2L1MDyfE+urQPE+E
zRMxTNGdqAo3BOnY0fbWCalW4kXVT5eA9yG+okZOWHMYnWfunZrrN9GKjsbMuxp3SSUdYwuHO95L
UZJ4+BQGt26E6g90IA1jr21dYtwfEVofP6ZJBGTSaJMhSpxoIuryL4Qa6KG+wCWE/C8oh/drJ3AW
5ED6wRDJIckzkwJ1FZv8EJEhMPuHzqrRglnpMvA4oyQ9bkhQPYdgfwRnvHsBAajFChRvGFP82y9B
S6K3rD2TSQ6TPmQEkurllcLKHGtfJX8e/usDOoYApVtRJCw61pZHqI6aRCuTS1iGdRASMGrRa2iP
Ko0bI2siaxlrEzvBXOMlK7+vbaAd53p+OnTgp6n/C9SY9zZUT5bXoi9uQRBCZI+4uPjrob66YeZ4
3c2Whx44oCcQJE/fEktIViGP3ZeJyhuSm7X8yovMKESnTgcQJsC92wpGz39JCbcBOgET6MSj4xFx
9FiDoa3kIrH+za90NfFZN0YemeXRPk/0zLXaW9ZH+/8jFNCqE4eeg0ROqy6rpK3tvCHrzUdSJyP/
6mYnwYoTZnppkme71s8plw19nn657vRmRfJtviq/myc9+PqqYBw6cbk16501MK1b2KoBewfwLxuW
F/LMTIVzcMrdHE1zVu9UZfYX+Vtwf6cx6on71hT9k+bllmhkcTkDVYRr1HnIdGK1touoM8vsX1Gy
E/xsrPMt2RdjjPx4pI6JVKYgXSaqFgRH7kpVLp6joc/cHBsHyuIGAqLieFM5OjLtSRdaqLVOE5po
ABY5IP0SoIq9GtwgrdEFatOol5nT8bBvXnvHEs69sgJIrvz4R6SkMel8rYnFz9ydsrvkSNcjatZQ
KDRhBNC7UFErETOUQfi3ugajaFZz0dTv+sh+w196a2MXQ4mwsoRcPhbjbqBceLe5HqnR2VBT1Uxc
NUH2iEaEa/0YGtC+iQNrHAkWIb5fwhTbxMliTf8K1D9GEpjKqPMiqoP0mvlskish0kbHvrK7FJsY
H5VBvm8DjWKHZmY/QyRDcc0tpg2Glj9QVyWfXm1AL6YAdemtEs6lYKjdD3tlvwupoSjeBUCEKqha
3BYboyBKlx1mhATlR4Xzy4eNLbK5KBJcYGmqQvkQ7NlA4+gJ31tkjQfc1qppjd0TySfTsuTNPEr3
NUxe+Eh6eS9Ve/lBgQXYfg3SSeUCLluG+U0o9KpSvWTgStA6fmEWxl7FOIGKoyE/5Hj8P54a2T2Q
QUcO3FslmxzN/emOFfDD0eMrQqHVf5ngQg4Fxf/nqrABfGP9BQCuP20+9aghkX7EHAHGXnMfYt6G
3N4RLkBSC7CVffccpsWjMgj9IVaE8LeeLrDT8zLybEQd81kNigsaNN5PFyDQCZzsQoA7QUDExnxW
wZexmG7fAjWB2GFYC9/1QgU3N98Ah7O/+weI8EVJVc2iGR6u1pM9147sYiq/cyxyjoD6H+204aoC
nkMF/bkAD2xpzO4YNoKqYmzwb3yT3N65x7zQA85EzZ4TnDSNGZH27sc+IAkpprjLpMA/L9oMYd1q
/VWTbYkb35Drrcxv54A8FK8a0+jdeZ6gqbSBCTjM2AKuPlB0zjdRLi4MTf/Bd3wwudwdYtRDJHQU
zTEW960jkzkEKYNDvrlwBHsuFqzQ4K2b+0KBntKh5cwFJkcaa7KBp6CSySjPTBfkL/fpBMROLzRi
OgigQzwuMqMoywSU+I2OxObSZcPpE0Q47RBpv5oRdF+/S4bHN+BKezJj9D2kGi42poEkxSXjsEyj
709+HyCnPlm3MbPyODIp8V7CKiB+4rzSL8yS4HBWEeGydRLbDJsKD2la1gz8JoAD8D9R3IZNebXs
p5aEz4BAe88axmFvd5GpAFPTEQXSs3/w4pWYCJKVgzNpeKnx1wF0Vhx0f2ppbtfJFudGqFgQ4AI1
Y9PgI+Ein3FW4aJv5TJTsSLtKiSzzc0XwGEVwAGNxBV+abFW2/sENhFl3tm5oo3Vw2M3tIBYGkP+
pONPDE2Qwttg04YYym3G58zdZz+v1rlugKVIK/J7xFNt12qbCJA03B/B1dENgAMovvGa5grIBa7h
QD3Y3bbxgJH+HFUqh/W37hPCbLuJrd+WPdDXoU9dKf8AbEs2HlcM/slL0qNis52PTxlX/vGRwuGa
lqlOEuCx0nxFLOtBq3Et5GTXxhqfzYjD6V7xMtdhxH5tWiLa3qHUyPnA7fR8JfVQLoESBnn66kHQ
QnlQSI9g5/OxkwBOW0iPXEgL6LSxOYFvBdMLkPyKyZ5IhbzZPgFfO//zbBLZf/aenvY/VNiBwR5J
BDuJDHLlSRYvYfk56+OGY/cz9URmPdEZWs1Ou6Hox7rFIrHN94MCnV0CweMBhs8355mg6X8FH45T
k6dvL2pNlSFUYRrAIyW7ZTEBshmi8VwkE+KXS2Y17D6UkVzgAj7wwPG3/9UFEVC8dkBR81M9c0zq
WAQmRYqWU4b9COiqJHsTMXtgpqKFn0iu4POKAtyJMXapuxL6sfKMVQuZcTVMZ62/Ljbg272P30/q
3KWi989JSqy6bOjxCuobcadNJ0udCGUgTI3MOxV0IjBMwnRRRmazPHGgl8F0gi8RlmjrkYmbcJ2x
f3q+SYnYHVxkvDYM9+vJSwj/Qe7B/6maT9gHv8+8j5I41FAnh19SwXoZLi/Ov3twsnOsG8UZVx1e
/8w7Sq4ipNs4vj+axyxcfhPJ1dUfpdAJ4lJsLQ0TGUlrhuqynZ43AHtYpPhtghv8ogB9m5T7AocG
X8+krDRvtfE+C4luZ6iaDRct1vc2HRaUAFG2L1qVh9Lyth/OZJizEergOKkPUdVO0JbB33wm1Ztm
KptwcIXu4viUGCyzBPueDiWgSF+ZL1gNlR7O8miBvwgOwoODvNsiv+2SZiYvwHu+qT2Qu5PtanjG
wEbRyQy80RYbxEwkRT0/NNr0rY/7vGeujXwzEUgyK52H4BiXwP4TW3SLSx+IsSlKgVhson32xSbP
SU//sCY0SFGhEveXGXhFMEF9HGxzhSoCB4o49H6S36ZYeUTiy/MuPf32ph+QFv98crhxmVoav1IV
6JJJC99rLvnLCmhUvMJbAWM8EOwkZUo5YQdeJgTmmprKpQwy5sojY5wRkkML5D+0E/WQ+KGRRs3m
8X2yZOvQmfvoiQrrVeL75cgA1UCBOwFgNiykKh3QBUEsZboJ7IYvpJ+Q18M7ydyIv4EvYQYr4dQO
EaUPEXCymWXf+S3u/5Bnmb2COe5r3FqwzDRGBp3wq9w+mmhrPmsZycEFMvFH3+YwJnxf9zXk/dlP
i8OV+kQu24pKtn5YB1k8mBVAqKPWgVGmiC4nAWRnBlxdi8pA76B8l0AfWaJ3z1ILDoBv5Gz/nOfk
b818r55DlYBIglet1Qchs4UQsRzqXEW+41cMHYWY4C6EuyeOimVHVRGtNTy/86392EPEo/aPsDsM
tN0/DqNvI+0P+ZzXKKEanw8WgNyjGUu5CXPI9pX1CYhOelSS9TYYN9l8kHgvS0CPi6bsK9zBPFCN
jcbEELkokhV+0WZIK3IApmPj9iHLk1+eUTCWhG6xnfIXFRYsvuuzaMrm1l6/j2HplX5SeL0WVt+N
oQk5A22x0Rs4NLoWxvEGEqwl8L7ued2XNmRNPqF+QctIUYyQPxZi42AsY1oNMtvZvPQTPRPm/S1W
jKTx7iNz6S0YiEMhGhFZhzuL65ppyYxHcM914zLIFG2nSxAUZBRzbFf+ujGpP/OOyEpN5WKYYxoH
NjIsGbw7wqvOpENBIGF5wPbDsBw6nfIqW/rBJ5K4U9xqBpiYFoWdgbX3hdy1atdXXciDBqXEK1OU
Ujqt2GpipsLxb8UMECYQdVi0BgUnyZ0R2aTq31bc4WN2DIOFrjIXI86zK25VqZifgrrdaLBeQiWj
N/YO8detIpesefkND/GakkNXmlLbCDTX85Xh6u4Nt5tjJyFcsKHNyWBbin0l3pCFNU76A1o5G6Mw
He2XylUTYGKetLsakE4Ar0DI+2cebnekV2AEX1kSLQeaG4E5AMZDRSxARwd3B4voZ4AnZkY+vZUu
nWR6BAFfh82uHerAW7v2uHqDno3fD86kPdheA0HnFNTTNZaskEkp4MEbTiUxRfMCQgo9vXJ0yAXA
gTZ3BDf+01BU8op6uhSwXRFMNfS6493Hr5wjfKq1O8ORV2Z3KfX1Ho4uONDUIiIwGRjNVVZMnfvQ
Pf7pgAxoSSIq3NEBV0qfMnhiclov1p8r28WQpyyT3pg7TMYM2EBU61GUuFtHJnfU3sJmR8fEBUrF
5yWHRWBxiH5Updv5S/D2aP2WKVd77VCaY5i+KvPcc5y2SZIjwMsI+0dypwAdtN6GIu9R6mKmmCXP
0vPyE6knWatxswdixpOP6N205Qhtv1F9XXIBBgst5BXw3yuC6VBVbDN5LO6H3VUxysMRLAXBQUgb
839Hc1x8q8ImGMPNgAiUZC+JncTPYnjlhmcqrnDe0Ky2WwJ1oDqfL8/rsj3DPUC+WB1tQrX+HcYs
Pib09VtLdL55W76KfaBR4aOD3OWbUpqBfrbPYA96/zxh+gJRrs1kZ3RwTK3nnRIL3lCCOQDNcKRj
o0OOD1lNQFr3gGUt1pGYWsPAyqIs7yUuZt+3XEIhtfZqt2FukXlQ9iuIcZa+obyi46GNTVsjUj5g
KJ6GeircaY1SqTpIIX+ZOg+ap0I0zCUJ92aP9VbHeWiQY64xPa8sHgbMHNCxDm0AWZYCndBzwfWF
1FBY6M5LF2tye5cxb1MjHRaRSdLjLSdQDI6+2avhfWIACaathvz1AW/XywhGOVLZ5fu4hscJxOBE
W2HmxH0IOgS30+b6g2lYCqYD2hoExFZs/ESXkYCY9zAJSAkBKd8GNB/CH+txiNjpiYss5kQfQLob
vUFuwKfsRcGh6admiXMSQaL3ieA3vUR3LON/byJqeNTSn5pLqEy5hkIs2RlnSOLGJjakoc2OJXN8
vXHgbznURjUvidffM0ZeJKNCjcseooaAzAhCj2gvhhv7kyjXTpsohAE8bU4ZZJHW048vZ8ud2/Ba
eVFUOQMRj98B/nDNRnU2K0dU1Hrqkefmc1KeCt95zyLb2BdA1wS70MXdRYau3mMockfGSHUkzY6x
7Y+H33MUCxqX+UrnOUXV0YIr6CJmBm9qbAwgnF4UHF8l3wtky45ayiKGrkAiY+LwGu7H3HnoimF+
q/S2/4mf9pGljVtZIg20wUCbtENezeUUmgvtcug8chfI/KWqMQxAfBgpo0PdF00i0HAI0sBETMVd
7Va36HNBV+0zx+WNy8cCK/QQHmiATqQrWs8djGL+SBUVdaYQ+N0mPQQlbGrbvZVvl1AT2PMgjuyF
3BeRmaRe0q5OSdgD3nFB0fSz1YXkiz3KG0W6M6iFlCql1ZZsq+t3vX/UN1Ij3ofKoow1OJ60H3UQ
9uftWCeL15EYgaxCEW7B0u7W/ch8cn3K+c1KQb0sdkCNKi8Q1cKxZfIAKlo9rhrUDbPHw9+TZwFr
3Q8SHMs6QY/lrnqQHO5VOdtj8Dop7bMLW4YY6UCxCMCisyt4kki/tmw37fwBFVLK6KthUYNqAGKs
aU0FUR29QORUb93napY/goablSYT13nZwJ2K7Vf9xFm8QbGOX2YB8VnHC49yXLFeSM2Ji0pDRhzh
hVcPqR2Hy7qU2DYYhKF6lwgvYcFU+SoO2oPZxTwM+D0FV+GgcTBdA9nUxNx/FNosye34RpEzmppk
GcfaqFvpI9Sub7W4VF/I1KQhMJ139m6oC9aKjFx5gWGQQilPHfOZkWj2eefTYL+8zsh5CGDiIhIV
KFsNsAIn7TKYAtqrR2K9sOt578uzRinb0/YmWUlbWHaO5A0AEhK0C9fTi3o3KUFaC5aH2a+tkx9D
QrOwh8akdfuIjCWlKWQWMblnfdksLj+0yUxE19MeGpdLNuSQdxTLxaZp9L300FHvbQdbuhll3oo1
3Ivy1Kis+8zwU6U8EkhYfeRiss1VImOuVE9JXPjWQH/DVEjJoZNwN1xEJ6grjHK5l0HfvNPjcmyx
dS9wJW8s6AYUVDTcKlDMUkgtou5nJ1G773g6QqLnFRFWrVK1MUaJ8Q0ZPHZdVxGpV6CIJLlUfMwp
7LBbOhfZtnTQe/e2rE+tLKIa/lLq7CCg69d9G26DLP8RLvVcjklVPrgff1JhZS/PLworGsU6vF6U
4FW/ozRQxkYlqUN2qQpAlEV1mvrzB4/OdaKlmOaHtqHinzcFogoFE818n6bdvhnofX+/WRfGAaRO
bSgiwc9rAVbdz+STrYVz+n3/Ucdzxc4K5E6IPy89FaM20UC3Qd+DCn9R1MeIiacNypjuhk/j5K/b
nRmjpBZfkn8TzRDli7RJxsn/B4ULMiLQASntvJzLhhn4ds46vIWhtn36XiIbd/AtS9d8D1XxsAul
7JIIcn9fQsrTN5jC4EdiPduxPYFkXRrXQvRaPQ7J+sKkEzjbIQFxqWAkp7pBX/B/h2OmvMGmcsA9
BQTquFA2Az7Q2+Ep/axNLJ2EEGn5yyb0DuqQaeDKkynkMkJD0TWvgZQmzTzMiz66GzVGvDjJERLQ
H7dBE1pmYcl9ILkRZouxd3zha+QJyillGD5yN1xrSnUA+AFelG5UUXKToI8zmJxv5dytwPN7cMXm
mx+0tczMUbfRUmQA1xruWLKgCD21Tif7fA4zllTQzvNoIuiAnM9kFZDeH3teGaOHpg/XNkqgzwiQ
7Nm52DNTmfZY+Usv2BAnYhOq1nU2ozwOgqR5ppk0f5e04v4b00emo6RD2aMMT+ygobpMXnjIMGBJ
W0AQZcQQVFjAZjivE6yZN3W7IEjRYv2P3WKNRP07G3njoeYe4UPHw4queTrQvfYY56Vv6jxGeR7a
cG+sgOslQiPiVkx6SckFYhMEGme0LEs2jrG0dlFlsL0hGtzkICaERcZ4sNTcrNk2CNIBSIU/Lrup
AMptdBOIPGVoaleVfAf8YlpUhXQ/xB0ZuM9VLlxCFYzqgONJL8ciBTs3Z+mBiH2S63JUyXwyDMy7
CHjEjMLtN3jYMOuYK5HvmB3+GjQDOV4pSxvp1gBEjE93faaylrc5tocPEZ9yETlPP4Xf1kyPKkoY
C4g3XJ/iSolk83mmxKYWnVqOHw5jNonS5XD/eIn+svHGF9gJ4RnOQeQA68VO+jgLY6N0KXdvEuWt
w5LqK6gJq7g+dG0mf4vHz8V0dOnaf/N84PWPLlVrXUg1TjwakYG7sczOBIeWTy0YCHw6/f7f6NT1
nSEJyNV95uGaqzUF1KrX7kCcLB+UNqXIoHqSlpEqmokylemMz9efmmKVlzRjNAOAT/wVgZyQ24XZ
ye0lF+Wc3NjRY6cvXq+DfjsDtJOXsxhtCfYSX98ow3NKvF6h/N8SoqC7n7g9jdHlltc+cVLZCS3e
fuBj+sxH0cbXbjrHpBdn9qOUDEZzQcvzojT/geOkvQW9ZzdNx7l85kpDgnxSNnJ1N2y9YX9ynlGb
vXcsWglfBr2HXC1nhfB/4GWHvfdlETf4zshuur3NN1s1xVkosn9Ul0E0dB7Gh7kv/JQaR8U8xZHL
ldGTBNmej/A+SQPLz2EACOtwzFPZI8R3dl8MbemD8+Qvs2QVEQT+cdVcLARkGtoj28/DVKbqEaYh
nCvJIViHE+GlhZNewFlAXS9259eOVTkwuJulvcvCWgrrT49RLJugy37joiTWxv3S+Lj+MR8HNpUh
4bQm6tseCRtPT8G+WFNtosxPScTbupSLJgwOuBGgEPNvob0gjTdDFhtux9/fCvdf4txS5nUlu9ue
Oj+bm0gPGOaHLtMOrYBCJWGKWAMpMYY58rbyWTtAZyuHRP+fmCLRV6s+orUR7wdFgH1J5O9mhWlA
YWVkbOgfhNSmVApAWluJ+wmmIdW/n7xNgkNcK3dBRXNQyago3PElj8ff28qOTnKV//PWwRveJGnI
BTHVsLARkU0AzPOdYInUslm+wpEXe3bzaybTb+R2eTtt7eFZ902aI1eg4E0jYvGrjdE+s5zqjFJA
Xw49E9fSy0l1DKmbqTmgNm035enREMfubhPsrZ7ay8bbyFTwtbBuc3XqNpL+nG5Hk4e3q7YwxXB6
ZThbAHp1psXDCa9aDirj+VNHkU3S8okhBUFAgx0SYxRK8ad+4nFCX30U9X4gxlO8KNkLpdD1LDFC
lmtJy4U6WrF4Z/nox/XxF5Ab07yOs+fywGuVoE43KFEMh0ydh9Fl+fZGeSDQ7LKV5ij9ocRSSA1s
otVsqe7CGcpEBWV2k5Kj+TExLEZiwPj3thx4o3wKmwAsxqn7dZhb4UtIo5D6JssdHJGF5A0K2oC9
OXzw4qlhy6zKZhZMQFlA/o4vYwiACEKi9TSH/11fmg53RIwDyaKaLlFQ+Mq9mp+5D1loJlN5PW3Q
daAhuXHhw3euzmrmdANj53ShMt0VNsnHQJ8i8uCY+DRDDg1C2N9MDHlqZm1kCr/OupRCGiiY1u+C
AnPNizPaxF1LT51vfcJnBOs3Wsu7QwkSQ9R+eRoAkjG3agxB+aVWb9o5U70SlfqZJDQ3JZbMBQjZ
jsHO96KNQBbNVciuH+BZZ1CEZ5jMuLlU/3CsBnV0AnHsG1vnXd9FY9Lu0A6BL9Glb96+/gtW7Lj8
BLg+tnQavjFkDJx+uwIVAICP2xmNu68UoJSL2wQks/bmyetSjclbjST1REQgYssFzdnJPmkERH+A
bAgp0I8vie3DflIkB1+lGh9nh4x5XzTLR/97Ph9ezrtlxW/Ee3sz0gFJiqqHsfTXCfvKmhVORfyr
ADYjnvJf66YzcCEZtB9HegdymhXYZCEpZYFtB3/Ia8B93gxfXmtENoX+IYd2Bx10XKnCexA6B5NA
6W1uu2nq8UxkjTNCeij9d9rOW9tYNZhTA3gWuliSmvD96g3J9CWUfzXuQBWHOU0cMtLlt11daJcz
r7FmilXhYOy453ves8KFdAXOruyJLm2hytuHgj4RHRyHrrXxXC9n0cabqmJPyBhp9vgCJbf0ix7a
X0l4S3nbkpRkmUA2YD1tUXW6lWQFBmOzvhWaj5CowB/7QNWvSoIi6wz14m/eDsM6HlygMwlND3qR
6S6HyuXrbdKDjy0d2L3sJHCep1+JE4eX26I0khwynXJZLjDTFpzFH7TPZubN9GMkxVMkgGbHlRdA
hflaXckTziFCTU3w09PQ3Kzw67aCRtLVA6UhULxa85/9jnhCs8wduoxFXLRlvVAuDjx0KAjA1pCh
PXoO1b38PnZkdD5Q/GVr3pAYTVmdr++cR6BpTtFykK4LwfJ72bfHStdYN4TxFYjexG8DQ2qhcKWL
hM067iclIGJFxe6pBFBHfO+PvprhIZWdO+6YLwuKoG3LAy2LB10WF5vjoJIaQ76p/2BQMUhQd8d3
F8R4sZ9/0HaxqyFTBxGRTW5VSadF8ZV2QgwpRfNeagop1xirep21dL+TS81yGjisMNW9d/Sz5Oti
bS3gRj7BLOYOAn288Q6JhGFhcKBE3HOm6nTEIytRdtlHcZHN0+2GbonYYJ6r6V7cNGBRW/14HXIU
KnqJzOi/MXEw9XwvLFTZNc8kp/gRJATsS67cgwMFG8nqJS02XY8Akw2H/uKj5Xz8q9LE0vLVGTvn
acWGWloUqlMHfOtDTf0aAkRfKseXnGfa4Ked19env6nBNVQJycqQkaX09LtUKhnxX40rPid9xZKq
D/Lj5BJVz0OTZ1JrrvGEIP2eCf6X+wNEedMTQa34PUdAT/YdK6mlrX4lY8JSTlc+HwPwNvXEM/5K
LiAX4elT+8Q9ychPqmB69fDBDPRmpPcp6PbYu4Uj0+8Hp905g5qOhftkcUaU03zBuD8QbsqPNi74
Xm+5s9waJuAJ+zabGERzrtbMESKrLTHYIBv3hCC9LzOMs3bNlZ7CZvhYtpRt9m3LoVo2mBzI39b7
D2/UWWbxa6/mZvsMP2PvPVnWTcnQzhN5tn8VlwS8n9kgLZW9zCNh4T675PlLuqrh8a1QWmZcRCjm
J2ULRQ0niWbjVbJOws3+a35ZayCj1gHGy2ep5ZybiCOE2b/AMY3U/Uh9nKBGv3EozBz3iyXmeTeY
SDyc692+FugM0+k93wtjtlooN/B3F9tEcW5DjC46//ZV8v0mGWJcI64iK1WTiXB1XeKzGpbKgFr/
KOBVP0yeLpR7wU8+L2O+ESQG9TZ2EjKg4pSvF73MAtSMOWGwU3WVmGQeTM5dbOP7gYBSVdUXVCNM
aGiFg2O84DPG1etMIZfqlUX5/J8w+LPACGuFOq8SeKZL4R+ni8grShofSFiFGFIPIRjGtNIYDDZ6
8AUZ+3yYCNwA6Nip/5OCylPbUsh1JsZ+r7rDZhMkvy6Q1VCS2phw2KRYp2llOCF9mph56AQ+oROP
HByR6aeYDiQlvrBOGJWRhfKpcSyKKPrxkEkKJB9Qoz45IqQ2psGfxLKNWuYnnDNO7aPUCBnhb/bg
7uEBdWsMnMUWKdOXZSSgqgMt0aBIlyyJL0c2PBne5FIU70Ow6PET28Fe780CnHvuY+3LgcxBsZ76
CvEdO59frV/5XJxr9k6mB3alvX1cX660tajJNrxNjmknIh38RHo6CklEk50DyE7wbeSZme1GZmii
qbM01rQSAbovOOBxl9HawSLgUprEwTAbfBmydwXSbkCzK2umXRPY1Hsz/K4OxAEcbjebfKGZqEa2
zsaJSn167l/Z5neKqruIEny4Bh6se7KDYLasGJ/Cx7RbBuwGi/9/jFoPV5hPQICkzzPAKMRxqJH8
5VIPruVzwUJIvRnGbFVR1U4O2AsJ8LvNU3HZj8idH00UODIww8y0Lpb32ayzpHezGfEIFf7DxJvD
SnCOoL0VdR/11OCZ4LIbG1gCjnXw+estmd8U+9Yi3bG84h4dVth67n2LfAtFK8x/fohXi0qR8Hso
6PbZ/R5Y6fCWfw/gyjYupKUbxYgn0p1vCxpcAEkUYW0awyP7uZx0BXANPMbmAts95mKSPoiz0EbH
RhQclxwoKN7pLHgBNdU2xdZRw1ioukIDY5ow34m0r66UkDaC0SZloO5aS6DWuby/CTH5lgUB8lMn
1MDGbzaY9vUx5JDvlgwlo1GTRaYwpywV39hYonIKHnPo1EIqbGSA/EHen/KliOP6r4mphujHKNoy
5T5bGRq7Ulh8B//ZgDMZ6xG6nHHgwL/ji0nAS0u6wB3zGpoiUVu4rywEjznhZlp7V8c8dDtRcCP5
7gYAZW2Mgy3sHKIl0SzkMLX44+o29S449LTO2WswF8LDxeWJqZuGriusB2mPvqnjJiNv7bvxphzf
NvQk5cJ+9CKEYDbCOqo3Xj18DJbeDio0s2Eu8ADsmMAbrEWHgVmmmdI89KEyZPTqwN112vslaCCL
dN+WDFDWXdSFQu6aFSIyn/nUyE5y9Sh9EvGJ1TbvRY3MgTSL1qclYPK3KbJ3HAZVoHiK6Peaws55
BApItPJlV846Y65ZIfr5XM3lb6dRq4TJzj2CRjlExuHlJSP/y4odrb4wC+/JbOgQTy6Hj9uQHAm4
TjVMRVI5t3GTWkbEx2QuOP3oewx2/F6xdWmnh7+Biqw/gAAtJZAQFaWM+g0YZLHIQCE6h6b2bdvX
9OAvyt8ww5MAaCgHJdcdfFyJHhhWFGzZlpMactccnPYhfDuC5YHj29vzlv2+fkaN/GDpdE/UY3E+
X8EsGRU6qSPStY8wbxoe5QJNrMk/E+GDOswDWI9lr6m/qG2ZdnqNpH7bCxnkYn8cS4ocCoMceJto
BfJIV0XJe6Ckk/8kKxzH9+stoV0x89dKLHqBmNpSFua609Jr1SBC7q6/EEM5PhkPzQG5LX4M4hZt
N9Aq84+Ica5EjLunddmLJ+UtyczjeqU0UGFg7573qavlj3W/CaexO9cYBfj7ODpMdCka1mb7NHzo
eQo4Foq9jHeZ/wB3pU9Kat1e1/vKkhmX5w/bxEAXY4pAXltLhqaPuSQuF+I94JOp/IWf29dr6qbn
lCeKXcdZNHt+3HJsejmdg34y+gPVZim5pujqJOrlFj/PtutQJuaTcxaJ1LwZ+W59Si1CuNYGn39v
YfDkXtKGxjnpM4RkLnHoiP91+87qFDe3A1hiuUZDsT5TI5K7vu94csaG1Dz7ipAHqKBRBgEU8+om
wuulzSTeI0UPSEQadnXpB0HIVTjnRFIsU0+XNoxlcENHDFa1e76kD8c74TAMsmSxopy1TgLbnOgK
fN4H8vTTfrIOxqAWIGWs841Hlauptm+NbGGvH/KNBGcRjdCyMEonw+t0ej994QoYRtfUIVvn68DM
eSLYRb+BeiYWHOQ+zriK7oVNObuCs/xOWPDN4fWYO229A3GAFagLhAydW8sKPEGr/pFtJJGCUT24
SaAs0Je798DKipi1M2aBKXOKtguYPasKSX0xopKRDfrg7NFF/epC1t0ArZ9N8NPEZIbV8fEgSJP9
fPvGIzL0D7IjeJnSv8eFX0HKbdZWRBEaGS2Z6dyukMng6oDZVWx1AAkXenFFSP09Qg6Dyxw5vl9Y
iBI9+g6j7eUdKh10PD+h8vLFxZV0CcDSGI08yymkHxJ9BNfrDOV0/UUx5RDlRE7Ui6cOU8oLXRkq
4AMzw+jsLMsH5K7j7zsTJGxyXv1s4tGcffDWX5sy+noOyKI6bNk6ygQPZJ8ihlkkBWE2LhQumERr
XUlPaDbDhVKIY6JgucY+faY62Jv83bL8fewUmYV1uVMtCJqxuxTpbSu5qaw8zrAl/23EE7N7a0jM
zYANsbk5qxAijuLaM6ZmLzAUX6jxHp6qQYGzMmZ5S3SSHbFv8mOwwLdvX6DtfoINN2at2+96ydpn
5dyUJWPAiVvSaop6brY5IuWdNpTVEcXKexnxwaPytWbZBIZq2t1ZaPY0d4xD+guDkgR5pW2uRtVi
qIimO53kA76Ut7y3zYk6HsN6wSXvU7Rc0Sxz6H7YBRcszG6HyP3M74Ywh8IwEzV3vqirbo/YfUr7
50OSz6zL2PhbG7CUR+oj4XvZjlEKn5ztecRCiKRR37ggsLYnroNpPSOoLgyiYWc5WuyAmWmTQFv+
tVZdFpB1qsoeQ5ssonBiOSi16THz3XqqzcVVrXTAK/dmggZ2KUhywdYHpXd6COAIewnCR00kfmYq
2kxHzReQ4/o01WEHHhS+eW7MdvHrWLAQ1sJ0uQ6uf+vm5deqGbraH/pvJzy/iah063WXaYYzDuwS
005rFLzcEdzb7eMlVEN1YbsQCqsEAGpNfF6jbQZAKuDmwzVZ/lNUlRE3SMPruCR5Hy2sVBCSW4DB
xcHJm2/ENJaZqubnn5m41rPpKSRlMiK5eNFx44f/56JXo+fFy3acOlHbBJuWheTlr3PgSMY2FAsA
Dh8puF4o87Ljw3Z7PJFdKpK8BDyccvnIztzOkGgJXJ4d1SG3jKTnpYuEyyqvlDwl8gqVSB1KSFQn
3P1w7EhjFJ8rZSru5/NsObui/31DYfwE87gERmlJuhGvQrixyGD/j6rZTiVCD1um0wTqDIUdPja/
kh11yUVTMQ97YYqZqF0FyMFRuBghY1JvmtaDD+r3FJceJL+WVsZl4aE5lq8SMROtHw15Ma2py2Z8
OjANrqGaML0bFrX6nnarFl6rtmhhWmK7nfaBCK2dWyNHESiZnQW55D1abSckqXSJJXppYncpOJCF
XiSl6nI/rmAJizoSCFD+bdFRvBqaUmes6RGTEOq66U7aDJr1bEywtVYyUAZhmuTPS6buBWQHzvj1
IEwpNWTV0NU/Aq64QpJbfXypCQFjF1oTKHHlbz+BD860H93OpGf1d1GWPFm5Mp7usu2B05kT1tou
za87C3uNliVwBu/DldeT1UkZaRtqqczIrUH8iG2qbVMkSFDTkXwX88/QskU4YPufSOoIcL/Z0ujD
SjjyF4T/8lMQNNlM5Igxv9RQBSUEG22s9h8Pyhq2gecEBBMUJHWv1cOeF8JKMdYTRqC6FEaVpylJ
frmELN2ESShX4+5tRXMSQKTyCTAos4IcG6WO8f6oclq4Vh6cTF1SfdX3rWpOKsZGtUyNF7YhSMzq
ODuySfzK1KbgvCxcZ3SUpeflbJIH+pkzU3Xtnjz7MXU+ngwaRvOcZBIc0cv7j/s14/aEbJg92AJT
eaVsmKbpOijTjXi7ouuse76WCfP/qvNSq0NOLwMEmN7uOOJ/JxTvMk0l81BEH3tybZX4iePnoohw
NDMWmy66rxo1X0BLGxK3jF6BwsG8f9e3zxulcfNADBTQuLPFG9OybbGibaUJlHQIDJqkCF8yA6Q6
5VG+DRMx9WSf8j7ZGPo9JkjmtAcM2KZzxbsbHzKwShAvxDgvPnseQj+eaodVXZXzEKliQ2QUqiCR
5BCTqJzYjYDfZrQPqZvJuoT0xH1rHYb+j5JkmN3SweMGwgkN82LedsJ+whPgvxs4wAPeLwX34RQW
fXfYA2oKBcCrnRdfkbQaCxDseU3MhI93nzsCOQYKwbhdCL17pNHcbrrzynlJFxT5ILPl943MntgM
CqAR0u8Vvclb/OxE+8tn5mP+JTw6SfTxswzqLV7UiVQNijcK2LK1QBfwV3YvBmmZpsauOtgvJgVe
v2BYoUFS2btdvmpliJ5uX1oPBUx0vffFJW5mhUi+uKjJFBSCX5uWITAKNX5693a8I9BTUFy3YkU6
hY8oDwa+8M2ORr+v/4a3RYHKfBsv6KJKgsazQtuP86+QWZoSswP3fNgsZkYVhpMv7c1imj5YjN6H
pI3TDVFg7L1uca6XAmGZbVPKxpyIjiaYN0nPQqDvPzYXP+BibJ+1ouJYPYQqfflYk6iXVRm/cFJ5
YokZpp6Qb4GDPf0M/gJwsOES+nXjEQJCiw/ITOvmEhsbMPjieFbAlhB9KvXokSeVoJwA7ca3WaCb
YrwNUUNC3K3vVB4rmBl0djW1IvaJzaTDc5DaTMuMQgxP0CqBY91n598S/htnQBReFsbVkQCYfwi3
+qbY91TzLLn7RUIZmDN2Bp6k7t6LpxrF5bKiYmckT8rlDnx9l+U69x2hDprX/UPZ9kea5PyPQocJ
V0Rzd7gpoU+Qd3nX3HANyXNaUIntzrRRw/KXfgJZu/FMSsrMeGLYlfw7hYI6mnmHgkEM8RWk5z/W
u95hZAD3jxD8j6DikU4TBveGbb7H4rlCSYwZCvkckkhQg8OoPAWPmOt0GNV8ySVSAZql7ywlxsY3
S2AOlhty58lDr6vrnM2snG0nOs51MMm7i/GVt9EgghW12+v1hrIxccPOSsRJplG4xxhuSd2mGNZW
s/ZxB+9qw5K2QoTk5CqGKXzttzd5JdV3Rdvy3yznnFp8RP0Rg6KYMD0hAWnPGBxeYTVbY4plLOda
DzMPnDXzo7eDwGQ6CgO9ZUeLa1p6pvFNHGggHmtpb1y40dKiqYhBi31WUZdpA51Eu1oWK5Ttbpmz
2xA+9rqL51wwdQElQwZHPSgaYmEYxiHJKTiBfr8tOBEyAjTzjDzFMnNXjBP6gCsvqn8Bl8f5QCIU
vxMLraSqmNZHR/OU7K3X0ZRGtfq/Rm1IJ7C5HG0PBymI6BfahCLjcehi6M/v15bixkBDQUqF5DOJ
62MU3Kdn7JgOuswgtJinv9YTZVixEn60BrKWvRFybNjfagkrppPiiuXadRZ20DqmyS8Vu0uU+DM+
p2GLJPXRS7nlaleW3ZgeO/ZNpQ8F3sDlWjhp4PjQTMWtlvyEdbZsh7SclqlMIIEdbTH6L+MLwOeS
PuOoaNfC+/bIbCpy9iNTBV+7Ka14DvzHKVPxncy69NztzUw7XIT+K/vzT0I1DfEIgedh1ZLih5DD
NhxgEINk/v7KiIZm4f6TrqeDfEmxmVa8QOftcEGFj4ZsCpii8bgDhKomTuXayyfrEU81j0F5hoTC
/pQFiXpG8P7V4bABO+gdH+H1mfOZxvyw6ghS1NcdOTBzoAAbsmS4tmhmMyHAivH/Zj04xQyN7Vzl
ES9nvKQTAH6S6xDspPrkUtW/jvZH9hxf1PmBVFKWnpX40qq6T9F9B+6IMNiJpkyBi8c3igy0t4zl
sMANxAye6vvJLKIkZ4XGZbBIkRlPwC42aMdftU112GPzLmrHCyzRebhkLkeLTgDzTDobFAjfQp16
nPJRh/x9FDBIjMpvusNghUSiLIUBmwl/Bcskj0DCigxAG2oSC/qwyDje4oNm47r0v+rNJkXwPnqE
Z+32MevhEHFt1HMaftgHUiQ2L1+SB6mK9U5PkyHZsaDQwJ9fkLZuNvWhZ01o6KB01iE/WY7sX7M1
v7GVLRCOIX1xCTtPW7JRDeAg5ODbJTnVExQRwz3V2UF+XlsFkgmA0l0GR+04898phx6gnUno+/Tg
F4qoEK7YGyMnj18HW5T/j5sT18ee3P4m77g5mGL90E9WhUYc2dJ+yuueFuuUGwgNWYTWwm44w3H6
y5Q2Hc4fA0PDfMuC2VpTDkETvOGWDtBFPWpyyhy1NhNSZacGNRVv+cZPnmxNY3fPTuYmlcNFLuhq
OMFavPdzv8gsJOEwrsodbKqyDkF109ICNeuPs4sTyGzGEWhw6NyP0Krt2VQt4kOQYea1TsQ0Ck93
5bFz2cyDhx+b48WJ84R1k0iSD1n/6fQihtNXm8fkHHpceibNmfHDXlhgegxOr/V7CWwpuf0XpRRn
96ohFuJcNSMnraCamAWdUmmbbEDJDe2h14Pn6ubLNXrudPT4yot6u986ZcLyy3KwUGrdMH/t1Nqa
/bNbUJ5IBycONPqT8QOgnpkPESlEg3/66UOa6aNE1u79Gl4s9uY4k+XWs6m+hfKXSpVF2yK4LjuI
QEYkk+KQyNqgfSAdh8zqxYYJpFxtNn+5z4wa/ZnlPatunpmXCSnaGu41Pd3k7xzIfSDL2ubVZti1
oAPGQhOlMT/BtDzDeCEkwuWlGV9zklocys96Tqj0Y/ycBNJvuQJqVwaZIVhQakbLlDAUBbsXNEXR
+7zDtoOCdoIRhJGLaOnMdwxS5mO2dK74n93K9Wxy3Bdy0u1/2Yb5UPXQOHMig13UVHUAEtx5Xkek
i4EpbilParV8XjTGn3fSCfzMjfTgeJd4fAfya1B9Riw1hd1335q8nkWufgADHRr9wZWXmzd4C3oB
GnOhIleS+VYgDFEdAjwLgxD+vjVXhhVbbZCTyh/NOTeDSBwx58epSFBbaiBIpKz+RxR4/hhkNYsH
3ZwnCa8EGOqztbCRxr/7AjgTl5uJzfkP9OcWy7dc9VkozmTQ67EBycLkRCT6xmO4zgyfnOHuTKe5
ximIrWeK+z/9wfjs4VjUnxkQOp1ZM9Set0YT6lsAYI2xqGuc0biTz2Em+J4Dht6BPlecyBZY6QEC
d5g1B3PjD50SI2U2AS04BNH7kndDcbMdYNBl4f1TcrBUk531NBuLlgkJ+HlN4xN9gmnvG4GicCTs
F/g6fvuW+TvypL1QSXHzcc2IueHg0QBJ2H+8n0wl9ZJUqB6bCHuA/hKcZdf2fPuRRGGKo9wyE+DB
MoYzIluAqwsTc0VCOghUGghLtdvVuV5U8bEn41rtPAJLHOQ6a+6Yz3+KItdqO7rfPZrCKDCsIEFt
7fyHM57udS0JkSSazz3dugHoq3VkfRtU2VkohwWuVLnIww2Y9P81lXciiADjYu0wJP8ULp93TT2p
LWFipDAxB29wccOG4Loj3g3leumD/9nYvwy4UhQhWlFCImucLvfrSfv1iHB7WUg/85RN8DohUB9T
T2HBabFwFLl/Bl2flswUCkHQSYmapR6y93xY69XpVipL1uD4cPaEwCFyKcG6iax4sKqs55SLNTFY
SEjMFbWHTSjIjEy+wwrDnCoYqedbgvK8wzygq+tWvseg4Mfmwef4mVklP+7nJpHc86mS/bYHB035
+sajlyYCVeBvW8euigf9eC5Tyo8QHG3nkXnQi33Kk6vdMMEHqMhH3jOvJM6x6jRzyIT+6KW4pll2
kFonJNeG1Y7boPmtc5JlwWWkDsvxjCeVVMHLiEN/mxKEJvDS/QI1IRKSTj5UZT/8xS0UKVuGL8bn
dYxcWcn+r9kPpRxibfPL11/+x7PgeDRIAc8CbG14V09mEEyLi/DnoBv1wWxIFyfrxDbK2dAsk2W1
tIgGAlyfNSAArmCNPq83DMjkujtOgFA2DERYO1G5hdhDJQJFjO4LftbhoNIpGXSv0nV5lVgZ/w1p
vwTwrIsmSlkC4ZFnynMGLgsv69R7KxI6P7O127snML5kUA1RECbCFLlkIdVwpr1L2e/dCG8w9D4C
a+TNzx53oYvil5ZaHaf3tlWP8tSnxGpJv/BrtcJyWUKGIh3CqnKkqI4yTCZNN+NsQK4cdaLTDtp2
RlVY9uGhWlrptz/pfwrn2fo4owB1FNf/JNipAc04G0xcmhZAQfM6Mi3tLdStJri3+Gd2Qzk/Gn+b
i81vwEfuDfAdAlXlCn9EV8LmOnoTH3myc7qSstcvWE8xXZbFqtFUuf4r+cNcyTrG8bjAsuyoQyaJ
rA+AGrYSb8Oc0CqbYWtLix12/TtvZkBaeG8pBSl76xeRcg5V5dMb3sPK12uuk/x6DA6IC86lD1T7
V94QMg664v0XFBSWq4Sy0gJJpFvFzaUywyYshUGgQeC1mTlOevALSqRNpAwuZ6priYhUYaVIZG1b
O51Lnuo91mT0qgPMj+BZkR52MUJekEtMFjlA8obi8ZkIPWul8Ruqp4VDNr/4c325d8AgVGyUyMy6
eMGtxVTEKGdb4pcY/nQlNEHv7T2u+/x2AA4lPBLYp7hcE9O0PLwYM2gb5M1gdyZ6qhAsJf/K/2B7
i3zGBkNhJ5VMab6skvB1k+ZY0fhF7atcLsBpgmt1c84qRT0lEM7mkq5wWng/R7TFpDGsSOngcXjl
JEcyyRSwcGpRqqH9Lw/Unz2F8H8ace1VJz90G9WInetOy88Pik5s6YpQB6FYtB4SQK/R3aWkArp0
VqRrHG+GgiDPFGyZkicSFSBuktxAAHWen7N0WiJHlCPaI3mcA/UD0aMZ9LafFCiQ5rn6e6Uhc8i0
Ezimbf1axO6qxYRess5ScMzUgPwuA1f9++po4ar6bIgw7hBg3zHb3iQiY6DeLGMeBpGKg5bewlVP
TuUrTc1qYADRoyLZbMDlKtOto5LysxiTCvi63N/23OEsYS4nokjsan2Ey+7u3whnmIa7FgvpmkTn
pqYRz06YuO08v80hOadPE7jAnL8xsV7CVJA2Ujs+KuAmTatngzi6OIomic31t8Jv34FJsrlNG026
WH5cxTIB6EBonAGC+zY+TgMfwsZB90Klk983aTgM+iZ4DVNDmwJ7fxRQ4UdcKTM2q6zBEyzq7gK3
I2zKmS//+ndEonsXaWcBISVKPNajhAm54q5iAq7XlEi6FcEU83nAucV2eq+DvOFtQWPDSIWnJMJo
q9FGqAgAPKulM8sZGzZBM+FJoLzyCKv/Z28Pqb/7MRJPPztahHpCS8XNvUbiZcjmSpqyjieDsClp
fql2E8LXQ+ZqtiKch/JX4hGF4VzNOMcNhWC85cg+tM3mEZlR5VRGl+uno8xuDH20pX4lG2gSifM8
4RjixNCThKs2J8A/sYA9EazfeSvrnP+hz7MoMwDi9fxFJgxEr3KEf+bM+bf3ls4uFgMr59Dnw0O+
NHAurjg7d47Igi94B7Fjgt7htnh8gLq4+TkILJ9POeVTYLlv6BtUhUn6gUP5Um/k5kdZ7IjCeteJ
BFuhJ6TwxJEnUtjVXMIO9+M19vWqZ9zM5LuwKlxvs2v+DuLWmftVXRMk9PT4NLrJ3opaBDgaNCai
Gd3ZRlkB92JBSzSayzYlA25b6v8pDZ+KCKOmkEae2wmUV23+ZPVsiiawZ2K5Dy9dB8MSG6ZK4Wp6
Ys/nCy9oxvMkvkZuHe6VewfK57A/vcin5WvJwfraJA9CQxKv8AHHmHMiFY5o+QN3OgveIGkGU+p6
28w9jo5wIxLB7yOrziRDjxUeHuZlZY8es1VfwLqevBWjegkeRObUE16C3OYnZR1SBXmNZgyLyPne
EpSGDNcFFZlWlpQ9yuaSSGMzshTaQBBIpStOFPCy5QZ1auFtUcIsx7JDlph2eo363SqUexwaOcJT
cQb+wWqPycq6AXwqzlEK01T4RSJuqXlr98mZ+E+BtxaZkuv6oGscZHD1GwdYqqODAN4AgkPRF7Gc
6gsJkgoIlQxQCLq+22eEmhQXemikYcEOfpHuQ3tlnyPVOq+N+kalTrVoqB3ad4qQ1PesGPYWBsHE
KC57Ja6/FisTefpFZ8oPTZ2hVVTZhAWehthn/UunlX7HO752F4Vb6nGKndRdyLJTIouqu7uM7IQz
fowA2x751Gbu2JzrB5DcRBvp0m/uQD22YF24YuoxdkGEjoaBxFV4wBtFRLg6xkba0PEA4plLMtCK
ksau5mxtPv6vV7eNXVFWMyZBJ+qXNylqmV1qerLw12CW5Wtpd1nxN3m0hrKju1I1MFqma1PJJRXi
IrHVr9KnpQ3xQsPwM0Ovm7gDLUxK+os6Eeg/pfctiwrPf8TCw4TV6bKx2B8XXlG/vvlpTcmZkojg
GnW0NFWUx+7x3R/fCipsOPbcf65GiQDSvZJ10ZzUpdnCUoTuEGZGyC7L87SQrG9/iTmCHrHyAjXX
rPayXHbLl6KaC+ULM1cm3ID8EOq7Smube5tmakLmt6DXzqRxXxbZaHbqNTDXxxxLPEHi6KijCD3F
TGZ8fZbDbaP8QVDen3+bszKOFeG924nbJwfiFBpIzE/oyHOHSwKBijiQroOBA/XHUA5aiDRCXHUI
DUfQC3VHh8LPfzstXethXjoAHkZvdFSF/JEigFp8l8QvI5f311InDTIVX7IoHDiYpprbXSW6uNhM
zW9BbqSmXyGfy+GIQ/ddPvQra6U5aK4FQVbe6Ly5Kmjq8kv2eYnT9eIiWKXpR2h0t7LQPZR+ynzi
ylxaEuHU3ZRs2Di3NF358FjhmdDWtSJBblS8VoEqf6xILOswi7fq1FHc68eS7GXjFkpWTydfdoZP
N1sqQo/XekeO+oL6+kONVfy7cdrKgJ5yg13HMtgIT2dQ6yzbJgdSOF56O4kpaR/JZ9V1GFpC4B8+
cHGjMhC6cdI2ZN21MqvzE75DibnelkOFhzpLz5C6s9KQJ+lR0r4Iplpef87r+U6xHGNlhwjb997Y
wsM9lO9cg8xvbk0i7Er2zNyPtHfFx/i0N6sLm4nlaHghH8R52pCxS0/osA0NLNpEQaK3KQRgCGLl
DwwZBsR/2m43lF/c2RFIrliT0kpP2sFZv9idYEduOCPFCpnPYRNJjCX90QCp/xwqhM+ImuJ9x+Fe
CRQH2pRdOlguF+9IQ/S7WUh/GkP9VLLArIuoGSSWmz+RDmYCTS8W6CqYiWCJceSaOoeL/hZ6P7Zo
nlgdT5ebpn+Lua7Xd78uHbJxJhm6bR5JxuBlPvyB8HX4wvcOEVhcLcu/+eYfbX7cwaPZF03ggGeJ
jBoShTnyx1PaCIdWkuo1zFxQVZ/oo4Rq3dibdtiA5OLa4BJFKwyAOsj2BuBspn2Uq12c5AwFgtQc
JqPs1JmB/XzYT+Hc+dWrSGxQjmFkTQDu3Aw2sGDfMCLQ7DAXpud7w9USuyq8dSQYWWNb6b88PI9o
NK3qgIhFJu3ShKqBbQFVONinOCr/j44IPIaDjqwI8TwcRZVnUmrRFXx28vkHloYqs20TaGICqff2
z/TubUUr8UlJ/pjeCP76ANuUeN2V2VdV8sqB88lumwpGhyOIWx0gwWbRazKkFn4F7B+O7YiV2p6F
CMiNnwJT04dFzDXoMCwyo9flQYRZ+OdpsV2CDNd1VeudlJ0X+jYHY2nGdUKsZpOW+0jB4jzDHKDH
yImn2fqQf4ATuSx7bqzfeq2fBf9ySE+lX+MliEfQEbdSRgz3I9TQbqXf29fPpKoRVA0tiOR5YrNw
U5p+/U4ApQqOqIYFykWE46ERl8Ux/ALPdWTnsUP6J24TDAYRWUwJ7kkIyAw9nPJpEBbWEP9Zpdpp
x3q9JOBMIF/jRgT+9jlSc76RvvPukjXaa1frXowyX2daFr4BBIcvm+t6qboEP3ZqhRCyKLe9N4yw
DDF1EfUGq4Ej6JFHprZZbdsyWndZlwAibIFhCVpeSo2IzZYwgLioy6gaPcl/w+Rjr5yoQE1vC9dU
dHhIghPFC3dj+zRpw6prqQpK4FSNBjWmjdzr4RtOvJdJiuHyKBLklJNB+TLfPEqC0Ps5/mM0007o
3OIvLurS8NZebBO2tyw603nsc0CCZxXz3YMD+FZOim/fi30XjrSzTTsp39KshFMhU+hNkHzrP011
NUl8yyZn22QHFtN8POAeVxcj4MR3H2MvMS+G2n0JKRLXPyBW5HT1sR33P0buUrwa0A4XVQYGeB0Y
qBqkF1ixASOEHelN5bQyTrZD4GpJky0CSc15kI2F+GeoFaERIDIX5KXgOO0ibP46fEGJxVEyZM03
MQuf+TWGGnVjAQohg5qpdm5qCc+DcFFBivaiz/7ntyEmi54JR/Sy3W6u5wPFnlbIuA69Z3J04UmX
rr/CKbndq4VHWDX/O/c5qqT61lUGJAuPZg+QY9131/wBiYtwPlBqMdMuKlYkTPsLhEbfhI9mL0fb
/lHRjIeOFzg0Zh1NNkODW7U2q7GaI6eB06QGgNbWU5QbPRO6wMhAcukZRFfzRrWTWbp7nCLkm8Vu
zacfSzTFrrJr+b6PpnH9GrwP4EPIQYKzckEjSuD3ouwux6L9G7coXMDuWM3QNoiHE4czqqWSRjFv
StHRWo5/bjcmYtUXbQDc/1CbUwgM60SJ16bLuKWZan0FfmgQSPad5LWMw5UTYSa5m7GysWH/kZeY
VsLdLiFqQajB1H7nIJnTZX0vu+actLSEYNAIGfxviFNb/yEwljn/KCJ0StsukZ+8+hvUwmH8jDlY
SIz6UDqLSZZ9YlqSKrJvCenItJQXB16VIBVvLh/AHsGpZjmlu9NEHH2mb9k/tsvxByOpATWNJLCu
MQsxyxPMPDozlxc7D9SXsa1Mh8Y+GzoO9UEo5FBkbFu0ZXZ56Gw3V0bbaKJ30731U7ahH7gre8dV
lPCGC4I8HpgXNV+mEoMYrDiF1WVuSpFzC285bVt24laYyXwbILfWPPlsWfgtIIvRrJALMZHlhWKA
UwTu1DQQ//W0FajahgcjW9Bd/TOMjVcPzoSMktpdJprR/48LNB+7ajN/ARwA1BmVycBdJ6rOneCE
nmWi9BLIom9LoOkRAlqKvs+8OfmcBkpR1Y/06WiZTQ7YHURuRvdg4/Uz7AziQ9CYmuMuXqrFud5x
/I7WH/HAtMhjReIi3Nb03uaIH1iJ/kytqBuq25vciCOKZFpdeDCrPqi1LD9HCuSQIXW+yTIMY8as
P+HbCSVpFjelmgxWmffYYQbxrYSdt4SS3QrEMdNoSF8ymtE7CSeiOgdSo2UmZr6Jtw5EnT8eQDlv
1GdkqqLKU0ootSs2ZDWRSKd6IE6PEEvcMVmqrY8PsvrTy30MvV3h3+Uxtp3St5tTGGhmdgVytEXc
egdgKF0zJMjiR3ygyIV/v6/OVUoXP2jAJTabl0NCrSg/jhLNd8qht01Q8LbTsVajkgx5HqzRVbDU
D8sUFgDg4fmoBk4Bba+jcFavvSBKcs4sbjtxxvJNh7E/zHOBXupJXMESZgVzEZmO1+QEib28nZc+
arCzPPAMJX3rQVBF8oLNrFR5LiKehVJHAYSZ/9hkRgMYDf+s+pS/OoeYz11wZ7Yt3XNMF3zBij5W
4d5cYzlsJ4d2+IvxD6m0HQB9cz3LYX+o0QBv6gam6PSg50Yf/FfQT+BBSCyglePUnZsWqVYkiiBr
Ct0p3hWjnA7y6n2C5O9aRE0hAcPER7IrDZGS6RQZevPIXRiCLI9KFWvfEfxFLMYXUPA/R6WHxaW1
F1KUzRY9FmQxZ83k1Ui1pgxSZJJHnYWCSBHzzNcF4w43gn5dQaIERnru5ah1js8bGSwcrIr2DI3E
b/SR4sxrGZm03wBXXUErd+APXOUmUn0Oovew4aPcq/BqA21WodER5h62Fae6ZUbGM+lVu28IQ+XU
5aMIgdyb3UH6CHqxOP2/OmDIiWEiBJQnrjtGxzXCaIi7q81qmZzPvysCOmQr2vCfu1R+vqEXViKK
PA0uCRug9kO/8G3Godyi8Jy83VLHmY9wHpAvIcWJ0QEKkayC0kElqWMIyCoOqlPYxxs+BCnq9ZUc
kkM9YcUfc7lIl9hEhHmkIfrdYaWG1VLl2nGuaeltUmYxL58pVeMObGNt4p4tfPq3FVqrul/w+Jht
wPKYuk7cVKtYrK7uS+sQX9oYIoXY5sn7aRxIsbDQBtShoZPYTbUT1gqJABkeXfbAmj10Lzv8JgKu
B7PxrvT3ssVx1LgLK49SKS7I3S4M9fbiIXXQDBhx5pHLeeSviJxtdiCoXmE78/Tu1m0MsmlrQbvO
Nl5W34ieeEpCBxpF50Ew6RuZtZO3XGjs8gnODAOJVbAjWJGKOVIr7e9p95TVJQS89jWMwYXtTLnz
ka98SUnl3pT+eWNs/fQSyvxRCVsQIJqykyDHsVoG7g5bEVYG8VVicz+N0OBlzy4nc3fwEmIvZJq3
cTUD0cMza3LQ8c7WoYQenTs0y/1DhYVCARSgN5j+HWcpe+DDuXUSo6NsTjmZogxRbg1cb4tg2Q96
NkzXxpd1gwa+eLgaqecZkKnrbmQ/ESaNaCJA1JUuhdhhIIA0DlvlND1ja8gwSAEgwjQdDGrTnhVq
G2a4deTKQqNAfNPCyXQRQPGfVAvIDNSyIdpiL1s7fWbwJFMOQ1IEWF+tKsurmAbqKn9ZIwg3jRq+
iyiou59ZsYkf2dP8wMfC09pkvbHTcPiy3pXcIkS2ed5p7vhKe5utT+URWinIbQnpIAjh4ygx5rMn
NeRmCpW8ay1aXDFDGASXHGNda26uMx6b5f8HGFvEmkHwdDZPjfoT5DG3UOZDtZa2Ae9Jsk5e6s62
6HNesC9dG+1pXAtC4JJyQtbX8WH9I7SXQqS3hhj5lJMsNUJ/dxwQD2KPd6A8XRtJu1QxIjtZwgQA
ivmNo9+/Olg3ihsO7tTje6++w6n0fvdNKCopGFWc/ta724BAmf8WdL8xcldKIVII4SW7mBwgSArc
HEOML0kwlMm0w/x86VTI7YHwNG0UECRI+mn/yCWhNJuGhL8RMoPbXA3l1M9T1YtSsgwuxE8nVJxL
ucjhzBU4N86Kwc870j0y86ZCJlZbIDDx+KS/saBrJ6+Q7juxzSueilfi0ZKEMLrj1/QKmAeCB7+j
y4CiGg5Giguk+GATl3TB6m5s2R2p2GMWilvBbZMuzx3cZGjvBlYL7w4vgZXDfFIFVc1S/ED4WDM8
M8GLJTWEg//D/jGGd6guIIPcuH4oDuuFNdKpUgNDMcygpo1k2bHF8MtPAbA93yGsvs1OFU5yay5h
a5n8RQlxrKnw+iaDbQM243tl+6L4CM06DWUkPlJV/7iOSepnGDOF6R5HsE9UXD3g96HwDLR560/D
vwjFBYnwwOyoc8eWmjKQ36AEzX29Tn1th91SyP5ZsWn51I8EzsHsWxY+JQG8fI03Lwv+U1rTsvRz
C7l8v3lv4LNneI1g1AhFAAocKOb+eIQ/JWU2E1aYLM0q7z/aM04vhQrFY8Dow8w8Xfpavi3ehcf4
kUgUnJYMisEi6q1cGcXNs3BmcfZdNe+H4z+XhYW/hOFwN5gNp8oOrmgFeJKdVea9zszAbkRPN2ss
XviYxgo0Ibzv4PFFMNEDyW3ftRWQrr91m3MrXid0EhDNQ58jrRXt0JWnsbm3MMRF2b9tMX9wFrtI
oIo4JBgd3JY5EKC55WiQUlPqBQEseQZMbA+7OUFcY3V1PUOdGWWnx9ZdUDrSRmrv3iTpK+IMcwk4
0V+WlM0tTYDBu7Up5cC/ktA6CuhyuSb1F1ndNEs7eRucx5ykU7giBYAU+pz0cHZorTu9s9bJWZyj
u9aBxpyn1dEzD7OyahdJl7KeasdsUYF5AcordSutwm0twR0D9VF4tz/ZypvENBMXowZSkbHMwOsi
HOqncdhwWsCRn0Ze/+YpBMbIppc1n1fVlpo9vV7haRix5nEsJtURpqvdUdFXihqRRDIBHu5PIkLJ
WdFS0v0fC1jHMwFYw9Yr0zMlXNg4v3ngkUzVxClCzDCmVnQcNyyE1LTvwlDP4Tq2KQbusEDAsVeD
+Qc+vjOjSU2ByuOORUn1RxPwNEOmd0If+WOYZ19Wz9fMtF8+1V2VitrrUK+wGceH1sI8EDNsQFVv
nhs8uqNODtvpsF8/ocRL0upURuQhfwNb3+TyAZM1jFzKUrfnbftK/GLT0i9QkJUnlO5t4ZY6q+/R
0TraAT1Qr1+lPPkccrXJly++PJCppFan9cYOxWQ/o6apXpQdDy5hkgRfmDrMY4j0saGtd1YEPexK
NCEprcywmeAz7pHslIl0MJ7XtQDwQldvuMQecKb8T0AlU6cRkuDrWFTNBoK0Znqd0tXNfAY9Ym2M
oR1nTZ+FI2toggGArk/FfeleQnkfeKyxGqa/NcuFcZiGb6BjjcOH8+jEpO7EECdRYZoexXXtmvpU
AHQOLm7ka1SoECQWZKI5u5z1UXPtuIWCsab1tcIHqi48TKeAeTyAgGJr44AORmxN8QXN05pyE+ax
dG312lIDBeC3XXgWxcpXuFcPFd3MOUDXzkm+gZL678VlVGam+2C2sFuoi6ln7Ev2WeT7623/ZthP
RY8D4O1LDq9AH19+DuboBUeqJZLm9gTzxSlnLdldTdlkIAmEcE3J/6tJrWfR1sejrYWwYBGvS6aI
kGuln1YTmnXJmzWOP0yTZ5bdsWCtuN8UXNpmcQuTf3xQ7dW23k+KIvRiwK4kX6AogyfpT6AHI+4+
l40v9f0RmADY4T5HRlUFFteVEcVpW9EaJNpvmEexXAe8ArwS2dfBUZkl9IkurTvelA/r6sNM0Hr8
9j0OTPZ+SkxfLhqHzLrp01KOEOuratNu385s6NlnTeexz1wHF5S4vPpwzSpkSnkjxPbCOmCgzl/R
NWEg117TLZFbE8m+YTVFnNG5qlKiJvXN1qsLJ5azfR639VhKOrCNxuQj3A/ITzD7bUpcyj6P+MJo
R+P0A1grnDmYHvAcrgXF5LktU9WIduwcbTwfWyDcVrNJtBcaNyQlHMfme+Axibbwd3Z9XBWC+gOm
sen6Tk/mWCeGGY6hLuhg5YyaneGMvKZMNv522zCdhrfmDCRfngPEVNldhmhSwUbufpdir57tRyK7
01pN/wP7V/wmAS67fCJe87E/1LEQYBwAjh9BYZ3gXuDBWen0i2P6E5eNoXZ1wZcKk6p/XZzQHEex
hJfsLORlJsGj4TDjnncYBhIqXg/cKkAl83n6b01/utloieYtv1azxq+ed2HSiFQtZ9ITI3UtF7Xh
6idDeENmO5RFgOHvcsm1TRcrFGCbOY+StlTxmEbs3020NiMiuM+G/tZbj9C1OQLqY103oPDQe29Q
BkApUERI80Tn9JnoNZ7FBfj+9lRcRw/OSRT0RFar+m76d7yRG3pHR7pBG6FEiBMm6Qh44glalRWg
dgfOGblfEjO7v5Pt89FE9vRJb4g6FKVLAd6Tga8+FXlKUJEytPTWTsTkIuzjfJLArf85FCpxujF9
yNFgPve9chni+0QlUnRQylojaozAfV7dcEPNbUtRbfN3J7C5qywAcdLmIJfW8QR9wImTtM+h2O2v
oxqQnEOKgniJR1ud07iQp+9Rj2pxz2kIbISP7I+T8uhwYOGjCFJAm1SJzYUkJwtOaP0c8zRdSqrr
ci7zhXtCeIKVB3+30/SkVV5uxKvEX9LVVFpxdL4ZI4yNgfGKrX4uWk4wqGPo2Kghtj1mzgVzii6d
q3L8q/7mDMRx8W3o8UuRoxRQVWYuK41UExi6U2KQfzgfh3r4x9XA43NnaBbtu0Nmtq1BXq750xI6
IAUwWunt9gXRVMGBTsOPpFy0W81VBwB25QohdZd+/25ayUOuO7HMu0kbsM5xVKfR2UjMZd5fnwYW
u7MsqMfMF44sIZld71EDTKqssFa87HrLlAqaooGccc6dhtWKb4L6jQ+kI1YPmOgLiP5PZF+GtsGc
n8W7fwq6Ub/Xp5U7s+kykMWjZMv1CLQAFA+vzVxqRYiXE13OEqf9AM+tKStM/dnVSoW18/SZjYDB
+OsoZKkI2h5GPYokPR7andYg8f4VmMUuLIIz774S5KFEiFkD1pBJmUNIMog9PUdowA4XhZI70/GS
VTCJxCcoHi71b8AJFc/tqYY7newj0+LFLC61Rf5tJ0OUoVspJ8o/JkmZ3w+h83hTMItBhqg4kMvf
96uh7KjwaWQ3eX53h7+ULga0N7j3bHqG2NuRcWr+NADyS4Ye0i4oRiIqTcphHUj/dnKtz5GrAduS
rozTbWjIq8aDO2MxB25lemooHkRW/74y0SOL6peleJ1/tsUvsayqLfoWqEQaX/mwd9Om+bQme42J
8r4Xrr4VxRtHoxd/h3J9qg2+DyAgVtXffYv3WRo3+3YvePWKQMlmP4zDJm8/5hPQLRc2TkvULWl+
LZ3UmI4UiLIbg7ewyJJ4YZx/AF/gwdsHmViP6O7Qq9YHk1K8jX9XyF/ucOXrNwPl6SwySoZE4UM+
vOMGR+x1aQEhQTtWYH0hNhAL1DKGwlMjkYWpYiW7m20NCE5nhnNA6QTssyB3TuD9W0IDnaLBuMzj
Kf7pnX2dJRv59fhhNUIoyix+jAMmBOS0IWggHWIS2oJpDd8TxmwtrN2UHoaldX70xCo7YH+vMnHX
0eVBY3OXX0Hf0hPl1qBd7t1e7MgGD1i/uNdNb4sK4KoRHEKSoOf9JBXcCsbMsaVHkXX0nURWqGf8
v16cKYZzJ05IZYLOPx8SrQc0iyXuAIHRfvK6+VRLpvysVfiUw81KuynmLsdtyWR3MfcfLfj4fsb1
M/nS21Mr+HwfogPGLz1RJjcRgzTCj4ulXqfG96S0bdhat8tSJguEK+mdJFYSGf7sW1rKyFJmfHFT
xsFUfnXGTFAirEAquNlp7TvE7Krn4d4RQ/kmnCyQD6Gsa0okL3zCmyOCGmzNL80ZW6bRtVeVKWpA
+NbPpFoX4NqyvRi/LPft1TVF8AePnPQPL2Ky1OJ2KbZhf0JV1JLfWhjC8ltGLt/ERG7bquZRBA77
6zVYn7aPKxMvOWtzJS900eGIyb2RFDtdd2sqU7xpviZlkt8FsNJFeYjaCJnNBT2jt21Bv8AbPTcE
JFuJj4HoWOifX5RjljPHxG+jyRb3YWj4Xb7ImfcJct3hI9uL8tP94bvaw/L0puEBgqMG5c3QJlDt
cDCmealmc9+IlNJKwxlIaQfiOeuqma+6lo1oVyXalzxkITjqWqNiv5mu3Nrm7MhXXugKa543w2hz
CXF+q4AmyLCVljMEdsy8sY9SgiL78tnaPNPK55dbgWWNWOtlTtlEVsPfB3mwhLL5HtcUQ/NmCY9v
NNXnWXIOHb4pTplgeBtFanEGUFl/sRyla2E+3oGD4K9yNZyUiktKFprCBeTGhp3pL6JHsN+9TUjT
X/UnJrR3n1OscvNhVI02amNTiIXK7yPvKEoM97yXiG9v0MHGLPQVuulOopZzuKv/jWfRUqkwcnn1
AoBIc1IKv+A2tUlGOnm5u6HLc31ugGXgJwbdJHySqAuLBK/G5sGPsiVxRFw1W8gMamiRw8ZZABZm
TqEkNF4xcJl5ATrT+Z9quPHHqR6yP044CslpSUDVQDSty4CbRQ3L7b+b+9zEmwplLJMayi0sLNTP
lFx7lwbbQz0OMCI1wsvJOGXvUp8EYbjK/sWw+HxQR1loc8z0IPW5GemOOB9Xd/L+l5u3krYgw5OW
5Enp4fOXTBebSXX0prfxtLQTMbs38SRXynwUCxq1ujlyJFpts83kqK/9JX4FZpk68jOXxjIJDUmd
04oNIqfj8DClU5nGBYP884FtwTtEWXCR505Ns/cP2ipS9t0GUGfZ+0VHOqZOIf1t8DCeZ8pX10yl
839cRoTjqoDEuLcKtJ8uv+wfn/1ANvO7Dr0pxK1tSzEVXBx+ZDMxRNVFEDFRpplKXpbcnGjdLrVC
v28kOZV0clDAM/wT3fhVdkdSUK4lSRVxcy0k5crpNcZJqWk40F+75S5PUaJDJR4bj3grILvJPa3H
ix0/mbCm8hwsg+/9EIV72CvuiAOAyykVREfQj8cnc3csSEwc/QZYeP7jlJp96IxGCpzfno1MEgqj
0i3AE/TS5AvmbT1/5/+vmPnqNPbKgyiKBwBWgd/z5SHhwAzQ9zIcoK61+TJB5sSJQ9+vDPZ+w9Z3
n6S8Rfj0VfGgcnXZKR24Xd/aLD9i1tGmTeRDrf4dEP119dmC1lTxf7dnCe7pb292R2D8Oix7BT+l
UyFYrebwrcCpgZthWclBqiUHJS0NKg/xk5aJ4Xbny+IbxZPklsCtosXesErOh1eYuoFYf3GIrSO2
bWfJ+g486TOR9IEDXwTJSmzTvn4LlvfFsZmNRow6qURcnaqyQrMYvm7BcToNpgiGeh+WD3TdRmXj
qQPdF7N26/bC2o6MjxcoKRLoztz3v4FqcLwDIDfmv3grAm+Ml55zH41HWws1IhhXpSl+Vf18IVx9
HrZ0qDD4RbXKWJT0kOy3N6BHbjmMMjBpsHW3exLVLOrylOxski6OTzHKT0LIJyWYy1RGzLLl7LL0
t3YedDRqe8/x69vWMrWE9A0tuBDCeQe8FYq+UFp1ZZlhlFZvrfdJpNbZYvmJ5UNNn9RTBHYCSC1P
BVxKBH4wTasHmp6Mq8xYoxFctZqOZZF1U4ynKu0hd4+yD9SZRLUofmfNkOlQHYymRfflxUhu9xbJ
EQyLh6EstI4kIY6YAp1KuKY35HCF3AZITnxwncz3SEr1Y81SFsFlqqscKvZIJeo5HFfcXV2ZWsQ0
MQi6J9HiAW3uVOsuNd8imMRMFuO3pkSCFH0Biin2Kyco3urITEGubfQ72YrT1FODEAndE3UfxZ68
XUG7+yfiwi4Ge3S8kLVNFnK2FXMR6ktnyR2a4OWepLq4gEZPFqC+LiGuqid9TqTPM21cRPK1EBul
bWko4pHoYRtJe1nk+uctkg+rbUSwF20/3Jvu3HV8VdHSouiu4HAI7Wg0mlpDp12tmzY7VJn/Ry1t
ASV0UkLbMiGXWx2M8cv2+IrttZh2sN9UHnR42QwafmKunlUFxtMQM9PKndZHLF67mj01Cn3UiqLa
l2CDcYHVB2ikciQXtTEmehvmfnK37SP+cuBdpW6W8XvAMMFvTLqTTkF/g9H3cF+AsiI0suRektNT
0R7ZSOtKDQ6tk/LBgkaLLX34sY3JWe4wBVo+8A7+SIjme4WJSr8b4g4nntBgeIM+L4GVtrUjwsch
npYwts1DMqLP81b9y7wJURyHKsOrwcNUOJbQ32iD/snrBr4AxK4caQlei1XEZl+P3BabPoqmfnt7
hw+yNmFyvzbHSkLDQKi+6qI0yqG3HfnTl4kTVQZhUJkqT2a3AgHNkzLYGuKw00mdUw176MojjkBR
6lau+wWI/Yi8kipa0Ml1qscf3uFEqtPVR1j+MMSq7/LQbQZ2Y5VA2mfbOeAgjodpJnb8j7tKuS/j
lDCONX8HeP01FdQZJz4sBEC7roDzMNUVJ9HXaFb5y/8DtI1ZvDMnHIttjXFMUUf43FQ7MXybk5sG
m/2dtEyreHrAAySXLncqZcRyynAzDUpJPzngH4YAiHQLRQrBC9Em3F27h/qktEbyw/SWzTLGop7N
q7z+GLV4QwIWMUEOcijkAcRFr90ePBOm56xI9sIuyOfeV3BxKqNBbtVHt/ZVKmdZpN6rL7JKdsXI
pWnS1TeCrbrR58S/ghcoZlkatL7Inyf5AtLykfwbHHYJncbvN/R5y/LsoVG6fHioLevjCXeh4jgh
xkVzikQ6/MOTyBwzYpgtq2uZ6gdRds4QkZCtnfZsiG7VBiZ2X6QpK0lMv/lQN+qB9I0EOwXV/dbI
DjfA1/+p9RCwKKefBQAtspSDoXYpwWvPZYGn58zwITtET9B1U3ccOWYaGyP5u+GL9xN7Vr7PIgLe
oygnEpflW4Y8Pl/ma3zZF6g6nIJYNqPPPtA8DWRFCK2crTMAFxUCkKBlMSh7iTE/Zp/mCTPcaivT
KUursyTLTKMT5g82KQXTxxS8utMGwRTulpD7W8vlX+j3bNkb+CCfdB9BH2UjVySlWpk5NK9/MUOj
tLvyB7ZN9svi1NiOiRE4ZPNy6dZ4JiFOKwJ7Eu8y5C/OLBvIGLVIIGQOjPtBn66Q5EiW3cSpQNGu
yKS4V6KY2kkLg0JW3EdWTJWRaxB1j7Z+bbM2bs2C8MpS/bAVSdh7AKHz5R8v5gc2XSChonnUMj6U
nc4GVshUl4GNH5Oh4g0LvePfdMGQnAUr9jxsYBNAzkYXpEOXfUp0VrDb9oagoqj/gPKSQSAfr/v/
5rciXbejpYwNagM2C4FIHVinPVMlNw51h0mQyrSBVnvuEPgbbILKw9lGi71HJ5OHXrMdzSAqRAZd
0yYQn0LhKg93IrDMgfa8cujvIhOAcLbv0sK0FN8xrPmNx6uXa2my0p0sIx7inbd4UjJtYFHJg+SD
klvdbPmRxYCR08RSd/Ij4rMh4pbJ/QJdIuMFnZPCUqt/LZh122I1qCIoAhe5xCb0a8eSMQmY6sf1
+qaJXcB2izdP8IZ1C9mmQaWqcS9XNqvYwiJD8rl+EkGUOPAuaLZZqM3oeX/Fb7h/3ppEuKtFUCZU
FQNMNQqjeOsgZ5+sdXq6KhP//p60Foo6S0nOcKSiPKeHM4MK97aJo+NMj/IKb/OnlMKwY/oQ0x49
Kdrr/wyrFgF0Tgd73wDAXrX/KsjFbEfPXpTTQO4TTF0oZb7R6hfoDR3pGu0toLCqbZQptUna4F2K
B0ZripZ0LnAISSPXh4nRj3OFYGVHfNn32tuMnubX+L6eIpCY7kxlI4yxwTzaEQXJoZMTLVLN9AYd
WbuwNf4TXe8wuht13dkk9cd8+v7g0WNOCtXuqKeShIuyhkkrPJ/k5/5TjOIiOEYQWV0Q/h7kqTe7
iviqm96oPdXxO+EFKUFeBioSeXiqFR9nIRuRN2amyp78AzNjEJkckbQvwS6RwVHkokEkwo8sZCVi
WsBFfQZYznS6iEk/h8m8uquiMUrzic2XV8BbZeIgvEiNx1NlQbDtGEbKmymx5pD588U3AcMgRdre
WQIjtObTDG+cUcUBCf7j9rdIU6uUT/HPiczyjBF29mSNUFU/q04Z3yQSknxEVFrVrDC0FArxHRpy
YJdj8UHEyijnY0k12trur7Cd7PllyIHZi3nAqZgFfuqoTIJaHkw/WH6SAyispIf5Pl/CpF3wpY8A
SGJoglIHe02sKm3H7w/LZvxQLGFBlof0eE8xahPkasH8DKROADvsjCnYUVDpVEKIc5YkLQn74s2H
NHBSNAMwugPadSf6ikOcJ9TFBCYKGl5JQn/l4CFyatdPMX9HVy2HzAnnJSptVVvLXmUDhic4QoUM
aE3e7/vX7cF/rkvdCaVozfwpu+4HtqICGLbFYtVMWC+Uu2BaIm+p0doPszs95nj5WB8/dtVZT4fc
gytuTSpC6I7p+YSKwT3n95UN9RT0HMER+reViejUY/XabjjZ+ioMUMmUBEloL5A2C8yu2+/1iTQO
dhZdfmWPD8DqW9jW4En3Hwd4BnfZB0E7t2QPdA+2SopgjNDBtNjEQcjiz0m4bvyWeSOFCQIB2Lss
glPn+FhXfG065h2iPFlOAKzOlOag8jJyxwLDd1tWHBpfmGSNYHMr47RqpFcEj5pJ4VLeTmSqLt4y
AQQbziYNMYKlVSFEMdqXsQP2WZ/t/ZBf+irL2IcjSTkIXGneQ4akCF1LKAYMIIsSRSL0p4s4LMAu
x7K0H+zOfbLwiSRK67tguy6bFQWoqYgF0d7oC498KKDSjrW1+gg7HGUPfxHwFlPJ9/XpzNWo1CMW
lYtDh8B/RDhMGbmanQAZ1olAXSdXWQNiVJVQELpvkvFYFeWaZhPy0udf0wRK+RI/1UCExsSSCpVB
Y9vrkb3tLsNNc3u5ZclUUwQg14pwOq0De05/JIDH3PxivCXhZVXz2HIbSu7tc6v3vt3tqqDRbaEE
hotOogjFu+rYaRrvDKAkJdYW89GySRlmVcCShHuIajnlB7xbm4sAhRqPIYgffp+nR6qvWZETYINk
IqrLn8Y0FHmqLeeZwyyD1xBKKit+p7HZWl03QSDler3u1F07hRMPFOvTt0fLiF018lU4zqPRlw9b
IOIe7QsioeF2T9hfzwUO6YdnTuUjqntcmCt41vP/8wqNHN8g+z07vl4QtmwFfyvh/wHPr2b3MUhE
jwOQ3b3lKcTe9JuLOwhg4JodNZbH3ddTkq9oDI89MM5vdw3AJm9kLaoG0kgQZ4ih+mHSH+NNcNp6
0i9u1y+Oq7SCfMPJQ+fYpKEUIHqx410FuGDsWA3BHKhYmGYGqaDev1O20ItZ/gKaVUO2viWlq5gb
GMfPZn5FFNnBgJM+lwvzS4noklRSI/MgznRsU78aJg+QCqz0HfDa02B6gtNrDgTvfrmYhbSXSib9
3NPCAodB8zitMnx/EMx5pLZALP7z5ECml2VvyLO77nC0gwDJyUjBYTCSdRRXD0f/qJSk2coHdpjY
KEthfkemXEzErDdoiBICF/xzYXL+LsHSa1enPZ9ICVpubClNA33tjoVzfdxrAmTfwcHEThTYY1gW
jJgKDSjjNFL3AHYD1asKhP60u+sDQqCX+CN0CHdrrdBCbPhJdv6uKzs5T9cQirrY11HSLaWMJw3r
JLsM8657mxNhJqyKlEVqH8NimOYH7uK2VS4oTrLavLbqrNjNPrM2wB7ci4a1jJZEMdkTi7vHM3vA
MFfSG5GHi1X8vW4u7dWRjwF7ASf4nZV2z2wKztA8RgXrd6Ay8+PhW3MXrslwO+RBM8j6OGJmvUqq
uMMOWUBFxcGoPdb+ffVIzw4eixygxdflFLDbi+7rwiIf1/xQavgjsLdHjMLWgcmT9kLZxlhgznFa
PaGyO+D75tZx4MEjv66eyCwpaZZjxGn5CTGPzAValJqEYQN5IAl59baL7ED7nbMc477oh0B+Vdk2
iOg2G/jhpWose8BK5byJrHBkz1pWKjMXcOkyPFQJemQoLrEAekutjAL+AOOtHDThNeFsZ/hBcYKM
AHqR1OBRlbO0Ua1VQx7vAkhjOTDJjU5DpQxl5WvXL9/xe5nHQ2lgZ2DOPsyP4uYSQPr+aJfyY0jn
6VccOy9exJTiPUe2RIHAVNv/ksHz45hm9r6tdl8xbxWP+b90plFAZjARcmiMgtTnTp/HUqjhonuH
U13NtjfGAiqRn/72tTfYqzAoHG4F+p5N40MsPiBco3epldqOt6nXW1grcs993zYR+qkUIjz5KT95
Y2K3IglIlW7/BlgocneX2RFYxLMjMFhrPS9R4nrsxnZ/jFIfYlYh3UVIL/FVZMOC+NNhYb2UEyHV
gt5u0AkOD8rGudjfzngEsrir8eRbWSBw/BllzViTvjmxpofGjJmRrA1igremzBIC9RLGP9Qe3LOh
5CsJPUjXyxFLmVwKmO21GfjOpbGpSvfLYKxB+BMeHHiOoeUNBZvkG7rNgpeIQQcYreQMJ5L96el3
+45KZs7LBDSuki8ga//74bwY7DarRRnIO+x4k/6Ya7WAlFs9f4K9IluV/faRqnD49yDCJr9IF3V6
nZ6jPEF9aN0iGKX0CKEaKHxwz7RvXEiJimGLF62KiNL7O1/XMTcD5qLUtU3ofOomiHlJ9+XWRx13
aJ3ZAIC0HiX+7+cU6Ytg7zxpecDqWv/M6Wmnhf7LYxHVV7A7ocBrcSJoE6G7YGD2QVPm6FwTSY78
kmeUvbjVL+nYwX4zC5fgFWzb43tBQ9mB29xTAKr/fi/NdZbBICJynlvDodIYQ8I1CsTIMVOG3QkI
d8uBDTZfWJkuMhZVaYTq9P6NKfxIWOJfM+MKYiLgpnGh+utOi0RCRB+ValF27lVBM4Y+unAFHekO
CgS+YU7G2st/IJ/3h3Lb14gr/fR+0UzPnZT/p5BcDF9U9/7JEfKMGd/ZPoC5vCQ1VttFldEL+0Lt
WAvnUn6A0S4EO5A/bt+aW8UleGHF6umkghqq9qSDcFZ4gMT1hZRogcXBdrYOyvRTR+GT7aCbUcfx
OjnGoBLvOLsdCSCSEajOqstXOH5y9QCjkWCC75rYswDSt646c15EWrr9ts306GVLQqtQkVmRxCK+
d5BiDxY/zk2/KlFKKAHT2PmG8rzepS4epm1hjnea85VN7/RvZ3otd1jkWLLvVVWChpKhjpkP0+vZ
9/d1Zz5Z3jviU6IbCi9vVMiuK67uuaQeZbvdgh3SaiJmphOGfrXpdN629GTsEyDWiCaWk3QRJoVh
35LpA2FegC5n9eb6tiCNL5EIoKFWi3ho7zMhboidfBlQDSUjDOUTpsptpaO18CUQbdqTHhKRXERG
RKgzKrv5ZQF3haGIFFXZ8z0MkdIl9lPVlfmW3BCo0ZENPlRy08FPNl2ExZgPd2nr71H/DPIQr+Fs
vaBfxucXMQ4opxVkIddZgnKbGhwi/t28vPq6QLPn+h7yrRik1NFNcZnIekhAmY7dH3QmJfNeSIjH
AWpaDGIm0rcWBp0csd21PHLvtYyEBWd6oAEtoIjVPyrhcmRjrueWJzOBjv5seBqwD8yuSMdoL/sS
goh2HO+6jqBahQuvQv/AlRUZOn+Tg/kkLUHZhKpGbroyB00Hu5RHcLgU/0Gd+V3vMHeCO8WWj5+4
nSSlZfz55g9cVADN/4eaF1lcqqar1CDSHJ+g2886P6A5T4vq6KiSaerTsCgSn+CugwcXXgiufl9x
xmW85HC/0wpe5jvT5O08p2GDYVs7TroQur2WdCP8HNnDhHfYNiHFbAset9+E3cGhDqpF2lwso7q6
J5geFsBe25O8OAs+EoClUG3cLSs7N1mQE7L7MUXWgh+/vRccZunSaKhNcZOkkSZS9QalQKoY0SCt
1iPhA4IcWu/0LCJq4NQ5rFiKwVjzIyz0ofzLXANBVx6S1AIoHLlGGjjztG5FsNm2ma8AoqwWx1QD
yVB0+Mv4NZCb/rQEhGCWhL17bxzCnaUArgzlJY2ua986RZHrALl7KpI+/WJntqgRRu0eJY+kmKXd
BM0Z8GKWktsXioKr5OtQU4sELtfeUwIORP705XZ7/Hw++2f7mGo5M3rGrMETBxxxBj/9VS9VudBc
Ahb0RNj6YqjBn2jvheqisxcMkhZD9fC0PHl++XbFSdzlNc7lewkGmIPFCETaeQ1qFuMAhoqO55Le
7h3Ft3iyYMgFKpkvTSMtFZaf0mIOeF/YeNQtw2bYPYxH4bi4WhiMihPNvbv3uAmMmC/gd8EX7xRe
0maC5p/zQoO2fcNJW8n3Hrk97bRd3LAFs3A4v9II+dsn0oP2kzNFQ5VeLWZPSqHleBBoT1WSCIz0
d5zbrMvtAQVpEqIxKvs2+UHgWMKM66CTmloFiB3Gq7TKGY/PwEvAP4J7Zoub9v2vfmTMGzVGhx2F
gynG/hxMPtTEaC9F+ISNnJ+LLQIfuM3V+O/PzlCLJwI4cvHV/rfKSoEx0S8s8mkUdqPAcP4PJTA0
XQ4oQjrVRc3RhMwpf4PIE/Dagzxh5pmnEHDarB9OnNhzPVc2pzH9IDCkGuffBFwACjSiaPG79yqe
CF1W0TvvlQsA+j3nDJt2oTgDtrtj7GV74QgNSjUBVhnMA9+BH7Hm8ZaLHc8ohvKWoiHKNV8qQ16X
NU7pOQ4qpRLCE32AawAjAzJqN7jW4mBI3kfoUGUZ446aN/EU41lpSvk87u+Kc9WNTXoXE8ydXXtK
rJ8bIQCim6ZY0SX21NHZ6h7woklT1D/iQ9pnVj+VAsJLrOCb9pjGoXHcNdYIajQGOrE8jQMgzOoQ
/sJU8RI6n9qjN/ThOxYzT7tMAV4WI7W2zv3eY3b3d7l3XKXxu/SRoia/5fa/XcwD/Ggpy30y7zui
O+94nGhysM9cuf3TYXDZfRuiNmvydcHbYe5Qzj/dIjus2xE+I56SXkczOsh2TNNtCRpcDMVj8kXt
p1VHjqr4it0oeK+R4A5PrCly2e+xGXdt7BMNpOLKx3XXl4IvgWqajuiAz23jYwEH2RbnGs9b6P9J
q92ttRRJ+E5CXFUIn6gUToHqHy0A1+XQkElnhZ5NtvLNOPNvRcLIuEc+llCI3eA9F+R46c5HN0bN
le7iJoOKPsMthq2gdUj7C606dl6igPzDxR48HNUHeXMXxIS2ytcGfZWpLOYNSt5E0Aje34q6SrfB
llQ+XPmBNwwHnE8iYVX3FBEOTvlclC5zDfyjAMk8/iLnSxJaFhyshdXTIHibkyTcvtfkjLIlbbi7
kExOh0MTzjiEEMXz8Nbk0FsjaAy0qbH+P+YlV1PLDE7A2TZC7ZopOWKWGNa6N/T3D0FAPDL6W0Ca
XJSGldH7StSbWXKWdAFWl8zy8U9rLy7Tvi1btiT35jMN/15QSekrTWzaPOH6zAkev2NqH+Wm/966
YMr+voYFHp2DTsVpv7OhixjwJvRP6BXdfdwhSuXhhckjQzz7K5Y6r7YgSbn4+NCHdNjF9ZmIu4aL
8BlnBu6vjP9sJRXY7lZ1/kTEpnmcB0/lLzRf5zJzoaNnXSzmmCPZ5NG4qiDSEIMtOFQv1BtyjWpI
v7k8PcoGGXKkCY/kvBwbFI69yqOgnsnPSvWwevkh32Q80snFbCjNTA0eHLx5OVhmne00dvtCqm8j
KR5BPU2qDlRPaAr47ChdTbBSl3IyePtr6+NMBvrjz/p0h5bYFq/wt4zhrrm2cNm8ONbvoauquqZt
vRWfOOhRyJYHGVDG8x3q7wR24uGI12OSjeUJWujVieVX4s+27If53Gdi0lrmwoisk7QrvgRoOzA8
4xAlr34jAzxYXVDb2U7vjAk7a2fDzY8BnITNO5+/5v4J8Gxm6HQuD/RY+y7rz0ILTB3rs4mwyHAu
vXsfLpi+scAZfsTK0gdPmTW7EvscdANwwAK5B9epaWuVSxZ2q8SG58LIvhllwhmrr2Y7Akh0ggPG
1Ur4+xX4lZEkiAMS2File6F/YmvDLu2Cu4DhEa23cjVGLX4OAnTPlZI4j/lV+CS6ZeUkIf+nfhSF
A6aJ54w7xmK6p1RsKPvcFDX0vtL7SlPoitS4K4KbW9XFwxyWHfTJmafG39wxrfBeR70mxNYUaqSg
muvWfuiNA2rFN+XXDBwa5LDzDIznY64BjxIFWj9t19UKOp5dczMxtav50LEDIVOOnq9KlglrJIHK
zFCNTCzB4wWB+a/nKW3aStqtBK/fcE0PjnTyNv4v+uJh0S0xNl38IFKvCuPKXKtyrfK7hA+c1rWR
ZrOzj0ktB2gjDGFWvxNrdip6k1eVP161xg5jOg91CuoqTc7e3Ob5lWmTHpCh+vlJImsZhaYnyV5d
fVnoPZZZvOhFZ/TkxSxOVsmaWY22qRUUuSIneGrJSQS+aSyP25ju9umeGe5qhEaDKNp3rp0KC6c7
MGZjp5D4QasLRnt1eIYvOtm68QUc0mRUXmNG3Kqyw0ORCg75fcQY0GfVQw0cCqs8sppeQK0+mB9b
8ujYgUYIZmBtZdCWKIn40f9rC/FJTWfZ+z7BM2y1LNAbpGJAl2neNquzqW1QEUBAejsC8E4sGoPT
uZnZQyP2gYHs49j0PHbIZn6KcVUb3gPCiZ8Km58Tpd/4wLm1TiC7fp+YE228RN7z5HvvY4pkO066
T3XIhj0Ct4nQA1OpZvYczUQSxyS8tyCy5L56Zi4OICEHJd/il5AA5bBuF+839sC2F9FIdeyfFuC6
tYhMRcKJzVDcT5fXn0ncLPEjY4yQludcw1MIqXAt8Mb5BU1c9eWuK6dKoo16lPz+Z+OlGlFW1e3u
uuvP2ofFOhwFqNfFoV/m9jMK+RGCrZzTF6wu8S4iFtlf6klNX3DbWCBrwqOJu8I5vLAmYzFh7hS9
LrKDCVb+5+DOzRtgC0drodaLxAUHCUtyNyTwTOa/vFPOY+/XIKqCsufii93QKPoalW715Qpu2GTi
hcN7ap4MfIzj/MHiiuRYL5bXZKKtGN9BXPC58fGjy+dTWv6tvuB5U2GpOi1QZ5P+KOyD2zxYlMVp
4JLRAMzskbCeX0wbemDNkrFbASjUnYkJ2WP6debg4myuS4GwkCvgZthL0n/MHZ/hZVwe9FyW/rCs
wYK4KQdUHyXdVwNym4UF+oJGkKnNd4WGEzQGRXtLm79liHOk4J5B9sr0bWDQ53luMYQro0Z/Oha2
yIzE/e7RaMALvxgFeiTMaTgpWuTkhifiAJtO8zl4rZvxjFgRZVtj3DtuNlD8N1UlbkzBuyTOhYat
dYfxxzMzWdoVWBwpih99dq35eWlayVPV7AcNsPQxYVFKnItRKYULnyjxf/ZJT35Im7SUT9wQBVLu
Bfrx8Y7TpXnGn5Ec8OYvChyplqRu4vFRIw9sD7B6mZaS5JSxPlG7jbCECYOYJ4Xu3HOAabqKsp+Y
SZDTxYKzresF9fxzjA1cO/eF8XHq05fRi4du+pmsFa6XvlspxH9mdJr2Gx+xp4NostX75Vjn+ugM
hoNYd7264ChW8AeMP64+0fIsIREtLnc5HzTgpikVOhTzPn1E7gZgD7bX2RkbW5rxh58sbMrJOxY8
YZhXdlGSuQw7C43wN+LdfhKFQliFIxOXlpcUyy3x/PMczEMTDHYrc+MeuWfCsjXVexrVQmG42sqt
96u/cM+tm5BhEgo3L6MIwGdb0xmSVfyIv42YxMajsQa8SOrm+6f5xAwtFAKNldyG3X/97u/vHdzM
YWQAtmhSoVAFSWfFBSwRTaO6Nn3XFZkT8XDGrE3bWpA/8SgCSeJGbxHDif6lHPmozP1EI/f9EDoJ
VFWwdMlFoFZWQ53H2ysXTETftxvp0yIv5f0zxKOjbWy1Wg8h7IQ/9sjd7SVlQXNxJ/kf6t9F0+1/
PhE0EPfQDlju6hWC4urD1Fh/ITk4qdMxmauG9xwUUiz69xx01hSloi9t0yoiVVE7DTyPZnFvzy5G
zoQBl9YPW7ofodTcfBIYJFW7DjlDGfrPJkeMWJ+WTRH8M+wv3CViaxxTlqXUX8AUdrTo/NuSGJvG
x3f2LdLPoSInAQILgWZ8sDMAL6s3ZbyVhRyw2We79RF10ix200wE2Y+gW6RzB8oFVqoD1BSfifGq
Ry/iPtTCwOGYW10ITSHLhwsNZAPwvkdv0qWFvMPaLeREp9YXy7mkTfgrPqbFCz2j0/3oqg8ELakl
TKm2zudI92nKl0moktVxLEcDKCnxQLl9l2yBjbv6PWZEtSHOtaHJY1pwcI5I5uChjxpjWeJkqqIt
WfvxsfHjnKJfgJkZMXpuU7jQO0bYINLDuvfSJIoAHtP1T1uG4RjxPKiNsduHheprFX7RdO6ZjFxg
OZLe5fzj/LgqwCcoZThMNXmKEVQmYw2wHcYPB0gz80rFFou1E8+h6jIuqjSUbFMdUiGoUcAqkudd
i8pB0SvD+HKRkIkUuJtQ6VjHjR4hvDvuiUXiw5rumkJjtW8I0svI/x5G1wnFc0vMGXHgLhYOQz7n
ZuqeiVZipW9d8zlTXysyVYymUq/z0+5jiiBTZQYnXyTps/SBUf/WLgg2IDACC07m7I7KvFsIfXXN
Gvwfwmrjlt+ehENnhuZ+2A3LAPgelj+Iv8zvPHaZTrXAdKk/Sq7+bBLBPvwu2ggzy1/yjC6I9aFP
kd4nc8YcVbYUBs6fgiYCmAM1RG4k+bhuYod4fDkS0LMtbbEUHBo9EWv7bygTUk1QhS64aYou7d8j
W1l7gqHSA6OLC+iFQ67WGZ6OE5Zu4G119oQORCozfWCh/58FczWmUiowniHDqToRQLclMfqkpjxa
7jCLMZlv0IIwDiq1zyY3xy5bfIO90vaAd+jEyFJH5yP37kdgw7g8PgGV9CG9nH/HkJqmz+GiEHHc
MQP7QadLZlBXUYXORNoKjPyNpbET5DDGHVq/iJzJdTZQq0To5goDkFtxHij99i2ZXfI7CujnKA/o
/+qUbBXWu7xO4gxHoWJvZOsDwvcZBsGdbCmqKEimZMuDmxUawO+2Q7lLwOvjRar0e3KvFB625CPw
jnCQZF/GLA0umUTnahuS5ERET4nMh7ecB5yo82CBZwdCre36JwkH92m49nruxPeZMK5viM6UYtGN
/KqCqCxtgBiW3FG6dgmUYMsdVTp2gg6z7Glz8CBhe3DiVwXelyl3vVX7e7L+Q5Ha/d/Izcpt9mLZ
4NlFS/6JBWX2niz9q5ZPKFwKTT7ZnyovTBXdYeA5gK39OAtCvB1Xmgr6Ui44S9HyBdTXzXx/gNu+
nh0hm/jd3aUfn5o5a5z6lywdyt6emYLGVRWFPU5Shysk4+0hUvMU73fOqVbp1fEmDuUk+iSzf+D6
rdSZmnkJ4TIlWKMU/RTgWpF/wjseSxXAh5vz6yu6RTjCmh8/9VBXjt5efHqYtkuQrGxA9t3XCy62
YtiXgbpvkYK0iAn0NZSTn+wMrLYMV9STZFQJM1FtIFCcz0lXXPOKVnWjegLlM7G2Ky+lLt+7qu9j
pV2YhN75YAETHTm4tkQ3L6Ub2nR1em7/Lw8RlSnykg8rtMMguRh0i4ZGs4a5pfND62xX48RyHx0o
IQ1FPevDJA7+jgogE7nAZuP8pVzQTZyHJtbzSkw8qk3KhsSuo9jx161W3LuSO12IHznha2vxW/Mv
1P2xU/flPnXKq/jk+v6rG1yVngRhRwKowRaHtvPKZaZUPO920uy+42UM4WhupX4/tj/xurbx4XhI
+zlqwvkwUt5pQuc5stOLFsRUdz5vOJ6Pj17m2DsURRifhBp3D0YiUiVAwlcpXHNDYpZgJBN+Hh4d
K/rW5XtnKdVMGYLaFHPCJdnfJoKRH+pr1UiVh2CDjukeZuVWfMUsmb+DsBJ7EAmeDkPwTvBB1ImB
mBnQ+oyM9qBxBoAueZlWIq0zyY1zRnaa1dF94HWPG1C+wxCy90FPkt2ddBriEAuPxDGBekRWw6Sw
698Opv4gSt/ZCfEno9J3ml4mHzFmEoiR1od3QzSHj4p8Xo10O1U9MvU1uOas2SRJPyZq5KCTNu8c
3u5OL5BN9UAdLS/8zXu+QRUyd0xeTaIqKJ/U0qTxiWfb/h1hR1yTsmRze7+3u2vM/GkeCnID/bq9
dNBt5ZtJCNkUrMUjywPB6x1Yk78jpsJH9aU/ZnzhF4Wj4QkwQMjxUqIOWqX8jn6wCARFzkWbkgTE
RzQ57VbcsKZgE1dGHfSXfLOP/JjpFpZRdslQy9e2BPjxro5zMLE/FpEdjuBYmzCTziXjfp6jnrk3
CoGXf5jM8WVWbWdvnLdfigJtTrLbEkqdfX2I9wX1OGzrGveqhyzoVuC8l3GIEdfEJrrtGZyMNIDV
DQ/9Bli9rfnLTSgLJMHOGC2rl4a35z+hf/nVHpxjzqek0yegyqq9QuqSUIMWRN8Wzs+Fr8RqyBqB
qAwEBbrsFaKJTqr+zURDbI2lC1CYDRuUlC4r8UbdttXsk8UoT2Plj0hJ6zjC23YOhKxVeAGMdwFs
oad3SNGiuwZ/ibhZqOBGtfcl5dcjwhUxu5Y2d1x9mxixmRbqhlt/mSsB9D5TDjM/QPngLXZq/bYZ
XDL8I6eTSNYBdJzNgYqBgDGbuujYGpY7icspOLZ9CvINgBVvBdr40ACimjTyijcWdv+hlKI3ZTT4
fJsPF0wtlUAhFzf8LJeFqmq/uYU3PfcQXysbSKJ/dUZ0Hqf/YK3Y2Qv3hda8xOiBo26xCwSZPxiI
kwNuP+AnW2/nJq4bSPX09DlRgopONd7iKb5bi0WyBGSd0cCtiBfbClDpEa1J7R7uvT3pGbVEknbZ
h5KbRsaJMgBZwET96qLTPIFXTVEMWpMgr9Z8jBa55u+hcIM1JLPfgy+q3W80TVycrwjocCGCoSTj
Jm0tYZiyrDp7KgPgIQOnZQR+I+E9XTgUvhIskLsB4OyAZc/sWHr6fXWTf+IPkT42OE1LTU1Za0B3
L9zl8HH8eOMWt1boiCrg7EDUa3k8rGheOJvj1A0IAhBb7TrhvKLUz6Uu0lfQZl5lCrxj8bBP1qq6
ojv+rwC1OQ3fBuTzlcNkZ50CsNp6hgb64eGIHGHSXad8SYMj5UV/bsiEGHLhx1K0+93OJgsAsfO5
dC0/1pxbSywbwbY10TePh4tN6B7jY3PNt7z3IgvS1PoujF+4WotWdux4WuIaoHDx7ButPxKXeczT
1VAVvWJC17YdB427E3lJwVuZSf+/AM0GKmBkTqJxJ5AYVY6ENjPk4HZHLAJygv/Rr20Y+/VSdRqY
fqGwH8NkDax/bXyu3m5uhFzu2Tb0TU7JeQIzSwb0yq4IXJaZke9Utpe+HPLoqNCXpwtPNKh+7hSW
lLGJRHYFaHor4jcyUUC4ufGwAHhRnppQc8yJ+qRNle/I6thEufJo767oSu6s4eC6AA3Bsg0mSyEV
k/rRDUHABZQtI6TH79Bszkk9cG0FpsmC37Q5V+pYIeBdjxGZdoXls5lN2vamdKPChtzMpdr3XlD4
fYMp3Qn3Tb37NK9XOiamtNOHsAv9kfT5XTGbpaPF7QRcul6e8oRU48lprb7fNT7hFb+wr613Leys
BaLi/M9RgQcmv+JtS9NPKc9+ughST38RR8VRPLKCHBEuLHnvtSAvyu3D9EPg1//p3c/eHexcoIfE
hP5pfD1J+klBJx6aqsDcVzsDR/5NvB0ZhXUAmK09/FhP0QcZ+6JWs4z26r8MX8fc9OHaNER9XgC/
HSPOKgbvZ4p8N/Op2a9AgsecXCT0Wz4WoJ3gz8kG7+UT3ZaRJyu944qMyXK89KriUFFdy6/AJzMB
gSjojqZW+/wcqGq6wJABVk9gjwdilEc3qhC4hoS6K/jP+B/aOxuQF+aJVnZm+Mz0BxT53LFzMCvh
nK6o+w88pweZ11XY9kXF19bOjzt5rjfBgnqRtJ9u+U7hY0aK1vJBGbzxvMeARKXYb39EVlj5j2Tv
0FwgJJAplZ95rowXZvU7oNo6v047BNkvQcJcaMmxqkj/4n7kZ9yjAMeyB2u414ji1blIh/sZjKAy
ne8Ho4sxDU6V+FrVJMi5YT5S0a/BmfxLP4IXdVhT1pb3/DDPmKj25KtAbzQBgUqawi2le+sRQHyk
frFno8fiYIYefP1tJlZRyldGnN2EudhIeEQix6jmWyNlMmS3uKdjbWnzzAA1Wpw5n3a8Ofgmlskw
5zVeqv5c6FBKMFMUREAFVMkgMOGbG9jRwRHvuy3RvZdCGtf/INoDZNjdEKIwYCZcnAfXdjw9SdLF
zewwy+ULKNxxaoYTLqf24r/TURJ6tV7aWdlvU8YVPuJ5Pbmtf4cu1nf+MrhQd4zyHIjb0b1hSXjk
vWdKn0ZPOV8diknu+pVAx59EypN9OYDcz4eacSbir1c7TRsmqXixxBLRLxOxrYYbb8yRW0+MLIfe
85/1ncIwcXCAopTtc0ktG6AWYIppi4NWBriLtFT9yBNpJSTyESFSVtKSTVPW5i4UgUXRecRWYTBS
NBxCUz76bYZx78ATEcqB5rEOLJKYeE3eidp69dufIVmDCNAagfj4lCL+Q1sL509zsUdAF/pMkhKW
0Ozgxax2mwrrR7ChoMHvkRLvah9duazTzlPKpuX8SEL8awMyx9eiZBPjF5yMhGcDNQPe/leg0Up3
FwUYhd+8NX71he+PeAI7UQovfklZ0rnXruNK398eMFZvfSH/6aIGXf/FaYqwuVrywrU4HEcOB6u+
mJQuZu2R4wqHlzI6Sk7i0DCBV91HJ3YS1DzhRF1c4FbP+qgyxjnpTQTAlvofuTxQUujLTzp33Vjp
3CRA/ERg7AmcOCdRyr0zvpY5RzHGYj8oyniQm85ZDWzGvZJjMvP4oRGKHjEet9/CQMtYDEMl646N
rEcAeSTAcGPOCpdg44E0BokHncfLDFFVoBKK9ARZ4RDGxMzF5+yOk/0uEJuIc7suysnGluDkIDbZ
f4G3RBxn8CuLpbVJqxk4eKrYcmeAxr/Awfbb1Xcl6f8G8+6xxVlm0CUMgPjCu57bDgODNcRUfbvj
DDrJM2HPr0pNskzGx6MYsqoH2Y+xeDdL9TSOGAPX7av51ryW/C/8AYbkMwmQLTjw2bLKG7lTLXaN
CPWtGTS+8slJrQi9RaWWzK0LcKINh+Yv7g4ocDItMiQVctbXT2937+bFLmeyL9fzDnK/5fTP6dL3
w+dVKAKrhHSgwqWzBokiWBXvfXR6ydvu/OoOLAA0vYgYR8PU8gx/XQF5pJ1ZYaEdwobRBrp8mGxh
cTi+m8Lg4J7wSIWw7I5rIKo3o+mVZ3dwv7icIurPWo1m0JGpXtUiuDpFOY34qm1sgDbOBecNWJX4
u3W/kZj7yLFOsJvL31jbQkfnawcJnYc/gSmC1Zp+jdB7F0z0LPRxj9PJnIFzKD2ZMGn/NVbjdzaR
t60frj3ubPQZANavYIvi4ad2Aji7VptOoTwhOA1c2/90O1NBd2ocEITS1hZvc+K1xnJLPo1peqSV
0GKcL55lUkkzC+cHnPq+c0LTGD9tO6PJ2oE08zsCIYd38BGXzLfr3Y9PQ0yw2leUUuMIidjWmOgp
FfFFcOHGirkb0yR8c3rBmoJGM9N6uIAqPd7eCZSbZPX9US/a94QjGj+bAkkoe1ZYQ5Udl9KJ64dN
d91EtETepvqrYx7GoZ6HzL9maExDgZdPO7fqR/xKXcvqJVWZUGzJhqvDcxR+j7rZNTopzGIeYAD3
RhM9VHN8O75ELf9SIHcKPpRdf0dBzg28T+CdLKjkvAs900e0SU9+MM9Fa19ejOXzZgNuJ7DamNZB
h0rhksaYbUXBuWhjDnzw5Z5u45nt6/UPb895cj2JU/kzeP23+G3jkfS+39ubzYVz0ZQ1UOYIUmqq
7vWwLQnT9Jqx2tZT+gWqKlIF8ELD/uI002/1jJpcZTl0g+KlvWw3nDLxRzHd5QCp8j4OSLXmEO/0
fVkIsG9d7ThWjuBBVJwAIHblXM7RUfgDhIwAF5XPyJjgY/vn1DOQYuMCxrEPJVcWEG2hJVfKY8pC
pcsyKutefTGWNLuXUKFhEP7cGUajfK/TMuk4jRW2oglzZLHwi5LWkN11VTuEizJbuduC0fFuDPUp
qo2ZrppkJ1Qs4s4p4fuI1UKxYAwJjZzqNTA2CnAJVqA/6oldMmxoLmJHZgTNWcgMuSBq8gti//10
AM7BcYSew5g6hU5OVj7tKmo7WHIjlTHnODh9YmZDJHllGF+ZMsA7CnB+EvUx+1ZIxGLSQGs+PfqZ
kYZrv4JOrAsxWuqtQW8FZiqCB+ai0l2yfUWWBUPmiDh8Fp8Ks6Eam2mOa0XcX8Hi8RrVSNvRQFvH
93zxdvb9MsF+2DV+urHJkAWg6g5JadD0cQjriUArECQuBQ03IbreOQwxNxROAZmmOWj9cEz6DE3g
SVq3V5E74NdiNwFswyuCwAZLnhbLuJ0JzjxN8eNp6Sso/Qc1NcQWZpxDlLq0VghJ6BKT39HWL/bS
1+NUzDWS7vGXVrsdNM1KfHBskuk1giSZ641phygO8zSQVMa0zmJeuIhq54GG9lkDiyLUCgtoHSX+
3+vMGVSPU9o5wCpwucW4gU4tlC18FJb2weY/KUpCQTfkDIibDRAmV7mmVu6icMTPHXtOXn340uxr
Bzbw2Mw61S+H30Lml5TKGUijuAUh6jOXOwxwsXC6Rg5cqvZ1nw6ai4AG6BY2R5nTZ6QTBtoklV3u
raWQmDpePGWoP8eiTcivRd1ECH0i2uy4FsyqzScXweKoHi9u8JHoJbqiZzLiqkL3Ir8mUz2BbHEy
00kvsWQQ3wTh3zPa/KqfMC04B6oOlBIFyE5YtSoOP/ynhfPLRMvGw71/1lfSbzIi9GAISRrY+SRG
L/3V4bKWw1eQuWrT5WcHCJgunMwtMVOpV29d1gWufcCbTtF0eGn6MjhhpcCwkN+n3XY4BsDM11Iu
hILtVmLHMjipcBg9Sqrgv80r3DOrt0Lqsv6NliSiTlR7Sb5lc0NGbYk7DbPu5Zp7L8wF84mKNQWn
n5eO1IVz3riXDGgra43/exyCmW+73KYuhDVV6Ydy6dwgDkgfH9nQMG2ovhoGWy1FRQksXaxDchrV
rWkt36/s68EO2F6A0agt5Zzq4fF95eoJ+fH1tam+6mOgmjPpqdXZYSGBZBQLGxRmrevTV6N01qud
y0HzYxqD5oarWX8iWc+w9c67hpxF3YQ4FvkTAHGkcmuuS54D9o8C3wkPWDStfdZcrS9p2IV5A1PM
hIOwvO4PX44/iNfJSRce8blPsLbjJBWTkkYIIWMKWJK9wunCAqsQgg+epHN+ZCg45aSI2VPYRFWC
GuJ3/l4i9XYWJpgyPE29U9cYVW2mfZCo4YREnuHsx53rNLoI4W/P7My22HZdCuWSJhk5OMhKA8Um
aBhvj5uwmAKgbZwIjbyMfGijiRkEVedTiUWb7dbSqwIcvnVBkUrx5Q95rMsdC+AvBDIQmRStdTa/
Lo04uzKXVpubJT70dpNslZ0bnHqR70jxkSSHDauRvSjurnxnFSYDjUbOBzMaTcEzwb5gIDtLj2FI
KOxuITH4+ibcgi0iKeri4B0b0GSuxfo7f+fvYI3sMC2EYujyPA9CPbnrYwiz5LqDGHuWJKBKdSrQ
YmFhQuqQKkm7ESyNT4XFfPw3Ao2qt32EGzZfEFZd2+tcSt1So7F+jk/BQTPF8+Vt6pzhok1qrZXD
yz+YskTpwhxxe9RoaGedist1ScAPrqGCvTrzAfcI0O4NB05xh5zvIDg2FL+4/osPbvKhjrQ3QPbk
q/IyezOG32yKIPwurCG0gsmb9hzPc9i69RENp6Bdr4LNlKtANRoW026+Xlpf2uw1ik00rK6UOqbI
YR9aNSKsUAhynIW+o1IGeLxB26IJv5q363S532XOCSGK91yT0AKjnp4sxQgAGks6RUsfSNnxx9P/
Yx2O3X98yblRFpHOjT43PhpluPpcjLsAH2OeH5nMXaIVSBsXse0jKmy3j4ugt3sUTOFgQSUmKkgB
TzhgxdWXZIIt/i71/q2eFbCZ/eIB89fxqHy3LRWkIMKrB779L8qOL39CoiIoXeN+qFOkZQ3oP+6Q
ztfW5CyX0Pmf0xCUKLf/u2VhXYCObknBhKIrKAIGIGKpX168gJGMl+x0ReE5GYr13u+0Sr3OYt6Q
DYxEERH84gPpvBbdwpYQKB9/3s8S+VAR/N5JGvnN6V4CMMxtIkecEJZ5ksWRaxuL9q4YWP+vivs5
7tTwijFbMFvY1FLZAMh6/nO3yYNByPhluRsMeY/LDoVYqj6CX5UASfVxrnlkwCijrwRgNPw+WjAb
+USn7G0VPv8uyHYVFFg2WV5vBwPhrRaSAdeO2IWFgYWSB/qEpe30BeHONEBCQG0Q7J7t9b/uOeLH
2MBU3UT2eO9j8+szS2dIQrtqVd9FExBibz5zjMGdwNazNgKPcYhMrojHI5sZaCJvOIUxnC9pu7wm
VVf6Wh7rO3o52B1H0gWnfIgj/OWTXCGN6LwFeAqHEKPXTpVx42fi60+b7j4qOHZMPXog03udGlI9
fztiy/exApiLyGqo9j3dPXgBpJYwxKrUXUVXthsZDQN35jBTezw+c+k+jUTvuvB4a63I76TOtMWe
yEAsbU/AjzARsFxZQllZ7ri9SCLTxjYqQqZJ+dHNxQ0ojOXV7aZI1rlBymxbpwKIJoEJcGyHdsY3
XeuGoB9+TP4ZvqYzOEdKTjH/W+FIRzrb/gtQGoBnDs9op6iPYRujJL8CEVttsM4ngfYSTgG4xMGd
+BdzbryIR1l8G2yB4p25OzqxGZbtutZc2H4CTTG9kcyhsjsr9aEt3lROuRULbXR2tkMJTR7ozsf6
ckMjcCqnlpYX/LeNmivg4Xx5xt2OsTnYVCEwIi5ITLvHHlg3KUEFxLtaTTG6lmXdLVrgp2yTAcW5
Nd8+u8CI/TtqZQsJzBVgD7AxXQzstyLNoIlxRXhGz5bnlm8wGZxXYkce8467FNvgNnp+7vauHP3G
N+2B9iLxcPcLnYZBNdqmGWPQWs2FxaOv91NlybwjKER/xRX8aQh825N/9iBf4WJd4JaFP8J+JZJp
cQAbm35CgCK7x1L3wjsIYYbk4urNlHBbIjFe4+KkC19are+x4R28nqlOVvKL0eSpgYc1c63qiMbc
X5MgyfnxqCQSv56BqhF80F5TZb8N+BLUIf0xgrCnIcfJrZhvsCt5CPGl2zJ5fYoOaaBo5bjmqdeE
tZJNfGXcv2ssJOTyUffP62fiiZAfLGFPjum1gkobpzkjQV8/GiRaIJk7xcPYPYJV2PQ/w3g3M27s
CSz5+cVH9fShilf2gPnIC+GPZ5jlZFxawn0EK0Ey91VerwLOiPMY/H+NtCnEypp8j/PlQo6eAGRU
mXgNccPM5pVrAorg4a1DjnYH8lcnzldBIbBTbRk7OWT9+iKqpdWMzTSBFKMtfD+edlLZIbz1khcw
d+r8/RB52cu9ZBYKKKeNM2ihIoiNV0pKAU++dYMJjuZ0oDZ1E4c9By8xzMKoel6B2l1N9/GOM1K/
2cTFq54EYdJvYEZG6yFAMR22RTkTWqYCcOk0E0zD2cnmAtLi3DPicVKKSCliRjNffiqtPi/twf6i
wa0fNyK2qT0/n/xn31cqx3WNQWSSZCjpSdHczMN+e4AD/2+iXqh2fz07pP2ylgmwhZh56h3Zdin1
B353ZhB3/Y7vw21zVOS5Q0UTNzIfy+HjPgF2KvLlgROja0nEEaYByiZ3wajbhE0qQs8pcw63TG7p
s0fYq+NMZOff3vReKXn7qb8yk917ejFH8SDV2y9McrwwOcKnXc2g3WDF+CbVAFYIij8SwhL2chko
O9gtW21T17HzemJgDoM7/opaKuM4qQd4igNNN9bEtVygM8iJHuWMv5WMN0FKnJLTazSctwdwtT0Q
enRt7L7U84IrN2BdSBkh9yOykd+6qseCKiKlLAYN8MW9r7OtKKM6G8xt10kR5+jE39ifcITHgYaI
s8VvntMdXgT1mssbz3elMXzBQdK5d8sEiK/cVssaQaG5seSpF2VkfrZTjw8YbfaVlbmDsNDg2/T9
JyfNzrdN7LacvglsGZnP5FtPd4bZhi0TD9xORoeVk2arCK5+Nl0M/DbeE4tCQGn/LzkrhbxAK7Nz
2+Rju0eSPci3k01RH8o+p50eRxPx478ML51QdZ5OIYWoP/PL7pL+AQNa9DZzIuQO8XgBQ92iOrMf
iGE6FbYekE2oqk6jgjER4agJY+cWX0Myf8ZOA170FJdza23lMEIJ8yHvLJmzclHfF3U+BWTt9U3F
/7qNW8TXFnDeuWl8tTBeJagUGYfhXf7nxRGjJAGsCPLpD+KdSxc1Bz37G8paocwjPjaUs+oa/Vqz
yqEW3uygR6e9H/X4KLBSdnDONDAJMbeBubWSe0hdziJIEyQpUMObiSFncf+goEXnLXOdN7dBDGEK
KPd3WIVdkH6/9ItaRrDC95XS2Cuqmv8vAi0ZwKqn0aD5YDRMEvjmEtbLEqI6b3EoOLbvUyT/aebU
YmTshYRkKQ/bHAGmtX7GtGpVOyxUyCkwXf+6q0Z1JCYme9iz2mxyjGWXi/msOuWGWrKUcubcaP1R
kXblU1+zhmBJTR4HiirWarVBeEBQQoIOyG2hoB8lYAWyvOCOJMG7T2ndHxb9tCOFlaDZ0z+axzIZ
MC2niFbErFKgCAYnJkm/P3kEFP5VUfwM3sH0ilyFhfXf1Us88Zd4Tvf9FC+9HxsnofVLbBEdQDqk
QkVGb2xftHayD3LLveUpZ9y/sxyLAAkwEzNsTng1B9S1tLhCk5EpU+yPONVAHahLJdQbaNDdC9KG
MpbY/iaH6EE0fwnivd5qeqa1lluF3q+MgCXNkqSjssTUiA+rGAdtYcKIHTNwskEODMvdxCdcYHXQ
SmfIVreemZrvYSQp50iAg9llTXkWB0IeR/Xo0kw04QPf8um7pT19HUaEOg/ET6/FLjzEvOGdsMN6
a3+zWBmywJ6vztv/n8OVDu98vkpkONSM5pKzwwDUIrjlLHrUdtgXQu3rq7b0TfxX9faKS01K894e
4h1d5sJHN/SoNGyWvgz/MonUC9/9wJHSwYY/DUpzrSWXNlFSAQsBsa2/RMKpVUWmO1qKoFaXGmPW
XZA+ErZ5ug7tcl8twWT4Lm1A/sBep9+LLj/1JeHd4ZSJhmzAv9kIx5jaG7DkT46edg0LYoVdbIfs
5LpvdiVfVUXwjuG/jiMAu7YfB5L4uHSl9RtQyi5E0zij7H5QQPBuIEXbncLj4A4tML6iRXUpJrsM
6k7H9qUjKu6Xhw7EYVTVGp1w6+3CLhYXd0VeSH+sOCZmU9/yfDtKCzKELtS//iNWu6LafzV6fhQr
Dtna/7/pzCeCW+N+APDlxFzIrt2uO8Vpc0NLeb17Qc5w1vzkwWwNpAnWYgG6sKtUMvbBCsJU2PgB
lRx8rOg1nd9Sk34VAyTyF26KluDTLYF2IFNW2QSm2AiAgFLkxyz1qnOdVzTyy9rUMDIQAsksW/Zy
6QQ01CNrhLcBg23E4kRTzLMXM3Z/IrJmkN2/xoaaD3Z6C9AMEBXQULQqy4rpTM+XpiBPF6MfD9E5
n14++Hq/+QGthR/jXKGsrZwFk4+8jxuv1aiZRjQECQfArPH7Kaz+41k2kNRyVlsmLDwUi5dJmVA4
3rpuPtaFWsuARhJ+srjpKG6zNj0ENKLUqsY/PpSW3yFjJiKbWCOR7E2zFz9JVZ/kiLGfUz3G/osc
DDvFAnzhUekRL2bzg04ilLUeJulzNmwhCW/cHezBIBDN9kEVeaqrP4ly7AvKJsLnFfnTnQWoCoLR
c8l5OUlxc8ptLtR2bl1+a1YPbQkNW18VpA/WSeJKmIKSDRQvRkh9hhraBq721NiHcYmsZ13add9a
OuYo2F5vOOUT95AQ3X9VRNr6wspJjTjRgQQmQusmPJ2yPaeviZ3nr5ymYbzLelZVF3oLqnd+W4RS
93micMfyxn1A9AOcoGYezEQYTRRseBUWwmY9Gs77i8hoiqN62ZbF602hj4ZIm/0JPpYNTMDH4tSB
I4TSijLaqCqOXffi445L2hWr5Ssk+eViysAKL4Ku9zSp3O5tSuc58wPuz15oLkrXs8ZGq1yhOs77
JMzh+Ubcy6BvEErlOLK0m8eLjNPK6KpZhIosQ0O8HDRdrz3q5ABNpszMcjhblzLq5NXnrU9vtukD
THVyntBD+m+OVUp3EvbIeIRz0b2dWjV/3yf8HU2bH5sQYZqX9vb3Pw2YkXYs7NvTh608vD8uA/fa
cwbUhtDtGKRc+kDISAa3MZdgia+hL+Nh0401xXMS+QjAvDk5UHJbeOn9Kb+DmI1JMnTD/LKOgpOM
87/+cZsd1p7iuH/0mt+F0kWhk2b9oUBAM+ilSPxH64RhDg/otaA+KQltJ88lukd+8HJJnJS+lBPn
D4FoErquSlfz9lWXLe2wAtDnmRj5i6n/m5R+HVKd2UjQQtu2VYz/fe3UW9W0aZft4sOEjBLrogaR
2n0GlnGowXXdebOgT3flWqVtX+aOZouSObPxf77MHuIm/cNzbgK1XsuSBECybMJZs8fdAhYxm1lt
6b5nbzCuxn6BUe3XlUW0fKkv5mql6ksV73qwiHVnQwRHFoOvjdaSQqFaYaRQ6LupEsTRsIgf5mma
2/KnPMI58LCklKTEAMeyzkF5hwN5CLRFW6N2t62yTARUzM514eOG6XCRh48vK9yaejx7O1EKfS+S
yYb0JrWbFpMX/W1TXmCDFhgippiGh4NXLi9Oi2NvZd9pX1gunrEGBWp4lXm5ZngxMXinYZWArEsN
HqwRBQRharzAb0g7SMAeryPOPKDgB3YRE+CTYsIFKXIHZhYJJHPhfzXQG9XKJmsZw/eYB2GV3skZ
j+4T9wC9d+uuI/3Sifz2/EjIH4pqhzDT6u2VoSx9dL7cJOtnlh/iffujQNwEcXHWNA+n6dCoT3UB
ariUL1TQm5rX5o+PZNT5xEK39sVRWgcEpftjAXrdFRbSjKFCzxaLVXM2H2aLIcwkJpae48KGNt2r
fbrXUz1uMZIpAR5ubgtPBu5sL2o9DYQpLTKFdmJpbcoavfZf1pkUN3zfws8UlsgwFZMSfHWEUyNh
ABdzU3N90IKUjo4hphYdJm18hdQjrAGCz97aur72dIzSJOndczfHbAV6YRt1BPQad0igfbvVHOmJ
rxOr0DWxmyjkwbIs9+N0jy4GZtrojRSJkSoIGud7Qh+H9I9wp2autBQ5xGVi+8+cNHllSnFFDDe2
dTiwFw9Klon14VWup/mVJWeIEEzbzcs5IxSi6+580pJKaJKrVGHcmVkwqTxpQCxjrUbGyyUAF0NL
D+o/ns/3ZB/p56nNRka9ZP41qRV5pdCVDVBEwG/U4G+OPNtCUtpdAwnrUbKAJDjHLD7inFcL+kt3
CE4JGnwFtVcw9lq7gb4LWe/b68YEw4wEGadd7Ijy9jcPMPnWv2XetQ8Xndgq6dp3gDdFdbURWiCH
nPPPB3Dva/moj7hyAy6ZRtfQFALwKcNmfIzfbNKd7Vl5ha7xRRw/MmY4Og6LYQMfLVThb+gdfFCX
mLtfbVKEY+fKTHv6zAWtx7H+eajclPnV6Va5x0MdMTIaDfTdDYGoCSKTFTIYEa9djIamdbuBU+WD
sxLyRYYbp6i2q9xeAi/WkQhsD9h7IJ+4cgsLUVZtTOSOKs3fCUFj1u/6ALKoZ6jbnRVUdihbMwc9
4SdFpVsqCWVgBRT+DemIw2GbzP28DSn3pL9D/9aIUo5EPyu0bhoG6wOvs1dQGuA3zofF5C2swjNl
8AUqhTMdujImhBIlMmeCHf+4VhSreC8tzggr3pmtwrwts3BWb27qDFxwTiq+S9/vOW1VWXs/Iqtp
8N0Hrmom+ARX/bIsnqnhXTBvChekkaY5SLq2LbyjHeVG+5RH1t0jEDxn0EybkxNLaZB+T9jkhhhD
w2zAHImURMPAyHlHrlLYImJalxonlavdeZV8I3hKjQvI71TfkHuVZ2dnf6cwYBZDJi2JX/nV9YZh
uGKMWPCZgvqSTfPc2CwN4YrNOhwrnT2nJG0IbgRX0wR1N/iAy5tSX7a7CxyX3Lqo+9tQ0DKN6bF1
n3bXFeP35smf/v0UxHipzx7zCkXDYtvHaUycHc6w+aFBVzvCiM1nMAhQd7JD77DyThUqrLWYnwqx
S7damUlJeVAGJBjA+RLjCZrSFyQuKbUJospoGSL2H0vLynedGn+T1OyJRpjhxqI0FD7VBDLWsvIt
XSejHAFC4CVPRmYeMKTkScmfaHsas/KXeZZLBIj7k2LaNO1nEr447B6soBWKkTCyDFxxk4SAn3o+
2tg9frNxbX1u+Vq+ALVPDZ/C6oQsN+OGcttl9G5vMDNtHkzu/qsbmmTiSI25WjxIBg5UCrTf0hHp
t7PNRPhBtAOK3BidNdknm809XzmKyzyyxA7S3S7GgQ3NAshi6ek41zV0NurRLRwq+ayqUqAF2MSV
64/dH3QiMAQtHeXP6A8rTz/JyqbSo2xNzl54jISJ4bHqIk62pv5T3zLFtkYiq/IPPEHO9GUNVcuQ
S87qgCpwENBGBsqAALvvoQEKDX47MSIByIUXhFBIW12f4kQR5uAoz1qGUxBqwpQMqG/8KXQ68Mw2
f1Q3Zk/skQfJNDTkIqj/f+KGKsb+b4GdUZhWDyYSpJO04O9R1JISLrM7x1ybyOgoVQGq1KUNmFlR
8t5Hss10TllokNP8jJr2B/uuYb34VXBgDsOdRSzACtrl8NAMdGs2jt+ZfHDl71oWE1Dy4XckzPuh
yOB930XkbeJxomSbSGAVkCpESXmirpRmq7F2pGamoDBCv5VXn1ZsPgWtL/mkt7Wm/UZWtm6fL3sR
A7q/HHivBXtPgFBqV96vg7RcU8RXOPaHsFg8dPXIJ105jRNB+8hJ4clI/ayrRURTbzYCQhnPElvl
Waq6ICB6z7e3aCD8GYyvE1bkpw0t1YJMzWYGR7GVaTlzKV37MPl4ELUOVrMgCvQyN4uDgu3RnFS/
GaFp//16AdSrobcX0YViMUyNnHlgHRrg4gT0TROcNTMbKxMLt2615IunwXgNH8zWlEMFAGTEyUfM
6yW74UX3a04QKxdv/wF/0mjFzPStfYuTQ/i5CxJH3NX6KVnj0tjbgLDhgsAREF3MIttYj3QKReWW
jUFFgWar/s0qhNCmWfidVjkm573TTGMcaY+BfoV3GRQivzyXOEw5oBLZdWncOXFnSxgiHIaX0etz
aeVNugSvh9nkltvGrgOd7WkDbtDpdA/tju2aISVJtP7zL1t1UwyHvr9aqRdCrj6OaQxJnZ7IEQ4P
24YK6yP7Ana8jPY+Rv21zN2qSgEbpApuRTMZxJ2KgCfLQ0tKZVo2JwHOmvAZWKbumo2fkAc5wudr
pcvJWbTcgpbiE+HPOR6nxVPVLZeqdgudaYGbz3pdKI7BrAbjofEFcYP2bZFhJizsPZCBl+THWOgl
9R7VHNXQ71xm/KN+fsGfA8jl39frDVHkoQKVWu2jsOABvNOuuv+j1zZgoFllfMVmUUHgnBaXtcO5
tDrvZYOUEyqT02gMGOxwUQu2rOCa38vp1iSR3iej5JHX3iWkBvwHaTC8pgvNezyBoP5oXhZydCnb
ApGim3/OUsgAwk/rUY7ONCq0PF7Nv1zOL0tPWM9F/bwXJhtCIACY9tv+/1aKeEswRKUzOUrXn/4W
U8mWrLn0owKPyI55o0NcsD3W6l7K841i8Z8UtW5Fu9gM1RpkeC9fpavL/gmZU81vP3VmfvgcR6NO
CJZXUZf+CZ1g7W6yBJkcdKztsD6ZExbuxIIA7c3kau9/Nq1H6lTnmIjgtA+GTEWGIzA+kIe3VsHx
JCQg44Ps1qTggLNM2PYtrBxBAEIxwHbshUpUkc0sTqMbHhGxsiOrHJ4jkxKiPOfHSCOFhE3vJmRj
4fEajuhSRV58yF2Hhxkm5lRHHaSXIqoHUQQpFWAVoZ/cAUbgTwEStql4bnozdXoSBD1fhkGyBxoj
HSCO8fpHSUfpP2JNpEsCugQ5gNGYnMctH2Ce0kp1mmjuzpCDeCGUQcsJCVkPl/QVWRzYKpRmXPyO
lho9V1cPI3RO4uByNRVS1ExWZ2pdckX+f0lHLWkU3A21R5j9+MrO1ANVhne3Hlq9u/16c9PONkmP
+fgqH/dVhZ90dedzAIPzkoWF9ssnAnC6Vk66LlQJRzilJnnCBsBnRLCHmi8Q9U8/jzW5AkpxYp70
NWikxwdnCR0GfNP73Sm0K69HCXeiOmQqTtwdD9Y/2RO+hdLpY44C5lSl1chWvmnTmRCMKa+X0QHB
IcKuDW7Qju2YkCWgNl8Vgm8yR4tMkvYZHmRn2FZcekZH51Q14ObfI2xzbpUIYAg1Yy4QsDTm4itI
8jJCkqQsYvISSstac76AOHtovplybEHRC3+OnKPpTAc9/Et2PcbrvBFDhLJhzh1LTjrNDYTOtfjQ
dktcoWLU037A1cGNEaj7JgMrjOlbYt8f4iqEDGCtsj74g04B5pY191EOkmR07dJKd2vC7p2W2Fku
TVQJLwDh3+zzzT1RbJQqRMhLtF1KYmzB1wsvmIdvEiJYxRmJpzRn8JusPooZNKBFGHh1xPbX3qhz
B5wt6i8MTyi3DRf8vssPBbIaINfkkqdpcaPqV5+NeTrJIRy8++rg0pfb37O98SINjn4hhj1M5sLL
yylNJhqNaO6Bm63JFI67fanxeMTdC+8VG2UbyDcSdGpgibyIxUTKH40vDQrAFfTNaMRbClsojmQm
uOO5Z8opfQQHaxYFPsxFcmndRiA3UiH50x0roo0qX8gC7xEiyKtqqG4R2ITZRFx46f84ryThk7Sh
Vfw5NckzB86nHPph/4tgQFYytiIPh8t5hrHlke+xxVhFNOA2mx4t9qkLbfir4alhPJ/iIJ7HU+I3
yfSZq1ruaiHcEb4jA9andEXmtUpykQiuQlNNjX62zcahqhfEH30q33e/r5X5Rd3R+gT4E5iwd1mF
XKGcySDtFeoRJhZkBtV9FI2j5ksCiWH1A9CSWx7qqjjc7ngQNxUQJrPthdRnDJoPvietb20T+s9s
MyJkxkCeSukxQicAbapyYrI0D+IIUESDbPbkkWA6aYOS1QfvJA/7tYNvwlDopKlJm0cE4GyAqa2U
Wc/OGx/FhqK+tLZP85u3jCCIgwhT8RLbRPhk0DU88y8HtgezxJ2MC/moGBXa3BfaRkT8wvHOz/k9
KasWE1d6R/8Xvye9M3Vqx2Q/xLmn/r/NSQGHwqhrWYYBd406d4x1ntrkFZNUaEj4JBBdb3G35igM
fMdOyagl4lw0rRstYT//vOuxTdWcveBTZtY9W7LMQO2HTuagRBIePTGAWtNeYL7BqTgugY71Kfkl
92Xx1k0jcN8lR1fm4JbYG1GjV6MQzT5cVovezbUTTevr6fO5Lv+qvBja4SY3IWtfRTzCHtoWFVLl
6ZUElMjRROyAb8I0ZT7Z5aCRaVJCIt/8mi3QAAmJHt2LTbH9nJJCni6yDHe1OtG6Dm/uJQhCcTwk
R492OcwU1/0Sa3rwVFr4KYaJAPSBTaZVKIgpXZtgvNAfYFC5KAx4QxhRRYEirHUnhaFWpaf7I6DN
GqcDOgJhHx+s1AJRbh73CB68joxsARrHVm/KlHGnjEktp42k8vZ/zIJixvxJFTDWXu5xzPOFYWZm
LWfdAgvNpraBf/3PL/9IFIb4Tby/metbyjMMOM4Yj1xaqJCFoMRdpaE5kR6MbaHsDJ+cAJdF70oe
6YyqzT2IiI6/MrZ+zPaC9bZkYRggFQun5du92rNZDSfYCw/Z05BwsweAPNFHmpb9abfDgWxW0oUw
Jm05Tn6RvG4CaPdnAL5LQf5bVw/wYkPMe4CoDRDMr4LWpMy/Jc2q8XrKJMbii8YBifRk6xoy14hU
liiMlqVuK3ZY5OMhD2fZb5zZsWSL8cA/N3SCnJ8Np44uLZCT/LWI8O77drYKVdzQfJkzgbutw9gm
WwZxgKs1tMgfEmovs2Z8xWjUPMtQ1TDln/ZBv9h2PZZ7YVGTDCgtS/vWZp0l8U5IAp4JVs2plVAa
pKuCzjl/HkIove/RE2aR21EBrHUqbrQZ/SPnX5LNbXb2xmhy5LM09zCEoWh784PWobAeZcuGgWEP
vQ1EXZt5kuGMm9bfEfYH6c8n7NAwr61/100ujAhla1+Os6G2XFykd1ycN80sOcTNcoArXaYSvIol
5oLbBX8p9rWvf1uJVc13U/jCQL0T+mfSQOx/QaT6j1LtNKmZQWLDDkLinydQNgzc0jPty++58cyp
+ZOjYZaxUD/ldvYwlNOLZvMSH7KHZR7AkFg/Yt0nETqbQFMbkUjT3JnVYbvj/h0jcmsDwzJ8QcA0
4fMlua3LVC+FDXJ/4VFNv2MMOu3GBwOgtH+hCjjc39U4ojuC9YGYQkm7aZMafPtdQf6jycT6Ut4U
WxIcH0/yOkwzHSda2dvtecVVkhX9sayOKJ3KnaD1mL/WiMZowf3sYPv8NQa4EVMRrVaO9ncdO6fg
4DYnR+NX+IenxoT2KvFzRjdzEXN3nlsApB1wJ2ca9m614Xwl9hiNre859qi35Bl6MpSpvdZJNRA0
O4/vlAd6fN3mPPxwpM1PsYxBpRnOXpFjLfJZ6Rj2K8zYLhfxaguaFI78Kr8sNumpFpOi4RXpLmwn
8rtrzmuesbOIr6xlXVwRo4t91MLve9+3WwofoYiUNP49wsDMJtdltUVcA17L43tbzdZ/UJbP9yuD
TOyk7UkhDSJV4qwCcIxZ5rRMd3FsL/uoGUIeVCbJNVG58BQ2zbF2f4CEbhmXXed5bS8QV9gG9E1h
ZiuSSkwtmgrNqq3f5Dls2A+l9MY/k/IP0hC0kFXcGFPs+CTon8AUOuModmpj2N9wjuNpEfFDYWsv
uiHFEarsiysCytTbu3cLzlBDgHlp8BlpffWDePZfJJ4tIssUkzqs6yP0GyTlLszn5BxpBZqcxyp0
tJ6Ir1Wot0ENAVDlNBJTdFtTy7QFEv7nuz2MfmFekfJYJ51JMqNa7Cd2d9fQBLB2LDKEj0bdhu0U
VsRGtQb6PcfeBp4hWxSs2vy/v6Y+JdJ645gx+CKzyOS3Bv73+e+tnA5Bah7sMaOhQX4YJFxNMWkC
7z2ffUS4k9OUwXNvVd2lU0ThsaxD3oXDSXqfo/Z07mCenGXJ7MRnot3oXQKO28zOLFjpoTsRg7Y1
+ADsN8SBTMkViA7Liu4oXUxwa+21LCDRByFzsRXcGRdjL1E2kJWMnSkgpFGlv5geuA6BnSQEBBbB
0fSTayKXK/pfKjhT6iG8ObzMSdrRoV3DTzcgEnVdJL11E+ge8kdBO5nb5DVXRUd5cOKLbGf7Bxrt
7IoKQicNzAHTNs9TqyfszWarIo5on/yixzrvFpf5N7IcQ402l9mtYzUZOC4M4XQzMoeoT6dzpiSK
TOCztaCJOmppddliJc0wVjoehfdiXmuimSLu+ew6AcvulfzV7GdTrv8qBTVgfQeI0ZHhZIaEFx5Y
hRA3ffDLMbG4R6HCeCP3spqyZ5eqlAsY5gZab3g5Ad5TtKa8u2+uXplAMiIdcBGMMJFO371t/taP
PdqlUnaBP0hD8lN3ZWjRbRm5nVmJ0XrRT+8UsiEHjjTT0y93Z2nMeSkg+WGtgIFXXpD6DOzg2ZFC
0iVM6KTN25CeZDIipdqGBqinzNVNfXesRIDw8HJTkrdXrsS+zGVL4wboNpURYJ/pX3JkkdHUodmo
hkW0joVNX/tRQUtd1XpO8tYI5cN8SsaDUjFIEYanjRZQuBwarnSR6xWa8yNPke/Gc2TwlTdqrRys
gcHQzUPk5iCNbVnRxjMwHucX52e+0nTDztBU18ne39SV2omT2nv76yJvo8gJ3eAkM+99i9lW+rKq
NXgj6SJShPNERLr7Ln53ffR03aHP7VLIn6Un4OK+pOGmJN71eSzhCYFn22w4kDidtWoZmieCRaa1
VCUsJ/4DvMnil/3y9a+K78mg69zoKFhLxJrcoTSahEnrwlEak9EuAaVvW4/dxsBy7/oalVWz9ISg
l8oLJW6lFsDvZjGeeYYfr5F02ZaR7woJnF0Y7EJuAeK7+Y/c6W0QoFJG+B+MHtVjM92NNxofhi/m
bfnTNcIQT5YmjgpUM5UGV5fTBv8IAVEcUFDWg0AnR7vqEv3JH+2g3WAAYM7OyG2HiYzNGWtIBu/7
dlwD7V5RmjA+oDOREMq09byNvg0/yqx2BjDK/O+s/Cezm+xNIdWc2egD7CLo4dglfqY/Mxns9xxi
TpwEc9lMp5j9s3+SEjWvyKo/p10AGSOQZnj0xENq6MV3MtUQ3C1yWS+Wa8LEANcdaaSBI8sI0GVD
TTpza+TubXknrWKgvDmSIKyNWZm+OJQm8pNW5b0avgG8x2T2ViRZy5eh3fgYniHsCKf3z0Hv5AfU
9PdLNO5Cuw2hAU513IvyiJSdn6PxBqwMrQbGmyZ1aMNTXHXv9sCd2wP4XSZ8k0HgdhWA11BRwOfj
rbqj+/DXYLXnVDz7AoO0HUxQ0KhQpCdVD6dzPl4ZRsjv9ibfL0LseVp/JwCS6RCoV+R4gE6HYy8g
bokTODVy1XONKbRqUhtguAsBedsTCMjU08SUPYmZg2wB4ZmUd85tTCFSk9gr/rPm5vtWj0rU4G6e
lFFv923nmHtsBtTZBeFDNY9Lawto4VfAz5i+WCUi2VmUGh1JQ1EM22sn3cj0QHo728mTHgtA2BFM
SntNgqX/K0+RJgcLd+zV0FJIVESx0Go6WUpUuR2Uj76IVpDgTccMf7dse/a/9/fOdctakOCQWNmu
Sm3avEyB+XbQtSb8v1q1cFN+iMOJNZswFtOOz1z5/GhNfHRe6NB6d/3txKmiv2wtQpqjYR5B9zix
kIcnbB7hyIxELL20UguQb82Yi5eW0mcNkTE+My8MH0VRhVZnWNltBuIlvxShSi0zNgWP9ImPqPEQ
Z6MRW/r2f7MdFCBVze29qZ2+yHLIw8WeAeWQUuJAt/mDhDF9U/SXyF7HvkcHBvgZrkYKw1SpkeyH
Y9mf5oET+iXBRtnznq2MExfwDD8QqGsXNxp4HY3hUvtInvKYYn07rGDqJlpwG13rF/AtPnH3tgw0
3Iv0kWx0pjhty2YyjWDmbwlF/zh7EeVTxFr1yClvMZ2h/vVjnVOBcPgsmRL8E4QxiF9OPfm9fH6y
YaevmhfpqtqUIQhsI0IfAz598yStZyarOGv32ixGcZPfjkoBLK/DcdzvlugFs1U28L3n2IOUxNa6
72GFgfwI+PdhgsjiE9BenS69rc5gWNCFy8wJHXrhAJycqj32OeMeBQkQpEsxRhvihxoP5XMfYBL7
bXgwwZwNK4I7rmRUO1OS/O1y/6Y7QS3P1YTM6JcaaXVGbL1857snDS/9FjYc90NI+z7m2o+lDOdq
xqNlk7sosGPZL+y4IzKY8k64cFYe0dDK2grlqmmJ51GbBsEN9nWQdroE91Q5OlguHi52aWfZ+5Y2
VCu1FojOzDCSQyu0y1jr5z7sdbWjx00MOSGrK3wGD+vTog2KMCR/KgSH/2J64GZfwVpuMidhj7cD
U9uEXg95nvKAweN/REq3jdATyqRk3YaNSgZmv69TOT/ipo+/o8d3ZVERyswNOvOeT6GE7s42KNR/
PKgQxNNo5ve7Fi73iU2ps0TxO8rxMHlBTp1ogVaMmCRJOEPgLLvmRD5S9O4825iaQfeS8+d8y74r
EyzwTiyOyNSsvY8WVyjfhZff80bA1uE7nbE+jvWFXvykx4kXudUKjYQYatsCN1Cu16TheZZlD9W/
ZEKckpBCxSDIyLigUBY+Tef0puOY3Z3693pTjziwDq6CyAZS/q2tX8uwp043TykzHLSggdz0f7yQ
UAgxCDRSO8w+w7dcnfYVD0jy7ykDgizZg21TjSd/4Wks1Z16fN4MzjPSed6cyH3+4B4eaYwjUVNy
/CtbF/CtY6o/Nryp+QcmiTNNnXrYiLu/wuqs2b5ybmddkAC6EOh0j2//Z6gbGNKEUU/LD1rscK/x
AY6CG3GjVtQprk9FZEWqVgNC4hlH3lCiJHHcbd4ntY43DLAjSzP5N+Y7ylAGa0jYGmVNj6t3J+dg
Gv0uGN5/XimMGlCGuh0E3s61UxPNAlo9ttiyG0Wn8s43/xD1B/wfGzh6qxx/lF8CVUfVnqVfBLQ1
6F+DwcCRbNl8l0NzBT9ehWORUTHPBGzV3kE++s25rDiYY1snoO9GvodOv3BTzPDaCpdALv3V8Kxg
0QE5Jeuw9POesNalIqYWIj3whCi4TQUePzx5/0yitqIxLWssJqT/IeO6oyWwzWv108hEO8oE9EGZ
7plQ2+kwkZHHVmUTm1Drbz9C0neVKzXGiTW6iO9hnMYTbZZeFmy4gxo73orsEGPVgkW6qXIB+WBv
5dgk0hySS5gxYyyDo6/S6S9UFhfqlad6Du9kToH+opzZFCY4ogpOIs6iyREwbYAjbE26pQJNvhzE
dgoBgP+jUmHS58+pId/h5AdWVpJC1X8J4OnTbd8w6wtec1ibpRlZpue3OddHbMKUZIGAWAWAxNhX
2oZiTCiOFNw2d35Xb0NkDr7WSUEwIXAoV2yS+6dw6utPAMDF2CsMlHznjRvIb93ysLQWczCyvWjj
LLV6mvv8de3PGcKRtRsQE8TJbYFaMTDOaFpyLBc+aRG7Z8s3upldxUlHXpNedTilb5HIr7RFMoQ5
XZogaCS4hyZ9U346patr5Q83/t/Nqb3NGM+TSzkyNZHGtwY8W1J110+3Vk5+Z+JhULgXLR9GufEv
PNTulmDTbD/Ml7GDeKn3QFGJeVwR/F4O5VzNB0jCYrpnE9rRFWPxFAL2OFrg8s+/OiH9V220a2Fg
xii6EIKieCKtWlnjlO+Ev5067MXk5yEW1fxaYgauJuNuMRwCZEloTQX/1nuv5QOk0pJR6pw3sol2
nv01ieSnPITcaDleT8PDXHs2uhMPs1o1gp22wvKPSkR6Ezxv7xq2DVSrVcg9/e0tRXCddglWhbtE
QEc2og51i0Rq+MndC88m6NLUbcdWYCVG/S4vMczbFJlxwpZAbylZslClM7p65DWKOcs0Lpx3PKjE
gMV1TED8c2Gm9iQlSvksRWoa/Ds/6cYKChvjLt3X0wouBX9it400gheaaaQCsck42C768WDpJCQT
EWx3DI7azsukHSK2HKEsQWPXc6C7SwtuW5xAyM8X20Uidp7o1RGSNEkW3Hz+XNMliJeLfNNe9vy7
COFA5/BJwIvEz2XfXkB+8b5//KH/zKj9tMYJn22e/hAiAmhCnac1yhKcqux5JlScUq1e2zHKyx8Y
hbNUzH1BUPhH1LPCZZNUmYZs/iu1ldggnTHJDX6bLNkrFEgJfVMcj4vvggmKrlwI+YYfm6JBXSlF
R+dC0i8gZWXHIPkFio1HKRH46SKmqSWeB8PENlMNJCpEJTpJMnirQeMr9NgKcdvCBnd9dYiRv2fO
FMdvnclEnJ2KeHsYxtOBTd5D5V1eFfb8yQUahB2/F6A/5lr/AAfB2L4RuQLEFmLXpw5n0mc1YWCz
nx28eZEzGV2VtzoAxH4gea6PTiqicYEYJE/zkpMBtrwUb3FUqz485463RKQs885n6TPUiy47pA0G
rkr+7ialD3T6ieEKyNEktr28UF45iMesI+zfiTmzK7XPFI9D+TihvWtKI/Tadpqp5HgJBoI/yAtx
uzUjZ2tffzTJJ6KyGoBYgL74ltBg5z/6kAJprWJa8Xsknul1KDRTNWdUqjv33SnwsopHT1QqX5et
YrvaHkijTxCl7RDR4jP4idq+DL+LBGUd+b+xkLdzmtxY3gJ7BWX5/J1zfcqORewGzm/2WmHgUW3i
qB3pg/iZPh8JOS9O6XtGVDiMOusYDPwx/8xIc4r7mxFEh0B/SJp5+zfMRpDUz5iSO/cbhWDpXA/U
LoPbyArc7HB7at+yx4YYk7T+OCcX0toHu9PCRI0z7kXX2mqoVkQ9cgF3QCFdYHaJpBrhIzjOoYv7
qnLXCa28amJXE7P/ivVAE4nUKtA32V4VzK+nkqUxLl3h2hee0K1SqRKTd5LXSKPC885hoBjoatvm
lDjhk8Dzq/GzZ3jkAeDFtAgB98MjEsncxhJe+VWljPP1gzqrGV+1cgcEIgxus/n76Ozp8heTUfJr
s44LohQi/V0E8o7loG8n6MZ2gTq/FX9NF7tD+TPrCnEdZ3K1b25ImobFRIlUuc7dyuSCB6gW+U7+
JF8yxHzhrTlycg1CuRJ6TpldEsRkSVrTIUsfUvnELcKX3ENJgfgA5avy37mA3jGmvOaEkCGA3eYu
JoFWIKX/9eFouiguNQOXSB4a3j0xdMaYAaniKrbH5xn5CSZalUY8a4aLifg+L97P9ist/dNOr+Kk
FreFECyBFUwPjk0QRmJUxBegr/wjsUezh+1KiSHukRkC+LSxG4gC4ZGXRJ0u1AmtwJlsxOaUyD1H
uynjeRTFw/94+/dr8XDrBJNbc7tlhTWbFFQTnNUVYmZr1SR7906Hwue5x13CK43ulDwxqHhU8J4+
cPUFGJri4SZh2xW4rfSIsfThvEEBfPiJbyGuK2EHVepi7qFDMXRbJGFToH8zfUjiM7sP9/+OaCyZ
gzPKBGGeclOfoPbZc7DeGHYV1zjFDjh5HU15dMfpoND7KEY7qYufqMMsD0N2yFPfBqmfTmx8oINk
IpvKd1mdHM7wwgXy14y7mA042etj7un8TJAGnJ6NN2TFORHHo/AZVFIyZlDTWSoDEDNkTjKaA6EX
OWqCGG0nhVW+PR/y2+RBj+Nm7VBGUMzVA2eXC6CHBU5++5bISxE4R0rk0a4CQDGVeqm57y3nO1P5
aO+uFFnowJoDu/LvnmrJ8ms93czXkRPJR6tCc0cWLsK1OQTXdS8fcGZAXzyIOZK7zeUZp11I3p4n
iAUjym+7a9arUxLg9EnhkijG1xfciAW7zpnlWKTpjj723ijypPV07x4yGSY2ao4PxctR5dXIKynm
WTjwPYrdCUqS++vDYMmLNMq6u2u7Ic8iSEHCojDGZ1GegdakVTe9oqoKHeUivCH9JcgmIUN/Dl+5
77Ub5LahUPyDkJeALIQNFJyjxtGOzdNc9YSnoCEf3C+3YWngkpWWYHJETzXTDM0cVExvZZh/VaA0
BjjwSCLMan4eEPx0O3v9qo/11bgrKg5OgfmR3u+RkSv1e7i7UVT8I6kLL/m76ElQTKKcpRVSLRT7
mHWcE0ynFbcsqu1FbJINiG9ck2Erfo6BmUF5Vw6tdtZ4grMpJC6ftmC7sPJ5vVg7QE7r2DxfXggl
kkohytAi/iU4XWewxlSiUQlfmPrwTMWjv2fXVacT4RhFcYkj6Xg/9gKsGECseRy1OA/bGRPwySta
xdzFFYW3ib8MfOPPxPjw+jwNwcu5qJy+/yOYct+D1tysIqCzFahW1RhrcvlklYMxS0ku9rGpZgEz
GrGGnR4Gb4dqQG+LN2fXth4dd1FwUMMhQTMpOvK2knJe/T1A7tqsLYvQMqu6XsR4fHHZuWWzihUM
kZnF2DJl3eRqKCaGXqSPiwsB1KrMPVQAChPrDVs0osLiBTyibFkynN/1Tf6L0vEpxAmsOR4JwQkx
zkpMVDsG2zZ1rokzKsdyB97SDCgTHGWkiNXm7EQAKLKRaM4ygyJ2WXzi1g8FzBSRQL2xp0EJdT9S
BWmHsnjz36P7v+1RxPu+5okCg8ZJ/jKk+p9+iH1MBxTE/oorJDFF+rH+R3QidFYvAClyV+JjN9GO
5iyocQN2nlD9o5K2F54+7isxExZWeqz8RcylIelClFd4bdcmnik6TNcpM1hHu4pYHJWQVqZyI7la
hXEI5JTJvWQGxKT2dt5UdjreHKsJ3s95+SrlO7tb8Y++1p7k13NH6CbNXcTUnzyDrd6wbD0Kc7Cw
lk9mxP2Tx3CuwEZ4uy6mSsP21s4XbXyGIrVw4w9ClPC270mZc6feiD+CpBnP5g3Ty7NO7br7UPjH
XV2T2L29wNymXViu+T/u8zbKmIXvMo1WKKj1GTDGPruHXOhY6GnyB90kleRCGoBsza4NBisIiPcy
qB0H5c3x3SP+LWSk+ldjjygx2skrdZtlQSWJDUf+x96yFB6jRaf7cmexFd3lLGkfTh/ixlsMZ5W4
t2bs4HElBMp22FtAw0TK2+UYgFvHbZZ+QjASbEhFE/RJW7h1OkuMQwY3esv/K7JIP3PF2NAbk0Om
ZzzCGjcp51DQK9QEMVWybBpiMJE7bBN1hcAo9kf7BMLhxa+vcs+m4Aif4V0KE14mC2FxSe5YGGgy
jK4An29DXKhVa+g5bkpxWrG3ziDF3uF5GOEz56fAF6Gmq0fgCPzQKTwSEI9sT7Sif5rLy0gnWrf+
75+H8CaxusO1kTbgs74ASzhQgvC9nkHrXZpRpvjISx/S6HCkTIA4V948vSKHtX6qtndv/VlHOzLi
jcXWlHUkLuyJzOdtS8zyw2DnAkRP1CSmuH4SDGidxejFdS8zc6hQO6uKmP/FALW+4DDtd5RHWZWO
/acYR1rGtbJsYstEL2irqBvcBiSahNes2ir9a9wStCyZQwjgi1KE52AjUnR7lo7k/65V/yskORls
yg4nXFHvdD1d4osjgiEXu1Ha0GhJ2xKWIN6hub9tmWVd7VZxtiPb1zAuVI/ClAS8VJS/uqOlERVi
UMPLw7NztzJzvwyJAV6S17HIEXnF5hx7PdMZcxtSGHzLO8ptq96Ek3J6H9dW72yq+vXS8Kysck6m
ESTZQ72i2bFW2KVLFOFBd/aSJ6lH8XmrzG8O1krnVbEepE6KXITO0ko07iq8C3hP5qF805zQu885
sY0RZIMhmHmfTRCyJ8MJC0QjUWKSpes8IMhjj7hQhp3pXL3WHVVHDMb1vs82XWqSTOGmWos3dh5r
9qVMgvnWkhJo0yI4/+o002QPk429x1hk4qh80sCmFNKffV/Zbt7erZhQXEslxjcQcUPKXSq3qZYN
0Fi9jPnfVdeS2G1wvzKCVZ7ovwynJfA6ZgyqkEQkBm8I/0jwUNe3gZpMQM9pFJcS25sWmpATLhNR
ywKcwjw419ifkjzVNDl1vRB3gIsxF63cNTjNFZjy0xZtqtSj9J8DeXTBGAh+VzulZH5+peYyCF1X
5XCYwSmZtqupI2+/iFyy5zVEM4sDqEdqRXxRYcZ2T/0bRucvy1UWjW9Gp8GM40XMJubC1J0sUilC
+bb1oLVbO4W9jFr4x98olsKSXkEGCmRQxbDUN1IHZtNKZwrq8p+/+/kxNFStVC/H9mzqsQYHr3/b
iQuL83KZluB5pbTBZh5BevkUKGCbt4X/T+AfjzXojLxnijE9fHg1MVRjTb0GhLpYpmvL5XZs4liU
t2O3UzWnWtIgJbC6bkFpSDxYcOLvBpC/F0YOTJsY9VTU8jHW+iEm08Og8ZX3haAZ5IJFSEEN1Ul3
Pg5wu9cYJocx57xnCWNwhH6QZetP+G/8xRCsSWgXWp2LxT0EiJZN9v6uN+DgTT/npXwQ7biyMGBR
doGQgZZU2CLtpW40dsI2zCt/7PR6QcELEFd+neTP9PFGeP9GQ2dsFQrIKzbCTrbCviclZShZ+hlD
5yid0JEMd8VHiJrrEHTGsN3Ha6QW2d15X1jEytMa78Z+0UYjkLErJl0e2VwLA10zEkoEOXEQw9Nc
l85Jy6IC1znX9w0aWTu+jTTLWFNbdkdZrk9McsOzppZu9jqSdvO/hMhwR/rqLbCILn3tc3Obdo1X
CnnOo2EhUM65GBqL2vK2FMLJTxMFZ4sA7hQ0HT1/Q9uvu8fZuI6FrRASxrCDStW/VKkXWtAD6wgz
TOZE96FbYYbWpXpthsqp+xConneo4jYdZb8fLhCV+1u/4nSpNyIS6JmwQS6CzA+BWfBjYdRY9npc
y1JbKICIKe60CYK/1Ag7M9SE7rRFpc7tSlYvY4Uc5LIReULZrQehfdhJ+xVdQKKKR7FjlJLQViHq
JU1tKUqX5B4JVoHadZok8wE6iIIbGsOPJDbq8r4Qcw1WWKguGJFGYcPqfT6O3Yn3H2DazTtdrzAB
s8miIi+ryDtpxj74K2pt+YB7tNZWdh8AgFIwVERec8jc6e1Qv7UQ784vzdb/VRkWLohh2aYgxFMQ
JEIPEQLySO1zJ406KPiaJkO5nScYZ4Jrm9swJV7PRZMA2/HUOYV6+KFQ5iNrRwbEC1MRFI8io0uO
NbcDq3OHoBlejG7pJyh7KdJfh7+gXhEXQGiYGg+84ZXdDOLbyEVQ+Wak9u47xvoVd7DDVggoZ6f6
pNReAby1cYZopHuB4WLF02YVCxL67+o2+B8HA6L5E9z4rKpi1EviNtx/PmilEGLSBXJ3P5bVqmu1
cjHt0/biXaABEGepFMf791CJfQNESf54US2ygtTaPnpsXfngFrKZzRG3qQqzyX5tIC0OE6ejXer4
Lf2O4b5HONc3QtvbDvdL3ks3XRbmSZbqfT+slZq0Xsr0Agn/McnuPemr/Y/TDU5X2TM/m+52GAa/
fp2Ori9eSMelDCjqX1JtKqBMMF+yU9D60Olk6PAD2SER1w2P1csqlxSaa5WyDjRtcDcDm3X2j4er
Ag2K6G/nqbOyVpvN5fjrfooPIvpn1II3xEshn7LidnTex0z1CKpbJEirONLQPKdS51zGQglZHgyl
/q2R1zU3SJ8ahCocUd0HsYmOitepeah0OJFM+G5MPIOKjHZ4Z4qFINb9jZB5YeMjv/bsboDFSWUZ
92xNwE7PioZrmJFo0eTm8Q2Lb2sADGNPikXm4n+fiKOx8YXN9PoEyqJEisjT1Y4FMhqgBL0RR4V8
S5MuGKeBADczss5w6ZFe1FL+BTtmdNlyG3v+qICA3VCEjSsCwjA4wro2Ik78iRKrlfknAqo2exzr
/BXqKDgvYFvxC3oyJrhQsrbLwiIKwuZA485EBpjmEV4V1g8moWAY2Uacmv6oCDPtUa7x0PS8h4l+
RjjAVAo/R8Z1e31GfV1D1cuN6W0op5r896xRCJKp0JkhjRBPXoOk1a8DezPsKJADl5dC92sjkQZ7
7ffUwr7zfku8wObisXAU7KY5VEVAW4zV3DZxE+Ms76bE+w3H9lmJKzka0RCkMsB020PQ9tLl19UY
EMxnA6fYJAzOOXtNFYBc2jtD5NhOi4QZao966XBq/A6/KI7NXYI0/NQo0BT5kjzl8UHANJfP67fd
TPmpr1et6auG+1jwRHBzNcFMwF/SpKmThyX6sYwLnPbvySuqQOummPggNDkKEXWoawL1OueNksbK
Ql+9RGxz9O6DATq/6YN5E78hQDvSB21C6iEiG/44uHRbNLl5p9GUFfOZcy8CUN7U/niVeTnPeBoh
a6onqGzV9s/aUcdDvxkXsHWPhVUwsoK9ENfJpgt68Ydjj0W2/OsTwmb3veYrrns/U549H3pTU8+c
TOAHFaUD4oNoGIAbJIgBN8OTZFJ7yFHbNQBxMBNDB44Q3SN/0zpi1cfEPF80Yru2SlU5nHbNZXss
iUd5oOJl7pX1WVWecBhjvTwPUaGO8QB+GMJNpjQaXpaWwglYe5fRkF3omQQdt4gf8oeJpei4zeec
W/rGQeOHiFrMXmxuEsw0DuBAGorD+8VFCKtczmEha3AMXvKXSsKy1kxNfQeTDbXoq7DA2AMLg2Hn
HDZjx41TxWkutuPPornk7WyEftBuRjY4hOapbJDOc0HaD2mrMNOtAr6F9xkDly+cPRiiqeDa4GtV
xcfMtov4e+SeWPVyjT8cSjm8SqEjGchvcjXBacHeSQiKWWNtD78RizZYlPYb+Jp/vHeEo1qNEL5S
FHcnUyNe8gmQxrRPlCbjNTf5Q1VIyOOjH+A4LTiNQtFUr46pwKoVhOHoSYa3nHJaJia03Hi6T+ov
CsmgafOR9o90vKoUv2BAo1uaXyFhUy6/qXj4MDA6+5kAedgEWBr5kFmsz2A0v2/eFG9Kf4FXoy9o
KhH1cB1iGdQBLXroMIKOhhKs6I46IuHFGJBdFxr7niMUJ8Q0wMZserb90LMGCiZaUnJCB36f5eMB
nmUQS87TqVkExhNmEGUCsEaVmbGEuLFFlHo/oLK8PT89FBoCRIGevisoY7lrj6Yn1Fa8K83TEN45
keOS/yhqopeO/8Xj05zg8b5gCJWIsk2ORa8jqJXPIFPaF6qymkYMRcPLCitidiztHwbEDwMs3w+N
KsYsHQ+pf53tSU8Gtv57iBxFc2ytbcarw1S/sRc9BRD8dDWdtEIzgrpFEQg5PYZCOdMazHatz5GY
TAJ6pgElnSrUFz/JpRrUkhZUMFt9eoZxwQJyLoCoMO1YsU9MDBO6eEjPG7q5zNl2HlB4NE6I0YMq
Y4VK1mX+HCBaNwhhEQUjcpUzxjQwjrGOH+HlHxU8t7sXaOnCwqr+WGp2wZRbV/M6jCRpdsrK4cj8
e0xoIGWlHmWkappR+JVzar7pdysQtUGhQT9WEjyi15CTFb/CDPPwICeMKqtBjXIOnT0y+HmZx+Jj
5tN2O0aW1+yP6yB/WSoAO5VTcyxSyEUOQEhF7hHisbdfvTnqmQLAwjGqFgqFNy25X6xM0yFBsFJP
OYlmLLATp12OBQlEkAKCzwXiYd3tzVeipdHc28GaJgtiBrk2CYXXq6EG2p9PFPz+79Bga17Qyom+
ujm/C764gAX5ekXhJSYQxgQNQg7tB3CoD2AukseDXlW5rUl1hY1Mt60KUAtmEP+eBSlQVDKTNavx
DSbWBYtV/hLGbjaVpzNxFa1zOAytHvcXDoUX0njTKDyLRMem7ep+W0YcFkhDpmHVTjh9+DRQRaSd
ll0utfCi3DbHuOgMzGMnCJaWSI9P4gubduRdRy+7vX9UfP7+LaFqU4CbBZFb/FDfha6Q7jJUJ1yp
Ct3lm8a41YJsDYYOSum48Ts/o9pvuurlr4zAxNX6ERj9Q4vNpzfNlGP852BEWGQ3lgKvubfCPDka
cDqPwRXizjzJBdMqNx2sDyuVnRZA7t2B0K57CROtmQKw1jEl09xz/gyu1iUa880jzuPqVwjNJDQN
Ez8jMRcB4NYljdgKvXSx8TEW2aQDaAjzb7EPxoxEP/MiU7Iv1nOWPfoS59LKfPRqjd8K7OR2pkD4
xJT0vGv1RhRDLtBGpw98R/lLySjhlDxug3sTrkVkAsw1AmPiDazSeu69E212NSnd//vudRIazDc4
Gn3k7SObz1bXdxzC5MtPshhS0ChNotiDEEU7REWt41Fk1xUK9JpDokPYV/bQV780HGRxYvGBh/A6
UPVyKJGH4RbTmCN96zfFO0ClfOhMWqVqje2FtN6Q5GvkuozrCxV+GiGUrK64esR+qs88AZ0zCAkZ
6IW40ixm+5tLrlLu6ZxUC/Bil3Mw1rD/6FLYaUe5vh3lCyxNA8a0pDKbYYvHsfjEraLFrxixOUAB
1LkWMK2fYhiof/1FG9hI+PtG0QKh2tFh6k/Gp4zGIDdW4BMX+Uwox9o2f9WNB0K3JqK0Ipy+eEuD
dK1hX5arFyI6vp3dPEaY8EeUkZncgrrWxQa5M5EwHtHR75xIb4AuTexI6685XWWR8wrL2TnUttdm
jSijK51MK1QK7hJRDsDVUWu0cMlKDgGsdsiXj5KtWD5nM6HA3H+z1GecC9C3Mv1iC/mjEGhR9Fri
BMOKSSsGZj2ggTbIp0zoIl5y2fHJvlEke26gq7CULW02ReM4zQ/iSOYOa97t3m4G91nHGrx3iWd8
6KDlWzmOKhpN6d6XXL1Sduh3xL6z2h+86UljDv0BjxkWZq24HUT2U3ddQjcdMaerYmf0nibTUqZH
+4knZIpCPT3103vFFEQBs1h5W8g05oD+92f2fNqv6FjyX8XFmAxEIQfj5Ub0jFApWwSeFi16uuuY
G3AT7PHBmqldw3XTRzQTABVIfh+XTpCBZTZdcNzWojX08t0rr4va34vrcvXHehoSWC5BlT4ddSsG
88+YZe1VydoyOAqjRSz78en4qnbERTe5ZPlNA12+SBUvTN3XNDxF5LWEY3ADg6C3e3BBGHJ4jmDQ
ZPoi+qKwdpKgyuCiKWX67iBJDwLwpDS3zIDWNA+fF8/hOdzoECD3AlS6D7bGkSzHwi/zBtz3PY5s
deuaabWeJT8JHZYgBIW0E/jUms+u6VEIKYGNWRNm1jBm/zbo/GeS7rUMrT42+xosb7Eo4nLkUmrw
q6xfsS5/6fA4v62srMexAMqyxQ1K4f9GJVxC6zw+mDKbQBLVr1kGPk8lBhXCuNQnnQVCbd257VN4
xOUoIbl/GPeZk74I7V+gv73WiFiv6MyB915P8RIHdmjbr//EY2Fum+e007uOTyq6M25+K5axC7AB
HubJ2yuZpqhOTb8o0AIAXo6eSsLLxJ/7oUyAXHb5z0r8oaSXjoUhIvJbVmn3rE+mffHBmYCNZe0o
ReQ1mjlspqMhHTU4DSvM5qIaoKyIMCM5PjHCSbWl2xRF34QGkz/SN5UXY2OBgoFhudGfRJuKq5NI
5KQoF4q4G7yESVSsljs/S9F/LU+hNcBADjt73rDXUGABNd1wg1QgUNLGh3s5lEmN5j/b8ln/a0Oz
tdcm29gX2PhfE59GMSKr2OFcZFlX8jYVwf3WoM2QzZUgbgxLZTOvMdJ6hdF1QMGhKXYXm3TFjDrn
CfAVxuNoyyxpy9Alc2F7rkw1U/8vMUIxhH2kxmCdUi5fK98TUgCdIGm991fihHIuJR+ynVNxOaIF
JwPihbZ12iF9YPVGjE+qE6znev0ul+Acspo2xBkkEBWQHgB6Cpxn7f8DCoaAHTtvleu92FIrQZYJ
n/BN8r5RLiZXNUFgVyJmsrTATF/Jxzv/gYLHg4heqrJfZzLncs9w60xvvlSRUcRsrgp77ZHCePnq
dY4ovmPIni8ElD/SFNyiSdj9CqMIQMUsXfmxWOis9jysz0Whkcnwphf2D3IBYiveSupTcSoTunhC
9sZwZlEggzOA932t4xTlVEM2Vq5ApacyvRbklZrbZgWZeHk+S/OuQH4O9N2A2g3HoS3sXrCpNTTA
r7OwDuP9dhPO64B8jidp+woEzeXVvEQjkSnSLt4BlCIF+fXR674QRh62ZZHZL0f6Sh8Th+a2WZHI
hZPtSyizJlhnt6e/U4ZMgMC4SIgWiMmZ2Lt0Ur6HA1uOIGqWl8OXu2oKAqzA/FbQPolJ9LUsRi5x
elBfe3L8zvwI0SBp2igeoKAo1Sz6AKRgRtB3fnQN34jD8sNGh5yrjJo9mqjnoxfnJ38HR4K6WRz/
rbM066LSSY9drm7bOOou9s406xuCPiuh4GzXNg6Q2CygWehDh72+9eiGH9Fo+kRyAatJiRKGxg5i
7r9H2cXTV4aPszuT2d0vE4jyCgvrxP4qSvKJ8LHjlxnfrZ01cORONjPZSpznULRhOY3rX3KgqFfX
LqlyRnuIIxWg0EFtq8fpvruMdBi9bg+k9JfuWw9BlQDUhn/xlMqVa5Va1rO3PIOAYFjnkoAAUheI
bs1IcZxCtnArVGSTeYSlZemgWQ5ZCWPTtKiECmzCpJIiiohcKA/yFVfAN7yH9cvP8E8gQ+W0uXLV
ESK17pEV7mBKXYHVOdVutREWIrh7ciRZH2gX0dna915rJEpliMJmU29k1Y3OdJQ41zWRUqW+/Ysq
KXxy7029b78e73RemPE2XWb6Dbwl1hwQRm8C5Iw6YmWZopiTHyDjz+dmYVXeufB5ppIQBajlbe9T
kkBmGHwLDCIFJNvJctCKyB7KQvrtTOE9hRNalIHzBu79cGbr3QXx8OMmT9YN9W7nsKAV7oDMrDMv
boT1Yv6ibVubCd36qCde9Cii76wxfP8ZjQ0zqaTMGTHJVptH9K+1OZqF8VJLS2a4u3TFrYp7Zlrw
YjqgzyT5W/sL+CQvVQCnJpAobFoExszmiL6iQl993vOrJJ8y7+BMrFU41oPvGozwiM+X0xPtM2rp
Gn8UWIj/Lmyb8eIDWjHJpAm+YohPoCEiWqDGdor3qLPcYs0h5myyjZtY0LFji/CLlx29xtH/M/Rc
sLnnUnodfXH7H+hGqEe6Th/4eEuDwZtQV//JMF6uU9AID14qR8HjDc+uzLIMd3GAwFXAif/n1EFu
qBOg8lz9WGIB5hz/7QmFUZ5FrtfFe9tvD9G7IsT2We20/MKPWobIcMGNTM8kIG1zIHriuJcToDCP
zHAE54gBgbkpL+YKShQoWdbqqasAmcJAzHmVKKLLPW77KQm0BUOr4lCCiyBZI+kOC6qvz2ZhFRfp
68WlTPEB9B3IM0cz8a9n9pSaqYHtguD4mXpxyPNMwX3YugLXu1KG2hWpSSwVvllS523aK7bRi7fy
atrHsfgfjvXJUJmQkjm1HkPP5PAtGol56YBZwm/G8rdQ4xlY5m6Xj0s3Ycdh/p99NH56DCteYvUr
7irggWHtlKL/B/IIHGgytEXMTTh7/edoE5+eyZ+UvKdLiRv1BbOuHB5eeO+8Z4a8KWaceqJkJ6SC
AJo+6schj86LZxrx+cO3z94rErEGApGCGxJD330kTY6vIFEy9O6Nk/MPUEKv4iw0P1AC1Tmk0yES
AJlk1y/K/ZnO9cKPaTQwA4LUnH461SRdyKIkZydz0O/nbEmTPDYnhLYbS0193bKD1QAQbhFA266Z
ipUzVfwPKqE1xtlEgThIhuSnMOKXyBHvsWUl8oUNNA7fSFGlekKLHXHlZ6GS3t2TbJkog5sWb5/s
lsssWUwuXMo5CNLfgiOsgidIaXqVhaZF+d/FGj5BAY3KUf7ArBdwB/ZUXy96cMuEgS8cc9RGSv2j
Oao7kF11RhoH/qfs6x1JDA2JGq8VC/f2V2tY9rJjj3N0Xs0G8EK2PpNsLa/Z/afH7Z+VIGOqsEWi
BcQgahMvSC6HXHQO3xlKd7qjHXysFJEjdDLIAwlyiCuRF2lwJm+WIdIGqU8PfzPcVmOoWRb+xTBQ
TEMQIYRe0Go9KlFxU6Rjqxs76aoryInlwtZHwvhR7KQHR9S1pWD7egkU1I/phcEnCD7KsSJu7pEs
axiGQ7gPho8ZWIpFK/dbyl4XJQTJIYkPSWn/0iMymDHSgFKGCQ9+iYBQJ44TG2Q7Omwmd5llkDjO
+XRgb169SwqBEPKBTW5jmcWSPBzCdk4HjGsvEHG0e9J/oT09bQB/Dfu6E9HUDJ7zX0hcZOAmEPlQ
tlHS1AEjgDHoJ8qgbosc2c16A5ItpCO0jY3LLFhowd6iEBhK9bweaiMM2+PVDkWNEZh65plF0Jva
LGHebyUpXXqL36oHZZONldOpTfC1B9epo2vpfdzObGy9+VFdiFykNlTfnnz+hJVZ61fdAnHf5iDj
htkMTAiTk3X6BLSxngXwFdMqadkxqFuj9tNELuRje3Naa1NWIjSeyiDRnCHbTZriKPHTD4qN+Cg0
mYHiM8nkAqDA78CFuifUeK2J/sDVfPRHCEtktl/9MFbxm816eG4mb/fSOyETWBgDN/JwJqaT3xtn
9Nu4xRPri2p8e0bE+gSJPeMzBj9/nEKb3ftg2tTUFtFcrhB18LyS3EMNnwBO3DQiUs99DglpRw6h
WJu3j/z8FqzmS6wgZqqfhCtitB1QvgCHdb3lQBxGVoavKOt7ITNpqbpbJJiU7S03AwPvY0779C4r
BQZceC89vLoVtOcNvokHRQ79Ykb3jcoc5047xWDlBT9wfp+h3NmGJYJcj+6y4D9XdjddO1NHpcn9
zrYx0UNXry2fcxoc0qXYkbcVvqACV3m7XWqmyWSrIudNvGGcxh06ZrYrknbAp1J68oCNSYCySJZB
IUsileFr8BtOpsYoZ3cORzOBDA0fHbxn+iiVDxZGL+Xwq8+XeOgI0jsKpeevOHvEl9o+QZ08rrsb
cC3Dfr2Fl6nHWWakGiveAM28pavBq0+S4dIo3CRISx+oPi42C6UFrU/7d5S4pyg7rUwwp/46gC2L
KDlytqy64/zTXq/RZKjBvWp5+ja9ExVpWrYkNiefQ6UVKxUZVVLu+CyWtydZ+sjgmHFNEQV0oxP+
HEpcEUrvkNoZvk7J2CxUwHySAZt6B9+5wyWjZLF3cF1NjZuojnnaSFygF9vX1Rbc4FVepzcZLDao
zeSqnnSZS5dINVe/uYX/i4vIj2LNcAYMrAagw/VZb6mpj/d72yIOgTIBfAgw1K90l466WWhpUfOc
R4uTbUdUBNuGNNP+K+AoiqtxsiBDphl4JYBbnwnaE2wZzrfPxYw/+uMBAhm6t9fVyXphKq4cRe2N
T4Am2Ejw32DKptKE5Ii4AMGa8DcjJ/RR09fK0x/t06+U5X1HQnKDTn9xzREjKBiohbMxgFjYBNC5
IEreuzGq/FrTrBAfjQfLwT9AgUQSVRJmqmOAKUgBL3DXPFNdUdh6DmPKjsTbNN8vJHaUOTX+S6lG
8gmUN5n60SaZXf5u1LltThUsleFWM+S1rNZTixq7thjiqCOdtws80En9WcNx5iE3s8Fr9hNq6lMi
b7BdNm8vsN7ALpZIfZr/Wea06bUCf9PkIvSvFvOp51Jkg6i6gqVOI1ItwR2XbU7P0k4Ig67VQt8+
LfD4ZvcQJRr0IShGoqjz1fwJMYb/47MWDypGnqLDjJXxmLZEv5Zrx3BvWKbodYXrM/aL25f+wnL7
0qeHdDi5VGacjyG2iGgtsFF6sEWWNhrae0Xl0dZKsOgLSSZbuBAMrFssMjCV0ayop+zDGo4n2sr/
6YrrjYfPUsfb1W2uEkCRf6gip3uqWTcoSKs3YsXZMlB35dxNzSi0vaYglrZvcl1SY4aKp9C/u42l
HbZw5NowCgc0Vblkv8rGERZ0KUmRbiYSrxEQOMkyEyXcBTZ+5xJx9AzJ/vmckUn1J7FydBDsMO21
JyQ+Xrk7fPlMdlAPf8ozOhBGrZtmscvMPt69ZXumonc9KE6AiSy0cRqLhyWO3sFmkseXf8c8Jhtt
p211vV6klaJaW4bmAVTQYRTxcnr+CrkR2bX7KmhFsTY6rXFCkFrUcl3183K5DsalEfpkIEOyUV6g
Xx1h3SJeBKVILhxu74OMdmBlnmA+OUJ6sX1LDq4ffTzDrBLoAz9Ob8N2rQnuqfSmJwXUiBCP5fLu
XgD85PCUqn7+C7R6MUESay5MyPjUCljzegN7r8zerZ2JFZ1yAfDHxSZaG2eZTh7d0BcCyy06XwJD
MUynbOxKeNAN787mcqEUHETfE33yTb9wj29C0wZgS/nmD355yGg314E58RSwkDxvpUy5TCulP9B0
eOdWHtRASMBUgjPCHVX8oOYLyB4TfJ9O44Q9p8vjFUnN4UuT9Up/Sa4ztE4Ad5xcnAvFaEGhImUN
ZaAHK0ppgRi9BzbXLP3nkNdiNQTWVFZHnRV7+qGQmalmDVjKB+MlWU3stY/f9vgIOvMQpAfv+n6B
j0YM/XN7rvpNnGP4KzT2IRdAOYvNTcJbklpjf8Cq6t4etzPxXlzFGQLqIyMSqi2JL1oRFlcIzADM
yG6tYN13I12wOPwdn0Rgf2hJ3zYVns66oUzfiF7VAyNwGwSzPT8uX9ML5tWt5sxj8J9vO5skt+bC
Ux03Sfc410Uv8wOz/1WOQymvKY9RAqNlaPRLco/cDVNr3auNAs9hgJTXV6SFhGe6WwR81f3tacZg
fMUyT6LqdWxUubXHEud/0h+3GjtTMxt30T5CDuOyuL7ObzHWibjtSKt57Ip+poi91hN/i/C7CKZ+
xDPMQPT1+cNNxcjTW04p7ez41B6eC+YV5sJndCsjcSOxbcyp6ldDC2b+OG2YIN6LHUyT1Hr9UiSi
4qf/iLBIJDkYm5bUBduhoyUv9Nf01tvDVMN6Xxw476bui7mUJoajGhuf6L8Y4BANyqniNV6dV+zD
nLa/IFBCsZKhog6rSeeZ6zaHqlMbgRQbd4unr9TxKJck1pLBTC+rmnp05Ah68QwtgPU2WVGes4ea
vxDx9XCxWS5OBk/UYQfwi2MRPAUadymm0cu9A9Qhmkb6nY99WZ4vKDzMiayAMRmJ92wI/ledBLFE
XmUKXqWxrRJtBqXBS6GWIiN1QepfMeXIQdLyOUge495FMGEjMqrNb7bkBB9aalX9AktSM04+jQqc
gmmXngTsSCr0Suz6b7VHp+Y7mk5/APEYwsfLKZyl6d1USKqWkeryE2Lh/qQfAzFm3GC515RV9wZQ
oDpFK0DgVCsCQB5gxNaeu8Tv87ukwWDPj/cQezu/gkhmLwomify2spSS/BszTktA+PT1+CHNoWuU
9Pp/eQD6viHW9LfF31BbU19hFqhDgzqRGH+4iOLEDUr32D6r8cMUJ9+UuaC6qrF77nG4zGVEXIWH
EiE+lZg0VMjLpfwjAHbxkOfFlzXV2nSjc1oq7dD2mgMTHhF9SbVbwDrEl6mE6jFyr6/VMLAMJ3cA
OfJhcxL/4Sga3Cbc5DxXBS+xRZokw/BR+3lisI5SCx7bX4nr6FErlQnR0E4YZ3fQbmCcdrKWpoxk
K+felb2qIXXiH/tS7xXhWeK71m1ROIUNKN4mi9jOcuoGBUJPiKCHJb3EogGEvQUJQOMcwKim+HdZ
lUAJGJ9jGvGKuphvHh+JwIm7ZQe8lTaCfriE2/1zg9c4wfx4yFNMErjNMNSA28PcrwJ5OXnaG/uu
7nyD9u59x2OazODObdAa+IO9guCLbIisN+U2SB0PBrxWPJI7azDrV6NxWQUCMaYEikXAM/v6LU8g
Xbvv6shZLZizsgf4pdfqzQIaQd6HYrY7KCqmSZLy5Fz5jWJxGKGCObLODOqvL9FUZm4gp+FvB7HJ
gwjdNbNxhzMO2G2ix4nX6hOyG4gwHIRU+KS9A6OUVcRp0uoPrtvNgNDHTohfwDA0WMBxP5/Mtzbr
A22wx8vmIJFn5Q5Vn4XhQ5hkh8w6Fk6lIODXqAPwGpZ9lx8LHB3tRTw/ygnohE2o4qCSAspjhF4K
ObWPOojK+hWjQ/iSngVXUwFvLTvAfdMFWadnlyVUX6YfhnjJbEfUCi+ah3f/mjooZOgSi0J8oQp/
K/rOgld8iiMKQ0HqrWYWls56ucXjq6boYSRT7rD9tEV49X9KYQQuFPItPWbJCmdc6nBMN/xATu8J
D7JZOBNg5QT20rj2ayKdbf3OWsTxy+9eWwoUhP1OJ5YxrCqS7cLeSEBmTVTqJ8dxhq7rqA/nBzHC
gd4MlcAcGXYSccy91X3m2gIoMNpe3D9NgFbbzbHywYgtxmHhWBdCGmtHT1laf5+D4HjCkYQGV50e
NGnfXNwmhi9QB3cp58FBFFLUljdP0GsNOZUclSm7G3Iq41oor+Q4AdBve5sU2dZzaY1XXHEab+vH
6a1Og9rapu08c8QqR0plk5YJgevDwTxFnSvQNdFcAb0HHmzBs/fvzlvVoWAk1S8R4ANSfISkFq0P
3LPNFz84ojD8xJEsHPMqUaDzD6H7QJ+4tFg4UO5io+5F8zyRQ2Uqi+kgmUqKCe7a1gtuV4Pt/NZ+
5nDxhDtkM76KCsCkTiZuO/NbnZ761tiKRZ3RGo1o0ymBflcjy+cQQqYJ5/re2yPZRdIEqeQtfBIl
YGZH3soAm4UMETxssKejhtAYU2Y0159rIh0fg+9zYSz9VqbIQQd41Ze3GvXzhFEMK2n1X9ftVrQK
CFwTRt096ySMtru/FPMz0HIM7nNiGMCA8bknVAyP7O50HJnhCuekKyYoxYe2vC5F6KJlRAu1lxg3
5kbTCLVG0hf0GVJGlrKQCiAi28kDXWd7qR9ChybedXwu6Cd5oNArDtTztOo7on3YciY5+f3VD5kj
dD4LilapkCC8gXtzsGrVtGOWY/7HPY5vXnMdcuwLDKscCKVevCnkLaH9AJM+CDCxPhebXFGMqrbc
e+a9YmK3UH4/yWxo+2Q7It0rTWYRxOf+a84+TPgMIkTrUD9nntRWEbcECvm3uZHUuza36H6a3anb
MlokajpCnulhE/RJegFB3UL3JZ45uCCoQjIN6gTji4rEDRUVuCYPIXK3V2FeDawg8LfB/TwiOX8T
bRjt6psxJt26MewOM9PAhQOtisdV4UL8g8+AJ0nkvReOo5RNbQEjgiFZxg7sFQyu/yd4DDaLYFqW
WlG1bRp8RLWxrEfAN+tfDMWa78DLeS7a0gJ2giXQ7KGLuRpcHfffergTJS8Dggne6I2jFUikxghj
fGuiXyifLMaJMjM+hznLr+3w2LwBkgscJtHa+fQipm/JnKCiUQ9LidPWbHA+nxqi68Jt6XKshb8P
ax16sQA0GcI72ivRmmOtc72r7C+xAFXiUkCiLllw3n3Ci0QxhAxnx1NgctNLet6QI4eaR2+YDj23
KMdEsz5hzLtiFBSEkA3ad4sACoGwSkyS7PcLRps8imKqXUIHTjInKHd9qFRea0Aj9p54fqcITcuU
+vUm5P/44g/1xAHnSdIjOit5x+FO+2Q+SRZ4VG94/zm3zAdULmYe/q8ykm1bAfuPweatc95UABsA
JG/YG17Ij01I6Psd6sexHOHNFOCjGARxtb3R7QBaCH4AdfLgOmrgxiIY5cF1+Ufap23X170mPOMx
WZ2+DIAwjJ7IKmZvYd8iFpdIDvIs89aFTBefcvJeVHKX+JKcXJdtFn7JerrfIu23xDaIp/MPyvxd
F2fQUYYIIHaTQXfLhtXRo5dI8VN76/s4gkx5X8t81HH2Ksk/b1qOh6qDlV0jKh+Yjpoyun2FYAR1
i7W22/5AJxUVge6eU31hGnOHLxZG2UhYEJFhaiXEhc5ulbS6Kn6u2dGbYVVkW5LXeYj7mb4mqLK8
8ZalooxlNa1sZsQCmj0JKDfnw/QfRnNlBowF9xYm7NwyoP5UF0Z3g9qn8j9a93Wzm3J1VH4KHGc4
+0M4C9NUwLFO1lTSwSbzVJLFsZGJqugWRgFeGfOyP4NouW6n9rWApbnL3X3ivTgB6Z/S5lKp7+q4
FE88M9hsWLDbErGj2wAeWB4KfLE6PMxt1Pn6TYQVIFMWIrNlqRfaOBUrKc2dGRN2XHx8CdcOfNd/
c3gzcj7JvybD/XOXGQhjqffsd3sD1NTeJYU5HmIMYl32iZjhG4GMXMFr0ivq8y2YxfPcSHa4/EKr
SVl6fTeYPst5ZQ+CjHfb9haBJpo/drbLLO3YeRpN0rIevQujXiQ1gdsCBdld+SfbDF7Hkmwlv+08
tP0EqSwD1CLejW+JVk7v9EQoR+J3WohbjH+Iz71IDZd7ncM28niS3aHiK0y9RhSNeDMIq+O1sUuZ
k1sPYt6ODx+QD3fBtm62WfDEdvvUepZmVGqQJpcfBqKqomDN8tBdwUl7bGbO9EOjpAcAQ/2b2FRa
s9RF52S/TIQU7Zvu34jY5VujCFK+uM9NuMg262kepeXhK+ngZ9EuOT6fg/R403Y1rUeUFs1gsGuL
OqQct7cwusZY78J7ZzbxFU9JFJWGrRE6oVXuSNSsE4P2LPrll2ZtiHY0x5hrQqrdn2awbHO/LZ6d
1n+Vj3NkcvF0w7uZrcVq4U0Mu+J3KQkx5ekBv4w4LAcIIlnTJ3T2EyOs36X/yhPrzm8g7QTH5688
c2ZH10IG2I/OZ0uAh/uG9BjlwwmW1ayDvDHqGv/eXGcDNTqgx63l3vyAaqyhDY+6TZgo4u2Bcd++
T+7rmrCgh3zI/4X4H7TlbfzYLctDdlGhxY9p2xRDk/5cdKNNXaP3F1NJMvW0Lj1HnD3/ZtEO0S9q
PcrSdFywI5x0XLHrUqQZRq4rFfW75uYY48V2rhc5F4u9Q0AoZd4DEn7BfAsfHqSZrxgvB9SyzTTL
UiVxaBlz/sMsHHBpWrrx017KiROmsOlFsdReFgAu6X1C6cHWJ63CAW0Bf3GhKIEEgV62lC0hzMB9
RCTgG8R4l2AXlMRLbS37G57r8qsOkEtnBXYIs+YgWtFHKWf/B9kLCQkA6qoQYky9k06qYXmOaSU1
YoiFfPswUZJWkHI+D+uwrEcmk2tSSQu//ibD/yx1v3bxSbs6DotFNtvEnxSUi6AuIAVTWe2oYFGh
QclpmEvRii+iLuX2RbXYHksVEhkEH/zOQdNfixifcBI+HYxlKWaRpxp794MP8Hs3RNl5KJyMBUOK
N2fMovwJ9FzD4kXw9eUC3jW3rSp/yUPXraIir51StP0bs47UpFXn/QEdIYX+9qwLDZ5OWBGX6C/i
X1OPLDnxrOgbV4X3UVDLsq1rzV9AfeI+wzW8o1s0GWVhS0xrltsux/1MSSbX46nyW+V10qRBOv7D
rxYqlWCH27Bmd/zsS8LBCqZq2RVYVJ7KWsn+Wcn6+I0oB2nesmpu07yjYPhZVmYohz2q0ldbSHXJ
vLWJd0dYm7BukT2N0WerT5wdG5qUChP14XgUpDrJ9SBOuuAdI2LCrJEXhVBDnrfKHZMDAUrzu5kL
sldxJTLXjDu5JtMgndqljMvcdHYfXjUYXFnc3ND7SyE0F1nEZSNcXmKmfTEuDfI8ISC1V6qm1E5l
FqluG9MumPiJgIDXtzT42nEhA3oGw0B+B4jV8hI/Dma4GywS2+G/Mkt+ESIZ/O5X8d5px8BDL9Z3
sONJLnLZNLPr1ckLjdFR3ptKOcgqLWqH88PBxIlp4bpQO/rjjZRkbb4WJ+CpGFVMcCCcPy+4FagC
/DG0YZcsuLsFbbF795g8P42+eVhjrLgNonRBGN6dXYUzHgF3xYBnwcrdfJtHWQU9ruFp/NDL4enM
voJxQDvMgC62YbJC715X4l3t05wLplVssysfb9KBlSBKPeZGK2ExyvBo5BLzmf8ePpDx8DLLdkD6
usHV8qj292nkPDc68g33HkAeyKhIG3M8ZZKMS3kikRxauczDdVr7o7GRdu6afGvcAXcgJKnc25Ei
AJtrjuVH6gTvpF0pFGBSpRzLzai8r+4kPwOaRUhunp2iM4RcgXGTLt0HKa3p+WVu5btcTD8rARIX
QunmvRxhzyrXhyMoqZtzfvqgKZ7afPB6j9uJoMqTDfNP3QQPBtq8lH3V6OSf24Fq9xPJck6LUKIq
dAMAzK0wylgID2wzvDLdwjK3J+vOOGLyHy5J2ud8/AfzOKlZMSirh7tnfdm3SYO+942UPx7fAHLT
8A/GzONHn04q3YNyp040GQ7iXDF2vhW8ZRYO6IMgl+sZnDKXRn8xzv+RNSoCY2KZDgcGcuySOSF5
kdoxPbo8m7lkvzO2egM4ksxC1k9C0SoxRMOct1evdcWQXMYH9FSpCh8Bg9JywI6+DdXOgoLkwFhP
b9AS3+PNcsPtGRW0nEgqfR1tq/mFVyK14F4W64kSuWc58ZN0scNNE15CzkVDwQ5ENxObLJ3mUQY4
xnF9oZ/o4Hqpgs3FFSPZioPJ+4kJine+HaSjhd/3oi9YCumeTdX3X2/RnNFOz4DTalYP0ugkAKQv
ozLQj5lNu7jAC3STDZ8gUudzKHYdKDJxt4ryFfVb+UgCFE8IEINEe0Kl8tghPkDt8Ucv1YwEKk+v
AAbIcvA4dkJy856BCh3qUgy1R5+VHUfTM3DfPAcrc2qV9/o0r0cLMXXW1q1HxZoXOfjCa55kJeBp
+eDh+XDsofFs4qRa8g0DKF8zcbMxgfP8MMGympoD7zi1F81Y6lj2dO1Q6aIU1ZvuynLlefx/E0CR
b9AnXnFX2ngMFm3e6CQvIx4Vw1n93DpGGYlNlGxwm0PW0aNQeR52asWtLBtfECNGBIWwFTzkDVik
gnJHiKjzKeAVS/hYONCxn9dIWL4dYlceqYBwdW7EjyLVUE1GUIC4cRa+rXSYFxYEhYgFL94xdDYQ
KylZE+dTCYCaUcTtC/6/xS5cJ5IJzcubeBoyrfH+JvonreRx3D3AyjGDWSC3+mrDaQRWcUtOw2tA
jXNja7othfii9dID2r7KS6rYIUDOw9ZSskzpnkR1akNq4DAejQuM7o45A4Cf0SHPMYAyEuCRDZEn
+dGbE6lSuUNqaoei+9rXJL0kyrFLPIZCdJ65lwoSZhQL8pqhNzKpiY7D88BJi/d0vivyZ2OQECUG
djpvonuamKKoeLLCd9+pNnwZ60lnWGL0NtpcBojHhRL8jOyS8I0clCedlGAuZkX1/Q0VfcCrSte4
vbtI8BqaaovIvFxYy5JkcpKODDo5B33K5m4bEb1dUN2k+7b7iPcRw0FzTTiHhZH/U+i9yXPABdZR
SpZ0z2E/wrk0wJAp+qbkkTWhfJLswgeVH8cSGeCD3BIWbJmQsJmo3Tr/b9jnOjkW/06+DlBQGOUN
qVFMAMX4tl0t6YBeU7StTF4j/yaWh9qyQ00zHu8vFIOTcgz5FCKFrlh2HjnywiYWGhYo0ejwPPPW
BUGVMYu7PueotRa2kddIDMEfh4zNUp04VwS7fnbJ/Z8ao8J+ckd0Urucrh9Khckfp/S39shkefO6
JS+C4eV2sOdryGAtYyrTGzeUY7M3WErbeAUOfJZcoottq8/awIgyQ2a4SG0ByaaO5olH6y6vlyAk
0gYmPsFuE2SC2Clff5gi5YuHe9TQjcV4CcTYSzD/LwOlgkJwr47CEcXjIfgZxD+PdVwhvkUHMrUt
mFeombNsv4LxZtb81DTarqw1ZMgxIhQT5GwJVusnIFbWVDgVxJN/hJvvexNU8+TKHQ/hTmeKBzRn
0eLO9GAZt9ZQqHi/atvoix4AIJ1k3MJUSzc6eesCvbx4aeGfD5iE3c2SWV0SbZ9YYIsB4Yn9ksZM
aBq/KUGTAiOtq4fs9dz5f2KIEJl9RyS1GBUZjW1Po/jyNP20oVqJgNWl4DHQoVgninUeQiqo+JX+
/7cIaVVC21Fp3nk6H1zxBHnY/eeSWlf1hXI8S7lTe+aeNZqRaitfNzP8uGdZGwSP1w9zh6t7widI
6xCvHlB//nQEoyTV45+HiLPwfNo9BSxYKQ2E5S/kWeEFKqvHpj4U/zOQVzyAxz4p542Vq3afBIbM
rm41Xa08SCQLZGrE46OTHV4Q9RegaecrtCZNrVnxM0OOR6qWuMhcs2X6N+IpuNj1poYrSb9uR6pX
UHNE5bf8Wr86tETYgDB2nDWTMOh9S94oX7WU6I3YrmF1PvkKOPDx9rN9RxGl8eYrJNzHZd3qmyOn
0aOWSiresigaT+g0QLdu4r2M+K/la7w7ja9MC0FkRKUFZqkC1UCMUgC83NN0i8kSLCgWMdm3MNQ7
oBEd+1BwwVgoaYvax+pZKFkCFxHyaSednXFmPOia9JC8lnOoTnzNS/8H6pAo7i7+9XUjRXTXzAex
/HDTjAAvelM2F8flomECXUd8ZyW2bL4ypgeoeqk7/EYY3l+5Ky/nACNmqDNsIimwQ08x7lTir0Ki
pMbw7WunHAD4J/nAvn1AGov+rRcLZa2V6UNrCFRTyJ93HckoiTqfLIRR6kR2vwLEOS7N6b9TnTpP
wGKKJ+cBIgIF2098e0w+PAaB2iAw9PFPj1bzGPuCpE9MacEwqmR5S3p59HyAj25083ByVyscHikn
ba4O/h/eh5qXTpEf0yMqmHnsCh1R0oAL8smxf4dwnRua87RE0v7atzXU206Or7vDtRY0Pd1P8o7J
8XVmCaGyb3vMurqYO5Le4ahui8lhVMJCdNLnvvP3kj1vA6rY3Fs7E3gD1Zg4bo959TsS1psmgiK/
DYI/cZZWFy5AnJ5076QbnJIf5CMSF4v1DieCxbKW1ZjO8w0hnRQcUWZ9LzMUBmgdZsQh+n92dpEs
WneWhIsxkAP8qtb6UBQE8ZO5j+lhTC2qQPLWPewB7tGQB8bOhbVmQkIgwgck5v93dJtfEcCu+lvK
wZkRrJDiXW/PuNo5uNNXxv2tgspWQBWVNG3MyoEX/kOclu5OK+l/C72pUmhZ9v3sXURRdrax4OlF
zkXCHcdfU+M0s4YhTe4dajcwRmKIiWFOmAIOxYFmDUwSz1tZ30YURnoqPklX1Lqq9PxqZQUzYuOM
Lj3LkRo+sS2CkOniSeIZ/8T340lxk6OYxL3ZwvjC3HvUtrYUcc5uXg+8G9WI0qQr9qccUvXq2Oci
Nn4mMFGUrH8wpn0D3JjIX/znpq1NI2wrsSODVrK3HLMIyndn7CvtirCmcjSpR5ejHJ07+SfJl3OL
amLauxEsoKQJV566LOH/PDbsg+XJW52JCgAawieJt3rcmaFSgO3dlunVoifk8MPSOhFvpu/giLeY
kQhEYgrHHQxiSaAGaamfUNCOoSTJiU0/s9+QAtZJVb8m4LPXOAc+wazsx89pffhSfYSEhhh5JULz
NVFC7VseHi4s9HoMu6AOR4D2odPKVyVKCTEaMCQUlCQ8WWGyyMI36sKVxPG9o0ZP+wBC/PGkl8Xa
QGHqiO2pA+RKquEOgEUdvxOLHjGw2lpn5O5Or2xMfKItzZHTtxqkAtAzmYHWlbsWbNvL2Nxx/u9+
6j6lzzWHS7w3p+T8HoLiIjQ1ljNtIuF+AFSJ2Q5dQ/Mj21ZowlxXz9kXvO42nCvhg35YpRN93Tdu
2+7v79wS0Bm3ACC4Rt7yoY9ieELs/4DGlNxDfrNO3VNxPH7Qs6Vo78CRHGD90fbWX+JHrgxyQEpf
pec3p7abmR7fE9IFVAD1H1ACiZtylMwH1cuvAlaKSkmfhRKqeGzSY5JJYp1JLQ+iMHcxIrzaAjj1
iilbxvs+Cw48WsvIPoC104ME9avpMT8t8eqlh4oABiXKWUxs3VilQGDaF9Fob8UkR//nIxYURk0i
ycQtDBgjnzr6gmNI7pyOBhNNQZUKYMxHCZ36YEAK9Mnaqtdki66XC7UbbG4KFoV5YlbuDYfroQzV
4AufOQX7S2FtaPs05SucgXzVI512NUX8f2zbj52UUK/wMH0oI20ZiE0wvfbLxWTO8yKDuWbcrFbw
S/qaNr59UiQh4MIrGooDxD1J6fy+aAr3fcsHFE6yelyXkPX2YfR7byQxjzU9uzOpSMxpgcYOB74c
byLwrFqoTf5B+HdBuEqT9qraI7cyzMffhCPUJ+BpapcYuN0aZL4pBRgn1dpurImBUtixhjLLcNnm
q04EVlr6ZmMikf0MSUzU8/Dqc65zjNUesBXmGXkTFm3LwwwgZrMwQJRxyHf8e1b11jM/woOpjoK4
KCRrYNeMESptSakCOY2Q113cNhqen3W1kynCec1F8+aaB4ov4v09Zve1vbI5gu2erwTQaRI/bUgo
ARVt9Q5yrggst4OBMfLWZNaLYpLTLC8cWxMxneM502O0iBR/y5XsbMkj2Au381+5LLTriwjyE5ZB
yn1IeBbwsqcfRhno3ww4961aBqFk/c3zbLDm0YEPCjbrKIbbGU1uIptccayMhIQZViWV1Ys0VSuf
irLbydPXKFPv0ms5jS9Rj8yek8KPyEm4ikx50e3DdBusXVgAKQTXjsctM4JkpCZ1Fj6QP0y0oLX+
EeWhGnJELz5Csn691qAY7Wd+bUGMBkMjtOompHJ3G8o3psR+ZUDTajRf+Na8TNBJcOxoSIKdJfjC
ntsCN5F9YU6ieogA+Ds2jOkhpRcv3azoHepdgKolRlfq+ppKvf1d0vSRtcp5O6ashTj4147U76Wy
Vv1inNUDiChUSQtYLoCa1NS3rJ0mPFg3N3lLFjSObikIP1kH4HZidX9cPZkWXsVjtpCns0SFUELf
o2HNfX+Pb8T9fdyBq0p/aRrw5ez2Z8iOfspSSizENq1Uu+mBKeT7SYAxegL34r5xC2akbJANF85a
OudiEytqHi93gqv6T8YaxXn+umMWZekK3dqey8LgTFNoZ3m112Apth2Pqo2m4Ic1LvjRKHtvK0jK
3gPCcvQ9+/wYnBfDkh5hZYBoN8SHV+2caY7/wu8v1oaZoHZ+tXLjt99BnsDWjAElOy6jn8BzO6iz
c2Ag1iKMR/mArhzpjDzJjwSa3Qix32/Be6OFj+tjH8qxyuhnjQDncDIlO3j7PEJb9tFPuzt4z5nR
cx1O3YaWdFeFS/O1NGMHXXDhEvBdR7sFNV49eNgpPWTa0ZxT1BEEDGGk9tYrW8M3kL248Cg5+VzH
64ihK1/GP/jwiOhp8ABeADPWLXSiafVNYb+auRseTnMQKAgDhjF0OjwJk0P7S4457wIrzg3kE9nE
Hij9eDb1A8QRBo7myzPvsQBGPXTwvQ9Y+V5yMHy7ivgiPbGUpVVpvo9km+T8IgJCaELFM0hROsGz
NyVdZijKqOo26pBJIWAe5mM1DibRsNuzfr/RynNJt/pMi7T92hITMZxpqrwoHT8sMpUfBvTNhz/o
5mFs8rRlTVkksKkY+P5OmJF2xhb1zYA65eBdR3JFkTEYrpIJttPjqqtVrqRjuAmHESOczePfQjAA
KnQl6ThLAC3BQZsr/ZmAodKGU9U6cmCj21AUZ2YTEEs/7uWs+2XhSkMOKRi83KfNkgsH2fdY4vfc
w/nHl37gzUzzrJSsqQBCZBFjjJlrq7994Tdy5v3nnkBT3salZvJWEoSRslWbb1CLUih2hygeYivM
xnFjiun7r9QayblbCWUJAy+EjwHfd/RcRCF/6AAjzNijFkb4UYA4xVidUo26ze9mDao2ZPNNnI/N
vRhV9NIyu14ePC/LP5Zh2fPmO+9iJ+IKIHOyWCtYEnwVDPJ76jSPh5cWEMWl3sd/ZU2M8WDd8oiv
LvlkIXsY1PeOFeT5yBsFzuVQco8J80bW0eUnB4j79Wqkq2sWAlBzKELeLlnTKDC383zML+VRjuet
hPJjfwwh59+pIMFZ76XXRSsQJdctPFWjonQR6Js8wCH+rz3tKtS6ha6VnLgkYnhSFabyz1Sq4zcF
+WMkLRG+gpE8Xc9u5JR1HghSrQj3b/R834z/KuAwQ1ELr+YjEx8lm5TpvLR889rnFIy8+pqi/0lQ
BWau1WA6HLeLpYgEtsB+tarvXClhHy4LT9t8y6OxYftcoWSh8di1h/11oFAJST5ZBXCmhPwnGirj
SAiEHOeP//LQGTLcsofPST/l0B29aFbb8A+1KeAfCaRUGPdxB0HixxFosmVVNFFCQSxe1QIgwS+z
SKOGCAwOhsWcyXghcFb+KB+98gfQ6q/bdKw+Esd1i+T2/jQqtPIxrnWRT+aIgyaoXTbsZwDNblV7
PcDXoe+dtWcLi7OJNse5H/U2dmh8/zBDmn0v997ShN1+m8PBbasHEgJUcXB4+BPRN/lDCNLlOQpH
C1ufKJPr/lYaJpfnrk+WUhKgXARWaRCWzm4BTrUuwBaJWk+pFH+iNnMn/UPLdnM7tAbURLaYx/t7
/uUH284kpnowNT69plT5UDzNPPaXuDVeYgVtz1EyXYBr4945Llz5hHnqjwfzsR6p+MScKjn9b2SP
ivH9PvIeIk1DlgCbHmzlJ+hUPdiNqq4rMjB2v+UuSCiNwgOHgc0B5vbruZKAIY5Sn3WIDl7Fib6F
PVCvWO+m+RqurApEY2AMnWgzjfPqWls0/leKEFErrUueopvPEgSxyZAck2p8L4o8nqT8ua+jIFCN
8GR1/C3z4P58gatjYl44PyKGFHNif2fhS9Qbna7nREx7lPZfIA/xuAYZT9LrSX2lZ9kIo4s2OLHC
5YL0z3y3+p+epi9lzNz8TAQiIu2vDhMRBAGWRho4h0+PqXOMl+P1Hrm7WLZ21cFjDlU4xBW1CyCL
n/wNBsbaz/Fz5kEWHl/pR51VXZPX08WftQ3Ip7z2LzNHHeZkvoxohlsniNwhCMOL4+9Zrkk26pi9
8hKAOmmEyRcwoI+xWAb5wgSMw05BLpP+03zoyb6JMf/EhuYpCHtKTgwi4ZyiPHHXs3NVI3bAXhQr
AJNpJ1RG/S0XJDo+x0cWlK0ETIegki8sFhSk8ukhD9FMIWmmiSvUsG5BOiBxA/ANiGZ1qR8OQmEm
p2F02JyMA4/7CsPfPJkNpNs8SvJ/Hnoih/PD0AOWTRUwg+TBOLywORsylmJ79uq6Q17K2/nStCFl
7Fsx91loJ+QbT7li0rZTZgDSdrmCgspq0OeMWz7cWmatYXz+CR3rhWv/JKwjkVvxqfNviuBUX2+1
PwNO/KyM40zZhbhFGPk0rfkC5SwV5zomhUj1jbToZUl2cp4Ngo1rp3iSNBSjvKgbzPCtNKgrUymq
v27UWLHtiWWB1F4520ujj+Qk6x1hjLIY8sIVjOGBIo7iwcJT+bP30Ar9h7HPx2EYGxf33W/GZHHX
5L2CYzq86Kw/93OSn6+b4LCjPGBp+NjvymdrCguxq8qdmCSj5K8j4gNiFDp0SDTJkNbTNRVcvOUM
3RGzpADSFRIaO7FF1h697bLWmZnumFRXsPZnd/QSyLx7361cBsWVTP1rbXbqQ56FiyluYd8ofTr0
x+Z1i9PpqGSn86VVb03Ju8K3NqIi6eAlfM1NIipMJhhb7cDiOlUoH92uMRY2Q5tBDqm1Gk0lxuRE
GB+AUT8sl+2hiaUpCB/ruLgF28LPoMurN6+SQagCEtSrEs1QRU0+qPTtK6J/SNml/Lj0OePbXH84
WUQ7O4PduhfZWZfsy6hBgYkZSb/jDfypxXew1vp0az7hoB7IGVefFxdEayE3sGSXubc8uVnQaWL1
XwDsv/oQ7dXQYz5Q9RqKBECe2aLjAuQvtK8rK9e9fke4142FiG3lCNYf6RGa3a4Kc/0Ilwar6rvH
2JtDatNRnmpRaqhHC5SGLuQkiHyGTFdTA5tpwy17UQU7wvm0JWDMAaYq5cNVpm/MxjAaJbC75ECA
AlkPor8yS36uLqFd63VSt0zcMxx3oVwfTHCalUzfKe2SMu2pndSNyyKRfsKxAU2aYDgdgx04bPt0
FJgcz3LV1ipHWf1ug9JBYg4QezQGGAsrFF0jDasCDTM+c1Nst2cIrk4y2CnGUBTkWLQRKbl1oMS6
vP303qBW2eNgqlI7oJjrH7BM5s02vxhz/Sp5mE6lDR+kJoZPEGDzeef3JyD3EWnhyw3a2eN+BUHl
jbMZ02UX+6gcCvnD4y81hkR0nbnh2T3T09jgjSeb27q3ImxTYnGBh6XgX8Ju4rOK/F2BDUMZ5r/I
KYVNq6XnW+HOLozSb+RIBbFKRd9uVsDoeWIyCmc9n36QcpHGbo8QtaQfl8BHP8K332X7+gEo1Nk4
BDyErZoE09YGX+CEWB44OdJS5wwa8VAoJTB3y7RSdu0tOT+Sdt80Z+v8ptunveEWz22ZDXmXz/IM
WcIU4BxYT9HHFe2rlzRAAbjZFXRVlgvsKye7f8d/dyxaxajTJL+8F03gxz71g2plUKkUEPTSLScN
TnYFqprrnGy7o/DzXJBEf+hGCHoHplTkPCYpnQ/eWMgQKFKyWm/EIbGvZztFX384bqSRY0Yo1r3F
AQODJIhr2lxkORTORTGWr5yWobD3WCFCEDUrD/QcLIeZYmm4GzP7qFxKtBiDGQlk95ffNgFKeRMX
BOAre20WPlh9aiV2pTzMdzVv7fnoW6yHl/PJMVLoZqVxRoKSh4ghlmTjRli86T7tv3NYzAPFIhHs
DBy6/qEtz5aGhcrvGObPga4yfRJdFB/hD/l6eqhFvcvZAv34AgLivkuYlbyjN49xf/IyNT4YGbC4
SPMLUvMxyMcJRpg60mtq1hc5Tob4rMrTnTwLSefqLNREMhntBygu50m5CXAPDS29tmYxvZ3mESfH
gF/1/fr6l0ZMQlp5wzT462HeKQqFazJZug8HMt5BLJpY3nZ38Ess74oi3HxMyv6BYmL3FTM8s9W4
HOBjYWM5/3/fHw8dadK3dURsGw9d2tsFyuCmgSY08QLz2KxkWOwgViHqlis+Jr1hdOR2MFWZKTMs
xGLnt+NWAtINM1dJYy7g0T99NsPziaBaESMip35m69CsAxM49EkmxR57fFdlg1uoF/ckdX7yQ55S
d4LkQRsnrXov15j66vZ9GPceC1NYpmtIuLHKqfB/q99eiyuuO2/C9i/q1SHJkc47uke9/PInDiCY
xuK9jqIgLWXuY8G8iGN+x/2QU112uLvyl7jxmcu/DgE5YI6R5nCgW/UI444WzeZKDN8sukVfQsaD
KZ3ODibHHIRCoeYIfzCSA0WtDeJLnkIhL+H7tj2QSdIKbtIcM9ZGG+28PMAC4ATqbqc1AOrqb7Cs
H6eCuRpevmrHZmow6BfjpIqjkknSPYAjsd/WsfFS94D019Gq5tfHYA3gdZXjGn7m2JiHx6E0Dlp2
1Mye9a6T/F3QUxXe8vjILTbFodDvfFOJNLEgmYayx4DQNK4jDtG3uJsEZY7bSNUSEmEgU9vkJPsz
qMaZb8eXTwOCKvahUF6DtiicjXNGmsBslSzvqscGsT4VO1ST5fPOPvalgm6Ivpxsetkue5AQPQbx
tIZJOBF58f2xR6MTyfnyxp/UH7qO4udsVv8jIGG7Z8U3HVe7XYc/faxZ4HScSGdMKbIAVXgfCpLl
mUz/l0BxVH+fwkj28sLl2/IYaJcS63iaf/Q8ykF5qNbvwYzHKpuN6lkLEdZceWFvsqtqYITNdsii
6DnGqwdI8R5OhXByo0j9hbEPjyyY0Hq3jmd7nXYgC2vgeSq6tzbARMOj1bb8nxraGwxVRziqFyy2
S3vKykSS3501k4YwRgs7TIItP/6O0gSHNhIV1DK5w25xs1JuGC9Pd31Vc37ytAlBLsfgMCAdzaRT
jIx6py2Ej0J0u40cnsXLrbfxcY0XN/Gws//gKdtXSidJn3IZ9wqthpqGgtfvgGgkIwkAXJFraudG
/sEvtTQFkmsMLFdgsPqA1PP75GAzI3y3YdJMlDycIbqjS6r0kY2eFrQM7bCTrkTznxtfJTP1ughP
1hLLJYugThwHLaYZ3D25ZdT+fA5lwfDsaG9CPsg+9t6whHGVzdzrgWbASjOGhb+ufgn2Mg9mf67g
GLiusGZ928YbYQ6OF6ZWmw1JEXNz+jDE/VoB4NzQfoYwEo5V61PcMbXc1Q810ge3rJfXPhKRLjw4
b/GckQzHRcBodgXpPAVPSVYkztEaUvRhyMJhy/iglxFT6XcxjaM2njIsJMkqIM43JeicB4yLP2q8
39OD2g5nvAzSBYj6ki6Yskg6mOISkfnD8i4awS3NM8Jis8Yp7G3TVTyvFuvVT4TwEH/Ji7CxsDKX
UX4sY1MRqWwkeJdPFJ1Hj2w9E/h9C+ut1zDK4GsvwTfhgdO+5vL1ICc672X3mXvZXyhVA6ra5fjQ
5mVHawNEnshqVINybCmwumqg+JrpWhQRw4x/AA7wSz0uxZKUIjKk33e0IDq7NHh/uk5J9+eHoCet
//VXL3wgXUd8PebjI8o3A0r4yQdgJD1dt4yQNKT2scpoONVU39+vY/9AwnHdmjHJgaXTkpj0WER5
aXAqzcLZCy4PuDuJR9KCyrBfKV1gtnBgnS3skOrR665OBNpEzY1P+lHnl8FfCxFXZpcYIquOjxeU
yhggxe/LY/RwAlhZkmcLWvg7KTltJrDDwFcNeBtT8IW61kSkypf/qRYiSGK1SmddZEl6ehmPOQTA
Bb9XlcDI4x6zhkXE0YIDFpe1kkzoY+eV4DYaD9jMsBQUizEQgIjK2zIEbeequDhvVWKNfjRu6rW2
4OOsSSMQORVvw+zeIeFsmfNHjZ2uzhbK4ZMFio1ex5gu21yMLlHhfLeLb6WNASp4oSiApARqp6bb
DsSwE1parRkHU+tCL+iqJsOnksFTEHknIb92++IjhOaMzqgFS5WaNaTC8/F09lzjeZKIvZliYzqw
gYL5Az5rXHL/IB7AdYhTwSsEqE1cbeWWhDNyZAIlY1xGew+kR1zmjckqrpi7TwTPDOSWXQSc3tHH
Ebl7ANTj8AgUXMqXNaTTubBEZrKDMdunuExIgM+cYx7u88LnxGR4v5ryoExGDJhSU/XcEuhc/NHe
BSYFSErYHAzgg5hbiZSKhjpHu1bQ+QUcihj/6bPNDOfqvH/aAurQ9tdyIxd4xE31w3ckl4IyW5c9
yJDfhvEDi4CYtAVZzgzvQ7DcpYglbV2GJs8EVrxEncP+Lp2xB89U+87lRcu6LYKTU0tOsDyo4Bm0
EHOJGJfX/jarKUjusIR2pvdV/iOj1/w5arFrhVvLELN0iAnAoOQZWeGylCFRxGlj9cEiPlVune82
R6byIW4WTWdEMmkIRsx8HaPnx7nPmc5QN7IZRQGfogir73+YfU0XYVKjhuY7zaqItWgzW55B3jT1
IHMbpnGsZClut1A+niSkz+4I3pXLu8CujDsC04LNKqInN4L01xaYeex+YZhzWsWVEuUjTK9dGzjS
G5GtbeBCIYBxOo4oBcfLDj0sC612BMQgFWKDuzjp2q4nUBe2kVqnvh+rDOaRfB3mXbVMGu4aynGz
a5MZkFDE0ASAG+GNgiqvPSMz7FUO03fy7csE7nXtCyP48DX1f0sYGWkWlh4y+x4DecM1AEEz4G9b
mnMl8UsOQLkiV01Pqw6md1XYl1KHCjaxI4sCwjphdlpCZp6RJJzorQqSewrQwiJKZbzn28j2Wvf5
ipPtYoixsofljAni2qowUGOo/NBR6qcTQkRw0Vk11EqqcXqqI48ZqGLvrLeBDIKS/QfW+e9n9iwM
OKp9qjOg0GsmflOPpoF/jGsCeXxYl+xFr8q3K7UHfO+Q7XowR8l0urkRQ+Oq6j5waYmgFUj2UnPG
+NMhqVRFq77umBLvns9kCW8lbJLkYl15fFro1apfdGn//gPeXmTEibDFVYUO01mdr3tIwuZlF+iu
R7k+vWZbIpzIkaFMNL9gAXSJEZR1PCw5tM+Ik09DKYf9EAi4d6MBlFpHQNuFiakENeJ9Tr9E3Fkz
dw0IwEjdY8tcHsyYrPcEeZ33ADXrb4KEwFe4qPK1/7edwIQGZQ3IDO9uPrlZRb1iTYTfozTI568j
IyH1Y93nZtID6AYNoT6AMXVE8ptuYm+tc9LFcFEUhWraSf+NyHeQr0pw8Ek7mufJuH62gmQQeBkF
o0tx412RWCFIzS6UN/V7SzSH1ozVKsHQbsWR1ui5xmfrbqU6f3IE5Zd0URv5OoHeybBeNb4Eq7YY
sHnPwK+oUrD5oYLVzKWLGQ6Pn6B7onYfCBxEsSZJlDhQdM0hH25OKfeVpv+AfbR/iX7cnaYBd6DU
qb8/MH8nX4F7YR6EMhx8duBgpmBZxDCixsOTKV/Uu1mrjiXZ/fc2G3Zm8a7f3wF1CdR7+2ufjprg
Fz6nRh/ZIHG5qO3GMJYNazxb+2lkxz4rqwWyoWMXhjHHCiuB6A7v7FHwvD9VcEHR5AVwQ7HufZoD
OW5yrF+h4SyyY4u0Vg765SsLP73/4EBfhzT9gNwcydLlo+5e08O0yKiHNNNmL9lSFR6vKPA0OEko
CRMoyq5slC1JeUrn3SCi5YPxbA8mwcQuWiZP4XFMO5Ynq1aH4Q0ihjkoTi+nFOqI98aqVsYaFUz2
bf9Ex49PJp1znu+Fkbcai2H9YLOeZcyysoZSpz3IsJBjo1N75SXx5t6/JJ1yprL5EqqyxaMWbty0
pCgFa14QuEmXBpIIaYN8NmCBEVULq+4+FDS766N0X6PtZ95BMxK3HSREyeWPBRfDilAcro6sn2bb
4klCVh9ghDXXlVNXp89WMuXCHpTKkvKSAGpsA2MiZdZjqdfU7Bi+uZIlxPbptht2vbTufmdtouED
hzIeJJxH04pfTFtoSoPgV/HwGB1j7X679XRPi7guRgT6efqamefVHLISrvKy0745ObxrS94ix6/8
1iGnXP1Cwzg9vdT8eDGSFrg5D1pcBdeEmJmZetsowNRrmzZDklC1QoMTZ88Ei/uJGvIA9GJiSPJU
Wd2vCnkHzueua2pQGd9u994SQo0YQjHnsxXRPI9WfIGFK8qlYHUAOw5tKxn4qi9NYh9FDLyeDz9D
Uzmf4YL8s02XPWuMTItGR4tZlnA5gbFgRKYDRoGehe/pAwClUcryUIeoL/G8Lvm7w2xi4OuRBCyl
A01paqjoE0XlKZwjzUTvogY1Ee/sQrBmqnNxemINaMbBG0YgWb2tEyFtXsxdHuUpWS1b4c8zzG/v
I7CG+j9aeWJhVTJEheR+u5oifML9uEafZI2eFDRsnEj6dKrTR5M4qnr7cStCZ63uaoSN4biMSCIk
HzoChNtqbqS6USeMr94PU9b6IleORHpyZ/y+Yi/rYupadBytvfIER6EltOJLHWFoNsc51pklZh11
XZC6GuDRNMSLrT7zun33WBvvDXTlnEXL7d0zJqW4+rmMXCsFToE7uWKrhm5K3ls9bv1UaChdfJQ+
fRM3ERvy5B0gPqy/3gIbXQtrlN9vR4Knss6TMkHQR+mP5nhl4w/x1CUTSBtTuHG4XP0dgbuMRdW0
tKr55A2822Ueh8dNf0aF1I2tdzZGYA5UJbEtEeRaqg+e8Nn7wKX9uPuwLgziQbxO1c3iNLpNxilb
Zx8OKbmIxnLnWrTzvQfcLvU7SqOSebbzSnNMvY9pbj9hg8I618sVVr80HFt+j08rx/0y7KUf4Wrd
wjqO7e0wHi40fUGh+2zTsSwvgEaWITT9K06KtGiluD/LvzSyUMnWxktBD1ngqntB+jX03zTLCtuE
QHQk3kBJ14mHlWPFW5sgv18DqZxmhwWLcP+mghy4b52AnevBdpEZmApWsJ28f/C1Zbw2MMZPJvlh
io62XJWEdUYw2QXKuIWnmreqJThuwBNO4dJFBGnzndluOXiOITLwe67NWj7QOOGevCRoAJSNKdlp
CsrUB4aF4MnErP1qwXCy/QLbPXB23cTiEsVL0gPujoKCKv4Fp3zp6BAM3xZNneCBkYNNo7q/p9n/
60Es6QoFlYwcj8aw9Z0pKc1dey9nS1vORfktaj1P4x+hLkc/Z5q7CzhnySWMzNYkaSMUQRYvyjND
iQSDoZEpJVQtGQnRiyrDBkIRjkZm/peeGMmMW9Zqne5gjbZRchN6SzzKIckUmbIUiE46nNz3eLYy
Bg1J79J8pVKrBMUQ9bOMD/V2jBxJgKTeoOkEke8QjNBZZyRT9g04yEfuU7zwh3VO//ApDH22beWM
V9YlvePkd5E6GL9R5IoTurbAldG7Zjr5wFkQq0JLTcuMoSdvr6NpXQbTcHIvaWfEE3XT7cNltuyX
ovwXD8bHGdN0VE9JarZcfrZwHAK+BiKDlnYFjHqpzwEuEaVEBIyi79uFp4oWH+U+IRNe3xpEVrcK
cA1uOSizNMe2kWflAvGLQXww+Q25j83nQm25FKO9cxB43UpT/y8bUDWskfkPhDM7RZt9Nx6o+UFr
UG/Rg8huTNkTkloeLC44Y/siQ3JY1UrPZvfvZS2T999DVjh+ImiwYFKc4dn2xYoHEEj0+z8SAZ7P
q7++fWXFal6j2hxlwVAJzncOl0pBb0kH58SLuZY5V/2Apqo7jjaowt47ap7Yb0HkNeoFlmueQFaW
+v/7YuLh0pUmJlRt4Xna2NlytRLaef7nZClKpdcHsso6v61fkbSSdn5jgY0Gg6kcfjDredSXTyRs
ISgIfKkQk2RIQV+KDDyzVN7zd+s1lCGxISjeL5pkaXuLGL0rXb2sWbrUl0m7MJYpr0kwCEOsashQ
DiDJ8SrcXvpgQVjKHSKaS3JJ9SPsbnpdYQMGflLtihEFxQRosOtldSeAUQVrqRoSdSse7oKe4Zxj
0eply7kX2TD2/5uLwxe6eGsWBvENlJxB03O/Csp51D3NFmvpsmMLfiW1YqioIzbB8Fj9Ou4vJ+sX
S8lCsVQXrMtsW0ehsCQNTbOlpTwpediQscT7GHvS2xDai784hmZ65gdgXMzth76xO01Bfj34DI8w
BJb3sRYzRvSc1lK8l+s17H8Gl2l8E3vO7pMG6zXH10VXY0KGVjWV9LSEY6OCEJxwpBYjRVxPC2Qq
U6K9vEbsCx3jDhO+Oyy0PngZ7CMy038n3lpede2fFKxGnkFcOdCc9CZTS2j0KQQggvjc62l9YbIU
TY4UIgvHV1GSawm4kHhi8FTem/kSuOZJT7gDTur4HKaYCx8esleHtMZLiW7zraJ1MDgu9cMEDwpb
7tSlDVK0g/5ECwuExCXfHMa3L+/c2HAhlhyOlckC/P0ove0dksM/0Edsu5GACI4wbutMjF+N/C8X
wF93r9PJbden3HlCw//c/PoY5vRtQVzAEWgoPWtjwpt3vCi1Q3Y0vhaF6UL6PrHRNrgfH8JWoddV
XylrJv46bNm+ghpfOQ4FRBH7uuct+sDrF2yLdPl2NW8SKx+AFBHtaZcsaFzd0Qc7SJMc3X3KI625
QqJy7hZgteaHBa7TxCyFlXravR3hSqf2lVSZdX1JoDADObnsob748e6U6k7SBJziN+DO0J3/KVzv
GDY4QlHKr2thI4kmqG5IF6fTy5nlxTVEv7kaPsQ2aRMhti56kfLjOPQdgGvi9eyKZTr2EwEjO5QP
RQcTflmvheJSbzT1/NUfVDxTb6cqRx+4l5GkAodhfhnE6DP7dvsvb9h250TVn7/mdUQZLzom0z5N
BQ0aXGB5YOtR1OAzut65N3XTGqtXhxI2HLpDTt1vtpz7R165ipbFwwQzHUJVYGReBNnxptHi6e4v
9NwSH2liiv+cxPi/XCZFfVJrmfjX9WGf7yq8N9IEkhwG90SEpU7rAuByKCOE3fbSE2bKb8Sd/cTf
f0YrCNwk9L2163W7LQ7HIavCDuNfgR/ulixhG9F3J+kDDL7/L+evmQxHWFUJFVjoBxNFdPADaLjP
qapghO6WD73j7xRRqvvT4pd5EoW7o/6qYw/07eAkd9XtFBqzs7dq9TTa2oaSWME2+Q2XwaTPLsCl
1xIcnv5Bngi5cAIxAGqqBP8YVhYHSfL0eO2hRuuHgykchD3vhYD1184PvrQUkFlZGaVbb3k/E1fV
kXQmnxKCmPvnPQBL1QVwlJeqY5y0DxyokNWonCQlnDLxrCYCtVkxt4yeyI6mqLiw4kF8zrY1VvtU
HjGJu0vv5lpFLyPfvQv/Bqj95TUvIxTkha17dSk3Azj7aSEfsDOEIFSLng++Lnc+APMKiTCdp/O3
Lvs9YQHo4Pbn0Oj9kPsHljAnNf0+xcEBrK1cnbIn+Wc1QjAxXD4JHnDy4g7STbDQOnVNgAoYUyCx
R/4qCn5TUzrERXAJiDYE0xYVKWfplgGTgYVJqHaGhUFApWveeDukhOVFFDm6K0OLsTzJl6Vsl7SB
A9uTIdoav/797jxrwlsXMIfjlkW0YgyNvPo4vTY268/FJffSVehtaD9OyiCzA09MvPqtKjZ6FXOP
DWD/g/BDiuDSUvjFVTO28ClAKOcv43g7oSbiVGYgivCEQS0EIscgh9MXc+bUES54PfiC74nd6Jif
IBHJNCM5IrDT7vAuoUAJEp27qvXBL3unE5UpcecZPAzsumFckQcaYoVwpzXm7AGVQNgklvmk9v89
S5MRpSjuZATccFwZL4e1VR8FhH8ZRZ7o7Fph1tF+l+IZh+6cvqbavK2P/ShR0G1Gcy4hPaypQJ70
Qb5WG42idwjrmBp11zdk30gfqOsQWOuKhzAI7TH3Y51DRk/m42S53PMpETIjKUOjITeS56DObpbX
0B3YJy4K2sUFVOZfm4OJRJKBr3aG/ye6UxdYIYiaSkK9c+ZuMTFxGHRHZ1PcklTo+Ph2eV5dzscl
Fk1a9KO+ZyV6OFz+npi/I+27ypHWP0GWi953uxt4eVgdozecvo7GnpS+1p2A8E5oZDYDGuHi/94q
s3f8vG8/HmAPq+V9CWiE7YRCib1D2JKVPftC6zz6uQhETTVxtERRe2wDJdj2usMywCqg3BqOkmL4
KfUXjG10pF8L8eiVqtKe+bg2D8hb3WLVoZyo4cheQQKHHQw7pFForE5VmivgUH8EvZIO/yvFI2ji
eU0a1hID/5U1ZFZmNDEuXZq7ZBbE2oVEkP8cW6elzTIU32XjpEJztL4OCe2JvdlV5QVv3w4xKbK9
46jYrZHFSbZxWAkn/zQhAqE1GWsNGYCHKpaWJUxiX1x2AE+z8oOg7agpmkwUUug6TDqhTklWGO3a
29NvizBfafnnLMw0X40owwfo4gljTTmsH1S0W8wjnXEqq70eCVIzXkfEq/O6CYakfZHUam/WKBNW
kcI3pdqLDIc5g3+gcXiTR7vArhiAZwmNQBh2+nUfK//wjsaE4YcTZMN3AlUhEl213t8D1g6AvREc
uc8A6RVa7fQxURReP13ZkTFjtlY+UPX/KJHwd3xRQpLpdK3QMpeN5oDEYN98JfmZpkUd0Uyy2mwy
p26YaresPr68/hmRRqhw5SJsIEn9Glw8MYsq6+0tAmUSybVTV8y1Oac8qNo/hIaI9R7Zl7OOk34y
GOOD7BEz1X/KQb0bRyBe/W58MqMrsgICFeCwfgtDDlpA5sVFOVpesbYg2/HQ/XOBC7ZOUUsG9yVM
biU+iqbKcCH32bdjE1Wsva38izPV/2KGphluwHnDfEbL784FM/MEucqNpDu8z7cDG/Si5MqwL+G2
0M/D+MIpaAjxmzv1VTbd4keE4MUoRJBhs5F3C0Sgna2Xg1MfYC7bpMKMtCDTrhQmioyIY/wQAaWK
EMfb5Z0ywFNRWU26eg9aDRHNUVo03+NxIHU7ddUbXLv6kWL5tNfk/m+JIxc52RySnHIEEejPSJji
Hf0IInXZrs8vCEotifzkPifKkYX5/lVH4HjQdPCfIeszj0t+wpj/tm3qiV5ZOfGZ/0DZg/oOdOHF
lMz5vCIDM/Q4yDhgJGUO3JB+TnGDfocKU2RQ9sPAMzXyharSIN+6I0tOO9Nw+SeihgJmuAcPRAVT
FJyFlyAIbAdow7rzyupfr1QIxzdIDP54dVNql5rl1+uA5zLJCb72laM8b7w7ydpR1EcfzZ50z0vm
O3dfdyILiRGPL7pmzpEScC9HYo3jGzg4RBynHgAAbzr3KHVdHhP3Xmsd6fjsOLdYk1MR9oISvTOv
YuqOzNtSpsWdTnJBIvdHvy92+QRBXY/EDUsVvSkjpMOFywuG5Aef+hl8dcMrW+MtvXKc9Et2/hQD
gnNMiaWhjvwMjiePjH6DdQiGkt9tZFybZJGn47SqfBiuOLu/TJMJkiXDoqKU9ULDiR/UuGUmoRII
SRerLMKP99cL7NMfw36H4zZ4ZHlV6pHSrUY3O76Lr3dU31Cbx9lKYC3EtHLurVskeNHZlDlKZ4gr
oD1XtBr+3uMh12Hpjqd1MGa608BxkA3+jmwere8MfYdS/f2dT7Y8/ZrsNoiX2oUOK3n798hXHudR
ErrUvdaIHkTPf7ew0U4pMUnDAo1K0h3reohpbLvRpDS239+JErIXbm/Q0gHSb6bekR6CDzPAkg5E
ewMj5MigHD2osEQ0Ts/wOB3HgnCT9ottRkDaTAyiDQxXt4hsKU14H9j5ohxuraE95xlLBclaq95k
niOGd6AxJ2P201kbdjz6MvTZWRACGBVdj+XTUc/2e8KDq7ksvk9wMVAr6SjSJYDVVfhvN2MMPrfc
N2RmvTZCAdqioiKdXRKOkrkIfjaiujTDk4UxSeioVAeuyf+alGU+fAYQY7v0WEtvVPlC1vGtn0Sz
OY6Cv+vkOygYlrbWMA8BzN/3ZD4Yd7+HUMgnvnTHp/f3NLmmc/2RSZfUbPRlRkBVIucKI4Vw5grL
hAFrpMUeqsaGN0tMcoHK0DyRFhfgEOJQDmG/sFJ61HGwsV0qKe/0i902lSwfuIFr8hlKZkWqvoLf
BEtyNdrSSmwrB2w4d7IjsbChcQfJQ+syS+T57NwvOukywFFA9oLcrmEFgfKK+QoKVLqOjiVJKQ3C
4RPhYhaD7/BqstOjZa3eMbgPv51I2UlGRx1LQ6x8SURp22NRHCobjyGH3RtDEmwSwWk94Gl5LHHU
FMiDEXCPNI35Cm264IXJFWgYsW7OOxFRQ50xyTIeWlAlZeWIY1zqKojGM+aUOyOtIIvquNiAzNj5
gM90jg5+mk2hZZLsiCHSQFdXA7aAPk7WelyPUi6tGJ7zmLYGz4ZbZfbMpwclRLoFHJyhwr8f4/m6
8Kn/BfM42XFTIcqxDaHyXgnFwjHc9yMpqZhfOQvy/Gct5E/111gE+KkEu9gH5lSBtkE0TQFGVZ9B
5kf1C4CtK//N0PzZjI+SQcBJmW5vJauGSr99o8KAqRMB9dqa4TvTnculnycEI3nUnsM7SBPQoINs
fzCTS42kuB0cQ4+aOx69xdNcQV/jn0ezIvVWJGIoH+31+M2hD1hbZCwxHbwpdFBIZVYr4icj5jRM
/cbyZ4ap56hh7x4DuL6H1LlJmYM+hjK30GwRIt9KiDRq0S4igg+ssCZSP4nsBJOXCVjTMTAfdH8h
Sc45dIYhMq3cJIgy8ejPgracRuSnxScOWAUUnDl7r5Ad1bdvkipGcHcmTAGF3SVqkRd6rmc1HbAp
KutQ6YNcfi88mokeIcol8WcVr8gNvtHfAQzFnVeucxsuGtafUirn8hItqSk96uQdC3rEXJCOT6nm
0LDLUK53H4z0hyWDbYovFsmqpGqbHdRi5AM7M5Q73GUW1g3X+GZZJRYnDPsx+Fbufll1NhbDaxSj
J4Xk1bLiLTr4/MVpTMGAbL5Ffjj8eLws5WTW2v+v7xgJj5Jk7KgpNu1EPiTNF0zz0+9lEQaLrbp6
0LV2YDSPOwqEC4jCm3zszzPxFUqHEjtp/bPKtJ8p33rZr8yffTq60TJNPc1Fx/T9sTqi0Ow4wd+K
Qw0asLrmnuEmOj2yfkR5qi2bJMLw3TXRDidw9PtChusTb9AW328LMUX5cbnHUcSK+Ep5IuPhugTy
vkqPUZvwAylLTyQtPxLKOllBA/9eBdz2jjH5fTAbHfGAxP09hgjnHdgvGaS3WQz4r3vvvNssmqHk
9nL1TSs7JA6z7gS2HKzQd4KHmZDiqIUteZh3QBTsYOy5eRUmj3eW8g5ahb1RONUZtHkHnMTtzbBO
gXAyyzZ6gQRAQvexEXgHhVaru7ZkPqS44PrEG5noBUwYPJ0fDnQtWG1qmUI/uwplnCYdAtB1dXHu
8reoSbSy/ckoeHMO//pqDwSWLF9ykM9pOvSeMhk/oeNpLqwdLQd1vzK4fQci0ycwhKgztK022jmz
uZlQcjRsPjSEDD9zXlliBfYV/aHhtBkekZCKDF430o4uODW7F3R6IkY7b181+5kG9eCwKsaILkBz
t74O0ceXNQQ2KXBDi5ZA8Ak9QZdCiCwsMoeVaTxqxMeOet4zi3alcCdx+aANBRRVRXweCJNabUT9
QYCYPbit6j4PU72BeZQhNORpyyP+9jZiSLya6L+9iLR6Wyh+1w39XfpfBcKXykTTHZjx64pOHHOa
FAZJaaMnFY5AwUS5k38QTbbV1RDL9h5Di+OXuuWRjIpfq9KHLMBo4YT0e8f/p0OFrsrFaJAt3Uye
LM4lYISVRVZyX7M3zd1VNg46ZdWJ/ee4KiRHBV1R+B8JfB5iGoHYPQOJY1cb4gciGc1XMNNXFm1j
Fm7y+7GPgG5aNJ1x24ux+andi+YAGB7kn+s0fa0A3YG2JWaAY4i0dM0xz+c1x6zXkkBJr3WvyvfG
dB8BcqwYQ6oaemsu2arRsrCI2h4/A0Pv0gcCiTALDehHMR+eJdBQpqspTK1xU+ckxrvBxc2nQK2T
NWQaohkJc3qsE8Y65yqIe1wuzvwigtcw2xf6ycyXO+/fjuNxkrd5eTNmICabDpMPZQSa3So75UOC
82G65vL0pWe0dsjBQaNZ6r52sgcZ+h68ADQKT1Mny1AtZP5NKoXCySeFbpwGkAPX5zLQidYPu+Cn
gJJUEjSL85fo4R07z69ZG8YpTa8aa1lluZeQkcCePQhuWGAs9OaiGubunzMrDAFkM0ETcNpEJYDF
O+7C+PMc/ZiaEAbsSN/Yq3XgHtgxFfF7wGqSV+zMqBtqwAg4WQeWUszVmGPvQOf00LC8QKxmVDQH
36PVqA9APiM7OSLdSCINCLQf1AbqC1rBFQ2iU03qR0gMJE3ElaZojo2f11WmkFvbTGPzqhOGMh1w
iGrL+OXbkn2yujASX8AnbdaQF8rndtX9654tyAI+QPWqxGH2RztLfAnaI7wqGsM6h6nuclYsdpug
Wpqcq9r3mBSFDxhhJLBgHHRoEg6Y9oMpdEA9t4m4l6Yj1emkkvVyF6itoIDk1qAyQyOKrpmGcMxM
ySDXPtfavhlcvBs45dEcYJKUuPcpgajHc9lfpHOHvDy4KB3B8mMkzl5Ul+yTxF0Ho2GemDClxpZT
gcrw7q1r1fxLUzUrP6phCkhzN3QauF2A0BTfHOalZfkij9ZRMQTQkLPtbZsItb6queLYSiFVdvi2
xLrMRKLEFue4KvtTs2a04YDg5rwdZe3mLiuDR8l0+w4RGolmnq0JLDW6C/Kga/lKSPf1/KXcSAlc
nNXR5k6i4susaeBFR19CzPCXSrc5LrPlN8Q6g1zy7ngcs21n+rqciCS8NrPu2xts00oGDMpkeChd
4Rh40H6HAmWVSFtnyekImXkgoqwKMDb0KPN1tjXzct7UpFwLh2Mu1F7LGD86REevIES/DECvPTOy
PLU33soLZRIxm5nbrcYAPI+xljHUGOcUVw6+vd1Pqs8vcaZoaCUY2OhPkAhJ1K8yMqHhLznPK3v9
ZsIRLrPJ8+6akaSoepH188MRXxaatuEfAxf8CYyj6mKPKzndfJgCIuWNdO3f3ulP9PL+jcAM7dD9
LGPEyDKVeLU9f1ps7PcbBdy0hWAjfjdecsxPXF776EXdrWT2QiOGqdsl+YG7qNWd21taopWs3iI5
wHAgMdWWCTP73XAEsvfiD60Dxv4KzkHlMQb6kd9NSoDZNakxgPcv2zcL9rVEyXvit2k10AIp7Q1G
BgPmFd90HW12OCdqUDrRRobXXQazXzKLHxLxIGCOzxKbc8VEjC3QtYrynyJwWYkgqRGRiusI2yU9
Mw/ALOdYrROD6McgUXmBpOJXiBUPPd5MGENHlpzTFomF+X1RypFV46BLvCY9UwrpmxNZCtqyXL/W
VdOZJowBv8HxORtehJt5Z7345I1zFTbuaDr8/S0M5yKs4jOn4MnPaemWix5LqmqWz9BZ3Wbe4IOW
xskEHBJ+reoBYf5W0tEFwgi13/LYmKtFC67FWweh3r7K9Q3cXp668nXO4muJYsNtiShP2317qrS3
BM0ESj+ZH8T71QbChr/KmwXUoD0CJ1Hi7AmfvQRaGUYggEAAbNTwQHMR5ADOjWRZKXbUo4VEQ8mv
91sg4HCDxeG+rHuoJQXC/o1iO2IwHiQZYhjmkeTQoKqGMH5ZGP3DciJFwVzmdA9BDyygDksLjL0U
kyk2pn6ImqSBy2/x69zSs/rcAN/JXZOCIvOxLzOAJ3znZaBElqBGLlc1yWYBbv3hfBaQldBkWhQA
swDBoMpvr8PaJlRdZ+A3qAx8YSJlJtjUUfSGML/jItaQy/4KbJelhJkVEZRoR6ohlBxXcyfXXF+q
c944wj6jyhBYqgS/KtXYGCcHw34OrTxzfIP6moJAv3xN3EucANkmhrd0wG8jzhG7eWPBUzIVtzoJ
OOHNb52E54kQSVGjoxWGAviJSFF2FTgqWoXXqlhUMhcvChzpOWhDrnNm59UIdMd96hsknYyLzDcz
cLS2CJcBPLBFT/Wk793KWP6o4ee2l5CuX2VTX9vL25OY9AVg9XvFlERUNQLDf14rnYEb1vlztDuL
uzicYhynkz33pBWFxxcCKTpmOKS7eoBvRXl9n91XQ2jchBGCHeuD0pAdJrpOnyWjEEZq5nfEunyS
Gi5lkWynrST3e1w+4Iv3X5pGKDppt+NXUxPGKl8mtEFKCM16id9/ihlT2BioQlEDdT+ZWio97uXf
7gFOOA1hwmMHsMn0zmsGTyB0yGvi+4LETMDOiJmGPugogRCTS6tYNboa33tr+QlOeG/gmrEQX4Oj
tgY1xPMrnqXsMSAC/HS60n/lsoF1FGOB2XQgHPf9t5Hh5lVHzEIBBrp038GUV9uih453sodJv6Np
zenX+IHtvJekB/2/903azZW3WkZc+5EkeBDI0q7lw6fH/nGgSv8H4ABVeqADqHUxB9x4HnUZbkVY
/3jVW5oJ0JEzTHb6qpsTowX6Yv5/0CzuycVtyXvMB1qVLkNgJqAh6iUo+06WYUD8ocglneDDE49h
QUtryRqRdLaPWZBMzXTLNPdyKvO6jfX1zX5S8gcAF9NcCpdHMO91QAyaMhde4pU9+q5adkb4/C3G
HoS+R3dHdX7lpPMZemc7q0XUG9zKvCsinvegWwL5It+YR4WTj4Rm1bYFrJZ4Tvl66JsdTouqEyOn
cStmWlGfMUOHAIi0r3xO+NOhz7+BVYg6l7L+QJ5A2MAMPJU3sFoLnzzxddstWE7/u1g3O+Qe5JAW
FYPRd5fwJLMgXYvAA9JMdHxfSv8e+U47BGOdtFPeDtOdLc1uPCpa5tnYMRLogW7HztoyYA45WqJW
9ps9dIH2ClL+pM0snoENLuq24wZwj/pw5mKkCx1pnZC615T6BxllOx3hCBk4xoaVrugYqrjClh2E
BDuNRZ3/QkkgIuqGZLgsspzopWNMkZ63SO2ciaDz18wKGrXo1/e/qRDnOTZB8dRKcNb9dDYzJ8Mu
ggcwMAeaygVNBkkcDsTTapEOJghOScCeimD6nf+xMUus2R9kMOnJigEl6lLQUW3KGVhvTIQQXaOO
B5VHywYA35bcumsbx5JDXj5l+TF1MRQVf42iVY2i991AZuSewDhr24IhUrFgh0ympKGKtphRi1yR
X0Iy04frb6otXObrx71wne50WcFOLqfFRWHHTgfGUeFUnxtpPO15piDb/h1K/UOcCx7ilHGnPNj4
piVdkle87ayLeEhCDYWUhbcfAPG0TYmtDjJVOHLbx3HVa0z/keGdBu+A/cChhR0r6/np4sAViY5O
3WXl/dux4bgPDpXw/Jn2deBS/cXZPI75Lq6kLe6L3TR2v4d0UOOL41+kOKhM1wK62gyIIc0sTjYo
59h7VpnnQyN7KTxEHol/aVTUxRaUhDWjTcONcqnp1jUSjDQnVFam/GdvM/4rlZBir1Rb63b1vthI
2WoerqXmiUkL/TjrGMWYOSVJcZ+9McdMfDgsZ2OzMsIOmle3mWaDwvtepobi8xYt9a+UdEacJ2PY
i09a8Dl6bX/ta/HEMccYo5Y0/Scnb22Eom6/D59YfXzR09H5ItJ0bLBh0NVkyHkbqAveQm8IN/Ta
/cZ5Gagm0uDRAUC24y+xP+wAP6mg2DJn9yQ0Dv4DjaPABAIlEuCS5DMztfLvbRu0Xk0HJVf7LJwv
F+rT0V7EmJcSeo+tov1E5j0hWgn4OfKGCii/5Vn3Ev/4Rv1D2XZsdOD2fuObzNnPbsTDb7N9SNlP
Nz5eGLWEVNGP63tyL1dXe3eyyCfhcNCJdLvmdownog20q4lC0qjNm+Q8wUM0AcVQYgyDv5HeTKqm
Fg0JuqR5okN6pOYbm9tJvn3JL40BC5YvPbH9la2eaBjkGuQFlpalzZGTSTxCm4mNHFV4PeXK6+x0
HOXtzBvzfLIewcae/YRrWgo24q9IkPFhatohiN1KI4s9K/o/i0j+b7yaSRAYe+S0WCQdio1Tdd1b
0XZh/VhZMxF8s2cIEfqdnVr66Uet8b6P3RB1zKotrpSkYEBnhHuqJlgrGgD8fUQOPepn8Y7zpODQ
FbymOQ4zBWsRjVBa+E1h45TpZEPfgLW4g+CORVFUFkPxb3rf1iYMYshILSD6dWjfeVKHyTtBjTe3
MIVlPKOwLEhEoPWu/30gfRvqk/SubpytCXVdfg/CwfvIkfGEgvSvRjnXVqv5JxrvmICGA4P5lxW1
0ROhGBXrEJYu0vuL2wnFg7E7vdfrCoy3kfAmCo6sstk3LcZzCNMhvXbglJGI1pCpzXfLyvrWHoyn
g5ypfWnDMMmv4sEvIl1i9RfSGuY7wTp2OdMvhvXbPxSriFO1Ek+WaScIgXAh7698ogPi0gYAHlXN
BI9nFKYFG55xpd2U1g3JyeDHDXPiShgxlJntMlRZ9pxpgq5PIpludrsWCZ1HHUnMjnyvGxX6Rbbq
RjTXrABg0VQRJSz2mnGou1ToZgJjQk/NAQZPZMFpP1MUoLg6pHZVm6MwZIcWnRVG+qGWBnUfKiAc
M1FizXJedDRJfXv+M7HhjWjY42gNAtxiHw+xcGpNy7gBKqSCfY28QZBLS7wFTMbOhjSaZ25rgo5N
kJRZH3rEivN9ZEACLlo/jQFH+zCL8/zeEQPq+XxsrSUK9l84lY3K0JPijTyfxHTZHJBG1daMl5EZ
NyDff0NVrPtJQ2ZHMgwk9yJhQSdCaP/y3UWshFMm4sv/jrVo7I6LtWCNY21oiHGihbQiBGNzV/Nf
tUQlClWdFXVFYWtEnNiFce9gCmjdaszTQFaIdYLKhInCdxEh+zDChiOOifG0OPPr6CZlu2fdCiOX
8NQj+CC4sau1ox65l+MLV1EXwPSqFkjgCJBLBg24GB+UTZL/HOJiWZyQuvkJql4S6w4WzvySoIcg
UTVGoRoQlJgJXNTjg768OUKNY6dCCqOHjVLyMVCMci+eQPomxauw9fjKCTBA7C0/v5N3CYnqZ+rA
MBT8dmwSsDtwj66l7UHSUJRbhJfvNw7o3ZNizQWtv+iUKgZfzAP8RChXQ319FyD3vQYLwWATTBLC
OMin9RTrB1NCSQ5Cwc0Z/Uq6rUaefk8/B1DHf/KprnH5YW1gXH2+WTJ0vOM7mVeH8fVQ5lCw9vRx
KRssXr8ZkMybE8+TvGPQZAjbeyQb6WNJlmjfQ5DTJ9ntTMbLZKlyOqmTqu5ZFXKHSaOTJGAG1oqR
in+OUizBYtLb9vQNZlDnzZsxerGbSpc5VkS6I6Gh7/NYEoQtM+u0zKhSqvobJ0VQnksShaBsi2bl
YXtLLXzQPWn5+9JBwMHZA+3vXNH2jEbPj88qFD2QYtjeWZ7nxzorTkWoEtXk4ilpmxDuRoPQLSqB
QntSkTX5b5pREp8PDQnDuR20OX7q14DYnHAr3+LsJpo6YJGjv2xpdOGXRkRyUteqqbn5EfbShPV5
M847bpl+zTErHzl/AJCcd1MjoS65tnM6bDA3n6XM4eHQT1JIDGXTXrYYoyaaeeRzsjWoEfVTgvKB
KREgj6YdH/63+i5B4zJSB897vFXvHgcc0BqHcoyPIkvVhpkAf/F6J8Lh1flJ1x/0Ij0vHbI5oO+P
YxObnFsskiJqi9pYLbNGcikHYMfLfANYws3d2Zl86wW5wb909cD0kIfQo12p3j+XdsmQkiwcX12c
6BhRLsuEWxIWmbj6xGuoKJlXnmbGQ1deh9Pn0DHUlI+jZuyhs+KJ06uBz91xmtweDKvOfOH6vWBX
tHM1k8GM0IDqW2Ko8QtZMEf/Sr/gESDsvh878zyhnsg7SKTRW2zYVhCKrASBypokBPxcGHOA/637
bhO9r0HWi1eld40ha0W1juzkKdD1Q/vlcI7OKL48oSupUETCteOrkxK8mGLpDin6jg6hGSUr3ARE
NBzYbDzgVkS8bThq+d+i8HOm+F4dcKQ0YLBaNhC1cVhRKD7avOmkrVOgxchHyrLiJWqpe4vzsHDk
ywbrk5RDQJ8Q55F+JdI+jF927cR1hq18hHsRKxjy2LzoPjNXbRgwI6+7LVKyfn+0F/FRYLZ3Hd4O
EhNZaqzmDELf38md3uBFXo2auYjhxB5+7z1rA0ztdGAPl2zLAVQOcAAdmBSJWXbBIKpuzv5qVRmD
mUb5+f3nOXXeK0P3t4CkPKNkWRdeLrhgxro5ThdNKaN6LCErrybudTrZvKlewWBcsHIbheqqAlzp
+YSkPNmAbG2xFPEhU6URMo0owl//YDTDWPp2w169KZ93PvtzD+/JSVI5MoVLQRAGADdhIWklXKr4
32OInOwyahj6Mbv8MXQrz2osUbNjbTpYFr9fwDykbOMTT4tJxa0RJ25nXIkNQjaaTYRb0syOEgSf
6TjubdFr5d2M4yxgKAMG2yKeCEO+b+vFYlDCyJjv1HRKxP9bGpI7jNFqIucdw4pIrbxtmYlPR0iy
e/sbi4LE0uyxR2S/63HSeloQQQPdNVagt+bIW9BnFEv9xkU2obK23stouY8BCcTCzugF1d+xndUn
mapYBP3e3ZeF8iJ+T9qoXS/A6zjqnQJdx+hKWQJADKNa7IjtD+H7UUile3uwlyQThOgDsKHgEI1V
ZpYGjMARczjIUHM6yMNThghBkwDaAyGMcR6WlJzgA3a66AUGQT/VeQ3bXt8miDg1wZ+deRov7r2h
DEhaxsFR1jQiw5nYnUTmeavWTbBuS++e1iUDADbP3itl/z82MeNgnh2CQjEYtdvxxk5vGJe5y/9h
jG/SPrX2xg4upJsLlGfTl0qtlKgtcud8fXlz/0I4OEFXPikI5Q3aBUiPUQUMvUWv1o+QZ/8CcOtg
/dbf2HZpmCxQ4pCl3zFfSIND+7D0UzR5Fsq/sBBFqM2hz5NcF0Rm8b8uDwpD1syMHG/JvnJacwqP
RlJm8/6DZxKuM8fGM7OTP888p5LqaH9HCXkgvi/DRVXXakVDdPT9rpCcLt51A8jy5h8jC/1b0pCx
uVRWYy2ssKUy4LhkB4u8jvdPQU5s6ETJKDpsZHPMr4czNEZfVyYaOnJaXI89g+tKYN/0atPnpfi8
/4VMvtANRr99hvoxnueQSe+di/Ul7A0OluOIMWrAuaNYO+PhdLYa21dXmytEJs79fy8vPkQq2CND
dCU4iEx4wnkbTn4XzJDIvD9sPQxVmQ1+vhjyX2GNK4e5muGOuzr6rvsIMPwd4eB+OWpCdbnG/+K6
gQGUFko8KPbM0dQlHeuQpxFYAvsn3qYLSJTRxhDMrfXCzQSq8EZRWtF/TQAkteF5TWUVe2sRNf/V
uXFxHGmcr7548NCyhE6Q4KaK3p5xCM565FNyZpAAFyhlU6tIkK+kU0UTgPgJ8AZGhc8ljmQfDpgC
wOyHl9kGo1fOZTMTRYmQs8flETfNlVYuyf7sRo+C5cwR2Kz+Y2zXzJy/RXECQV2urOZTx7r9RQnc
erNmHdWRtY+dhh39pEW7sQza+YbpTKhYcosVq6b7umTeiDuxObqjGsuim9hxxxa69HIo1/qw0Mvd
COd/6NPXEHHIKMRp7xoONA3eUSFY9s+KVU1LzZpKhzYjUGYmPg7zPlR4nJsnpStQn8wkBPsbXk2Q
IzY9TpMUCX6s/9bGdeRwwkNLw12xlfX+528kT5vJZEmphXZnSUKPCZt1QX3X52Vpmn94meSlAEN/
lDXIZgz/xcQCYnwXDr0aS+wQrWWSxV2Wn9GtCkvQ2xKBqYPPSZI0E52lz0ANIkqNwCYdNezT6qIn
wHYk4euSfksw17gV1Vo9qa4wBxzE7g2gOCebXBr638wYaSlQ2XJI1eTpppuCSZTqQBMpzZo7wm4m
f98kTCON/lFBmyFZEGV8BrRAZ20BUoPQiRFC3g9RpaT96mcBJfazo+e7vYiWoBFdRVQyFS2XZhbl
NENgKsB7paGV8WVSSivKaFMaSlsaHJ9k2cygPGEVjOBfrAVe9Fx3C3LAN/nZ8Ll1XMiTzxMb8rcf
sZWakkXakdolQSepz4fZd9K1MgtyHixCXyLVlzT3DmsNW4dtkWf0axxYfjmRAaGMZAqzVtX0YAFB
RrT2W7WUV4Q2/qIBB//pmHPGGkVvQAOaF/nMngMshW+O3ZvM4n+SXI+Ggzf0z/NIlIb1vz9BhLqf
+BKH7AxswBd5UnmGJ0JTB4/Qsj//gtWI4HUd+TgJMdmPUV15n6OnOssqQO6EHFfUxnsGV/OwJXyE
i+gSUuTNKeglVXWrAoYwcTOvMq6dQ/qZ8ZFRoiWXt0DWq2ApoKVhbNko+CPx7WsgaD8oEUXindcv
Cdzg7aRG5tHsvxqi+nOEB6nqaANqZKD3RJ0rXFyRu3PHSuC4e7/xH0Wc4eTfD8yxF2QRscALASvI
QAeCNWp3q/NdgPQ/o9Hw8N+y5sCVrAuyPVSKZxIIshfX+WF/I55SwgLzuJYU5cS+abAf36RnV9dV
QU+820w65rk5ByySC7wUA+KnZpw1OY5P6VzUddTN647VM8q6pOyBYj4tLJjP2c50uHhvwsAmVebp
8Vkzk9N2MQ0tJGAB5Pewz+wpsQlijBrNCnvpHDXpIvEMTDwF/KWKjQu1Z4V5y6HrByKZ2nTDzwtQ
3Iijh6oLKWyCXEEPAxswef/NwkVeCGje+Su4Ll49DCkcM8D+b63+zfWLOIwu08tGw96m2SSaNlwR
ow7LUfZ529wV8Y26ktRUg4fVa7c+xTaVJdeCtcMZjGpVwaA1mzKuq3+sy4nfsSM1CUYbqBDaKVLu
JMbevugyGeKZUHhiTZzpKjk6ujc5UlIwdJlOgqBAoA7otxTg3G+y3c/A1yUmp1NlivptYt64MMMW
Dz6mkoWaZHeZ7IGH1a4xXEkapFQHJxx90cKP0nF7nAIQKMCJEiqvwVXnfCAyS94Se80d+T+YZI2M
s2Rt0Yt7xRIWUqfTokkC7yMDYX0FeDmZJ4FX5IXFcLh3eHBMxbNYUxpesHSv4Lwp1N7QMCuiTJ/P
SkoAIZfHLhSBTLdHtybIAeOfdVZJAOmLCpdlqhRwoXVBcRNUXX2i7a3uI9pY8dkkNy0j++JcCj40
O8261CMa7SHUTpbXE+2tr5iN88Zw7c8dkNArbAcjpHbSmqAZRDVBThxuE0fyuJ+f5npiqxoSg2xI
bRhSNUhMZ2aVM0rEinmzGgKsEMRXzgIHfh7jcf0g1oHWLYIjV/tjz6O1aI8Brtqa2KbbxfFwg91a
ZNEgPUw2r/odIdtYmQYz3zI2C+wFZA10Eppl6qDqPpF4to3QLG6zSEoCOMh/YSCeMzZKpUwFTnOT
D+ySBtY0h/DMMC5nOWKRQZWqH2r0P3VFmS4Upi80clbIwJyMuWBlv3iDthi/HpT1WZzXWwXTiIeB
hqDToJ5J/PNRYrnQ4+Vr/vNCwUwqhd5G/3mbMlsoqQIVpUA9Vqqsu1xd+CWJ5N88I2HB6yG8pKmV
Cg9efFw0jNczgEqjnKLZF0NelP26xdJEJwGiZSe4A7W1FIxYSFXttDRWBuN/PFJllS6FfX1yZdny
JpgLNX7Y+WaTHrL2FZQjJT7vBxAgeYwo9T0HsPArNpuzjv8ykK455NcKwk8MmPT7K2ysxHyYoE3V
3aFn+vxGCBFNjxXTx0MXOVCT0/tVvxXYpGRfpXjdiXZCzIhZxWnZhj9W+5nArrLzU92X3Gx9mJU9
E2bjhWFGYxEqXDJOu0HdZn7UavV+M0Vz57tFmB1WLBWyI0/EEF8BCLTS5xTBKdYUe0ZLlWJBfYCl
WDU/rG4DWjnMCO6UFDkh1AVbimLERX1oFIUCxJAqtkuSi7aik5urf+1OzRYdiXgPOzBRxi7JJqm4
P4fb/y7MBmiEj/mHcx7gIEJQRDTgLSJV4KZAzcQI1WpMT1sm3P/3zLZLjRwGFn7xbCP5qo59FhBN
VYriy+aND/ynJ2uNSEFNnh3e7E+W2uZnLE2xqO1shFwAoqXNmOajt4ZnaEdkqf5dY6X74wv1FZdF
uewypJxl64afxwWud3THuq2I9T6fKwUknsl+y3SDfRGDPHeM6e+1f8OkquwUgLmpoVBbgMcuPgC9
kz7ZrM5CBhCSup3JtD2ZOk5MW7922g+fTuqPUkoTuN/9mToLdKIRtBS5kUPrnNCnLcPvo3pfLVo2
FMmInhpYkXMlZEh//VxVbip12/P8zNijp3B0ITmiPxRdYBbb0TdYTWCHAXVHwOkdW3QntjmcbrdV
JUBe7oHBN/SXCePWWyzCQlt0HScQ3qJrs8N3jWcsQnvLnNB1gXwRRoWP/ubnk9I26E1KdUNwqqek
gb+ZFcBN4E9IHk7SY7VmPKp+NJTgE2Xx4d1T6QrsO4YS/f8M3VLPieP80CERx6I3Voq4eXFrlNOU
B+9DAup3Wpd3bba3bsY7v/K6zDhRLK1IQUX/FfC0h7AoTBZT5wsQKttOSix8T0K1W9e9pXxqyzS0
jJFArpzr2ZCBMmW2lOp74+ZmHlIJWxHc5ZxlImLWjnJCsXb4rmXv0Lea2Z33KC+fmmJoAniB/YDa
8KWoa7c4jduvXZA4tEWgHtJsvKRtL/2Y/t2b8Hx7hmy8TvOc4MTKDexvkSECkkw3wP0+oWY4koqE
LI/hJfHgnv2bPelGS+pL8FmElddRO+vHSdHYaKaOWAtduFrgaY2FCMaCV7yF02Se57/B+kg12aMF
38/zyjNxb3qlSxs9q6iVDV+2OAk8WEEZKM09sWiKeYb2LlC8B70jvlbv2EydupP6jSmkRKozej5V
3MwCmJ/rsnkQ85ID4J7FyepeXLdAzZ0Z94QZAI1Rb8tw7T3BWZ7Cw4nHTkavzkBld06BPq8zQ0e4
//8CP3T8zdNZ71i99RCk0uOJtD8ZvgMyWHeZk4vppcNAgod9dAM9ANjxYhj03+43IdFwd6Nj4kmi
gBFscPDw7FyUcdSXW9vSczi8DhL5RUHM3AJlOkHFk9ClLA/UnCngXiJlfvw25qwPOOVEJvl3ARVP
8JxejUGCHQUg45uMvRWtTkE6OOyVnvZ03h2yuqEu7VyqrWtBK3Su5EAcqKx89srXk5RZ3xGIZHc0
7JiRmB4+ia1eK6JxL+nf5+/QWbmbysSI233hTlwq0+t2fqLpwdGafD9LCRgVLQQpNg76Uhpv5zjC
7qd+PNXGeaSHNLt/407TREcZ3VhTiiNMhJ5oVFtMCv0fjmONfrdcS9240mE0+tHzaWgHnECyWjEi
b6afDwM6SQ4UFRa9sqMqwkZnHAOJ4oHgngSK4RrnnduQ/yoUYDUnXFuv5Q+MFSdpkv6BeCQIyQUd
6JMxgJRpgOl4Hy6EsPAz35d9NHfrFAsvT7bS1iriHMwBulXy/xQ7+QSRVmnjKtEOQcpanZGLIqcc
ypUUG8qt3V+gmbdMqzcPVHtQQHXoEQRmzZ6hR9ShjFwvwk4W7ppEvaUKfCMYqnlDL7nZ34LY6DDK
djIRLsYHv+khSPsBicrBpFx6SK5Szoqcf0sXxAdESUqmQcByDzTIbOq6nce0xHrYCaBbUjDQdIlD
Hjsg5TU/lNh5E077WmRMbohHF7gqn0NTt9BD1MWjUBZjo44wNtngZQs3sh/hClvTfO9CFhDQQnyN
cQl65djQaBdSiBW1xw0rJjxbS0JAMcPq/bTl3gBDD5TQoQ/obCACa0UXB3tdmYbkFmW72sJNhxRg
L+B5mQFV7O4U9FD7xvLZdJUrFFrA3Oz2YWLo/g4f86TDXu1j+Gvo2vL6E2OqjYFlGHymd7acWfA3
nzar281KxC95gynNHzPd2OOM4ANK96S4QZs3qV5yOe9jSmrvAHc4sSC1jY7/3YiBRBXLaLJD98dM
xoNRL/n7mlJpyrC57QqfdbAFDqKliz/V+gJQJ62P/EUecpmE+IcXypb6ZWaxTRTGvXbvDUfF03ay
LXMZem04gSLQ5L05trr3pEi6ThAxPlvhJH6ek/wjM2Ix+wFA7FJdRf1Cps2b3i9HqKz+KW8Xh1EN
FY7PozNUkEYdmYtOtBERhrgqYogK2wrMIu5tX0nAHjuYJhNbdW8GhGwVZmfI29I4nrfBCs+WQwDq
Mzc5VOcOjH3reeorz90gH3o27mI/pQGQgcYLJ/3rexZMYE/4ZonNh5DJUvGOj4e6HXDVcReAjb/Z
ooC9NBlYR0FqJFBbpTruDTtfNK49fip6coJV7igD4CZFKi50qPzgE6bvBJB1ofvIom+kk40v2/pN
3zoz4WUunRKEbk8+Wqb5WsKenxgkoKqcTx4DpQMk4JXMziGxgag8fz3FTCIWAuwsDcU9/m+Z993R
oMpLO9CH89pk2OfFHvX+L4dm9XKRTyzzwuMRyUC5qWU8d1cubf7b76K7yFq2h1sPh2RTAb7nWPlB
o7/57t2zCufog2N+meXg0BFPZn3l/a8+IjUciIzCY/tZetb/S6y11bPTjewJoROVK9mF5K6Zvn7z
0baCz+I4oTj6z2ei2rCHMkA3p6lr2Yk7FEJyBpe/YlJK+8HMLljaOkgeduyjLv+HKrAb37tzUA24
Vx1NWR48dWC53Dxt37lRKoL761d2f2oHvYbN/a6B7JqwGFRrzjStIH4CNiyxVSakdsEidOeA21e2
zYDqsHFEX546lS4C8WRI7GMsfSDL5E99gTE7Ztbeg2xRSJgfF25UwXpc19g4c4DW0vpDYakhc70N
q0yn7M90uAZT4i+8snPtNCbzeX9nomxr9nzousB/5CQ9sTD9kYmxMJ56rWQhDTDhC4ik7GQDwUUE
mjFiOzRAFNvUpVWYfAGPLSrzFmux2Gacz4YWRLlECn48CUBrV3GZHjGr9ztv4vUXPqzLCRm7E1O5
IMours0R76obz+N6VIfdAsuoAtaJ/WK1qecXjIJ28dsrysbr193LL44hG8mzOvpzYFLD569/JtxQ
U5piOn9uMjQ6waNx6wUDT1KggzfMxbTE/kFRoBuQS9bLMJdVeZLHCkMSKlb6+sRW9UqyYFxg9iDt
EsK8FkIEy6NiodF5DLTw8n/gXG33iKs8RrrT1g/cveJXJYV3T9mEye5jzSUac+SEou3TBQgJHUA4
5AsSDfp/uS0OvPt7yprkIAt/0cP4E5+7l1k18zdlP2Atlzb7AiUQtafANeontMqt9I/ik54Z137m
qJMK1VQchW883nHjZ3iVLRybn8bym3tRH4U2/xGb6iYcdnO34rIxj+Gqk7UyWdw0QGKfHo4MbBwg
qMSkvYk1383CBAekOMpSoOHSJ+SOmUlv5dbp1TQxlRM7gIEtWFNoo0HRbw+Nua9/G012qgCtY0L1
kP68COL6zYS9ayGWU0wWlw0w0ZVIed/H88GPOzcl/Lz6UQ4x0PQku36q2KeXc9p67th7ttzBenwV
CbFSwZjWPF1mZrl62Tu02lPPbI+yYjgTU/a1OyWOY1DPp1uBS7TxE8v8c/4FboNU5rlF+jU2TFmP
ME9q0Bcl3wr5JbPiKYxjWKE9WnEiQHxMwMK/bdiazHev6S9B1YY0g7fsvMyOjCgrF8i/j57R2N5s
7w9sp0eEIZ68kSpLe5ocihYTWme1n8k2OEAmzfwUXc+CW2aJL+JE1mjZiQxUCP0GkZRKbGmnmUJb
1CrvgGSutt0KzLX4KHCQNqBUnu8GprgZmZcScT5y1e16X4jbd4qAj8pq44R51O0P/fN1AVak+r51
/SGJ3h50yapPpv9JVLdPp0Vh7Ui+6dSgrWZJ2ezZWSW1k+/XTkKWcZTXdeLBhiN+KaewJ6l/OFXy
AvPRK1m8HrWejyCPdTqJF4gGyF64H74vtHa8ojpGeyqMG0a8Zw04VliWSUlejtiD8rfCCFu0gpo8
O+i3pmuSWmACRW0hZXj5fO+qCn37ACexHaiRmSgYuzAwr0EaJZoomu9yjjjWa9bx2xdCoadXh4fs
zhbUYVhiBwzJW6SHGdoXf/O6Kv/Ca9v3AziarSoLxTUlQ09QUoCX4pp7+LtYxW6fopLpJhn0U+rY
IYWU1DDQj0wfB7DpRA4cdjvXyXoVi/FW9XANKuTZbWbb2/KGXfp6bCRiFbAyns3Y9en1vpZ1ZXjt
JlVuXJxAyC+r7Pi8eQ29XqwtuEk75/JYB+owjSr6qVICqfDac/8C/6oHUHkEvs5pZdlcNHUGpgdZ
aVFEr6+5GFiZieuk78gXPdILTpyvVGJ4uO4aINEYBGqxcBH+lxwHGbx2TrcYqzeMHv08eyVhP9Pj
fGH1OoVLMxLvjZyDK9PTHQHz4kssjjlq92PnUY0y55HIeJ59fYVobreiSwuALEjx/I0cKowASbaD
fGGEViFKhY50C19jjkjFh21bKNXF0Vwv0bMt/kumvTY79uS/pvf9eL9j8oEGcxKoJAsVUO3LeUfo
k7YxuS0yVbn5y0sf0SgyDYcdECALl7N+wjtHMCxb7JS4mdZs4od/HMc0h37D1BuBpQjJgCem++/f
RJnCYqAdG4p74L+n9seoIbIZDrF2vS4mgh7XcnPQWOOCaizosMZFwWB+0aeC3sm1qwMvGKKUpEPl
1kh9TVdTwE7BMuPCxWvX5ZC3Op20GaCZUOKZpnO934iOeH4WLkqi9//qq95/jULpJOl9TOsiU/fk
hKxnBgg5XH/KdmdeRZ6/nDNB/lBdiCjDlLVy5Pc/tkkdmoNbHU3EKG/OTbnd4EE+HBzhWFEbM5H5
nEr8wE0gfdhRm6v0y+h5Nu8eHe4heFFqSi9eBM8NcxLr/7SVpgHy4grD6UMHZFW4HYkdP/GJbSND
oYYDYW9BVQgMX0losfglY6gtnmcxFHIqSR3lz0/PZC+ZMCzRjIqHeaTjNbjvqf9yD3hsteIS1i0K
xTom8ebDIyL6Pl4TXUgZIPDvPsqzUb7Jp2hK4lCo+t+52bx2qr5vbWNFj5ibXmzOzUP8VeGc7xUj
cGVfW56T7stdCfqyFbfsMNc5eQu7iqAvqQYXNmOIp3uC92u4VpfiTh5CoK4DZXV5UwrcHEHeZXD9
gDJgVxXsGS7XSO9e0CczQ56hgaxCM4Q5iEGMEYpBys0FCBMT/g+wH73H66cCFH9OO12sGs8ObvHu
ZBxfBS386FvaEtaEkhx5S0NGzWq4/Pi4Pa16TQJ2peWKDfq/q6vkhq+9jL9L6qNKwzGqcg2AADwH
iSTi7uuV/vpDsKBMnjkdesHPsw8LnfaUIl67z18FXKihO1tdrFVU090KEsyb6HIWAG+lYVaM9h2G
2dLbkg69DwL+akOCE14tfZh7eiHrJtZw3RWcz4B+yVS/F2STvnCyLfJO5gpN+0UidKUzbJyFDIJS
Rtwyx9lduNLdTb3aeHC7G/YJvJJTN0BSFWyMD1e4gFSTxii0IAUQGrEDWA4T339N+wtP655Uuxps
ueloTMoW5n0TvpcIThE2XEryAlfdNgDFv7C4wd+en99cQMGDCaqIFk7a49wYewc1pDA3i0bQvHDD
ZohBQ8h0piVT4svb8EevIfNm8NpzVxvOMx3y7ZpQMe8NKL/YK9dUmU7G1/H99nvQALY6eE42MnJ4
rZzHT4D7G3NtQLOaMKv85y6E4OEfloxGo5I9p9LypAdGsCHHp/npVRV0o8KmuuI8Ofag8n7VLNR8
Inh5rc8eYYrubdS1mJOsgQMkY/r6YcQiT9yS7We2HvlW6uI+xvC3Qrcq/NvrsoU88f+Z1ytt5T83
vmDR3rWOkdp6PVuEDE2ObGdmgPQ//ELmaYtP3rRjtkgxLoczBtqO4Q7F+mVbc6H6bntPSwcYs062
ehOo24ObTKdTZStSFiTBhxG2LhFRR5W82mFPm7vE9sxRFBLwMuMge2t4VOMQWOtqDcMWV6GMzell
71G2ttb2y1gqcQhGMwE81OApe+9Kz/LC9c896uQrED0kcEVW12FxoW54nuiGWbKbJiM1PPaGvC19
Mf7cCdEToDRW3pLRQIka3ltT7sAagsMy+4dB9+92JRfv4rEg5nYS0MpcHgsOX2FmJCIdcPr6Zuzb
6+BUpILsL9TheUfzaVyJjArvLndnWqrcpy3NPU3OCHJlgOWLtDKiq3ttYyGXqdmxpcLfy3PFEbG2
RYsoUxUTKSRAqoAYKeSMLNChNssAEi+kjvlPchl7MDiBcTnPddBXsMdj5/j+WHcmtSujfXwJnj4l
bAtIYXccHxhEApGBwHp+yqqTVg6Hai7fKzTLHIBUkQA/2RdniyrlC/ytweubwKiiLvJ/gFcnWXFL
c8h1U3tfBe5TE0JyPetIwwMSApuI0dWuE5GmR6jY2cVxpvFABEoirSwBImyvZZv8FioNxkowkcGc
jB/bxRz++Axk9d9ajCkEfhUN3GkICE305xkfgXYpswoekzA4HP3bSguinMgx6Zl8BdJB9QwnJAdG
JIQa2Plhkwx+273yoXncfNfPkG8GS8ONBNLxGz+ItbqogZFHMbH3uxFjLCPXZR3o5dxBN+9uHuJX
sajEGMMAt1+iGCC9V+TEVmGqct2TVgQxxSyy1N8PKHpplQg92t0cKGgEv40VPcKVqOrsDF8aadov
/CWwudJPUE1qo652+H/WNiMIUs1+pcXP3UpIy/aljM2WhcWRUsfFtE0OZ0x32xS87q8qZuiug5Lx
kvboKiOr0m9dd43rxrMDWtv1yWpMgTsSU0S0LQC3kQVx8HqZNsz+TDWM6cPUYzBK932EIZOS0PWA
YwaykEye8101SLgjjU85Ms0V3iNiDY9uYcwB2QNc7gQlaHvbxQ6YblL+PMpO6L84WecvSAktdFkL
cK+4Misclqed+KeQ0kg32Te0t/zkfUwsNXIlTtpGzkwQIMopO9JullcemsrAPywNzi0uhU3+wssk
kEcqhU2cHOrAU1kq6/mARWnCO9ZQgCxIg7Of/+IfuinxcUkOh204CPts0j6tVzCf0oTRFR8+LUoP
el0aipSpX0Va7TNh1ZWns1Rkdb9nKX348pA9NeG3Ma0ijBlPb2jZKbWJgJmBIQk5O6hDzCTtYWYF
L8F0ZSDpZCU0q3ybp1NyRtOTjfY80XjBFpxlW1gVj9GY4JhiFvOUei/b0Lr0ESk1PsUGe/uIzie/
fzsqB8lLBibLdvBnot/dfrE825Keu4QtJJ6un8LiVNnrWo4TjmCibHa0qxY4cJiaaMWc1YzQZdXN
d6H/T4lm94x5WnmZuhujYh2VQpVCxCXPkzaFq1FMLfnWU7uwJqrDIXXJjqVBt0VukFXkOEG3uNau
D62ISTPHGq5Jp+2xNreSsYXv3UqL+Lv9YaAWR0FkqifWggCcR6jhydL/8M2KlHZsJD3gHO83ndkN
YQH4FRyF/hRLas2CQ/6hphrbhbda/QLZsVVkvZv/+KW/QMKUpyo2wUjoW42usWKQrIO5ucWbjKNz
IAdNXoFuU7M9A1qIcxIBuWtTc+6MTK8307br+xegbVc8raw2TgTJakGXIz32ljtRpmt3JluXHI40
aDEdsqMauFM7H0FQlGY3fqoLGRkMEAz0SuPRK0LYGUET94fbgGBRxJblJJnzwLw3oc7ARoO4gzCk
/fbVCFUYdv5HMJKcEy7J08hZso2jpIRmgfflW7IMoEMg9ueoC65DkZaYxyyYgCvIJzXNpLUjMrhJ
XfXf0p1OWXjvFzRCVMdo4VgQDFsa7EbKLQhNZEit15TFEiWhA8ydP+z+6el5tXOfI+cguQ7ztYFj
NgYXcRKgIFDHqbrBkqiT4fyUVHSjnxZftWQohIF8/OIVopJhNC4H/AZDoW7ReoeRV34hk3luHPOP
jx7A6CY14bzTyyhgqhR2IR97eKjyJjw0hyAMhhR/AjYkWut63Ccc4lxwW+hDekJExB2O5Ny6r6jB
0fCduXtNIDXPSu5+0c2ZGpm+C4HoyeHUjdnNTYydA1B2rIp4zGVaXjfM/xU8TZHK8AohezhlMW77
tB/Gi0N/Q1aI1ZDl81V9BfsK4jj/5nErNEGtdbXA1Kp5DMcz/4+pwlZNgmSAS9orcwFu5+W4wlXQ
ak+fb/h4SRsI7jWh6eX6shRIMbqYON8AVjx3hUCFKJW9CAU/+irA1PqKpw4Rh9a9J6vCkY+/Pk1o
oyTbIDiSCuGVwUCw4woZCITU8xJefb56hj7jD28Zovep5RXRXJ258XiMeohlWy4AtKx665kmYNcc
8Tmuc/FH+wGQPK1+VmKKAcjNJGTyjITpqwGDmCE4g6iVofd+IJN5ec51xlToenRxf7Ze76tTOII6
E0qPBeDms653Pk+0Eh3hAFXYpFgRAiRUigwOlHnGQ+B6VTKt0ghIOsoK805OGp4a7vkg0NW5qFBa
KK/ocl+asjkXiXb6sQsIN3H8nqsK5GxHZ43cVtw4jgls1Gh4UEqjq8KrBPHIlbfPxoHjWVJrF4hF
6mrbffwx4dd6hKLVKkoILng/UJPf2ICx43hnX0Y08y7meFIz4+mXoIFe6GI4NHaOBBWi1G4bHCR4
rerQ0GwJc8nHYIx0kaEiHM7OplWsSXuOcjgUTX4SWgjOqapGTSvIPRBI+8jdHwbTlbR5fuf0voPv
zeDsbRb4aD1v6FW3UYgxDPBjhtiVasPPhVkhfTyMWkFIktGToNa0a+Bu2kSxb23WM9IiWVHcvUBi
+vfM7J9PjsOPHSqltE/VuK7niGW3ETFzQIZDJxsZwD1tFIJ5tgiZt9Ye7r+gJ78AbF7eU1kaxrmn
hNZOY7RCiZsAUIiZSQPY9L5foTtGhZqDabKk8IgeE2OWo5nLrcVDLWkF6u9wZU++DzI7eCiqhEUI
3lyspsiaDuZPxlS5AIdvGrtAweJr0MS3gF7pMBbn7tNd/1J/nX5iTe8DbqbMzZILe1QEa2JSuF30
5n08f0hzePtUVLCuBZ3Woo4fKelQOwO7/4HPAHlPrlNJy2/Qax697+QF1hpJO88lLSO7Mm2OwWCw
r9Yylm8iIVaPTP1tZ0g+zMEvab9urmyKEeiB998KSFJbH734w7CAyu/N43YX/lXvHcisbv5+5Z4T
o4AQDcHk+DhiBam6aoZ6vEt5O2DSxUWNs+zs5JwuMWIL/fNZXN7W0rFI6P5TEEDfl3JfdMKO2Tue
e0mneCp1nfBzIl8/BQ7khJzHWFOgfbNYeyiHVmJr+zjHVgVoV8fyWsBdjQyV9lfVrLJWDAvpnt25
ACaZgFRCdPM+k3xwUUfFFuSZmg9GgZffmvcCt4ylyj+iNruhvDrIA/SfjqIDzdDx4y/GkIYfrWni
bP9tcDvONLNX8PACNRy7fOU/ShtJv7YdpkeAxrbGbys1gKj/NAZH8QFmz+8DUrK9tVynco5y49+r
gr6taxBs3W07x/s6E+BA5+eJdBVzkiRMl/xxQ8xFLdiItLyg+glQ4pnK5kSkXA/iEGZsW723l4hA
kgYz1QUvKhIvuhfr0gAkBF/H/Q5pd6VOHKCKv/GqZ4o5UHYafiuya4yIEP8nppWPKynrtY2MCEGz
Tt6oQdpGX5r5jjxpdcAaSBdgG47xYkW2tR0HlIanjC7My0uiUUtVEHPi6FcLOAJZ7QM9Ql/WTdKx
rQbwmfOnLospwQ/1Eyj10eGA/8sTCLYGqET3zAHc9hsHhxMgzNOWCHD/H0doxD7jCOdFYmvp8yOF
7v/c3vOmWc7yNOq/ZFiQcyFX5TkkpLU6doluiS/sOv8rwcVqk6dR/uG/iik9mKlMVHkOeLEFMyp5
deixcKaWVwkS8Dx7C/IWqtin/AnvfbEv6Y7IZFI/6/DFN9j/VSy4ZIWdXASpo63r+i4Mq1RgBPvP
N4evNHmPmmPwirw2nQ7qkKwxh+XzTYFWhxscdptheFZuGzS7vktkpDo8EzObihX52DVL2IWc0zcq
kklNllDjD1pE7NpGld8t9U+1/ubHzaD5MiNNLzu3lI7OLitgh9B9kyoadunEZLU1FjfBOki7Wm9K
indN7wBMgPGjuAaJ5e4hVXoB5efc0PI7SMMyNoDZa4gO517C2du4QPQSaEerQ7+yItOfbWHz/zSJ
2+r9JXAI5FEVmZmvpJu/X10YP8mGUg2H1EN7I7armvhjzrCF/U9fYNa1TAxQmzw0143xqiqLeM+1
srE5+aBwjBfWFah58YX5dWgxCIDucdLUZK6lsVWfwUx99w994y4LxZdFSgp1VdVwDfxH+JttHEfV
9IAwNQFOhMeCZBwKomBKNcvmhpmsIjz9X+uhupf6+4daHV0l+83cbhC3CHM01lbX0N/WAxWUYrT8
IfVNYewKDCrXTKFBJxUZ18oXwrnW47LZ+DAy/51z2QP/+Ex49VICkclv9Sdsm7oznei9g7gKaxkL
ecmqilLs5wTI0l9nC5EWpcoSfjtiKB4GbtBjhMfkr4AnMe2YRKhtruVQwzdbxD5MabwgabqKbVC+
2CHkixNplucdX4OzjgLsnelIbtJtKuOX71C75fUyBmHySbD0m+0zxN2EoDwZwChyVLVUobzjRZca
JDC+YeVR/Uyj6OydoIWmgML7kCXiSYNMCN8sIPoSU4omzXgP7cL/nUkmm6OyMa8FdbBvKDqoyxDL
7xiXqx17rVUkbp46b9VFjoDL3R3nUFMSEsknJbkfHE5tVDyaVPIBLtV83f3ACK6/ThLpUJGqPZwC
nyAygxbMdAIu3/pAtiPf4IXgXxxNCpx61fiQ21wzOa5vU9/bS/NnXM/ZZo9u0WOBEylr83k7fF34
J3FSxHSsOGWhBwsB2C/GDM5aOmgTUjbKZESlu/uyzcgXzfl86WouHTB4OnJ4NdNxpz/MRaJ6/KR5
SruRCWfkNuKFnotuYjGa+bQp1KWwL5j49kPQ6ENLwDWMy3Zqa82AHA9E9SDwxl3SRLxerT40p/5K
NmxoR1qwzxTnWN6ZQ/oeQk6P4h45LzNP51QY+DK3GMebHZfaRYsx5zKrIaLLnJr3aY3XaqhF3/63
6PYDHiqmKqGkwd2KYsLD5iEP1315VNx8ofpds221pudLECQiT3kiexF5QgLyqPvUJga7ZzbcXQCB
9uK0Wz9ZN0CKKQJXzPxc+qFixvr/AdDd3v9HLqGBwi2MKwKiEHoHn8OKHQwmmtFmUGubpqm0R6gT
QgEJJZOqXDit9CAk2oNwDTCNO/6nTEc/euJOovfIxAqpj4VQLfFgqmh7e1N1VKcJ5ThUjd7spqI9
V8SlOmMsGv8XyoQB1LPnZRz76UBP/FjvhG2iitQzMXlwRdEn1j5pA0V69o9a8Ag0W6x2P/kQZR2Q
XwrVxWeAdMYcjOnFDrClrthxHvoyuaJCp6TVKVhjgEOzDwRXVVzicaRUOued1UmVkAE1nwmDKs1x
cAHa7i+Ne0d0U9iNit6PHJVk8Ae8x15XycGWg7OacPT40d/GENk6lzlA9zjzJeZgsve/N1RxxtUj
RiV8c6s9/ArEoK0IPB+IkzXp1KF79MGJ38Gmez1WXJWncZcoTo1Og/y8q1VmYkuf8b74OwDraNuJ
3sIbA1MFbvIdCIIWS9v3Voy5OhwhJ0f++TLFeIRQnLLdDVn4jXgrs89MF7UjswmgEzfstBqC560w
DOQ8WNyWSmWcYRY81cmD3lvNgvwAccndntKxp8iCrPRvNqFk1rfwzuAucfvjjVeV6fsTtW5PdiD2
xQKMe5IQ8lDCJiLtfJaOyTyN/Q0k5ncRsSCf8nPQEhYRCfeE3XwAFvlub53sp/FMWowxu1SJNZnN
fqVSUVwZy/mYvotMXEGqW6Sfar9db3H4LOa/acZyrreXum4bT9UHgwN0R8ZhMHROQzmxWuHCnDDS
fkE7InhEoB1Rs7AE3mZx/zKezxDzRU5jm36M/Pm3tKk+qJXwBWKr0YQ6LvmgvoYKbTKHdYze2AEd
pSPJVQNzZqwQUOhO+h0FNLahbFz2URMK21z76HpNhr2tghMN8Re9Ic/pJo8N9v7q21mM3YVW29g1
/iYSu1Z6ODCygI7klMOOVzbkn0hBDMYYyL7nFyDyssnt82WKcUJQYAc2P579HnCCy+1RBOtzN73Y
sYHmUuZbBrsFtWWWnkmfx3E9zsrzyB4USlqalM5tPsXlJbcQlkM6W9avWS01ymfZ3OpPDiVmepm6
NryRXbo4wv61ApMNxb7CogGlNHqDhFFigRVNiVY3EFiA8V98r0wZknK3sSLK56V/FrFVa9WZTZXb
ixxJQeo98cnLdF1IDEgq/KPlqPaV/avuEJiUMLenK7XMv9zM3pve5y13DCTOwJPrr4retjhwPjVZ
tp7+Plx1k5RIFurHETfeLJDSEoafI9YmAuojcyeWADKY6SDODMS0S/Wn6XGEX/A3hMrCJFLFgO/I
nRNF5cGVIY7HxP+KNPa+1RW5j106gGYn3qf48eteMaoAdijFsGpooYrywOLrklQlQjqiNFSMWsjN
j7gomg3HLpbtF6+gm2HaB5Z9KSRLpiq+KtjG4JouxDhp9TgDuVaZVCQf9d577tom0kqggQSUNyat
vgVGxDAa7bdjCpI6qywSxXn9hcfUVywd2ZtT600KvNObqQ9TaHN0vd/uXIX+ALmcFXdHadT5EJ7i
AkR+p6gqcHTAO8oITNEAeRMEwl7vxW4FSRe5ElgpNFT/iOnkekEYAFYYAMJX2q1AjH5u+X9xKMu+
Msl0jhPBiBHLkBPXdFUxriw5nCFiDLCuIU8FqSCa2b6cH8N0mDtBU/ogp64/LbC238hD75Tf15b3
5nDit2WxT1JzwFYjQ6U18EbO26ronW9rfap18NkGkwroPZigIAP+GGgup1R8L2QgOcec3BZwkAb1
qQKu/5drLFvCE1id3oTWCcp4V3WhTMDiQdFhCNzW18BKJHOSDzQx7AaR8GOHa7UaLyILJUoZf/qw
YuBI4U393wzbx/2s6Z3ppJf0lwoMDTwiQbsByMimUBWT7pRkx3ILzLU4bNYyxN0FZjT+qS11F3mJ
E982Rf1M9aPhp/OyT4IHmwc5K1dWqhf7ddWcGFvdRq0iVNo/GuBZ2hXRsvuuAEqc+a47Ep+prAuk
QEoHe+oZDPwNIAMzsv4dwuZGzcwqDEwlm6BRkuPGedRHqcIGwjRiI6X84jacvQoy0EN5eS6b7qTH
OCOaRY5AYy0qt2SYAQOmxypEEZszS3q3G0fxQ0iC6RedOy2Zj7PlVhEIVXBHqotxCFd1QhOKYhw6
2t0XpalKv5dbrIuXsubqsmkWZ/9ZskYQDGC45fKjJ/cTkuHvA+1yJpIzyhCqbKdkl4nj/2r2Q0Xo
SruLKQEIELYr0kXrO1LrGTYqaFLmUL35nnLjD4elJa4QkYB+pFYZUaeNjNqDOA/gDeeGgaafLKE/
rrpjvmlJxZCsAy4oARgdNB2XdtxjX21WVrG78jeH1Mni/pyHIXVGlxfe39V7aM6EoPzLfJaZQrZ8
3Q0outIazDlh8j+0rPBgkjrX+K9gmJyDdX38dHrzCD7gxKluukQBknu2R5mxGnLTZtRmTtgWaTkK
c3VrL5Nte1kgw/95m2i8dzPAj+JP1uBnjMRAitRPXfDHjB3MIoCIXz70hyKIGDabEZaumW1OmpDK
BbjGr4wXOOiL9fL++ypZAPTJD4MdHVltL8R3DfcKRUtMg7Wk70f7KLVd9EL+SP1R7dp6DNV1vdUk
3N9/mHYufrwpAjX1FPZlqhOu7ftTzpLnvfbZmpFUA6BCV4qPZf1fsmZuBzD+x1yqadHdgM5WVDaj
epC4+JEa3NntKboAKmYQ9MlW50LBlEHwoAg+0YG9/Zz/tjr/0s5J/q03Kb4haZmqqr1F6i2OfNi4
fXoNEqfNAaAH4V5dFlf0X7rD7C3IkipmfLwtu7B2h2qcq8/gNAmu3qTTqHDbO7WP69XB6q9RMP2W
a4SqOl66LMpClVqLPhHu62ukLa2OkjIfIeB3cDkJ03LrjJUOPJU0y/LS9vLQeKcl6AQvT+BCLUoD
crpTNAhikGOGyFz4WTKDVcSHm98gaNz20Dbo3uTn1Q8iEGpRIxx9Z5RtSJOyJK+Ldq+8oB6SwFNF
BJoD1KGWDMmbgyGKu33SYiLK9UJxKVw+MVQfjJx3g/PivMlXycf8oVAlj1hUptU5pU7qPcVVxOqY
QQRky0zcrya7R4nOdUrtJhYoUTf9OXfDf4IkygzY0j6z9gKOSXWxGYl3KynO/cp6bR+venllJazV
z5Xh1iDhqdljBcwBB39neMF4b4EWWEKvKblOCw6BgZGP4Mo3sUYJ1LyjAuYW7iRI8wHOcUNPz7iy
diwC4zY2z1ucHx2kFuLnHqcK379lYWy/jclngkBEW/EcAdhnzlXN3wVAbEfrXTnZWtk7wGSqOYR0
KJ3cM7NYf2ak9lj71d3l2U/KkaHnopNai6RpMimLCtHgmmj7FUroY7y0uy58meUEdhk07W2dH4ZG
KH5fZqLaJpYlyLZXrNqHJoGBormb+lDpznqZQYU6yUjKIQZHKtDgd/WdKOwZR9t3re/Ensd6Cbja
jfefAS3wG6LB4KfQLxaPh0P6HLbnuN6uNv4jIdgZTPwHwi++E8ucEnSsAff3X1OlvbpN5ULBG/iB
1yVDF4VS5xxkTXbfJVFENvi9rjxJ03rSMpOD1JzKMdbnYa14isf+LK7iuympU2IZqx4+LZBSwPSP
9tDtrFZP+vXHOtwvvDx9Co7N9Dz9Jm2Gf0EifsU2aMiENA+TD4fNUm/PV1viWBTn2xvycv/gU1S+
yry5Ujccs8uf6K3IsiEdjkDY7eA7vYe2A1a2m7a9HRB/nLRI0j0C34ZuSauNBaFJ5jee+/JB/dtF
PtcQEXImJdGIBHRUr/3HRsVoXVVcsJqDeOWOqHEDasfQY9IJur3I7ysjq4WH/xFY0Yzo5LeuxGic
JrpJ3+Y1BApgvC9HdxZg29YhObeRNYkrYRF1AY6585dsX4KFJnTSRAepbeg4zr0nHtFXtaHs1EDS
jKl9CgSWuHBMn+rwrq65Ct7eArrws4dogWfIyNvJrUUJCnjk7bqsBLQth9So6oWy54+rAVQVpUyM
XPvSsvJS0OmPff+bGtU8mVPFMc0P7m4xqlDcaRR2mVzBGbY3f3/jOWflVndAke4XIQ+5bWvunyVG
xOmlLyXLvptNQBwdraxPlFB/DeJWMGnvabt0AhlTL1V/4jcsOSkRYAbpDw9dMBBTJgxP1eMJhXby
J9sbnxIZwfqDJoFh5x/bDYT5Zk+XbXAKWatZIT2MeB7msnA9eRtMsom5U4cNpfjlnQALglnr2yJq
IxSnkgU5XRcwSuwTDnxeT6+ym+a0DRiZlsZmCa6ff02QAgG0LuPRMYmV3RT43F2gfSQJewQ3aqRd
A1r4bCqteGGFa/FqCw/6N/nogpgwzB3hr2iLRWunt550gcvHTp3hu2ZT8Xeg5GtJFEBmT/OxyPHX
wNikXUWJXp4RS/VD9clqgXL08hAKbfLEPhMx8FWLNirZVsIfvAlyv+vIueRwlT4WMCFKdU5NOe2f
LGNVhjuYrk1x+A2nq8FrXRM/qRf/NJ/NL9B0ivq/iyQW6ApYvotvqUURQkJNkjzB/lFRo4nCU3mW
3ubtBMC5tSG+NEg+yYPrdA2ExZ3aGXFlpRgctGzexzWVpSheN29uU8aFcrYP1vsasVmnHpbs3Adt
qbdg2aDsByI2wfShwSRfMnbyHc+SfoU7w9mA4neZCteJz5tLg6pKCtrfYziLJQ9TolbkF9ipOznj
ChMsDxsC0hRrvtj8/Kxl4Kb1Hd7xn7xrDt7Pqu4x7Xx5UTATimAeIk+hzJEvbIObHwgfXG5YtCv+
B8xFolDB78YafNQq4/KX9ajsJ2QrhQs+96Z2lrxJNcWuTj4jRb5i8PRSCgfld7799tR6gY1Lwoue
chVeQWS6YRjRvJORYcFNTtMz0DBNVarriyaSpmHk3bo0s5zjjI7X19FrjQ2UO2DQQnnWLuo32zch
Op+oZRd+RM6ZqAxd2EJRyUMNjLWJ920hxcB4gcKvj4Q14zBmEr7qRImyoZ9iPviBYad7EuT63VLb
y6HvFAOwG6xP810P8yZsz524tGKHtRpny8j8MZSC0dUGHanG4onmiOboo/GGzNjMET4VI97d4o2g
GssmnzYz0fn3FdjNr059ycpo/Qe+V50mujtZEDJyGV/fnC5gAWtBVn9nVvJVW4ZKK1FJRz1MH5mE
rI9AkqypqyCVGrwKpE3sEuBlygDFlwIA3lvSbaMIcco1tuft+Sqj5VzsC1oxgIQttCStdFpaGX7s
X5iMBuchMAYeddbvSX4czAk0Z0m4WVc3U7LDR5hpLifGB61pMdCcyljRWX8/aIuNCbYOwGkl/S4E
3QA27eThpWE3eZk7M6Rbu1K+aF2FubKZYvgtJaSV3MNl9WUGUrU7Czftw6BN6Ct4dde2Zso+m8fd
XilhDKMKqgvrLdsJgHg+wVsEnibo81G5Pm8clOyvjz/ueGkOJMpfsROXcYHZxRfOvQbDTNq8QgJa
pqLy6Ju+LR6tLefEEENABI7OFK5cCwQtQtERuuKYiMut0CDrpxFun7nrEOpxjyIDViyhEHw14JVR
qofRw405Z9NjAPKTYU7TMS2gv4v1LZLOuAfYk3483J/qDn2JU996Ax9SdIFy3J/Cn3rc5qfb5PRv
mBOlCxezti+TD42PBds0fUvYsHAwTJc5RMjuVizmgtGsAzYjWrYP00cgYDKDMx/lN2wlnY9/nTa2
DVqA7dJXtjdQGuSI/dIox3x10OcnxHOkelL/ADkTqaX3q1XO3tCHtLfdM/1MK8U34m6vOKnY2Djr
J8JYAuguEVXtUlckAp9ikzgge3gKVdDy5X7iZVWSPX0Lfk4gxY1qCTciS18OiFNvplkOKgvn6YGp
HeWd+boKLyc9qqdtRz+ZfpjRAFTtZNOauT3N0rmwUnxIkwEMfH3h0X40dvSJW/XG2sgZU6MbyDnN
+ZLoCG3iCVu4XsirhE+Qbt2pE2cObWbjlwWaNTOiZU39HAMWqjjC55nwCKWEO7ZWzY9yBC5KnWUi
dhpGyO863p4xMZapyQv5Mkx9B9RnRMSJTj/3iZv+S3PZGUrqAfmFzWVLyLqiOLvQbnzj3k/LQ4M1
Z7v8y5mdKtOJpwdurdCdoqpKsd8Q+g+gm5JHwBud9cxAR8k8XOGO3Du87PhQG7zjGurTmjMn3YaI
ZyB5irp5ozpXH7vMFTJmucgEIdyJseEu2D+MUXbRO2hqxzdDZ1pK+r/Zw/fJYO2UO60u4CDfJ9Q+
arDph8C0JBpzbP7G1pI06N5gbHsOamDjiq11lvo1M68TWND/PisgVvHksppjp0TyD08dvmEmJ2ZN
zdnLWiNvOToIDgPMfpV8v/Vx4Y/+pvrrHSv9zDrgTmEbyzTVco9qY3RnyIRNc71fv38xCAUf0nmj
7zZQ078JjxUF4n0L7bfcgVcp5/5MJz5J8PWN/RcFWKXn7qi0kow6Vw7EHVEFiv9rE+qzbmwYpWEU
7PXg/TkKUeXh1xSPpllqUl5HdM549nuwOd9fRRKRL3MVgZzme7IGm3wDzLTBVrOFttITo0HDfdu4
7PZmjoLGCgX23wqp/bCQJYDTN2fgyyVRcShNMgyqbo12oVD2d4b2PktdR/2IKOWpHJ3UoGUOdXKV
faHk40akqVhNoXkLw0hC059DdzVfmLmCcZSmn0xAHAzmKLa1bipUBfkM+FgNbJlk2Ah23B7qRIhn
QNbv4HJFUssb/Po12d3Gqwj5M44GPAKntU/5G3MD5R7LJpBVUPRub3JdOb31hp2tvO5w+nAl5n+W
wp5SX5dZVmA+1j6h/z8UIWWThxqaCVvN8MeZQbqwqWnnkjiXg3/K23QJQHkZvF4WtFoZf+ViaMVd
TXFETzqpmWdCXxaY9rL/tFmVggmPCO/pIEHmjVuD32O8O5W3ONDDPr2rKTpPRg8GkGbi2TtpTeSy
f6Tx7BZOQYJiaeUx171HnE8oZ8XVGjgWame68Vy5ROOFrtya6o4i6/qgIDmMJjVg4qQJ9XWLWFSU
Sh3YUSN0RPhrnYjPwYjU+13RrpI5qJ4hM4ln5jWZGNdnzAkYdaj/T0VPajLpzVJNwQ9VY6oiCcgv
WNSlnMnNgVXCcvw4bNAqeJp0e2EPG8tPG/lLtz8FZ3Kv57RPLD3JwZQasiJxN1/cb1tJHWlPLb1O
PA5HWBp4ZUOg/PgnDNDDg9PDnSTln540B3QDRRgFJWLL68wHH74/oGhMTqSq5yrG16yG44Eh3ZBE
r+pWxXWauw3yaTUYb6uvLXcCVwwK3PnFdSqpDJXDs0iIPFoezzEKF6gyo8q4ts04ppPGL1Qgn4cy
R5baN3tJuukTozR85vm5N3D1Y/7HYccYIbbSawDH29QwBRhDNvpPzkqJg46B6kpikSarU73VFSdP
cSngbptF1p1hW8shtNV+2V34QdCmvaQuC1DliAx9WLigzJXVm0bF/8ep5i+Ozd9yg54Je5jttkMI
Bm5BGEXhfe7QvnMCTPj08BeBaQNrcT8At0mRVQEoRj/K4wOXE2q1SFDPTfQ6zqSvLe50iriYHQFt
vgzxLWwT5mraN9p1EJRmT9V+i71558ANA+j3uGFlaFCntFKVHFt2jjrHdgHhtBFIZamNsO8RTZIQ
njaKcmZ2bD1dy2EEjtlQsw1LTvb7F7h99s3Vy0I32rrHlOuSMJe2KPXNS8Dgx+rkesqwBaGVzIYb
O6XQj0E4PkiM9Qhj+IpVbEUcijoVCul+OfwAxWa9wVThMl0r58CGJXP+z1iouzfw8KjncF1U0L6A
C9iom+9VZdSzPNy95OixbgnP9gQlvD3IoBXXe+lWJiXvOk4QeLWEqb+iCqJGmWn0e5+NIO21BnZz
FulR7A8giiyw8E3XY3rZsFpNNxRw2tLtV4nSoMTIN6Bli/tx+71IGsqipQts6VOFLqTHXFPQPh2C
WnvjEtKSw41zvE66A38HsiR/rd3EJmpuKtA1HtuuxSdSHDOVMPEfldmrquQtCd3B1pHnrY+llgsE
vVQrOL93HcqaZmpnq4x46mik3JigeJEaaMd6O93n2v5GHr5iX54OIUS0AKybOGOW5dgbigPF3l7u
W3/JQci263VNGlg80WtI7vj7oSkunPDJbTCSLQ/KmGrz8jgw9Wpzj/dt0SFpn9f4c/VkVtjh7yRp
6Ms/hudZzMtsqMz61wH14hYjADL3Mm8hyDYWc1QWsaj3ZxxP88BRZHe6N7pfyiTcrvkHn9yQoo/d
WJRoKr/UAz/oz9yrJvRPZdOZNJNDJCljzM6JnCqC+cz6XqHt9Bk8b9ewyDOMVSZ+z+QU46qC1YJr
M5OaOyIWqNiCbJyNheAl98fntE6dLUzfJAdszVC0YL6j6TLCPVINX/otMxldZYmHkJWj0wMwAwi4
rzXJ7Dy51pkzl3ZtR843ezGNKxypsUvJwGLlo7/N607HcJAz7S0PPpSsefVthzjjxs5io8hhzB3T
qDgbisTs9wIyVJIzRt4dbvQACPKo5WUOfuWGLgbif7vmvCTTt9MbhvW1GD9EZG8Qi6uhdj/yPx0R
ESnJqwY0EwJ14ebun2WFcQwC2UlmFPVsUTHpW6yx9glWwV5rq2+YlS4mIZH4oLyCoiJtOrlI8Ibt
73wD8pTpNJcAVxPk3ftP3YDDt6707OtvcWw9KZOhCeAToF2DHxvrbQzWPBtwKM2JBHi6fp+ilV2B
/yT9vMIB5HCKv4AFFM8a5FESpcEEEvZX1RMo+QyXL/Gdvy2dO+nR5pkCQdIuxB6XmtXEdyIp1xHC
bIwKIadZd2tGHLXE8Xnr54ijW/lTxi/woWdD/5BIXedBXVvGixviUf9fNZGlj2IXcynU1GoDL69M
wxRCLxEZcBfIJ1fOHmMSGVKtZqAR1GgZqrdKeuXcNKWxzHNEo2m+g5/9ER/R8UoZ4sAKGBq/biAg
+WvwDVWwh5GbGi95d8mXZYOJnF/76jFB9chJQJi0QE4MF7EUn5smh36M92DBxcEGCSXATJJO8X2P
xqRZmO3qcphSaKFyAzA5MQMbXkQzhRimOmlY+CLB+vBhSHTwdp9rDVVSzRT5mp+wx1jhuoRGUFK8
wH4VdtCN+Jjc39eYBPaCFlzxoQlGFxZJ+mXmxR/sPVT3D/DTmDDvDuEcegF6mZ3KlXkd2vMTralt
buwY8JG4J9mYvHtsPQ7NqYvrEPvpwSwrm9tm1aKo9EdJPiEKAsgZIgHwlq5R7OKBQFPAACcSM67V
xE5LJgHm7bJA1D4is85ZzqXupwfI4V8y1ky+Oovua4yI0Hy312bfpE04naL2gtaIzdsMKw0VXR5G
Nn+kmGaJGsV7qApKM2F67gq0luvLCj+/MAp3CVJTFZsa/9kW0V2v0Y6L8mnzHvRyLEu1KL8oQQlV
mH3Grllcw002P2bapxN5I0J/uW6JpnDNYe5t0+9OPNL6egUUK5FGRkARjlZCw4L1mhSEEaKOsAXn
5JgjHA4rC8aUxJ5tMV+gTmWF4s59DU9VH+i8OdwYrbnF5q8s6AceHdNnQTRL7bgrPlBSo1qj9J+C
BU47au0jFBuk+tz3/09SK1kNAeAV0A7TDbdHXawRNBx4CUJfk1zBa8vmX3uspMrExzThe/4Wikmy
MTzmPkGkI7d3zxGuxfUWL9foOihcTnsJIqE0jPYI3ZPXPBSP1RD88o23P25wlZFdPlTuVQD000ro
giRFc328ot5l37hAL3NUVIaHqPDOhviO32s1Nm4syGJzlcYxoOQSE3Ow2rCYjruxhXt7/xJXi6cQ
U3Zp1nKxIfaEh2M8XJXzm11ENtoUjG0qMp7G9P18AE8SRJgOW/q5xfU4PMWIrjeb4U9gmI85uslB
/hD37ao8f8OVl3X5F3hkWe69b8UWYD57sUbgwb+Bg2tbfFqwxSM8umTTklHyt47POL3ajtdrYnBp
PnKmeLfG55fZp3RRFb0+IvtdjoUV71CFu5q45GBYebXauoIqIalQ2twnPgBshGmoiWYXjtOMJQGi
PR3DTT6bu/WoOmONMjkcULBDT1c6aGHZMYlvwM82grx0MhV6+jVnCPKgcdXJ/PgAwr3yDXAJPB99
nkKq21SGUZaztKchGAw8YSNeRorAR7G/bqFX2hULyVh/8r27pqQKk8jgG0aWM0xp04E+P4OJSXWh
bf1ZV5l/PJiWsGRI9CpW2HP2e6sTunzQLJiqnsQ+JluJMXu+RpNTxvAT0xA6puOYzXxs+cyPEKDa
CFmDmHZH70ynGv+qbKApyTIzwp7JffaMrJ5IkaQOrvZpD1uiKUw3lcZWTz9uRWFNTyg5FsrQsplM
DGEvSdZCwUL9mliuRZglFkvrzEPzMxr8vz93XFPU/OmwRssB6wNWUTt6OC4gB1oSyC4ynLyHPc62
oDnKIaUL20ZpPRa0YdyWbzGBKoXkZoHW7xWM2br03vxHMcefglfEXbDxl5pOydBHBe22ir0+PaME
tUm1Kk6cNj7sUYZrKcViF71WLcP0aq9vvpMIehvbd1M5fg1+IYUK/8FQiEO1yRxodZiH6ZjfZ9/4
vLlaum3psYJom+KyYHr3kuhTsu4PgP8eX1paskZVXcO8xIONz9tNmhd+GknOQlDdkC9cm9MfsUPh
dGB805o7tXDkLBYcRwGiMaetc/qZeG/L+vFi+y/S2W6aENoTPHkm2etoxrvmXW4oNhe4vU6vxqDq
Tlk2ga4bLGSSq78g0LQbujIPlSpQ7iAHRPI06DH8lmZG4WidK6LZ6CKuAQL6I0K5M88WR8Vhe01h
iXTLPbc6q30yKw6RYAGUihWFxDWltXoilRlbfQYOGHDYPsIEQ4MMBZc996Zvnx+K5W9bbp9+SoGG
7CF6+DsImFm83Fu4y9b0BkyFjsuVtEWbtvUtpEetcjLJ9vWHEGKvNCh+ZuXfgEyV597pyNHKH42R
Ifjyci+eh7215x7zRamvvzkSa5Ghyrzd6jD84xVIvuRdZcYyIG28IZmpv7sqLmLgi6EiMAH+wfBD
NbVMsFP56brQV/0Kl0BwGJcKClpzRbPopbdmeI8O58DAEoMBnbvc4lV+sEi/I/pEuNp/Wkp3tgF4
rQ6C35RkzddPiWMGqFKM6YsZYWBror8mKS/sunhrFXuX62CeFYTzH1KO83ByTGfloKr1uTJODaqk
7lSBgSozClAmV+qzq0Q0S1hAhrP59pcBEyxNAH5tdvjq69npzL18G4acgeNzkqz2QsH8trLM3Cwc
90FAumsJheiQ0nSzw0CAgmykIr/SU+rbdrFjginC7uxHDQxxl42QizORw0OyGCUNfkzcp3wTMd0J
KkHKKg9sThgab1ZPP3W9RAKDgyWCCnfIAemo2euohWTCudzSYJeJjxafLJEHNI6YdEAl7IgT68s8
ziu94JoU73+YqWI5A2owR5EQDsqIs3HBvcIzZMLPAcRE/1swEACFycTy+ugrU9G2ZSdcjP4dOclY
buUl6QP0n6mYMxXNnnmDHvJZGss4+ZyuIfQBxlTUw/JrNMq/DJrQMitKI+YYzsI2JGee9wvpzGC3
Go+KziiavelmFxMuc2If0WMvNGuapebrcblH5G0kKYWWz/jDxMvFE/G1DnxJTCQkCx48tU0q9RrG
L9TmS6G7M6Ev0ZLooVjlpetga456vNUTnsgI8VA/acIsules8km9i8W7v5MVJNTvCcqkwiWx2A+g
G8XuLc1LdwmD2DzwoGmvbE/nxmSLNb6A6b/zbd/k5AKSCfeRwnYB9OxG9aM7D7jbZwMvilqpQO+7
rIj7tdlEjNWq3//TPq9TVt847X6heAWdiCnwMM8Mst8+C5Mclyy62aLY/d0l8koUvUXB832JqV9R
AO92frKTjXoQOMV1/YC70iFdlf1bpplYEbvEB5HACzru7mDCIHbif9YMFfMMrmgFdSdacHMEUT0W
CKAEmrJHLbiW9WwpJ//F5/yQQSpsRGXh0fbONk31sYQR/OpOXFUhtz7mlg1lowMXLTRlBWT/1rIA
gbFv/4E4Dyq1oWV2MCb2aCnfWBSWMFt/J3XSQzx4I7FXfp5ALm5kzi302ePod+2U7MGRI/HcjtMl
jV52hdUvaeCU3nPzm7fLkrJhKPZ2WpScoZ68EGgaOGuQ1aKyDG+sfsPjN5SJSTfLpTYhBeDWoTxv
m4A6wq5kHR3pGbIEkNT/VWMXSzQiqZZQSZ+t1RLJqPAyL3sEeJAK6AN9IxZewqbr2gKMaE1u8wR4
IuI1Uuq5oFkUuyk0qhP2MniL0MRRfTZdAFEEH7KwT9jd+imfCsELdWcvziU6yQvBFBx49fTgbYhj
CM+gWrAxxWiXu+NV35Zc2cOgABByr6NzGMEKQqUPTbbPEGugzKEbWFu7tlxV99RTwKq0KFsCtNfX
XQ98D8r+k+Zlm67fNTcQy0GQ1SXrOetSSdlzBHqi5QfpNLWmNjwKTTeCpFYUfFczko/apqbwkGW/
oOqv7VII5lOCe+4271Lb5fKbBmIo8p+z+xDSyd22wfzdWJZU40x6SysuNMb+CjX6FJk/a4w0ED6J
Oi1BGMZrEuMFmZ/T2JWKxHpOxe5K06hDQcZ414QgBKyNmFducJHvFjsRMz4PahFw5dqzKJDBlSrK
Jbt0hkMb2G+ByJChwgHs0o3d3EAwbMI6kYzJT8KNibsBwy0VT5tcye4o02Lw78v1owTiprIEF+ve
GuovR9hwUBzDGeD2R08NbDowSQ0pBIRl9/K+Y6buxTJPQ1Os4FbnfpmEZ3r9AONYallX0SGJLtFo
BnYRcl+Tw9K3Ywfo5r2zHQvYxJZRYiwGdTYcjFNPrV+GXSADFNmrad2dSQxMPAwXZ16P3oRrc0T7
msPRr3GyrO5rzyzC9V6gXdHU+zuzIuaenpe6E01CJYWJxFOiDD9ccXwB9bCRbAs7VpC7mqMqEtCQ
z7I9nBRfTyRFT0rXq//l2uEeVlcoaYwJ61/6rqv5ToLLXEuyqT1lO1yt3SL0OaXtnxqaJY2VtjTv
Joibu+R33GAyf9S+/eTcTSvAXYXC5GbCdrbf1bVyszITilZkZFEdD5jt+j+4x75jSrTXJ7iqpbNT
cyYCKIDpqimDxeLnuULWPPnEYyIm5dXkkQAV2f2N7kNwhDwVW8Ra41TqssW18q/Ib/K1IOerTW7E
eSozE2QdK8FqcgRbcoHCg1si9BeHJpPYUjkkJ+cDGFcQsYmaAaBrMbKsTbjS3gHeyIyBqOts4yOh
phCyH2JyiWMrnnm4sJKdaRow3ePU9dTL26n+iOIY+0R6TrVk6nilLOzdaah32lse42sX5mg2aQF4
RxkJOvzW5JXIk1MKQ23+ErJsjSt2wARieAw/79bbg/5CBvc+mvmdmtnHO2Buao0NDSAKHnimrSss
jQKgxNwvBXTiGsYJ1SA9ujhFXnOZgcAXFLjba8omlZsQexjgiVXecvx85lkokUJvrvpwiyCsISlg
CnyqnMLEXC1yEgI5gSxyPvZA6tMwJ3M+lkxItd6PiZyp8BouCHpF05OWHyCKvz0wV/9goRIMYmbc
op/a7ST22yCLq+FLW7gDGCgTGasHXTzWzA/VnzYJKFQ1Pz0MCvlnr0GZBRPRxLsY43hOvKXZG4fM
7sDc/v9R/tks2SWVoF1j2Y+xacZgQURXRZNeqfUFCpUA1xFhbyMX+vmTaamYt/ZyBrxmh8/fa782
2JReytx49w/7sQd0DncYgEuaP95YZDLRP3fjPljY52yW5Dqs73GROYoHK/C82vyjkeji4dFlKmdy
xz9AKBYx609MN+v5ZvxSksT2AYY6jo2FM8svIskE/DlUBpFAsMYAzWaRixtuGxwRq0nf3Yi/8dAi
/iA3SjIDgdtyKhC4vWZIgnMS9l8L+eRVQk1doEsZoZnmudaouwq/iJAwIyZxXK7IXyyUrh95q9NE
iAXrMONLCTmlh3cOTozUWAaV3+cbhDX0avlJ1GkU4eRBwZMrDrpJFJD2sLwQMKuuYu8DnBSQiwxg
6fWLUhraOpM/2TlBcylVoMC0boFhX3golbRFnT9v12GSiUHEvcsVjEKMoY+c0phuj3juyqENl4t7
1lVeMrRzYUskU+41YkVEBPC7Ydu+/iR+ERNwhfYQSo+dhTpsEqHnPiMXvwMBmtnwPAU5JxrdDRPt
FCWNMn9PXx8fYd0YAUqCAT4KcqaOksLgdp8t1hgnvh5N3ohlh2lEi8mdR/Fz5M7ySCLH5Y/rqr0h
HLRR41axOfj1XJYlZlnlAqMeVLZAi6mvRHuv2xdK1ULW5pRDudpQXC2bBvo87gxeZFAi3cDQRoG8
JNTshgncY5uqzpY8InqFVeSLNqE3lNM70ChSQfn/B2RMrisKn1PQ9U3qkeaHHP4raGkUGXJGBlKi
yll+GH6ga3Cm0INns863hmyitRQEGHBR3UmThRH4HP4vio2vBFPs/k5h5/DUc5eYOqCor2dIOklb
Iug9D2CXzavjfkNkwz7F9CVJOVU4wFuNu9ni8tQIdN5F6ZO5sdzpDdLLNhhauM6L26N/nxhHpnzC
50CrP8rVvqz676+YPlxzcZ7M42RW3hH/Lv6g5bLueLFmvnG2pKuhCS7/rGma8B2TeRgXWEz0CbIZ
9Mdz0CMR3+Wbr7Y6h970xA2bkWnFF4ku/vXHvtKewrqRSYzeMHtfiMzzJEpZyx5yglJb70RxHtRB
kM9YqwMt0aZ7hxZT7/2OGHA9mH+c4eKUzfYjJbmdy/Qiy3QggBknIk2zFgCKObVflU+isHN+PjYr
7xG4zwsUa8BgVAnKZDbyCMeXis3JhEkA5Gu/ILXjGqovd+Hih+LSkNFTswNxl1BDfRJybggpWb0y
hAJYOjgECxCyQM7hkWz/XcOjttkR1EwmSYhTXd+dpoUGEDgiHM8kGObUtCFsdx13RYPZlzex0vox
MS1jSndD51KPYUevTaBeKerWr4DYPZOXcyZz0t5KTZO94tB8Hq1Qu8HT20+jxY9OIt0QxGIyc20V
V/CGf76qQASKswQI1XHDESpzMUiY0xoagyjjyAT1yjntI2h8GGlf6CNF7Dl3ICW5eW+jINGQ8ysf
JOP90OAbbMt/AE3kRDtj0mDriYF5xGjmYNlyy77u5q0rPktjzp8sbEX1u9uCVvU1WTpTeIakQiuH
M/9g9mn+6ZAUdrjQITKApRr62Hqr2csGeWf+Fz6ifML0LEM3xLp+rBsW/UEKCjC8iYti3AWImBs4
qFwNcxsH9HtqY3nUhdFZ06aL2GGCGconIJELpSORGfCFnXYjZ7vfWC26bxrbOTS08FbipbJ0OiLI
paR/KmmWr8L7PPAB1HOIzk3cQ+MrforJMWBudJIM17vVwqZBNbPZO+PG75jPImJAvkVo82aos+Vb
M7F0T2YLBmqqy71TTS4HTO1pkhu/GvF4yE7jLInWcOwiJ0NOZAYf8Vf4VjNFRzbx+rdX99cBfzYf
K8TzjL6Qaf7DBS8hlLDLfdAp8ijWjDqkh68N4gY5MYdU1TMJoatud8oQxM1FEIARFql6Vj3IG0AI
mT02vxDJYO8R402WVpWlZ2CQsdeQQvt+PAWS/GYkDr14GRwxr1ovuFf1xI/XBQXFuwWT2K4hctG5
TVNIJ5RhVP213VGqV8tWMNTdpTfnn5/AHoON4RYILJCi6qI3UtphxZWNlHJ3/Jr7Dr2XlKySogb/
AcPfRnX6Vsm1o1YwOI955B+LXUyPPCxw7vEnpjN2xTrz6HD7TQk9kAfFGSDOwcfU8m/UDMzbIgD8
BJQqbwE98eKCJi6kHCwFswb33OYE+r+Tr0ZE4TRmaUuwfLtR7fcBw6HT2rXEdfV3bJeIFpsGeckO
YOinZR/fBddJJ2FuULWX/0Tbl/YmLk9qbX9PPEr4NSfE9Y4VJs5WLoypkTfZAwUwM6hNTvEupWkd
46f8IuREr6fTgQ2IbV5RO0QNIkPKiKkxqmIIltblf9ALxt85MifD3u3yhR/RRfokZIVV1K4yPIAj
4Feb/2LysD0nBAT2Nle2r+NH03Tk/3gFbCtWUGxwl59Zp2nNATBNpJvU5EmGA8rp5SUWHSk7lIpE
ut8UK40Rh+ctMNW1s26LeaUTnfujtKbxfjSTcql5CrrPUZ7ZuN2LWR5vSobzWMd9lEejGJNVv9ZO
3l2gKkelUg5EgmuFYfFUVDb7tOeCKr70iuRCev8tU4Hfvj6wr0kaSAskgJoRf+GRksL2Wkwf/029
t1W4OB6Ai4Tf5nNEntRhVhb3kKNCqGzDunKXp+5z2pJ2HybJDDOnefBk+ZN9iLqvk1OQJ0c+wd9z
RXYTRNos3Lth6sDxetkRcv4jpe4Gzu8qdWy4Px8DbhgOBB/7WfMXN+mdKcfpLxmTlWM8r6QMWr2X
KGVoFRZeSJWevxIHFaT4f37XF+hDYN5fWP0u8fAl7td8Ap2MnlWZxnNtv1M3xO/hDSh3IlMOi1mG
MIThbYKjCRJiyqLHC/jOSvS0FjcTYuKWNulzfrF8Ob4btKkwv192EAFrZUuigqORwSV/G+TxLdTv
XU6q3p39Wfc0TINH+qUxFLTS10+0iyXlo0i92ZjMcecUAZda/jTyjoZFMVVjPZ6pjTeN3yjwi4To
kmMqi/lmwjvnTKPKKf9FHdGOleK0ThoZZXLCRXUTGjQ36v+uw95uUHFmA7jtpbxpHNVz/wzFm1j8
P+9RU0aGMsTV2qFRvSHPS7w54rWLkjGHaRaeG5XNB7gZLzU/tT1yFg1zjm3P6aS6ObhWREarZ0tR
2G1AiXqLBWnz4/rzdmfcsW/i61s3iCCLme+8W4a6nv1YVDtI9pebpJ4qPgY8eirsuW3ra4GmNMhy
LbfDfEpU++/SiWD6JKikDccmZjRCfS0wyY2u2AUolOajy9y7Pm9irtYEBDh3GSrnzNCAhv3KJO1b
vXXulPWzQAd0L6H6zL1uverloba0Chby2yETu/fDhgkwJPS7lKUdAhvy+nJ7Mcq8zq8eX+/kJkzw
szTsXjFfVYNYYIovbAMS5GOKnSO5++yerSesJA/O+CzmDb6bCC31qGLTzSQ2TrkDkFr+BOC+a4X+
qqeSqQJy8DcGULh/ROe0+t1bgR0rGf6eFR+AH8PclM4PNA3M2hL1wDAyTgdMIvyzSA3i3LcgOYH+
ztEVcl2o2Pv8eUlmESZiVpzV6EUQPAOcCKbPQI+WFhFGsSzgVLyiu4WdxbH+BY/gaELWpsMyUFS+
bekmes5x+UlLmcn8TkrzfY96zgrqgPelGs2wnJfNda+IBlVFfuzH0R6ZBYkLf//btVQj0ac8Ltbx
92ZYAIEWMNQU6EbfXkP79u88QE/Q1wEYuDwIfEQrfa2/mHUkhFdSFcbtP4+m2hocf83OcFhQBISG
9OB4HwtTuqTSjzLqCw6ywRzaJ2pjxy0ntVb8GKvS+wlVXtr5BUQSWrDMtkrrSYovu43dSEo6DcA9
KoJaQSekp8EI8T6bhsHwfaX3zVOzl9IeJ3v17ptu5r4nLxLesmJFEaHBhCPK9cwvgq7ExF1E9/tU
8GW2/blo4/N7j8tCIEzs6/nmjLUfqOTkwiiYfphVJFit3A4oK2/ZU61xw1ZALiAlLEwtCrRi2yBi
f/KV9vLU+NCIAAMgBxyd6onuG3Xvtl/Q7IWz9FqJkToNeSzbe70hOOaKjo3a7aGsSkZfsL4B9gr5
aSQWVsoDOn0ptEfuMDaX9LcD+6axbkaPWFai+kBcuA0hv7sxY1SkISM7JlWPfS1wUUUQIJVKH5Df
EXUtwPimRCEfN1wHLvQHXjsZQHZlywTkjEc1qGd/xwRWugJbwkNJXIWfKBl4sNLWUpolYrFXOny2
nS3hfVgMZaXt2JmOsGQKxguDMEsSADCNCPyakEH4kcgGm8EyoVYw1bW3rwwX2F2xiZMZl+oyOY84
eE/IkHtU07pYmJO9UF5Qq1csYqXiSvCSGdbyDXNxtyDWhqmA2pG/NKA1ZaazdISbMmK1rAxAVNZK
hKtusjALEmghYXonFWotHHRe+IWEsfgORlwvr/5j9urX0s5tJo2DCRmKddkJ4DGFXOiSI2hgDIox
bnaSeYyop7ZTAE5jHitPjxXIH/rvzACS5Ilue3sxG7tBLjt0a6LMdQeWbPcgY5wKqipHLjvwGZyJ
CAESJHhNb55uszRD5I60TCVDvDIpjaiiW6yyev02G2D1ffJMIMj9LZyGGuZLLDz6RahvX8VqQsWk
0pEnBieaQ5OB6ykL+Sb+gh+qtzs3iOqhcrrr3bDvsny9AgNRGQcq2/yp07h/ilTl/S1tToMKJvwI
oZaHesGTobV7JIXFHAmmU9n+KbiChUZq95fWeEzz4wvO4VYqeGS+IjxOZAZo1Ue6C4C+jrBg8FV1
RFDTpkdQJJD8YowthRVbKDWxu+1AjwhZlZ2uxi/40cO/iwptf6SsCJ7t3pCBk/qKV2WN7dcpx9N2
1seSV7FRJScDe9hx9QMjaqekRryRRUaUENabL8n18ZV+f51bCCYSVcR8aphZF5SMSJmCisf/9+oe
Y+YOG36imIicOSOXXCd+O85+dHNSJBAmGLXOZ5qzv1JcMT38HEX5l8P+3MYxA2SwXc3BS84GqQb9
kB1Ks0mVXI972cCVVMZ4d+hTBu1SnZBm1IrywAnk8ikkiWe3lKtI7jmvigw7gNOnvWH2a528pgG1
QH7lNWk1litmtB1xi6nnh4ZZSSI0/k9gsRD7J5ePrmJjXFh/mNx+lycJXA0wkzU5EUwctnKFYJ3v
FgMv8K7uzz6ZZYM7jyP3W3gcaLh/2TwGjx9flLiLEdOnmg18h3NWLpJwQkMTH2WS2PsNgEqWf+7n
5isYX4rdx6BGeEb460/ROVwmoBoX5iz70tiE+LZEjjXQ/xW9g1LnQfIzNLsAWiLrnptR93LE5UoD
EjX8FlOcuPs+0/icAFZ0ZgpnNkbzHz8jU2XoGiWzC6g3tQDRJzPMnnnkeRekUsk7G22O0bbuKnOK
7BHVRm1p2n0SYHGDYTjQIBK79TnpFFuPjkPt3o8pWm6n57kyJUrDOHlbrk1fi+/kVI+/t2hgmV1d
4UcgDPuQbjVEZu/9ub+cadPh4vVgeqfmsj+Wj68DNg0Qm3HX4I8frW6y8JB5Q3mFgKIG3Abctf8e
wdzRXWfRONwju/SaIB5V1PgoF602fg0n+s6+I8dBjt21FyipvVspblmexQKfflv+SHMPZD+EEyX1
5GCCTknSbsi7xz+SkWnDeLN01HwDJEvHJYD4P437rP5HzoS+T/vF9bVX2M2BudQTX2LslYrxngj9
0ZLed3ap3XP+UC9rrXZVUeJ3EWOxy1sJfmwkZ89UWzZodXLBqQMfCWa7VsM0TdHDKjOkbQOnRQYJ
M3QSGYeqgkFh1zCj6mdnrfuduzIq2UW3HNt1t0wgNwEwzk65sS9LqI3wxKtHnoymyt/XuFJg8P40
04WpceGiszaqJ9iQy9aTh/juapYxEmU88JahMySKjp0oBKs7QtoGCYlEZL2u1NWdFkHeukYqh5hC
q7rAVPjXSeGiYQDGqHP+aQBHpELx15mtEjEDJSlKmOufOZAzu8Tde4BpdKAmsg6VagC0e913IhuO
QxYPeZuugPiGdaSHJHar31sqpUj83RArKPx9kXx2j5O7BKjYWBeHzzCR06q8gwPWeNdFiKOMhKbd
XjUqWXAHzjpqInvkTI2DAUI/9iluneiIKGHFQB0m1t3YDt0GC6ltJxeIqSjCQJ7gYzGVHhX6FxZ+
1Lqjd8F9JrcYbPtubV7gEIJj/o1IV2VhG2DAfiTwdhmjPWLDTR9ktR5v5oQyZp77hexWMeLZeuOr
F008wU+ZEj9I9Yckf3618j8vRMOXek7UbHSSI8ybuN23vCSOu03x3eK1kg5HvbUju2o4VVu4uyps
dNHn4tulmLzr2aN1dqHKggDjWkd6UXU4YZw8yI2vtSZ3Jbm/8MCj8KgUtS7OD9nZ9Yj6mH/a/Bks
mTjb7Oy0HH2XwJvq1cyebnABULPPAz9tvIX+k5C0GstZwy9kTC91+Mry1TIsx0AK5VMJz/S9ihWi
h2WSA2ChFk9PRg18NX1NwCFECr9a9T0JDe63locyB++Hf8v0eGZvA6wjyZQHXeW4lDVGEwzKunEN
doo9gEuGDeCRb3Q9USu0n/8HuM+G5jO9uknviaa9j181q2S+wLf+DkYTEbGpJNAl3j22G1wti01p
wMJKhjAtvLehyzZmkMawHM36sFFhfoWjm8Kd3vYTJKVjdKfbwhw3GJrinvv+NBD3OIV2OIdZtSkG
L3RYgtD469KObTFXKZHfjBq1zM8SoZ4OJj6FkRn5bPWja1FZZHJDY3Nkk7frniBrTLEl80ZROnzf
gpVPGdBOcdQ+6MrZufDz6q4Ww4277f09D4GnjLQ7AgdlDx1/FDi5CNIwDV/BAY5ziBn2TgPZ/9bo
1dTfk5AuncA6QB3oNu35yj6ZrlnLSLCrTsxuuGMRD/rDFrGmI6i2gNyVJVnLIgUEaWaaKwLHSaZX
TcxSDQW7OK/TXtyogPpperRlSxqeo0c5db8OnyEsedE8rGhfREmm0LASAFX7b29/+5/CqocUmdwN
1RqEM4MvbOnT9g3ov0J8dotFpqEwpD8hTB0ispbd7hJIwD0jFDRUJkXUtk2j76u9OjoAtTd38kK6
950a91RR0O0n53vpoSc6fn78BGdpoSgwCqLDfh0SDl7qbHG0fLbtCZhfOckH0FaqkkcoiN472Isg
IXa6tAffcZtucLoKFKDWBO3+XDKaoAF4N97rUGeb+DRVDi7+gEd+F5KluvHlEo7pND/99oeqiE1r
7lLRZSPuMOWDGb+PYuZdFn9vH9iovHkyEIsYLIf9o9K0rJScee7M2vPq17yi77ZWItxAw+fWxuE3
hQ9rrMIu64KiGZ48Xc2jAklNhxihf8n4xUTNLWws1Y34bg2x6q54uTlxE1psCsOK7JaFWhcgAOWX
WcnHJ/MDDtc2mXaUJL537ETVMWnLgW0sCQJ2VZUi2FT3XgI7bhHPhAPN3kFAs7HBBzOXgzKG4O5/
3MQuyJnBv2S6+dIDjzJogGRQI0ZSI809XWzrirxC3Brv1tUb4yIaHIJ0us3IPWU0Lb/t1+T7wVHU
nQEV1RsJ4q6Ueh+1xxqs1fFpir6QAw/lPCrJ4yjSDAJb68PPeWNsAbeqe/jzY2EmToWlN0Uv/AaP
PBg8PomtoZmMA9m+VMfqraoxqZPo5bUJ2hCQs6uCMK+QkI/caBvoA8ISIW7Y+PyCIyJWa867yyjZ
xznVntPJRpkC2jPPp9xouabpmcjnTb4e23ewDZJY9Iw568nH2iehqRwq2q5NDfmK3FZfeb9JlU/o
zWEBDQVqcnibgUlITnJlCI232WKS6+0AUTwyzMndU+b99hUB6R6qqNDgjfKYZE9XBwV79Q0RXGxR
n6codsLb819G/xlQGeLu737U+GBx1yn9bUzxdVShLuM/SzZogY8yVYGGSAVbdukQ/PYqN+rn8bAU
acGsj+KOWYwl61CGj4/1Y4Qc4REDm9/kmJBYDv8nmhFVffzg7kihCQSNCD3Lf8/LBNY3ix3mbCVx
HcHL7CK6GhnQldFveHImgM8KWBTUVj2+NPzNIo1QmWFLBjRSAoVoCZZgGAWoLispn2+p5dEW1Jy2
AuZ6dzqd8k1RC2x8hqp+/fFb4MZCQJH9FuA48ERB9vUXkQ8BId1Fl6zFsXqvTzv4cSvJ4oFvUo5W
iYJ2HgTXU7xu6i5fsZ13Ljmi04+Efg0BwVtIzOSjoRTTQYdXAg2e8Yh+kDT81y2vOK4plSnCImwp
fsrYIQ91yTmW2ROLWm4SAwOy8m5TzBAvlT2JUvNnPD66GcZllohzkk5dNSq4Q7hIZ+gxGemhKfkN
ddLBnt7KBvuUQ40/dMtHtbZ8IEZcj2esNt63PygrTV8E+lq3960/YfRYlTP+Ebc1CUYZL48m5LPU
HHg8S8tPTkD9lIEY06TUsOKP3Adb4Y4oYBIdsVmOpHUWdLyQQYp5YJcK018RtIKHZ5HVm9d6k/+I
krHWzFjShl8+eSn0OZCmYRMPMgRhaTURvNJKtpU+jEq8dDSC6m39vFG9t+h+MnriXKY0vDaOhc6w
FTMMUcHy9nlU1HO2ntyztdAu7NTLQ1pCDeTUQiQTBRIEZAgA5pZth/PXhRRnuJQi1om6vXev/pS5
MKWbowyArhYitxAQ/Toep7fstSuk1+Rj6MaQT3Soj4hl1ihMQ8jtBzqBzGUbhULDGnPlLaQqlWnt
i7J8Fm6cR0kxCSH7n/s9dg9Cy72Xvis5KI1VEJrB1hHjvmmD30G22iJOcik0z8HHnW+XMIIirdVq
IstiUSh3EW+fTAwwbb9CKSvTDZuCwJF8ecoLjXGQPwChDdMfqn9ctmgC6Q2UOXWyGvGoAJQiNndu
gKvlkUGGN3s7KOidHCJPPm+iZWI3vb0RPKWh+8ZlpEAKWP6TkeOEwtKBuli1vQXjcKxR5r97cowd
mqCqSbVTolW9XfFRaiU+r6pU0tF7iTxa8kyVh6Fw/5Kj+DQTHe/7+RlTTitbGoXGeKxLgeKHuOdE
JT6WKzpyXP5QpHiB+uUIXtPTlSMPKETKIgw4CGl3mPf946jpPUhuN+TmLRh/HDjvZf3eyk6MxqKy
aCx4MIjGbBEJOPISsw0+oK7tVzNs2c1LlPqlOSSt2zMqddvNhU+roLx7QCXugl5U+w60n5BcR7ty
mMZhIBp8IR4hPf8j6QnIt2toy8cxD46sfc/y/5FjD9kgPGU4hU0bMEnJ4w2v73PMa0IST7CMt94w
5n1APa0GD6Jp5ukKy4PTzo3uwjNrBsWBQH8QVWnuo6Gq/d6xHIUEFs98Y1ntkbhA7WcF4BF6YxNa
bW3w6MrYGrPr/VSK7/Im6yYXLLc0ODcHUe/WIpuHBiXImKWaC7ugi1qvaHkiNxPITiQbXA0dbJWu
+Phyf2OvBxQ0Csp30OalvOtpDmbj1xKZGR05TEd4zQ6Uit8RinCXAcNUIeIt5r+v39WNKmVrBUIF
1G3Q2aentPoQpOn7Fz068x2uhJeQpav2SG8N727mvL5Wqt6msKwswPrjgG602cPiFE7n4ac622SK
U62QmPp4lQGzntZvPpJfkVGkr2OfhpbR+/KSBMeBNaZ6HXuPttO87oBFj5YUeKNtCR892YaH+fng
wnPZIiey+DIjLvFrL57jOUl/jnTcf65TvrpR4C7RzBFkJMUMB3hQPG6gmCK1aRT66UX2RmXh9b3b
02OZur0R/8xTBlHu9HdRDB+kkEqwdXe7YGqnJyk4s8sffP+GhNhz3HSUrUYW5Plee32o6cHJlge7
cIqTS9QwmVbB8S1JNrFnk41qmEGBfp53b9LtjzbxEZ6J8npnKCdfMvSRP/cgVIORq7j81x1ksFyD
nrOs3Wnzxr1NRm3Eln9nvCRt52MW1wcpLBm73M5g8vKQc8kqCQn3YjlGbixIuA5F4ZwTCFwcINSh
mZFBaCOnwlgl8y86gJ8wXVIFIFTpJENSh2A/TIUAuUvOUHBYhE2U2/j8o0OBwUYp8tJ5++g4CPVV
YEKBwUYbiIZ0uu5/k1fPSSS5mLx5n3blIHons0fyVE1TDdu8RMaOh0+0N3FnKIRigmwDNvCmt2JU
hH1oq3C/6zyeL83EmFyBQohKYB6fvqjAW1O7STL6XA86SwGvky/Dy17Vu1hh7THQKhuW6HngMuMA
5jW39z0npEF3RqjjcQZ7WSnZM3+YvQpdHnPfomP1IB6DnrUl9BFiGCph+OaNfjQkpakyUmSQPe5h
L06yvK2qEigAD7aZsIrYGiivh0TgcrTpvL0uc7nxj1sScd/FLK3AldwEldF7OIYAhZGFYT8Tcawa
BsVaUZj1nm7weeCBf9hFTADKDk4BDoSebz9So7QyfQ97+67djIHA1+ciEEopkpdK3H2JPKeIbJQF
ijOPFjKuhk/41vLMJmleSgC3fdEzQFW3TueFI2UxFB3keRRnWZChiidorgU6tVgZ5S1vzieN++Yj
VF7wkdJghezbtWfz52HDOLal0lDXUfUC46448ohyES0sxuDd+4kROdQHbL8Y+NwtoN2HsaxwRk35
SjaRemTfLCRQc/Y1n8aFeVRKQgjU/J7Bt7zbbQ05GCykn8F/S91iWny0SDrV9vxWI30pLX/JnNAK
OA7v2/LlDLo4PWKbq6FEy3rW3kuFaMgnZhWrHyAuAFNhdw4vGQjbmRotBX+l0uNOR+2W3nrwc4pv
mhuhFGAT2sZ9GZ5TYKuah9BnM3LcJhz/gT1xr4s0uQfMhHwwt034uBSzleyV56y+rHqnghyE7Whn
veQTGeMy98uTu/UgcYgYUbqrHxy05Kd+6iRUjtXuGdYSfC0ujsxQtuZDG3OCLQQ3BYANusJ8L1R6
mfNVNrLrvmnj8YU+0htTaOb6Fb7hD6A5Tt0Nf+zQJRcCCERzAePSutjs18OFh9HKCcBsHbkp7pP4
L3wCz50Edof+lzT9jNEkDQcnzZpc5YZar1ZhXR7J1hNrf9isI9hb6yB+uBGXJ6yKWeYQI0xlInoK
NEDdf+mJPz8ZIemqYVpjonr8o3IjXSGclLGUpGof93nw8F5kSmRQyZFkHepB2nNvHV5iDVae/8/k
G39F/Q1NG+N1bj67zk2haUbK5kKppb01V9KX6N9oBVemdVtG6ldIG8aNFJTm4MV8Q/Lo1n+6p2mc
UTp1PNQnaBnKkrbPWki40QCv9mHgSPy7SNG/Yj/pU8JKPEApYwPsiTgk3HvBWuTuVsT48cdN2688
DGnjLapOGkpma8S6vkZ+KDgS44s+gMaJlozgiK00CHhcnSXFPxlnUuBCB1CiqwNGrW7z1v1dI+w7
aiUHhxH8Olu+1f4lFtJDTPUzn2p+RHwsMKxcXEsGScOJdsSIIaFL40q2+49QMfDmee14vlzgnVar
pg2zZ/OzuQhLNhooTQIzqA+7u/ZLUOOBk4jk+3hDpspAJu9QPBrK2U94IDO0iupiEchG2mL8rnza
gz5VPK6c7y3NkDTu1q3sBwD3GMHSdHoZRVWZXhrs3JQJHiMIkUex5QCS2RU5b6H66zuAPx9ZNCWY
2DUjtrhRjNNIeWmqYOyKGwpXQw2kfIy5FXH7ywcvI82xr1B4qqHQzFsR1iuAufyCjVz7Fy8Lo8EB
6Zb8RoH/ajkR3de3e61pW3K84T121LcKA3f0v0nEkY4Nm1vdaAXO2x+46EjOetYP7jnTjHS/2XS+
7eT2eO7dgNb1Wui8fUc/igiL7/Vk4jHL8FTG+u+JIn5Nc3q9pKZ1/X9QzTCp8074X5H1ZrY2yMwe
YKk8JNEqZ4jkeqP7KZXvovLFYHsS6PQrNt1iwcFux/t/bnouNbC11WFB41qI7lXh1aaK0FBcC73E
WQseTZPW9ske7nXKPuuQZ+zTqxmEeIq/XCXE53hnaEGelJ9Gm6O+yUqAORaKmTIbv2bOiIZiW4Kf
fnTXGWv2rwHaWFre8+DKkDhpsQHw8tXS68890E4ReAcsXU5H85oJUzq6+Ag/Al+NX2fTIwNsv2XL
E394VbCEB6Q3pD9SmVFjy9MYqVj+Q7lYuBoNurKxqdXQaYefpqdeD9s49TyH7wVkJDTz3abBrQDa
lpTPc13av/T9g57R5GE5Fsrp3uyEtYy0CWk2Ae3x0R9kuyGvi3sppebL2N4nGZCm1jGJ4V093DP+
EpTa/XzlxwY5trnP8zyAJMe3Tk7kZHzBGCwpKTP21ltbVmalFVzPKHtsSJDZYgjVuzC+y7J/N2q1
Wacc5kpIZaA3ea+wK1WTFQmAMKvIHhi5yXucSB8pu47sScgWLbMauIo73maMtL1JyGczx5fa90r0
UHno3oD5F/On90XQRWJIgSGjZ4pE5ed5WU9iJHYMWBYuAxNU6rfb6QfuGL+2nsBkGMEFWK7iWaLS
SZocEXT10JWdFuFIBq28+NKti4SEtxPaGoPvd+aCxKXdrpdwUAjzUVEiubptooiPLOxFvQmoSDAA
C8PGaW58Hflc+RINRZV8bQ8MhSRqwcBP/9DIybcTFpm6VzYmAfOPaT0UAr+hcBIBgJng/nO8F3jk
KzE5CRKn6Oo8gzMCfEVVK2362OWJrjBOmSQAEoT38oPNpwpKb7J39qM7NqGVtUcKhXRGxXb2EgFO
kQLivUGckwu5QBTv2mDfkINCX21nG+gUJOA5r4cFKrxuTPExpNRD//tZ8rkU543yihhJ/FYwyprx
9ViDQBd4/4P4+Kz9Bsu0Cv9w0+naLgVz3f43lSgH0UcFXVgx/bcaQMo0fJF8UEQkNJyOk8UeEVQL
Z4u+9JcgMOKVAvC1UMWuPWIRQQi+QNBdktF6uGd9lFMm8+/BFp4JUKtDxjqHct/Vis8Smgsj9Z/W
eCVTIXIa4tH2wTEFjBgEOXpuTVUf+qSUhV/OEu9mDVkVbklvsH06OzXTKq9a7qfMvXE6NItQS9MV
67G8Zl6A08hW+moriOYFf998L64H9g2c/Xe6vwNdRqnaqgNHWYCK2uevUbiAKJ5bfYAT8EMgFo13
4b4favcG8NNDBvMtDm0zOre9wyc91al2FiWdGrN0lcl/qof9OkRGUV49Z8MJ9QXqZUu4WtJGbI+a
8JcEZECIoazpyPCYL4xLMM8vH1y4tmW2qbQTl0GiZC8KIyaMR4e4Tm83FiJe9r+9RVU/0Kx/u5/u
8o3hTXPI0SyBSvp1thH0nHKa7t+ZDqb/LGE1FyZsCzkYzvNu+uSPFZJhncpknwl3GgRLuzw+lj+v
me3QjNifsgMXJiJNY2EtlkwWXS9mrls8RH6YUY0Wc8uaT7w2y5KVtJLNysfRcqd508kNv3cvuXU0
EQCAsGtXOd+iVpdgiZ0eedBQbMgUEBvuBfsAPS0Rtb5hNtoJZMrDPDxQFyg+KuukwO5ZFMdTRXQV
kLlJPPhmEJP8ti/ST0KfmtDt6vfpNMAvMI7QKrt/poVxEAwTWl+Fk4K+HLfzK3adhgyn24Cnrukl
GalcqAkXxlr7Xp+NKxJbHQTxKP5Zu933wduJBEixllHvFhQBReBdvG6CLx+QC6aRD6BNWMQwtyrc
XDFgkF+B0WyxF9oiO4o4fiM9gIq0pxBHg7DRsDutTcHQBgl62uHfQNtyYYgkLl/rQleHiUG4aNLv
J/5zLGlfNoIwxK7oinniMFocxRbYyqG1hST6TqxUB8j2mUi+PDK/m9RdU5z86pmDIDARmuy4wbyN
2V+oswA3hBIX4l0zlwW29MbBduuGaTiEogxD3KUcHUttvR0/KeOy700usoDkfxZbGk8bnEnDrObk
V7Cw0yxUXrhS4Ppb+SGh/KvE9eFAb+WJ1Uu9KV92hT+1vUaWh91lrmIPgJUi7CFE14Mv7qdeLRLj
b4DVQJVKsZ3NINiVjZZssM6DmFLOpHQ+CxigU4khcszHiluvzHT9E1hahqlxQMU7rkfVF626/q6U
frwPoFHCu5yNcfS2Y12WUn5XMDfEPOVEn2UxAUfgtObNoLfhm2bGIZs+p2bjpKtxbe3d+QbdSmON
swRGGchT+RZJVW0v4aA8t/aliws3PHUtbjA5GXnuohFMf/S0uYfw2PMTl372CxZQpWfJ6eXXDvst
IMFsnzTpCakUOU6iAvQRB5qP0OGXckjDfWQZNCDoP1JvlOwen3Os0CoSDejBA11Qa1uhQJOrRndm
vnv7hCLetP6PFTJhPL7NlF/Gt9/LnmJR5fNzoSENxvGGhUngZA4xuCeXWXj2k10hEjZLH6Fi7C3n
ahgZkWIASG75ofUdXON2OjIDYPV+ql0C9IHtJ1ACH6Ak/2wUTdzURtYhR80640+C35TXKhCaybn4
pfNxNDO6lWSI4wTYbH5ojSdclF/Nf8oaj3G0qtTeiASzYppjjXdW2x0anF/pPRFIc/tkGx/2xE7J
twmd0Pcq2mTCtbQuvgq06yTCJ0KCwy1pL3oHVYrq5DyFQHxBTKh7aw/OxiBYH8ESQaEWo/pwDPG3
AXtgEkskOYo2DraIzRd+PUeEvI6Hxh3ur3hsij0YEz+MylI932WImSvXD7mjTZFSM58Qpz344HyB
liinqYfKoZefaaAJplUUqjq/b1NSFkltNsQqB9V52o3rJwOlkjfblwUzYjlpopXcVmd+c8PDqyY0
nY0KF2luxX9f0ZJH+RPqlBKw7ZKT3YlJjBa5JWsWuNCqicuU6p3I95I0ddC7crIaxtldY1iMBqI3
qLAn4Za5NJQ+q2rxSI6iwewrgo7TR0of5nClQPDDQOD5IHzNWYsEZwGsJ14OCQwgDqWPADpcobPV
n+K8oSGatXeo/vRjljGKbmUm7JcnGx4wkh3npb4HH9pw3aztEyD3SYr4i4EC04MaKJWmbumeKqQs
C0YO/Ak7gJAAkMtMl7LNW1R8gW62vv/0v36eO2whXcWZik3SaiPCFOIISPB7JfeidGO6Y+9f3TZQ
N2ijs61Kej56tJ6l3khw3C1zGmxBYwkkapQH12a6Hdae+a9m13d7fUPYSTi10htUkc8DCtKS2n2N
94g18gOJdRGG8EPsy3doYbnyCUexKDiZT6pKHLFiBQlOYR9nhxHLWRsb3ODAfYMB/g9Ms/95HTBK
v8++/BZ1SZGyYzC5cz3LuaIGsJF7koDEig+1IuHBhHUmTw7NZvkSAXrRTNBLxmFLCukCCaCmzjkQ
le1bQ8okW2vWrO3y3DeoJXRl0MV87QROM21WOdQ9tL5vlF8yNS9IRDHVfQEWITQdXMnffbqyixYQ
54TXBLvhxzO6mtKxdhHarWM2Hqsax1WWWLDaGywDWFhcxBGL4Jg6AvbLg1LQhryH8yr8D65lN2Cv
Lw8YWA0jJZks4HG55J1kXn0qydYj7Vy2W3W2zTlaN7F3hzSNLSyUUOCfX7jB5DAnn6ZMJnsj8J3a
vs9IVp0AIluVlboWU8ziODFUdwKC5W1IGlqjs895JQeTZG6RP/b/ApJxnA5ee6wEHkJFEXqEza5S
DUv3nUTbQmPawtfIuqPOulIb/lKwOsKQ/fkKNe874Xo/XH9SAxxKJp9n/GCoHd8X1GUegOCf95aI
zm33cG1Dn9UIGYQ9huJrsolqie3ANhaYEbIWylnEt2z5SG8kbE+Irr6pYb3iR9hA56lYvn/erOjC
d6TRkZI9g9jGSOnXjmyzWLjsn8pPZvRkUGhgZxAn1Gt8YSNmKWs8m7pckJ/Qu/YFQrlNyGHJZzuW
NrzvCxvVTiW0x3i5kYwiA8cekZQhPpf5z4roYN9YVCZvG4+kw2MnA5wXQGl4mFbOWI9bEugasxHV
qBkInMR4IZFgnHegqZS3eE7rjwnnxOnZNQAAeJRp7sdB2n6dnO+suhEwd1qt+sPSJBVNoLoodUbM
vd/jJccMS/x+LUuPYvboSQbqe1cQIZ1kl8bo7e8APTgJvkXXfDYppfTI6ZoVAfSMo46ajEKkd5G8
ChplT2C7RiomcCANFj7q+LfG72eeNejMU1rTc9TtTySrjIjNznY5fr9ARbIBi6sKoxAXEfXjcdE6
Xo2k+DpyAxl5OGIIDeJIbBdR9FV9WSguj0Rf95TFvpcX6dcx7ZBzHvQrAat4ssaLWpDRjfWNuXtU
85clvoNfZ2ZdYJyhp9v5eP5vwfl+NzVW/0vXzkWpw+R7HYPTy2uwCJSI34da0pHiYWCNmIkiI5cX
v0U7V1Ac4rGFWOJt+dJF2UGZmo0GLhJkhcSaeoTOuBFSj/8M7Fa2/wEFlX2kGSvFrlezSfpTWeSb
3TMY3QFaTs2pG6A24wpuyJ2/j1OjFS2fY6n3z8zpAFtyI0OHhzuA/cm2SsKJIW6A1TzF7lkZWSY9
LY27b1oJcmTHA9+uxLLqUX8/j2vdy9sHBsjdt8QNWre7lJp8mtBZt3X4svFwbxUUekyRURcMd9LX
8QRjTrSo6QimjxOmaXIvLCFi8BUiSvjVjWJUNSUdqe2BlpZbxBekwEk/1OJE6lFDvFBUqURemcX3
wDNbLwZJ9GIUqJakhqJ2dveFxXoijStP+Lk3GycI9eJQuXJUdjCrcRbBuMFlWO8Lgsdy2kCF4CEg
eZWViVCizTAeCacc3v7K6CaNlptCrce0G2Ng41j4VRSnpQIKL2g+530Km0s/xph1wSupiSsLtPU5
MfjRAAutSLF6JEI8ywa9CB7nY4L/r/iMRz1IQH1ghrR8uwBG09n9ajWxaLEAt4emNEjgZwJrM7IL
nAbE2N72ZuVoTYKr3A2zLjkPk4hMly8EPYXhoYCUa7EkF2ntBZ6bdDwGs76MFG1pJEZVljx3OzBS
luZ6E1/VA92yCd/A+KBc/K2tQXVEZwWvvRjaj00g+a5qCJtxcsmYZBxcoLd4b81NWQSPk5oYIua5
HiOWvB2hJuFKSjSmuwN2Ia2S2YriYONlEsZo4pJPPMH4pOYGh9fT3MgZ3NGdVnRboysJ/ZrXbAMi
vHohxN3erHlmf7bGB9iE4HUqxgq9C8b4Fe6slQ5CkLFcQg0OliPmGtIewzpF4vph81iHJHFr1QzJ
aZ+9a6KbBrkNLaT6H5ta5mbgZFJ5Q0+VPXbIHrHSfQbzgmkl1tC4ixEK/VclfOi5ziGpkXw9XC0T
VW+YIUrjluyML53Ypbet5LN8ek6wRExuJ6pGRocf3NkdFE8BmelZAFXPmYHjzRwyRz+2Krxu+3Ug
l0LYWbO5Kifo7jjwDM5KY4bxuj4kb0IkLGWAmeUc3FM+Dee0iOFYZyGvoJULYKDnChbFP/IdBWYC
eJ1bGS+PRFDeKz6lZyEJtWtggJ3HAJeYODP2kACZWo/P0usGowYRp2wC1UG8knI5Q5y+P6MdEsA3
1pWGdkUyHHOGxejDT/BRCRE3s8Y5tEwFVzpcFzVvmpG+wWu7jU3H+EngpzARU/qQfdgCCInc4Vd6
p+wEqMb247lUyHmTW8VrYSYWNtLw8ET3TJTH8zoRBPsmdlnwLLeOHfV8/mSvfbFVEjeDXMH4IDIG
mI8mcWRfB1iL04nN7vSSf9loZ2Bis0emMIMdUxEwYsHMEtCnQKA1HGS+BBYGDajFoI7km+98h+f0
G6hx2rYEY20M3KCWDb5M21CTDDNHlFIZ9/v0okASw9ONaZ1ShQTFeg8WKTj+Mv/VL03RkJzK+uOD
ejke11Jxft5GhZo0UA0WA3V+mH8sFPEQ9YKEjW9vN1VRz2SBUQOcf/VFuYzFwbvRJjIMmPovzAZX
J2v0pNLXXJDefoEfbdaLnlUF96dclk9D35scDa29n1Z0ms5NvH4ZdltKygzzLlF79OVNn8iHYRV/
XttxHlfoUO5wkvM2FwuvirH9qt1v2EdznG+PZ6+GTfpK4tESQk3mgPuS0ovupTyb+gptzxWrIoSp
YyU4PGq+EMD4GB4glSXWNCFTIxqAjqfZFZmQCFdxLfwGS6cbhJiHzwrnYiU7dJCcnU7/bRzH36mG
DJg+vORH3tmktzgEa0UDgtIHsPlowqYP+JO6z/18VihneJMQyj2x8Cjr4lsG0BfPlhwUDYDN0VEG
hHqQd+uPXW7Gw9Va+V9soZV4DKJlTx6d4RamxAqpDmM+0FoJrgM3z25yWXJv14SWHQaLW6lZulM1
sSxhQEDIy8FD39wtryW9fuhui8o3rq50FRY6oKWQkgQVjHvJ/thGoxJ3UV+uo/aP1qrOVUPRB4Hi
H8FTnOyTd1QgLGFTxtThjzNuPRuTeJxo2h9D/LEXvJ6H7A73zVptA7X2sWS0VYbJqiPYPEmvEXrZ
yfPu22tuVH7+lkVJh9I5LpOy8deSGA0/MZ0+B5Wl+gdD595/RDBOWFIA4AiHPbdkLGvQQgLiE8EU
URGcrj0sSkCjbn3c9jRYLws0eEaeS/M3nvzXUl3JgOzzvVNG6YRFJGUcwK1+9ZnTpOnrk7+7oRHz
ML4Ig44mUmiXSGcSiM8ya8DBfcR0AZN70c8krpuXg3TyJnLiJQZja5jkozI5NbOfYGKBSJPBXgPE
63MIxrJCCv+mT4PfxAPUphUJY6wUSW4XZ9GhaLNKGxSdpHXjH0IF358bViTla1n9xUmZdBYrW5Ap
VHNwm/T5zTJynRvwSOa8ni2ndMCHNs1s41eR8ixQkcdMKTc4C97OzRadtZ+p16asl/hgphY+fkHo
71X49NkBB65ZcmFmGPz80keWNiR11UjxMuRRlQgEy8k19i+Fx5IyW/ag/LKSjaZ6IMzzxBoPUniK
6gJntvlZS8pf4fwXuQcKR7GdUdTgNrda9v/AWSKygwwpHyq//prz/eTu3+JoZFQWEb3ICY6XUxe/
hWXeONoNhml/PZvP0vk1AyYkKiiosFE79oJIXc0yKvI2inw6vxDB6tT6iFXOnA1VBv7GqVLNYQrY
xMfXGDYNFDAl15hsk0BOJ5NmgZoUfU2pfBBk3QNQJu+dLsQwhJ/9unLXkSGytIH13HaMHl15ACsD
/DK5zDk8jttACEnrfU4gYMp7IjPeabQwEhQgiSgwws6Llfp/Dkg5MRP0pMRcvL7QVSw7tPTJjLZp
SFun+qI5yam6FllPc3M1anqIe0HWACxjoIS1PIuDGwmRRzslgQhNxaKHKLOXpRm9QUB4zFVty88G
HVooNWYsaNZR3uP2w2qpkYIUcZr3sBLWrW4m8s+EaeQb+BHYi3NBM1bMHeMs57wxzxTPqgVk1zcu
u4uuaO8uucKizph35Ca9vPrCQPDvAWXZBp1a1kRVezzf74DaN1X+Ai7g341+W7EFlxnUkjsPlPwh
sgBd8kFMWawTyP7GRo3l60xxMLxXbUzQTRrtXzmlTHimkQHbxjq5vWDzt3LXCFBSj08xyvqu/0ax
E4KVHjeC6aaObe26LFEwbU9jx02csByCtCcvvx1zEGb5ZYurluBRwKWp3BEpmWBnWPJAtqFEZm7N
mjTbgM0A5jsrNo8RUo7C/H0aChIxj0Cm5ZlG0OYbBHZqh/FhQwm9m9KFXN1sYdzlJNSf3bxBTbnb
41bvjauk85ZBrK+rs4BVqeiMuXFHcua1xIzTFfXY1N7bd5gcVVwzAPQdg8L9V9BhW375YZm+C/M7
/o9r5c24AYRt87mYYwEOtKuwVdqTBNAyf74ervoLqS7kUIRvBVnhZWuNOKp8jawrXIrW9/xmST18
dPYfjaI4bt7KOXsB/DqAr3ufC0vHdBR/I5L5eNcs5eMGe9R6sO7REK4aq7gz6K3B9owquvZCBSid
h81OsPUzUWDEjdSI8AybxwmS0JmP6t27pP+cKUY5nT3nggid1mWPDMXEaG1aXb/r/WHglG8IxEzw
AMqBDJIJ9j2Tb+cue3CMP1y4OjDGkZ7XT+8HQpUmRX2v/sx6Y6gPS2dIbnPxb8cOQanlPvq996tg
oGLjxqbIp9unXu24+1O6BCNn8eo82af0WdOQq3UwnL1N4kLlEWpnBsXxjj1qqoy9NHABPeOsaMDC
AzpTcQE957OjW7J8hHQx2TO7ip5StfTMEsA9+5jl6+oLj2PbRm+zfMasEtk7LRVZERH/Ty6b4iHa
GzjzRBd+YbQt0GJY9GbPr5VGvcVlGRDkPP/lMY79x6rbKp6cFC2kHhgnFATgYfH+AAop34Bg32CJ
W/2MDICp7IM6/BWU7uvCPo7TozhgQsxhCs/a5XCOqM26mvbnHtZW1WcrKQ2j+PhWWXPDrqsneaM9
CWdLzwXnag0Rf3TfiEj3bPTJkFowGxTBDTPJM9yPVtFtixdLK7z6uMZ4mZz1BUK3zyMik2TugiD8
PUJTzkuHpukSf+gPClL088CZBSUXmzsq96Qu0+IpkrmdzKEyIw+ZwGsrHxvrjHrKL/vrzmefe51I
nTBCifdsSy/ywvUy+UhuPnu/fNTO2Rcfu8RPM3j8k5yx2+ngDsN3n8reScZdTWep60oiLyd1FlCx
0t3faTqr1TZz1XJjNVVJM1d4zGoareSYEeMsXnoXRxsbE+2siGRyZmP5WgQVsTLatXJ2r7geH67a
LwZF7B5VV+cER1+2TUsc38VDCT0x3SargaE/FpKWDWiPlg3WeWoFHHMAnwudLF7Bk6iBB8RcX/qF
6mBBpSZo9q/YD6iBWHm2ZXnDQ4ACVRGO6c5gYsbEhNf0NjHPptL33+Z6jUTlFRBSVpgzTPWHgelK
Bkfch4+imnIvbDSbc/MSYFQ13KehReOewW1IeRYABZH5V/KjVPwL3wscruYUqhksWzFRK/BT1VJo
9+xHcUwiz5QN+wSbleEf66nNoGrQ1p0NYLCeFiqSciukpOM5NMCa8jtj19dJC2jcYtYh2gIlaMXK
dLKww9A3uvCGmGOWugCMwDO3RGWOixg1pXUuBvgBViRsyeM7PEPVWbdaqWqgFqcSBqCdKH9uH1Wy
EtflKqTdwUU/MiZ7bKIESn+FYAu6IpIXVMaN/g9oSpS0I2rIbtpzY61Uil0ZDatNwReYl2Ve8ASE
fGxHS1/8HEWoFV95Vat0SvWPVw2Y0ptGyKZ3aF3safRglKTYZRisOahp5KwxSadjjx9K9rbvm/Pk
ZW2PFH2Ffm+hHok1ldESKt7uSMlE1dZhhZmFuSGc0L9EJtqJ3jXEdBvpGZDdoSERt/CIBaTsT1F5
ScGgV3y2zYKtlGv3A+BUnY6DdFDkeay0GJTEc923IDFygctqYYYqNeLkL0MQGyqmhxpGsl8yiQYK
MBsYIXWT8zMwpF/10KSIDEkLHq1wgMUC2D869Y4EdH3m5B8F1fu0nACu0y2ZuzQ/RTjek30/Wj2B
3VtMPVFhWHV+SQZfHxCQ+tJf+zHw5T1ob9g95LuhUaPlmD6piTwGWF7aPCc7LjumVCNKATSpjLxD
8uoyGAC0FzxczrtCRW65+kZaNdCKzUYAIIaHfaIyWdeyFgyDnj24o5CiPNE+6RZycqYKn13/ZDJO
g6I9YWRcEUFkwjIbvahfVK+RtVVM2BNelyWYfKwLMtQRJfmzQCsPXC/9p8ER6tigrVxdNo7IuOsu
lDv9jQELS9mk7UPFtFGUgBK2x++VvdPcK+/XaTJvBW8w49RSUYJuKJQGnwMpKdgn81bPldbjPveC
LBNbcZ/Mv4Qlp2b7VrnzOXFY2RpZham6DdQMFwUnVL+HWM1oEC8p/Ymx888SuAGejaABTzhs78i0
L7Z1x0QhCoSmT+IYAkuc60MVLGw+gK4VtYmu0edkF8Bbm4VSFZDXZB1kH6/H8Dufb3vJdpFbCE+1
pb1+Rbcv0tw6Sh2w1vuc+Vx8msoCB55uI8VITavZZoraQOjOmXCR9PCvtK7kDNJapsFSUUJ8Ghtx
ilO0q8yV3TmRfCSODWRbPWteU7lYdKM1HumL0xzStmphnEW03gxmVLcXjnG2MgKFWbATVxSn+6CN
LtjVm/IXleRxX1F7PqSAHjbYYGdRJhLYlf8TkrDzGkzhhNFdKL/2S/Cv5DggMQ3erWtbBSOfHqE4
EFqJR/zO1aWEuMffSy5q0rrgAGQqcaPmk9Mrk5IOta8/orHvc6osopf+pbFUOix9hCvGZj2cHnjE
ugSp5R3bmzSBfUedIYD26eRF/5nIZqZHfncis8SRoJ0dSOZGy54z1UJCeImUwddXpKurIxpJJoQQ
jz02Z7OmS53CGvvyb7P/lh7tNJZ3N60nNkWn0HzH6piS8UiitQbDj4g1dRs7oJ5NJsWfUwVaH9mx
We98kvpDesLiwoaHVlR/wa2tRr91H6BE6/NEVp+Xub5JB/vscuhP7WRL0PePq4KBnK3m4usPibXO
cqHFo5ftHjEHyDmzhLQRIuXc1DwRwv6lgfy80RCyC6DpSDHM72+NAiFZ2P8k7qweGaxDHFOSu6GC
lrrmieob/BvG7J7b9iDFJnMY4jWfJsDVATrEKoBA34U9CP6W5Yqrd6R5Ow1/bNF5H/TRzRpbS+xQ
OC74a9BSY5S+6JJSoItevjoJ7Q7sKwR/FEAOlhh0qiXKazmzb+5XUJTDT88fWpzWjasQJdx6XbDc
B7J4DgOSmSXCuk3bxUUPDWDtV2xX07aWlhXNWUsQ4/cr2OpD1yASgTG6aVYhd5kowupXMjXfKRU1
qeGmYECirOh+onA2ZguWLJtP1nC+iadZA2kKpTUkFB9/UVzpsp/hG0fpp8m0IJYaxx/3Va4apD8O
QnPg1uFTl+LQ9oYCJq0nKOvqR3/XmzBnrSSCpfwFxNpwtOrBcnOPCdhncIUVVjYNN8TCRGRgeONm
8qq5L5BcR5PPom9wj18O0e8nAyqq67rpnmrmzp7nAQ650hm/dD7hEmrFAfl2in6pWI0daA4HF6wL
6fLeutwVQEphyMMMe8GqqbOCOP2VNoLIh9lLkjLCLpbVYt7ZLE6Aj4tOuwzfc76yYzkcbp8q+31O
oSnxYOiAfx0sJQh2hariYU+troDgc5mWbm6h9HMtvdF0ZX5AhXRAVS2ZUKobhf3vtqx2wIzbrTz4
oWSRc5XvvpSuJ6EtaADvIfDMAyiA69kd94ckN3rqnCg8zR8UCz9cRGQ4jBIQ0Hjf+9xuVu0R+7fI
2Ohx5iINO8lYCmEIkkjEQ87BKl8nXPqUwPC0D23YdM0JW8Xllcv2XMFY7MwCx+iKnwppmzMCnQPv
ZWbKTl1+i6Cy5XQNwP6gK2vV6hBlu0jRbZ6y1HuDC2lRZRY85EtF+EsTh257x78siDzgU8+WA0to
nPx0O7RQd4R4mFaTQ4KDrTmcu1TejvUh2AlQaAtDhyQ+VfWuUJ+p7mQPWOmZWfA6alvnYO1cCimO
gAdGr/gTBxIrUAYmez83SGYeAr/UEd6eAdQ/Ty5+4Qka7bNxaOjBzemCRNv5+E5amJEZzYhIaBOO
+vc3/5A3SLXDBDpbXXO++5Q+1XgiPUPtkjNLoCSNH8h1eZmj/oLGtgeZeorJ04VDN6lOjps9v/sM
qt1eyTVLwvSnE0/GfBrHiKZHZKe5N3drJfHuRSzBN6Cu7dG/EXFvB22IzDoOdo7g+/IgmkvvBHgO
NbpyeGa68ieQsihtq+DpltDhLaCAE/EQKI6GYX/Y7Wep+IEJ6v0OsbRgAWFBIHEiaSQ8Resgp3Xo
B/sH0ZNMfntDGMkKb9HrAoDiQslSp377Npl5nGfsX+HIajd2/6SegYXTJqbIDF8XqI66myLmhjNA
7aSrOeuORDsy5vmHyqxAP54E6nmgYTldWtMnmkjzmiL4/xC7D4O/TARJR4BAU3Mn3uJhLCNlqO+x
cuLyu2IubwJ5kWGzT8wz8QZ2opYhlJxxwgPpmWmTwDkh7mDyc5a4mwtTmbgBnSUUKNEMtwyXZrEV
CxoTvBUxDdsu1YtlIj4jRoy6Bs+l2LOirXDZ9D/rn1Q1hOXpvr1KCxO1Zet+ZrsxtBayQo0+ryad
Zqlv0A4AhUm1tj/FEr0AdQ37pLG8VjM2TnvLuoDrVFtXd2vfQaXGw4XYLnCuIBJrmzJmECYKA7Uj
RPTeUt76yQUjxms2Xb2afTA3yx3wV7NtGnZ6HE5UCNSVK/C1bmNuX+VjP/ar0WGUEC+V+Qxq18Tv
W4LKNA+449xT75/rw7iZ8LTYsswOD5VJXKHE7lyWlZhxWRqaP/KIiwXmBfbDXiME8HOTMCHKRsx2
7oOAOKPQUhuC1OytjxS430COWYvSY5c9pT5XPMLgjoWI9Y0m+77HB/k5Q5EZHBKvya3YVNrMjn1M
TV5rIUCZPndSU83Sx05bH2PMPQjZ3PZwJ4Yz76yH07CoTrDgK5s2nILo26UwxWNKjMR31jiH7A3F
G37NgcNtoI3JBzj48s6VdzuWrfaDDU6f+ej+YXhSKIgn5wmF20yeModvYPR0+m3bES/oBhdYovMB
ljoaSRj7vBo+Yfzxt6jLFc8Wbm6DDB5YeOvzeaklVwAH9hu+OfDSlIi8GrhfVAxxgx1XirXIehKR
zjLmIlbmgoDu5YeNgDQfufCZMQE5UaBIhNWA70EFn6HPM7fKDz1CpOVU/oqO1lPSJxH9ELBY0aGv
zhjvcNWaMbo8o2F5B9cx7IN+gMdqzJeaKzn89yUDMyolmcY16OYEeKMfF1ShVjsjG/EV1Nw4w7Zm
Ldb2M9wUUx38sIcs/9Zf8O3vOm+2mxwYo7zkgFvXVV4oATHMo5mXx0uMmXhtDydP5HrWgipr4qcA
yZYGo88D4wOAs9jUUsjVR6qqhCOnsTocr9sddnn+hoNgL0pXb5tc5G59mKBF+wXz89MpydWUohYI
xFUhS4UCzpehgP3/RdJs9IoPlyXZRQutrrtfXoBwzJQCdPgvG7G+hqsylo/jFE7ijHOGpf/aOEtL
t5hB4GGCdgdUFM8ktpig4L/rr79lczIedO66lxGlBlsyWXVMfwEtaURzOYnFMF2dnZ7UrqOGVahe
hxu5sIxeFo3YYKuPwNPROnmx4MDzSYb2HKWJYipXIristEWzejfqUIFlxP4zDeA3yO8shnWyeVBs
vPdW63SLyNunT0FxTZ4PLrxIC9K5+98VfnFw3mFtMOS87CNI7HBeqnGAPvRSoSaTKowokPyvjo7N
KLItgzapdd0fJIWmsrMym8XjqyM7jVhWcOqrh7IBsUQKaWTrVaaDje6FdfPBHt5/RU7EO+DWgy99
SBaaKQnfX3skUgsfTKCUnZcSitHmvq2WBvADXvk11s7ZKTAdHTTD/jnoYxM5kLeq70wOHNDFkdxD
JnYV31M9ouz7FVgCxUF414ZW6sYq8z5FrMcad8tzyZ5UT4TyuyQOJ/NtbKD1WTGj41JzqOnTZ07B
ylyhmCbW57d2I2YoA7RkajosGAI6etxXFIJYG8xukvsC/7wHYUgxUSj3KAHpCqc4VjOuGMDAI6SG
EI20VG0qUlafjkUUA5UQ2K3aaZy8SZ0l61x1BcwR794OAOEC13sxFGMVOOjgAj3xKOECuLbZ9yty
uXJOyE2IOmuLYMB9uQOTOS8u2FFz62tjIsRDMbUxqYrAqw0ojX/XmPBISdcZbZejZBI9uuFIw4IJ
vaQysfhuMyC6OV9mk1FI+sGbRC6f7sdppfG6SbL1Kd4D+E24Nh1gY+KfpFC+25NXHYXiGdC+rw6L
DImbKDMrXtU20yGHG9AUajbRXdIwPsGcKJD9PHB9limLVPIPovHrruC4yn3gMhCNjX/yHHzReBeZ
OX+LBZ/17b9l0h0MG0xB1j1zgFxxMwUqse9j5iteQNNV9lQYIq9ckLetirNRCCYoa2/48a3/XXPV
0RBzzw3d443x65NeYysR2oSeFQZLH1+zDvw+Gs8mblMrUS1+bLHbPxBkiPoQDoi2k8y1tHms+PVu
GhyYz6manETwVpFhsm7b3le94J42arDve3/N7lDucDGranvxhEN+3x543vOiguGt0mHeYZJ/nhA8
dREYBL6vhOHBfeMtcMRAgT/SQSqwMPYRSrj8DTrHEfoEdFF9ceB+sSqHItxwhiZZyqskZHvUQEP1
Aa2NQxUTSx0G3D333yh+wED+NXot4RLu9FXQ+4nTNpJg4yP5l4/U1v8JhA+R/zQbu9qEgcwpcHZY
1K2d75yyReLi1mGUOdQP1mB8pssqO2ZK4hlUxrMm/ByWYRxIm5tiv+pEA/p75QCrDipcKst5d104
XImzmpy5r0LFccUT2iqEJdXj9yuS+vR5tAisXZx7qvo3MeRMWGKWbYLcqAhnwnVgk174wV3vZ8nK
3Qg2E8BUKArnq8b29fjhFtgez1+XZbkTfdPkagFiSQx1IoopqqO5eKKx7cPfSZ2iIvomyHNHCC+D
lQGNgV8irvQYdL2kmrVit7tI6+zSV6wCJY0ClFSTNMlDdCqeyXGygjVQQGiiXmzw8pR0ZgCIhoCs
BZ/jJDDkbR2gxCkTGD/I2Kq5wHmzL7LSF4cbMJCpxUl4s7EfSO8xW8iiQKcUxtxSPwoS30ZFW7Q/
vePmRNcuu146TiKTHlheQ+TTnYnjuZmxmuS6an/OqTrf8hDGkncithuHsoxMek73pOhqjVMAzqFi
8rlS9C2ml4w2nONBKjHz9THlT0pf8CaN8MXnVv0tRqLP7KNTxoPKKBS5ShZCUqol0dLm4wo3mrVm
zC6jXeiednmJz130+xRCdXxHfsmuPUP58RuxXjIKRNr6Oe6Mff8axzo9XFsibyHfUKmpySxVQvoD
k8SBbN717LAtz3D8YL8G6fIrDhmIJLgU8h94SF08QDQM9Jc5fNyGWwGSJOqAZCOC6uTtsVaR1EEt
48rPjYSF9Gqg4nskGPrYQXoB23HLdCyhtRXSPC4z33SDMbvED0Ar5QUg5RnRFKLn+99k+rktor5h
ysAndssovWYDtgUe7VYQkIBmsIy1kJy5TSJ+brmAc6gw0DMRdY/LUMxDLE3fzHKJTseGWyejNqFg
AhBfxS8zkskxahliqop4UQUvdBlhz3Iu187YVhpfEieyvBkT/JpgzqFqYapFpnUQDOKdyeOvk8Z5
F89BOukwwI2O8oITbEDN1/3EQ/PkKA0BNcPjk3VkuFd0l78wdH/zsDccifqWP+D63yMTI+5R4wG6
juG6G1kBzb4AaOAlcKSd6cKt5S/40SA+hQRBown+bUOrkoF2Fn3IPxzQUOjSuVMVTqWGPQPiSTmW
gY2PUD6H8xZ82mJcbJqN9iHRA9e4uBFWMZ2p1bHcy2nO0QN7kHnL8CGkD9boTw1LBAvr83H3OpIe
vmU/ecGqwDu1aXkH9ctoj4V/397zRnAqD6osKhiJIZ0YieJxgyVxlAG65ZJvje2n7vrFsFzQ7Mix
T/Uvdp3Drx/qlw/mf5gYcqATuvMMw2w1l5tO+OyEnGpdZRA87GeFJhs0BgI9fAEEIc0H2Kvn61fY
BoTvxJz03B+7DMQcvPeX+4aDOcC0xbPwiwe5Obt+bUvtz4j0rXl1OrK0kj8s9ldJwoy4tNOeuCHe
nMWgTCZeZ0h/RiukLeRBkEcHGfBdhroBJHINiKfGnEqdaN7kLfJhccidEiVrckQvQ1GWWWIsuxZm
cPsB33oDMASeWuHfGlAxmgQwinW5TqC6HKkl+eoe8552EmQk4tZEXAebtduwKgJFrkzTaa5X2FMV
J8bp2V2JOlcDBEyXlpZaT4tk9BMsynmG4QsrAXZaBjQRWOdS6Is0Tezlbt5upJjNjzlEi4ruhlnk
1PgmNLt2eZ6BDZTQkB6zpF6nhqwoWUzSEciCUM+VuBcBWYfAOAbi6rUTj31VmyETpMz90UsH3Loi
04UxvbLKb/boxipsfvO3lm69BQt+ZoAryFRZYnJ8gjetmQSAChf+e/zMPlY4q0a4XSnjQrv8trE2
zBrMHHwzP5FAsnLC5NuT8stsn3lcxVpoazhMUYojXWB0uEHHj0oJspPzqSyA83/xb9BMFQaYVsVL
hWtqYsI/ve8n/NJmK49IbSDVSiWHbXU39THWwktgYRzf/ZihmS1yf6i2S5s4JoKs8ITgcSZ/2aW3
L0BuIUUijqrY7b06ZqQPMyAJr2OSmQuYnlsSOA1P9jn/TSNNmuG+/oizy3/4ty4v9JePa/t4lyu3
RcoifKTtJqIQzJLsKRqVYUZDGZEMiLibIe45z+GjgLMSrL7A0Nu0PeoMv4kuAWPMT2mkfOXxiNYz
dgqQYMEfflY9c6qYdmlQsrfxF1CtpVjPPrQCnpI+xFyGcFf2AIxu6YR/SPwGowSZMQYwxshnK8cv
mcjKuMvhWMkMaxgL0fhgKsRw9Sw2O2yr/ne5elk+dV/G0K6HdnRUZ/GeTKY/odqjBl7WD19+qZoI
2UUvEXufvI8MOy9T2VzebyBkQaWiFVDQIb9IAbLEyI3aNb8NO3fJq80vayCNPy5ALziKAlrUC6vh
LKAHRYimERS0uzecO5EJgxET3QDNs0EZEoqvPsWvY5ISnmRX2H32RnkSSECiL4PMC/+JIdHpkXGh
wtPqbO+UncHoZwqVw2hbWAh1ifonHbGh2eEYope9ziYT9fVQhwKxOiaiwZQUr7u56A87XWQvJYoC
LjEMzlIRNurOnXGcpnX2vMWgCdMyqRvVyT9++N4DDiJz4hXYpJz2NUy3oUc6dFHwDA2ks5NqW5qH
onRzqVLwAGsM2GTk46OFtVIGv/7c8j6ph7n5GAn8GA5CFEmzzXPTguvVJOgRj1ZZANtSROtdrdPN
niyMM7UhiERXUYZCmdcMhWU1GxQ8B8TgOuhMrsbb6AigPxTBLoD2g/P7RZEr2Mxfi4bOlparL+xM
w7HvN0JqaCRaOEGoHd+Wz0Ek+RV/O0lHLnV/OQsUZZTLZsjR33q4gMoF1e4PU1d+AyN8F3uIoDBa
v5HwjjAVlgUOgn3uVk3KdTdBRyg8iWMe0omE6pfhvwycwMr87cBazCWVYQzpQjRiW5XKK0O7hIC2
xdSo3idOJiTo4Hh3/ZOQ5rbkqEFx1Qf75f6UMa5fJL1w5Qp1F2OIHhOqZkb3b+QkWEzTV6XmkD8w
Qc1ILHhlWbLf6qJjWOWURKAbJATzJIVkL/p4YIe0JPMYmeN6OUJJ7m21PKVj2tP1bB6OK9dhoDHQ
1QmduH/3vHI7JClhM28xWe6RcdE5ThqMLX3h9l07LImLZ6j4cX/3rAJKNWwWmhO5V/SMa7fYT6hI
mF+2TNOlJmJooghkcLnpNX1hR1JLz/rtfD8qoYdL9mgENM4xuCI+eQTjUF353RzTwgA9ZwxQ/jts
HkLZCwIvZpADTfNrRfo7ORgfDd0Zd8yM5YkYgAwbvuyKOIITrsxPlq1ffHcv+TK6Eew/Ycs2D8l2
UyF9WN1+cpU2/DXyjIl9O6mQfjScRHCDXxQWU30Ay+MB8uQB4JPRtscEaelLxiYBjhFQEK+2jLuJ
NefqCsNaBgjIFnYo/bSeIuMCyUjw+JdgQL/UDHotB7zY1R2/iXly5x4+cEyhftzkkWNVppkWRWZi
oIkxJGib3r0/KEfiVUIKY9WDxEZU/AkJRMppxE9XpLbgddSOGxaZkVKGxBWH5w8q2ihbJAnyPzbp
HtU9mXa8sDFIpghy7gdi0nyaUO1PXElYzTxPrfwBjZCNrT8wiWxiz65Tgtk757Slgkkkgil2VDxZ
qgVp1Z5EiogEvXvTLmuLHLp3aFAovLy1LZ0//EEnKe4jSOKctu3tLry2q8vz/GM3gPdHeN86cOu3
K+kHp/QGhVquwLwju5CW/CAMwG+zI5xuGFmmGMDkqsVP9GJmOjuRZpOM0+1eONKnTYe7HoLXKPFL
ee+hyNF77f9zXlHsVcHEqyyn9BSvC8t0Fd5HNXshgUUJzN2WpTuX5luZ8MTnxPnSVItTmmJFLoFN
z12N1r1Ucm4sxWeFM9QoTAHuXnY4gtVjKY2J7j+XWb3P/kz+9uNEDEbfAnCh5X+dwq3UsZS03HbL
c0wKJah+lHwW4JPDJguIk+HBewupTWa83mCByxgpcQYtsx6eLtiHbawU4quEaKP0AwutsJQKfUM7
5I4/YbRqheeoPv/x1jG/RFh97dUXPH8AW2MvlhWxASadhnVCnf4GwEo9pxfOHPAd7eFAn3Vy+gm5
ljH2od1pXxeYZT4iAgFZjr1yZAUXGYMYXQ+STA4BFzgdecMmWcM7qNSSmUIafjCTG2DzVuL5Qg0n
XZsvWICgpl/kPfmXOe2yIR1gxn6bdSihRs5jFMTCk10rWMxo4SRpnWJ+zjdXaMcTL+Pdu/9bJoAY
dRKREF3LaQs3a0JauoVmd9mFTDBDraPhc2g3JTA7O+MCq9yY4ughed0RLcQHdwCL8LUQ0ix/FEUC
P+Lel2WEDKp8DQwKIBz6Oi/jEgO6vSiGvcNUfiAzL0+7FOsXxNIwhJpd1E9vahKxgOALYVaMmuqi
FskbYMuCPyF+bUlWRa+ouE1jt5kmtaUWPjAWEJo9UxrrKbdixAofKEzepRaUSru3fe0glHVKY8mc
I4fEphEl/F9DFgDtKFGGO5N+LsyFpvuRg9fHfl5DazbgWymxk6OGLFpRaaWiKsr1FoKOsKmPsKyA
OD5a4OiaGchyBEjQ2oS/8zmQKykBKxH6iZyjMKJG2tC12WtMd7qDUvQJXsr0E6Zv+ORhNXKvqFD0
Mtdzdewo/cFnU60W751byfdpesp8OtdP22xhslcao4UIzO70dInJDapFlmmbBDsH62UkQQMrK9Vb
a3bZiOiKsaCu5EHognnm2hnPhikCXW5t80PfA1Q2PiKM1QwJbMeXeYgSqOImxMiAXYbSWe1ObD+R
ureBMbveAWuSH1Ou0lUTdG6zX3iaNa3ctaQ6w+58rV/GPhY2aHJ99+IYdTUnA8KUZdCWV/WfKezq
OkZU7tO135LNVUcSdateOQbMawmIh7YYKm8KujtA+6gt/guDXJ3XTW3mUAoVB5ZM3trGVcpfkaeY
Ifcb1DLMVbnOpwAp7/GRekV44nBDvhQNaAMJPAeI80VyUQII2OUFUHxOui3CUkEHSL7QlU7rBHF2
SvEyMfQZtkloV6NiT697fbgr6F7X8fo7OKM6UtBfb4KtE9/3RmTRF9A+31CDC92qBogvkRSY+Xjy
2lnAohJeIiBTE77vdyfYNFvh/f5lzjnqNqjUmSznwDVq9iHiY2BrYh+zotDHliE13Z2no6M139S9
5VCRA/uFSOkcIMmO/zUZEl7GnuMAVTpcu1hHNrH4F8tLC7Ek4JtGYExHVKYnnThheDK2jH0km1Yt
R3kmBVRzJd7qAuLuYALdNw181Anye/jGvxAeTFnaKOIKpAWR+LlDp19AHCAue0iU2J2XSDD/UKly
p2uH7/doHLc7821x9M2I457HotioPIBnljzeNP0sFc/YxBnNgGL2K1Bh33fmtQJVQcgQDqWtMyUt
3NRg2OM/sjsyMn3KiJSOuKYtHuOOYo6tjmAUVZ9WJ2486oJEatoqjI0uWP/5ecBQup/DrQiE0J8n
vt2Gk3W2HrOBHkMZU/BJyh/EjTMbJOOXbETOsY2UPV5qPfbDuZZjss72v7fIzE+LqPAnwwFkM1nE
gkfnpzVOng7HFuAwDqaz6Zx0GwqbmnMfrcpmh8rABCIo+WOohVgompH6weSafVuFPU1VwfsbeQ9b
FhFvDGsoyKKR+62O3cIViADJvLaxTbqBFXnaez0a0RT0TBirzwfFp3+Ccx7xo2BcK0qo5yhL/CRK
UwDiao+Jqx0LTnc5NFbAxaYmppCsLOOVTUxAbZ5C/WRQ9dd5iPuQpmjYMtKq8GyaR/gjXIBzq1X2
d6d5mqFNc57wa5R83fW06eXceTaSsSu2MdiX+qK4gLlVqb6c9PDf5uD3T7fp2YUrTWhTNwoM8MjF
hxgghz9/GCUv01Fgi+oHxqzMbN70he3MCQCTsiiE44TQqSwGicL6H3XIyINoYAGbGvLC+ynQqoGn
mPHJ4GjgOnwwCcJ25nc8shYTRyk13fmRlqc6Q5qpduMR1eZvWu+631iQc8FG84WbsDBOS3cj4Jix
yn0mOdrN7fJs6isdEILPnxVkVilf1QF6wEb4WWcen0eK/OEgWDRs7qVXPKYVeA1CxyZcFMbTkY1M
dotPG6TqcbfNAVGy7xNUulcqLrF9Mo9/PiV5ErqDIDeIRuK5J9V0XIeXbWgnqP9rQBOWuZd6SsWa
01Zq+H1qSyIxwucGGmR4tkQouIQRJASLO3NShCCpiXdAl89knNnYZ+XENrznULxWPtm0IgavYKoT
juITPErK8W9KJb0hWak2WC0Wf0eprbrB4cqW+bP9AVuyVvT10MJAGuXGw5wybXc2NgR4TZWvq/NU
ip1ScwtevK4clIuRI87GlmJwI77eqgH+x4XMetm8LDzEU0uOoqzrYipdvzHX8w1j26ioGYcz93Kj
shY2lSV+xq5vRgenkBBEuPVZKcEyvHm0fL9pd8KQf6xjkuloTLFzzGb1328KOEom1oQFhvKBn8kr
YYRh3Rwn7BEfd6LLgf2qQz/JZYyLCAzmrb5a5aPGItLow+WtW/qmzZTugiRdvXX/Dxy0yqPYuDf1
Io+EMEQQ7JUPzj5sDQJtPTpzQTBEGjwfFwInT0rnh7lWp0mTqGtZ8d5YlCUi2PNTi/gFtBzXPGkI
iatTMBz1/sAXfG9GiIbqUn1K1dwa5eCbsxSKOQPJFza4roZo4DQn3W88WCVGMmJqW0nEUkt6NYoX
r2UvFJBZ0Q6VnSoBbzT1slIfK0LkQ3PPHno7Rl+GdYl48sgCBUwZRB94hswBkYmVQQEwEEEC7aFU
wE76kzr12nJvlI+69gqcKFSzXreGmDTfATvAsa8NMCOJ/BtTdZSxAFC2/aDwuH675TGKZ1Gr+yV5
f6osNguHynodHa2BXZ1bATNxeqnpguZW2JNWOHy1qzT3DM0pXv+pTC2CQO8Nthk30QaoI/P8NnEV
arLwLXGdTwQQAw3h/7nuha8tE0babZjdpeHO3DCORJkgGzkFdqk6twi26xFQ+v61sX3slfE+0vn1
W2AemJCee41nV8sxleyWBeCTgnNe2Jp2TkkAj/stDNXYP3XiEKVYFn+Hv0urQwUBcqQX+rVLny6/
5n7Ujey4ghbNb7OXDkgd+mN3DmrXjaRHXO5I7A97HhgqjLXH3j5bHNhIUkMdBHQQ8cnKpPTSOn1R
g1X46T4k+d5cFBdmCR78AwLNunkzomArsKMsliPfZCmW86p5aKriqXFgR2JvenXUSjse4m0O7BPQ
Dmkt6VuS2E31jkL+x0z8cPMNSJYL52zEUN2ec13Y0o5zh+GzUuEdfsBY9WIV1HsRGrkfMgZEHI5x
dVx3vC84Jp6Bq2zIx4Uo2Shg+LjFXS9gIX/KE7ztaDm72QUiFlfjc5FgeWzCLEmXKHGNnhljNN1i
4n5vWDbdOP4c8jklkqscRx4mM7ywwwqR4520vw0ubRxJqtLw8g2yI9XlfYKnQPoaZfD5PlFPWho+
xDXhk0LofAnM6JgkMsFnZYEI7GFmqpw0hQyaw357SymUgDgBfQV+nLb1n/gior9d4bdJpXlgDfNF
xw9Qyo5R2jwl9ppqCgalduiYgKVE+HlbZ3SzydCj6U4md1rLng7piuebosP7BYYMUbsUHXNcYhiu
bqxU4HeucnTgSYnH3q0AbEcSk42OVrYCfl1abFLw1PRApFc0bVEW3R7l7jb086cnSIsNT3J3PemE
aKmPImR9sCvVQoziBkCsNRn7pPWfdxjW+qebMx2tI0WzfNIRe3GAjKQYcLtPK5vjAiNIGHEn7qqs
xjU7jfSjcnqgwnNv5YMTd0ow4UBRsU5cpxuLdj6uiF9+z/kDZ31vz14gVjgMq3HNbYZUib32qofT
/6QRnKUIQtl3cMe3v6+ZcW9LQbrMCuCcvTrorzQ8tkrzgTSbOF2V5/CcX0/jNaWt0DJXdgLddynI
a1qCNaxtCtKque8nKgGQ6/lphDRGYnPUAdLDV+p05q9W7+GY4qbHn9NSyx1AwHTqINGO6UWJuwtR
u5FwqxMuKKvXy7U/5C3Jg5rg8QhIf9HRFpIUc3wV5Qvf/Ffuvwa3bd2XGhVqIbLGAfF/0Bz+n6e6
C3uezBohzk1xEe3c/3ziW602IwdU7aAyEnp9YZEw1F79IShE6uMlKDzGmG61en7kEPY9rZI2z4vE
8zRz1KMdh9C8Jkovo5fbIejlDt9vqgB0Y9tjPousOkUVSMjpeSOdKF98qrChCuLFhvOyitJdVxBC
gv9UrUsMUejyBWWbaevEIjgnAbPEhygGTbiDhZbg0vS9JEJHJTCCRfIwk6AwgLy4uO8hgRmTVsN4
oWOLXBc3gILpsCXm7GKcjn/vW/BoDlfS3GMJFSnwC+itxNkMkaBdf4c5c6Dqy3XsaqXh+DYIH0KS
NL+qvf1TibFGk2HtI+7TyAcAAXZ2BLYnWwAg6sC5elxsNSe9YpdMo58qtnk21im3Hx9zaF1C7rtx
pMS0TZP084BsZcRInbpJxooo8ztvyspKlzED3a9QoiIZPD0un3djdCUmXdG/uy3RwJP7liIaB76H
k4nsTT8qVazhUdYFMDUQaJzM5mrb03NLxtA3SNWKqsNhhZ3b1cj44jPo3DWcwOW++rad0ggQ/vmw
ql3KPQUC4/0VkXlTQCCn8WrcBjgyAiu06rLNPynsjGDRSxxKTNaGDU4rlA1PbdSizCTbuv+WRdHi
n4XdJwkdk2am7Xnc3ymrJF3P8MQPOIxmR0EiXdvnqM3hVG7kEE++Ue7uo7byR0kvecrFhy6ZfYw7
STQ770kP7hlGVTRIJLpVBT4K4aWjm+UTT9ii31vrNXEHIhrLryh7C4GM7H8WZmWzpmGWNh0i2zLl
RXgPk8rlR2LebrjsJhHTyu/sVKeU1biFUxdN38oRlqTiE72jL9Ym7kmUTgdlNf+Eh4Vw+ZqOoOZN
t8/J2mmrXsESMHm4lyR7+HdhhnKIPfShyTr21Hy7Q4qJQ4oLuXo5vS4kS9NnK6R55OXD/1KQGvk3
K8szmAgZyp1AZ9CsPt6hB0tBMJu8NHQkXIeuFIfCcqV/T3BCvYF7cY42s9ki2pz8t0ROu77NEocC
WWFbQzc+zfVqoRwiiW+oAYJdgzHjnqhaiTj2MIvWVXph3mNaTTSPBkeSn778InHZQOeHrj9NvLOk
aVl6JltGwA0wZtRQr7o2TlbppRwU5eAvBiDNCWuM+ADt8y5lYaw2B1Xw8o9E8tB44V/BPg+N40Ap
6i5w33RhUosQXkwrWsbJVRet49kQaDFAXtr99naCgVfigvyUYGqUcgCHCFsRxWy0X69QS5dVWVAS
J7Cimei0CR55P58j8JQsBPxY9W73uNr39+1w9HzfJvip5iPcAI9+UZZ17dObLeRoiXe7FoPdmGQT
ee1xzgvVs+W3t3b6O+xvOV8mIo3TuHi3G6K/QdxuhqLlYCij569u/MmFBAemREWUK0Ri1ueq3jm9
EvsAySv1zz3T4Q/apY8Wj7LdUP8pjM3uFsm7LWyUANkpUTjKBmK7DTeosZyCh8ENQs6SP1ngyuPF
6y+b6u9pqDK1m9GTGjl6bjoox7G+trPYrt/esU+9/ebXClW+RQm1A5/zuHhEt1K143rqnjZOKo/K
s8GVBDYID0hzHAZF0BXmkCtyeyP0McLiE/h+HN+Ch792o+bWQZm8KUOES+KSy22KSRyxkNZYvqVf
Bvy0yN2HJWvJdeOM37IzrJh3tRxPlEMQbrIMeYkpD3FuOnBC1MA9R3XHZLqwM684F7IV2c4Wjw7z
3uIAZocsif5Dj5eNbIkZ3CXgLOjDDowBsKKLhS5o575SXKdyoEgpRE5Bh+9dTrDrJCwP0eyIhRtr
hEeKWf9kBcgVt3K86Yy/yMGy1lXS1UWoiLyhJ74AEmhvzQytFDpRo1zVuJFj2TZ8Cqo0UPKWsLpQ
S504N4HNgDXgx56/jP7yshtQRIoYvEzAvTQtaL5K/JPrJoNG1EYUl4MwYmzuOQjPF45RFhqrp6cH
YMSSVxnwzTAyaAnP6KveJa/xqaSb/ggAMV3GUE8SAZlb/10nVOcdvMAN6OydXuRXPYf0atw+pSKy
zTKNJmmMbCxQ++rIGKDpDjFFm9Ak3Ecqmlehibtir9q5+GKCtYH7pPau0XyhBrW7U61BT3+ybPpl
62iVwmg9Nj4g2Yp8nMr/FhhfIB+xx/H9w8A/AhqCqEnjbXAN2kDhu+52ozBsBayo7AEmqQ7DeG8K
dgAAUcIGI/1xXW04RIxZpwXKxQZdu+YmdYPpr6tMTnCBz4RYtkamOIdzJK6b7pF2OSZEjXJ5pt2G
w5RbmxzE5PaPqF21dQNWLcOeA1VI4NM4KdcSWsair9HfdUgS2/zSVw06bJ/klH/ONBnD2Op4ioim
rWE3DhXs97lELD2osE6vlwMBDqVWIbKNJ6yOIoR16ztevxt4VyyqKt+yLRn8cCJa2yydpudz/jjw
tlNFDb4gseln0J/Ftm/CD7L3Wij9G6NOrnAXdbu1JQvHT99dhlJmI0Vb16v7i8xpHFAfE+P8YnAS
AAbSWrqXH6lBhzDK/zC19rChg3ovZiVU7E0qb8QkPWBqWo77OnzcA2QHpEa/dcc6FpKr6SW4MGVK
C1Pt+2mFa35q6gc2dOnaFJz+GedVcDNFSuQ4bciBExbnQS7b7EEyKwemqU0HsrjhnlQrY2O22qUQ
hjdV5gwDbM0wVtX00ME81TYQVjF6fwzQmqW1Fxh8LEnh+PtsKH7Nl5axWzXf2RkdiX8odxNp5cqt
WbNcARnjipT8UUyUnGMy9WL4lIxMBGV7+NqIckOwWnXnzQOCCkTOIuw6qe+I7+orfuoHMPFe/rxv
N5thki7/ORhgF0zKszWprrmuvKDm/jdQ57gG2b54v/vcxCy7xvi+q2hyhArPK2gG44ojJQe1yg1Q
hSNr3VN814o95W9umkJph7XlthCblD8IIf5Qu5kIueTn1fPiJGBRzjeXSUlrrGHMAEbc15hcp65H
h11uSb+VuvqxNfyMOPMdQBURr594H/BL9xLfr6hpUFbKRyqOdrxmsAx35ce5b0eGvp50tlzMoft5
gaGT/py1pyz8+otdecmtjuctnYrtam8AZC48kI0BmWY0oseLv9c++LU40v3yhceXj1/+U+pfAyeJ
m6ts2vlYUkH3yxC4nbgOTWB028pNeHk/h1Pfdyt89gZ06RTSHfqb/0VohK+5qUV9JcPgfTzB9okY
600G2zABzAX5Pd8q6SA8yK7rZTXw9nAYgFFcMDjbq9y3QcIaOjLbEsDdLSxB7gBskvB0tatBOv1h
vPJo2hoKeYc00+ApZ1p2fcgWlzOxgTOk/J+1akuKYeWC+B4SkwT0VpldxV+fvzUtD4XbQSi39oZL
fm09bqPF0sIhcMxnpD8sEc6DfRnSIqn/ajM0Dy6mSSsmsPRiNxx6wfTBidOmuMJtGa4C4Zc+CuOl
FNYlzDaiDFeYYVeiBFJ1R9bZYsRxgQbii3X6Pareeh+WynOAzmd+JeGTyF6BAzh1+N2XOqZbXunW
N8+gfUYg5VtGtLRoZ+4R6ty0F+KmzH56AARkN3ufQviepkdJg4FimSQZVSzId98rGx65xcUP9Oa7
MXizCw30R7gN/0uV9PD+Tncae8zauc8v4f1Un5Ym2/tG+eogf1cfci9HGXVMZnOmLGmK1XBqIm1L
yLNthGgksvIOSF6KdrDhIeF0+ZK2J2+86eJrjjqiMQNiBHYfyz4Gx2qfPd9QNqLVcGdyjNWU098P
5hnz7+DMNHhiVaoA+b3RTHSOkS+aMNvOGJgnSauMh/WFSdnf3vNobxolV5qp4SAexYloSITY8hyO
eEoyRozeW5M31FdQ5jgvl+9HOKmyzzse4EY2cntr9HeJjmnSqEGCQbdPm82ihkzCQaQwb8nfU4JV
8F8giqrBh0aZxAYvyUS7EkLkvTmOrLT1lnFfbjtF7fMd811pOuaC974i8M3cj5ig8gX275QdcUJB
sOJEQ4VBEO9vuaGZrzKjyq3exKbVGq611locNmtNyYoRuT0IcrMOa/1PEdVZQvF0lp6lPCwsCntT
1WLHgRgnx4iKHfQt2/nzL2Z+kNc+50XCiJ7gt0x5HaBq4YnNhApyrEoNVBsbA7CnDA8122qGnhAT
5OFK+vdyBts/IYnHHVeXULZ4NHmHrhqgTmkQkqEjTdp+NZUihEdVgkakm9Y05GWqtbmnPsdzjFWO
1o6oIdNIuf36e9X083uEjnxmbi80ezOM72dGKMaaX65XtH+GAMhYAXAx76cZA083EI1jkclNJNij
dvR+rVzxZZPuzYCEOXaSW141Gq2yn1F5Vov9Iagc7vkX1jdlHviJ9q8LiN22YEnRl/OdZiC0po3i
QaOtc/S7GrnuQOQeXd1EWNGbWooumnOE5R6I449tOofUi+vSjXz9eTEU3gVkezYcYVBKTRePfoBi
p5bzeTCQO8OSIbs2E/H/cnUY9na4DzD5g1wSc52pqb6lVBwEAU/5LNROgj1PnnsfRh0bSY+hGLnm
z2jaGSuqucw4rv05OxH2dyShuieguMlil9B6FiDEaeQ/YMHYMlIVehqpw4uzNNviTzrJPJa1AGN8
bOrNUQ+pFHzJCOjiGymm3BGT/gw9VwlUfNdRgWzJOMAg07aCZup41JbCxQJyyyK+bonMWm3vj1Kj
6xRzgsz/YLBpYXngDrNuT093xErHLTAAv+WEGvoBuDW5d6pfWnwUsAMUy1actwPvdeYFk6lQcaxe
Ei70xrqnZiwpHxeA+1zKGgV+oRhyrit9p0/A4l6C658GPEmAETwd8euyGztudyznkaRflbtxrvb0
6bfxK2PlDNIEIi+D+4iouWA3b5OadO3TuZwCEHwnlVviSAoIqXmCy09OZKh0oqKQNAj6RZW+ykvo
C+vKG9SgddmJOCY2OJpGzJQLh4xd+zT+8wnuq3+GVkdEcyaEo4H6ZImDLbrzosNoNc60Mz5nf+3o
pXO5A2i8ym5c+d0YylEw6jCDfDotncDDhPrjSBCiQgVrj3AwPVesjIsbrXecLcZLUwj46p6U703l
VULybsVBint404W1J8keUJVpiSkV9nTYmrUBarxUOIuSegI7YgBxOYgJjAPzr99H6YSQpjS32EVQ
pLNIKf8/EywV3xtgzOsbOETWV8VSToAIzj98Z3wHlenXNeuFmVpch4puTlslNhXTXc84NwiOBdGL
ygRB0Ffa9O9/EK9FAuRtpThd05+GWohXQ31RmAwRL2PBJTNHqskn7GyJVTq/ovMttLE/orrPMpZf
OBvTpMHja4nOPBHNKUDNpFonoOW2gcf5cKnu3OSHDBYP7SAdqe0mNJIN5QJ71oo4Ab6nIBftqOd8
PUTpJQ5dyCfIE/mizSGeGN8AsCz1lojsJUXg+yffK6Iz56Jl+l7Tqn67aoxsSxaumjvBILeUZV8B
pIsfYaIoVYvaxlfIT18Dwqyr7Rrc3q/LqVQGG6fmQ16UfzYS834mSoNtS+lCHUVoEK5rfsGYxkPC
A78nLkjW5nlCIjy5MoUHUeWCdg/o+/zd+a6AURpvZjKTGo1UNI0jQ5IUs+833U2DHiwtvHFIDWM+
wUbpUMSRiv67bD5UBemwESfgYXJiZ2lRtM0NRSRx13xtdD7d2dPTVjjlc692HcXw7VIjWHH5HH4F
RoVZO2htzOYjVqBpIGGOXO5HtxnetB2ne9Mm5vutjJwuGJva9uYhlseDuyZHCGR9c1qEwBLwLJTR
6EqN7wLkUWFWP4gRxs2t5A7YZWORVW8wsjQ0gWskNQV/YjJTzK8sXjB89MRSsjHgxy1XINkzxQ2U
CHISX7Ut9UDydFaAB9/CYPnlLDOMukQ8ZOUWaBiu6NjVIRIpEdm0QLpBnwfCSzNGXrt/c9FnTaYY
QvPRLQNi3gZZjT95nZtEfxEZnpwgvOgLDDRHsXJrhlVW4RTG9dujt/FCvUSBGUaqdRRJQvEXjSiA
N3B5uVg9fvwkKW61itF+ZaXDcWtX/Mz0lFFWuQJf940F3RTN7NgZW8aLCz8xZVgyOfi3kwyUXs1A
9qCE4+1lY672PSYIq+8JlvajslVHDD+TLf1lwIsqVDDhT3vMlVzow6aZF2Gv3zLk+xTpRgVi5lBr
KWp2LaS7WqJJmiY3CGzfhG7VS/OIyfwgJokbsOPJtzwnpDkm+g8aSSwjMIqGXg3pQyq+KIdDz+AQ
WrxP+qUQ8U6/Yj2UVE7g1loSJUIQSZsTIAWD0qVYMAaQisk0ul5eoaJq3x0xW8jDudmf6zUzIC0H
ugifbK8gDC2+LHiRNMPSScLiZGL8cqhswnXb9UpOCW613dm0EZg8TNftC1lK14BTuRmpj1DULZAP
dMsNApn412FbfshqRCFDtUVxh9BjuinqqrogYkLg4oQXsmYQ71ngMT9ZwXgZXFXr+ljUoAOkLYn5
y8sOJait22Rc2xO48+k3/k5Lj5qU88JmmkrUf39zdj5/RpSqMCIMXdR3Uk3X/Rxm+jgsaQwaK0n0
X+aXLNID2y4YhhPTkNXrFTBIiw4GEPb6fDI2ffWBAHyc4yFjtTj1Y0jaj+njhAmMZkrckBz9mzcf
uaAY36fe9hj0vhgyFGMuffktL9bFzWFnpoK8OPQ7l6lURZ9KqEihseLBuhFc8zNyfEq24UgXN65V
w3Ena8ijhsDO1N2n0NAFm6XGDJ9JrGLGOpl8hlftKfD3Xlic6uyoPuwhkK9KunepS7SI6sdt3J6W
7QPZpWsl5Yvj8yFer5litNcozgQjHwKudu2qWrpT2QGBqRS3E53/YZdB9RbMaU+aV/FDfFlt5ShR
KXaYt6e/jLxaMqk8Ov0KP5HwItMkXSan480asczL3bOeFUxT7mNS7XiLTRa5Pis+If2UJThS+YtY
Hvm2htXOuTTqkZNRjv1RTmWLHsozEWUQc57CQfJtAG0esv7s7D++dZdwa6IYEJZnoptpXgZZmrEr
EaCzaxd3oMioAzl68DwD0b3boNBYX1xekLhYT5RGUCd0FLW70FSnfMZGEmWnpt1OhalQp7y0zWzq
8R5GKOAw+9x7AzcVS8u0ZPQ8rMHLJ8IG0UO3RWmUO64YIaQ5hQ/nvhEuiqhGjktl/70YcMstnIBJ
R9oG+g1dxNETJtAwttW3t1dolyz1QjiPTuRL5VBXH/qNwJ0ZzeJikX7SoLJ/fe6kY4IECOrdEzIg
LvYSJbeejQ64+skscin1qyNWyZacDQqjJptowtSW99/ckIQwdx6FU+/DFY/41z6It4wnxZg3GBbB
O76x+zRoEF7GS4vMhdZeyUdIIFB8aZc8vhfN84qKBwLNUwiJSoB1FEnPMDmjH2xQS/jkU1b43fVc
KVZCfCtX9l3OqCMd9bk0JeDuoAKBxajvI9Bw7PxnxSoXW/1JeYkjLdNmnYUOhGOM7aiznvJJuPgq
1fUI+MDatk7sar0XFiR8EXPtaepAGimznWu+VMafEij7NGZzRwprJSyeAyG8CDJ1Daq/vLG6r0kh
TEht4hoeDbg6wBfnsovzsqiGOOMgvIMifoFkW1Q7Jb5rhuwq7YO4iD5is/IhS96OO7UsN6OwVfC2
nlFUlTDyz2mqmmhgYUT8+0FWsQyTs7IE35IA5Ss37ck+zcA8qk6tDZDq0IoooXZxZCamofJsIOGa
a+axZMlwSY+d28PDKqS/wyUY2t7/u+wO3rugaTiMHPI9F6bWInlbi4WmR8okLprj3VVyHrzAFyXL
mbU15Q/Ik8hSleoxhXHWr0RNihXNyuTj99G4MrTkXHH2g4esoL2FEtQIdPZ5gJkacsNpyyLNudb0
D5FmYl+3H6ZKto9HumHbHg82c8+t5iouakzWbeLCfcNnyWCE6mFbIgDLDWaBTjch3erd8uiJZkwR
cb2Ir5AaKrE3zTWG//UF7C/n3kFdAuwwQESi7yiG28PkXN/Hv+KFW/Rsnftf/fC64as4KQ2wXH0K
+JN2lm614VZ/u4Z30sVlIKMXv2ri5kSOUalN9UL2APFxVjeAeNiDHtrv3Oqgjhc9ffLaGJa0MRFr
cePZn/hEjSbK9sCSM+64eO1owPP7HzF/xXVlJHMl4lLcaKwywZsZSTKOYgbt7RF9Cb8tKoHY/Prp
SARQ75eAD9nEKvPSftz6yh3saRy3i8cZSURIgt0oU1hw+lOeDk/9VDi0YZfNl0s7z+xeQ5vT1+Be
GTT/fLOyPhzIHcKzUhYkSwZ1I4Gurj/EdbMqi1XdGjE5GtItX7Ua8J8Ye+MqgoSfVTSRatYwPT41
oX/p4bzBmGX6apw+3JpOIb2xf7bkXxagnBCim6HBxKdbMU//cpzKLXooTTD57eNFPi874ZIseLB3
TU2w81jydk9Hb1lhBLNWj70IZfLDDOhq6DBoFtO7Xb4ZKDyqohUpbkloHDgeGuG1kfU3/oC3MgwJ
DjtnLnZUwhDVYZo4uBzL1lt89fW+Fkv4aNbXVFUe4N6GlhMr8NXzH+NdlHAVuG6E8C1zONtJlsf1
rBKB7SmMLVFd/e45IiBeZ6NHNy39oTLyx0SSIk8M2ra7rVOcxD6rnVRemWd5UjpOVvzDSD8LTFgV
kkvIzOqhiMOwwwoI+DWIy0alkFMZI9FkuNUEH88pItxa4NHacq3oM5R7ALsvydM46aeZW6sgToYT
J3nTWpmGFEjwV6IhV70jjhH8KcKBqa0DldLo6qUjFDoeduRr882xAFuhHPPL45QDtwVrmPq4HDR/
Db/hwxaZlQKZZySRmw6KwDSy9BFmiervz0CYGtrcMuTvcEAjPvB7KN3DMaRL/jcdDv+2hHjVEohE
jxvazSU7/eCuWcuRTc5nmXmlxf2L+S4jRaxtn0YCPY5I7dFTeQ3zOvuwT/x4LZYFcNmfjuDrZ1UW
s2j3eGNxg2EmepQhGXFDD4PVRjn5l+RVyfNlNERgj30PBJBVLpIR5DDe+Q3dj0oWznlGCdJQ/a0S
hA4pPA/LMBPeCA29TCwKLj46EsBN0gcAC5M1Dl0XcEbkwI+8pmShkMD7XiN/TZ9y40wF5wVWqgv5
rnnoxhTtMmC5d2hYcghI2mbrFQblnlHtBljv4vpQMX6n2CVmsMvi+iGa9CVezGVqXC7WrJ25A/OU
TCkHOwPDcKl2jnlguxc5ABCg1kZIH0v8NN/lvrYsykX/vF7TFDN5M2MG0LN56Sz4aQb/zFcrLt3F
XHcS6Ydg/0vFrkhejK1kCXmOeq2Z4bUj1S8YN8/UIY5NgHL64danBTHaost0z0ELXE0Qg2lAV9zH
IAhxkcIBWMX6bH/6VHU6rCF42tlfkCjOTX3Q5mmERyHghOjlZ5VcrPwsyf11oeHxVAH+6tMifaDV
bfTEAP5GKIKqAFhATItLx1AB23tT9rCXAXnYzkXmmiQJBkYEekt4S28vPaLPFr55ZtUOFWQ9IMBW
zjUm+ImztgtDtDwiavku3v0+4ck++EfujV4HH1PlVCB+jvGb4LcHGJXR9FEUu4lqUJDnp3MElQBO
dJP7ajaS3DNfe5jkh4ruDx6lRhG8f+Pb+dN+5MBKYnirN827uiBcGC2m7+Rb2r3Q0BrK/dGC19yZ
G1W5/a4CbVZn5Q38gGEkU/BfCaCTTvCVeq5wjTI1tS3yTCNbeVl/NFRt6nns51ltGR0PakmbS2xZ
F4YsgercL4WnLklYX/Ej1Jm0/2ADc6ZKaC3fi6K3qWpBP8qs75R+G0OzWEaW77usr+JiAt/UElbE
d/h11PvkZcIfPYahS9I6pcLrrtnMzIlXR9ZVz2+vJzZdG5NpdDY0lDuhsulMaVWIitdYsKF2JBsx
V3hBGqe1g0vt8pEihqV/p7cNhlzyrmu1niCgNfEEt7I6jdvtVhjCVf0wzufF36SEK0oXX33BuZpf
5M0yB6ERxeLQltdp7iIAF503xhpy0GJ/sJeOID9Ec3TFWc2jrwzQ+W3D8ItKI2OfxQg/Vu/O5r0c
iD547wVcS9KDD0GH1UPaN4rzEUJcRynP13FYzz+5d8EjaU7lk74xj8g9uWyW/HS+Je6qy1g+nyhq
OdfCLnrGYeap1jseMRe4cUO8AKiZeoFTpEG856Skbhai3WCeq85Ali+IMOy+paTXBvlFYMvcVaMp
kxesfIIukJEaxFOM7YgykxiW3+aPOimgEPYu09lwAom/yX+11lm4ZPwg0zLk0D4Mwd6hHE9NOxRN
jTdEQLqAYhPauqsxaGiOijzGt+2l7LJRZ6VNQWj6okKjF9En2xyGtk4Z6Gb0oGzW8gX41+mxZ5l/
TfdfJsXsksISvMTpiFRdFQKU8Fa+Z/t0B9fKNL6aLUTGUpJg7X4gqYJ6ilI/h5Ck7EsFxZdEbN3q
e8/g1h2W7EMnrTf6a9IP7ToLNzxCOa7Gr3ElXZZ8gHfwQULp84Bz7uBE1KVk4xhehaq5QIewEwPy
FNaL9sr9OT/lZiUxuKP5bsPaUwOSnSUl7WsbkI+qpylBAreleBbb77eE8OMeSow/fjfxdsb60YaM
OCdkAHj2x2kaTOlTUZrm7xqmHmBTDtQT0nWKuihqTtmsl+Wyl7edrm/aGVo32ldb/0kdnGirOD8Q
sPx1jofahc1Dge2HjIJSBhDPPrGoyQV7E+cP7CjUG0IvBgaZ0NS0BP+DxG3mYrMblJA9xBe6N+js
8R3JvzW2gbSRAndj9s7k4MUt16GO0g0O6y3ITCKArx4C3hFg6Czw6k5s9Kmk72oDf16mypbCGRrs
MqmTplJXGQWqz//XkReQ/kiPGCir6bMjMxV27ZTi7ey/3/cfZEFGj3UrFkqo0umRUFT7YgUzoYf3
380Wlf91Om9Ir8N+4E8uQIinVHNS2+Urx9/5N28cCoG1R1jBsaBhURw7Po66t2PGjCjjaDlyFaxK
yp3dS2RNy4g3YJ5HW0H5Je9xGqWLTo1Lh7bJTgVEcvo4ilMt6ROx3ksQOzkUTzHnKAiaxWAb238y
FdnpuFOIcAVzzL/aER0kgShtht59xKDemz/H4nF0iSHW/SVRzFjO5RC9UyJPvalPLVs6f3RiRKZj
Hut3UZS9hyhvvczE6Mxw+iFJIRlyvoJgD/W+QglI31R3ad2bB8fsePtxOW88fq2LwFbDWoSHV0Mk
uTl0g7kV6RsUpwIbJQnP5sAQO05GrWRXT45PoD161ta4Xh/Oon8iVBIfVB79pHZ4+zevkokJmwy6
dkpfAdHgaIGGWNFPT2Qnnn8Ugy6j+B7a2rZTBcEDd9Svt4Yu9RzkF5W71tuBW9Mh3JTmAQoPogw1
eUHbxFMH0ssf/CKWyTB1gXoD433SnH9iUDBxaq48a19yoRecmVoOB3XY9zbu8LTdA0FzkZo0Q+lZ
ZnJKXD3TfCaJQcusHlc5RStRx5MUMd0ImNobGBjPOCxj7MW5BnQOcJtOF0uAyqR7Z6mbmB7IOJfb
RRQlNOhoMY5kVxqlUErXftgOyrENfIqJpRrAqgPbvSZM/QUz+t4kUEA4D8F5sws6rQO3YahWBuoi
tFC3V37OuLl0grGnfteN0itB1Az9fSxCfxphoRK2wmweqKwrYFP9H66urtWEavwmxIo/VrAVG+s6
SwTgALuXEuASAbZ3fvHyssKxgbl7nwQjX6Zvzf+1gKgnmSrrCuWTj2KZJNR4Kdc2a9cMqW9mxZnk
VJz6ewGxatc244ddXdlRLhzZ9K/8Fecn9EHYL1k4WzYtI+YlfFs026WnAq3eKyEUXSIDMmYK4mQx
CQqlwiu/fp/sUJBbZ1jnFUN/1py3BmYcq1vgqb6JS9Ax2DX5dQ7Wo7lEM72QyqX1rxaQzE6l3z7h
B+6be62pAe23Rmi4JRbpr0lDpabArrezhrbElY+nfokEJI0mSxpgik4dR2dQEi5tS/lb1jL+wbZr
w9M/xBRDs462E6HIH2Hpk4WOLIZjbvLC5IA2Us5tcA8DEqzm5/HfCC8SowgQgaOMp3qGtif6EiiM
8LT6M5xBGlSoKkPtktD2OvqHW2YPj1k7oKjYWf0rv/CfRJw8MT9jV1m9Yp5nRClus+aqgKydVYNS
71HGnrkbt2tdt32lns24NsrDX3ZOcmxvBQMO08XjodB4aGiWhQefXbl6lD7NwbC0c9ve77fiA6cJ
nqlrUOQBP4aUrhYLJf9At0/Py4JQqON7plxMHeM7jcHlbE+x3w/LvjBhcJ2s8AR+oylt42Yj41e5
hT8fVA/Z4ebWAG5X+PygI/VpKqw3wBH8C7Pym4mtIOSNiFSS06pND5l+pSht6uXcvuzWgucLrXxN
i3BTKGExRIsTIXAka7SYG4+FDL66gs9YPAmH4oeQKFQfswZsAmQDQN0jtM/nTh1kkzt9PuV7Apis
op00SjmCzH/8Jrq6c/VfLxUYYUWLeDWmCLsBplGZ+RUkyCDJ0Af/jB0YI+cobMzPiEy5/7WgJU2H
5TaK5bnfaM3tFsS1Wf8BIxCAj07/vHYM5UPwNTKfsdrst3oNyqoN9kcDNjr+T6Ud0H+D8XzldKzR
3r8+S3yf7QWc3vA+nnBvZwIUjl56MzsSH2YNgczWxkd1uReiIxNmSOgIVA4IdlHEJihurvHpY0rw
WHsb2p1LE6R7hAOWuFDJbBM73kw11x+DwBwB5oIgW+uuF5IbPSLAzpGv2+/1z6xLNhkykL4N6dCe
vMIvrN3LzxIckmvkyA1Vs4rcAGt8yWh9HbNzGDDTKfev7pqH2ihnMYKRaZn8O26lEoD4fXkhQ6Ie
/j3bMDH+1D3IrxUNG5vnbsip6EKKcjdFmP8SA+P3F+BZOGPJwp+eYnN1Tqk8QikSOJmbxq52IvyC
B53cU5+XyRvKRmAd9slxJokocGHY6azxcpyQQf1bQjHTzketg0FwDmsjihRvO+1SN8VX1FbYJXCT
2bMOPeCIC8KBAGnXbL87jG3q0kYBUNzZcZ54F8wkWlTYI+7y1V3IvmRShuIuPfzvjVSm1mqwFukG
6K8gxfwmnWbMNfEsWqMDItHD3aXwhE8QfgjS5YBOjJX4gKAsCsvbqGSJU6rYMoBcLxbzPHeOU185
E/zcPGiCzDmYq2/aaUnFSCkAFCcCBjfGH1nyiLYML0kqF1YPtLx5BZnV6o9UPcok9ulOsf3jWBrz
At5dJdkQYCnQuvcOZwPmkQzJiVBMmF3ERMFa/Nc7zSGyaeddjTMhUdFLwMo16tnxdCWvc502A7wF
OdRRy1MbkTW/AM538WXpOxFrgCGT5FSepDDISkS/58SdJ6y5B8cmz/z2/XzyiJ9gC/+IcutmcAO8
yzt4sFofOOM/dtPMG1bIRIU2bkGp8pQFoSHdfvzgdT6kVUixf9vpZEULTNUa1fw0J/jQtCFErojD
L/mBow5UYbnqihwZEQygrAZwqk9Zo1fOeWfilIQB3gcnxd00yQUS7HBEC/SjeaVaCnACQQYNYbg2
eT/jPnyYnjHD4vFz9iubcKu8niof72laUftIlCCJexejfdXilRn8OSEDbnzQPVDxoATXPnoknVcl
WnMlUV/8qe8D/+3rCS6bI4BwYSPnC6LvaZ3dmf5k2q0f5ZDNB7iHmxw51XnJvr1SPWFNVj/ESERT
F8e7cOaZJcbup8V6GE/o5a3EfHiDO9IFXJhpb27KTzISGln1Y/9v9DDGkGN7Vnz6eZJ07lMKpQFv
DK3MVbOnCfAkmo+D6cLjj61nPdU92nAvU+ueuBvm/1QE6QqlsqdqwjWE+vLU9r1lq94E4WKhFveF
APw0IFS4YJRSAcmlhtfgCIIq7RnhuxfERFZFJiP1qNx1z7RMdRGzLjCoz8diVaJzFkVoh+8Lh/mI
XfwESTqeTvHTSvH3uEF9D3p5X1OwRv5V38e0eL9josMgX462uAJXD8gZ/ljnq5xbmpZUJESdUmX+
a0lrejBGzT+Hs1d4LFY/MyCsl/4gsy0ZO+cr9A/6E0uasC/SDwu+A4aYR7fLBp7QwJDc3VEolJBG
NBhqwdmxDMSoUH6OE0wlppHf18FpNvuWuK3wGfKr2FR/s//fnzENjAtuhWrYBpbPFKs1fkM18zfN
MTMqkSXfrVvOUcLqsW3dYr4uUe9m7zzUg0OKgTiHzSUhhmGf/yypbgtg1C5zBwIYy8EccMu6h2cQ
y3piFfX/cOL/RWmGMZ6rUARw56FsxxQQVM5wP/09zbuFZuwFihROv1x2nQ9ve+qAILc5ZH7+ifFL
OoX1pONRTvKBt4PYgSh/1IJY6cNBmiyavCbs38jr5C4qmm/i01NnautfUHcBgtIifuazHJniqXtS
figJnO+Mzeye0XqkI/Sl9FnnIk5aI2wnEHDrSnwem5JCTCLi2K07wW6k9NDGxaAjwXzKyNOag//n
YlqQRFjq6rTv2pKo+zng0Nq1i9ousQcx3nhCzKwnVxKDCwQCA5lnuzu6RaBtq922IjlVhOmg4ivu
rsi3CV7o1diPqZmqcjRHRO0HQFCYQ/6Lu43uZCkTC8W0uKqVyGEq7rcEIQJRAD8zQwKTNY03iS61
fhKv47Lt+eFt8377uKTdRRpk/L71mHAL1nbf9EpvoY8D4RGVsGq+ioK9620aNo7kxcPJ0ahISBSN
K+WKfWRsKxNJ59ESFuJna0VQyM8jNoGYmkVibkw8oxOyADLNYs7HhUUsZzs9b/U8r0cWndTgKGYu
iAaPCLOdsYGQo0e+E3YF5aqpRpotavBuQBortuiQ3OqSK2yMVt8xjhIyduZWiaW7uhFSpSxYwu5O
ynsxDsW18+nwbPNVmi98dSINrr+OsP5DdH3gadI05fhtY6Cu++oLvCtKHA9cfYD0TI3bPVbcZqw6
1/jj37ZFGTkW3GkVNljlwVuJ7sl5eMGpXHGYb4cQ4ZvrWTKtvzHzhTk6lJz7mQ9qETgl0uGRxihW
ZTkw6DVN/bk2cmI9XA5HmL9A4m/FyJNtaCZUdyikW8arsH6nE5Z6TOnr88ADrcWTajA+YpduoTHN
4DJ5aJcmkQi2T8Uj6IRqLRE8gY4jpxHBtNMgxNO1HbN1fSWvOCOvYBG0TtT8hJ7/LxDmGKbP87jR
UlgSzsvUsF8O0HDo2pIllrxp4XywOkuT7FWf/rmZcGq/+2Z+Bpk13LNa010gW8RAPRVZHDH8K0Vr
/LQgCeDFpMsk5QFQTq+D6wEBSlI9j+5Qm426+/WDOxUbb9yIC6tmqGJsSwIf0H9uyJzN7nnLcoOp
ErNpxCngeh7RZ25kpvsE+sJgjF4O5ToVA9tU/6lSo+gb8xvYC5M3r9EyYRpwmygSW4Y8/xYeH1xB
2sAXro4oDamFqx2qsgdhDy/kMxhk1TQ+Yk/NPilR6APaFhOC9DzJmNWmLzp6EFWMLceBf6U9Trhb
Wyj9oXZy0DGzdD23iyLc41D25384ySb5L62a7RnBqb+qk/XTPHPvrokg6NGoArrs/4STXz0WXN+5
WjsIh6OGbAn7G64XJmY1jWn14+stIIyx7CnCxxqcYKAxqvqiJr/qKp8fI74J9590tfK67FQcDL21
NCC4ooOJDz0Ju9TWV/5iE1Nc8nDHe1clCkOJU/hEqAS7flCNu7T68KvE64qo7WKZKeJpYfgK4to0
vlFv/LoCdaY3mtE3+Kh6Hc4t1ZsrmrWaGLCyz9JvBymVHNwn2/7PTmBegtRtVdwEATOKSeTdEd22
z7QKq9QSSDG8BM7ti7W7vFpPu3thKDak/0XJy2pR/O7Hr/2BMKvFPbEB8iqIKGiFRWjfWN5Es04I
IY5vf/e1jORkHAJYMMmXtuxToZwr/1z7hUBkxRpRQi79MtnpxCL6uy/yRZVeL/2Wxll5qnwhnGFn
CtQvRjOHU0mkDVGtgF0b28jRAF2GWbUNFH+SXWC5dBdBjKxfy0gveyXVJB75ZTZ3QATNj9eOJm4a
FMRmBxi9af+PHlUDI1foJXra1IuVnjbQbs3nSm6145JdzSxPEWLhyOsKTI9FN5bsTtpgIMpfCqVo
TswtXd1Gx6STNTnlnZp4VSWsp7zESF1Fv9BOIsSFpYKiZrlspwLZvtJUAa3PYDq16NBQS5dLe6AH
o9MaHM/LA4RBTDouQTHC6cxYdd6G3d1SmatGJHWhRZwUSDeHCeVl4POeAXkotuXcYXWhjlaf6hhK
ihOhW10DFemlPxJDBzjZnsnUI5uVPIevA+x9+rG6jL463N64TdOaroxA0BQeJ6zKdRp/kMFOxDuE
fu1HuusdEazpwEORC/VPR7JdfZw3b5EzBG0N4l0m8HeHGCpbgQ/QwtSFb15wT8p6zAfaQGOaz827
WazK8HVnjGc++vT4f++Y+eNwvIHYwfEn3Xjd8XaqjyB4YQMyl8PPV0JCdZ1rvufSyOEzn0jxtoMm
zex4dkPzKO9kY2jjm2KXPTB3W5+775nOAcCgBOnv76yLu9dyd5TKMLsyKhAxyF41cuXExPsi1oCo
Si6Nhil+LTQyWF/2YrpiCUPkPwRYW8lYs+nWuH18tDoDuHlmjvIYiCHPoGzyYZxpQ9dVpqMQ+q3T
mJIKm01wHCDL0aViKVeacoMZh8jmAC7lf2L9iSTHNh87VtYTlhmIvl8KVsbffZaMU2MHL3eUJi3w
oqyBik8TZCNc4ashI6xiHjWJTPnf32UFaQgbj6RjleAwUhWkf9FYBYqb2JdWHe98zlH/cXW/3OmN
StN6TIakGZjXL8hFloLyzolEyD+jmmJ5f6Mq1PgnVGMWHgI2HHGFCvvY85gn3JJgov60Bv2DARRQ
giGoDt8FnAl+b4h6Y/w3jYegm9KHcwY7TvvTFKTV1knNzY6uXrpuYRUEHTc9FSkZMSg3Pxy/ryoo
h5hFqg2qHoijuYwnB8q/Te5L7H1cr+73PmjB8fpmCpRuGRzdn4gJ+6nOKh1OI155LHXD7MSdKrNM
xkIBiVbX/nTL1U0wO07HW5jaiIYsHfyRCvbXhkseYRLSJyfLVCQ+rpuTiwhWBTbecXbKnH6ItfLj
G+tvKqClOww5YMh2WEKZ6nvQF+cByF/mPnvRVmFkS+cuZYBMS1YuQ9zHAv4GJD68wQirCKTTabxc
8oWF8NsF/V/hbEfUWlXeM0sg73ItKXCY9YaqNV7cMlgENLm2vh54BkwEu/8P/6wojdruFQafT0f1
o+ntpv+AQWyRolzif1rrytSSVQuUwKQ1exNspHLsjCNEvv9VWxJXzLZEFGQR58VoX5IVUMHouw/f
AQUNYYS36mrXsGxMcGOIGR5IZ2zdxvzeTwauMJxXTwSCRxz7v9YbU4v7xLZLeuGhN0fKm/qbNPNz
VGPaUp9nbh+86dFBWPGRNKcj83/kgtNOkmTojoy87lUgfzdoSjMfdebZFv4H0B/XnpeY5uEwRJvZ
oWKNmXDtuojH9GOlskTLSLs/OTHxxtR0MZPoXnBAgZy3mBp3CdEQtAyn82khLQHspzR2RdiCanfo
cnto8WcreDHkFUg3jRqVvIzbiKtUrYNEq7QChUi9DrI5+3+CJH8y5gtrPxAtCwqMH3b0mtJiJ7Oi
LFRlgdK+h/pU24u8s+VJMmqzjl+9rRp9+iQJCtdD0FjNmpAQIHyR0EVwKYEte/LnHVXE1eNZSXrU
EUahpadrWCqPqvKKNMT7PR1UzSdAF02x0Kuwc099ad3okezsY+R5CW1i/vXHvz8e6EXHpWQuwmZ1
a4bF8Fg2JTc8Vd7k6OtirusziT74RtPYv87GCxYiZBw0nP+oyW42O3z3PA4syoXhKFU0VA3wrivQ
kQMgJjgZdpAPypZptHgx4eZ/kHjv8eTseL8VvoIpGtzmi1Fztd2iBMby0jBKYzyWWFTAj3WEwO3W
FNoDfRsygQ8Cb2mNHk1r/xYElEbHi+7eIG28qIJbBHA05QJOy1kuej+j+KdFjUBkagkLEpjvLM4H
UBcbSSohUvlSTIaxkT8diMAX3RUFKfWk9k69YOcSyToN/uLhbzpuFwAQEN+0OCM0lTIwQx31YgSa
WqKYJ3AjAvayB4ZYWqdPfAzo2TM2YiEGt0uU+vxAPeMun90YB0sGN46KAW5ZR30Ckbe4rDUtO4gq
y7gTtGbdvoCWvNChlQLk2xyiozE3/inVX10n8Y6yfq6pvp9lcyQ31VR8ZCNuIcLmbM+h42HAh7Wm
YjBEq7f1yMdWb17kt49LXPSbHp4xrg05w4xKrDdH+SYWFiHRnhwtCMFDpWo6ZfwxFRlyDHzZ2YGo
1se0UaUU+JXcieIt1vGWY2vrQvRXZPukAO39IqEKrTDM15T7/Muwe9IPjJjA5mI3NQ5fLAaq6O9n
Whf8SgYdHkZUOtTtEpgG5EQOgGo88Tl9hXqb9a8uQTpFl3PS9/1M1O+l5jkO3eK4FzurRJJo+qGd
9YzBj1bazfNAaEIzdO7krU6HKCNVVRkqLukqk6Lifb5DyaS14uPaGyd/Szj45nLqP5kGQzrfr3VE
qHZ/cmoq4SfmyZiukaALmDauG/RBvdCsxSlaXOr1QiMBc+vIsdVihlDRP6Qcj0G0nP55tHmUbn4V
qLNDvM5ndu1GADYqK7VT9CUy38QE+wMJ87I4Z3mHNN1mY8otUi7W2aNqO5Gi0WwzT8IJjzFXqwBR
rrdhYirizQ4OF5xqxeQNf2SZcAncEQDx3uU0sixuz28wF9RDlb8b/Bkyuj+PXYWdB96BujMChkRW
vIdziZn5kJFSJ1YE1Oc3W2468ydgrFgwkfDg3VCJc1yHan88KylQl7GnwiSXaCkruj2J0cFoXPv/
3UFJEDe2US8gfo+hr68MLv09dqxl8VdJBm6PfwsYv4lYibNq33scJocBozFIZ6+1UDB29wNou0r9
Q2jTL8xGVJntHLZRaNIYFe0sTT/de4+4ER/JzvQnejo+f0eBUqYwKVqKE19rXdAEjWtoxQUysD/M
OVFtG8c1mVfsqkDilg0278uzbzlsXNI6WviLQX4P2m+Pa5JtQlihsP4WOP7cIsFQq1rO9Bqahmzk
Svsyc+N7nIsjiTEDpm26N20pbIte+G07Yb37vgWR5Q0fs6bge1AqsEvshRa3gQ0yhptG2Qe9t29a
Ezr2oN4TWprmt2G6yQ+0QBMHFSSIrcsRobEA5aGrGMyt6/EE/6dp4idBvQ0FCEWK0JwjdFKGm2Ix
QR/vCdUKu50m6fqofJPJWPypmIx+Y0s7WJaRH0d3uyzBIlfbO1StoIFfcx2BYCCtOSekvMBfdR2R
gJqFgKJkkPd2RaUb1rPuXUSriKkicWkuGI3bJxJtFAESGD9Z578LVXLtnH2H6GBrO61/3F/UoOOG
Az9VCmL5EZHQ/JZQv2R9rkGDLHpTBCAgHGTWTobYXoe2WhknumGJoIUClfrY9D+WhE07/XNQ1LbA
Ro77JaRl0nz5vfbT3ciHjtSBAaaFV6xnPb3ojy80YrAu4uv89jse1jzBL4UNIvrUwlHkId03UCOr
wDKt5atcFhR3pD+hW5DP1XntNeN2AcLdNbSdFB5WCbVssLckTESXfg+VkpgiW7ucSnpIoYfRUseG
p8Fm+PbP2YC6QAORUDNc5IFXvDbxsqY5HP+XRAMfe0DnNBanUCrl8PcpVtSEDNnY3YnQKI4iX0GZ
tHAGRwDRVBI8tbkQYb+GQlfH5YDVNNyn3a0wS+PgKjgFMHWkh/EXLpvoRn2PYbecojJ+dyVi7LD+
HtQrjk6BpyOa5hDP/7+b+2bY2NX/GXQ1cvTWnIfmB/H7/BabAca83/UqtsuvMt10bTdLxwtrDlOx
lpRgXTsDKqqTAbWaj0kfBhTloh7CEYUDL5obmDDUsbrRzmOqeLRgEx4fyUzjBcgDvh8Qkrnz6mFL
oTUcpxqiQqto3g8mOJSGFlg596a44E3O3kqlViSdgb0Cl4nYTQd4b3vIiaUeRMghcmsdcfRi9xOc
5r6QEmPwMNAt3LkydJxrmUOJqtMBaBIvgLU0OEsk4cc7ZRLYLEPr9UnTXezI8I6HWpxliH7jODEf
2QnXE8rXR5uztggJ8XVuP+GoPIeXaM4rGOcbORola0ELzDmR5uOxCYm3sPZLNrg/7Mdasl47P62F
0Mrg4Y4cfG5m4oX/pVxYpEbvggpbgAPHa5sunBoobj3jqNZahrcd9dulLsjrhKgILLTIZf6oJf+K
xAuTQLyPvlbaW3klE4aMuvxc23P8eKS6H15hmuOeoAuTU2bpHA4uUniIFk4aXnFIQPUUuMx5YjPw
bsbZ1fWlWAJv04SglaIFY41IhB2ffhpPeSR71oiTPjC58LgSziv/8xJ5ekL9BomkoGF1s/bCBt6E
PLGvAQHk7UUuGpol+IA+LQkW7CnWaO07AXnzGAEC0PDljy1jwHZIqp45bwY9BdBZvCnsmCu1/XnL
5O17NPe+X5DJRSEOAV8STyKCoT4shQeTSEMTq7EECQeN29YCgFaXKXUiqcoksp3aOH8tfq/B421u
Bmh7cMnWUT05UsuENT35Nf7lzfnxKaBMLQY5rwhkx2BYElQM1svIg8XcC9F2VqZnnPBqYiV/6Yju
//WQr1ave0ZLHgxabYK+u924vBDiZgBuFO+1ljh3yfakwFPZ8+Uj5SjPAVZ55MfUHnEnO1WefhQT
2IPXwUKXCsubSZq09PTMYa7I9HmRgC/vkVTIMI76DvbbmPTP5hWcODZ75q5+O53iPquNSSC0ojOd
90y6XeOYD0kjljuDiFwxUzOoCjgj1UD5a7Y+B7y4Men+L499D74XMoCVrpn4kIHvu8OR7YJyZe0h
LHFOs+Ktrb0S3ux0XQME2yIfK8WLW4q79UzMQx9lLswqenoC/HtEWabO1nR1XTyq4eLp474GIeGr
6CseO2wD6RV7ug84D492nqbPbg6H2l3xDYRtarR8H76jgHs7hL82LvceWG/i2ZH0AXtElXmRZeQt
+XB5sk9hQ22+bsEO1hlD0MZym2n7ZlaL3ku7kJnKEIOHNT3sVi6znu6RYOfq8lOpUIynjyLitwht
Y1tb8mwYGNhKCQpSVnPYZcMZJtKXtHgt9Vh9PZDXw1a5oiAC9fzmThcTUHqzYqDNUZX9r87qeoSm
/L1LeZ756C2o3lojCfpCj/5EjOXR722qTm45CW+bsTtruJb00zWiN+UkZE7v5fLG+1vDegDoCIcM
iLXofzIeJK3qr5VP6AFsj1eVcIS7u7/EZ9UReWzPyDbdg45VjGohRwcrzDUsASBa3XTEt86b9H7L
73vRhJ6K2jeQLiZW15yPOQrvuixtULASJnTtNFXFQaklTzBqneqPrGHJAHgDEc6lSNRg3+J/a0x/
dUF1+xTir1wZ/3aLVqahMyTyR0uNfzAYr7HrGkt/ml7iOubxjoYgTL8j6n7mqdxD75RciHdr/Bc8
F1ZVp9izMi9CB5vHjQey6LDXjjq6QmU2mUuwyW5FW5QZIHja4nq6EM71MyWMR9NUXMnoUMzAv2tR
6A6ODHZ9Va7IJPlJsJQzSFb8nA+r/fqPkv3X4bIt92T4tgPqB06O7/4havmRF1JFTGWSGCoj12Xy
nUZVd8FJ+n0lLejNsTmfwH+JmvgvccD3wYmKcnGgCbBqpyacdheJXWqXCQmI7NhXgofTTXeECnZC
paxLdIY1GnEfVWUhJ27R0Xqv8s+w6sYDWSkigZiA70j+SRlnqTQ3Up29P6+f2u+5sBa9R71mhF3P
1fHTBNhZvTsnd5GY8uppHr0Ocabx9u2PvADM6yBUiQA+nEvHC+yxIQ4TWZ9ogKg+Xf08S2jMNyEP
skAfAs86whQ9V7fEuUJjk0tQEQJTcgWHQ/e9OcFPLqxE3qiZrbtbKlOCXo/N5gic+YhKTIJSBqV5
Ag7uaEbdyEhROPbAz3zWrZL10flmsYJFvYuH3SRdWiuM8hNefHdIa/E6HN5QJiL3PMUrT9PW981g
wFJi1TsPbVDuuoIIxRRWHQPkpDAKDK/TqRHZtUC5alfCOWr/jAHLtbZypKHt2V3f0tk+UfsCNukr
TVrqU5ag61cCzHvAhqiJ/m3y1o4+auOAmpAJ+/4+6VOY7UaNg0vvH4ylJgRJg2ADbuDO9HP580Q0
cBZeDwsrX6BFm2sMyJoYPbgnnlbNk1+qrFP3lROnstr7HoZhKuXG7qY80Y115GsEhHKvumI5Ic2H
BdPLwkgEbolSXxrhRiNsACmAksfpswfgLAT9yTphKeoZNrRGX3hC3MLHVsMvVL7JqsewcETaZiEu
y0+uL2OOYmFJdinv4JjvFdb08TSIaxShuRiw44GkMeDrnSZQA3E8ahNfF8tChws5BShDLZ1s/ZrZ
Tw6iJoAyAxLnYn/2rit93T2fgSNmadHd5V2Bi9Kl9UJBMVCBngXop888E7BEqtntVH66pB7+Sosm
Og1sRw6TKBMarsNeB2oJbMC6gGdPbM00w12AZ24AgxjjRa/8/cctnuw9nZ20CnK4Uu/2S2Kntwr+
fDzv2VlnPCFLBioHU7yvHqT00lJ1K6wpSkkIKX3XBqYUW8gcN+sXU7lYdnpUNN4LYYXCwqRkvdsP
y5RfAw/OjJoVmXESQx1o+kVHlGcwi10jE4bhm7QuHXGNgAeGbqhtLEpu+/0l0olaSk4smpeAoLBE
CPl1AjS0ADUoFKiI+WOoxxjdmsoLB6Q485VEwGk4EjuRzwKSYPoggbpg/ediCcf6K803XbzT85rK
bNA3FepPFtUlWEvwNZz46SPy39QvEmjobQJ2hebrCK7A010Vq69/wHMJtyPwVU8ioiXqrhR9lOE4
vEc5bcDwWcvcya9cDsE7Z4JsEHJw2t/zuPejn9YGO1rTY+GFzkDcrVgLIhJ17Q6MRyyp3FwIgsST
55jKViR2N8lGXGiMVYwadxgRcP9Cum/waRQoSasnuS07oV061LbeSROAJy/bd3pvvtc1HPVFDRXD
mXZa7R340JZq72C95QWVVebnY3hY99g82SPRvkhmiRPm+rYFK1SvwSILyUsbkI2PcQorp5GQD76x
4sKIS8shJ5vKqobFxn6Mf+CZVc4yNLxEb727RQhrbDD7nsmV43+icTv93cZbGwqj7OT2IuZFlCvC
Unle2iFjpRnyFG8xY73mg4UzLcV+GlyHB/FYo9qbN80saSNSndQ1Y5caCAmJeXsi3NVEVrbxILkq
+l8dY0+Jvp1w42ueG6ovbOamQyli5rqFAVdyTz9yWjHDgXePzE6x8iX2NOQLoeJwzligNeS9B6Ez
Ud0u5Cu0NIsVXd6x6elMJJ4g8puhx1ST/+D8FJ8oy2eNy5PAhd6Pixp420KoK3pqjdfz6qTNeEhV
wKhElhOktZxsHttXHrpT9Xeaz/SiNR6NhQ2TA1ZHTnwUqXsDOFiHOqBuVuXOvHDF93kvpq33TaPf
w1RTzQFPpsL1gPyn65IYIZNn7SrpAWwVMgGCVhFBy1zqulXgwJubgC5/x2GQOlkekWXiHTYjgijm
pOmN0HjDkpol85qBoRV6SfW0BBGxFm2RsG0wXPjNMt8J89rD4lfZy6IXWFTxwz39S8GZpwXynt87
OVDH1PJCruiruXvPr5CTYTOLAvQtbGTNwThT3qmHH0C0Hzj2a6PxALDTQ+lzt3oFdkgPIbF3VDAT
IZV3dCTzIy3PU3fGXQax7MFraCNGGFj4Ij42+XKecyVmsoS7cgbe/MBMpElTokSg7s9kEB+s84j7
Aa07H4KQwnPUjKlXNno0B/bPAR66hq6ppngMC0KvdG5b//R3bmn/xJXis34zWmTK3i44Xo6BGYPk
pyrBLMv1Y2wdL2jF7Z68NLmEytXF5Uw36ns2ZcqaOpCTKfETdXqFvBIT15g2qttEq1dTNLpq4MyW
RV7BY3Mjrw/83yhSiCZiwUDncryJvT7WCIr7gFraupX0jyU6BfGfUsLO0xox+bEaV8QqmzKMZ3fk
pcaQF4w7M2C0Eyg9HVF3qzfMdvDxvOOFwqhGWgVcWjPENh3jZW1fbUQ6hiJerObJxIU4B/c+sOLG
CiF/cX8a+vTZQXh4NsGWNLgfp5yzn6ZeeLwNswt8I7xE7oL1FEEkx0TisnbETaWN6r/gZuJ3AZcJ
3KWs/QuB7kNSqjJ+42mYGrDW3jjG3+kpN74V0IDMh1Kd4oEdAuguWfkyWz+INTT1+f4bvQSr1IjJ
uJvde24csVB8FB0uUhEwSCoozaP1QIpat8dcPkDtb/NwReSWHTG5V4U+kTduEDl5E6Bc7MAelwpF
w2FaNs1UIhXDYzZ8CJ062KXa7Q34ARLZf1AqmQBR6yo10juIz6YM/WgbXTvf0ZcCmyF3QWxcdXv5
0vIYE77h7hCkWWiVh2qRsDhOFDeGMWwZnimuTXSDUZNERpEJ9e4GfCJfwHjwfRXZuJsr7Jq4qZas
nHOKhMEbSEg1PAOS8aAmqKkUrqU9uLGEBFFvkSOd+KCmKloplfe258CY7heib+rJSYbkJOOvy3Qm
XWTybL1P8yCPx/nPJPLBJIqABBU5sE2Ofz7+jczZ+VxHd6FTs/ier4JLyWP8Zeja9MaV+L/1BI4H
Vz0HfY4pnsmxJXmsZqH7hfzAD4ktwdxvn4sAO8XQVK4iH1lP2R+lvd4BdiWjAlxYJlO63mpmRsjz
jJOMk8z2BI8tvfYGhaCmF+nUiUdaB5g4wy3i09R8Xoc018JSApnJog4S1HCrJMQ+FebrLbhjqzvk
N4XPc/suv4Ze3VMR8/TiE4dULAx0qHzbCogxdsC+twnfaFgCHhvaR0TnzTefB+KmxEqMFmqTaPDC
6BJUn9WBgkx9mdT94w/+2irXfLTMpU5000GLBtBcNgl/h/512NCZA9RGC4WDmSDMHuI2Z54ixfdg
2YnjSgHrGO53moDuQGzmtgqxFCHyVu8mYGeuH/WLTCn6xLqXqU6hx0JVnxZmQlEJaXjuTtsNZmji
QncE1wrcHMaJRJyqlPu/5wMYt+m4vx4tyCyiTuu2ThAeyfnNc/yPEHugqLskRkyQ5UO11QQShQBA
4vbC1N3KR7RkjEPZYa87lVqOMS5dZEtyFuZwf9ejmQAIh6z7Vf8OmoZAeEO1jiCPcvPDyjVh2Y0m
AnH0As2wDwwUFDffr0RESlbMa5Q4U+Eeo8K57R2uHOIAPxIY25WIxhgV3ZSAb9dSUORG0nvHvEby
VneluzW6bkj0sSOwvawnmeTF7c1ATz0tc/VxmWexqM7NCHeIZvMpgyO273wM6Otv7PWr/LHS8pUP
z/Idgb+0s2fU5oVUr6X18ejbMsN0e/agQWt4lFkDWu5IOi1Qd2uj5rGQy0RJasJ1w8IsH1MZTcsg
ceNhIKHnhd2tlnWWuVIR6VOdeFzTU4d+fWeVyxGCnq5WDJurYA5OnhcXi6Alap3VELdLjJB/cfyG
fJ4dmmwtNZwGoX9SaZaAFbBYJfkWH4h0pTvSleNCC/TpCyWK60gEBPFYu5ds2p9eWKs61oel1oZ5
/BlYcpvvA4GokNLKQAoYvH+JY83oN+N5uLY9JTKvjTRjrTz2oQzJes32KtE0678W1hnLSeVSCKSM
DWh0+agxXCGVxRJwIl9FAI298mKcZwQjBKCAHFyto8I4Mh4Df02J/8/j5zWumTXB5RxCwooLA57R
FLqIbvZEfMp7lTbtubKwBWazs0c0Sns9bFnEeemfXHeVJAZLlQVtCdbVsN41NkbFVPE1MTWGf7WQ
aqhT0J/+37uDABmLjbuWAAg9EHQlxWJ8OBNw8lYfO7OIEN75wjRPpNvkjkWWSfNkdkd8fmlKTCqn
jfRQAv2CpSScGB19ADJs1OQc6v76l2GA4E2G2LSD25jZhcJ5C4uHgKcLkaOKkBAtxjYfhVlVuWhb
+/FtDEhH7cembEsokPHc1TcJSlkuVOdGrNVdgk1D7qBLDD0gW+Ln4060jai4+Ho81F7KJgTmsYah
5srsPO+BWKR2R+Wi16qiCXgZqBai+4rJuu/8vPhcD2NyYKHV+z6G9/h35idUGu5YZxgEqhtrkLbR
64AhFE7E8ao4ZLKojS8trbUUDvArS5oxNyScQ99sR7eFHxojn7JJxJc3YdnA8bPbdp/0BQ+JnfGI
sVulp2anbAzDK+NMcXdrvZ/UB3Yun0w+zawMCDwGBkLOYMTKLG8YrKELLTSNNcMyQxMZ09ubckqz
V15X4aeF+9/EyZZmZp1EAB+pToqUniitRIonQeBM5vRzdgZo4cafda4yWH85GhlAc+N/lttXUTBR
ikl6LsHkpgKTi3YPhZajYFBoLrh6Pc2KGfIJ7FCZ/LBQlim7v05PTqi3dVhmCvcA7cU+dhMruBKs
wdGsSVBhDqzDHjwkFn/Cofq4z6ZHS1H+SEXpdTnPwA7QS7+3cZDLM9uGtNChTUkmjMY4+O8FdFyV
w49jGUu1gMhq3Xu36eGQGp+Ym+HKh32R36edMArJe75Aj6t3YwPqGXKAcS7koOe3T1X5uw1AA9m4
3x92LxGsjiO/uSYuPlUkZnanqy9dOL/PtRtalaWK1HC44OQiqkssmfYprtV9g3DIxXga59LcNqOE
L93xjdv8izC5H0RmL0fHg3v35yTA8ZVAvFdnKSX+1bZrAY0BoCYr7hE73ed/xU+xEufPuTlFtwt/
qRskkCUejnnKMno1uQKpOUGRoD6ITZWHkctznznB5OTauQzCWricpRnWP7iF+viIjyG1PmdZ9P68
iAZsfeSYo89mxGDES21+wvQpkV117v0X0sf3TMiZFVF/44AjsAPlvF6tsSFAZA/e8sANcg+1j4Z0
Jwz4XtP/gd8dVVGE4m/cg2cE2TnSaZ8BMX3QFcT9KuDYzUq54OCc8V+nZtQBXJw4uBySiIeG3gDi
YtBssm15YDDYEXP3i3DKkgQ1ryNnf1hNEC2qq0uzvj0GuNGg9AysfMMEvk9LFjpArQIhnqvZZa2m
YAIzpXmdT8/woTFr29+5gmvepoH4r7dqesrLOndV12PxISG1Xp6V5L6i+uQu4v/2Piw7wChd/Htk
LC1K07g7gGAGviiMa++3+xIVcQhvUhqO6ddcLsuGSqZ8nVk0smWir6P/byDzI2mWZWWomcf63iPT
a2DssZPoESBMGptif7q5JHOUUmeztp0drBuZ5y5DPaVmBXt5Qpq8ZJWC2HD4PBLi83uoVKLhrQej
2QgKDw4fGSMK5FbRpFz1qNmnmYc8iUKXWHBRJD7Cd0sf4C0mBMwDThI242uQVjXVItBBEtHzTLyX
cxsjYDRJvEeLvP+BNYeVimDc0q4tOWSfIgCCfCKW9o/FqWx3UtVaJVAKkAiRjziazIMqnzKZFUrV
ZyqstiyJFqZ/XYAEzqZhqKD5mzRSkWK6BnD8g+vDWDPduEqXY7Iaxl+YDSion/eKektbc8uQs3uP
nFiSulZHZD+F7+qLK3yE4TddsdhQXxbYIPiZmDn3/SLeZnLO63yRzUSFMsjbjKo7x3gWwaiht4U1
kniegnFpE+kZX0hyQl8tKDo1yZf9Ot5prkZrdxJKGPv3irxrNyL7M4TbY9YgMwqu7g/qDCmlZiF9
bTf5YO+r0JznFMjDDWNANVkNjICFC5l35RKOkHpW14zVo8PYWg3EpY1ZgnQShFGIYQsSvQCApc+u
9UaLQxiO5Zla2kjFC1QvnBADlBZzAohuLNXPXvLMqFflf9rK3hr6BZUcM8NjJmk3SuGx7rl6oZ1n
m6yZokWgAS3OXN+FzPN1lncRcO3B4iT0opCjcOBUCnT34kFilX85NwK8mi/ayVkABniu6wLteSsG
/HcfxKw4a7vgbns9xmEQL5Br0TN5qMqDd31SmFX+Hxqz7l/8pgu/ZLWv4LrNGzov/68CVRY0xM9L
tpbNUto6DcIM+5yuOjCjBbYD3aYLqWdaxWymIvxrM90zSs0seRurIYCv1C3IcFCcDn434ZYZMuA8
FD4lFP2dTRDZWF9bkbZNVeGQyVu9VmQCZfYylDRkRRLuAJIJSUZimc/t+W8uwiJmsY+05JeEwPHi
WcWUzLsAVnq4SlX2E2CC7KFId0Qh/NvxC+zNmdlDulcDIMop4ifFfqT+8zvV3tLtkH92zmLyXPyn
IqUv8YqMCyPJyiwqcr3urxI/dNj6tDfnxNr3D3aQKs8XR+DAHKCV+yNJTTEVqKtNaEdKFHdlI6nc
zRJgVAkTR9SXEqkQKQVA9YjPQkGhz7fn7kp/fXunk+VVWLwQDscHnHBo/vWlZj+87FX9zAM+pm1y
F1LRw+dU3TR4zCQFewb7nlCodL/ZEtkVFbMomeFRVGLAgMozhcLbqtB8tkszyPwpvU845xRjr2hM
qhrGlzHbEIhAfVus/JYGBhOVXhSzTFI+/kjgadyya+HuePZHzTQiXfef7uzorLP68tbiF7tslir4
+3pnzjuRt89rsypPcMNpTlliMHGaai1Jbt9qgqN8QAf1c8DNeQ42rBa0Ev5w4VB+1YCjdy65zU90
T6rWCViyBttTWv/fu4a9S8BRrny0FVcWzqdSnVNYV+TH1FO/OR8dR/B0xONA/kYECvhpAcuuEmYt
oOwVlnTbwmQoy2CiTLvtbXtv6mP05U4a0Kf6BPGir+XAc+ARKBn1jKSrvLoYwRWzc8MNyDcZUFyc
jpL/0ou1HjFmKqzwqoT+BAIzW2+07vHHY/rC17JcJjW7UcKUFEhqp2RYGSXtGmbY+3R4O2hqJYwN
UqZEhxrHt/1Kp9gz3W+zAXHZ2PrxEB6LirDwDu3w6OUP91hyjO4UJyv6E4kzI0OxpgmppZ16mBH+
NP/slOYl7zbTzJy8GEfQLtKcy38fu8fs/XFNp9HHu4JAC/r87GNe077iAVx7VaQ3i1b0IIhCPMwQ
5TE9VE2XJVPmpv7BDlNpShuQ48UhP2oB6yjCusFaWEAeQpxB9zIFXgWoT4tZZd5ltilY02eYVbiY
EB3NOvGPd2hleFGCMXuPRADa8aVHLRcatfs7rdHIUXhlfmWnX1Urgo03VAazEX8wR7ar1eQhmMeZ
LmRTjZYUYJ5mUJanRKxThhyOAgy1RJbQjhI2G1vRJNJUCABau78sqiieD17DCMRj/6WVjQa4mtq+
ztXsTSRyPfjFyZC2yodC4x4pghDtUVLUJkdZk/WeyqnWwTHdMYdszsic+L0Q4T651K7IWgX6H0Xn
gy6ulAJ+RmXqpYTZsKy1rkSA57lxDcgQDNaHbn9Ju31yasgxl25BORssjLLeDkJyVxhRcAEsq8Ac
N0Z3emVC1wc7Dv0LGjKsgosRinf95hc5DCnRRtW7StT0IRgjUzlkH07DOGJz1UtWQ9sDaB9Ryd6v
HIT2ZJalhTapQ246EdkEmTn/axxVU28Wf0HVQn8ylYrilt7qquEepNFBkpj7UqM61ypnjBw3Urfn
W6j7kAU2yIflgrji1cx7sdMy3IyEnZPkBoJ2vrCJL8EsmlzOKarB3zT6M86S8s/LeOYvA2AWEOVd
WNp5AWv2H+evi1bWGyqMbcyo2nG9pCUPvKbg9+EjY7XRo9mkyVdNY3fPNzLNVrFPwqBtvpOltxM4
AQofvdi8yDpNxxKu/o1tJe+GTGCkszDVCkLi1EOgkCf1O1nDYRchRZjrtl8Ov2RWAIlLpYjm9j8m
OxCyl6zS9PDp79hIuC3mLJXYTg+4YMQgCXCm+yWgJEOic13N8EQNPl/ebPnPlGaBKM0I6b4gCWPh
Wp+lX3JoFECkOpxfQlvqi7pIvEaPePcPhytdBIKo/uZ3vxeDlZizgVH/TiyIaKUiEeJhRW1PWjqb
tFPYuSHtbelHW6/v2U7VeB/+AgiSjdMSMjMXZahRnCBO6OaZHNs/jPhEau5CSdjCd3M0dPwpZfzW
mnJsVDphCYqXbX0hyEdmAHp4VFftUWm/jQPHI89ldnJRcR5TbpsXWWTuqmWOybndBJO2UzNZk3mS
MTioxWdKqCRp2wE5n35EZH1cEpNQ4wmt88CbQ88T3S4uJ3kYT1wW7k7/0ezJ3+Bjt7WGqCNv74fr
+ZarJyAGgUnNHRBTDdWeDJiAUupidVcVxKUSxM5S9IApUcpByhurzb6z+bxFb5wykn/H1GvQ/mQv
x7y3kNJ95vsm4EVgr0+tZjRkVMzlWh22Fdlt4IuYjCtIo3Gh2NVGSfzP2Ta5X1Vq3018pLXR38eZ
EZjqcxjab9/1pkXUxl221lFIvhHIRGp8Gs37A9sdeJ0pZUCUAtTRkHla7Xb9tz5Rd1jydUPxjwL7
qJaoGkNBOF2z0BOnnT0sAp+XR7qZljRTzQ9O8BkeyZ+CuV6QjlNrjSk4Vkc9tWD3ZWexM2AlzyyL
bt9Xsf7QSDBRJRlnrmEHVLl0BFMvGKAQBaxgZKVeoc9f8wVbUftORXoKH4G1XbJUecvnoA9BG8eY
Y/1U0Qwd6vzXLLBi8hzJSU/1eVcXsfUJgfeq15mA5pzx7IVJPN4S5A6adL3xpxWV16yFlb/hO+wS
LBs39hoY3ERD3rp+6cnZaznzKlmn3fdvYrqXNtEozju5WeAnllRZpZOT/42nOgg9sOMA/eE7PtOi
wcS1y5lP/RXkZq+2LXEPmtvAfsBRUqXGWTxt/Xh+wGMXp5K159x8GBB8xv+EdMEiDqHmeFDBe+ku
j3mPBzqk/MtoBD/AUBdvF/xy6NZG9USOUBb87kJG0at1O4tOPvDm+4xSN91eHRn/dbGVex+aFA/5
A9bhk7iXrsI7bSuYJTJH4sYQm8r3Dh53gJEiAQoTT/yT80h5tjLU8cNUVHD6crQNVeg48oxrkckE
zJtSJMVScKvR9Uk7FT12ZtVB18UNoFp/YrvPwaQ6uEBUKD1dOHo9ixXDIC9W8ld4qiWf4Hd2ctah
8GoEk6i3DqoEaCMqD8hRj41KM53CsCG0254leuRRwkkUvNARsVKPsYJgGY0Gkc3j8zzpD0M9HvUS
LZRCq/G1Qk7RkLMQIBI2Ri+n2UtPWVm3PAj0kor8E24BjkO6bj0d8G+LU1RidMLeQJISJDJZ5Aah
0bTznw4L5elzzobQuNdOcMNL9xiMsy+e9D+S+5ddm4qLPb0LkDyYxb9ZBwBwKvKPFwV0rAavR++h
RL1NEs3e0cjgCD7C8MjMiqGaJkO7AWldnMJXvFc7AOy/Hz70lyHfS2FCZxmLtGyzTl5po9mz7UwL
fjvVE68mEBqq8yYwXA6PFiv1OURzHNaZuSY59jnNJ2XhM0nWCQ2vA6CqdcqUvJjqcRvyjPFkGoxG
EiYM+SuS9Orvz1yeerT1rlhjFzVuvwbpiEP9pbqlABWRATRPQEO8c/9+WX9mXAdGllkjt+wF8VtY
Vc3hBYw+pyaktJYhW2VG3wc/CZx1HVzOLWeBgwhg21r6ndU/8t+8DWuboNrG0IlYrnnlIdXiD2vF
MMYPybi6duPODUKjq2k6swwKMx2SYnuvj1c9LVirXL98fSYllzxuSte0ojNcq7M5Q389U2kFW7HV
t+OSWgUM29H+1vtI9VL3kHYOy+8+zXDGeeEVEauW9MxFG2+tr51kYnYC3FDtHe09dfPmWqgeuGHP
BSBXzk8QQbMykcJ5BWoyrrLSDk2E+hOJx6cRRQigEr0W+fLtBTHHPM8DuhOjXnITq2zMLSFo7CSm
Sl+9nwKqpSaAZ8ZqEGXB26tKRQlsStSPl2n1ox3zmJr6Ix0k0hxxFE/Z3eci4zO5AnR4Kc01QPnQ
lWtdFYibHagyt8AYOYf+2e5VeY5wr+u9+nR7oj9pMPsTqYXlWj8OML01oOOiMCv3x6i9b4TQCJqY
W+iulLEsl8V5GEKwYleyT6Jv7sbHwov+Wwox/h9omABBka/ek8ydi+/PApo2rjmzrBWFN+5La5Gh
n26v9HMmvSjComvSdRclrtKbwzBCpCZjP9C5drrkk1hmwBFIUv3RIMbstNH4iSMoV9I4g4SUOLnY
FxrLc5NXNJ9Pgl9j+VW1PKK5PiiJkk7OWg31Xju5cbJNU8SdnbStyXdDwvF64cPh1hThGXtFsENV
OnTbyqGkrBAbTZrQtn5J153qvezdSNsTHKZq6jVTM4Rx4csSLKxVGhhtgp+68iqPDLewACqj6DfW
OsfMmaqXcdaDmp6yHf8/YTx1Ze7mWOQM/Tl+4a9sSfzogbRKBzCqzuNGaJnH2Vr37KLNVTHN5gJ6
EeYT8caR+E3xKt8NOOtnpPAuf4tbKG0EOlsshlmHeVbbXcPvBXc+NMI26DGVBl/bhgC/zr5CkfZh
EQ8LzmLKWAOn2ySt+Fu+nFihMbkc7+wvwY3vkWfiRPfxuLeRj4ZBdHZuTzti4ATCOmirVu8es6to
MT3ZLZxT0y2RcTTeVQocG4wsNQg4WyTRNY9zuanYyVKNHnDVIhrLB57MgYRUjRYHkwVgeRBg5s4m
VCInMbtjADRFNttAEBAOSYhkauBTNxIYplhMdJMqCO9iKMZe0oaFeeVIapqy3WXMbeu3OJRIDcL2
sr46Xj9hhGn6XxyZmI+HdVgf9dIxMrBaw7/jBiI6cLLRoeq6uSUXbPgKnZktey2Biuu17BAT/kj8
PqH15/fwsZPSMXKixHSivrSpBrisAkUNeiKxaQNc8sxcEsZDvgpvLB1z6QiOADsnqvuAsfowTsVi
0I6BBo9EmrCv1TrvotbI6CXKqK2hFovwPH/8okJik0Kgshz+S9oGcEQuWprQABz0NXt4Vk8fI7Er
6OJ8c+CUBgE5Gt7teej2uujIIexxp7HcJqLm5akbWru9dYZwpbRmQg3kSR03P4rmTHv8R+obGVYK
V2prM2UIu1Q8jCoyNq5NMI8oSj0/DTuw+XoGoNapwiM6Tq/p+gJgqek6UkyAog6U1c2+4bZ/ZVaa
nNdDR//+e+5oMmhvMO30AWrsA6w9bc5xQ2NYzsqUwO3VE0+DeyUtkIvYt/sWQqxEXqznxakcE9iY
w4kUvJwGYZ1uFquGRH67obnUiiSz+00bhkPRM1zA1SIxAEPwSGhkamp5GR8lTEp4Bl7tDsorOCIP
dO57p5L/iI7Z9zly7FjBjyERshQeGx0J3+JoLvzVW2smoS77ZJ6bYLAt+pM/2+avcvlSlrwL1knz
AnXXGL2+hfzo+M3IGB3AeVQfFkIX6OKNnrs9NhxTjRYlewFTvis+xxifBpr8zxhr/O/xzka9U7s/
tSG1BfgTU18l0FasdK/wXVe/H7YbtI2sDfpJZHc2XHs3bzTzTEzG4Tj/2gycRSTB0qqEqv52cK/Q
4Urso/I602N3uNu+cFqtec3PPNWYGSg1m0gJcMnxIsfzC1zYwbRAzo5wVDgFT0PKswqt9zlHYC33
e3NKJAxNm5yN7ao8ufUgscGx4a8N09dIaSofV+foHgVAzPllNxOvwOpaI3jNL5QogHC7Pxryj9kD
Ix09WRwDVwbx/jcbovyIbFlcgd5lW4OL/3gt4JoTeGJDMBu+hNa/jgSnDiMOYbsQFeOxIVjTgP2n
g8rEnUbNlvXqWo+wMNjb4PY/yIJuYusNQ0P7/xQNicT7/8fvcdmWdQxdTr3kARZzKPu/dQNWgHnN
NTjUjFsJEP6Tl+8L/HW4DONH22t8T+qlS5r/ql6XaSTWym2SxYTelm9u/U9sacHSGcbPe8UiUYAx
UGseexUL9xpi+JQSdCvDfnO9iEVnuwmn1iBsvN/oZtN4tumN39UXPNsAcbSYBSy1yE0C/7TNOpCf
aA0XyyF9Yi4H/bZFLJ/SvG01aHOkK9DtsOgWFB0Q/AjIxoRUIZb51vGnh6CVwaE2dZ9yiS2W2eK/
6nHo/If9M/L2B6q+e4tELBvKVHSk5YerVKqqLGDjFhoprspHcvlwFifH1GGkgQdbazbrrZW/yTfv
MBveYXmCKmjiz6m1ybYv/HZnqZkvxkezsrcUxoDtYgVeDOqFVSW7QWRPBJy53vuqg9rwIdcl4Fru
jIR4eCghWaLC8BHNbmkMyDCnvHr3bvP2FkYiHph2AFIJ1oV1F8w+ILImyPdGiymRJFMXZQpu3BWx
LB1MUd5saj8LxmbvYkxUE+GCaYVLUnHjZh1doE0OmmCw6HwE0NNBkB3eXfCnelBVm67G4/DVzfbu
hrYAyUao/ZhIDLwqTR3w+zbjuhT3zhqbxOdDOlkBMhN8vztHz3YB6jlxfBZbYeLN/+o1Ox+toJEB
DxG1goNSCYJV47bw9EX7WdRuTBNmXkHKpGD03azKubNLr+p3a9QRl1RDWJm1obG4TXmgHujmuXzK
9lVg0ePKa6NDbtCG/1NrVNATnPQw17Ql9mSGEImfYfv5XOHjgFp6R5M67itfQytdfOQ+3xQrED0q
BJWww2cTbMuis0UPHT6zP3ePnQ1lNQNvONz4B4zKY22Tc7wE4VXg1lSPZRM8x3AMhz00Dm0Ntq7M
YclZc/UPVEuzMX8TIWYxXZ+0l4GFgtErC3wt0EAYU2a49lcCDvOLycbs4V59aNVjAOtXvGNw4dww
XZ6OW38Ad1WRF1pyNWM88/dLeBa1r/X5zrOZvBEmHB2MlLoRGzcNMy+F3a1X9FQmglurzCmnULDn
Ys8+Pn0X8tJ5DgQXzbkfoxPXkCDUHtlwFX5F5xcd8z+pQFWgzIzLzJUNqFzXwj3it0F6/xdMCgsQ
Fz7GacU116SezHHbcceth9uYY5HCzwQm0vABqPGdYWmJ1yzJ2tZ+DlXDgQCnH1aBi5U6W0nvMiVK
Sx4yAEMy1aqUeHhbyB779vzLTeROQxpECZr+lFfUjH+wyfEQg25hK2c3ZfzVdLL4kThp2REuN0+C
SU81xRHDCXhmvpYJa+rtEzBTWwlxRdfHWyGexD593/wgcm8jIc2OYkoHYg4V8bO4Kgv8gf1L58wj
4H+Jx4r5YnimUa6sZqVmIAwv/+/73Cu8cjpy5/puCw1jP4T3Qg6AZ82MScFRugYU5NCaCJtgCjVZ
ROVxwVhssuSZxpyzNcYYEp7OXbA2ohUkfgtSpKxz41RmZ8IR6fIf0yKyOZs9i5DNFcdBnY3BYhc9
IMQ0XnS44iX07n06Ull3ZosxN8jO/ZkD70EWBH/GWw8YRhakXJI1egCJ9oF0b44gGmdaILh0QUHn
pvkRvXfnuL47b0npk3riBzr2HkWywCLJvdg2P/ZlzjzB+Kfe1kz9rVwA1q/C6SubxTr17clqdkLz
QsoQ3Ky9GRNY1Kd20xMft4Mn3oA+I6bz/8noN3akkiivLWAoHl05CU7jYLOhp8vLVyf2k4an9EE+
ZlzLTg57Jci2b/cvymhIrYrI36yLmjd08mK08/LaJjMwz15dDlVkMGX+aExUzME13elxUaNd1O/B
CtU0J0ehgPCtKnUWXx3NBXgEQ/nQzmUDDnmdB5R7C8sVrUPGYweVqcvWWIeBi3vxefAJ7zrDCSdy
m4PDOJzfEiZkluS0SmDug8dNWfGovAslGm8i1SABvPJJCj+2+U8k0tlteZsIHNTojn4kvg4jcYuT
jHwg54ZS/I7n5Zeno4oqaoudTNr8vcAkDeRxSPKcarXsHhkmRjVP7J+QzpIwq3XDXIhCGkDrYnd+
SD7TaY4awBvIV33rSL/XAmKG/BUf9orstQRostEbHPU/k106sz50p3YCUu8gCYDpShS1tg5qfVyG
O1a+PfkYCO6dLpNRZjklS6YSj9IeuhwHAorRIjPm+pHpID/JKe/IiookG7Me7Sq+WzD6PBrUFFI0
ONagSgGFF4YtwBsKevMF2+yZ19RD1ZE4Zc76g1jTjLaDzV9cOuziSKUGLoafMNELGveN3DErJ0hC
264HsMFcDC5rwTfk4lwZTKArJBUPfL6FBo8KYSjtgpGpxfGmQwxLQiYF5xAKAcqT2wwLqMBLN0jC
+ezr5n4ci81Fb4VZ7GHyuGsqdcHVRjgVo6VoGzAme3vaKUxPxdcU6YG7SJExLL2R4ZTw7pBMPkRQ
zH8yp0MBHkiJkNxdoWOCznDR20uscvF73NrXHxzngNI0ZwSE0lDzCnlMalOMrFDQxtBUA9lnT9cF
4mjJc09As/olmag+Mv/sg/SeMg+5xbpgdlt7GgSlnm4Be1MwQNAM7BDA2q9NxYRR0In91gLND1OR
bJpDTnMDf1p1qHzAuN3wEEGN5KUwUnH/eHT84Q/skJCHuJ6wC3vTfbKs63wDm13SNTx2WZj0Cy1M
w0/odO71prV0BfMFk4dpc/jn2wK4Fck+Z03Ob5LhjOWj8IuD12Z3d0jngBYIW6k0Ezw+mdbD536+
vii43gKuDPwAo/xiL5P1PAsR8rISp+TUJoxwsvm80BFD3fehV6RcWs7UQxl7/pak772Pm+wGr2nv
4m9Wwu+9gut+vBUZq5pP+44FRf0qvNUqwI68vflqSstOBFXmgiIDf5g+uIpZXuayJrqp+7Ql5BsK
rmx7/y+Fd39UUKMQe71XlHB0C2bafoNchao1FVnUA8lXv26xNUAQ5b8zDiBpmNIY2lSVCCeoAm22
v95TAxoYTRvesffXNr9srM+4jy+e/gzQ8TN+br5K0G/drlU+JUzkBMX6sq6nC30nLGb69uBRo1Ey
LbMQXktprGqxSkOltX5S6RxBUKByYO0GiBspNQNVzPIbYB/yr2Yqx/mLLS3YNq/P+hg24q8gOgy6
7d/3t0OQDO1MvUfs9nKcn1MjP6jXoYAER1GQ85Bvy9oP+H1lDegIltJUqAujv46h0qBlYwjsJ5gV
VT3dqg9diMuy1XmER9QquQDJ8yJPb9zJZ/nB2eUFi2Z913H/ifSA42CyFuo2au0MX56mS62YNofb
DfNbddkqBWVAIs1mZ1UlfqY7prKQaOWl9lew/ER07SCz/o8LMfwcoCc3wF2+Coe87sEdoM8Q/StA
4jegUg7MBHs6WhLuAaxfRArNqn47rMpY8AAqtnfkHmjR/eO39SFtg4ABjM1BjdNER+8pcLukFjN/
4jHGJvduaePGnMpVUsyG4R4dk+Vs36Z30rWonfJU8zB9DKLZopeMW1mX4XcJqEalsf/iTbMbUjek
fva+qEBhuYcYsOAn8oGssAUF9VXSJNy9XiV4C3p5lphbiqBNocyeII7KeQ5kbh4s69HtYmNOYZpR
0TZfhANj7SvVqHfYh0W8jlP5w6FDcjY1sDOTVBQw1rLTL8NBEGZPJkQ0JYoSKUkO3c+ge8nF0g9K
OrIfOE0/IXvpUzVwd4zibTW3t3LDSTHZNWPcz3rBQuoTKQ/GdBmI4g4XYtL++nKPhX7BqdbpigKL
3SY966V9iCbX7LqK9XzQib7KdCgL0JTOH/aXfHEU8mrtXMfh1x5vw9RBdONBvvbEA9lqVQHikUax
rPl3JOsng9KZ5r/jiz2WP5tQ+IjqGzT4nJi1iTJaGGFeNoCh0aq7PHZAQTseQRSmBuGN38s+CNnZ
EWXjQ8UAEB/LTjXX9KZUxZEhq/Zk2sQHVmiArm6dOyNUJrQLkncWO1SZ4g24LKgkulJIu8kLng4M
4+0C1tvBqKUElSDmFLnVTAI9caH6XJK0CQWNli66iOPvCTAT9f1yw18+POW3CwDwTaj0Hpv4nqMC
LAPkvy9TrqjPzwnN15l+jY3khLQkMOOOQoIezndRR7WIlFs157By/b/xlwJ6yPUrMI2+sOapGjMQ
+MzcO4M3sg1pBtK2wp9Lt8q0NywFUh/hMIcE3m8zzBU1PynqKyMxiKfVZ0TR+NSVK1ZrhwQLSkWP
TrUWLEc4e9TP5XbUrU7F6Cyn/Rwj5kFhZtdjqycdoE8I6ROwOerD8XkDnHI+ZoykCOCDVOy5Y3MP
CvDVbCGSAOlN9HHD/XDz1enL0ZFf8HPv7UYukdGAAkUcrsqAFNLEfKxKPFTXem5ihh6pkulNDm/G
GSdFESyQWsn+UbTa3AjDPGo4WkZ762WG3iz2H3YzmqGFUDD9wQKiFwTYDH4iOxY7mC6VWUaz9GR6
yUNT8KrCO6TgR0j+5oVbwdqNHgYPKveauib8SCaoKW6NMX1y/mMkGP80qM2gjgMemunGWhA/6upY
EjyVIAs8+vxH41A6pit4fmI9/n/g3edknNVdfdt8ZW8W7qz6gcj6SzVki6t53ZexYKqlcv7po3Ul
B5A0zRZcVNCbcIHO1yoj6js153RRD7T2798Q+VPe6gPiknfTQDj81xc2Ev8zIcFSySIk/S+O7C2j
te/6eOihyHz9pGSi1HokAQryq0z0MFSaBOW9zLlycaysT5vPjuovhNKnJcOoDA1Y8K9i0HRxZ2HF
YNoafUX//O9povgMh24LRVVFvqRs3WsKEmaklhsTS4YkY/oWqS4f/Lpl+tEs5I2hlrUzkjkpFeYf
5wReKGWoWingcm4J71g4aybL6SKMCJ9kduiLlrU4XahObVxZbDBouXgqcB2xOIjnbh68ml4wqO5b
GHpFldR38N0H2WFJovvbrPkyQnCyVjDWG11B4qC1MuWQ6zxD9IxfEMp1wsEiZPapK1d4EpiDssxl
b4To8Lt07TobPPl3fykmI9GYJ2yWgNpna/zPnHTSoiNR4tLZVgnS8sx9+Ia25GWS9SI40DdIue3X
or33xWC09PswptB3yB9Zx4qeoZziwc32LDDWDx+c6GSdrI9VmFateeNsKbvJWSpVfqDWGVUK/ln5
T9u5xriywVutFJbX/jl4ShBBhge4Jcm8Hefajpuey4czY6N9+FaClP9hDP0i0H9RC8laTzAZzx3T
PnuXvhh0AX5WnAcVkDW4Je3l6G+aSYaL/NhrBc2albhX6x34kGKh67tyEpdgaLO5AidjirGWVPf3
4+Zm9irHa0vmSNJAJSzHz7nPG0/1fZRsCO6tZad9fA4LUEyR2WxANWgae087aeMVXaU4Ku8Gtzkk
qtX4Rap9e7LtkEvOFdqp6rSuiq5A6oq83HvWzsBzdA2gsPROpHDO6/qj0Kk3Q9QdKInb1EOxsILe
fyQcR4kfgknINrIJvFkgDYsRr0XjIL376NVj6XV+paUaxUOA/4j1WAe0Jja+Abhr/CDgjfR26Z4w
NKLwJ1PmQwd8IUb3mvLF+1XlQVmwenidgqGah63OeW0v7UBPxJdrYpDvWlrVpKaCU888d3/b+aaI
8OGDZ81zBY7S/ZeyQRG/0NJROD6aIecDViXViT3hyGNZSCrcDkEZ1Rc2RUK7SFUQxe5IOcCpwpFc
TDSTqVJgm/bnBmx59GBiWxQy2xFiVVOu1RmlOEBxKbKCTmwIEu6zNvYi1cNUGYBwy31IawxUHFRF
nYEyx58KwYkVLtnQ+Rn8/mr4mTmeDbXVSYJ/87FxDsu02k7jXUzQr/XU7Gm5RU745rHxoCrrrvz3
oMvpC6BrwxpJSWydelNaEDT3qi26CS261oiyl4UYaNgvQp2Kmalz0uHZF+tFwq1pmUpqp1h6JUJX
33jdUYwLnte1rRceXnT+zvQySl2RwIIj5wFimQ4vmRea2hn5cKkFI+gYU0+bxfT7ss2WX+hJpn+O
4hIG1wHBtl/cCXAUitK9LitjqlP2TG2HinxNRltjcttln6PRqFN2Ew/jTKRYRl6d1nPLjuM6ki9w
JWuQUlUPxpLGSebjb6MslcGYrtgOxBnF9GhLr+p6UTy81q1F4ySetIKWbsAvFBz0D3hYS0hj9jMY
Tl161jwk9xUlavL8tAmYmXn+R4Xn2eTc2RldT5LfmFFhAWoG1+46T22IX38Tr0T2DJzrvkFQ64op
L9HZy8KyMjlM83PJlSjm/nEzJ6LCfcdUAFv6cL97MCTEidkLM8VajQEJBnR7hfemqZtkJy3TYE+A
sV76MWQjj3PHuZC5t0RUSW1VE1i3B2S7X1GwRr02SkoOy8HijPo6lkUm80b9eUF/4M5o2cPR1L/L
rl0uOq+2da9DHUAsMOoMpmQwH7NRNTsfdiul/RZO00kM+9ENN+VX/iLk3f1qlaw5lLvm6Swp5lfu
RDbtihvmtj1jFzqOezG10JAel4DdeWRWU2rmk27pfrjYMp5t/flDPXMRoGeYmsUi5kLy2isnMU3o
fTThnySwRQT3heFWhEduEUFrQPrQIPPrNG9HL+/Z2i9h9bE6+a6Hv0rVJvjEXbF5iLl+4daUtm7d
eTG06HXo7nr5C6ZMik3NK8mQAfciteb6oiU9fe6k/yEvfvV0S9aoePxa+lotQ940LI9NNMDIwuky
LR4vumSSckrNjc5HSFwTy1WikTXTSbNUVhFwbJt1S7hmRI48Y4pCcvyHcbBGPD/WBQiUzV6o0TaW
ZwNFxbYDMtgKD+VCE0UawbqoCoC2ANBcEBuC4SEjmwh5fNtfL0MSUW8q3EGGvADa/xvoESPHKDWM
v+DTP1Q0gR0wyMeta7kjJG5Dd8S5/H8I8dhrlzlhNIP+aiX+L2f1qF4ZQceDgo/CwSYlZUlc9LsE
5jc/SKh8RvH9xh/3FOEjtHJuAVwof43RwmSpNPSwruNpi1Q8TEB9/kCE7Z0nVMcLvMhNLeH6DiVC
+BYBmSkqpLnojDHcHdy+DaAdOUQzzG6cYEJWt8pzX27KF5eBQytHmc0mkMm9x4bRGdbgFy/zdrR0
itQLsAS73+ZJBVTIqM1MgA2344713IF1wIdN08DG4yBAw1uDpUApPIApWitA6iOPMRKftZl7oxg+
DzGYPUCBSH4MwOVc8tvai7hU19GP4ARVE/Cd5VNzGbtkAe7DW/9bjwlME0WsBIlvJAC90v9QfHcQ
4MreoVuU15vdubfgiEoorjl0qS4PqQEeyHLmNIsdupuWcbMuYKh0K+T+EuWnYn5ags6MrPg6Og84
KMew1cUQroHkAVr1L12zugZ0e8M1OMnzU8PKQbcTrhMqHgrieznP+1laXCTpQTqH083b0SvOPUVq
lZLwlRpZGj/wQGeAuhZOhy3fOVlFcGty+C9xqd0rreGcgvNvRLeP1XpBe62I5zYh+s99uuEBeGMV
pEvIE0VqhIGGprhwi/KIeqAlQ6jVbx8U/yWMBhjMtTF/yEsK0JIlYt1/98r1MQ1JWcem0inizb4q
aw1jLO9cAf/jirYgfx2LhKi7gbZsSXBLd71FajmjzrVZgotiC7WJCTqEy7JiHZ1WCwxDt26Gy48H
n1DLaab/9u3OHpOgI9gsDj+7bfeGfQoqK3MKci+l0Vx+8e7jt87qTtq+sJVuQLqDzsHkaEPW7eFM
NAe7qrdcXoCqyfPyCK0FTLEtsKDDVsffzAwUdeka6bYDciBG9OKOsQ7oRwEDCdzH60cWG1/qIFDK
Xr5w5bHg1l4NhZ4SlwrE1IeiXASDQAtdMeG+YYkMXBO5igmERqvVrj+Rp03XXmtlyinb5Kyaj4zP
QPtshs6NeIjXkoP2GfADWAfuIJ2juu1vWwOo9hfn5quhNuogmAKqH9fYB49FZ+ZORe8fi4KctnRG
uf9d8yG499s6HtQWGJu9UkvF+oQjttBkggKNiDr5CSoA+0f6SVGX0OsgCzNN5VFhsbkXAS82ONRi
TVP18+QO0+4iTNlmT8dTOpDlY27AXGsz1v4OK5jWgWbx56JiFPhcWibBPS1rPyAsmEHzuqtOHbNQ
H2xgqXhRbfa4+1zNCm6jqbK6sEhQVH5MhqAPPwiO3C8vB756UNci4oGD/JPa4s/Ui6nF2dKf1TNu
v55f02c2TLazWSGt0s5tmRUuSAAGqMS2gqeLDaL1OA6dYrRh7gInPfDRHFeegguLYBmv0CnROfnx
YjPWhg2RG5MpaFEkjleXK1LRCtrsEXOExNGf3DqcopzOZFsv+1h1L/co9LWG299uEbzE1bX0Uzk7
T1SWbu0DjQiLO7ub2D4mEmyI0pKx2ty/LwXiLA5pKiwN3H9mINv/WUh3lwi3yqNZVgIrSWJojMFh
CooryFcCH/bY1uPKT1Ea8Y3CNZA/8OX0c3x0Uspe1Gc58dK9LAgGM0DInCwTyEapaLJh8QUtWnbA
r6xRdHTum/xr3HFDbBvzOatae3PY2wtybyKvGPUkaFmVE9qRUYQ0xUKi9H2h1IMNaYzJOkixAuWI
yvhY5BQIDSWfNkSywTCDKMhSeLkCG5p7zUJ3XnHlU5AnQPVHTkCCYcF2mMZBsQKbT1ZTzlLkEvVc
Go2oLGAG1fQ1mKMPy1B4p80W8+8XggazaNa/ijxm+K0PrKHlvV+Zg2VEYeDoJyx2I7e2k+XeY3Uj
h+MZ3AvdG6z4Z4cW30Wf08ywjHyRUTrzH8hw+Pkc2QuDcFXP6erhh0Vk2/bySwcXIB/r1j09i2ko
AyD4uhZmfUDLGXTsJF8EyGkd12aYxSw9XQLxNI7uFZbqowwRjXRWsuo4Wy6Z2RU7y1mnoAPfFhjk
QqrWuhLLNl9iVA9U9npeM/74ywyigBshcZCLWp084hV/hlZhtIqxbLmPhlOEqQpAnQSzzmusJV65
OmSSoP1m+wL8cesMshj0o7L82XAH+/cNMa/32WErXUWr5clX6V1X3rqUiX1T29S9m4AlRjeYcYY/
9tQZYOWTFmG1Btqpl3BaVV6EWbzmD5UBHnsqLi5WXws1kgvtm9hyVGRoCpUg0ox4g88TioiOOU01
rpFJzomLUteayLY3F03YrVh9ndHJSNIEP/KgxA33LVZU8RdOaaXB9+LgMVVfusMS5ChyOM6gfBUb
VhUR4mpLnVVPVF2BoveiigeAYHImTBE5zHJJCliPxl86b94vSQ582OJGAuSqy0m3X5vXKJGJWzUo
+XgdWdZ4EGZQhI7czdczqGktkQraH+dgU2d9ZUgd+OrI1MMRRhXEk/hkrZ3v/7w6+3KE7pbaF2BT
hXh9e6CJOPz+X70RmzqfHqOXM3pUkS/FziUDj5ymPmk7uAzuvCBugEsSOqG1eHFzPUNdbbCYUV7z
JHGkeB/wVIOhI3008v9MRf/V35YspcJ4OpkWLdgOfw6v0hjgx+MecWEYiZLPAxz34TEv+34A02Dn
amTkE0jhHjiJ0e6WEA6sSKTxO3civlr+NnlpCbWDi6En3oFLFHadPKP3snxyGOAkjjLUfwZjk7aQ
N13I8a4sQPiSUCHiMoqnUqYElcQIED4ONrHnY35Mn0Cq87Blp+ISIOfsERHAjSnq03HGK2IP13G2
k8OreOQqiTtc0sVXMjQxUe2YY/K+/eOK68DNBlg46MtpaZ330gOR0spy3HfUg/TACBJa8giWO+k3
nO3xPQjWuif36Kes5BjQHe14pGq0Ztr1IWD/D67h3adZjzzk6k/no8hYa+3G6KuM2O7mzBAZu/fg
DTxUcrTGpgdG+iP6PIpNBi8y7/wgz9oyvdUJYZsiTSbzFEwQXlzHm9rmZ5vUS75nXVnyHz/05cNx
ADWIbylMpQ5XH2laiMA+GiHpMilhpRVd8PPrGaTgsfCGemHN3Bnmaa7qHMtQYkkt1P4ZYm720Zx5
imKFPu1m63kbE2x4vjqXMGUkUjRYN05nxS0e60Ob5huE0rRFjoWneAvt4b2GNsCv4GviiRk+KToD
O8FA8/9aHc4MONNePNElc+uKWYDjZSf3VRa+lwrJE5Axf07QLqND1ueQYrgMZCqn0nCamplXO0M8
ujj86+kKYFQGf/Bf3Mq+Tzie1tYkr5InnxJzqzAxvb+mLlobXz0PVCnV6fLHO7Z1+m/h/CE3re5b
FsareuxqBNrUn+SDEag1YRz/IEhE20woBaiRrsqb+uLEpghsafbb0kA408ej5k9oLTgV4WOpJyir
G9lmZJTNeZckYyJei7M3U783b9jyrYmiol9+KqpWx3vkFJSlnAu7kYA1exo+ZRdwdscxD061fZLO
Qxq5ikhRV49uManbeYMYxh3VlXfo0T8fU/rvZNkdSBOs4l9oPJMxhW6YjU07IsZzngYXZUmH5Ozp
Kkc43ZBMF4HAT5cT8KV2WERRKB9LnA0U5Uzin9Rh/upzRB9UL/Iux6FyobxBKbjfXAumFgOjnbQi
BdWLqlWYaDUj0xhbzVFZYA7x8hKgIyqq+6ksqQvCqkJOApWSNxgLxZWLvv4zu/u+DacCNArmkd7e
z4shUbW6uBcY/DYqheVG6mPvUVwBfHtmHX5tGfUTERHC9fdcROei8Kcd/Ld1Es8bCx0usZm1tSY8
zeap/HUeAnOpJLVMsbH4hL2Ily7IRjrMfFtXfnzEKYUdrC2hxnKb4CnSRaLHWXSHXTWebG3gZeZH
HvL7RWOVOeYyy74Pz1su+sOnckxLQBB3zwMI8R01ychXfZhn1OiuGe5zefGkj6j54kDTvvp/QimF
K9Wk0Ri+L5FZo0TdRf44JrFdKC0sfHG5SWUnU2BMN26dvftkU3MeleGOVCbn7HXr4hU9whiiawGB
nbv58nmUygAkhz27tfySHYnc48TMifwJ9GDWmMlqGSHjfinWFMSgfE2iVBEb+utO+SsPIhRg1VL6
dlPCREUKxHpkMgNIpP6Na5Y3yyKp1iNlU2DpIYKDtusfFkdAJ7euD3Q9t8Fq3x+D4gNMOzvs2Epx
IfgRztjtA+ZwzEGy0PcqwWR3hV2Bf4Q/q8JcS5Xx8tJUsrPfEjACmQdDrlSRzYL0Tlo7/BpNMgGd
lGoFdvCUZ0be5qhcYN5Z5tLmToF5iAhaYhh1nMqeFDiyTnlDIZST7SQXATsOYMIqqy1r+RXCKzUr
WDQJJhenAtpEBGOuxJ1pC5McnXNRuJcm7eFJrJpFREj0vZD/K2wL+kXG5EUuA6WzdmquMdBVv2wu
PeoBpWjoJW7MDtmE6DfuF5TIX7JrsvZT9wl7NuZ1iGLn3kBRRuNItQWTcB9/svXXuqzqvh+w+/4T
gDIBwCklAG420VXexPyJH0hvGrIipWVryDVFz6XPENujOpE+87LEb7eHIImDwNkaFncqdhbY4r0v
3+P9KwDeltdFlynpf/RyK/YrRv0LtefeEWQmU+GAmmxCuez+weRST+cd87Dez6m/fb2CPLgn/jWz
dZ+Qo0J5C+S1xD0I6ZmBlJAUCWWoP4YqLsW84jaF5zvVRYf/H6gCo2beWy5Q4CbBZSbjHtB+t2WV
iA+JrSv9OM/SPlNkhEfvCiw+PSOvpUOC4tPh8aMqfVDtyCIvG7xtdK60X/Aj9Pc7HTIcKdxqJxNM
fbAZgCU6ZtRl2HgCHJqPfEnm9M4iDRmCLle55BONdNhWGPHiUHsmGTFh2ievlbc0CMakeFjXXdqL
fQB13J5CHHRrqNNmECoG9Qvnl+RAm0kPQtrHrVoyW9aWkSGKAYBAJ/ui8XDyX5DMA3x0Ul+fm2K6
aF6+xkANCk011iorx1AC1XhWBx01xe0eu29YRkewifVOsMYPSmeAaADN73nLZn0x3QlIt4Fiq0a2
x0w6cXSgODBy9ktHl8fFbf9svyvq9TVzAjKB4MgOw2r6XsV/OcuFchb9DHbdawm5AC9wUbKoXtDh
x+InCdWpfayN6EBf9OtXmyjTV3C6bSBa5ue/c5mRpVv0k3S9jYIgkDnzNoQqnyPgBEZhTaAJHSPX
npq8BTt40Ggn7P3AAxRg9sEiCfmKGiBugbiAtfLXuEqugn9og6/bPhJa5EBXv94ZcxDSpfu9dyMz
5LohkuePyslQJUA0xLvToLq3JcVWkLCD9vvI4V8W/8yPtHgEkZGn80jKbSPboWkG2ri4Q+oIjNJW
0GpVLPWJCHt4dILdD6pTjVAaQv6lFpSFioadU45SKVHEzl/jkozbbUCp56UA6FWk3SJirt8HKzFr
eBkYwAcjeTjf2YrsD3gVwUy83+wwd83b0Z/XfN4nlQHWypWq01pwHqnh4Vc/d3uf5EjbB0Mzr1Wy
4Q0EzlqEU+TJxsZhlodaGCpeYhyBt1tbLQEuOJc/4gT1hn8cLb+sUt01zPHpIcHwf3knd9QaHx7i
8sUBFKlzy/9s0SLZZ0UAyiydLuIOvDi7wGX6InLjUoyEl8WJ5OnEKWI7vCOpgEIOxLTiaS3SJ3Kr
ODBvnzZGWWqR+yab3wYDT6BOmVWfuEERXfgfToFDH1BotJXgBYIh+Jb0QhjDr4GwvPQ0WPLwdsNl
DlIbD7tKaVQbha2QydtATCqRkGtDLZ0vTEzGOk56cNwuTWc8yNRQleF2R6qTJBMgb1wlFRgjKOyy
Hwpd+rB3vkV7gFiV6MwbjLkq702XrMuOFp3hKXwD6JYtorfFDS6XmnbbNcQTowHMdAbAMvYVep7B
WlpWy9YiKR4ZORA344WmcBWwwZJvkl2JBfbdKUzPjhx1LUxuH6QmdsNgiQ+yG58rqAi13Y/wiayy
+7FxW3Rb6yGLVVSfR6xqycRNdcniGe/3sWORLUHgm1PYTqKsHe2yXaYetcoel0EWxksaV4w95j+f
MqJbl3jgI43yFsqeT1u2UCShBxEgXLvTQSZFpcdguvqiuqOhHiDisp3pJ2kxNBDW8taThrgCp0hr
YMe2TcgEs08oZf1oUHDrGcdFjW6f8XsWmDA2kcqK0IQkPLUcEj/iZuq04e/auTuMXY8poq4+53Wa
8IycaKgcMbMmNAieKpH+vG2z0gPbUIWeKyVpytfcA+sRTsoXCUFz0NpxW2vEP30BI0DddEmM8JSi
T6nvdv8LZ0rDUabHbAz/l+icH+PiYkl25jHH/jswWuxqqktLTClp2kdDBbnvueJaB8PaJAWqcAnB
1NwFzYiNx92+m3oSUY11MwrEJHk+Dab8IcwXpZ6hcEPPZWgwD2flGni6cjuqd5WVDW9PF50y9FmT
SvgYlBWA5yTHM8tdM9ec5fg9qjxCFwuZZoRO7HGJd85bwGS6NZNuFgagiGUQMfXpTWwfD0NzrEGL
l36KbWmxgEyrvt8qz+/i6GQ1KyfCDkNL2lOQ37XbLAq0riekbh//N0/INWlyltugVHDZmy4AVeId
ZSmwbRJ/pQbdNKGHMfASKy1jIwzMABXtylESQniTZ9a6veJHsYDb8Th7O/3jIwxI2X1OCOYl+EqQ
qrDJl8g6SE+bor9vCWqMfwSNPPQdpK5VgXXsUcksXqhk1FSTalEdW0av1Av9LxVrUHE6/t/lVetZ
xmg7paAoC8YLjHUnaiX0DNRn9/2pp1YIRBKhP2sfLXwgX3pgNBXke0fFRf96cN0ym1R+tfVZHrYf
/SmtGnclCkg37pbHep6k4ooPT5t2HW6WLqKpF2mrqsCIwDgnUhM4fSCF3Ui5iYN6dII1oCGn3Gvm
kxOkPGTrERkAmpQR4AOzPmTj0/0PwtYs2gUkMnsG/QzduaCwPwOnjxYGQt5h3uYmPVhBh3zg5Hmx
jMQET+DpMAssCcC7OOqmnwrKvhotX4PSKec9L8Ppwgm+RAyrLxs/NuLHnrkcOcGDj1JaV5ZKYtDK
H+C77QyJmnieY78JC4ot7v//764r1P8QNCXIeCVLNCxAwuDOqEO63+hrIt2hXivhSeXKhF6Vpv47
iHl4W89hDp+EUIpRblK/2wFTzOyHvN7taMFiirVwFl+4025biNjP4SfCzulylvLbLgPnRFXh24Lr
pXkZ7vmJpVfG4cSM89+hqCfwSpA7VoJMQgONlqNp6tH+vglswSlGCDs2hxfFYvM8lZBRSnbSqpSP
+GjbuVvQDdZuCtHvO84bKvZVt5jagI5gZELgdJ3LTMvrxD1FXEuO2UlOJCis2uteJhChFT/e0ECT
1SQ+7P6lDx7t2uvow1rncz2tDEm3fiwtTDZAbzeVm/Jy5bKgnIYmZCmjp4b2DGysmQ42YA8bwHxn
TZGyj0l+/PCwrdqUnmPQmqF6EyAZ3yr0A+/rVN24lhcKJK4A7llcSMmuPMu0JtH9kVXdTy0SKdho
vkaOYL8gNrjwcmzqTXiW6AMOaNLbh2ptRtRS9EDC44GiAb7XUAEfgBjKrW1hpFrNMvbOI+lv4mzC
1LDCHsu1Y1Btc7J/JNIhukekzAITdiTHOW82hthnV7PKDRfDTW3PjJfxE49rS9z5zZxmYHiuCxLT
47FK28nPK+fQeU40jCNNFJfi9WLK+U5QjiVi/g0UIyv9T4unZpq6dFFmI385RTC0PsVUjLlW8Pr+
D+hQPAKaFOknt9r/RneaUk1Av1EFzmEm9985YnDCoiAS7xEQc6VHSvkstmi8UPh6RlGZUmroEey5
IEXAge6Q/qcsYHMxc5G8K1kEx2ZptPftUSWlwU0pb/lJPxTtb9PhnIdJzHDRmSbx29XT8ycXQ3ly
xSTaKRBCZdjK5+oMnQ2urhvkCy2ztS/KJkDFTlYkgLo5Fqooif3sy9XbB3Zp8d7Hkcyymo3zKdGH
reoTq6OPI7cILUc7c8239Y2xN5iudeD0ojuvMvy9bpAcQK1QNihGgkG8c6ilRp/smvdrHkfqJPr2
VbSySngkCYVwLFNvrKVA7KfSbLihJdQ84Insd9mkIUoFITTB8fP5Ngm1R0rt0K97gwYtQXf39ua7
ebQeiV2HDgq6bx/mapQSlPgyyqaRvugHl4o7PrAtst2WOmtnT2kgYhEmKSqZ/CX/renffQBgmXux
R+UHe1do7ehOqegsNDbaRN0a4fctMgm4CoYA/vl/Yev4htnNt3dv8iH7QDC/B0Xdgkxq9n3cVtSo
u5AmEIU5D7JrIGuU79ITvreHULoJDT6VMbGMubSiiKR09EsfD1fRY3RTXkFaYjAM5NFQ2oWPfLlB
60ph9zSkv9uT8R9WFuu5/0yWt6xP9fzJ+FHzUj3c2mZRONmqyy1qgzAQFKPyOZu1SjN8aZeG2VKj
tjd4FJu5qGsh7bFZGLsDDD1dF5l0IbF4Wwk3akRTWuneMKZQfjQBiqtOJP1B2NoxQtzh9xIKEJOi
ryTz9tNwEraeQcTin6BMQNg6/M7vG/T0Xj9jInARncEEEYdjB9wIOLsnz+mCO9lmKUXvEk9f6oQ9
62rFubxJSokGJyRIYT9iKXg0Vulo1us2z7QufrVIwTviGwT/XRZ0MUts+iVUQWF4rVtxjj9gixj5
A9NtyBzXnekd67YBS+jvkEo3BSmp4vZt6bIGRV6yGkBlNv5HoXg2GqfUDJsUgIwpP7Tqb9Xety9Q
Np49Ayd1/gZmHfX4hZCDOAk1NpsG60sTAdortgkVmadPFW5Bvy31QoWy6K0PP8aXMfiCh7w2AdR6
TGXTRmRin/0R26RqjC8bCdwDTNgYXpANT3lpqUO2jV1SCRTx00hP6Hl1oZAYaR39bZ76Uuj/zICU
qRQavuNnzyNpZgsur+HLMw5+nzch6GiisTo4CHbBvFg92Vq9pq6zOo3teCASYLEog0PBjObJ4qJe
hGgPPNOhtAL5p5xiSxKHs83UtQIA/ApY8x3+FuFfR4MPLqsSpYMuBSSnFiRuJn4p/FjCbd29VPpf
0f5chPbKH1ghBEBi7zfPsBUFLOtmU/C4erEM9OIPlINco7MZZZ4RO4Cl/jGIophYijv7rjXXSfKg
PZC+t+P0ZkZRVqSQjqBig//aHJBku5c3g3WWl4f6w6nzHAqCCxflu4yN4M/UQg328iC/fbsxcBlp
kl9uNu2G8AES07PRRD5huZzib/IrH+ShxyDB7F+7YsnRmvaWTkM5eMr2EmWVwO11LcaxDr6Ztvjt
pRKXuVz9ppleYEdRBUzI8hmz1ytDsl7tCKivGSo+bjMIdYKdV7RKT0Q1NbMvTm0dhBKX1vFE07Vp
S0knMf2Q4V9yqPCJXwiMpnGaGtSpfynk1by1mRBS866zzurH7QXMqQq9MgeS/vcK1pDWuCDoNBed
bLTWAcEEzoVg8W0198aGcALLykF1YHJveRY9+LkhG1E/Jv/O37w9Bq/XFRfI0RCcJOenJpNHc5vH
JsWwF7EepYNFMn4mMZh1OjV0kin7pb7+ftssVHRdXi9Davk9j2fg2ljDNr+4+EfepqG9L1SuuLaB
RJT1gRVVKb2sWF/KMNIxH1xZb6Mhj50vfBFXIFJcb9us9m5dqIt17J2f4fRjVzB3uL1pg2q5jCq8
cGBroK9hzZbztdDx8IdizUQ7Qog0mteMaZscZ4oTXSt7iRWCrzCWS8HElONzDwGckEPqltEBOHZE
xzugy6lupdRGv0UstK8r9jHN8HxRrtR7CB3vFzvVA9Nri8YTPjWEcJW0eoUvFsIR5Trmo2kENNnY
HdZXeEVbHX8qy4AnGBGwFVomJYRuFYgPFz5Di/ieMb1yWhl5z9bgSlWdYw5F7Y8Sun13UY6412Xg
L5UeSDgih84NwCD2Z64Z5cn9vvxCtcoqTRypwJxy1AhzPPX3y9p2xZzfi2OtzFIVCOXXQ5YRc7uX
AJGZSJH0iuyB1zKe3sjIkcZ3z1VNNEzrp0JfWq3KOiklbUtZgvLrH6ZHl0wpqvRMi1GjA4ib6d2W
K3ROhkSlGseDpyt0Mup2vC2VtvMqYupTX6pUV3b7EZumgROe63ZkSjF14muXdOM0ETBmVF354gEe
GrxCfQM2zdRxWOJTud/ipAhDXiDx2KC/D/dSGBWj/bZdaI2X/aJlwbtoK+4ECqKg0soM6ynRnSXJ
3vahUGyfLBzOiaERvj5yGKnbdmRi5fSlblSPvfOjJ68DbjIienkOAbpQ67KqlNmozJ33J/a/cOXE
r/HI4ylaxLEILXdTL409jFnUtRUK3fXah3vwQwrVU3vHVRyPpLnJ+BbCzqbnyAyHHUfd1OMj4t5D
AnoQoOnuwnnRgWXF9//QKaCfpZSbFW55PClg2jnq2jLiFtm4PQcAsgEOESxKPsby8m3n26ERfGse
hf+HYu9v208dSe2ddOKZmksGPXMjY3gXmGcOwsTXmGi+07fU6ts9+6gnBnAROEk8g/3l28E6v2R4
2QpAypdC5W614+SQotiSSRi8BevIVV1m6j9qUOtfdpNsczlVGc7yLa70wK1hbBGGfFhE58UYE/CY
OjKM+FLZfnih2ojps7VsDIqaA6SVh7GkX4c9uIpbMTRALsPjZlmB6Ebigct5MSvwDoh2EW+kTWqb
v8bnzURNwL5sSTfhT2oduciV0KOIfthbedNr2x33HHdTbvYWmyWDTxYUeVTTPD2Vda1yZXbozGr3
9JEkrRiVFOlS1wnwnoKFVc68I2j32gxXTojd0akB/AoRFm2729kEfwuDWG/NjSqqNS4eCnmRmc8s
oSD05FMbbPMEnnBNfSZVH2dFXCMjyZ/FCOyYN+WPeahWqXq00s2kK//WWHdcJkuEwhj46ArYVXZS
ABbmdXfaqIW81lkNN6jbUGg47U7hhxTvfsXoGTIzJXh99ZBNXBcjO3nKTGptyD13/rwNQr2gVffp
X2riVf+l1+EINmUh9U6t3Kjem5/8XsS91KwszaJOYxP7t09MroTy3hQGmOff8sugOMfBWneGXo5V
kI/GEphUphxGEmibUNAGY0sDc7zCVPz9mESumTt3SNmpBl3kQVJAzo05ix+zeZn1P5qC4ob9hzVg
fyxBDV0W5c041CIjpSDXQNYU1pCkHzsQCfGZs00Zp3F50dmz+gFUBG7bj9d78FUVPcb8jag64Tdp
QuEqpbVkq2N0JTmI/cdmmQ9k6RH9aQ2bssaoN55xd9S11v/yyJR0Os1lpudP9DwnSHbvdT4rVSmK
pMYYqeg9vCS3j5NEOQ4rZu97QJw+3vBDwlBjqZcvQIxVQngAeM+6Kv2MY4YqEqHCccsA09JShbt3
Xig7iHLe4iOONTb1xSRBr1k3XGVW9nt8sA7coQE2kft5FpNg0yii+i6dWzvDBGj76YDYOv3nEx3Y
AWodvNLikminh2SA2DvFcLDMaM1zWz3Sv2DpXcn8AXNe5cTFBA2xCGbroFGWNS4NznfYbJZjRUZo
9pPYPl/eMQ4UvM8uC+9oTZSVXud7MJUrmJ4g9ph2/ceSO3POI0U5umummSUvQ0oj9g6+ba53wSWP
S2B1iD9lwukBZEJk9NQP5UHT+f0EGIP+oasEktm+ZRM1cc8ypHxoGE3smdkL+IjKOYJP7xD2KnTG
RiRwmdEvAV/2AvXSOiWx8RJkkRguQ+qMb78LUXd377SfZEdFKu6PvIYGozTtXduT5ZCAmhKAVzcK
IVXxvoGZJ/BdhSqDmCbnDMCM3caR0FXw7YHZX4T/BTWIb3mBDCiWC1IQTS8RO56YlpK+zijMgjnU
HOUSoje4wUUXtDPMnuc++foHGUMgDh7llkTyTXLcwu0XGFAXh2hl35rnhHJXsxMWLIPjzawxZv4e
2ZU2OL4tDqkvhXGi+xfm7/JcV4DxifqcxDEqNzld41JO2OjPPNsIyNc1x6a77J9843VkpHfjwUPt
S89/ibAsp12ws2u/E1EFnSfdlD8juF6KfOt74zurl27igzfDmA9d7xCr7IfHFZlm5/vvQbhbpELE
Q8N/cKg6j08pUkEzmWrrkZmBKjRF7bfFBNuS7npNZzL5PChGex8zpLMNGDjZoHaSuIdpSuB+9di5
gOYFa6ycgauSjeOnAbdGtKIlh4+cc0Jv09poViYKIwfLxxoESSu2IkKmT7nwdHSaPCNqkyqr5Dna
p4GYPTgOl0Jj8UjCsO4qJsgSB6d5tOKLO1ycveWVlIcJf11O795NPyAcW3axJl5weJLi0CtC1fEk
WPKWuNga6oVk6lN7mVGppBeklwr+QpOmsAoMdxvuNCS7TPevezvB2B9zS7RpHI4UQ7w/GMCOlGeP
tTN/pr0SLVLrdMT3AfRk85Q1YUSH/UDo5T8lq/D/aLDMcB7KT2n+r4ZQbIsUEujweNFGrE9aMfwG
QfRZt+Bhz24E8u8n83qaR9SGvYz9vAUHdwDq68MPqWlEvUu75Z/hIHq1akXLoXuEuQ1k1jNkPwo4
qR1ARSVDxwNlLKpNFfdlbzAycYs0j5vli+xY3xFC1ZakgssLAQWrthNCd6bJErxYFfM0PM6EFL6b
LhyX6d1sGjSDYz4T32OHEmZzRKCC/+7ZW18I7+P4YgCEsOZNniHpXZZ9phj8W+etvMOIqldt+zai
ZV3zcq6eNbKlb8uBlDOC35bm6r69Zis4WuSjM0r8Axa+K5xCSuuKt8/wz5nOWucHIe/PilAvAfkr
e0bfoXN+8HFEXqARYU5xtSnIbUgzszZndO0kNcxsb6nDuI9ZZBijqolLxkbyKIHBp8boVy9hqLRA
dHfaoJqk37s2qQZO8rHG0XmelVX7V+WcldR9ZatprAhGdTbcxVP117MLZmAInGVP6RUx/w6dfHN1
WhjvTjRB1PLD9VJJOiJJPRVMkQ93myArpSupNHii5f+9C2+iJ7HInJG0mN/GsnNscpWUFrpuRtkj
X4wybTsxM2sgTVCnlK3g/Tew6HJzBLXO1Ff4kuuCygH+AZYt5yUAOMBruM2bljSagEeWbe3ZEqAw
Yd6w7phq9pkJCwPPdX5aBV7yfQ/lCSA8dYaUtMT/9COmo7XjhW9w76LUTwcrinD+ecf9D4Dr3NaV
63amwdqj88jLUYDxnSRzr/o5W76EfkXVRrUjG7UudA8T66eq5Q9JIMuVrjD5HfWGKcWpiokLJhbM
ZhevwFIQIWjrf37P0zdpB9F7vI7++AIL0iRltWK1M8pWmAdW7EdnNGOxvmnI03ZOaWRIn0rYLmVO
AyTU4WX42UM3i5I+2dvmraBg3GT3+bv2dC5fv/yW3KPyf4YQuHxy6vvrXOKw3CCX1zkzDNTFVe/p
LaXA3kWHpgQsjNsiW5IaCAUbje18N2Bf0KcII/QwJcQYNhlcifBz+Nf7LaLZJVA54TTbXSuRHRma
lr1usmvkWtI+F7eBbogmyxljUeF4SYZOuZGLankGS2BakJ7Htoiyw2NUZW/AfkMKLb8SanG8MH9/
ojpoYiSFYhHNN4PHpAJgfnKkJJ1d/Psn1iV8WptyLE3YiF8IDQzhzlJkP8gEieKEc/FnZGStKTaW
IQBz+jyyPdwU9oyvWpDDOYU/zNkMbuzq+APbh3xVZZuAZFFc6peMcU98x11/n4uhT+p4ZEwa+B1m
TmPRbTIiGY7Jz1bPpIKxBWEWJ2kR/tMkAuxzY/8QunAISVFaTmkn00JuOFb8lnsWSY5P2a7g4efm
avlWGrpQ593buKQo08zSjMMke7Kqv4UZZuz1SGqqxF033qUJZaz75EmBcnPzVh1uP/HKCZxAnYaw
vgO+KohWzDQDlugEhv7faekhDiGK8Xf8Wcp+J6KGskrM8Xw2hTCsVX/2SCBFTIV2ON3yEwD8+5q+
ZEqvXihkRZxtaW94S6r/tfcBDuS0Y5S7OrN1jQh21LIwRTSKLZFAYx/pc5ehdvBFQiBILoLYPyEq
KrnIb9rZBV2pFcDxe1WuRseKXFs4mqaA0+DGfBUyFAhabirwOf9SiSOovojtrK9GkxWh+eAoJYkI
lqcFTSZi6gr0U7MoDLQmnCwrDKm9GlV7s31puGVs0TMEE5XQC24eTPKv1oSME5MuUeQStddIcBre
G+QGJHiTcSytB1SclKs6jkClKol0S3ehE50L9FwsGAG9rFWkvjyOISFTUve8Ww/a7tAe9Q2Q/OOA
x0lN4DFOUe/KnbwU5Gyp+slAENAixOdEh3dRRJAaGPfqeoARyqtLHEPCs8GB5z8pMhyojMJVOywf
dowuGI7FpTwmwbHG/UJ55i6TQR6r3Ah1xAeHrbfhCeRpBoJM4xzCwnKMCUd5fBrnqXb/hCG7wB2r
L+kMV0kUGlUkjOmCJ+MEDEBC/tE5ZwDecCuEuje3CVNu7bUvkc3S7VeD3oJpoHDEj+pdia77gX2L
OeUtV4p30RYEGRljKV8cXmmYTDlft76wOYxf2peEecrnbC3blidk1LWzxpwWPg0AHND3NQx4G2sn
yFndbKPre0WiCs8MZ7r+wtWi9yCQbgZVRTLLWmVLEfm7lWdnpNKjDQI0IyvAnfQTSQ+erlU5hulK
54IJnTBt04XvACR9QHRa+2z7o7hLghBM6W6WppRkfXtbFdt+5qw4M97m8++HOWNxNBJQUCr7IxMC
W5GQJDlfaNjdRpnTCXQYd+Igtga6HqPC/jVgy7s6v6TEJF7w7KtyTcDDeTudWTsSSyADyZPLlFvM
l3Ljl3NNSsasBHfhMNebBLP9Nitr7JnERXPZGiLYWX4gjJ/7EhsqpzKW9NmLgyDMCfjSzB8lCmA8
RFxx93A+y8DO6vvWASONG76ut4vS1qocyoES6Hx5N/L3260bqY3c+aQzwAH9LfB7rTr15hEWieeo
eOsYBjDe1zh2vaT0+G7SMjM9PTzSGusUm56O5hBcMxfGQh5rzDvJEbt9ul7V5qpypBJpY0+fo8Eu
dcZJ2yVITomOpTpm73iIFblQtXyxdm3c5k4lRB3VAGjhYDUE4W54+CCPfd+MaUlkgCexQoOAW0Jd
nHX0e/ns0qn3Dco0gYLOISSTsB3FidLQ2c6hR4OMfRoY77eOBBE6DqPthfkK5M9ZFjpa7H68jCAF
lw11tylEkSTGuHgZ/wdzClEImwVRzM/S+8AKuWHfBnaK4nRpGBMcepuw1YTKHXLKJbcRqqFtHDLr
hfdTIsGIg3q5O5k4KFMuRo7AEuDIY0HVAAOmbwR5T+2AtsQP7oIeKu+YZSDh+VxERyebTRDPuaoo
Tg9Ks1KEGoOTiOkViBSgsxvkkGc7HoURNagIofl1PkGe9OQxSBSb8F7DMjOyJ1UjL5uUK+VAPHgT
Rj8Xt3Uwc7gJMW/j3sek8BXztsAe8KXZVqglttl2E3cAKcKyrxO7pkenikAHfD/4CwA2sFJmVHP4
Nxg5ODmPkUPGqVyN9sdJEG4u1EvQmujXJFlGDP6gKSexCyZjIvD5Jz0e9tHOmFIqj7sv5DyZHZum
rCKRvjoNw2Mr0a4Pkr/ziETcIv0Rm88nCeGjHLmj6qcbG9cT6VaGlxLL6AYSg4y6d3lXouLlhyMl
2H+aHlLt96sgDVmWpTwjPkfUhR7ZjdYkXKXrpXe0zy9S4xPN+Qr2/mJUlwBdSNEWVel1xy4ykrYP
FO9G+y5yYYhV4/gwbjBE74+TzmYcujcs3I0EuSefWiIhXXiceqO1gmxcQsGAzyd6yk4FcN/Wfc1s
ZSZR5njXa5YSmCEl/uI4xpwPS2B1eXYKbsHRVIAGLXEUSR9WHSSHbyNHYdPjW82YQwU9p/xKkfni
1wYXNDCi/K153m6h2IwnSG2r5oXTH5Je+rW+eqts1Aidm7vzsI40iYX8H7VPOE6dZTUs8kAQXuGa
IDL4RMsaHQgH/f29DHqeBCaBXK3tzmoxhsXWu/PvhrTL+q4AIGjhoTR7II3BAp0IgykYIWLihvX7
fk9QTFFDJQcc+MQ/9toHPj/tWWDxIAjKsWALagKiz3rSBc0XmoqjyWe1jZux+9/cRtPvK2woY9Cj
DRbPROJfxq9PzNBqJUL+Ozsv5HmJ16AHU6Rs8JBNW2kfdq+WVqn2eDFHSRmNU9huDUQqDE+XO1Ld
WIy6PmdHbKMGNU6FW+zMvAO6NpqjbCgxE4AOhaXV5FCqr0zV6f3MBYuaEk12t+PZ8iKdKq3UJBJ4
w8/9Z7LaZxRQ6jiEQaFxs/BovcijeqaLQMYlmW60fbSXla6CjofN2bX0ByOU3HwcM/Tb9+EgHLFt
2mwj5BO2QHGpyr3ZnuCLsRppFrj2mTv5Qp2JJDQPY8czMdCny93MGo+LDasZE6zzimcfjaozYVL9
FGMxQD9TcsTjqxUdUCK5ZU6xwXEZ/t4a238a0JxnhI+rhLqCkNxc3/y9Q2YYf0S9CifD6NpLDOJp
AlQkYm9l4qAWbLM0Esv86lrxLIMFd/lDUrPBsSnV9rzAxaBVAkv8mlVBcROjEu7NZ3T29PeGdFD0
3ywHVD4KAZkHIrZFGD9LVg3GRNFMCTig8UbpMfZbqY/I1NsXH8rhsgT5MybGn7jzsj1tlXE2J87Z
3d2ElHo+QmPm6ybgBP1djV8aIS40U0tt25iejTgBwWc40vhl5TojriNLUIWvNsF9Pv9bZ8A7M+9K
Ay8wMgqabPDrr7SZRMY+xUsu062od+YKBZv++meNUkPMviFFu3sht+HTn0pUUD/HLxGg95R+XPtF
28KqOeOzC0R6IIPGRaYTJ/RJTy0GcBgfDYRW3AJLCJPCWc56W5KX+XVYq0KmrOwkbgps0Myv+edB
HiLzpTHExJQuS3kJoqb9gQEJqnLgbE1Qw6tIicaQfZOkN5jSOEuSB5nLLakeeywvyW0vDjhqDqSC
ujlafaLVzJyn79I9AqL/+UWF64u0uNMb4OEytddrAgXAMEIKB7KuVtFJ/DP11rGGdgzyfJpJEDsg
0iwfNsbOi3HCSQ42PhSBeRQS0hxqsrT8A/FqdMmJJEZAU3DfKxgqPJwEIxjgMq0xYPbSZ40roLPx
d86xNn+6FiC6aqyzxEsc1bEVa3TkXA2pmfZHhpLfiu3B5kI34myj82PdljiT+BOIkOrimrvPb5v7
+Z66ZNNvE9LXq6r2nlha6qq5Ysud6nM0G4nRO7LEnbRM9EXMi8KiLEOIiYI7Wzw/OAVRch2oeNBX
3QbEYJLhOp2rhP4dHmc1fyZk0hb9Nctl9TVjWpj/sfVjZ37zpp56lShyoUH0mlMLqxGHo1uKlN6a
gHL5+GAAaNbRF1s3RsYIJ6WN3qCpP+onUgZIWppcx9LpnUY5n/yvJLJe7AjrgIltPa7zFNjcvuTv
wd7WgRH9xdVuMoiOUM+KnQrdwRSxu4K63i85nBfs8V65O1Ku3KTz/se4ABqG6JDjtQi1ODXnd+lR
zb6bUgg31VzQitgePb4Xrl50HgHytRp68iD6pTv91LqX/r6nytOMIBBEdNKQEkZDnsMIjA8PLfMS
5xT8bfnIIDayW0xmvamzyHGKPiTdBZyAD2I7a0T2G0TE9dXBYy3oyQjxqgCD8HEtVxTvvE6KIZ7P
AFyWId1Koe/L2b1tqE456cHEudrAX+QNeF2Ns2146CQZYfsJNdfMtVZAyNmdfpgMRCwDVaJA9unV
FVGfxPKZtUOC7ACHLsHEuI1fuEbcmQ1N/Kofqrac33P+zHWxguWSRtwSb4tURJwQz3vcMj6jMf9c
BGHHwNjwrrJx7AKmEPBW+hdt4Zanddb9rKNtiEPF2jLnWk5WFRthWd5SpOAI5VXgggh5qNmFnjAr
GufMhhfU66AzK1puaPA1ez2jlZGyEBY/ClOFVw5scdZXAu63kY5zoUwytKNepsa/Rgyxu3a7GWlG
qPseSGqlzCJTK9Bm0hT6Apg/Yks+zJRA4mvTiF7x6+9atAXnSf8NioTHSZSpQ2OHXCjio6LMVfrG
y2gtQ/497uO1Zo+gA76i0SnoLOLBfnSc3ilV4AVPQ1J2iMDEEGWQaKNqwJe6a1fVUOjn3dVMHaFF
pC8MgF9/gkrpiqUsyhHF4AQt76pi00X6/qNV61teEkbR0bx8wvcli7WJI4lr41QWrYIn0Witd8IG
5/PSq+U/RK/NaR5dTHgNXJpE04+Ia/oHTkvtlBVG6ckK+vstZZcc+m7Zpxn9kpIK4TiUvigY0XiJ
wXUoPJlYCmQqXVlMRHmXgYQeJuTm82dteokVHj6PWKk8waiBWbchHbv7s0wKntEXInS3ng3wsAtz
UosmogAs3Kvm0iD7LbBQZLMwfmXKlzpiaYXf2keHQsMuEBvzsBidGBvLJ72+rLLg5FlAVz+PyXQe
1zJ5rNBHHQMiCIfbFh3yE8k5nWvw1CTT4vEUSTuqwErfyDt7d4i+YFD5/E4binc68rWhGZVl0bUA
bimLZN2DS3o3/xwMZogd6RWV7k/molmSj0i5t7hZpeS2IcYamyl5u5gy3NxT/q40zWldyqgoaJti
RFf7JeH//sieHID9sk2z2SMXi/WYMNUwSzI5W8YZSyDBOfWoi7qv6cYylFE5M+p7GU8czeYB4wl2
7EQHAalOeYR03VQFakmmzZs3RNiZOCaRXxe3phjn+BVZcKJvoLs88c0IjIvrZYHmPfkhMjITcSg6
VbPOcQ6iBgYdk6G+uk5mgMyAg4/KJdNsWYnsMNcMtaDda1hj/z0iU5JJhzel3Dk/GeLFqpcSzqVU
1mz9iMVfYAERvTxxw45RZuLLGIpN7BeFCDoA7PSvEABCS9Yn6isLlUeMbz+lmgkJ5EH/mh3Ozf7d
9Jb2WzRB4B6/IXCQAm/i0u7pVFA7n2fteejO0Myo9rqKsRPy87dSczMQAD8fiyJdQJipdGp0tHyh
a9bQuw6wD+2Qw8o+/njDz7MB+rOE6ObUkAhRhWRkwfEBVz2UtSJNxQ3eC1NzpaJKbvzBGhhmTznc
aMMv1J9lMYX2ZMDWTDzB9QCW8uIcN6m5R9UDet8KEtLY1mzt2LEUPi0Q6p0h6mv4ndgLFpH6SyfY
ma2kADJP6+Pmm/PG79U2m7pKam/aoMpRTmX8kjnhbDZvym4BW514Q/c1Hc/J1SDy9IRUAba0BgKZ
S6A9Bj36ebzw6kR+q1yf3yh43BNuMIZywcAZEx0PJd4aYnY3wDTncXar81QDTIp4OzD+cvZD9Kag
kCJWwZR8TXGSxHO83H0qmmd7qmb18rr8/Bb8N6uIE6YjWLUfVmhnhEFCqiia88X8O87hzEUj1bfR
dcVqsBPsukf0hPiKz/0/aBzaIvKulvqya6syWCepTOvT/BP39zp4x0oG8aHY+K4yMB0oMmREc76c
aNfNdp7S2uWpa+KoUJ247ZIPYstFqe1TsVWbunES2d+lbGxt+xOH4UxzCdWIERvI2ZCKJHZ/gxoS
ZxkpCv5JNfvDNDb6E5v0I27DC/1DtXUCnHYnBmDbkIPMlDDr3bf/lwDgaW9mldXKzvirZgCPm+G7
B1+WDz8x3lVbZq3PfV4MiZ5v8A8vSXfevz7WkIF8Z78SUxPojXJKmmN7y4X266hxaAjpi4ib1pT/
lSUJaz5xNe7PM6HzIpcsqpKrS06B6sLKyn/U7pCScI5oaS6jmf0NzhgUy2kwbsljHGSi828OAWe7
lLahsTRjt2BzHD4lDpHbrNgBkxDkzBPsxmS0AhJ2QyuRMdtT7KUOA0mZhREotbERuCm2okQHPF69
ar0k1j/n/zvtgG5qEbiMuKg+rNgPh6wXJkei7mGs0dib46APyeVVzVNGTPvx4WOW3w6nczc7Wkoe
bvRWj6A2vUTePfrGR9CxRD5fNBhtPNCwgqMzDqkLpFF4rbvc65UBPVU/r1c8ikkgStI9swK38UAT
xoOep5RWiz2enFL+viBRe0dhApXMU59fF+HsZPxQ9DJj4T1pUPSpGJZPR4uPiiwmvy10biEQmSuY
oZXKGSb0QA07HBf/oMfai0us5BJ6Ch2hxzUCaD4IXtC3TuySkCDSLzLHU3+yJySxHoh93Gk5v6w4
548120bLGhlFFwVcZ4fILtTkAnjh3iA2r3KuQrVOMllF6ohN6ChTShSWcnd+iylT+XZkC8c+wgdz
SjhSaPfzAurNdrxzgCYnfV3UEtSQ+w96BmvaFA/ktAlfHVWmBJUTtwTyRyKP/1Ha/l6rKh6RkHno
h5np136x4VETbQPVU8FtLn0s2SBaZUA8RKgq31T9IXwU89ngbVZ3/Aremzr84qwb8x+5LEcbud+b
i+xHxyyz7ReCZZuPbq8dn52xcOpwv5JJe7t1UHCkU61gGBbA775xQVeglVdtQci/UDyyC3rzJqMx
u318GyidGp7zojWE5UiHwsLhFbpblzafYGNXbF5DplUTCqtDWHuRRu5Tam32p4b54QcY6m+qqKgP
EmD0Ov6iP1xDXN0a7uCKmC5dBvE2SnMhHNY59wmvMNHENwUoFXdgTb4OsG26GMfSG+KcYT4JLTZc
8xS8xDqZiul89BzVHC0EIuYxTzwjOKYTB4juI2/14L5yGmCD7xCHvHihj2w8qPtln6LvEwubsIkB
ElvNBZhrywWk3ujSAFajwqTmi0FVnQLjXnnxX0Y4ZJ+fGgBZO+a29Vbtc1bSqEZIqMhmPc/wP1BM
rBPndVsgy/o0FAZzI6bzLuxvq+uXT6V5/rKuz7Q1eVkIv46hfuWl8tq8CeBZeHj8zOPv8SwAfPB6
9fUTInPnZRZ20WlM5n2fOPt0nOPibxM25W/l7Um1ZgLd3K0bOai/oEtVgKwp7R/zQn/PrI2uO3Ny
FYkmpti5bSFj/WtfzI8y3RsPLqsokTPAqoGncpSt671S+telxldTbBJ34TyqnIjiyHGTZkruGchg
zwE9RpPCD5oCDDp2eR54ZVhQ6pKXLXRNSb9pShmLKeXYIPQkl/RRy+pXlpc7rVtSi8mdzB+utBI9
0gnel/cbYdDscZQRpJc0yN5UGq0iE27+yzrnotohXhKxtVAIhLcwd3JewE2q3oA7lss+nKxYycD8
G6Tx5DrMsyWUubzPeW5mKS26hj0sKao5Z68Mwlh++OfOyQkNnsw4zRNwU7gjO3BCXkprft/P5UGt
9fmtatU5yrIPpkDpuIyV7OMdJ10g3lZrZU/5ForAgCcxDVbnb4H0DISLJ2g7WICGvXMKyrrRLn7p
18HjZkOeBvENvvLCZqBoEWwnVyLEOBAbhrt2/KhGh9dadM8YxGDg64LOz8v2LlFn05IXxiet6car
Nq++kUYl/0J+FQuM9ENzL1dxtV4F8f2Rzi00fIDJ/gIm1CdqIN2XCjkpzZbMV1yiikra3KTg7wu8
XMwwZsE6HLA6WPf7a2vcT6qI29ZFw/96zDIGk8uxsO7j4hywIxKU2rRHurUhJmCAvAqqyRXnJT17
+FmE2b4XYX2e9BZ+o10SKsxfxhhuR7aNgvnAMv8zP9s7VzNAkKTnctohwlrHdlaX+kjgI9LEPnbs
SuFvWSdc6o4oD3mpVp7BKW1bguehf138lamuWvkkSrAYIQG1NF+uAvojzW0wXDbfeVuUWKOyzS2j
bmx+FkW3vTMnnnYKzp9Fvvf8d9csPx+8Wu221suHDfYfo6t5aWfUdiJnWh3EyLdAoK/EUePziOYm
QMzquPk430bHccPluiiSjEdFkJvp5jcfO7IqMgL1T9LfBaPsNq6DMgKfIJxVc6EHHLNYG2TK79Pp
dg1hWEJ3l1UEWuBupyst/UCGYzrjNZuxDBCdvtX/2PQ4glGecNI6WCjXbUYmXxRYSRcY7mVyHzWy
K/YAWn7wj9Jng9BISvGukvngft6n9H864/kTXlIzOio+Cn6aaQepnP75vNp6bup1A/V6L+KrGKpM
Sy3ykhmTbhhWViyUuoiHSR/Wn1yqVumKLVSicb2cXB9GXPNQe5Xkb5vV+c6KID9QQPaOgTJv2Nwg
XQ+2OoRy55onY7t9hQ8rSkBV7qzpIWgSmhK/wIeX+/ihWyn5NKz1/LRsnuffH15Yt5JP3asZ1dpW
voy+ZOYk4KRxQ1zeLCSb0S4FYDvrMk4NgIzHkieLWNfVIxS/VgPiBr1bxGTenRLjhXszrF4RAwG0
OEogmvaAGjvoQrdulRdqeTt4iiCTgo5tasxlb1P3Otoleln3CnzRf44b4JCKsks6th5caHdZznbg
2Bh3i1uAKeZFCCVFaFtTpYWGd6Zx2ikvdLZIs4sU04e1QNj+M+NWjopSp9cml5hZzDZ6UX8sPs9U
IXaLrYurTXECcoN4EHqeM6yEtSu55QsGpwip0++ICrzfY5IwVFhszXKdLrAg0PQhwdZ4HrxMdZlG
jxBwlOdbtY6qTXEd0wjk3owiHXFkiuNmgvhKhB4Ta5YIc23GSS844KnxZraEq5vAE2cIhU7GGrZm
mrD5Qoi53BfacXJPKZkqZEHmEey3GKlFH90UHJtVnX3vWwVXuW8Dt0cTf7CvhdDhf+Xo6tPwBnWl
a5TQt8jaCxTwogw2z0WMpJzjVMylb1YCAr+Zubu1jyUJGPDQi6hz5nRkyxvSBXHNAEUes6dU9BwF
Awzn7Ks9GU28FXU+fdy+Al299LRIPU+Io14muaLCkzV3qTMv+EJ1V0xMG+D2CRCLtVq/BgSD2Xnx
xpBP7hoVkdohEsjirbfty0ReqsJ2PgSzY7f7qp3KZLg8ZyFU1GqwXWp5lbDXjmtCms3lpCRtwlf3
YtSrNPF0gS0shoFg0LRscvFC/u4CEB7o/0btIXieVv7lTjTaNBXN1clhVz7yQNtD5nA2Q4f0G+BA
QP95nGI/1Ji00FdOSotbIzxG80AEATbgMDCXx0d6p4NUfW+xa3HntUT4Hn1muRYShxiWKSGMgG6j
tgTdA9eAXDoZy1VbcvN+eI/O6UA9IGE51HEXkAapkOIhSAKmNlUKXGZnaHWDmNLrHsWW258VfPG4
lnlgGGseWkec0Nat7NuzHIhLIlzbu2EJX4pnhoDOJ69E2mfdr+plM0ktlz956YNy5gjU9V3qFzlk
fl8xkjldvsp1rGAxq88/7y0Oqij9EF7Y45G8yV5wTP3eZHHEZa5MikxduoWFp3xqMJAUaLL0r7uG
g+USanVOdF5pbzH1I3vqYFyzeb/dFNH2adKRhOuZZQtUH9VhKeuuX1NUXDk8kR4eBfJG2s192mCK
klsjWPVoamDL+cPL/yBudazKVIVHf/1OSvvsH4m4oAAffvkftMh+42lBoNTsgc1ly1n4I755ZNNd
6iRupO3UadVdwlr5i2VwR/KziJ1xjDCNXeWiA68w/vWuFeFfj9ur0P2Q6FnVMImszZFKaR170edo
meXH1y6j1COpryL2Ye8+069y79/xa6ICHQlU9F1RA4eQuahoXkKWUcwRUnCREVJlLd/BhzR6kHDh
fcaeUNGZ+2e/jEuYIrCGUzGmMcmmx0qaf25gev2YVv1WT4KQGaU46opGZ6mA3FK3DBLkRUlo6NCd
3Bf3DvftBK4zPbYjB8B/fcBjt3nPZ1MucnHyvQRbqGMaX7NdFxcW5p3VXDp+ux1VwoNdrPDx6qsR
NsPcdcwDpRVNJSTePW8z/8r2dhwmAWcwov2oZBNpk7hXEJZN0QtmtZZS+LmSuJMQ8Tfj9BsONnjo
KDj99BYmQEKAut0Hmy+ubU0+yuu8j1aqxoCecFEhSTTKlQO8pH/H6OIhRceoQnRxb64f3cphJiac
OL6IYMO4WlDuwB4ilGqab+9l47c/h93+ZkosbWiTKy6+aGcW4FOqwSSMjROQEokO4r4r1Y7Iu5yK
UdXldP1P9aKkM4OUTaTCKdhLecV+Q83B/izmwmAjo6gAg1wNTEnb9hCKHKFtPmSgmnywZ9Xfo4vP
AVd5DghWjxpj0hcVUeebl+mYu5ASvXcuLCOcsic5zdCKuDZR9U23Rhd4nGWpQqI/xn64A5bK6JUW
BKT1OFat+VAFpJCwy8bpUKxfcKXEAydEJnyzVn53Ng6EKvDVUp1IprAh5olQhgxxSpoqTWlSTw0K
hExTLQHJbjfp1fpqDhKAa9NZBOYbdVUUR3YZpORbGujBuGzPYiSqZuL1bMa2C/k00ZmrWK73Sv42
lJDzBAfSPer8Lk6HJoF6+deIDaV5BYiV8Eja9sgyqbMBEagAlIrNFtEdwip1iZvX9shCKcS7+ej2
UGax2YTmp8xulx3ietrXFxClZ5f95iF/la00mn6YlwKBAwjGjIoxwB3CexHMAUhasPYRSzQ5Bfnr
YHnUEUfPMCSnV0TRHXbV10PlaOE/TItnFASsl/tMAlXVHGe7bERTR7USbrsWXb7RfGow0O+xH6s0
Wn4lct/vl5jTEDnkcWoZYvkyq2gbMP1zNezI5JDoyYpOHgwah4N6/7exf0/AYjwNdcG/9CtCOeqw
mFP3Q1sTAUToFUorax/0T5Oi4PrAdg2fVc+p9XAUwXxOE2cb6OjI1cTUAePejOW3NJ7omcivx5xX
5MPmvd6ZRbd+l0F1PqpFj3AdMTeYiMHrVvjOwzByhwNpaypdwh9mRw+DFx+mK1afMaw37+PvVctp
TFvjY/htzRXyP3NMJjo3/xVLbditiWmATucowItw8miy0Ek9gM+Zs21AIU5WgQYBV6BYOeP6crYA
z3cAAFTRT3j2JtyhwGYmZ7F9onLbn+G3nPQANGm7kWU7aDOTmBZZTRCpZCKsDP6C68zepWHkbFnZ
Xnjpa8NDxghZD1PPHyqkoAYC4vVOJjh0p4cQAoPCSDYUD3FQaNp2Vzwxg81RBi62vVFsbYjqdb27
hruhHhix0WVCkd2kz65hljdmCgn6Ktm+FyLVRYSau5kpbtMsqccvkPG7n5K8qJjVKxHfO6b8YNvo
1of0/HQkOocSIFVeQZizqBQ1nl5/Oa/ojoG/8ef0nX7vlazFEBQbPoCKrhzYyUFig3Yt/jnfR283
MeOwSt2+ClC4UuNYPGwhK24s+R+nAfFerYsVyZMXAY/WF32rk5SMZ2KfS0vLQCG1MdTgKvWYaJkl
9xPpJF9JxbyQ4RSy9w6eAhX1mzunenC/EDjXdGcFbhDDM7KOWYnPbQiGc8iywSv62u1ahPvyt/LI
CxQaw6hWY8G0tZfVI3RwIW/IsJcuoD+A9XL/eo3fVB9FNtNnxHSr+grFdxwXjiHpm3fm/p1P7jZ1
rFmTiJUiHp6F7w4T8I7yp46Rg6wWqlsWNvNXHcl6hb/5zqWQSzQ8Pd9HNoH3sUFt+dZjYOAr9+zt
UQ4k5nN+Sw+HLmg/SVQ0qC4aqb20EZWHRRT5G2XEkJsNhTAWeoEuZE6YPFqGICMICvfT/IHyLseD
MvPGeQPro00YWYWp6Dd6JBROHLQE7CWWOFriIGaJ757cXjueiIj8Yy13k6APhYVa2EPiOhKL00YK
GHtRhBpZkK5IVVl33gCC1W57o8k6no54wXXXsUcPZ7V8O+8J7ZQQgJJotsu2+kc58aDWMutIGdyQ
uIBOXMMqal+OSM5bDtik6m5EPc8283Tp1b54OAWE7FGiqkUcK8oWw4PB0BfUHoZ+SOb7qmzT6bWO
KzWNqjZLkuGyDJTm5v3WleTV62+FCGJQ9ozYyMAzUwJsAKDaMfpKFGlDCq2o9thDxI8hq3/HmMFw
7sP0UGuJrtdSAx3Jsixs3eQSStJ3pSow9odwa2PT+ieboPJiIUi5qGXuUlosyyoMB0ahJSfk+4nF
h8Qx6VWaHr0JD6BxLb5RCueFRtJGneCuYwKqddgzLNfoh8FQw5jeXAwqNO+pFnq1kpIBa4gTI9bV
2ucJo+6CGcHArqg05QocvxZJStJMjH9M9TEjqkaKKJSvr8hQGOS9oxPfZG+StrumfiKlxFyDNco/
2fFx7NpwFl8DXwojgKyzubHuggtxzYMddcn3jJYXPihYdL5dmThQ8kpd61YIpJv7wKttOdwObpWh
RB00qFHfVIPjSvkaoS3bvoJm+x+LT1ylN4NuxI85PxYHMDVf5Wf3vtt8smFRUYGXCCGztJ2E9rNr
N+M6JSyvVqKttiRtGcRtB3ga5R2oqxOVO6hQUPp7Kea6dcxdSzX1a6Bx4bY/DJURIjREXxqKneZ0
gX/mZnctmZ30egZZIKgUtrt24/EtHz76MdKHxVwCUtPy8A4uLYkL/Zml8dfJXNdMkjVjkNMhhYUb
I6rfb08yLepMQuuAJqiVUPmbJXGqL2HU9yT8whhTTDOxKIaWutCGOJp/UB8S/3RwHPGe2R3fi15B
v5ZJjvjBqREmQFQepzFApJVadqKKEwh7OFnTLU515XdzcKJd2+VHX6txQEf6OgB3qUYWlYhAZhft
AtfRgkbZO4uQnJzlxr+bTaUQOandZ5r9fMfw4tkaiWqiP+bEouQzZUxaNpzPGdYy3Kn9cl0oy364
PsjDK4kS1l7oBChqXc4hUnDXiaKFWAdH1Z76uOS3iXvkbBR55JY8ytX1WTtYnpmBdWNiNmtOQW5h
YOXBETLlEXZKUqDOSrB9tCrqjAZSqFUlZj9JquOtDhvUzcTSedAhLDWxjjomYaoCBFySmTAnuvnQ
cFM24NuAzHHv8KTaljhIVsVgaHSxhe6bzw57+FO1iHtfflgDxGNUQhUnnpfevq8ymPdcRJkwQOd8
SNOGIU7pfPLELz98YC7jd5D4JvmkFZU6UWVPXrbI5FaDlV0f+WHRsNKsTBI5DEV0v3IhJ5qGfZRH
FhmfECHu1EvdW/qTRVU/iEdYgxgJUcRW6slu+cChlD9GgRqpL2se9smuQdU4RoFvvS3ixCrpmx2E
dDfunaCoutfgThuanSw23H8DVCXxxXdys+xS5KiStqAv1uo7o7PFUJnB0W8waupaFl1rqVmHpxlR
XObHfz5Ukk9blj3SBlhMUvu0ujxPsDrLo4Jv0eyjXTHa97K2uZ1KFQSvlRQjaCo0lROi/K4jtR43
2RGG3wjSqkEmw+iq1AdQJSDTGi8+aoUaWpkrwEn8eItU4VQXp9r1KWI4HGMq9Loz6IzqX6iUZSJH
wJc1TpwW718uWQ9WssIN18IxG9B50NhQsrVPugSSak66nQXkaz/jz2Mdj6zKnwNBbLDdzl1Jw2Bw
ZvsUrW3Zaz5jl1o6US68v70GynmrRijhoILd4EnDXsqsv9ob7uQnO2NgJqS8BCQzg4dLwYQr3uuR
/N7l9pasqWtMAFqPvhQMZObwcnhxyDoCKMijc8uP+vAzK1BASjWuqd48ICQsgJRZcZ6V56EYw/jJ
WsUQGgujQv+3joNc/aeMmFS5iF7wM8CPAyo+uofDyV5KiRsUYj1wbZ8rwnZjq4TPfNVxPlOLu6PW
nPKOBZvpNTNuNtt86cBdJ3NIkFH2F8jRTBLoF8R6/lE5vbykrVAyVraLOTpx2ieFXIlKVtTsTfKs
vUJnm14OlehwjaYClmHA1PH+JjJ9+aBq0WPxqVJCtZBx1q867qyZQ48GQJm68FdqxlOnEQFrc/df
oZAXGHSkDJnSaZ6f0ouLlA3nIupnJb24K6LNMXejXKnNLsDZn/t3Zy7pc02x+fPU3wGzr4nd1y5y
zFAFQUHb0SamvfP7026VvZvunNcmnouVlIaF5iInFR6LSU59c4lY+QbGcRqGs0jj308CS2lb6Emm
cNUEdXDHPj2cEYZzcDyi/1QG9Fie/Ax/4JOdw9E5cDni6uzirDfpR4fPqvFuaT5NB9syxjFAuEBo
e+Fq1sqQpAWVCbIHeio8ihQyUBBfRumgOtV6MXAdTsf2JxtqKYk9TdMzgFqyltsf3N2TUxH8wbXd
HShkm4DT/A4nr+M+szF+4G2s3BM93LKmKrJ6LrmlU7aus+xcxF+lWv4IRINv+JO80P3aLpymBu37
VciKYx5eauhSdLOShFqq3VjoJNbEL2sMwLZRhkS5j2F0/2edWSHxJTzpf2VtC1Gm8Rim4bNf2S8J
gZHizcfvjfw3gOKcLLhDKQ0+g1RZzG4PQF1UQBGpk8L19qdZM+H4vKT9X1yM7L+2qZpQmBCzbrLb
EOhfClUR5AZk1Qj7Z8bTqGS8vJJ8gApgF19Ka+MB1DWh/QdsvavtrWL6vzGd2hWbzGuLofKPs+kK
SPBuTUIz/T6d++9xyE6Zx7bcfq7ALcSvy6X/MrJdiQZqUafRReYhX/oXI20Utfzrth8h6vjWUMQ4
W36lfZtDoXw/FhjCeZioAKfG6JZdeGFI/DQsGDyhI++5ZEhUg4N1T1VJy9RmyMf/LgYYxpRT61bM
yCdyxiayiYuqujoFf4OY4ViG77qn+IneAtDQyWtug5dgehs0grh7wdxiFUr8U/gGQH4GRsOu2jZc
CnPHw/UWXRYmBk1I3LKnqmcvtmYq+ZN6FxLGDj2pE/hrdMF7J8i3DqAnTbQTKiEYr9VBVFr8pbZO
SWWnnzMbODuLLaiH/sO+Udmn+ATa7nCbZuhz20KuV9atOlmVIGEbBjmLhKhWgDWnj3hQUQy4Vl+H
mn9NNxJXoL1iQEswsiXej0CcXKBJkw/TwG1RCaTrTZj0DLJKrUAnEQy5GBFWie5Y4CvguPlW2MAb
zxd1vo8ZQSFUeSuMI84i/BQcC/2JgnPzGTe8+TTFI5B8dsEMnnlLwgcPt+JCCSoUVq4JmTSm1Klp
mZp1yIqwuTjDhndJ9NCQCWzZRB/+KlejXaj0n8tbNksMQ4BUdpWjUd8iPyJk6nBn+yfxOKU4LlTQ
fe0FjdHUIeGXWTetGXFnKwuQp34X5EFK5e+fhs5yQZBqtaeX/h0ofMeUpaWEsqr5xCX+cF0eniEN
INZUXdeVFYmV7EgS6ggMtLtFuxdHiK3gGUvezNLKktZpSHJZXBIps/gI5RRbyGPtdJFMwOFFm+Sn
o9G08FSXyHUFor3ChKi3IoYLYzvfCNR52j8ow5FvkfHT/35m1K+R6JQjZzZbpBkQQ5lyLB3XzENn
NKYUjxJl9BO26RCtcL0YqOSAobmCfWSRdO9HnilmMLyQWL2VXFcNn/FVuXSGRxZfYKbV7htl3f1f
djmUCr8DDMMQcgfVRMmiBNKKJFrvyulCspjGES2TPfKV6flXwZTg8YIElWveNFuJgJ6G2js6K/MN
n5JuKbS2jyYjyh8dbMoG/mkYoVYbHJWA9LKQyrJ544ywVCGljdbXYcJlkWj0as07nvsXpsi0jElH
uJYlDdb7QY5vFNxAXKWu5YfZC+liCvgYohYPfUarwXg6CTM625EtDv5BBMvYz4wG/ls+X3RhxtKl
dS5j1Rjp1TLls+mLSnJdAxfYX8srOWrMKur7x9PA2HLxpdU33LDJ81AvfyLD/WvKetXsxBNfeM7q
HaO3U1n+pM+ms6Ke4AkGQ9KiVGIvyOkLl0UIbukH825mvCLGOU/i3Y0Y96gLTuqG0odyTx2ROYkn
VNCRpB7bWFjvhlcINKrPXjlb9NyvGrvV7geeKDM/R1LyuJoOWkUVryXm641LY+WAoWaLI+Uyo+Et
0O8JBTcqOteGiGUBlEP01u0oFCObp5sre+TPzt5CQZvpWaFeo7hmNH5Q3b9ibADTKHFXugGbVPmg
DLwqcQtghL1ABpV0nDqHJmL3i7padVAqHofD+AlDxVnJuefHNYzZsBwEyCW3i6b6xJyQ4OwczEx5
XdCN6DJ87b/foVlXbl9dHF0gvKiO7kPdKaWqHd9mmhAXxWKYK4aaAmdLLJ5Rsdq8blcgXIMK6vJd
M78EP+d8meFGhkN9j6LbocAi0tBV2xWy+xPjgAHJf0iMr3zaA6LN4b2wygCXdvLRSswRoTJQS+CE
YJ81++Ung1ZFnUDhbtO5LI6Yd6d5h9Uee9yzJwSy5WeFEuLZIa4aNODpUNschqpmnuD09t5BFyG/
bH4z/FCwAHja5//2v4iTqLJN71bCh7EqiQIT5WZqpcUo7UlxsEx6Gxxf425DDGNOfLWu1emYOt9J
dCNCRgMSVeBP/9+UjC/8TxE3zEilbS+r1DfwyDyqtQGAc+JpHEUsVC4HT0b/g9bbQpobsCVQtNzd
eQ9qXG3q0y8fh1akbXQL71Amarpk0CA/rqqi7z1DRDOa2MXeu5/yX8D0Er26W1XqQ5C04EnB4UKj
gLWweDrkiUV/C50PQEqMK+5j6C9iPNZoFoQnXHUqcSa0ZBPgPPzMP7vMW6pvFRYYsxvyhB2p6yoj
Ng3GZj+By/JTKV9h2Dv9+iWt0M7K+kqmRjYCwrEUr5R8P9UI09aam12jMaOSInqMh3UrIM2i0n54
LTcbjpYvK/6Js1RJTnVEh413c0pXuKqltjWLoINUxp3ZeBVphfvg1oPIX8a+79fUG1ncF9v0A0F+
wTPm9w2byO87mYaSTqoRhOVF8yHpqotkeDsltdu49TjJ6Ci4Uy+6n6VmsXHBOpiuBp7EU4Cmx5yM
p21HnSFl1QgtmR60DumYDNejZFpEywXOUQaKWX7DBk277rAx8mFRKAyyEFzQhfsdUGPstKUlCmxZ
fp8/VmkImjMVZob0G3yX87hGqPJu4ERPQxrwBUX5QQk9KbIjoxyNZRb0cL8DA4uZ0nRkgoMn4en3
b+kUNm1M0ISVrWKsRdQ4p7YJ6x0vFOJfn3tjLAzeUKRL0O+RuPRJtkdRp2EnRBfNqX0Hn/SwvgYK
W5XaLnDItN2/c9H6mlzFnMfwmgz5Out7N/TSHZj4ufeEDctD+wklYezI5vzCGmdsGO4ecVdkjrVW
8hMcaO+9y0AedlmZuT9CjExx3U6JGZCUklhzQB20937TPW6zzsvqbksEz53dayOruOhd5jgLprUl
0NushpbNtISC4fD66ifxCxZOvH/h2DeTw4BXPAqlb9X49FdE5yPQZzegDapgdKuiIHdm1Yb2o/Q1
2VzndhNXgIAllKpVbrEEFRy4ikeeJwBozQSEenDMoCOKtT8oDIKk1Byl/aChSxm6BtQF+vYAYz3W
BM/eCZ070iGwjtaqjgFXcvUGk5QtWvNgcAOmYT4VB4IBWnFWcy1AcMfi0UpMJOpC4pnrk7uSIUbe
qnyglLSRCod2bI5wzRVTOUl04QXgatwKML4wjqwgBM0pwxa+D0EfLt6hQij/0AeZxjninEnNIn3K
saHk93d3bFJHxFZFt/WbPZxjtGJEKndRodFXoERQdjRbNxfZXeM9KGsGakGaK0bl0yUC3ojyYx2v
goiP4M3YudF+H5xkNiV7f9eiXMfDbgP3deCChEdX9Z2GUoQsuGaDaNXZFIIl7i8j1sMBWSJ9eXSS
lnfFlHvE10EwqFy7T4yVHZEue6KsGaCY1vFfYraaEUumOCW9rUUbCXgZkZTL0cvWiEXQoHEK/h1h
zSllZGzgcVpTWNmPTu/XChgqc3mcI80e1dtGFNstSDnyhvlDO8pSDASjqifxKPOJKCy0wkvXFbiF
dzlREiG9h+Vf28ciozvlx9VlD/E9Nmjlcaz83VMnBuNiOizD/774/10LzyE9j6BWzm/taJgMy6pj
3lJqs+DfHjrjEJtoh3ctfLh/IKMI2b+Kdc2vQICZQ92ZvVKu6XB2oEOiw16tvrzP9XfX6YUfjOtX
IMXH2As7oELVaMxi2K99QiqmG4V7htDEbecrzfb3HUZh/VieRjX5pYLIdO1pyGS8/WMctDfQsQqF
14oUcwVztQsKeC0LnjPu7IN/bJQZaF5Xi5SIFAFzYeo7PVP6OeKb+GawOtP2qr2kx1mswNTL7mWd
stgW9rMPp22R15l3mdmKH8m+1JdZkIl8ac8hKadsK+7Z3rL2DP2pamIlpoS6cp6oDVLjaUWx7sXm
OTmimSxdWmSR3KUMOgsQVyHPYT55b3W0ot5FQ02UrX523r2z50go25Kp/yU1xt5nfUs/SB2qnAsP
NjChfjz4EouCXqFYRBMi3lHOT14jqLp3UELMxM0dQtjIHeua/bNV09jAOuNrUeQVw6VracwUw9Pr
Yqjo87Cq1UfpcJkCU5mpLYi8oKS2h7kCEoT8E0JGUyTSqWEg6OCYhVUiygh3IPY9MF1yaTsTj79W
OW+SzNxG1SrHm2fOyaTqF48KNocdLIVT/DHkDSUfwZ/KfAL6EKenlS007L0/tae8MOaJnsEfbrDa
cWiNkk43RIaPPEoP4Bu/UMHcS4H+pwiVmxT3kUuqQzeSLtTUWeBOEmEKKOgjtDGaWV6tF1sjnSAs
rZkpIS8EW1G1IvrPvuYo3B+6IwC81AiZz4xfQLjWMcH+xUJZ99bbL3Fwgumo1vozLV7rjtkcOEgN
NnLaPJU01yOszEcQeNQfCveFEco/cwy5os6I1HFVBkUWHLWm0Eq2ucb4aJOWjQQ7UXQ/FyILG5dC
2DtS8+SQudE7Q/84q/KFOCS3tNjjoY3xDhBPgMUzhQ0LdTw8xoGlP1yDMpzhbviLzkR6iFubi5Ti
+30tVKAjzEcRE6LfIrIgtdv4nJpt5lwwsH8VU23OKndGQiuBuUTfw4tZiW+oOnoNRQCebUxCwBzP
wBGJPVMST7ji8i4QgjcgSy35QH2lA/gvzE0ylf1A0tpcZ84+vwBG5qDm8byOKmmekZlR75aus1mV
dObe6zYksNUNJVGwbyG+UfCCOVeUcBLAcze9Ui9sJs9yG+l/flcbdwx7M8rSZ8jXvPt7spAOqS9b
KahEGcthvKGniEiUUjgYvQjdHZsXwTmjZ0yYaL6gKJ4CP9HO1JOii084Jni26Llj3dtMaF7fqtFi
50unYovHVh6ViPTNSjiYaBjj3Y+MF+cIkXe2QqrdG0Ju6aGHEsH9II/0Whs32cVU2O82mlbq8b2f
5saWvqnfxme2cBxzGvlK/UMfbjuSGYVQAVrat3ya7HmXiE3bNcPulj7lKd+F170tJjtRHQXblIow
6iWB7Io6V70fLxRouLPeaZGn6Vd7XnfW38mbt86262sATo8c9mew6yWtnS94vWIjfP7fp46Cl4I4
8VRya44IjPScf9mGV0xRehSKyNc5CcDcujJ+FcjYiP19WIFxEWPB0jtLKSKq1d5+5efK611uvfIn
fjJI1wh/UqBrnhkrNhOR/t+r62IayyTiewrO5/YlX9g5o8JJccAFEeJOMHTFwDUDutQSedyYpAGA
toPdX5rFiSsG1HlsiUyuEN8ntKQXnm7NBsXkHl3EdwBEEyBuWVRTid1EMVm8TORvO3hhvV+IOmwj
rVZzD3XuAmJ7MK+reXVSe/1nOUIvtovl6ZwKKrm1KbrnVMoK1IIy6zk5Ds6KZ4132iQwJxsB1A++
Tlx/LdedlfqyWThp4BiBO2Bbzh1bi/DQFWEf0dZLCYGAUQUSRjGLFB7b/esmuKey9+bM4Q/GsIXz
QNN55v8pnEOsB2FNgi4EQFYES67GPYNiGRXiYO6a5X37X/bi4/oKOFwhXanXM9zX95eteOX1z2Iz
JOcDAEeFZ7WjVBMBMuBKB0x+IW+t5QnN6Vi3xs/6JGMo5lzOP2qoCWzupy4/t943pjD58zL7QRvv
p2KQLKmEy2NifvsKH4VgEOHom1UcIEsNzvO3MiV92zf0FP6D8mKfnbayZiMZJQO8+7O6Wu+ldoqd
SylqeazbVIOdYX3VQPgdUrmgRz5kxOAR2FtaLiFwnBXG9CFhN78wdnZ6hNzyt3sdWR5Mgsud4Av4
7Q8haIXKjfqdeF+NzS36jdPGwna+yXOTDbf32ji0xmWTGU9slmRglpWVvnmWckXh9Obl4xhhi7gp
+WGItiYNvWKMR9ng3QGXz0EvYiPShp+7Yq2Gn36hsFPOHpc1bix17Tp3H4BSSCWrNHQp1xTUQfj0
5jdF5uCho22YLDphqxvPQtXTHE6FTJxDasX6itp2C6dgKzpTu803dhQumf/5FwMTRV2RcOkvWv1W
BxbfwcfckGwVUPtMy95QHE7yyKeofEZiCrS9FkGFl9tu4NNr7djlMBAqwp42Usu/zIhVrmDQqyU3
c3uEtAnPgUyLbfZfSNhIeoHqe+DZH0nAqMQNnRHSLhfg6Z35hrkIPrx6sQgk56K8Iai9SX7JKylC
hBZiu1QvOZGWem9bRZllVUslPFI2Jnt9lKn4ZjJwvxqNnSQlmv5wbpnesVXIPtaSUwEp2YYH0rWs
FqXSCWsJyhksRNvGvPCncm/CeAIVtetUdwZ5QT2WR7VmIARQYYi/ASKBVAGSDCEz7YOfzbf8xm2D
mgm8pdpM/pqc7D/6UYvOZFkSWtS8DO5ukikjKFqnW0KmtFSNAVGNmOmbQabt9Vd7CZjH58W3U0VC
UqKAUsl2DkyEZfjmM2hlnQZp6i1oCyRuNxU5b3yx81rU8NxzCaIlAQ30LBVNBd+FWcq7E/mvk/Wu
wKCY2gsDvCiih8+K4pwSd3MhwZTATr0TP5hYcLh9dAMNZrp/sq098WYswLQmJVBvYacKL3OelOF9
WuhTxIjqy6lYgErRaWpPRJdcUeTHMzeW+cJwynGhoJsmPbkC6t/HHEMhVgInCg1C1OoAj0H3mD3o
1lErLfWszyPx/OkU6dh0maal5mE5oFcAN0CKhfa+hRxUjCoXdOBPXhmC3NQx1BLStvPpCn0Kr5+n
qOpyMIyBmU87h0W0FoUK+QDVAoflbl0opabUhIFNXJ9AqtcQoDZaTCudpJY7HKSnkmLbX4di2OT9
bxKf8X1iAXYM2eZ0LHkzpAQZEHzC4Kp/iMPEjmM3Sp2T7qwVKa3TZYqq6MkzyLVWU8wYbqni77kU
dYULlvZcs0otPLMmZb81p65RfpFnUoKBM7j7r2Y9t8sO4jXAxKZ4FiLgLA8K0a23Jf4zIj9i/Wst
1L6nU6P3GV2A+z2Qbj+xVh2U60j9hSND+KOPlpS11tqckUIm2mAkPjNlMmmiBLghi/e92bE8SjV9
qpFGdUjI5HXNvR+cpvXuiM651pyQeGD6xCrXQaWRuwIAvdGB4vn1QQalCUPPbIxJWf1BvaTPLxD8
d+4Ibta970F5mYwRkdqGtdQ7HOBObhKUnCLi4gv0Ha65c7fS+66/6esn4hRukbeVfl3SOWfRoBTG
5dcOC8llGl7zHX/qQi8uEieVV701cxPZ0tsIR3sPrzXYcJWOEAGeUjmPWo0INZZKmGMi5ZY9o+EB
qkQss+9lkPAov3OWv7CWabZPKsUaXww3cyXXa7C9599pKqSPmujzLYnTPqq5X7jHlwRY1gL1kJOE
6fHfEQ/XPPQbmkMxkL8owJRymYhj8KrnkYGPlQn1JA91YIFfAFBIe/4aBO77V6TjjiCKC73rtM7+
P41Jz4SaNQeShA0JnWiWBe2Z45iFYYceCSsjUaKUPPFFiUtOJkJHF/UgR3Q2xy9QhnWzdkaVcQ9n
4reepmVb3jDCSiEXVcIlCDqVTYWnZyo+XQ6scTjzWCateoD8yMFwfETrKxNn1fkpq4Jw50BQhnN7
q1cd3m1XgEJEVsn5ALvIOtXFzOKbyabjw4BjOKP4aMu7ig+j4UKIU+HvTfWQ5x9JfRnpSTfEspsP
Bjo82zjNQwPq+0pHvBI9qIAp0aFFz6LE5SF/wS0iW2uufQ+G9LSrVuN/xWz8Td1IzAtmKSDg9UEj
ssFpHuy4xq21QGE5UNVRcR1kJPEKjJhEiFr70eDxy8Ycmi+AuwhJo3GQv3EpV6W5fORLkjmuFVvh
X7dNTPady8h7UOlLdLyO+DZNmmYUlJy6cMPWjJDASS7DUzVGIhq9/Bh+Ql2kKz7lPbERwCiAHgBS
bVmU61EDV8PUQ+ggI6Ay0AuFZQ/d7bnvwJKnq5nGPluBr4djbza+aGVEQVG4j+B5t0/Ib+sNabvJ
3LRrano8qUVLC8QSEtU1+i6a8ar/Vkz2ICtLg/jAaxp7VxlVRs7xZgyCQqnSQuWb0FcISaz/5e8Q
+VkBax3NZYdiave5ZIxmXS4PmdTHo1sZT7JOX+RAVPjef922lje8hSM6O/81xT3PZaIVazZ4vXL1
maBTTWWj/SKMNq0aff1fuktREPgBfaIaQyUY8aHT8UcGBLgi+1xn7Ca/79zdDGUl6KQw5vy2mAr9
uMvFh4EsE+4wjnOiJL0hojq3T5WNr/wx/Ow2jXJfCQCBrr17DzhJBY6J9LvXOSwaTFTsLDhPHKgm
UJrgFp1ZLhnWbQW5D22nQ5zmQzhY2GWHCw2I5FHOTpvrngRfWJGoZsjdMGJTfLPpBbnVzlxdiHBk
zcR7tdOhKAhaXezRp4R9KGYQsF6PRhrCW8DU0a7BiH5lJW0JgHHBrvq75WyqBL2m3cJQoPIQ9zWQ
3YJTnigEyegv8yePi6QwE7O0DaxfNeMmv1CRV0DrFBGAIe2KqmAu24dSjg2maPcp48qZ+f0FQY88
OCxNIpK3iwJXEloYzLyvFgCqSQwNGMVmPci7x4DUAaeTf0TYjKPuImzFytKyVZHOriFjp5cq2F0q
SQldocgx18uOLX6kxqqdoURxdDhWYiMyUpL38KoDA/AUQdosmQ0Aj2yst9ZfztwZcXN4xwTJeFnZ
9X0Jdv7sPES4YXEQaNO6eBkBYm12rvP15trM2CuIOV5MgiaNxCc4fyBY6xLd4fQgNC42/PrXr6zU
3UxsMD/ipLdbaAfr4F69HM6YrrOXUiKbSPQBuxk6hhl6pP4uhGfb+SuZgms2xVJMHE/RaHD+gYvy
gJJgx4sjLEo0sooTLUvWpAxgZA3n8CQhW3/pfl7v13/IjluB8KC+GeVOAUerU5lokOI9fANFiL2W
s5hGzMJCcwr9+pGik4IJo77XEKOcZiau+M+IfnVT/Dg+9HCIXiEhqwtBmbepMeuMUQZ7SxWUpGV7
NY4rLw316D5cDjJYe9457xHvrpOxjv6seyAwshG6kNQlZQcxEzoMlifyy1IOybuiiWransBBMNtl
iTyHpqAyS+NSiueO9SeA5B2gd9bh7qoMzEwDluoIATQagVnAd39KpSf5+Z5UabJ8TRtiz7Fvdm0f
JJ9Z2F7BCQvoaBYw0hsgxYa+Mvagi8GrBPFFzGfj4hL5WSH5nZ557CyxT9KxjAQ8N1XzTmLRUU6e
sGW4G3qcTtouoeILIE2XR6MZwScanYIrUuugAUFVFhxko32JNojdcVuqejPkS01A37+4aBz8/t6q
PJiJ1g6zWDPed80fnIQWzjSY5qkVktYlYaFUbw9sZUtBtue6JLrRl/HkHBSe3UQqFatoOjEfata5
qJj8Zoj2bHDqv2Oc8NArdYXGB3N2zq8IX2vb9oYkurfk8Eigok1qjfIAsQvVKjRKsa3QauDD2vx1
iojOXVC2U3ihlAqvWisIcnEXl6lgYjyN4blwywvnN4DuSbWZxbBImIDRANc5/rvGBYlHVMSNhT4e
bC+31BfhzNxyWKAET7FaMBbat5aJsDDS72zxq2vsoFBA3UMVhhAoJWn1oFXjKIQzIOYdeWn6ecJc
G7VFqh0QYUmPOls3A0AxI7SvreTg/ChIiKFcCbDXSdp6vFpx5eNZLSKXdgL0ntEf7MWavrJGjfzC
yHR+hifgqIdWyFW0AKFnMq3UrS+3hYiKSbz8bQN+HfdqvFAmgD3f+p+eNm0Q4MbweIjztLR5G3Ym
sEjJFurn0r43Xssjx9CqCrs6EseJSwyljFTTu2jS395PySyYKcwlrAjQTV+w4GfE3FqK0XFqutKP
x+eBsixhd8YcZb/K7n8ev22B7z6UZYAqeC76SKz/brjZmLzGTzw3rfTqN5x/WJWmlja2NoBIyGN9
JkuruLKMbz6WcORA11Hc1RIR99Lb1dRfzq3lyYfJ0kvPAVLU8iW6RhB0KimuolYG/GXiQ686oA4j
bwvaScyGT/GJNn/LoZBK0JwxwAqmuugoDff0c52ryLRpAqROm5jJJbmt9DhLCs4/u2p+2bEmxpjm
IpB2rYYezaYgyRJCvWh9BzNAI63PUpMb50Th+oHSt7itIWe79O0ETqMx6AkTRi/l9ChRqwRydtcV
Rhix9UbkSojdOaYXX14LTFksmNs3Afx/5vWce2bFick7dgJ30f9+SSKewCFjN6nR5zZo8SrfdktO
jVwjbjqTcwlDxPq7nSsiNa0TPbnit1P2uqPN6dX+BWehWHpoXMb87V6FbtiPkMUhRKfToZ4aeVch
3es46czerAvx0oP4k7A1SD+sT69mFLgck9p6EanFMCrcVsTYUDfOzJoj3k9+8J/CuMgSZ8Hz8x5O
w/zcViU0EqufA0OogtOXg7ZOnBqEzWYOZVo/1iY+cTYguwvvCAPPj9JAw9RsURK74gd0ZSBo23nX
Qzxa5k4g4Kh1ubfrfdDkXLjo+oAHA7juCkc5dMqeEHWNI9BmvbZFcWY5YKUJ5nHFAS5/RYAgN5hZ
2Tbj4so83IJmgsIXxn5A2kepdLqjlCRnCHh13+ZGb5St21BWIPxGlS420tizBgyt41p7VG11dhQt
xk8aMeUuet1Ev3Cof78qcKB1/LW3Jdj9raFxqNPHoEV7+g3Xb8HXVJ5u80qnG3NcEwepydDwHLVC
q0BlFbTOO1eHnMKdNLTLoOO+cCK7ai+HkGNga8ceQcJAz/soNKoIhDyNGnxqkGzdYdj+XJ4hdcCW
0XyGj5J3AwNoUWr0O+lExV7vNamIKwf+uD8lI7+C42a9SXWuyR/tfvZCgz+bexQCI7HjRA07lGNW
RQNPXLjHzdZeWuojxbLDCmJAFkDmsMexoTaYF82HNwTC/N5cuons9bIkhX7T68xTn1w3iR6ndPpq
NRpitrlbe5DgoIVqjazwyZpfFHeiXAldMwXK1ibIixWhL0lw9y4H55V3eoRX672Wxf57ZXFvcuXt
IpKWUCAHW2MShrDG3zhYaRIacZUcHI5wMpYjliroJOSmTY82DrUMtLos9iEwEsSmrKYUMFwU8Q87
HvKRKbULc69AcMgWiztfBo3V6ApGmJkn/OtfDu0KM4cT3upAAoJqYSdcqCy2IG3c7vDtnScm5oqc
ryiMGQbZhpaDeic2kfDoq87IiuMpehb269IjNhuZQfI+qpBgzLlEeDzSRMvslO5gG0Dnbq41bXdO
TN9wQeGhmq9ek4ic9O0FBDN/zcB2AlPUzoM80UQdBYnHKzc9qcF1GLBDz9KDIs8mWmhl0lEj7o7C
4CxTXhPH6fa3DKx0Bklq3v4UOxpSkA4DUSduMyuo9rWP1+Mfu43VI2sdZ+TiMKhiH8FYmAbS6kQP
RPnHRErYYvSJ/DQO69Z9mlWUPB/xwlQxMYCgJwZoxUkWj5hPsKcOYGfcPNakdlC/NhU/YFW5cR7r
zV4cu+hzuzJhmxgYHjZ8LyNRL/0mqJ2p6rzwH+HqJvQqmKXJmY9EUa/GamWohQN78DLRmh0hz6GC
BaTyQRr1vZxzHfpajr106ETCCZLRW5rWmF+/OAij3gys3KtIn6pk/JpY0qZySnS6s9H5yX9Zvvw8
KkoaAM6lmN88DWvDLwFjImyEOl1d+VGVAoBvxthv3ZTH+yQ+vPi97bBXNAUsCiI8IogmW9/DU9fm
wQHBURK7goI5rhkNVcYRDgYfVwdb3aqTo2fE90heIA57Lp7I/DsJh3ayFURcrcdlu9UmSyyld89Q
VLe4ukJ92/9/9pY/jpBd9O7bexEwHbOfN7YwgWtUCb5kKxVq1S3FKU2ZyTlhbhoM65McoDm0X87k
7PJLyPfZgsdkky3wibUd/7TOiZ/ZhVQhRemHJORi2HO6gVtFPlyRbbGzh1jXQefHOJSpWIK5t5l+
hkNF/Zfj9YLPHrdc/yy3Lzjo03gGZkxnAeFD27fjn+qSXs8e9wXqV00VH4VrGpehmVD2kD3KcmxD
Nwp47CcuzeT9BUWJVWm6JhgYQwKCDGsKA00ufkUrQODIvsKCCteXGSklQl7+3nf6AiF7iz4P3LjM
0tEbUD5nL+jBFCIpsJQvLATsIKkelYNmIlzDnBdJRly9QiGHHbCqmFeaQsOS37AZjnd6DovyuqvO
iu4ZZcjGsftW7BULTXTIaMM8TnAi5YfZmtADPq7fHss6shb5wImKZFEn3ennHsFHpvYClmRFAO9/
3dwp5aLSxsbqZe0jTzcgKZVu0fsk5iqQOS3Khi1/aPL1oKkMhHd8uG4reTf1mvpkrfH8wj1RlXXk
CwSWMl3TII/wmg2Y/nPHa8y8/tR419nu1r25I1eDcVfikykSWtprqL9BxJIGN9w8agcZyzTM2l1C
EjNyrFDwPKdYHARzb6CcFpgOjE/L89iVXWVVGKUjKQKXA/Zu99S/uyoveS4d/chmxjTxMqICgEbv
Es9FCV8w37wlKgV6BZSnzEP4d6ggbpHCrHde1cE76eSjyx57wB0O90aUisNZr/gG9YGCQTVK4/rA
Yf9x2AMaavkaoEWVYvE9CndNjYg4kGEfpw6vQ5SE82vkXUs0M1kWpLiF2DdFRxuy6aXVMDIytSR5
2AE7G4LA8ja5T54l1tO1KI3onCNInQc72HeyPMQjlnErvflnk2ykMPQ3VgP/ochdorTZ7mbDO6WI
VjrbobalVhqhdvAgpjp6966v4bj8tGor/v09sNuceSHU1J657ZzM3jSLiNN17NNaVwO3HkdeZfvA
jGcA28bfZw1jQXEEFkgvbCL04F1iIcRCoxeilWQZ2D/sij67cTjUmXbpsB7VhXLuof6Wsei93VjT
ymdva2OO+QJ13q2Xi63YtPgEQW5T77P+LfdezNrwNTAXqqVpYikTzVvY4SDobu9NK4oVUwtqTHsc
Ejuruywimd1xFb1JJWd5YzTeVkdeTUAFA/+Uz23qmdKBvLKkdx1t3T9Yc8grGsrVbwgz06XZ/hjh
Bocwdlcde7SQbywmMbbcVLGi50oRpdKxLqabjCFa3q+wFIs+aR+2TzxxhfK41nUdEc7Kx11I5uPC
lMxtoRRcFYh9GRu/mfNPBfzGLykhN4qYyAIHy6BUCOkKIDjJM1Oz8CmSiW7O2YYqqNWjw+/OnDLg
odXGo35AerofHuGu9L4pBQuS/O9GWA4cuhZ32+8bqwwBnluZGaPVbFfyvgU2tV0Kk2nHEl0VBYea
1G4ZslkZdtydQPx7YyWhASdKq4ULJLE6/NNG0HdOahEHVYikZrJh0oZlHIXyh5VlYGmKGsALRfsC
kDRcHCxUKOq6SDnV04XpgsMo8akGWcr0gCvDOk8v5zUGfrpBDMFcPXFcsx2+6xw25HoIAf5vLaMq
cM7pjYtH18YkTl+kFGHBMMd0hNhVjLj4vUY5hy8ZLS4WbLmdo2/6qItbtp9LgU1Nllrmwll1hpBR
VZIYxT3uDKfJWHuKgZmitfqM4OajxaDe1BJ37LkyvFjqh1oEGBPHewziMfw1kWOdQ4glJKaV5Ccn
nZSELqwtqMmDo8OZHdiTmcor2i2StjrUcYZah1UoEXXRkOiz/Aucb3UHHjAFR7Q5JdhbVrn4Vyox
/Tg6ORSjTw6wRaJj4uKc+El/XCWL+He2BkG3Si4MJF8aV7tySKHRAXvKS/3xtLz99Xm6y0vf6Nrk
jUImAL1nmEL+2Y1/trdSjkKge7rUIclP3soiJ7x7cHYLDZ6BjRkKLl9R7IIDbrRPZI6Nf7NXzHSp
Lu0CLnppKPPD7NaO8ieEGOZ63paNysc7UAylieYcVCJNqzKixtvBoYLeV0LyW4IKLrAXyTY5ImQL
BVkqtjVFBzEhVOpEgZHL93Zxmj8ozvpNINEn/Ku3PXK2vII7dgFb2IQ+hgxy0GHQsXDOOC6L4y1V
SwbOgDDnMGlPRPoO9Z60CgD6D+heLr+xDrB7+AtnDR8FShEJPIsyp9pWrlKulhyieWTYK7I18I/J
+R+C5rum7+lSy03Ac7WbZlscndJLQI5vto1wcKcDtjG2XBR81ObX07W9Zd2hU3pa2oBmC4Clq4Ra
gC8oJ94mL+GecjscArFulj+w8ZgPa4/QSClOAPJQhpoSq5qKEHbVUyTyA4T/bb0E5cIGVpCeiDj7
oDFj5dS1clXrR8YNcRhWA49kG5VbqlmndhF4aEHGOxnH73CfWmrkYwC8AgwW2JdzDIuYOjKkW6vI
S5HmfZfJq9osXgafClUUuf5Pl0uKbeCDC17anjLVvXgsWQq7b0hjwqQ3Rnn2TuTHwQZyUa7AmW6z
jMImcOh6Yl2w5Edy8dw81dkht2QDM+L3XQGQDvVVTg3hkggkmxvb0ReFsNAjqUJ8Mmm1Ss/53RNR
5fUbnYJGAQ6OEjDgbhZGPH6nnA8T3Xvt0Y2DLF3fJgVvgoOCbCkAxgVBNMz42yOzZH8AIyOCBmNb
0vtp3UDzDA1d/mtMsRoawDIC2I2z9ssR97xxUcJ5ccG6TNCDfjPFrJDSEoH5Sm0ynUgur8fBw534
tXjPYmDAUllzuX/xMBSK9AZKOu+9Svb7m9qB3q+T6EnTOVcLkGO+TbKnflmXORYnNs0UkAEi3L+M
0nhweNwlklw2wot7O55IXyTFtjEw7BNeXcOuu3lGDPGPg0rYppc9FiM1e3Bt8FMsX8+Pr6lWNGks
5UxgjXU3dlZYRqCMUZ7o6WJJRR7deMZ7IC4pRFvXEJEcuIu+MNKc+9wCI5I6IBegwmlOMJEWZ/VL
VQfHQD0x1sBkkQ8uRggS7OFfwm2wH1YWHnY/X1wrwfgLeKtDxM/NuqHTaJcAw9YKz6GB/iYnuQsp
VUCigepqXrgMW4XPP6W+lXyaKtRgOvPX3oTTuFGqlEixzM53WDxy4PB9sjTd0w8dBQIIPtOJZlGC
kZrIGDxqlVpvZw+LOQrqXsQVd//8mv+YZf3Xu6hcPi47OgelIPpeUh+KuqthApx3XyEdcXZWbmsB
uq/02+6GxifIMU5gmST5CZMkUF2YCZ0Wzl1U+K5JS9o3JHOI6YRvozsJVbgaR1ydChGD8clqnRZr
YfFUX7q7bU46rTUPZuxQPxkGEdHtxHBI8aOrO9bVk/X8GJ85mCwI3hGZUYZWv5LAlRvVUr9x9L8U
3gvIjvQBHThz6ejluX2N/NBVHOmdcNHxDNjxhIUy+j26ywL1SAqY6/DZGNJoXy/0fx7le5OneGNz
r4mKeLZUrqSadoHuzp4BB8NMCk1ZG9U5YqgTbJ0/tVa3cUWuPtIJhjfHUcOdXRPcuWjh32j1/E54
3KAbxJNMixbeq2dde7xQBgqJEAJYM65wWLTNinNYEJPrQmizyu0gjHjcxOaMNvxwFrCNjqb0U8Ap
G/oQ6Iw8q3XbhctzbJxGSk5R9t6jyWI5HuyJQLeDtMeopicwU4JPzMCdfKKI60MfIqUcgbwD2gya
ZzssOAqQBOsEUWnWzZjVgBZ6q5VG8/syl7JICgcf4Mw9h0VU2ohHD4Lj5BL/QBH1X+OWLaO+Bgnu
MzcqH0s6j4ttq5JNFyvlIviIK5haT6Rf4+dEGQ2PSy15gxUX5LdNdhnHcp4zgXAKMMrx5p0luPsB
AMBV2m1kFCLrxE+1GHUm2mTHcH3luP3wOfofaCsc4uzfUw59zUO45pXUwAjibQ9zYBBBZhr68/29
CHXlNHfKqJf+W9AFzsM4OlbtNqrKPz6qn+4yNjV32rzoROFJ+4YU9FhgFIrMec0j7oE2wDfSNMJ6
VuH2dOxHxzCeeAthwhxM0q1Si6qplyURQ9S3hQg6Zt5T6+DJhhB6ipa6HfRYzr+3Ry0SEc4yMMLq
WhrYnrobYmrgYYiYXv39iZiNhGS6Kesq33JwvcrSQ9GKKWdt5xVDAhBvpfyrAS5fsEedNT9kSzOF
c54H0Nz+IEGHbP9B1lT+4j8xEc+lyCw0tGQGzXyp9FlwfaDBaPciRy6iwWnv0yGQySMcwPeHsmQ+
4CiqZtciIlSiiYpea6wf/oJZKzWvzKfDKfDvpSTQDYoEQOciqGSGz3NAka2sN1MuZE9BQzxvDNoN
EPyBtBiCWytlMSu8iLm+ONbghf9JENhwmZSpSgTsa8QrjGL7GCL+x/D/EDqnTfZUL7AXSEmz1mf0
PL2exkgBMbzFiX+9HzNNFDEIUIG0U77n21kuTAc5oTPNTQq8kWUtL/wQ6JDDZWBlWqOFXJJvxGt9
mDFMgzzK47O+wG71hHWfq1Q1f9MHQTdTgKAMWr1aEt2pn3enKxRmZT9Nn5zTH31vJi/bgEWlQiiF
fKNp5gSyTI40Ul1TTp9kleGXuD0clLLOjVuu4SbFx2lbOfQCQa/58kFfkrEkzEKCtOKHmvNAwyYJ
s/dbtarrz2AlMS1OKTQQljsICKEJsXzjNE/eDZ1mUPKr4Dfr+L849pX5l3KvDi2ncIg3Qk4KbSe1
Y5Geqej3puaVgvfoScFZZ6C2MWgBfQs5QoNpoNq0CdgogycDZof9aJqq0UEcF6FApMQwQ62p3eGp
WooiIfDoExg+fC6mzCNPPivLGADX/xeCeo8MrbC9IjRpgYiisHAAg+HrHQvqkg1pNzeY6Ao/O2xK
LUvcRCqXNUqfjUQ40GAkEK78Q3AqFB2jkxHRxuYgFDYeW7cdlhL3yWeEgX71Y0Ilyuzp6I/6fShl
yLe3eJf7NfotGmUlu/udQbjPNfayYJp1asejrPiJttBN+65lE+DVJ0a9qgPXUKl8h4G4rfq2La+d
zi9gjxLB4GKl+WpfUBD7PctIwTeeugox8BhCuYjGl4tZeXaIsk8zEw5Zm9N4Wo5PKM62GRCTTMQa
h6Qt6nbBawydRXid0yZKwBM7WG4mNpSILMtSyDj/zwKP2uRzfI58baz1In8S3s9VuZQNW9pwnbQw
XDYW0MADcr3lFYid/j0TJ1MQvSiuoNckCtBTNRyQVrnmX5PTLpcXJQAoubWiuTTfWiCXnPmum8z4
1Xg71Tt3Fbjaa3f22XCgGNcrycTyaOzEFu20WbDVYEZ1RV3ludTD8One4p5uLI7AS0iMnrQFkDPb
fhnHdA3NsYZq4sRKHIYjrcN8E6ZUPlnjYqqyV7viaiOr76U1tbaH3nvRYkT5dX24R3gJMtMbpaGB
WB5hdMw9KQ5xORmaUYxIThaBuBasRyw10OHM6vIeB6DkNnBM5/pb8Z3s5GYnycpl2KUfXSy/SLz8
cRHwslTVDCQbpmTFKpES49zTnKxAZxA4H02saGKDG7L+6DDdbpDSpSMZwQ9RTQTDD8Uhgg3QOEhb
TjCgdUPqNbU6veH/eFPuFNhZzQ7N55sGrNr+w8AbL1w9FbtEfbZX3cHJAzA/xEEbL+QxR3/4BLQX
DlA9CWfl9770CSP5Z4qVcJe6++X0Sjy6nzNrUGAoAGC7fViUjD4Ze7z5LGD8aSZedBHZzTZFTuM/
yeZINJv7V/pCGrULaDsQ3btE4+D2KGd2V8wwVV91xUt5lbiZW7dse1gV1hx4C+mu5/Qo1Pyc+buj
RWyUol8ALVJfn2Xn/AvLr2h5WSnqckAfMAn4OAjAMtnGui57E/azo/ezxuvLNHjvoPG9g6b9SUmC
/VL+Wwl9HBH4eiUR2msonB2w4PSqByPvDdkgKB8fBWj6ldgjfGNgpVBT0qUw+vXFs/KjowY+TwWH
87ku4eKLbe4sFdidIRTuaABxMA6MqZu6pKsHJy3us5arTRj/xq/dzRDgssANpptN7JSMstwvTsb9
nwsceE+yHa1fwWncZyDjrLIEFNGYcZb2IuYfZpZcgO+50kTy/r26US5w7E3kgSsPlwo44qz76TqZ
Mgu0YCicQWXGrLSH9exkX/AHYmvhyYoPgDpkGmCQCJEQX1+Dk23NOr7CqGFJiO4OqLJzCnMds3mO
U90mPJqYXlcsjyIJjGNx1ifKXqq2elL9q4KPoeFgUE63f0psQiaU6SNbwREkDeudSj58yP6StscH
fD2K55hrqoD9NiliZtPkJeAvMV2vZKHCJlQnERSwafAj2iGRZcL3l1M3Y47ftbRuR99+vNneW+U1
z3CcXKF5ahSBuBiMIjx7X9qHiipQu5OnEo4OKhN/7Jisk6EBLiGzhuGJssQlSZgHJmxZWW5k5dfE
yRxr1zPqlPx0dfDh06Vbc/MFA29DKff2zHxNeCBV3L22/+bT4Q4bvxaSkpLhEDrzjtoYeTbJb5KE
aRNzqfL/pkPMhTv8tUfXzV8SumW3XOmyaJoF2dv7nwLOPgqKHE1PaDkjhS7BQzg486X8k0+FPpju
W+NfS1O45QSXnTTl1xMRBbv6Bv7R27U42TLl3LNjchrZfqgtspWpTC3mVsrohIjRfGCt8mjRz5+q
5kgDkZOnwXAaUZoI1qWwXl6p6sQYHZpqgd7WnVPlgBegdLJg96WjeHZ9G///Epa2s5ZbSt44vevZ
BJbsWcDmFe8hE+Vfvjr+YZvYAkZNmcSubtKE47MwS0jGENH7uqtLXTktkn+aYTawowGeq71X468U
EG7+GXTA139qsKKyJpcEY/Ms6RVjOF4AWR4336VZ/a7L8myYVq1sEdAuNcFv1e8Sqp9PCduLY+J3
Q5GxnnECr7hOkYr0Ao3Er284vu7lko1TW0UANQ8YlKQdrAqtv76VrpmIPuauvsjbBv5rQU6ZHlLw
D6zfDDTSKtFDy6gMQfSlzAmShUCqO4p+B5utz4FPtE51QN1SfLxcB4a7Rq/oY6i42hZpczUgrDzB
3uYRvyo3wowJlwIs+np98gKY0YWC9TYWc/RJwHC1EcJziM/JK6luIDLw8qRc96q6iw7LH8lXiwgm
3riYB4k3f1LZGD43KOyuZOyNmNJt0E9yVvmFY+VjlgY8kK2da5XutfUs5G/6bb8tShcyvcsR9HLD
wyogwW7Meg6oFH6+Jf+k4YcJyO91PnyCwJPF59REI3ur3agRmma9TJqpWLz85KQS/ICk+SDPlAyU
6wAGtDOWwHRTMySPJu5vfjqBHOo3GKFZx2MqZZ4f/9GSxoK0bNey2ydtiMQrvWUtDPrnPp5WVWcl
3PWb8fKkAH2xAtakzfzxPL6Pc8w5W9ksOtldzhcoDDyeuzoSIqrVKOXuWZw6Ot1YafhzoERdMzZ+
WprsUAKaJhH7nAbudyqT4QurNkQg+V5PRa5eilTAhfin278l7/cmTcOG6W0rUz89XULuuSX5DsOt
LKOTr/wwdCvjtQUpLqhqZhDHTqbLptT8srehx49H9zYj1A1htq2apA2PY4WO0gN6rVpM+M+Yt9O4
9z+U3QPIem6R/GxMn+8eBLKQdM6FSIpfVb6Zq+P2kWKqccR6ZsFZY51vo6B6CtfgewKCVxfaHVYv
cQqFW5AtpY92O6VpN23PIUqPeN+cuZAuFD5MlnrqUE8otLiX31ywAvdV2VaqdWcAtrAW8CmKO/BR
TeRzP75igJfa7QUm5CId12K7dZ7LqH7wv2DHi4NNrVPzWY0dVfQlRE6dGrRPkYS365MggB7RUi/O
mUysrnxk1mcJOtIiI5Wfd+XLkwb/2vhb93cRy/VNzpU98lFr4iZKZ9MrFH37r4VDwL6y0YutSDgZ
Cl2A8oUB5rIOo8yYR6GH+Onf4qhcR/QyllDz1h+TRyGXy+ne9LplROhBEYjXgaGatDcUeTmK/ShC
3+mMnLd/hQBYPZWuEyTxKDrzEMSBXeebVjCZK00eYZwk1odbKNiB+78ur/0L9QyTT+zGXCknWyIN
C9jMDWjhaSTl19drGJddJYFhE9ZPrVGXvo6pbNL93FXzwgHRGOXu7zaQl8CDVSarElucLS9Jt7n+
61cjkkGsrVgygomIIKDSZ4tangy9FfVw/3vzDraCpWOgBd0cGhAWLp+M3YzsMdcxDu8E7bOj1qj1
LpY6RbQ9FeSXj9NOW6VkHGmBDMx8xOum0KqSP9WvIi1G9+X0mtZbKwGyu7pPyeBuo06tizS+ZSFU
jazm+i8GFgxIx2lDZtQBcm1zdvLzRxTsiEXJrbXH1YOPTVOZjQX5CGI9wdv+BEVT9EdM/7lklyoI
CxjX7g5a62wnDPt7ZhwjTkXVpd0OtvY4Zm9aY+igVYS/I64+eCa8GPpk1DG27SPDrqS0KUKwKAqO
214zUi/AFhrtIEQljmwuqvIJlaW/RxlJUN3fdjta65RqLBK8vE7G5M5IriP0HUWhzMpo7H9eOJ9F
xT8kcFnVDdIdUMDifsWh6r/cENP/DjZUbxtZBdDSWZaNLHEU+cZTs5ezPfvnkTaPUSAIC0N2f7SS
6Yw1kXewKvqUfNsoVZjiXy1ke+EIsNYDezkZQLZM85Xh1q7jErzG63UeBYN29icgiHr1XR6BcCFI
IqEszhn6j9g+DAlXvgjhGnonG21J10npVuEWK+bgc0xYNJ/BULQ3C90EFQYoldZUqFHerakT0au3
qALndo3Kr2tO/N4O+Cv6mXdfIX3Bqk8gUzybbtizs2HbxpIpzh4ASkwVroGcGQbJCvfRP7qLVluG
gKRHiH5nscysKGZ4hWb6W7XfqqwkydyTwZn/Fu8pSK6peCekPEr1mof1EPfCe85y7+sWOpOrdJpw
kdPsidg7usCR1cJai35jnpB/4Ng+BVjGWEpI7GcU1zNgrM7zYT741HkIcOxT7a2pi8qSqdJFfI/7
ICnm6AwRI7rgcqr24Us4FjbHTQvVhR7DDKe6jy38+lKHUKcyuhqEMQvI7Fzq1+x3Kv0gkXgg8mQR
vJoWR1jzH6kuPj5qS6qI1+9T0qab6d7PhQUQgAcflGXeFemH+G5Os41Bepjeg3bGdCO2n5XzTmzB
ArUay7nbaPAln19KsGcQCGWcbkl4HNAKVQofKWwa5NpPXVwjojOkdhF49HeyQxzS8Lv1DyMD+rBo
1xfpea504K4Jqei1/A5VoKqfIuTsLA3pti+AIrB70tOuMSZmrMVGPVCucDH/O7kVAUGSnls5ongb
FSpfehoS1jGGXLttpp8TmTC2juQcwW0Sw+7+3hVBXII3/LJMk7uXODnxz0C/qYzElWmmYkFPi1fh
HxD5oEngjWq9Dwf52GlMfRuGjfpBTWayEEJJzCI+f9K7/8N5aR9HDLgqqL7UQBIFMpw8jYRf1Ez/
pH9fxc1f6ElNHaLlX3cg6ma4+ai5//UXrjWHMKIGpEkfctbj3tq+UZjelSl/GENzWJysB6D2elGA
RB111dXrRU4GwsVj31ErLgqQA5PPYO+c/U8B2Ou3re6+ZgBhDQ/jCyYWMgU317tXCRYoB+GzVpab
RPBJWm4LpS0fASV//5e00c2mT6MbMbkr/N7n5rEixrA70YGYikgFSFFChHBbCfVrqvUkvx5K3aE/
zRwhjQjG94QsNgeosXlTPyqn+mWAfo/sTRm61Jd8eVkd9+1vKX4TjPRqsAw3g8eqC/lmq3KAcwXW
+JKRWM9SXoQyZhJTDCM6oLocj6Khvbw2+4tVCybG7mltskwhCvVGyRrRpXNFkI1uEsK9gwSkIanv
FeQHCX5B2u5lhZxS7gQp4XdJtV80T0TqBrIg+64+/+osWxWMadLPwj4zIkhcPKdxlLsDU0bjqvFm
M3TcDXN0k9mEPhdFbD8I5gSZSOGQrgjjPFVGTA1E1aq9KRcapwU0ZROFp3dQ3kOQ6qi9t1IF9NiE
2O5Z3a+ILYkykoiKMW8g+5HDS318CF1r+qxRSOioWhQ4YNpMeWEXZG8mNNJLFlHLwnDbr7NSwck/
KnTNwctvlVmVUsNRjQNtotEEtVvViMqETHq4/jiMJmrYL0qX6nEFx9HxOtp/15fmxPiNrw6vuJWR
qU0lWMPypgYLq4AacMyuWNXESggiwG88ntgGMN+WOiiqGiYfhgD0Fh1h2ns0D8lSK/pFs0Xs9Zaa
qMxNRD0hQx1zrB7icT5ip/MK0HRa2bpzQx9sY3I1CMBcz1RGpzC1b0sIwtoKq0zUBnVXr/vzxJKz
sAUUUl4Gz6ru2Lgb8LBHYQQ1lhSNhrCOSoyG5jAJbEeD4ZoUfDzAZbfoVqHZufbxMGCkbhlKs6WA
NlZ4FFsdEnKcPlOBiVfn5I9M6lzpbbDGTFcdDdB/cOHMSTd40dcmqCf6t4tSg/WkwRWmteKBJ5qy
HZr0/43dXms1bKTl5lUpK2wfsVqclWf8fgx5Va/c/MtAYE6Bq36WE/z66KnnlKjLQIKiTfsKHOJ9
o7KZN5VN9VA9puNtS9cwydu+XjHnbcmOPt9hMyqqQ4KoA4+r+bXDXzWofMsGyzLal+nNe4OkwRKP
G7h3McLYInfHu1EZJVr8aCef7QGQWbbO7o3MKqMq04zu5fNyGbORa7e8cNWWDFbev1v21eTpH4I7
avws6wf19JNxXAdMD/PEdBf4SrxCJ95gl5twLmXSLKd27+ndWbrjyJcd3CrTguYeu1CSAyuqCXzS
JLcF2C5yL0YpboG/lDsMKtQIPsozFQWnAiz3a81JCWm1kX09XTSegr68ua+xEQcinapZOTaQfqNI
0nWVl40OI2+sf/0U0ULTBL2TProT5cZjD2C/AyE8ZP3wHobZ8YR9N0MCkHz1zW8h0eE7VNq+1tCd
1GuJj8/EfS8LlK8Gndmoom2vJgUS4G+O0wthJVaX3mnT8P6bIj7HFDhxnww50wGC+zd1plvkIywo
2xEi3yc8wGhedPSOprBLKLMWoJP+qL2bZR4KBJczaTyMBLOrbg4Nq4Cz/mKMHS8EPbxyxO8zARc7
kVYuGfPiBr57LIO0ShLdt0mXpU5cptBNg946VuTofG/+ddO6UBUeaoGWwTRG4f7zeQxu7nibazxz
GWNgNfKPVcONppUuhHzs2FOlRjFExto19Eo8PvDwiS7CHApUBIJaZn6Fbqc4eQKyNER0CPeMpXh8
aa1UGMcwjZjwpekbB8hj0dWQiIvpL0ctSWbtdEqAHEANF0f9IY3s1oeZnlw6gYbqv9G2DDLuJRh/
YHY/cMQ605XcbhFeCuFJgFZhND54ADq+RKuz/xZ/AeHVCG5LB3pyJhLHL8yBOyRCz7xH8+uD/0W9
Lx4YotOdx7jb16ao/xoF9bxUIye5RyueSdEGdG/bCjMUshILfznqjfhox2Dh0jnRV4hqu2r9n4er
21QP82z7h+pVBwBYj5DSExdRXrGHf/4i3WVNpseDRcYNmJcEuvypiN8EH/+d1Nc37dysXj+nXgQh
Gdq02+5vjShZFt/Fl6zYNyTFmgF7z/6jiJJSLrxA912iYkfVyyisIWs2o8WPhE2VwxhXchksBnk8
0+0sdcEnnS/h8ZePfvVpJ8fPRn1mgfqiQGE5pFgqedoWiluN9hMIPm1piunSoZexJ2oEQd6HdQwx
O1w8RUtIBgKLHFrbpYU3Q19jgyqHZNH4L3pznoUMXsp8NpFI0y+xPn5l+JAL4l99dlmbAIQrRp3R
FjlRk5qDbuBIu27wOJydzClJ60fkZywtjmhFfijELNEaT+E9dyaU2i+sZzr1VTJP3v2lfnY/a6bS
mYSFLDUx0QxkwnrBN0wGJ6ROwM0B/OdBIX6RhHxU4x0YgQLJCUdQ/UW0XfsUPMxmRVKo5NzOTFSe
IkJ+dg4XpLuthk3Ghi219ftJBFXeaeD7akjGqLE7rt/rpn9NJc3WiV/9ruO6hGTd6ktqx3ee95K8
9OScjlw+gMHzSYWpo0JhBBvOhC6itaUYKD1v1Dk9cTP4IdX14BZM9yiM/SkxFAiZeaibq9Jg64SP
5eRJghjPsSN9Ndo0+1iWR5oimo8XAMidedxZ36kInT6BeglbG1eJ8o5NI34W8IBmxKxH8DNLMNif
cubjguiE8E5aGoaHRvcdRb/WXX1H3EXHUGaAkwM/vHCTYiol8F100GX+cIJqzQalhecwMg/4l3qC
E7ip2pQQo2dN3IgkJYDJlop0xPE1XqHqvrkNlHyyf+Q9fF+b6zGxGqn9vfE8m1iLPQJMoaHaOsri
Gg2NAbTM5viDyRcV1Aj0pY7YU3CuZDOsqk4cNUpO4xMqqm1BnCgafKhKRyLwGgZsmcdZ9m9rh31g
c2Uj7NhdslKEbaSfiQ6mwe+LkW2J8CY8Q6juATPJrY0KoV1+xyP8HANFIRR9VL1JWYALPRyz5Qpu
jpnUHmXDKvwRf6pnGhxSnifZXYak23t5YXZRwkQtBd9MD0aP7/0f1H9yZxF4wOLG9Cxawa0Fpql5
bu+Zuiy2oi+wPDCSaWLh7VnvEmAujPndW1pHmzfHWdUUpnAv83O/eWRy4hl+SECA+u8jbzT7vA0p
kJb6LXZPw6Qx8cVVyT/Kjl0gbifMaqCktncNctGDXwTpM7pAZ4+22ZY+q0xSTNHS3Im8zmgvgRcV
yNIg7DiJRGVwENyM77au+YYoSJTB4lpt1urwGtWOXaG7wRTaPZQvaV5HVFa9oH0KvNjojcazVRy5
fzPs/XC8eoXDkcQYGewH/vdVsSaoykGuDc1sjdcwFRr07JNHyalZltUxWPTc4mUSeqXdm4CiV/1W
RL5VP2hSC0OOPDRd3zsS7RssjiR0yagBFUiNoOttjqezoTqFQXSPUsNAls0Uqmr3NzLPFh1sJxro
bxNH/BAJC1Hz1csC5w7PgFTMRRGkMHPA8CsyTWzLaloMBr+tS9fqBZZK1o2xGbjZOtnwZfolgruF
mxCD1vgoUslmnBJfogu+/9C2rMKqxz0KaLA8flbIwA3FhhS+G50lNwcrl/U7BKNU+9m/8HL8Nl8+
7NmeZ0iGNJAphOCUwBBiu4LJLf8MRqpN44IevJ4Lz+jNm4dcLMT3KZaoaLASKSK8ZA15z2coDUu/
JZI6wYUeZfM2o+UR90n8+xH1qe9FLe+r8UcDB/YUTzgfgsQcALZ83UFhoJ9p4RHf8+C1+tL4doEx
vwCK85fXdlgLRiMvYKTzto8njMs86ZhDErsewwiTdB2JsBCRq4hIF+ubVi9YyLwqYiEwXnQjiv06
GGFAKIW6SW/knDpPd7PDp72DvPmQjVNcBl13vGBF3YrtZTLjJvkatEs6u2VyWSN5xU4kAmvtYcvz
zSkn9I1O+b0nUAPvkpTppg5X1G+fyDbBy/THETUpQQQAuOgeYc8XEe60qaismkTVwZReR9r26KOg
TsV5ypLznZHrp5qVM3tvDvugBMwtmVnMmniwyJeX2Gi0+YRVurVifWD2l4NU/603mDjUVDIb+5sC
OCwIhHAfijhktbr5qi1Sst7Mv7aXVUlynFN1q7AIjE3TpjhpowXz/e+PmEXsyVQEKw/Zp5T7FNly
iYXSpaU6QBurDL4+GEIPwkxOkd4v8iQ0pBkljM19uqbhc9+Da7LKSKvCiAel+t7nVckhERmojewZ
RUqBZJE3N8r7/XN10Ws62TURtiEwG9qpYEx7i48AVrKiLLGYcZsQDYKta3+yPYdKx1L5EQc86JyI
kQPnimh7f4BP5oxAB4QqDbi7CNRLJmiRPHmDPgagSwYY/6LFJ35RA9E7R6+VwbUHLc8LQqQsGZnu
c5oJcwPY1V3fF28RD8yr2ZCgkZkOyeT/lJljvjxayExhLPkLOM1F2UH6q7aT6Y1YkIU8fAlkwBfV
cOMtqwFno+kPJs3nt9TI0ix7lrrRkaw16z+XiXSCAtpgBEHugjLpyQ+hwM913IG/VGlj7LE1OG9d
p5BDDXn2w498ZSWJqeWgojfb+SyAnCgON9x4nLni1eIEvhmURWD6RpNsROm+Xq4ylB+r4YA72NrU
0Lit8Y9wJgO7JjNA1FpBh+ZsYruqjRxogX7elGiF4HLl4iBNVGHU0w9UC9cBkS73p1kmX4Wk7Cka
BsgeiWh7KPO2vAPlM9sCzC4d59uFgtOKlkXKRrRQHtDg8G2djeNu1wF3Syubynr4Uxtkl/kKqOuv
p3156SXQC3O5DnldUN8EhUQKTCwGXJwTQIKPVw91/rb0ckFtcPVd+UtZ1e56SfThOuxPInVmWR0I
dFIqlVeMee9VksGkPhIksu2ofarvmzZSHROfETfPFokm6hSwW1tXUJmc/WmE+8FuqaeIcGXBlbFX
85GrSQ4lCVe/uvORPG9KRvA/qwSzUKjcRVJdqIITThnuH+XvEBeONXW4C36dhBFukMwXAEjTTbPe
fh2OFo/KWEoOJ2G08vNqITQOfMcvn3Dwg98imKffDRZBu+B5bIpn760LtvRlBb15xn92UhJy8+3y
4QRNx0d4UozyxEd9Pjr+1Vk/xCd9sncTIxX4u8/9EHsXk2QiLacSYOCr7I5HqIVdNi62nss9xJzZ
j6E0pgkC7D2PFPM7wG0V0hZZFrX/d5X9Ah/XWQGePIGFM+44jMV3S+qXhwcGskN8cRKIY2R34rKz
I0C3SrRJK1O9xHTacAKWDthdau7wAYBZsTSxRyfa1Ml/ZX0NCgg9FsxoFLQiXesh5Awt+Fj6P+Xe
Z2ELlObVVhbZS/83s4gRuA744e6P4Uvy/GeTdZt7ZdUp2hpy5B4HZzyatTZmnfQ62r/3+gwPdbuw
ZYv9XHhD30cDnPl2xmP0O/J2FDbkFV7TowJbx0ZTEhmIdhzVAHfZP++Ab9yVyzJn5XYnz+kbVptQ
Vkh9zz8DCSlOAJwREVsZoVplHAW6SFq7t5RQ8zE6YJKpdAqTUIFqM1odV2HNbm0qjZ6HPV/MfRFz
us/wA1fyPwDBPKqUCC3au2dl9Pr254fr1hFrnZ3tKEGis+mrNIne4WW9LXht9R2wseke7+Ad+F+v
loKyQGGcxFElztVEAgK560U9aLS0/ckjcOeggUUywBtjfyqaS9cl5xbB+g4L8HOZwsCH3gbvmXF+
3QaP09CWcWfz3tev/IdVdWRZ+w+ruE8uPrgVoH1uT82RxV/MBDGdmgxWk3fl0MudJCSMJuNNkAp/
0tT0ryMA9VMCpk9D3xNp0Xn4+SweE1+ZgzTZTGIvg2bdhUbrX3lBplFVUG+s0X88IH9upC8DsE7L
nJ92TsIuMySG6C1P9pldYWXZxJt27iy1Dv8PkeGPTJZaau6Vm5GXRqGyzpHUcIhRe8RQWRiKfBcE
GVvrMWPyalQDwyXILhzLMCAxcL3OYynebE1YiKedhjbtRpwDloyXzS+CSVVqcjphkIkRU35tPTC8
F7nOZaq1R1+a8o+MRvyzg9odDCKYyeLpNI0CtQSRoenuaSeYcqDE8wr/TSbyjOTo9a5tKqkx+dmh
KTpjfl4imRElb15rW63stNFc6DleUSqTJ+XlJw7GkkJYoLhWnKUzEJ/tZmqZTCU0qjo7fn7Jnwcq
HAyv4H8I63BxDpwi075BADuqtXvw5MCyaA9exv5J5S+GQqVvWRg0O6gCn+JWLf94P0hRYoalcP0d
CTj79mXyWhU0XAnzyNvwtiUpgwnFf/ko7i9ubNPqQK2mcjVhMgl8cgEJKH5cRffR0TW4IIX8hWrA
g+a5dclz/CaoE77USSI/72zdE5P0/l12kMIGYVtMaZy34Isdwmg7GatWUw+FniKRwv/D1IY99o2o
PjIwBmlbAjhLCBPF5ydBWisuVFHh3ktCPeWlbBkGtya9V7mTkoUTkjeHAKXW/1So9h9JJ5oxeImw
y/aw6TMSLm22OGxpEjYTJwXIcMtk/GclUV9FN9318zJfeeqpAxV/Lk1awT8rshfZ7ubw1/CCewEf
XJOrO08HhVgC2XYrS1B8OO3sQu5UK9Hyive7gVwgbGNEyZC/pPCkF5xhrDqRdsuCLtRpFh+X5pZW
0vJ1kdxToV8ugZ9Xc9rKikNUES9Nt12Q5Xo0GXkLxjjI8zhb/uLAQxMjVf3T4GMKW60ccisLTKNN
qjnf6TCMU7bF0ELz1N2kceN3/W9wqMhy1fprXsE/vyTK93kRK3HSVg08LmuVw1tQhO2YjIj+3vaL
7n5qQT70bshHLr55Q5ax9VYp193zFihu+nXfnaIwH6TyJskWIlWRnhZ0eHg1hx2QGsGXdHuhRGJe
Qt+C4zCrISbaRiUl5nlfAt2UgsVnZvukfz2IVE4ISEcjFqGRCaGw/MNWaHm65tRE2EElAdD+bsbP
1dES93o5yLErnILNgeyAji9Vu/jI6Lq5cK8cGPeiAWi/UJA8aXm5CWkSuiZ1BbfZ+0UsNJDOqF3l
Rn36oxDVRGkFthr6nvnDfVFCi4OxoIVXY/2QnhNQFIF+T+bOpiH/+5VIW9wSiT0ukMs7YkvtU/AQ
txh5lTfUhGpZOreYxY2AwAEXMchENTPyiZQsjX04RoOgvlfjsZW7vkdZo/wl4QazxDF2f/qY9nr1
9Srw9yMxvdIuGv+MS25QfVb3y3LC3Ha07Qiqk7iDPv6eB5h7zlTPZ4h7au/57PqdpTtoqeZkIE2d
cb1KATFndFWOUGwFY7b5zbsA8rwA6ICkeJZYV1+AUU93aigXL+/7I4VD66z/2Abx89XZOnAzX3SD
usOsr6Az98gK3ciS2VF9I0lcGFT95BHVzry8lQ1M9gmaNnSml2ohwlgkbhMryH9XtGhyu6NXKvRE
ZwE4d/mWkGkp9uc/GJsdqws2qPnMSzi/+k65THnFIY9xUyxoQRcc1ZqVC/nhtPP83ijH3vmpMIq0
aBua2or88T+dybSVRiNOwsNKodIotteWNAaLmdoDVbHO8Q3unZ8lUAMdpf1Pz5VgtxzD4z6IeqV0
OvDmdmhgJMjxftJsiYGNML6CShkNYueLFs3rXKl3VlFfD5fi68afTIgfB+9s8Tbxix0jx3zE81Is
Ad++lEpTdc6vzYeISODXSqVSduhvIM6MbJuUqhe3c8o+DzzIaJG3gHnJUqHWiEb/fjmQQzlBaDmV
35kV2XkSGd/zm+DPZDu4ucZSsqUQWemD5Ib9vpe0QXVy8QMT2dwVezpyzAAxmLbHDEMjLnwYGfWQ
/1S17qB87cLR7C4wNmPuPpQEzBD5SBnn8Q13VWCpYlFJSc1XEzDICVtBa4FqOnA20j1sD6dyLJBE
gw4YSPATbicVFHkNRjDXiTtJm3Ncq+5abaLU0c6bjW3ORgN8AeC4CFRLDOHxe9AucA0hnH/9mW5X
ojZU0bd9TYNQnYuymGWlsY0bhjjH6AcOZQQtdSlhCOZ1kDCqZKqtsBOKm0eoCJPoPZEibBUsjoge
bV0uVuPkGiFwVUu9X2FOwlnT1xBQaaMVJdwnFfrC9goKIM94a4SvYFqB+Z/7ODlNUHKGVimVLJbh
+JIHbXjkXv/NHXr4xYLIx5eMAd+plaBQ+rZgUw7kLoO2kRKWBj/G/CseOJ8ZT/w6CUCcXhVzQySx
VNu0+JD9GVKelNpqpGeKZ2v6ahZq5MSqXy7JZnnXiPHrvzsrVdgeXerEt5ppdLcGDN6EN2fJdwon
l2ZvJLsF895J/eZjpPqRbs8ohi8I9NG1eon41ykfwcUptdliU9MJ/hYS/ESl5Mut5265OJYDjngd
bTDWhHIYsBRkhuGzKA9V0IDpcTve+Oh2Anszf2nH0KWHY3+oLVpNu+c9Ihza3NU64TtpSJ8MAbxa
GtNLfAv3BZ5jEQp/qFi//QaIvBqjoRPH3Pg2EeGmuFA6EUrUJx6DaB04tp8hFsL2mTPTJ9kfz58A
2Jkt4hjNdoLgqU1e6Xc8hOOxK/OZ6KA9Hop7RY1XE7z9G3LLID3m6pf+DNqeN1UuV8bIBCteLYLY
FXziYzwgq7Ymb23tOX+axVUvC/15brPexn6hnPXza9NaQUY3KqvXlI4l8yZwmR0LYBAmkb3WGNIz
tghR74yXaApHGllKnNqGFTM0yT/1PKjDG9MEH17lFngge6Wo0xahlo+1X4a953fbjrWnwc7wSsnY
RLBzF9HytLKba9y9iAti5gu+lAmj8arK+RQFM32tf9yVe3ucllxQ/Zmc5Es8TSWLMBlFV6//pFGt
YVpeclwIGP0FowQNfMM4BJBhWuo1RhP7fY2uR9QN6SU8LnbPtGGTztXMDtMUFXTy20Q+Lp1Q0LIp
GqzP+c++oHiaxG87mGgrxRWzAt8yXzE9FTgV8SY6hp/s9OPIoW1LhLT5yBiMZxR+I3gFG6dmvUGZ
BBlTTwTpjG7SRWCzI17CpEuH94gPpHhyTVdo4jHjifUbKGJIFw9UOceQ4bSg5KBqZZtzbueHLGTM
eUQK+5QFRgI9LL/JXkMA75If+K2gJm1kFRvIELmcYDTvxHDP8yu+93FikS7sMD8D/U3JNpOFYnpN
9Sk/972veb4v7QzoWOR27ePCGJBvg7korZn45zGmiAYLVVhZyS1/DA/NiMRvqS3wXyfIt/N7+pjk
p5Jxh7wQj2NPyq+7fiMFojzjBlZAT1waYbQpknKWfxdZDHbqahjUEKabkZl7uzBw0OcdoWW4U/Jt
u2ju+QYRs4M80p+JzHnB+q/4HzPSt823RM8h6g8W2nZ0CHkNE8+h2Am2/4y2xna8tjDVHlnNXgYs
o2PKfnSIKQ9/Ko8/aGOOvT5mB7ktIZnq4d/B5fglqxYLPjilZP9tRJRz2rg+5Je/tR5cQQhOHRkw
/V1cFt2dxJUmTZyHBCULM5BDiZkbfJJTXZPWbEUPCb8DC+ok61sszBENfkHulYrM5HDCWLPa73Xf
eQpdvURgIODjD9ShY7Oa3fxZzCXCijzJ5/pJZ0KYnN5YLICybXZlOuLOWpWsG8sH6A/yZlrKxsPF
q5HlVPZCT/5w/fvusaxuN6kI9iZr04H1w0Ovf+UQZb8l06hCFBO2fqEnw6XUvzsBhTEnMNkZcOwS
QyDgCS/ymhvV2DOWqJbj2nbSoxwbmShgi3N7J9Hn0uQF6wA5Jentb64UbV/6QmxdkvoN59TCYrTA
rziShlFw6tG24FevlZ82W2RMJe2GnJuAtvEo/AKIWt7zv5XTHfyIloCKYmPivNAG7XEN5ffu/bG+
2Onfu7uXQpAf4CsZKf3DGoWB4DFORQW0tBbw6S2UoG6AoTUCWACAx4gVOwQssv8mYii5usIvsnJO
yFOMkCFv0oHNVlOBI5MMIBLiwEbAMKFMcCLB2YSoEpVK84pZfEyYi7MZk4iOEXTKBN2LJCfQHBm8
pD7cmSZw5wUL8hz6EAuztHq7USsHT2jWp1BNNdw7gfCu9NEXswQuuad/1pJKWJeplAEixi/uXm4w
PwqRWpxeW+qjjrtL3DtaMMvEw+J5owsqwYSYdKe8u1k6eUHU1KxTjuDZlgfR6uVU7tAL/CHZKc/1
pN1QsNSRZJtk9d7L25SbqrBquA9Yj8RpoJATKOI6BFCiDWHGoQ6PrnOYi7tZGpeKJ6jg1I0sHYze
8vx03pl4PLT8cVNpU894fp+GfAzQCxr+pORi5VoMfJ2zMqby3uwj1DrZNnYnpaZBapz7i4oONHzI
kkKiemsFhP9yggxRjT33VhwM2QYmOuHvbJMdKGqoHtC9NGf8MHHGLU1o50VImRjwPFIARcpYPGZ2
SZgt9ZM+ETkNI3szq867Vd5tVIHunLXGX5x7l3FWnntZT4Tvjb4E3JaSxowaiYtolDaf4n4yzr/2
cdbf+wNUNRFUmqkytipjY/ZuyuwGWkt5lXtY+dlt1VNkFEcfWt0wvdMq13rL5lnggwL9r8hXKswZ
VkihBvD6eHcqP3BtnAqQ+PPmRG6RBDFpolP0D42te8Ij+sqfYrBVISafZVOv9sGTeKs2tF5SNs6v
k1sU+b0lzkEKb6QFPKVtf3mVwbXET6sg+bGhkpTMYVbf971XSkCVBuJJZ+bzFWaUX2ev6VVvh2tB
BtyUK+yPniRAVqkYzZYVkAp3DCEv4YH2e5SCRFak6b00NrvgOWQr3RAF+bgTgwvZZuktm/yIHeyI
3BQWVTt7pKyIUnNVAXYX6jv8BlLDprZlbakaZCYS2At5ryEdKc/34nt14tuNuNEttvmwIZfL0pzd
SmQCH5tSqrDWs3KAor7RFmAFQ5pcZCyJsnNC85bvrGg/SRqlB5+z8sypon1XCNkYY1jJOamvwxqZ
264/jcnStbXUFt+9Kzf22LvCa8sFph3OoPL63GJFtfmHac/NqAnsyl3rmObFbeUaGaUu5sn3Gu+g
5wjdPEZZOb2227t+rXNPIEU4AIztMTo9JGA+fsgIrY7oFpbIjC6ueQ+Q6kdobXCDJK2Rh5tWIGZd
VTFiFyRd+7GdLix05Wtts4KOg8CHmNyEsz/PH6a0B58/Zlz3jaZVhYE70yIkIcYvsvm1TdasYI/K
wLhUDlJopNC+g0N/rscE8v8hu5ACPT/avICpO05hVXpM2oAHWW0Bw8wqtFz2+QHYS39ebBlSkjkP
KVqeoFH30pOZctdIVqbwWYOY9rEyvua3T8LBJHBcTarc5rx2E79USBQCtoVjpkrWD8B/RgXJfRCD
Z1VuMyY5yohrYy8jDtlUZGa2g9O2NAJvesWI99/9UlWJVnlH3HfRsH1zSRHHSse//i+hRLGCtgEA
yZpkfjLr46g3WHhGPUrtYPsBSDQdT1570ansMmqLoNuoz/xERDWSa+azGEbyhk4cWKb3d/8jpC1k
pHJ3HDNYgdz2mjOIw5eXDL8tBYpEO1DjjIj/pc9YIPCMeDf9JYwvITlanFJlSCUCKHRAdYoqT3yM
nHrYtKBihU7uSh2ahIEyPayO3pzVSiLlVLfP8hE1Of+HsXn3HVotjth6A2R6ys7ccP3bwR2s/OBu
REufnvQHgbf+olXtkQJosmiaOlG8lXcoQBAT6RUgBhRrDNb6K7YFBjiXclgqlRjaGDH3r4EYbcLK
KpQyH7SDGlS1Sx97HA7Y8SDrI9KzjSXTTljt4pXCHdM0wk6hDSt895ucu0FJ8zfxQ/3t0QfaJNUQ
5SsKqOB6vF4S9eF36wUVYEiJSGb380mV/wcjjHNw1boSEa1ca9Hs+tfyGq4bFqOYMm7zNOz45l6O
eOMCzXJMqIOB/XKiwBMoiR7i+/dnAJacq20DYg5Yl86snakoUFNMAMRpLtSEaxgURqnEmzwSYfmZ
g7mtJa5SsHOUSRYmz0Mv7F0mXLVYPsmyjZMTBTvrXxJ9w35kBiEtmD9lT6pphYgCxUbgJsDjOtu8
ZEv208aj5S4rR9YxuPbSfpkXMDQefrpZh7MOyGbNCkZGHDwpWRM/z5QQfvW44QNhS+Vt0w/KufeY
qKtgLQek8h81b/oNUmDzAr7jrdh+B/F+YgJKHsIe9D1Zns6o+g+vLZfxA/3GT19tLJZpUUZLluNs
QmxynEuygEt+xmM9I2k7HaPMGinP3jGPgFKNgMSP+9356IQ6QYuKzoqpXelEwsApV8vnq1rMoEbx
F7FkxVY12s6VYhErYOv1BReDCwip/v0emZFWBXzVqvsTQMWfuzWfvQXUnWCaxWY4tJd+3QwwTnSH
21CDO1hsv+wbCHQ0LDd29iuw2XEJqmeHjJN4wILGPITdnTeJxmfBI0fDY94aHGwzdVbrnq/vz+d/
Z41V99JwRh72eS+KLZXY6fmHh/uQKboqkBvNkniQFdBrDI49zs+XvJeALDyxqm3nWKx4vWW7sTk6
ImDqvyvTUitkDf5GF8G2HEVFHdtOH/FFh+cHP6T2xpYjjmbzoHcmJ34dCkv42HtQJgahp4SaQo3i
B/HEPA5MMaKfNf/9AB6vgL+wuRRXyOJ1OxgFMGXhMTBmlS/Su5dEWXrVN45IR6VZ1owj2p6z9Nql
sigjPi3Dv3cRIzCUGQ7oXHxJp5bGYhvOaBFDuurmTVTPBsI7lcfz0g00vH5PlxBAyUy/OjXrWrqO
DfZnA8BmDhgHRgIcvUc9ohA8NRHJaD7kZbyFQOKdcdQV1vGdAJxut3NZlTvi24fQ7hs6Xx/3jvPz
n7j3SdT78/2cMPRrYEJp+T+ainZIxCC+KRXXG4i8ryNo/VrS+Pm18ltcOVkSOP3tZHjt0J0XAU5i
tQDgeXjgcj/76kzFPmegKKqKeDuv9ONjNrNF62uYqE2av3Qy2OVtevh41w7hxSgz0cm9rXlVimTa
ZwhIhzfh/Uyk1gjPNBQmv0LqE+tA+Imv/c7GMSs+GyWETBZn/h9OyL8rw+rA9hMU/KRtj8zjNeoi
vmOjfRvDSPxB5rx5oaIyfkT4nEycSXEfsdtqClhwPtwKEmFFGSa3frXRRahIylWcxIi19GzQIOAI
tEMgRUofw7IF/lmUTBz+dmlvkt10IGYYXX1EIituWvmnec/8PFDAgVffg6K0AnTVQGGy12BKPpu1
NlYCjKArWPvLIliThDLMJv9EqqpTVYG9Nr0T9C40z4qlSVX31hgslZmzEZM+VQt/lThU4HSqT8cS
gS7y+hh2kWqi4ktAYleDbwu5+kCjz3g5q0ct1lS4j8zlPMAo6B1JN5i9ymrBFg7gnVkRmXwDy8L4
Q5iQnNvz+78pY4HoJDLnUw0eZBlq8ip53/54/cH8InHncYKuSZYvwwAwqj4ro0AlYtEmDCck+8mO
+LsPh9Z9Hbh10WuWcOr7t+FHv10leLjYPyz7kL/u+F1Eaq9/EucSwQC7IDVJX1ZxtnrZi9/L8J4o
iKdsdBJLTcF2opT0q4VIa7A2uR2ADzMCtwfNQbzNCgNfA+ZzVaJQerBdblQR5EiBUXsnBikksIRz
bCQBoGCj4mJf/bmOLE8CE18u/BVZUay0QC66g8JaiAUC+r2Eu5jqC7HQFzDSrEsCddWnC7gZbCdF
TtID56bEd8Q1Mg7R+cXvWSgPTwH131I0235K7wRTRJ7V6X0tljLPjWNAuzYMmbn9fjsLNj09LoDW
h70mvchm4D8qdq53Ex6hVNs/oDgePfLS/zXyfF0uZVHFU9/+jzBRdutYw4m440zYCfwX2MWl2Xug
4PgScdILqOEk+y88QPDyhIfBjf6RFIiD/IEUMbpmJPLokYJoOrfQOTHSEUBFgNm4p88GoqaB8L4M
JtqTMkUGavkAUwfKxsXY9ldEAz0fbK7NC+WMODV4mfcKSVRG16sYpvxHjer7ouJTJ9VYORHtvdYI
nldVXGA1F7diRFSimQvprkoc/QCjsn0bQ9OUHh+0BnaORPeHOmN+V2+GgeBJlClXrzXskg7FmIKg
Bb65jw1vGty/lJKAJ6Mx374cGOwVK2cskgIXr/zBbxXdKXzbIaQ/zAdifm+8CvYV5jJxKzzP6tw3
Bx9j49weMNyMWqg4BGJqtWkqLU3PY4pZfVtWzgqsB8JjPx2SqNw7kAN13+IgLWvULZ/hzjS3BVAS
Ka0oapHxjxUhxHT82fZRLPxsve7WY80bF7p/mDlWlQVn2YJIpNRHGoy1EZo2z87uS8c2HEENiOdN
tQzEzTg7YfKyPoWlwIrbAlbFjzkpcX/6zMaWB2yEaJlE8vetRJh6bhoJVy8Do2HDpA9eherrDtc1
32lytnN36s/uzoONirZ41JcoKhz7yRxw1ICxrpWUQH+3LtcwnPBfYkyh3IrSCocz36763XbaYjPB
cuYrwN+R2MjEleizFzjinpiACMbhWL05smWVOD+3qG20quHY3SdXZGby35USiFczG3feAqC9UXxo
JMoOootgYQJ6Rxopkcw52RLSZyiNPPa0NN4h16oTQRANzii3jYuSvp5xZufeo/RZ09tmuanWDULR
7MjMTBJV50W4oErpTXiCpYiSXQFK8fjbsN3E9uRUCM8KHq6+TVGzHioJOlBwDasin+jLccjpsXK9
vvPdPEXGS37j8dy2BRBE/XqoKIEEU4XzbKEddJZFyHT/i0wbAwK3SZ+bgEfHPSsjvL+eA6QKHbZK
Y/vsYwrth0QmiUcjSWeSqV6hAuZ6Ft/0G0OACxIPFKleC/IUA798YD2pZGZAIqJ9j6AK5UnXkS0s
MsrRNWv5TVSd2C/8OJ0eeXr+lzxt1NuaRGze1oGbNUTfPgOuzoZ5QUCi7BXmpJLvkRjoHB2MdZky
eZm3IUU+8n/gc4k/F8lsol0D2HMhPy6d+cT+wiPcxskkJPv8EP7jjtS/B0yyZhOP1bfVxFHfZ0l0
aOUR87r+casbqrcivl5hrDSBuAG2boDLcm9+48QqA9SqWTvrgr+6/nl/aeeFg2LfxrPHxlcI8xBD
vV1paJ6OMcYoDHxk72+a+sdicIQhqki7Fiz54K2+lM+2dHyH1SWOTrTc6549kZJxxIY7kf2OXftM
NQocW0Gz3lS6MmyNIbZe8h86zfacm3dq++GJ0bsue1R2HxeaXTRpwrh3gBm9LwhJScLnzrGO/5Pw
hn/DD/RRAuGdJekxqzTvfksHEv/BzPdwEo1w1zd2TRZ7yMlw3BVBmDD4e9yg4KUVESPnSB2ey/h9
SUdOAnklR/w1n3SIfMXpGNpBi41UP8cZlRm0uZhr2IGq2YW9kwvfRwyeIaOs598uAxL10PhGHEew
Ip0OOqKctyopSL7TEh0A1j1o2en25anoc+4IrdYAdl53hnWsvjPM/FIYZCdVarxM6SzJdaXZnlC3
EoG1/T1y16d2QlryzI/E8CaO/uZcijZqPX2Fb82TLgmDI19DsrYdqh/L/Xx4p/CbGJaZNVcXHOgn
F+qYSe+5EeSSUprNck51NWWGnlHDJBC7IQ19Ogbx78GrT586UvVVHP6IO25tjdbhGS4sq66Md+Cy
8WsX4aHOIQmx80TADlfbl2/8DB7KwvtGHYCc1lAEHVvN/9U20rqiJWtA7lmRXl/AF7qj8b4BeYpO
pPll7gLlYXgLeKRvjq/E38zST8v5GerJm24H74jGl8b5Awf/wdwIPaxkjkCb6eRLtJ4ZpD2tmLyP
vrW9TlH6a12+LK692qpqynhMcl+igXoLyJurhgsaTStb2ekgs5VcZfCjQyoqY1EOKy+koe6ItvhI
WIrzbfCDV56/HcnA2mzqMgGumvrZSVgKjSIIAzq6gS1lTWUbdx86T40pQ8NSrK872k0i27S+1WLi
oTrObKi0m3Qs8/gPjTB7ogzcFZA5wymg5/IDT3+UnmuVhnVQm7e/b4Gw1iJUf6868K4S0PhcRUDl
d4/zD/ZJrhfefPPv5vAR4QZq9Yk8V2kX5gv357OQgx5sLG1tdIw4BbPdb5DnLp9KNPrEfgJ/dkXd
skojz0CzP7n4bf/wOw7EDM6Pi1TvqFepiySVbiVBAFVkDqud/PN5QEviJqEjZijOyu9ZbEKSut4w
PmdQM+Pt93Ro0y/OolntppmvvYgvA1mdpUwV39KeJfM/KwSvuqNRcLw1/VuK26CL6+OAuxx+w9Rz
QIn7O2EqDIJ+I6vyUT8VZouzeowhGUIfIQdh0ekSHBOVJCIBIyUnFj5tS7ETLGwQmSG+4tZWrPPb
l1Ve4FHq5dq6Y+EexrKmSVAA43EMTnvNQrLRkTJRVV0NadT1rTW44X4fkoodapCyz7QkMT12f4PQ
a6iCH5bWf2rCiaFy6l3u4wltZAIKo6kOw0Q60sG67Wlk1leeii8cLaGfriGb4T4oLFb07n3fEE37
n4m58JtnG4Kan0Wa5guRGdiAfhEyguYsrB8eI2apoItIASOjYZ84KC3jw5awKpvgLG9n5HLwu4wB
ugRNB8a9yQdm/8gRAuNOvd80TEo9X+8PXoHeRfSp5PRTojBsXhRMy9PyNezEBIiM5xhdjJi6fvVv
PmVc1+uI0l1UeGbyO7KTzWkymnhp+LCZNy+IfXZ3qTPeAgJU/1tZMt1X8JPoijRXGrgWOkvXxaMn
DoNUIDGzy6UrY/qtmFWezbe+/0b9xUdva9fPxzJYdSLcQINyiy311w7E/Ghat5wauSiU3LpVXnAU
23iefwxQjHcMSsRlXn5ZYxzPgQ8f72o97GOlxjcr5lrL4RfK1Vuita7eDhlWL2DEnKbmUEv0lRil
KHzHcf1IgDkxhNkhfP5E/QCqeCR+wL8qeCvx64r/yu2EOA9xPb04DMvjGpPp37YPf0dRBGO7vASL
RqZCgFQoOZeQNa8leM9AvIK/5Hw8+oSaV59yyv4yq/j5aPOv7IYKVk9+gsTbSca6PHAt1ZgbgElE
gb7r5UqMFiX9CNlnkR5VWcNQ9d6rjLb0DEGdVYGIqbDFeJGXU+eO5Pj7uAhbLvn5t/A88lhTn73N
KrRD+DwezddHoVim+kCEo5bdxVLMQuLah1ED4VCKDOHjltOX7ueMXJysiSmukZyI1eiY9OOzGktC
qQ/mq+X9Zax+7dCFDQ//YpyU5AmnHomVAOn7N7Mv2yFpROToOGwKlgV4Cvnjq+sQeNmMM/5FB3iv
F9D7F3MPOL4XZetkgLtb4SGu2U4RuLke9XhWdV8AiT1gbdP2NVGjPfpH7Atck63XG2gu4JmxkIHa
HWp4go8caLJiWZmNal2o+jrV5WWhrTcQw5dI4uKsoquQlYMO44pwprMlmMtmfNGdE65v1RT0KP+f
ut0dawxZdC9uW8b+z3wspi/9TGVw5Itozcismh5rUIAT9rXgCUvUijV+SqU7LvZCAkV0sdcQNMEq
K4qmKA7al8BAkdM6rRpVDQTk3mCDNPbWL6f+FQfLOvKfKVBm7mu7CGHCSnnwzDUlNR7Gmfaau3yh
0UPnSSlMxutgMfQoD7qmLkGJB+r5VuZm2KCQHJOdZyrXxZXmMVuQdjNTuvLzSahNuNyJyAA0CjwH
PDCL1X9o/bZnSokc8/2SYzb1PZm9QR5d1l8qiiKhtuCzAljC3EqKmA8OLPAm7f/WCFPK+Ays0Imn
FUUAVOcOqTlpwWKYXsMh45LJsQy2dwUlMBaQdgfw7spVJIcf2LDeNtDlQYiHgWo0KmNBRHmWMZPI
U3mvKCwujEzYJDz+orV0AhqUAU07Y8Vg1Wd9fA2Cw4VHA2H41eoM3f7r9KM4wrhnL1UQXRMU1gMd
OslgVZAjSynjUt69cVjPjxvgIJ6XAq0T0lz5g2+UPq5bbBXCVlGU8TIWS7zv7aniRo10X4YenkyT
xHk0l2+zIN7FXGEcNxxhoQli5MrNV65+aWsL1WwmLDszv4zkol4Qo3shQovrn8DmnD1855ttBc+l
Nss08FL54Tlw3WWxHUSKupfoTU5l4P6oEk73vffO7wir8zSSZReYUuaQ//BIHHFPhSvNEyPVjPze
QXZ2qkVU7KZ+xrVk+BsYToHrYhz+sOxSKksKDL9ZFzHVhxoEaaj5v8Kpx1bRL0pFzTLOJpguIrhV
DV6RaHxbQcSnBxRt+QwAAk9enhmOKCeyp8HmAn9573UcqyDnH/6zRK5CNkIgacWLgp8TGyoRRk1/
YwnYYU7ZFOlCeyr2UFpQuMNhMpHK3UzMIMJPQ1ij/GR7dwULZilUOlGs+Kq2l2BTdDNX4NWrvIqU
+qbNerqd8TC42/i9w2dXfKZY1L3BvuO/mXNcWtNuqUUby8Uzc9zNBO9+65An1oRu1YOJ5fbaIUQz
zRQUGQ/3FX8PrfOZM7Chg4Pn3r6ZwReco095BG+7oLIR+9AVySN3bWBfb5qde/ovkPO28pSzH2QM
JaUxPhfdiWW/MbIyAZI0X8hxNJ5iMBrAJi/O9VL8uip77jjKotrJyA9gvjOWMnTlnE+YBORKBxfP
vVxIE7yHAkN08lUx7baIMolY4HX74lrWndKneBIct1+VvMxOEhNOtg/KY4kT33RCikqc1vBij1Rr
SxaNMWCsfIUibZvO0sQx8ADBUB1KC8YPx6lmDX3hJzCC2wUF+fJsO8YdkKxiE2s/AWsBKHM+jTKG
5AI54pxyROb0l6ByOjv3hu9WY7jMTJVKdmaCCjdAposHPxgKebYJ/rUXK1gH7eWA5acXi71/Lo2I
MEXhg1xxO6+Mg34qXFa9xQAd3DFSih5r47X3pp93ngk65GmZD2oyJLKC1+JHf78RVJvm7W+tbHQp
L0w698HaHBIPzw8BJPGWJJcG1wyoYT0yOmLe5scz+1WvMGc3F2dNaK+i+StcEG0UJORoQNEt9gy8
nA4YkBY2aKTMkoUyYRigBeTpawXx9n6cA+7+5mkyQ26UZAGxVAHBvkAOq88DzOI5i4pabjFulsqV
aWpJ3IZV1M708b3djeMysQeGKtN2jyA2a6+AII56RqgpodzCKqTWEKZ8XB5WDRtFNqTXY2+qqkMC
BfLt+wbd/yc9qSswucqe8IOE1fTtsrXWBCJLzznhq597NwB3LfUoo4M4DG3jINsADIOliGGYrQu6
IqzXYc7lOs0nC/j4JmWL360Gler+vFueyyHDw/VMd18NQjxN/6vw0nfKT336DoLKNc9hLamyNUrE
6nfc47o1do6gh8gMohx8h15Lb55/NwjRYjNN1sa/PejF3wyez7q2BtTxWNRnz42pf5qWLXejcTP/
9JiKU/D2SXs+KMG0ay6djg0Hb0KyL389D3YdvrMY8CyRA3IFdBG2PujBsX54O3AU0aSQkppGVMWy
kBmdz5aISIcy419zbuvWMR5B7JYXMutlmxiwIEZO8lArqCgToThAjFFqOFOMfP/+vd2oKPKJhoEG
10CUIRe/rGTgjhkL7odqRTI075okXNKEB7c2hHtNd5oonaNpQsd4bVoY+KHgo5eaJ9js9ThdbQd7
g+UCOVvlEwdVIW6aAgIODNlPUX4RMDM458YvhAKQZl52pzglfUyVMpmK/FBgyWO8sJGonjPayTPw
zgFb9r8QoTJGH6Yag4NWc1V7E1ZIDA8xC4RULGNhxW9gtFgitcNTjU2uG9iK5lkY1GT4A+/4pUPK
cbgUJ9fL/BWe9RECfiPoDIfNd5juOZpJnWSc2rEAR/zFTpxQMaYHl7tFsyyf8egc+yQrk5WY5Or1
o62ge+oNC5LUiN3a+m56rDlNyFaPSLaA7Qomy2D5AICzzH2/IrBjnor/zxmkF5JL3+ZKvHUk8cj2
dmIhoQgvJxszCPLHrBfkpJzzMBJ8V/6VNVqbg9sq7C4vcQxKcVE7WugKAMT8SOUwfcyyNWt8RHsI
03bhQ0Lpqsrg6TJAoRzUlofkoU48AID9QBBjexmzgEoHM4gQyQCHFRfLOcmGByO/iSFrZIY1cDA3
SMEf/ZHY5al53cCOZHoxoO/BJy/Z6jmXwU/cl8ewgDw9dsqdNWe7tqNDu2BEtxUfafgP/YVgzaxl
wUMU9ueJiercxqV40xFyCJmS/1RXH1SPbQaNKj6CDlPOVQa8oyrAzaBckaMcZoouoCNOJcBDhgTl
fIKkrLHebS55hsPzxtx/jE+VTN9+J4p8qkAS6gkg1+n1CjHwWiQr03fHp/CRtA2nhr5CeAOxdip7
HX/Vm6lXtkZyIZGbLXLcMqwL0HjmWq7I9utYGO6oAvWABnoa7PBtDpLCdN0CzKlqSdInEwjuOTla
eJfrKI6wJb+0Ef/nDmF5diTbL79MzQu8Fti4OXi6Jyb9cpPDOXECyBxHuxR8I1q8qPzs/fr9kBAG
BTqGb9oTS4ZsBtjNNKO5RfnIJHuwABDyva4fE1I4+7atiC7KoqpCgRdGZ1H9Laf/SPYZPqDGGp5o
Lx9PjEl9DtjnI+Qlsokg2cpnJJ5UwwosO70BF4wImEoaqspP0QN9C8d/HzYNcSFrfq9TMBhREr+A
7nv5jJ91XkbcXcZMEptC0LTLosYJGEc/0NFMmdDUCvMoyHdtSuTKTQWkYPztdjHhCGtLDQlrl7x/
PorUn8hItV4mldQjDmy4t7y9Gogdohuj7dzESxm8aA3/+bu+39LVmo0EJLo3G3lEhyirm2WSwL28
q580PVsHnthvlMwuaf4qWGKooT1GzGWF3QyIRL2FY+hOEM0KHPs3YyG7mHpMu1DwXSwFKqcgAmDV
4Y4GWuk0EBI6onVGtYEzYHEi8HK7F6lrFvTVGdpcolfjNZj932RBEDTMMyVus7UoMhTlfb4zt1yn
/03KH3VjbuezdeUAKOZATNTSqJksL9BFtGYjTlWZP8vQlWM19BIFNNUUFEuirtQK3MYxo5KuFUdE
ICuKLBhXTRBb0GFGcQNlQrws34Lw0UEkYVI/sW6RBC5Y/7B4XJFhDknKYkzR671AUK5Pr1qjJG7U
sgz3ad9tP7BHhWzvsrOcU/GZcZP4bXxrE1WA+dHH3MteA415AeLdPQl2YXwgzcxaz7p/iaLtTWqK
46cPYjiNlEY3dSlu82RHvTMbAWRdkkFpEqDHwaXH1HRKNQtqH11c3/zML4zQrhoK3QAcN9F8a5Fi
Xak3GUQvrj3NVLw/NwNBY4QCm0idV/MfCooTm4kS9x18Ikv2EZ+b4SWTQfAodh8RcmqegZX43M6n
KBTGiRTBru+P+2ILwcntiHcU5Zkx64spNgd5cJQyBz81MjgOZMTaIxQZiQ7qjSxp0BqovNlu9pD6
/AJoJdKdENFBcKaZ+EWMjktOZ5ENZ9WN9Ts33SkJB/P2TZVxDztubvNhx63W2QLMYlv0INCwSQkL
vFDR+z3IkpveIOeCjTSm2+nRlLngKAzkCX6gsAb5DJYaUsEFkhSMQU6S30KZKLTI/opHQc8jWYdQ
CrDMuggDJAJKq1ATZY7UtDooNx9ZZCRaUtvcfIyQ7xP1kwZfeZcQX4zcBrmKWOpofqLk9tL0FtwX
H41QjVp7YGhPC9Y4HPVQMqjmrPVl0rnEj6d7MWwmgT8JYs/B2EuhM546Ela6+VUxh8KlPjyLexnz
LopvkgX97lzT+AxJd7RcKULO85WU1mW45Bh64ksh/Wd1bewQHfZxPeOYUdJERuipn438eLYRO9Qg
xBTEa4LUj8S8MDuCBipDCUGcCXnzn0cfqylzKg3DCDFPSrhQ5qesf/Z1ywczpMtY8YX+pkzoGOPZ
tfO1iKF6LnLSwDSUjLz5jZLYwDCSIibLrThy55qJqnef5DFh1inuyCw4WDMoPQi/P+heUpFZts4n
pDqbrzuq1go5wrKHOjsPZ7jnoHHmefJbgxY2wburspXxIAV1turxP3dWNtHYAoHmuPOPNf9ofyjm
rGXhK4sus7+rWGM7GeHJN2Bptv0Sv+nDDgtmZBy8MClvE393Q4xNnenPK7zNUQBBzK28tPMjDgi0
welpuMevcdm9UhD1E729jfuurGnbmXIFKp7ryOk/NEGtda/EHujvenBAc+wBL024x59hCRv4/OnP
qP7uMDXGSKEtNLHlKGUJsld64q1Kw0ZzLR8ipXLleMuvUJ6QsiZq2Oeh1DKh3zSuIOHIK9Pm4EgY
2dOfUgc3W/ta7ao634y0V6C68rgByREflHhpSPMvD78E3ss5WHQaGy37KwSq5A6cFvsJIxqH688y
oGKfWzYeByIhMAkfAcf/+DXyEct/Mxja2KnYfYGFsVNqT42wDsGl+T38hPDuuMY5RfZIYwroLPP+
v8l5PgnI96zYLuVYz5DE21/maQRP6me5AOfqOVn6UIN+yFHur7NNPS7ezL+JVVc929qzYS1ZtKIC
4PD2fUZ4dfvxGl/FXduqx6WrhMmXSFmMbrWWsLUeFCFQlwDLt1vS7VqULM72f3vCLG8QUn5QpZHE
Bb2lbZgamNnXhazpP7YGNXNYH9lsm84spIaEBX05XmoYp+ecsgTTT5M/ouxAMU5JdaTvNIlSJ7kR
cGXw/vPrLA60twqomzdLVHqRrb3mfmS5cAIV5FhO7nyRbBv9oPS/J2YPGQeJT4SjSzb84+ST0vAo
pYfa96nwIURvdrz8jX/2LiM8dK1KRgltuZBVVU20A9ctpEGQL7wLyHmrq39w1zeYCPurFfqVebti
wv94Bgjhr7kpUYPXFDG7Rz/zFtWJAJZvPArWLuYfrlW+v0KvgzFsVfLXq7bLwAt4jDp7FFM8rCcr
h9peAwV3a0yhwrRuszEHdg96oHcQ2xCFzFQ90w1bC6EpV+eRHvPhgjMcaXuZXlfnpu9yNH36x4TL
e4HUc6vbEUioGXO3TAq+7eq5fu0pWIG2rQdJ3/xGwNNk/4TbTxLBS1JfaF94oEdLMwEmcE7KdP6i
gB3KcNmhQrO7A648C+c/3Bk3EZBW5LRE7xRAzB/C5ZKyzv9ExonU7FbbXC5+csdTAUwvgpOqo9Ym
U1DdNL4ghn1hG17DQ7UCdaP+lIfjKiaOGnxAJ3yXA/SZi69jQsriQTWZtVvRaxieJmABfj52cueK
QFEzloMGSYYrggNvKE3ErLvQA5SFHRaOCDNPZ4o4uzpAu2rTKw42VDu+vsuNP19nufD5TT2yQO6k
2LxmPrewgIfOm4DbVAINyL0REfc+usOTSA9D1ndhstnhTyZ+g6eP+QccqxM94BePMg8udVnz88jW
ZCmuwvAk9tFttRL944j4N25Stbz+FSEMl2SzxwokJjCGQW+xmmJacZob+BNrJC13F2WUDQFLklnD
wd0shXG24tvhal7lkdIQyL+HO7wiaJMbJVQh/lYp5f9VaiHESZul2NSFOoFDyWeSqbXBac5CDHnR
TsyUnX2pDDJL+S3mrhcF3oLhZ63uJUH5EBeXKnBKJB/4jG4Vys3Usd+HfX8RTU3W/XQrydFx7dYj
cIc/Pg3e+4fDOG2aghHSwbd5d68d7W021+kiUVGg+IPAhGW74Pbt3NsVJoo3Mdc2IVLumqx+Z+tE
EHyee95rU0xTM4t1zt3beVE0M5DCuAj1/a2EFvSoh/uNbR4YqOpWovStVl/phsCedKP330XycDA9
Js61ajFyxDy39QXoBX4mVzywI1om3WHU++USOeL3mH6VM1hN3UYMEPcs14omkjNRxPCiC1JHVgPV
QZ2HZK4vnRP3HKf7YtXKmGPWhaVZIAzSLPVwE24SXl7bZMAHhytA1se+TVb/aFpsuRkW+bODDciq
DjnLBYaJi0BKikrUJrzn4to9EXP093sJ+8nGCBX8EsRWixXBrB9UMprczoyYEE3A++9xA7sUgB9o
Eu/r4oWzXErp9HBTFAdAb43w/ZAGBn8mEbbOvPuVoigHYVSasro8hEk58aTHgXv/A+iii8Cts8/m
WrhpxVrm52WP9BgfbhBvDiiDkagjbY0g8Sb+cB0AWpKMrhk2KoOVJsPlnncMA4QLTnRqh9IQ4vrp
Ebz1bkuPqXoR0qMqSTO2I4gJMQ/+7EVEGL9ZrNYpNjNC6gZV7aMePBAZXnfBqgXjvRnVc5rOiquS
Pbm/tITD7KqJn0aaclNNSX7ADANYbkdZZnEh26ppN6jT2Myy2McJsm5miXfSazAFYhdP+C6wND9o
tKkctQwvlpWcWiqwZoTrvzJMCNrPjhjZht6pyiSUw1p8vlFJ6Jimx8leyCMuim5vXQk+YpxxBYLm
SkscDyLsnzG8XJrf2RK4Ruqm43LgRleBoT8Yj9dJ4JaQcEsAXxHuBZKjdKmoqCogMX2WvmPe3xJO
4Wp2ssKQp30sMunnAjMcw/3Em0fGsbh1iMUF/zFrlNQlL6YZS71lcG5yz9hJHwYIz9G2IkGZ0jWe
18Rj+K6YdVqTD0embexn9PYY+vJIq/t5XivDvyycN8y6yBN6DFjtT4ChrCZAw29yKv50AXlQzfI1
J+a6HxiEzgP0JwcT6dQe/g4xrx4DqMoWGAH7Rl74hBVbepCKQmNRLIgiGnRXa+gLObFP7ZhYkQHf
kGJ/PTeEdqddRxOsHnMJ5k+D54tvgk3p8Lph3H3uQhLO8ZycytejRALU/ehl/UFNXeY960keZztU
zG692KTE6AWgUFtwHuk7RR4XvRb3D+/GhWAcpkcdRdMVQF0EXSc8ub00mVIgs1ym00p7cEcsyS59
yKXyTnJKOSohcdeZMr3DiV/NRkvw0GotLSn05d8YDORunC0sLwkh9E0jCs/pqTy/qdBmr4HAko3S
X4jpeyXGG99Oiq3eGueD+5XHZixZJcU+oc1LMKPRhNPis1/XgGyqhPqrzAlIfRkohnFzG2Qog2zQ
aVbF702FOWZtxuOO0deysy0uYrppiBsGgT7ccQTO4nB8kBxgVuIS52dUrW4HAdESV9wCOdKNYs6P
yaPfTM9WMDj4nFtqWZdywHfXKZOzZy2vUy+Jv2dvUZtoiA8+VAnaYvHLyMV+qcmxOocG7RZuQwQe
bCX0TneFDocaVYgeDqoqgBCL9K7nlyemAAifkM5g22dkQFRx0+q59yvtB6kJ8iiS6Y0C9uc6RDYl
sGWQqOn79Rh3NyyzsBU3b6p0C0xOqMbwlC8kF21wF5KtcjKJFLXmDVnY8cQfMJdYfYLAFIC0RZvy
8GvvOUsETYNJLS48w4GU46zjbWWbS8NR6NC4RvInT0k8+S9iEkfpzExnJhFCvkRpikBh4pVyfqPP
wGXDu3BzLFzZwqJnHBCmuASurenHx5F0mTM38eTQAKhorA00H1HjBRYQueSecStzZqY49sB2hGaX
P8XXEF3CeHI3a/mg2ji4NrGrWquIJ69uQUNANeDhHN8Aihl3XuRRJ5/7LTJ5/JXPMPQtczOyiEjq
kFu2FM1JoEP3i4Z+EVvDqyb+TP8Yyz+UzlbYYB1zdkqlpQGNHrRXry6mkRO/JY26IedqRjvwgsIJ
lzCMskXAdAUFu62E0RLRNzkDPMV14KhthRmptjgS+FRciO2i+xZWVDGGVWajnX5f7OFzSOZYLhWl
8Al0wLnp0WWE1z88jg3wkojoCGm8q28JqfZOTS6kSGGyEkd+Pfhc13bGCLqQgb1M0iBGDaJvfpVC
hsuBV740xGyfTC1kS+jU79G3d3OZC0NFvvG/f6sa/TjEFw2oFuOFjfA9H7s7aCSL4JS0bhkNLA6X
pT6X8+UhyybQqWR85SBIPH5I11tExmj3ev9vlon3YGtaO8Wfg5xmkaaQI0qQjH7aU5AkL1pXCNEL
BNGxB8/dOAQeyEFbRbeTCmcyG9zO30cKO+dRPaYtX/e9+WosfZSBPlxQBc6SURnNVSB8falPXxDy
NzBiDal9O6Xk82eUT8uuJCEy0fSRdIinKCiZn4G3SAFO7vIH0C+ZZmWlM/aL9xZtrxQ4pIf5/Ewi
PZKebFda5D83XNZatLLdYrxHDIwMPVV/wT+NjLfNz+X2Po2nIJOEsbSZDsQd9MVg16rn15jk+DPK
QUegFr41uT2/N6SAJUS6h2V3sOxJrHvsU0ttNVzaiVQCDWw0ZfKc4RODUCfiCUoYGeFcUfFfc6XT
D3pb0fvGH3GVi+oWBVkL6vVjnRgSc22RoqEETCQYVahnmT64aBtFU3WfBL7jPUpOFBSm1ZUawLll
gM+K+Ir/Qv51MQMj8Dg5v22Zak9ugstq8lo++eIJIqsWoaDju3D/+hA+R5Z8m59Vo+fads6Rmu9h
JZch3ZvSKUGo27gYIkzEB5K1UAVh3Kl08tmRbceRP4gAaoMnwzAFexLiXQJB4uQI5+t7+1zTqiBr
jx+1M8SU6RHdTPUuYFheyQLLdjcXJexyUhG3HEmVhiEQa/axXJl5exjcotgXr4+1oHnx9zlZFSzs
ID+SZVmkCPogYEUUQAZhJ6jXqxY4HuJq6TREp+XyP/qUdPVeMDPJZWEMrmg6c0rsk4h+9ZFXwIRj
senJiVUm31keHyOj9fbsB6xP+3r7XwjPRmpsKBv+QIyUiPuqBILFuIMOeOgU9psT6mY97nUyhUfz
x/jM97GVKTSVpKbt3BICjcptM3sn06BWDUeEzFWEXh18Sp/M8F8+QK005KEKKZJmS1Q5vF/arrIJ
ZzlAo+y72k9H+GkWg2wI7GBzmD2iuWP7Eo2GTlTrj1w/Xt7Dfb1mnrgkohw6OvxavHZaFJiLMsEn
R8i62yCcW/Rk5kgXMyd8nBoUH0bozMRc4Srd7rsybxcwHC0N6iZDwm3SHmBC1x/RVlEYWTgo8Tot
RzkL3L3OSG4hcOCKSpRHpmGX6Ug3wqI63N7tT1YTS6tz4FuQNy2k3FZYXRZ2o5E1HbCJ42+s5+T+
bCTtmomPaHCIoxAz/sb/+cHTS4wOpvPS+YR+EIhF1ubdtQzGVfU+fDXshd8ufGGqL69Tei7sNu2r
FZ1p2fCC2xnDloXnlGLsAWw/cELMMHqG+ef+F9uXa/j/8V4EfDWlhDMXDkIWniHg7aJ4GyDSUxnz
rk57c2kKWqfaf0/ja/kfFW1qt5WwbFdQ619mXboTopiFldE/eHuWsxcoBeixwsXsxYSKuswT7DxV
DCLZXczZqam+lNwxDLPELyVRfoGQshh04txTo30IBxAI/X9SJ74TiAK67BiK3/es3lpbhxuFphtu
XA/1SZaRim1CZ/vN8qqtkADAMS+Uw7lf6faUe04X4nQ0/S4PeuE+OXfzKoYxP1qU27Kc3V35OpvV
Tv93MIphsB6qavjbHom44BdEa6rfL22nW1uC0Wbx/sodnbq3uNa88A/qWEsBNJTfuHrptrL8hjFW
l+QJqDFBLdk6taIg/5dVoTimGz5IgDKixVtV03ZnVL/OUbDHbjkiJ5ee8MG+QDFT6Qbfgyd/0qOB
xJ86cYNX2axziqlp4P2/gID42R8hPnde4SbkKJwmI8dOVVfTNJY0DInRORYDRkX6ZcW0jmhF1S4o
xwvImuQULU1BZn8iBWXtfP6GuoIVc40D9MmXwKqybe1XzCDy5RCPCCw2Rxb4Bv6zxaL3Pcom/SV/
XAQIkqh82urUqRPY9eRE9olHF1Mt/OueZe+gecTHyoduCM75t8v80cslTPtT62SCojctcTRHUzOk
yQgB5pvK1aSc8TzfwQO0fCd/DrTtM1tbKEg6OaAq0HbSUQ9qABjmlcNTVqbObUia9CXxDUXA7uFb
d7hGpKf+nw9eSiFnNMZAaPznAK4dOWjLJTXPi/WnzLgep09E1ZkiRIIaZvtEPukSXY98h+9OA35B
qIpD7phtSpnWBU1JzwDcSfOfxP3UqCSYNuK6/KLsm77NeZpbo5FUFI3dS2GrVnAJsH/fsJPlBmMd
jcKs/yNXpqxDi5Dmr9mNZ7/42q2FZuQAHqHlSKeG2myG+SakjaCsIHkX3RseE6ldcJ5qU5mAF+It
ByvR38Kd0BNOBeZXZY35IRDEqKuZpk4Bn4monQo/yCf2cibOt0tDNQob3OnKBQYCtgzDl3CtxhHr
YAqGjFhtMUd0f2F56yHBfq/WoNuVATeyWjBpXk3iAZlV/isTqnqxcXdaE4DhGPyW6F4h7LWJSVkv
Awk8X7/2U8S0t0DnXjicLnGi9454NxYxWcRiR/Iutdzf8gP4Bx7Evnz6Lth3+7dPUxfZ8UEcZZFE
+W54jneKgbG0kzwSMyWNZLyhAAYe+i7cEUo4ywGV3RkCbMx7vDVIE9ySO8x48ynNRFhdwVSrGBep
MR3OY6raAf+5c5EqAFmGfoH9ceApQqVI/CnLL9TjOv9JmeICvrnhocmYMRZCdVRMytIg8W9LEc0A
Ut4m/xOmkSw0O7NGyQrJDz3kuB6fzG5GbCV5gLGYVmJ8Dl0R7CPl0YxDYIATjAVNiC+oJpG0wJy2
9+GgtkC3nP10oP1nigr0mGtOpmb12gXQ0YsVbn5mzZlgFtHZ8wJbw7JPQG/Lpl08DDet4DCEf/BL
OrWmJ6B+ZnNkIcHl+CqdI89aSrTjkR5rr5+Or4T0JoNMDHiA/8cZUkxmPiD8xZ5p94ku3C4+8ksq
KlB1NeQs9ZjJdVVnAzZlXnw2XPQovP6ZxhfLMj+P89wZaLfD0vd+SylMQNLIRhO5xJ/60Hg3/5yI
8kOoByWms9peuwkLPidgBfmeRHqLnGNa8gz2RBeeChIBcNYEpzGC2rLyMYfwlaCdl9ghg1X2+dkJ
G2KPi3xAswwvvhE8nv+t1VB8CJvn7cj6F7xRvwIoNkNLeaPkskf6Nav9l/iRCJcogJkD/KgZdG1r
8T2CPhbKNvhXrEvvpuLJshRfd4g1i7jyy9WPbTyBByblBV+eR9IcF7Pnty0/sq2C7iDOKqNjUSDX
2rVDilL2M9ryRaUU8X3OVSUyn/ZOrn6y8qvNysVX3gYI9SgCyShe5I70qeMAk44Qwh1PHRIOagNp
j1vC8AnkBFxziSlLPFEnlU3HTStKGfKx+pUQ43UbIuvp07PfFbNfJ77gBk/AtcXV45wDdxWJrzeD
gblEJbgcG6flo/WLAdqTUinU25FLkeNY5H+GQ7d9bsZjIvAFNYMmluwjT9G3y2R5EvZZMeLJ1kO/
PnW+k4wfDLPeeM7BmNse8eZo3IZ+JKLT7iDsMIJtSBiC4zajODa0WeCv7lb44zaLCfpvQ2ydVCHl
bXhMI2C3hvK+w4utJYYD3ZDFunC4hJY95j1YU5jW19sduQcFYO2FrmFPTTufuzxaBuBY36nzYOG2
D8w+UyiuR/Gjsg5ZwouS5Ndn3Qn1grSs4Lyu/REilocKQ1RtgMDI/Plft+jnX90mzt2PENxg1GRU
onm09DimRIZTs8gqsIcKPQjpoUJD19PC5lJefdhKJid6kjD59KojE/cLvat+JcQ24RHlxJAhK4Ho
+zoRZSkVa7N/2TDUADOcQ8kgvkiJfCeMRJ6jTUZqOB3EymFBsKCasahzEFC0pVwULyXagjGCeOE5
8KkpuC5Wtk/7RTrHABvZFDaBmiMteuZKeMwM0AoGv/1OblSCA7pMtdacDOHtS7HwzLlZfXVpZYK4
NClss0zJDMEt0KmZhJXDJtM5fVmgyTRJOJuF2FpRdodfNP0I/w/Je6haXFeIEIqRz5OdE4myME3c
QL1UP2Y5GuBOP0GatiyjWpkjKJK4ZZJuLdg7dHS4f4d7vL0l2/rcqe4Hx3sR39hNsJbxwPgzdecw
VsWNA+VPfQkgBXndVBMKoGlz6VubcUUAzKEwgcsab03d+0bgAQF7gvzQtx6sgSRyxCHQJiBks7Rg
RxDdPVaRIQ6vSQCsgmsyegUQGWO0hKa/bByp9YiHqOZ6Yw+AitresEpv/2bkNWTNV7hfMA4bnxib
9Bi1UyjWzzWfg3G4gtOdxrRxx8zOZZryfBLAX7umwUvXHkdaZ9bEQwfAAZHQw+QhpH8Z2wNg4TWl
B565v57FIc3MRxgP7u00HM7btiiGx+B4vEFWbK9CQ1MwWXZC4Rnsvr1aUmr528TgKwLCpOqOJvHr
+ZUdgQwRMnZrLrizqrJIC5lCW4ix96c569/+/z5ZLdVxc9NbQopffphskJ0IU+csoiyE8UlRIptF
yQlHNlj8eWE6SiuA6xHOWNbdAWOgNsqT9ccgRFlS5OD/x602C3Y0empsXzKEJf3NCx5rVE8G6NYm
CzmMdWdcl9w374Bs3Rtwgqtjs37/BWiGNyVUhsZHIHmM3RDbxOZkldjKBm3aWZsUnAPkFsgAC4Nm
3p1jh8wkWaaZa/oelr1lozlpxFJ8B+Ta/74F40TuWeqtXEcICXq7JPGgQ7MRHkXTNpfMnSZ4J6Mm
FYzZa16BAgmTPP8VF7YoXr6huWfhfMzlQaobzmBqO+2xUAnhmH59BGfLhQgsFUNZ+tbXJWiAFpnp
S2B/s7mA/bkVK/FPDi9Lg0tL0GzbxLRxEOs/NqRY5SNMckh1/M+fz8uqkuNg2D4RAoDTWMEcc5fG
w+ZdNXQlmONhKcBYQqTwILkC0UV2vgtYi/ii2vE9NIV6Mt121yOXdWJkJ/693kjyAWemu06XfAh8
Q3NKn/jChTTl4R6/WiQl3pHdU1mRn8W1uCrjKWdAXVO4qFbRBBZUZ9jpaOpHsresz7pXGAEorz3D
MbeR2WC4OkRyR8FMSX2QhqWqVTZguUXM7Q8Z2Nu6tAD416zBI/REVfi5zvQHAbNmnS5qnvi0n3lq
oe/jGe/VQlRt8Vefyq7PVY0nNkZ/8sDHWhUcqLpS7bPFc5c+0Gpn68jw4jIIw8ZMC9IRBd1RV1gr
lqWGJZDg2wWMnO/PXIs6vO40tWiRjv0+F4wgqjP8Hqw1KQI/TkWF+I5BElhuHtyd3D7V+EsTTbJx
Ig8xX4y0mRIN+x7fBba6H92iidZmuC7+6ZOj7kBEwE3vvJ6reNZTB7mO4nk73WbZw4tB6bPqY5cB
6pucttUv3eVnSPZkcqNqyrDl+d6ByXwRpCLXYxuqd4986WABftuzIHa1hHZV7IjucZjqrKuiCytk
YlA1E2xeDwNGo008m5mydkOdqH/BygLWuhOC8Ldtz4oc7a++h5EZFQw9+S4FnQsxPeDvOEmseHmt
XGUaIX3l+mhGs9QuQudG9XRzNJ5HpahIdLOF85ajgpz7RTIBX9KROfMt2bmjMOiI3A4adI+A0Pbd
YePFXtY4Gw2QKt7VgDoTz/DEoPkoklOMveQXGd8axLmyessDpz5Jdtnu1zGXprgF150oh/2V7Jjn
VpE/nDOXbYFdcxLxtEiPV6GdUehbiOETkkYeyR/dkjyd0lSGiDMfiO47zYs9vEg44+B+Dit0G8As
cGyBLj/3o5m2C5qAtmjVWQ8aDId2J+5plTE6YQRbB04MeZmU1+gY8koVzFGkBvLLw7fOlyIcclcd
YfUTXab3Xp+nMQoJSlEesDda+6y0eQo9EaOw7buoB8BNgkh6ReHeUqX0+7JCFKBywmyVilMHGFFu
1pbwSLowdo1/L8x3srb4jgQ02erf629jDUBh5YIImkk6dQvYDQOPSq/+jerwEexPsklF++u48L8g
kdiowFV9wKasZmQWDcFs7zUKRzzQIDRMppG/VbP4U51GYdE78gExruZdY3jrqHAUaGiUnpCKuhu+
QTZzUTFVg5oEvYAzYNzQJ8rvOCikCUVJXh2G25p6QZjw+s+cB5npX8XpebJ/87NjwZWJTI78B0u3
qB/V5RaOKTlUd0gqqi+jSFXdMkWSjgd7VK2kNczclPyf2VjkAwRsRD48UNgFam2Pj7q5vmzgyGZw
4sequmcyM43Bk0cZQKjpYiRqcp5CMhznaZqC+6YcuA/eDc8XSdqPbqiy+TlRr8hvQgSr8BzEKReN
D7sSfVxRINVG3HapEqnhJMW/E/ZNJ8tELZ0FBYiyPz3vDDZPrYUHZAvJ1QqpDxH/45EL5LEq1GqX
vhIaveRBJgBUGLWhSvtt6F9HZ5eyvbQ4uTnM/d5m6ORdfFEEcFwVOBYcEPKQvIz2utIOQL7mztKc
lb0UIAQy3eQ6f/yDt/p1oPMhEaTAGD6ni4RGRkAf02vi/q8OM5v7AkFYGJCNcgYAeL9RU+lZ5U4P
uhovAlWGTjnDxITYfdqn0UMRT3O4OX3az4RefldtU1VUtxqzb12duHBvGEblQmfNSmiXgTWtO2KP
QJ32ljUzRcnLwkqb2QjPto/zwNaIuXIsnw7F5HKoPC+d4VYLuXo4XsNkLHdwYohLmXMfecQMa6jR
sVFS5mGPIUf0OtjwqLHNOY0Tjj0pSF5725cqXdywwNLaR+fwHzAcwKQVoEWJfLo7F9V1Bziwheoe
riQNlxvvs/REapHInmIb8gq3oyhmdGXC2s7QP9ILrDmqGmXZVTsTG6+r7vxapcv8Ot3RtFb2eTl5
PYSxL+3yE09IfdqdznaEwl/Kmv6ajGegpKzGAWnBp5XfgpOaKhTkElP0Jty/p8U81AylsrqpQwtn
KWaarL3K41qNiiJ1uqVIKerXuq5ackb1l9DDh1a+e/CRaCPKrhVhA7DS2vqRudPNRyvefrgZOrt9
Lzhca7aDsSaql44D6pWNkxXYTgx6yTz9b4nzHhAr84t5zB8BU8D+BNhDdKCd9ZZiTsJLXSkNmvYj
GKgpoZWAwR6IIhtMLuBC2fTkHStJb8ZDBRtjA6suXVIdfkij5vQMcwrlZK6qbpznPEKzTK1c17nN
wCVCjvemzcY5jl4Z58Nw3fSssjuDBwAxcL4auTJgL8k+iiulzlYi8tPaoOqPoBmI1lC87SPaFZtL
/8ZzgopUq9lQvOSkQJJg7cfL+aAUHqUAPFc3G8YxFu2unS2ccxCXcct7ZALCIgTW6PSVs7W3ukGj
f1eTRXCh0DItw3Mg5loR8gIYWRP5dU0/1QxWCbs2GnVni70ysD56w74PWJ3Pvt1vHCOhBocEf3bC
t8kicmZnVZMyhOFtFU48RQOSaEbzxdvjEjV2//LY7dMQyEZfDakNI6Ld0m1Cxi/kJ2QutDpzDjSZ
OxaUA3xO4iSclou4f4owiY+9v5Eboo8VCR+Q3fVnCuA5nB0bKQzWZ8hx8mT26QIDINt4wy2q/3tp
D6gufx4ZiPYErKG7g8UtysSk2v9s1HX6ngH47DOKchEhmCmSjBzIsPGLcp+spgM+P1G4j6dErXcQ
7LMooG4HYBqEnR5lBw1wjkhFI10j3rnTJl1vrYoDXY7ENfjcu/PjRyhMzGFe4lNNhrI6J8eO9GsG
3yaZ+miI/yN50Hb5sC4VX1TSVFTd3SJNug9cWEbzWuQhpY+01tGL42NHu20eDgSBn5CoDzgn8g0U
w1/rPeXELUpKPmIPnAJnTZrdz0Uhabr6q1WNVStyJuavpgu4WStGGyuT4QD4skaB39U3HQQEhw8d
Gl7a8wWo0xtJK+6u13dU+W4lrTBR/tUbfyd27JbTWGFharNwJJT+0v3mUGMP7G3TlaUa0hHzKm/g
Y9kyYK6OhQoqFgHn7jaW0JuAJYxznl4CiGuSmIK7ZpjEgwW25J3AalvtbBIL4INtcz4fXV21L7uO
8jEMQe6vG/2+LBTYxGyyeRgL63+GGn86HfKOt8r/E0BkzDFCo89icyYvCL9DhW6s2lXzM+U/4QhL
dcsMvh2Dl0ZT5lO4Oqb2O3ufOQ3Kpwe1NsPlfX+gvjiuJYALpYdCqbfpE2b1L89P5KpqhBgaylfz
FUSU3TYrbY5se8eTQOVThMP6X9HFg2Hj+ONg7OTI0H3riYlSZeDeJN1gy0ceHl9+mHoZw15dRAGf
KPXY1Ssd8QYazt/e266LBrg2CPRNV43G8be7DbpuZNvVNrnGpXjYrvWf7+vyLvMJFmFOR5qljbD2
J2ba6G+B2WFZ44zC62e0CNXjGUC3ZB4FuMYN/7xHTZU50cZkAyVQaRAX9mo+Kz4OwsNjeRHRBcPw
YWNEylH3QbyjSxOvYV/xHIU7pwz/sSIGNuwxT52WKpKgBrtMTUaEH8MTT8TumnlEZ4ReycmZNmS1
YKJVE5VbQn8u1oGHgNlAgaF89aD9/TCvuhJmavLde/b8nlAtRJBzqlfTbtWpi2yb7GEeonnOQTp7
Uhew16xd3X4XBvva+1oTPRcv4B8Fb0H4qZEk9ML7BOkz8ti8I0C9hVdKBjD2SMlmCSXC29jfsf/V
IyGoKT+fmjVCbSn4vPHnSPYSystZRWx/UQlbN4w57uvxXDQNaBkRdWPP3DW4tx4fp9DAtvBKtlde
fYFxrzhivwqVe+dNwGs+fzUhi3uhcH80Q2s86A3x046XyCb1z1JUjl+33nywfe4R231dLF0FyZ2+
/h9/75DioJRnS1Cmk/Inh9atsqhy4Y/sQ/uHsN1MDopCbyL6O33kY2Sxi4QU8toikWsPl4VYJMQi
WIRKzTx759zu7rk998miDBtHPymuWnNcBqi/hdOU2SdGbWnoyk8MXAGa2Di+M81VwxLUfmbngeVN
/wy4MEzROLeX9PWNy3lJdAxDxP4Cd0HnbI86qeixFgaeKJOjDIDt6Eu75o2ZfHT7/I8z2AHL8UL3
8opJG4n1tsWgtTOcY977Ajt16EexuQt/EFVigNV17Fv0nSWAXveNov/92+2uI/4tBvZQT2ufvNkS
KtYz9lCTV7m0RjsJnr3mI6Jmy1z1xy3+TfM0O2DKSLY5ByLtSWYJx7PICaownseVxCEOiT+JJ/bb
J2ZYezYz+hxoXxoFPGH2Ej09UoA7EMFosgHiB41hNCrImoIaEaPStwPOgkM3Cuebc5VHgrQmfCqv
wur2Yyffpj7d3b9o/ta4oMvgr0f/LHmwJhw4PM486XzkLO98DFY4gofm9ZmG9R/pYjd4t1n6lF6P
hRDsA+Lkj46XPHebhEU4TM+x6Kvmvu2FyHcocIJWAv3yEUPZiSYCKPnhVga/0V61o3JOGvuuag7y
Y/zOt8Y3w/L4Mt28fWdcSJBSabHzsn5aDMMPVgnvvmzzwphmwArB7sDunYgIzDrcpdby5D7DovM/
n/x3R1QfCrBFDCebM0vwj+DghUBXdTj9LsOAcv1D9WRU1k0zueG47O0B+xIo/M79DV1qzXdZIAiI
c4mbVrv8++fI29ElC0N7P08d5mxpbjWCywntmxinnC/0J9lbwNEKZpOJ3DRkX8sgWu0UpeaueCUj
y/iQ0aaBdO35QOSvLdCIeKUEPkDYpIMc1+HVqCwzFQCgOL9rD9I8oTOvx0l3kgxVthAk5Qp33Lhh
HOjBVf8tm0Fev5XCY9GiirYeEckAksz0F3DLWs1VYQnx7GRbL5zZd7VUjt++eQGM64Pq/HztJE3V
HsLV+lxE4YUEQYP8DSWGolYtYoFHW2Nq3+EdVsy6KJF0wpy6SN6SP6xIJ1G8L7EGZEp5RWEDczgi
Jjb00hEGZbOYqLwY5/PVCLZK8ry6WcaMWLIGFAsRDDdDdbuN9xxdazT0I50a1F7p2GLzR7crBax1
OYlZTISd3IGRvxnlcUcVVcSMudx3aVe5LoIJtPMG7WKUk8VRkqXLL8K68LyOm7WlzLEC9ReBWtU3
WBJQVexIhVeE8DQBaZu2B4W7aiSNyfZ+cJPESiVuw7aZdhIicfXXyBVutSg/00yk4shl2tWryIla
VvUhnmDpX+6imHAOXzRiurNf1eiwqoydB99XL+zSqje2rSaA/tuTYwZM7z9iqUs+eaznyFi9vfMq
i4QgEJEj8TkZZ76nJRCJagP3QYbVpfrDt83ZURxLd13xv4VvF/mtFpInec7uRv+IL7PZlkMZQFqw
eZ14IeBykBjssBzkrphNhL2+DeOOPbhKdXaybls3/fyiI72kAwDDDdOHhtNFTlhiOzrEyCqKsLi3
7Ew33maUoIUk+9f6uLJEE1EyXDb0k8WU7Qo9gHw7EgypLd98J4V10huuSVnoMzv2R5FuvDtQVKnY
sKULVLDa0a+eyqOzi3B5MgDUEHNUtLxvW9c2EDATGgRbjJp/f7cAbrFyzBvGAsDoEN4SbSyjvNFk
oDApDI2l/FBKC4WVK0jqS5l27iZw7icCifkGVcXaYfhJt0mO4ff+Ip/zjfcUR8QwQZuMk5J9tEEf
UNNEdm2OlSaDkzTy9z5yiC88pbuZhc+6OGZR1NUB4Icmn7rZqEgorQAHsFwz0COi0TrITmEZv1v4
TR2gShFqGJexCwSsMVePlGI+MRaDb4UZztSzgsq2IDz4hYM0FVBMeYAvfKPuOR5lJcnpZLlJjxgL
AoV7vu8ZAjPCaGXNQCAQ004wv+YpQwmgNirYCsECKmQyJmnua1ozODbBT27U7XkdZ16gU4xW0mq4
OAFVLntuGMwQjzUWJVuC62q/Qv8CghaAEnlvPA1yZLLCLTEgm6Kocw0CIENDEQgBHMJXaA7e65EZ
s+Nnywr/lx/H6JqsMSCe0lAfOpcXBCw669ZhR1wmJyfqXcsy07JAyKpJvmG0dIHhwkC2RkPRUn9z
PvQvBTxc3vTMX6eRO/3ZKkqGgoI5XkrPNfPRjOzvlgCgj9/cwdJnKrDRiPytQsehMZN7LUQqNQBO
e5ufYwVb4meywTjXlZvghJuv0TKty23mCvKztIBlE92c6XLPrVKgyJuOkC6FOc5+ZEcacnwvbCB8
6uZpcmJs0WkEgZhst/VtYfs5YtZUpzo/4gk0UlNtln77AJ8IYziyl2QhwgxFGpN0pChvhn88BpsB
4EKn7vxxtVQb5SyiSSjgdUvsWB2QMDT6YCJUF8DTpokq3cgqo2mmk3YsHuqqnWXBKKMw602O74oF
g8Jkz0sl+QWBP9DQQo8fYyKjdjOq69q5aOgTGTIW3PTsqcPDVt2Q1j6IOm6zy88z7S3+T4KhMzGj
4e9ULtzluPaoXtDaOHNOQapiJDFc5gieLYeXQAdpe+XwpDxU5OfJwzpX4rL9j8bd/Ua9Ex1xrkOO
kVPvPUtkaOq0c9vGB2aQHLgak8iQjVZEN4WHtJ5H5BXdPIdkca/AOORE3blct7charuipPgeW39J
e5X2dCerAhABkKUJPAZWTN5csd5q1eTsQu5XrLOF8P0EH1R6535HIssuQPiORHKC81DbQjgWlRL5
kLFVd4d48VMoywqzgClZxcL7kJzEjJ06d4lg/cA35yYO6QBKPmsa7fdnZZqk1D85nbf46CZwBzut
1AuygsaFKgD1sd4/9jQyMOGcVma6+avUCWJtUbwOcBKcwzFZKBdiyUbqgwrtS8qpC0+PnhNbJEUD
QE7SyIzIbt/xynHHo7NVABu+KeJfePiv+d+nHCCkd5phYilKPumX/J5wl3CX/qerUu4MPrLsN9Bi
dDFCS1k1PhiKe67qkmQuGzDLnEoM0TGj3HWtu1M+q4h9o9ToFFC0vOoIDTj0MPn8AmoNTTgFu5EE
Rel0JUiB34AqYX+HnA040LD6ld4/gM5wbrB0v0RupzL/rQ2P86SFEKFufbOAslV5427W/WP1iaSZ
SoJp/klMWPmF6d3LZs1bs9cuxrZSKTQW8sGqgslmB0eDNd997M/BpBQRTQw91CtyYWu9jNyW825B
TE3st0wJFK/NjhRBHZ3VJpYvbYOP9akpPre48X+Yjb328dHtX2v99uE1DmB8ERUVJaW/4UXqQv5S
OiWvqWk58PugI+lZxwfBFjBf6/VtL09COwdbPEfR4xP7WdaTcVbAGaO5+RUKhko9kKU30ZOgJN5x
6w9YaZ/V9Kz6Rq4QRbaCXzJO1rmFw1OacVckvtId0exuTRaP9a1CQflTYXVkaQbW63d7utKb/XQE
hllxPynInJPE9lT8uTnhA4vZCftiRs061ujdtVNIkQcqFBYb5SuDJ6L/MAxli2jAlw2OL19wJyby
XBJPzOHiwax3wKjCFpC+7GIWvdknF0YSJfWOBbfP110lFLbMDsY+WGwvj1oo3oBvWR5eWVzkSbNy
zDOWT0WnqxAUz0aVoe6bF45ZYpIS1LaEurziwOfDQz4dsTzJTQhBgQncf10dW8AJ5vbIrJH+7WSm
Rvv65NhOpTPIy6WmfKfsXQgMQuCxHTig9y27tzKF0CWQ7p6HSCZzI0MiuIg4qlisMdIBHbKQUVNx
Ri+WvTrwEGtPqfiiQQ1XEnqP5Pu71MWJkCv7ANKQalj46vDvS5MJs9G6snaahz6GDcp7zbp3fPoA
qhBuvKo51BIDVlpAwQzIt+7IsONrBvLZlspdv70Fg20G1lLdaaUnCF0+TKuLpss1XKrlzXNzLBvM
l4wHa0MOhC/+wsGjoWF7rIkJvDP8kHGCbxHMKgRsk898Jx2HtbChIGQ+0RHmO8VkF5ryK0gl5Enh
7wg7b8p29JEM9PqfMoYntHOP18lVqHAKq0crk4Sa3NTj/B5dqbSpD1zr9y/A/kM8mA4Y6tZNat1X
1BQent/84AnXlehtSmfvvyND45UsMuspYIexfHRyiLWsdabvrG46+plNTErkc9T2yO7M18s7cA0a
ti7XxXsQ2gZ/BrwFLLEmgnGj0RdBHnvee28YqHAA5CyE5wXvLywNho8lbS3AX6BIQsCdjIvg7IdK
j7f2h+OueRlPw43YPjcqvGe+avvPqj+a5r0XI/E5AkCZcbMzEXa3RWRFlPPU+gQAGbUSBy75LpU5
y0rUlGcIC5o6QLLbYt6P57fJOcEY5wPLH7QkRoWOP9vuet6AfIYnkiLEOBJ04ds0+H3sggKaP0in
yh3bNWpNWTTO3Wd+m+ZsSKfuE70JJgZaVJVW7jHH4K3WvTooKX5UQRx6eQehsdYKX8Kc6Dm+w+kn
Ni1d+olJLWonjen5m5rICpWT9Kps2WjP2RXNMNNawBVi4EWwX8MzNlM0b1sXc4iK5FMmcMYWOmUa
mgkyc/k2fcPTY8XQLuxAleirnepSiQKdNp2xHcMgujsraybQ2zRmY/+irW2vi3OPBJy0RjZtyfrt
J3poZGEw/mTTn+U1rfKQwEUuEUXghjUX8K18/Kzh3qr7Nb9fN6wSIVjQpG5csCD0NBZEAqAllVPx
YzBrd80aqjbMt3QBoaT5QZ30zX+q7p0kKAcWVVl/RMRnewxml9qlctu2y4uasZpu7FfiAoCKgx8j
6GWWNvj86G9cARd86eKvAg8kXMsIutCAfYKJlSK7yycCpgXutlooo7UucavBCC5W5i77cb4Bvbk+
MIwAEzazFGAIVEB6Ir6SntJ+li7WPP44dfclhGokSY0Y61cwrSSWBNN+6mZ23YBlgDSfGBt/6j+8
1CddSmba5jkgnSw7A02WSDFBTBm4+iAwdM3ruZiZ3vRKfWNgY25CzvV5hWWavBx0zCq9JznZT9G2
AX7eGPECFwGP/kWm/w4vOubA4RytGTrgiQ8VAl1T31ZWc42U7G14mQoBeaEbOYOi+YeyDGPHVDfz
iAbzaknSikeVXcSg4JiGm40G9YnaS1vhni/R2pit6xvtjF3Zewg5jqfCUe/OT009x8IM8qh+ScbR
RptFwZoV2NPVPxvJpOUO2pPd29W3C0fpN3/GyFwKsIXTDFdcLn3jQneE7rdQLLqMnyajV9UIQ5Mp
QCmvBLAySSYmrNXpzUmSivNrinT8x1CocugNIWm3XQz5oE2tnLsHUqojiOrUpTWmufiFOGYQ9ixK
H1eVp7smiN9lZXPpprXAYe3iCHiK26nJ3mPTEL5XAY+mPdKiT3oQXllMHJ5rInLsueVA8TnAwKix
HYoJ8uLVzVi5FWbkChpQ5Kc9riw6Xqq+9ql4EsniUI31WZNiqg1YHqrZyObIlWGn9U9OA6VriKkZ
7YtTn2fFm7On0DFi9tjwMSnjFttSW+uC+m7LzvLB5VsqZ/CwuDlhxww6d2ALmy56faewHatxt6IH
6J+ag9RKq7rQcyuI78WIH+JXTQCc7VJGumXfLo1OOGWARccuebW7s7625AqARJPQ9jeIqhRHybJ0
xcbpJRtAwNkIm3RytuQEjQMGkis69rgHu6JDI62F4GSCPwjkx6+EDRz/GXM1iR0sjiqs8QN8WZJZ
zEqwX67TwNYgSCIzlc79zzVBrgimgoAoFNa+ctobvBDar5PbkJIMVGw9w3xgYFYzz/0ME9d1151N
28g1wryN4W7GWoubWARlJuzp9cnZlOk+9MlMdvWOQiDQB3jAunu6S4dBPxRpbGy6E9u85rg+a2gP
vWYXXLqUPiUJOnhrAFWjM4NLbw8YipEpssWo8XUR94pwvABlggWoClXuNcxSwOTPuDuO9RmpF20O
ptv0MHP9bBwNHVzETmzaXh86WnkdUS4lT8HyaZIalOa2fj4VQrbtKhue5e9pFBPSLymNZbb0yPOB
11voVwYCtznjeaTffSzZaxhGKpxX9JBc7tDpt3fHNeyaB42eyj2F46n/yQuuW7GvDRiEsHslXwsx
U5VA2I4TvO414PV4Bh5vgAeMoNl74087fnzqpiJO4LOKEpM//w5+pORWl4ZiWruNNv1776pa8RyQ
jshA1TSOM+M7h0qH7mnck2oL/NhCAP6i1ZRNdAwrSfTVR/m8aJl98WMrXPzQ2eoUqKy7+GCd3o34
pGk83sQOrWIrV8O3Dm4jXN1fCUAoVegfL+y2ON0EC6eGbWDWR2EO+9f1UVoXYgk7tcfGDXMSMLIE
BrknL08Cuzs0ZKl2zukt79kYmv5DC2JGxcHHObAWPQdUPaXmD3td/nUaseeNOsAD0i810I8qUF6O
WWHJk0WMKVrloLNVAKXVr70FZZ/9tA4Hw+Up4uPAoeZR0hzA/AeIFeX8HJzmKcp8lHPB+w32NPLg
TceQvnV7Av6dOhXDJeiTUI7SrQSMNZoYVOZTcYIMzy5sVWGjfQ4U7WVs+HLESqvHkX167RvmwAKy
AKKWNcsYWR4+OvTNVNC+Cq5dTPwnKFR9EiqhpNSvqNe7rHyVY57inP5mlkelFc4PG4Rkd5g5/sai
NoJwwRCsZ8M5TWO0xUetZYdoyLpacYHjIypJI7mJ8pIyFTvQ1jnEN0ox4WPb9Hlz7aAwcRlMP7/S
diIXZ7aeCvLjJBPoSuK6XpNL4lS///LGAYEGedTsr5BLoUC6ZEVhNF+LGx0lWFKm29/Wz1gABKok
l/EX7VQcBZJuRVvmRO/15zKvcUlmrqK6wExOh0GGKHxp3yo4gzzjVz0nxbLeR8lV1blxW4hDZ7KH
OI9r+GDp1n3EooY7xLpZVPN9IUj1wdRz0+x9ZFnxI8yc/gxyo7tKk+liNQgzswia5NuA3XtpOyeT
vH+A8c+hb46UaZzgTmiNMLHhjzGU3VRi3RW8b/GR5OnOa20cMMov4M3ZWEwsH15eQJn1vJ050arj
W54KZ1EbZllWxLr46k0WmCYUHoZB0TGTHAMUKFh5Z/n/QWreRtm4PnFBwXnBzt3Ew1it61LHllso
UP7qOO02ofJt75VtF2WooMhySxJNiL6r77EGLb8I+NAcvMLY6Sg8DtqCqEwZYohZf7h/k+yalnmZ
YptLGjDgeKxAi+/R8bhuzaptXdSwx8SDtk8+5bxge2C/wHJA6OvM8vzbB8tRc93oPAzULlLod1Cr
f3kwbjhy1u2cnFpWWUQ6hR+z0lbAmjuCWW+ZcOCB8YaCpzgg+xCEAMJ6+Pe6rYRpQ45rYZopEWAm
p1A0/1A+s0c9WJurCK+zri8+UZdrFbRd9iB4rIw4WwGl2uP8jDRaAFP83SIPDdwzGvQ7quzFnWok
eIO/2wbNUsfjmnhHvHvXFGSkV26Zp7f7SlJFAagB1nfyo3OX9miT4N2pvPRYxvL2CkfIB9UOHIQX
rn093Gm+WLY37D9Ypmo3EwRfemnsWPk25hB6B8QQjUyVABMuXn4l3dC72jQaRwWIoQIkvUoCTe1O
y6TCrS0F1zeom6yRFvC2Q9hR9RK6phqiDi9Mq3sV0JJdc25kJTW8pdd5S6YMxoyhC1ROr6cB67ju
v2lK4rZgdAM6THKJla1wP/EFVMurlZuy2kxsGjxoQ2gMyht+WS+x5M+n3RWm2EziuzrAlgWsjfbD
DP34CX7Ea8njPAeLlEqS2b5czcLhGgHGCaw7coYlJ7EJTxnF/R/xnCn/I9dx78eM+2OWDr4vegi8
d/hK1umn2m5QFcqaXIsLreUgPIDHdHrsMaL6r/j0zJyQke8LHY9O6exs3vHtlu3cEM12/GsVfN4R
GmVIyz5x3dLh8p02ey6o2HthWwhR7KapvHT7wQXjeauLzu9S/PouQ8UigqQ3zXt92KdlgFAMqSv6
XCe277ixTVvF0gWJdmHzvKJ23Hunr3YV8pgG3+g9b692Zz706rVh92SiDjD+4uxh0FedhcMI5Zkj
kD/ONlNQYZuALXfVgimuLqV12veBgAQivz4xSfZukQSIyrGwuj+NtI70sP3S7vzhY11/LfUFMgb4
WefPOXI/4KPkWpd9b3AjnHX2aW4AMnqLQE9HpSXh2yj7Vvs9adjHtXMpoYAjQ+jWYyUzILpovwI1
4zrokA5eUgKyM4QeLLIU48ezx+9vNeKou8A2NeiLNUzOjU6piBJ6ljZ67B0h6fd39ORNgUbn/Fus
1kFYcY9r1tzPtnUULOgU7/FsWl2scEH/tE3D7ms9oMmVTADafenuCBJAXYuuosKTfsDNwP1KWdc/
3BhDy3KA9tbjXpkIxtL8wURLR2Lol1Jr1+nrsyhMTW8Vs/mpv0Fnv9d5lXGw6hMKKEfL0tHlMGaV
iy/JYlPTD7mphpthdvWBcgZKtAOOELy8dbx7HFgI3VcmFqXeBx3H0Qk7+hChTQFGJrgIPi4WLURD
pbtUJUf8sEhdCBmc4duiDfwXBw0UGrcDuAbvxEeBNK93zfDr5pQHFHHjiVEZYEjP5Y/IHkgChBNf
Iv4a/dhBsR/3PJfGjI9Yk16OdP+aGWQCPEONByPFsf2svh7xOhWs4lGyCvskoeO7bYmycGzNPmmE
C/o+7GZy3MOA7STv1dwMWx/acTz4NhET65aRFM6BjDcQtNiHCbKFBLq9FV8YX1qIYndl0qKo5x+6
7cSJ1zc3uBJtO+/1gp8crDcOyvILLKSGQg/pEjnXnRs+/lD+bsYUvssofe1BeT99oNgmgZ1bf/r8
3A0k+wJQV1sk7l67kzB9p3fpEnbNPwlT5Yws9MawA6vluw9cFh+FtDi1ZsJCKB6lku18SfTiQ4V8
2JLj+GiEBoUsw5X3/CwUiUsZc0T3jbSmws9kn9W9mjtHSq1nRJTHKk7mMtCAkR1xCBAAtxhyK8Lc
AE2dPlT4nyrVlz2NeJfdEyvxftSntKajYe7vNpdCNOJtTgGbOo3Dfje8ZGbP6fZZIjKBeimgHdoS
+VDZDM3PCfpxyLsQtkDZqD8+2Y2VcxF4PrLvs3EH7x+DLDGXPpxGS8oBerya4Lt5spdpsgSiD30P
fDyHhafGyJWeaF7YVqImwTWjkwXjZVdVLHlzMy3AfRp+g1OO1ZQ88uZOfjKi9dYDPm5QRRDS8H0P
gJkZNy+PcK+QMHsbClYv8kv4TUHSrNIwITRPq0eoy7d6Ix5Tc58yr0CSqFNxs0yrTj1dvXORr+1W
XE5pq0RBh6kRlWCdjSmk5WwAYMQpwlueIrSzIK/Y/FCvPuUvJKMoqWW3AamLCXWVjb28aadxX27J
pVOe49j/AM5PFzkrlHTNSdY5uEQRq3NfZz+FrDz/ZSUHpSHJfdFodTzWulBFwyOpm9+xuu6L/F1W
Xyn98sNIJVJqrSUOvni1GMnUCzOeyyqSw27Om/50REn5pU+pG9t17PqTvUpoeHchhVW0dVzG6tDf
QZHO6lBVWLAxglf8fWwapsNQgM5ycr2lzDLret/rHu3tBVMuUeiKW89FQ0rq7H1dw+DkK4NIkwxK
c17Dt4HjPtDWYVId+bg6GtYTIDFxyk9INyVnpdgRlcwH8VZVw7anb73K7LcEcaC5GvqWOOZts7IE
yTbfJvfYkhE8oQnu6dLTOQqjlNC5zv/zNFBy4TCWcYt0fwIpa5wYB6C2/xuYBvM1VOAhQIu3fFIl
c2mIGF92Y4t6cwY5F/BAULON0JtrLdObZQIfG+n8myYQrzUecHO0QEXGaml5BMvxA/qZLJBgahdA
LfbWY+/lT0xbiDVx5FZjjXoKFCuwdh/bIKqyLnUvyYrJtwzfqhRh9Fy1eXai8dMHcTRZ7tJLRJRZ
dI651Te0RD9mtaLFeC7ZeWrYZdd8cgZET1Nsbop3pChZRc4AGpQd/SMJgbIxPOIkkkoUombwQmXf
Lr+TmR8J69ZXzr0i0iAloKDtvLhv0dVBJ8f6gKMjIQkSmj276AWzI8BlIbmRUB3tM82To+74YCSF
4CDUdQrMqDo7kxf6yYYbgjAwyIne+Dwr3P5+v72gIZQhhQIj7xQi7FdnkFywC/btEb2EDONH7BVn
7qv8T6aNb0MdU4D8stJ1pJSgSN6499eRaZt+JFJtSsG4oafm/tjohj1KglDIbczkJAhzLJgj9YDD
amxPf4+DDkP9HGKOCnbijUgf723ZwLZXldn5nJF8t54JTjKaHXgGgdUJN36PB1V4CeOtgG54jrNn
4KjdeZ6zqysxXizdP0Z4/u0gTAP0Ws3//gENnPT9UcDsDn4O5c/Cw6/h3CPPTfyd2iYcjriUmQ1d
JvrqYDtgCESPudP+SOwibejIo0OHUBJzKYxjjxCDC/C4QTcAkygnv+q1RqMIz/qs4C/D2lgzB5uw
t7eFRuvbud6gE3Oz25VRJ0wdVdPmyzPoCAPL2VL39YQuoxPBjobPKTl+cm4+ZDxSval0Qv7pirCf
iGa3DB1GLAQhp+RNCZR8/ESo4gDJYpoJn+AexPI+lnOK5eE0+iZ55cRbkca6MvJbDU6yU/1/P8SG
n+hu7emslZXxrxY4AfMXL0DN40N19kskBsfGub/FNbdagPeMsuT5ovIx8NadUKNVz09wsRYGzd/x
Z41famBMjpUTKBfBBtkSTOe0ZBucYo4W7I+0xqLEwbb4M2nIJBxCEq3r7rJso0rxWkdbjvXuZk2M
6Y/rXJVZLSscaOwyYkyfAAxbKofKQDPRb3YMoC7DTEaReNItQTQKyC39r0hFeEBIjK7ZcZe38iSI
uNmh07MkPay1NyVX3+B+JoPK0iNUMe5eLb0GvM3325ZV602aFkba9XgAKfFV/7YDmXbwbrOhz5ka
0+UGWT4Grc+v4s3txLg7fuhpzcSxgM9KxOwFknyQhLGMkg6kI8rbi4lzXDQHoMNHIA7DuPO46sWb
1emYSYEOrIWnH0PvNkJOkgU9FVXhV/Y6Kzj9wS61qridU8XritfWQvy8xvW1hj+qQWA3YmLAaldO
+A1wWK0UcSPEoo88PsOXxqwfQoCeidy+qSGaHrbICo276sw/CEi9fl7gXsvXpA9fp5A2yerjWKkY
z4Zadlwnoj9CndxsXhBiVppMYS9NPVt7ejYIpAsa+Nz/qPehw1jmoxXpVcgrzz2Ok3DRLGHES56k
v/BjYNVKc02y8dH5TjEBYt/KTt8mcymV8PNbIndy9RHgpagPqZDZLfhTZBuVccNZ3cBIAVQMPCd8
lS09ABS/Vwwh0bodUwzlTQeuTHbJ+FIAaiLmm15QJzpDqVCQnlinOLkWGLuNnc6VL32CfjkBtpCi
u1zueywm+TqpGVCniqWqbB67WSYHROE4QFwfj6EUT5Kr4HL7dgcp8Xe7tJR2b9M324q3zYNtxXsg
QoqP6gRRQu+kvZv9d/dbK4qG6tf4RMZ2XkoYXoH+1uKr0IvBiJJA05rbmnXytiVbOWIGrLoE1n6q
+u8AqymywUK8Img/BaKHh5MYx73f6GqFO5BuKMlGF9TG3JroXUZWvucfLshGT65FFYqt7QDKVEj+
XBe6mIIUy+OrJuBGh5VwOGZwPzzrwWt3hWhsDtvZ8JJU4QTtd/d0PgUp1yLNPKjDgBOPovrV0awi
uMyLLvvk08r3/pG2qrQKu8SuB+JFFoztY/i4T0uzyVeaw+38kWDF26YFuNiYzuJsEOyrS8zS1HPP
rIFHzzekc8v3UMClhcezlLzgsQaZBaSZejyaSYmiE6GaPBJ+uSo9vdH+PHxJ+EU0RZHo0WpMJLF7
MDIaMmbeYErAdS/1q6+s1AB3sEPANAn2Ojb9RqbIlBMxc/m2p034U0Bx9zs7RfeKA+Xxpag9iR/c
7tlKV7k3VMgH90OXsaO75ibJmdXCZXfO/e9X01s51XoyH7+Gf/TFdONGIm8tffzWQ5hLlYtVXvO0
Pa0tr5L9vi2i5iIDjkhHjWH2C55YipWr66zBAucOvxrTWjTJdFo+qesULDVcDi9941VR4jkfSbCy
/spQ1EBd0LxTqLP8wnfJHmu/IshBvyzVaW9e3XgdO1eNutfZLzbctJPH5CaaEBIxGFLwAtioPha8
u88+ams1U25/q3/MmdgOzG/QNAsxIiHKzAWYilAI4rPPEH4ECs/TNF5Dh3Ori/E2T0eRO3S8fGg3
TeSKBeARqvTUDTbG9CZwuwHX3AfwOZTRD0yYGkFg7GQXkN7zIe/f6qSs8GUpz+iL8/af6XVOw/Zl
LFAswUDcZSC73400cwkvGTz1NVpf2zZD/Uan2oQQIcGoM7m4cQvmeIoDPEuNev+0QeBGDsr8qUvv
WBN5grgJNVK+fXeGn/+3g1J9V73QMO/QOHzsbhwyUKIxUCIiVDsZMnby7w7j5asVvUFrjGeUKKTG
/Ya5WfVNJoUpcgopeTZAxVZ7GFXRmmMxiL7wsohD5llNO8FNOGst/H7ztyYmSOjs1aI1eaeLcmDn
cafqEskioMJ6kFvBTjj0sHlFpX4E61qzLDQCFifyFVPLJGwZKa+OeWP1PVAM0g6BgN0OCiOx9gnt
YfmyH0MovNBU2lXGjfFaI5+M+z61vFFENgYSVK0X64rahn8WJ1nKBrHAGhdccWe8OHiZpRRlWu95
yG1PrcEg9S/gx284/nLTChGYigRX8cAqNihbf0UEioFvAV7XMLC5CgwxXPOioGn2pzklPMaHhlhD
vzDQ4fEEGn5Au0VvFYKNsMcHUoqTcSnlQfnf7jh2i7De9+WXJsXRTTApZE4EesH2phkDhLKvUZ6q
JRtACWcJCiPN1QczW4Vkqh6O+W1vUWJbm97zrLcpHQZGDsk/OUzVsv3imVL27HevJbBeHL/XaEjd
DnuEOlbSdVJklDFDHskEAfTYhesRnSk/DdUrV0IJEJVoy/NFB6golnWqi2PFKa4rENInK+ObT0LQ
LKL/giLjWZl/swRkYsPio68r7rFNj6CkghWr9xGPkQLlsZ15FHat+PXB8gYhcVtjlN1tYD3iGaER
pEDRlXBLol4VVb2e1rNvAF893kE6Au2DZlineyeeejuqRCcJTsy1Iqs15tF21MPWrFNRLNQBP/KT
07r0A65l+8pCoorR6XBfAgtbBR08+BWDvXIMncLc4O9ABjVkdQh/TTKPRjA8PXtj5n/whepa/qe4
pSphCQwmCZ2c4PSgnMoso9sG7XIR3fmILo6f4C1jSE39Ac9rrerW/CZ/C1OJ+bVaR1iYPmVG875I
J0cREnkHixYCHk6ztlm12l/eygfGtTX/51G3pSOmziRP75fS5tHnsgDVG6n6DIkKBqyw6mveXAZG
lnBSZK4dxnhLotdqMlqzhpmNsbT7aVr8oMkv2V5FlPopyZlXXbkIE6aylEqeb5V1LuU7dKXneanh
5SKyyzxnyLvdi2aVzcsHIvOOVq1izisJrSxbZUs0A+HbwEz3WPEbcwa1kXxeIcw7HaJcwjffqTfo
AltQbNbV6zz0Vw+Wm78l8iuns9fBUt9RjafmZleU/jJx6VCoe0raAMJUjbQbjOccN0QTrGU/FbR4
I4/0gBTwRXTghWRVAvG5mdtTAGkvVkSef/p9cUggb9RHMyu3J1m6L7rBWihJZMc1mlSIr8S+sYZJ
d9vuW835Cgwbu+RnUzCVL2N/E97e0zd6o1SPl9Gy9TFBKdlim6FSkGkjrN1yT33hIA+J54uvEAV1
nNT25gkw/Aa3yjlfdqYvah5a15ryF5pL7qCOE+CxzAGDbUQ++D2D2OHdiTs19p5dYC6KLwkK000p
zBAfOZbHK2On8ECanu5wchyzFrnCDznSZopdfJ1dVoIzdjhAzlvrPZtZm+SrV1uNc92aBepgNq66
WaSj1QChpzwspjXv/EkMtjC+/tRc3bavqOdSu8MEKGLmkNZkBIGm7P4cSElCbYBLDBtMQWbbjijD
dseN1xotYuflXB84D1qmQqcAqe2K1/TSEhelRipTsjjUle+zFnnV/hSKBUY8HWPjjjhEX4l65Vde
ZpApqlGt4twtZDtRW1hg7wB3Towgp60IN+zOB3cRIY+zuXCDl/IQk1s8e5K57E47ijLwujbzyJCW
S7xde5QxQ74xXNkEM3cQjvOfUnxw/GJf4WQ54qSRmL7+3DOuAxeNOIgDPSDciRGhDuVF5IBOgsQ9
Nlt4w/jOrHGlaCjAEd6EhzY67FalFsUz0HesADAuyXpzfvZOm5uJKmZ6kQylNEXcqk7lmTnPM6kT
Oes45yjLdPtFQItjuXUwyLHEOWtUVTWpwtbhGsoUDNRUTCoJfXqZdsQ0sV4EfjZxdN/ucrA4U63X
3u+p4QKa1UecPd5RAsE2yQwVLzt1Mrf7MhCbeg1A3XlQiWBUlz2Ze8YVOniftLafdrTN6XS4EEU7
19Lu+EOPJdZJb6j+K+dR7i5j/NWI1SV1ey3hAMYMw4WTyeAYKUn6C5d/9t4Qn0NBxcrNMlC0uBpC
VeOpPUjZkqqV2pyVAdBdpd/d+9La6gQi7ja69QfVvYRaPlUsr/htsJn/c/wIkVxumkxPLtvfb0cf
ndOyH41zjQD6co3MsHmTUPNXbl2FgDspFDicuSVgbhaugICJVGT4CrAxHqn3HYalRYQIclkfg/13
7Y990SIHjMxWWOLRAkw3BOUaCZIwErC1JbBsdHFofV848AV7rBuC140IZAyJO7cgjkv9+FB1TKfM
im+LpDKCX6HeA/4Y1iKRTqSCbdjFP0CSVmo+Wl+6/GA4uN0ZDqCzCzrO+KtuFNCjMTJhd24XYMYz
JlUI51bD/m83FCUKQjIyUVZ3g3O33QY9Xk9XqHBvM+H5a6xbuY+yuaon+a2BpTXR+9kQL5iEDZI8
T5qEwE/ueKibSRkI8uilrQwPJKHn6v+tfB1syl6zjFQ9iOEFyNOK8ld188JLInVM4eBP2H4mm6vT
TJcCEWswqNMzSBvpwIFquFwrfEacG4J7vXwxedxC7kd5usb4FCe/FmaS9EBTfNqq5ZisvhnhWlA0
cqv+XyJ/Lsfd5oCNit95WKg/WNm94e5gSCc+ri030j7KwyNyNIzbKpQJkcd/3SLRTLIcnBFXop+/
JCMyqzAvXJuFxuI0QOSA/37+AcEN9RYMs5FEwVz9t36iJqJtXZGN9wbU9TiMNcmn9w42YA95sXN3
SBXUeG7fKeyHT7kht1BxeZTZ/ozdag9zzlQHyOaf4Kza7+yfSlRqIYogVA6nFIoY0WEbLhv2iuLy
Lj+XRa5qmF94nmmgzwnliNuwFL9soKiFe6pL5Jlccy3B9od/AbfZETfSfNRrY194IANO08za2kW7
I9tDvGR1QVolpKcfQMV2ttOGhIaq4h8g7e7t4588e/OdVE2eJ21Hzqb+vPC411yw16hm4LFc0S5b
zuDWoF+ijbk4kjxvTkv8Q+SdgjaLHFdoPxWPuG8R+qEdcoubfHtrEeO6ywqB05PGdzJujbvEbeso
8E4VZzIbebMRFiA/QA9Sp7R4ITOA4u5HbECL/IWDo3X4uc6VmSqYFxQdbCXGj+C3vxdTUtttzUte
CJLaRwX+R2T/3b9iYhFX4ozTh974e2Clz3rFxjMJF86bJdUHVE1D1PjH9Cl1WyrVqZZ9jSEQsxV3
CHAYu5B1NFI+Lgec3zrnICIiBAFa70RpJr72dzYU3xylsllY1WxlJPQYNAKH28LD1/zuILc5Cn3e
lxZEJLaXk4/U3+MUykOnPJAXO7ZtrMzcqwgIm3KRjvAoiuOINWF0cPpf9Ca6twWkg5Eu1QFkliar
gG577x0YyN9Uf+bi7Bt+ubfoVJNAQPTtrFxYw7dkG4/pUJANEdoirmXAUthCUgvFZPDLnX33UXu4
PJT91VHIT9q8YcFxAAP3IcfnRPyHbU3LfYxCF+W34ymue4OaZ67yUFUvnzkZHPXv5JcSuk5tUJp3
5oQSqEKW5678eVO0+9f6ghNr+do6Eub/zusEXMjwedah3Md021cBC4MqrX8DmbUeOwmjishn5JOl
N9EW853DwLfytm7fXq+Z5GkYnot7Pxq9zssbpy65Fh1TYwI04nnoqPG9HL3rW4iJOOwTxATMOlu6
5/9CVoAuYmgZCqjHoM9KH3r4tNcDd7Ywek+eltq49esGpdwHW5OcQ4MhjmgTO44VIgkmLCql939D
v3ken01o/2lrqdteCu4S4RP9azGd+gwWS1Dcyn1dqMnqGFk02g4nNT5TJNwDe8Jz34jFZzTrVr3d
Cll+ULHaxs+50eibg+ZzZUcwEnRQ0KrYCgT9RWBuRHgtxRiujsNVUoHeP3iGEACPW6jhBNAfDjeH
FTL0f5aijGsfCBq1/KTkai/q+O7LRAymIFiiKJB5v+a0PjdA9DoZ2iJYUXqsZnD3QElHX4Dxapb0
KsdQZtFsBPvEQXBjvBvU/4cFAOW/MhwOqNFEY/BOjSsmXsp0vc44v3iYOIMqMYyhitu+1w/G/V5c
OL7PBUzXJLqoSbVte+2AEr87Wt858+1yEk18LgpuhG5GaxzYHxdA6tIcQearlxDy25vl4Ss0OCo8
HCg6JzZbwabz59nTs3Dw6EKTH/TwCvBRupGUuf4+kXJKPcf/w20nlox1olk3N5y2j54/214oPih9
5h/GmyTDetXWVeJHcdX0g7Qq/eaz106PEmgRCbt7KyKBCrpRq5KlPfLQrjWfm1IW9iv742NaV6UI
Pb1GiBtWSw9tCNp5q+eglOkTFsioSNkK8pjfVNhuOXPDo66bNNhi4kTy3t2B7NGwhj19ccqlvB9c
eHecNjer3DmXwwUs8KSQDGb3vT/oC4OSGTnbAOW+oO7mtfl4yRkfrW3FSaCkmuHpRnus4WossZRQ
Qwm5H8tYkqvgmaqWCb4KB7f/1/mzSWGJ0GODlp4nm2UAqoYc+CwfEAUwyxHS04CBzGdh1AvkFzFx
oOOnsKxCkCWYh6JNHdHWzyvKQ+KgtAvUWClrTXpalLkZDWBtad/TtPh9sL3Yg/+OlHJwX3hjHpix
0uSm5HXAmEcNR+Izi2kTWBMFqrmpCF/ErWphiVXuzrY5yFzmKHpf6hUlPDvyX4EVKedKSxxiV/21
IklIioaT4Esobjyy/EpCe90VHu+IKkf24j5TkDiW7e6wIPK5Hneyl4EGj8SXpMqniw/1VlouKCkk
VYYyxJNXF8kiZASLwZ0Sesol9JKqUenhbB90R6tMbTcNhSfFer2YsussQVyNpSsDIamGuWBbt/is
WRV4cwvUFexvlaPSguYDB+HCe19ECG2xUh5dfwfghZCcIubcTRqXznAGW5w1P2ywQ//tZLIZ7Hs6
z/Bxhj8Rk7f9r4wpLzGavYZSgwDRJIASfkPdMHV1VhSltKE2kpVKgTvCn8hhk/Y0lKAQZ2phh8lW
f735RuzZqo+nlXV3gNmrA/V7FqDruulQwNHu4kVxhX5U98Gji8P9nFmNRj9noYmVAhZ6KFyjTftm
e3N/hulIqb60vQZaXYErf3PcXyWwGkZf88T1IZPqs9X8s1SFs5t4ODl0mLDKoKDj5Ouop9bFuYYK
4zjSznzv0Yn0bXa1CIPld3egLzvVl3rF+WQSiKFuCmEd6AFxEogFzWXhihVbfuLoerNS/sYNiVAy
0tMXJLWWjATu8OXVlR7v4UNV1WQ7BXX5h5xVkaioFKtgK5rQH0nyemgP2IAbQdyeWH2I7WJxJsEA
6Ya2oV4r1P3K5ddT+KkbVeWGdHeT27S0SUj8lyz7IBCTjUWLSTb/VraVPfxend9IOss9m+AdNiqe
4RD4jwC/zuerSKRFJ7f8Hxz/mFFuUdTLBKvt1PpR3CthMRl5TNnD1rjEZW/ktoY1cSjZHKDsSQl0
s7I7gPfNAjXck5RcrIitiWJ2YQykb5rTqOLv7c7iR7dd1xijtvNfJQtXFCmH/MqiWcXK8QwDTw7f
MOvMtTBC/wR5jIu4aqT2J1oJ8CFk5NW1uMc6HvpSP/c4O1e8RskeRYl4ZfXP+89ZOIntWF1m8VaL
LuUnZw329Zjz/b7QXwaiJWfooS46ocOTTrhgoSQoYoFGMrMgv2GIxhvhDv2csxmKI2jTYOBmv7aU
YrkNWOtpzFKFWtF62Yb8c9Ln/0WIX6UI04ILJkkleiObLqkYs7Raek85Df8ox89wc/2B2DbSANKK
h8rIVSe4gVUYmnzCtV4ouIM6zlZ8y1caPVDbMphuDCXelfSDtKahcNOoML0l64+gdLm4syOkYTo3
cVXPeNqmMFpcknanP5Fm1KsHA5QY1Zbj1Lf2qdgpYez2W71LwSVzOP8RWvUe35SlQAOcuN2Xsgiy
3vrZty6IAha78HbMNmovUnMJz1UKRKoHr50YZFMI4gh0VFLoDZ6rMxbHefk3I5ZzgV0QMyAwbqj+
SOy/UxkSqr0HTwK6sByHd/TRMwjZmnbbK8GeJmLfTELf3sW+Bspt5DjJ8C4R4I7n+a+JJkO42U4x
4kXiv1/KhQf5uAx81sAYI+CwC4Ne2gPxokjfGnuMjb9AqI4eCtQp4VA8RvzdccqSgVal7NJpMUr3
tx3Hd+LCf7VmE7VtACtC7AkKBrl7Z9dSKR+y6zN3+HvgEXTPxoV4rLgwhi2VMsbl49ukEm4Eml1W
+cTHswEkd40gg0rt4jhXeEm4MEHGD+zCffS74dWSCfHkhh58p545lliYIAvnYJ1h/ynqYbni6/VA
S+1TQmtltbnUQzDZ7a4KvJHMkVMqr5kir1uMHjm68yGUPK7scVkKJ/ptK393qcZUMpX4LH79hnfU
7e3EkK3JdKPQgz/BJ2iJLeayDJYgsiyMk2aPigTXv/cM+hqzSjF8emrIOxeNRHLuse1bK1/QSL5a
aAKvxQY29pNGsxajuzLEYdmV1D0Q2BkmkwkuyzXbYEj5BJ4ZVXCB65a7Bhcn9AFMPOCEackGLjqo
zeie7isnGEuScW1f9RwGln+0iWpRqHFHSTcq6JwKjF4y1MOqIFTQQ8a84levZzVDG3hhyN1riZQS
xeoZjp2t22WBA6tZ9ok1p7nlcZrzZIr+YKOXBWURtObZ7qL3c9nN5NiWgvALhtrmzSSiSk3YcQlA
LFePMz4ItRqW5JcEBl4zDGBLorTb9gopdYgN3/xkWaNyhkNuQ17U0PqP9AVSou4KQX9LoNET35PW
xDzDaDQXlv8l0aJyFdBrXjbhupxAB+1BFQLt8lCP8s+FWXKHnaDDerl+nhcU6DJlS9eTl/yhH/wz
CgwoYJEgdyJaob9Y92RRWMU6EcWR5AbyuoMGldalf/a8L8GOHrT1MosM+tqpzcKVxF/xYUE9d7e9
CXYV+DqJJatJ6DUXXjTNLM1naSV5J5GY9XaZNG8eFOAQmd7XHGhZDgTD/LHNvj7JVtSL+ToejcWy
S/IIeUcn6F4NZAVW4ir3lZzRYLGha04braXgqxdD8BrNsQxgLIu1+RLZp5oD975doYJTKa2loSF4
nD55NN48kVAKtLwdykOnpdBIiRz0OxVvbTBehINJgnPLRn+9TU2IgXqXsGFpvHL6Ajyq2tfEcSr4
vhIvnKITVi2JhQZHHHQyZpC1PiGgbWrBqmUgOhq+jOJC6KyDuI0600pEmmDHEjjAXjA3o0H+JQXl
J7lH60P/uvEYOcjk1vUewXzs021KI9xTQIhfIrTH37KWDR13c3AxlzgbXxXH6SNa9+uImVwKnQ0y
fC/7NTKdtgNApksWr4aYq2ZEFahlAXk1ABuWgM44io1bxyEi2/yXLwEQJnFonENF1yAGSULEZOYx
LuamwptWEP7dv9H9BqOTt672OoJeYyfViQOcX9YoL2dvz0rdzmcKZl8HBJ/oPXVjU5XaGbJXetms
AvQk5yuWj7XC7D1P1eUMn9ug/VAkNuVf3ZfqkzZPfMivYftrA7XClOeAcfo3i5AuzrcN1V0HY7TA
EByjgNGO4yKCuKWVZumkvi0c1NPx+IuLYxp1uycI5U44F5f4G0PHkrMgo1f1ddtiCdNedsSJ4hVg
YPRevq0htCCENXcKwAFfK87KV2et3TCa6LXUDhSmmog4qSfgtc+dQvC1F1y4GgvPZELOtl3EUpZU
YsSkD1pu5SVNy4PQfv35MnOyBkL6j85dADMtOC/FIU3AIMR1Bz3RSblaooevo1DgBvjyd4B/k9gI
jGJRPv2GJgxHEYfy/uNPPa1hXg9DlIcpmRTtlwgvxS43Aj8oJid8wmUL8q5zyzS0dncgKe9HghgK
9oV0UOraQJM4YO4RP8PecXDFwWnXwkq9nPCmZ+Z26L4iaqyGxAVp+ob95f0kCojzYw7JmDbwxvlC
mzB9Yl5+6A8akUZFJdBUAyGO+bHQmxl76MmktnfmZqGxtWXhej7wu5qMbc2ZgiC6905MX8hRXjQu
u9lXoun+gApaLbmKr/Re6AMBZxJ9o28P3H6gTKZvYLuIJFO9jfDoyBw327I/hC7Le+PjMHwj1osA
sCDFjiP3LvpysCSkj9Yj8xZbWRC0CYMJuyBtGlJMMVZY7Lydz9yoDBx99MdZI43EoVEuJYSF6afB
t1qKG42EgMbVKZv9FDSlSJQGy70L4ylOt0Wj4MaAmkp72ElvyzNfNNASZwsTh/rtrVt+fzBcjIts
iVcBEhcJEqMMDwHSvS1t/jmujIhMQMSLoVtiLbBXNI8bFtDbxOCVxmHNZgCUP+HyYE6aFqSIBgyo
EeZp3nVPgImfbYdzKqYRn7VoOwcmoN9SBsBMeDDL2lUdBtwe0CU4AUEw1qqI5+vANvRLFUn9KUFU
cYfB0LmnimvHo0hfJwWmMKNpg5RNfoPUzSMUp+BXZSm/6/7LQ/YQXue1dM2sJpz6m0hk9e44FDuZ
xUn8XRnOS1KwaMr5dPcofOmfX1HFeEA246KBOWyavVkZRlFNrOi/1/uzzF6yyEoy8IC+1Y8qXUI6
7jEkaqRl7hT0VA7i84pxnkHmnYuHhCBMt5q0ezjbAkVB8iIn25lZyQ+sdHxPT7YA1PQJT1+tf4b+
UW6iLc6RFWW3dP4n1SUzuAFnrHjhO76zqLy0mQHglIPTflrnfDqk0/SeRGYzqL/b4nlZcg5onW8q
FKGb5EsU+zuZ11JYffBmaixdHucMizWqYyPCTtKB0GjrGEFzuR3BJjEy2MvTEK1jqW8bKdfKg3oe
aTXnnAzh7Q9lynKrH81OJu8a2RDT6NdfA/swV66vjZl2xayNuNg2ZhK/FQRfUza9f4cGoQ+Ge/Lz
NfNSvQe8j7RzYkSfAT2eKDBMSgljszSgEOGN3xbFU4e54SwblN8zCgzRotQveyE1IQtgBhHgccBx
7rqqMWvEvwlvOs4MJ9rcJjJz3MxIkiVlE/fJuZ0/EyKDTEtLWi6OVm+RAgIXZgW7A2NdZgeYIRl3
NTtovaQ+J5iU0hiJ+B9qbiwIQ/QLyJOlu1psrkttsE+htxBL7H7RlYpj/MxPFcXl9HM3YmWYhy3o
QtfAKC84kFmaZmpFBMNrREoEPVXaXIn1j2ssBK95YucHV5N/A5SxRwhDdUgolotYEkdtgfOnDNdp
bobjzXLJAdqEZoKHKjm/oqLUwjrK9dM8FN+o5vx2XrGLTAnfbqzBLmeIytkUnkeVMkK8qEAN3ImQ
9MqdmKaM9Q37cJajLuGukMF3OG2T3VQF1deJe+w7b+aoCylWxu+tQey5C+yNRN2X5lUH7Jm05POi
kMGxUh+oMeYuN3ImWIsdKDJsQ9f56OcOi//n0r4rOuhkrWHBB6a7yWV1fHenETVzY99WnPN3U3kO
n0ihhI32boSxOYvR9+gm8cq8wEq5nf8nMK0g0ib0Tn/K0RbjSKJunkZeyPPbhtE0SCzvcyzuClHe
gxCdd2AKMUIxnwYrI4jSOR/2RI/3WB9WOScuEqK5kIj2iasPoP4l8qSNVnCbKNPjBL8kQjgO+sgB
cjO3osAJLtFuBECuVZk3vyJP8ZK3DyyUJdkmJBcw0wAWgfduOZB1B9KioUFCuwflo7HO5Sa44TC8
c+gFYAU+JSM4qUWH8zS49pAa9TLA/ST/DoG3VR1ks9hvRylIPkZ0rr8Hny5OC8+nbVr+ILzbdbc2
RyBt0pK0FbnvlCJs2fespgitggbdZ1413nbT0uYMv62MgbwvE/AujU1ruhFqBatmY58UeP1hqxeU
ggj4lFRgSygEMhdi0VNoYhZ2cpeQ/sKN4xrPFyCx1XDJslXLs22X/s0yYJ/tX3vXgYlqfn1YjhtH
Rj/0GE6iGFArVRhdPiQmWoaOPpchlbJA7TRn3/+CvxakWph1owJtPbs48SJvx7fM1V1pJQiBxDD0
IdnpWuj6a4Y4IXdtNEPlrRulXY9YU7edGCgSB6CzrjpQ8jCMvklI6HATiOOaB9Avhxxmj74YyfGj
p0xT2rOTB/STeqb7djcMjMRbnFR/Zv+UFeuTRZl3EH94THHXyiHBce8SoiG0FksAKwQLtYKl8w37
dPRoTo0bzr2myBw+VdQnwVJ7A0Kd27jBgz8KFcYHGQKJGVXTaJCNrFgQk3cKp9mM+FguLIB5ngI+
tac/eYJDVSV62RM9qwqWyXdd91i6+9nWu7nrxULE37hiYYpIFNbQ0koPg6d5ogtyUAhBreZvmiEX
rEDNYBnhSFe3E3JYuBmFTomH+6wRxEyg4zFbWHKzjoE6qGPNmwqoBazY5pRIyKWZ2VKX6C60hjOm
WT78aUy2Truq7Ju2F9P58OEFf8avfJuV0ejSSFFETTh8yIBYFvwF5iRhbOKAKvbWOUCfxofk9k2J
1d2dGdaSDcQ/Pk7ybatYLA+k0ghqD9oNhpq5YaK/nN7RWT8MvZL6N2qr81R53eFQEg5vfC2Q5+yf
hqmx/cwaIeh8IUJwE7VdjmdzNYxjRuaNLfsxTSUkxSuVjm3CK+D8tBfT1xeprlTkvtEAsHVTXD+I
pqNb30xaXSgsyQvwMOY0KDjSRf865LlJm7kMHUMGdgxaydqpQdpkaqa7jHyLZ+D4iHePoJopZrUo
ZesHyt+e9ZvkbqERyI6NbQB1m+8tMuGI9tagHy9AJswqKL3gdE1r1YeGsC2wxXUgFk/9518hdqpZ
ru4X3jP5Q6XocPYZku1xlP2kfmV6Yb6nS0GRXG4Pr+O6lfOT+A5hEb/NpQ+0YvgTgv9NT734y5EQ
U3FH93EH43NKMehaglEDYIdPThDpFoLofR0VhP5JHWUeFBCMGf5Cg3Ykx3iqVyc2dBynAyQ17Aqh
ixPy/pMz+0kxlBZDbada6KM8hYGQmo3JKmmM7f1w83mfTD6XoO4KDSDXCkDKjJN559mKRMSushm6
7T3Ic7T2wzZ3/ux/PvyE7MnvuTCSBSDl5/qJd0eciImiBcShVzlfsxI3oExTCARlTRM5P3fiMcJh
6JPNp7j4kpUlax3wQXDMzjC77vjWtAiRuFa0b0qsj/62eEh2NBwWh5thL2O1xNwu/jdXHV/1Jiha
TWTmd8WO6HTVo4YcLzw9ip5e5uLGwaGNR009rW1gtibnAteMIanERl3zvjllIXV1GFWbvAVwAPOG
oYsVRQJU9lbboC0XkLgVkc7mddbipT9tA7iq7DHLx9e2lSJuCma4MWpdlrToLjWInODQ3IH0So5l
A5AGaVdGNHrfhgGijsqbE7AsgRrb9ZxzagJTtpv7/W3Ksf4nto9jqC7EYGrpD1lbGwxq+ieCqokn
wsBBuqYAwOwb0iUxG3dZ33dhIDG2NM1LX/7h7ubWm33BEFP+lnNHAA2Ee3TqHneU78qu9m2NhduG
2uFKX24oUiznLsJd4n7dpasQBoAmJm+QEGb1sl3TqWQu1u9A8UoN8ORT7b8T+G8ALiAI1WCMpfPI
GSev8vLZwuyz35loku24L1vgbUWRwaa5WPQNeCKWkbVk3ftiYpcdTcMgtFjczgXUTRC4dJJtCtXt
TucV6KWDkEH5tIqzQCcEADn6/5x4HuCV1Zuf53JtqfVgzrxVt4ajUNyWQ50BXkMAmYqF5xRV9mKY
PirRmaOYD33eMUCAx+hrUU0xfTfs8DMOhLf5P3bY4qN9TJ0qXYiYaentwFxK+1vShzDAkqTaVDID
hX4SS5+tQOmOioP6R1qS3TliHmB8F1ymbo1lLwsGfaWnvDpTjyABNvF1h/EwQ1YEnX/rd5lOKTRs
11Q/dnIig2KGN01VUUNOYUBg/CTn1nhCIQMOd8sR6YGr2ZYBWK2WksrrN3aRX5g19GpR+SKag5uk
KhfNnaECNh7Wzdvmhfa2CtUUMn092IFGB7WKqerRK+T+2l3F8/1qNBKUSzoVWuN2zJRlPWIZcs4I
oLSiW6+rdS2mYMo7P0A8FSvBWeFPUR/b049svccXeCqdBOH+fhcQTLvA+pRNZjV00Q2vgewFUMz+
OqNKaUhfidUF4ciz3vwuAwSg6aq18ElLJAGqaquFby2z8RHy/j6H0l7snGCh/ZOhwwcZBwK5nG8s
kFivcQRkv7x1N52pvWjfhfRTLNOqZ4d8QseXDkPm/3d+LmVAG3CPfOtsZBHqktjqdb4hVn2LquI/
yfYLKRSrX7SZU1Dyt4Ie+8Ap11JCX0wCAMD7XS67DWLTqObbx6zsbS0GwKT7QJ9C0NmTcpr0kLS1
2FcprANjM6+CsOf13nIiOMXa7jIX2GNpeT0/p0Yaa4gHsNSspbgLc/c0hu9M/0ijDT77a6q5CkH0
yZQXYGPkdR3snFSz6wnGWvPdK3a37taEU3lpe4/AgFfPcorizuUwp5oJkiS1wTp0otpYLdnnYWfj
Vk4DjUWuDkPZ2Gqa14M7jXYvxIKyaKWNF4H6JaV5Q0lfC3BsAu06c0zZRyq95fUQcfZwZ5GSUvMx
uV5/020JBl5t3R0d52Y2H/MW+k+S5IlE+gn0vOpN83BChbs/iWmOmFSoBi5KVKvDkOmMQXNMEFNc
ZkHdR0qVLMhvrFZ8ZqQJtbzYpm2jOayXLNXtLGpHaB090N8lYDQhmnWKwlWmpLueMUi/ja4F6t4b
vuZo1AiK0QmYed6Eexl6snKC5efnkXWibrAk7ntMPBHl7Cw87aVPVuplbhx+wdcsOhK4Y5Op5KAB
r5olm5HgClBmMTkmJUQ8s9O6vc2pI8MfgGiLNXP+22FDImsO0VSyuy4FefHhEhalnrQFpzH/oc0Q
jnKc9MyaDVKXhcZA0y298vt0lGVPheFqqmNtr/RKGdfGYRoNLDUJWQ4I/dESWlM65T9lk+Rciz8Z
rbRZfgWxcjUnmMyFRO8VHzQIXaFCwB6t29laEukBWLh1/hcv9zwK3vDMfzpbP0lyG8hXr30a0PFL
AuCj7inS8W/O11GDf7QmKL8vAgWXONRa4DH5gzLmVtF2GxqD3Nevb2YDBqJ+VuAT8r04zvu9mWB6
p2k+oBWsAnqyApyTMWPIYds+12wCjTlA9cFojsy+N19Wq3NL4+bNDKZejnMLGG1Qqp4VwIegdJPI
FWm0xXnATNtR1QATBwpKpyS3D3FIR8x/Dxhz8IQTyOsv6kjqR2q0MpaCt2i/RoW7BJhj7WrgrRPV
62fz52ygxiahaOv+8axZbhJ9TG0426sFMlLzD8Kwp3hm5rD83HwAdlj0JoppLdUzHVU56gQMKZFV
9DnvzXjx+yDej5ufB47p2CHjznXxLeFqKEDNYWudfVleC2r2qcVq4jthkJT/0S+EJ8U/X2dFs9GS
LRLKRAZhmdeU1n6F9SbAJwgyuAfE2McG5xsgmnguXe98c7gi20/Bre5vzgl9s5rW/VmccltVsv0B
AbwcD5eXr9tBJnfnLTvj688O9YAXrFBU1ZinZO2kGIZ/Bf4FYyoDXIBULhVGDrwbcY0U1BZgV26t
V1gEni9SCMxPReR8Q/TZXNhlFenwuE66rrbInspShYA6UBw3j8/SpvaSeo7ZPhm6P8GIJL8mZu1p
VkM+Tuaq1yGvDX+X9SINbQ9rKlj04q4lESyNi8OOpiMzmE0nJllFpd+4j/HBF2g3gnJulHRY1l+M
GeOcyxDhpcogI606CLgsIsChkjlpNCATY/87v10+AmFdf1qTe85FWzMVX/C75COxvmmGmR6B6AY+
vzimC7FPySpgJ2WaozMF9wnwboSNz2cns71BsvQktovzYZZTWBZXkimUzSHkVqFV6zFnm3o2sAep
7yyuR3KmTuMNcdRxTDuWOxMGb5qITXo0/foUDiLAUq/cD/FlB+D+B/CO4YLc/WBdEYK3sjL7fQDP
ASUbz355M4I4crhHu5+7X9qzQBKXsDI8apt/qtK1ua9ItvcX4IGpuCs6XgRvm7/3zhduDGj3FNyB
+F1HYOCeuUE71oO7bEmgB4zskuBxxVfiVtenHaUEscBWFNEIL/p9e8KQ1xK1tSryzB1H1o3i/16H
T3Q/PROQw0az0Vkdq+m83DQ5Hlz5yDKwJRSPPVXxNq30qY/PyGFgLNZ68Puu7cG2s9qVFJ/VKbYH
wWnA00nc2B9M+DTcKWWVsog3Ty6bCIOEaEq/EGAkY8b0Ud0CqkNji59AzSRYPZfLn+wVMZrnIlzd
JFhCGJ98lo1u5iJJpA+Wl3UurwoPLjX7NKkGiMQ6utPHp/ZhNrL4UnhXKEYQE/Xag87NcbxR/WmJ
VW5uwf+OsEx5jpnGhu3fR7K+Makvxswo/d+0r50mWJ9mCt94dTHfVIY4CgJwaSwM+l3Bkx4+yhwO
6Ws87OvOGOYZnkoc7+5u751w25g640h5b8FRYZb7Y1RWKxQywtx7vvdy7T0zK39XzMTvPKUNaYPl
70T8CXsYAR73HlhE5ma3xM3dvvbH9M3Vm2TFcd+a5DZoK7qOQZSYRl4B1NQctDpibsGswfxoE/yH
DZJFtp06xtUPFhrhhjgo0D2E8aUQPjheTA8zddTicAqyqR8THgsz3jZRunZKpc8Hmt7E3aedoOxC
Ul8ZPQb6hn3uz8itHi1BuMTbjmSVlcwreTtFxgBdWk7vaDGVTlf4wvWIywIcz87oADQwsuh6yHV0
o+Wa1s3J0e8SGUP/PNlYAhKcv/Yc4gZSxOg2WJy50OkZNnjiz25Tg8gtekHSqwoJxPF3wGP5sEpW
A6j5pXILsbCzWFqdDg4lPN7b4+6zUtvQ5Li8cXne4KxSovPcAR6mckBP+0799kiZOnnOYwLCckMT
eHppYZns8q+KgqiqF+KZkVEKKaR7+adpkxAmNxiAou8evkseP6LhJDRdIMSg5TmAUZ9A+go9r9h+
1LStKBRYIYYgYHGtNtbH4TJ7MbhRDXsAHPLmTGG6iD8aFobahAAsD2C8ZKbMoZqelo4nMe5DO2XO
NifsUef/n+CgzhvaEOktv/h+B7NcDZLpaqiRBK0megOWlLUjG3FeQX5bfrRvtu9XNkBFOca+vCd9
XMIsEk+sJBV+moOHWVsu4AFCSlatcoeLwrXh1vkdl3OixXsSAsT9xu9vmV+fAyIKa4crZCkpx28p
novVuRdpuOEO5g2Rrx0VflBbVsLJvw0UHdLIVmpVJjqKRZuLwOPY7Dv+aHsCDZCbm1vMJWaBJGey
AOz5Pnv1YAEzNuSkx8zhutHYno5XXw08KgijyhNs2Bws7Q0bCa5LZm3LCNRpJ4ajyB2sEThl0amS
2v9KQ61RYps4Uykv7PQf2MAiEJbtuTO5GqZWlzpozuTvWIGwet9lUq5UfyoP4w5PtFxI5yvhIw0z
hTzzaUOTdvaJUnfyVZZnElquIL4LdDAQ/qZn61kMevuELuddXtTiTe5nLhBaFpt6Rv5OjcIPXxN+
/IfKdN73LWr1IlsjXLcbo8UKaLi6VSMuFJdhJMsitn+vgeLy+ZDms07lP+2ywKCKNTWljdCShvoc
XymWRJNiUTFDBHB+xg2RuFEkQ7hzOghg89gIo4ZmnQhDCBeBamggLuQFgEvhO3HBotSRzmbg48yk
FdOAoe9T0rx4pOd5/hUjivnqG9QtBndGrtkf81RFsL01NH0trp1f3OBcuTLbKVNWELb9nSAJLVy+
AFVRfIaWDq0K5fWmnJMHngiXFhTS6vELhTeum5PW+CPOF/3ZlfvWBKL6v3VG72PeBr9tG1BA+Gxt
SAbwGX8fzhveeqyJahcnpS837vY/JjtAdZVFU1AoMYjvDdPk13whQRu5uI7nNfQwxCMm1xGhfNjj
yQ+9LDgn6DijjoArPjgnTHnZxlCe5rdzP3rmO7H44lDOCxuISSWjViUvYbeUwOCf3sOXEO+gwLH2
hsEZ99MpaPT2D4vY8BiEko2U5gCheufMxiu0Zir6Hv3Ycut9MEDHekzpBqcBZuI6G0NQn3hzzy6o
oIJQVjtq/RtCzz1u/ejnvc245kgwreEyLY1qno7n6iji8tRX9P19zsexDnkGQfCV8eitLX2uMElv
Epw6ikrFhzI8XNCkO3yS/yKldnlQIg6carb6MmBgVqcc6sd/x3ZXi3Lx8LB5gd3LhewaZpEX2kYQ
HKWPuLa8U9El5E8ADsVgdXFA8Je9UMD+Bq0PezG4yHLbRbOAVoOQNNCWPa+yuLd9pbp9JwkkWlLQ
VYqGmhnBAnHz6VV6KH1Cn5VvuYI6rAEwUWvpllFjZVS4Px/XrTP3RcyOKZ336Xa17LDREwxf678O
sfLMuGJ4mCUtE0/m9VcIiGmW2nOFI9MMNeTIYWyqNKoBvxPhg80p4NPXRKmbnUc5qlAjjmgCRFt5
+Ne8d9G9kezBB8w7nAqegjMdikbWcwTImTrXFPRD7du/OfLnuNN7sdOXwuF3EJhzYap3SmvSF9xf
8KXunA7p2R4iVS/5/7Zlz8hdmvtp5oeAgaNB9TssGUbbSuneWiFn0syI4bnK/SgscFFHfer2FuGq
fx8pZKrXKQwYbUsiinUWE0GMl9ZzC53HGGDx8lKxCjQ1ECcaEJi2fS0MGD4Tu0rzrYstMTx0eqDM
wwee2k/KSgCyMly9Kz+fobzw7N9HovDUtBntkpcgqCv+/zEHhv1KdCORlyvCldVQmEFJUEdzOgRX
Z9TaWppiUAWVwGSMFIK7ft76VFR+rih6m6BNv6mqQdOFch9CDmQxHHDmEtpdhGrfNwNCIlKtBLty
nKi8eveF5tAZMiRB0crThDUKR0dRlmS959BuRQag7sINnGxBFeKzbOlnIb6QuDTiY7RT6vF2YhKj
V0Y4x8Xq0wkilOIkyCsCkm2N8uXzfuhrL4TqbtLejPOosHdeNvyqQZanCY2HmZ/NWxFjAHib2SSa
oNfet06JljnJGtany565KKof//iy5SMrrcl3helDWIDxy7dxmz1xnPmohBBc2IVaRgJldyxZEm9f
5NFF7eKkF2lIwkl9wLVQX59DiG8XuHerUocrjGYBT+AtLV2l57n5uPZ1BTuMWPprlSs7t4CUx3JO
QsFY3+LnYtbgwu9MOk+VK/KK28poZix7Q/ujrhbEu+IFqG12T6O6DFeYjFaZ/pW7EZ5sSXr8zejl
kOLfom1eVgrsY6GmrdgrM9l9EPXWQCcKQ54OOdX1ESIuvB9k6eXn77XxdEJPCOVGEFY5NcNTPzmu
obJH67DFQwYC9Jol+RVuDjLEYPzuN2k0dynYQwwR75yGK0MKbvYQtSKGWUI80i9jOIlQPAM+liKT
j+vOxVa5EyXItNP8ar2Q1fnkjvH7lTToXKcVd9LvN0/hy2/1jXDpkj9ZB9xyztpdUPXcSCnbd7r/
R/CRC7GRb08O2iMFrIFFCZlFnAqBtPmnla8ciMAwQ9O2pTjHwXJqhNKpLb51oFh9s9eCYyFKCg6l
NM29uP7gC8yaVM2qx0q+sZTXfwkH9oRq6Cd5epRsBs0ldzRD6jP+AHwom5wCu4CUe/UaBxCCyO1+
wY/Qvf1EsMgL++Mx0Sv5gc9KYtQIgs3zqM8+42Q6ZKs0uSrFzcrcgikSber1DGamGtfVT/s/U2QD
gxtLUHFFKBtO5bEiSHP56ff2AIuSoUgLTmUMe/g27cYBjZpdFDMPdzSST6C3nVVZgRGOxZHXB7pY
9HzI5yWrlUT12gm2B6Oe7mIvtpzewheCEwT4rrkBGt1Mm+CIR8oNA7hZxa0ZcOXZUjAggMX6JdZB
8leYFBPIbnqN0dH1phSFhH8mKzMnzzBUiu3w9mO6WhxoNG02F6wK4BIrYAQPb89vKoj+j2aAvmWB
y85sE65eYhiG3kp1sbUi/wnW/hrwrcV92H6c3XO7AgFQrjQWfZshPIe4c5S1CsVCYGZEmzscUkcp
Nuo0Eh5nkzMqy62nV4RjucgvtJsODiqmQ577GJ3vIc/wR/+U/XoTnaEEVY8/VJX+cveGtp7J7ykl
DwR63z/ia2SuJCW+78QkazFxpIxA5P4HN3oexsMjoddrWVizYnsS6kG/JF259yxwIKV3tvufb98H
tnfxBIpm82vgI3Hh4d536nqeiE2vgCnnIep8vEg1daRS5OLLzG0fdWvkmZzFimdRHunRuAApSUZU
qgHIyRU+B9kYx3suqfNiXe3xdYBBBVV2O443Zvzob2zoaRNwjfgG53w0KQCHFtYr61OYyVqJtWBE
ICJ/7M/ZX4g233tDg+ZunAY/KjDLiCn1dj/S63ed2642o1oHGKFSHs8/NxVLVjKjtzOHdCZ1d3U+
Ry89PfCbFxUbb9ByJO4A8GEwfPRRGXcuXRZGmI4sPchPFUQppgiVNA/Dcmpfdqk3B+TE9w2jiRb0
BSNlkEH11X+6X6IYVnX3BiZasVecJ5JiT6RAfJXN2xsEWPK5CEZcmnrpNEO7ncL3TuWsjtyeqQjO
NcIrImvxGZhDRlYNQvQIg6QyucnQkogjmEdX2L3bedV6bA0aWaFblWo7ge7TQwrGdS69zAV5eNIr
FWwi9wlDQzq370bR5Aw1hWpdAIBVjREpTMvqdRtQSR0fl7tbwbIotlXY6g+2kTBzR1zuzjvQQuvK
RLO+7anxodajrz8/VK7UgKpvojPCjeJl9uJmTBwVbIR4yp1m2sOZoBsFmd4Nqi9wAPxtH096ed/5
LfQEDqBYUCZ11Gau5SxP+N79UQAtg9i/ggch/gr+u0tLUBE24izTb4XQ1e6lTBf6tKHbM4YD1H+l
RFhu+eDL1GYsw5eJQCoj48J+hYHj+Ao4ehKlMaCeYh8tQpNPGuifXRODL4mpmhl73kgbxSpB/jVR
lEIkNDDr2cMjF0cSPBV17p3WqsU6NipjfOs5AkR839ePAtptuOCzEKdSZZhS+HSWqDR/4u/P1ouh
IFkXxXlw8q6yQcgeIbXXYr5Km1QTnb44jjqfWzJI/tN+bitlXXmVj4xFSCozesA4VSk6wCozBnZl
oTgqTuoYzMjHX1kjKyXW52eL9rjnLfiRsjMN/1W0DNsDLeP9lm4EVlHq/rTLoiCXZFUDtdCbAF9X
GXaJkySpicI4ZmZVIU0WDf/zvjZa8yO+iUZ402R2y/QRF78fOH0ajz/s7IO/gL3vwOwfrMmjkbKm
kGXPRKNuDDKOgtPFXr2J3OYgZyqlInvlfGp7lzvIbRnzOxRhlt5uypXmy7Uqj1h5fmCCdbHhJEWj
nwaosSY1CYHhCpwqlvcPN2bcEnLwwcSL32GxZ5fLFI7HouHEoTW+2wUsHR5uTS509svpnRUUdn3s
uaEyZX3r0PJ2h6D+2/0vgeI7vFjEPZj91UNdAkX5PExNdo+cIcfjBTtnLDDK6AJaFK6GqywR9KVq
LbdIEfc4eE+oEcl0o1ANhUi7IMQeTR1+rWp0CYkU70RWn8Yri8ZW5RUl3yvrwNk7h7k6kBZWDRys
Gp+uOCiSz1Zl1eYoQLuV1/nGRDiyTnXV6QXlXq3uq7SJHo7P2kbmLz4X5ms97fginmQlB6EDeZeI
9SB0sMu7V/XnJGYqpTA8LgEemE7YBmdNvAdh+wp60UaxtHbAV3ekotg2TAFr0NKWWTwCEDsAIy0X
v3+Zqk00Jt8UdOdgvBkVu8Gnu/XEs1qulELYvWXxwJ3gMOeMLyVdNQz/ANSq5AwE2dW3WTv908XR
MQkdbwra6q7O2mrJ5Pz/JcECbL0zGzvO5hD7rMnA7e27INswXh2FRhBHuJbkZ2kS7zM1dlsNljPF
C+WdIsb7LJW/+lQ7JwXJaX2C0/VhsfP22erFRvazZ11/GBtD41hU3O8XuE9ruu10vJxrjExJymUD
CsGi6cG7Oi+24xPH6sLGCsHl2htUWlFwTzTwIbEluCbH8NrKvxdf2s2P8FNTnAfsGVxXrs7IpIBE
+pBsxQzFKhNWTxYBGMOQgqJ6EdKiIJqg3LV5K8FU+MlxmS2Qkr0+8qjaPiDGwI6Cqr6Muwwc6xvC
M4VZYdNuGwP7NUhWz7Yr33iTX4f7ywB8i7n+zR7dJxsOFhGZnIHGnNsSiRNpkVFSryM/WnZMgMUV
euMeLUBHFsYYxT31hU0nmUtJvy85ni6i2NN7hWE4/EtojxQ5+aOHVGLErMG08H8XWgYDCQ6M7YJr
vizBMB1xml668eCly1nxEyHuzbh38JetWI9DCew0zPsvPEbIUyhCBExFZ9+AXK5xIgMSekl8VG0k
uhhuPWd1e87vibAylo6XGEyfnUbH9fzgsUw2TB4ASZ99g9TE3n7/YItQG1uNaO8+vLOQrH2oSsW3
hf0p3r2c7AOMfxql1luyusPZhgsFAKY1J5nZQiDjkkY1xOAn5v+VbsQ8e5AiFFc3cSUi4lgjtQ0S
MYmCepYB92N9TSCvZWi7t/MU3SR1CCYHPiozNY+By8gIZImKhKDfnSsUj/IaKyipScn9sHqP93sb
6afS1nvWe/7toL8+juZa3owh2CJQ6Klg9vEJ/vdEDltCLKdTzlpyj/q8WCCXZxMAIDLWZcNRdZV7
M6mabuBCsgVLhutFCj0KwOrvQRSEmcQ9jcRzAlfIdcsB+XHrJ8sXyaBwANmemGNdNRbdJ4tIlxeM
dydLngBtHK/jfWb8GILAZg6T8lQYQ9PfWch9f3dZ/F/1noUYT/3HhxQ4aUHKR6f1zrbYQ8uebHOk
JwBW3PjqdKAcp9zN/ZL09Al0dWyZK5UhvGVH4qqu/+xHwVTO0caR/PFVAh2g101skrxkhRGdeISl
HbJKEXro63J8XgIRaWTC3upMe8J2Ry8yXqmC7O9WBtuflQnRVxD8fk07PqY8fsjNBOISvqTDkFin
DxjQrudLf9s+voptEaw0tu0l1JEN+mhyYXvQGgwOO0kzEZp/KvgSy5eHoiN0ue4glbaJU6DRm953
hs5htZEBTAuleqGkB4P/pUVB4KRYIiI2Z3/ks28PhYDX24ME42jdYNCNtlzNHPWQQ41hKtNUqVQI
LVy/zRUG4oStk1FrIb5Qu+4UuqZReU9Y9oFTS1Js0QiMJFHe6x5ccjS7kTTm8D80C1ZKId/4uY/a
46+NDJBxGEByhR5Yoo0OlILSOxMU6H9M9PmvqRFiir9f1+bdyRv+4Qiyfla4eR51leUnoQ/jV0G8
rExqUHI/5iKy37kUibFf8H5UArZtFG2ppaDlbRUZhKE482aDbVva80fL3rtSwWu7TamVDMutQT0V
JHnqXLAyr0RvS5IjjhAAgkDJoUoJEHcv8HJaIaF/rEFQ3Vj0xCTsH6AhSPtPaRUc3P+0ShI1jv5b
EDWooWzrKOsmAcDfOqdRjalvWFCN4CiscfWJfpyKCKQsg1fAVTj6vk8QmxP3vKZIxP9xMg26LZbe
9MPIFq4O9NPS7Hm5JfYQy4OxDr8I5w+DLGynyuan3icbDfY7BZHpS+CutYOyuKRuQLR0kCOqOSXT
6LFCV+zbVSF5DRncVz7VEqROIBquBpR0bEIHu4afbzrQsQco2ORJSfwTlaEKAgbAURAdMdy4U+5Z
xkS+qEfKKIyeZKTlNMZQUHPPd7/5T+/OiEwmcmSnWY14CQdxaDb7NLU73Bl6CIfd5dmseU8PUfzS
m/iHwiMPvgHFdN263qoIE5skMtICt5h2NranlhlF+b3k6xX9QKNUykSF//SPTtwILR2W6HcAaTxt
uNbMEk3S0tCydRN3wZ0H6KJKsaiUZwOgMKlga/gCNjbUm9MRYvGX8yP65w44cGy8HojGpWWvVPvw
La3pKWFkdaJrtCMv6autzJRakpyxpSVJW2Ka8RZ3Z45HxIuu/zm7Du5eWIVSfOyX5g51kje34wzk
wuK6dTJLYhHP8joQQ2naXrZZgzVN9tMoqUqSWRmTd88A1KPM26rHlUGpUKRNuZDtGmSny+MpSRMN
iSHIWKt2JfjG1SCEhtjpKwiz+RDxiY6tdrAuBu+05feZ9pey6rVi08ZYSVI9kNgC6hAcnzrNI4fx
NY4LGIVihuFZHwhB/x+tqg7OKsKB81BT5wWBIvqjzi9vgp90u04v0QUkGmpEZIU8g5grBXdr709H
hy2D2Jy7hu3D4wNayFQflmB0noO14or9fPFi+RztA42RN0X5FUO/lIM2xlM3pVMtUkhMMYF0utxt
bM92kXRDZWECK2Bl1+bp5RHs5w7dvJ2UIZclHsKOA/mN1KMYtvrgiAdWQPd7xj5gcOz9mdC9ASHm
7IbseFoP4/9wqO/c82ooIW7R0iULfaRLGWf/aGqpUracJoBS+wWTdC8evB17hAiPo067OaoHVx8W
2zr5tjsW5oKzd3HoGCplFal+npwNjnEQgt3kHBmdsWNLWmvG1e2G/9brSVF4ispBOPDRqVUU9MBc
bCK69S22fDmXsOe9h3F74RMYzS20Zy2z9ONtj0Gk2q71qcBcgYWwRx9aSgP8Cc90efj5+r+D+xZz
Ur4iRaztCMMjgZgCA90T63WeWsS/atjuvueUJvd/wJeqfRyydCEqRvZRyu1k+jCxH8ZAB9rjyNBx
5rXIDrrGbLxLLJ4HmmD+BJZJfjJ76Nndzth55Rwvq9mJa3a59zCvPZm59soSicv81tEpuA+x3gmm
pcGAhjhYrEnssBCtDxIKv3TJkqfjr96peKLck3Z3IZdfJFGBchAN/YsWWSfB+iAekz6lMQm5+prB
jAPk3MxyL0IhRW0DASf6L8K3gFONnkJ4WXh1atv5cRIZFUYBkeiOYEhWIBEKvkr4vE6QhS81TBr3
1c2TZDJhuXTnN2a1P/ZytPDpzgKpXiVfgAXk4pOEq6EwVkbdiY39cccJbo8z7XE/GAM/catAl2Kb
kpcbWpt8tALhLUoU+u4PIUd0AD0o+/Q8zL6MPsCoPpjaquGWSTPWOUmbQrclwdL3RdcLe5wBU9NT
GLpteYMr+d2W8JW+GjKQOWftToOJ6u0+c5bFR0rSSLEo4AVGLG8/G4corTSkA50FaLqO8yaH5Zrv
reUhrjTuZ2eYJBzUhVhaw8MlwDweBjw1oFnX9dguMrq+eomUAT1FISaJhIPccuFB+6MpZkunnZln
mZEZZqZzrN6vbAjjxfY8+dJMaNZDJqjBjHw5RuAtN6VkpadaC9lksN9FIO1U4/me4GyXlJVtwiZD
cDX66s9bVKmadnyVEce6bMJMeFxruYmtgRtzSNNW8WqBsuwzqTVNVxxuYOcNTC+POFB24PnaiMku
ruq39rp/TVQDUc2pbVQbcvuMexWBWYXw5L20Cks/G3JBUSJKGqI87zqaSRlxozmPJc2WR75TqIyf
GMMu37qojbUxkGYNJaXiNvEmr8RRYXw8fcB2tCde0aDn/5lx/8sDTKv6aD3w7BXpelgtpgqVGBOo
nDk+sclaR4n387owoN+Dh4/lI9oMiGkuGT0MvCKXNL4V3mRosCBBwzqzStZx0ymrd0kVm+djqFC1
WFqG+tnaqjHSu3b2Cy4v8pjdisH/T69LuYOzZliMOpI14sTU/ZzAMgIBj7l+dm8F4dGlWL8PrpsH
8zP0bXloM3IUAvTrbLMjbdygKQ/meKHec7dRMM3eKbKLBPhcTa2KU29CUqt6iurZRBSsALWRsd0x
ItvG1xNpTrdHC3opej/25cIwT+qeW6RwkIcaIWXzv+ws19cWbhXdMx0aLvguO1ivkmE2ZQF0GNBt
FBdySDHxwiWfqJOw+7m6CDSmpqW6YFUk07DPt5Wy6+tCH4u19KMk/FVpIXnb3nKHiDXzn8zLnO0P
aNjGmXzdUlMChD50wsXo4+lY6wGTINghXjhhO4jyOp4Xo+pSVnlvAYevDuiQgF57f9D8MOClevpD
9IQ+0e8MBWwm9kuHFqv4bix7TPX8foDiiRomkuKdTL30Yn2mIDnT8ihQJ4eMiHurSWd+R0SBd0AH
N5D1Iy1iGenD1djHgEXhDzfEW55XRMWlk2Kox6gHQzXBLdibEH0+9Mq84a9kRhuxBW6qYUIAmNys
FXZM5mSEZT4YRE7/C/9vWuP1RLNR+6BnHr558a/dIbp2S2uJiVw3UbN4aqlIphDvqGTsT4aI5aPE
gSXcL69nnXA49xywl5Z+X1EqisoX+eGlsjj8pddpRSQCsHFHPhEjo4+2i5ys2WVGuj3tv1vK5snK
P29HCP0Pfzhz9aYut9YuZZZXtL3wYxa847vKo+/3MOEl+OUs7xSgc4HHs+GFiIl+J8GLUs302frR
ObQUmt5nWC1ce06pLwH8yQOdTb27sq87euflhuuXx5EO2DKFgotb/YlsEjx/g6wXdgYKl2i3fh9W
UAvrAVN/F6l1MyRk9DJPwBGTw+FMWopUajt77X2lMH3OOk/HzEamCDm4VBSm+UXceP4J335Lq1jE
xMRM2A7VQwPHdOjzRqHnBvT5zdYoiftQJedvUvG8EqrtZIdAs7LJVCZ8zBfNktrV12M+KVnQP70k
tZWRHeO3GSk9Ek5aRoQN2FhbN7cruO1GKNxvcHc2XYpe7V8OmpK59xZa3nTfjCokjpoJJRWYfqOu
OBiKxWASZ4TPMzBZoynLyRRG07OtJtt2wQBlCcvQ2RPAGIeXt0c0pjQOAcegSdZMwSILnUDfYuGj
/XvVI54z9qpurEpINrp2TAg5TVljUIzBbGgw+HmITUaa9SdBaSPja/qOPRaj/ej5mUIjVnRMMW/n
jHuMBBDrmgBuhsbV9gZ7WdqDL6je8lbhyOfFP6IbdGSvCiZp+mMIerpL7Ph1MnChANB3JE7QV249
gO+VDoIM2Gn2jce568AzghS3JiuV19RZpFbE6IcfjywY7C8WNj4hvmCIPWUkxnytkh902nm37UUY
kw+yINNIvY215YJl0YLdVKfzpA44H9Xn54cH1fuxRK4rdxr7Ylp/pGSOYgjHP4NyaeF2aiz7VddL
TfkZSrKU3gGT67c5IhGZ1iuKjQpKY+cfpqLb1oGIfHHb6564ethFW7UKEVddMP1wpxTk5beMNvWS
FTNLhJjC9M0hsWtapsHcV3u1wBCT7XXakiHwhLbuUi0lHkBMM2vSMXg+gDNYglgF9wfnR9Sgq+0D
iC06Cguw/32uAuPyVgvOl5bPG3ums+gzp82Dk1eUX90vbHgc0qj2xt3aQ4wzBgmsAozAuQfUuoy2
SLrUEKlE+i92uaIX4oFgKwkuppP7WOxI4ubN0IhAWjNCXRfmtGCLB3xnq8w0yafofq2/Pq8vdti8
O91C1l7ACb7DWtjW+Y40/fEj2cSx3J/iDNlscnPJOv7A5mMp4WeM0sWsryFMDdtc85c87c3wMieH
YyZ45SwCgwY8euUAAlLq77sDGg9UPbnRS224Jp2Py5YCB15FLYcaVo4hTdpnEyTyrznLCZTjepEA
mxhOkxX4Ni5SY6O+4ymCdTP7Fexiwiy2SUKvtEy7/+nSaSuAW2xd6Vb3X4vxDQyfZYCqgGfUUq2j
QTQSVkgejCHHEg5a728n4W5ISbqPUsTlXwfQzDoXcMH4Q7cU1ZjILwU4vrinohd3TRLkvXDOA1it
9TFEItULMjMnyCJwkCjUIl7CdWm5URa6/TauP16p6hKuag1D8KU20XXKb8fvbyPjI50s8mPWVARU
S6/q5R6sxeRRjSdOrBR7GknJfn6bjrZn1nJLzCFUiEZ2no6MlEoSBPaF/YkwWVO7S7lKxpoCkAso
ZjEQk+Eb8WiaiwuEzXOGGiG0NJ2BjZCRscg/vVU7c+Ml1rpx/N6Gey5KC+63qJEgjy72I9ebmdlo
PekRZtbJnesRVtgQY2PFVOqzlsWu9XZsZKPVvGecLoLV0HZIv31iP1Q5ibQq7lZzBENgr50JnJ7p
w7Ra9E8ISvl1LINomymUDDoNhs+PjfFvsTis3K1aXKv4H5KxANUKC49QpWN2UFDjOP07bfKSwxe0
qCWhuxczI64P9/nZyUaKswa2Pm5jXqtdVDH2zclFIdiVHOjpOjYOvyF/sUjAosn+J82J20rHbzib
Vl3Vc0+NaJ16Agv9yDl/ki2Vj0c5nTBREsO1UWtH+QZjzgvJGtfG2JcGpRC36SAGamrSGELukWtB
rr5AnWHnCZb7MThaDNi4AYv8VUiaSDe67JjjLEanjq/497H61Ld52DX813T3rBi53492tL+UOL8s
b0wG+CVPvpH5/YOpSog1zptW+OXCaVCWByPOunScmrmHhLjjmAqoIiuiBVhci/s5RHhKVI1cevOX
F6KcZNn/7ipB4nUWxLKsdwZYuTbrnDTZmfE9S+tb3LakAHBegDlozQoDn5fI+MCL37GixamA3CAY
pcjnnSsVVR/FjqEhjZtYbz6K6KRv6ezXecHMV7sKpHJ1dtXs+mPPdMun+D+hicZtw68HWRCMPSlJ
tl1a+JxrdqFfBBOvTANVjPf9Pd3/q18JKOcvvVe1yzuAhO5ZiCfWN8jOTTKJ+2nIIGgfinCZ257l
7HEDLX3f7x5kOxKUDrZ5wwxdiKx+NuOMWeo8GFQ4QElzjcHzTeqaymxyEs/C1MluMXZfthpHWBpj
3mGVd1f72AtlpLbDDKrxhd7B51FqcogkvZm7UnTMCQRvolQGlEaG3W+nbBHNB2rPNAKErre1KgUm
tADDtWHp6WKb6W7nxWow4SIsfqK5dmiOjvjJ0V9COv8lGCXHbeFqj7UN3PrbpQztO2AfheLEXUCn
tMjUEhUU4kYVpR9ujKk98752/i1r2V+9pyPGJrBbCXLS0u9SKJUGHUQz8a/bDcq1c8Gogz8QCfZ9
R0TC1uDqVOGqpnt+QHSA4aOvRTkkCO0bqsD3pTBJ6ye+jeAltcpYh6I+U/Iaev7xC6ooa1dcGFp+
y3/v7WMLvf9t2t050NHzrMXMMdTbf/h+bSbNnHPf9TFlifPqFrb2WlNoqrSe0p96bVPKwexArY5w
5Iz16o1TimfZTxbBKF8sjR1YsTKf5jEhH7ZeAuY7LdDtQDjeZE8TFNRvc+920tpYBvApdJ8QcntV
h2aQ5301UXfcHdzM4i3uLKKGryU4xMSnEYAHWBd6iwiwUv4prnB+XC1QKXU2xUJ/6f7RL5vcRrC+
LnNaDcChrINuSOQLl67tBKRo847eCAgnSSUqZQGXGjFOe+df+x3+FwYmCSBPuk60tTZCGep4rQmB
fv1Cu2Fzi7nZNIHnvL2FNmjCWAxHTG+qRGTI3LJrI4rpGb1sd0VCkVyp+ZIIwKKVMjyouYcwZDVu
JSX7qv6qpzcd5jgA1OCW832BFlx938vfy23UezZqYYoYwwQFlKUuQtw2MfD0HwlwYKw7/nxTd4rN
7v+pbSFUzAxqOzBDW1xXRbbXEAZETZ5jzOX8qCq/g7ZvQAAoWBO2k5+p6Seqj5KMkxc+jX4997wr
a2b8FNeAooVyvVlpN2q0lvu4USQKWy672h8013mDfYiUmybnIcP7tSBohD+iMCboeSIIi5KYnqEH
8stojRDMLJy+8Gvm0Gr3KGzI2w1Tk58s3ONeDYJkU8ieS6cssBdsxFFUDlfaNVhg+dNWXKmNhMlN
o5I6GrugQAktTMxVfpXLBydYlgiD8nw2JrwTGsHaZnlV8nLwKQFvZqLvb9/+vmxZEmHPc6fw0nPL
YcnFmNZ0DnbqFQstEqPUabflSzMbzG0r7J1ThXf6CX03yrfqxBTa2Edn6HlEORiy6OgwZoW0SLnp
8/X4B2HbK7dF8nMQo59+s4L2ph4SxRNAjBkZPjfuaf1DeIMOaEaoeo9/gcYZGT5z+YwL1Ug3nxP1
PzSnE8OiE7/C7f5melxqTjm9xWibny4i1bENZc0AYiJ0yX+CjOPQFefBSgtl9rIHA7SuFjVrqoFY
kvfWHt3whSqbsOE15e1VuOYaXwxogwPmpocbMX8D2X1XrAMpIYyrlu+l7b6yCVQRvlTvxC0L+0+s
BYfwoCtSBtzH9fWho8b2OhGp/403H0jIQ3paQGuJWtSz6cai4h7kflsx7leQn+tfIS5mQsAAbd40
MEohyjn+ZIyAkVVmSws2GinjtL8k9enAA82XJ4Eim9X4JUIIjbRgaSZb9u6+s4lYwu9HsBJxutNH
amDlM0Jg4/w6DFUR6DstPdJ2FrLa1pOt04nqjFPiU9iZORc9sQvwqTtWmu4FiZ+Jx210WJrQsLJp
xQbXSQ0jR5RjD5OynNYFZ4EmElD52AQ4O4Adlffv+eNuzgXgK+888k3HoMm/EDaxpSacyRlJZscI
HdRyzAeEqX6Kw6qlUNbH8mXKXF9+vGYvX/BuR4My1+a6Nx2A7FidLq0Ww/q8VTK1dx3U6BqnWx6G
XqM3S+/BE7r7u4bGtXfv2KHOd13uLiMtnPkp3CCvdD6clPZZc35O09sMiDOhdxDO2QiDlhSygR8I
8bGng2G7lLnc2Gump73GQYpZ49NR4Ks8rWHvpAhsWnQgrXDe7GEh4TYfkEWp9SbZrdHgM4EMySHg
VJDX4YwuFU3TrbbGU46XZ7yNUHFy8xZcCL9Utq5qgdnDs1RSbiK3Cs/Av0zNV2eRES7uccum7cKR
8L9G+vvHZiLtzSsnDYezErDNfrq9VZV0BwE+szobRrDkmxXwthI9HLEW3KvrfVdWZdgkA9KMqsb0
B6kU+sFxh3VKYSngHW6/XRppZ3/8ZMlvk7AsbqdrtSfKpEc0qtzmIUEBgdnuEucmE6RRoKROE3Fw
0MwExDF4zK/Dp9TvhomfNTXR1CYBKHcdJaNnmeo9ZT1E5U8O5cF0NzbRJqsQ557gp75ox8K56Qlu
A3rjAPBjy7G7gJ6HEVEdVOOGylh+CffHNuzF1FcV5QOJo/yBrrNsGHRyIIglCfu0UWJzG5XheW6G
wqAIXcFK6sjG/t75JB23taCj6cj0qTryYLmd+Jrj71tpX6wGOw7AG1J3+e49ituZkaNFQXfLmoeV
KukQm9s6FfYvamI4opvlbdyUJcNPP+qsYnR6xeLPZwO0aIf4GBmH+nsUSUYELFBuUuXqkxmHtV8f
Q6IRIqiradjdiRopFOttLbCxxACedy/DKtRCGydAJSsM9/xyFinWaZhQuIVC0WiBl4I6UfkzxqDo
rvID5uS5R8nD9iA4R/eUcriCy/xVpo1zDFlRm6xkGuaO0DN9sOgIfIwT5nS5WC5pD5oU3Jt4bzb1
I0V/p6Y/nFEBQuw0oCC2albUwcSuarBdjcwn3qLVdFSf+sS+K33kdJR7Ia8itw49gHZ4eiaUVtec
W6OVyzhhpbbG9QwtJQ0Qa0yWj/qj6qIbk0k1s6m3qUUFubq60qGfYAwLOZMeX0M7X6wmwP61BjPG
XDU7dXAx216HSEQ7iG7sFClGjrMkrbz8cWAmfgqQsI5wDfnz2q+6sCj4o6Kpwek9AcBgGgQtwacE
7gVh35Yy1TxxjrBmkXu7hfjQDeEF4u0EgfNs03To4nOtY9LcrvuTGHRcx5uGlCp2VU6DrQk8K4Vj
rzHvuc2g+KoubGymaJPv7RixbJEjmbwdUI4JYexYi82zMhsv3Bx1+IdZgzINVp8C1HgVuBOMWr8s
tqjbNhU47XBAXpj85qNqm7mO4Fv9osMuBRY2bybEaKK217gzcFgJFWLpmv0x1Ic7Vq+dyUVjdmEK
px3c0t1VvME9NTAyntw8eOtuznt8rqguiiFdB6ZGXg0RssBGi854GM/VcuKHeR1bS1qvc5de/SRu
/Vw1ddxqZ1x1QIJXP8JbHCQtVDCRAoHzm5nUDGZRJB0PahJPzeK3RkWDF97SBGPrPWOgkBJbC/CU
Cx4xiysNAZLbCtlSWQQV67K0f6L7IsN3wNB3FABZjcN396dyEO6/njwy30lTblDw7Hu0abrX2Sd2
aBtM6aPu907BcNtOwZo3dxudqCTQmtZCMlDRJK2B+oT2bliyCRLaPuInLGY6E8donz3g82+9ROQK
VySgt1IbAW9umHqQSHwhXVQAf1kv8d6QgcdvYBqD60SKZfBx08yybHnA9ouYWLtkTUjkL+u5admf
r7cFHrkUoDi3ZEoX+65ddp64wLVn1LLKl2CDGu3cjhVAj8KziddVVbbwGsGCKdUNUrGUvMba9OFS
qp16MLRPYE2MZSHShX23fo4roPEh/i8siEg6Rv7rOn4O6Ah4oRaMRGz8KlYODgQYCELfdnDuK9mF
5t9c/7/mdPYcPU06aXRetDlPbTbUXn/U1zJ5NfHYP7q3qfZvwb0BKyXiPhS8o5fgWGfVRSyaQRKl
EXfxSt9zA4LiWn8mN7Mm0H3hCFAfQr+3jcjgu1xXCl+SgLTiaID4fwXFkxz51FfkQyRF5FsXbEON
/f9CZzCNPgQdlOZUspDriFVpCROwBT0RF+AdEe+4qr5Wd8AYwraesAj/yzm/StPNyuE2bzF0rePU
9j+fta04UA4DDEO3bYsSWtgGIZgFJz1eLY/gLuGmF79w8Q8CPZd62FcpsCT4rD8Pv8gUrttYx0eC
64ZWdmw4e7U0fnxg0Kk3H9BdrQaJv1+k0vSBJ1WTQCAKAeuAA49aTF9atk0QkMTZfUsQgQoCRW4P
WYjqBSTbo74S243+sdE1ndhDsasuSelE5g/w8pYmc07m3eueZDNoxCVmrWrPp2/GKGyo/wTOuJF0
bDywBMCcWf8QuOTNgwdScicOUGr5vHvv2xmqDPETV869FNZmuTrzMA5O9I/NBbr8Wo8tdjvTymwP
idQb7mCINHxIiPCsLzlCN7AZZ4Ezy2MSVjJu72duaOM0wbsdxjw76pM33cRpf1LcsS+nQBw2tFCf
zxqb7A1lBGw+dkFlO8KRbX8cf0VCmhtH+rxdUlqwB4QtN46JnlIkG22ezOrRsqe9jB1QWHVunu4G
02m3rwdshTEXfRpevenyZ+D1s9pGpO/X9clBJX3KyAQZiiJeAvBBfBP4RLZyW5yXY8i9dqSMvI03
6lSuG0nUGSFqFjyYL9L56JrH8uRapqnOIiS2vg0EI/Y64Dn9DEEsIJC4Qr30iaUJvxO8beabMML6
QD2SiNUlGk++Q/XoVuXnrjSbv+ct9ZrmVYWmLkm/Uz3RwNSwNtqCwCg6T9nTajV9y8Gs1/IqfYfJ
qJ7SQLWvuGktgoVMkzgFDJIYXd2pWNLQxC501GQjg90OQZcYB2QpjpvKN2dYfNoXl21VwLBsrkcO
U+Jx5J2jWqFqt7o5V1+SWnQDTuHfjEnQP35OtLdqOcMFHVr5JLQ09UxLIFS8QOKhTfhat7dYNPHI
KTnyBCYHy1xBbE6wRHVYXTt4FgYajM0XRConbWt9ddCD9w1O/x0DIYtqf775Lcd3SOsKE4Wi7Lno
rRQYcEiO50oCtFZBR7HGNO8eeQSDP6kcfnHq9l9rqLyvqgg7k6GEzNPQt5eE3o8Vti6UbQpsKRfA
9p+x5adOVuPDqr1aGyT27XWioUCUqNoiGvm7JiZX1JmyxKziKGZW6NlAAucQy0nYxu0nQ7biH8Vl
4cVT0CmlLzP+FWjhDSxXFvk0uWBjZc5v5AzlFvUkorr1q5WQfqeQAJuKgubCLFyDYYS+d5nH/LWP
jN2kPWUzHb45sriSkfaWbRgjklllpKFmR3Jtnp8caJfJHsi433dzSQBSzJZDG5YAuTqSqWp1SG2C
X427OdEsvXsEuyFQjc8NMVCBtCgruNojMEYezeORSxIxD5YEFsnXOnmNEPNP247KlTK3QCOmUT53
piR0q64yv+jfzCzSWvhCgmXbc7UUzOvb05QFf5CFV9sVbbwAQLIhnNjzJAdIMXL2YtN0OSbwKXcW
NkN36RnGW9zhymAnl1BC5r1YLrNwksd6DJ6V2BkG8Unsvotlk3QUW13m3ZzqPqCOWoY+uzy/AryR
SdmOLjvCsEHTZlFWbRtHr5jw7skpHmYBbvRrJJUZgIsUqPaPLDL3fJIWRira12rCbENLEcazVjPz
pZujiKg+pwdohTBxECACaRMM7wXW9Ri/G9xyppYwqBX+JAI8pxxLEg9x1sTlqIohvabPgf8vghcP
GMnipLBMVmL9s/D0ZbPd6HBjQxOoHycy9UoP3buC50j8XtiB1uuqQIN94V6EatQLHlsL+cGnUYaF
U7vnbY9ardc3pGoFuECyLu6/il9o4IklABp02zGufg0n1xcyh1RzxcJ7MM9SmhVnNtuczf8meyyb
eWt6jBrStnGh7Ipu/05c8qmFtg0oic5F7tsotSI+nL+GZyg0V16kKAphX9CFVbu0u5yZ5npTytZ2
qSqGc4PkVptEwMbq2AIJOUdLDpykDQBmqc4wjRVXTLgsXOvb11YAzFkTLiFNiSQmRZkMS5sW2oPk
xo4PIHfkfaJNFCcszSlmsNBdHI20hZBQu+YAGtiu8PVEtYvNh/OJ1fj2gYhf627Rpg0UaE3WmYKT
QlKS/2jc4Px1gh36LwvInnI09KwBGgC6vjvtvuCXFPbAzsPsN+/C53RonzKp7+MmPj/YQpG1sCA0
dPisRejNzW69/OhAL4nfVJwRgtU2zS0UX29FrnEwLQryBcQ6qhOqFrVbomh1sfpqxtskFmTCfKQp
iurqviOWcF17o/22LamF+CPmRTablwdDEaT41PVyH7sheGet0p+ZPxVmo7qmsk7xzR2KOE/8dG66
DO725x79VJ4K/BhGncotoE6rib3PrJJtEE8S59zFPjR8gxicTxMIpsJpqFWHGBTYM3PLxhXgDil4
AS0flMRTf6n+8lwLPeyd5pOFv943gkiirpa2alW19+yInHIxHaqqNYYEhLfvhtakwsnqcpnC50eC
ZYNJLa7J3Zv9Z1mt2xsckd74KxHxrOj2Cicc9XIpFJ5MS+d6MT3gl7K5SJDfNacCTWDTksMn+A5F
JgDVHZhaUD5ri1z817rVkdTawXAoH7Vbnpc/9IcwqBi1QiJIvuRuiXkmK4Rj5P7d53rSGAyfbhMS
vPG80J6jufOtVuTBNCrB1aWspNNtkm6J/Mdh0dzt9r61ZffvI1wOzwi6+K6tp/KpaM1ia51OR9DE
wDyUCA/sYQptZgP0lBr0HYd74gmesOma30+CCENm9NlroDYSb8Ur14dKU+sSQ7D9/dDvPilQ583V
W7aSycODxpdAUpG0NYAk0BQlz31lgpDORVmiRiveaXnLznBWfogpm9x1x6NChSq4SQIR6m8hy3p0
ruvMo9P8nF1Up9LmCE6BDS1st3DxHt7i6Lu7B3VeW1PdqbN8nqnN2SsOQ+ieiC9fTEytvt+Ys2VN
Wts0LfFwrEWBZHgLO94uqBCYMNxX6r5okNuK5DM+pdrUBbAh8AAjGc/N7dxqQZ6DckHL45c/Ti/M
G8YcafiCzn7A+q/D8CmrxlFL6a+oonuBSIXjBBiMebD4VIe0qj74TA/ocqvFQGSTHwnBpK+d9D0M
gLXlkXB0zMgY+i9TcCYN1P5VAFjOgVa9rZWfXH1fnOv7RCnjFFAtHHBEvV4MFgoxBiXTMg41SRJ9
dnml59cw6toO836W6sjC4uC9xR4CTirUWOKwvYG6xixn/KmFzVyyfyTIEH2FoMYhVgetp/QZ7P6N
LydhPA82HH0ljuynHe9k28OJpQdlSvdoSt2crYOG6Ovk47ZCnnXqA3PUr7qmR5k1+gYU8gNehPY+
+YDjxiRHX9j41oGcYkskJpGjgFjwf7/9gHSeeEyskZKecX6965UO2bToJzn2SZOlVP8OHf+wdkCC
FclgVHROB/P6SqdDOKn/b1baAVEe26zozkI5hqFr3vdFL0iMajtedb0qzkuP0MQC2tuyWtcGNVvC
DRAcNVGBoU45XMFKzdnwxD3WgIpVHbLKzfHgV18Wu/E2saExPETsmqw63MZ1qbloIEqkiG9U9DOk
MiUO3RCUlhLZ0xYjXEMeQ2N9C2KSmtt8mGdy7P5zH89zwHamkIlAAgKgWNH/f8UcHa+m7RBazit7
+LnTE3MTLZOTyxAWVmTJPVd0UAvznXVHXZCzRYyLDDURu12pnrAjqZdxcXzN88KUDsjGuYRBtEmm
IGVjVqEVoGHjN/DqoVoqWyMywuLT27aIae0qc0d+75q+ZgMnS9kL8TNG5nQOVpgSewARgVvdixjp
Z2amvGl6zfyUiuh5ggOSIetUshmC0f5C/4sy/7nEv+k61dU6IJSbvU4zcgipBLnycApkpPy005q/
uR1SFzI/g3y3RKdMTisb5rTjrtLfqYUqksvViGcZoAlFhybVJqv4OkT/HMEBEAumR6ujcHK9G2mL
Y3nZx+Xkub8Yd2HS8X982w9cp+3rF1d6KsCsN4zQxRjLPKFHWZNmOZxKXJSx+Diyxsp8+D5wBJno
Uja3vVdDnvKVOR9sI9PB35D9nQQx4K5DmM8v4zwtbjRdzOwkRHqMPDDyuualBAPWYUc3RT18qdeU
umKK5i+bv9612D4GJIuwF9H0rme51FxsgoR35I6vL0HciLYOaJSuCAp+TpqrOzXuJKU/Lw/9l052
HZcnwfC9q7BYMT9znivjUs3bqTtJ/tD56nmQzVLSETKCwsYMvbX0fgI2KUV0j/eebVudMO0GbRNC
2G2oPfr9EfAzUDbqrOqXQIIlRa6LGziVwEYya+rHpvpESUS1/QJpSEDyKXs9/wzm7xuGjDtKcx0o
AkBBywbTuBD9Kw/FBm6ekr7ZZd+GzQJ2Glk3dW9q6gCeel95KFD8Rx364VqkKWfLybMNy1NSbnrv
LhDT4bnbw30XUIDerWR9vkFIZpP1kXX+euDYA212V4LYk+pwT7NMy/H0rcxCoLogLBkWU6fwRjEx
kW0E3Q0lPQ5eP/6Bk/M//lVqMREQKczY22Ez0GbxcrjUhhrANNDYX2s01clv/kIIR3YbtTFHf98G
Q9B8C7V0QM3h6rvUnuMMJwX0Quhj4lp0odEeJ6INXsOE6G7xQ0VDqkDvXFrQj5IaNCpJsggF2eBz
4GrvtSh+J/+nQ/UTlb45IFDFTBXndA8WxNfUDtzMtPc9xg3HrY0CwoqwAJmpjAqm2jEkzBKRQM9l
m44mo+Rvis5uB83vYQwF9rJ8lfkaKDQFFODYb+I2ICJS9IRFU9+HDWEa+c8YR9fUucWye8GfZ7sY
pRgiYBZ3wYX+WP3l2lR3AyIP4TwZoDPB5XvgI/GQ+uTjWb1XNb6TV75MXtROFV1cOF36QHFflIq2
+GFVlnx6kN+3QXOYkJIqlD4rhSJO/aW9yrngwGa3YqlW8DsI/kfgkHvFeGqaA1eigusaBDomyq58
/vnZm2G78G+oevGMpWFgy9SP3tG0uVsIVDgl4y78tA4zQ9iabzPU9zZY/8TCNRpTUi8iFXDwDoXW
RMyRepWHPL2hBvVWjMA8e30AU80XEBZcZYLao38+ttcDq/sn3VJvbpfMRW0mKSINPZlJt3CbKV0Z
tz74JSDjIlcIUhEYBJ0zBTcVFv05KdVa/3L/ICCy7nIfn6asIGrBXnXjnXLBlE5mEygoi+R+yI4a
nfHT4Iy60lHsp/jNPv0l9cGDdNoBCfEPeg3HPX2qifO2km+ACiTqKVchwda8kZ6NUw53BElmP8d0
CzYM6g68Q64h9OKP8Nc/X7qGwZ2bA5H5s21vXL246viJ7HyRleKYuiAIhb0qQ6ZhIEIzRCPx2rd5
561kD4eG/hXmDFMFshSzevFz/0NORWPGf92od8xPGJFCjaFb0Ey4qHWRr/p2VhMB11GWkOSesCqX
fHDnYtW/2DS6vI9ik0YN7v1T3xgwcgLrPVFHN4xySpVwWS4R1CsIZ8p1yMlhDFDn5B0/BWtjwi1Z
gmW3IImGPl1NKRmxGzcI/Nh7nqyQSHyabK9jQwi48UP5CBZ+79Uktd4FGVKBztJ9VHxKI9BoY+a2
F3lpbIcJY6B0+HuduFUF1k+H755hCKFN6tBXlEHNG6Ez8HiPf5u6krkaFiU/hcoJd0hRrD3Litlu
KgsglXYxjJIq9bxrs8IPQe0b7SpE2FfOIpeIw5xXCWSY5kaVkQYuECjWuYRVABEexD669jpGrQg0
6HHgA6gdZ6OxebqeZyyXLTDEtyHyJ6im1j13r+VrNkAUJBvtdVPWUc88jlHs5LBlxgulz8UdIcvz
im7+qtH/P48EdaN5RN7i//aBsckfq1JVmqYeNnfxdJauNlnbtv8D45td2BjFQArlcEfE7PfDZ3km
gsDaSrLV3wG/iCM/lPts0we1bGQIjRWiFZ7U9i1LcykoWNA2YOH5ALimhn31nYenkwVmPFwMSm2t
7Gogm5MLxf7VsxTU0umNKCELv4JPPkVXywy8MWemTZuLBAf7+k03YHfXQCfrtSXHY88AiuFCmfu5
a+gTokYYvexCCmj4nqNx333xZrWbdmLtsVW2DeKAs5mM+9NqzYP9PbH62r0n7VflVVEZO4yiWwRm
mQzqLrZrvH96+3qjAf6isEN0TcSLW/a3z+Cots3/eJExwIi0RwhjnIZtqCJn4SQDFBQVbT91fqxh
l07B7b5EXtSPSY/gSXgKThV2zp/qhdn1MWp9mtsHikDgovQfxe1K1Du4DMpCKU5dNmU6UfvLSOu9
SOK5eipMto8op4l8lFNFV3FzZ9koX8midQQZyy8gPr44uSS6uO1UvT5zjFr7Y+gV513iujHPtjWW
v4f0CpDk6atwIexhb9Ae/xn+w70FHVOM9uu/L5IC3c7IaCCOq/4r1aBRzSiKRoDA2N4DE5KouUSe
kdnWokg7p1VM16mWIxcrUYkgZqRcwO/Vc2F/sTjImdCRXc/KnU0uCFdWhpNhasc8L85rqc76HIoq
6ONUmFGLZEtpH7jP2bglFNzEfEiTdL4llkDGnNrrDB4U/y2HDX+hM7FrXQEdUcQF0S1BPiU+fggm
dQ9nI3uEkRqv36SB/3MpuL9+T0Gt5oDhodmPJaHFZ5OR2cVGox8C+ypa69g0fQ7vYjkNHekNLM5s
MuiMr8h4n2ckUlIk8Dk+wlvnnwFPWjHRV2r8p/nOz0yq7Zfoh5ivRU2b06oagSiZOq+P+LibBE4i
2g+AK0RlqUwEvvyz7Sud+bVeDf6VTPf0+MYHD1/hXwMRZB2FXFZzuh8gsKboM58Q6t2mihkDbKJr
qguJJ1J4fdviedCJbp0j/Ujn4h9vawN8wGn2AnioiBFjCVPbk0876vxQoFhgHGvx405Q2w/5wD4L
FyvEW4n3TPpmWQsPLU3i7ywQOJ/xxYjrZZ6K1mZjRxWFvqEogqmxjas4pEZswznDiS03Y9Haa0FV
YKMud66w/Q+GMnYLTY+ldNycWWJGpCWjVCyfp3BitqOLQqR1W4JI4FhiBif49a8EbiFMjhqSDAgP
35Kw+GZgFHEMy5CEwg+QHPcgVSgOkherzl92/WkJnYNubN3QZEr8/4deeWvwf1+Z0pZpY8lykXD8
xRMZmaKNmiMDguFiBFmC5/HJEqpbCLKpPD0oUHJQlHAeq4JJPlGxKoAZb6ffPqhLvgSPGEa1ok4W
1LrpadHXJ8UzKRGQEeyk93B4oZWCXLIjnu2E/K1JYc14WHxdCaACc9xs3tF//WbkvF3rqCyDXFAh
nLgYBHE/pmf6uvntjFWSqkJcxyCcYpf6cSOryQfNbp4osiJxfLVMGV/5hJ1SDdN+j6negTDisBY3
G0pAb+JrQitBZcRAGXZDZg8Qv+nBVyajY6fRqRK1PADF8L0t3HmkcFXx1Dk2HipslWrECk78uXGM
7EZ9QjrN8lvQa7o+9U+bTrd95V/uINux6X4fTEGu4kObeoQYCBm9/kGLv3pocWzPs6uCEPEcPpxu
ytj+cg+5QOSnQPtQAyuqBv3BxrbgLAdZ4Y8yHnJZ1woHuqS7Q/qNi6kvb4TKjOLzxrL17DEtZXrB
Iew9AiWI20wvAQmaodF6uXMIH3aHZTrMX51oLFQA7Z/4LfZwzRPT8r4yPUlWY2FMm5XM2ALow7Cb
7yJtNm9Jefv82xvjr79CixPx88C/S1ialwxNZulYXxZy/Ftz/DWDrcAtgGWPIEfkEzDCqtxE8gs3
KNkQCIhH6siIoHNoPlyFDZrX+GLvPu0QMuRO8HRBIhRGGuuV9CB1vaNRdOVWWIdZW8v+l0s65/MV
dWqRLWNn6CP3OWxrwlJAGr68psOuNAb+1J9P3U3jrltLZdUf99S99wVzIFK/fG/zHE1VsC6fuxhl
kNF9s5iRPaqnGjRW9lLcJP3/UUbBZeBdfYLsCKMMl2TgN7GK8cUGFBbqmZkjhHZ20QYIdE8BdXM7
fpBmdcWpM6sdDYQsokjyzZSN7YRn3OpChzV9YhRNNOYZH4e6zIrCDve3anYYlfXXo8kFIehFLR0U
sNPvuAhC0vRAdaJ3IDw0K+Rhna0SrVhq3MnSTXgH41upOsLGk9zXiKomc4eJDaWfXiANu8DsUT0p
5+57mKqXkx6hfyh6ULbRGBbZfcb8m/JpE/iVVvk813a6W14GsS5Cr1ur4mnis9zsnNnw2nb36RIJ
Ds/DgBFzr/h/Qk/uMSajDV3AHjQX+pve3xr+qB5rFbNg3dOzMMs7EuOcNhIhmTdDeL7Te4Grc4GL
SsVzYShsid5Bko7VkBdjMSi1zd8BURdmsWWOEJwJv/ffqnxYLOURLsmtCnod4YLSfu5XkZATLegh
3ioU/za7hjx+Nf59S05z9oMpFuRqdxoPmEJqCZyvujGFQuYpXj799K19KCxb1cpV0VkEDcp/UVtz
tfdr1PrfVFMEgHcK6gA8zl0JVr8Izq4ZEaa3MZ/BQ0ragVl3il8/FeoLDVf7uhDZqFuf7W1pLAaA
7UqjrF7hZHNX2a00MsOj+Wu9A43+jJFOHbdssFEP/taC38bT66oEyLhvQbd99vM9Z9wRxAY1RZOg
so7TNOk8wectS1rEYrcWdeIndZculNgO9WEpjGYkc7h/YFtu2Y4Fb5xP4KmSD/avBGBcD869dVm4
c81bJ/dKr/yqFwTJuIrKBtghrctnnmClZP2u+niAJupOlrNiVv3LNg9FVCBkp6q7SBLU079MPepg
Dm6asZeN8cSnKlKqQRJoD9DAQb3ThdAPK3BW9fK8RxOuAd1krtYu4kwvKSJ4XWH8TeC3fx87lBOh
dfQ+VSoRb0dNc3291cg2u8uqtulhjcgV0iy24FYzhwMijYBWc7Kq+EXV6k+fgfoI9HdnS7p7UhlL
7LYsFovSgqkfdZiSNag6DfTShVg4bLXa198weJOtnjqtGiuMMNgF1dz6ZMVpGG7jYFjoMSYq63OK
Js/0vPEHczPNamnbxg1HUrgoQ/hbydpcMwNu8nbpEh3r4caBDsNKw2XCMPthxIy/F2BYgE+JJaA2
Ds4LkIkosLaHH44rGxwXv6YeDd/ACP5Mn/sSAFlDbVq7wIrdHNAMX9cEnZMtBNT79NN3mmgskkOR
Z64sFHjjiDb4ZxdilZjYFvKVDgQxZwh6yGCe4JCZzL9Q+yOlVTBsn9pHOZ3rjs1wLK2nOUXh4Tiq
vqmwEaryQC/DmbjizJTNuTo6YgyZizF31TrLUyKJQ9x4Ec3BmWhq9yn2eT+X+Afg08zQNt8hriR2
9WkuoToKhK6FSozGqVR3bVJLkIE7gRR53ndCir2pC7bFUUKE4JzIBzKU4DI0qQGlbbXKm87x0o3q
jjVztnmGsKGQdHpT5Eg19d/wYbGMNqiPTQqkSVpIJR6GLPc0Kx01IDQ5hmkCahdmnb9bPj1CHmDt
vZKGjd/DTsuVIjpRSOh3kyQIupDeD56PxIQbeW8BqapyRa/PM8P6kdcue2AQF5dcNkffZfRE7Lyu
1R0W0hd96FOMVHDZomYbdTbvaFYovrAirb+gdju1cCZTBCoUaxmpSDF5gd6SKZ448Sx6hkZyNH4L
LBoIGi65sCRjzGL/p7VI6UglAKcnoI7s/MGQ7/3m1/xMNsMBzwbQ3ZJnFmdPDGvR5vPzAz93krT9
8g6Mvcs5TltFCpqGuXRh5RhxS1DUVMT3nOmjDg8Qs8Vp3qYRL/aMKsrE9BvwcuFOuZsvyCr6DIGw
GQwh+qkCq4sDPLAdXPCl5/+7250BQrMldZr5peP2D+b/l8IN/k9Cl3JV0RFHVUeUfJI8xI7/X+ne
X+I6miwE7X3qnukCLw7XTcYSxD0dtij3f7oMVVzT5SY2DgQEu+zCFeNz4TokwRffV0MgaELUiISY
Th3xWiAQNAuLNfmeBEbGtJR9gGC1lqvpi3PglOopRCOCs0Ei/Lj9QCiVaJD6P+WJB7aL6ATpgbTi
kOb68QxNsHut+hFUgHkw0PG7LQVpzG5le7L96sLDmxkH9lv3ENTf1las7Xj64dNkOz2gR5zm05Id
hAo9/zuZktZ2oWQurh29VQVVv4VQG/3U5Sl8PV9FiVV2iuf1rUdRxeBWw4qdGgfRfZgpGPyuI2o7
kZti706G6cPHlkXO3ZU5OvMmI+TaCqw4lJabm3GYOIyDk7j4YhUNGAUrdFhpkwfC0sMR2TBaUZaF
QdXcZ5vZ70yfTQWBcs5iNY05nkjUjVDRs91KTwp+WthxreXCmSDe0V66rD6ryr3MrTk4Id5eIsr/
pBPwLwk+pL89X0/layM71f406ZuICvyxHUmfGDQQ6QLs5MQ3g0PSqfRyICTijcH8s0mhfhlCdcEW
v6UoyZBI7JtVMuGer+htubP5FGNf037i8s8uxCA4hn+38eGR4aMw4D1CI+ELJwMx6nVg9yK6CEfK
M4Ct4IAk0JiQ7KmgOXSC3BhpTfIAntBtX6HZD0jbA1q9fhlK4R1avbDRLGr2+AVnWt7k7LezZgb4
tvndgA7b2QJR8PSVMV6+LM9XHNnc8CC+MXsRL7pWjbf/94xDJ8bNlnDFjTSyaQdUnnvd3TvsTnYJ
MHWdIC3Z4GBaV5AE/TMidOM+KCz03JSbJRMriu0bOGooIj8aLpZ8MJkMTMUtQ59+4kTDA7qtbsWP
/K81Fuxo6wzD2a16jU1XfO8Hbbh6/4M++0fhjhcl9LlxD/z1SJmvtB4BgQfZugImK5q3U6Tz4kg4
MZyoJs/SFnHfRrHmomPNnivyMiDv8ddjEPeVTi1P9yppZ0dd3xPmA3/fIft+7FQ+uf9F7hrSzg2g
owlxk4yFkQGkztxu7KESI5pdSUNTMszUzIsqVkaOMgQo7Dyf34j+sXpMOCBosFc2HRvFwBUL+SO6
K2etFp3ByvivIxfxTCewf7lPTL8c2boZHDlK86oakMMShx37Dz+WfQ85eOXja22Q7BsVc7UPZBma
XV01+5hO6uqlxBSENPZKRf7KRN5DxElgc9nLm5zs86Wkytguu4AMGRPILdt9k5EkRj6J/VpQdN43
J6YNXIECwW4I6YcTfySnttKAGT/DOv6gnu54SRNN5NItfALVuhgOTGKkFmVtT99uIUO7oTglkq3K
1fnDQfz56HLuk26HC8yspaxkBVramdy6/Jh3z7tA4NkNMaWiXm/lot8s8qjpC+zTDrPImzdlOEwn
i9BPHBOuOq9zVThuYy2uUYPqB00Y2lox7gFIHvsbuPKa25KMbrtmxDzyMkCp8NhFS6HZfXtUJAdv
aOHa+h7kEyXxFHmlo0FHOLelF4FqPawwhKaFCUsWzJnQ1fXqxP+DQ53kIVM1FhOdnaUeAu55TLd0
Kto2wLxcuItFvJn2WitPxSIvy2zrUq3PnbMlsqsqWz9zhBc5KjcBbRE6vy1vEdysREaJ3K1GKLmM
a74Fv/BxeEjXf/103dJ/Q9QXFwwFNqEkh+iCeaQsar95akA3UraeqoDqGVb9gsPE7GjfNgsTEfgm
adMRE5EbaYXTEldSgvNokf+bOur4DW1F9OSTbbG/F0hxPXMfI84RPXI5t6oPtOgxl17TgiGdupUq
cqtHe2bGhR0wQ9F8LNEP3x+0xBOCU/qiIMlbmFe39qdR+VyLz7HVDZF2HVLi8nPz6Lk/UH/+wt+u
KB4jMRIXcLHzWfkb8aq92ppZXJ5cho3T0hfnpZ+YMMwUt6upVbDz2oB/v9Ex6X0ZIKnEnmwZmxij
RVNfvW4e29aHf9aYi48745yroxmYbCA9zX5yvOa/2Vz549dMCZIxQ7mUD+m5TnFBOLGX3FUine/e
iUIpCZy7/MrqHVdM7WYXIOTInUfRDWtvxhIMpgSm2KPMaVPA1mA0BesZyogtZfJvPK4Tw1OqXxXX
wba6t1s3oSgeCA875cg0ltwkKAfY+oCeTD2kfSgffoMlzdz66OVeRRdrYSCcBf/9xkTcGcPKEQD+
NbA8eeaqVBGT/bN4byJ/WcEuCfHRs1lSGGkDcbpZxiVm5u2Ab1z8thCYtw18g/h+lWDDaO8h/TtU
wVghWAfVoVQ7xhdlYt3pQFXE5L4EHsk7KKjpokiHYWyZW63qcZ5TOheA8xJDeOICkwH0xrtdc1PI
hlX5fOONxNrM8wNvnTFugXYGZ7Fj/OuG16Xiu10Hm74QqO5dBm2ro1YA2T4V7jJX0jBQTdD/btS4
4ptXW0ECRYzcPlBNE4ISEeBe9t/QSmohSNdsmEH8MKcf3DScimDEhOg0l1/DeDvRNOPuz0ebbJH9
Hkl8lTs+2f+ZO5YMNxtNDy9cWkWtIlqeRo7Tq956SZr/tMLyImoLI1azDzUVCeC3fNRPxrTCUAL7
C6NXBdkAYmJE5oXMJAE9y5bks51cMcZmvgXP4G1mYNE4IYbCSqAxl6d3fBf36a7JQdmH7PPUHvoR
tcYMAiSIrTvHw0zkfiKBPtaKVPtDbch2u+4ezvTdsl8US5Rmz3bXGhAlU5sGz8Fs27RjqU8pDKxF
Epk7ItlMqGmwqMIV0zYam6z1d4QCDzr73ec/gjISIJX5YMMRq8YfjYKvcfa8fOJfeZXc0aGRBU2u
GegudR6Bosg0IFsUvl9Xixnx9rLNiXWwsmWPDkLauxkAKgyleUlui38LXZ74JQ6Cl7VpPiSQ6KA8
RIDecJU7Ltwwb6ZactCeExc4JQq8zpXNNWpUDWR24lEPpuyclT0HoxrG8pZeuCctA76YQgMtQ+Dx
EgkF1ldRozBsTtAua4xsHA+15T+A0fl1U/QXiimt3lU2qlKRBzDssjqz5XmYhl4TJA2F0J4l+7bv
FJaGFzdzzcZQBUSdF9WLkDLnRvb7/D/xMNy/dkXzv8cqiUAsAeXnNaGDH5mzwoLKnP/8/6dLtEi4
kbJFf+t6RYxDWz/W4/7hpQzZ5dXc4TnpHLYkxl062K+lScXzmcBMKtA7cRY6jheAaI59lQSQRPnf
CtMy/UtlrERZLmhR2s+xdMEqWCbXGGhixDdz6YPR9ig2ak5wmPfrnKswOh2M58dLQOzzhNdhnNrW
SlLnZ43cGj+TW8vY6cgU96C/AwofYAtNtplL48a0eAWl9iAnhwg9nif/vpeqckYQE7jrifbRW4Id
+8TwvDCYM2HWm/9lVADCnPqQN96QF7v2DLcOv4AbINHAnD9xb8O95PZoW9Gp+ypPW9XN8ovCVODI
t1PPQoxI5la9hBcoE+CX31ZkrO0TZpLbgCvkGhE3vO469+9/roLNlmWjstVs5FbS+nO/fWQrWSFF
hbEI6DaPk+0lqfXeEhwGVfsP5QeQcJAGyw86IVfyGfFjzwjGeqi7wrDp5TW4put3xqPQK6pP4K6m
t+qjzeiTVZyoIypSU9tHynAOYO9AIllzTce6rQlBlTv6oCEOe8VpHIsq5GVPSKy9ymDnpv7zOZo/
9gZpcHaRb5pvNw3RdvasjQcAiO+6g4rnuZueTOo5K09DqUlZeaDDlhC8o1rtROp/9GAJXnGdyW6s
Rk1yimaSGGOTg0uqykX98PtYIgB/VdrkdD4S44Eoy2J8YoIQoPBCKHtukt9MHCGDEfInd5YyjP69
TFPzP7CYRKxN3iiqyJ10x3ooEPYG7qp8l/9EIXDuNSufV03a6TS/w+cBIPWBHxK9y2cZxfqjpO+7
XcBittzuZdulCp8YaV99uBu4axkPNMVkBF5ukefLhUukJROS/B83JJwccmzUjZqRswln3vkGG3d6
a0TXBAcO7TgKvMoKSCj1YuASzYMa/UNVli+iaxsgxZOEUYotmLGJKezy13hRrXVTm4y+cp+5jTW7
3vsBhVSNiKe2ikJ3aX5i/8DpP9CVDoHiucRPDcGCD23IMIO73bnM5Or9kEl35f66JcQl3WavYHeM
5RgRTtYl/rnkK7dX70oxiYNVosXxkF26mhraAdJV9fvp1hs1HgSZHPHhax+WnL2UtSyQEGqu8wkw
WmccffSccvPGyRy5KWVQShqKCHv39VaSLbNnqzz6oQuB1AsC448+w2A4CWdnh9n4vhdNsoiRIfK5
cKuV7tMHLCXOt91CAgwIAvbOOC/MxrzEPPbeaUY0oPsViFI59VA90IxUam/O4x4xlN5XVmP8LpKH
BdKs6Rs4RBUJ9QqcgLx2L8uAcNMOALSLC85tHMbC7PPuE3Cgwf9XkqGimO4DfXtqW1YUJeNdGeLk
4/G1Zkrq5CZb9UyQ9r1PCqQGk7Wo+x1qSzTwIu7Fc+CYXey98vsXV3MG9jGaA+pO6mM14PbLjO7Q
IdQtIIKyX12pPrG0GtEMDoOmzHZmkpKuRb9wRXW+4UfkVKxo6EMUMB+7htKqTk0kHCgM/tckmvJ1
lI1hz6KEuKmh2luqZkrrFnumy/xeZYN0U5KMPwjWFBQDnSygupQAy2mGFHjKp8z2bdEMyYe4b4IC
JxwTpbxx/q6RINOCfdWxvDeksyAAKMdb8Jep7zu59n2XDbHVLieZ+ucGy6jcdNcThpWDTNqEZg2d
PkFJ6Ya34u7R2NZGKHPX/Sk/yIWQhgEDUdBVt0usxzP4y3S/xC+zNxJynuzSXHueRvf8EH5GHOao
rl99/QFGo+estQOjacwN0qiH0zeTnuKTzPPxiIjnfY9Mjo6MJG93W/6drigA/fxiZTDbqM760kCk
lDI4GRV3gGwTL2f1cSDV7muACW+X0IH3mJYJZV7C/LoEbeM99V8EnDY5A5gko+wYcyVnPU4/nILu
T8rSOdByx8B/NtF2N4uNdx5e+ROBV6J7luq7vzGNqRcAdc9T4CpayaXygaECfkJtFnLn+BsrZ2WY
dpDbRsSRPKEj2rnAN8x24L0t8hFJStxRoySL3sw/1y7b9PdgHJllpnZB6L2fux3BnunPDUQ8Rj6C
Vc68gKtkL703831ACd7BPkyjgTx2NeIvM9YsNvKxsRkKiaY7HAFqMVffrCwFikd53eA0ea02q4zY
SGVsuDvBWAFYq/P9LJnn1D7RmFprRZrEhAIeISh5XLjubIk0fh/xBvtq3WjhS4BRbQVxmgTSXXfY
f4KkR2aRXxz0ipBGwzvqb/e5NYPLAkonl7zU+hZSYoc1Eohw+UUjTPfX+G/jIDACx5R8pFLSNG3a
ObgrENWF0qLrNu6UMOZUvHc9TTc2CDYAlux/pOKz2jVLz0TaZ2c0hUDVnhd0DlRJiADgwThabTFp
gPu3LCls2q+VkwMidmS/HAL9bwiU2yYiDDmUD4ReOBonvPFnOvN47l4rcXX29kCwU8EsW1vjF2QI
DcyepNF7Jhm8I5+2R6WacdQvi+zYQlcL4q9IgmHVkUbK0lBVZUVW5JISKe++BrAVWoSStqPtPK8o
FH1IWliNrrtnHQpGSZGn2QsFZsz0dBiPbqMtfoxyKLWPWG42zCrpi5YYsmi345kLuJ5RtWPVXrM9
cs8uDGW73WlGlvwrPFfulLtz6iZhZ1z7rAm2ZoHfnUwVzNt2t8uP9qGgEq5JCgvAibA9y1FppJnB
9VR994FrKwkOBt+wTz10ClIAkm/PBQXGiXLwPw7i5NED26HU4TFF312PI7k0FSbMKJJVUMLwSu/j
NvMhzfkwByGF0lzv/kUVIhWHMmr0iLglYcVVUsM6iQn3yDCTkMT0+fVCjVuDX5DldU6meDFEzx7k
MaGmZyHpfHHRiNpX82O5LhEaV6Hu3mFXoTmGwqLc6MjLRe0/BNxvwee/AcQAqcXz/EZHmyGijMoA
UjKD1vKIobHrauV6fMsyioB0C+5KdSrKI34EgvbVExEaCgU4kOuoV6T1udJ3iFLb3hQKEqpf08AM
15RP+SKnWQGPxsz/UQtyzABIBLzauHIPpsB7HWl3N0PTtTp0PTPhXW/P9inqP8PtzEsiTnaikfVq
koKMsLJQFw0n/4IA7BSN2OO/PFY45od3m/5y9/WAFd3QP+dnYBNydfsoQx1HnAE4xEec7AQDxD2x
zpG+y0/Lz7qlE9du7iV5sfk7PTuAuU0nhFaN6kn+99PAfVfVZ+ATo/2coJ+14EQHzdWTGOnryLkW
3d+bXghxQUPZJgZq7Pms1h3AZK6449WB01L91BDBD5yZFH5B6LvNiqyR8b8zaIGu2URE6+0T/Scm
3/+G06FRxj/B3PlNiCBHANhguk6AK5x6FaFuoUE/SPPvoNL6/ZF8SdnYQg5UpjajqllDaskGwwq6
csRzPbGTc2RRe0Y9dGadfzGiBiIID4zF1sTVc4PKKwD820A7Q4A8Et8GWQ1gcf9a51WFMQq4luWL
K43B18ziG2Z1f1Bmbi4K1C4SWQRgbzpiTh4hOjK5p276MBr+a5vnelCMmuJ7ykmVbPqICBeEZmZB
O/Iy6hMm7mzIzpaY5Qt9Rkf0TsVLgG1AKNx8ORmZ9YJhE1oyB0h3sK+ipOUQLoCVXv2tEq9EWYRe
AIuMaRMSIuEHa8MrzOnVTBzW65uzL9yKCyX+Myo2f1oHy01FFenSKmhdg4H1QoqQ/AYkp/F9kunB
vgkPeVqDICbiCRL9sNJ6TsU7+u5/VmBKMy7BEufGvdTQcvQ4LLVOnOkyVJukSD/pKWQUFeYGUUqa
Jz/y4s67nt5rTVLeJYkDGhbdRI0qDhhwUXBBwCWSDLSy5GYWm/LTujwbWYRHJTUVT9LnPwu5NV7q
INh7SIQKSV5fuKryvPK0qebwrebe0fJsdUleFsPTx/Jk/kTUpvApPxfZEfHWtcGwHCRacsV3oAdc
AQnD/t6eYI/nxK9TTUz2NDcg/hqq4egLNQ4xHzy4xc3ED0kZA/MYnOgsiULiSMaJVrb3GjulDyIG
NgGc7yCeQfMrdV1RYgMm5HBemMfFfVoA3w6/aFAdFh7fplms/Sxyr4OxEOLZTqTDjFTc9OztsP8O
KfRaXjN745WCM+6NXsFHm68T2eZhCYCm75ZALei+5G5l3nazGkSXOzoaTFBOopiYRnLqkkimR1XG
ThOkHCDwOUf7NjbIzhW799LgZwAdQ3uElrP7QEZslKe5U/pfd4Xl4VTeQ0rG6MRg9LOYm2LyTLaE
vL+NmH0rHgXHk+dh65qKPnIxJBCxO0eWQyTQEMR/n0fPAjO71mzWOkwdSEPomGgv+XziOPJZuox3
iWQlku7o3yRjLd2ywfCotK9R/e/Mx9UMDwCS0HsbhsTi+Hpoab0qNQ+SYtVkHEP2WwN6W6zKBxIb
9mhxOXp/n5oP6N6fjk+dV1amYIjf7AkAKuFGOGtleiv1S1cQtwPdxNcZKCF1dafQOdep+JtcLFdm
yPXCDV9TyvZ/2fxgXrIEVSsTnu4Dkt6ORhq6enR+zkPs6cgBOQ6TOjhoicyru4ou/GQFmAclGzG5
0EZQ5+akbSb8wxDFtYXZPhDuKwNWXK0vhpmj8jcHNx4r6kV3ACAdkZ6VHqON6D72bt6PcMgMs7zO
/Olf9hWNad7uoncX975gWTGzcWwXSdldli+Zb7XbISsdVu9Jf7+WHpdHEwqwL8rCXraX16Amyy5U
vcpzf7Fw+97wS4U9ouw8MJ3ReAR2+fkiAklqwqL+g0jET7Y4OYMFPbKWBNEcwk6myi7qhgBJVWzW
9O2BxPVSGGntI4iij6rSkyHrvvpyYwGE3huSEc2tdiVf4WyJPmH7UvF1fvYz83ebRgnwnR7iBy/j
VSqVK10i1XiUGnxoXxisiA3HYWi+wktRYZnv6yDB5BTtLINhhdbTsbhxbIKF3lLtv1QfT5438ZYp
Gx0jlS4zdoK6ZvwAIcVbAglgAPlHQec6qJNjC0Ts9WHOa/XnbYqDpf9XLnlwcMghFsEv20BHSG4Y
D5UiYWbbubHPCMxrP9Ww/5DSPkmXP/cqZ3USn+6G9GbmhlI79xoNVo/FfVxCFshi3ef4Tr+GLbXU
3hOyh1woutXtreIpCllDq2E7JHml0Op/pcgN+l4ahIRRkfeQ/EdXrEnCMBGLl+PgRoz4oScYo850
h2fOb/u2k9y/48klN6RPzpIYxilINyr0euSCoctODJGgQWbl2oHhHsiMKwRwy8pVflFR5X7EFNTQ
8SM5B5qK5gRel+OXflMpVOEJHyq0828Zzj/6bIWJcapeMeuTqfcRd+Xxfb1QO6M0w2XTmC+Z2z+t
J77sS9KAHESMUoDAS05C76YkWL1WprfxS+yNo4Go5dVD7H6aMtAc99yfGU/SLCwVzh4nH6vhV26f
pUcDHlRwCrux3/85+RnRkvNTwtvXecvOSDOiLzj5WhPUxQAW+nvkOySn//YSBKzSEoU0/2dAXiGh
bJ5OH2V004RvJHZyrbNQZG1alpZ2DkBgQiIk4kFX6XBFpVWYkylOS4AZZm1dchyoavBNrW+KRdjK
6UvKoJyQm6D43dJvFuGt1FYrUTnyk8OoUGqFmeEXc4mEtYkdvJ5lPuAccXageKMxaioe8UnwheuL
k5xJ3jXbo2GErUsxK+D7Rz6n/h/ClV2r7hnYpTMF9WsLKhwX3Pweb+sQdKx6Rah/rS1isPhPuCGN
7g/cxrqs3mwOXShDjaT2B9DctsEBm7iTXp0A4pxYRYgX6liEa6GTGxgwta4efRYEku7hnsnmgc2a
MXoMLOrnUr0n4RLfaIZnMX+t3dAt8t0OiW1ByOHR0v07zDSwsQLZPoC4Fxf2+kyoXHUfKGPym5lF
WH8dnl18+T+vPoCIukhqxZfmA6qizO2qzkd17dl9ak+eGkmXYS1Pq/cZkKwrgoAjF2h8ghht7010
L9+fOy1LdCFDwGrU7lkhbRWx5OEcFnOXSJD6cmqX0900WOn7U8T5+kg1cbCPTXSEOyQUqeRfjFde
l1mgm5og3/PLKdUGFinxHFCgvgUy70kp+80SzGMDn1kEIfmybNu74QJatwjUH4pmYyK0/5oS6LBM
ym1ai/y9B9cfV+5SWJLS/fBkz4jg01SZ5TTseDb1/qh6+6WreHUWYQKcEwUfLhxIK27vT7MelSCQ
XSqg/fbAu9aJo74fS+RJguhz3wDMteymOyVFF/kxprXtMDzjVcd4AV54+pfW407U57SsDElQZU+H
G5/re/3vQNi4trTQ51ZN6D3lpo6nElk/+nrJkwta08rdBOdhkwQQibKmBS0beWSfjjUNmmjW/Q08
3zg/0x6RHUwQ5pQGaD0F/emmehGEjhS1i7kXoB3AtJAIYCHQE7kOuEgNuWBjPsOCElifEh9MSK1T
US7Hvuw66jla3oPDDBVzAAwnuu0EtQsnPXcfk7dk1K5KHTCadQaKNDug5ZhPNOghzPbCSqJfBoUh
6XmGX4L+TLHwZvLPWVZiuVNKlRS5r0uFc3LCAb0PFJA4h2tv72mRDJjQmAZ7Y1C+aF8tw/wo2I0X
HTRn76G3cddKeY5nViIjTniOAZ08xylvL2NcafZ9RXdNZoSbI0ruhSjlR+XW/1sWVMTJCvs42H4b
jwn4AUifibYhO1MN/7lgDSotro8co3+UkqwXH+A2myLUdiLbITesdoSySAgjErqw2exxqInP4Tbt
sF63XnhjjBMD0Vg4lUi/R4wU37GIeX/Y+BX2XaoDnmJ8Nexa1c/89xa/N3Kec/mklXifK8swrucH
xbhAJPju3eK4La93K64Uhml/IrJhfUe36E5vQsMjsEE8WgrRgO/yqPhJxbBKAtJyw6eU8pvLBfmN
d7nct2QsNb7FYZsLIHEpaKBdWXyoE8MeKk2+kbu+KJT1QZ1h3Lk2q29TQvR6k/vOQTSr2Op91HYm
YNchzg35SWSXDUgVTIwiry/BKYhlI3wzjsjnKOYbh8qagTY2IBkY0kzfPdFIysqEISNXyt0gL9Ul
L1FVyT8dXD4Wkl6B2MsS5r6b+ZNCDcYdqfN5yp60Zlom+D00fzSWyJaD9XElj78nAzmRBvES3mr+
xGB2njNoKOCoWW3g6vAkvIjauoqMDbwm/mjGH7U2aWhC9IgeX945eQZhdAoDAvqG7Ti6HKXdecGr
+rSA6ifvs5jEUOQeOR1a78gv9/C8dM/oFyIZcpVPjMU/YxhMhGGfjH59gk17YXEKcGg5Ftqekgsn
pUVCiERIc3tbqQk0TGFTmX9VKKBAa2Wy3+hwgzbhg4KFY5X3wYgYVSiz2byejsaqpYvthAIrwV2F
Bzzjd7J2zyLxlJ+18W3vKg7z4oSguKfpFiWGWebUsC+r6AMdCiRc2ErfSnY/hoTiQoZImcZy5kD+
y4UYfJy+nFpParUMsyDygNMjXBQ5gDjslb4ToemLUWqWjfkEzXqCLwTJH3OzAN4Wc0U1ce/94bqy
Gbn54MaHBZZY637x7OgPSHO3bd0+8Od6F6lkQBDlZxhgpcS14rgG3Ql9h8U4ZuW6Q39/HRtxW2SF
5a1zlYZbxax5+1Z0GE0TT01fzzReL9pClUf1ifaqTbIb2KANAVeAAabaQglCacgmYIvUB9yRTvuN
clcIJwM3zut17/J/K+9OLZgMcqu1AEUWUPJHBGMVHMvM+DXijEq/Zht1Wk5p/DGpCpYHXiTDtGAI
FOBBjyaq873CGJtdfMxXrrG8tkOjTdrRWGyLYIEVFPC0Op4H3MsXmGWRyUG7AD7bat0ggxUAS0vC
J3ocCOlN7zfN+yiaFoDiKKMSk+eeqCalBuwoBtfTpCCZVLKk7iP1z0uXzUJHcWaxmjvviOfEGmDv
FuLWTAOPYNJ0ycaelOpivHRRyfgitf99p893u0Ze7RmF8X1LYDuvS3N/GhO9eB9q9yweFqKsLgoY
BnkkhFysdIHZ5djAkvsmAZXDKXGfd8uKj99GtCVoMluUMr2Ui++UfhmHZpa9d4Gp0I8a8707l6iT
V3hg9hW53UlfrUkjJOvRcNLzZoXjO1A25BAfTRzlKbF/ny0ukojSS1d/yfgGJN55TQafL/PgK/xZ
L5lNFkTMmPiAPUuPwB7pjOxj7DGbtKODMeMQ455Rm+Czzo4bcY2GdVWJGaOFHxachsM1guUxOk+u
Z8NxvtpbVHOx65bPUnY78hcNLgBmnkS1Y8lf6GWSOk3t0H+N+CPQotFxAqY2kDbtorFefa3DcLUE
lQpB7KpsBUoqQAD981AjJ+e0ms0XMR5GH8MIqwflfIc+nW9RH6NRHqK4nk98UQyy8rrqxW2YPjP3
VcbcHpWyzhLdByaQWBYnMciPPOW11URMV5HDaz1hyvOuu1sd+KbHq3Mkteg9SCNYCEf45tPi4L4g
pxwT5JPi77Sa9345nqYukMrZPIxnXyy3e76kUi+mlDtPn/qeL0VYW9DgKmLeYN0c7HIih+vdkOiC
bHlxuJdqjEor4ZSqTcqgLTM7637tL2MQWxHLrGZgsn/QWSeVKq3CT/wtyHX19tXO17sgPSe/OAfo
Unm7kPC0VdFgPr7PfdJAj9tdJB/xI/ivoAWP6qm9/LPyZ9pD6dhuwVgtNyDfJeakD04F/v74Pw0h
ciTifpSsbYe0mIf8nDPmhKGt/yzaHge6eqaP4JpPBwnMksg8IyHkjjkq4gX3//ZYg7LJh0JYxKYC
/UICZtyOKSR73j5ViB7hge8V9YI49QChAhunBejL/x6mLOXPmOW/swTaWLVWDWYSWAKUtEL5HtlR
/e3ajN/KC3ShzbMu8C0lBJ+BFL4hU0Xu2w6yZgU2VvNdk6JmyGYPd2Asv+lawfOMC+5qS95vYKoM
i8k497/vl4GbnbwRURPCSfhGBxMkssdQF0Fxf3hgVHW0k3M6BLgsIZ+sDXUxUYbei3yaFTolj3it
ktqxd1W3tsKvBy6Idnvop8RYltrUPQFznUIYB9LHEYMpUcwdSEyar1T038Dkgz8aUOroDi9zfk2c
pC8kAAjmPtbXnO3tdi08rOFF0vZUo5qriz0fijqYRVGipvUSYcORrCJL19E80WdEwFG/whCasiX5
/xN3/ezmdu4RrOyp/vcxQCpI3nS/1FgiRGiAtFNFb6ptdd0518H0AxFo7ioH+X4abt1qQo6cHHBa
VHDnxqDv30nB7DCDC4KefhC4BXTzLFrSr42O6sQpsrgZ4FSyG9Zl/h+AB1eEZ8KD4kZCXZYNM4Ck
QRPy+BIP5p1G/e1zbRrAsGqaDAL38sYP0pSvCeoFobYEvKy06kMdSj3FQngPVxJO8t3Ihfny83UC
A6WSDYRt1uwN3gokTyl440sbhyFJj1jsj/aJAdlrMXMC4ieA9VHSdlLBPOU8eSYRBPJAONHPWBMU
R9gSBzvoEyypm7+SmRDSHnGRiLY8unqEjKBIIOpTTeFOCop0X4HgEwV9BQHzNMbGqbZCqB1WRWo+
1IG5i6RYTy3wxFzzYHPtSlDopvzWZVQj3XXcqSFn04+Puj1ggJMUDHnVz84/a1E8K6myfezFgJOK
bc6UYGxyfExJz4jAjGAGyuhu61k36qubWtSECqSKsUF+cepiBtBYX00fPPdHstN9NkjvJuQBfArB
uUK048n28X8KYdQw82BdP9XLZGxzLGMpuclqFknoTIyFBgFQcZrac6eWZQvjhKpDKvxGM3MGOHvz
a1lFKYdtlORZ0OydUEGqcKqLIkng/37yYx4J7UtDD2PCjpL6F0yXnEjeEWyP6vUZR44bDxjsyvuP
Xef/16mxaUGjw+B+t2TpmGlMN6wiJPqc9MGzHx8hF0g/5+IkStylsw/5BfI53BOcSzN7PVG2jPnu
aNJU229rwNyGUgoFoCoauj4ny/IRGCDlWdXV1xgpR8e232Y5GhItIVfW0ynSiS8pAEU7kCWnFQiw
lMZCZG3c8XZfcvLfNebl63Ky67a1qUoPfxMntAdAb15fJYluC8VNN6DUN7WRlqig3gB44Clq226c
rQACSEdSnkSoOL87uApqoy1MKrebG4gzwQ1OgkdIZyfGxl86xt4IpXqBYd69zXxjzVCsAWc3/a0a
zj6Ng6N2qPhUxJH/ztGEIazoDhf6kSbNJNlbHw9tzPLGBfsPEpHRboPaBDmizEN1tEtyjzSOnLd0
YZt5BK9rt+JlUDVl33eCDKGw8aiPh706fd1sHluczP0cnbnRcioW5Ra8KNEnif5QcrKbMlanHumL
GT/HtLszmVjcwSls7ftUhf+4SvRkIUOsX7iHeJPOBIwSFzhXXkQJLjC0VXAwep7W/EwXKBJEzJHH
keq/o9oJKYjAJixDiWtWgmcld6gSB6mUuRVsTbRHpkq5uJC+/bVUhI9G3MWEpTl9peSKIpiZ8cVL
nbE8Gj6B0n5OWWQQIU/obY/sqznXF6507AVen+fRhS6+UXtGrOY/q2/O7OoSmUMHCQAPUvZy2fTr
wYzjQnXPNqx4k9FAho1FDBmSifRkCUksStritD47EYvJPC36W7SMTcdt18PsrhIVPb+zFAp6yNW0
s2Sgd7eOhgxVSzC7yu7DpNvrNV8IPTKPKC+1zoo64vZVQ6LlnUzn+O3l1aQRR4kMI2/aZAel+aEp
yiVO0l0yNeQYJkPQtoJheJU9u2y4Q9awjn2TxVx45/tKXXlsE5BtP0lFfndtugDPvfkiP9BJKIUX
+9W51nnE15y1CUQ4jOhgDLAwJdm6VPY4n8Vkx3v/xTSLJnuocOLA9z6GYWxwiECwQ5uOyjHi4VMA
7xOjRZ3PnzPHMdCe+IZQmy+xVF9oXoNVwS0e4KCCnMEejVCS14d/FfbS41iOGSXmuWtx7rJBe6Mg
lNMp8lpqI+GQ6rVM+ADw2scTeGWGPdYKLjRyN4HaLO5uPaE5xpoODhRqFyLO0UT0O35KacIg5GfL
I5Ta/o212Eo4qCmgg4ZtbMnz3B3bSq2uswXyWNADCaha/xooyUew2mf3bMh5dNcjq+OQ+0EWkqvv
0P2Tl5e5bAasmn0jRGudZZCfgvn19X5sZaWrsGNcI9gNeRnpwM6TTMdhynUtXaLJeeL1w7yv4LPl
lEGtkU0DIo01smbaMiLYViLX5ZlypWEKxILJNBxMWHwRDzoi2OYTKXkbu8A04/ZFnAkO4d3xBVVt
KGUwNhKSxbjVBDEpYwCDxDlSEkREo3s6aSBQr3Ij2qNNvUDsBJap26O+uFW647UZEXONFEUjc8mf
aOJMSr9f2ODKuuhhFxRIqlfg+o2J6PjXUjTg5ljv9ykFLJMc4Y1qXkT8eTJH2DkDFuuT2UgCEhrk
hodDt+/ZVgmTJSsQnmKZuJU+wmek+MdlkKJ/yGoF3g19y+/S4LD1aCn/sYixN7jtGDHbSM2OZi/N
sKVhjyFcrzq5T1MpKz2jCIfqnVfP149jFM5u2ks+UkOXs2OsNYef9GtX6OXShm4IaSCMKCCMazlL
lFMXvH5Plx9gulqU4yq0aP01Dr9aujLly7j94JfKkLIsm6JGyBFC+VWULfaEhY7vdSBYmDSNuoef
ElX7rXa5MT5jIwKvunswi4373KT0Dr+DQoOjB1HVQdvq28ur+ANCMxIiZE9G7016+bGZiBxWgDrL
6dTDmYFEx3SZ9bIVvfLMWxlqTOa5TZgcgMoCff8dd4hGYDE7oPRRj4t4jrkXnSzKbpF8aUnxwvve
FVOwUkdTH+YheFvkByHwsugPDhMpxjpCyZAO5eEkWzKKnJtZOsU0L4MpWOGiPUi2CsG277VgPwyZ
wjGNAxCiPuxWnrltQosERu+5kgxal+vAgH+AyDI+AOVOOdPASItYFrJS8rlUoNf5zmfMDTkGi2WK
w3j8xPBJWFDAqfdkT5qvy2nzKoe3ljEiC7IItBYUiXdtCYD3oMvKznGjIWNZGzLMP6ck+wOKfDXD
IZeERmvQrkgQ1kW3seEg1JXgPjZe6a685hzA+EGsJyzIY13ZeN8DXllP5vZ9TsRHJq1LXh1zBxxH
3xVwES7HqrZOOq6uikrjWtRqyBYRMiJB7tjeHuUNY/U4Kygh3ovTnX9ryLzTcWPWZFDsLZGObEnm
lO62sqIIN0nHTTnTX60sY26r4HDaOoUzpbIrDA19xLrCQw9t5Wz9+FSfm/3TFUdQducozp1ZCvOB
fptVPIcCULdZmd3O080hsbGaEAv61wsi6V0ODw84z9j75O4EH9DkNw548eIp6h+n2Xzp1w7gPB+E
W7Y3kEF8AsWDApy6skBQ1YtD7/ckswfT9tk+bQox93zjWNjdwJ1iMNRXsitB1tw+dhtNzVG4s3LR
6VpUyvy5pFwgz7Et30ER/gdiEFntYsIU4WPRzf+Rx7B6XRLe+uwuJuQH57hIO7w6LWuBxIhJ4una
R4Ux6JjRsx+n/lGCu9YVWtsh3d3Y7olWcRBsbNwMJOOVvfvdZLU5IxXk6TmFFkFqG2AunPemMqnH
cA4Xk2khREaJt7xsjHz8xK4fSdeESMuwn4hxsX4RDo7nnXum9fcaXbX6aa31xv/NdWkWYiqjfAb7
tE1TL7HkdL25CWYra0b/1o9CZCEyURkl5nDr4i3UWmWcKzCZ1e5M3Lx1q5pT57Xyk4oGGErul+2S
oEaG7m+DYzqz1+44JKtxihZHOwdg0/BWc0F0upgkFxoFBcEXI9NAe5fslp8pG0m1+hLd+jsZkKzS
1zkLrjRc/Qg+v7ln7yqkkVLEnDm3eLWBjSG1NEvgB3nJOZBE+MUIN//rAgTewnYWE9inzZhl4h7Q
sBPNmE6vDZeT5z3McvOr/xhTiqnxpkwV8EGYhPmty7XAXY1Nrc5NhKSNxr6BMGk9TgqRD4FMefh0
wKHhRlo84pgje5RKBDPxWEZcockDTBwW9Z9yg6qoGNaiEXb6D73bskSpUGyxA0tpHIGwkkaj8MNb
5596+qaQGQie2Bb378haNc6mFoB1xNoPMLkCmPZUq4CJjBiNS2VmNAVrz7zGsZC/6S6pNfxaFnF0
/e63ADksKmA6VfpsSNOo+ly8Up7F6CQPGNnjGBMdfxe8T88miGO0KtmrAxFSIKDO/PE5gNYc+Zh7
HBVqKeXpejrV2cGuP/cIbR5reDXpl3IPdussDOUOIaCIKIDvyDD8UF/gzC9TWKmBGrQlgamU3jai
iViM8k1tbeMXWcjs8o+oiAi8kRPLWxX93BrVo82LFddlGnK0NFiQwgaz3g9DpLURBvaYFhsBYtvI
nW3hnLMFx3Q+6NbnUL7pLWH8vZpwPIdO05FhZlk2qdZDv/ElbzBV89uowZntm/PSmZpHGDCIqVvE
GtSrVjeSEP8SqQ0ntQNI49g7UtXaFS3ZkxbFVkQXPXbMlX2TUhqriSIKor/FnBORFmIROjRynMrP
YfSR0pHcr1CvVAqtupx19YGRKoo3ZofaleraSc55SPPlrd06a72CbagZVg3TQ6uQFW/fg03pe/xr
6GoFVRR/tAsf/UnaMAf4F9cIm9/kS1+cDQHNK4NU10dY7hCAmKlY1bPfnPEksfNVTvNfcWxwJL9f
7LNvqAfscjlqPXFQRpu+JOG7HRTZPG5nyXe7lD/ZfL5/QU/zOhVezSX2UNob+4xBQ8GzqvnmIUvh
6Z7QtLg6cMyYr9qa3jr9cvVuUlHAVDXyOYZhHvPZqGaDx+V5gm+fI7ZN76cntR4inr8CofLlRerv
oo2tqxCOn558uboch4u5UiqXFO5IQHVKQVBmafaCk5qg9NJF3PwAus/hEk75uEFCyIcFzf6hsEJE
2xTWw8aiu/B/OczVF429u0s0maSiKtdXyYFA597EPQExusJARiAx4elv5Mg2y4dSLr/4rSMChlYX
xeIn5HnDMt3ND50X+DDcQr7MRGGk6Eaa0vtIxD0cVbXwQIb+A6NF9EzaJQeatkPSY7IGpL8H7soe
HRb2BEB+43mnkv0eyCvxpKMvs9auovJNOYJQ3ck8dKXejL0EmN3rjV3eEA1q72JwI2qGEQGmXBPU
7+YtmaaHsp1vgON3r+urRFanZ/WGpHVP5cQYMTPRXxBX3ddU5v0GrhmuqYHiiMqfiWJHBTTvIas2
988N+Tbt2CgnE0xnGcWZavCOtlyfb7rqz5YufJjqTZraf4H9EGXVa1SHcv0tovffvgcnZlo7zVDE
v5wJ2eNNYsaVLoiQAQD6dbMfRp+FcpTXO1qecPDtAcZZrolVFDRmuR7ktWVBHqJ9wcnoEBo1Ka7d
736XDW5NKq7K0cRsBF0C+G3q//37GX+tpasz9zb3QJm46v2kHO7VRNL9tEaVjygL/CxQjmxEso87
aW24QmCBH/lci8z5nBMzPeVSgUy//JjQXCGXoKaVAE/gx+rLyHEZkf5I9+FDB2qg9mUKVzi92IGv
Hso62pIsNFg2yzhMYDHf9/HdPo4zd4Wy89TiadkuyPuBGMDiYMrNnAsFXLZs//FW/VEQCEatBM0l
qfRnYfmGMQDXOcqecJzWu+yecF7ejRdv/8Prf0S9wgpifISS38SGxEstW3UMrgM5twj9DG7orDdi
rb2P+rEq0/b5yBNWU0XFEh7CHkekdjIfgle/e0HZZKzjKi1nHpHqzYBu2wuAZGaYGpU5WmOeABL5
CfQavntyj5aKpbboeQLQtJJOXBfrmF6gsCKtRzAacUdExLS1V32dAsIe/AqouqK7xDWcYAnxE9OQ
PTSce8PmiUjVySxZSGF5c+9xrkQ3AiqY3Qzjzyo0pD/PlTZOXrqhBlwBDhNWqwF4y8Wf8v3Ym/zf
2X53/XqmGVeUqNbn1lCW835oWv1zS24Xudu3RRlGo03Gq3c0m3kc7at1da/S6wQX6DxwBNgXZKfT
+xdRDV34NDkUKSl7KD5H9JMOFumzYGjXYSuc+7P95jmqsCqV47S6QUiblNME8q//uNHpBUjw0EFX
6I0BdKmRJt0PeKYFJ/kQLCfYMWsgSswO5sAWB5kIoCo1iqkuLizTeGrVV55/TVCuou1adZVe/y3Q
LDOhHyGyAaXFtUrDOU9L19CMIr+9PyFAUWnPfFGHJ+ayMy9zUV+WXmNCtrBfxtkjEanfvT6zvT6C
Uh9XhPlSo5p/zgToVFUX2rLljQYT6318Ww14QOcMZE82jJ3466bFd830spNv1I6jV6/3wr/wVPuF
dxmfP4Nu5gjwJD6IieYWref4jMW1YOp76ly9xNxU3SX6HcK0noF7C0Wpliru4UfBbo4IS3QJfIor
O5h1hz4H1FqCVwnb1WQehArN5FjdNSR5FOBZuthUwLt4hWgBXULa2UHY6wmxPEY2GSAMp5OtcDqU
PM3fGuoaic83trKPiFfInoRf+u/KBdD/UbSiqFSLLHLqmJ8A/V/IvNd0t13I9WlLVMUFHQ1Gw0E7
QoYpNMycQtir5A3valnDQ/h+0RNWdkg9PRzdMlsacG3Y0+PjdYuaPk0CWboaEPa0T68uKDYrG5/+
WzafK+wpOvAgKpjhN8vyCPGHghRogAQ9Ml+Z2bocGmzu2t9XB4YMycMHjQ6t7Leo8ZNI5Gv2PO8e
Kr3Zi551cXqxMBnIzF7M+QfqvQExaJbxe/StaOrk1oApkVenhMX4Wm5z6S4Ygbjkt5WV8/4zlX5k
lrHzlVvgiLoDzuYuUuyrCuSIbPe2jRukb6sgJne9nbkUKozI9XwUUU1IaPNE9NVQ/RUIvGQKeetN
fXGFkzr6nfs9YyV1q7RcO5Kx6ZhDAUnflGj8jd0jOnLdLyQB/QB9ha53Ts/8JH13xWJLnlvrPF+8
x7gVf2IJ8V8TqpacJ63XCx3MIa9QTXcnPtlbduSNxwpKOJYn51fktEM02LwQWd1z2kTGD3byb7ua
iE4zL0gAOXduQkyAhRAaPQIXCpDu1fDBu+7NSxHG1/lnVrmNY0j+EyiA2XdTy7sVqylID1QOTlFk
mH9f5TnGwGmO3fqC6YUfbI9g1/1vtJ62GRzBp6EeyID3hUscp4Jek7j+5wYpvo60H06WhG+9T59V
+sNs4MFZqF6uvo024dwvax2vGrRqHJRAI90b+sqlnd2QAeO0s/bVdiV31ccNtiWdomwAvJID6Gda
9UB5Bkvqbo8FujPWQr2juqRX6gzPlp8LK+O5qdnPP+jbBEj4P+rknv4NSNM7i2EqStDwueo2I4Yq
rpnqoDnbk2NPgw1Fx9JUFD1V9rUcn10roTUCxsz9A6ktMvk15+tnAB1PJPCgiawyiNP1J7tDZyPa
vdj9CTep/eS9msVGTizLi8X1JBvUz22tKH5SS7KAitv5YZ1OtDTmGw6FGFPjVxATQ9f0I9spWhrD
61jkH59pl9+cW8z88odboOwJpK4k67NqW9Vcj85I2BtkUfC+lYmgi6VAJsplj1v6M8f4Pkaco4Bj
BH1Qki0lc2upYqNpBoi8YSKcFfm7Y2sJjNbh09/AXPVmsEl+qowNb1Lz8eP410WfZOoaQ21N5C5R
5MSOrLyJRP6M/zPIp3dQycXvbOwsy5QVCXDNt1NFkU0R39Q46Fh0D2p3QAV8zgBXqMQ1LMhiXNYH
dUsCUt2ahC6HbdUdjAYTLg3hjNKrSVl8ggY/V55QIRGmPleZGvlSCaFKF/34gnPNxzmOFhzWl6Kd
VSPPbrF/f2IurdtJ9UZvqEfuYkPREy710ZWPtHCv+KUaaKr7r8R4nrzO5pkx6NMmVMB4A5gikNEV
p/ssOF3lKqgwvZm/GlSrPbOP7KsxsNH9W7IISJzZi2Rv2Rnh8bBMn1QKdHDu4ITUJU8XfOkfWU5K
0+I9JsGVsLIDeHgG9RMcdiN7fylCDNG0NsLm19nrOxJfqPLUJDE1gDCuWxkycqbfv84jhWciincR
neBOfHKNXjSV003S+1h+qSm5QmuHbJkYzJB7hlIicSIBYizMIqSix81AzEiJf4z+4ucv1H4SWqtg
AZFIqidKTUeIj/1lo/ZjAakghrO/XwfSnhcxB8D6JDoBFbClI8NeNgHGIkSmP7YT5IFeyeEICrKw
s0+sl7oEkDFprGxw4AXvvfFkXNrcVg7vX9Hx3af3VW/X0/6cZGKmUjIUhBhqxka0JORm/XuMdFvM
3jESEGSScYcmKoZ8P8tM0F0Yv0OThx6WsoMbWlfkFFc0iFGf0op4suNn1TVCAdV9fVso+H7aXcFC
VaWx/NPWwe8voEaKMojDyAa0mJP2LkDIpFGCKYUImuMkKno7+17N15PWo++pqC8APoRUFDtJha8n
Q8Nl9KgjaSF+nSHHZQQo4H/BZycDc8qVGH5NizofHmB5KNLBwU0gSv9myL1eeQfrUxjoTM7fES+O
23JBGvKH0MvfUH17XDZGDk+7j8E0rggXm8YW/hb6KPoJXlZIM+dITZ3fiUbTPULpw+T/ZiN4eTMH
SiPLqyzsuY80F6QVSzNNhMPq/XCRuWkHQ77+ia0vGh2ku3KAsnKvb7O0azGcqL26VFUE3zHnBT+z
isgYv9kXq0mv3rsa4PHq7va/xys7opjuc2c4NbvBwzpZAPSJ3QcuGSC07zNx5cRYk+y4nvz6cUs8
xdtaSVpQCeqhlo1fHRp4iwI09LloZr8VGhF5D9bZUXuCcV6HTzgrrb1RML4YUk6FA1dKrkd16jXZ
NsZxxK4qJ+OZYMnRIWHEUW/vpybQqehSH9vY2Wvigvr8den6wOl6kEwvJcKw2uLARftjnkLFbUFD
Jxr5ouEn+dCYYKNugM5kqar2VS81xMXBpW+JEWrPBisqQW6bsrrGa6Vm33S0HEgeS2u/EYc4LfCt
cwmfSwzUhSghX4Vt6TqdjnsS/tzd/PcZjD/Bx+L5A8gkbbwtwLDAFRXrkg433xJcEPBMl608enM3
a36vI+AMmQUHXfOhrjVaNL+fwizyPCXJXP1GFB4LighkXwMGniNfB0fCbade6aDO966tcqqt//Ej
a4UsWtBZb51kK/vXAnRPGx5qhUHQFOSy5QUtpg/+Yf1sSn4hsw8vGyypd7rnmj0Xd8tFFfIc82Bk
9gxx3XKHFgj4fnSi6NSCnzJdlh4VWBC6gKmTF0t5VcP7wRbNa+olqJSMRonqjXLvtog+sMyXWUJn
5J4fR9Fv+eMOuB8ys3THqCa8X1XM1I9l08j8Hd75/6tndFJbS60wM69Ft2aJdInuvtJS2IlKZoKF
RsZAd+so54tXiXs297cHDhpVTKwzrC2F3+1z0Uj5SImTbQ1hMdQQtNfwgclCeljalFGRs0BhSADa
SQf3IyeJz1cQKpIckWOJiP76FZ/TVLAyf5r8z/sdl3wBLqdf/2LMF4Mknz0jpSdqT1LiJX1RHqae
obbpIj2oqD5kIvKekochR5ZKlFTANRNHg8ZBcOTqXjweBLpI1MVk1X6sfmnHG8nLYPxEphj12oYE
s5n1Ai7cmZM3DR35LSQ6ZWLWYGZms3g2RiREIc/qYqLKgCaEv/z0SvoDlhS0E3OMkhgd+lHJr3CM
EizywaV3vsB8AxQwKj5sG5OO+w7Re9trkaFpylTARUVj5FqVX9iEP2iJn05RMWdi+gxtukHx9uni
+GoUdfcnxOleVirdcKSO9FkAdrk77zvmYCERi9DCLhEyFqDEfEcaNrQEtr17PBCudWe7+VphBqV9
fiyq0OngpBhj28HSuYcC8euFJt/tTAefV1asMT7CZGXtlxkxGw6S1ZDYpgZoAa1Q1hz0Qz4IPskk
TJFyfwXnQz0vAJCfNvZbaiqCFiCsibmP2+c9tq5tClhbz4q57r35UDDRyCtYxSEb7wzsECEKi1Gn
+xZwfSIM1Kfy0Xi7hHBZb4hpsRQI4eHkCbm3xJS5Wc4g8AFszdnjh1YliTUcxufkA0PG7M2oGziU
eI3amHaJlJcKHtxtlVzD4afHNflKdArI4bX4VE0T01lniaMsq7plDAUfBNYtFqBhlkftNE8ECF6U
Qr84+L7sKvKVvuZTWelO1sAf8uK9Nul2gUbL2+xqZQF6Ddpyyps5OdiS9TJ+kTxpmwPn41P/J8CZ
+k+YACbeJ2HfjTuUg1rmbdahlktvwVzZfeCVkz+bNUQM7ycY54ModSaXyb7wx4GoXBajhyIxqLXy
fOhRl6O3Yzn7lU5dvSAMmG6gTwItYeW+F9rfzrUEM+Lo+vi4iIYfCIXBVWGiSw9CuTHRCOnzKdFx
jgJ2BKXXdp33NJDfQitIuwnlxZksSMLbqpWrLDdq3ukxLNOFjxoMLHRdxhx00P3GCe9eUDdD1p7/
EVoDg9XmMhNMtzlgeak8s3/2/wOdG3ZwG3sOufst0ZFoir33S6bdhWTIk7vmqi1k7K42SC0scASF
PL1qMsxnKIXohR6zY9OiOWncbafNiXdIlOeTtBR+ZdlipIMC5H5mdLrwbUT5WSGvyAVxdx1G2lJt
3Wso0Y4TSA70karQek48KpKK86i+rFQchso8Gc2+w6haJG3oZJQELZJyK0Kbf+gJAUN7dOjaCZje
sjSgO3DWYgCcvnJhfEx0jCwK9bFUzl4GuyL+K41ooF4q3l65DGbDTEQTS3Wn1cnv+uu/eWsdl0zN
sy98jGgRna+Ky4ZuHU/5K6GTEhJOE01JJVOV3IOs+cHRDZYgTx0qV+SJ72szp0FmMI7nzEaT3i1H
CAr0XAb8oij9ibDLozivQ379UE0DA2axcuzsogCSqKcbfJghpwZ1VrrN4FAx9h1Vu7GZGr7ZpLMn
qAmKSs4FMCP6vdj0BEoKdYIDOIGMbEhMZE2H4d5Lsq09TXMiDztCU+ZDRVnVmxXOcaWQuKQ3HuSc
mjMxxcUbQefGBOIl5ihynuBh//T3eF5p5c93I4c20FtZiERxNEpcTx5OKELnOj34W8EyLt1OvkOh
HJAi/XumuUiGTl0q4Z/Wph+lAr+MtG8yaMx+E02EwzeXFxajCzE15aRHLUEuW2Wv5o2KykXBNXHq
CTkjaQMN1rLnev4SMny18r4TSmKg6iJxX+XKAm40XA92rTFr68bTPxUE84ZUPfW9uFuLqcWYzBKA
/xfrIXNZa/lSVc3RQdgHLh8sExWBg6nPxllBeH8lAp8S+R06hMnHUkEq5WfyWCVyZkdRsWvU9UvI
RhcN8R/UwjL5yY9pDP2egnRTC1PONk9VzjsusrhkFta8MLHUcHN9SRcaz3gG4jmkoQ16fFzEByrU
8/OggTLyl4sqZQ2YVM9beisbw30x9Alvu7hczk/bRb5/2zisovS42nZyEvsEXn/4UDuy8ObR8aeP
IS4LqxaeH4/e5cv0JN5/kRBkeVvnJ7febvO6AXjsCFej2bXnfj9yNQG1oXwx7eQ8HIoj2W19fODH
RHKY+rscgiVTDoQUN56T8jhvCwrsyoS/uPCAZjZQBSPgSnutqNRp2TsnPgbv0PGIM3LFc5bJHyRO
c2JCE4IgwjNffX5vUHf68SiveNCm1Y4vB9FzaGROTsFVHp7ac0H4QtQ711/PrPURyaRJjqxsJEU6
IqxgQMXHom6Bz5oyWJJCYuuCZOkl6ZqUumofwURE5iaoC5JRKFnZtjJ5Y3+lPZKDPElLTb0iIF0i
56xTMqgC5Y8WCwjqrYk28NkPKr8T5LCf1XHI28VmweJCvIMBI7wdETQyADgxH07WioDkTzc5aQa8
fjBTvgCbRGx2nyURpRtZP1kPbuZelGe+aYtxGpwyYK4CHJI7v52DkOktTJCKUYHki06hMQnf6D4x
Jbkiv1D1s9pzqzGl2kwJ1TxR8MiQ9IE4Ic+AAW1cayLBm0b+p8VSZrCTpmJQ76N3bGSg3dRqM9BD
b+v+E/DLUbJIZ+J+4qVa+pr7/k8tnhInHwO5Nn9rBWf0PoYXNv6EjL7bE3f5OUB8JCOzyWlmaE0N
uWy+ZlNzGN/bTLcBbZXVhq/LyCr4adS3Fy1+I8K6lIPu0WHa1L/lLlhr3EMvtYFrhnpnbAHufj44
UcaRmt6NDy6lhAMBjsoiFc120eIIwZZnhP6x7MpVsZusBlRTN2smQRaAAD8XO8TBo1oOfJjYGY+M
0cGxLEu9nekbyGV7UvS57upO+nuTzXCxMhIkmoLvBkHGixqqbJUrdLP1z5Nf9SNDLimefIKn7eI2
cPmTqsyK2UvXV6Iys5AevQkhmrQXFSQ/96bjSqp3R1BUBkwMaKsheeKtSDamDv1to0rOm0CJ97ZS
8bjzfTyHpkr/ULIs0mgAJijjkgIEGphP4/1luOhQO3Z4s0daKs0/ePOd+0s2EcglUptsBs7skZPP
2f3IjJ725N00lB1eUlRScQtKcLCjsn7f4DVAkgIdPpXAoTJSLLy+xFGhz/YWQnOpBQkSCYmKNSEm
eck/N/Bo+7VrKKAu+6mIkr1tISzsIfsfTTsHc9hGFWc6qUzVAS/sWkiKcOcwIJQM+5DGu+xA+Nhy
GUpXRfxAmQeV9m2xXwAuiQsAlBpMc7x5knH6Rx8wQYIwxuJspum+QeGlnYmqQYDTafE3i9o+WNgk
84xiGlfbrW5y88BXLTT61maXy6G4tlaXvn/cDEW7FnOuVBpY+YRIJ7nGESPKf7cUb8htPzOFdcxQ
t8pAlh+4QycQz0hNcfLT9cxtElPEU0IsPN16i7cGoa+jWWY0YvBeBDD3Uy+TkkS9BkBNFhuU78hL
eHWZNp3OMuDqSmAQ9NOO+n98V0rqt46Lu4nR6WZNoZ0v/z7HEPPQZ+3Yn1LJcx7U2qWWtEoesoSb
rB6LZ2u7YADY8/vbIHE/NhAurbkq0OLAhK+rYBgRinx3uFbIfs8Zx0hvr8AkiPvjso2wK8WqC+aQ
UrUjNDHFji2fBbPyubQIUlLsImj/i9HZJj51q1bLpGCi8onB6MLL8AYeK4++JqjHZ5jFCqOSixmu
FmqPSuNV1Juf513P2xc50WkjABT6j827kz3iLR7vkV34Tg02HaTDyvO4KFAOlQYpEEGPXgiCSavy
8q3HwOpv0SiU+z9RUUJb30OWAs5aatE8YcwIUHI1WhQ7H1c3PbqTzIo8rir43qUUzKibqm4cEGL+
dJ3Yem+L1KClwvaXNWXeiwIGLS3VgTzXAps+3qRJYP/HTKWmTKTsr7jktHaMxwkXm/9ERYU5Ssvo
TargLy+kdfWKdXXfuYfa+xtEj5/FdzgaBTR/48B8v5ojpM+IxJVZTpxYZWYcG0z9lzpXhM21exnX
T3q05lOu0Ch2JxksR14NDLQFSKLs7e74D7zc8R3hKJAyUr2Ew498EoPMLJrzZ8jkL9wZCwvKgYlQ
aM2ZRqGskTz1SuIejgTT6lkX9mYHFK8KlwlnfjAQ4gzSzJsk1f8aoADx2KOjcBQrV7+boEqPht+7
b1kyz+L19/p2JfLCAoh6dYLoJDG8tMcrboMmtutgCKz8ttl3/Xr6nA3I+bwhGhJz5eyLIqyHjF9n
nbkoaVbt9iuegMheX3r5rQ61A8XrztW4dQ0m7HUNP+nd766ROXT5gSGWD8bAj6UkFk8DsjupaOOI
AoPSb293Fe11BPDKsNhHrcvmvyw1JTIPfy3v9+rI61OAX3zxaK45KJygbqD5x+JFnElNuUiuN4sQ
eBiTFsK5J4cEP+STvIAwL+7EZk4E8J39WKgAl3EDwMy5F1RULwmKu6hxK9qWOHkq8H3l+p/mpZpO
SHTgP1/O7qSCsgrFxlRr3Dh1xBSVLS6S6GPhZszeKwxPOq+riWKBgcadzQFgGXwuVPCgk74xFAFE
TdeE8PB4gczN4EdtkX9e18z6s87ComXmY2aP7wS/3kFRwTWTTYl+Cn7SQGFT+tWVjssVWFVydRoj
7vX8wwrbVIxdnnowR7yXcXAnPzoxFT13C7RjN1PT6GATeAIEd2rpfAHNspvDQTjYYRBbwvBnBqSC
PpTt1OG1FEXDMblMaHySvDfCTU3jDvMnvdaJvAsFzoniPAfre3esOZzJPIuFMkMjbGWJsn3PvNI/
LdRij3POCiXJHBkO9W5Dsp32Wd3bntXPho4PHBScxlEzIvXPGn3xsNBQORAvKgDeKrTIHX0+7QpG
nq9+kE9ozF1oP6gqXPi0IiFVpB9yNdb0DAvaLpfjXufM/llqjsVEvCFOw/IFtjQI+Dfhm+BrHrHk
5u1/eEY+wciS2Qp9IKWppLv9kNoxSaXv3/sSr1G1fKXy7Janx1ICEuJQcOKB8syT7MrBQkDVL7Br
vbRlbW5Hq3gPFGCdJZzKJmJ4sWvOp9BgHhtN7PL/vbTo5Ll6jrXl+WRKfQ+6t1F5ry9BVkaF+llc
w0yJCqr4XQR9OeEXHMsu/awhUwC+DvuzFy6YuV/fz47rPEjiOz5VqRgVc1HuEvV0fN67yj6HKJRe
96vYElXssn9bwu6yQ3g3iYa32xvRazYuHmXEliTN/BPokYsBFdjUQz9zyXB0OQaLVIxezOgPYPxQ
+wM9KJB4kVaQIaOvi6sdbFcxP/jONa8KALU/NYfSEEUSMfNKSpk7QAh+s2evM9GMTBHxOSYef5U1
2HBBM3heBKukrNcyKUaMh3HnU1KLevdAodZ9fHuabK+m04x7jlE1hBCjPvhEIs7e7WQOWTkFv5+k
+MGCVnvjwucKXWsKd3GOmOcpQgyU5kwNGzGRTWtfVXL9wn1lE0F7MjgKJBNenCR5mb+9sNfdkWFI
TJj1ZQuSwLZkn+Bw8wyxiRkgUd3ibAh9+elEFv6BpDbw0IVGT/U1DNySn87/X+1yUJWr6dJCwfKi
CiqjoqyZHh5/EIBqK9msIUVkaDbmW612fKnRH/LhAbDP23av+YNFQoWy3PQj97v58NB9CbWEUxu/
6xO9mubMG4wGveLDHixcw+Hj/ZXbAYuMzVURTTq0at84z8aP/yEIDUXSJo02YMcQtuwghkZ+0Xdk
fFHEtE7zUBPD3aYJOLNBflJQVvahGi/k3KTayebBHVxI+vYHbrM3xJ4HdZ2c4Mt8FHndq16n3AS/
Fn5Y//HFV+qmjFRcPoRYdP+/J6GCukPutRm1W/hryufc/p5g4j0RCNHwFWb1hu4ZpLdWMpmxhwnd
HhnWjulervYm5OAhg4bWvFTC7mtIuwqa77T3Mhmo2sijvfOsyhQ8t+jBPP3SvSmxFQU8TDzMGbWA
5drnHdwYBBr31ulSKX7VQw7P6e/kbsz50yTyTKR4PwniyMqabYO3weIDCoG52KXv8PekKeVnqt6V
SdYxc8U3iMM9CrNqADQUgYgwcB4A58Qw6mlz3GRUrL0kPwvZAHGR8kXCx9IAxr0YJi3ZDXi5G6kJ
agm6VCh7IhtdjoqOPVm80xJUYFu0BxUWhSswUlPPysVyNlk8rOtlLYhYOQEnE5oMcN9KpSQsHDYM
qKqagSleVikKK6g2vN2tlPJVhqIday+MTV1dEF4zEoFEeEZdbbyUMH0DENTPt250wV2Q5Unt357D
R7Azmc1n4LWHQwKbTqkEX318JTqRvhsMokxXNAcX+3Ta9Dq0VVC8pvBwarkQpfONJmRt+IxlqdcH
k8XcDrLuQU5HOCrsN9o463QGAxyPiD4aSuNO+RUyG7CYgQd2NvOsB0p7ZkIdJ6a4WAIMLnWJ1U7y
qBU+Ll9njZXt+pC4QkMc66GsDH5rkvcw4lFAlEpP6DnASyHc6/KF2DQjLPNucK5294CfQIl+zPUo
F18IK9XUtsjGfX4XJyjUNr8MWSxdSfbVXDVi+oLP4iEAQU4w3vNg8cFsf2L1s0pZr4ureXP/0/Hw
W9EeMN/hhlRV407jLhv46XNM8VPmq0ixsmrnVdna0FOxavdYOFnb00ORBdc5KSzoFoPmj1E2REA9
9fgcA0O7og2yjgxtj4ULoNNrJqVWQ8Q150pq0lXwMpD0+5P1U9SgGhcQ+eSXoXYKuiIkSULPSclh
Dk2qiykD6CTwpGtj4K9k4gYCySntUQypQgitFwFbDAZ45Z7nipM44tGT8Pfv4Ea+FGfRxwzkjML8
SBf5+7SUUSRAeRWt9P+npNCfzOtUm/FCU/NE9XAyDLp8MXHXXbFoVPljFibjmNnRLyzhh3slYTOg
VWIEU5WXWlmInS13rxrWc9lTnJrbxWqb040AiNcoAKkJEOaeRzWOuMlQ+mLrvCy8nIb4DAiIrRTW
4DD27UnO1y/n4BVpoIIdLeUafxyovvGjylkZr+W1fpLtSivNBai7LqhTgnudul1psYuz5bLcZdWw
pj22juFJ5yH0ywDj0rO3oMvCaKNjBBnHv17AIfBVypOficerSqFySxqEeLdqvvITe1n9DGNiZaWR
myLuuMqiSd2HixHfEFmyd2Kh9sTxQDJveCtjI5y44pXHB1dsL3XNvL3aaZwV28TLAu7bIsGZQ3vU
m8dJuTfZ2HiG0LttqSzYqXC1jt7tL1HVt6VWQVocFVig/QOL97TESjaAJdXfLsHAQ3dIAhXP8u+1
gEyxsT8NNk8oSJQ1+Swf3vTT0BZDij8x/2MuR+O4Vge9oOkoTiHuzjx64htFHWvGC5CBgocdICqy
QrIZ0Sr/SUq6L5pV3WY3DdxaR7hxKBfZRV1+tB3oy2n93Qmf/2DPR7rh6aNJLF5O8V7rykAsXsB6
VOBrH5/6LArrd91sWdxrkqcmIC61jiLwcEHsGi/2EdClH6+JiXwrreywsL/plLeT+5SGsbmzEQsz
b8/1/lcpIxa5qxyG4T8Yz6iak7bR3+79hxTT/OtXxAiKma7VKX2fEOmfFU6sBcg4fhOUGoZ86LW+
s0G/vzrwiaT4jeUdimh9KQ0g9IJn2tX0pbMLTbs6WGHL+1prV8HGwcSAjcQHXY56Kw/q5rVKjKbe
gV9p0wKuMGg0zC4oUjmmSM8mm2JRNrY39LZWRAr28Z1D9yzSp2oqPxvEZyl96KDwmNGiPjqw38EA
aaqbcfSQUxR9+EMXuax42srooKoazQitCotpJia4JtMtHOfjFdnKbWktQS2yGBjeaZjRLmTv7WrE
CwntPc8FjDZXlZ0YVwz611JMNahdIToHebeiGLmp4N1zxCxvWOiuhvTbZ2Cin9ynNdwNWVvRcA28
JUxoaJ6dwFR2BqFHoscmGBVG+FmLQLjVOas6Z5OSoU7z5VP+/EGfJIEwkBfljbdTxudqN5eEkeiI
okOtX/3J9lhCOxbwriCvOO5rpWOYOVQzrp5+4dnQIMFxO/pAtnv3y+hj4n4YuPjQBvml1WEOeULw
PV8Kn0G0RBs3zZT5bCkq21S3wsQ19V2FDveL7Ve8btn97vxPYEWC7xSs9zKzIjM51ekbWBg/LOSd
nWUqxt8BeD8jDUHaPoE2hsRx9pR5jVrOikRVU04i84TrM/ahQpax92eb/HNNUrUh0LO3CPSNUhcv
57UeUfZCGGjr6E5fXaaz+qlPKxl9G6Cge5XIzRx+9ThRSJ/2HqQBGxcysFGgqlW+kWDPtH+SRHZh
oQzOrWM4t8OYeYtEPqTvNIM6t2Cd/Q5FWfEwu1oidTTqnKVDONglS2IBkuFzC08iSJ7Hn5UU0Bwe
ocTW1Lfa3I6WY/miILmk6XtbF1PxfxHWrjQ0N26C/ux0say8nY62o6z2Ic6uONjS7F9dz6/HxDu6
lfcnJI990NDp9N5EefhNDJqLfI6ZpxGEVNyGIoYsaw6ipTUvbt4KPilhu9yeI9pPfQ7HiF2BQy+C
Y+cd31OoA4WGc3hpLHxA85EL8eDZc2Ii4oO2ZzsTlwoTSOzbTAgkK3Es8ivgLM4YQS0y6oojQHnR
DR/Es7Eba/DcqYSqlkaCjK7G9M/sKKvD6Ndyd+vnhViX0Fr52hpJqIeKULB2z/1kQvToPz1SGNar
mzk8g5wtnxLwkkm4fIESNOsR6ri5UhRUWuXnPvFbmYGnDswAjghPffrpT0MazvD2aKew0JUbU0Ez
ZZkuFxIHX8im+iCy6cDVJtLuCVy9aHIu7k0g5VSpVwVQA41yPmOT1cV5uNjB0RVXKgUFOfOh0bFQ
+FQ74GypzBOYEA++BxsbwzAiWcemqR2jxyWdgmFg8u5K9w7QylwqFsVyGiZ0h82pGWSQbpM7u5Hc
Gvfy1je9R96dA7mZiDz8gW3DBSPGXHK8XLQf7IMXG6PWlw4hYDqlsgbX96Omg4vwBSuRlKrxmIkD
gTUXjArr9D+nNOLOauZSXZT+Tqdl7J4BqkVfOEMEWiG/mNaUc5vyW/DqffHsKBq/LJXsR/IKW27J
k2FQWF89bGQzUm0kAm4++2Gv2Ooi0bW83m0pBy4panfBq1nBKpKt++syCnweLnd7gsD/H24350wi
ZTzGbx9Z0BmB/MYjvzKvkoJVF+m2+tdj4IBW1KaygRKlfw3go9WUL72o9S9mMtBg68IhlwlDXRGX
IYYixVtbfCb8wWX6gEobKwlR8tlpULCqxoFjKcHDPfcKJs1B0eejEXzOJpEJnTb+7hxqshxekc3h
NeW+vFdCZaNDS67esySt6KlV1tMbc4CmwST5ZopQJ2KtLkSmUCcRqDKIMaXOUm2jJm4g6uSxgPGn
Ie+PWXW22BWzx0fts2MfCY6H6xYa3rTiStiwsmOeNDbvWz8su4Yjr3hTlzWMgB5fXEF5N0TLWV+Z
2OeQ8JkbTTTocmtyRiMb5WxH/3TQY5rdOzu0r+M7C+NucZjAkgAilTGMdxJjAxmPeJmpg61l3I55
Mla+mCM2Vxpfx93EUX9OR1OvWUq/u4GSWQgVLzTXY5ZZkFqHC14YdhiR/HcFOOKVOiQi7HWjTTvH
MvBpxU2I6b1YQtrx3CxkPE6UKQqii/FzSgUoajgSNqF4qTvfkzDJAM7dbQncZAaWwCVNeYLPstH2
g+somSLi6hLBiVw01y7LkX4+D2ZQ9eSQtSkmgvyJdzFoHsIm/yd9aRFca9L2M0tFcesjdXXauSaa
QC1qYU+kd6oiksLP0zY/LmQl9DvheBPpB36PfR1xii78P+qpp7491UBhSwy7Bv8m3qhMAkvwYnAU
+nOYOJreKJl2KPUJv2YQOZ3/HOAVXTz9NTVDuWbC1RBd2Wt7nIH/DCY/mooc6wH/lrR8ewoNcpKA
UdnoQCeWKG8Fd4ZJEBks95lFSJQxE6kvvvbx3BY2XRXUNl9Bjqvfm36TZOlSXXjb0i7t7a/UEsDX
GywZznRGGftufpe3nbJyHcsOvaYTa2RRHv/u0zFMujpUMYKC02esH1XcOLJFb33WqprR31u8xlgj
VllZuno3fTvrLH8T50rVdQ0nxQxJt5utyZBzyQvMIzIAgedULA78xkEByIu50FNkMqzChlI2JfTZ
HtKGn1jtR1bnZV/Yw4XkfnbNp3fSOM1lX3fJ5wwxOQm4q8k2TmBjGBA4n9mKR5x3kenAnNNFocq2
mkM3BqVkTRHqzyYv6QAo57XENUDeImoF8jKjrDPywu/ysstC5JA2cUuq/THqV+G/LHa+r/o5e/VQ
t01XOt6RThjoZJnH+PP3MWB3CbK9Bk/Vz9Kq0cEIHdOhreg89s0UsE7SipfWq2KMRS+gLibXdcea
JZduUnv/FKuCzG+ayP5OWnFd/aXShHM6J1glTKlWi5JOgjYGuJ+MHL0W+uxkFjFxUeabmUxFCIHv
g5m2i5KyM7Oznhrk+qwOhzGxXapOfqSVDVx0/DMhMsT/u+zb45ABhQJnA9eRSF3gzR5coseRdVKM
ex+zrmKiXPJzqc/AF0OwK7g6xB284MsRHYCHgPoy3FFUpioyWOo1H2CSRbBAd5BZGpEeUb20Gpxv
GaV94O6x7YM1CP/OfHKoS/vPCeWtA24ARmSmEDMAszJFGp47Wjjs6RU4i3AYMhm0Yuqi7qvlyUES
6svL6KJ7eCN2uWY5paQfIjpmjYh51eC+LlkScf9p3EKfsHm0OmLFa4ccvF1FzYIN0BBdq+ZgiUNc
s7JKg3W632dspbwO7awTipwewt2BKVYv1xecsNi+xtEaXWK7rXQHxJi8mjjSWhvrB/ATXhObwUfp
VkthumaTK5MjA/3yrgJ7KJ1BEO6A8JxbR6v95UTs0v0fUx8cuJU8pTycz1qUZMX6twwVz6ka1n/t
wX59yDk++jEh8DAcKvxFXAUJDD404/95U/4E6goNao1dwy/m5NkgElZpQxORtXIiS5cBArXH6I9P
JCxeZjGnsDkyaPvmI3YEjKoi+veSrA3P/GRA2k9gfzh86lAo+bw9gdFaLPksug0xCejZtQ7MZKZT
cpu/9J9EVdh1tProCynLwhPx9TBu0dtiLxgubEwgGptwfqSY6FTSMNJRFAN+HRg+1eHoTjqqpe+n
pSY9obh5k/oIyWbwqhEiRo2ybQ9LR+D2vH26lp6i50+WJw99NSAVMu1n5beRw2D4o1f72nuIhiET
RhrBOJgXeI+R2ZMb1XUOEFXRHd/W94tqGBqiylg2b2IBlmZMgLl6AUTA50/IIrbmyAVI/lvgMs3s
0yUM4x9J7oPsf8ksoTM1e2F6VCxDJMv2VmLcOqNIO4MtSrKZM0IReMbJBwRCUenP/38OECNIhRB/
alIWy2T/2oN6Vp00xbN+Rp5pbXV2JNqKkqYCqD8yTUDis1Pf9re7og/vEYdNOpAGcAJb8lqe/EeL
TfYRasvq+sST/QLqli2fbRYDcmsQVMMBGVA8dbcvkyX2fVKzfDku5mTX1IqbdgN5IFBfZE3NXz0L
snutexqQ5ogPekvvlMWM1Lz4M8j/vhpx1fuF2TRE63ZW+kSLl7/N9dtUGjLRZ0+9OQxepr4ANG94
OiFAIswBWGTZaKI8PhAQ31LG34XIvdoCBkW9atVSpsy2jKk+IE0Y+bnANwdYO7z02gGjMSnC5Qlr
6ej7pC0uUrzE8ZXRl0jPWbzIV1mftxMrJBbkdFx8oAD272ywbRM4BDPhcQ4hhv9vgG529ZYo29H3
ZU+f61YSdrzW93V0j0STMCTscglwA/flx82H6c7vTrOpXGkx4yJNd6c+YX63uJpf3VRGEjZetUxv
V9W+WPW2wqcM3s9u4S09f+ZDQxmLmb1StLhVwIo7pjQm4o5K/DNArbOx/xC0V15FwVZEaU4PBUqr
iAVLVCruKy0B2bGMa+qfvjXy0yMm+iI3ar7FAL/1vhTfYt3bYgHH8lRHj89s/eeFMXcthqGzPBfG
M7bmBAtReJ6m3c1nK0RmL4AKWxjoJOt88W3Uo5fB7FqUQrtqZIW1ifmWMUQvyza4StIDdVbyc6ib
1swqPryH7CNyh8jY68jv8WDbu75umdfmcJekPZtnE8TGQyj7jw+md0FUxLcmGNF45fruaudu7B9b
/vtCIaK7X1WksM5lvLQgOziEZjUZaY3sx+mGR2fs5RukcoAc51dBR980rdX9ixPtilN3VQhj1u9Z
85ul5ZaRTKkN22L0asZRh9wHViLQi5XtlfM1SuTXiG1DMPYxMJx4Rr6JlEKiR4kwBxS7bn/U2R4a
MuSlQwKmhvMiLfSqUGfykdFsEbJ+zB5XU4UB6Gf4Vhr4bCF+wBLqax6aQ6orNgAPW2jpQ7msVk0B
QmPGGLPnmxSZZScbyHL9OkxWwmfr8EvbcHUf5ntHbzhDVwUuOG/eVvRLSsKG1B6E9UlBe/z9W44t
pk7/gJ5j2XuEVtnu5ILfXmCntlzz65LKR2h6x1tpnCA/sZWrdtZBIWLlKqVpnA7wLkxh3lmeSarQ
hUubmeymw6ny6psmsYA2xSyPLXVBihFdHukz+PZgRxoHQkpnbDUWIWlSMD4nImG+4POUNw/HrCaj
7TFHAyrHsImrI8ZH6rAbenkDScNQlsaU1IKWXkNSbWhToCwnhh5jVdZGgTzqBfii0etnFb+oC7KX
1PQztYDWkr+rgOytx/pAnRLqTAhxZX4SsYjY9wAY5EU6vL7hJp0O0TH5UgWA4kEBGbE6lyU6/++B
oD8L3ifZd9jr4UmcuqykJgZ1VCb7bk/BO0D1twTfzoasgEmKenSye0osXas14wSPdk7a9nEldeWF
lLonWPMIuvupiX+Fp8XIBLMZfxGwkRQpHH6mitLveukllsl9L4ZSbDPXrU0Cr9pUn6BwAffyDsd9
3hWiRd+wTdHzU7kpdHbPXLCynqAKhx2FK/IWhXh+IVeOMeDjYC86ZKHdM2Zq0Z0EwFGTh/RBMX1f
EqLs41PJ/tcBenb4+TW3GB8nKUcGMJL74liVfPI8gnHEbXpWh/5+CoX+CZ+DEFD5f0/+A/8tX05r
NvxMmI7G3ApU/ZqYh7rU+zs20tLrgjGwqT5RSbvvnr5I98Tp524K6WY/zBRsg3zJBOducYDAy4Mf
AOzb+DHsjDdCihSoXddDwKpxeTyZJK6bps8fNFwIY2XqDz0PwW3d0OxF3Vw/4yltxMAUPo2SNHC7
4Yk6ohrQhk1AM+8RY45+Bt9f8Zr0axXBIN+ekcz4rfwCr91GfPoU/f9tg0W8OPp9zq+8sSozs9yb
rnarNHjNIcUVKyw+82OJTfcSluoCZIIYWM4xcADKtOcj4Lw21n/KgXvrMFUO8gNkFzZYxC9sa0vf
UhFX473E8YIvN+YixlOeK5wR9R//YB2GGCyUA6Wmj7R+IzXjZe5R4TJPY/49/77/Ft5EuhZeottK
tNcD1L7vUkbmkUaMevM8TmUjDM7K2kGXbQxSi3e8jCowOM56L5c+lPIv2nDf2sVK8/QruXgM47vU
zkirEUJnWAx+OcCp29JEYP0i07RCiNiB+0q4eF7Uh+MJIhMV6vqMCtSn54KbWR6maDH+Xy5nomcl
DIWRyTB2cCbgCMrObA+6izXikMX3J/jBy6QNQWv7IlF7u/CrMWbbT1u2N5YSPTbA39pwYhLJmYim
3uB4SENJOP+Jm3k/TDGaFdhOK5Y5zkEPOiYH/My2ga2hLcZj/qWSHhBXsBBIKNfwwVvOttlchLKq
+1tQPSY/wN/Nu8OqZtuCbHKLcQlXXVfJT1hQNJRigvdBsMhMEAoy7U3zXLXhhZXsCZHmCkihadhz
T3MRBPU9kZ8IlVC7uc+r+jloGpp+zbNO9Ya58X29XiuiUi7ozg6xhE19ByxH9OQa9b47q4NqfgAt
+LyTTSL86vJFowqQBYmQwnFMYGfhE4kOUm9cewDzReI6pkNeTK7Tnf3VTzzBzJzIwG/sFUcmGZS8
4SO2WsBjpuFZa743pTkx67BfP6TPBrbTNJeSZX46dS3FoCuLYMIqar+uhVJousboPT49ys5jt7iL
S7C/1wJVPx0D1caXbbH2FN1k7bMqRGJKvib5ghM8g/9CrTWnlf3OolQYBLDrBSKFvLJ5n5YbZ6ue
ntwVQZCjEVSpqw7NTX1WkyXncLDKgQ23RfZAbNzM2/gZ8WKNY4Vb/+qEdtqq5sdghfVh9AUQeY3r
qphs9V7Z+GFTKWEWmTyLLUv126R4RaNbNA8AKs5HeKDgELXTHTMzBgEZDT+Ye4Nu7g8Uo2FbEjLz
vr1SEJUUmqbaEJksWeSkQQtLhsea0zKkTkV6P2RWPgw4B5VrZbC6Y0QHt1nv08cNDo4CzkWAMRqD
lGtOkGvm3lE64BheOTsS+AdmLdWXNCRUPwQq+3LS8IJZuptLuT8xFHBs9zE6l7UTuIyFan///VER
Z5EcyMmM6vKTf4JmsyS5dlBLbsyLVDT0lcs4aKMASq3Iu8vsew4ggubwz/Copy2g/OAJgxyJ1s5u
okPrM7uzqd2g5jCSeXw1eLnklNUohPjTa1kZdy7Hbdhsg6eh+n5pXvEyNT/AJGKc7ST+p0vbIN/d
PVeDuPrq7UeTbAVXwnOaegIWBkP+t6hvZfwTUAMFj+D3+G7QofmDyBYhnufV+KcpLMezS3AbOOb9
J1CLomDa0TT20l4Atn0Qy8UyF3mWUXYF9EW+D+SOEoTJ4yDKpYdxnQY9TtxzGxlBwbBO/FQq0AcB
GOlLO8yU2ruCEWsDZrEcTWmliAwF1B5RI6ug965Co5rTGmpXVKtWqrnAf0qUim7tKT7J+PGINxG0
2K3yxsSsJGzqX1HgxUMCGB2gGsTeo2i4d/WBCH2ZyTGEdZ5kWq4N3tV8vPuwWd1uze37W7h79nGf
mYMLbqdIO7PtA9Llm9FzaUgfA6pIMHLPr17fbBIcBn0LOImuZSbvSymo3pMGM2BbntMrjt4b46Zh
VXprRKHe38HO9rO9jecE5QFCLRBh2gN8r1ToXOUCipjmX4IiOHx6cZx3XFgUH8O7DBXj+kUaNXZg
wFa164kpn760QeiIkAO7p36VPen/oCk5A/+YQj2O740otv65lRGIdvEtoT90k8M5iFo4EriNq5qw
vXQap+X/22j2hETzFGa1q0H3aVKxb9KWjyq07p6IDPCaZwmpN3VY52X+LFqzjO1O5JWxVdjHX0CH
/N0MUx+bVpf2qO9d82lKYdhoiHdHHUBnjTSOHfDwGTa5DGUdbQU/8jvIBTxGRdCS598AHwWmZz8v
qj1v7fPnj/7qdVomFq9GCXXJsbL7AgAW3H4wVZKNzjvCrdLfhF/9d5MkU2idrfxoZg45/A+gH3mH
Vev0dSqBPgVm/vZBoIH9tbuPDDzkD0z9qbfADhi4y3V0jAnW/h3wlUgwAPW4jkRDNnrZXWPw6DdH
/EX4blyUbPullPiyV1xhAUfL8iQ1zbGKZvBr7HaG5+c7OqdhHVhvJ27e0uY37ArYR2GFVlhX98Au
wQK1uEo604R6eS7Fk77vGvQAiQH3dHoT3Gxs5+kNxpInp+zHbySTku5mDN6CsOuF3ao21BeejUGo
UUfmvCwJwFmGTfk/UnuL09x+ovyehstC89X6rz6mdmi7dhrGIf8MfEkjlSdhfKVAeZ8fiDZjs2MG
vCLeo90X/g153/I0+lEKPr/1CeUR7BooZD1PxUBe5/oGWnFAuSvdSgN6Yu0K3EwkV4ugCLxJZy5f
YNqLQoqmr/dChUD2tgifSj7YIjUegZglCHqDCj5DZuicQf2TMnopUkF/o03KJabUoqITsl9R1vjs
DXUlkBSpoxGOk4E/N2KUHlIv5CxXMCp80kH2tvcD0kNRwOboq9EkPw1ugb6SY/OPMgdM5BxFIEpV
mbeAmEG1Kcn/i0ZFmgYk/2rWTSTyguOYzUthADPsQ/nOclPIPg0slTnt80kDDC/+WuMkBbRhi3H0
RuI2JjaRdOp3Dr+TM33+Q+yyCw4/EfnlzJ9oxmU4RQJS7110/MeGlKuiMgnlqowoFUL/YmDgRgOc
pJax9YZpNL9D0AOJVhr9TPCSaoUFqsVeAK2e3XFUePTMH72vU9JxzyFf39PCq6XuYiZM2S8rhqJ4
Dr9KTW/CWQfudSIkegB1nZFVklnvzVES1nI1RV0dCdrOep+kXnQTtSna/6RRjOvEmMl8tKTP1Fon
x8Ly5QQPEuGiInAi60x42RgSvmH+hrkdrdjJeMlDbcBq3NsEO/FSKGm4xDSTJBpashiHJE6Xi+mv
ZmqXmQyRp2Xvpa43X9zSeHYxEZOm8FcePnBn1icTe+rkRtrXEEEqNE6nXH6qta7/+Lo/74C6iU+a
neF65tsTeXX+DYQfDHHpB/8uPI0CGG0TdS3LAufsFbJ3Kd5jlgD/qGvqMA+R6WKi5Bw/MkOR0Bcj
zGdKmrkmM+BuwOpPTU5I01RCrTsCsE0h6kkxIR3TIBGxZr61X/f9NinMKg0ZL+xwtDLqL3hqqhap
DGdTXXc6tAtqgyEdM7lgY7/Gw82AVeqE/Iv5uxrzse+6OuZ9Ul2SJpweR7vB06dWVqHzSPfL1clb
lhxymIpFvVmL/mjHo1SQzxnm3j3MCZy5wBxEZuGQY74isEXm9tgwBPVTcbm+e3a0fLhLgdUCen8I
NBhOmW6Lwfj8vYDuZil2Go2nObrNNeYBZoxxwPz3D926jt0By3Pcx8enQbbfpm2nxbEba+IFjlW1
VvbUhQKC2bUmiEhu/nB5eCiD72Y2VvkJz8N6GBRtdYSMit6sEsoCBX3LRJbsaBSk9nRTVlIiu4Eo
ZIGN1uvRtpCJDfpomzfnEr/KE95ZAnV7MADnC0gIIqiGWTza27yuiOO0yLPXQvyhhj56jlYU2Pw0
U8oqIrw0aVKSVtxmifqy4E+miQxJrV75C5/JrO4/cgAwPuMPCPWG8dOMOBYGJryeNYtOiwNrHIK1
cbXQ2uo80AUlzFBTivXy51oiJgyFHn+WGwJg/xW7cImOlyV6rjKy0mqUvLhF2oZlM01RdFWQA1a9
lRhCs/H/k80MPl7sxtwl0NrxQDxR2Y6TfnBOsny4UsMe8K+U13ajRgU3vBfyDm0POblOy3Eor0My
dPgfZgG+4QoWlZ80due8h8QaFLqfz93d5RLFhXAvqt6my9sWlFUB9j1RIsyFgbVGcCEBgbp0NZgl
/2/iOmdKRirRCAoDwD9J0Ei/RR5O13Abdf/wFJxE79GyWP1JIV5ltCSKQV0KBcilSF06e0s8I99o
69hJOw2Qhsn9Xeto2rM7HCPnzxS0hDNZsdFSqs02JwXM6ec8L9eyR9dhVPuw2/lVGfAvv5fv98oG
uN6zfvxU3UPwes4H73tFzkcZk1qe+tlfL00cyRkHToL8s2x983EjHE7btGf8laTf35pqlakh0Khr
bnS4mNwYrc66zpnfcoL0l3zP3NEltUSJ8Gd40/WJN5oPWZ+cB9FHKwUSSd3AmW1Dokc4v1EMVOus
FIZfFxbmPHujPXy64e+fP9J9SPdA6BhBZOzTe+wXYndOzCPkzfsfI5sfzU1Og2hFqmpJcFEZCt3Y
MWGffeSiMuFlixq9P2G+dPlHLig4GqKI+ayeAq2UUqE6bui7CbnRXWYS7wLVFNHdlqxAKqLLYBXp
pIrdfPwA9SkbUu6skpLLK374+eglR/B7iqyi2IJk5zymjSxyqH0JYa6zud++mtF2eHIVyZ/qQf/v
8gIzggi9euu6J3lzRQ8hIh2RXLnELkZUcl/tu1zbTjZ0lFPbog0robQtQlUSU9jNndFNldZga0rp
/Ot+RdiUi+KAtGIWd7/jsZB2HQDooxJNCJftIfDOlpk9V+brUc1CRgTxgnBTUaywagSoxMohsyxt
iy3kUCZSDd6+I4Gjj/ES+G2Ahi8suNPXWTbR6pVIx/PfEiFgqhfz6G0P1TcuLddcqZ2pGWP3mgxU
fWHmsXVgGbXhKREcTvsuHtRGuwIQHWeY1YQpzIU3+BU6saPlxxQNmwUCJMP0DB1IjihE872w2eKu
H84qUGnNLLYC16CwJgQyw4sZoYu2ovpDuzEWrEFrdbHGdlc6D/uXSucVUJz0H4/cadt1BPpnWUOz
t+5bxsVCy3FITOVSA/iUyvxvZhmcf3pDxq8vGRH3h8IbxKx+9QoSkehOsc4i43ecHMSMw6QalfCf
7Qeia6a/L1+nZFIj0WJKr1vUtitO7GrELW8xWzX67KiVIht/peERTZIHETI2u++BUXIZSCO5CEHC
WSccdmJvdHQDGb3AQbtR8rnX0oMjFXQ0aK6jnubzcD24Enp3k0dOQOBg1BPDYpcB+8oUWsihvMVq
sosYr74Bd0ToCGhka1MtekcKsMy3Pien7jplDMUl7ZipU+q94a5dtZkzR9p1VpAW5qwnexP0lMQx
ABHwnn7ZlQwQPdjo7lM9umF5fWlmvWtHCS4xV9coacPZMiw8tB2Ug7zhYxbUVwEIzPeGLLPdayRh
+xLMZkYMtHRrKvVCOo14Gl7az+538lb5IlPAybkrYqygjiXWNarAVRx8glDLURFp7T4XbNJy1Rgs
3NLexSdIXVld+P95Zc0r84Rqq+ENtve6guAAhKGmISuhOSvUt+thNDMkInK8DxfaUFaNXs+gKdbw
tS5gGza+cnfk6BHpb/78nwqH9vEn2w42dJj2KmEijBHPL0vK5mUakz6ElT5GvbhC5KC3Oy/Riq0Q
8ZR8WCRK30df23fuXsHsomBwdAA/vGBX9FYmU7wQ0haQ0csHWkrDt9vg/OJaByi/d2TB+5ETS2/r
afkxZwBaNRBdhKTPdaQ23flqI/Sy28Ha90mmjvWAorxCwuV6ht5DqSrwzXzCYA9NqQ+OlbG7gqeO
XlrthLw2YOdwjnNnqinq1zFLwKWkECaBHXmyqMm/EnvjKSwibXJ8rqBbRYpNasA3wceZp1O23up1
FbBGvlAP4Jk7eZ1iq+fMah6xaphlRJJRD1xxM4cZvZHm8hdqKmMzSFVCEiGqwRbeDHvb/80HLKpq
OdBcdHEX1798hnF1sIjBD08+st3lLHQyQk4646gFjwnIDXYHWDmKPUzJdgjMlc0IIKf7YafXY5hO
/cQh1xp7rXbRAEbJB4D9y3SPObVuSLf+tvV6I6uxjMR4N2D8+Vz6ZdJYjN46ITT+WoXTcC+kysP3
nYNy9Mas+Yowa1YV3Ake1RyPgFba8k3Wz7BnAbydN74ZpGxQ5coASFenGC5AX54+ddUXnYtrLvAf
HQwS3TTFKA/La/chC/kU/ioac561yHZelIPwEpOSlnyhkBRhr5dV1x0+9Pzrc8pK+OYtkpX+++ZC
6h/GWLXfpQc0KskLVlmI3Xh5Bemw6WM8i7fy7cMqjvM6jY28xoUr0qyeODq+34C8blwrgNMvqAn8
59Wr5xCVNu5iqmAedvutqby/xwcjF3y6xHzEQO+3xhjD4tlrYF03xuIpPY8iatf0mmq7gEKkxa3W
JaZ5GHjvSPZtHqcPA1llf/1ifujnzcVMM+BJiNhfHjPbxQ6tkLof87Ngr8EBFALlMqyF1rWLktaM
QqyUQzD9gJ9hHToiYxIKi7AoZTcMSp2RVNb9fxX2P4e/goNNbdb5WyjfQzl1OphdDfV//Bl49SvZ
cXKzkkeIlk+moObK5W5iYIVAsnf9AXxIcPbM0xO/ArLf/1Qz/5PWTZB/jFNCH3MLghdqg8+y0rrx
x4waHRFjK5eunPt+52Vq65lfkiF+QgQDiFk0bN/FOs5CSGMhjIRgwbSiyScrUiDMVYqxu0XrSapp
3eqDW191AjafDPRycPxg/iFlDOX5G+dERT7ObTqmI1wST+vvERbeZEWGwJubJ3HnYx6rN5eh3NJB
f00mUPNaFMGllnshCMbRiZq1ZwgELj5N+JAKmYDAxdA6xQSm7etNK4SC9lQKregcx0XRP/Xqqf1F
q3yuAUlwzHAQq12WOz9Zu1Ev/3Wnvm8B/4Zg/Umv7Enjx9F2alVDJ01Pr0yxTYAlTI3dug+zhmUI
UVHSPe7rok15I9tixxcptMGWCmX7fvzJwYrqhanTZdJBMc13pJjNPTuo/zI6DT2NRCW5f9sqhoe9
Qz/aeTa9F1j+eBBJBfgL1paUlw0X9IGWYyGbVB8DKc/DbKeYFd19NK712H4s8maEP+ZYDSPVTbzj
IeeRhbaaicTMq3KDZmSAlOlXQJx7Ko7JdOflZj1TvbAM+GPH+ft8nmJAZAXsUSZ1CcmDBCftbZLz
xAZpoAdlvYEGKLR0YKtH7FvUAgwYvD+jBiheUaE+3c1WL2BhIoWGmVTHVrMihxx55h7kqHutxPRz
5UUcdWkuLjO9THKIaCnugr0me3SAAojkWi+uuVqWTWs3vTtoWK7rRjYpyj0ieDji16J/MIH/atNW
9GC4CT0Kc9j1ofOLEPtpici1wS2z/w8QhHhFNjD2kxcSNR76O2dZoCufKlOHBSebWVj+VSbhgn5X
f8fIJBP3kc+U6wzFoHWCNDeFLudQrb3PLO57B0eg36Q6TGtugdFyka1ZvMvDKVbwXbmEb+S+O9Mx
b2Xd/UGBfmCOBn6vXbAuM8vrJaBnstWjA41h1tYMzod2Bzfd1DUWLNDLL2zg7FrfkDnZ3SJi9bA9
hHi6hHUVQxk+5WLe/A5Yrtl8M5ju+Uj+s2rGInkSKtKnbu1ExH1fO5Kf+3WxI6OXpjiOVSSeXGHs
Xv/vv8suXFm+frNItwy5ybTTw939VHqsMmWzVml0B5bmVWrtMOvTs4M5zsv8kDZgkL2rWWBB9zBL
Q/IrLcBb+iFvktmKmZIO/7Q559YV/g9nPUAmCYe6/EIXhEo9djlqZI/xmWfg44Q8viZGBVMiLsmf
yNLzyWo3GpIIePeQzH7e37/Ib8rgk28x13IfbBgEge0E6PQCHwk6Vlqp7/MsLX8QwNuT0wxwTmTE
mgOsJgKVfneJeIhmulPt33DWsZLk3HYxeRC1hD21k9AFqWbi94/s4c+EWF1XDGZQj6fCoyrGG+/h
WJR3IQFTwozV8Ha6KgQVPsSHcoL4TTUY9Ieqr+w3yi7HirwSjOi9G1a+AYgyVwMXEyDrJC6uHKK9
H8Je5/A8uO0AdmJCoxmYELr6dwNlFcVIiOdygxVL4FlyR/vgcC4dQBHuG0TGiHOqCmg8zIKRRCup
xToPoszrjQ2V97l5xUsqdiBG9Ajf5zkpbV6aFeMTkd+hOm0ApTYGtIL3ZDFzT5i2Vn4rRr45OEwv
mJXadkuJGjI9B8VgQpFWJkk0jxpkOg5qEDiQzobo4UvPqXRjDKGMflllKU92PboI/28m13xRgNUs
zfi6X3LQQmxH714xBIHbR8FlVnn4MG4xSv3gtnVIGrD6i6MWJZ4PvS5w9QXdSrSoGz9+FhNMbIDZ
JpUvEQLEnCZbMB3Fx217I/aAdF0qP7DN43ZwovVpXb30P7AGHkZpp1BRDYsIKwCozo/F50H8DIeY
Xy8abHyA96YFP1wiQNVC8lg4KNOGaR44W5RcWdhr+ttHnDwPYhIriO6yOMvgkbdYan0ZfVn/lfgv
f/yefPjA5U3tmpDvQh7Eu4L5tUmJxU4ZBb5sbKkA/KsPv5jZ5XJedpX88RfoJTSh8BHl1Yw6YeGX
gxLTSbrzCufmgTwIIMVYEvdwtfn8LePLflHwnzhe7w6xI1+RKpeKLtEWPfdpc1M6wJbmfnFMVHTB
Nc0kbRvsrLNRKekAR0f6DesG23egceBBOPYZCqliXzLi+345GSUda4xpGnXe3UyH/rpDx85blJNh
DW3bFesKTSnNl4ab5CvJnWXo/79QjIEAG+cHVOW8Odri0xFI8kNwehygzujv25TNyM5GcNaF+AvV
hq0e97GIetSKQABpvP8Z+iCxVGgwDjQoT7pYmHK6G9wHu0idAAxnQl58oGJCcwVPN6AWwF19g9M1
f/V4ZwlvYpT9upiWlANK+9Gn+vKCFjb6U9r9Q1oISlhMI1UHBXeeOT0/OXvo95/ZRTlHipsJyFeH
a7J2ZuIE7NWAtQqM2UF3Gv8QANmsWXHgD3pfIou6bRJ85gUNM4haogNl0gerUYOzB8Uc99biEEyu
IKMUZw1uEqDnhVqYqeCY8jrWZFPKOU4rIXO/daK7gyDkDQthypmJiqF4u2cQ9tbVIULo6RN6zhzh
1vsCxdfuGtBYXCoqB5kNc+RD2hVNEyurT++X6JlNlaHcmGPQg0S8U//+tRuylHs/LFzO92HHX7VU
6p1fWn3V7gUdHgFUzYyRZfDDAPgSY1UBjR+Cc6kbgiEyW3EMg3SwLFosOvjXEQHUL5KPd3y9mekv
TWIN4hmvaZmTE6tU1lOsek648LxpfunDv0+YTKJaNEuIYsfwdLwTpL6VcLdFZIYzqBwpLeMeCGxo
S+Hwj8Z43HGJZSTcBvSWfB8wKSkBgBKWJVxTvAFV3hZY1Uers9GF2KRGuqITM94aUb1ryCdxDh3b
FBJ3WxzBsXGJLjftvg9n8vEg6H4SlAfJzpsDUnATje24piv7EUKM0N9HJhOFn74gOqiaP9UenjX3
+JDzsG4hxDURgprLxjNFtQFhxvq5h3d/NkzkNz7oFovBNHUaOGWYWIZhs/dE/tgG3boxqCL45Lr+
HzVc/AG7iExfDm0omlHrqsdx8m9GYvChtDfoWf+4XYrhgr1lvhlniVQjnSraNedA/n20pCRMFD0/
A1mPi/iNryyPetNRpIj5xCZ1/doImpPr0RNkgeqk96L2pX9pnY0nx5YSVS52Mhfq0QXpUKu96hoW
i8qnNLzqP4oU0Tm7Wk5KCwj3ssuTbiyzEAlnO6J0GKKcqRZ0PUT3KDvGLG38sCrstXv/EvrQmfTv
FF4RU4VZ6SzFwLZHI++7Iyu50a3vSwSyA+FWdnxbf1ze+Lr3PLrxGwH2wTLVOGqKIoAopthzQP51
Qb1I2QCOife5oziSvzY9/02F9bjGmvKN3SKwg8hne1Jgq/TVt0ruKjkT623IJYJdDF9TRDl1kVWB
Td8iyUo0/ehr0U5KByZYzyUIAehh1kwDj9thL9NbX8w9UmYmggvT/k0PWoO5/5ZZj8kmqZ86PXPl
NWr/uaZkslQo3qM2eGPX5/BOeZRBWtR2r5+Ahbmdq6j2pUDYGeiqFCz5fpaHL4kbJ1rfemf+NpYj
ro9+W4ij0CtkVLPupOwlfN5y0N+OVQVaj2+79yR/3j/RqUxP8YmNI8Fn62e9fw5jWspke2DSEVqM
/T5ZQy7i+vrmaakHTghvf/FxG8wrp+RNLHMeoghADXv4lMId9Nr7YaSEgX+qwXpq+0BAoSXrJ8ac
yyQSzQZt5PlEIsRXEHE4yHBteoV09r23FZCQ2UqgRmT05luhzJlNFICcTM31yY4BO2OKZq7EJ032
+sD9jjK1n0zVjvdaIrJ8vb82csWrBynpaEg0grEhUbDLnjUHoSW3NhZHv1C2UIRPL3Ui4/uRQ6c+
eI5QkK634R5erTpJiI3FX86ewVAlXLoGEpYsNIpXEQm6RWQvJO9d+a1YLDnCbc7AiI0Va8WsTtMe
umZBvURiRx/B8Evz1CXzm2qzcbXEQfEZWi+kv4thNpSv2jL8eHa4SumxjCZtXDc26XoKN8ON+zzw
gH3YJeltAEQAvI5G+yPhH9eEOEEtF7Dq71YY7cZwO/APuVWoHhfba+8Derq9PQB39uelFXjxG75w
Bm4NdBsdxx0AF8ptLVXs8nZUxwKQrIO4T0tvdw6XK8bkUaaAzOQ6wM3VBY7VHokzBWzhVjd2MOZI
vrIOJzMPLI9lJfJlnWaGPlDMpCtYmwFGO7A81e7bqeWHWN2/bqSoBA0a1FLMgrtOuIIb9UvWevvW
WMIgW92yO6nXws+VYjAUBJG4Dsjh9USgKA3nZ8vLbUI/jvnGt/nTJWzVejGtB55/7OUnPs4hqpW9
0ZvCuwwGCqTxNG5mrxKZnxJIZyZ1c+S050bei/msk1dAZOQnP6NYwMmpTbLBXvZuJaqmWkmnMSHb
0x7SkPRYlYnU4AGRMqt683Ojtmv9sus2Yz4Bjp/fLuFIBe/L5NwYpd7V4B+ONl+k/r81f1+WLYPu
8zA4fp9+zC7Y0QWh0GRNZvaKXjAolxG7jF6tZjgJEL73Eii3EwIaXuZeC9fXhof73MrY0qQEmlzp
sH+0fK+JjgbLl1iuJC42ttAqooFc7GDUbgzQDvpX6BhxEDmOUfxKb913m00H+PRrrEajhiFiPfIA
93R67Lfs5wGXnToTv4zrPHUuSZUfT9YSb4hRsmiqiyqeuxUfWbwlgumj1ODizUZt6Jkpjb9LUIRY
TtNr53Wj4L1dSGoKWbpdP22C5QRD6qg8BVxfvgjAqC7Fw62bkA7EoGvJAt5oq75dd4p4FTSb5EBC
R8OLoG/GM7pR9PXTBZwZ1gSovlK37+QS9PEk1gkK6JI5NXYxyq3F0OiJUcDeuDWkbhk3y2HATLgx
lgVQoxj8nylEdulrO6pO+5rUcDbu4icNJogIxOM+/88eqXuHLh8PzeGVi9+RQElLCrVMM8bptkLt
t1hdNfyw9MqSrxa3aa97syvOsIR7j/LxGAdMpkavatGGp2vdOO2Xn1hRF1bw/pHV/lP3M7n9wIlN
jGZWeBoj+8tkj9wKS1rui3QrvJmpR9RcSPeKMBAIoV6gp1err6MXlZnM87de3LmlxClIrbfPUraP
/R1Q//4xIXEN3bFS5g0WGJMoEZBBsFayFlHVp1bl/tQxDHNSqw/8Gh7ZjkArJUZ/oet98yM7/pvI
3J2KNEzvluCOlIoeOXNFr/KIbkkmviYtM7du6KyUZm17qVgpv7BWxfOTzmLwAFynJODLM1nAgm6W
DkR/n0iUoeMcBQteL0rDqICPQCWkoZr4oejjRtQX/RlXKa7X66RylBW3bFg1lRc9n5UZWvWIrlzm
TXf2ky+2EqCD127CtM+nRzu1tpgN8xO5ehnu/+lY/q/ll04h8E2jfxRNOAXdgHk//x1A0jP/Om0K
RUN7FvsiX3kFBl6LD1ZMoc/tFrdXGLvv9MuRu8Ew01lSFMibdQAgB/0jfQDff+I5ZCeHzAdsJ0wL
38S8JmTxdYqracvWQE8qcVbUxVKxJLvk7N0gt8is2oHt0gR2Agdna/W/mBC8zdzKPxF2Xa0mjGVE
ZV/STIatVzAg450p0SqfGShWnTCve44HXAjBYfyi1zBrGqNAODzKmP4OVL4/V/m9L6oURdV7PMm5
HV7TR9xr+cI23hcrZNgzeOgN7+f2I0bRf+9JE3hX7uHDEPYReWhRYMdQlzxCGI2rRM+ggb7/Dk8X
ZTs3Ob72TvGu7OeEklHBVSSjYi+jkjX6BBnlzSoBe8avI6Bue2X0mLekwzNH3tPQRc7GLASu4yYx
KQAK6SyHotF2RVNU0gP62M9tALPPCteNF+3pIYKPf+ePyK08ssoowKdm75UP8+NrYR4ysqV/Ne4n
pOFmLlvMdU+FuxA5QLE8sqgQL2SYiPs9KEq8g1BpbGF4Msr+dzljKwGlkNoPf+mJOZnxuhI1ZJ8w
fqrwYDlXLHUdAKU0BJHG+tIAbNXm6S7A/uoAK/eTvCM/ZlPWJaKC/uwD7Vo/Z1/353d2uQIwTY44
lzfyMDz5FspjtHyEWJuzZmsPASjnRT2IbRKO669AYhKjrNdrp4pRyFHZzf9DquME3z1V7fXWKbTE
VPIcYABgTVhJA7EJNtNYihgE5O/fvM+m7B4adpHiqwHVa3IHT8v36szdjjSgtSdD3M+OXv3VS7HG
y7GKetbbnTtYLqaFzL2UziX7sOl3mEOiWHqFQj2UleFRhspJx5+Z1AjKmqZcH3Y9jndDQHYAaiAU
X1dTaWSotDT/FjtAJ6BE7tYa7aoTKPxQXmIHlgCjKhANA85Wv5u+RhAkAyKLCkqyS/FIPTFPT4MR
hRlOTm1Dyn42XM0DQrpIKIb+NEmcF/AcnKCuXuyrMWhIucu+q7iQA5V7rMf1heeNOIU6gZcIxw9j
GuvYyrjfLmDF7dgKxWbEhG2f+w90XL8+fOno9gCOeKnOMtNqFX4zqubbN3IpAzLH/eHgYBEZlwAE
i59oFMFMEBczfBQFtuwFZgDSq0jkFozx702re4gPe/lJTX6pUN1BqKQZ266U0xRyJ1tfdvebxkQn
y6wIgtZIMcL3lgXDmy/Chm0nkQxlsFi3AKi6dV+A+RnqqHlJCfMSDWKpZKye8fHvwdkwip2oQJuy
3gEVepSIjuFeFmmXdcov6QesvE7iktFkpT0pTmrRbwooFcMx1vmedBB7Gs/4pF8c8xApR/dcGH1z
narbe0eqTXdIn/4wp2+k7TRPIguytUxYyhqaQU1KandMQ4RJYzfXNXul+6FZKVHA4eP5YVCkdpBG
g0ctuzYjcNbcaVmP4zkKsT8wAWEtPKtSyd/S9QQ8AdLqkPF2ymD0AjXDgfLp18mIzPmjzrXG2isI
uXKFn5DYMF6GG7OLq7vPvKCsUiJTmRMywsET/CSN3tWyfW650C7x5PyCJ7Mcv1gPvOvyBQxyiKPZ
26f0NLkIiGFw1hFk1w2A6CZ8maC+vGzra3gAPEy7YruK4WMFyuUVOj8QS+R5mt+g9zhqR4Eb1N4e
0UFsvk2C8GsGH/0Nh5vITqIXQ1U+X7/mNFtibbodtxwqIZXFGJx5ALNnL4P9dN9OFjTobXA56qxH
AjzWRk9Op0aaUFeLsxrF7nWDVUKoao8m8U+OG0OWpg903SQmuR1HR6O5ZQn28erAvGGU7N7QctEk
kEOwx9NumLIXvXX+XodAD2+qXzVH8IRmH9LoDuPZ6uAJjneM1UG7WxVtsp+PR5xjr2JC0mOa7Ud/
rihxdSi402eET/XnqYLR1iyABhqjWYwtAOfi8bxPVURC4OtN6xetvIkgWndHThSktyTZd9bOPTWy
QDgc2FZLcLHAyj/jQRESaxv8S/pKJhnGkmYEfXtNPlfUuh1m/UIzcuftodFysSzASD3fLxNomY/2
8bIaIz9SpE8w5ITUyVZ9Xawrt0AVr9ZU9qaqbZbEbJkyKmi0Mq46xXIDGVwwyPRQqh8cFEY4v4jH
HimreGBQISZm82YG91TdhPts1q/N7klHAAEnZeIMwjxGeD4HbcLAc5OAKZ23B+Ekv2VqaAkKhCvr
YMqxprg7RyZPla311ozBnB26ndHW8ml/zT9zE3SWfDNtGUWQXkzjNG6rmxWgTugB7gUn2OXhVXCo
+NJ4xcX2TsyVwNILfIGxGLxe9ce3133zTxvQiHzldRNxy7Ob3R1tO/ny+EYjqL7lSbbZkIADLNtZ
FxjaLo4ilFhyzS5R5veFJ2DQyVHAGAunpyf65GKLOU0xK/hmjxYoTCC83z0IjZl58lVzYaAtQHOt
5/0AV80mHXGg0ISaIEjzJa50vJ/xlBImoDW6zeFKjzMnh/urbLtvHX0UG4BRpnfFfPT/cbHBRXHr
xjJzwraQcjtKPoshM8HxM0KdyKabUzmwHPyoG++B6GAvS4xY9b0ivR8dbRPUSI8SH1NM96wzChxS
Iu2IFV4mgFcFv2HwBAenClZfruchlSHnG9u5P169zAZMFZ6tYbUKAiR6R4iNkI+VC0UWMVs1xFei
F0VV6GFWGLnszanA6V6p4/8MGQ144/5piu/A40whB82sAAjGLI/Se9SYDJpGwXxeY/S14xsUsW0C
JbQl1ptmCORHWkdx5epD0oUJJNLZs6P9gvNxuFGkPJlAWv1Qg9FkMPWgGRPzLUmyKf5Px4OVGTbE
oehTGlu40CynuDs3XtJWmKYVcRmAn1qysunspMP3Sjhf/e30fJ7lpuXtqf+lxbBoqw/+YjJ364sI
5ju/LjkHdR9q9y4Ou2Fk3ZH09uVRWDc1Q9gF3EdEKnvCeJ4XJMR4KycuXI/dqEebDODqFGMQ95tW
a5zQfqEPU98eM3njGPkw4Da+sl/hYz9ZTna7m8ffQHAZ+J/hNC7OLUhTWt4YoQiamivuPO3yo0TW
xheOr9chOlSj7c5nX6ajS6zXB7ChGLbbT3IW2bMTzaikcf0JdhMe2i0Fa99pyDV/GgBdbaHQ1AaQ
Vx34d1gtOe5p9qt3VOJAtXkxUbg3uqrkUEOzIsPs6iwgx+a3f8ExbwhhOcgek6i683jc1MHIGFAs
288HUYiEjC0mEDl+Ez7tRF0UbKsQdDktwLcboiL0QUWm9In/lnYHgw49cRVcuYqxCvlQNzmxW3FI
Ur3pRm9Ov5WtnvSU2QgGPm7FxuckzeETKu6woGBrJbBXFs3eM+kRdyDdqsGWBgU7f45GmJV2u1no
AdWnnXcCln/O7Kb0/HubAaE13e5XPPjJ3+W3ngmwU/WZECjxz6Px+t2AjBWHNDAozd42zjF7T8F2
1t5LPxi2ctD6I0FyDwyvsUukzdLgybR+u9LJSQUlpvvVo8/INOc0r+ZiILC1TvTnT+URTauYJCwB
ISrlfxaXA1HksRl6+645sL+3d8nsiA9PLtLv6jTNUKlc7JbmWW1k/59dlQW56S7BxNefuv8a8DVL
Z+9XDZaYpJgTKcRi4Ytnivubk/nhUoX28OjZJNag7qEj2b2QJx7fBFb4SLgAndbUcjnlGxFcNAB6
j97VIstMtiAUHT24fNfnftICmsOBCvk4efvsIcuqgTEZWgd1/+WyLC3ZcGNPHbYFVn2hvebTHBnx
db0QKeZyBVA/79DreBcQwunqYBV+6QBsYwhRSuqjdCsaoE8Zkc29Cl+kl59MoyngjQQe2WnVrTWz
UkrLpwTHWa3RkGsxVo6I8524WKhAc+FdZTIwWEOYhAiKQa2lj5EUyxiK3qCcKTBEt1GbdeauMw7X
DPxE3c9pZeVrZ4A+4Qv2NvscvslTmjrz3AqPcohhm/5oxCggI5M7K2o9z+SngoT0jwgghKJbaWaZ
x2G9UKCxckAU+Svd5qwOqO4iRrIrFDs+br/kYyTFi5BV7YQTGxZIC59X5pDLHFul8hc4crPPgOSm
gFDBJQ2tr/hyZ2XaLr8ULAs3DcsuGSRz4+zHTBjdEB1qF290EvKvCl5ewb9kRSwe6DFugk02XVv+
CEJEYvhExi32cxbeYowRkfa6uQOGVoUmjj4BZUoP1cxRcYhwAUVW+vKYZvDq2PzDNzfNTiow4nH0
vF4WcVfgt43giXVsP5/H2uCcS7qM1xgJjUUptfHW31s7WxQyVOsJ94mCeu1Wg7GISVxyb3xn4ifW
GOr4AKB8RjMRYw+JivuSsr0heBlgG3NdQfBQkcsdJfu8gV8CdGkpyN+hipZBCvBnVT3LNkRFschY
a8OPYZAe6rcWTIxmaCJfIqjJkAQ8gXCF01y/SUfhK2Ys4U+8FxoZF8U8zW8Dez5pehP5wXAtB9uT
o3Tgkm/HC02X38yuxGiLrnBo9tOpQ7RWhid5dEdfViOKXFWQ1PwJh+nHtdv8qPs9GIF8p7KhVaC7
6XgTPH1z2A/nUOn1W9DArH19Wc5qqr+p7GQNq4WI5/Bgf01vPTj7S9tCHnEyS+AC4ItdGisL8mNc
hotWwRp204w5e/JhTusmCgyYOQI6Y60dkT/Rky0El/GObF1heYUXG0xjMgL5DzYtE8kihhNQxpfX
l3dBuwRdMWXFDq3ESZOM7Lc5A/CZVKiVKVcvAlgLbtHlJ/UBanUbOqQ8hnQg8N/SlXDrI0CSrMJD
4HpH6AVP8dQAxmKPgBYcqO6Y171YDoyDUdbZMyq74YfDZ0lVYY0e1yz/pn5chwXej9SW4CTX7iRc
Qwu4FkYgdlqB0ZCD2QNCkFS1AwCy1cMlXhf2Nfhr4XFKOOHXOEWLjuAZRsIQuUFwyhtRYfV8kdfG
KJJ0l1pkpF+RCS+iJkUIeCkal07IQxpnMrM2oxisno9tMhz0tNPn8F5Tjyv5zsBdiJi/FoNpq5oi
nL3EZKY9OvidAN7H93fFB8LSSXIgYP2PMQkbdEM6Ka4wcbOIcfWfCWZGpQeUTKOUSYVHuuIplLbX
OxvnSbLBCZTeATsBXxUmYl7cRLO5WdjjqVasmZjSV2ElaUD9GA1n5uSl3gcxbbcS/39p1XTvy+1J
WaCW9Qklzna7KF4FjdRbjtnjhzRvY5YcRl7FQ87UrMDH700vEEBVVMaUdfJ1lASyMZPicLczgB9L
ce5FQ+4B1SzF9hhbFNO+LMUrEuCvZfBzigU481y7wa62SxE4J5dw11B/M70YJoPh2n9ASD1SJJWM
NGpleImBvvMc0rXUPYVBA5+gcFL7ENhhL7zEmNG4BX6xX6kkmGOdfJjjWS/CmGvoSVbg4K7wc1hW
Of6fY0JRlMkEVztGJIbe6w1SpaNTPWyrwdO8eRmNB4GNmHjHfcVrobfY5lgsakj0TkWdkepRnjJk
zDFuiC6egEinlaffnE5vAzqvGDZaDIUme0jLlm1sUGXLjqKk/MQGJGD7fs8WdlG+XXhpLQ1HU/VH
MvQmTkvDtDCVEQQeP0kW1rOMCjoHI4uquhAcE/7481xoLCK0KWYV9ysDkY99p4pR7dPtM/EmHn49
xczEyFN+On7So3cpNUPUirOzVVWCP0yanhoge4AV6KFjuazoIvyKFXhxu2z2w/ZVJcS9b52KDmkq
HgClqw0skdByu02eVc5xwDdfjsMvRKGRIcIZD1NplgHsJv8u91R0S70DJXVY0ADkVRea+h5VpHKU
SpcX9+KLEFd4SLh69JpWdMfkFBiCyN95D6zpNYOxd6Y2j4SRP+F9KMbZTrCWQY331ODARS7IVO8B
G2B4fREU0ejr/dt/lm4DjbV7q2sVNckmlosc6lQ4Vi7Qq1UhOd+d1MAlodaOBSLVBn65+jWhfq2X
F7hh01WeVQWTmbTO/v+xzkCyPNs20aVfdXs+T6gFmJ54pznWFrNJIaGWLWmbp7Xn0iinSEHDedVo
tha+29qG5Ya3a6H4mJHmhZ+/u9LdMGunsAAF9ZtChBPvddnRHTE3k/4r/rE7yPqYfZKcjseNeMnu
GmMaB8benPDQp/2czueCEQxZHE7kaib75k2VaFZL25DunQmgFZhABMHi5q0wd1gYC/97UupWzmwn
EFK+xsIxOKAuRAxHuZ8DJSeyEtZ8+xIt3rvWjHx1p6lYgXBdI3fv2PXau1OeTqb9oyPXkumcDgGs
Yokug2DrsfIs9pEKmlRy1mjAV/cOyKUUzrex8tddV5wTBRyS6BDg7IVZZnWCM1YFhzx0FQoDxalb
kHnldIIa+kgV9IPSw7nLVVTCjKKWObFiIO5QjffTjtuE21QBNi3mPtWK62RdPRlkniayU9my5ZRV
q7QkVKeXxtrmXqs4UsrQz10iMhTdZh5mr+H8IccYZ91XluZXaITIMGO5i8/AQceAmFxwanGxGd04
iE2tV6aW3ynWaDGnXxKMODQrHxnSdgEToWiF7EM+CmWQOVKNHwHsgULAEC4mGcY8uhoukW4g+FxG
XksHXVnGVDKeaQymmqCIaGEZ+IJDaOhyvHowEHTLRURYK5n4YBE/vMrAZRGLU3HJi1ZVJgoFTiLS
3yBP7x4gzpN//UteZ/PzkCUO6ryzYeGhvmp7EISsmOavLrJIE0fTgYV/Vu5d5Dzevc2XqDoyk878
MPuylyLWci+GfapkMqA6xP1gXRmSV3d5QFE2c6MTN3oPkiJxhaUUdq2y7IBqdUE1Y9Jc22pob5+k
S2w7VuGbKp7F9bk9Qz38TSGcgJuKZiciLWFs9OAZZyAIF9bsDYR1a5AWzCVLUSg4mgKdndgzTApn
qR3zYpr0QoV5IqwLtsFSCGr+RRd2rmLiGTWxT23Q0tSM+ljwDeSlI1Kh2wSsy1uMbstUz9TvQCcJ
mM+Exuiz7bbTVbKiwKIEDHmhAzSaP4EQK726pHAxJLzylVc/YHn9pNWCjCi3dp3QkgzY0TsmnZAj
Tgyv7s2dNuZulIzRSfeSVkG8/s+hqBFV5MnjrVISe8erJ5lXxSfCzwaNdv7dpIu9k5ThPAWtjWxR
rKA7SwmRpKeIvyBBS9fjAFqwScuW/EMx3hOqJK+3wK/U6jiFuW2n8s6YfKG24hqrKuiFJPPKJVl8
UNcyYiSLT1d98BEKbujM7QBL7NHQmqkq1fGS6dc9rDuho03pazVhbKscjHwlA79OyPnLFFpV1HK4
vUEEAH+mREXtIO61l1uaGlhotL3fW2LS7HYEgLt9QfViuC/027dUx1vGaRCQpl16PjULtqqsrAl8
rQCPpghYeVowLFghIUZcTGEROJlqgBtn6qek0EcLyjRMhkwpY6uFVEwJIZRTxlnTfhwNusvbaVKV
2N7mjYTPRLkm6AZ6+LO9yGifx/jfoCu7fUTVgNk0XYLlRN3NjOi44XLXQesQdsii3GU5OC6gRjnw
YWAop+6XLMyvrdWu4xsEUdBJMq3UqOedWiqydQerza3MSqsmJT0O4myEyPYmvcpiyzGq7iW7Gxz8
/AUVN0aLlUjoDJurLzSHGkC4QBiIxpRYoISIXpfJ+nuMCTXq0TjcgmfvMX9XaW1jBA1yzv+WiKJU
nwAxpEcPBQbNd52VMF8T3/vVU/GjfOQmg+um66oc57ILmhdiOms8FYZebrFSrWOOzfvOX57YQ65P
Ow1Xu7znv2c0xcTTC28Wv9y2oKc3Q1Qaiy3Ric3PGZkaiVBAM9nBwSKnUROuk3Tru1oRsjL91nK8
uEbOjt3fw0TARqY+LEYPmtRGQ5dv/5ICwe2bfrdFDeGC98G4OC1Z28YoDABf6ADnzlja+LTR4tnz
M7diiYEsjl+U3Ifdj+i0EgOKkxcsjfyMRIJw7Trg32bv1oVNDK4IBSY/tLY4DQfdWWgdt0697Bu0
5lDcqkKh8ksJE0amDppydIvpP2OqgEAE4QKysxYfeoMLHq1nP9hGEk5u/K07ETN0/FUJLVFv6Iw+
mR9/h22/89q4Wdekbp7jiMX+TMBI6w/QqpXQbI9erz5ufHNHP9Wf4rZ0QybQdJl8NrfUdUFuosD5
tknzRXAcMoBbHkbWa5Grq8fA6PxqEqzaZ+IiIyacwwoi1UXTImNrMAug0eRsSOZLu7B4jj5R9kxV
ivwklCNp2McUWehZf/oo+EsxWE1y4PRRZwmQah8qDZDk3qa3eQU4pUTQM0JUN/2DCM82OScg7pRO
uMbYFdazGCnUZXtvWl94FUe+L3/VaxR5PydnOXW8z1Y/ibI0Q8hhJv2ON8M7FOKfpkri3kNeTCe3
nHgS9IfySSidCyAYSTxojldi9HgDG5a4xMKot4U6F78JGg5MryewSOhDd+63WoCuwt+6LpLlSAU4
caq4Ptts9cYJOBiZR6to8oqBEbYfHA8HUz/Iy2Shg0SQrmDetAhQxsQZE1NQsTYILuAsXC1HylAE
FHE0x/zxHCYlVQniqNoi8lyuzr/TybeZloIim48N8LTCWUyaoYatajjQ/iFj9r2YJJAtIwLirX6N
Dm/qDtz2blgRj+iEqQA0YvjjodybULy1yXLSihR1TgGYrbh1e3jQotnGo0/pGs41LII2aqxZWjak
NSZrPmK4jzwwdKc+0GJ6gEXy6UKFwUA0dWHzf4dg7LGbuoU/Mdct+NFgRhDT0JwHe18RqZ81nu/V
i3dehkeeT6ty/QnfnvrjEf9xPe9srwsnrqm60z0qpc7WZnbM5a7r5vFBIvjJxnhNLa7btYHJWgGS
3CXANvt9ev/ZeWEzSL2jOOceC1bID2syMOEKoejSljVuXMtCXQAIqguoSqd8A/7TilM2RidXO+SX
VMjGijX895N76pcn+rK/UDTcEeG5Z//xhD4sEf3w95v9VW9tiB4kW3bvBjwa7fpHXpDp6QdsC2f8
lrnXxNGw24T4O3Xi40U0GfM96IjcbgZUPrsnMneuDYyY4oyosr13H/YXocOGKWlW0qtYWnh/h1CK
Ht89wkKMOchm9O+FnDXBGl79UH9KmQ+ZrYUiqcr09ifrFAugpqdXNwLZXbl+OIkzVvVrkgW8ys3y
0Ih+4TAbUkynOK87jSCHrIBSLYVMY7OwW5E0D5C737ShItzxPlkvM6gL2fHg26TpEVweziQjjBzH
xaUhApV+iscJ+EShen7UTEKAR7EwhjL2QzAOceU1tS0Cgu8ihRI66tqKfTYVlTebKHy961A90JP+
6MUcnR1KhFA0EveM4OZt+Lj/QhLIHT6O+WHfMP7Ic6u+bnh5b4aZ0pqn0tl2CbPY0dWve5kqT5X4
x1TIkN9+nV1nN92n1Xrnqu+jJoB1xz5hkvRHVf3jDjzBEJfXHLqXegI9B5fXjwzaKcvVC03N+3Lf
+LGRoeYsKKfPGzPJYzRzoQV1nTbAUcd6rwFAPAuiHObY/GQBk3giWvi20JLTyFbr82LIJBkSA4mg
zw5g1NaTaCy2O7gyKGHeF1bR9IdupwZoJB0pa7KPjUg7J2ktyr1XNkeCgOsB6CfxRX8V3a6pIwgI
MMxTcIwvfCusKleEeJ2D3Q+eG63aTSgkaZmVsDZTUJQVdHd9yXWdbo5PO9TPT0c3xLq5ZqEOJUwP
FKzygH94vg+bheDRvyCEEYPWX6fuv+OsNQfHsT20vtGwcjyt17V9pbP6R6tVdj4woxn8qCqZSTpF
E4bsIHECUuAMOB1ncY9+2nJ0JuyFHv3WsBlAS+j4R5gQRmq3GZ8ED+Nh3ZV7jqE923S+xGOzyYH7
QeUxFKMCwneVmMDtNtVX5zZ7WleOSw/FkbX/w+cv7oFObSLD+XMYXvgZPsbbPci2uN68r4Hw91o3
9vlryDj5yf2JfCeAPhOstPKwapuY6Ds6fvwpicQUkvCFqp4/3ROWPqGqEAQIuiY8hqHlVcJLr/r0
pxwHENhFSw31C4K8sYminMwEFIRopQ7TI3d9BACysij1eU1xskfSOLfutt6E2UyZ4CqO+B1Uwv9y
0LRLLuZz7fUkQyodbSmobcYg9SS9ayQkG9JPxrQJi+qwXk4Gnp/YYH1doxJ5uTlRggi9Q2xnN/K0
9W3tY3p5y1v2oQYFnDMm59SXOkiGQw7hBRZ8DWS9cFAsSe/RaqJqYFNxwjp8socfhebnYKiP+qak
JIMvHFc1DmZ0ZxJLbvY69OY39x31aatDZ38wyacNinVZ6YYyuqFq07Pj7gmUV/8LQYleVvh4tRt6
xKqEPIQnNc9Zi4m8fMkXgRe8BkXjnSNPXOCW57ak8Vu731IwlLV16jBKjkKdOu9uhFQRreqWCu4S
FZUyTJpHfdGnPS4V4M4w/c4cpMZ6aauYkmgiVLFkvp+OMRYhuejsbLILkyxCpgGFBQpkUoUYLUGP
OH0ruXp6VGyZ5SJxlmQ86LpP6+xvkS5HhnW6FHFKjleZz88PvIdQu2DtpjGGuLZqOhb9GKBRCIei
re3LR2afattdVKU5HSlHArlg5pmdOoHNtKdArKDCTvL/K6YcMV2w3pyKK7I6I3BCTY6RAnQLa+6G
lOduFCAOMM9F6Gn0uopW2Cl4ZjmBAypimZuYG+ZQfeM2fROljXQhfD4XnYhbJXOMx8NG/pFs+tku
MLCGGYIcTAajoBjkqlt7HXbnJd3Xq9eecxqwfYwYreagAfZ4oYcuYk7HZlEEdhCGsu2/IR5TOXWi
Ge3FI5K6npYoKXPKDZJg50VEC9WXadqQOqmSPf4y9pq2dtcbGh+1luIIbeKHTrs59Llw0i1Kve4T
c/IY6F+C3ZM2fZ3Y9AMJQFT7nV6vLe8rgfqi9Z2JvSS6LKLYeWjKlr9ikz+VKENCFAIScyplIj2C
E3ZSlncdJMvuul0pZ229aebRXSRd8HohIblDBfu7X0mDSm8AabwyAu1WUBjBIV1bRPx6lhkCty4Q
h3/HOLyZlNUfxo172SPIYyI3I8BqZAKUucxIsZnmUEkMFvqV+Omf2HHYlf0CYNuRAB4NU9eELON6
WPWfX6Tp5hs24LvyRnqqXxvpKRAZYg39DDx7DpMzkIwqV7G25RqimdoBoR4WEREXWHaK+/pQbRfU
GxVe2ErDgQ+++7FhydoOXjRcs7Rgl/+p431K1QoIpSINAOcZJMuYkztPJ+MpfAoZbdHh4CGV7HDH
YSMgDdLaPOPAOPf1QPuIqRHeld2JdC5jLZuOJx1RxjrR5DPxOBFdwY4ryDdK3ITAWlqiMkqonDAx
AX7oYCO/tDZ9Wk5cCR+7y6PyD1bZL+m7iEB2OyXBTnSHUhrd1/M+Tgezk6MLrd+JQ/pFGyeHuc9x
zl0NfRj4IQSLcsQJG5FzyoyNjt+t3tIDATEcz4D8Y9roAS63+GNvcqhMSvwbbozZdVgWeQy+l7cW
LU/etB1UCBrifTm88BzfS729EmqJJgrUdSrrKkcdKHz0Z8KKRsBzlUBrZeDvYl5NOIeix88v9Qdm
chL8MxOoF/77Wy8H7ymeYLSG22+q+/rYGCTKLdY63jemzk3YbQHQT/FlHXhW7Bh1zGHLPM00MqDc
aNLUbbO+iIHsfYK+YPxqPlA5w/NgnjVTB4mB/RqbO5nsZrR2gm8aFMD71RLVielk/KCwrUVUasVT
7kqD5TubAOO5/sZlh5BIvrYBkHIPu7BfdGAyl+tCaygLUmCw+Ax0BNCuxYcvg3RIw8uYfzGoM5d/
faGHCXo9E8i5Tna9vRyxNNTNH9ZVmfqssTMsc+4PoONqKAbWC7tplkjHBT2phJna9n2p72WhWoAC
jP6Y8fjRW0wXycHqNDk0JOkalaI70IuPyDn5ckegL1qq7vlgtlJk/iT5JtonCfJCYlMLkvNnl0EH
OC+vWVxJrdnn5AzNm9NJabagMhx0UB1nP3BT6DDeYEp627JLBqAovnc32uFWzLgwkrj11stpPo6j
HOnxvvB+dStwJA3WJ1rbghqvXelj8glamCPqFXDCCROEOyv4O7Pj9hrr6uKDTnC/rMcOMyz/1R36
Hgv7RgAiyWzSUqQGNtaSZ47wekZeAsDHJYAypPnN9fhnmH0WXKgjsQldgILb42stOQfxKTfN2zxv
0OHlcQvRv4QE+XtUDUPfkAhLoepeZg6+t5eOFFx5vRvZhTAfsjVQ7MwRJtimlhaaWjgXpaIvAw3J
+dW2CV56pR6/BX4Q2xHXw5rIPeAYO9hwTemuuQl5wWEvRaRYoksf84eF75aYzGsF2GWk61KdoUIn
XNxcB+81XRusW4kl7dpI9LIFDT163IJehtyb6V7y4lIH1pOewXuBbW6wXsWwBG78WgzK4YnNNJGB
kBZeTOKQnCI0y/K4TUWLUUQt5hrZxB820SimB4xnuwjhqB/MyKgonYAxehiMipV2WpDyXfdMbrcq
4kRfbVFaokeBVVZauWAuXD+z3XJEikOkO1VKaMvSSI8JZ9ywVgNBw3UtM3SzktZjtZOakz4PZbdU
8G5DXPVt7VeQ8lZAnEN4zJILI/p/q3FiX0EzsOZd+X3MJpQYrLZGy8iM0+lqlCRMPnkCyPLDGyYO
CAIBvbmqQR1jOd4IkpLqm/Z0avodsTH1tJA5P09gIyRV8s2I7+SB9/SRs4fasYTHILk5gMZGMiEt
fPQm3Tg8FJVXxJ5kwrIUeXD52wbUvrTvhs/BL0pjRV/XQNFX0nveWUvlW3Jl7FzTH4vXq9R8vF2P
waOAIXo2Cd38T/315uqgnFnqeDazQMsGy1dSWaYggfmRUBZQoi8npeM5SUR/2UWdIqjdVh66i67B
xfQkb6kDNHwCWYl70kXbOaKJmU0AFn16f7BKQpoGU4Zvzn8epCpGDb2f+BwmZIGQCnMQWzkYFrSK
jjALF+yxHqPp3lNdx7ZZXBrhDFAAafrrBbDU+GtXUR1pAJ8jwUfw7J9AfiRr0MVEKvpQ/iZtLNG0
DpKulYrWU5UJe6CkbYzfY2gdklJohn9kJkcqTMiTqh1Gn6ksxbTPp3przlRL0BffQL7K119UD0O3
/037fyZdV9LufaZvV0//gwTFFEJ6S6rFXCL6hWOuQqSGAJM4PJQ8txHIgQbuGiGCLm8kWkCVALKf
/DwPzllOpNmRLM0Jir1OeE+41hiybtWrxEZ3S/B3xRmxCLADdHSwX0zgTgzOcZj2X/36gjzFMKEd
8PnIggB7+KG6Ku7KOWFzjd7zExluXEEckdr1nvUTXf6vTtZBmZNdxw5kymwwEZaQZ2ST02hJXb//
qbT8r80Hk2HdfK+B4N2d/MGaKgxmQEmwL+lDElSFmOShLNQw1XaCqnRqfNTO4MU/tfPw7Id0/iIH
8t2Q+yf05IHrg1uwX1Q2wdapUjDoFpszHRqKaaWkl67iZ9CaIcptoEZHkzbkvtu8miQiZMadPrrM
lMh1hTBxhbPiOl9is+byMXaJHielGmF7xqo5iKj8KeC5j0YAk5BqtutPHIYuoK60d77/s7PWyBz3
l+eZf5niDdkdUaYtN6TOkpQaFWSFZHFH45MLP/h1UXV+OYxF5OqpxpxAUM5ikrSH+K2vJQAfjzJ+
4ZEowWUPMYjV3+/dJEAA4kaGszrcQs8KoYYXwKjuan73PTPxcY/qDZMfbGZKX2BORj7UxLVu3FBz
6mf/et685EP4GTxVv0MVAaZmkuAHWMfBx9wUp6DUbMlKWJ67sw1e+F9XiiqYbuxS9npxXcLfHHTL
uxBvILRdcndoKueTg4wSvAeEmqxbt77F4QUjNmweljQqa0eIdbqVg60vV8BfF5VYnpAP/TIv4KRD
oVimxVl+t6VFfHaZfbAFXRaLqNtUBQahvICXIqqvo6XHAnVInkMulBF89mmVv2i1KyG73Hf+etrH
ylH69KtxnMzrKrYr1UO4EXn/PoxzlJbxM+zxL9Z07fVsZwi2+TcKT7rBNKaQJ4BEjRYM1mbAwQvW
WWaZ+6hr6RDOdyKhT0XIED7/0/0lky6q0WcbU7s+9i9/CKcowqWnu2KCGgC/ovQAtr9R9HrCgu0J
q/3vx2W78ZLEGHlSD8Mqv93loVJCxiuju4dqp5utJkiHGFa/DQ5wqL12o3epE6Ve2V5Ej7+moMf/
HtLNkaVS2S1YJcKI1sqQ17cbbQFc3jQuRym1LaF0prif56RcSxD1MGGNdg66fn+N5T8Zh+YpIlsL
Cx4RucKM7h8dbbiDQfE+/ZjTWVYiD6yO+z4GX7ZB2wXkazx4NWegevKtj5yO01UmBB4Q5TdCAPjF
YaFi0wRe8106GjdUsz9/QlMquluBFJvFz5qdekHxD/P1Um3L1SArAZ3qNvCwfY7uiTIob36/xebE
FWmX+yFKpPLgNg8q/ojwZLhA1TBtVYFkWjeNOmCoxT+WS79QkDMAdvexeJpnK4DnIE8Hr01eEWBc
zbt8u4Cy5jdAXztiTH9FXZdAUuoA0vZiDMW5OcuTqyChzalzRU2YzLPRjMS0eRxCoEzByCfPF4Gt
5VtTWULecwOnzchDzCCtz4Q7R7wwbe7LxCc23IjA5YgiZ6gq2qrTnq6EPuvsP2zUbezdOBlE4MYl
1xYw5HI4MjTq7DZKBdle5DXRLy6LTTPh0q9twho0KsC6KHKaTx+QBONFrzzJi8LKBu5XV95VwMLY
0MECONreMgZ92WbbZfz5+6vNRLKKzZfB2a9LP3VcS+6jPlHx6dFVYczzDBGMrVyqulLZ/XSFH3xB
44RX0PmoI+GH/7Ye6hPFGHaBDeTRwLSYOawveHNKAmEejrHhnLBBdj53vXkxCGtX+eY8OBufnGx6
z7tXLYrWmWilQVEampu5KyjGjH6fLeaqnz6FFx1R9xo9gkGXHVIYoJBg0jqAN5VrarK4FOSAW+g0
eLmSm+71ew3UGW2QDej04Qi9K4G0yVHxOGrXr0nJRI9LEKNut/oOEDsZTUhOFeM/SP8SsLNLpq6P
bh4qXVXZMxZFka7VHvfCKysY/K9ACs2EeRdUkFSaLUXRgF+4tfcAMg4zKcUbUPvpDVCX3loTNiZK
FzvanNyW7ADL7fDnGXF3V025r0qUBVHSDISsxh3V2hzhbmU8+YJVtqThHg7YyLNInyDb1NzMQQNU
msP8jf2n2Sflx8ewpQkmQJXVLNIxz5Dsnw7m+HyPNrDyU09C4O/WC9ntQnYRiuJjcS6r02amesC7
ERFiqcjiMcszBwQnZ1qetlDiGYD1cHCCTpaVQSvejOTNESWTQ4ipqGm3Mc4jl79acKzNk+0LY3BG
nVN1EHjy/NIbNKtNs3ZA1zGFTgSrxi0xll4CRdKlnbjJjbYeV0188WUkvjAyDjJ9GB5psOI8m7ig
H2sIIFEMwZd5i+UMs+Irx1Ma2LQNk53rgV5JBcdFudCbTSMfT585De5akOyrEeWPGZ77DSwOR3ud
LFwQMDXxjskg5Hln5YQoAIM7c3PKz3XlJCRpVt7un4XUNYnyxqbsvQElrutpqXcInIPzWhbgn8q7
00in8a+E9tNABSOg9hRgTiNNxFzqN25KpaQYUthBjWEe0oVRCPFLLe2bXpR4/B6KIEFonYhoKqOa
fpPAW6FEWeT2Skbf2IpBzUBggqD63Hp5ei+MPQiWzZc7s1CnXS+OZdnycDjmfOMvVpBfawMRm3aq
/7kYvAnSH/jn++RY4vjT3Bg4EORDCEcovGbQAglBBk7P/wHCt9iybkgtUTVVxnbxm1b5facLfgm2
dn5tc0jh7WNQGWpN6qIn545DZFMCvG3r7YLSZeKo3IC33vJhESXMFDcbBmFLtgC1Z92uH3Jyp+vj
S3MU8IIpByjOVwdS6eRaPk6qmud/kyvaslPhf8y6U21GdIOz/RgzyJGfrh0Ao79iWAABsJRu7EG3
6Spj4lRQGctR+ZacOEYrfsxQjvdbNhIZtVqMGBEHg3nED/cfg53kf1UXEwHOL5ENB9T2hVSiNf9h
kVqrzSRKf1lDsdreL0hdQHf+AU1mTmk/C71iSdBA2dfUlBjpG2uN9vIojEvkgaSd1+oKp+mfXO+M
Yj66J/oP+0smxoe5iT3dYEIDIHX3FKNR04IAaTZxssSuqeU+xPs8K/zDaIYzCj9CoqQ1vn/wyCGC
HnHNQ31SlrdaMoaS453gKcsGS48jiRhf3kIrMgBzbqTgg5LX2s8x2bCn7QZ1HMpbTLGMjsv4WmkO
4u5mk3er2JqEPiY4qxjGHGTzRgN4yZFHZsLIWed+Fc+BTK4AW06LGcLs/XAGMc/t2cXByq5NVRXs
Zg1PDvy889qY+1ZjUu57QjR9ceaVgZ+qcerqo+pF7qeQwGm6TTlVbRLy8WOLXTK8fs0pV3inAWw3
VN9ID0wCoLQ1BL9Y7ZU5z+WcIiNziWo82IsLZQSmSkm5o/gOqJjQvwOO6Zp2foCUN38bcpYzvGM3
d7FcIX62OGZNxFMpudQiD2mpgR9hV2bOWerc9IP5DtdU6Ug2kEoRh2vyjEHc7VZ8hI4+GjdtDPHC
1hazwd1414H6Up4OqKd2g+cWzFZZ2EMReymtF82XP7R1kqoxDQ5QZCPqvsG+hhM1VDvteHrdZ5au
nfdej0wCILNgPuMCzqO9voki7gWRxZiU1zRONPai5I8qSemFXXwGo5/2SmA4GoxC66y8kAq8QgO6
U6r/zcOrDOvmEfLhfheGiWnxkp2LNIqqDkEOf0+lOlPAg3IS5DN3FS4xypTQ4edVfiQ20FO9rYCD
yS6QoGOMyuNWpeoaeEXEkB4NtbIGVhLD/2ilcFwvFFyf96a3GjDkpukKH5syE+DoZAvwABQe5dDD
ZJgzq34iANNrLY3rS7zfdTGUEjgufJkenJHtyLrx6bCA0zr0D3kJMBZkuxURsuDwKDUQBFh+3Z1S
60B/JdTewWti5j+OH51lbFWEXSf6UtqCOOFr7j5nvDlCPjOEVK3RmldMt3La44O4kUuIoqo/X0Ke
AU0AIvB7TUQADYBobmVDShb+iZgSSmeN+QSQ933TMNLCHAs3LYTHxydLw5szGWlJsxrzjgpD0C61
fneqJ4MVL/B4S5mnamsTb2I3zTUbAnYnwOZqhcYnfobAxKfVw7KTtYQrnZdRrRPfeO4g8SdaHcC1
UD+nUTTKwTtKQ922KpsGFn7B0FHZDrG5hMU5NfL+gGj7v6qz23hMTKPiYU12ZOSkCVlOAZoH2fed
WS/kZHJNY0STWa80mcMpyOnMpOmCTRXSDnT2gDOYARZjJottfacjRAYuBbvoSmsxcaC+fx52yY+v
RELTvyeU0VQDCuTeQkYNmoI1yBPcTKYn9/W8vxTNNejFYTl7jlhZ3KVmbsYa1UuRJjy2Sujv2PE7
oR0uyi8IwQsU3cQU9b7cvwl6eAzktMBipeJrKavj7AWEcXMA+DVGvgvOUKAK5EfMU8HQyTaUiDT2
IkSIJcmAW1lzcCCEEzDwW3FrCCx75CuXq9P0gW3hutcB6Z1QTbJcLSdGNtzDo/sPmW4OdTtzWS+r
nMqw4mSLtuP/AdgnlUlAhjxy3k4sa2x3fKPB+aid8K3AJfIrvNhf3/hX0JcHeGFrIpB+GIxy7INT
Oh3qesdP1mb67MhtkF2L2ILAcyREeFfEKHl3wu2LyvzzP4V8eQT+vRBoMCxRktFiwNH4xpkUbaK7
/2DWH5CIGleQlEOkz83Af4XemE37W9cTh+MTKwGPniDEy0trpuCPrYq/KKW+EvtdA27ny3ftvSaZ
VIqL4E89cB7D10ZMfIjuYa/3B0QTFz90TZguxF/xw2O0/UHkhlRb9NMsnql5EL50AWFGpGjQCfKG
DwF4E0gFy3iafW7aUsdI1nmIke2phXLmKAq5RtL02JxhTidu0nkdYL2n2UqIN1dDpcwT8W/gAicp
vUH5ALwE9kUybywiO1vRltafF/J/SyZ8nIEI+QHWJgy/wHgtl6VTAQoO8BhHiqohA71g7AHX9UkD
bzIOR96p5ZUfzyed1aiaTvLQybU+YRFUUWlwCHxpz5U55TkdUMJq5RwHaEH3mhpCCPmJsr9P+Zm6
vOcwaBpP8mzy25aa02jNYqhG7qTIofRV8S0Nje0aO69BlLoRScJRbHVvKTRKvRrylF0GGKBDvmaY
CLKk9nns4SzzbyRQyQy5w56OUQi2HGwpYlVGo88fNFsDmjlLSe5/rbTDZg+8dt+N/scvqXrYstci
ImxnOu6J4+ca1THvMvjv8zv9MNdqX1sBh+wyda3h30xnPIreY1iLViB5M9fFljWWKPz9018fgR7T
w3hHUK0oGWYoyPqcJR3L52rOE+5C7By1PJKvW+RrwfJg9qtHzQjFOkdY71v5PkxXqjWhxThOnbrb
OiKSkks9wS45N8CBm6W91eJgXtzWsL4i8CjfPGDcWfDCK3FhSrbEw69HWPWDEaISubHAMz50hMP4
lYkCrF7BTqWOoq0E1mhHga+8/YVsu4QR7exTdoMeJswyMdRGHC47LuZST87ySIIhc0QEDPr+SntW
25WyByqapU8sy5NCt+t0drmgqDoSItZSqDRxHg8gYwTrwWUOpshfxnKAS7sFA4fvyk4EwVn2qEGc
Dt10goV3kfBmIz8YLTPlldyCXBNz5jH8GaR7Uh1dKLAaVNxniCRsvo1N7Oi4pSXyoELHj/AhImQu
Qo4wAsGTUsFUEFxKTCi2l3dkRQSUyzq5f9gqIjlEPuRQfUxwQKkWU8JO1Lj9gEbu3BJVPgy0zu1I
6S74Yl5dUoiuuAs26XgGnFf80OoUSJzmGhdcOgFHj//ok9SqJ5CVqlMlRe7S5hOj+t/VgAtHSgvM
r742qkgWBnl4skXiJqyWgUHdoSQx8qI1P2BAXDFbiSAx0lGvXLjBkBUa+YSrCjsGalg9ybNVzmH/
dEOtufURlUIPSYglNobNlKp6Y3qXw+bgc1U230ZQ8Ocb+n+fZR7h1E0zYDBIHBuf2ODEMC40mLKK
jMJNJOm+jzFwgM96zHTej2r3JsyVx5xze1nSGoL2qUq3ECOVaL/ocxvMYkLt2Cy3ztbhRugdrIoU
WxvwbZ7dd1svZ5wtYqiCgwd9T6EGuUiv2+iRxFq/Y5fxQiUgCyL3ecn16Zu9NN/OzuCAzjb0n0IU
+wbwqQLK0UypHnMCVFZdvGGTGBtlFiVj+I5C/wUeFj2MWYcFGTk/1+8MTDSvfp1lWwkEdgtrRKq0
Yy9ou5WrxsbyXGoRXkDfVmBmfxh4k7N4ZRSRuw2j5l3bgTXw3NYFjdqa5zNhr3MgXgikGGPCk/6U
W8njHbEkioPrUS4B+qvTm2Ht1kA2+9sIay5whkeGNwcUo9XdocWgzaS5P3RW/WUE8TsBm8GOeb14
JNrP3U44Tcos7y2QXaCIIgCdCm1kYVkhGRf2/4fW6I5F5NKuLrvrFe05MjPVfH4kg0Y8R+XRQ/vh
YJqmg9gGwYZyxQDKli5aEUUcCl6MJLDR3VBGtNTToa33mWif0C2rGGkzkVJrC/d2b08+V/Joszm3
HToGJ57oAeEA686bTWJqRD79xXOf+QSv3kXJIOSg/a61Nt9CNJ8DFNpPCMREMKMQx5JzkPGPuxc2
sYxZz/jfP0WJRao4pUjrKwVY0IQj1f/w2rCC+BlKE/HWpSAn5rW6vnSrjBlW7BL7uH3z34UMqPFa
vsK8EdojrORu3m1kFAMjLlvGSINeKdA2sotgXy7rMedUM5fY9BpGpKg77pZYVbNedkP1rZLY6vRY
/zz1klrGIB5NkCip27e1Dn9DPWSBGwoZzFIV7I/E9UBg50i/DZrfDtIFBNHiDS8YR3xC04LoOfwf
x3UvPMMMs6FAsO1ALtVO1Jzhy7/msiB88UmeODaDZvDWvZqRNWvEZMMYX3+OOt142+J8clgImwNY
xKkUcxN3M2wZzFGJa62WNzKCAmb9xjefuBuzIpsHimzEDHTpDXFCJxec6CZodnXxhWArhr4g/75x
H7jANZR8hE9owqkwWkl7U456BPr/fVY3hYERACiwSZVkRTJcz/RJ8B3QG9W7LbhZ3vn+JndpiJCT
dr42rzPDhJfKMfTrc3nv/XiaRtc3FJIfPAEwxwJCaDKti+mxSPKZnfnaRAWK1RrWk7eprN3UqFxt
ZGeLp3G9yz8it4JTYBh/PsEZHZ+77Ozf61exSNgeH9+U6pMZYCbTGQ8wlvQruiz0baIcH+KTeTfF
8uJ9WUxZ3usbkVND8Tqus1eT9M8je1DouCkN1+TJTCRAgpESJUbnsOVoWzc7Et0R7IhsKUcCRQ8+
MlcWdefs3bkbERBvaj6Gbsy8hfvKA7UhJBg3+zWf7izHo1ln7oIsx5WAbf+ijVvcx8sKIpUaUJim
/EvTO+3/VPMP2NICeW5Tbdugtqh7uorjoeC7T/utFgCqgSdzZLxSUUS0y9xKnWBdlFk3HNiyQYz+
RMpaqpFDAyuO4y8jsMn2XGrLCrdD3lGyqZpLUazVXWTHkdRBBeOSwTC0LRB5MRR6B3MrXgLeLMsa
MIEqvoB5qKye1eZq0byOABzimDA1YDUSUjxzoUx9cxBCiTW3d2dtBd14waRCAuMdvdW0npCW8el8
qeTZX/5r20mOTrTXPWc+dim13sU/I9ms9tNAIUFRIkZaAxaT8ugXHJmt9YhqDIcVYHlsf1V7zSjV
4lGauzDqDXhXPbPJQcFTKCr2dH11H/zOYCZ8NF9SpptYaKSkTFD71GAacB3VoKtOLbykX3SDhlV0
de7NaklIr1PtyL+2IIoGv4C6J8uV2nYeA18STI2zLMnRe8RLyQVR7AoGkj+tuwI4OiAJzjWmt8xJ
Eq9ImYtjFT8hrwMkPdJmp0xBUK4goBtkeECZQtBqGSc7s2VVfiEvLzpDksCp8C/PgNccF5m4L7uF
Ydvmkl++eWBRjqo/K8RPTvf5kJE+2lwfVWBcn2HBPfPO48tYxaf4V+Cn90EzFExCjQWy3aIdwUxS
3yn6c24XyKskZzpjNSLhEtih5wuQdLElRefsRNwRM3aHVKQ03q13zrK9B3H3EKWP4jvKmMjPO6ld
zh9Da3mQFZD/EDJv2ux0E8xSYrJytSMLGe3ihLJp+8qriiYpn756klajYmrCi5LoT9pUvZzgTIy6
fsMFT7bGCp6yqBbGS3nQbFtf+syXNjNGwFs2eUZL7HAY4DdVub5fz5kVM1rBgX8fWxlLOD3eeqff
mQQNrhzdR7lWWMFngPT+XF0zhIPB87CLfwG6Z6d5giriHGGwmYhkq6IB+zMxVl+bT+7g1aYMtlMa
VShNQ9S4PQhzwHNtN0mv2LlEE97xq+TL1vwrKgaGaGfsRREleEd8V2w/fmEI1+CWpNWWIezltFFj
ZQ5UtushzRbOXhnGs03SrRoDMy4HtmGCYhOsdjpLMBmCwS+NwXLdYwks3sZE4Kitieyl6DIYHzmq
0Eed5DBdqVpOPFq8krHGQTUncF+v58aeSLH1JU9u0v+P+4Cw3IU8i81yCZJSq5lb+80T8br2awkr
tCs/tzGe5XhzE9zS+Yco0+kkT5GZBui38+Mcp4orEHZlRLV96cIqVTgJxUMdc4rIYM1hhlrNGyKs
B4DiudxTwf+LXNy892r70s45XphqNTJtarn/fgPjBGFNVhAnui8m1O0NuORHW+1BVrX7PrViA8Ex
J8723VAgTIifawjn+HOBBpYq2HC73nHeOiQS5z7t4mC4PabCYNHDVr4CB11O1na7ANYFFC5iTuXv
0Y+spVnw38dw/3EI2MU+zq+Fype6tEzTOYJLrPFQTF0iQzrwjqx0YjK+qxUJ+6WgTj4PZBf1VxVZ
u2CzFvxdcPTv9W76RguGufEYV/rMtsAZPJFWxeDz5xz9Kq0GEgbJVyMzSZCmBwixEIATO7JekgVh
lCIZkrkyFj3xdV5NicC9nj5zk1HvSsa5mnPHeeCSJqLE91zcbXC+DZFzv6uU3CJMMWGScWEadXQc
Ebqljn7rmtWXIidhsgaDkmlezJLjCA2GJyOcwRng8bLuOsV8ZXDAw9y28FLbMkJJRul8Zit2oHKF
GpKa6NhMYE3BIlUlhsBkRoOj/jiVj/GYsi4KO/dz5ejCH594ONu60jFZjSv7Gk1DYFWBZOCfwYVb
hGd8ExQJAygtWn2EidwQhIjQK0KVmSwK9aVfT3a7Hy48EmOg8PmCiBfumin2u5mU0raYV60X1ZbI
v5IjjwdCzV+4A9DkXENoaYTqaqEpeag4Ja89hDX5M0W39GZHr2bv7w3FYdklZOGQheQZelkesEWa
dwabZj1Ci2Enpe4IopfVcTLH1LjFyckt91Ll2kyReXp1Nst59kWUSv7oylYmwD6cp10N/jDA3OxB
beLgNiU1u2eQwqETBfg5A8FPCZ+LowMmKexKrN601QD4hQ1aY904WwNcehYgmuaVIHrtZirOnS73
iIq7mz93mHlTO+DX9mdXJrJrRr3M6OSqajUKnjlqPEURlckps9lXxuqoQvjTSjaFX/PcxNCsj+PY
hjcgHcxoGRTPzADEk4i4FU4phpyWZrHs7UZ++oXshpcKIVD5t/fPisLYcAohQgFAfya4KSe5VvBy
DmaSDg5kS5LUQCxmqaDzcs3kp3qpgx7V4SewGQEX0u5GmGY6HsRsrzoLyspTulGrUT3n2jd7+Zbp
kjdOZXeSs6jxIFNgz11wAZxmQoSMmZJlrRsYRVoVLknyJtyIfyp46FGoliZwKrC7h3i3u3ZsPBa/
hMPnY+DRc1PHn+uSkFJQlQfPHTKtX5Ya8j4u2bBQ4l+91i81DURT+ab2VQG21PyaoGmItsgd8Avy
NCdKRi/YgmiaISpn9JoXebH655Hss+BGHB1osVp5w/yteuq9Nj/ofwozN9wndtYGC4hy3UzodW+5
NvivUsEn8DkKadW2XBfFPI5qC9KKf22K7AYN4xCcKn9xWidBDaONLjEYFax/5qrSbqUkJNufXiGB
BQ4FuSz7nPc5COmayqxC6mvkTK/h4jMZPyMkrUm7GkDl0IqR98MgAQBw3vLi/WGECYmCkbgLOXdt
HYEMqhiY9xOT9R+UKjo60WHQ3Aq75E6PWVqeULIkrz0Nf+vys2+akRLgkcBXPm+IqNBHmhCphPbM
46tjojp4mzMplxPVNTosfS2rKmd15iujijGLDALW/Y6ysX+NxWEN4xPgG1QfurRaXEcbsqR8EdTR
UQ+KOMN5JXfMqfOP25WUhuSDQgldyEql21oK6R5qVDUqtEwJSphhhmlRixuCU6Ok4E1+hIfRpLfd
uaqB8WqfnVVPKl47TpB2ipRwRFCDljxfQpcRCQWxnfhwCqfuD+1QlfrSK79XXS0X+r8bB1o0j3Uv
3nLm+fPrtAArgwnXq+YEEF+uUrYjwj24JwBzblnmh2XqiXacUIpXMB9xzzWSCcXdWL7Sc0s6m1y2
8L31cPLfqMW4Ywgtaw579nxTSDZKdrv8w7RIMhK2/zWrnrA5xu/FCJroZ6u94TRLNv4+/rjvFpUD
10RdtAX9N4muyF0PrHkBTv34VL3JreAeFWuBQ+zU3/54uQgG2pCluvUuGAcbR9gzRrkegGeMba6a
FBer5/FkADzM/KD9Gio4455wqt1nH+9SZlEuznbJrQXFjUfLOVzsWvaoSfq54iP0OjqoccOaOtRs
cjKgtiDZcSuR89s+Pj/R6gEF67e0xqgKcauhaXyHKIBKlJ4ThtWx9OidKZd5IAQu1GCOwuBF5bnP
6jNMdrnjLACwXysOj2UHVc5BeRzuzNSaHDj4n8m9zamrcn1FZzx3CgcqTgTS62cr5u8Ol/ME3CaW
leTBYVqmLMLOGDQibs5xAzppVlPo3+uaVVbnsr1LIfu6pQQvELkJSHmYj9Ht73agGK/dMiE7XOEW
JlGMwY1VtlYx3oO02ADNiRnRI50dAHxOCGqOfEA3+qU1w/fsu97KbPfhbmkUZDj9CGZoo+ATdem3
+swpGXH+iryDDAxHEEhBWshrJD4QLC6wcwspzky51+UPB4oS2miTDuqhkJMHjbSSeBQBB1EW+6S4
sYeP4m8Gi2yw/8qTUKFmZE7Tm8AphswMVlCoWZjfcsQP/uuymnd8Ygbc6JvDVQk0+LJ5cXPyQ/TX
nmwm6kBTk2SsBWqwwzMFDWb6HAOHkFAdXMMFRIwiT+j170GQd4qgE4wITjcS9WEt2Tf5fjHyJuQ1
KMNru9WaYdyVULlOQaK83l6aF2XK4+agGrTcdFMsf+7WGl9jb78afJOcycZaUFu0Kr8NJO7OvRHa
XbJnAffb1tK/r+SCgerzmmR/WLCmToLmGLM39v2oNvG0g5xJQnD5je8G7G3RB543o4tRHoIs22NM
SeWRq4zel5xF9NA8oNIkqTVxBDMnWu+G4NQMqpPcsUXX6PNqjManlSijGP6tRDFYCG07sdB+ip2S
7DlIYeSQECdRi90lGcaCB0ZRmpJfpXb45sEPeLVkQqUY2ruCe0ZNb3ZZNwufWYn/VmFCKGTaEyg6
uaojbVlJMEOwFJj5a3uReizTnDweFF4jQdaPDNpaSe4gzKwnhUxxq4kuR+gOmHICFGoBEMc8hb2B
sVUTGyXvvSbT+m8kGVPD+G8xYjd61qnR4ywfukLZ/ddjl8M0f6oaLWCDwvox/zY7P+r24ArOMoqy
JJ4i4ElpOPyuCtPvZMf9K6MTXvSjWvYAH4rgNJ4yJhM9Gr2ovdaraF7fBURvczOpaTRybmhTFcHJ
DGVzoM/rHypXGX6U8rLcmswolMdUY8JqMfXpuumclcEiT081HRNHVSF/URkTGR5TFVRuwcWbStr2
EyyUJaxWkLN+Ij9KCKEPKv83NoZTbVkpWYlj1fPONp+u5cnwtZe2Xw7pTplPnJ0cA9mj+6p/djOi
7ymBEUXRhap9yyggjp3RT9ZXRnAq6NA2TuxB0PCz6VhfwozGwF21JvEqS8PzRkPJAQXOjA1QgQmm
0DuXUhCLDiQuyUV83O2iKxOgnxNYeRaeVPMmO3dFAC/0cLkKk6cUDjuTVLq1x/0yeZTjlHTVOlUN
yip7ywcISN9MBq3JO9ndjJeyXxz3xLrj2VZxo/JFNZueUY2Ta4J9XLsk+kO4Y5NVBV1GYhs2jrLH
8i8HhPqJhWJQ/7td16Rr9WJIDMqHuo8PpsxGzT2bLEx51sndRx42fWlaDmxViE33wn0/YVsp2P6X
fqWAljh4uMX29MB7QDPPZf7KWpTCp8YM67VuSss6BIzhgb/e4GY1frkx3A6SG5eVXhUE0osCg6oo
wjmL2k1ZJ/6UmwTXVzTykAAkLow53denFyw8h1Jg5aO5tfBIPJLbyuv3VkOaj7Q+UW41qfds9CUe
COA8mScfFTNXO1XL1kP1DOZlcF97R2ndkMMb3C/X+RYT2LLucURh0Ildk7OKJabeiXitzOBbCwJ7
8CJAEFhZ1H4JljnLGzK6RuV8kCcks72j8VyusNd1NpjeuTicTMF73aM8mtdMaxAeVVQcjXPFnl6X
tENi1Zh/xkL3mcWrQ3f825ERFM81M2Mkoll7LfhrTc7UIpflePPXtPS66gtyu+GOvUXYgm/XRWuq
mg0Fx1cxLTaiMz6MIU4ngSsRbBEsThptkaTkYqEmUzrXR8x2DuGnh7z5mHg6MtJgUr2o8uMaH+1y
YVsh8l0FXoZpOIX5DDd57iryHxk+ptG7Bg+hRF9roz5FMKHXaehDoI8/2/yPV5GLjoohXUNoPFy1
Bk9VOMqIGye24ijNXozLoV4vACFSN+cfq+48YOO0Oiqk/vzZ+FLKu6JPmjwPApxh8X757HQpEIg5
uHImsF/vDhxX45Y0a8lroxBQ4q3MGRZVPi9r7IICvays6Opb9yq6iTpNU9FbJ30sU7knLfsrjyMi
+Sr8VelL9+8qDAIUmQCRdXmXLwZsUI1zKyd087CLVJH+zV8A6t0K6dssuM5tdffAeEvUqBmC05F5
sZbeOlMg4Qnr/3UHoIcnGlab2TYq/Jr1WOjgTfm5uco+z24HzO9118Ck6YTXqpomLAA+2jL/v6x/
y3zM42MXC42r5GeAbka+owI7bVoZZQ0rEePg+R/PV6cGoO3ZV9S23jKRHK6NZsgPrtqzzRO5NMgn
jR4irwtNj/s20Ix8gsEUqn2Vld/LaLWjhlRnL+ZpIg7tRwwM8IycQG4R1z1YSQbW/jxDr2vQhoU6
PG0diKXXU2InYfc2wYvLAVBCeqqEn4wK21UC10kW8ITnCrKiu1NLS7iqyv5CBah6lHXB3Z39Jewk
buwo5rtqyc3yVxch4xkqzzuyw/snWwCJeEL8HFBTDLwgU1B1nHwoLYDET29VSfxJTuhbd4FC31KN
UD2uPGmHmDwcCInnnxonz127v7kzZKw8lRXEABsatEvDlH9ixqjq0LUNDx0WpH9QTbdhyd2yVnB2
l+iQ9IyE3yYq71ubYq9XwmdConA3JtLI/5yxTAixpuK2e36FYumyL+Vy/dxSFkUPjhK6hrVaBaiJ
Omq3NK1kCZFqG+fOfWbV5QEgnzIiVp6AcRdatUfx6j7MBtpsVINXfleH9IorwX67NmRVTz4i/3tj
r1cxp9R/4tbJNibK77Ig+9qjMUeaVNr9EIFmfvDMw+qDY629TdL0h1/+lcSQfbxBiGKVjJdYdlxm
rd0m7fyxqMUnD8kTQCXhymkOkHQgjLMbVwzLPjQRbEMxPP3hRdScQ/TrQiOE3AyFqz7S3RkASs7P
MNYQHhBDTBMHAn18sxPB+cAagzBjQT0HvSI9woW4sZn/vN92Sw5dGYanZLj7dyXN7kdte8fXPtTD
mnluRsS100VG+p4nCWRHuVTLSrnPilDeaGPToahejVLlOiUBlagyF4cfrBzu0PuLQ/sjA5xFF1ks
6QsMdqrxVz3YoR81MetSx4y2UWxuvYfsWGzPHc2pSUpKzDmtkfsRnG6xSun5okM6/3tC4WzJCS0d
QEB9gvXbMl5igxCzrYgeRCeVyGw4uZdK5ZmRaVflpy4u+IxnoruQ7nXUpNJFuuXmvk8tsvKTDee0
7iIrf7FQI3FVfnEP/ifKRDeSMZTI4NvV9RY162GwSZbUFYd4KJunfcnjT1WvaWY1avlkCn1IwlSk
5pfCTq5DFR4bj1GT+DzV4N+2m6YsZt571J5MJ58vpsxW9VGxSwwYLxq6QBCC5FlVYsRE0VqRsB1K
SChEpdG/atzsrG4Gg4D1SmXf0S8jaAFd0+ok0SmPvHutijQKzPjzjSKyppAqaLCktp5FxFA+EQ5y
d/75vmBLdM5WsUdGz9gybFeLmkOkCsumBLevv/zrhEZcrvK+jmJepK7WnV8BNqOzT8xx5km5tLvY
UTkfdYax38AqCQG/pL5vu5X3jrLrZXzDaYIY5WX6pp3Rdj0KJUGynSEk2dSAJ1Smx/UMVKh5uf5r
vJ+Y0qeT+qCrPYFpGHnL3rqvXQhlXXE8MQ5gfrHU/kT+/uLw03JiugqxOfPvGjR34ubWCMx1YENr
8EprSXRI/CIuwgQioOd2pp6gxAkJoirRcy3TjGREubyrdwDSUwcJ6/AHjHPvVSBRuNC2AR3SLw6C
2Bkf8yT0Jo6H2AE2PlgkrIFO8yMWJTto5E0xnwmSbYKiOK4NwBo2Hd4e1Uo3wHuKmgJdOKG0tWFj
xB3DkXZuTLlADRCbJgUbzxZF7cYuRAGHDMYIAQHwzX4+UIYqAgN7lwyBawK71lnbe8hKuVwD16iC
4Cz5VaYbWnQN6t6ES5zneOIPXVUHCHTlHc/avqtLarxLTpR8oqkgBuToVAdwiV48Xlxary4DQDYR
hkvmj4RNjvzI7I4JhLyDRh9uzHXYYcGHVxEt4YTylmJ/sbWPXZ0p2QX7DjdKXTYLCIWK/uS3jix5
5S/BGKsjVBNvhVQgQGABSPwuegdTUotURbP4P/XsTHU+SR1266SvAhmTwrMvw9LVsJLPnDExn3To
FBHICIQNJrZmi+zKpPwiq1qbgAxJJxEe2/zZNgCyctTMZ0MsEDqF6AK/k17vjGvMXft9ZmxZItdL
PbssRwrpIUhB3cqWV+7QYMdJHP1VOoayP77RWEco7JXcFAzH0Zjzk8oN2LMl3rwUo9Ugfm0u5Lia
kgdO2AGIgqQrHOhiGfdTqxEr9m/CLhmdzsls/7Bm1OS5DJYeTRhN/3b9Q0AYKlLNj6e4GRV3PrTX
fRgry3KaEDn6az/Xk5gBq6YpHFEraqbC2aotPVkJlxcLa3S3DHpuo3oe5ewPa4OeP5nZPL2TGZkk
o8rmxPxiKPHTuq8hjA3A+fhh7EmZrbZ5MUzJ88REVp6V9ESjz3hIj+h1/DTNbql+aHntlv9e16bS
jTmhTUkVH+Dn+CgCCub9p37lQKgiKm9Z7Tv3L7koi2QFXHMcyCE/+kv96xl5KmDupJCQ3extaT9J
SFVyDXoIKhGnysDoEWjpWQWtMKkQEIJ1maXFeFhWel90okOYvWqdbJBUjhDAZu6QyMbOYbDvJA+1
Hz3CJxB0u7KSwCA6vyZB84X5ocWBYklGgCucW8tcWabfZBxEUXDp9sMQOUoWULWgaqaefk3jTkdE
3VPo3zgO4dvY6wLJjB4mCVEMWN/pkXRLp1PUM4zDDb83xVb5AtqDZ6B9lYcA2mGlFYjFh+DWRb1I
f3KMkUVdxdRfn9Qd1t0J53oH+CAw43TIU+XlbWD+KhZGaHvYZmDOQpE38QXO+JWzeHj2qOopbXtd
f62rxTQB7YU7ucAp/VrU9NkIeLD8WqvlRUsOxLNaQVKManK+K7VncZCJtb1cDLgkfG5qOXK6hqXG
2bECDGj3XjueeUW1qWUc2bgTlYO+52FPnzfjrq6ZQgObg2JD8iUVsMeRpjVxcZwPHQYox3Z9+Xj0
HLLHry3sBpoXu5KTUELdzBELkpMuotfEFNk3aJzj+ty16M8SxYDtksv2slsX9OAnzzwMeM7uZTPS
AACmW4pz9ycJIBd7o30vSV+OEyB/eR6diOxjxxGbkpCqY8eLED9DFO8YQMXiVfY9iSbU/LGq8qMR
YKCxJX6JiXDEWqMI/IjLuxbuR3j75xRDQ1gmiFiIcuLximOVlDj7LoxMvzZZjuHlyJ7U2ca1NLns
KDdlJ6kHVl+Dh0RzbLW23qRu4zj6wJyA34H8suIe2h0RXhVAjQh8M/W5IDla22eT3Lnn3nGyn962
EarquGryZrQSOqhpDFvvLkWKqxoU2zFU0bjlTCzkMlnG+y1Bb0bZKBH/hyxc6joCWDZWL+5TGmbk
5QKlf199WTs6Cc96oxTrztyiZpLlDuuu4YJ/CldM2YDvHtYNF/mfVBnSBM1TN5yaucxSddsYe8cX
4By2lg/28hCaa2LpaUysUseGptSIJDzyVF+ry1zeiHcKoReB4atjdkd2NNDm5kTwdt3h9qfD9Vl6
GlAbRsZFVEy+8W3osnMdToZOuRQPTvN03OiADWHkykUhuFiooV39cVz0ONPpCaMYK6IcXLmtlY30
SvGEMF6TX8CMUGsjAkrn/6Txn4UdHOul3S15J/i78sZLqmeuFsER7HpmtcOChMWNGP/hlmWKkmvL
ex+5wsCLayAQ5PyoYBrOkYsWLWisjpXf7djn7jP0tb5yZK8si4iKGhKfVDlLEj8RmVAVVk+4Ai0x
ealCKpwanQVg6LZzU7rO4aCO6Hr/o2WvE28TO1qRZGmC10LtaBIrq1azzPnKLDIskGDQRMi7bOXH
vE4PdoCYg8gkmeuTf2rSG4N7L5jY4XFakse1Qo/WaFH8D7oD9x/Cpz2zZv1xLtE8spteRTu136hb
aqjbNMZT80lRliUNi79+a/Ew5DLbm/odeofIn04wj0q3KGke7pZ3NxQwsgN2QpI0FiBWRbLNntc2
8/c6NTn4+/91GWwf7uxTdxl2S5WQvN6H0qdIBl5HQAUEC1aFwAW2R7XVgb6v59Mug178buFwPyI0
6WxBvMcYvI6wmoyrl5jlmvJP7Api3YwLPOLtEYzJoQyevWTO6pY9pT0yi+QZM/iYlLb+3ADYbspY
ymjRYqWvI13M8sBfsJPVLi5ccUWyOC59Sp1FgEan7J7Zl0JcVoyNBPcC2Dx2fwOx8zAkjB9nEfwg
K8CAVFBvftej0nuyMDf58cjstHud92fibnvWI6hKsaxZ/Kh6gSWnylwRXGdWji/bzCiM4zEbnOmp
dD9/fZE0UhuDkdAf37WjhMR7gLPL3uZFEB0Tri/qs/ouQOOs4vCZ6VNJui1Lbz8/rMD0JHa1oDU4
4lC3pSyUe7o/RioENXUbUyLyBYLe7x/6PpQwEa98RKBl7mZbnTQ6ACVog9NpV2Z9c8QwjdHvBDEV
aZFq+aNAxREGFOv4sLRS4vCBwbM5EZMulyS8sKQzxcG2AXL5DwkeYUMd+Mwz0ezwFArKckXwFG1v
pshdpO26OWsVVIvwge2Ee4DMvGNbXxlvaJdD32ru8RRXJPNzkVy7x8I/eqTSgkTjMhCGT3PUB/hR
XYqPjewbzQ4KzRjjW0aLTvyxTQT3QtWfFxRibnXuj/aeK94ccysmZyD30B2LKWGTrJ6RAY6XLTJN
R6qg2ZsdB0WUAjtp3iKWzkg1JK1sT9lzkiMC3T2i3vECEpR0MqKtfkhyKkYxkQwMKlmc2/dGnHcI
z5wNMGMa6QvIEWo+tpbhncx40lWaTxi3qieeVmnzltaoqeM3VmIeMYWtUWg2WQtp/agopvZoDaUc
171K3gLZm2G6hcw/Y8i9ogK1zJ3YrIGLsE8Ggu4xthhY3YHh9/eGi1HEI7ZzSWKe1omZ15/Cytft
/YDoV7+z658xbJhqX3+VEbJy0MleiZUgfWzVHm1s0ofTeRRfqtN4JbZaDxfrnstzvLXm1Zvrz/Sj
spzoI59yJ5im6O+AmEQjzSxm5NkpdPPk+1rRNXbEVcvyggr3dQYV/IGoofo7UfED0QmTiKKR3ALv
Ra4jLgmu3sGCxVZnMmLYpDENJ6wR27wuirRa20pzxS/mcIrQzNY4WSz9S4JOokoO8F4aD8vt5TNR
B1DWhOLDajBAPv9riie8fy9uCNoLOt7wiXT5LXFSVpGQCkKDbJQ34jfsmVnZseeKJ87svTWkHFNu
+uLJRVVcuKnYq7r157ZmIq2MeM7f7vgC988Bb1mhUW8RIsnlm81TOjJVvKoINUnPOGykPXETzB8Y
/AwLu2bHMtDnF8nXI1isZ5kd+eEINqowt1yq87VnTpxnYCq1N0cA3TavqNjrXLHH8rpb9B+2EU3i
uDsE5ENWnDCzpno7bXaNRATp95d9lzeHLdblcHgu0JpLLE8gN8F4lH5r0xRnQv6kXlrlbSDG5ocO
O4BXFYvL/igPSWzZp/3kyFm4H0muE5psEjuhbLPuOmns/2tdYvY9pPWgay86piJP+6UBpsrDfShL
pwS1JL4hI315c6AZGl1SZSpB+oIhM9bZ4T+y4hiEr9l6yauzt9IlAL4N4IBED0AVrdyhkueXdVIA
geASguadHRhscCAThki1B0olgvC1pLJu+HRPIBfa4AA/8TqMafvKVgKw7kUZih8re/qC0/KpeAfp
qgr0kCt3odvrsKhqpwgLE3WXwwfwHlq5N0LNUOH7Rp6PFBDIo0Oc6wp/ErcM7gM1SClhQWD+LXoF
1B2p+6q+qtvqahu+svYPz6RxgiyZal94jhE9Da4AfVly4RNmyLjuVTGmSEoudums9Qk/jkrYIaEp
WJInUn0gHQMcRCOkzUGPhedNChOq//c7BZprvcGRlx5+ThkpjCLEOfJiZyWtrnpOy/VPdSeVAdr1
apnkmhAgifflre/pSnX7n9DIuNeihd5Up1YBbOczbYTlfTewSHsLA0C6GmXSFzuOksQPOZVjdhAB
Io+UyonIr1AvhKl6FOyLPaNCpUNIdrTjftM2siYes5oH/RETVnDkuvJ0VYnfePnGEchqaMgQWQvL
y9AgutRtyjDW6+rQGGmMRuM+FEiK75O0ER7obDe3+Q0mfEU8SI6Aj6fxeTy/yVr0bLflH03DopZs
GqxM+NNj5/oSw977yjhgDPEW3fI5lnEZYgAtAAT5f/DKSHfZOQBYffippJvcrGOOcTXbmWsdKnw1
VxrLuLd+Xohf6Tm3tXddwu2G4sgGQDeplIexGu3MdnEIbAMeSISb17HTL+HyGnUZgIJTGermIM2y
0lGyGBfRsrrSEK8nslBwDuiQb+83RniHeX1y2XVIV2Cxv3xegBfJWO/afA7WUz0Abu5AZ0uC9sv+
Bq2XU1VRsB5YDhQ6it8shZFDKHrN0g/03XAgSij3i4v3evZzrdoYlpso0kTP8o26qPs/RAuRmnFv
Qd5eBjOWItggBbP6Vq2wvyrv6XTMvlMujY6+B51rX8YuNkw0Z+xUYG2+ZSGTb6CkL6goBBFL70aL
TPelQQGpXWrvwQ+op0PtEYYTt49iNK3ASjipnC3fT0O2TvHJHo90LKYaW4cRhTMuDlwN88oVJfAU
4GuefN1A7HEU0MC7H6YKKM7I+ESrfPd7wAW0+qaYz97MQ+SRLSEIMAal+kWJB1n0UKc8RD7OoJv4
ozvk/3ruQaSGgP5rj0uIpjcFGk0tGcYS5ZuCg7mXZkiUud+ZvXDLRgz6RtayuX6aM4mp1rgDePW0
kWA6BQHTxT8XVn8zOb0XsVxoxrot7HronHjxBXgLLG4Ykb5mn4U2Z2Vncuqoc8Hxrlu45FFD4yGF
MEQs+U6M77D45FUFAZJRfCc4hwlHf2Q6d18clkxMdv4CY/WL+PRSkYBVFfcKbAMQZJYuwFIIOtz5
WWWsJuzKdEl1zuBGAIF3VNAmDly8m13GoNjb69GrBNOREc5Bx5YSasjoxk6yu1eHU0o3M0Pl7Iiy
zpC1obOwiMHjsJaIZqx08062lJ6zQV+8LW5DAq1/ubI9S3hla2WNhSEVP6jbR3ervctIieA5YR6I
OsqlKrA4DVpweSJyJ4tPZAGqnAARdO0Du3tUCbf2jKa9NW+L6QKjAPjM5d5RsCZIcRwr0cA2TkJp
Pu0sQpj2vDMDeTcxNdUd1ZDGQ3vdTLyS6MkVD3NGGPPLrP8aSDGUqP6ZEpB+x7NRhNR8qfCcIbUV
+vfeWkhKlE4Bl0XMlAELrPB1SBg//dH1n1YC9JAcRPypOTn+vHOi+hczI7qcndreMQe42aKdABEM
x/oG7jK70AEA0U99OY96KaleuUHZa25ng+KKWIkKz9rCdxbNcQkpX4ED8tkJslSx++Yme76NkFix
9M/j/jkAtAfMirk0RZQdTZvkrJUdC1ASc+NR7muLS5/YwVeVYsKhmjlfgaOGXctrrbDNwg9M0dP5
5wYcfjKhIqm7X5vhNCeDzw4O/fX/rUuGuwnV5KhyQyfCTyvIXTF78/nTmuRIxDaEWvm6PZbMStto
EN4oor6u6tYLczZN4SsRQ9Xk11tCAL+xlkIb/hsAuWdmuM46PaadNNrofPKbC7EzPKrFOzcd4v/V
HRStVLHkGf/hNoe9DJmJnt0KJctUrJ4mroNBzrOSrVjn4Beg/Wi40CMI/iYmhXo3Ac6aadefpwC8
d/3MVBrPJff7K+9GxCb4nFs18oeiS9GjPFjOKO645OH85cbmQgVZSluJZHlUO6EG2HyVlhQ6yjsO
Di+OI8OL5HSaSXps+8haeQojviRLJ8MYlNlq5jZJWGVRincqUIhG1GfL+jJY2ZTsIafs3Wghs3pf
WZeV5zuca4eA9kixrW/JKbXPEM4Nk3oVg7LGbPM5WYgRm1/U4QWA1zh0UDF4rfqquWbIsNEp7R5I
SCE1KouB1u/+ZxCHjfgWTOeS3mBcDjpwtr4M633uglLvh2o0Yb3aEvRAjdkF2VGnCjL21rMd6Dpb
dpr18U+/Zo15gzLccu4F5iArlRwYa2QlyLtDFE0T4335STrb1wUuCiD9+7pZwxznqxdow99TKVpb
+VRpKSskrB7bCW1n1I04EAdwlKG1dKaI5ngkOBi73m7kN0UD1D3bD1yRqtfrGicopxQOUXUlHEz8
73eJGxcyQSVM4/rO5/84BQHQzVASMJh9kLXMpBvDU4S6fE8NdQlsDkoy+LX8Djpoc4kO9ujHzz/j
PvO8jWNxXfkAm0qz5uHrTO54JH7fVB5Bvc7ShVYyJwTi4azwKtDuRVoIt1rOFGpwaaU0C1Q+Rlkw
Iq8pewcVGvO4NR7tBDdIIaAvm3o7On99prHjSuq+s2Zj/cRmCSpVS43wV38veYWn7EqfDlJ+1zsj
xOeagS5t6+vJjILlgkNDcM1rpzEZfxL9046iVt6yglirExpp1f9SgE2x7XGmyZipM25GeHzomvVs
wUiASTck4vGB/fVC8RC0RRVJCR/lPaG22MOEHnw+YpXrX1uJNYyVo9D1nHa46Tjhd73U+2kFT9RY
KyzAMBcvlVQLL6xCLHR7q6aLsgwpYwysjEz9TvgJvblC06Dp0fSLZmY2Ifn8JLV8n7P0pVfWwCJg
m+jjFoYrEL2fyaP3ok+ZmCAuAsKv3k3b1G1mkLOrmKk8WYe04ilMr/eJRWdrFYwNEQAnlHFjX8nK
hcjH1TzvbMNzboJtoMsaBbYdF6h4IzULsVJVghq++80CMql97KLKcrfhC1j4L3TK//l/969vmL7f
FK2IpDhS5h+9QIPgxW8dw6GTQ5jU0CJT/cNzduJGEN66+k3Pn5OIdGQvXNWg6WUj3FMqLd238m/d
+C5xngaLT4gU3BqQyTzrhfUwWL/Bjn4ueKeUwWpOnnBX92U8D83vkojgzhelTprdxae+OhxhuP4l
7q6FlJdtAdvHBviyqs5oN2ePlf2MXw/cET5VUsmQQS0z5G0a5WfwuNfS8cdLj3pcFZVM/KCNrUq0
mLWYJMLdkH+V0jCudBvcwi3vFyVKYXvAmYnclywZPXWejvYtOfnoHum8+naCQUzYwiC7b4tlWaPh
/Gbiz/hzsAEjnr+zHTYo+GIffWwCFMoeYBb6GRMH1hqT6c8Vf0UKO0kO+CyP6NgI4AV7t6sIQ1dA
q9IfdAiqGs4bUNvSKKiV3P1fRRaDM2PBcWzE+cCpQ/Y5Ww5SPVhPTs1sUUbw1ipSj229BwA2jIGS
IRBMWFoFx0beJiwuoX+2uLLzeQbIUVYFtvz8VZl06lKjWdAYtlRP44+gx4C0lDXPYZz7/sy06iwT
n/xxMxyAmIsn15XYGuFb/ITSNdaE4TPkZoKWqRTDZ85sGIcmnzX/YF8HrDpI0Qgyk0uxxYZUrRrK
H4UB9aD1jInpgJKJNX05RKXaCKc5p9EiQZIQwNQWUmEBC6Mdr3cROPe/TJFizsUUl4chG3PCaGod
HH+BGN7/2YdyGCxaAANN2SVIj4n7xqG1CcpXmB4+IM/iBUtX8naxGNPMUg/0uJYvkW7ZXHtQPuP0
vigHL49pl0DY2M82vpRsmoMXMuiPYHP4sR3DHFcqjV85ir/ZS3nfqMUStyD5CuENzJuzn+6VdG7j
XBRlxmFD8bZdMcGjUW420se6dCAiqTQACcsSNPMxojgpJHp0cImpLDAv6UgUzYj7LqVxVKQAPclr
mdcdk8yNNolkpNOlKd0UvaFsT8ZXobX9vQA86hN6GVMPRxy2A99evncAjSURjWr6JgLxx8X9Y85g
khqtxIhIb0nFYyyd9dXsqJuqtbeFBxMtd0wUXs7ANZrk5HrFI6aRLcdAkhfwP+05wZfc9znYtTeK
V5czc1r7mnJG23Fcm+1MPg8Ti+dqBFaJcXh3SL/KservDF2y00QfcIyJzB2w/HZylIwmqI/nfoRj
R+W2PQAb/HUxTofuJRPEJfU1dti69nKaHqN8hjb0S1HZ4wRuMoEHaoo/AiBp4HyZ9VYYnR3E/Bha
WCOScpWH4lYOs2Cx3i5kfPNGhOsg91E9Qh49Hk0RROQDAhpwO9vhDsOu4h/c86XR9pAwNfDdf+pA
LBAU+GKm5Rh3UQaGw/yPJgpGKDZtl3MGjEQgaOMMwU+1j90pbnd93WZuml+6azFATjkQPV++rxgm
UD9zMWvXMbMCOpRhdvR4eploqYo4JXCVXCpSDA1XJZlq4lPAAQsSRj0NEVll25oCFKd6wg3BBSt5
kN238XSwURJQYrUaBd7syl76Vf9KFGKuxgpypSQMKf1uqpj1uZCmr8gvHJ9fj08B3DWyTdBrzOR0
n8T9ZJi8YSBQlymYzyWm87CdSprOSY8pz3VeYc+auQkUm2rT7ZDH1qTfp+uVGamJThrAqZScrQ/z
mWot4/4LUZFZ+hnxLPv8J8aGJ/lkx8oBBTFODJm/UMgPsZ2X8lghRlwd92BcUuFrrnZKJRFaNWpi
gyFUGgXU+JelkqxNwSGlvD5KgLwqbagNfrw6rPNA+Fu/BboKsI56Eb/uCG1g2F/5kqKkSpATGZol
NQLKJjR1R+XUEMVQY6wN5F2AYbL1Ym+JYEJGQc8MUVGc6YT4Z9YRD8z/h87zFHSd+lgIGx6MZaGA
Ppbq0WavfB4wz7XtVaUVj7SXWqiJn2MMGkQQ02y7L0l81uYIQXxWmrC+BBzW8u4vtDNUXahdXXKk
AYciPRigu8rz6yq5iSeDz0V/BwM+f64kVvutVrQ9HyVRboxyFNS2MgAM6BDeKCjuJCORwc5PfriZ
cfwPnFc5VqHlY4pCYzukpTlrkqHB8scVHX583DSSOhtq0bo6PAf7JvhwauCxqW6AVYCXw9EtARK3
Poc6H2L8BGaT7Hd18Jhoes/AMXmkPbGj16zZNTEe0wW9l/rq4xm2lboLI7BwZVGn5zJG7vbqUWn/
lTXQ3IrpJ7nG0MpIcnqgoNEODD3T7uNAWX4qUOaVKfLE9K5nsYrvJ4FvTTqY5YfsQ5zYU/Mk23s2
x0HCtJyKGoM7TrQXk4bSPXsZuHvgZ4oR4jgWVz+NgIc2VXeLYIMfJ3U3Z87Iv6Ph4HPTSZGhYpxq
TMLnS24V5o5Jyn3qiUVmqodnHnUlhH8MkhrsGbt2P8l7aYcsT5EyhhuSGB40hMYJWUxV6u8SCsBK
m/yf/OoF+wAXNPvaAML7wBt8UaL3jBUQt/VcMu5/9PG0Bdm3F4snY/CSBCwO6NDkFHOn8CvYpX/W
9J7A5aKRXeQI49EmgKciGtsnLs+1A2j4baJRmpIzDzDK+gBur9JuxnXNMobUTaCx8Frj+mRGzG32
gekZJfOsVAl275SFHGeq2AIyVQcAL+ApIj6vgudppbd9OW1j8bU0qaOvAXuj6t4r1gcYbUu9NM2T
axqeZ7umC/QTRG9XMtNeyO685RyyMssbBeI+rclltBpiqHtHvCzWvY6E86LbaiBBFbOCCOdgJfcY
SoE2mi2hecOO2Hw9FY8ZfJs2Oi47Y5aOPTf87BYoqditNsw96dwvoMqpgS5256s7PE+cTEf4Hy/a
4mygufkewG+mmJt691Qff0yjF7kpu5g28wtTmQvNfDSxmTb+FwyxrdxzqwlMO7XwWNaHYZhrF7BU
1QEF5dcQSEUyTt+EcHdeoF70sOc5fEBHWqYWZUjyX81HfOrNNhZCQ2y8zOh8LLsswLK2pk102sL2
9el0VJjleQF1nuxn2heqepfADH2jGIBvgVNiRL3mdSXZVeMQ9fQiqbJdylsVUQ2iohHEdVJAgXfK
50Yh900iwkXe0sidO0YUfbhL1ZXWM2uTe/FjQJC1lePGt8g7W1bYW5ekoy4eUXRUlOVkCFxN3Q8j
4n6NQllqDPEIFlEsj1xgVuE026ujrgtvY/TYmBvrEaoa2cKnYHLSb0IHDEY6t0wHzwsAfCUvaWph
pApMLHmUnI9GNZe3NaiIty+MV97GeX2lbhM88NJuoJkRGZOit21J0cWWEBDH5cyJ/KbvziGa0QUn
MO5/Ln2gi2b+7klJtlJRjhOUnt8K7QKzLrKAGzkS0UAG4NyBg3RhFRmWqABQ9M8U0CDAI5RsnMI4
UMi1hohXpIRbDRgzbyRTGKdRmG4DP9PidwJc5/jTdx9jFYtGESfdTq0QJLRovL//nYrs4iFzdWyD
ToLv5SMyyT11XPktEfrY8JzbrYLZx2aocb1ijoi3m1xvcEtwG3RfByiUa54d6BF5ELVeX9g5vBYp
zCI0hpOtqHg+aOOIlAEzdFYi8zY95tkapnW8a8+7tYBHzmHNQb1Orfi1EEgUJ2rdPprS1N2NOYFC
Hy/0ImksnQHhqNdMSutlTS8FyaqHbZXlL3ktg6Q5tjqfBVcsttclEDLp/kyo78tx6ZOr1Izz8UB7
W4+NYdlmLlTDLfXMCdLA9Au5XqkyOD3f3UVFS5Ec+Etz3BjEuLzQdDFZ/gn5WsEVr17JZiyi1X3T
t0bUwKY1wIDyeNGQtUGYOv9ZFeEmmBWcKi0to19KPZEzW8L7spXPrxDO44xzWzt8kBPa80F7GmtI
BdbqgAVSoal4X4RlSeRNk051h5prbUQToVBx5ui1r6bXrhkL55m2utr8KqpKZaEIEu6I6dzFGKuX
wFhwGWpFpF2FsK5IvWSfskBxaMrxXchj5wm/UK31yxRrbFSmKbs2A8ZKmt91dah6gAS9ZYecrd2E
Vu2aNwzCP+JAQufIc4S4Bddn0LYIGVQQIysxjQaW1qDfZKXcqSiOTFeVywdt2mIRboyHjPesRZHv
xuJrIHU3PObAQek3/ba41CbSBAyWhoDl7sWu0zslTL0AuYKGiI3gdIzy8yfBs7Gcrhg0hWaNgD7M
ETsiTGB+aSPiOu3cPFFVJRBrAIgzJGGz+4tWpNbS3rWCWQjnlc/NvcQVq6u1v683cinymIpP2IzV
DfiKLzQbWn6BLjeop2aZ2rTKuboW9bZiDed+Vxdk2kFtNpNqVj8h2Zki6M+AE9P8iikYco9gnO4C
B1DVV7BMYEa2NKktFjf3jx9l3QmmP5EcMA3pdZKkFx0cRk9Wm0dF8Tmk2tClhhIWEeh3pCFryAL6
PMYtT+TkKvvsGzEiIiR/LXh/wtM8fZhG904+fW8lQexzaa8B+WFYzCadmLrid+v+7QFmIZObMDQW
raXtWy5bUiN5Praaw8HsC91+ndODRgRJu7El8F8ZiGUvtQ9R5AxDvIIKUgX+cIicnMFVuvqWV7FN
cf80J/35+hQxY4ETcCIMlbVmGJR63Dcz8/FqRs6AKal0e/mt1lqx6OQ4iyJuT4ERm/6LRwyuDGaS
wMPED5ClCjQoGIA9nlayQxrbcEHU4VIjvDJY9XpH5MMwyVze+cX9XzfONSlZANQYRyeKWi8viB6r
m/Xf+/rP+QzTfcxH3g++DqKQAcLe0XW+ml7Dqd65Cp1AbH39cVeHYik6YG4oFNZc7lwpypu8h1MA
Z5cIokLOADN1Jew6fNTSHSnQ9WbVCwPgqecJkbDjOzRkHN+uEpFCm9YggdNh4QpslxP9GAMjn7Hc
b1Yw8sIqEBGnC9P/JuiVohGJSJcXKYphSyvAOVUKP2XRH/e/6SmfbmJJtAQ3qGA+n5GomNBZJN2Z
4oQBBvVM4V6CBMaAeNKtMuLuXciDCQ0DsfbazZPR3Y5w49veldxsWc/xFD3lZP08HnF5l+IpLNeU
Eoxj63xdzJXHSWGTQmGgFsmOBsZU+TiQaoZhXlBmCvDP2i7toEVtJQcVua9L1md5SE8D2uIMv1uO
+IXn/ZF9aynitGqq2v82rnwaxzKPubmEVg4oeynIMqf1dWTp59qxJEJwWdT6o51xbeCK9t8gSMn8
ogRYELuSX+PtuAah/zkFY8rfOLjTKHdXB3RZLvnq7/S8t8/SZAoU7fcaJ4cAYeX/cXBIai6Jfl9M
vXLv5LTwv9j7WoSmGfy4dHeN8aUnlWVSEWUFLek6hIl5p+DmakgGDfGuuKou8dG6n9JqPLd+VRYr
Mkq5979XMmpw3on3uOdpfgH3d+9w2XX2jwd+3REiC6LUGJB7Ij6gqAjdib/0QJfXtWSue3A5MYTE
zTfqaVDdkO1BicSUhX/quCR76n+ra3no3UvOtJ3cTIC1VcsOnbdf4LqclbVL6vLRrQOKNbdTqevb
nnyOwku5yTAbeWe+Bra5VSYo7eBCOywD2AVBNsQ0ZnUuiHYbDN0//USGoTekU6N8MVl+E51irYI4
B9JRce+LT9hqlqJxFTHniMavNpm2B5sKHsddfwVxqA3FtA/qPA6x/idRfUNBhpv/7ggN2KebmnfF
1vYyYMVCM0+eajO9j0G4f0xvWgCZUKzwrIvIIbounYUR8ksK2T+4C2jqYNQ0y9UE3T2hLm+/BJYL
VRLa/CUreUEQzfxjdKWM9PIgPzIVyg8WVvmxvsxPIeb/ZLYNxiyb+GT/qTItQw7VxVJxBLRRpgUl
kG22lcR7qHKOWzdbLC/gJUtIayqclOB62vHZhDnLgXlzZ/cqk2yaZkvaGREiB2Rqlt01ng26MlTj
Zha4M9XwG//nq//cm/yD4/uP75JHeSte2vMMjY8VNPwxhHdgjsgPu7jdM2cGxoxhHnKCUYEDHrXo
+54NLJKpZmAzfYatIENPuQlcOUh6sGn9kPxvmoYjZ+pOB8cmQ4eesU66K1FhPoLXtODtbMBaVD9i
8IeBm1mLaNFkpa7DOtuVXmsPmKhwQc/fgzlUfey5YqVReK7deMLvxEVB+/i5QyAOIn3pA05lo3O+
OAK8uk7inAPtPOzNhIRogO79uqnjtMf85ywl8nBukf/mAT1mFXx1/8pIFD33flSwsLsJu3+gdZc+
rKR7YpHEcdMNzefSMARfmgkR04PxshiB+7nAr6ba1eZHQUI8097c3+C9x/Vhx5r4iyhHfBa3crPS
kc1Fg+LsmlcKz1a8cUwfhz+9mr0d0APQzszVLND++Db+ktbBQNC/XCI0nu7bPEemTkqzAaIEVy/3
kULjzkC3z4hOi4KUKMwXfu08dRSv5X7ibce3bzCi/iXDsexbKOmW3lVq4gl+l1KZbPjkFkeQVEvS
AaRrA1BESuF3PcRGG2JjCeZy23XzGJilc53+kCPrdRgwkWxr5Z2HY1o0g0v477E81xI1dR2FWZOp
663oL8cr54zr5IELvm+yus7laeQx+S5k5VICloj7dw6rOWd5xlItG5OqpW7nS/hIJUuZcdVxS/Nv
z6QHtzip0eHywWvk2PwHGc19BuIhKjH5iG6d2DNDw55NqzwCfSXhLBU4IALbNIVTZDa8E8W3UDhv
ZpT5JkXmoBB5GVllL6UIOBrlDR/2waSNmG0LSgQQ8stwvv1BDp0agoW2tv26RhKqP/YnfV//Jn7F
rdpH/ttyonQDr3+quaa7I2XvX8nP4qdXFeoQSUtfJiqEmIJ2sSbx9MsU2ahnCIzWJU2+k/reVPx9
xPZRyX6ZilD/S9brIb5E3DMz470GcmYtLsCcppCrEqnT1dRkWI4dXJA6iuMRM22N17s8hZbb3gnB
Z/5eraCAsqquLgnhgkbdv0wvo9TCA+ZjcRiIlaqb5pR2Lu9T56jeBzdp7SVDQE6D4QYObz1cTuqE
V4Fes9L0RShcya049AAJewWa/nET6RWFHQgSClkUzMcciwJ5XDot2mfTx7zujcAI7vtQK6Uo6/Hs
5eo3t5tPwEYCCV+7zU3BcowdDdZGx7Vyuoi44C1/d8oVjR18yFFyYUA6XULMyXsgF15rcfsWTEJL
UN8eWzapxOf20JbJgGECDVB4r3G1vuDJ3j0Y6CoRk0huphdSzWlojZr9aG5dmmynsxRDf1gwFz3Q
QCAY/V7IKSr5louK3KpAXSeXsCr8stV76bxl/zAVvFuU67wQ3xEnNxu2R/Iiwh8cRdIn58yFvA1u
geMVhqgdgP7ed6fRjvTAwd6y3AFKysopLW7olVekUTdRfiF9bQvmcyjGgx0AJtDn6yCkuXCuxSyH
zqCI7z6SCnSdotiERWdFY070x8mOT3HPfisRsyvXCw0Iy5FYkTaStenB64jPrX4JslCli/l3UdYd
W895rsAXDWaCbpuWAz0oNDXXWIkqR15uuvXlF3GhS/we0ItAZpF51iVBqZUzRe+LmqeS3jGlRgN5
+2k0ujF4Z2srfzYA5ximlqpU0uMiLAdEcVQvyzmiAqAiawfJ7/mff3Wbl84R2/Hr5gH8eeF0Wh2S
SQKHmYLVOoX/x3bKL/rP6lqjoe2usUXHG5K+QnN83yRPiB3qyjk5a9NaD1iNzYig06/mLHGIxn36
Vii9RkxmNFFmevb7hgRZD4bfO8PxSWnT1uAd5t1Gk+NFzQx99yCigWDvrj+h5NfZ4bXUJvJyOy+V
6spl56jxyL4wuy3Q3h8b2i53b9LUIBAlN3ia7E5p8r4TJk7PzYDZbdchroUQw0/VL1RXLdjDyHWm
rrTGnFAA9foSyMddcu2pGCVr/kQFu0wQuQzc2rRY/dn1l9vlel0UsNcF/VvYAYsY+nMs39xk6RiW
0Ad4F2ZZbCQFQqqYsHJIDfF87MshNLqJ8Dvye65/skKS5hQ3ex7BH2SCUATT2BOnveJSET+JzLcI
5PdzV4LXhT4a3tWjoeK0e1bPSNf5Y1jhM9A6Cze/NTOg5O+hqYyX6b/Vt97Rle8dXoVgpIALzNXZ
zGy9iGK8uwDEdIZPM/+GW98FggthxtMLuZ+DMvX4BrPJNSG7/rBZK7EoOlAl/jVXALDE5bCGZATi
IMEZmi/eC/XOQpfIjBNhoVc1kUK/ptER1jP/7fVDGVYDfOyZnksHH2ua0Ai+K2sIpkODSOwR8NOH
4+UQMgEn8P+jw7HD7lKSi7rTDn0uoElS+B6Xi6jPR1tExOghmx93cCZZNb86P5/+CU+A0cth0EHQ
bSRjts+/x9ZRwYHUTFqfBYb4GMZMu9CkCzKSUYOm/2ZD2/4dEkte1RgxTaPnNb3QqiC+UQr23LNe
CDmXFDiF99+cmiz5Z8n3cAxcPtaNvfv9Ssz1DtEaePmpwGo/TFYrhoa+qyay+oRnETr0IDBX5V6B
1tbA3yy1G6dYNtlNqb/rRgdvRS7uuOx7ZEevt4DDZO8hn/l5pUTCzpd6CkroRuYxsQgnqTBJKUKC
i1XYdSN1dSPU9V4JJ+hfQv7eaVa6307kXAS79TMUuzb2tv5UF3tS0TuQgiiRCdTTcKxplAv8ldqV
C5+msF6Gy4ETBhWhcnw06aCdkVsMg2+zFWsOJA66yXiTpbRmiKdFai0C1Utv+mTc2STbn4WYzpVw
SfnFXR0ZgBds9xeqvY1lBBoe99XQMrpZQqOzvAK1TRgE2DT1b8kmgboLmn2lex5gKKXxxvbfaCio
LlDA+4Xjri636dNdw42dzorbNrKwVX5RpNf7O6RoGCARWD7OkcTVwDEEqET9ktQyQxTf8Xbulgdl
g/BHvLDojaR4aR3XKnTgx1x1GtvjzWzqMyidYi4g2H2ozPE+z15u0iKhZYTdo+FQC3iHlTboUACT
nbqoFIfb9ntIeA6wdK3gUkJLmIzOs3GQacYdEWJdIzGIpGe5h2XJS3nHCxgEiQz+Y9wH8mKpExJ0
dk2kQACFcsCegZr82XIC8C2O6ReFuwW8wsrq3Mb9Vcjrtr07uYksxY/2ytgjrqCfyW4DLJZ5Xxza
JllcrfJytJCCSseH+Pk8RPEJYIxYcPA3FkgVTlPLZjQEbvhVG+n2TWXdDSbnQwc/H9pQcKHwgdyh
CQf9WXu+Su6M+ClLYuW1JBwSYg4drWYL0dsMYwFBdffwG/mZOq+B03OLK2kybFQTAl+GhCMAckVO
Sb+bGxac2VkbSOqqfgwY8sYMRwLjvAqepfCuRilCPwnCeKrAlZ9Rk73/xBZgL8xcdHjYkOKgRBF1
vVRiI1P7SD1E88StovmZyL3fj9az10Rg64NroVkOc6CU+AUCCM+vdaZXcY2NNexQJEuL6de/hqDo
V8psNf2BQ1sA8vU4ANw1nG1jYq+JpJCGrGGeK89mTBj6USsFTswXIRUTMpt5zt+QhC3v7np4D3WS
8mFxPtvSic0I4rnFcBFjSW4d1LE0ww8s1Jl1XZ98L9b7gAkHVFSKoLX0MSoVxjN61PkA8F0Z3eyh
qhyi7iIcDHT+BzgujInnv6SheHyyVhoX2NK8TTk7lgmsWGoivwqVqLSVKOe0SD/wh7k+sW9KUHRj
CJP+RX2nArxb7a7bpSSkV+Q5NrD3CDOyDNmdWmFPo8+UJ5AKIjbO0sY52G17EVY+3SL9C06874qV
ipa3q6Q1uL2V/LD75qll0SY+dnF2ymtUf5byEfubtLW1mBeNSerslZwWpkTz7r3xLGGUfr9R7IwJ
MbLKkvgJl6cT4XWk9nqQdTFJQF2JoYxYLleNXzWttAqdcqhC6CXH1q8FEbf5tkUNCKl7VbfEUJrs
CzmtZL8MTOsK/LHKl21+DcUnVk+/cNKImisXGjYcZBb2D4aQFpFUWFb9WxoZeEMHa99p2TX+7oaC
WGoIOSUq4MzdtNMxYHXZS7KpIVyetLjvrRH8jbkAWlTKUNPCxWwOqDW9LxcA5zwncKDAxvYTfhb5
DCsFcYX4IPdebcK90JFePVz31FC7sMKrD7VBz0FD4IIJj91lm/tStEx99Y7vkUBKquuvg/+9JkOH
i8yGbKqeSP53f9+MQH60Oe9dlb4gFJRgc9GgXiDT41o47mtjXSXpVrLVq1c9gSTThfBAx/Lj6bLC
83VdA/KWK2u3Xsyj/zJvdNKEr0vBLdQk9ETJNqHj68tQmQ2NAsBjhxAetbCiCUnZ4iV4a8+Y7Q/J
UuhTXQdonBSAAQalv7JpOOa5GJtEwSkUaygK7pjdImLcgj47kJsFWUroYlBSH8veegKOtcs2emz5
qsaAuHzOpt3TSET1XFHCX6SGQfBZIX88cvqv/6sGIP9ike+4bpDw3dPixfm5J8UqR1HnKIrhw/wD
w1/+HJVULSlGsj/6aoSVDfr5wIC4frDjV5IiGu3+4jXHoZnaGdmJKtMJMLf9MgYaylMdIC7JYFYB
GRRBvz997KaFp/xueSpDmgWy0g8X4EJyxXWpVUgm3jaMFCq0YyaprQrRluUmJ+tKn888teUid4Gm
/RpEB+HVvtNfxSfKRii7Bw2x2LaAje8QSQUsAqALKc/oh8ion7etuvIOzf9Tpdx4Up5hNCBXu6mz
qugXSm6uhBuxB3Cok+FDV0pfJPB3BmtOM1IA06nQeezc+27ub6BKdwfpqYBKJXRd5mbnd7OWhfiB
RLyByrtegCUCh3oRoj+DlIkkR8svza8YU8cz6bEle7UiVTjdQImz4QmW6shqyrehjYv+fUTklITU
RTEF9t42ZztI1IwiTux2Lwj4ZpIq6D+pfm3v6HKxnjjCpfZWnx0sw6i2bDMqVxYmIbuVMKOZMGiO
jZJmMZzSnOUaLJBszjU3anqVPJylX+yb3mQ067ClNhltWigzaz6Ql4cys5oqaCyurbt6HqdtGftl
ljoosn1VHv6BLpJvINAUmzbMoq+EpPaCXiVd/vw+sZONiwn+/JdiB3Mno01ftE6HIwW5F0F+cke8
ZDZbKCRTMvmG4y724EzFA2AhVnkpSu8nKdSwP/FSHfBBRAdfu2g80IgP0vQCNW+jJHHvvYY5K+6Q
WT47sKHlnfrzUucdk/xR9igjTTMHdiRkhGscxbQNP736I+Li5s/NP6988YBDnndAdyTDtB1zShi6
L5cFoiA5yYF7xx2VjCHhN2QgE16Z6O/77hNafhhskxgZUuQBbet5x8Ed1Tke1S4iXXVyPkZeSnjY
VhFnQFCXr4zRMtcBSPEbgnC0r+SjG2nWokkhiU/pqdoUVezYuGB0c3sVSyI1vJ1OZpzNvSUJUSi2
mjpcG75EArK0ldbtMuCAdpjJ+olHcwXo/5thnAY5IJclCZxNL7ggx00LV8/o2FFC4mXJKpDd15yN
yqj/pk43bygxDJpEnvMgiER1Sd3ckHJlPIu9cchclnhYvrOoGPOvTdDtmEgt1DmSke2ZOcBZDTlC
OtkptDtdum+cOtCxlTsxw7fNYfjvIGrPvcBZJewsqSM3g9Sqca5X57+jpjZpWtOKs6rzj3rbI++i
d8yTY3wBAGXoq0NWwU/PeWWGlpi7QT9PoblxUVY0KC4LQoQ3uEqLD6ngLaI1cHq+knOVIaXkLQ7B
JTEVHBQwBVvKPvder3BgQLRZJaTtwoyabR4oBGC8P/79EI2ImqWF/tcbvPuA/C0IeNHJRN8reLQp
sY9rpmwJCpWqHcTPNvZ5MxWbgMK87DMygGcIijCbI7wohafUALIT1ponEUb0Ou+VF3cTpkWKBbB6
UMmuZQpt4odX2GjT+YIBMUOahjijG0c6glp/iQsG909MN/oqMvOUwrw01o3K1uq5dKAymJ6CwHzs
Z8NTXpj0bC5V45PlamBU8D6/ItIm/zLXx338alu0KMixykQBcBSEMHA/qXjggFdRFiXIvAWWo1Lp
96rulaTdDMMWmpHFV/PqNoiZJIyksN9TZ7koukL3ipKISuNP+ujr4UQP5jk8BvvxvUyUpNLml7o3
BjxQ4ildFXiRzFe/BMP0JdfT9NtUxvzoXVN1DKSm/DI4NJfmjY9m0PS0yLNtK/PkoSAwTE/oukgX
9D2zIaTmhTDCWS1xlXW37qGTm3npMXZ4o/qQsgMGHh6KQvB2OxLj6M+ze8Xh4Hr0xu1yNzzF3Np3
6LfDLSE0WRVQ1R3k10AzJwXBtnJqqz4ULFZgezK/D2SsDyxA00+kUEnqwGP1kdaylMEDdG9eOuC6
//U2RcufDWoUoonvXRSEoLmxzAWsB+fr/GuY3O6bwbMaG3LAxG6icA/AVYwzbw94lroBmUp6IN4H
ppoRsdFrhA4Rc8gJgdaQAAnDHVo3pDpXsfd5hc9l30+3aatof2/KUW6rD7gE46Ux+zz7EXLFry7+
wRrvaSuNSt4kZqH0scG6XYChEsGy6CtHEEruwOWmttnybDpu+tsGLqDYwmq8hb3qUqkx/td8Xs+k
fOuP8v0cjal/X4GDOjs7lXeaicJ75wTzvw2R+37xQaQ7wXZYmFf0pYf6WcYdBsXDSbRRbzcXVG2E
cyQdq7rkVhqDK0F1+Xu2a0y3oC42cWiJoZ8EUJCMOzX4jzOfW3kPFoOMf7cwEf0+t1Qw+6zoUIki
iA762RKgRGqoWoiJFXeNIeZ1+EXW3JggwgMcAtZ16WYhJFXFmdz6AhgrV/Z0ZVe3VrsAms1EN1OL
/HysI0Cx80om75wWc5SeYZP+3AhLSlKYz/P38h6zCg3RIZT8HHjfCf0y1SET/hhWr2bwOhY/qMVx
yqImE9UZgJ2If4Yru+bEPMB3gqT29X2dT9CKqEusi6B/Kyb7Ki4Vq0R7susitH5wzYjYCWcuiEC6
Wra3g2yXjFt03s21akGQPsw1k97VPlCaifAimJdIFFPEwgCzKMySTpOSEJ4E7brAxDJ5rpksbi0b
d7Zlxz87+JCGZHOSPeW+sSCHpcaB58PIU2+yt0o40VQ6wfknfO2RSXtA52CdEORqBI77jDPnZz2z
1spKGwunpW2NAWegfb+xBOVvh4j8XFBiUagidB7UQ/8gA9Cp9tj74QRRh1Cqx/tCsvQcbPjtTDRi
TrX9fX4VJXuAv9eXWKyGD7nFrTSLWe6YBcdc79FTo39nXNA64LZKTjjelLpY8r33XTbZLgvEhCY4
ozcOmcNxNZ37Iz4UJA7xCPO/Hl7Gdzi16qCCYgkhH26v1Ba5D6N6o3lGtzi1F48ILNkGQKA6UaaQ
XVnawXiZ4s2vgoqWRY0hJE1pJc9gKpwU6tyAmioAtaiI4F0NnivXdQQmYVwmJOfUTyEARFH+ciYs
LXVnrnQ/jeISelfY8N4zkVaNg/n1OGWeMSuZbifZg9xjdOk2VzPi0sDmkcwHCBtPRKLU7Ag4NZHO
p1F5xl2beXU/tMj3wNr2F9Cl+/glIrVupDf+3CrxjTI7I9FWBRnLtMM5KzjZmcYc62f6W7sNQnBp
VP6vwvhwfu8e6W8FqcnSZusPOfT8oA1nI+qD3fMCPUJhFyCodVenZnZgFE2vAk038MO6poDJORXt
NeFNApUt7+f92UVlB7zYiEdPb5zXvnHBKkp/0K0y2kEhHxOXoaQjvzkfG3kg3cEIE+Kiwue4CbfY
QOuxy7vG+zQq0/ANE+lvdvsXwPH/aT0Y1B9M22/Tf5i7i8FIQLB8YIajfV2qulWpiYfIMUS0fCik
ik85Fneden0LZcGi0lySmWhAbUeY4x5/XFvXnZyjgLYQvLmetwWlmizKZmrP3ySIwB2Pc3X3EnGO
d/zg0rmhm42gOLT8jpJPytfanDfm3oiNXVHOG4PYMI0vWsrVKm/Mp5LUPXGKnVFt5jVJIU9eufAw
Ns/GvPuEtv/KTk/6m5GWzFCjMUpL8LMtSExgHdpdQo+aH8bP25klt8jLSCo+AtX5MUq0PPXob2y7
k0GzuNbIsR2wk/2LDS8Q7orN1EXz24/XPs1Hq97N+u4xXlO7QehU7rZOZ5MTPz9paF3XHu3LrXJh
ykF0SUA83eaH6QSLyd5JlrSTFuoDgYw4Mh0sXH+OXv03j7GCqG+iKHYXdJJJ1wgHYIT2Uymh/HHf
vq9/UNtJBEGRth0K7/BAJgLBlhPwIYVaTF3nW5h7nqGMVtgRPzU3JmRGc3FsZ+9Pex6LEnvZFcU4
d85CdCSm0rn8WFeWFnOjvh7EFpwDYaNHa05yoi9BGWRQezfli5N+t40FmrEAxEhW/9+mGfQc5NjP
9OGPLvTrwoMGA7QonBxLWe9FLrsensLXcncMTIry+gSyju2Y/VxDxKaaLp6xgyq9xO5SI5RjpdkK
D4Bm4n42QAjUPQQzsrl6hQJbE7oub1TC3lzjVs/S/ESy7rT5d/1fitwiZ70AqRLEvTwMFsHJ22tz
ilmA/+GrE6A4DcZPqo4KPTLsK0HynktLdRUu9l5im254DbCcwEaJEKF1D+VguEhHbMleg/9um7wD
CJlxnrPuodjjVaD4+SR2ViY8rQL1sjFCrzzICqNz9VlSZwgQSgzi6UwSrLAvFFKXgbyCFPsTta1V
5oVtHuv/E5YxMv4xFL12iNwxcWTujdn/15Cka2SQ8gwJBmwxk7qtw9LSLrYrdVgrz/0K8jSJGJuM
3pYKOS7eLVZLvtjnDKrGjo3iv/k/V2yC+H3ggm2t4KXBw4q98DHK1/54jX7xXnzbKlL/KlEz8GBL
KWupuDgMaJyWYXY10X1mU1Hezpw0bSY5yik5wntpDcfUoLbnzNjB+Z/cJrjNu/2iHfETQoo4CrZP
VBKu6pufYhCCwYzhYcB/wnfLzJu0xgP9AYr+GSULLI1XNySPCu64yLylGps8+y4rUvReNhBBAqZt
ElC1wMtE14DE8dMG7uMNQhf8SVRDXqAT7IA1h2AMFsIdSXkXOnKeIXFdJKKFyrgkScPV8IldUs6R
czXhs2+nA5Q8lWJTDSvXWuIgn7feCyuM+1Q5w86Irz6NnYkGMD73a8XA/CLVAjJziazT6JODdQMX
nFkXj94kOydJblEhIqCo6xu55xQq7BKdXxURlou1QwGw8AMZE+1sAUiR/jbpaLIDg+4jmqtum0ax
fajT0I+BTCtBTY09jf9RTUD3aWtTj9ZNtsLybZbQrr2WeYxRoRG64wfrPUFpO41yaIkPbGzdwiSD
tmeVd53GLl1npoZYaOtktXr4hl4CzSfR9yIX7dBRcOIQPtjWVxu4KeEe+aPYvP9aHD7m7VUxt8Uz
+AZdDtA/2D2ZFnpM6vsiFVAfBF3H5dqAtJ8VjUmSDooaMD/wrdpG0RL9f2qSUv9Aw6823RPxPR9L
t4LNdIKHKTKM/rUDPCS4HdQC2PlM1ATk1j61wu1HjyxiZ9vXRYHfurF4oksptPflrJFgcBAFr3Mr
GgyGDnx+uUK5ziCOq4XH9tkl/tBSo9RA9+FIrg3mAPGNyBzcKvp3jTHqDfm64lsDNQYUvqrrw6V2
k+dPXUQsJhTxNlzxjOZUcJfhCoe23TyMgrRyzjRLKfbLeP/W7ME/yLSzyVewR/PIG03HZzlIbe9P
MHPZVs+V4evbysR+K2wZZgHRkOOreNjW7UCiXA/JfYlw23GBau5Ps6eV9ET4s6Pk5u2VMPk4zHSW
dnOO/PcmTN+cjc0lwNV/QqUq50Rs7p1dbkSY18fTrNuGk+DCYZc/rd0cdMJJPxNsvUgcW8e1+Hui
vL3lq7DLr1L4P2sJXHQY77Rim8y+VEzO1a9rX0rUzA2wrfLor8qHFgs3rhXA4yWUbFty0WD2LW5R
DW8TKwp8etQLVGyCSuUXQvbU5rSyMZaYTreIqPWgAcaRBIQ5RK0tUVtt4EqgJKyZE88qAcPsSip6
XwypIaNAu/b1ZpJ5m9BIY6NGpthyydWpdl4aufn+64v0pwkFL3Cv4eukZMmOifyjX0EME0OJ51p1
xa8E4uiNniMO3+YjTIYjSMwyBo/8bufHQeTPMnBV7OX37Vrnl5oN5c0JBkzSmwr75AzbKgOTTU7V
iwX+ueq/kT9DZT/wlOLlJm3yKagAFqFH70h2ptgYAQlOYspUsWMj5M0T/gFzfoQx8TXc93iWLOW4
rZlEjVVcLqXoCyRfmgRGJ4x++0cs3rww3JQQe/ns6vbhV9nqBamBkyWCyY4Gd1LueFrIqwnIt6a9
hfumpWBpD00b8iXoMiWtYJq4u7Ua+y+FwsSPp68R4wUirH+WAcZY3r1a8uCYWHdka89s5KGMpRVt
KrgLXj6ayFCJEGeAsvl63qTSAcvYVoIjBDKQ33y9KtxLPDWWw+DM+IL2A8/xX4F4zyMp0SBLZ2RF
Qa9hBYVmoNS3nrKY2JtNXDrIHWS3LAwl07/P68E72G8leCZ9FcnEByceO1wZjUWo7MzSsQOHKfWB
zQDnsFpqUmW4Xls88xmxUJyVE5pkoqtQjSVskAxVykCNP+KV9dkgWWzKn6HelO2tyrbEkG67Bxk4
hgkSMH8T+5CF6b5DjL3kSythaJ2EyCFYfL1hfhDWLlZhTPN2CdgA6tk/U0dM8vAoKvcCdoEYNI7T
5AbHtZ2YtYsniZqLCNoGzcrT4idHSwHvnNOGUHNw9TfjG2P2JNRlPznf/EM3Pe0DhIgCzUIDkhmW
yid2+QW6RPn8IDpvXWF9wX8SNOyVcByVZiBtjXlvdS0BiWc2DPjx1xmbCjAnSERphvm4fOH1K+VK
ffXqzn2LCFq00lT4rvY8O3cGdeO0ovC+8mO9arWD/4vF532ikdW/Ezl6Fa1zrdzjVTSZF6IblERo
wgO8/dcW37CP20aEjHvIwVb0YU0IeOmB3tGlehlREmj7OT0bCJaPKlyCv0BHIe5l/bQ5G3Sd5MNY
KzYoknD8LLr8foIc0CZfgI60O6Wfae3diVnGD/k1JJtlRSpQHbVUueMvkgKUq86xb9zkbR6xaFr8
xP3D8Ho1RF6dbhInywn264l0XhA6mdskdgbl0j6t9d9/2BKfBQpqHQqupiqVUBpah7qOpmzvjFsR
C0WIk3CWPJi0HpUARRY8xBLrg7Mava3WYVBDNPnsRRpENacokbCsFbHIgkytM/Io5SeDJYCz+ojf
m3bFFhk4S96Uw7DkFGNC2d1Dh7ky0UDgsNZc2dljcxrs6cPtHWtDR3PbFjLnqHdXCgRY4bpzGJ8j
WMyuOmN1NZHC/xZ396Qd48FtY3h5O5IcZkRhXi7QCo4BV/QcaSCMzPGav25Ukp3plz+aIrCJj3SI
nBqD6fY3QRvcM8PI5//CLzgwMblZCW1QBl3zbvXkrX0dZu0iwHQ+O50WxYz1ceE3FIEkp+bn1+hG
tOfOp/nztOU7zYmSWVSF66E8ffuQhZQVjdlWEL/XK2a4Fd8s4Mxomy8h8PvutnuShylgXWAI7hL3
d3620ISqxW1UiMChnxJdhUZWx8d27IkYEpQvD1+eK870cdCTqeQFvGWVOrC9x8iFhShFM/iW54ok
xwz886xesJxnIjc9dH7cfp5HFGU+Z0i5xfUyXu+uny8OoLvVX84HEfx6n+IXsOT0Sgjk89M3lkJR
f6tYFb21u0CJicqM6dPgyBDrwmuDHDKpYb5ipuoFZwtDzrleEp3Q9W9vuetW926/FykG+d99GlGA
nI+3YG0YVmd36JDJkSnTdh4dhKvx+ROBPr2/OGRWsR5ov63RHSCcPuC3Qo+bDlHNzftG4opj3VV7
hYMtDdVXSa/q0KnkF2+Zfvutk18HybjBpP8kxRL8gnL7pnxZU+NSld5cQ9iO1xo6Vlgoq7HNhxQ9
cJyfqfVuhfyPgm9k6vERbNDNh4Au9RmQuT92uA1/DV3HbHLhnbdAk2ANv9h3oT5PjFvDFPDp1iHW
aAYticaIJjAuTUNgAP1RWObAG7lcGrroVEY6QA63KeTgIl1XJN6Hkwpy+75a+YYwE0Hh9RQfZJR0
0KbtOn3J1OTuiEUExbEtM7LYfHe4NjaZ1SJ2yxOPWxHSN5xGJt8lRsbRhyv3S6SfqI8I6wQcFuwz
WMLbbo3ZCe4UqkByRVJc0Sr8nUVC5jTxeZPWcp7PMRF+flrLoIlFFcpkPkjGriTCJXC4RpR/9+NW
YbozZQ4vLB/jKqPHFv8XwMJ5nibcRmazYKVzMTSD3PShwLwu9ddbIfqlCcIMZVjy8EiJtwjIU12a
IPdnPDAlvMKB6D6YcDJ88f052lI4XTw+ray7N/1EcUB9C1zNCmFJs8ngVF3rFFp7GMo5mRQzK6jg
87kinWWMffdoTvBkeRX26USjvlyxeJ5cZNUGOADOcnkaWXPXznj5bi6U6NDpLgdvDD2B4PIU0NK2
soaj7qbr9OBrzq2gNdrbUaXc2K5aTpeRTfdvUyd1WG6gTWkpUcrCJ6Gv/tw058Z/MI4pKkEKgNrC
PS4Gp29Q4NQeKWgQpGBUKQK9aWTUD5GNi938dKBS35hbrgHuxQfDiytrRyywqgniIgdweus/b0P3
j95llFU4KmG4fyWsGMw6eCi+rm+rYZSNxPDRjz7O2uE30EiYWJrthW/iiSSF+Qbm3ehvUtaSiW/G
2EHqJaH8GkWZFwXu1J34rSejkgkjHTnwwZzTFS8175u2KlyElR5ZAyWNLPFpBHWl2rertC0S7+Ve
tpGVLAqNuu4gOFoHdEx6Z5STxogtDb4kVEIXF8sjiQYpfL3DxSo2yNIcwG7fctdj54St3ErTyLlm
+lWgxYujLAVqjpC88KQ6TTxKXAcT3jaDwuB31bXreXJTJiuNiNpxjarwiVBU3HJZgmsWHgJsvLu0
jm/NH/AIjZyq8ksUcwZRcEBoXpI5qjEYgzR66kaoaPWR8Q+IANeO8gbB/iXJTb0Dlx06vE4O+Vtu
OQH7JoaLtWBn3stvik/dT1ScSQMI5mpx9309bOt2F1scocZaG+9oga+6Evmp3SoqC+yiMVseun+s
Bncm2skCuqNIF/ztZ4wnU1fj26sXRKkX0egHaV+Rzdm2WDmPdDhbIPQw+vx9HLf2YBZfIQZbMC2j
khwIhQ2NCORJx8Wy03YBdqcK3E4WzuuNPnppn4XubutrdiQT7EqH6btb97wTlMWLfDYAPQKqlXJG
yh5vKSsWLhBlvmgIOgwp6808rPWTcPAlmZwSzJ+ThAJkPQpnCesP1AQg/IG+hBTYwm0USgN0BNW5
8oGksRH/s4hbUk2T9n0DQOLZx6D+ObGjGKmFE3bPc5Bf334zTNCe+0BYhIDpJNZCPDk8AnvO3aYh
9Ul5T/xUcua3AO5fYplywfDhmUfp+j1o0KxqhDnIS2YCREvmhJ4cbS6E6wTao0kuck4jCQ6JSHNh
9/oVml7r+gJc3HRp9J+pTw8kb+n6nj8xw0hYBc+IfO9FJb/nUFfn/ay9IuUs2boRjuqZjxeymt2X
whAVVZ83u1RKHECdFSDKEA5F/FRX8so3g4hg7gNcg5Gav8eM2m1zuu1zbMLvxLyw4J0GA9IpuVkR
dCPlIcZ+dOYATbQgFXL0pNRTdTajZiKsE+DRs1xwewFcmq27W0wlHf0mA6fYBlpwJBM7LZnGlF0T
7HE3Gmwm9nj9vkmYWAPJpeqbPAnX1tDYO1ev0dZb9RPdy81Kywl+cKZL63us5LbhmCUIi6aexaFT
h+UCw09xEhz5RSdEg3HwSB2/wjhfUFEyDPRqmFM05SssFUz7OD5Z7MfoWqeg9sqiL6ICzNhs8KXj
ydczwR+vXOSrNV5E5wSPi5XTu5npSdHP0SFgqTvILIw00Os0ZwoQO46FNp7Niva+39xwFF2r5feK
8cjtakZb4QA74qKDAZOIir6YxPCBNVOfW0031NxLXaVghMOwI8yTWOSjcnY+cnTzf/lRWP9khuk5
3VIA+UBJzYRN7HRVS5VU7zYbeg1+u3TeTaCp5CN2HYPsMi/iUG6BW18d7AVzx8YRzSYE6eTHqg1B
MMbvkVCESwg+XvSIVS0PplbVcWoEljpDYqty1O5daVCKtE2uULEIOPNJ/auRHMVIsQtFCaJTmZxz
Dgj4XOg24YlBCH2wXKATVB0GDzMzPvxUNDjGN5kOy/wR47KWJpqEgD9hbLJpJD6TNY47481V6Dry
i2P84BIxQSrxsEk+uxGkGB/ovlwpdJ8s19l5bePXfaAKb2mervxsW49E7qTOT1Q9u7uAe9eLa6OB
kWD0qYfOFLZLj2GScOdIAVU12SCFMHg06l7Gd3dVgxVdqNLB/UDzXyFnlvQ1FmpZk0P1OvRREN7Q
idTslGmBMZ6xFJCFMv+8dkW0kwTwL8kkRV+hu+yelLn8kIA7QCPDmYZTI3qPMYquW/BIRNJDcxDQ
09jiZrSg9Kjtx5TOt//qMO2OUshZsiMN7UNL21WSU0FfYsgzNXiLTT9Gh8almFlhufY2SgxLWVjs
RSMs93vaJ/kHh4KEFzeLyxhZp0gaLolWA1M39QIg9EG3ueFPHSsthRBN1mkStqBbrT9OyaIaEHB+
67lpZuMVMXz17Eg1H8nw5NYDyT0Xj+Ji069oU9CNsIbqCZrnKq/43aOvn7vj9uRoTn8FEk10lXMo
TpWYM5NazLbNL+iVeDZvr3y48KFCIKORfo4cETVRgH5sU40EnomgJNDNJo1HvNa8oItV7Vj2+g5o
4DmJ+p1xyF0xBrsbQ+/kinhUDBeOh3FlDxR6GjRbVWKrZNt/HiRofIxJ9/Kxn/DcVKN0jqJeC4d0
xF7ohyid0IAf5CSB9+92YsRM55rJ4o+qVbe0Vfu+62Gm9ub5eX3q+E2lLOWVPkdWqELueKplcgqn
F+oTomHkB5lN1k4Y4LV7FwEi54HsWxVornXZP0qTJtdMenQeU04/DH476oPbE/qplKJE3A7YuFiy
9PnqYEFOd6KzyvJ4e4Yhtaovx+yoMvRguUEJkuPl8FYYeVpj5JY3Nr0+T1wc9BHCzEG0/T0WqEqI
xV+UYdyO2JsKWAmlSGPI6ARhp1fuxo+Fh9+JaqLY4LIRZ4VhMPOX1A8eYpsMrlrIjf9+3mCK0zgs
ZmQp+e8iUXpWzp6s0c80Y/Co8BBXWmFCxzc0oeID/6T/bbPeeleyL5DXJPD3nIHWWcqKbWdi81A5
ihFaazcpJQMgnE2qaLc+QspUw2xWlffOO98croUZOf8um+OGECPyj/Ef54gxcgHmSrYjUc4FeIhY
A6pP8newOpeNCMjtPGIchbNLSMifOh74ksyGuULKcOD5I3xMcTGP8qo4gKESEaI7iFxY/BJotKIJ
ekXsXjmnJAHH6yv18XrnB+X5yKayzFehlMuP08JSswb6rq+P5wtjO1/6zrlWgQAyPU3rgSkRpmQw
mJeQTuO+L12MvTlYMdkWzXrRs9+3CXYFWHwHEHg7u+2hmf6xMUtsmIvYx8tQm3K9qB93lUU/6DG4
8u1AvvMdCaVihmAC6wb9JNIw9sKJFV3QS3XUoORl269xTcNPepllgTGwbP+51Co1vAy4fkHZsq0P
6BHCht+xASiZeKsKu46uxPenvY4F9qIowyxaYITKARZlxxNCdIsuv+cWVZ7J3jEKrk5PcJqVXG8J
rMO2IkmleW4P+27JU0gLjylxP+071HTzUGxV9NYMr+G72WJL0cpf/VrLWSFCuljA/bJ/NvP/B2Ph
0snC4VBX60CCt0adqOvsCbSDY2Hg41+gaVFxHhJ0PCYGPCjcv9WDU7RenlSEJgtGnvuUKSSKL1ax
eZ0C5qFYoYGPVqGWGTHwUOZI9yMFUJNoI5W1VxdaxnmGetn9uEek9GOlSz3twTMUa8rr5V+gnEkA
dBz2u/8pJDS3lKvKptiADoIytOgek0Ptt8Kej/jM1krrD/2aAQQvMPSg5fcwMHrQBYaLiyw8+r0G
BteaXSYLHOgPhug/R1UVOJH0h+kfUA/Pug831fAplFGfiMuIshPA9B7/Ve+I2P5Ci+wBpopcB5sY
+tTQMum6ybGW2WMzzNkc1p5Bm3st01kSjwORaaR2zloir//PCtlVhoa/rApLt72vYkUyjyRwZtRj
vTdUCEIfCyQTUVfoYHTfGV0+Oi9hFBO5pFKnbwVuuWDipTyHUneBdKrr6krd01KZGCVkkw6ZC4Si
B/We+iarvj3U+WRtYhBmB9inO/eJq1UyRsrLDaUipvcexTv+7koVCBQ1JvT0ch3GUh9au7iETZw1
5BgmsaQh6y4efdrPUQp19g9Q2u2jzLJ2v1fLPpxLpCD3QCEyZcyxMQKSD623316iuL26vS8L/cJU
8ZRrKdKF3VMKrCdtyni4oFJqeNV1z9jQs4ffQYRH9G+gAwxf27R7AeDxrmcTLssccM+sdke9GOii
3doCp9Di+HJYc16ecC9/IvrrAaOzw3tCQyvp8EzvzF6BZSHAMBqOItThzQGCsq9BtMUV/sJOdVad
zy5++8ALlYMEEQgDECfCrZqe/WVhL+SMOCjc6Lp4IvFChAaIH0YqJB3v7LyjwXY8jkF3u827BYE9
2y+qQb1vRpzfvcQrXERmgG9bDtbaGwofmxSFBtxRT27MP177SfrS46+xZKOw76HtyidqVCNHW27N
biQ/s7G14S96lJVRkHB0PWJINX8TB+aOMH7msCFBd4T8YGRPJJBHCEPQ+02vB57LhbEBZJwviZkS
jFhQcSknvmU/0drBdv9dQKqRlmoauJWMQWERL1eQznH8IFDBqvRI8fY4QVosreM6luibKi9QHm+k
KDTK1Ce/Bh28SfINl+kLW0PRCvQU0ZAfueZo3loE4ofMSytOBKxGC3YlDpidbF3jELM+5oa8074T
SOkM9LukLUwKJdBLvhx8GhyCiGIjGsaYcN0vyOUXxOy67JZloPhjGA++nmsEKamBqhuaqTdVec3G
Vmyhn6ok2clUM9/T2eg9/KkCUy6QBKoKYOsWVO2BwVD6/Q/46tNybe0MofZN+TMeR2B0vzBqrSSN
+FbQOsvYkc1Jo3xX13nEPVlhCUUqex6k/7KWULu11VSabJVOMwvDW0fLh3OLeH8GG4DlRk/BXb6N
WtWa/v2Yvks0zPNU0VyMcsYZn+TWmeOqk5eWthQxABXdC4pWwLkhmr8ebTD0tW569o35gZChiFgr
4AxZY0Y4UPiDqu/FemoIRzLBPjXuVOhs3F0R8alaMEYLWbpCKPMONtFgWA2UJoF7A3Vv+zr+sNUC
KJXAgL3owFjhAsd1sDlEQ261ft+e7vMc5H4e5LuePjstr7oN/2s85fq+RTevTwXHwBYFLm25eGXd
HT0FsHoT+xCy6FXZznO4eSqDPEhSyk3sqJQ/EN2oI8VcOlR44BYxL8b3EHQEX90sG+LB+ppGAZBO
AeEzim1Et94VVEynuaNoua/RfuESPgDIjsPFN1ZPVZwArlTWwBnIGT8//waMouI4hqWTXOfViZdx
2CFqnnGTt5pm+MRdKcqQy/sWfbXDT/RGD24KfvATNuxerPl0E/0YXDe3VossKivnlfR4wwy/C1IM
K3HqYoBgpNFeDRcVioa7YmTwYHkSpQO2z6v5fN5HN6Pv/ykHUterLTjSFgerzr+xwBbht9RZ0qUV
HCOkjY4FKXp8vhG3QWEh3sKFE1Y7ZYMZBxQOU3OE2JsV4PnWBpDXTsKHQZJ2Wq9S8/zvmx0zPIrr
RFQkJ3kcRmLBkI2MJoOhsqEKJPOWBLl6ceUg7mmBcp66roDeoXmAW8qCPFDzAIH2ech25mMgoLss
MA0ivdgE67rzhFWwBPPHty/RtHTHrw7n8ihhvqi55rHgtFQDqgtpCYW83c2uCKX0zRcn1Bi7WIgs
gx07HoEyLPAxDCy0ai4CfdmRKfD0lGT8aYsXLMiGPxv3ykvgqxzbIt2+EdLO90RdGpL2xCizEsnu
8kwMBWiNq/29MuxdUY/KlKYAqLAXNXecRKyH3415Xhq8guo1ojsnRQFBv7e5GcVXnBrLqrnNCM7p
5iugARWE2PgMTsep813SRBwaq0UrgWJBEUgN2SvmkWH9luvWde4sexiebmD4a4HpxBwiqbhqE4ec
r7HLOkeSFKFWnLmDTHlEeBw8CaxmmrwFby4ES+2pV3hg0cr0saCIybx9v8sJXLoy0qLbx5zodFKQ
K/gLDvx4PyhqR9QyPt0Pgmf0byEdzd8MuDi9Ise0DIc8Yb6n3p4WbYVj33octKOCkPJOdcRxrlHV
OSFqfiV15EQPfm0i9K/B0uyN3LArt54J0uYPqypwo8BzUkEcrHGrvx9Iq4clWU7vDMdXjIhYvDF0
+IiD5wRZjGX56S0PYqW+NRidciZ0KKMbdXomOD+H95xs5MZXpZ6faQWdKWWIm1ayjdp/DKjzf2Io
uV6g9Ckwm09rOiH0X3wLTCJ2UEgbPpDFbgCkz/NRE0sio2ekELiiILU9vHN2KpAwxnN1A4oqqJC6
y+zBl6gH6UdAwL+yBmSsPaMf58VMGC3g2j34YqpCHv8SJa2/ObLQnDuTjtiYvtRE1zyxIMgTcY45
ef+B68Q3FZTqBJhVaueHUrV9WPlIFwcob1nKskmog98FpAXwLW+iENbnavAr7R3UM+59WebFU6Zr
urZQ3YyPm4O5K9Gstm+apUK8ELzg8sHIIhb1z+OdBaSgxg0uml/DRycJvXNyZFYbkWX/1P4spdWt
lxvcy107C948vE03/BsH1rgatXCLiWjBWAAfhx+8Xpv39OUHZA8VB8mPLk3Z0+jH+Y17XkJxF57N
lAcYvalRYAmmg+9fdIh4+4oyHwfXJ2ardiIGfXfxz2AJZraaPdfEN/s/2fj7tH4dS4jwmFZkJnZn
CQaFZhAPAGygGnFG2HY0C0VmK3pARR/QcCe9kY31XbSUlK8dvnVo2hdI4PvY2axe+2Rf3J1G46OA
SQazAv12fqOOLZstRp2TcbYCQ1OFPJwO1tQlcT/PhNmXUk1Nm9swAc/6jxaBz11gTtw3Xbxe+05i
h8ZYoxjjzdiUP6UaJUuVe06wduwrX5v1nA3Ktr1+lGQ/iE31wx+iBjAKhbFAtQWry2o87b02mAYR
ZPrYVxPgbH9uEvynWEmYoW7xXcb5VrzzNro/KgOLokmCuvHijeNdev2fhWcTFc/a+4NSEh2cnZ2N
IrdvBJiOu9q/s9BxoW3KPlocsAYAzu/C2WTEA+fW/txPyuuz0X3IL8+r0AFjlYgDILIX1fZ8yHac
FIxUAaqhhOhaBLVfBQVF4kYHsnOjZgK/wWh04oM+UI3oOHTpbnHeNWtDBKP6Fcv4El4cmZinY+nq
uKw7q7CC+uuGSyqxxPjPQK6MGKUB+8VHiCmV/gUh4fAJ/mPrgAm0irNP8klRxYQjtwvfu9AbXmHv
Obx9Re0Q1RgPt/i9SijqP1qa8XP/6rzTeAh33OX+k5C2MmKQ/rnTp+8JxTDJzwPN3jHA/gEMlUxM
y4eKhWLJ4pm4E0s40+kRCN2i5qWoK5XSCVHv1fav20HY+hdWX1xKUOKn8XnDQWpECYpKRcgEBKGW
FDZfhlNOUDVdurCTZQLJ8YI85zVlOaC+aRnfDdJvVDtaFLQ7uXCk/F96qHcaUCtHke5bf8rnlTZV
y/pCcfpe08fR0WvIkjA5sR5MQcsMfuW3zTXVFLbaw1FYtjk/ir07PXUTq7pRU10v11XqHv13BJad
FEvH2KNZFnY97cjkd6kXzrdjUjJRLC1ScmeSUqng1uhxFhkQcr+EqIdKYpec1PXx8Vbe2EFRCck9
7NrHOUYtWeNCx5taPHlwPMIurEbT4n3wwmV9WTvzKRmxum80UHkv24IAeIJOSO+DuMLJli4treLB
I6HsTyg13Yg+hno82A80DemwIWGfEWVwCWB2AW0A402U6j1px4RdU8BP8OOL9EIPpNuom0+YuSPW
SaZ4Le5X65WZbVY+wJygOaRyn7KcB9F6cvcnC7NkfyqAWl/Y5hEbG2qEcKMUZ9ZPQ9y4ehQmtLYE
4lGfka8caHDY3UlocSh09psIg2H9G+A8MAJVlNclIyEYecKdF1gg4S++lUUg0R4bPZqYDmIMZrdS
2YDBB+aZaD0dnj2DM5e8yWtN90X3yEgD3NLM4Ss4DG/gYq1PFwI6+h7t3BcoUqKJ4AZ7Rw+JledU
Vr3H8DSneITNEpscJFqLqsagbVhya+xNukQDJxj8U1Gm8f/iQo4gKmlB7fmM6fUqolKhv/diQelj
oWqokyxjC0Xg2puyR/zEHRdiO8JY4XyJZhvwH/6ED2/Q0MDVmrVRnYojZFi3VqH9Ke44qqjPcAFx
19fUianIN8fROEH2GWbrtE7lGitaKCcw3lR3n3wGt6AaPPsfZ8Cj0TwxH80Ot72LHB4nZsPmB/WN
KoEDjC1g+hpqqjWp42AjKex4dwawS5LI7Qko6vJCbsrYtMVdTOsOvLz4+zpC5ZxBXFZZphqYdBYm
t7a5M0xnHIqy90PV7it/uC1jKeXjEkP7sOGkSq3Ww3hBdhXyt2HDJ7ubyslBW0CtEbVpvdWF1yAY
LIQJm7GE6G1AzSEGrStvcg9emnFSrM0XmtSc6CQDPg8vVuNQMnpi9K8uV+RhLAiRXLZw6wuFBSmf
dtE8cPg5107xkq2bWlXgJu79OShTD0d/QW0d1F+3MP81V2NIkuFk29DeUAMutlTLxrnxC8owOOmF
2cDa4CJ1cyAsOxqa1QKUm6Vim1l++YnIsZ9KUcGk+1dmomYMnG8PmgAtjS6LEfl/zQBjxjDSZziH
8mlR+FS3fmQl/ikhTb0IrUiR9MLZkaCi7gl/3O4CsA8tTYhoeidGGUTlKFsfGZS1NFZhba0PzWWh
nwOYknUsEnonmU8o2O6Nnin78AoYMAzUVpUqcmfi1J59oDfBHD06fGNez5hlXpX9/BXFHG5CtPra
/gK+eHtpEjwPxZ8Gpbwfozs2DgXROyy74p7OzOKJrZNnj2H4FeOoNmQJgbcVbfMNNsgcCHqrXnU8
tLNv8/IDKbzBns4C2Y2lMQr6YllvW5091JhqAGk4qt/1isDqjPuIZofwCuKNeY4k9m9x7kobUpD0
rCrwAK1CW1zI7V16iT/UzrOLBxzO6ZpJKcutO3vbRJC+SiQ/PXnIIRPY37JdhcwmDYdzdtPpyEFP
Steecbk7BPfVUQR5vCGqlj7Oy5pvqgiw8UPY5kn+CnArw1RYZ/aqgwjV8q4ua+dQoUri4yUZ9rxr
0kP5k/cXeBc+LtE2enIk4xsPz5bn6AUhsCqVZemhS5jrbMT1AR/wM6ZNPCSw3MbP9aMR33mMNvRy
1QZMbzQ1V86SLXKAU58cjRb8eWVTXJg+ul1qXnZh8W4uXzEq9y1ZCSLujoSHyqW3fsFvA0VFw/E1
Mu7Hc7P4HV/g9jMy+f54Mgi0nW9jFMgsyDCFu4VUZgMo3+2fi4rWiPsSCrf0N/aaXsy8VSPLozLD
iXwJsqRw5L/36RiLmesxDbF4Pd2pTJm2rm+8fGJxKKqjmJC5HewqDPhJtJ8tqf+ylFUTi993AVg7
pEEF3XrlRq4Jckj+l4ykTUm1w10KKzYSvrexTd+gp842+lwqx8xeMyUJ8CEvaqrwRNPqkqp0cW4v
G4U8Xl5xImVEPF1Cg63tvsqJUjmHpUQAimarqO9quW5pljhHKRmQXSj1ABqU4sAsd3dbebXhHuqc
8mO3NfTGNCsLlAUeLkXRUYgXw7D6RS5Gi4WSSkFy0foHtLtDf4Y+JORN7kjtzDZKnpPrUgozTxlQ
YkSgXXAn6RH/uLQsA84xd3FC8Ry8hrG5u2XeHmuAgikKIz47wxbuUnjQXZElz5wFnFJEuZmf3T3G
rHNI6NCKCUqBZq7nH49yFD67Yd6+RieY5EkValn9tC2dSf/559pbkzhUo1Wk1rQsC9tJvA4/VKio
jOOjFaLePdAcIZiJxel45MMWUOPufPBEPjoykLpB5ny8WkNJ5+orOGFP9UJK6nQeXxA+VTdqVPju
kjwls5fFhnHudfp/FvmygyFcvbBLc5Gpfk4k1UTK9ttPNRitJnwdVre1VLkjhcHZk0EfnNaT85Mm
n6GSdjp9WmNN5BlREbD5wiWnytz2bbAPfwUw87Le3HlpDzzJ5pj0sx+3Us5Mv98i0uvZ7B9GFztt
m4HQkTpdpr+2nlWzPeyglBhU9694EBOBUOAWlcjtx8LthQE4j/9K963GTgGDuUduCHj8avWWP1iw
7Mm+eoyjeadynrBtCVgiXCaamO0cnd6IqJj6kT0gLAVb+quO8VNPQd9lZE05yH2N7CZcTiCn0Mn6
v0IrwTbXWvnxQhyOx8g16QvnO+d6kd21wKiYY8eaQyiA9jSxt5QgVYqxuHvlmzUfcWPjUKsvO9Xi
VuAi2RBNKIIn/TMO/Ns1CrVxYfjmhc6fBprcc0icdveMD9Gprv8jcWI62r10kgbUAKMU9kVg6ZAL
SMbdu+TIF0bJWoNhNxH3CjPl6GMozR6Q7e5k/DLey87OxauLHOz65CK0iP/ifqpGuJJu05kCx7wB
BCjKZaaUoIBnyWKBXzhReG2POXqib/Fkrjyhw1JZiqQq2Sz8eB5VO5mKwMK1m/7ux7L5UbnI9SHk
Oxpk2b/I6xfkQTgTCNoy3NI2DpeVva9wRz7pVMxNM2MgXGz578h62ylA1B4sI/npqBZGqQ0Rgz/j
s6IuiJc/3dYMdmGQGySUR+xuCYaS6WvHjjMYUSwn1LUCpBsAgcSnOhMoTl1bV2rQoDIHk6KWsCi6
wQRY0va2jMpd/qRyfU5VoEi7TQd4C8RIlta+q0scY97FL3ZEzPqVdaxVon5X3shGqmV5uMaLHAQU
sZooU99ek7D+1RpNUmFTjEfZ69f6FdlfDUttc11Bt8ttShzI/RXMaljSmpomQqANLbXtTazS6+Tt
jo3kA3Gep71RScZdwbGeku4dyI9mGLHSVreVHzxVyto2aZhMruppjnawmViXynRgyFhlVj/lUOjI
MKgjZzU9MCigfOpyMCyQ23bn1CdvaHcH3LdnwdfE29szp6lxuFpj+/tYHPjfrOgkSAsdDXedh0mP
ZqV9L554vBDah2DxB7PUdXQpM+v4LqXQuR0qbZhN7b1jqqlloTiBjRRnXD1xDK1FKojsE42mLE8p
4YFZ8yCWxsin9FBIUDyFOFRsovrXs0TeeHu9lPNmXr2NAm5uM/K+3wuAVz3lwpREVs2ePvDDoBBn
GBnjfDdt56990koVCBQsqg0x+X/OZx0PfepqHJgrKIZNs0ZrO9FmLH2VAIFHPOTUGHh15TCwripm
05vvrVNg9OIak8srPeX5S0dyXWYQEX9HnlRVehBxqWbmX8Deg72oXqKHnu9Afm46VUQhZOs+wbz2
5SMrIjmOZSL1VUykzZrfb48jeKB/Y+6exivsGI5ZUCHFwchrT5adeP/QQvnDHVt6tV8M9BVgEL0N
iCkYulzKyXcWLk0xD7hMVo4KPdGmEkZXyYpeu1J3y+bJ13kvwVrwc2QikYovQOz7T9xT7vMHe+dE
84CkP5Qzje+L7Lu12PGiLpjxRY+xpVnj7IR0Fe3/n4fTRpQqCaOnFJ+QsVORwWaHScAzmb1vvfKj
m+U+oVbBNPCT93iaGYLU8EvSmnVqIt4YogegfEG0SzoVE7UZn8NXiTId3uVTtJ+PgedYtd6Mui5v
2xrG00qOUfGbMTVbWf0ri/VaBlA23ROkXTSfOAD5VjBcdEIyEmLjoGYvbVwQ94TcPvMWo9nxgslC
luARpyhMCw0W8d+ZBwnC0G26lhQly+zNruBMlpS9v7Gy225DlWdinB56AlV/h2DkRE4S35FH3Db1
ftUPbaYyeBLL38MjuoAc4D5EqxaeUOvlVM5PzwSskBuUysLPSy9iL4HOH7bccaYmKliAkmG+kFuh
LwsBaQZYKZwlWUwPhW4GRXV8MSs/Wumfatdhvg1X7occ3MslwB1sPMZPCaja8JBih3jTxApAPtLg
x69LUomcgLEoxVsgdAJ+C4dNNf3hv2Wl2gnqKe3tJjW1dq4yqstDVR8Pq+cS0cRZRYKk0ocriRQD
9HzQV8GQYZ3r/7bgAU2KMBkZ5a2b9Ho6e3kc4S1e8kWenciNZLeg5NOt4Pw7SZO31xjF/fjHu9fX
OWqwDWdQatLBQMsd9BcoHA6iljEsU2AZZZpHUvRzqoZa6rg312hgT+jjRZgVThhwLe3vKKkFz/zr
+jiZhTudHUVYEcQpM6g7Kxj4gitKBa+szqwEbb/15DXceZZ/UO6uCNQ5QnR+UnQcODpeMMfSsyih
ypmrlz1hoiaiIYTuv3cpsALcxn0OcDlwMZi0XD7uRaJ3mIHlU5ocRc21sHLRS0Dq/tjCv0Xs7Owt
grBveK/cYVpgE5SnUIs7MW+AycQvDmWZw7xmlIW5/cSN7zasslQBkZbDIl1rI+NCff6yQBdIQN/T
IGyw0mURr6JFxUH9XlzrCxBUrRZeRKzaYirJA7hcUPp5BKRatR7Ym472kB2JtCRNn8fFSKFaA2JE
WBN7FxPfPFIagE1jIj2Y5PAkgMGzr1aWYYayHGSfseLsApyf4LXwJ69zGTbh4D72xFs1dRDQtxex
xpXVZjfsnLZE6JJdwge6S+5b0bS8Y8iS14e7s8wITUz6Tg/aTRG0K6Jp0RHkQhR9JHVSkyGDqi7p
LyLhkwj2/55DSZ+AkZSeXtfZcblKJZF4pvlnG2Dm/afFGTiWTYSb3rdQjkZ1dwpky7CISqFPMhSP
F9qoKHt+uD6oTXZfb1XWq8IAo9JUqFkFn3QFRoWFcYyPOrxlXeT9dBX/7ssoEkrdlqG4wLLxeSR4
M4twEirZGrQJJ0SEEhz9L65ZOJnQhGLD/axVvnLcnHUvy4OvPf3nzZisHL1fAn8GK8O9OP2692Tp
wd50Ke8gQpGrILknvysqWjwai8+F4cBXgaLqfR5wjHrQV0fjSSSK29xQwZ7NVvhl8n0r8lesv4/G
ZQrDvWaAh6DAnmbH+oprWtZu0VvTrXH9Oaj5KurYWSpfwMwhWJm4jFsSm3UL4Eltof0XIxdGYzBw
ROs8Rq5Z8ru1kqrH3Y4qToJwlvAGFAPu/6zNluZH+RPC5vLZKe83U8UAzr5wjpeFFraFrTsprkvC
4ttfo8I4kK0uOIMlS7q8WbT1aS7LzQ5xXdLkvtt8ApUveN+5FQL80JBjuAXTwn/TGzL3ySRKXE8F
J3tCK/aNaoBxTQDSGL68PaaDFgTo9vF1rlCa2XcMbMvL3G1lSlnpTwipcWARJ4OisM7fGI2Cleta
aBaN3k0WFZwdwtpvQjjF1lYtkZv+Yy/eTmQgxa5HRrQ81coTmvvbgBPFw5uesPx2CNRpVKyGFywx
1NF7XK4ZfGnJhWQaxr1VdAohEiWD0O4dYAilKm1Rv5zR0FzhRigRJznD5Z3IPsHbThIhR7TolO+R
iDmykusSHOP3VGTJslS8pYUo4ruSky+6Eu7Ny1O+AV3Hhdn/47p3VdzPdDyjV6XU14rxsebooiKY
wdjCP2+Frxe9ca2cSufwKxS8ZEI6OR6S2vpHqssI1EykgL3N1mVCK18ApKRut1tto9zDFewe3/v5
eNzDup56UhVvSuiSrYUlRS5q15TQkAwOH71qHZAmsNZpK3WyBaharBbOAebFTbKAVgWPTImErX0W
UdUI1CrA5KRzOAB2u7u4ENlq774n8uVoWIl1+Kt0v2lHH30PaTdAOOGTO966b9z/bYmr1Rd6tr/C
i3P1+nzM1hvchfpOR4PfsLjROmGAM8q2UxuzoCqD2YR+l0ne0gtwpIOjdlZ2Zb0sA/6ZJYmBh2VL
G/wMoAaOABnqzMUor6ioSbC+CBfTyFo9rNVVm439JX8XhFNxWDd0DkmpezgNjLLkylM0d96EJqj2
shciY+lnRpjmFJchJP0+pfghyrize/h+eC4/0cbw1N6XhbDbInSOcG/QGvCdyTGZrChRVRmn6KJc
A21raXGgyLa+aB7TqVCNy3VstNHmCBeqYPdyLZYLHHaK7DkWUHIege5e5ocAB8NmTMXm0m9qmoSL
9pVv9speVI8NuN3xTF0V3eOCxn4iR0qH6hERZOAVnCj/vprQJGC03gMThtMKWMrS42yo6bgndSpF
ID7tldjS02tYPP+kK/S6eVCBRwyDrrKjxsOWfIXnp6AkvUydXcU4nvuYZy6LxUtfsbZYN8+B4hO6
JQTXHxrq4Vsh2PZPAu9CwCh30UsEwO9fKDIOXyL0+IlMgdI8Bzafs5vTPQXkvV3bh2fSBP5EMD4Z
SPvs1k2o7w/0WJU5uympny/pbc3eXh0oLf3SYM8bwbolrvfbIOCYXqffbANMVB8jUYxffyWA6UoQ
GjRBLCNX1SzAqrAPipAgMPcaQlt0dIUe9bGYVbLu8skWW9IJs9cf7nlpjC+UuE61Oxck3oEj+NKw
5xFL7ZiuoJYMWwLMjFVizcO8tmFbW/U9Vk3sZf4aivn6/O/FIb827uih+ih9uFUlKMLRdooXnRjD
Dw76OJOW0Ip9qLw4oOWn955ZZDHbwjiQuSeJi2skWapwHRMjiQ5hOG7eVPvIAqKHmchg184It1+M
rSGjyjPNTGNlkGTJxby5Njhhh+f1OtV/wxHqtcLzobHZ8HLiJOlAlmIcAqzvmVRrMl2kS5hAF1/z
pSGr0XmI7xPXxI840nYZ2VzQBKgu46lL5H/vNP+517ip620gv4K+STKOuvI0bOwA/b15zpNfThAJ
OEZIf/7QxKUYX51Y8wpLvcZ7SBeD5fhTiwVaEDhPj6Vnan/qR++8M8YHvPyYi8C4xaqMcZa5k850
EqDA1VGai8XRuKOmtzNxr55v+y9KRAkG6Ebc51XQZr+jb3YWwu0ZHXKyC/pN1ld8J9ZuM20GGabg
7sxRFD5ZXrV6qsyJJedEEnTWMJ/eJcduN+wA/hDCXWuG33a9kdRc6QyS5eh5q4ZEL2iYjzzFp/Z6
ezhSJ8gnBfSGUX0pG3EtCZymGTM4HBuye0t+V5jJt8nOtJubLIoJDYbY1hpq9IS80HfracMdbgfS
9Jcd3dAeJQ8Fycf8hi7H3W1xUmoQ+1v0ufgt3jGaU4JCBFud0CsAGBUEYdj2odcudJv/HuSDKTwu
xvNBUKGVXiZNBcOpjUHN6LqanJtQ1Xlr30RQ6skE3NPRfrigMyqxQcx/bWNOcahkdYaDNDDgqWth
MxI6j+g0HeQ7ln78RWt9HKpNaqFvhFNlzbdST2xZ9BC+MJDSsIm8LEv/p/zrnlFCP07WuwhJHtEH
DfV4WyHwr/5I2swQETj1RA9smlRJmoBBuMKXz/KVwhdavBiMDEuFoYJOn0bdYkhy9++VMQhJRprg
i1KgUYYo5a5zAXa2vbGiHkikVzvEbuoASGUi8bi6BnCBfQeP/cc3PuZpXrirNq4nBeWlHDGtZg3r
qSQ6EXzgjkAxULv1oH6PKWlf/kqpkCBtb2po39GWpyJI+tLkeNtDmrAeqmn6HIs5EPK4WITCcCny
YNFiGvLUme51JjsVX4MGn5BQje+8R6ZiEWIqx/xK8ZXG60f7msccYIxLi/9938jQ8FCR8v1RGlIL
SOIPgcAQIQwOnJoZuPu+/LIVxKH2710BTtiLzLDD1xMwWk9WxV7zgkTn6MWJgbB9KytBV8LquQPi
Fos9HdaI9Vv3Kxtv77RZlet4fFHPpcHUXfPSItiAVnKRYMJZQcgNpBuCIcgK3mEhEqIAglvkrqT4
fz8nLc19HfDLzFDJ+G49MoePmazGj2pq4CfpYPoUMHv9chsSN2EDJk5/3zejxrYVTNZgGpOJ06Od
jBQIzGDaM7GbekLxJZ5NESb2uqmoWBZZg9AxRrBr7uPEOheI34jJtsZPz6C3JgRe4X3L4C5QMJRy
Q+jVaiQ80zcPodKgbPppaoynWivZVG0OmLqRUsN/4Qnh71wtnN5ZZ2ZhKA8+a7VO4HfG6RTlpyDw
RiVzauI/Xi2YiJ5177WznCBJAWhDC+yVmpBpmbyoTry8z6ufzVjzSlBe5yA1VAWQSzvR3DRCIKfn
Oxg2l2++PF1NFggIxxmcVWwetDy5e0UYBjh+JU95udGtH23AmZ25Sm24rfxLWyVyO8k97rXeWmTB
aJb/jd68Nj1NMGgVgUaMDFfiRYm4PpzpCVRa2/5jOeZJReSb4H1NNnFl5Q/W3QflwKg41EIMf+9r
+ZNFmpzwblZzoWbDqjCtfzH8Q3oeJN4UzoOfpn1AOsaDgFNqppY58Q5CbRY6m3OWJ99KkqAsR9iN
u21EqMMFf7LYUat9/ViDqsBhwqeMpxJQGx+DDglk98eb9FPgB8YTT9UplxK5z15ntGIK1lRqv3jI
wDstQCu7SBDBdbJdbCKphtmbkuwvqFpysR2z7S/UxuFG8rYF7PGWcTqGi4Mb309wZSWyLPN87Den
/dgzanlTz+KBXz0EtVMjgNu55tLli9iw46Az5TXoxrETQ+P7AnOMmoPo2np4am5MKh2DiGT6yBZF
axGgiEraxvXieNpcTC7tBUGoXwgt0OGRwj4VFASb+1SWld08sYAd5V8+JGFWVyJrulXRQmbhpgja
ocaswK/zEnJ6G7IXEE8UzGyc1/i98UgX/NVM1cIdV+cG1juppDOTHXQH9pf1Uwte6GsPHy8yvcAl
YwmhAIC1PYznPCQ7k5dmXg1fEtbjtNYwHs63oZV8GknW71GAGC4TDDvj5p3M4PcsGYFHFUqWLeyT
LWjfCQRAjdv2d+lSldXQeEAr5tueUxOyFZMX6oVYafPvJhGSKfQtltruCnTKWBHTfmp5/CE8kOx/
lL9g1s3jAwBLJWMp0FxIgQo6Y8ibRD5gnpMnvzoxaMA9LVERjIozbDd+5nkgv4FXcbfICPOe5K2C
8tuHWcPGkDtuoSIhv8XcNBulW+o/yTFIuTgnj9TxWgh34A9++gEs6hbrRkv9WyffmWk4cFBzHBs4
UlyeRg8yM+7i012/Yt6WOmTW+TAC+YaVJEFvsWGsDDRLe5BzpIPsweNqu6jllwfi+LRkiMfsC4b6
F6OTsDoWmZV86Qx/cOEhNoJUFi0kwRglwO7hHo1dpWJXLNvc9J5TTHetyUYLbe4npD1anlAu6g5b
gvqYUo3ELtBaS8dlBNxx1gxN8rGdeExtpS9+VPYn+5rPnGMRSRJ4fDiKhVRc/uPxEUFq3/lobrQP
EWEEKbgWjnjGmccoBExJrFLryWOjcwFq8iqG2gLX+DkONvKSC5bAq+cZK0JnF3ba1/ywuHo3EzOk
AGj7SQOX1A0Mnrs4jlYPIyu0RODIFAr87WhdWF8VUQLqEi2naWokfUXqKJYElJpHKxaFDsrLqDjs
P46ycT6lZ+FN/oH9Xe4i6eNhcIERm4gxqKA5NltuvcY8dJUI+/xvGudLtFBnSoSSrVTwWCI6rqkx
SXSqz7umldKFL17yV3YA+E/3/x5F65WlygMFK1XQUWnzmCAn4FGLo29DkuE1bdEqxP1C5X7q3sF7
A0VcGUTsb8abvmh900xXc0vN4Ir/uNMTBcwFXD8Xtqj7q9Brqe3v4TVqI9XeCjsu0OWxs9xvu+tO
vJ4cA1UqpAumcB0mvICHT2e3EF+vF80uY4FvIfB5DQTHO2QLGuxnWgAbVobvU1OnzQJI2/Kz9EBR
J9Nn9Ngcshuc9HR+hp9n7J+P2VNHI4r3Y7YdFDlXVyJOC+rFuXAVTZCxi/Y8OwjRRcBeTGqRcS3d
/ErCQQ8HM5Xwcj3HcZnr3R12y/xGf1gDJXpT1bBBmRr7EsLpTyvZERLUyj5GAc1qTp3EQ8mLE2V4
kNXPboQUnO4v9bdjrkN58nrsQ1SlCx5e3mPM3blI9rTgHBtzG+5aYLWOFRCSCgasdcf9ZS+r+fk7
MazIaTAOikzHydXsbCguJsq/si/mO+/StdE8vQ3m6zy7HQvGQmQUaqBTGHpyjXvbCWEQEjNpHsIC
KbMeo8ZU/Fq3y/YyZSQS8SlXNeaZon+ke2rtRcl79cCeiAnBZUiBUqojfQW3kh6fuhUU3fhDDz5H
cZvNgvZOFnL6sV3l6Afhk6DYbqwzb+4SWMnorjzyiLwukls+6PD7Fck4486Ks9Y03YqMpQ+8XJ5b
wCuJFSbtQx+Iz3YnFBNYgSDhu/MDzJ8PqJ+s+e568d64/PcnOXa5oOL2Bi1+vc3ZgOaBBpmG3Yis
pyXUo7GM4zgarcdCH2YOoH+CkXrZEn/rioSvilvsRSql7mJwSRbybLpLNcRhEsJCs6iEdIXn+C36
B4GsX1Xn67fV3RYIFCH0jeAmiCgOmpc8WvC38T+wuttRCVJBE737Mrn8K+byd88S70mW0r6pz+RL
OOXkc4F0z/EeKro/Wy8C/14qDr7EXzhzizHT1DUVmdpxgJG3q2d4Bgt8WMhdFhe7mILoRq5XdVsi
LivaAf7vBDBwDgoK9ms/ePFboUQFgBMz2wPjgO/6VcDXfmArtgeE32LsCivqTr+DyauUxpTMZnzm
NA5j6HvmTCAzfP5u6d95T5z5Qxd683xk5VoD0f0cjiekX7Ku8go5kGZs1h4WCfU7CYQZRl3aIQw+
HprUUJ44j+rBmmdofQVjh+PzzLoRzOK27Mz9TPanGFcSi2CqwCaHKnmkK+gzcjcs4V8l2EWceS03
oaYCvZ636RmFu/EglsnMzFu2lxP39C+05QwSpJWL3+gPwTTDGBWwMepWr0LFdp/pWl0Hevv+eA3w
oJ4bfTv10qSzMS7XVoZpfe0l4Wk6rp5XyVUwy3JhYdmc7dQ2/FJcvrUbX6DyUa2M4r+6piPQFf3Q
WVPynFBC9snvvpJG81ED3QbP8T6cGEsJyWEwTVMARQ0CpmrILTDAFTakK9R8RyaKmU5TSsTO1P7Y
N+OVBKYmtcnogy5AphabYR185xK0z4LVIjxoNyACEq5ipti2YF0CFzsZ67fDjCD2R35RQs0cWfw4
Dkw9X9AWZ6cas18GcmTmn5FvKguf7InBiH0bKXfpyijJvKJS1bXLBH2wBvQOGM+Kj5DxjmZO14sP
4we3+/CAKulQeeZXsrgfT8rVAYIkygC9a/R9PNRnbNx/eIPEQpfxGCqj0GG+uBfCfu57kJOMNAOg
yUvuhwdXlbV7pKE2QZ8/7gYrIHNPhpA/24wTXtyzlKiY0noIJ5FTjuwsuAALDWtgH8XLR1Fg3N+v
c0yTcvjZeUJj0/EotAejBnCxGlEFfR0dcrpBqQAyft7hTwGPw6Cfs2eNheYR5/avWTWnEVRnlj6E
PWKrmMvrbfZ94Dc1XYjk7rN0dmmHrSvWtshg3hOe5sK9y99XUubCuaTSgMxNU/FN6+Oskz/XKxyn
DfcsZ+kPCUXu3hF0e8wd+gEZKHtgor9FwychUkxwskISacx876k0gEzEsJjEZcReA/b3OJg8FqC2
vQq4Ru79yDnc/vqXe2d1MYeI0F27Es1FdQ95b8sLw5YfTB58pOCmz/2cXNdkGvwaffAO9KPLEoaS
Hpdm7U8IuwWXxQYJy6W9TrvCDDrUscOrxDIns2dEsFjyfUd1f8skDNN8ezYMzzETlb483GJHF5Sv
KVHmmp/z9gZt1mxuRcPz5s4KEfHbIlGVXC4tzCkt8qRwTO0/gwwD5hZLSRpONcspmVQqQUCJ2Ps2
SyWJvPtouHC6Vd5lAFTV287EbX0v0iYdFNlhjcPIlK7Y1rW8VafA2eRSOzstxyOGRLTtVqpC77Mw
lBzSVFJFPYKCRbCFNJtkZyjduMc4JuXfI0aBpWuJO+5M9S9rG5et6gwONdTeeS7B5xkf3mkbb0R9
2uMw+/bkZLBSL7pb5T9W8+KYvHjOW3zOZHPvcvFx9VTJRBn5VzI0zQ8KdDYW/YQ5OXVnNqTR98DD
VXFlwwKxc+LhTIYZQSogJN48fK4gq5ZbexVb7dwcFusMU0mSPyoYfQknUtAJOOczFuI72FA0ZGoD
JO5W0iDgIvTC+s0jY7aTYtshA3N0+uA0kLkhub6cDs+QAzWTzkLBofEazS3KENLNjewRl9UvGFAI
3uJQpK7yU+063zkmEnLUfUgi3jKpDibroWYn8+jIqquJuVjo4W0qKTwUapP4ZLncc8JyzD/OcfAw
BKcfc/+Iw/gUM5/7wHw27zPmNewIkFKn+pX2wvWd6At0cuXqZOs8sfkNiUbkLEMDHb1P0+bfDgiv
a8LDoTdnWeOipCR8d8s8eK948XzN3ZpbBRR7qz7OStdQ8RKJpwkK2+3nV82QPjdLAkOO6FMXgSIp
7maA97Vby+nD59myIkrofxrU5KjK2zO9AJZ9ecj+kVrTVELgnzWSJofh9OpDzs75uia7r3C36wVq
MDOUxgWE+gzk4E7AoXLcwpUbRnmQcawu7v2+9N0qsoo49mRijiz97a144O9F1rMZ7X09otfaNuMo
XVRHVtIGJq1TiUg/+ayM7auK6mClUCgeiGoY+Ncs9lrqWjo+iX1QyBHdDtpUdXFxMRWn3rvrOd6N
conqCaCHXh8r7f2bgNX0QacUsBiz0iQ9dxm1vCOQOkXsEB1SvClPmIlxG9a2RY9fd7dW3usWPcCU
IHXwDfZCX1UZE2qY6vdUbQ47KTCAZlU7DqmYHDDJ6Qa5bm1jVzzJC2fGIJlds4/wrjPz06NWmUvM
LiXmtWMG2qkFWnOU/zcWc04S7vuLQAEBt/MjpK4XDo6+rjKgpHpHDzjID6CDxwa2CPOtbVhgT2yX
37Beuzyjgb91FMdvm85lVLN2BMVlJfGLD3/1Pxl8Bq/VhpMsG4EwbIp80ZPsPxeYLl8fBBeiN8Uw
gEj9HSxZvwrgh0Qy8enFwB4xDBVWnOkOlm21oNbgUyqy5Wk+fXriM/RNe/NiwjMTq4MFxjk++eRw
tAj81w1xXAyhV+KFPUqm0qk4fIIQPWPaQ43ATGaZUFgQbXqp9Xa0hMFRFji4W4nfvXdgjzNdZkzz
xevZ9CGTFHEp0nRdDoHfJIR0v7IwrWi3bs3hu1jzAf+MgbBMzuAdubwptRjzfhMoq4rKQ0g45SGf
YdSP5zB9WAr15cmoEFIaHHugg3EdOWGAWZILSSRwtZB2Dwyqa5vTnnCARFby9Ijr5a5VoSWcE/UH
IpMHXopZoTOMbCilUb4Tov5IWtUQRwKzm1mjoyIfaceZ8pdzMEoR92qUZ7UaDLOZKaLvBE/2H+1n
ScGY0f6ck9JdkLqclLjpBAf6Yh2dIBCvpDbUXAT0fF7a7Xa4JVwWLbACqx9li8P7F/MnWpu49oI6
oNFrLUm7UCgwKkcgzMGEOnS4NwpK7G+SCgy26dotk4aaIYZx1TCSx+mWJkyqNK4Qhhs4i8skQFie
C22HngWuXUAa3Rmm7CPTf9BwQrOcSqMJq0g1yndhxttH5P8mHAzSDa7aWQVlbFB6zhsfyPFJybqf
w+yiHpwRas50Y6QwPZuhgslpnUgU7M7hOGqd0gmISNGr3bEhza6H1KwLyormdTtZi3Hbojkcwh2Y
+N/BBNh1nPNPbrUYqEbsmrP/tYjAYBivs0rLuPy9ONd3Z6K6DgAyveU6EUHin86xLd8qosfjSuTW
Mf9qBaVjRWu33hNpIRsbuuNZ2y7JaGmEbTv+mKnADIAxT2kDLAn7V/Ekh+jD97QebjnLsDr77aPv
7VI1/7xCIEwSZFn+o2fBthotfXo4h7dfE9suZoxYQrrP8GhgZ4e5c1qMB1qjDwDvivVPibQNPnt6
EJwUmrW431ko0oDvQEknqwjtMjO+3iCAmWjAmHyI6gF4FqGbAeAHhK1yND5PFo7/kJqpUHNjXHJg
jMQuiC6zBTg23PKYT+TeobQYutX/GGVVMOzESlrw12/u3l4/koNafKFJ+Z3xlr5kLOuqePoZsLu6
e+mmX2YZJWKkmE8Kl601xehxGwXO0Jy/SNR2xpYACeefS3qXeDzYyKOuqPMOoaOun4wCBNrJp81G
Cw2aVwdXLLFP/ZbDHN45RFRAYmMpFfyZ4tIBSYEgtQ9RFae1FuuBwz+K+ys0KhCSMrI1WsZWLpX1
wN/NdpSw6ka5DTnXb7YB9KR+Lhvjd2nMpk5ndVgdEIsc5Hbe5/62XdukD325NW4BCm4MTGxGipGX
QVlXCBl1auuucOSlL787yG6Di/5TnVXAmJ2m64POHc1R/cl9Sl9YAH8vdj6bYv7w1xydOpsud7JP
VoSIuwCZyFfHtwu6uNn/UlhF8W7MXy51wmTFXwOvxY0Jz+Vfc5iD+WveVRWpHLKMdlp5VSiYn+3a
VCCY9yE0Gm+h/UCiZuDpiiKNOx+apk4G0PJsUksrGPT4A7W2d7LlDy9DLfRGK303O17koLmsbt0H
yrEQGQ4kt2xwdzD4MmomcminKczQxkQVullrWet/Jl88/1b4YdT1/DqtVhldKBthJPoichCkq3Jx
OcApGY+Q7ULGjzj5uayktuf+FzAi0M87fDT//E24tyivF2KdGqIOVZR249wNm+gsOkt0CpBaW6GO
dUnokLtitEODIHgYz7iLzbub9H51cF9m6lata/u7DDv5rImGEDUch+wB2lpr8NSjMStMwW4Do2O0
urvys08ba1nE9phREMQgGAx7tzzW+IalUld/mIYVjsu96r6kJXABQGPzFz0Y3UWkfeKSMKQUnQ+3
tHnRE+q1Pmgy4oGzbBNz+eCaxJJUAMKa67Vk+h8i/ZTgIwwuB0gnoZETHVcKyGwvMQvMsvaICGNr
AGbvnZWHjdN3+fGz1KEIy7Er3ZmTtpC/s6tiTuYoNhBmFvopRY7NvJbrstIYI5v9TOYTWGrhvJHd
rr1lmCwOD/bPQx+IVZV2/VSZW3YNQ8wF7KKsxLyPIBl0+fGngK2EbuZlvcBQ2fTUP8VqVcROW16f
cqa29qRNvqdiIWRdxYryrR/ek33luwTCOYjtNSsA4LPnQkuDdY1I36V1Cz+Pu9pjmtZrkAw6L/oM
8L48L4gVZKcDAlXNzJfcQ6lBcNZBkSFai+rWsh4X4nLObpmM3FBUEfhUtsQTpebh5tV3aD77mbvd
1gYOpU7XkpPOtEPWnJ9mw1djAddXn84y4IYpwFF4MC5I/fx4J8WO5STp3frzHBrgzzyvvngbaudz
8cgU7ACi7HiXHeg0HbkEQX3voZ+tLwM905pigt05EHzplTKvkVsX/0fT/8VMKI/OppPp2kfa4rPF
jvporXbniyhunBhn1r8/c1ot1pKCNDupBuOuQY9w0bLPMGPjev0kRRlu1X/UgaxzwQ4sDpp8IF1r
O32kc6drZsHN4rQmfgb/0dtD8H0dCyMOPSfzL9PMdJbyja9BeMrM8vuLa2rBfo8EjLEPENFOscmC
zHi0hL6vRRPtnsp0rY2Os62jCk69E2Jle/EUNqVfP8yvNx+XYBNBEtxBbL+67jgHD8JVwvzhWPBJ
A6KtKPUTolnuCF0eZ2UDaWgYiB8uOmIoaKhjgf3jDw7Ut4N5lVlmiceyIwZfMtsYtxE1ghI1lSmR
YoAQ4WvG5XcLeZxX87Z6ESUwn9OQWU1eho5YDoafQpVg2Hx8scka2JvgMTy6crBcMYEa8x6fwo1x
6Xo30fFhaBswJluCdcf1Nis8ochtuY00Vx+gtwDr+/gPruOo+1WKisIYONJRAfv85Ae02nTV/z/m
lvPBqVJQ8xr15WdxX8syLG32+XT+gdsBOUSb6Y+jbT7I1mjDtUxpOnChL4mKhLtsN50ehB1rHyKQ
p/QxoLTNrF0nBt+jg/OPDfg0iRG/04OEjkZiV9ckGP1P+mDxp4jNeLPSKLVbTzIwrgKYxne1buP7
USTsMvH2n9Tk1IGLNFViiOUEg3D5l86IYe9rsLkGSPv3LzzXi0W+ob8XtVI8X5UVGtujJ30NjlUN
sky2V/yq+jT5EpD4aYB1JRI+xYJRMl2kur1iL788RM8pNZr9dvC5cGxGslNhULSrRjdAGoMzfWnB
RwYa8i9EEJzkAfdmhRsrnoCfKbuAbiCqZTb5cxE6X8tXbkLIztIu37nH04Rx0Ku83G9PXvxy0T1I
fCDpQi1siJfBpUwNNYQL6QCqjyTpOyp428QenXde93SeR/LC6uU86Vem9UMrr+kOVK/mPqR7olUU
gXARFp7Xq6O0VzwCYMvV7qlaXNFWx0vgU3zRtbvBGHK9/qlFt1VfwGQLbaubr4A75rWcaH0g3L72
TRAIg53R6RTVI21T/dr6kTjR0TYs/prZvDcSocFNMCgJwto5pztZgtkaSBibsmQPaXASoJB3PnJa
FwiHTvfW1NDAgpmS7IgZpJd3JekriOR8oXiRwez5NyGySfiz2bxwiw0vcQWs/NfkU9/sY49JWfPY
BP5wNfE6DqTtlSs8Sol5coF4/RELaV1FFYbboBpWHXV6a2Ymv8YsPOWu7jOHSdAR/RbHUDis+fYX
wjTO1RHF5moMfacQrL+Uy4QPhfKZKioSF5doto9luy9AI1FV7T3IGcuiRsz2/2CBD9sjdp306qcr
C/m/7aMKANRgH0vQq2gWd865oOsPIg8C4D5NBxiwCXazdAi1CQcXHiTYTbb3JHqofvjZqO+gXm7n
tscmjnplFpmYq+TiUpTvJzombx49x0icoGVPtj9iStAeJUSesBJFaEToMJfz97Gq4zqPh3mMkmv4
62WT4MzBXxzx38hFcifxLeBSwtqaqvpKAngOovUhWoxWaeIQ307SQUUaowM893c8goLL/5pwZB87
Av2Wgr3JDN3fLitrXnCKjlmnDBZZM+3U51D8eRaLajtc0WCyWNdyuHqBmvokzR7sRIVnzZOuZeRz
LEr4RDM0sqN4k9txvIzrNXF9LhSLG9araQaNvKKAsO/H+Bu1ZcoKZFw4bVbCddB8VvMCRO+noanM
1hVLPKGK5+1fF6qb71QbmPUZTnqoI1w4yg9HkyacUSvfA9epwZQ+aJrScWAj/2s/dOXxQm1g9ZYL
io89aX3AqNXN6F3eG0FfgSYymRlsZBmldZQQ7EWXVG3zksc2lDOyabtNWgO6+6fhckYzHMIyeMNG
oupAshcc0jlEZV30ifbU+q5H6FY0OW3tsTL2ZUmh2C+IAUQ6k8j+tu1xFec1e/9ABiPDThHQ6X4B
+DQn8/ogthBIhCQdfescz7urod9Jxrhr7YkSe1FKH+IRAQ0pG6Q1KPjLFTBuiRM2f0cAeFZZOwEZ
a9mkUvUF/bpDRjKWmk+0emxyMwVchNAdVQrH2EnSszzZ11C0YL76pWPpabc2msbpPkWFbhMrFG0G
oxxMWo5Jcah/RNUR7PVImvHuxfwHTluyGLmKQhpHn5qfqqxRso8ZpdjAufTrMEUcf9qi49lDn9LU
mxcabnguAgXWUWf014am52VpnMPADZhu+WIufj5U6SAsW0/Ya4YA3oHB5TSNfbIkodqmD/ZmTfxa
S/yO5QQjCff0+kluT4BSPTzQnajjdrLRvPWqm/wQwtYN0FezuA6Y3hWTSLnsJd3luIVQxiGVV5rM
wZoGY76uyHmfBDr/x9ZQXWJFMfGj2CXg5HFolLnVwFO3bqPBu7e+w4zw6fUz+empTFd7BCR+SxBt
bmCJaBIMA5/9rpWuPF3bQjXMzzkI+b0fDw0cpo9FpKPAwOgatDTD/byMNfCGL1J2FXC4uEdCk8XU
zHVZ4rIFzUS+iFKh8QdeE1K1kFWE32EjOTfxwMq+VvUiz60EA6c7qfgP1sqmU4zqk64LjfKsapeM
UAWR+uf7TlJXXZZn5Ftlz5AYZFG3ro8kkQkKqCDpiFTrHlOs8JxKJIGlXyOAWGH+D+3iiPpSiiN9
4upGXsG2qbXkQPrN+rGxy6IkTH1N+M61mWfjqJvBn5f3K2f3fiZZ1BQUNOnuPwRY8TDrmtey0RZ3
RDefw9a6Wc7QCuIxrGlvsU+efvFQuDFHD2i1sJZEImzz/5KjWpH/GGJ63K+Ohk7FbQQyrrG9eWNH
LFmijo3QAHxBrfJGKgN+creVXneXaavga9ztOTYUMsH8wcgMRAbspAeG0he4KINR5FqezA6Uf3xn
l1TSRX8vkLXcKSJmWwV04LXnANidVC0Q8UQwFkXePK8XHxPWmqASMQS/eDLM2Z3nQjH/C7GbZZ1u
MyPEvKSpGf83WMoHnwUWU15x1+RUSVtRV1ZnCQcl07wP0aCc+3t/26qcqTt77OMj7YRwhLUvyWJn
cVHaZSiljGFzlNjF4ToXiIGDO2LO9vGAdgpTzrJgc0sssjO46lz753mGfcWT45VInRAFWMyQ7srs
RYDhYBQQ1UV/VQLWB2bsqhggpxskJTWxLen3TQnQRJl6B4xB0RqB2WU8jSDJYfWH2oXBnhOq6xPT
E5t3cV02FFFxKciGAy2cPjq62UF8lBebkx+4bUXbKGqh7lqpHzCerYonPcv5pTQXxFgILVgtA2hG
cIPbC+EleWQBHr6Z9NGdq351uf51inG2DVwY6vtIK/khExNzI/QzQuTfOVA1FuwjSlQlrSIQsIUz
erHmD5hb9i/qFTzLBkSRuqbljyC9smHu3vZGeVp5qLZk1st5/HSREmHTzv4KrChbd3S7ZP4bi+nM
2mBCOCVLIYqBoYV6WPNEroTM+hKd6jpSNrboahN8NHgGImsUDMdQYjK5+kn5DoZfQMUL0iT4S/kL
2DxHyILTTwrDPxYVbHe1JxWkuYQJ1L1G8Y4JPepdGnP2MWxvG2XNmUtNyC7priK+3xq454uXhfBT
FgOe845w0f3cLf70c2qYlb+xNMD0QBOVvhSES3H2JnwyprykvF6HTExn+ouAmzs3P1FwH0c4gRy7
qzwbqcgLBiwttHfQJmXO7lEUXTKJrtedlc/oIH5k9O8rfK5peNoAewOHsFlc0LQC4NtMud+hV43Z
IQw4+/RyxIwikTl0kiU0G0M+PMXjLRYQ243LfGSq4niq4SwvQH2KBHs/R0GMFqWcrpjB41Rae8FB
X1B/fcKSeLQyxWCSRVMPqGXAsN5KJcJ0imo/ijuqJx1bVv0rItB8Fc2TVrDHhoUzIak8/2LxrCQE
FchBU0LMOihOq50ktaVqEcDoAibs765eMqs6ZWp2dPpuz3PRRDdtbDONPNnqUnA2A003Equdb11G
g1xaSU+7RD3SJ/MGokf5mLLq+BA6E2wCAzl8BSoxi0fRIZhp8eIqNtc+NhUJSr2z+zCtHYeXbdzT
fl0kYFUF1LgD/QVdWpO/BngRAgnz/8Uv5xoeYcM0CEMTDWeBB+McTcxljtU3cqPGI9BzdAgq5QoE
M/vhZ7NjGA9kw7qPjbzb2JQndtwJhrn4fU7WZ1TfZlxc8wBcn1ri6hje6HWqImuizm9+CAyVucpC
awwwdOyuCLKbE5rkqoAFrNboFD9n/Ox79bk1jiBRfKQbn40UBLsucUI26VdhVVpPSIhK4zdVmFvE
U7mSRhmF3/Su0imWLcMXRJQBkzdL5J1Yg72fOqbxxeW7oo986W2F+qRmONqTJ2ThSrdRb/2k1WCI
qR0jrnWFAGMmdyU52q95JO93T4nxlmr1WbapjgkLc8Un0EKTBYNU0ODqKFRjfaxVRMACK5lN7aX3
i2m+bEocREYi6EHVBAzCvYSFddqlrM4cwX+qML98m3zuI9FLrumsdqq707oD1X7jfaKiav1NPNyQ
m0Q+MNq+MBI1o1hRM14AifUVhO0uqmD3p8WmzfRifAYFkM0xPGd9IavohuQximAY3l1bIV4bT/up
qt6Ig6VfQl3vb48unJW2nXWphX+nXHRAGXXy/LL9J/CrvPvqMDYaTefe1xboxdLDzhVo9kkjl/Nf
O9e8wneWKU6apxDHYqRYR0hZkyNMnKYQP4bFb1zDCcUyKhBvT/RyL6j2WUmphwfx0lBYrxgVvGvU
+qCeh8s1lZ3AP+7teiA0BjFWpYEjrFKDY08DDfwio48Npmiew1IVJ744SVeCOgy0nrqi4fFTa4AS
SOlYAKEcR8D2i6ZaV/tEMjwlgb9EFvQNDAVzXFEIOF6bXuQYL0fEeoYfo+JgNw2WGy+rhHSSIQ6J
kWP37jHEZAyerO7X23EcFEGA4rITH5PAuJhdJ99P7pavZw43ITfxX39TEfHsbpQJPNy/tdJWj/GZ
4qVXEQl7kTSDTOjE9sd28ULpVIhYgbtFDcJuq3YfaAtVME1Owg4QTM6rVM/WmroUj9lCnxo5M5wi
e3+mK9A/F4g63wvrJBjLuHkff9K7UIfuCOLNJsI/wx10amdGOoe79tnClnGH8Qa1fEq34Kn/0Kyk
zb7HDg40iHydgg9cX2B9NfyldocPFxnHA3UbH25uMgDHqZ739Ywf+swH5pNHt9xRgOlr0XALmbf5
sPWvvrZzjCxrDBE/eH0m2VVXxQjdU9ipEC1MemIxWqQRGtaefrUMVd/6Z6hDcENT3gbAYFQeTpHM
mhup5FXw9oVWoYiG3DzRALJIbq09iUuA5F6gK7YFFR9POHKZ8wRbBilWMmutZV6asw6PBriXoK3P
XBOfruKYkuSMAfgU4qp5v8amiG0gmHMDIE/9M9XcGwNCMIatUn7Mfz43uiu8qES6dxrU9z0AsEuo
72hZPVZyRfTw5AegTpCjKA6EvHBiPVABWVhVxx/x81gsdYN2CTRVFiDTre5cXqlYkyaFd1Dt3gVy
PizTxa/9JhYObV8zWOwIJONiqDLEW5zSe306F6t3b13w4+KCEbKc6W8UD/hyqcs9kk5Jq1ujigJj
fsoZFuuUnAgTgtODY2rdR6O4VnuCgRnkZo82CgRR0utPwKIiXtWRk7iN1XsEY4M/UeLDeHx3pRNR
vZqDxpuUJev3CHJJyzHZI7bkHlErbq5X/1dATNT8WxOFLm4JBb1VtdMmweXuRNUpWQtSZZdRFMHc
s85k+d/amhHj/Mhoia4lkY/3ypRfRflcGHurw0ccTe/bK3nDU+2k3MXEaqnPh7M1c3F/k+nJsxjX
65qNm6d3Df547HImLIwYbgycA3PZhmQ/O/buaVPzt6oDb+0OkkwE9mz2a64rgJeBrvkHZHuw4qKq
ArP8T7fUh0i1Sbm2oxqXoQ2Al4gtC8w2QpukWg3HZxN5DhRW8pCTgJtr4kFHDuavu07UOBFye07s
+eGn54d6raaqekW2rhcAuR30DvbysrlJPeJ8EEK8PvuDZSEYAbs/PJOiv15JOAAHhO4DN+qJ2v2v
G35d2s1J1vtTN5iDJMkRowoNiN8TlyCOCoIzNv2vRrNTO8XFhRdHIbEyGvDNxlE/eng95SZ4T9pK
3gulD3i4xTuMEoGXi1acq1DXmDD7qBCuLZ4JRKQq1oS7gc3nALyZXbAwSScDNapsN9QFUnOj2Fmk
yagDE0ACG+gMGYTouVrfyJfrYe/RMvPrsvpa7DWUJKxecZZRSW4p4kuRLU9EliuOokAUwTls4fQ2
3SP7pzTORI09RCVMoqHL46UQ1d6SdurXk3Zt4XdpT5lVLWgQlhwib2+Qf+9OiToGKOreSFCO3Ze9
ab3EDR/ouJmV05AheQnHVvDh4Mufp67NiUXRMIvHP1QWORK62L+LlZu3VSpDDjkbeh3oShfO7GX7
8klr+F4s0iZYrtBAjlY3ESYB1WdxqrfL3H38Tw0sle1WHQXmKZ1jh4mo0FoX5uM/QmD8XtViVMVU
9Z6P5wPk6s4jfT+73OW4582i4aWwJPCDyJ4na5F2HEmn25IsLGWKA0aztPATLvqdCRDjSKMn7QxZ
MSmyxX3hFrlyy3QNm//Q0qn4SPtyEVMPI8rk/zrdnSFsejfF10i0OeUUlNbURzh3DpuzYQuEbLpl
PDivD3Ypvt66F3NGyc2yt6VLETGp6nVYG8dmsoyH3FkNdEsZBDZWXs3ZENT1C12FFlLcLVW0h/KE
eIEhFYXOOh9euFmUsrRpOuDxTNiA+RJS3j3BvxCtAz6J1iGW71G8SZsesBvcS7wI5Hvgn+5wZiH3
HB9SuOd3eY4I8Yv2+yFvqjMXh8dGSH2mlaEiNhC5SNbOr2Dp7EOiKRJDZGxZRuVefNDHlw9D0sWw
l56Vp4Ve3BLtjueJdtpveN6dEY7idRNHlUm8HvSxsJg8nu9dQSwYrtPfNviFEO4NAQ2MJW0hODWf
Xf0Xge9UoeaMP7IBldTiND0Sg3gOd+zHI/TjKEv6Wnhsd3dAigG9ds3HxuYmD8re5/Dswp0wCOps
TD2i8BK86kvJ35KC1ipFmnKJU/7BU8uf47N+fwit8y/cNb78L3htmw0heBAw7yUWyrKxiiJ1dFAa
6JlC6NZ6gDEe1AhAAzIOv32lCYtlJDUWtx9X4Z8z1FRHKxVPI88rLPSgAIes+ipomwhRamph8kA3
S6IzKOrHNfRVRqf684Q17LnaTS9NGiNrw48ocvPgpJGyvuG+GNbJei/NCyRdYW6zZu9LBlfB84jL
Kgfh6X2Kkg99VFFvn9OiHMJRLDIsAP85zWjanywhwdHvBkyKT16fEsBWd67Ltl03gBIMqu5XMMyq
euwSMwy0CWhM4ValT1lWGCVN5UroAv/MOUuZ/rTpI4uPexaY6IITV+tDX04t/BHz/ElzsRnE8qaE
yuQua6LLLUfPfK51ctm45TJNFQ0r0/1/BQijjSZOwHajtL3gE24NJDM58WwoxyIwDMMH9DBPBRle
jmrqEyk8sRgb5fhM9P3J0jiVillzF/u7LLKcZYkcpDLTcpawgB60xRYHnhH+iTxZFmWwZVBRhPbn
jJmszH4dFhe8yz1GBDZORM8jLSgXqAqUrHNXcUa8BXTWHDUccUKGseNJ5lhb7kW2rTKdXpyixAzE
ZjSDBJ9tknpi9IyrMSEHk9HfVO/lvaNR4HEFb/oOjou/+WmAA+mMRGREuwSspJmOp9ouGSQ55zpM
RIqabuKYehUUWTqDv+1hbKJ4ja/IfFOeRMpr65oPOw/Qibv6NEMQX4Ha0yMbPVKXId5zx31kzK87
L1R+baQ2jcfTGRYQ76A8siKrcz520EcYyBVfpkq1hU9OfTtvgeIFA61d9NL2ViJPOEk6rUpVMvK9
J5GsAvSNrp+fGZOMEZaVICXLpCPtaVW5WVM4t5sGxS/RQ3TWUh9EGt5bKW1RzIDuMpX/y+0/jdCq
N6w2vRdFXDDCrnpMXEjrjK1d/WOQ7Goizud5GGuoklzH2a/H5oYzEQGMYEXpaRDf0j18WCs5Z+WF
qxjmZgKakh9+XFxf2k6IqvagQki7lyfOLUNyOichyh6N+pDZxoCoLjMVG1saS3h4pD9Y00oV621d
m8zSs8tZnCY9V4NHwP/5QH/kKbg4uK+wBUyEOnCxP2rP+3HpsZcnyJJOpT8oeWtj/MiL9UvJpPkP
II+J5+4fNZ+FwqrUulaa59BRi6eFjxxEBpMQG/P0PHfIH5802dOvKu1AQwErfzquSj6DvvXt1KXU
ruv6xE5aqxQej70F4OUA9wjeAaY8s+FvtR8Cf4n4IyPXgUyTkPqg2NKTy23z1/2ySk0Y2nVvQpkf
xdiFqeWjZ0NELR0JrnUdSnYHApLNzx/Ag/XlQP49Pj40AhWxxlb4Iw7sSft0jCXtx+KI17Cbu9Y5
MxNMc5DR8VFYthIiwehmxcyTpGZoL9IluzlFutXQAZaHJ+3YxrbcEPyO4UndEMVdYqpELIjcAusl
+C6HDxq5tFwgWcF0OD6lIpj5nWSc6OE5ljCjpASs+JHaKNJOmGJVfgHk3fT0fvgvRgM7nCxeS3YJ
gScbfVvM8U97yET6LWCOlhHhiescT1Ed0GXESmXLGdCuv4eirfX5xX05RSH7GdcEGFkl4yYu8evg
uV1vum8biH9+4zDFqT3Cv7Zxz1fblgRGwrPgmx1diWcKFkYuo+Xeg7PlnYvCrxf4B1X9QaqF+ouo
tu1XDCDGOSJjo7uKA9QWmng+TuBVjiAOg0ujEQDfYePtRwluI5qAHaAhQ3lGh5scf6hbu/BDRTS7
/ABYq4vm65SSYSViDu9cZemAkmwqnMdMLxaH+YJAvBZ0nnzwlOCoZmF+qnWg9NyaA6I9Hb0jxLPk
igGtSm8Xw+hNV0W8muuROPZFbwMw49PV424pRxjlH/Os3f2eQPuVwk9j2kssVohXLWo6fDqgv/BZ
+accMECbz1LSznZ+AyXOjA8fSGYt5IGmkMtd94e+8U/XRVeXnjRlFtxHtZMXddBK+d308BVVODC+
R3qoDUHsQ8eF0oT97VCTnOayLQrbosycwdnYPXzw+yu829Mkhizj/qbpBxhdlxp1hehVh2wUDu+T
6bsSVfoMIW2AtlkKa2r6EpP1DnSjqHt5EznIWBNbpqF9cRffbghND7g5lQotq5gVx40YCFjGeNv2
Gxrfgk9esoONbgb5l82Wwk1xJWB0IMNj0a952GQb0D5ObrRUxN79aIJpdl2SjnVL0IEU3lvFwhQ9
v9Ej1ss1BxFgOSy2vwqyCUW+1+5tdDveWO7vLJ5BvmkYhuHu17KuD80ZIC+5GPYfkRElD+hSRgYn
Zq2chLw/C8Dmoh+MXM+X4P20H4RIqzOHf3dXWNNvO7B6oEMskZq3TfV1tMQc5bu9WYHu5GOytsGt
5Ug3tUempIA8dWZBSIzDGkxcI3Ku4U1GRNv7/bQWI/yKrZgkqYg1o06kpBa6UrO4ym01GYLwUG/r
BIUrTImDvlYD9ys64q83pOyJNeSusEgNAH2MPpT2ACRIWcpbQzsASCC90KEgD6SNvqUeRAhKuJ/5
I2v2Dd11odsq40oYDeUNtws4AIGASCX5bwFW9FYw6+GYvexQW8KD/A71EAqKfJlVMoCGmjYw+Eh8
pQVQCAnQ3//xs5EkzZrbFeuyzvkdI/4/7jW7RYczF9F+MpXzCHSn/L0DAmYnrF/rJ+3QQ2rMYXKr
5+3qJTGdBj7AceCvKFWAnscA2275lNfQEK1CdVXcgBJ+SwF0PqRCJ5hbQOVvOToaY6C41q1tYR5T
SAC6CZp+sihDCrbR7M2FDChuoaeNQxPuLyIyFMjEc44DaCtp6mEKnc8V0rUXukDihZTbC2l6wZR0
zzTd7mN06kyA9xHTRqmmcNir+WR/QQ89lPdF/5IygKg1RFThFneOe79NXJW2EztkHSUbdq7xRsjW
ASpEw5pND4A/xbG2m9ZVFe/swQFM3Eyq4skdlSBgF4dygyC+On+85Yz3jU9pxWo+AiupF7aw0h3d
7E9uefYA9Cdic5RavR3tLS+Ti2itqRt85INm+Kf06gDuSRzAc1FiTFThwKdDIrkRiDC5nQmgS37V
89RU0jUmB0ieDReksodBD8Nm2BA9FDH3nBvuQIsPY4c+C1dXy0AC0sMsENKs5KYCVhy6k6hbUg77
T8t+jumwdOtJuSg74284ZGmwZabsy8nyr5IAX6cLpByYpsrqjrVj4n2PgXFSBR6fuD2uZglcbIfI
85TZAWa+nOqZBDtMMf4f5+M6Kj6Ta3orQxKoAc0pE9rmLe5GtP8Aqi0guxZRbqNsSyCyLyfNIPDu
UIiZMS6T16xp7wSlupHKdpm3vhzcs4TR1glRJQmJUBUbMNu7IejM+iXEQRqsJu46rElQwuyns+vr
2KGAItXpVTmeL+Cc4uDd4K/vot2dEGQlAy76Cd/eTJFuY5VCvy8huniMh8de0VrRkyCjYIGer+8t
OZ4zsqda8EWqFstOWxQDYkgIUJeCWELhJAM/gtn7gs7PrU2TCqsa1zcwMQSwiIiOzyw8+7e1mMAV
UqyJdIrs7BhWMF0UCFz74mHGt2mFWKU8mkTSHBGURwStYPxuyZwwD3yg2dlQs87s/hEq+sliU9qI
OLqE1WqTxZEsbeR2/z4geq8bOq9u5V8ZPMSI4ke2NU1gBpLgvM6uQdqfpSOwlvlPpwjOXXmA/Evo
titGjIf7FgAct2N09bfMekEGstqEvv5s3h+E/dueDv83xHaNXaQq0prk2lBAb9h7bFMqbdFmwbOM
fnv+zs8wZPeUyzjvthnds5c+35GsHSoIhglalZ8ER6AyyQYD39y1AiWyQjwRJbJDUFTqs1afPdQT
K5ghQ93EzSNywIymqZjH2Ed/4hHJ7PEPKJoXMneMNTS1quNrxG28Qt5bf2CTP7oxxn1lIbrKCc3Q
p/fPDGhYMHY9iaWM6YB5cFo+ucXB7/qgXMDRNmlKaZtSOormlSRthRXq0grADGevaOqUvQKbKBMp
B1v4SxtXrDaMf4GpmGCJ4RB5Vx4dTpf+y5NG055B0/4YOXys5Yo30RR83FFh3n6KPNCT1/WORUVV
NMcSjsx8jABu6uv/jKDzmLsUrJwGaiJnzu3H1H8GFVXHY+Op89ubiOmTRDziqBYE3oBUNKdgRUC8
KWspQX3feyKiafXbwXPdem1lZnOSInSEv16p6FBm54Zpi3ScPZ5S0v1QFd7/tLSD/Yliv2PYspWF
+u4idzBULRdCG4zHvkZfANhYPKO7VQbEuEV99omm0IVckz4fXmVqEA/G7FNMBEmaE1WgGv6ArQCh
KfAFtxWf1on35b5oW5jbUN+EVcETxT2sBjtt1ZazKa9t3OrhUYr14bvrtdOAng7/+BYWd4cWqOiD
AodE3ChfrqPzQ69kF6SVXRQ2OFRnWcz3Xh3kRgSUt+Gha/PJJFHTg6Q6fLP5P6Q7077TEa8HqVoI
Rxguym6MwU/a73gO0Lm2iIQgW76N1CzAYTAZBvOzg5Hy/tk1Str/qiik9PH14ikt9nEC9WGdj0Px
A86wp1jT6wOhXGyAfnUuM+7rg3BqgnVbXH3TGVqvEsBJ0IuWLvZR3SvZHGPyUjUdo5y1Dl1rWBBL
CNiFE3B6p5k3zrBwDiigknnNnS9Xwg0cGQKQoo4Oj6GytoROn9N5ys+JOfRwFPMoxvcukLDe3H6E
zo1puvtFojHPNdB1AKXgBaVboCKvrpgRGbZx9pkYb4iewPOk8FKaORzPL8OBnO4hRps+vZluq8gH
NvQxhCJO37CjVHHVBZ+nlS5MmDlW1SqMPW+0DQwxg8CIhD9l0tQrLhMPF4ll6Y1JX08mokFH6Y0m
GM2WlS1VtQbjvpBgfB/NhjEWNJuY63F9C8W7Zj6zDtgPrdfGNNtkla6Spz1er3KlVy4pCoE0lIUq
bd7RVshdijVGsAkxqjwlzl/EJ8/qSAzrSUtWGkxkv/8Ha4XTke4hGMJfUEgoBEk+xRpRlsOpsc6K
dqUIWC/6zIG+Fesqi1zVqcERvRsVTOI7sy86VkkOZrDKrLE40t0DAVjs6qqLnuhpWn5EspJ9kV2s
CaWn+4zpUbB0aTRFtQtUmLd3e8rcfTVJTs7RLhT6xvpKBiQbPc9a38Nh3i6I0dDRdgRavCgnxRJI
zSzhn8m7drM0Rx/V6YwzVydyRlg3bxCwiS1Ufeb+IMczgeoZTX5gJ7w4Dwrz3KG45FrwOmNDqL5Z
VSCHPT9WUqqrfhmvP5f7ORhqy7dX8Nyd0+knulSvT1RLStd4JzCakK50FFV4+BDjlHZNmP3E0G0H
l68L7YcmB0A+wg1+MO6fPnIYFKBQAG8XI4czGRudcCFM6TiTBiMs4uJnvN0WfwSxCq3rz27IX1r8
YSAEA+d1cToNtcrZugIMXWkjdZtbZ6+WLgGgJXS2Gk6vYF8rmWuRO5BgJHcwKdQA6/mvtCJyO/PW
0YZVl6kkS3P4kASHpRtAC33bNRFNDADUIG8G5DlCVMtZarlmqPefIu+WvKVL6CgidLVrDBSnzK4y
kR81EpA3CJBOAq0q66KhG/ubPeFoMXHxPUNKy37wtfuL1qYdKOsnluzMvJzS/s06OlOXOjjdnzKe
WfTo7PFNPWaP3Av9XAhK7EiPjh7HtwhXx2aGhUPMYlsjsse3D+04I/IpS+FN90yWnsJH05tkq9WE
02D11CPUxh5zo+jj+zQ3+tEY7XndWkNp9QKKNkFbUWngKQdgoXuJVRg+oGiy3Yn0W3fhH8+hUJBL
QTQBnqCLUwN3EMuzSbRunKwX7Tx5R1r7iHh0QSlJVXEuKzTzFStDo0ujWguqUmlhsX1kAxySt5Ou
I+bKsW9zE7nRUuVasD3B9zKbHl9rKzORdt+PZYcc+1eH16TGRyhEHLM508O6wJGLrZYRLt+ZeC2c
nTvusT3f/xThZohabaVgcApp+40faBONFo40O/VTFaWVCmPFAQnNygVnjWO4H66uiWvyZ17p2pFP
kXrbBjj1Dypt0ZHjJAjf/Y9sATjwp/I4H0edA+Of8DiPdgYim9g5Wjve1pCgeHFiTNTFgfV87mgV
JHs58wlX0zDQL72kjAgp85FBhtWHr1ZwQwmsk3k6Fqqx0NT9CwbeygZ49dzUGd4yy5liPbsvwNjQ
vYFHUY8O/m8yEIOaja8tXy0maHVNlKpEozp9h2kHkgX3DhRuLhuc4PAHaNHAW5WURYGEj+aonMJL
8DXObXsiAiSnkKeMLkORdqXZnQPzr05a37rbwgQLDuoE1BgPuvCUamcAYsGcbXKejS0uiuu12ht/
ARNRITM5U+iyH5TWAUnveH6qX3fTjj4X1qwIQ7tXBbIEkU/0TkyAYJSxXO7ft5Mt/w5dPnCT2w34
j2u5ZhMPfy2zTXP5R5JYOZ5u/kK9W6LKpPk+p4c/sgNolg2ZdYoY4CDMULeua7jqr8AOA/GvkOWG
Q/mm9wdfEjKYyz8xIB5KVJjjT5E/tIvoo1RoTNVkJv+lRb8vEbOMBQ6X0/tVzVGEisySNOeq1bcQ
qa/4r1KVVBV5UU2RZROcg3OmzEjsuuylobmUxzaAltyw2tlz/UZLqDjk7EDV9DQ6w2ca7tYvd+1r
NZNgXOs+K5gYvOZ2iBSoymQs6dS7n46tKLz0dn7dzu2n5tHg/75Y8hFkNwV30kfDf1ewuH+Ybqe2
G9vIKXGsiZdS3qBFcgyyQcQJdZjjL36JPkJVpy95Fmg4bad+3XV1iBCMagWV2hwNlXfqId329TmK
Vr7ua1cf+9m15BUx/Q7kGF7kGJML/I+92RgMbxYarhpWybzR0JhcZItmbhhUeuFudT8VLwLYTUix
hEPr13OL4iKSgdb7VKK0jgtK+sO0xbL9HQ6qNt47TwnCQ6FF+IfBDXpqKWs+64wPuoz5uCgRegcZ
ebLzCPQGrCnTgjPqVMNeS9kZKXlffcVOWV1vV0SigFpU+F1aXJDhKq5DVyoEBdkwqsLxiGBc9U4Z
DFkg3sSRjPS2TCXienetA05+eqzjN2dwkWxQgnYytwsc020QHN4h+Clzi0NuwHGbGsaTJnpduZJO
IJYD+GvOrsSxUKlX1E2mkdlt454BkjSrPwphXZ9VIRn2lC02lLPBIOTyDNmS2DEr5TC61M9Rudjn
pBn5Tl/wlkY4YMn/hc5A0x/Vf6JoEXQhBELB3Ku9fbQxPXsh/ijr7PtXFCUvqkOE3NrhLGSaa+hF
Yf9yfJaItvoYyRUUphnjmZBo28G5y/5/eYVyegBCR07Chi8+w2utddDNPPBoy1T81KH0+JEw1n17
w0CyD5sLkQAQoF3muxCyG983BGcho7CEK6UGcRSfpvBWl52JXm4KfEaAoDd2mDnz0eTd6GS4YHHQ
GG8ceiIQ8U6D3mML0O3g9milxr4HgvTD4q+4XEn8SqRFJEPbjiPp7ngRhzEAPoS+qDyfi6A2jzYV
Odqxnamx8RS9+J2ABesLMD5q4R9YnARpOp+3DVsp75bts5emgQcjZZu14FjhX/5d0RqbzOrNyMlE
RcAJIfggw1p8/5CauKX8Iog1EM1qtCshO76K5Xv9UtCSgUe3wm2TkAqGetwKA9jQN0qV4DL8hiQD
GTJlJ/vSHQJUjC/+N/Vt0C3xf8TyLHVzKxksBk3yUKj0I3BG+lFDDY+FQBufV05BsY/ISR1oPZGu
IkgBm8uMT/uncHHDqjyx/JoaLvHbjOdyu1hW2jpJTcByMJl6rxX1LT3lXqHgdv57qhp+xxbyHh7r
T7bjJn8DU8iOGdP6wv7PZRsA4q+FZ8Y98i56oxH98r1g7eeTwl4+Ay2yrswGrUt2z9tAGxmUwkM4
dUPnP6VFN35n7+p+n71S/9hxWQeEv6hNpTT5rFpdXhSCr13Aqoc+hxzGZhJnNQVDNE9DtRbw/GfJ
Oby7xzxMnS3pr+GMDInrdG1v+RF9gMK0txScdZHDYBP07A1XI15/yGon290/PQVYU9IpfEhgmpLX
pG34xDdN92TP4aiEHVJJt9zv8LK0Y2OELTnlowcuw2xXHsOG2crkCqbuMy105jXbGNWImJ3Wnb4x
GRGTLx4T3/vTR8RLeTYq1aJLrI7dk2AtcTHRDvhXQlGx0eStHxm2VL2lHSr+kHpTJhPsJVi1a1ht
8foKUQzCoOWubcWzaedYIr6M7UZP8nYQLkl2ezb+r/i9XJp5uNNQHN39Q/EMwD3KSPD6VcpzoWei
JY1t14RqI+bd8XMUoAWD7iy42sSYZZG+VIVJ4R22SieWbOjQuMc/tyxBRV2AfNWJ0R6dmUzJGEGW
AvWT/JHN6GmgJUA3eTni+6fUuxrs2HplpnnYd9EtVs0XMWnZTCFF9eJht1RmRW5wkIKPrDjG9ZVG
OJoi1IPHD3+e0E8Qb31PGExaucwRz4D5iuT72qcfy7mXxbEYsMk+jh5E3K1Qg6BIR2Zbx1mGpidt
/XEuXCyLJFAPP2lb4Agx8E6lzH+Mo2H0hmoV5ixOERRp7GxAc10g5iCqPJeffHWLp6fk6uNmLpeG
6gr2Uj+9XRGZJtaRcPVxyi0PFOcXn0rMjRdc5Ib3hYAc5Y0Ca9762dSECwlh7WNV3Q+J8tAQO2ik
3ZDjaqnB+s5qKqcbDvXN/zr0Nc3ypJ1a9vsRBRmZyRUD0VOBDaE2HLfUMnAf229xLJa+JFIBRor9
mirRoyBEdp6Um23yvVuaA6iVTtr5xY7ovs3/PLZ4rGfG5LykXswTvGgDrj4L3ftj0qx4z4Di0HzZ
HVQXBxCWxjYNHWzhUK12XCPPts+zsLB1gnXFiPDhBjDB7yrbDwSM/zOrPcV3jQk07zZnurS40eLj
TjBSbgNweWRT1sN6Ph9k/HBqdEWTLBqDbp74qftQHG9Gi7WrdrD975pO6Ij6e3haNS++VO/G/8Cd
0YQ7x5wh3bWml3eutj7CBiJ3UFakZgDgaet4WvQBTild0ftIt+HgVEMI3A1aQRnisDRnM/QFr9fX
iRUQ7+EdDPuV2Jj/8MRMyXT2gqJW5UmFaafw9hmEG9MIWRrMIKBMaRpFbXtpm+719JokyFiaNpHH
n5t0avMxVKLmTldlQ3z900FBC05JIImMfO7aINXNHEEmScsb+iFtgbDJXsTYtgOTsHxbgXzBk5C+
Y+YtoanO0/LNa9jaHQj0eOUMa69wzgHRmjwvGZ1gOPeT2+VFHp+8Eqy3C9jytbSNJ3qKH33cwXKE
ZijnQm3FvT8T0uF8q7xJEFBy4l28Kobh3hKkc4Pj0c+k1YGdimNoYnOneiKwn/FhvFnvsV3qQqlx
rKeZr0qrepmVItVwr916HDkJvA1f1fpcSe2lSlGeYDJobIjaHZc4p6dAnI84O9TlM4X7pYW4Wx88
4vbHljFF9RSySIDUr3bTz58OCg+WnPd1JvwCMTPIxVuK5uO7qVBKKy3CUjhXHGW/2uW9W6Fqks6V
AkRWf4SgVhU/m4i04UOocf059MH28lS79IQEt0pFTleyE1QfU/m+GSnCpA05VBgRuwkP+J1g5por
qs/1oHjNxfkfY7s78W3HQCrZxtp4uzD6APSgjT/pcNCaakAupYdBytMXaaJmlRam9E/9ZeQwklbf
OyTVtlxhXp2DN4b3E33YaRhwa6K6omKPEZwa2/bpHiMR8tzOb38w+PP/EPclPMGlGG/mKNzXQDa0
Sx0/w0P4T8n8vIZVmxRwjbDHPZP5dTFJHfIeFPIaWXbPPPcRYFrSpISC7/CdQogeZXPBV5Vqr5L/
U6jhNn9TDIweUMXLsTpzAr6cztLei6HxsQr2liS/om3ZOIIx2IVF1Z5x/eYyfcBPD4IJ0QUAPPdO
YuY6ILLfqiZDN/zV21JzbhF90g+UlaVFQkCKE73nz8RGisHBF+oiQy7NFZjDyH81BkCoPFEa1meu
lI48jhoNM4H2j85v93VWKdPwJbsyfVKeRO+6IcGe/PqMC0eGl1od2DZ96RdzPnKAckk34fc31GYb
qovepkB/vudW2LeUPbdM+MWE/SjbpwmergLi61dGdeqODtaaANTV5tT0DjIgwxPoQ9ntVU0LWjvW
wSKp3r3in+BTPgNg5BgcOvQkrsJbFE7kK1PgNeJ1BWvAkWGlqyTNGAQQA+Jvm6gXp0cbxSm3jxLG
E8PmVhjdgGAcelDfpeEu1MM09oGWLrl6Yojdg+IujYXJKWJqroiphY47TcG3vV/+xOzb/AWrHZJq
phcKsTDjThjG6NHLnrMctA7waDNGOSidC749xNob7ERYLLbeeiJXV8iKCaLTICgoA7CfFqmjDDCi
njlDEN/hYDUWWJM9RZNqWKv7BuLyndZNCEXr3YlO1y3RU685dgS7oYLutrdQ17KXOHWs0RGG2I7Q
S5NLqnujm5Zxswko/Gj+VQppLzraMTtZpOSCxMrerkWWnvG12ttBQVCcPDBSmVnpNBmcToux5Wbp
aA3gRypnE+Rw1iQbE2asxpkSsJyVOmVyyRoxSvkhnICAoUYz3PsrvDanst1YJ//o8yiKKUEMz3Pe
t5aRWjYJ4Pt7MFEdz23OtcXejTNUgY8mbpTQO7ZiNDqirx0bMaJF9eetfui3hLGFhlzamT3U+rL7
nxM+Mmjj7s3H+tn41yAGLwbW8sCDoGbnW581YglLi7GqW9PNqfHttL1tfbqub3R4Lc/oAscrzG2N
VsZHeegEUda+8+ehfqseV8GlMSu199U/wd0noZ++E0Qv+T6O3tNOY7GO6H9Vw8XrqXfthosn4QSQ
6dtmZCzRi5wzbpQi5qajq9pQxFS5VHcwQtvpBmy1AYvhvy6gZ+093n8HjUbJ25R6dN5G4+BDidKg
Uxn6cbhg+MevpeuESMVwchvW2A1WYYodflqoFZlRUu822sS2YIUCvi//5eWvp7Gdyl7rxldrsEpS
FiK7i1LJNJLEldrk0fsbsyj/y7jRM609Do/TbgJ7bpAayqjPttuyG3JC5+z/tteeV8PT4U9t4t8t
xVKCfXh6ZLsz1ZqFM26t0yIW+kkfpJ1xPKKicBrggh0oCwz86ha7FT1+ugOAqADdFBnnl7BFBbMo
krdDW7tnNHzMDJXxNkSZwD86zwf+1gneTzK3zfh6sRUOZvxq5Zaiu3MXL3JFhT6mNQTqUVlAVpsu
kSxvnvnQJ+6Qf84nh9ogflCs8ySgN1EdGGU9byIB+xaTkkxx34wzjzfbDayO1k/0CpJ1PdkJmNic
oTVlHFv41+fP+gTee9ZfE0IUNSP75vWA1KO3lkCuRom68y8ia14XRZhnvneA6V/ZFRA33ZLMKXKI
nqze1wSwv5wQNUasYo/yd0sO1lD7sv5Dg4zE7iuNyrWWxr98+WD1wklqAc+e1iEXm0ySZoP7yOR2
WQboyVe95MCruHumz6hs0ZkhXissqJLH+0upeZqibZZI/DySC3rimaZFWa8dGvFtinCYhbBl+S+h
N+QreMs8Q8/xBAMA/KJBW3Iko1ke5uT468XDQMHj3WLnh0OOUvW0ib0OdQIPyVO+NbdDWra3tWgy
gaUWaEtHP8/YXn5lhEYFeRjnwBlBtkOFPRD1DPVK6nvK6o6JcSl7aUowVUlOWQiYCG9AXb/FTCFc
+dbClLMKImzL8Ar7H4w5vbPz/aiQl6raiNnClMi9DxoONhVfWm/BzTQdR1OMlrLRlET3H5qFqD4f
lo1BP+WYRcgT1mZrMi85TFcf4pZEzibDmg+wAiA1kzcREJC4XJaarWa0wAK1PeljlzFdwnWNuyJg
FZu5uE25a1Y2i5UVrKDUaap5YBECPZtewBdblBL/Ijv4MBUB6rCvCf694w+mBXvAn2FGMlOcDN+7
pNi5dJoQxwuo+MsUvnEzbfW/JakA0YoIVeu4+n3sgUTyG3QwQGTq4g86QUtGRJKZDc7YA++QrI4N
LsYcudeEezpcxr3ueYvqNa0vAtslQ6U7JZhGX9+/UifJ52UjV3PoSa3DHg65xX8LnM1V+GSFhZXC
A9EzpCXOjoYkluVXTrpTUYPLnZ1+YbQ8SHzpQzUwo9CCzI6LtIB+HRGj7LnlWgw2pnwpbGjT5Gh5
rZAp6lx4xqtMmVNftZM0FJhezZ9uPpVnibjRilk7czgL0m8jYnGkhvMxnk87UwNFPrm5McTWTrZ4
eLRxlLu1QCRAjXx3Bdb65gVXF7bSQYLELQiJuchc2mAf8d07fgpwjGTHPmpqXap5paLX6wW/0kQn
IQ1MCuRidspYvEFsgyAfIoupw84q5YfmG5Ri26nc9Bp/SVOAR2L4tzHQxwPMIbXbkLLEjRGuI6n4
uVHY7Iw4N4YdGRnm0Hs2+ng5auLOsOTClxbCf37Sxriyj0e4geluEqI8rzsekzTLgq5ydCeJ6PrI
s1/+33dvTBtipRfrKQTYLJG1uZNX0yuS3382qki6hUxCinZnkmsugkil+x7kd2QJxVfafPma/G0T
SQsUazYNs0jk1N0S8M/KNGS/w/9Gay6UlCr29KPYQ1jl0snWguM1XYtfTQn8jl41CuMAwL5kbc0a
paJ7OECXueA8vtnQDXTJrLnVHm8cPCFl4C8o4PriroqHkkmBxg7Vf+FwXj2Au6FbW+Cag6x07Xu9
ibS9aPqMzsErFR0ob8I/wZ7ArOh6K8gxsyn66/vlPSZS9UxQ6QPbGMD61GTa6CC6tbb4egsQ8zus
7MuBuCKJjKJ59Q+iFUPvXhZysZOYDSYPStHfFlsIkQ4pWuEu35vqCWebVQ7NkWfR5QccdcezXEBR
J3USyNRv76lbdLG4lQVuaV60+/3dtj+fyO/CX9XEcZGfsDFps1USmVW9xOnc/63Rcu+m6f9/dFi1
EOjumCrSeWPwWruZoth/SfKlRaMbCUg9WUTRM6vj2p9xioA5mu8Mnd/YKKtorwWcx/OkcSQVFcye
bXmC7v3gZFww9pQz7gPBc5B/cr0XOIWOqWHipkJov/0SHU/ZBbg7t/51bkoi/xs2JWD3nOnfXMlA
NMD02vIuNKaE8aIGAQnYY9gMTxWD0G9qJvLe5xjZCn8elAllngW0wqtSKplKrijABHR1E+ZfYcDE
YBTpxlGTSqLGrIM+VhqQExNfzmghocUGLxZiBy3FFoMIuBk9bbig5xKw4DVZzgne4pTXvrMzlD8Z
G6Qo7ja5O4JUbQeFO7kWf1K1VfQq8D/bou4BOF4qUDl0LqmW9Vc/y3PDprZrzosPU4V6wirgl+Kk
yrVKgTbaZj5kJBgqOEBYjEu57dPSFRHPl22W5XjYrKkAASET0w437pFiXVqGbG+QaQaKIIzbTsbc
R+Fc7UdruC1FLTGKN9V+eN4VO0vBblB9zm4ZbQGPIEU/Y48B/0dxr0Osew+qI4XdxCbSCYMgaen/
0woJ2wSd3BC8SJxtqrAeu/m66qm6dcn/GNZ02qgJeUPlaFkKNLIL89gj6pHAgpzWopBTnfi3iYxK
p3yeV4QWq7yfNsCim550LMYwb7iES+4Er9+SVXCUrgt8G5iLn6lrKrZxvDtuaQDP48dU4gTDtsga
+kpGDpdyEkQLwtBVzVe9ZByRWHkfHWrsrBpL52bCig4Dc4KATddygIZCZYZIcui/Azc76PFgSBmP
iTd/g1g1d50uLJf+hRcOD8CQxWBT43BzEFv9VwLRr14k79LNtArR+R5QflysRnBE7PvArc7t1LIo
OTImLsEcTymxl9v4PEXf0MksVg+T6D7FFbBTigjMdFnZ3EJE9+/RojzzBuc8/VjIH94Sgyxo2nDq
f/XCgE5KZZwn9v1Vprr5skR3k69KlJyxvD+lLE8ehX0HW1+CVn3g/GQO8m3dRfVORY14ryWPAKOj
lxDNXci2M+PrKkL9fiYJ4ufLKEYKK/lhx1YaLcfXJQ0nucDbw7tKv3/lL6aEns0dFFwPHv54Xrzv
BTMLR9H4RUFNI3vfvBYiP46ebAclGWM0ikAdckDRqn39rjhw4hSmwpL582oUxasNnnAXtN4rGWK8
SiNYr+QP+uCaie9ywI4mIWJGsXVQtqGSAAvZTqTApkgT8oiqHXZELsMAkXVv867COJOKYBkzwY6D
adSTF2ffMpkcFJoB6DeBKNUK/1cZ4VQleWuYrtrfuSHC4jyh+VAtPLuHiFSZkILFjK75Wy4uOYZo
9xx9q4Ohk1KbUg/hTq34gCf0yZM5DfEmZqzrVcIpsY647ecatE/VgoDAo+OQ+EVF2MfzfE/X2Cwn
cJ0wAwOdcN4muTyOrN4Jpnycuj1lSNKR4BXjDbZ7v6uVjUKZK+X8sV6WzbPKwiO5DwLEf63mL+eK
yeSZz5+bATQLpBBtBhkeR2nDDLt7QwGWMCwwbsikjsPBF4uv3nB8Un5HLPC5GHWmSCQ3LLwdyogI
dyt0zXNbB2hOG42Rnh1NhyAh2kKEMx68jnO1LqqAlY/+Eac1XUJaK/v3ybghHXZ2QH/jYmu++h3c
16j8nAcBSGkCAxw2BeZpj+PWFQwZmyclcnH8/JnuNrZH4BAs9zDxvCRWc7iY0NrpBm3tn98FeMzs
VsHmF5WUKbNEzf2re6M35MfKj6DO1mXuI0R0O95cRYI7VUk2lCtVd/TB7nwSXyFPGi7C3VRfmxk3
y2RtSfSZwT6yD/VhX71nJgSlpd1+kOCuYoJCoYezCYM/RKQd3Jf69fC5+Y0b+jRSeExrWvma/PTh
MGdW8fXNhTz17CRB3dCbB2BYLnhUMWz1ZjvnI6SIOIdDzvc31hl4wSlrHCngcfCk+ammbSWqraiT
rzoG6If/rinwGxgi/3C30e/Bjvb9D3tbnVCmhQrLIFsDpviQGNHF8jwTWmsT5uqIEj1V+SvVOhMs
FwIO11Z56lgde6VXuNRsPrq3Rl8/EMLl1okU71W28zMn/LfzZ9Cx+nWqglRy0llzrTEQQKpcNRUY
ZYiJHlVX4VoQ0GM6ddYPAAT6gqfA11OQwtBdfQQAIveSUy1WqDcYzI9ZZURX22u7E+wFQJ3AJtbI
EiQItH2Cg1kOO4cMI9NVtHwqfOz+cLVljyCALEraHq/YU4s66+k61osZaL5QxPnm+4JYJQJ7cMuI
bc4WfOgpacRchLlyFm5GfjqSRjtdWjdjdeuyjQv9WpX64ZBGFnvBKE1iezgnyA1sDVyZhR/kceYF
zMw4xevODZ+LZy5xg2+Xya+iLnCAsh7SqD0rbRSc9Y/49OeQWTZMrb+5ZFd9KI6btJu7E9v3+rzy
vlKxnyOZa7rsTcq+JcUSYD7rGaVUihzYdXAZezrBKDvE7UsI29XEuDSIgDMtlyr/UHK/1HLdj4ip
7X5T8lsqlONUSGzoIUGDU0XUZRE06QxsEVGQ00I7qbKykeyqQwz/9ZnfQwAL+233xGqzTKkNoIKY
SdqKGhsp062L20GPK1NWw62YUUjKA6TJKl3sPm+ZjEJ/TiDDvnu5hO0gEq6inwcAr661DGmx1Bv+
DB89eQc4wV/R8Zp2Q3+GPUGMaxZ+WrFAVFaGF16fGPIkcMqdYHqbjBAQgsF8mTEB5GCJyayxqpgZ
TlsmUlp5exxLSaz9363yZmoKWAHjMoLLI2X154LVXmRu8UPaZEkDyKwdkUgekq7Y8HOEdhnDfNK1
ydcK6IQQNUfGpWOUZ3Fqhs1GmXjNn/vtBoG4x6Eyk/jwL8f9wKW0H22GUh56Dc3+E6Qkd6FWLLaZ
XzXgH2Omaw7gljAEwUVT4zWUubVhs5AcOtoZlsauxxgiuLmzOr8++jk0Aec3QvZc0Uc4Uv0f2ML5
1spMgF60t3VxwT5tIAnb0EWNAvM2/+c6IAAJ7nEtijLFyQvothiKlKbSVTBCYYvSfQJEEpWQYMv4
yoVPvKEmLddOh2bZoE0lDD5u8Y/tzV+oSryfH6rgecvEUsHJWsaNKpbnts16g84atwjm2vlEqAVG
R6lXUIi9swQDWUDxQpQJlyY+Qoc/Qs3TghlOSyqkdpUm+e1EzaRrXdFFktqCPNOn5RuZJfsj+BHl
R3siU9AvpgfKJfXYQEAPSk+hD20XWsev7W1RY0myPqN0DrkBMtLGVs6Wv1rzLYeLdSmwBkuVELLo
H4ZaQazzdVkjlMnlBrYtvEovLUbVh6WQZZvlZegDiwjb0bSeRxDa0rlpyCUr67KjJR6kTITrbDRx
4FFMyuFuj+GhKZIb2IstKrBgbPiL4XzCoft5Lkz+/UhAlMqlQER70agTLgM07/j7eG61hz/kCC3B
KxAsVlizBFqSFh0C/FyasfBsseAAVcwg6gk+NwTNTbaNUCaQdiILCcLb52LSsUeI6VeiXoyEQ6q+
JZk+uZeubA+v2iq4SMO4mr9yjFQ1qTkzCLS/rDLmRH/F1yuNmfoZd5aNcJ4jwlxO3E6Kyyx91nwM
q607mSlrFMnkVFJwAqu4eez/LQi0OlVgwqE782QLKD4IlTN6BoHj+ytRQlzWBXWiTUzocBJsPgo4
4mfniVfbTB5v85tLx5epymuFydH1qiOnKI5e9C5gyYThiatQUqT+R4rmFJcxbzYQUcYTWq97m4n+
cnV7P5HY2uOCp8Cf3AFRu1Epobfxk96Bj93lBt1Tq5uf1dYfuGEHBImMofl9Wy68dEaW8lA/PGzS
cD98x0p6xYBrOqkxc/x1iNqaY+ac8J0rpmKHkO4nAwxWMGPD+sScwXgLqZFsseFOQbDqB49xQdVQ
act1lqZhb8sgzGG7dystzd7JEqTxoCiGuRh50fSu9IuTOBLUnAcsR9uc9mlzt5u6SnUpdKOmaSUn
UQE9nL4PzonsVQYUkfs0p8ptu7hfSqQM4XkotNo7dbUlQY0airIJxY2CQtfzKbhmpqT3viBvVjyK
hSDu2vCJziaWztM8WZfwaqK/Y3tXI86cQU2tOQH+WJQRvlcybFCLpKUNTVmXxJ0wf2ZG17k5rStt
AuUldzE4K+Ln3de47c+4fU6PuoXYGJ5VIAyQNcNr29C6X4DW+s5X+olUqvK2Pm+IR5DN13672OSp
ATrkGeFbwgEpq/ZRRw61brN1BHKgLQa+Hrnp3dAAoRCCHNbCzBgoklxOtSm/kbDyYVqCmFQdnuwe
YGz9cxkyHYTdhXAmLXB9JSRZnA5n4GKxD20kY5Xrl5KrFCSwqR3fvjdGpoY4zDYy3c0zjNG6a0zK
EvTrV8dJu7F8qCxyZoATSrSt4N60fKJ3zNzPfEsX5b4JOSdt2dYyGaLtSHFRBJgwoIATcbyjTBhW
rgK2IoEQ6WE+AFtneVvPPMOcyXZ1M+v3Wvk+CLfsxtb6KJEk+ovpWrgpUwDqcw/VxaGI37xlgqtC
v5b346YAKoiXzU65mpzPXSPvTuMmQCgHQg2nP6HMfLXrs51SblivTv62GUOxL5327eJrlVFUeb3P
zrINSvGGZJ6gxa2CEAa0uWqgACpP8kj9XG3s0lvdm0rgbAcaRanOqhyTgdOdjYxKW3AAMFH8/fLw
5R5/7zOHzKbGYZBTgQiH0QstqFimJ4X42P1IFHa+74Jo/+MRkweWD110ZQEkFt8kTxVYuSTYkqE9
2a7Eu/FssRnqtD1lp5VUDUKwTKa9+Jd1WACGHrFzvnbDJbi/UzTnzfJ1GNUZUR1NYwK+0C9q+wbR
d2qfAvHfpDOYqlc+T20BJp4KyF3qrSG+HvdDmPHmqHZ/iQrXkHqPlIij5C9wK9BS9WSwtOg0Wom0
W85bEisT6fcvfYqj4Agj06dQabEAPb+sB8t6zrV882+UD5csieJfVJx2SuXIh6cKh2+K5+CS9pB0
p+kUjFWTqubfL9aKap0oXnqBeWlWzr6tDHnnPDz6ai2nn9MKhfTjfiIPGJiwl3blpXb2PbI3VNqq
F4sdaFH1y2Aw9mXejz7rfZ2z8/ZfChO2trIY2vq1f9/R55mfPiaMedGyLFpm2io7amqALQb8tAti
gQw6/jVzDyhAybnPtkfOLXlLBT2/Eo1lJWvKqWwtLF2WW6fSh8ZFajJk6j3R2IBcy3fw/KdmkD/s
FNXMsiA9VVfpoEDE4xiBmi1/ZUCJc6Gh4rujmshv2f+D1JsdumvdA2hUt5i5+hQzw72H7xaWkzn7
OKyUHWK6//lNb3BwFPtv9eW2887D8szzllGspYl5KQ/dUTIByuKcHVutfOz5UYDvG6TiIw5eIabK
jTqthsOrtR6lhYjsWc+2dyNklWKGfdV0j128kBls7v+79cx6sdK3U802Vau+yG72DW6W0dQO+LIV
coDXslDOVX6UvY2t8SXj2Xysrc5nJdjNBW0k06WI8ouUzfVjufJwF3sFgGA3iHa6OVixVRjv69Nk
S2n76vg5g8ktA7EqxjR7D6CYznHTKwgheLnaZApKdThwiZ+2qPy+qZPNsqUQueU/QJi0ldoHeNGN
bVRGfrm5oKqaf8Af/Gl+cQsMJKzIu1iuA1rO2jwBbNhAJU8yS6g6wwUlXoUdDWUyoO7aHpxdHE0K
6+o+XKVKiDRRkn+5Q6SJYvQkHIv4ahSPSl4hBcfRbKP8G2sOleB7S9LlE4wPjaoM8ksJpFabHO2X
Kmy3Qhrr7BcuGmf19eln/H3av21KeZkq/8yofVN5n2L1Yd/aAzlhgLCZjOtyw10EKlnXKyEcSwp/
w1/b4aMsRaV4f+2eH1DcIlgydJALadw4XlwXb7Yh5Xb9eO5r1Ttu5K0zthiX6/csXVgPJQ/pkhlh
yl+yV+LLG3mIeb7Opn0VA4VzIEccrdaVpOhEIr5gs7aLlCamnc9YAFhiWcIr0Me/zr7Dy2DqFo+s
8zProhLjhFMlWOH0fiFvOdFQ1dNg6IekA3jdL4k/TmBuo2dhZDGWzefj6IZKNbjeTMC/WDLj1boV
Dwm0/JqpekACoZ0Gp58LGAXUJTL4Zd0wy3jRRgvGGeE61kSA3ytNus7xSquTlNgPkuCgvCcK9glc
0BxGXub6yuCWnY/LREswHbGJ6bW9vfCqBCofhdvddJ+Zu6DP/icyuvCaXAqyaLSG0qHTiAVa003c
jqeurBrOo9iaTkLXz965g3wlQiMkm5jMIW5Pbsx3nbzSLRpH3KkTZpy4jTfQPQ8gGTWgF2QLCtAO
9BC8MMraBOZps1UsKiZWT1iiVwbjTBS28yDhBUAmu3VzAv/IMf+/tHVAos78pPbVo3Vdvou7OW87
lS0JrzSgfwnjXiXYwuPuu2iyukFEMmzAAjkEVqWXWk9+vBu8ADUIzVe5sa5153txtnjJc/WlM4K5
lX/NZgUyY+1mo6IvwQ50OVR066E8oEY+atPKbzFOC0kMW3+Ce1EsLTb0yh1C72wE/adk5lzvVJPZ
QXKlimHzXzqGLDiMpqvhBAjLZ+5rjh+pVFumQ5YhAvPFlCBEsFIzMbiF88KGf/3fUMs7sI+jTb2m
a3BCYSyisJqlTucwpU+oavFjRos+te/DNEJwnMbN0nkiFkNi131O5ZuOhoq4qJNnLC/qRfmN5XXy
cAQui/l2aAow+w3X5A+x7JqzUboKQ/a8ZRAgGTAZDm3DD31KKHQfqaG2+x3MBGPsOg/wkjzY1nFd
0+H82FgZ8y97+zNFf4glqq02cqrJJhp8sRSD3JAQEOnnN15I59gSo/9MIpqYFAzOrSjEHFDrNk47
D8diO2HcKGP+4K7YJbMxKLzwCQ5jW57egPVFLGMnVcsbl+uZq6xJvzGV6xkvhgDs3JaAA+QWtHxM
cLMzuPhVTo2dAhZlu41ygNSiQ9UYLOwJ76mjZdhk/SwonXHqmMYivA7kqYDcE6F7KGEjBvGl3syn
XL20jrCCfLdQo8RMTKeG1Gorha6WJdmJBMpi/ebJgZemizaR6QYF/jE72Tx4SQwLaFSj13pSNzrT
elJ/4MaYFDELfUDdFpkrZ20vFjVPohPBcJYtVatRluSHQDHb1rk02df0bEVzyv6Ol0Gw0opw5rkC
bsZiCN3oUU0sbc+gFqh0g3vJVuSgDL/JcJZbnfrDChy/+jnVOg3yah0a3C6VdSobOWfcRFYLrW/V
gC9zncfZ3fb0rtDkOOj36+56bPwUy19ODnEpnjUr/nFbGF/qLFzdu1bVLd38eWy4Y+30ENRX0b8A
Sb/wgYMjnYwNpV+vxLIw/V/SqL+n1EvZ/ufgRu/mOFirtMYjG2PkT+Bq/YvKkf9y17qt6djK6uK3
IoTO0A5+sjAiMA59TpWMuHGVkHKW5gigmiiejNLg77DUQjmEiXYidIOoADaUlMYkZe6t1ANZu9MD
D/HQRzYXWQ36i6ol/R0ewGm2aAP7L7mjh3v1sYrEtJa8QfOKVnNh5sUXGSkfkigTXu/cGAmzZVWU
b474RXmy6+s27+cwE9pWbuQFAXgf+qEa4f2hVCJyqCwrh2TB03IgFYXJ6fmsmIfoxoTMyftOyYDi
aU4n2ICf5worllkyjFZozFQ0x3DvHFVissvTJ1EaE+fQ0VianCEEhLDR9PMCFXFEUALGb7B8w3cp
NTbXYnAkKIprYxpaPlwrNn2KjqPps5Q3YJ73yaDnW0IPk0P+ajz221+Fr/qCnLG8jRCFPSqMlY3n
C91giOtfdW/ogefnjjTkdQLXkBGtUbjU2sb8WruLDpBtVYmnQXlI7PkVWqWGbeEIjRJwAR+LbOR9
F4oD740QWBcbrFAIqLwDKb1WHzYXnvOAnh/wj4BfB1wfXRttP0zSd3uCFHKGeEhhv4AQf/pesP4n
g/moiD/dC/J91q3IjJJQqG51LwcJIxLPIzmzyTNEjyYaDNr0c6KpKvYdFLKQY6oCbylV/8KGPnIm
UvrRFnq47C/d4CjmB7ENyu3K577LH0VwS6YT4vpe9piRZMfXtrP7sFOqUotjtyRvkjxscEJ/d00I
GmZ+kdoqLcMV/vTEsOfi6bwwo5L8ZSmjwFp54pQBea6bv8FwyOQCCasAZcT4P4HooL/sXfzNMDib
uRXWwGOiOK7XpBLyymjveC+I33Ogr609oQNTDNNFKPsVfwFH6yKGukryJRCoGgCiJrvxoR4u0RwB
rlWcPDZXUsuvwSPOrFCcPXrdX3Ws4Ga1r//5skFub5dyjscnQAZNHZEMJeQ/DnX2gqA/Xa1FhMQX
GIpFkAhOZ+idY+v1Q5t3vwbrG28IgXRSYQIMG8EnkykGsrwJPCmkHX2muDOiRXwF3eol9Ys2u1zT
aUO4/R6e4otvQ0bHO92wWDmmdkd90KG822MLFZVUkCIqKIlQJqj7NFLBs0Su/zDMHjFCDX/LaMJX
IYAKTqmfEFneHvTvn4i1LUkZkLHbqNO0ZzzjWhjEtsCTPgZ9OvwKTw50JxWpFlIF+y3Y+qUseEgu
vPQsNmHuh7krVxzv6oV3v6j9+4ZT50luI77aqTw2u6PpvXkg7l8MlLMbR4eTk1twGXIpUF5BSrG5
sr9BSORQwmlGvroiJUJO3z0yIBecpYDdmnrePhKdcpl3yKYDYVdCGFhaCRHBBEWdQXMYw5TwzgW4
D/LYONWPSZBx57xPRG/1+5xI4FnoktiBcGNXI1hgNmkST3t2iA7sPzp4L0ttJZQ7OYUXm8492iIl
PAaJyJNzGi1Rt7QpHk6JI1sTJW6g/x96l+Q6xd2hYtRZmljpVrYdVtknDnTIJWBqVEXte/3MBeun
udRZ5Ku3zN7jin+zqFPR0ps3JG2GpxJlJ0SPVgu7hm0bmGYM9TPnhqj+2RjiEOQiMhvJRIZFfKbS
Q0TgZS9ZmZ4gCxkiFG5X8u5w5nxn0RO73EgELITULjonii+wkkKrOm20l0sR3zfGKMrv2IoiG/Bc
FG4a7pq672xAka+iqfkH2QU/sGjpvEJJxCdZYW7aA1GCsHQjWRX9K60wjv1ZulHauwI/YvrnIRD9
r2MpaasNjDSa6gUHV3VGciTGuEzx77oZzIcqfSq4evUEDO5qMkKJRGyrbniTJUAV8UmDLnvZEPxN
Cvri+4I6sTdxKnEh6RJ+StCc65TO886NDhIVUNVd8NwTL78C6FIFfFueFQMc8oZfAZSDUNjrdRxR
H4OnaaScA/DkRcCUkHm3Qbcb+nJmNDu5mb/9Uxsw2f6RB+gB3FFaK/Hv4q7ucyvZtRTFJPaLxMX5
jhTZMIRtOm+45EYDbrg3qrdCy/yt3XSsJyyXRqsJVmFtSiRAM+QbC3HWFQVVkKkZjFqH0yAjjoN/
ToJbwrz1Xw0GLjdn+iSNlbCyMzIrCvqz61uqbY0d4Vo84+R7kczJjtX29tzHJY+watBjLvYCO4/Y
3R/u8l1jkHxHS1rXb2rKsSYGTIbJ4HwUcQYJmUtoXOmrBeuLDuizeRg/wGpiGTIrbFTniSVFzw8h
XW0atn6cSzNlHZD4Cwj6dI6BzxCFbMxCLsd53cV1EHXi731o/a8Aqf91cNGwdE/Oiu1rxUtzVBA9
B4geg1xqkufk/9exxGdiEWCjJdhJk1WM9ozV9t9lHJIWDvHVnK75Z8FNwAdAMSvvCkHzVOdwsRuy
iAiY0j/tLHb30XaaN+hcJuacoxcAQpVf1u+S5Cn8ET7K8Fi+AWVEGkr0M1/HpSgu0TKtg4c4tDgd
CifdResceCnQ/avq27gT9QcKtz1qxjC0AVn8sE9B9qKXCJUCpZfORkDv6aq1LEatdzbZJyQkmQNr
xZUb3FjHOOo6TgZkde6Lo4M19UtyUMA4z85gavmq9b5BywRumEqYt9zWHt1ggHGGhMKuIhpE+bsK
iSYIL2xX1jkzJm80Y2TA9Pg9jQm9D/Blfl1Gx93cqxGBFwZHTaG4B/khMgdORgXaZD1R8xkbKfVt
uZQIDwgiaNorcNEycZtlxw3/HMxNvN0H4/38ynRZB2ktL++d6SBT+AZp0THlIdddsR6x9OqzTQ73
6fOVHv3GGpwqtCgfW8p4FI5uDWkuNF9QcmhxEsOwZQpQzttWAdjebhYmtiBy5WvZ+0bW0frRf/QQ
HqbYMvKG4OZti6s0Ec/iaydI0NMZxsXctH4NJWcw3KLPmS/YD7SpYk1D5QsgP47gPgV7VzziY176
QONKaVjgp0COdgHQlIM0K7OC4NDFqwGkYlzm0uOzYHzI8M3WvF2yfEqfFbhe+l21ukWDnaA5/zm7
8B/S44ABeBQCq+DF5bw6xCCAQPdg2R6c77JZoPNunaGE6XRRdeLGblUWZ2MhL/m4L6Vo0HZEFfbJ
ZgDljJokXu6TM3cod9PmLkXdLOGvN8Z8li7XTFhYacJhoDeIvYK1r49IMLc/qiAxFPhDYHz23sPA
oYSBffQZ+Vf+vLG18D9jy8IeOjrwInCGC0arxA+1vYiPIvLHvXWrDCgZYrgoX4Uy6dPoYdfLxr7e
TO1pf7u6nWVQxvm5hggCusupCWx7lSr4SeKpMJi7w4Zp3zQg0ifjXduH2cIMwj2H0/bAayvgwdTK
adZqdyuU+lU4/pddOwcybHzJGneyLPOOcWykmewwG5JItTRo4d/c82zgFHOjr+BbeGxBTRHZLmdD
G0OLnj6eRhOOnRC6KBkNOE4wfxOngoYraUkHd09mGlTsBucYJBOgWCzTjR2/ei72PC0Oxky+E/R6
8IYr2V9y42kNGlJkx9GIZ9oE8pNa5tXlRko5K3Rau4rNNSPp/Ye09CvZc9bobpXPOA+BIOMoYmpF
Tvg/bku6PcEsgbn+9Xpo7NvEhFan5F0p7ahpPc66G939iFsHluSh85Userhg0TGvL2KJE9PjBaX2
SZ7DCB8QVuzyEgyVZTt7p5NMgTdCKKT727HNVaX7h42YpYtphZ8ovQqRjJH9rC0rxdI7/d8hNIUY
B6pVb9xLpFGIIj4G7afnJxBHyeK87GQ8ecbBuKM9EX1GE1KSZdGpQsLTfeUvuLNK1g+baPUgm2EQ
W4jjjqqu5Bo7MMHbkp0jqtwZbDsHD1UQLC0iGnJiS+0VAqRnDbMLy34+BnAb7G5CU7yvr0w34StV
tb/7fjWwk8U+j8vlSPZKiJjULR8cvwY3zY71CY8SJOrsihPTTnPjgZr2GCUq3BoOX6kGp5oXFAX1
uk85N7iyON17olA59Pf2Y1jVA9Tlq/S26twnamIf7ABJ/DkRINbnhwv/CktTJJAGBYskL0TP0RQ1
meTXTd4cgfruXsZ3jkvP8OSu7eYV7sZuSi5WiNtVdLNfdpw7R7pR9vw2HJx+sF6QnEb1RkvVN3KI
htolLhVJXwP7lj04Yu27oiE/ApuRVLXL1OcJ4eEUIA/5JoSPkWs7Fl7BpGX2tHjQPGmlyMUcN+ar
IBLd2WUzN6mobNv1zmuB6wh1DSZM2RbI1SRKMrxYD1tb4wZ15YrZf86vLR4QvIoS8SBhAT2T7S0Z
X0X0gl+aaolVEjWFBp2a8XmwULA5lWZYB9b79NDuDbxehIIm/SMepIAu9UmS2ozDVrsePEtCwSXI
HVORglxZDEw1myymmoRsS0Sn1MKkZKe97qBo9E9br5INqcfk9w77WacItDjptHNaK+Rc++OFgj2B
mVJUOhnc2W2SewNgQs3nyqbkLMKrM0UJ37ahQF5+bxAB0a7MEhOtx4Sv3JcZYYO4rylZIfOMJdAv
PCYE6zZMcg8t1lfw8angg/SuTo5UNXvKd1oLHL9jXLPFTyBVmPqoDfcTf19SLL4Cx1W+lWxonwY/
LrkBB0PMGkPRkY14Lz9ct+MKJx9+FFlFSxkyyxFioBqibCUlI5PBBIeJ8+EEWjJmggreFrw7IY0p
z0qW090r+bYIWlIT64hKTyb6tz94pYSdozfRSQfTFWR2sn9g1MkO0YUFvAAbktLkOPxURBp77nT+
GN8RfjNDxCOpMQ8NEPlrYCWPPXNkfliMII34B/JaNSfODKOlt9HQWFBsqiB3juMo4rO5hJGr1RAJ
M3rGh+LMOcWSv2RMuTFSP3+68pi9dCQMXyPKIky9Tugmok6vxLsyUCva8hCHJwB0vLNFnyLVdFdw
72m6XS+cBEY9BrPcibixTQFth+8TORHoEo95XLtf8m78YBf/M34FNtktgDCm/IDswPVgay0pLX32
G3rr0BzbJdzAB2laxPlvT2rkUWTGeszV825lPG/KxbKRkTMYp1Lh6Ig2UCWpItedUtwvEdc1AFqE
NVnkHhp5RFGouiBgQmlzfk6V8tSyfYKU8TdW9MEvEDITU+vPFM+gOe/RsWheyF0dneyZ/9S/6g/d
5MQyt5QgWAyBcqw4zwsfWK+bhmyNkVTTH8zNFzL2fBlbw23wvZQLtox3eRvLxDelNhfXa7dDoWEy
BBWkQ0VJFjELNhF9sGE1M3xvyw8pmRZy8oOB4ksCDSAli9LJur6e83O851H5ZhiyC4ANb8HdEl28
EmsTSEhAe7oh1U2UyJjlitabDn2OEOON6RugpRE6f4ORhucUxl1bQ2+s3yN49+aljj5yVE2/ISJ/
+o6Oq3RS7WNjh3qVI2db/m9D15a3RaE6S3zD8RYdEeJJKRabcuWRMuFVgl+okx9Y+fkqujciqnyI
wF6s/59WS/u4B/Wkr7lDPRUwXkNCo+5V3TkmTzHaG00qZlucksAOMzfBBFYD58YWP76kzb1gNwEJ
nmyEusTv1Sh4mviIdEAZCQV4N1gAtIuyvGsUuRBM5J+L7yPq3HsZ58UpFCp9j0d/iDy+Wy1AD5mc
vmJcqhcdFaUxYYFjn3hxMYB4z7sSZJ9cuZz8olAXGExl6fKuYmSLhThJgtujjsaGDd7vOV5DCNw3
LnjdXKfOGeQfufsvG2uAlMjbwKp+Xe0zP7W1kc3zAeVipBIG3dkZIC2J86PcKzvK6WRT9sN0Zc+W
nAXHybCYYhQEpMXo89nFPtYdoRsHz8snsp82o73PopfL79Ko6bn4MdnrWQ+tH3soLssuW7wqwW9Y
r/bBHuOtFRNiCJXPVoAVHAzbN2XsCsMro0geErRc3QYflRebUC3mknVGGWNzr4hNrF1MsIkbhWTo
0VbbcVXAb9EeUdjfP8tzYXUH56PTyHvEcLKD2V7KGkMn0z+CnpGxqiNDqyLLDRLSP/0Vslty0XAV
3ppOLnX81BmrLvZDZ+b3ey7oym1mup1goQ1fmw/rBAp4ZWTVmswnIePWPL66qHzW3dJpTkhj3Upi
RuS8RexhWx/C0sjZaGIwzxufCexF8EJ07oVNzLB2K1nWfgYcXXASbjp/d//ZlToREB8yOYJxGIzt
JRq03p77+x/hkgeKJLQ38CevAkzATGg2aTPST4i7BFzZcmJqutgC81JtnNw14hKAXaaemiCc6vn8
SnmHMHr+R9QSoV2nkQoUUgyzpFjTo9ukGXwp8bYUrcdQZfLtmZSoTnf/nq/wrdbrThp20aZpBB4/
p6KgLKJpiwTiaDv9huA0702mUbpwhXAcc8zULWqCrZuZzjHiDVSalGSfJP3OGJl+kD+njUzAxSgv
f9KV4xNgxWpNT2PUP1z0ea+rN+whx5xdhHJdhMuQBPUvgY9JTGfJze+VqSYFISqpP9kMI0WMM8e+
u9fmw4R2w3Eg2OqGm7SDIdwIlN2C1pDBx+5h4IesBpyyD8Y1dK1axopsbxO4vsFk6GNti5sRtIIh
F4Ce61NoafRZy0iW+vV8dDhUysFieKjvnvV8hki6C3MyUA8RODX3sA0Jd/X5unLrT8PpseL4rS80
yvxa2BjJh+ykQMSqos9tM6kyZiaYdlLyavlU/osHqRaY6OohjKonSOUDDCqLgi+d6gId+Wrwc5Vm
yVS8ACu/NQmCjj7RvTUmXygxsmLUQ9qfR7ID6ZJwkei7smIMb+1I80CTkkkJ/+sJul404UI+9VH2
hqdp6+a9S39VrHEgpNxI/FigkMnyDFOj0gwQ1g8+MSNXbVSYD+vCCKfkFdbZKSo5/vtBIxAHwjdU
T6ZanHH6DqpCcBzhcvivUzh1notyIrn/Zevy/E21e0lH7hHJsM6fjO7LBQqeJeFcQgKMH1EqwJZt
YdkBlv/0L685mdyquS8SSJQncLmHVy+ZpBiiyIvoM+RjoORWjrQRjchxiO+HRTA04cBPahu2ag2w
T4r8X210zqAQHdyOQW9AiS0AfPoHGrAyK6E2tDxkuK0g4OXGmX/JepYwEE201XpBmBLiSyPYvkIP
cWuSVxzT78xTxGEgz7h5WHlYMZF4zTXrU/xc/5mUTIwA0VCD+JI6X24GMPIQFtyxgRhB6tMp7fX5
4eprol/5sjnHot+ydTP8/Efh6WVpuzvN6czsI43qNPosaVm/7fgB2V/gQkW4WVePtVeejQIe7gPN
z7uvLY5sdgmcSl+aSd2fLTF3/chnC6pycfZMOnKUnqg80BAEu2cPJlgMOE6TUy0+UjVi2SsgW/DJ
644WFJ+f11u0y1k2ZsJSKW7upXVH8cPcsuL4FKubnbNHpSpsaPRybcwfMTA/09rfSUS8WXNnVgWj
F9uUNE6zD71KTBxreohyto8zJXDEUOrt6jdMCskxNZwXVnki5DRmQPmhVqdqFt8h8MNbMn5nUrJ2
n4QKCPe2yYrNtgWSor6y9fWHeLYcdItCorocGX4o23sPgIVk7V+fNE7mYbuST2P+J42GqTmgESxA
6o04okyJcD9XmV+aUljltQ12EOyXFwsdpFXWOYPNDFzW40jqmydhBdxwm/baYHDiDTmTZXXrvReK
aTPlzjub1WMtCtWpdnhd/dbJVmSC5hcGt76hptbN63P877vbD/0vQZPUdjZF+Z9TT0Q5t5xgXjCx
nlw/XlvXlWANXYrV8WgkU1UG6/WSfda0S4QrLcQebGyexsVbAnWRzyJ3xTCrC5ua1lqg5+59i+WA
okemXXkcB0EXrRH3mNoQTwqqvF2UwhXR+iRgYRPopEJB1wjCg5Si4q32kyo31XGdbdH6Z7IPuMnu
Kt666xh4ph+dfNekl+L0bOlgW5nFKryQY8oVPLJHchqgLTuRt52rAKD3Apn8IyJfcUM++GoBJfho
YBUhFNpP/Q3HE0/21F+TUFzCIVgpKfaN0KFW4WGw5Gob8ia+WFWVlVVwuUt51J3NQsTUcfTMKLQg
jxgfVYqSLDg+Ls6TDCvMOHJGRy80j+eWMrk5Z+xVqRlphYbLu8T1iWvdpJ1thXShD+KkwJN2XHh9
IuRlTLCdbYBCVXucBFGWE3Ly3Q8grFkqFvNLx+5GwtBBp4qzZ/u5nPNImuiMyhCyAGW46Io4zVas
j3GOiv67pK9JfYuWknQQ9Qk8uiStRXE9Vxif4Lj7YaNTgR0uri0VSex4dN4jYcWoBi71c5HuWIN2
dJslpEotPTZE11TO0ErFkZs+VTBUIkG2cfmmVRQHeuv3Gl6JRbs1juv1+Ol8FRDclGCa2aC2DfSx
nL2OHHRTN4T7nIg0Y0jLPgy3R/q0RNe81/+MygkVyZW1tgd1M2CwrFKqHKGq7rOsdmf7A9OM8Rev
UpPnMdpjGq6cnQSh5DxTig0GPPdLERdUqneihYOjuBAbCGhP1pFXFYHMZ+ggUuUms1YwgrRbUUui
pfvDNoPTNhXa7haqwrBCEKoTKwNHRptDwFtqsc0j4/10lIY1F5Q4XyhlZ5uH2IjmOQ/7JFm8IQ64
4ab9mHl4ei6AV9eBHaETQcr9+t7ITr0qDk/JQEz7YTKdDQSGcNw2449m0N2mjmN5PLe6mikvONlC
oXVPN89jVOsJlREHywSrdAtcmPq4DbbcYtNE1L5/Ak57Gb0zNMjGsBk6yELmDWr06xnJyUDv/aB7
ZE1SKw1kyzoqucYNa5chMujAKkcw1Esar7ly8lwAb/YRjqkoZy1J8BsitwvGKBdK1kSYE3o8/1cz
aaLrqC2sBr1B8Q5cE4C7CpNrTnuG3w0XqjGVY9zbZ7nWoYjr4eHOd2XImQvGqO2XOZRBqxBbwl9i
5kM6gn3lGxhQb36p4NBXerZG5SBFAOeBrQLtsAguzsCIljqPYFn0QbLUL0f6TGBxYMiyXaDf3Fy2
nzjVBm0mY5V3/MABlJ33X4EpCSKVAOD11qB46JCZAMffaGtX8QKVnnaXH5t+iHgeKzWleH4qvXv3
up3DcDBfucC+FoS94Gqbi9okVoUEVfO3EFWCyg0vrnH/U4jokhhRTPXN3gGQ7zR3vpZGOui45sZe
ntEpK+s4Mi9Oi9gHekA31BS6hpEAobAVJ+sc+cRONk0nS0BSPfu8TF0HepIkmHce5HH8MH3iRr4D
Ok5tfpOcm6wOYL6s8v9Ol9O9gZ7qgacmDoLFCTqTNFbC4VQGCM+xAV7vOKEiQm++qD8lqf+pA0Ue
WF2o0BXRD5tzNH3aAbKTPkwPqcSdy5sDKnNhocFhiQF/I50XEAstCTYdPkczsJ3BLQKHc7IxJCJJ
sbu+kOade9dp+manPFAU6BFPdf8Y0M+7SXeQJIWc8gIoPrxxtW+GxVlH60jw7tt6S4Ly7u+NfHw2
FpW0qZayXUqHy+eWGVM9EyadwnsmsLM4WvWGyqFgipjVYiQZrY+QXy1Juh7qEAUR/q2Z/7/taBWO
lLW0Y0mm8qJ5Pq4p3qJEerIYmfXsET2LmhXehL3bQn8Qgh7iYSMcwHycntQzEr6d2nniYOnAxRe+
DTDxW7zemJU/pViM3JBMY4DTMq1SbFGJq+HmdPMoHGy9rzDdUNPjJMHnQzRCYjoAgq3UyNtq7wHH
ddNrWLbeTyVL0qXOxHBELDrR1A0VKA56cjJ+1U3E00X+gXVQUv1aTdF7c3B3jBoKd6tH4BmArgE3
Bc3+xdqHtvkSR3ZSge5Nrr38b2wPhZzpFzO60mMo5pFyjcsmaLLDKMMUazTinHiToxW5Kn/NLict
4wal5PYlrF0WmZG9Colngk/OowGwa63DzlktFRPMFtQIHqHnARmCezqZ561akrskAaKOo4VQHu5w
zaBKhk8QMKYZKdjNGi4lFy3qhp4k/ORVgiRnQ4kggXu/7hSY9omRnk9QRSbe5xxoEKLJDiZX0DT3
Um1R8Y3CytNZmDcBj92OqX77XVAsNkakRFwKyutqOc/T/T0QyRUsNHRZ2IwWKMa6QDE7ID9li/Zt
LasIycDE7uDg0JcKcC+8c71TdCCqk+sElG5K1a5IQrQlqe9O1T9HV6mhR0fLLY3d1mXTmpD/m3fe
hLw5IU4SS8un8wfBTGVZngxtDMW12ydDeRfx84bXLwuduMhfSTIzrIJxrgKAvpoZE/DBnYDCkWFb
OLtpsP8wQ6ttT699dlEoVfxDaU47ur0pgrBXF4RpCZPCGzQEiFqBMJozSeZ1D0YpGZihjQd5nLgx
LTHHg/uSaRTbzt4rGBT9zVIKbfp785pvjkh0ZyyKWcpZ4n86EIG4blgTXD3/HlnH0VkI5KcV6yAL
9/Zd/w3iaCL+5WHLErP5+UNqQpERhEdhnYl7cbncBrhocSnhxJ8oV8utkIymyP4oGFSNa2rY/K0i
pwWwkMcFQdZ7+IqBJDaFEl6nLFCDS4/TdqfyM5oXvl7c/rkNkAZOd6o1E0wXHGyaJmkMvRPB6N9Q
FrTNrtuZNPxh/p53+NFCgWME+gZN7WG1FJBO7V2IUi/iWgO/brPeDuxx9IQVk2vnCtRWdFxwe9KC
LEGFQxpTTP0afXXx3o+hfTav9l3U1mFWMA5PJCnJsXynh+jNgtPXjrQQJiYXcQoqHFIKR4mDDZPM
I0ihnhA+VurzUjwpqxqhGBSnpHaMYUVM0JavDkupwFmgGEbW59UouCM5pvQkluBVYvDD+tAwDQBp
bF9xMuvfAvieL3pHSm9kIJa4iqfbKgCK+3c8Kpi9U7f9hU7wEhxGBGO09iC0JnHaamP76GKNSLsW
mGoPHAQMPjFtHboPDrJmzZQZVRKpzFlPLKqdEiviDpHuKfBKJPqoXeyxvr6Hfdr3M27VTN8TjRnQ
g43rmaBG1DZIUYq8VffER3Aw1p0QdzOWCCx+kZi0bTmtqo/9VVK/sZ95oh4PsrHM+GHEzyB4Sq20
+d/aerJbO3sCQX7GdH6P9OLanIc2NwAq0z3u1QYGkz2q+gypqDd/f0Z9KqrMR6ujR+7npwuTApI0
7ZB/e33CSEGOaXVGtpZdwGY+BbIvm0E+Lfsz2e8DiTMEaGFq73MuGr3jPQmbjssWGRn/CgWB/xcF
iJhU7CoUft3TsB4V26/VoVLSlY52Hy71964vilPXxvWfz0YfVIhLl3prTiR/ixnxPLJ1VaEgu26P
7qM0i5ltDDAekIXDf1OXAtZyHjfvT0eofn75SEN6dZNHlG2oIJBEgPo2rrutQGR2wmd1E6Wk1p/9
K8ZMgiiPVNKaLbyh2B3fw9uEzxpcdhRbxu/a7jUhpZITy6TSRx349YWCMo2Xn6sdUn7Vzv/ALY8A
+fmIRPhEEuXqBRVKZNz05h6OSfawPb8SL7K+Br9lPdaFfoE8dCJkge6uVuJO5hmGXGDSqtccBynx
KUcv9K9E2SWBzmiO7j1oca08Id6ybFuorq2MlM+eil8jEBydWXsgHtyCxN/vOQGn9PmqMvKEMrcg
yAk3HTkuWpizvpXw4aKgwU/xVVIK1HTs2hV1ncmBdogWGjznha2xb6iLRa8ui6+egCPxvtEAEPs7
6zU6Znf8pgMWNhWCcFVWmr0L3PbyyuL2vH1+c/u3EGr+IDiXQKpzBNmvFS01JMxmaqCvblCC5jC1
W0uyTWFSDrfEmuSX9Bz6xGcLlVvnz2yDVFI64hJVSP4cD5KlBzG02J2eM70gXRrEzkQ7+/6lMHrX
mhspQw1JMsOalCCW5+pNxMltOng+WmL7+kyec41p2LeI1avdo+FMX6yP4UWALLnF+/kv4jP3Ctky
nhK6bKdbSuxXsZEdmmz22ywBsQMEnxPlXh6mp/eWZkjFL3qnUNOnOGYEfJupp4R1DLLjhGVGS6zp
p3vgb/tDpBvRRiHavpS6CUF1ERuOtuSf2WhlLDtN66ZktajvxncRlB0BAHmGQ7ZVvFVp2FB3G/D+
lBbCM0Vgmrm3p4jVkZww2iSY5ktZUNhFZzGlquOxfvSvU/KXsXnVUPwGZzgoI1l8vpPP4UeKVP7Z
v7YVbz0D3zt01oFwKGgt+viGVKS0yyjTonstK0SiCxU0nsVavpfhFa6jQXFYY0HV+BAb841nrt4q
g4vKN2/2tGUauXG22o0w3PHkyqi8vxhN6opBzJMNd6cKzw8qUNVXy6ab4ybxe2ekfX2W5H34JtDS
JhnSWJPN/fD1ulz3SciYo/D7Ux2WQaTunSqT1vBVVurVaA9a2eth5VWCBF2VLxxOviowwpZiVyzz
oJk2FYos7lyZB81Tis6IZvolMBq+jaFyIrQzDMa21fVxeqa1BCvK+wBfiZaZXQiD/KwS8+qCoLmY
qU+/bRrg8iDfEUfE9Jv4Wso/QM65n5TruuEXMsqeu94cshtf9ha8wuw55OyTI4dJMEYZSNCNOmYN
/ArxvMu35QQX/iloS0kj5Ck/RXZTQFx0gPpR4uMDeFv+F43XGkdUOGV2Z7dfVH/LOFvRiBzz89ot
cVLoR3phvCpTZNHx+cApkpl14HvuyolQ8EFXGwQvlsUYB7SEuWquFkdP2huu/wLroFiFS8hN4c0x
CAfldd6WTlGokNaCVHsEscZRrBTBQH37fF9SFgkSpQVbsIZ6PwVi5w7JoSnP5JGngc4rlIk1aaZy
xk5b8J2m8GPRn3J5Wzy3xWSAfo3UTKVLK7650coH1cb2HK1iFWblO1T+QuK4wOBIOp6lwCT2p6P5
LNTmjYIqpkU9ZUilycubFDyEzFoTHxqUTWwHGnO5qXY+/cEkxyF5X1onZCOaRP1gmfKlZc7ayR0f
fxgdYc0CwDXca8tKW/G5lkbIs5+Ge1pasy/Oi+pusQAZq16O9HAYXdpwLrp6AbDG7JO1raYDpWbd
cUGzPbgTdEE4pf+0ljMAbQgiTqYyKp2qz5R8ebIN8W8UJafwezWb8FNT5yHe6VTc1fRfrk20vUPr
MIqm1c/7fb2qaz40+L4xujY1i4F2TaoEq6uWs4P3hHji4FcDtA+U0Ulfq2DKlwZCxHDLBUXnfl8M
vS25RMY6tFhwFrUlmiNoG79xKZVxrbqzO9tJtQTzfXa3G/xXMJ5JAGQkG4fQPW5UUlMwbjzhtI0l
TXqmiDkO563IA3kUqOL848bmMrmaVia4kh45dFW/XAJCgdOC+vXuiJ4sSua0OUi3nDrUVH2dT7wX
z/AKjOBtQqIVaS4NhWndsRTaa/KzDFLWSsPIYRucONnQDdMey4vRX/BYAIIxggcSeq/VAuUbfJ8+
732of4bu4mVWMJp+vx6m7J1ixW1Xhf4IJ6nL+ePzrv+3LWSPp90ZTjmtJqIUSOhOEeafJX7keyBh
PIBnlagLWOg9/WxmVu3oYCtiOk5FYrfDZmaFZ5AWDUgucif43w3t47izXXxTjCnngYijjSQ3okB6
OaedybIZcVrny0uzjnWzPe3xmGvHVgzafhExB9KulOmSQiVZ9+A/SplYKb45kn7PvIpIgiqI2tCI
0vKyCqIjBOEOJ00NCaeQYIEal0FbP9CFMYggVHTdy5b64RUTDV+wU20FdjbhPsI8IWfIJ9LZxkNO
V1+//WwAI1AGCBR4W5dnDz8n0Km8+2QEXg1XnwZWfdOGwFn0yERPR0GDPolgqdtQKi9ThPppywLf
Y507woJUv3UqpS7L79wDCscJy1jKlqTp9z5nJAVHHpc/416PhFIMQIdwjxvR/NuEmdJqB7HlDIz0
3DTl6rZihCqj4/IahJgPwKnHey9SEqo22Eqoj2cde3XCjJPVvwnZS11nimA7tM5vxAJfBlHjt+e7
jCTGW+OAs/iqvDU/llWCCchK6ZCjrmbZBSiziPFasTD+qTx3MKG37UHdx7OTr3pUhhCOS/qDw9Um
Yh+owjS52lZkjQ/P8hQWN0vnmj6QPSHt8kQhJOp97MsdJ8HXUKcHcAnwWNG3SZqrMUs1dYQqlaN0
ZVlK5piAnRYHioqGuMdzSG4w+E9AwC1cH0c98ymUG99FbH1jSaDmheU3VKrpwOlO/wwXXbzlaWcB
KWxn0zMNTgPc6tHiak5qR9QspSfsOCQ6F6Cn4evpfHKNNrM4sdJhX2iCl3v5QYWBoOKSkzLVsodq
z6bTumSOh58vrwZJJ+nldu7WQmEo1Utr5RDxRp1YVydT+nnFPn/JAq79edtXB1wPudlIW1s3WwHc
Kbii3y/EXzGGz9nb73Z9UzFg713ah/hEeYU21lg3WaAXJn6KMTJhSXfNvk8yWtAUY0O95AKdB54C
ILnPrDEPMSi1qS2a7Fha6XtUtvZSqpbwIlMoH9DXLSxHImp3KNohA+Cpns5WoEOS4tD4Dsv2mW63
etZ9KUAVZTV9g3naAAAt/z09hHuiwz0J6/oS2XpvnMm+74VB2Zedu5pc2LYn+QPk8ULP87an2Q6O
bgWlbbtC9RaA3j63zuSTqI86LGyxMP/Toc0OyXeaxpFR2FNkz3hENsIPxhUO3bx/Hu3qaDZWYUG/
LobBOvFGNA3ai5B+ysDS3Wnb856MZN2sVHSgNeGZyV94tPslcwPrEEUNR/4MABRjPpnYYWaPK/K6
CgLZwh9hjcxq+Opxr72fbIgmFd+OFhda2oRDFlnE4DFVuLcaOLARCv7uJCvZDPnCgqIXnI9vGlOB
9Y8/uMJWbbDxaPg9NTpwlCunSpk7B6Uimh/IoAAm04KhcKHklP6fhK0sq5bG1YFQIcF96LA3QHuj
+6rzLrilzC35wNRbknqmv5kgVtQmcDC7kdtQNdxzE1QkwR116THtIKO7jVZgA63+tJq7mdtntEnC
sJWiKbC2xzVw8EZaOb7Gygsfd/b7MagF7qPMiVYiiWrB3HRwzCstptaXpIa0rLy6sP++gkcnDrqf
VkQhuEkNSgG/+hwbkP05qwxpEa+zLvto7dG1VEHeEpH/XjS/+EEbsYphr5q/vkmD8wbomRLdi14o
DM58i/ZdEmFT04Yoj2vhIt7siBQKus7YGMSeXVQI3CEMMd2zekCdSSBtmyidsEPAJ79Ufz38QyTm
tZz5xQW0qhngW4Oph9X+0RbJ8NPpSvuDGNO16kT19JKULgKIWHXHNr07o52pYrp5t+wF67L+7D7p
I3h4BdTeMO8x9sGmpnRFymTeBMjkF5A+G8EB36o/+YQd8XawdudBeC/CiHJoczOTDckQA3oKJ+3k
/rN877gvO2JtVz6PNsHr2rDfFtw+TnYzbyRIQs1xt8njUg2bjvAUhw40slKsil711aJ9ybIAwS7C
p4xbYKNazUqGNLES67LDjHhIGV+Z6/czUVC7MOb0BEUO6Pib4DAAq5NcYbspDqe+Q/6Z/SRSaStE
0hnl80VQ/BaOdmWP9jRdHuoGHSjsNAiwNBWNbe+x/C+SfwmaMUiUl/SI4ElqfylIJa0VMdx7rvC3
SzHteZ2spCgQjeo+wtOixXY5uLpyfMGQDqHN3VqjxYgqKEyUwpAJ4CLSAzfe7+8LEcs9b8fEMAsH
E3cPquboK83c7+2XHHesL1c1qRaYzFnypSSZiUqmlMeovsTW++hGLdKjYE7+p4bGxC4SocFmB1Pe
eBRWOtXcbXa0dbwCc3zVL1V1M/zeE3ZrjTO0CX4CpioCOsDPqqBpFsa2t97v5F2m5A7YyjVv+oKl
bWQMBtrSy5og3LZehDn6klgJhf23CXI/mOYGLda6nIJF+72IVBs/wEIQ7/5fXap2ot+rZaWa7OeO
zSsxkwrf06YP+VXhC5pBlYRA48vhALJw5uMKoYPtw3OwoSMh6Zx+Ws+Hwb5+L6ej9VHZEoPl4Dye
noVr/tIAQ5v/y95Ph4Ms5rsoQTIuDRrsq02IXusIFtjPOgokWVkPZQ8ff5sDhBo2N9JEQBUml8Nu
oAh5jQhLtXoVlMQmAV+mlBlIbIIhJ4Zyf4ti4L2ku9GQIDWfB1J7ojuvufVLAmy2FscimhZ8o+8p
XASxO+Ib81CKex7e8mOwafEpT6S3o+e4YKauHo47vGIZwLofgP/JdXtx78bvzTfXrWFdYu+xZ+x3
Ma7fy2lDZ+fwoUwZPiwcTcQLqFCeUo2cMI6JnnXXF7espNFexBXqYfBx2eYTVJXVq9t/ZirQrc8F
4LIBuCM6FOnTXPg9nu8pEh5WIotNiHfZDvhXp8HPGPYCw4EVxgMWKwcQ4PsgQ9sIpWuoSXl61BDZ
XfRkL1/ethcvjZSVdS6t15ieYRMMLGXKcknNpDuF3qgpTzrMj8l6uvIHXKzMDlVsfbA95pLQANK1
x6pGDMKas9JSqT0IPS2RER+dIBdiIXQ6jgv2XXIEAweWZHnVzyRrOBGjynxFO6dgNUvfFvAjN2oX
rMMxSX10cJaDWBAVA9xVfJz6KSTQ4sSRMF4OTA+1L59+/EiBVIKdOx6EQPAJ6Bt1mYC9WM2mRuji
RxPdhLw2g65tpe221CUEKZmseqObuwg8i4uC+kq9SIi5DxSEDEbnAtuIcFaTjoSEv/1lF1cLPhI5
9Hj6iaPLg6N8BbvGqfM5pMYOjqqYpMkCwnNd7+dniKOYRLfPQfUP/kEtCMwJEn6DRdUqnqgJoccu
Adr/ODLJBr6SYyGQfI8xvXMPJ/pP/MzAPjQq81roHXvBYtzvF50PcP7dP95kHPWeZNHvgj61lfON
EcQ/KEyUEQJ3UA35pFJWFNatmPdPqa9RBcH2/EsvsnPssv2wzeUslbeKng7Hbhmst4rHWtrd1W16
pROKAbwFVV3wnW/6N5pesNtKNd6LWgSf3sODobwqkc83Ra9j2QalAKY82HrB9Li7dqEvi2IBZkNw
Kmg8hqulrVd4kvDQ1GVI6WW6p2ccvM166FCyqGb7BKSwYLElctYu4Lp2JLpgrj5OlSLzQTqPSRJz
SkWX0VV8UcFG+6Lg/vlqFLfQNhOfgFv84OlMTJbAq2Os2WdxwWw2bikpgI9vRQY8n6HIoR5ZkaaJ
H2e4bUbI/WBVQkBFlRpA+tURh2CYzAT42896S3nKQr0rMeBtumLA/+jehHS19Esa9VB5uvReTj74
S/aJMjJ0qGX4ZRSOPflCa/aATA4vJ9a/UJBJoWXbof3lWmToI3nU4wB2tsWhf7PzE3hjYI0LzF73
7RuzZwt43Bv1d0hgEKmcGZFDA2yFDL6S0Z+4LX/LXFH9QyMLE0TVZliBlqKIDtLGYjSXogIyVeg2
c5B93T4CvxqO2R/GcIxCgttHwHf4jkVrZ8lVIVapy9DwhkkNhTOM5i/mwnXCdEZZ90nQjpXxgq2z
tDnm1WajFABzD6zgVvRdQvB5iWqIARPx5Q5aR8h3F9SH9e6Lo03V/DmDZPuQX9xC6OwGfhg8+rgs
M3wCR35v6Aklz5eHfXJ5hdhSCnAVvNbAceisFmd1vvRYJ4D6O352WbR00ZhNhUsdXv8uWoEdKaOH
ltA6sVpFcZvloln0rN+W0lzyIOyciS+8Z+z69vc/fIrk+tsbFX4ijGJZwTBdD7uMaB44X08QqJM2
bvmXAHkkQSRyBLzSQ8scbWG+s934t+5obYpaG4+e2Jt+r34hLt5qGFIsX+U9O8yCHbMoubSHmBXV
B1MmPhq7TXzPQqzjOa4cvy/gSNGjXafRLsSb/O/DEKnMjjWUnOcX5TNEr8eKVP6g5GfLNErzz/GU
/AytPQ7YSntaGnfKbXtd/roLGOmgxE2hEq6tpDan05IqE13iIpFmDSgAve/AuZdYC41A+LulbHm1
ughZZ6JTV0+d2HDTN2X1Mz/ApmVWFzSFEHStTkAfDIlAQAouSEyM5//0k10jhLxe4TK3kv8RBDFx
2dhgME9to2QI+tj2rYlR8s6iR69XLjEA7FVrZNzg8HmUiZgdyAzkP2w5wUkcP/rPyPV8PQf3i0yI
uzPMJqynujvQcaDHGSNIOOYg5oM8ZjQUmm2ubt+FJl8b58bOBqLLh0Fp6d/jsAJ3d223cO0lQvPJ
ZfZkGtdNm8tmcxYtmlZ3UFHwQwAvVhevz4Xco6Sy3S4oOGWgwVveUbmWntr2vy62Nup8+eu1QeZm
rWRID9orkjpPPy90Bo4/sjJ29jBNB3wkvV73KPybKbNfc3el4uX9LiOLDG41HhtXYGdsd7nmEb2x
7YL2F/xLwqp5YComGCGmKAKqerLvZyfSuurxwC4V/0R9CLJEp8H9+SkOcO6a0M+NkxczH+uqiqz5
FYYSJh0C80/GGKnN1Yq7WkNeU1IR5xnd7uaJvrk9zBPszRyItByyP5yOUWGcZzigb5GHKvfC9WoG
8VhleFwZLLsgM3MTPrIMgYd6MLY1WnEqXHgR1Hk81SiVhdt9kPAvQprcvd5pULDjnb5MNszlqPFT
RiDy/6DcZQyzvZzGQa7unbT1VIG6r55OTBE6bcGAo/MIh9di7OQKEhNlwS9Mm15iMm7RR+3cXa7L
KvnsTNj/WjZ06d6DWHuPpFz0/CtOkWrtr118e34oaZcW3CjTDwGFaY9pi30gg6c43uwtFOkgRtjI
L0M6FrZ1JOVkmhZJdsmB8XbWDxVK1lxUUPiZK4FWPH9NeJwBEKWwY0YAu84HaFwgUwXh04kAUp/N
pD3/MKO9VAs7PNeTeq+y4/VqQ+RrCgI6FpYZ2+/da1V5yyGhcNAI1QCNW7UljIX0zEWL/yamDgiV
kTn0sc+SONkJp7gLGNIzA426zOvaDDsbNYtevwn4DkeJvR+zyG1QqKjEdK/tbNFZTlXqEQttCv6Y
1E2Ni2ptlHBKnGdipe0kiWYSDeag/ebG5Sx9qzyFfyFdzSnRCegTJPZgnvVA27kCCRrI0nVFpf7H
hv2xBB6cAfaTIcMlQTpw/ycnvW9aK6DlX9R5QMhNUSkueX/JxZH84DhKJpczos5Jghyzkqg8aYKV
4C3C78/6j45ZXz5rgkUlA02yMujYdyBgh/s9k8/lfCYDJQFLjNtVqfKq+FL3pt+ATkJrWysu6aJg
MbCsWkdkw9rBjh0WVeZYsA3EAYDidejQPSICkkI5yFktklz+i/iALZHHmVpOStaUXRpGBwzXFhYF
5ONgT7gper35WX8eLJU8637gik2tPg/3DT6DRLYMo6lXWg/Keytoxtw3uegHzozuJTAPc+ahQE8z
CTdqH5XporvrOFuzaHzBQSGPJ98fQEXo+Tscg9xvyPdvXSp2wKBpC12V1MBQfA0mhKV2OcKXmfYT
0qJaP7/t02tTGSSpGPzBF8qi88P6hcolqrYDzJbQ//0HwLXo8kRTlZZm3fwTnUfWlDJH60gY71AT
jpPXOoKVnzKQ41JpujubWSCmt7lDhxV+sCJc523rgCMUe5MZU0nK6KPeHe5UoKu+sDXSxcslKofv
qU13rcgptJNyWamMkTTga+m2E/VR/f6unA+bgJX8dcrR8kuJnkPrpxyPTp2vj2o+5MXxstALh7Nn
rblD3K/KpiusiJeroI81WvoDrQ7gKMiavMyTAyvM1qhSOeA/bYW0f8eyUndDTzyNAsGopl5EJw0m
TbHJLxQWpaKN482jxd/HkIoA0URgArecEa0te0FdihVgrNg5IhCV6afHX7/6XWpEYruS75QgylSn
ZFZCMMVphntkmTrQffDNODrC9YLIF6o+lz8QHMBhEmv30xk6OXp+EHVqGtm57Q5K/n0iPMQDsFcb
PLmYUY6ynFck+mfyNE3CvxRkhiRVFgFH6SaAui8CNQAAnw2sPOdOKWG1D4tC+dFftfBy7kXIxSnR
0jZ+HPs42Dqp/n3biJfUcgIw4t6dVwm9sMYWRDLBIEqw3RxGQ94DXZArcHbsrdcsgvVTov1hd3mm
mCOzuyGhmQQ4e6YepaPMHIMYfm4V7ZvrloTX+VFIkPz/ANXfGnePJB9UM/N5MLXA91i4iLU+9YWe
+MsZsl3ZhjNe26pUqkEoGkjsyi2wayabSjL0aAyNZVy9CNJQBsWTnmvGI+BPWlLEjGAaMe1zmWgh
Vs0k/JbpjCvsQNDycbGk1KXqzF8lLDh64Wu8v1PBA5colwRYC6k3hV5QUa2nqziFD5XbFAIfzVXW
vOjooUvI3cHSJMGKXjCkEiMsqE6D7Gr62xmA232/Abwxp/yzMnH/eZ24sB+SPVL6XZ+IGowhAvyW
K13idNYWGutwZSDfKLkuk7YkdUsxT84Rsk/6/nyN4Jle5BYCtKk2ePK26tO1Sq1C1J5dvxyvPztG
vzWSfvqCAh5hYFIsjVkhze2Dk2shNotxNi5SCUG0TepZOu17T7GeTBUxmmlvFwJAocLNoBoNByx+
cyVnxnesEDpldNZjwDy8De90XfXTTYda0KZlw9VqjFE9zhYW0Re+VNUG/OeUwx991TWD20HDtYwx
4iGlLYNhsuLFIj3IOXZio1UFn7LvzavSxAqIgULWrQSwkJtD59oYsBCDST6qUVNjKq4Tm4gGLCQp
KWaHtaBisbqc4bNV+NsiMzXTyn9hu79l2bOa4CHynpt00TYYf2hA9GJMqX5/lCcRJZADDRWVo2DP
zxhNE8GVz0UkHNc33JTlAeFEf5w99bDTcaLsIOK/qdgFbtVF6jKSaQzrW/dQh+58Y9VNo5AAWDrY
o/sr0CAYD9aKW4VZgmZMp7/6jnyuPTnuabeACUurDWo5NgtS6gdZ/za40vEUfmsxSbsD0ubINQ5L
qNFkMMPmOWnJCFOkZMcvxpnbPZOXU3b6t+RNeY6yt9nmNQ8kHA9GQgJBAPbrurq9gVAp2/g08AuN
e5yoHhnBkHnNqkXJ8GFWQjCCG4qBU0i8va8obfdufPaRuq4E/zHISrjqRotchCGUNwhmCU1t+Aec
wc7M1A3eFRazfo9pgM81f9LagSi21UoICwt1OztkAMs293Yga6SPtXyH7nVvXo2ExS+vhTCq5Prk
Hvf8nxujtNALYGmp9lg0pjz2cs86is3yJHqZFcDSNvF5U1gpJx78DEBYZmylZr7cc/gKwHTV7BAs
E3GQQvogxK98vTWjrUdkAV4gdhHb1VtEgZ9VnAX50uyd7QnssUWDOMQTSycVBbTor5rLFs059OdD
s4whuC2RIsx6oqS5V8xwO09M7FK7AcQl3r+tD0elb6CfTtfTzyZcWYaaZTh6hqtF90RCfd2mo4vy
3lm87/EbBg9m3HcaSetaNeoiZG1s18mZi1bBABX9u8ox7YFRXjG5btxMlE4fYd9w6ThhZ4WVBhO3
DMh2bQBLilEG+yrJLlF74dSjr1nWPQmDc8MAX6laGtUuuodQJtj6Meqp2KauVDJwks+9jJ6KnRl+
Rit5sI2HIfW5+//z9UmmJs1gyEfrD31y1yRCVBm9jAhVjrno84vC+r3NEVD+GCIiM6Zy0GhFedgG
ZnSqf/YE4Ysgj+JlYqS1dulaVnTDc/fRG4JWcTWW5ifr1kcL89ztBCeyH3rUFiUxkylCjhuRKyJ3
59m9c0weAO1B1aer3VNX6VDk86wHCH3+/LH2Ar64nrOyce28IFEUAwGFzwmApTFV2lOxprrgnt+V
se+gj8QK0keJLZri//bCxzva3b9257f65kogenMsbSC90X9gtyUnL0F9Mf25r6C63g2rFBinrf3y
ggf1zLqzT2CTsUuyarR/TYkWIZcrf/TFnDNC4Fe8qE6zlsWG5m1OB9jmJvAfl+Fd+FPnBiLIweAR
AQBxkqVEQo2GQ3gTSHMa/9kQH1W2g4Ldj4xIa8vDfWKC1QbU+sg4oKHHizpwIyb9jEmC7UzeYes9
zMOFoo52zkYzNGF9teS6qXolja5pDi/+Y1iPhuTAHHyUzlR5gwl7z4dqFHN3OSZD7YFaWyf+Aft8
whDQiQs54n3qE7ZQgVrQLUk0vJjO+WMjPsh4NaI5zQI3YQfkSAlqmfyX7IX1o9n8jh8Wik/OHRdE
Lwk1VW18UgfexZIBwfXYV/p72ztwA/lk6VxnC+5XIDZ5Eeq9ZWcQF26NncaVqdSOM5JHz+3g/wF8
FEU7R9zOm64X+jZXlcVFkSiHVvRnjBxy8Hm32iBvhCkjLWfqjK17EoUkjfBMzZyKv3N7xOA/YVWw
j69giLV7hiFsSxbZD7QeyzYXauFHAgnaVvwa4EG4x/uNqPLgJmjlaARPFffmiD9hGFyOlbtPD/Ec
/cWEHPUpMtiLbS9S1vPPdWZS5igWX0nl5IIe5H4kEQ1BsfHzFNE7MPGhv+Fkj3lVKnuSDr5QQo4b
t6m+0tiVoTYeJwJR2PH0zjP1b6FDBZj+xvHSMfSQR0/UJhGF2imtR5wHDRZG5j/VpraLUqRaw8Eu
EKvDNde12OoWIhD79RHqaOej2Gg7MxsT8yJNb+ZAV+ux3h6HPirUgD+SsiNNEPG5NGQ7x9lPqLmx
wrV+KRYe2ykLgFW++tAR5bPgITmMQjmCmcANiv3pWDOu8YlPlQ//yQaa1V99XX70uVGPSCq6z5f0
Fg9uDDOqXYG08/16VffgTx+3kOuxIzfDf88SW1s1ZY2yDidR8qtH7evLzGAV9oeo+p0ZSzHNDTb/
yMcHOpbZofW5B4w7+GOV8Tc/pCVK3KJ0bUqrrZ9YbPd8810wu7G6qwnZU0kAAgVHNuOZydh+wuh2
31XI9gOUoH659NqyZcu42LFcc1Br2FEHDxQfbg1t+Xo1Pl6+dEHz6Ew/b9hwrY5i//gOQi1fmZ6C
+WzcSvTS4otX/u25z7+B1iB3Z0jAbB10OuXCh5rYqw/Tuh4o+oaufyowUccZDYjrqJw+Efy+8BcZ
Q/qFDrhHMP9vuRINlgJOzm2aXZZhYcfcasmlRgGj3d0xLE/jibwsLmngAgvzz4M9yFPJFKKARPBS
+hm1QQ1+ClxBgCUzc4FhYvsBt5HL1FRa0aDbi4OTIVMRubymalKWr6TOFc+99CS7nuhnANEjmRcn
S0VvQM2E64/tIq1JxzXkA49Bkcw3CGNIkN9lb8JKhPF6HQ3UMzGrBRBrwdfUTI6dV269Z0CYIprg
+y3J4lv4v/apvVbBp/B/Xo1wOOn7uVbvWZ7uOgY/OUa7tl2y0AZdj8rfxZY4U87F7tklweFo28VZ
6kVJBoLAqlODgmLV+7oYukVGSsDef6c90O54WBz9R1P9jaqpLrxw2yOnzI8LnZwmRuKNjFu+vKUW
hV6wyU7cCHESIow9QyHQfICJLuWZx6Z+MhY+wo4AZVhEWNfssgoQrH452TVmgY3fHaM80SgfV4Zp
tORQIH01eaUNwdqCnpkokcX4JEo/1L5/6e4Nd8yLE3QLmbaABxr681U8c7N5hx2XdQ9WdjM5RqVZ
zyQMInGNN5g005wnwPZJjc6puGqf0kTSUhrCvRcirmABmVQ/7oF6HUlX1eMPVdmSsWgKPaW3nEMB
SWcQxgDtkb8xI35XE5hLOzYBH22zQhiExhR4veS8KKTmTQhvlbDXdzFygNfN8FqrRReq4ZMLdK8O
dbboS8kD48fPH1tzrXZpS80asrET2eeoKorJcjtXhkEO1zjTSbQFyJ9ANxSaW999GJB/uWr5S7Ol
b6tEwSBjGgL+oNehMR0AS+syjz4IXmESoZh861YXgpGq50hRQEE5QH3Jw/atadlu7U00XXZ/ioKa
0y3m1Tf2kkkPCEmJPcoUwa19SSbgWs0nT7YkxjPhmd39tIEWdmTPjTnhiUJXlyD72GHgqnOrxuQV
UaAVJw9l4YQVIv/7QMOTUoIaE2K6mszKHkWTUorwuYl2hMtYateAhd+RKACGZLHNlvLnNGvrQR+9
FxetRXrxn0MV0pE7E7y60UJXiBr6cPeeQfxOKjv7OB6BEGtoBCFA8BzCac96YhxP4GgYy2VwOdKk
U7yGWngi1re5Pbla3MxcYyoH+yrQsngFO0lWRGG7CNIPFsMO19QVfpON+mPjYzy+NrsMJkOvKwTO
5r1OeMtMcDjbVpSrWU9ZGso2Y5PJrXjl0VhAvgaxpncdEhUaahbDJ6alMIFImkxOPC9+1juuskLX
CWZ4N1jfGhFEjNAItAr/D7DMkKsR0jBecuIn65N5K54xO2RVigZHSdWyKH92QNFRWVGOzsy/hN0E
hc1bbsYSqM9IXeALjJTAuc7s9a8S7dhQAoJFlkLVSUCyqYFtkLWt8TVKUD2XRI19wT0V3kq2iUPl
PNW6YkMbHeHmFIKVG1odETS0844ZfU/yfIHFk4s/jGMiIZgyJyZXiqEO5tWrX+TbErKKRmd8Xmbd
dmmkC3+wp199AZgXgPqZXX0q8pVA5ZYY6w9vdt+Z4HTejlkCkj22JctmQRvf095Tx9R+xWdl6PD6
j7PszEnA1lBX54r4Lfyir32FHBNKKOCXN7erUrqXEtFIS0FenKJVriH2+r1Y8Za01S65g+K4QjAs
bRD7ax5oSm6QXhfHKwxcfU3uYKZSmtcBi33dLcoP2/AcbJWcv8Yd/UDh3fCb/xYtBAgCu15H4r7i
Z/92vVDcojTS1K1UVHfhEE4l3/ZFaC5Y0jDhk3AL669DO1QOc9d6q8ZIIEyeEtGNLSGVIRbfpLKN
uTMkr3wcA0EaDxcNAHOSwrXjjqTzW3ftcFCPsr8P2or0YpDqTuFklggA2uyvr6ITa1cmSzsIEIVO
rpD8mBqIOGt5U+p+R+kFW6jA3QWgBoAmOtlu35TNa+QnEPwKsHHmPyyTNnR2NiLbG+64M6yqN4HE
juJBE2I6c0p+ossBwSxiL/rjh/AATq0kSplzP2n6k37PTeIZBR9FKtQh4ABbxcu7nlxUbEvQpNnO
wt/wnZoYzWrNlCI/jw78kAtNdZFt2g/KRDUoF0HNW9TaVO7hEQ1A+aritT86xM7ZFu5+3hLKSFFL
VQFHxoJT0s5Kd43ad5OA9qGqqp3Jpt1oC7PCtYO/Gqjrn6JCqLMQnDvAsLOC9RLbfs9fQGH7PhBP
4SCThD0LYcwrSGSiph8OYDs7BfqGqT+O0e+P5fK+Rb811zugZ+q0fc6DrCbcIgv6iiSpvFL+fn7d
Ff03LjZg/GuHGdFCN/y2WUpEcKBb7LETAJihdi5hGIJRiHLs8xSWr91a0+17a9Ua2bVrd7tBGvrq
44C+2htkUM+HLXdyPj1h39g7mPUq2Gva6Fg5Ug3r/EiO0ZniBUKxSVJWZ/R09Tvjc5Nv4UdXydjy
xOSRQm+UpjThC2ytwze+Wu6sPWACejAyV25k96NOS7klkOxHYq2Be7Dz5lEkiwlZy3VVrQPcexun
Nych4jgDVg/dJ7mowTBhacemafGmu7FhahEGTP14wkNW6taoWzZDWmu11kt1wwydyuUZf/k4fjvq
JP1z4aXnpD6VcocvV+muwj0tL0GGBy02YWv92s3aN1forNqRDBrah7UjK5xMdPX+W19yzwAaDtsv
gBXxp62ozp/DX15uS2qXODPw71YReFT6JpkkBafzR86hPlopynXDE0mBOh9pMiT9/WBVHFmvp643
0sv94KBxZPeH/RUAF7yY8Qr8CZttn/Q1KM9OY+VO5HDRHQ8besezSGvcav3pDttTCbIrCBaYqXk6
P7MBOKIg99ULNetsBM2EfugHRq/CncljWsH5fMB8KeqxVUQoevXoaYGSVMhCQWy2fbIPKrLRLG2s
ocUjqOWUSwobUrnP2xISvJwhVjhlzTOz7RHK2EkloOv0MrrMkwqxlmE1s3aQcBjUrDKUP9o3bGGT
hG4gmy3QIYUwxZnwyIc+9iP3Jru+FIPbfhLjrAMbulQlvnrRaDguE9V/dUn0pme6yHwxcBIMpq7I
o2CCGMsH9TSfUKJ8Waf7m9FU6S8/5OC5hw8RQjl1Z6Km2vLh1TwJwNQD7HGgylCR8zQTzzF7gSGl
mlrDGkUgoYjQyQ4FwGpwrLf8U8U/KR1Xf1TnSYeNiIE1FA6c6kQvEFzQpZmnRjIduzLwS8uapYIo
Lt7sShVfyU/pTMCC5jDi8wj+qK2ZCgYXC/DElL2YTgqqsonXgTCxqneNyOdxf9+UsNZJrWX1t9IG
PSyvyEThBfHXXhUTAFsVQ3Qglxx3AdY89L2VvQ3N3MUmNyXbiv7SwZaZQcyrd+4zkYLYIIsbJbtg
7VbVlVBQQRPNWLebh6g8qWdGKZHcvcO5oGxNPzQAgUu1iBpDEUXNWIZnQpzDgptR3TBwk7P4HYUE
siG+BWANOWbUpGatHdsw5xV+mzBfDqUUWzzXjVfjBAFO/Z67OFPjpsVmN7yRfWGf/U0S+w8aIs80
HU1LUedqJxjY08kLAkcWEj9yhQFxS/ncXx+yDv0ZWXLxA61EVRCL047wpsbqLOSLn2Y6ygG3Pzjn
J2qSTpLfHVWY8nlzcD65VNG5QZxlUKDid3Oe/AD1Ef9W9pWMH7NebzmKXpsothiQEPtUNKQeBDgV
A6tSuCaisI8vSoadWCZ8FAmxSps4vFR1ov8McdtqC4mPAtFm1CsfuobZ+InamyZlJXiU4jXqJyE/
fNRVZmHONaI61pHOmzS0b9SFvZ3cNUiVmxvvw9aQ6adew3dpWjRao/lTrtAbnnjgGRkpe30ZNbyO
adihXvRoAme4oPCeWkMSP5lEoXTrCK4y+qUQnYv2MXUB14/a6DY6w9xjhNrwxXnnYfygd1/PpRt8
UUkgs3eznF1VDDyq058ktc4N+z/EQH1btLFqIbd4G8pjhk6ecv5N87dwPfbyjnw54sqK0YOpsVlL
OIH287TEyb9pLQH6F1oHbGRWbipIdORABKvIbJGYrMLYPpU/2BlygSNEcW7xrbnONJx+L1ahQti1
H5iiZ/IeZBz1jfIaOrtAhEIhrqTDgX5zhL33aKEoQOOkuA3cSjzVmvGV1ECnwn5xOpTEfCOXIloM
VAy6tyQmigsJXhHlslcorkThR2Xhv+IbeHMFjefOibj9JaZ33gZFEM0P6GxSv9mdlVqJvMhmqgt6
hq4JQxUq9OBBSIcap1PX95cItvpDpHxvxEMw5xk782rGUULwEggQaHBK+hRJKl9VffzeVh56Z5pb
PZhRk4YRtL8kKZUqkRGTkhdr0xGRo2r3vr5nc8YH/sUlRBem1pKN7XpOuKtWQcGfNZp8tAvoTmjM
dnxh9nFX466/0H4AH2tD4ewxc95bgJGWPBk//4QPoXNrcL8CrlfEMq/QfygR/twnpc4DBFJMxdWi
OHgi7mdj4yW/9w99vWmhzI7zYDo3p7UP4nuvhXJg60DmM1xJsLzTPp1gNtgVQrZp60JEsjbe2gja
dCnlUkurYxIRIwmBjryfjC8FX36prEZEtjbxWn59jD9SOZKa1DP5CXt6PPMkRswIRGwK/Di2i6g7
9E4dpHMeZZSSQWatXNhPPqSQVkIqjmxkBVfIkzmWCEIjXQO33Bs+DSEJ8ytYBXKFZbdzlhGBi4CB
C6ywq36UobiLRvkZmnIdHliHDqlQ6ZNV9wcnmHNcP2vv+dw6+u/rnucUoA8r6TAT4rjYWET3OFnU
yfxApA98XRsu4nxjLQgfvaUVVr0vuuiprGzqFHy+M3kot9+iwQGzXQdCpXUGr3zDsNXCbPYwWdIv
b29JNcOMkdNnJMr3mAxzMgmJy7DsJKjxtfBQflWrinzzo5JbRhNYXmg+QE2Hql105Pbpwq2EZ7bl
5+n0lMNMEU2jdvXZ2NdPcvzlMtTMpiZJjzry44qztGU+Fkh1R7mYgzNNnWJ/NWE/3BTki3JdzYpC
MpBUuTpJkr0P9RmZFcMF2OlDOvn67EFw11U8ZJtaOnEEiTN/phgLMLhhfdVUUcvXzaI8RcTLBaYc
RGdT53yU0AMj60ooENYUCOvYSBBjYlEB1D7nWkKbZXvrDPpAy6nXYqOa1nMOPju1fySeitVPmDTH
Q9aNFVopKV+QF4Ezdxwk3sr/Ub+2Awi29JhUfpIaD3vb1/WRDBDIxNP/blErbyOXjObizlcoU5UI
aeAxvidW/c6PFCDwxBsnRxgPJCR1VxjAiDZNr7e/rwYGpWTQ/wrcLry8Hh2HoWgrdoU9TTrubg4B
0l0RZzuHy67iDdsvLqdK15RsZmrbmyoFTGZxCXl7TFUQPF+kKmnJZphGUU5d4nSxDVbnVl9JdIZp
kfzqlEYu/GWovLEsjR55zBIpFGEGEbZpJ2XA6gB/zXSbKmMaimmfSxYsXzgf4NFZguev9fQNmWHl
ITAswuciFoPkU8T2C6DDMvJESllu6ZqHFzvOUCngadlw2DynaGo2duCxK8c96z8B/q6DNekKYXCe
Fw39rLsRqnRWYIKGseapqbxZU7JZlQXt8IlX4hQNiblMbRAdzGhEYHv4sHLgX/pEf9EvkX/RHTGf
tZ1q7nmDjiLfeWkZuJ4LNANd/P4DA1UgOxQnN6Bf/oyYUgIycoOkkkTatHtsPv/SV1055Xu0yiKb
b0UVlX6IanuwksR7x38Ji0x3bZgq//65b74aQDL9UOZsH3ZLO2CBzAYt+AMsoGcLxz1SkliirRCu
iGc780YmbiNr0JNMvbCodLabguYcTU/aMpcbCPTRcrPSiXMsVcDCysidmTT0ST7uf0bem6sx5l3t
BpXasfyiFHKYaMRNymoGdfA43Dk7YhqJtJb0lsiAdPFgvN+WLy6LsQ7isu2NA1k9FW4nD8Paxhgw
ziqQQG4lm6pNCI6vHC94IyqeZxUEa3p1yxY2MPSMrhliaoR3djlE+78Lzkxaax+mMjcPA8nGmn0z
QY2RsrHt4Sj3hpl0n/fiFH1dwKD4O88Rwg8+12Bcr2Tz0kV6OsN5F+IgiM77ERdnwDS+/OKOUT9J
Mpd5yDtcakUzXdMfpPgztJPLC9RqC2l24Tbf95Z5qTXp0SiSAyqQTmLtgqiAV2a4UC7QuMwnzs00
QDyoXn5lP1LWKzLZ3bskpsnoCMgb3V1yOZdgE03wfw/hyqTwLnWtlGZps5hvAt02Kc/KMvII1SjM
t3sY+wRRfynMqp7urgrfkR4xS6o5Ndqq9Z8QBf8gNt4Ncp3RwAL9ZUrdVWZVF8ie2hmggirLfkfS
OONNF6k/qIU9FQOKRfe4lH7P/7p86JR0ozdhq2liS9VRR+euP5KD3gq7rpPpi4XP8rrWbjMnpPCG
IXETBXSRI564s1fz6Qbd+MktiyUkEo3nvA5dC62CPQYjBJ/CzKCkGxnV0irwEDUyjZB1lnxPbhSB
TQvh38Hu8LIFTJNEKTp15kD8jCGrdX94VrGrFWyrvP/XLApOpRUuinT522FswNnu0FfONhXqHgRy
zn0e3ObwBx1Vnzpg8cn35y1HEscjtQEGOJWtPf3SodSPQTwYVY4RLpv/qW/hysjp7WjrxqmeXxjY
S8D+3I+4DtDHomQTQhbcioKhBkLKaZjWkqWBmr6zpMIfz+7iHG1ogGmIKTCt1vFrNnJ05fSjGNXT
l5Xj1Pci9mMVGAwkxw9uGsyGwxLQk4sGEUlxFhJNhNOdNP+LyLfIK55jGZoTna5MN3HaEy5ah12f
+ctpPF5tmhDc+PMD0advKApYuiXNJEUc9UkZYBIwm4733CrNRx/KyQWaF9/G4OI+G4qEpvOlNCsO
XYwBPHwZ4JEnHkjaxMJxQNZtnm3V3U9S5vtOJoyXI5gUtUAosLCCKtMLDV74GW/51MTmu8I687dB
hR5AP8DS37V6TzJewJsO80HPoWR+x0DcY21N3vAImsBZKR3Ac187/ok6dRHU2eydnPDJmsuG1DVH
1ruhdAXnQ+Qe3eJE9EsEux4XZd5BHuhiqEJgFHhoPnZoQ/O1yEnUezqw6HM8YTnQD6kNaWiQVaJd
NfjvCXH9aNsBzfyWW2tbGhD27sgZ0FGU6xeeJvRoN5fSI3MCvbltptfE/+cKpsFmpXm3cCzAXlkd
x5Y4qPq0M8JilEe2O/wej3doTNMbcYqe2cJ0Y+GjtRsQIlky2n42coJ4Md0hp+fDcqQYBgsfFbvM
DqHNaJ0mWHgmnb5DBGH92EJXKPzdL4eTFYYLWNoC4onezi5eD222VyikAJOUoJykMwgrHoTMYBLN
4vQxp7ioTWkl7Yok0Yi8kK95mUr5jnZbCZZdUuf8T7Yn+dzJSwBPA8OwtUGaaTfBjvL4bqfNdGA9
dMUm65vAEjItIJ1zKDKnkeIsvrAstu0Z8sc5vpDALlVTbJe+iQ5XM9fr72LBZkCOsA3jslO8wF64
B24OpzEDq7TE7s2jTbYx2t4IplO4QnqjluqvyihIBlIFICOPXzCrpomwZswiaLW24hHm5DNuaY01
mXrGnrhrWasM2P6J7Jk1JRKNufcpknsZ8NTQkY6sJd84v5cE4GpndqBlFwSvd625M78K8yPo8rDb
OiBuRp/Oh4GOHzeyDudkY1lD06zEm690hR6kNNFvKU+jbwaF0eOBE6+pDXXYTG6mZlnz4KAMriKi
l4lfRbhXCSI/McmD0c5nq6w7OGglvRQHpwM5OItcK5rdyg/eRg+kDwQj0u7h67FuDuA57e8ri5/l
7dnVNVvXFcZPrIUP4kKyUVbW1PTJaD+P/3TitXcuW0el1GPB6Ndwc7jcrjJx9KY0lf6whPHQQ25l
syOM5aEPyjEpu7Dy74wSm61z9qiUfy2N3Di+OdMimBvFboEmRiqGAJVQQ2p1/SDGzrRgJRu1oRli
ubhWVYGRuMks+wfVCZTXJvJo83rObMU2I5IgldqIzsnpAfOguDPtS3MMmToZTkvD9pSFbC3FZYLd
yQI5dzSsyFoCHbgAQLqOOahZvPOZqsXcc005q4DaKgSqnHWHlmgZeOWaHljUpZCBn0xDHaIxwSu1
QOb7aABh4fW8fCLNv+t4iTiBix/Qg0FhVmPY+LkGlSLnNmaMRwmoBg4+Ex8HEXWhIhjQRAR47m5Y
/U//xcOiEZL/BdrfdcXYRKsdK/Li+IUhXfK3Aup0NAuVOu3uS9W3eTrUBFy1xhJG8nU7AkFa+9Ar
GEJ7Oe1wTIU6oU3ozLZD+SMnuvoPqlaZfyJnv7Va1Jv9ehDSXDtZf+sdc44TIkM3t4AVI7q4B7zE
EhzkyCdZ3EBmcGL7GWJDVmVnQit3mFzbtzQJyscELWmBxEq3WxMrbXV7M+iH/eIXM6wrmcM+CFxQ
FCbCfMjg2mfregw2Ix1J81dL6U7RkCdwkDXq6CdJ5rB3Ti9ZOE7EMrvXgNTrafT6oaMrSCIi8hp8
/zKE//upIX+Z5bASPlSB/cW5FQ+PSNQPi7z3joc87ynXEw4RfFowlldEJu5ol/aum3PQw/NnY3TE
xP/I5xRmy8oMyrH5zC78T/TxnjWHxaeF9IbNl8FOHv/MPARwp5VbpcW75IZbL5+Qa77v/1MS04ML
nhmcjgSvbpcNkcWdx487f/Bu8GvRAiFnVObZz7nvLd39IZMcXrEq7j/PHt88FeQUgTLClcoyPLoR
zgo0lKTBXoFGxXX8wWFBKdM5zCIu6w8X8E8kr10p0Z/rbVntWONJ2rjulIqCc2ZD8eoH5RadfN8q
8kkZSLuFAWqVUoMlH0DxU+deDhfxdjczJHYWQ+W2cDY9yF5yb51YY5Wuy2r2DcneRr0cvWVR6v1i
pp+65ou+aNc+gwtWiZqyt+oOh3b2ImNftM8+JnRAjNyyctk6HoVF9mHSaQQyBbEDmCixO0U+wG8k
kjZDIBFQ4CEhNnX7MLUj9A2zyooj9EZ9yCRQT0HT0G425jyRIVhjDfPxKEGF+86P6l31AfT58QCD
oC4VmSOYpffuvC7E6QPcQ8a+NJl8Qm6WhAIzvL0B4N6LL4BFnDX3zgiygAnUiwZK89bCglMN4dqW
Y6K4GM1WZ7ta0A2YGZ1l+oHnKwGqUU0skWZOVyI4a97XW8uUvPnd1Ove0oRvYV3deSypVeC4dRs3
9fduNJa7vW90kS9UUGLSUCAReKiglRKdG/7MMIZm/PXM28J0JuWbxoIbAeCTOFIcX7ro9t2yFC52
bQ57glXOo7zPdwdxdMDirvLHjJIJP5Q65hln+UmVX37nn9s4ZA/d59h6WcjFmMPB5WEbh3BI5xQV
hI9maTAIUiNOMQHiWIakiD75LHP8Z3b96M8l5+aX9ONWUAmu2o6XbIK/XpcPpFvlrG8fIkZ0s9F6
ZOLy7/1Abzow6+jCNIb/GH0InKGkaBr7EcOmjQ5laMZtZol8iCdzpt2rP3OaKcZBhvX0TYO2y3sB
jWpsjTUoz6gaZTqmQnKpVvXEL7SVDTZAJqpxoPMD8Z7eUeHrkcvh+rLHu5Io3PNcldex8UbXOMWR
lIL2FhXSYoPnhA3bLCwBwfX0MpApoGd3OsTWr4nKQ9VE1O0wytBir5CsEzGGSLmj27MPnuqD1hVW
LU8m3WZHyd1vz5YKR88atDtOYLWzb/lEHzGxKaPZ/sbqKRvPz+PomXoOt+DGIIBdrx24JoKaAN32
AlY/Usc+fNqC/6tNfvDTYG9GGBQhMjvQ9mo7bgd1aLOZufyCq28TCZLFUyt6GXIGFdPmwlVGbE5Z
Db6fVEEaSb/jJdTPwESEd9GP6r3BWT58/BJ6jVimf9OimMbSFT50ba5iW0PrT65dN2s89NUqREYB
S0qC/X6Z5yScI3/SJRdxh4uzLciCyVtFm1mC3tIB7mErngG8kWkd0G2OfJFJ+RsvTsn8IMHZgZLB
SvtfqUZpWCDLkJyt0h2IdDoXgtqsj54+S9Yb91UGjEGAb7a0d8pPC86/tSiGBGH6V6/FBaVbxqM0
JWssHjtDoqAvNBMHwN2f4PsmHnxefBJktoCuiv/ZiyaqB5V4fitAOBI9R4fIfo7PrnmcjwBEx7NU
oNy2bZQoLvZ7Jnibxa2uHCQmMs6TajTSyb2gwgbgw47vd0OotarcC93dUl50EFbMxlH7kT2A16A3
33StO1cm7boGYKT5q4vyAioEzSEcCWV4Syx0nJH02oLorOXYKVjyk+tsZaWryJR75xzhhRFOudg4
py4W944TN8TszMwOVPw+VsdqEvCD6T75q1lxDz3EMLY/4bdyZYITukC+n+FWyxm+8fD5Nc15CZfA
euzFxLOgAIC2lxZum6s+zeMcbXxuXnX4Q8yxGeARq59njBehURGhjN7cf+H+X8sMI/F9jQXZ2p7s
u6r/vZ65iIqQnZ6fX06vuIjuGV+VpUkQkPrtHBd9ObR7obRrYKhZ7bIq+r5n691wxgqYbDqeWPYI
obt1vHTkEXEzX4ttmDZ2+TfrvEPP/XWLw6Kj4Cog0d6eX5Tz5XUvWxysfMJxozbJVlFgkALduPs6
HMcTWyh1MWvgFMuracW1pTMX/Z5O7MvlNbMy+bln0S7j0Rheo9SGrw6MSDQlFI2UC53TSMBKtrCe
YyqDDhJb/o9qoXumMfM2XgZQb68mVf8eoyNoYTor6U9yecVW1k13ALZCoG3bx/MTUnUc/W/BY6eF
DR7qO13l1tllQhzvESsGeyWKUc9X64hpCFS//UtlsjH4Y3V7+8TvK9jqjpXtOs0sl4p/WHEReftr
bOFn+uNZY342nk08yaSWLYOGyA3AyfTlNzqyN3b9jjMsxvMHLitg23qfsmljZbz58g64DgrWiCCX
ZhkVRs7OVrs/h7W+XUkt7jvK/g33vetPFR7sGguTmizwXGRJchkRHE7I7d8ewUX9p64AMc6RVZJX
0hLyk/ft6fTNRWAs/X7Cirb1OCAltwAuipVCwgvV/sex2EOmg59hY+J5UfC31el4v+wTrNZ1/2NP
SG+d8+UV+EEFAfxavDP4kN9jCz0kTdeuTxRvXGu3b6AgtomaIbfM4kBQHQgjlbog+7NU91lVOzeV
5A1CEX+p0jd2e/59JImsgqJXMoarxZqEAnNkpBGoBWc5f2pesUHm9lTbIlw2wAyOeWbjKjzSMKHU
+oF3BfUvHAEbg3doA6SMnbb5z4cuGLUiz5epfJeZtoHBNx3ag0pJNZttQ/ObNJ7SYimcCiikU3pP
QG1yj+VGfKQiunwBls3yn+a/oYRRK/wuIBrvsBaeanoF5CcIhtd5sYJUZIZ6SHRm/NEZICPeD4Kn
zyaah9bKm6QbDDDvlLRtV7GXEEpQIqERbQ0IPcwLSlp00KCxXnxf/hFJlJfwwhq1vGV4LWRg/B6z
LZP3rg5peSurUyxGGS0F+ji/ZaD88s/iZn/ksZRvfR737PPs/CtX+MvxK7eIJm8CbwRMpGlWTYrS
TpFZpLxhzirF3+C/wwEjvxQiUihKvosz3lmGEXNKcZRSodNv/e5AZfwWJ3q5XVZ9ySvNsCXauocW
8xBh+LEmFIk6Cu7e20f2hmK5/3rrAjeZFEaCH+PYFZtunxyj88k6Cthpa+BWzHIGDK+T0iX5EwTB
+kx0nCzNrYbuCYRqMzVqJJlKhI47o7a4wdEBXP5Q9ISMZvBg7LCg9LxlM7L78g+t8kPKA+JATKJn
Cw8ScFGw5+//iLkVZKYP+hlF6AjMaeVhhijs3VTyOchEc76N8pLL+iNKPVUP4ameCyqFoDxTBSVC
zCcIiUyQ3JrxOhiWyCcDcPrvNFX6E3zz6KZMAgzevqgB8FOASzbrxtgQblFzEBruxTGmYDlA8gQj
aAigt0KfT3/mxsxM9M6IAYTn8PWFLofEDkyxRlnep0hokrBpJXblCukkcSjHvChW7/u906Gq/2aE
KMgHula3H/xrpROqYBbylNRGnGP2zTEMu3CGp4zW1MUfuUhgQUHUNXRMnAoAmSUyklt2P7vz2Vmh
1QfKh22R9w3MZEndrWGC5NNPBbBwoc0Jnm8tPupaoyMFg1KqW5MSmp9b8yJOcObUvwceDF5t1ZVV
8Pl3JgKaEjCbHxgMFwrLo1Lsnn1QHB6ChpMH8B8OABZcqLCbwokdPUTyDvtR9VcpmVpDrpyM8PSD
p7kv6I6F83t3hPjPyOhTanl9gAu+4DU4xczom9RIvbq4Qx31jKYKbcGvcXS7O1xZmeNxlROmbWFG
Ox10M0m9RSOSKd516Mrki2oQ6eq8jWGKY+JNs+FHrzj8L4peQGYTUzikE0lt9nkdZE3CaO690e9i
9j+uPl4tZU7YcoU47Wlc38AFtohYlfrFQ0ZEqunNDLgxh/6AnTWu0G4Dg+GZOMod2JGyGBacpWlP
lSPUogd0MJ5ZFN5E/TSaze4DNFgl6fneCjg0V9q4LHySgsBysfal7SJb/3aDpnA5jv0ghQXIUSwn
KO0/6X+cH5inRcUknsVqzBaM+JGZUeC1I/MPXiYwxmyLxahF1+CgrNq1dJEVyo6tfwCom6+kb38k
IdztxRZdft7TFfqQXMzQ+n1ZUGe6exx+OPcNkyy6gs5elqqVzPpwAW5rKpm2nriwbdx/qqr+SMff
0AvHGuOgnWBKnZv9imkMsn2/YMSs0bGHgpMjHV/1cIaifx8X+hkC1uKwBiIhEi2V2csinvMxnf9X
OM94BGSC02Y+bj9NaUh9KxOnZY1RJlypL5UTJIA9DZxleO+vB+kIuSp05eALp6tMk7PDEiBJg5/n
Uvsrt+44ATg1p9qJKTjYe9PNGvxLFtuRLSS/04WQOcjmHDRFMBKbM604ptjMTGATVxJgyL1v3JKF
pEDz4H3b94VMTQpoGpqJHFEh97bszheWV7QurRLBoo/q3Yc+1NtHKKbDCa9dnL48rT4LR040iR5D
w8YMN94yeIiv0F2jUDJbQ8BQDyouv3rbp9biMFRq+5rZ4h+XYm43HDp917KWFxa3qt6/2kfUjCiN
h4XvgA+Rvd45zrIGV2IRPemHUVMjK1cma6c9++F604jPT01caWlWF4GaO6znnDx1wfvRbxEmrjT3
Smy/37bWZNxrBYGG83B4HtSNXp/2tn9GrI5zJgeTvuH5hsusJRslU87s8sOW/Vd0gv6pCslwyGAI
9Ns5QO6tgWzDy1QNHDboO2WAJ7pR0q6ttCbnJ+RD9A+rnbaV23JtEG0LYAQfbmEDRBchh1EktX5I
Vr+kSO3/uaLFbXzqzQel+/DqG1Upnw4pXeU364YK+E73JNG47msKkfWHiohhScrDxAoUMCgaHqkS
sWRE+AptPJ/dvKw45jICfL/1tAxexJ2QlVe0rhpnjO8DpQJ0NkD5lSTqOZSYFtG0W3rF24wCq7Y+
jGSUbgPQGVJRKCp8lD9razpTKv+5iNJho3w73m1rHzNPCE7qYt5O57wrCeOFsfe7iPkcYGlXDLWL
3IRsLbtUpst+rXnrD0oRYdGcjBf6kx6tFd6IsbIwF/4L59PAeBMgyKDE/3NSKy/XbtZYX/eGi6gy
4D720kKJCL5ZkXaWULnr/C6nZ9sIjWuCJmWGH6/miQC0DNIVILYdJhbOaZIiaDbFSMGp8qROMPWY
YsbqghGCrXk37cnChT+1QC3z8e8/J1RkVfp8L58Ql8aSzAYxszTqbSVsEj2YLgUbhnSuotWpPW4f
SMDNf6vHSOjEFzNONoO0nyxNOc4k+N3pCcruBN4+GTuEMV7lZV7eam3InQZ2+ONVFvhWXV1QoDkQ
SZfQzmQlSwuMLa182gDKASPiTsppCiwf2hz3qr4QtZOx46yEp2grhKBdPi1Jp2c2RhUXEEiesvM9
wcycoXiHp6GvpzRtVceAz7G7ZDylcHrJz3lc6eq1wL35NM/HKSWeyBjExX8gnS8ywe1NcAu9WOXa
qDvy16J8cU0o6UWCjfhsgo31QWsWBIQ4nKWmftf7SITqKTWYvli9cgBjSHVgknhgrNwJXzXcefkc
fZmu84uDXj96p+uNbbMBB3PRaQJqMD7+P38UIV8wVi2k+33FL0Ht9nJvV+DW/t0aS+SSHFwGyZT0
bAr6t0aR8eew75scoZKGvYylQ1+z0JslgRPZ3piwdIW26YLwiddSenHX9JQxlGyv4A57bsCVq2Fc
xLSdaYWaaimaZniBz04Vhep+ItzFuteeO2oDKrugUg8mu9c1Sx+7pRxmGe4ME244OM1P3TNtxjAc
fGTF+BVbGSAYzEVTf5ZhG3eqgRmEbnrQf/axwWHi/EwN5mKA2ctgGCRY+Uihvkjpzk+Zr/eoB0Gv
o6RvO1co3+mJ9hUPAhDnvmNq5ONflTUFWLd57wcfz7Ecm2VjgyruJ+7o0gVReIK++FnwwZvULugX
5ImvjQJwnt9K/uECJSxjv//tJaNgmrdMOQ3iQzbMEtTGlUCfdiPcaxgVYT7KUXOe1aLQWbMo1nZr
8lh8qLTSDH+S4nqFG/+C1rLiE2XOFayLpwGGRaJTXC62dQz3RKLmodj//wz4lcwqng9NDKqW5BXg
16BfD/jIppbfsVFOPaFIe0u4OMAr+PB2TmV1nbtR8+aiHypJQJGUqkbCgjfPnCCyTjwhp8mG9eLG
KmakkdYmob8i2KbRVcSXewazxFzJVOh5pweQLET98OWmaqBXJ/t9jaL63NuwWwRBQJ31ee4NMlcP
mPXjRcGTU7eVP0H6jLyDFCVGQnFvwgvKfhAfgGdz6MGQc9Gxr2OsifxWhpHOs7G8gsVs0tpOQTvX
AX7oO1fvfuozgqMCt93v7h2lseRuYMpx6xnyd7Yy5D7w6Z1mnjfHZICK1kL2+haYUS90E8jtABJd
52yVGAfltiLQ1NbqAUdvpf5dVLv7bzYHTbjBI4C7/jU4EPndKxsH06m49WF2jSxTnzWa+VNbfS77
X8Y8f5fFi5FGv7EFty4jEWhHfcv6ILKLaZj69Vfel1SqoEn2Foq25KcEaGEnpSYNJ4XOues3c0a9
w9/yOgOW5ejtr0Dg22bVCucm3wi6az9poV2OC/Y3n2ZVY9tTz+XyPaO66cR1s0N1eSQANVz3A53G
pxd395k67uOqzocanhe/EbyP8TarlS0A9FXW8dcF2ZeARURdsXLLXysk0i3DOPgpIxyrsMfbSvpL
5vYf8wTLkSjaIkmMw4cXpbr9kGDiViMK90EDZB0igkxQEtJIpjWEwVyd3vVA899y/UhY7LS8kRIh
MxebuSYDx0hI9Knljua/V9KdaOWoDhBBVsWzS1fPBn+PbvCl7aVsrN/a6L4aga8emFv7Vqyk59+t
KXYTb0hX8uJht6Bd8lPBzaSzMjSA5639jUXPELE7EsFtkQs46SYZMH1bsiY+G56ANQnpVk/qolSZ
FjtI2BxqYt3crQY3cLcRDM5UqoGtz4AcXy3tFkwnaNOMAktQXtrYXfwKmxtcWp0lWo2yWy/E+zcQ
ZmlpFDNnxy8P6xaQTen7EjWxNqTHebveBevY43iXMSJ92UQIlICG7eFMVrnDwjJvy4cWuWcF4h5i
nR6B5r2VXwz7XEo8dgvRuv8NPNBB9CRUOPp6s3cAIs6/U4Pf5ziIOyMYBr9vZHO6CeBW171av/0T
NUIJOjw8OVKheq/sJ3EG4Dp9tpKF05gLns5vQDudIEbmL9IJoP1yeQFS5GbtWoWH9sJPH2Ylq+yN
4YBUqbqKpDscZ1mgpN9gxrOzV4eC+kdoeiV0ijRuM4SoyLBhxMQWfH8+HrNDNoRvoOGChNw29h51
XxiMgvRZeEj8+MUg8JEE4W5ghZIAIM+hqo6k3WO53/Lhj6kUFiclVHgAf1VP+qupOszj5uvUPTqB
QJMLawzVxURzqpUp12st7Hv82zcJG8/OkZDjfGuGW3y1zYkgtU6xq4rH8lDLq1zCNzrgCbD7Q2qr
23rWyewNxVVKZPTpaEx62u0OkrQ8A9ghedcPjQIWCkvIU3WxcvCQD5KllXoBYh9YVe/5tEpB63R6
IIcTfCXzP1s6L6Vi3zufLirMNlfr1d1+WnNkH1sFhJojPhZlceHnMgGvRsEo9Xk24OPLqIGb+I+p
tMyr+Q4ZTSDWKA/QONRTMOoh4POwPmSrIPTmb9uOHsz48haXmvnP8ImDI0LClqMTUxLgUSuvHa93
QJT71C3midhXSd/cuVNWYuPtK+FmKXOgzxMZy/DJh2Vbyixx2q9ht46lTviDE+U9e1WnIC4sR+k4
S+Aw7N2ZNmExuwPAE3/wAG0Zq1MF/4wpZBXnAB2ZZqDT1KMD762zmvJUCkYINLQZM017ql+SvQea
WZCpcMuOcVqtbQ1LJhZ56Wj9Pz0SVXC2Wv0kh1/8mnaqZG0MYNhB0vi7hXuSq+FtQrDPNnniP5uJ
zi5W8MAORFGrf9aF4zuTSvSt5oGsZJGaNp8PdQGGa2xXHbHfcpcjZtx1Z19OVRLKCT+XGgwGn2+z
AMnoGRh6Ot7+MmS41TS3fuBDJqaFqApegH8GTN+zuARrNDW5yjpIegvLMqLlAcZ3GUQvu2sOQDmM
lULQGlZ4YYBWFkZv4oH9DldYb6SbopZ9dAqvtnEBXK2c0G1/P/V3/ei/Q/4keucKw0RWDTWkns6s
66aVmzdFlGn6O3YoeFNRdRJ59uAQkfMSNCHtWlw7h5RH3NQqNQ+eicGzaS1p3M57IGp49mUmqa4l
sVBktYJCoo0+auEzcsB5wwH8KhPGefYWKdhhwtsXeZgojByOoE4mTRh34kXH2yXQ2vJh3ZjbuvH7
J0Syvfh60coJ2mOZtxVtDCWBsMv3rIiD+L6j6DD+YFeltSBqccpif33zjK0fxAsjELFLXz2Jws59
oJVIKN+mT7gf7dURlrHTzMp9Eax9xMZ2feW4N9c8DWsP0sqK+63cepOmCORmnTTgW7HGGXTWwcPD
g+HFO4r8ySuY/ze5i6SFco/IgZjZJlX+fvmwsRsQuY/L0+nf8mA3ENeFrwEcnyouyMB8TJni9BzD
bFYV1aJwcqEzvUBtlMYdd8n0ZJCnFhtVDaYfPQ/bywM/v59CNhJ/RITknLMlbCFSz1HArO2TRHnh
FQiqfppUCg4MyWHxDjcynFR40xK6MmHjdm8R46QVlQdwo/adYS1r3JV1DujRH43luXI0se1MzKiz
Bt0z0g0CoYDGlquJ28+RzREKhTC9J02/SHoivuUqysCAE9IH0fdcSKxtqFJmAOVR+oHrJidc3nRa
wcYZYSsOaydFZYds+mEq5OOxoSYBk78ELESggCqh32y+YQ78BSilWuYtFD7mAUftpGbhQYn9olbX
2TXAP4b7bBrEbgpgsoqViRbmYyojiNmLs1HjH5v+nrxKxn69P4FFWWt8jIAcfkNZDZqsT6Nh1UYX
QHY2MVR52afroMwMroOZ0Y++yBuDikFTzxaSGnYkxFOsUxe9+x0bPCRhOolOs02KMR31PWQ36ugx
ylr5AwJiT+T9kpnh0gN7QgVG4B1mTGJjIgfSozbLyrulGUz1nemtiTtrozCqBvno5s8ppwL8VwbJ
Ai2JClc97eejFWDGBhi5haZYYLIHsJmpsEXmqupFa+gKjhb2tt146vZLkYu6nb6MbKwcZvCy0ZUU
bKKq8txSV/RJp2bAPeh5USTpriYzBHX830L17zwndeqJc+TBcD0JB1J35T8aZ657KieWO+6QqWcL
jADYRoILNWqsyDI2mEtzdYTn7p4gU/MgoPXxUXc0aDG7DnfAqq4EHbejvjwci/kNUREnAJLXO+G9
3OTF+RtxY6XAGV5XR/BTvPOQ8gzflWV6UFjwhbMxWUrR25YXryiMWfxNMj0Mt6zOQjVv1+zFpTab
6IPRyouna6wrdqsHTryyCMdtZGyQOn+K6oEjMEkYYFdL4hmUt8Ndbwpkyi4je8PWP0KhFek8ClFf
/g+2fO6/Od+dG8M5fxFUZNWvL5hq3OT7axwN5qDBtRV7wageY0cwgW06+qnZJKEa6G+jkpgJAR0N
NfOxhOdK/hpTTgs/o+ypWHUW2ZVa8wrtsjbuvzUlbXB/Za0+Z/6bw1pfq2ktKxtKrrO2l1e+D27X
hsNu9lqflhZq6GS9lsgO1PTzFPWbORVKwicT4ImxzmOxfP1c41qtNKiHIMkFChiiGQkGDziZBZk7
RA/YUsPR3vxHTAAyhlsZIT8YhODVHi1bwJQSFhZRbO2o0zkYiSM/bCUMhj6FRisPbcnHjFFc0s+m
AL0BU8rG+0C4v1ioGyCu/fxyAL5PcEXd5tshAR06d2rYl/ypmG3TrjLCsVV8EyXtDT/xo+qfQzI9
iVgN1EXEnYcAJUY6mRJ+qbzod6O3RdBVcRNO6LIFAR1OIJVUmS5zO0JBwBDiSdR2rDYkYIE2blMA
U6/SEs2L+ekz5xMAEnrLHogAlgLRl5qWjC+48jyP9sKIzxi50RV/TBR7TcKdExE1y8EuadzWjoBI
cjW10Ogy2iwtRgPMy3dYbZSVmjoQ3hrEUCbC79AcF9/urSF253ttZLtWDhm9heh9FgZDY5G9J6M3
McK6CzDQ/KBHBO47MFjkNkq8RMMo8gvDjMLs9hoo4a7+2AvuovlZ905E+naqAw9HZlTXNiJElC3z
rbKgVEZ62Z3ysqGqWE1DSBQGvNrb9MqnjLNT+JUOjyKvTcdf/lHj/2vdz37pDUlkSswoNfX+h0lo
coTq+UrWOeYaKLXRncJo0UZn/SQ1McV4Kxk8O/RP4ODjqEyXPRfNQx4Pn/pVZInameG7we4uQHwq
Hut5NqQjbFEvg6ua17Yva0tZOOQAEYM56rNWvpjjHIBRox9NI3Nn3HrrY82M5Hq3XKkYgqTn/2e+
eePcrpDXLFumMD87fyUQi2JftKmL2QDCzlt1JcU2igAfvoEtuMjLRU7bmlVYb9IbB3oeEDU31uDX
CaGNH9g7e3xVr8iPqheVOG5Xj9Zx4CiFLpTM3Q2y8ZhWH8cUxjXg4Z0CI0p4Mjy6uEqHyuAbAm8v
R8102N5q9mzKwyVJtu+ARGPENj31gZ4LpGGZFzWDeyz/wdlZ2lLiTqiOKpvsgMGVriohRY7CQyav
sgZJyjF5U/GnkKa8O6sCBj0Io/2GSrxdvAAfP7Tt5EJ2OtpXHSg6C+14dW8UXxv5qdwCOEIWTcLb
S5YHVlulym9b/j7CqZiPpD2RiBVxh2CN8+Uyyiap0DAEKLmBM66WU32d0VruDsUrVRdcV+2NUBi6
JukzvocJHbeICWE7+NLrqYTOqvglYvSmQnfq4BE8EKZuRIdu0SCplb2AWb5qmE31IhpF1ynVMPLB
fltAfvKlg5ZKuhW65pL2miY3Jr4qEGB+3p51SKQEhZZb4v0w0x9y5lBH6sfrkIOkFB/6LI49SkeU
wFGdl7QGppSeWAWNEO0haAhtK4WKV9Ho6nDqlo8uANLROhobiahmmDtHGPtEuwyHFu5Rd5Pku7Rc
WR2leyVXiZCe++ZX9+CF2WWbNYbzq8uX1QgCicROk9T5iGeb3TshmQb2Ztnf7ob2nip7muGN3u+V
b3MJ7hxnlfxlR+rrEICQBAkPWVYZ79gU8mKIMtIY5V1uapTDnGnTJyvLstl4P2+mkTtRFeRySnIC
OUdHqWOPKQaycZCJCdjId1nUBbUVg86LpU+ouccGMc38wpUVoZovQZ4kPUgXq32KbcHte+F3oMU6
e58OoYqH0wnhDfCqWb99eUHpB3oUxxdczkO6T9csy4fd02whjD0k/gocQesuW4Nweis647sEdffA
S9geRrIc4pgYXj7+RqwtCIimki51U6w8ew8j0wB2ARKXtZCAgZqitjH90asQHkmkzK8hqluT/DTW
KH8VMQkAqne4/DvloBPfi6CGaj6JmwtD9nPs1vyqhX5ivX6L3e1xdV/iXCTIzZmsHV624ND6+lYL
DLY+l4IeGFdJJRxHHy5drp1yUm1Dbvnh7slOkwn8GgT43EOWSleGLuveabNgO1/VlO8OOLM3mbUM
YUtmGZu9az0p+pEy1fbOKBAB7VwZY+URqrln1u53s0pqFXvWM52WMvJ7u20wIqSSr7fNIL4PtGxc
YocqssIh1mIs7F49k4GKRXi/0THNJNLM0iMkUpXRwjAyEMUJ8P5qWvQfz52+UHKV9ZNYmkPtN7Cs
u1y45oqK7FVNfDjHbulCxo+/2CkzGON68UYkYiHQI/DRJSwZFPpFlaKcgd0xiUwGTK5RXYTNrbV9
Kct0DkDwwur2FejCoaRcVtmK5VSRt/WNwV2gZ54dilg9i4a4phZ3MCH8XEbWmxvAXrVrYptccl2j
Lpz2x3dfXqNSJK9yCZpvYWtgLe32X8xKWXo9LYU3QPwtbIz+aaPOJsUOqGCbUznOmeCITJ2wzPv+
dMpwnoIt0GI3JG5A5+dz+9rpD6d3jp6yI29d3O8BQi88cuz0HCzd0UA11LYbARxIFQfqYVcqXF84
a+McfjMwv31AC4NQkfEw3jMc+cn54qgP7h6xVAuM/5U96qLcLw5eHX5G0UGMYT7AL3UyNQbcRfn3
i+KJ8A0HX2qroprdiug2hXTwQlEwIqAEbqDhxDC4WKGwAKmezxqvM/jg6UzQk0SqmTFC/qdC4g5n
BwPFu0daDdovLbdYmi7cRd47sBDjHT2KgSHCXnAvYpE3dFuoi88dJ2jnOSV2ADMEFZS+830lOdbR
2JLgq5R8SfllEQ6wkNiGqe0z6wyA731bK4AyfhqghHCppZMXCkgNP+dLpb1rzrXHJo/J8TTIxuBF
pkuVSpYf709v97o6U4lOTz7QUOLP1XX0G2Dz2iuxPPnj0vJv0dLNz6J9AfjbrX9i/NLtjwLSR53K
fThhVOvwn/EvhY6ImamUgn+zrGoiFgiX7lme/QeDyHOuIJbtbzjCvrAq3jYwznTFglGN7lOextMb
rKuAgjaooyTGOC6rpBInUX+MkgA1yqKL8chcnfIW90sHaLvKLoq42X3ifhpd0SCLmJBZqscDY0Gd
4oe2309wydV8FEZPgMzX6aAa5/9vc7NYjM4PNhN+fIOWknZHkBTRODKrGWD5hLrXz+rGe7HctitW
7Nq37F271DZofZcUqs1REspEvKPYR/oUg5lVqgEKayAwQqoJkiDWq6qTTFGFiNlnEHS8Fa1ODDm1
n5UuzWyBwKuU2qK7//hGuW/IU+/pKZFJJKhBa4V79Nt9g+vFPq6Ao+XIuhLQxcLO/tLhNDpTD7Tt
4iF1PNpi46OEZjfC9hTNwFj+63dfS1S94RoKPkI/13HCpHYAHvYmz1YT0CqdYyv6RtflokUP1Z2U
f8HMiXSocyNahFT9m6aDiIQOeCvh6RvO/eF7chmw+YQw/z0ZqWD9WjKIeC64/Hzp88ygvjK/w4Hs
iSCTLonaSeUSLGzeQwUpH2iZhPiCGInMwseaY2yPpF4AEVLPGxUML/p/0R8Mq3fMa+S+7dGHKrYx
bocDzprBuYqDbPG8fSNEbxmg7xU1QjzXn12/onXOs58cBIDnGcQfl155tR/E7vR3vUqYGeL+4YIP
20GdkSKx7//UdcNSGaA7EYoSuewh+0UwJJLtfoOWVugZtTUGqpwuAvFqCn4Y4KtZAjxDDm4oeAWi
pAwn2BOz6zL9nUu6QBzeXUL5IbCDINrKip5AgpbdXVOi8RAsq5WrSH0VnwiL7W6y3Igz3blNflMZ
gK7eWtWlmSIlkJ1D9vsiRdbc4j7n54YznrN/14zvvC4ngt6mhfbVytLYUVZS3qXh/LLQWkgH44hj
lrkWHQZR4KJcsI9nWBqo1LqFHItZ75bmzRYYZ/hzB2afesl0l6nWVew8F6ChEki3lOrTKHGuoLA2
lLMiBXmuyfMW4PCPWTjx0yMc8nPToLuoSxS3RtqmjVdS1FcK/uVapSNK/gbuu7jI9PO9kvLhNS42
mOdyrmm1nMIh+aHlT/1qQlVQAxq3HxfU10fX/c1YeHC7OH5uAIRzpg1Y/L2vph+FmMxyiokyhMQP
xX97Rq71ujgSeqCK0ydWDv+DBN5kuv0HCyZK1ckn8KqFuicO8bREwbiSJpd1oz03iG9OUK9vBHJq
HgJ9x7zOtV1gmcmCqemXH5fXtOiAbTRjvp724g2qhEvqFzctyP22gcCjs2xRBjEsnc7Tfu4LM5Ph
4rz1qnfHsPI7FeUL6UVrBvvwTTaJ/YJwUBmisNGtHwnOm4me4TJr1OLZjLKOjgDyNW+aQWxJlqn6
xRIKztgFWq4RGR/d2hLse5v8cxPLdlA27i70TT9iaiUIq3y9ToGxsZKq+y5DMBRyXyDMWFWd63Qj
kIh6NFGgPpVimZnPO6Mm9/FfTS7jFmXyNZp4FT+6MJElCof3S8GHvuYgZryzIak7PtZ3bwNEqJlz
uUwBjPiOgnnWmJRMMVmjSaK+abSDC+2XX2wniNiGuHJp/wVaq7WbfgQ2amtJM9mU5SS99jp8u9E3
S73lHH0onCY9zOsNSBrd7ih0R7zXJ4flPdsimGbYVlMX4rzkDddnyiBXfq6Jb3vsUPxohTuED5Su
CNZoLhGtxMvs7xzVo5nR6eVKWL/qP4ysQc/L6akdMjPDC/WBvGNjyUXdV8c8hOdfKhI6dj8/wZtN
FP5nbbuPfIf/DAk0knj5RwUsO3+eep53mjT1Sb3FcUBNp20ZOskaPED86KOoBgHQHUX+LsgYHhpb
cLbIaJKGQ0fSpsHAbFjtTe0ZAAHAhyrNMoUUsQeYPe8sdD8mCc22DGCfq9PEgdevrV+JN+moluEG
FkkDFmi2mdY9+e/aft28/Syypxlw8aybXnN4vmeme1+SNtiyDW8menXp1YCEOX1uPZqFnqYVrx69
/L7ps3Sg6KN3kAAevJulw6aghB9+/VjP5yUaJOXE6YAJ7JJ6oq0twnuvcUehLThCHFVdSfnstkD5
HWjUEniH1Mz6iaC1mW/IJZji4gWuXrvXUl4dF1nd5I/Fg1thWkpltXnZOyBOAmRAgcmRTcarD7/8
4HIyTx773QWpyjNrzYFJaQmwEWmQbcHFVV60CT++0h/I0apPTJWDKFbYlFlxxhTcwlmC1wUkU0b9
Ul26u3vGqt91/Ttx8ZJ5dYjE80xJvMaALFKwnbpKNPBmzep6cZrwNW6hlHvlSgrvKP85QT8btK8s
N7Ihy5F76B/x/sOz4HcEMTon8xBeeQXNvhsVyaHLsRk+KqLu8h1/IRiXIr/g4fC+3x3KbaRtXxhX
5ajSkspe9Am9hnCx8wwIvMiZfbDK4ph3siiVz7D5uB6aG8FNmpqZrYICtIcf9v0pD6/QXh5O8BgA
NESIcyu8JrJcD6RXe05XR1ersB2RTFxHYhE/87mxrq4S3rvOZxfia9t8XZkeg0Ez5143H8E+N0PI
3VshRWJDNyOekbdIqOzDMwvCtV14tdisuyW4VIIj6jYruxPe5FOPsD6npkW+KAn43Khmhy/C95Bl
mFSw4vUBNUn73V3rmCIx3DtAiuVNd5kc0CdqTrM1bMzeXNAoVwWK4zELsVn+05OvTf/fnzn2OrwI
pakTeYZ4lwDTgQYMeG1gdZT25NHypPqaGgPWExf+Ld8CkYsNu5IBOrTgGmC9lUTz2DhAbbSvmXb1
WgDPnfFuovISzCUYEKykrZy7cQkvgghsjZy0Z9utVSgJME4IC/t0t/OrtZpA5v76M3HPV6nLNAOb
7a47HRtV0Eid8vhVl4Okf7K0BZCKNgiy0Ktt3WILP20SPTXc1ms9+g/VrE60sRsFObxx1mAxVIp4
LImgXkvReSD+ztJ1mdxDIeHmt87AWbnE6KTUnUG0KsyQGt8HD38OZzO3PzToVhj+U07KTOSISlej
cPnrm7P1P4mct5hRMGX/4ihT62m4Hf7LqQdHSvC7jfjIi057HQUsuiHuQc9nVBk6/fzihwO9n5F8
LxK2iCOkqiGw5kTtHz6EIqFF/ekLyY4mBS1k4JXTTccpgkoIx6myyEknWf5nKCGV7UMaKrAVvm5U
X+AgllsR51QHHFyJPmUapggvkXKjlNl3MVvkoSMrFFB6vSUIRPJj6itof5yP6RAgme67t6fsAtTl
wGbYdDTbJFfKOQOo0uYt2dd7lUS0ot2Y9XbkWhHFpZpjuMF8PYBSyw1WbwvgyfWHyofipEtw8oay
5LNN/BtvmEwb+ZVp4aS3MlkpX3KVI/ujHYgaK9eMVO1hOjx5IRRz7fqdZawBZpSlRBq8XAma6O3X
fJIQlryoKElJ3SEHUoVmqTbfz3efpOpmXca6+8c5vL1sy3OxArRjaIFTUT6ypRLX21vQiPt0tbWI
Um6nbDYzhQjHt+Y8g6WYSxDkHQReO283vFvsHtMtgd7A8+ckct9EiLIwdwCj4orFIN3gnWFCBOWT
sP8ACNMx+tkkgG7srgKfLdXF3sAI+ZZ21YyAxnoAS7c6Mb25x/4gYJtPuuQ7QIEJCLmJg2+ejUi/
7w95tVKvtZ8TPa8dlPZcgmZKxVhpm8RMri0g701A90p4xEBfjYnsK8YMcP5RVV6T586ZiBN1+XKd
TryxwKoCgE0ZYvvFbWJbMc6EFuK/+L85j2iwzMM5yrXWUGi4kLU96VCTpg8SPTPxuRttJnk7Osy/
HGqe3Fav5TBTtJl+KTKXvQsaaqLoFLj8yycwVC4EpVZiD9Wl3Hptg87BC9wga/v3V8+ym/Hayo1W
TqhWsfMls3PRSrNIcEzhayVCp16ysh5bfMheVY3bJCzPubWqzxNFMpVGm5tMy99LgX7461ed3IJl
bPdaZ1Lexw5w2oCdOP3avmIAIlpXrjNmIbR9yPovbY7UFI9wMkDc0LSSd5taNhskn5J3ZsScFhc0
p3VlsQezJRcGJviuS8ULmdH7Y3Zs+EUr82fX16I44MIe++FEUphK0gEEL8LeH03fW9Tj2arexl+K
THw4tFwRwKTLnaj6vpmrmoZsw8HVIfdkJ9ejNY2L6rP5VpsLi09E+ue9gm6KGkEFskPE7aIiV1fU
tw/rkzRFyxGijoXrK8Q+51HqP6kpLp4x5NCz+Au7dOpw5cazDBkLoF+lvYtz68Tak+2guWDRpvG3
X0UBHW8XjRfyX55PcWDJn6XUddfSl9qeawphZrZFNGQAX453kq/pVYKUGDDIK3ie8801i342rOIg
wYzxH2mgJgR/gm12k3a9BAJdKVIJ4/0v7ZJBxHYxynrCLse56vDB6R0X5vhMEoWZq7JgMAnhsTJJ
/63NKA/8nGxw+pDmw6tt+ra/eqgpZLmGIQCwUJztotB9EHi2+/Qlf6myr36MnFSYyehjzaX5bS0Q
fIi7pqW/Zvm3Vx7sWLX/112wSwdu4I7N+qLeJsh916JXmGBAH/uWYOuHACRNs8w0p89iLnXbUEJ8
l/Dlqs2Y+vUXyrGmu4aEzZXjBkl2dZCv3nO9fpMRAV/pybnpX2LjqsMmNR5kXu/LfagHhlM1g+vE
DFer7dWS8C6V3wqxNF0YiFH6Iton2adalDiOfpQ2p1PeHLtdaW4B2HATladfNc5zuVRy6q5gsTTI
OQo/y29gWzZuEU+VmBFy97jfTTlh8x8QET2IPw88wATfBcSu/jA+QumjwY/oKo2FSPCvHvwqdh7p
8sKiQMEKODbhRgu7RGtzj41V7ypy74oiQWQKdgf9i5J+vslDuURHK6GcA+3CCtao7OlgNBzOEdBS
QqG3UfoQ+iEqTjc5819715GSoLRAldfCHyjI8l7Sq3SFVbAmVMS7mM1qBN3RbO8E/66scyTbiRaN
YQu25z9DNobsBBnapCi4TDDf2POB3TDMjMqyw1NcRzlnQqxL4R2mnwiDaAk66bGgGrb2s9iHdisj
HjYunWBCzXfpqhnRMn4SxOht1Q5x2jFo2gva6Qd6DQNS0Gj5kU9ictt1pdYgmEUwkvR9lwqPnkG5
Lw7lZDnCYhHj+JcEa4VKA2katgk3a/pdfzCYkjNhDxWhvQ283AWy3jk0c4ACUstylh90cEgb6BPz
ckEulMH7NmfTxaTHA1B574AVITpoMvtR13QshNkEJ6Li20slUyu6dHErtzfIH+MKCnibil5OT1pA
OcwJerH1GlRUzOfe457q0ZK/LWHhdUo95XpIj/sUqecsJIhrVaDp6LyuySfXSuAsWdb3/01EAv1F
BLrOiIK9qqLcH8/R0bTMDVAD04YVwvEv0wQttL7Kg9njx2QlTuKUAF99NNRKK1/yfDF27q+oo+XW
HMtz9Rn7gu9ogv4z5m1p50PGUCNKMLyaXiJrh/kMCECpHuwMqzvx2NUqdhHhDR9+IaZfKM2kCqnG
w2YKXKU+FjDEzhORU48pY1BMUeN1MKPJ0i2fpIRHM0pWK8IuaR7Ta+AwEst2oUSyH+6kh88C0TlR
kdGAPJV0NyfVMpMYYw5BNUo/Q9/56fHJ8fP3i3QVFDzPzx6QscxX45feO5PPVgty+hpzk1o7OKJa
ZVkxZDUMR2dRMTppGtfr8tWqazYT2mhW46LJOz06RJgr1a2pdu6N3Owsez3KbCt+f1POMqmWx5LX
nlVF/RP/TP/2zjUT02W8aoLu363ZASiA5L4uliZlYyd2z1pmYvOQj0LzVgD9DcGD3Izo+BxRzPSt
pHEy4S9q9JB9zoMenUuXFb6qz+DVKxlQluPHndpg/yJCVeFpkM/rGrnh2rZ7D7p0hRtNmBItB64m
Wnm+p1hVtQB6sa2wSfxKb1XWVbjf5o7nN8w3FDRpav9J0K/pVHvDbCmwMFH5aC4e+5/iVVqH2QQs
PhfnrIRmnh6Ci2K5L0phdDUCW4I7VY9W6Lkjtfhe13uzEjRxoifEt16SYT4Lg10/LWZwKvafmFvO
MoFaQLwVhFWnlKWZ5ZOhve0LUV57WT13228qy0CL2gEEkDmeVRgoqNvYmySnE/zXTdUoDXERp2kr
jUa8fWhAolp7kDrSVNu6RpPFgzg4qVU9wzDTXlUlqbjDf0na/gT7YygyN35hBifPwfyuKlLURXT3
/1U4IbUt2FjWd9e/Poq5BJfnC3gg04k83m17g6trmShmdOSgKJwTVkKEBvr9ST1Fg+Y/KB6Y6sOV
Z7aCkOMZhYK3+siaSceRanijDjsC/6gUT33G+SUEz9V8X4APNTJBeTkN9zbLTJBRt3NM+6aSs9NY
9KDu07XHKKAtLQfIJ3WD2a3z9szGkTsROH+dLKSzJHHdLFGycdNWsnIhFK2XC2J6K+/MZ+wCj02m
WZfMVMulKvL0/voFQjhggXPxRzJMUCOS/2Yq4hDD0/9pgC8ahg/ByLiFlmyga7etciopUhSaO3/S
u5edEu3HW9MeIdpTwZunEwyA8aSPNzTQFC0lLexXskbHYdQcwfV1Brz4POXUIhDiIpTKYdeQorKO
l1cX14VWSnrFhJ2iNMS45AYAJ0ZbfJrpGnYCL+ktwg20sO29jmaAHm7t74VzLc1iDbWg+DvepNXt
lvCKRp5Bj8J7I/hGxw/5Z3/XLbGAeblKDg5aX/hMC/gSpzAztlaR7txkasOeAvvqnvOyMQQcuyhZ
ljf5HJvqEP74Y/YJWa4J/x4EQbzrH7HHQZBOe94wFP5AKGYZVW9DiMl/Olva6SlcwjvmRS6NTKLf
MJeB3ctTtnVx6YXNZrPQqHey4yqLDhlpVpLPPP/e6e7jfWuyixugmNCc8tn6AV2eTGQkdUs60Ifz
42SKxeFPEkkmUTJFrRdUARa9uYB9g29NVthLVzED6EWuQ/DSJROcoyJ1PYGZAgF0BDkM43Ij1yOk
PXiD6Tw6KbLYqqBFbzn7bRwkBDRlLYrdhcySDFdI9ln93+99O3cWd+ZjPlKL3wj0sxqauWV1GAe9
sgRNx5imJxfotneVN5IZzzAWbIHLdt+kW+db1XyMivMdS7e2fP5o/uk7zZTxCtNDQW64CwnMG8Ej
oc4FIcLbZDd1HLD+SPg/47UuDXlR97VGKyXizsT5f0y/w8lbS5leaEBhLvYMWEPtbTW3Z5KZ5lGn
Ta0Y5Xqpz/hcjnft+yT/FDw8TqB3D47w9s3O0sxedOhmuCPF5WDjGTCq/4fO0ZywLfl0ga39PY/R
DeNW4vuvHzGHWjGFJdq79hkz5IjZ5EJeOhSR9cZq0c/Avkdz1Bhwhxs9EJ6YFzxcsr8Q8pNNX2vV
SnUhoQjj68vsKqyTIA6z5/KEkRjVpCMPUSbjMv4ZecYy/1qNXYNV/Evu7SWZ8JLjzMbSzbNjiWBS
QSxi7Lko3ZvjV6yhsbbKVOFh+N5JRL8YKcMp5vZ7anY6dFjRL1SJiY1aVQxgcGbJ6K2eyIjb8Du8
p/bwFryNwh1OZgNjRYwHlrUm25aVG6VoZ4eHwgffQSxDOq5mQnQDFUh5SBYa7IwttfY5xC26faoO
+2LKOO9B6XTKfAjEGAZ9QDVQD6XIosYqlKWNd5jPsAfUWp1VkOd7670kZuqZavxI3O8tB0YmsZ8i
ivfbB3rMLFyX8c0zAsDQWViplj8DXRXehJ4nFgeukOclngRcGWfuag7cmMu2E8nGql+2hDf6j5s0
lVF1WxbTQRaP5//yQBVEaXtJauHcMLAxe1XHDilf25q9RVkiQyZBINlP3B3yMb7eK2RxTUgEQd/E
vhhEqymlb+DGDU4nk8aXlWCSn2Qe6BQki0gvjkS13dgS1r1y/YhwW7ViWjfqPX/BdFnWp+e/2CiC
vDwmfoYHRI98HLRyDV+SE67r4kUx87/uUlz1lCUqxyjGNUcR5PvNukeJmTetkuOITihiy5AWERRT
56usnhq4W8II5MzlaEaiwTvwm4uXfD5xLgIiBEf9s+moeE/8C+MAx/CFwjGK99aoWWtVBI6KI0hN
JN8hdaG+3bWk/hPHzaWGcUzwdZYPjNmaJ3mHANhPx7YEObzhhrfbz8Gd3g7nO0K/30VRufRlnRo1
JrPvldsA1aXxWsNB9Y0SV8Sd5R5OrC/L1dimuVo3BsRyIusjNRJsS/2qghtVDWvwnT6wkFbvqEQf
UMSq1NYvFqWpMxVw4Dv/f26Hh2Qr5GCC5nhIdR80WiOVgtHz9Mg9jG4l+mn6B7kOw8fsnH8JfmHY
B37kb2lMA220IasR5dEMqal6N46QDiu1++rTLSc/fxo2M5/Aanu3sG3qHEMD35GxxVKwTrPRnqfl
0kavV1YUrHW8QBXfVmVEud3DYyzLfC0aGo0pfbLwVjqs2AZsnjhIztaMhUHCrhPLb/NUiWiLlpAb
8RCg16+as7zNK3N62T7gUk4sRCtOHatsKtl9YLhi/Qxl1BSuKIT9ZvR2/SarfJbUzy6HhioeFRJE
PxvX/yrjwcEvvpepJGaA9mKLUFOd98M/FZG7BTcI5F/1Dzeas0oFfxMMkzJ/grMF5/GEpOighlpJ
GfocT8lsIfBj8V5Je8iIT4fHhOy6GCgXi372v09OAIOTQoxV03kwx+cwX9s6PVK951LU8uBL8hBi
DtCEwcl5yyrxIQOr+EXtW4TIA9dOg1mQdhcQdijGIjTOxcxYa8q9Jyw67Yb6/m0RwOFqe9ysOeG5
HZDwmLH+8THznkmrsYOvZh0wt7jdV6VtCtmmdBHDTtTkmyCylQ9PC1/YNjugAvrxcI0+ztbf/XHh
K6xSb4Lt+WJdWhGIR7Gukpw3CHJ2cfU5OdHIjhJdkiUkrmlXLvxkfZCfZ9LrfTepXyb75Ef5AIaD
SXtVpLxGgSAxErVLuqOprSyAWNIU84S6R/rBrqwQK1q8dMRKGYSSYHis99YjKCEsqGIaWtrqr1KD
wv9iwdQDDcv8acDgXChmhpXwnIYPi95HjXAAwW0GQWrf9EKqKZsIgUq966Ka4uHQzTALdiXwyimC
C0CfPV3y8obK6dot6VfTfk04iZ91xni/q1dadl5ari+lvoPKyALt6SfKGbDDQvTkzduQJNu0J+dJ
sMyvTN0waqBTCsjeRjaA0DTKbxWcf/B1POo3/eYnUanKsl3HdcC5mm8pBY442r+dfF70ZIXMm+D/
XsQb28olYIcjGq9lMk8J7mE2D69Yy6yndYUxwcnZpirImhS41nDej3doA8rPrsCKJ6t6xM6pYLFG
voSv3xua2+XGoeFGKdH8DvxQ9lpqX8rPVBg/RbEAEs+kPCCJ5Ex4uJhBIGwtdimB0yKGZwHlcyah
FxhyDIEMlcsNXtPDVzQN7RMdp+fwKDZs4FxaIwJyR58SeS5wEoYXuVM5JSJ0D8prTjzE4vCvrDMd
tCliMtztjFLSGprVvzE42TWfA2uHAU8TAUiYVByJR8+kfGJFDq0nqOSlhUt4VubmI2kqo/NC+UYg
PvrDAVTIbifZyXZUmccQErYbtUQOuQfjhNsTtq5quiuj6pQI+uTnpUKD108VkYWzsVN1ZK/jx1yU
U+le2DxqqX48Tbe2U9XIrZw6qetMJPoGdukKtNSaGNTskRw23IhYlBcqgb3BovJKJ8ar94XhfsSm
26Hxtml9AwTuK3AhNo0A/n47jCZxFNUmkOGAr7qxkZUO227tnbOb3s0bELUtuIimojhCv+oKBcJu
tI/27CRUPvqKgQ+rEZV7a8iRdNQA/qiMMCGNDs1SVEltUHUChgMdbygEGSAczDO8fBHwpcyI7wWX
0HfvKWHXHgzRQMOebNR+EKS4xhVvs1+6BA9AN1R9qurQSw2GqhZZZlAYkHaeuhrx2DF+l2pfKwSa
gVaia6tV/eFI+BONtcpd/7mtpRJoDiQEie97nDPWqS/paHx7TORE/QBoyb9kp+6ZUVQ26bRjqC58
+Ptn0BTXEwDGqpktCLbJrgTINXg0KWiKjRWWVG60mUb5zUi9//vXhHhD1CmeFVjS7UEay2IYfNKr
bzrlVIyeuwQRxN0IOqV2AqWAIetNCB+GuiAQ0G2mM0FkqeTYWwFlk4Afh8mCcQSz027lWoyVp7dR
LFzWm3IqtEGyavnNnCXfTSDrcncQ1GhICCeu2JnaLaXK1l5b8qoy7zWMy/5WE2Y9QP5maZtIeDEZ
ocWeSyB5n7FD//koiKvtw3b8xuqm2HhXAVZ7aPpLiT7XfoEVRD4AdBoXPxgmVZAIjar2ZuB4e1FW
0nqPmuRSlLRcqHX8eOKmD1ia4YrYak+lvDMn7iDgI02y41TthnOkWVNNKd4IMZIKvJZgGoGfl+Ae
C+bIMRhc5rbvajBHxDpCLaenQLCBKrgbPo0CmjzoZGRcBXJ9Q0hMEJIfYZomdiw6v2oVE4F3YQkc
t9jjeIzQIhUBzcIpiZ2fJcrby0BlpUogNf7xYq7y6zAR0kc9Hj9IyCwvkeo9Tf5TwXVvYGuik/Eo
RrO+sV4pNXZeJCiJphU2ArXQ6/enjHuABZnju3kUDts82lHfmUncFhSzf0VnFuCYREjxK/rLyLYQ
yID74Yhh0lz/n/IYnVa7jZSoU83uYafFyBRYKxrSRHrgLp0BuLmoQw0MnLZMtuxW0VpdcBVv16h5
dp/1lKrtxkDoaUBZbTaS0rUnFh/8mMz5v/ojlFS/09KR5sZAf7Po1v8z5ZEYCyTildZW94KOMB0d
7belEDIJjodsjJbji7jor6dRDswED/WKEDpEvbsLzRT15PnZrVckKD2uYkeK1bxoMYOljbBWaQXh
kk2C8IgATc3y5qFc5u8uAq8RWTpSaFaJUr3SlLVsrRiLSoCTbP/WA5zUj2a6i7+WtlEyJ1b4z4m+
E9GixhluSO4dls5TlzJm+yq5eTVq8+UKz1ucIBRW9LDrZL2Y8PTZ+AT5g1c9sI24jTi7nOzN3ceD
X07ei/hAxr2IF641RB+FJodWseooFd/o/ygUrSenrY72vDiVRwlz9AdWsMfUnK6S6hlGgDCbAFuq
Lz0ZwLnAS/6KSGwDVpZSIdL26gG8k7IBQ/pSNONM+VklLcMpRdXIQePzm7PPJfUEpFo02hrh7slZ
TiUtHmUUUg6vQDtLd6AYPOk8n6KQvhNKXV10ALyoiX0RyRi8CAsww5/oKhLfqOuD82bJ/U8T6xhJ
bwqAT9VSbgNtPWxo17P7QDCuJqRqAlq/hMB50q/h04gV0XBoByAB6r3PteN2GfAMLB7xNsmsTrQS
QwHbkBPB7oVCX5NrL3FHlJC3tNilAs2C7zYJhdnl1gn4VjXE9BiDvlQ+IfWt8isqW/us4hrcTHoa
jbfdRBzcWCXAi3U8DvGAeaRXK6N0sRaJqBqwQHVZjXyjo8KDicVqDW08VOmO0YKqDxwPdkehgol4
eyuBfbjO14kw1J1sv/z/vM/s+cw4hKJ6gw2OA9YDZI/sCnlZK2daf2kNyA3OVPERLfjDQFs+uENC
xlAmQm6QUZdgjq62rwNyF0Y1dHNx8Ie+TJwunTqucknMBua46HxxNtUqKOlZhRU19HlNJGQdx4X+
//tStQKnxybR7h2Q2tn0bWhs0r2ubBVKe7PSCCP/KCEN6/Iqkb8gwvbSzz6ZJ4N4exWXcIyN0U19
dIy2tpHWm/MUJ532nHLGW/723WHnWdT+Oc1AxMCW+Vl+A36AY2sL2ydB1hMiTerepvq110qkJ63R
rSJLt/q5Peg3e4+xm6Y4mUcT9ZWenLPfVFiJrRQzHiUjp+lCGxG4kMYMjGCuZnE/EbPMUBdOucXE
q4TxtbLIOu8QuOdT+W4j7AzB5sKD0BAt0J/bBCEqju8+WlW8cBJwYHPfcurBGmSpy0Aa5dp8IT4/
JWmFmR8mVMBIY+e6GKMTc1AK6N9lpn17Ep+NtsWIRnFuH0YWOkIUVGbLF1AQSqKTbFOlIVdHiIRI
e8rGcFobNHxEWTen+inDcBNM9O7BEwIAY9TGTr6uNbdzrRmHsoZyhaV6tvGCE+xuAQBoLkJeHjS7
qZg9d4Benetk6BYGFvIBxJcVsBK9f7Ko++Pmqc0GBGh+NrsZEccZj/qu9tRpN8IZ9P2yKdf9lW3O
wcN2dr2rz7TK5qcJYj2sjEhcPPOQ3jCTjZe9gmoYX+R4CGuH6wJ9RJxWg7wvvFpgPFzUUC4E9p8m
CMdPB6tqZokYdUOCMdf+9K9KOPDvB49wWB++KHE2+Qpl/Vb3zyq2OAihmepFAd1qMAMmooAbjS3y
9E8EaIfUE0A5Dr25TEi4+IubRqQH/TWRllLV+nbpIU4iZXz4M5n82nmxiO0aROvVIVujAq+nFyB0
TbBdaJqWtDvcTvbokuU8BT7Tt7+DoIK5kCqoVAlch6+UW3bg2MQBjcRgIoE6rTAvguTb2DLI7/dh
JlNzRt8wTpSAHsBTnnaI2iLCAp+Pu8gahWZe2YO9ztQxh3UX08cKuInOGqdTwFl0o7HMMJzo2gJr
tWJrPa83ho7NTDKUIX0n0A8Jm3Ma7qcUknzvWWW/ek2CjFNzhD3sp+y4VaQuRX24YaUKSINgmQ6p
4+ujFA8uWh2w6A/Tuj9G+dagI3ue18CBT2yVNmAiDrSjPv5Y0fBvyA5Xq5uDSyqG3V4ytyA6BHtZ
/YAQBFLxi4y3QV7syw4Xb1SsK2ZIONm2g9V61X4uDppgmbyqqZnohNZj9K1s8UR7LuJghKSECD33
tOS2hDevuVA8wi8pjj6C1GiiEykEFcXr/QWQirV04MBK89sDUxDishM46T4wzZDFi2Y8PHQGAjer
Nr+wOjbW2gzBknbUhDHzyNzGzh2vDeoC0AQxTZY9PipfKu0MWi0oXclvfBWB9vgNlAavjG/XwEFt
yTIuTO1eMZlRPlxiduq4vPecBJA5cvNjfpilKShI3ToWoQdGqol5DtcE1tyFHJ9nJ8jDDW/kM0aK
pirTRzGTLasSGnTwPSsGUbVtual3rpcfgRp1ofPBJaDmq1IrU96NwA3Hru4oNKClVhyf5Uz42R2O
v0c3tvy0y7ngt4K/ISNzk5EYlrD5ETJhFlreWGS9xy98ewV8SWwqAjUuP5911B186p9dwBwCcT8W
tnDqcgtRBkqoEHd/Lq5PACRTDvwBgK4STG+wqOD1GdrwOfKo+kJxZ0rZtG/sWcoYBljXbSbyls6q
rxKK8gb15LtOQlpIC0hfnHJFkyUKbwasR9gXeKb1xnRi2C9HTjHQGvj+XiBqvBGHzwSo81d20u6e
kK6mUAeEdwsIneohVRsQlMCFwTc7UJuvmZUTbtoq4kW6/QILTJcElcJoz+O4rpqFw7TNGFQHly79
nNxHazhQpXW1S4HDNWckiXXWNRRcrYecbQjU5g7P9NpSXX7qAt+syWXWB2SR7ClukXRQD3OCjNok
klXl+rVsahpLhR8ng0UOkB05OylKYw+8vGtpeao6KZE+Hikup7BFYz3mKiqv/4j2sVIpCwnYJGbP
0Pn08Mub7oqPBKQZ4BpIb5VmnkjVVYWE4Blj2zacujLXyZymZHW3T1JW4zF1xxEO0H7hnlS97O6t
LjA+tG+CZErdwxUMPk5fuglAMu1wst/vs4bJFSCpRiDWEXGztdgSHRHqnRUHelN77i6uYR1QUoHN
pUhYftnTSljrgAjGbIFUSz/mAmYWwIYAk2o0KNc8cen9wutp90C9biBhA1Mmi+Fcp6vUXRxvgAff
EF4vhYa1DG0mq31R2lOZbx+3KihhQ+qS5lFZRKEuvSLnlJUh7OZwzWiKDWo3jbndBLhlsAScRwtH
BfRLnYz1u68c3xFEk/+YcfHtd0+ZIkjACEd485fRtsJQDLftvCmzBCj7LJaYIuDZbnzGUyGrSSOP
s8vMzVg4X3P9zBX3PQkXrEd5+pM6wH70ysvfsRoaEhXO+nka1axdGzCCQ6nwM7ajaeb5J2ibe03T
uTPJMC1Y9TCfmIEwRIDXi2eJXhnB1dknVlvIF1NHooseC2hVXhKxeNjds6Z3n6xOPgKkdP72h0SV
ZmW4MGKHLRxFt9wWHOYE+vwlgd1haLH1rnKavW4ccNqvrpo8/Aps2/IM2aq2362KYQH5M8QRLeyW
FdMH7q5UVM2+233pslRaIOYagI4Md9gmS6v5mkqRTEQqM1VIuxE8UQAzHtm4OqGjgl+Zvbg3mJ57
Usz+JDQdnY24pcOvuAv2GqJYOYXbNOKQDcteqtkaGepH2WEUheWRB87fAkZ3eQohLlwi0prYU+OR
r9J9tut3k034HNsDsLzBoke/xu4brQ02fAmGdrqzzqnQs3qiSKV3ZJVZ52f5Yl+n/rBFXwjaEAyE
R91OnSg+r5qWJuH1kBhXcKPPDcvmTP+/vrEo9SNyoooT6Rtt/MFoyxJ6ncL3neFqEU32ZVt4G5Wm
Xtb62suwV2AhuBEUbeJ07lUCqAOP8As9TYXdqb5JuPvHPeP77PEEeinIWhWEhgoSYIIZF8rkKlFO
EZpUY5FKaIRM/lv57CRoS4FAx+jzwZLgxLrHMDIBv2Gyj+hKM2CCfBGuTE6z2UGXPMu5Nuft0ayc
MJ+YG6kZWR6fRKTsVtPXScDNRvoLd6US8K/a9R6TBbcIpcVkd2obdQkrs5EItLQzFY3mYdDBveiO
FxNVCjLu2YZFWK0wN5MqqpCTq4LVghMTtX8pIBjR5uotZMHdYlnMUbfQ3UCikeR6VgMVFNdA+BqS
rNPJ7SYkFFxSCHLnhosm7CGczbuSaXw9KWGd5UoLKNznKL9oLIlHXL+CCS8ijckHtZYu6xq+GUyf
1y8hqdzEVLrvWnhlfPmr4IyfNYhQGnSsDnXIXdprXIyHwOjusgFXX2o90d0Wh9ZcRQXoT0HcLDLe
g/WvSDPg9LNS/9E52EhI0YCY3PexkmIIJ6b0h/B7RcI0TYkvJg5IAIl3lf+Co56O2TwkGDDOKjl2
qezzsBswYkPpin1IgmRoE2D50QHOAVE0CmrTuN/2LvMgUvS83Aw4KwbE9lHlUS1brl4vxWdrDwsz
xRNLZZBjxsLXIfvD3arTr3q0coElwNN0b1lV+y4asBZzvW6SYtXXklH9PnZ7Oq3Jy0ChKK/yBfzX
UyfTMlqqaQmG0HC7zeFpgoMEWVMXsfZgtT3et2RPTDJfkRzjclxzREqa+mTBmoL8heHpXYvSXPUS
1s7y2TXAbaU0/cniv3eQk6qBm4hzsqaUOIuwrGSdpQqBW8vuZ2qRwjEFzVN9NSLpOEnC/EOGsyWg
o8ruBFPHLeoI4/eIWvQCbsWBtsT2g4tB2Wa3NEKncePkxdFSTgIjJQQCfrk+lgcV0GLXQiu+YcLP
h7+nYXuUxwnO3bQ8BpJewgLXL78FZSFP3ASBjIhgg8NfMOXy0ZSXXQn+EUxBRhHYqbysffortgpB
dJtXYcBAg4q0fevsWGoJZAJmlWDTF5fQKkbhGPfCwjrcRD+MeXWcoQgZG6/eh/jYmK9OD0e3mNab
iSIh7lJFQVFg3o1U2YqnDTEPFEfTmdTGU50WEX8twJNL3T03qI2Z8gCVDGMLE4fIYyfelq4Md9TV
h9fQ9ixAr1xEtcblf2yBnclfuqGRnUHJrDM+OlxrjjB9ad8g0qmfIJwE35u1GI/+QAr0ZPGpfZvf
DF/dprcufvrRldvMdu4DoTV3mq6rVzZUuZCI7zOb0Nvij0YItrqIBuGx9tsUImpvrsWqNtaeVZ8X
JztRvKiYFEvK6ecyOq22xkOLzxEHlbXU4xbTN6C4hEquKNBaJVDsGWCRJoPc4YwaWfbpCcUTchKj
tn8/MOwI1wUUTEHK8eizRNodG3QcsuP2MX1PyarbIkWAZceGRkjpytMQxWqEcAUwBr6DWwCwxCyI
3kqPH+VwkLiLRkUV1bt2IRJrKes0wdOVmtRAIOQEWCoM1EDzR2UDdrC/6XyBLyU5JmKxEg7YSLC1
1qbW8HGaW7Plixqtf335MOthA0pX9moTAVJXcNLOnOXhtdOkj87HQ24n79VDQuHgWGBr/XJXt1WI
1sUSO0JW0LNyHv4cJch550XnZdjgX2mWMBa8MkgJihkSnI1x0kXYLN60NAsQSSKA0UAryYSmFGOn
xDzFD5UtVGxmM+3xTmYx2OsumlSm8mxu9YDheCSGzHWUdQlwZ7MG0x1N7ey5Z4ikfGTowv1hlW5Y
J45sABjQ3fP3uuNFrAZpv7xEz74FrmJgA3nkhmakgJ28ox/0mm+F6JD64bESPO3pkF2gyo54WFt9
p73icAPhPSD3M3+/U+dyTZ2KJLwKEI3CH6R1Nz4xr8tvGspRq1sXJug3oL2bx1WPPPv03l8ZaBOV
9pS0KnLp19HPgAAU1BvHQk8h/s5z2mI5P6ZhQI0T9Mn+yT1dc82vLS5bzlcDpTLLmqBpt8VWksa6
DBVaL9+UAKalopV4SgI3V5kgMfv3t+9QJJYNr03gzdFXTOpiW4EpZeUwnq5tWj6d7twExkZB8kai
x9LDKbSLL9CeHzBaOjIG+MlVmduGQ76EvZKuYTglWJ7emgPzgo49G+PBovZLwOYBr8Sv7WALDTYn
1/ljdLrOupe2g4lbkxdAOastEPg8n66DLJBSz51wgFF7x2TPdXsfBNmThw8FKAT0Q57UDM3MxsaR
442PR9vuTM8jnOHANRzjtinJJ+AkzSlnJJJF7GIjNUVM/Mva9a3QExuCezvGnZinKMvFbcoHUugL
18X6Pm1xlRvk6sOLBVl9SOUZDUFIavbD4A4dEeOF64OkTjI+u+aPzVL33VgkXT5RZelqseuNhSBC
kJrzSMog1racbEBCfpcIlVVVz+LXsu6KFtofAJeyI7Gd4wMmc4OFhSsf3MMZMaAQq1Wfs5Yisgue
/DLL+2PZ7N1LB5Z+FXsgZOig/aiTskZ9klMjKrLzNFHKREvbzmpBp7BbsouPvipllE+ARTph+bR3
riOisFT/0Psn2iQVxL8iq63QmY+ldHREKapRGI96ZXTS7EAntXbEl/aEPfnp/ZoYkQT+diX9d4GK
4vqLj9jr5KjD003OV9jlBhta/jwgDVUoLq0JjglZdd5WlCJjYndsOwf7t1UDkraJAyytCqJdOi9P
Pf9bgX0zIvqmuNQUgJMYLZ2Zy/03BldAIagb6aWdhPq2sa7ZZLGKDnwgJJ7FugCsocgBrioJnnE4
iVflmNtGC2ABmfnJj+kON+xPLbERdCYEyE8GV1+GWZGGubmdkLBoa599IGuR13R8THcX9AoPtz+O
JsDmyBWzg/87xopz0dvoMP2U14PBioag3KrwUUYa+dJbeksPmetY5ckLwV5jIpz6Xi/hu4IjOJeu
7D6/B0lsNeEoIRid+zZix/E/8pWBg4bfS9xxzbaj9yeueDY6S4VXS9O6WpO/6KHsJqEkrrExvquv
aj6hpdfKkIKw7Jh10jF2kO5dnb7qSLKduAa8zs93j+lL7hi8cRoqg4PlE9Bkciqg/0ZEi+BpjWy1
zAwoeKCFcHlVf8M21AkAShNO8SV6LG+MxNwBF0rtWgZQTzdq1i8K3H12pAruG6EcY3QnJPd1doYs
92K1v7UdsueV6hXcIaREiNUYl+nn8hum8vs+bY32EEBDttS5c3NjmxjZfQG0YpWUCc2CE+BCAos7
BvcPevkAFgqq2b0ikpORIzpWj5ypcBi+uMxiB/fUPqzFXwz6yNNai3tslQw7fjYin7ysbMIYfV0Y
/+Kvx00fQoaFS5lIo+vicyOdcJrnOWwGmiJNzKHMtS5Wlq0mebgkqubW6qakNOpY354oy5AJ0lSE
+P0tr+hDql0ORG/Nk8XAjqC6XkBgwhI0qQlH2WxmeNmUdp/puyjccFo2nEq5nTZCeIX3DPvKqYWh
3/yYcMdCItqIK/+hGPvCetWKnq8uVwSNtWPsN8iREgASqrFgwRlP5r3K8m2QGM5/YH5i9AQ2rNjI
Ou/Mo9vKfvCFfMKyYiBEHmht5OB+weA6poY88ZqWxEJQwCzGp2hRduYkygwf41bndL7o5ok9cQUC
aahbjsYkQdsTW3M3DScPOEXHjmrVoTTln9LfacSF5amxzwhgV1pOSLdEagPmtPFqGwcO1+OawBCy
iaQ2NVaijumKnEEu2ONyqC57oCZDVtTBeNSku+1IzLqD2cg2th6sMVnqXBFtBLtpds7nVUBRwgXx
tz0BWibJ9Oaay29cWnDBMBV/FGchykFI25qhsp75zGB4h6SeQd2W2vkceC6MKDo7WohXRMvy9bch
b5AKcmNu4jntxC1a7KZga6RezgkZDrTXLpbfh9WK3RQ50bpAz1dfimxcOcmUbAEnTX6mylM1mtc5
GqQghz7pvl8uFWEd3p8/UsQ2xnRDS4XmMx3PNlaFyZzgRCD0yKT+h/KNOlIJNz0thZiQQ6PRYO1n
Q/gNSmNjuf/d+VXspY2jD1yzl+spDzJm2hmS320geQLVhdR8NqcCkPbsiXl3Iq3Xjg2DQBVSRYLk
lflZguV1XPazU6G6FFVIoTgUGWQ/9bGslbjwt0Ep02QlzMxVRYoG4YrJr3uiVSraGd7VOIqmZaFt
chKuRbkQ3qSag1jl/nLOtPzSBoAQ+IynncwS8AtTM+FTNA9iCMTh/SyIvtUsORfTDhMFjLjZ7DcE
c99jfqODWEIQgaTViSG4y9KiFbLAhr2CjqeXUWrL85BMf3qwsfLP+aT5xCkyK0aHj3UPjaefspRM
hlKLAyuMTsDd7eH2KWAeYlly6Y8moO0swSVoyYOBe0bgwBA/hkRfh5jJS24zXajoDYrSRZPfO60d
j7ZEMipyRMkmU/ci+Jls8g4g0LxPbJkhoFkLbX1HB+Ki0lZwVD1Jb9hs5XcgMMDW4vP8WgKxVJhx
Vz3QTy2XvibubF+PFoqAHISeO1w2/MmHYv+4fbQ9W6mZPz0CCuANIh5nJx6Cka6JWJ+FpeXxwqvX
8K4npmfUf1VDjFfTrgJMfRv/y1BCiGmFP8l6Xmbc5fzbrKvPry7+N2odJFXxosMtkCDaNIxzxmH0
bDhcuFC0Jcxqz2D8IuTU0jKRZ0XIf213OSg/0Q0UfU42hm2SRq/qjHQdX83qYjqV9NDTd1O01+/O
DPh74xhOqYhmKYvTaPJ+fap8WoxYiYwHjhYzGxv/yvjqEKkz3wnKTOOem3JiC67KhL1ENOlN3Df0
ZSwQzuMtSo5l+FygIApojklQXmWzJpOnQY3mQQ9a+tXNDhBkuWaDLRKyoXwhbT0QSNzNeghxmRGo
hiU8HYKXGpegVdjdC40F9UUF5eXa/Cnf1evdoVn15LJfFiF+BFPo3BaaTVASJCWp6Wt02UJaVmNm
ZoofZRQGarLS6mS4gtJZkittc5kaoFfEno6mLpKkkYzYrGBvOiD6w4NjDCp4hQFf9VYVBWPdig5k
52ulqI/z76IOiRtGWpUkM+y6l8I7ukhsYaWsKM5Bp0voL6qMs9rFmdFGJ/MLwkYFmZNE6/Fk+GSb
Jal5dRv66ClXZcv8zST93DcPOhw+EmxhyTQq2SucXMvwngrIHjQNwvIK88qznUWZ/yvErEcnRMoP
O2nwVsyn+qoSgMzmx0PNtxJqfxT3OHKui+UkhTNnNUwqtP/GIJxXqh8eykaiWWM5Xk5EvZkp8Z4f
lFwzwSoJSGbndZ1DMQKOeJFb7pb5N9hCmFZ8P6LZj657Z9UL2UZBApkvCASXDBPLqTx7zVSfGfMK
t7a2Iy3RMWsCd8XYD7fEzNp12+a0VpFYPan+PZGKd9NFLmECACVBhKfePZANUONbncO8mOIxX81e
WzLuqwF1V0nSOhv/LJV+0BaZ8lSGG5pJ04+GSuDSYI4ZI4jGjS4P5xhoeCO4yMN3amEc+seOumas
o/JqYyqQhE4hG8oAAeScdB8JK5KRvUVZs6uozjqkwstB+T6QGGUnFgTzXgJezp60CdQPWakC1oLt
rDEf63MfxLe49kgbrBQRiAUBALG90Bo1+rnAnzgex/AV6uXrp1HwYTQ6M0I3KFi9nFW0fz7L2FGp
c/y2Rgkm+MDnEmp/wIOkFoHmcQ53ZDmGs2atUlyOUQ8OLwqQtC3HY6/BqsPyEPAHyaxSZoSYcFOl
9bd684Z3TbLBo1q032JXHrq5ZMyeW96WH6Q3zhoQa9x50glD0qmbNJY0p6QRNBnIBvIh5Lq3Tzbl
3sTwwA7gZRodsCKsrhbAxaBvuVHbVnzcozMTzpprydEJveo/OPPPKx3ivAbEe+76rtD8aVSlIrfh
eqoJCYGONaCjrQIyxIzNIYbusy2d1YyCXyt7NSK0+G6DMdCm3t9c1bOB8f3Xwt9uDnqcXewnaBRc
ybx3axNVdd/ZLK8idcs59zcS20dtZmrADGUhJU/kaTjIPlJ2v126Sl7ZA49sEs6Im3YO2tXG11Tx
F3lQz4NQTnVasQuaLgJRBStKfFW8TGdNrMFXIeyTbjPZTZCcHL5UZcm/GkWlr2YzAbzklyMqTF0j
76X3mm5uKPrJzZXB4OJ1kVbUWGNCfsRbBI2WxdQzYvmiWtrkOMZ07H7F40sczCfycbFSbqMhF6kN
7WcSLw29TEeJjXU0fZm0nDCvJPSI3zhtxude608mwW9pTLS5JikIZ1Cw5x1KG+/2Czqkc12axEvn
zRrTPPRN73CahrpAmSTVXp8dWtT7INvhieQ0G4IHUhE7ImXOurOXt8JXi+P5YdyYUlH1f1FiByAT
1buiWP4wPvLSDa2k3BkJkGuqjCWw0c8dBlCQea1KPkEoE9VuMQmTAfqrSR1M+v0PrMJpV5y3UihN
7lQtgpWk1LxPwNTbDH7LZhJWqSf3kFRajEheGnidMvKO8ZBJox5WK566Z9vQEAWdFm2puqBIkKcB
IcEfd+ifwy/qBdl8+VAKeNLDNNclnFAkCxlHelMgMgZnEcyWBjYQia3MthVWHPGKB9LQGKLpv7O6
suE2NRnuLrxwu/sFEbcVyWVWDpPVpXaH7fiUPgX6FpkGECxKEllbIYLt4WjNkfd26FjDOauUwnPF
sC8nawJkrDzBbTbl87d43c73jV0XOH6H9DhZ27ZWiK3j+6TNtEA8cF/JQfams1Z68G89yz2ucAks
oSfhsl9tj92o9PUqno9QE9A9BfoW+3v1PjB+WVVHNomvJEZlU/UFfOw/cNljtlpudfoL9gwJz7tT
u2sFhUBSdgEiU29KXEcQ6CJ+iXatGPjK64BZU8lGapBKmosjcF4a/tWjYk6IfX/68uz/OM5FJ99n
+gb9+csDcb+wbEv8FMJUAXdJSEZYNDo6gfJ0n1TllP+BqORPcwy3fOsNipDIQNzZ7t8w5E/p29GM
05eNWQh3i95/a6Z1Qgw14abrfSsi/TU5qBLTFzeWum8C3ENn1p6FXwFaeYCi5SEq5fExCy7Yv+vx
FhTLsjhLU7rHGQZHxJAUyJ4/e7ot8vowxmsvQ6HixISfR4ByxoICFydLj3t65jKy5Kc80wCRxsUp
QzHhg/qRwLLw2L4G+/POGrgMwZRQLFHrvtJVwDbsej+DEYU/XGAFtG3s0/kf/mpiaVR5ZUDKyqdH
LFn7nd5c5+oyz9rZhPMjDHpTVf1XGHqwz1vxDYOrb4BfT1fogbZ7c8wCRhj0k7rb33IRfK6J82sv
5WrH61AdDUvXCC3H/U7GM2rF1iJDC0W0UE/iMKOeqBUeL7JU680Qyx8Rncjidn44y1wkhBC05gvH
P75Xm9xa5/d4wotDmnO7ReJvSSYIt8c7J+UPMyd48VAug+q0cI+JeFKyQ1PyQKLHwz6vQiRinxyD
E8lfF9crfSpmwE1Zs4vWrjmHvQia25x03dKrinGLEWRnkAURYZmAxk8ChDdWqaloq7GvzUCaLX8A
1+apyTGjSsdZPSWkeDBmYoJ0EMT8I1nh0lQgkf5RIdxpyuqgAi8HhUfE0zc6Rg+cDDgI8b7kVMoQ
+U4V0wekjAUSatVzlEQ9eA5+zGfxUttxdAhktGZTaQvzFlusSSSxSg1xzhG6WS4ZcxQT5EnWXMpa
eIqds7pqw2keWueikg2OWd2Q2gIcOvbpolxzhQOAUGLiZMsDOFTJIPUMuy9jBUmzNJeHVFsJ/lLU
PLVMrh8YBDlvt0QfC7chDjPoSwEIWjUUc9QS90iGS1nbssaehHJXMg3aO0ynzzbsA7r91UIBdvFO
np2CNEJ+8cK+vRPC+Mp8g8R52H6Xdc/3wNN0Hxg9sOeJd01Tb+0sbtX1xRUk/XMP+g37YMslPeG5
Tz8icyp53HENsLzBrnkQnn7ewRRd+pQsaN9pNuL/JqN9EXKl7wEl6y3nW+0jMTrfpRzQEbeFtTIH
fK1mmHfaICW+nP6530rnt6HfYL4sxguxlOSckkOisj7tMGCwzIY99GRAp1/bdBf0F8BOkrKQfpkD
Q30qH+Hs675FrSdxR1BaGa71qc7zLCjWH7WLcnRzsuLxwKXpyKoQNLkXI/bdDyeyzSRJMKGHoU2V
oteh4edJXvl5wBPs8A4hKqF7c2E40AfHNXBfmkckO7CKm+UffTI2hu3wnbnh3vGwqNdlYh7KTrnE
xq7TnJOIC5t7rsnibJRDLGAm9ZxueqbuXjFY0SPSaOx3RTIgyIPXIcObWSEa3SQBPdiCo2dRLZOQ
K3I6QFDxOVtau+0vvkCq7y3Y1swvR7sLq8jXaBjhsLEkI4Pz73687sHDlNJkouMVm27CmO8MDr2j
UrHoTO49Qrpby+I2sR1ylgrZh+7XxqO/TDOVpSeYF+RnB9lnOpx7PU24HkX/HAycmDzJXtAJDqeM
ol1qFTzw+n2tk91p+GtpMukKRD285BJRlsCe76kMWAnhwBIsVL9sgRj6WqEmDST4Y0ECCiB8pzmD
hvwBoIgJyW8u2nSE5oGZT0rJjH9Vb6O3DJqOi7qlCQfL8tmC3Rg0BCb/EWkz9ioPQj2PorgBrOgv
80ztnJcwRPF/ZnOrcb7oTSbkwoGnGETc3xP7PfsbsAfoR7Xa6jTw/f6IjGMAcLxStxtAB2/t9TVh
3FKqgHvyKDlzdkTJiU6uZY36VZu8qIjZhq167+9QDTSV1xidxAdA+1kc3oFefalZ0yn8+fIAcr84
JJ6nUpwKnpV5LUvTabfm2LM2LStPTnDIJjeYlJIOOmrT1wZaWV69Bgianl/O6LxFEv10GXBBTaJS
k6f5MecFXHTqEXKTl/G8f/SmkyQnVH++VVsEvSQigLIZ1MRylWci2eqNqCNWbc7oRvlULt4hEbzE
f1HzkB4mN2bI4vJJ0V1zfj4tNJvBWNuQkyxOkuqwSR2I+VObGcXdWee05j8aEAizJXqSDJWeux9A
Mt4nDBLL0Dbc6Lbt46F2MiN4oKoWPYhWeFTMM+G5M4wJilS9ZmsPK/MfRycZCPNcopebIgqrc+Qg
wdrq+LYEGKnQjpjRifaoCdVzrzQUiuyPyboWPZ3fwz0N81O2lY08qPiAMif+oH8rS/Vc8b1XTI8Y
yb2QMzb9ljMxnDPNWxIS2gZm6rIfpVo+i1Dx8PVZhDi1mwDRGE3VHBpjoVrrVECtpRX6wyEfjgri
tuOhv3XoHBu9/HQsKH2eFhBu1k/vs3cMxT30tF4oGGRNsZjjpUtRmMxVeueiauzrdVmrrdCMc/G1
jNJmr/drBxgSAI+fZ8ELCjP3hIXsNLi/LUoRKU3Yq9H7kVwy78HuIPKMzFWeaEgvrQLJBBCPNfOy
s1dx/GKVJUCGW3+6mCcYJDvfQ8A3cDI2MGRcsgp+dcOzR9ZtalMilup81vJZ0A4A3+0KNrxEeey2
pqxvlnOB8eTgAEPDY+N4uDAU3d4CZJLLLiZgAIHCfrrKy2VciGtky8zhkTuzywSOye+qWFZV0+i+
DgHVN3sdRNCNVkhKmkYN/D1SjXKCMWRb5nfxb1xU/WToHNYihhjKvZr0dvToJfRzS4LX8lfjr6XT
6xFk0gMEh/iefl6mI2DjK+vOVvYZeNkFXEjQj2QHpV5MotEok4Jpp3hVcOBC+FT/tEtRtozKbGAz
sNJUSMmU7EUr4VkiJnzlQvpvosIXXEqvwlURWk8e3rnHB3bJH/O7Cm62N51jnsxxuu4bDg7Li0ZB
/tYr+qF8dnVve+QRv8NHcXbKDUs5ciPdDivfqCzXgu9VMyCjIm13MeyJm1VpjMh+99m81RvQWLRk
T1kOcOmVNJuUxmp8dm12HgB8Q0XQTfkkzqCbwZ6jv5hYQU5IU76WGnl38O/WG7qjTyOe+BiV5uAf
elCPkGYn4Z7AGqJnjq8X5w961VW2mivBWvqXp6kXNVks0EIyuoFZ9k8oc3LknD2LC6z4X15/cXox
NTxP+YhBVt5bbJjCW9Gyb98/wxtobGm4JDKzEEFDZNNcER7pb03BDREarLydp3PxKOgjswVvQbA1
BMz+OYLiNNTt/X+UCR4cQWS0OI2mHqQpgok4n6tdtI3yJdvtA9MpJ4LBRDIHZOfQoSxThSRscJZR
BfNttwy1341HMvm9B0wf9LvWB+zAGQSlXCcfU9w5fsG/Kpga4RE1XGtA3hDhqI2Jj2v7v/NOMFgC
E2On1Ip+Hj2OsSDggHhXA7rJg94IjkGdaa/ufMI3Y8elLuia5vGkNnJSbjm3kkoaAMUOMUlHoAES
nPg1eqlU8tFBy5zpDkO/3F5tYpLCvJEFm6ekv1UvvpkuLRNL1VdYgcKUvD5FUTOSGC/cUSF6ySnQ
DW7ZHPOMPBw3oXLBVFXRbYT1/sSi/82lfg2JQFL3fXI9amNCzqJqGJflV6MCLX+3WAkdRFsbD8P6
ApppmRfzlJUH1aphW+Y9OY1JgF91LhosEJIn8Z1LE8FHBkSv269phlrRTotU6SAW8TP7S3kXIc+w
QjnBePY7ac/B1uG/4pDoJsj+kndSwTNH2aI6tzLMnFf3qCD1Jv/ju/BO8wiW5qTi+3HDJHOnY4J0
Iaxp3oFlSuYKDT+1f+9NZRA+KDsA5q44om7dUh+4hFZQUxZCySDmSjToD48h9g0fZIOwQbWG1MTE
XQFdhrQiQwuibN4tdtiq9oqGieH99ZJQND9pKz0A+lUN4n92iKEgjJbTNUBdgFb903c/HoHzsLkS
P4NUN8MdxJ9lLAtjAcGFS5sAkqjHVdYMiM/88MKTeJ0cqS52nVdVByv55DiobVRV2v08McDYuyjk
YbT4PA+TZ6058OpXK7pf6R3I5LWR5jNF7opmfOukFqmzt0DfllZ6FH1xV3Z6CUKRX/MzOKAqIAV/
3RWvOUgWJHxhPOgCx5LOq7Fiz+u8h0eM5PZ7BgWyeKERdbdEZVybXSvkcIV/0Q9Mp+0si76YbmSK
0jOT5Cy6q+xa31++o86l7JSAxZh5xZegcYkVNZBSee3Nwc7nVVCYltwZQzbn4b0Qo8J9v3TzpzZZ
NgmMUQ/GJ/6I6zqCRj903iydfP9LlGgyAPNbT04c1hhNY/pTAFUdHysTyWCzdbclvPo449WFy64D
KSF6J4emKm+fKVZ7Udu/dcdNVMxQq05ZhMmhxIFWqgB9zjegbOHUj3SSWoz6ilETsnHeOejNu4sO
P3spDcq3NprnnE/IlGSNN3JRCsfVLYCYUA3Lr+Y7AfXoZ4WVJF12qqIdbWxsOfMh0Ue7sMoajQ+P
7/M5RXeiWBQB/GTyHKmTzqXBDIQfJE+mddvCb+9oqTNgy6Kzzsa3TujoG8GOovIj17F0ziKtP0BU
lrOByYbuJe+hn+ZxX8mxGFdHX1sfFXcfVbLlPxuugtEgaIYwW/OaEd4D8XkopqS7M0PN4Vevj9GI
vKPs5whivLuROqHK40MpU9opJiZS3X7rLTmBcFHhx/N8PlVUVklsObTKuQ4lh01IVgZ0NOMDSBXU
2/nQZxuT+8G1ADiDfeCPXuxtOnzTsCyPt6WUjYvuxJzRBxknRzoG5t6OI+RZ2r0hgT/mpFDy2um6
aiYO48NGx6GzIJLl8VY0nlvf8vjJHNVb4eodBmMQCTIvEz5a9prWrmId+gcWgpghICdEBZ0eQTbt
MDB6hoWiAZS9eytBtT/BpzxXTcRJxiaeMVYGS2RYGMDsc/NkfVu0+i+5hvtFc1i6S4zf0vKHxZ45
teau7KoZ6e1p614aa+97FniGtBXhAdJQjI/98kBz4D+xK9WyNPc2yJ6igSfkFa/diRCKjt/nXMp7
du8pJc9MyWdofmmrf/0Jca8mCF5X6ZO5KRkHiN5KnhK4LwjUnEGWVHnL3gGG7RTmeKFPeNFBZseP
D8Kr5THcc7REbEdYsRSn+9KQCk0Wgjes7p/trWV5HinEdUq0tZZ1r2mQG9PJiVy/A7iaN2wKDaBh
jJxOqeDd6IIfBFtz/aFq0weAD6L4R034EG6SP2WRRQ98y+tlVRr9BJucaqoAIxj4O8u53RYZmT0a
hbVaIz9pXgA8PTniR1lDNyHjKSg6XjqbrFvs9J/yDHfsoAgPG1yzxRyNL/H/xJdfUdmrlyQyS7HK
mIaUVFvmVzfiMY0oEbwW4t7PDQZqiCUkzskzfz1cJsXBMZwIkdWuvjgSOk6p4f4OvgOt9slSts9l
pi3RIhbxtv1HragLoOZvqkUDcr2UBIjvUdWdCzGeNodDcqJNWpRN9A48+VxTr35V0quK05OF2ors
Nh2mBqkVP3MIZ8k0SjtFQpNOvR5K2I8FaWkL8q0aWVXE7GvMg5F4DCEjqbki5gRwMZYX7o1D48Xz
9al2u0cFoRCAt5y1r0AUDCm6k93ye3d+kHJnxgEl8hgQ8kAjzaYZubDDBu/H+7ciBe07jri4zdWN
Yov2qRAqQSCNPUBMM3AnCh/22wBQwqNSvx/3RQ3zCBKeBl9UlSQp41anaTX8NBke9eGo87Z/Nes2
TK4a4rIBUqu+n668Rx+lDNoaT1DRcUG5RWzQBh5ZbRmk17HbjwCdv7IoCHDZ+j7tV3rs6/Z7nJ1I
Zghmb4lKc43sUhwd5krYY8Ft0jDwTl40St5aIfPIy4QxyCX4E9CMq0p8jSLZCD+mWc21SFgLBvbQ
giLUjh/tM5ciwQI7VDbBbMKgd+fyqhGCiKgY/1DrBF6DLZtP8DQKFCZ+IlnduXIjTypADE5dTFhk
8mqLKnMYdRGFkZTSHfjfVy38AU8D4Iaf4r1biAS6vucFxpsg0mPxCYTBlTJTKXhAzv7iR7KMBt+/
cvI1zw5eai4ILrf5yEwTnv4NTcdztZfVO95viSPWjmjt3C13apQGpQ3qEgy6lTCgyQM3pGQS5xcX
VvJAXqlNBE5wsn8POHx+x0wWS/i1eiS+oNsrW/lGxY4t9N0y3mOYIhJY/DL0yLoRR3R50PAoWavR
bnTDSEKqzfnOXHBez0KV77+raXgVGXYa/kdxZ29E9a0hjDQ1ThrTaXjNjuvp1rI6gahq83Y61Muo
HqwtyvOa1h93k3gXj84X0cY30mkIGVCSn+Ybha/ROD04RseY5eNNoih3/t14+1Vm0CwXh8aE/AsU
ZaM4qetgjds+27I4Pa7V/stzU1LVWSMoPMkUPRakBUhK5nHpOldpSRI4hQmza6wAHF3xCZ3h19YS
RcBMMoBkSEtuQAtfho3+38qMn5Qi4110TaBCBaFvXncyAf26N70EsBv2mSE+kM/OpEllCxyb3SnZ
TLkhTbpNiwozcqeKKwPNga3QzUoMg35X0TznfcP47Chd3UIpvSNgYfi2jfrklJG7lsaucV3wCIev
YLK0h7uQtBqH5NDLSZkt0aWpkOslHwwjhWAexyLUR+fWb9DlFFFqKpPW+HU4R5LxxrkeuW8QVOVM
sHwV5WtRCyQwQ7irNAEgYzS/qFQ0AoEBRFBV8axOd3sfXrWxTuJw7bwbQ4Bm9jIPzxIddNhyZ4ol
GIkmnmF4hCb6mc0kzUD9D7P8dbe7DLh2DPKjFbRhjzs9u5pYgFpXKJF2SbJfTJLz/jfAMg2l1Xnm
fu402jKl20CTkuOGWA8jNfroGT4ZZnlxTgvlQg0i6Q2YHG9vhvPzjKHWbcShD9I3Cm16jzQydPnm
u4q1/irmtk6l6Rbh3PljBMv5xjLOKcyTJqPtiUW6suF76j65M4SFkoIvSZMREZ1Ztavahew2Yrzt
GwIyECgW74oYJCP8Iqa1AQEJDX7TmbfE1XMKJscchj/yUh8EQ2rjEwrL6PTjv929dkMkCDutPrTl
xI5DFZ8eQ9fIU7NElkON3SsHsiJ0skvf1wCMcmXLziVBNvAH7xB+ff8NzJ1M3zzjGq6EHOTRxfva
qMBqJNTbcv+OebrcZGzQ9tAY8pKgNrfLzFpN2Jt/VM2FZbuaSnixqi7nAd4IXQ2gQFKKM0jTRFui
6PvYWUhyDEBe+odGRVhfHHhL5N5Sn8cGsqjfG5euDs9Mx9joq2Vz679lbHE/UO8YQE4MzBWS7Ch4
T6uxJqDJiaqCfP3BkFbfKq/EyzSEPS8SDU3SewxKVbkh7tTWElRIJjXkWZi63/6uZkQNMtiBDcIN
iTietavwClz0HG3wgh+/pAZ1mF92fgdRZHWe5MCgnd8Mj2P0DnmSDnnQb76B44fvCXt8wl0pL3qV
scfq9fxMTQApHSGzGiZSx7QQfQcIHuas3r+cIJXggqOJ4CwieM1fickB43XgYMYwZLxNNSA1hWt3
0FhJ/tmgipb56KPJm74bl/jf7aDtFPsVvMr1PHNTzLaU0cqZ0zP2WAWxeKhib1fFtDQFefM0fw3Z
5M+32pAkKU/y9EuxB6CO5gPM/J3cAk+u3Sd746uPYF03mx/DiNDqwHDCdgilZ7j19PclgZduMGHh
280x7VPUdFrqUl9J4wd9eOEzdf0lNPprpHwZkgh19XlYMzvPO267jXtsVcIQ01DcseCf8Ck1hcg/
fhTBdQwbCWTpoUXv3mJikoNEnlx9/lyRrX8wyxarA6Jb6Co/4uFlmuHvtE/essvrd8gcmYDr7ha2
tzeJF4iF1U1Yhm5d8jJarK7VpIS1mDxc3I8C0CKrLuMkGQ8vTfxrK/KbbkpLr9efPxExalf3EpKH
V7Druc0hRjPueh4CcDV1p0HpBo6ojRuYYZTc0MoJDbn6HTOpFN/QBWODJ2B0htUb1/YZrlGeJWzq
8ccZkTUxORJmz+9xoR+Sjl0IyA2VfrRQ0UW3cJDxvAQ2J85oOkxbPDmtsyrkguwUGyCrmuWHXrqa
DvrKOVH5Xa3aCKVfMYurpv4JCo64Nr4SD6wxUSPGw073/Gll8rJGFpnnDTL7/dYaKSIbyq/YLKr3
K8ixLmp2K0bxM8TfA9iMYx5r5vuj3NVibNHBLC1kSRPQ6IUG4oVm6VQcqMwimDe/+qRbWWtJrjQU
MBYkjidZVl6WRW72x3QxfTwZbIK0woCLmqf4cyRMmJza/va+W1f6/Fm9VRyd8MugpWE5qaBg1vIj
xv9tDj7exGsLcu+vpSxdUMgeAqRad3RishWF9S01W2BlECjIn3m1tPiilCpcZZLiBfi1c+uAVSYM
jpBglm2g5d8gtpvEpy09PsHHy2PepSxbAhHiySeGKy1IipZ6N9mHLmctFT/Acvx3m4Nsy126NuAB
HsLLBwweX7c4u3eVOv28Z2nrYxURpJYF1vMws29FdW99HKHkytSYKXrcYXMtVuXEoHKxfa/5gUOy
AHeBLr+OdMG5Mxt2Nq3UCbaEO9HkcMj41zKwYlDcD0hkQnzK4px2Tp0WmmRwXJ3cCR1ntmJzwbnR
IxaxsubuEaxqAl1BrbBv0UYMNaF0FRDhfUKUenSV35GTrE1URN7tzr7IV1HQJ0nQw6PW9xibMQ1b
s3WnnJ2qnDRlpCfsj0Tbsrhxo4XM8I5qbMxuEAbPj4wMzDfLgWB2t5TjLWl4MR3JXdP3ghrY2zlR
4rUPunLlo7VLbyZVOFLn/ERLfe67/wYSCa/cv9XePWtfKxza4mB3QIPqo4ApPcnT63UiSd+mP9ri
yKUncmfuLnOpwFsZ5q7dZmH1nSSJJxykimNKdGI5f1SFWkQarpeOFd5XcJ6eBHH9p+kOWm23hFf2
g22B7ciK6To9YiCA1hMo4wBpnu2Wwol9aNoKtsLpMpwHtMDKxMhSDWWEYcJARx78CoZHv+NXyCvT
q5Rj/eUYiloc7CznfZA7/0FvtQg5kLfyShaiKutwOiDi6ffhY2FpaLZakJTTcq1rdyGLkBklil78
w/0KWHrWv7gfXzvIgUf8JpuWRVFOQRIWdRrZi0F62R2BaXXJJbQ5iCy1Gjim0kcFgHW0NX81lXZk
DEjwZVTTZ5gOrEtFMK3L3Or8YP5jQBcMIDz6jESN6sfUQ7olVNu3odCcs3qjoUdoghTfo4NckMI9
g5yk+jwInfNmvh1KgXeU1eCGojQuu+MJcImf4n0LaQ3jL9dY1EvaKJ06j2e2ASDfMjG5GO7Nk9NW
meH7GitVI8jzt62yL8XydutL+Eq8cX6MtwaCmEtNN/9hqO06F8habFkHESl5lagy/AsbaJ2dF5DC
V9HQbinWUMoOV4bCH4etND/cLnTLyw2kJEDxOh4MSZUSjp1SLyiavIo6SjZOU/aMbLe8MnTG8vNL
bmFpGYCDVWWybPuLzOf3pZ9tsT1q88b5Di0TVmsreQp0MbpgMnIdKEET7N3tKbxDcBLzyAz12w+o
yJGiNiteNyzz5OmNu6r1Xb/KHkOp1WwDZr89IuKRdLocuq4tjwrhv6Ozz9nViN/S8b7S0RezIw/u
88bP4rhENQH04fEYItFWUF1DNTuUxHKDDtKcfOpBcwr9sO/FVr9wBCJ2RJ0YjN6UeEjCvRCOeZW6
y7b3sTf9LE9G0OHeSGkIIDN8yBil8ZLeeg5aiuBQyger5QMnNjbWo8bG+y0UduGxW6l+WnNATlse
SEzilBt5BApz1pH7Ib5z7PCaeJ3Q7Qxx5rDYtgPJ/xuIx29F31wkL4grD966y6p/7wpCroy2gM1U
9jjp9yYo5We4h+KfWTe0fOGAJN5t/k53sZwaIFI5XaNrgRw5MFTM94Z3knfv8JJY6ksB1hAN14FR
zZD3JZAohEeicirQrK5pUmqTDvHvDAHVu+s+Lo565cg1XKRkiDWhSs4SfP8bPIXHIqgfovolO8yP
o9MafboO14+zX3W4nNGgzNAv73Rop98PBQswSSGiAB04DeOOvBHb6b0fNsPb93NBRsZhdzWqQYad
5eo6+st2yKx/3gPHvoKv7O0bnRjPcWj0aliZQorX1N5tknxn4UgGyj2HaHpQb48nzVCjnIdqMt4k
jQyb/pixm0WbVUPfsck+oUzg52zWZJmchIPEiYGIZvC/eAknTZu3TR6Uewy9EXVvMcXe0ETjBQoH
pf7UrECnuYWKR8RgKBT6QiZWLM62Vo6g4a5orqFNHhUhavq5d5nat8noOOIImb4YH/vPjoDPRuto
FgDh2yADeAxwqZm3GYiASG7v4hT4ouRiWD6zNYTryiPibxB11iYAGOXxCSbY2jIbpsPvTVYmPo3F
LvXeIOxapheeKGDqzsJGqyaNQVHurZfzWfJpD6E1d1DLPMAV8JWhdDIwCaz5dc/Gb56D2hJNg6Ef
Y4yX1JudGhac907DBPBKHNFTs63FaBawZAcwdCGX8+Td4iSLpTBBJd8fSAryZ8OlhhYr7P0LL5xi
J4TPNffOcx1kKAXnGinPYu5hgbl/4GkIxQJmhIJs4WFybIEcdqphQ3VRGtxhoEDjisFfsI7Kc1lL
6aKDVeFkQQj2OE6B+AKdTxWPh6jnPUP+pglQuCNoz/9m2+Y1THhFugAWlYXB+9oOLZSFmy+3xBSr
XsmbGVrrEpaKDdBjX0VMoF60d5kEmgRyJIjjSfmHO6OdECXWuOYWphrmF8IYPbngN/MtPl7wqfEQ
1cyyBBAfwsTf81G7o19XpxJyYqWygt+xeLEeCYnHiSAYg++opfbhgBA/D1lAotdMS4/j/OedEJI5
dCZz995dE4LXkYguhhk4esco524eUREPLdq8R9JRDHYunD4TQ8vqJlbg/Bs7w89kafslPGoGbx4X
TKAPWw8v/xq+aYC2OOksc+Mzj1Li8r/awQXXEvsa65nTyzyK3S/9SInLJ33ncS2aa3nEmdp9b3rE
vMS6wxA6BfPvrn2ITzJZ0a/Ma77M5Z7/auf7OGFpbIs5feJoZkPaJG4OqJRub+R0+kUQO0VPmA0+
F7zB2RvCISTE9FxGrPtVisvI/r9yp/v+ECVjsOrf8f/7jujv8DWiPrvo1nKivPF1pLpU5I6UTxbc
PRKGlzIHjoLxasjJ/9mAav1e8rNir/spuvKUX0QNJCeEBOdx01uLOjsLthMH5u3uf5v3bpiNjBNc
O3frn8XsiRtsd3pr18nt6obvf48RaXI4tiJorFoi+qh2lJhrWSl4exdQ3kEFkKl5jIJ0tU3+6KZH
Rs5V93RJYDXVEJq+2ssV2WdWBnTtSobNWGb4rg4kuPjc3rnsGaRk57LEcyDI0bPYDZgDNX+52kyI
toMxXU766xaTa8oKEa1h6BI22wnifRPiTFGhAwmH8AEzVlcawhWeqy8r+5CIKRnnrxdaeI8gdsfW
GwwUp7D6wqRGodMyK7MGPVpUX989wDilczzbJwojd3gwnet9G4u+p0N+O/YRGyXoFBGuPXGMbNzT
mN6QgAlQ/cgje3SknvfykzdFHjOKmr7wMORnd9Tx1BcGgJa7WRqKUcXR4t+h4xCyVlwbXy+e4aSz
SHmwfYwcfcmt+C8pRBK3EJETi+gYTDtqt3YqieiLPdRQF8CE5I34++R5D3Iwr7jjYh9bNahJGIo8
sRdxbnluTNLLOQOd+WYxiwscuZYBPbdGwf77n92gAnIXy2+Oe7WBnpF0NyeRGe8h7krGDDgD584S
nqWzMb3XiDp6J5lBq6kEziRsnFOT0lOLO4oEFBBMO4QbTGSJZ7pjSzr6FfyyWQO7lxVq2lYodDiP
K6IEWSk3JR71g01NC0maSWZPnquvB7ak7Cq6+aJpAV7zQdbGV6eKD5sB8yRep9ikGWF8OoY/pTdN
82H8PnOKDmc0dhYMa/jfgB1VapOMi/faLaVwRAmDoNKCBuGGUsVjTrmsvC5TPK1nm1SJOfr0Hslk
yp4jHOx1LPF1TgMJg/UXps7AtIwzFGafzlKhe9vbUNa++ZSCsLR+urHXE1EodMCKpJfnaMZtSI8X
cThcIiC7y3r1YTm4M3obThMTOI95hJQx47bwlhBy322qZYsOrkFRl/hhTRJU7B2FvLpyaL1wBH+9
oOyuGb/tlJ6uBpVwIuKj63KzgEXgsC94R/Ke9yqXZVFjafO3lYd3uIpLM5rWnNUlb4RbbLMcGMzn
jMCuP6tt90227ijwqriQcDIdyjIpZ4/OQwM1mK3ixx3F01buxmiY8zWJ5IhMt1hwgcqM8AOdl8mZ
hEpJP0JluuvJI7MOwszToecxE+bwsbWTcEG/xyWTZbvoTFJ2/mf6cNOgoqVbQwoeUks6TsqmLBO6
1EsLmM+bbj/m5+xJRNo6B9LsdRyTCBJIAyeRzOl6+Kq4gskKAVeVsUMABolmhUQCsi+SZVVkCTLU
LvY0IqgKADlctYAT+X88b/2T8sUUt+SCgfl6vsfo6BNWtQy1cqir2DFYx9G3iaW6cmnCMQgt5okB
+JTvtGz80QOaO3/BQm1e8LKg/oi44kFQte6qSsrBY+B+Hak8F22e6NM2vGH8XA9wTdXF2GnbcVY0
7bB19Q9+VhKpO6EsLkFSgecSUUrqEzwI2oA+sWGl7IOjGgjf7zZNZ6HeiN6RpFNlJdH6+7rb7YJJ
ejmo9Zdu0HhZQmljmddGjvLr/g8G4lLopxfxOdNgdSMXhzRotHX0yA8ZmnYoF/k/8C7QgXafTJj3
2cAf3tsLF3/OcBx/aytJGR2L3qX5eUP1K1reZjs02tNf4dInalV4t1CAjFKk4d8tmwWewBn//0qq
frar0bJW4Z9CoS/QQzYlzA1WVAbISYuzedocZea4Aa0JbRamDAj/8RRE7aYnz35s8Z9AkAtMJYIr
oToBXGExQK80gJ2fa9/rCjv3gc/zgddXdN3QwXaWLvkRUS1LIDFsACT9McVRgBCWTVfHVytlICEc
OKlmgA1t9iuOZ37cnWdxENIW/BIgPP+smr0692JmrQdiLjjZk40zod+W66V7fo2zcpQ/9hWPNIQA
SxTBUvGUQPX62QCCmtjO0hnjt5f6V8u7Y6LV+sZoqB9yCc7Ih6nmedOS2YlE2dyrEHcSVvbo9t8b
cNQtDkoXCbv1IQqcTciqoHdzYkNI0p/8z2UF1e0AlXcY99u/8PZGkwNn62uGuwwdtS19l93k3T4N
G1LTz4Rq9tcw/Wu/LdGvLMC4nsMbIALknXKdBhWu4mUa3J871svcNmMahgW7gfXLy0DZc64T6lpA
Qv2ndMmGiMaKApVigx7D/AXxHjsxA8PuTTUyPgXcJpzB4PrhmqRJ3Jvap04Qz3FLrBGVnsOQ0N3g
mQUWVdR18jF8Rt9C8EJn/f44U8VYRnf6Ka5vj5ucLNO6eWLSaPPSrfMxhN09Vs08oBx3TtHTYq0y
gYac4XeikVHJRQXhIUTiLsPJ3fKX6M6JFpAfjykIco/69YysMyYRrpjb3Agk4Jn4BbwXbzwRJzxW
DN5NBqrvCIBFP2FmZr6gUmOFt7YhfSMkBQD55p9IYDO68S94eu3qyTV30ZAEIhk2D0jg+bR3oIqt
t0pfPiyB70slCh7GuFDV6WivHyKTOoNh7EouwnYp1ggAgYTHujG+y+ZERFsQpQ6pF+zuNq0iUmj+
v8zOj+V3xVmLk17AhGMyvoFblNAICARtf/rybozCEoTI0ZoaTbNTosVoKWI9TzxRgoo8WgF/VQP1
m+nSsjrA5MWZywdgAKGCMlN4bnrKN1us4J1tAmbkVoCgpJDZ56UOVYZqwIu7yl0lRpbwHe+OCmZu
MprkjNsp6NPA9j4Jt92u81R0GsRnqOygDCHKBF7Qyzlv1poUPufnlsXk8WrdOSZFvz4sil030AQZ
KSCRj6jgMG6W9Iq8Kkf6s1Ad0/kKLQiwsNcpp+T/Isws/EznswJEY0b0J6kxpvNs4bjRIVok9E3i
T0ueeGfHUiC5UdI0k7WMEv0gYGf2E0gQCc/EP09CClBy+RD1+vIOS1/pT0ubXhYZYS7tYuqcftmW
Hp2bmjANkQ9SfEhoVPJ4DcrhkgClIgaX1LhuY3FP9vvlYxWEFWh2AxmlM9uR03zDUtlpWaNFDbxg
CG/lJ2Xtm8ShdgUXQzpRZH5Kk9mrReIjfBwz+m+TTjf4jhFhoxJZm0NAw9pzrvKbsGJnEnQqAIyb
eMQuAPEHxAHPhH+uFM+cMqxtVZjTVCvGi9I9kL4EZM54+2cSmi7afjDumAQsanDKr39Surgze0uy
iX0cq/5LgjUk/2tB6xrH0w6JIEuCAvJV7fNSovekldm0S6xfAi405usZINeO5SNU4iLOEW7RAUjY
Lv7ckFBTJ7jpWXnPljY6vzy8yFQu2lgmbLFqP3C+Nvf58oAc4Ml05Xfk8hSNkfQhA4PbO5uQ4XS7
XB3mZAQHZhCrs9UAA0vWg42+BDQu2hLC1jIVj2ZknITGL7lxEsqZ/LjJXZSpiGvNs4nYfbueSb9c
TEDJxEoM7jmt/efm3MYdm4AOxPiuVwD6P8LIU/eByP20ammJdxKhTYyAShPXfcvOEXaTQe8NK9Bb
S5E0FjWLqZjZNEvOS/x+qiURki7BvVfEyrNkmHTz68BW1hrdohrqIZeLgn+2QtdbhjOcOEwnCFCh
N29MCokVjlrTvwUXyOQ9EGnq3eIwS9UFVTHtJIycJ95nPp4SITRYzXiGdvr30G9GsXqz3d0ouj0X
OAuy2xgaE1AkfW1dC1n70VAX4/89BSWG8ODDZRID3NLWgoThTIzvbYqKlSlnQzs1BJg8PAIud/O2
h4tOa1yuQgPfWDoQtlesFzFMw8AAglevseCudfW11Dk0Who8sMDE80uIsGTrQ8Ct49UB2R/4FuBx
z08taWPIJ3hzCUiufvp8J7n7AFwNcuo8p19eW0RyDfNdN8VgUR/XOXwnDikk1H+hnrdS0YX1m7vH
09S0EVk7hJGLlnJuHMYAK3teHjqsPr7A+bMha+JMZiE4fNyMaNmlQt/RQlJw0+G1Ds+AWgorA2kY
usX+y5wLrhW+mrpxA1m33Ycchz4w3tFaBiLFGTG9A5onsCOtGTF54/Ra6+P2bZdb5mReHtov1n2P
Hi9qfAHlzkjHcXK9KMYkLAR1Suf9DXFiPna8IyvbsT2D57yRV1ojTmfExeb/QkqLpP3y8nf9fV7y
0lhty8pe1LfYQX9bJ7jcoaQPou1AmqzcsUzz0oKnDk/8bVk63cdE135mnRMvhM5PxfUuwAg+1alD
Cd8vJdPvMnzlTn304CNZm/GPVtwFQY1jAV/uevGXoAy1TPKa3nCspX3di3o7ew4srQJU6fiFgZ4L
X8IhRHQfilTGIWPdUQArgZMpVmcuugtRqKCeHW9f13jE0bVgRAafs2gL++igPokoO17rIJDSXpow
CLdUHekj6cdft7BYFd+DCkznb8ZYfJyQgC10LjqMHQ5th+CaZaqywR9MNXcnH8cTNEc6l8EnB6+P
0rOMvxWQXmXr5d7NNq2p52pbez3SzzXGVg+BiAND/8iztcu10xvm7szp9RQgONfDciODYe6K/IRv
KhCJqw44KZS6QTi2G7abxA7gIpzooNYcBev0AZuF8oYIXvymgIhouf7+m0X49HDiB3LK+1DVOLg5
AGa3oLl1XOdhb6OlT3DzPsINd1rrVMLtwMTaqNWvrVmGFhrXgh9eGPAXkQ/NBhkgBYmwmhC3uT/+
6+V8Jh2+FY2pJP/1givgTMgA4AsuLwdGKEaNhHwxi0gi2PFxPcT8/wv/ZHx6JeixaDuH72PK0NPa
5/UyRej/qPfwB9irxyhkfGI7BT5K4gzq8bRoCH7QHNVoNtoGyAQ8L1wpgIIIyEMaSJUGe1ptNYeD
vLGtgaHLQXeSegSgppV/3XMsWyN26eHTSQdNivzr4ugdqrbbyF8MvYkdrTHmu+VanAu6uvd7l4V1
2PH16Ac6OwsJI2fvoD2W3sz2FJu7HvxFawXz5h6kggyIQPszToMxOC4NaewOSxyj6woNYiiOw9g/
cwIGfIHScvrvQjkcSw+G8Q7toXf1oKnnh9K5XwNA/77i1lXXLJsOAfjVNGj+o1Muuo+T/+ZnwAEz
pSQy9YNdx5I72oyUqzzEFXc1Op7QBpZWypbinwSeydITeCuTIiu7NcuzYx9cvCO7+eKzEWQrCcNe
AzU0v7BRG7epV7xtoQudGvHhqaSqgDJWk4SuU4PhsL0ThFMAWyzdej3Ev6I1sUHWN7YrGIwOQaDk
CjihUtjTqLq+c9E34TkE6xygQHsoOUt+lbdcJg8lIWLP5yyy5ICNK9afsKJn9SIhBS1QWuAfIRD+
FwF7nn5hsExXblrSqLZO4KGyIZrSXga55HDJBJKERQamISTQXoRAMYlpC8u+YJMQ+Do0ULdMua+M
Vs910jon/wp21CfHzDDtiXIfSV7R9b6NKkdA/ykRJcbwvSFMaMNMwNIbF+IOcC474Lets+nMzeMk
6j8fa7L5escw1m+SwJIYjqOvprhPUCFjSCJDKf3LrLw94SjOPqQayqstl+ePDewTfNpOCoE2yHrx
J05Mbr9qEdPlZ6EUGYv2ydtmbaMhmD/rQWVKIukRtLn0gBrGXIX7B1wGWw71v7rTUlmkZCNkYsbi
ynKsIyTk3fcsGp0Ma0xfeVQBjjdMyrwAvL6Kk1HNZAzeVema+d88aOAyC/9NHkU8KbNkhL8Khz2X
NaTRYyQmZdfSLAr96z1h06q5XVbLSQXZGAGUrhmr02+gnz/Y7N68+omtvPYF3LFix+sD6bMcH25g
uF3JRM+WZv9+D7Qca12p6Qt+yatume+SuBqRX2PdmovMBecVfsqw5HHltf5fU6kmpfdIyLtgfk4v
0Cqd9APi6nr1drUAjD0pVbkUlLcm3AvHwL1Hpf/ghSrZqvi9L/yadzGsh/Dj8x6n+0e4F8RZzEq0
CMN2zjWEyF9Ewo3F6LqPjh3U55a7gL4rrk+gJqdwZ5EvL8Z0lE/FiSTCSX8hz/zG/QgT9ljhXjpf
Nifp8fYlwsuzSmTEjBcboWDB+VAZpee45BQw9JP+BozN+VbMKHPyAkscJc4M5D6BB2ffAKkgBtg1
B8a3LwlRQsXNCVtx/5eC/YVFM1auqYF+W6ZiXwd4IjJ8icXRjw0qwx6pq6qk2kXUzQRP7WHxCd2T
ye5MYVZDVForSHwD+/bamfpcRM59XHKruk7tWsmptiirm7ewi9+3OjizpN4voBpYEWfU1Vma4ci4
XvRA9e1I1vkxM19VphWAkfufbC0tKnYEMl+KxdV1In2KL4ZFEibqmTsKRN42Z/49GTO70ZQOsEtD
b3Ci9wQfohkwNsjmdFG2+tO5neYbTsLZJwM2C7maIws3GsjIzjxTpmXya08cpsEI3cq+fRHpNCQ8
PVxiHuY1lkYxsAeR8aNEIPUCVy/Q5CdSBkYingaYTkiXqzZ+Y55gLkHt+8BVuLPf+p9WyhXRwhzY
GEgVQh72KSRj1+LE5RE+AQMPN/gsyrtrWvrS8uJlq60kyi1IKSgLRGfyFQKJ/wBjo35XZf/WwX+R
ei0kcmVB7exl/9EalP6M1a/d1xxe6pzgWqb4m1y5HmSjfgAXvynxqzms/YYjcZkLvt8J72WgDEKw
WMg5oiNY0XGH0vPjmXgYwLO4Oo8tGG03EV97aXj3QfGWSxDcSm9KDFKWu4GkRt6S0FKOZS1var9Y
BtP3bitZi+XyxlJs8LDOeP2mCqH10X1cgJXH+id2aSuIdF1k02PlU7ovq1oy4OwFdz2Kph9FdA5F
Vppy8X54sirapEDk58H+o6Bv0LLeXHLEa22Qjb5X3c5KZvsWTsogwZZHrpkTWBg4MTtWW5CT3GaH
9HwCPsZy/Zeh3f6pSLPdKYMVvLsTTl4dMLRYDpRIqJZXGV3nEEhL7/UDnaSgFi1x9qTw0/4Z8r+t
3/xNKAtHvrRmyEZY26OGtD909U701gLWM+CjmTufeJqDxP78QihkXDJBuOz9RD38gFe5Q0nHl1Q5
nVOFJ18Z6ciazBVw/d+CrrY3cJjGz+PfR5aSv3gmz93OwkI3eh88SFMaCRi+x+MYmzCvEDl6BB9+
zPeopTVOAfKjt47MUjDl8vE8U9llZ9zHxCbD2GtDq9eZiAoEzoK8IYULTleBSGnCWOA4ZANnr01+
ppHafBVEmJYxEXbbTcyxG978g5dxOxyWQPkVfj2gFJBsK6JmVM5QujavGvtyB4PtWXglgsbaAcEV
RR+4D4eVAz2TRXqRrpN7t2T7HwKyffUXxuCmLtxJDH0d/8aiRXW06OaJfvHvTMJsH6mfAJwf5+Ss
rY8W2n+tzyTaCA4xGAgcaADeWs1UbUw41Ph7lFcjirfeBFi5SckBEIsryJCSHwUWYg4NWOX85Bva
eakbnu7LiuseeSkA6L8y8pGZN6wsI2/3w3h++TXaAvOndD4rXmrJOMYtNX6VrKY6JlU+2QctzoLi
+p14hwR4/PmQq07MKmXDhzflnhFvET+PI5slfW6EfrESd8j/JhcmZmpnvEYoN0MU85Xo5/dY0N8t
y4XHKzwMLAKM7w60uzJiIwoOrZ7bURTbiw1/SUDGsH4Ta/gO/LOVidpyDu7JAdVM0Jbgh8XdrVza
e9N62ajXvkNDa03mdtGlqM70MraUinOGEF9/cpPYXMC9T+S1oDeJde28kWP4VHnitZlA1fdCwVsA
XbRx3RYFKv6tIanDiN+cFR4nzM6KTexl2PhRwdNQrt61XoTJao5V/tfXBmdqdUmXgaNbxnSS5Ev6
2aAcbMf0kpIMMXeRc0rMRo5KvTXiGriiALkFFDuixiCDWidrjkwXipsW7xLRtZX4b4TgsdbzUb+M
xB10j9A5pxd8xGBAZRuTAtej2Q1c0wYrzCKkdXDIWEeZY9AFK7I+ygtNZLdzyPk/Ea2Muc5w51OY
amUa0B2i06eHIHMyhjgcOHyNXToS+H/V/pB2boAY19IV3UKnbZVjA+ZKUNPLT4+jKlNE/DceoadV
7+CDOMyyhH3q4oTReqXTo/db3tZC5lbm0lxpF3QrZ5sE/u5vJwTk1exxYTmnMriPmjcYavGzYBME
YMlgFQ2hx0LHDxpAjGdcaeWKnngf3xkfOUt2PlMzL3pqkP1lTbkak4wQMqIUMeO0UCicvBaIKGaT
yGSRCre6xtVGnwC6G97wt9Rqig4AoMPvCrC1yNVljzfHHGnM7Co+I9ycEsSxHWoEZsEg8bRh8Jky
05oKiKn3wzvv04l98AYh2KxqCqpld464z9dYK1bwX+fkEArfALNEPTcvTwQuxHms602Nlw3inLWR
+uQaSWjeCgUm5WL/8Mmkwy4opwLK7gBisyMnhj60sIWw2vRL0FcrgXXP3NYKrtxJMZKnlrC7rXrI
9i0xxyMWwf7SRNBIBEsZl13NFQAEvziuQrvWK4YX71WbkSwfOaogU/4TnXpxVTq/lvoBw5kpFmo6
GFEBL4PHkIzdcn9JaOo4EyG8Vdo3ORn5rdq9r/ezxiVNKO1KgTUCuQ6ZAuOlvFH3p3/vV7q0dp6m
23zHHlXrELD5Tz7Qg0LU298RtcLHkPBVUL7StpehFPKJL4/wiovkDbah4VVYyoXpx5ZSTp6Y7Ogo
2hPoKUjmaKFzmEqhFY3z1HKwhZO6XjZksH5lYCc94WB4Id4qLkToEHqL1hZy01qLEi0tBF0yrf6R
jvnNnHSdhSr/M707cet+vyApt0sKb94OK12FK6E0Vlo01f1MCvoR3YlpAj1WQTqXZQX20SM7nzYX
yEWL7k/QjTiaAc2D2nxmzJMFBOIBpf/Gair5RuBPxqqJM9QQSJq+z7W1q+dW1rfZ2f9Hkfr7YNOU
fIQapP2cSo4vh0dXOTPDo5H9QAEl8tIWLd6Rq+NuVZBelaLCi3JHT4UeJ2Kg8Puwlb6dulMc2NZT
owuOjH3gNFGqriCoJTF7A00my8IHfO7tDpUq04jxoRt51jcyktWCMaHeJh6624JDrpmjl/H6b2oY
U2fDR7ZywlgH3L7SAD2oUrX30Vf/QP0Vu1hetz/xTpghDl7/QgihG6FyogsNJopwSXpasPtWcXxF
p31tehpRnihjtN5fWmuoBQbCQ/u3uNNSA7RNVTTGHJaiHDNkmgpl4oIeBGFwJ6mpCZHQy9Ya3yRR
kVEdDvkI8fBC//2tFp0GuLuQ317VHOVpXjyD8kedik62OAmheUEEk4im3cpApnuaiIVQoMOVe7Gw
ocwrMEzXdpCHV1i/+AFkYBOwHch9GQ6wGacgtJLBCkeeEGC9tyMwfNj8PKPfeuz9pn9ywbiJHPly
jBd4GK2T/0FfgE/wC3q9MvnoWz9ekWB7SBx04LdUeKMY799tyCpFfmNlewR7DjkcUuhqucNGe9aB
kVbByhADqadYvPfI9rbiiUgmvM2qRgPqQqYL6tTxvIe8u4BWdK5X9BpTedP/+6o2OzCFOOrb5Afi
8zzqgdGGN1WC06tO9/6qledwaMQ5GQRwYl4gpB4LWDOg/8yJFVEdokr0N46qPkYYRuxRr73zX/bx
Q2+0IkUNkZAItpHpS8SRm0yzzoIwEBMO42KgBTjP6X6joU9iD6y/tI94WOFKjdnFIf8Qo4sGKZIJ
F5P2BFYsyx8FM1cgHARPV7jZyQV24L6Lu84hfV2Qdeh1oPsFn3ewyyz+T/ixGu+H1oS7Yq62mYkL
aa+6ErnNWsOuWOZgqdkwNkYoM8mNpIgD5GLB+VQzVf+61TXc8+Itl2rsRd9jr9Gse+Q1v6sfyVJM
3lbsz6PGBBwKLC9m+zmnrtG7lB6wBEJjy0WvaxLIX0tIK9cSZh0dLIhycKVrh1wDXcVueA7YELVe
S4Y0rZgdKLuAP0x2u+qRvrQ969DcgnV8+kcDrIkQkCEvqrEtph9YBTVnkIAzKOMzejej/gDqhY0K
399SLZZvi0goC3rawJ5mpCbx3wyeF7gOOdYQiDHaDQjVRKUep31DVMnQhQVEuXn7d+zQk6KGmjLt
As1DD1QpMUMqTu21SqRpgHyea9s+1+298oTOi1d/tDW0tD6e4XeoISfD+J41UE7qpg94eOHTtuXN
O73qUtvSe0phr6V/0o3NMKkGNDv7JGeH70X09zD7M923lTHCYo/rsVYSbLolQO3DVW0QoYHDUkE+
s4yWFKUUTyRCiq21mehYRvMnGCYrJr96an86OmiHPMx/aHkwHp4zl3QZDHGcRQdDgpdHLqN9ap3s
1fUl0PaGAPCL7yDjw7cSJi2hXkqP1YrNoNoDMDnXYvNeGvx15VcpFuc7pQ0OfZ79TIFg/hl/mX94
b+ajBdUE0K5+tUZvr7mvkw+JzuSEbjPILeXiXiKgneQYAayNSl1ufRsDnmQMW2oHHyNB9vOJYljQ
scKfwKio6zAeWpz8t8383fDc21tGNMPs9fYpJmi9L7UNB6ZwoHygEB+H3dIjKesHtqlwxhVpqDSG
O9AHp5zEX9uqiNp4d44gfmDzP6ZVSSRWOMpFpCWeAEPa/SbdtCqUk8VRYAi/zeoHNQSztALnyBOI
HCp1QSQ93/E4YMJfhrfRbmbFyyIogMmp7CvbCh1OOU9cvmMJlFQOxYVvhyjotVdFHTas3Wlf+DpC
EeH1iXwHRluHCq2yaFRewH+oMR4n2H83Q0EIYdMuSDuu/WjWmg8+4PBwE6o+2irKxQlMaj4NeicN
LGT4f09L3pa3hXBKwcbg7IrxN4P4s0+GCUC0VWuJHMw/DDMOtnazWVYN5jxWx+8m4EZjIlRUwQF1
q/Bbgek8HlmiQKtrRg587s35DP03J8TWNN9HD3WHbGAlDfe+teE41yGs61zRtcfBiClYDoI3rWgD
YNi9kdDl5BV7mlWS3Aw5oBX5J0R5q59dOfh3w2mnXbUcDtyw4CZY/3Uu79I8rlYhgpKXaTofuMHq
Lmt5Orfmdy6B1HKHArX06i0xsgGeLev+/J0GTOuZl6Wo2vgslKT3pcPP8xTtbpNU8HYkq6pPsu03
JeO2iJek8AaMinhNHzzGVhOqE/0g7goXtx3QTTbmQurP0lGHHWfDGnHzAoKZctQhLFnGT2uX409c
afGtXXscPTY2/8hEbG838WjcyruRjnnF57NS/ZJSZi8hCQxLbwiugSiEFBAHBScTHzrqU2SiTCuk
aBLDiLNbhCzGMIoKZcIgEAc0Ta3FewU1fegoxzw9gSu+RNYWCEO4pl2NYPbqaEAlH+e3GxiilHg7
obZXhsrz5E5/QbcWAOJ8v/qxExzlAA784B5SJlBbuXLjf2M1oCMpqfUBhS6osIqiS4tkCE0Ob4NF
sYcGcw1VYVE5hC5Orgh5YAJ/HZuSIKsalhbUOj0GOumBlWRsdKnuSOxSrMCnHo9CWDfL8AREp5px
XUx20NEsHUZ8cX7apo6AUKKc+1lvjXD+ciVlgaCzAGxlB07ijkpIPjgRhued3UsVYYXxODkWD511
x7YpONUnAlaGmprp8NDGzJOcEJwHXDzE64euh+hlXyVMxXBthGNXR6ghUPv8YEmpt/xj9rgHHJxx
te4pXhNbTPV9932U1uWzmBycyZdMdmPBY5LwpA/Ld2i1aqoQKbKvoHpqSb54YXMusOjMGUxh1iL8
eMjKm+XCmb0YVVoKYUqSQF5K4jOiAhW7mjbdcRrcv1smi/v+jkRnse+RgP/nf07L8NanGVPgEkTE
XtP2cQJwwQ2WYCiDCPTH3c0zUVydIQhU2hvkiwlQFk5T/FGvp9D/FK9CaOLgBGV6pOx+13FezSA3
uEF5b9hITnKpwRb5uVyc7U7IW3kViUvZ/11fUmwQ8lSbLe6MSVJ4MP2UNS65nq5iyQrqjwwH8m8E
7RbbEMu/88PDDyLVvUYY7G+SI4pitJ6AiO+k/0oHxiqBJeqNG0Zr9p6jVovVhOqFZxs4sJqjN7dg
hoACpfkERjEnq3dJlBivRtqHKfrGM8gnW5skZ4XxJQHOFfqSNFAktRRec8cBzphbUD2ni2RIFw0t
UzsZHzakmvUjtHP2Q+wYTJYPN1fF4HD05uG7fUsl1CNnmxJ3iB1N+kLP6AMX24kOogpLxC7kZ9al
iB8FsPaqrQtLUvWXY/ofQQvwXYVK6gHY7cKzf7ELLndYp+9k5LEzzC3M3LKR65tkK2Pt/VO9fWlQ
sA4fQtQT4cGZ9FrFrI2+dkt4B/jRJoFtPgeIPGyBLUnrFDzCbuzSQxCgRhYKVuJ+7GXe3ltqpndX
e/dFWaKPmIcGRINYnZEC6oYwhStQLBYck0ipBKIvgj/ESl+CP6/OK7pJTkPhDjFY1XdO7gqXbUjx
W/FOYVQM95CldPygtTRivxs5XZcqKTIChkEeb1Je6BqlWh1/XRpdZ3bsB+G1RPuSsuMO0pETwysB
Wcf+0dIiKih03skRYQd9/esbPGzcV3CLD2H2Fnb88GjT9pTQ2GROE9iGHFKEGfIkXXRdgmb+2ZZO
ezT84hadMkBnFAsdmhOUxvp5/5O1Q1iXz4pb210tTnlXB0ewuH2nXXIytYv7GaB/ALinbESNkdJf
uiEAsNxEVfTx4vZcIp+fuirQc5cytt//N24OCDgOUxhaKJs4q6ZvOefrlpz5L/mpi7zzFuXwkq0k
TI5f2aXlgQbK/W9oPF9DsMh8ypqHrhSq+2a4T7hu3HO6XYVrp0k0bd937ydvWqso/uKdMlcb1klJ
Pw7TLcShgr7bJY8lOHfntqbDciqU7ltbM2WsW1HIxN78260VwQRrWdmxoLqyYXtKjBwM2TYjsZvL
/HxtNxBto8n13s/KwR5qHOCaletkGfda9OtRFn0O5hnuohuVHZNhj6p2csAnOVAoRAKh8Bt1fOzx
Xs2uHVvORE2HFvt5kkzwERqo1WEdVW/1LIbku+UKnIWzsTKc3x90pd6RhQhwjOcxRP2WfJ+x+0BS
eVfz4Y29ql0TBVa8CzTmYGT2kHUClwHNzSNeOEQQFIqUHsSM9qRMzky5aghQrEubkfqmxbtE+H0Y
uhYfY5OWz/3QQtEDLxXi7/fhJ6KsHDBftYJgfMR6FeJ9e1B5+Nq6MfPgGvGKJAgZpwG3BFXMcKgC
taYEZxxfkhvnAgiS79n0xjxtIvXIrU1oAeV8s51C8yE2FmADI4OZLGa+PqXXnfuOm2cmtnxkLfCV
pDFN1Q1AwaoM9dO7otmkjGy2SVTav9AYzlZKYsKhP9cnN54E8vURtNZnp6zVaJ5+2ocW4tTdzmEd
5DAnobpWvd2GpxY3s2guQBrs4JPyeubU9OQEIOJSbxmlnKngGEeLCpdPnhS6b/O/uFe5f1THvH3d
nMrxKKsKkUNFH6bTHTC50G14Ja2UOf3tEj7dI7PxlnsrxA6r8U59U3w/3WJ+cCHd7zOEyycUoyKj
GCk0jlg846x4GHc2Zdmr1dgWILr1WEFcf6RBT0oi2+iO20aXIFFUgIPVyHN09S0C9ijqYR7K6VmT
8fEpgRZqzKusrToB4DgdCT59uAqPOl7X456+OC1kicj3OG0QS3Hn0Gje7wX7LngRPbldG/r91Fak
ub1aKYd52rUr7+bfWawV8VqVKZFeZzJ5GGS6vYvrCIgdRAsZuYV1/qQYJd+q/t8lJJujYHjOxH0q
cFO9uUg1nhfc9zoV3+xwtiULPcjPQogrRvhaZz9AzicxEluGLUva7v7bgbgNY1SQ444hLJqpRBQW
KgVWFe/EHFw/elgSiytQOkj6VELeXcbbvfus991KOeNZ0DScDzy58ZaqGa13fx5CrYALyd5MTato
j7EKEDdO9+Bdlz+WohCBM1C19lShh1U2rfUVTFVonwfzHtubcgaUvuXwi1N4aoLokt2AntIglxuZ
nCJNa1Qa9cJ4g1l1o21AEz+aL9kbivUQnSeQ1STgHJS5itt0XAU0aP3K1cZNqMwZejlTSp7Tig7H
AMLkJUwjwKSRXn16yk6ZANA64ZdeUa8p8al6tEpABVMKXeUL+XUNsSfn+jWurnHJXKhBKvnPNSWp
ETrjxYyaw12jxSF8PnHzwsgYW0ZRoZByVpMAqUiJmcphkx8eOrYRLWATqKbqddnSFg+exy4mEHUl
jZJVD6vfDRf2AvlA6eCrZdgpm4CFJHbiZiBBzu10pz+WFE5dF5+cVcnU80lthTRSHMjGkpG3kQep
C4RuxLdp1ILBNbqW9XDKtzSDpKrXvMftzYUBS4nalJvMDrlfI5vzZCE2Etd4atIuNpbsLDVcqqLe
LtYLKzOagDJoA9aDYOQVecym8ZjlGmHGzAPo8jV28WKTNxQjOnLJx96K5lfokOl8Y3ztrAOS/a0m
mSQ2N9OXKbawfUVRHpEPWXF3vjtVMcggdxPXC4a/tT1ZT1fO5azhqzsPfDUZte71n6lkM8xzMvZi
Rq9U2y4nhju9HluM3WCnQHJW8/+CeAzX2+vf4/CdfTTpvgOK3OMXFOfyl2JU24SUPQU+F3lI8o8F
VGjFvjqfpBtZ6a7jdLp/MUAUT+dStshVVni9EGAsfOGO7yOQNmK6BmpzLP4EzYX88K1ohHThmoS5
b8/HlEUJu0giBNuqyejSxrUHNfCOKnpw0sh+VK4gW+b46AUggVSPkUgKFTFx57trE6/SDG2OZqhy
lxwPmveXQh0FtYe7liv3Pr997/fDA6fF0GZMiGPh9FD4DWDEakLz3MpR2e8QNQ55CS0jwjROqUut
IhkLLqCGkfyoFFaWJGBSIRxunz+JZvxdB3GqevF+xnnXdmyWXzTtC1ZuU8pkPWKr3/K5CkkYgjSn
z1WHSElCxEykEAIcQL57PhhtWQ6jz+qRZM7B1V+j6RzZABp36BJqMW6D+N5WAjV7v2A1qSMJwg59
gZvaNPr4Zs4R9HWf2H1ORczCxR8KsEY8o7SKkL9FoC/M8EGzyw2z5MfOWpl5zFTd5yetsL4uIDAz
fMZ6Q2jaQ39wQAcx9hJ8mxM99oHaLYrBP1vciaNLl/R5aoUUYKw+S4YHIxh/6tCA99KuruIxoJOH
3+huSI0jUaFgSPVQ+MFoMKfEAiVXFVM6y64nsl07wmaW7wjQp31Kc4SoKtdyxVmWLOxcEjZyE2ru
KEz/94Rg0zAkM3yQoEEzRLMZJkqIXjc+Y4eE+/UFq0rxWnMc8uB/WXCVBJp3cf8gzk1/umCn68AX
zkTqCat81fPtcAwRPMslBvtUEfGXzKEquKOxpELa3WIgMj2znH0fTgWG2AHY+Od2oS6v2GQP2QNu
uijesaUgikd7FImbAGhBkcxmQYpP3gLitAdoJAcX+XXH03JEJr+Y6eok86M/rhe5YGefZxAYRXmp
rEejiPOS82dqqE9/RowW6RZQ20FHfO1C6BTQXZzojBbrt2qtLnEyCcVoIm0ToKofjEsCGw54gZv4
zQasBkDAqPEGEruOWnKEhoyQSXt9x3lXZEDfD46yWCYBLtKVdf2zyKFglpKIbepl/cPsPMFTyF7L
t70gf9tNDOr8ygHJ/aBNv8DAjYRHHQTMLt/HAy8swWrDTRV7yLTZOM7LTHUaPIekaeA+DQ6x9TNc
a0bmIs8Mx/6S4QeI/x/J2EjFZU+aCh3Z9MJAwaUgYNdU3sWMMKTNwU+/Bb2RIBnmEaFxczN6zr4A
XtnCZRR2mcDmnz6lgeA83hTyQS2905MWRV3VP0pz1PY2ntGgVuVq/q6vH1kAgB975yxiBzC/AVYc
WQ77BY+rtMf9mskenQvhcirCm+TR6/mnTnXo57s0mihlJ28nqHejq3yzAs6P8Nigj9uudHoNMrmP
jw6eK9s2M+ONNm9cGaj3aUpIwDb/C53iPRK/jQlOStU92WVbkT1yRcQAssoNeZjcTiCAwkbt97gC
oNGGNRAgt+Kpg/CyJNPHZIzlLOY5Wa5Ab6wPkPNaTOkcyNCIdx/5Id2ukk5PmcCY/215EteesqsY
LsC41Rxb07IROOdmmua3pbZ1u41j3cSXp3rnOgAXQEx6l9Gg02uGyPtPI1O6SYDJXFlO2rzVPLfK
ZMzBTPGmrgPEacbxfun6pUO3qSoQweXV85nD8LRXl0C5XsYmCH7BQyaq6I/X3Ye8TCN6abGhifxM
AZ9EdXWZrFbgFka0aIZtY+EHbqO5uXoj7/ePgLkZCAQyLgHoJV8AZcwWHkkghEfmgA6kBMeiRwvI
9cTrZDrRpakbQw5I+QNg7ZlAzt+7GcgwfQ2MNLcird7vQzOb/B5/2KU9rUzYYebez9WCngdNaTaM
OkzH4OQnzgmIcvw4MWHKLUbUQFNIs0LfKXgB7rQ6MZ3bkGW8XRsPYjkkoh4SEqyQaHjsIYRabl0+
EVv3L77l8kAAUyG7S51OHuQuU3jg5OPP3wzK/0sN8Jtt/pST3u19zTn2NCR9ZanjUxnYprcg3qt6
47CYu2DJ881PUq+O/qaHO8b6GtiIl8+ne8h4b0qR1T6AcHBPABDPHvPo548rB9E5XnZeCWQ9s3TH
rx4GS3dVmo0o7tNtArOdkbpvkmM7WFuawoZ4fikBtwtAbX9cXI6Cf5Q5epSNEatAMqYGmOM9B0CU
wy4bh3h+K7oD6YkYfo3Ya5WAPxyPooE1RTGk2nCuQhDEOjFUw9Yhq/zsE4OTi0ovnztaMiofQ012
yIVLC8Hale9Iew1U39e227GFdm3fqdnsYBW+3gdUoJGkt/5sXZetaI39OmOfq47qRnXgHUCiIvs5
zHJ93bBvY1m4LZL9pwct85+ZFOs/XTfxaKNHaGZHerlZp0lxYgrkwGb3K2CqA6ZljfgQ7QzHdWN0
L19x3eCQsmMnrSS4631RoBVagAKLdAnKUb68V0sRSrjzhNqfkefaz5xrWVFtkQDTbxmsNARS8ws7
WKpTv4NpUUG2wDF3rtPRqcnqntSAOzAxC7AHZ0Me/AD07zVjP138M99NC7VmlLazt5WshrzqrQjW
27P3Y3XIZ4CW/EGXs0+AglM5b/MkfvqqUhHgDRIKvE9v6jpTIhX9D1KcE731u8MdsuwESigD8qP7
y0LFe6rx06C9ObU9feU3ByBLKGfPEKhgECoODtMl3Q1c0I3KtedEJPrcVlZpxYctP5HjGZi0KXa2
qUkU1FM9ekHGDGGmbLXMUC1R/ghR1mCo9HTZszLD+cGCtkATmVM3FCVQnJtzvsHJc0ij8It3Ad23
6T2/kuC1mlBdW8KfSBFnOi/6ShvjS0jUBQtxz7heBxmfbx8Sal8spDc495LvxWNSvuiWUdJFMC0/
eP6cBO/CWd1rHoYBpY64yYFRheP2Uw38nOqGaAQI1Q5Wk90J5uZvaHP8X5g7+7aZIFpt+IhGGgum
xoSJeF+FbbZB5AgmmiaGwhNTLVhIXjkwvPSiOZ55xMBIv/H1Jb2eGHOKNOMoMJPabQyu+OuTqz5d
+9jw6jrKkKMCgU7aVBCwL3rZPywSPkTSS1H1wRhxJMY5ygd4dPe1S1cbvqIlKoquXcdGW1j5YReG
Cs2zp7istUdNBCdBkWkgp9om0E12ESY2HZweZsTYgxgFqIaXubwo255LaKBpOBmYWVJ05DstRWZ6
cXNWcoVMLNxg0QupXQSu4XFcbJONnTIutEvYkaH3hZF4/SAuQf/MCQNWNvgYV3PigdgCwq/OVVtD
JPVWWVDFqD+Bsg0GTw4+0Z+S7ceaqRQCyBAeK9k4eLQ8J0fcKHabZJHYysNegmoNeMM2Hk4OGSwO
XTmd7lXHmLj4tUo1WihQ/2TneqwCOax2Uwd6BXoOVy7LPxcyfGDPOnSHQ3tSJnuaH6jwN7z1cyl1
peDh+1w/53K9KJ2eqFVQL6b44wGvs8J/yQjLw/5fQ+NPNRQrDZG+CebmNjbVeEu6tU83brBl4a2A
F2c6TJe2OgScxEgS7IRJR6mv8WIW9R6ttaZZm7/aez6+fF0dytiW/400G8OoQUyRIRmE9dpNG5vt
4bm7kKa9or5T6W+VAuQU2/KBjNy/tVy+5qeYvlqfOuGhJcplPCMrJzeQvSilYMbDd3qEgkYRjrDy
WkxIU1E6g/HuSUVVqX994L5L6pOrgoG6blBIL84QHK7k0qfZB3vwHg04z1UnIjTkh0kIlXJLAEC2
Eh5Ca45jCpz5JTxAvsOzyUcq9FWRDyReZVd9k2CVFME9QhL1b5bUwqoM+TPf+eRGnmJQKBG9MBKC
1scq5cb5LwGvknci3TUC57rqHP3kAbclJ2MTf1khZVH0qpyaWkTB9S5KD4hJzBGPEk2GN0wOXdlj
yZ9CQdzyf0yzh7DNMPJhWd78IpJgbHR12KkRP2BsB63Ra8z4S9Rk80coGjAQbO59tF40av/viVvD
6Xe2sSptP6TMooJtvAQhAn55xiPg/Hqmevjs5E1kTuJfibf1AqELXhYbXdJYGNqlaMKBusxqdv8H
C+WOvUUpA8vIRkaBgfO+pYOy7rkKEoqaA8pSOAJhgQhQbkxKT7cTFku1cNH51MwDDIgYyTtuYhxK
GBEb9yPUc2QCOJoWTCoyFta/PUQQO3pMV/6x54ddQVguElV383gjW/iApaGWdQw6JWFHDJKMNjUo
DNJLMk2MOgcoBOJ8uiFOsw50uJWCXIIac6eBONAnLa/eihb21iZ0Lj3pcoY1bsQ+9Td9imnHW/uP
J2g+F+ENEIkk2jSqzHdSHBgOo0Uh486IorudYiKIvtWQHMrFzQk3fhu0GnrNpLTNnMtPy+exVWAz
gBXNBUyqk7WacJFQ/euH3kImXWcB1MuD/OPMCOmhvw2hvGbkz7Ttb86DTftmIOI2aZ0lOADcEgMv
elp/1BcFOmOIeIP+Z2Vf+yhG8UlasmF7aucnX9v/quVklU4bcP7rMv/iQgfeXub5szNHOO2gtxdG
T8lYnededUkVMfunsYWfldpS8xULV1SkvwxiNBEWcC0uANoekJNFXFPFYtekBB2Yildmhl69x0Tq
Jv2M2pUk5gd0xx1eAOOc7J9cs1h6KfgpShY6FDhMoolsO518gLwBzHJkmqE4TptFudQXKKYmdgVd
LjvhJj8Z1FhSpO9shzMjjfIIJA7uHocmWqCflYmBHbvzAVe6gdP3SUEx9jy4Inp86ql8YZ9ti33D
DKlSg5jGcqO2yJCemCl7gfwKDcWcOYgYxNfPElK0093t86LxmsQ00xiqxkZxxbwgsHqgccY8PYVT
NFoHpd5NydyuUDVorgu/WhUg+DftSF84/AoX2CEYl6x+lEE8WrNIr6dmYRsnLMEX980197r0gOS9
CIoDIYtVYaHxzIGSkFdI8tjj8eAaa9oA+w2HbelR8Mh54AnIutSIimiya5gSyVX1kxur74kebbjQ
KmRbEa4j9+H0qN3WqHmNoIAXdsZuOWlI+Gs/LNcXN1GaYGIRah25H5HydI5NimjgZ9uVZz+YhYxv
1mX7yHxS9UFaq+JqYrk1/ATDptXzji0AkaGUAKfcNFdWNVNl3GpcJP6luO3OT+mNLiqf2P8eMJof
eCwRsXJMokbUARYlYMU62DpxNIB+SUkwuqu4RY6/Q7tuE+aGBkDvdiZbnUGECXDylQyfeajNK4pJ
fWsWH4lt0AelZaiEtOE/B7WmGJpGeZC61yS6NgwFlmiU3pYfkoqwclNYVIEgRNc2/h+dyMARk525
7OxzGgWIeajzSToqzaJ226lzUS6hist/mh+El/8fsS4J0egH8KFCv+jh4p6RviK80wucKuai15gK
ZQUz1zonPDnJVJajkdzQ0oZkA3Xys+Dy48RAyPHLd7rTB/1M/4sWACDwgcfcuW1GToUtp0PG2zNi
A2uqcD7MU1yUiBi9BBCo1qqu8f+gkfAwUyeFfzgbikeLU+rR3j2GXa2Wy9QwiHoXACuPuAyRKK0z
kM2VYlviCEdrRMCoRea4nMQGg+X/ncuwZQ3iz01HPOIVAjVhp1tzMaxOj4UgO0yurEHaZ1/WqpgR
5egQpyU70qLHM3gVIoUafaDSZ8Wbf3Orm6282IHonWA6ymXxaX1zIAp2Rb54x1OaXbsC/OP16LX7
ZGTkH/id6BCRnZsyS6psj/Gk21+IVcL3aP9d1VKZh6ZSYMzJOgXQ6ywrzIm59GpOPeC5/ROoa+Gx
pmsvH788Vvntjuw7V4mp/0Gly03us+/M3BwT7aXcxVIR28kpWLfEsfvXg4a4BxBHdvd/Zh8HwVxs
R1NV7kZQPcz7sXGrv/QniJoCSG1pNlbsHRdUnDcUtdcvxsgz/Tr4rCr7pE7Nh3VHGX65/+WyoH/C
1PS4hTQlGkK6ZaayWxYhmHIJ0yzza7s0TJDxmn+9kqd9DehlJBdzkMTKxGpZ0ty2m6OsdjlrDT29
fma2vmXwG7RIqckeymAYsoIil926QZNAnR1k7Wnqz7C863zST9Dc8KvytUt+bZYcdHYwSohl+8In
wS967ZIUm/Jq4g/wPwz3ajoeHZUbgkueVv+u7XDDGB2wuEo2mIluKWMVseMXpvYBHolK2FNBBH7B
p/ruh1sgN6XpJMUC21Ivhio2iZYMnIKc7t5pvbFAYz7RFdl+daAAx7pN/PJ4O2u2JDJ/qMrQo3oP
1o/KUsMEhyPoUAmKgL5HKoZSxkMig9DeokhiYV0xy50DEZcWWDs164z+BYPFczUcwW5XCLt7Mvv8
OmGSI6mFkZZMLV38GbRoef5pL9Ufr+SaYZRHe/ksDn9XAUhk/NIMjVLTH6ez6NSFT5P/2P5EOXxD
DMUVltW4DHI7wwRAkCd4MWz57u2aKVdHL7d2sIwzKltunbhIFogUVzOKyBsVVdMtx5lMhkPua5Ir
1PJLo1nAiDHqNzLGXSY13jnj1Pov+/SSgPZzRloJOGWl5DYjzNCWN/wVDDSqWXx70Z2b1Wh9asRU
8GLrorHZTPxIHBjo4w==
`protect end_protected

