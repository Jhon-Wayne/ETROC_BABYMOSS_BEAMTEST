

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bx24XPMbQl0ZuYgzgnvmK2UJsn5v5rHRrHaBzymEsRVRAjuRN3xRCY+goyOwSGiaL5BZpex2sDSK
2sd0nljSnw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CSRfZVLMWm0HJLEB7NOFzWrGIhgXL0zMCnVPoqKjG5Ur0+RK898D8TnT1vzg0/m9z9AJo34CsLar
7ajBwWmQaStI2T7HakgiApYlcuC6de1XuIEH3rZRMj/RWcjpTLbgkrbMj7lCzKzQdvZHARVRsJHt
n6KxqqDLGxMs1/m4zV8=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YDR4T6HZUUPDmkJ3uEF/8DG9RH1KIm/Soi0XWVOdqKCDBSgk2PKH3QgKdeu/Ygc+E4sEfsdQ97ZX
ZNKLn57bC8vQMoMyVXHXP/gB1IkATHDtiORbiLIN6gz0rbLre/0AWJ4pnD6+ix+zJ2ZtVx7uSjJD
UeDwmSaYOZQhEg4QN3w=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b5TzJrebbTGq/pRucwAvmRYTRYSTXLJ31UHhj7qPdtWGaTRXaKbjtJHLK6r2fdEku+xRcQgb4iwR
VR2WDz2dfhkKseFS1Yxa2DFJTK597UszihjnkRHDocjQO3cUY+io6Cbq8kFDe4t/wEf721IVy63Z
z1z8RoAbpBZZGG1+seGG0kHDtkTe8wOMD9mRo2qsutfBPBsV5sK8/fmf9Y9E2sAlYwKjVvsGOjpr
dIS4pkfWNQ1UbQXn1WlPTe4wXcRDxSDWm2NMDLpVsB7PHxXe/ma6En4gcBeXFN40LqU3TWcyfbF4
Fgd267nviONJrvDRA6uaiECsHX40iXKsaxsGyQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LoXyfjLEjXF6IqzWN8H3K7nR07wwyqyXVISYV16h6KsboFmbDcRTEPo0gH2rwN+AX6fpfnjiQCDi
qZVj+jq+3Jpyaex4T6xZDGqASKvTFZ53Vog5975jRBzfQilhyEnt1jyw4Z0UhtEM8LILdgabJqA8
cXdC2MS8KixvDgzWP6ABnTAwC9pDqbLUIqs+coqVvcy1nM4qt9WlS3/X4SHWNrmKgZ5d/HUtKouY
9yGUMGTi2nl4U+Zd7UaI2yJjVCW8JLst+BTCam4lPyVXo4ebpoEbDK6tTwa5DlOxI45b/ZooNuYE
Rpmlrdz/peCtaLTTS4+P11HF/WIAxGHuvcXpOg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
splRKPjEH+uTzvqD2tjFWmYXGYcB4TmcJH8LhGT8ueKKhMoa+orNkr7mpiSfxGo4nOfb4ddB5A74
rXupMEGR44uXFXmGFms0uV3Mo+LAVOswYWiSib2qqWdsJAVPQV+uS8kwf1pFIhgSfyhJYccE2+LN
qen4ppn5nmwPuAnPwhqNoxWgV6I1SCeKHMvOOim/bGhWBFyFuI4F9GeL1p+BC2DYSvijB6DHJgjd
lmuMd4WuXe78W//Vv2jhHriZx5nGgRFuRWE3VBR/38AWtMEOOrO4ijdAV2GyHZrphPmDHXfSwU6z
9JSFgLsD3Pd9zxwPDkqCeFOIFV991nTMDEBaMg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4032)
`protect data_block
ZaAS219W6bcUidr2opI6O8Zw0EmE11FQM+eCJT4jozFYD85GpI0IY3/ZfOAvWVs7ZJb7GMAxibpb
cq5wvqFmp08K3Vk5xvnjZU4ahmBWRSnLACNcsXPON2eYNUqlYxRky7LphNNCvh+pLq7SsTz9QNZP
1i4c4HKEo/a177KbQ/aMvVtEXIT792huHoU7/Jc9g9JjHnBLE0qDyadtuMakwsixgzCde0Wv+SIx
ixN6K8tMy2SpHs4s1N2YqMjl5LZFnMhLm8wroz0ZSz9JWd55YvQ4AmFK1Omi6Ow6kxeUcxGlLJKU
i/+xfugXmH4DRlN5TLYWaxbFG+2l0m1nfEz3823E5KMxdSoxdStKVaqnlI6sXZZfy4d7RXCqFgR+
uc+Qi8A+yfGBFZ/yQF2C2eToOB2yYudRPVAIxMlGEZa4LcLDq9nrNjX0nxb0ZINO6Rehz94ji57w
CR9rqu5fPgutcU8x3Ww4L0ci6EuCd59h3XAI8oEhKmG+yLJyVXHnPH7SdEYTOgB/zFmOwhsbbHz8
rOmgYeOC3xzGS3lXoN61KEW3s8YiNinJbI2dkNE0urdGH0vFxquohYKGWiu/z9wohv+12VQialqJ
zf69wbp1+YkoUocTeApgvHMQuyqx+53TSvNSXrnZvtI8jUn6q9MED/pzi4PwEy/M67Oilmxcwg6r
Kb3WFnKKRGHfO9NUMsl0CVTIOtc4bRVpuyVSf7Bmcv+fEh2cgdjlDojrapaDxzV16MFKEzjkNAcy
AX1BjWJ13pM4rWy1b0PqHffQmwdLIPij3d8jVKRgJqj4eNaNB5iZsCXgyX/YzqfZcBfV3pzJ/5Zd
UjaZJ+8btdu5M9HguEHvyPMLjd5+jmQIq3tT7poCJ+zB9VGmj+D6jAhcPkj2bOsZIMRSGjqNBXSw
ZDAMV1fEUNlVRt14UbdstBXnwaNFkhRfQmZBtjAYFw/LvvKYK1tT9LydSAiIO7BFR6oJbmjd4wBj
n2Bp1TB1rwqAZEjJKiOLfCj2c8Y6YBIpgSGWsd6jKIYuNtZBs1p6/VxFZQSuWROSAppEMV8NLhyE
1GVFAYy9R2O9uU/kyKYOTI6QUjG+EK1lHo6iB4IjgExQi83mRZSK6nuY9f1+5SbVCsdaXfNG6CWl
XItzF9J6IvarOxxmec+SnlZngl7VLBVtFwBUkOQD0s/DAWSdF80gD2iHDYX+Rwlnr2CO+Ym6TSb1
s9JaUopBZgLxLGZVNS0UCez2zxWZmR9khY9eBq8sZu0d6ZRkhBj1/T3SM4Ykn4uHZw5c9q0c1bFT
vowYgT+ns4JfTepiAzyvag6DOE6Kw408O74UyjHt2Sq29fuIWKEq1+/DEIb2YACb/Bcsfgg00tgU
uJOlH6lk7BRBbM/DtBpzpDUd+fBh9dmfjGlH/ZLYbKFYpqmUvTCAfFeIh1MhkU09tfEDKpT1UZRV
3bnr6MNTmYb9MT+sQ2uIJLzM36+WUm4PcQFNQ3AB1kX6Za5V1bsn6NWrC0RA6GeKIKPPS/kM16Fk
Y5uWQpmXnmA5Ih611T8/6QfUQ6CufYnGzqlxVrcqbF2Sx5IpwnXTW3XJtNglptN5WcPk2JGvyylL
egaLJSykubQW4DBHFPgsJXpn+WhU899MWP4TRfURGR50b+R0apWvFW9FJf71KcRntAB9Ifz2y4Tm
aC79nZDvbTcJn8QPYMGbFSX3XY/sFFRRKxf9lcuFa5zZcKyQkShFk5tlMpGw2waSqOUmhFMvhhXx
HZYGMOpg6TtiBZWejTflxoJc1jXN+BkEc0OOAuIb0V7e8Y5N0QCuh+gMkBipre6lY0Gt5gBGnTTX
7qdO0ptcTr0Y3Jlk25SKrVr4U0LdlAXGhXR1vRh0UThwwHVl8NcZmRT4rtrshhsNkSblhxIIwDui
4cekviPo26s+H+/cg+FvkWr9T0Ac858RaeayVheljD5oscNEaOJK30tIYpnaxwrwDdca5FpgIjBT
q7En/KUxYnoKdCNxROMwIfW3Zg4M232t7Aa/1+No0MIw+WxG5ZZJCynr9zaFweK3rXjFDfGnhJ8k
7l2ulVwUDeH0CHEdUEQdexyQ/SawqjBMrdd6PlwkjwO94BdKrAol5pPZs4J/OuNTtZzSsu2XCf6k
xKSwdqqdDDh2tAHJQ82HQu9E99femDCAGMZxQWqqR1qoFevIWsXlevU1WKsc50d8CqJPiIFSUKY/
DLP38OHEF/r3e2SNfx7uS5rL1W8cgvuixJH3Ok8qcb85Eng5H1aEgPdYONhYt+0c4GV2quX8iahS
RUXxuJUykJhoz860SxhaVHoNopS8wPmLOjVp4RlYUUuwyyn5FxM2bCYFnIdaaRQTstDDFecpvidy
CnLlOOkfEkFBI5HjI1TwYnAdffBM+9qn0VtXSUVgGQaOnzWEVtaokKDqK/yGgkVfuMlkC9Cmw6Ak
Y3cv4BPBai8S4+MD5oP6ZuGVDfjtOv6FKPxPjr4TWgrXNHJ/t4QAwxwoMi4zGQI0O555mnkgZ+aJ
qSmX8W5J/jLPL/L6sQ3rBLaqwqqWFqGzF13mNKdj0QSjISWzUtK3CNuI4MuDqDLrs9uCgannZM8R
QBwGOlidqkqS2IL5afJIGJwNbEIP/mqLxaW7K2UiohcqBdgxillavH+B9p+dPPOzxId4x0Tbj+zv
YbAZpXx3JRu/A7vMVGLxZXD46rBgdjEoDGsye/xj3JoTZnGpT+Pdt6G+rAuVCWhwq6S1UKO/5h5O
pm+H3YmF/VVnphJfwys/Ek0sL1A1eOzkr1TLrm4sJKdNvWQn/INKHFyf0w5YT/etAh3xBjdf+Eg+
PgWktnwaThrOiL0QJoI++spwi4RFEej9nI9BP+WtfX3w/woaAztmaxdUxTV6DEKrSHYi4aEZMuiU
p9CgJgumOWOKWlvXWy/6JDh1Rp097NtCfg18t89mzif7cbS05NHcI6Hupyoc523LuPfX/UDTLALB
+ToVHQomWbEHH7Y6Ts0ifIhvMHxkG+GQyj7a6f/6Hrx9dLBVO6XdUoR0u0RXQ3CZi8PHhJb7tdVm
JosCsxUh2sfYVFOiYpP7I812T+SQ7UFbe61h1vKV/Q1sTO8xMx9BX1R5m0QCYfiC0BuyWi0vO16n
ikeR7PMIDZnLYUUYRAndf11enzII1S2+e1eiY60x62NCTi+uPsHfOb4T5c+cyLYDVPKVp9MFK6qt
faUgbFQEcj8VC+OB7wraOnzBTRebZttB5fUt8NPpbOPVKhrnyjwv933uvF8bfOGPRKseFZrOrveM
iquf16NloevZVUPCimBYc0naXEKtl5q41vRl36IRAAObB/eE7lx+InAJm4oBK8DQV5+DDal+Uk42
dtj7yt5fyD/+eMJKaqlTB+RPXNgndW7bPu6RVtZGzvciFD8Txod/TKxxgo9WV2htG1SNyZQGMrsb
aZQN4estNRyC1W2q2xnWkAX2aMIe4yIh+gmbkqpTa5+GucWsRcV9WYjK7PZ1AN9twlwqsNbeUtdO
C5uPkjs2Xu2wlydhQQ4N6sWDSOR24A7jUCbR08aR/7Eizzk4OBv5p2x+oaEIvIKERbV7bUGF/60o
d6cwc+cp9WJ94019C/Q8RLCh/CDRUmSMxeb0AVQsWukPNr/iFM2JKewNcrRiseIDZTim2yjX9Gqs
9bwmfWtfdmeYH5Ldc7OmBTAwZ/pUucTvSQZ+kosSEvC2S+p0DcrfiOCw+45lBvI/xuY/U/Th96Iv
yO2MHWwtzQI7+TlMWRM9yrrKiJH87lSddryIL8qp7smCduYYKEBTQDWfLrBPDvUrE1Mha+bCiH1o
JmLiBIJNDLNn8JWBGME0L2N052ej1rxDAMMkBktVASmSZFT5Qehuw5G1FPw9+fTu5sKgTSPQxgRb
iHGGmHnczFN/YGhqqlJkeYXt3CCeYFV9dbPczKgjWUM3A5Q/6SoOHxr2j4chcdRjPCKa6UnF/3K5
cgK00OgOOO8GBbyraUQ/TzpFrs/PtHCpsKcyAEPHlNf0CdTjjYHVSTnwWLwkQ/LEsodemgKP465y
bg77QeK6D3ho8i3VGdzExcrGJUBv5cRsLA6N9TbezFkIU2MAkYysB0fqp/vjCnmTchvNpR/N2SxC
jmvvm17ZfXCDMxI6ShQGPCzdQqZv0yv0NFUKJwzaqTmNBGrFgmw3OD8fIARurdtc0PTz35JiqZqV
ntWFe2aRvV00Ms1Dv8vfn9y8wFZQfGDZxlKcnlBI8Icyi0o1WsML8SvZ+UdUEb96ejCRJsPgzV2n
qih+Ha23XB8g/V3PWv8yLoZpjoO9Q1cjcJ0UYBsBJuhiOuFFF4hMDTt1mfl6jRNu209QVp1dl9f8
JSw8xbPGY+n+6QTWSGhQNB5VfSvk5XfHwJtZ0hIMwuiWCqZlpVRESdr/FrKf2V7F/BM7/0tBQksy
1ITLqbcg2Gc7CGv45+qswUtiZA8nVfkvTMK3pGXvNfwyJXthQoSlcaxWZHnsXZpjkS4qZOhJF5t5
251Kdu25vwpZ3ftIgcnidzmtSdx78NDNBbnY8sw+9raB6WIufW0Rg3VXef+HDAO5JUuQqQFbPi+W
GjuLAvSyneLOKIJCgRoujAY77AFEZurssMxufYdPediQpfGboGf2nJHxZ+34RpyD14SFlTj6Gmgi
dM1cfKgWKT3PcpSYnwZO/LNFakuHH1wLo86XNAuiej3caeaKWlVGIlMKeL8GCNznBkirOxcBXqHb
TKg4sKnyM4eKntgDQrL9LiqbKZ7vSvLw7PfTQqq4Cu5/sNbYL2f8drtnPHEdbWa+qS1MXe2Crsrs
3Pcu75ASuVwEdvLKfV759wflTs3Y/zFV7ZXabwhAhFiCdDx1SzbwuaZ2w26XGPABtHUzvD/Fa1o/
0Z7vsx6DCY3aigYnjKABV4TQ2b/dtgmBkq98PsnG6nZcLUpicFmFAO/17ydO7arZZJZadlVTdsMQ
OpiuuINpiFm3r2ztLYh2qgYe6keDeBjLDmZypYDI4UJC+7lAG0d7X/Ry0+Ylv/sWdJ52wbKsxO4H
1+FrW1DIIcv0VfMYGRKPmtF9o6yzhFwOLUaNyvsgsU8U2HHM2ulZjC2HM9Sfeu+ht2+HzZ/Jvu92
8R1EdNXstrP4Sgm66RbJhqT+j4trs/1deM/CfFG+WXIJqWzAoO3fNeCeFlbju9eoHdE2X6Lajloe
RLp/yQmDL1vfT0MvVnE/ZeAM6iDneF/TiEsFnnrA9KLWTliEE4bYIlkIbK8yBpyPekx5GBUkqDIG
+kvjN+vMljSInCzdf/STFaboM/PluI3VF5VyOL4llaTHILms+R98avG6Z6pL8rQq1DjuAqxuRayM
HmxUEn1m0AUjHVYK+JFwrlBFkfqtlTm+mMdftLmDWpjxIK9GcCI/0Ij8
`protect end_protected

