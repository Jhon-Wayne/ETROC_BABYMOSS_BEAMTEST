

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p7OtZBpltt/h9CD5IsJBmAQ+bQJxazkQVbRBjNJ7LWO+cgudo/XA7alKhPL+qAE8nYmt8n/nhFV7
1FHJnU9EmQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o0V8lbvMs2u7Pr48iEK+soyjigqgrrzx5HsGK4k7Ph8gI81XWNRtIljFPpaeGwucYu/H+gPVGgh4
LxNZUBJhgeC8kZr5P0UJ497gR4WHGLQSo0hvtVYHYDlrxnVk2S/+il/2gMAwvI5YF/lKiRUCJMb0
2mL6cpx+2git922rE9I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hIqrLT0Q92Qul/GeORaSvJHHAIqLk6EmPwtSD3Sw8K7TFMN/pzvjFhA6g78oxGwtYju17YRUOAPP
BxWjMZac0YPGSx1A1AySaj/jWf8/sND51mJS4hxixMPKgd+iJln4gROFDpToYNAZ0eBhqGsKoRPf
Exo4YtwLGOksTW6jkb5XyScrMy9eg1uc2W3HXgQfQg9hr9gpWWe4xqhKUCFXFb9eiIDe3eaUQ22t
Qgz9S0YooH+uhgkKhXgOsKoG8s8RO9q+oyyLd0ANkoAdDySOy1H2+qKDhuJHoo8oHgkWp+t8x1nO
sbVK5ZibMfLbKeRbGwFkFsj+EKfWfOy4ck2AmA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O+omGGx7WVLIBeJijOGvFCJZ1IO2vxCm1x3fAW3H6+gw883MkRTmRZO0ddVzk3pvzQaBPeJUDRsY
1XbF7OM1C/khYSkVv9TjyhihrgNNT2rgkTkWtfQNoOMnsmtYkK2fHBBMyNXzHPZRBh+2VgTZHxjv
olfJ+wvlLAdf8BqZKWo1gutmRCut9sBqwVpKtMbEKFGRBnt2pETIJcWkewW45hEmUxoPlXpgWrRg
sESpeoKuutTTWJor2paEV2RoktNIWs/+x82raY47L1AIZ3uy3vEVemolA7/fyBhQXHdXuWEXntN5
bzesBXIrWmoZpCMSf+IISz8dywoKgC/dpdCKGQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pc9IPtPXrLLm2VmqSrmdhsB2/sqloTepqxhS9rXzXINDRuCWOADiBYd/5aw6fJ/PtHP6hvfQmgPM
pe5Rbb9vXhfZlTdZe6IYAV6ajOneMnpE0SRKlyLpgkbpQbwWF8Ta9x699vjybNfWF62AYBS3D7DQ
b0t7dD7uNK3C2oBkpBFbB3y/rTrUlQxN4AZtlp8BUDmTdKIOwvLfH64R9omltAgRoa9eT5fKR+NB
hJulrR0XnMdnz4MTDv9F/TNStcRrNIf5MM0b3o9Lm2heOPvkpoBOr22fj5c2jTQHuYFT3gyiU8GP
rFykj34Hi9/EcnhfJs9E3mtp1Tszf4e89AyXHw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rp2qWT1ngiwszVInFfAgNDsqirvFBRH0fhGMVLdTcJjuZF6cagj0r5deSp/lHSGQXbQ6hn2NE/pT
sVS4xwCY2B03TkdpZqI4G+dZXB8686b5iwRUQ7S4WwcHb3WXRb4Df1OHJ6dgH8h0dIOxvwXXNlqh
PKzd3cQ77q4ZzFc8bvI=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JmHrUUSZT8PLNYfmwBtqUH6qJ1p97BdaA2q40RVMw79ZG2/5JMAd6P3xNNzdIISzZU+jzu0NYPxL
Z/zfPbolJrCwAck6UGljZ/OOpPHLUDGkBAu8BIP536kFNfmsl2/w8PHTByudSnwDI/YKiNqfsxGP
M6Sq3+TkXml3dJEoLhHWDNi1mL1f4wADZ5vEh09j4ryxXNWZ0T1vCwLDq6JQfC0fF5S+fWguWeoy
y4GDwuB3WNo6v4nkxnIBm5jk34GhklMVorbQQ90znGRfAejdTRlBiH1jH/CASbqnXiNzj4+1wJ6K
83Kv1+Hi6TU2vQtu3O5wYTXjTMpJrASuG6iNvA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
WX0PnnYbLPETw4Zld4S5rBXAmm8TEONJvi6KvKR5bsWQSZTgAG9KWwplTB/1hrBH90hh8bnp3ky/
Ajz1ueHsO+6x3VCdv2NocVeHs6MEOoP2fYDLsKPgP0kqSJhYDvwKldMAHRE+vS3VB8WYNqkpIWbp
bBta7xh+n+VPPr2wKIxmH6b6Cq57ayyq82IvbvAivhSu3xR4K+O2IdBjnxygS4pa9IsDcZTFHHim
qAJbiVtIW5FbDzA9fagz7FEZMsz9nyXi4cZE7c0Bcd1Es0LYleQM02l9gK5abBXK+JLiyoHAQVvL
NmY0KQmu4x3oKirYYKdISkers5zBYCoBs5/kOARbuOhhvenF2kd6uHHvYrTV8KrJ+2PleCra3Rxt
bDUnZO1jSxnRYZNgw5g24MKMWEfjk7IzFn5qUQ0HpucICCJn2YbN3tx1/niYLiK3q7lelSqoBO+Z
/GIY4hPH/5T8NG2+LMvAQs0Lr+rcFKwr3VHhzQzYpj52W2LQxwe2L6GQ2PPOvjSc9N32EIdv08SU
BmRo2nbWA7M6kTk5ZjUsxEQk1kMdOe/WEA0pE98YglkF19S47R5OdcLymwKgz3rxri85TYAT/q6T
rhH+je5K2gcbtjDpFLMSNk7M7vkuujq0g/z5d+nM7suA60CTGXfN2/TuvsyGCa+ruqVvFFcqHcAS
yyLmMo9QAgbj246A2VZENj99pRPJ/mp65ZdwaBq7W2iNo3izn8TCi742tjSbCDRxA1sY5Y1PzPff
oYz/XNFRhMhOa2/CKxbu7GTX/2ne49+rTfQxpI8nS51tickqlkH2Osbiqgghmr2TiuzvhyrG2kjG
QAsCO6yguUqAWWf58M+zWVYj9mQ8RAUtJ4qA0bmNNoyWDsXHPQ9dNQmBzYi/M7NDtiYuCyGT3kzD
wH9cQhQOz7FXIo/WF2QentqoQjkIgGAqSvYM+bV/jHMLT+o9o7luqpVOBuc8cyS2sbU0nWarfJxs
MbeKXL0T2R+ZZARbnSpWebvwCnOmVJM7DZLxQIKI3bzIWL1Y/GEokOHNKuoyO9xsoyQcG7Df2tJ7
EAR/yBA/aHDBNtJ7GeY5aytSmuApRq17Qi0F11YxrFQOmw/xG3Fm5dJFnsV4a8fZDQFUo5XfOcbc
dm3ekwg0KZ1jDSS42ih/2BjSlFCOgaiR2jQp1sOlETVrLmiU7WaRtu4wYdil8uiPHKDFCD3zmhHq
+NzUd8gZGM67364Xd+Ux8yxbiXYLkXvYUaWhAjJhmV5j9i1Omy0i8651Ix3xmOJNpahcwPkGlG8T
T0VGuRwRBM5sNRZIKURaCUZERPYCNnLw8d0PBFOS1lnV8aC2a+gA7tSj5wl++cKV4hqReDBrFGbs
Uwg5G5ThqgzJ0Q6o6T9KHHJO2O+n21OHkDopsL91Qm7UxgkHSqeZSzf0Nx06i9GkMy/1oDUwYhWS
2zBO5EgPCXbe5h9GKsHDEGNfzkjuoQ6KakYnJzI3JR3kork7qY8gMmsgClhXlUxgwQam6RCFWlSq
9WIHbbREpN4CJivCQGyKTjWsEnpztWXrP4KIHFCVuwYRoPuDmZEXhuZy9+chYtHLhrUSrgnIoEEX
zFP8r8HzKqKjRBU5ohSSUwnPsk7q/Lx0nbXa9P7Fcf95ol6N1WDiN/xVcxAcn+jXog1Px08aMaTw
LoclxWvhXT0KQOCvBPRbYvowly4qSPG88igXeLKcju81VyFggiuky222ZiS+MXjQlUvRInMn4L+0
KtW1LHIeA4Q4kJdA5K45SgPzs7WW5aPXfjMpJu8oIvz3lm0cOn18oOc1u0OADxq5fDA8z2l3ogl2
H0/dglRtLRnZGZh8zKut3qdyqL5jAueXeYpzB5DGwhlhJ0SU9bjOE6clG49DQveK68LqOxe3MJkT
VJR1Ek7eNzC+WshmL6KOWNS9xiOC5Ny3LF4+75uCAELwhHB1isQ1KuZOabwcIABjdQQqChzj+vyR
bc3hB9LTBABtkeCkRnu4rDpFXF5tqvWkef80zUgDXEltxM2KLq7n2fRVDQWOuTz4L+4HR3deIGbp
VxmvJJ/06b/LVnlkTIb3ibqwVLCEMnZ+Dc4o5Jr/oVV+i73nN/Egdl+s/CrafLGfHJQDOujQMyWG
EMveAAeajUM8BIJEr5kBWNY/nphemYtQOkVuNhUNrES7NrbmVrVhocbhEDcLCU2/wsPciUczqVMg
tPUExRUkjq1A8sepOheKP2kyL5Q0qb3d5+LdQMA59/Tolk7CkOPYUm9GF2kSyX8QNIFM6tcgVl6S
zR3clVht0V9xyLzuVqEZq6JpNKSIMKO3geoLeDgwkyUb4VzUocRZr1NApuuvqsqmdS+KgMY7Queq
m9ds+oPnUcCkjff7bHdsgSC8AWOrqv5zdrwGFnrNX0tnACjofGLKd+SoO7BZnGB7QeibED94SV3f
GaM2WxZNQZ7D/40dGJdE+soBL0Ta3JShEJkpJh0sECEBwiZmaRypPGYZA5bXVSZAfxE3pZ4mOjXL
OtaTDGhBZrd+hwLQ+5v+HzXI5tLy9pghCsgoNya9QK3aDePIsu8KPSqXAVyy/9AhFjNkTNjcZwng
rPJneiNQBM/8I62picMplhmvQ8AQz+8EnP/X/gC4qV7lGxlKhTmubjBVwVajwWw7Hgr/qhH4Ag0l
J3tbVUHYyB1L+srtSXlKmuF6SRVRxdg2uki8ZbQf8IrRLVhK2FbmYZovoqWXUEc59noCRdoknE+0
awHpKDaViHajwqOlMEKPgAzaHmEoZaFxrj82n5tZ6B5xMvHwitIdh3I8PaT6ebD828Lt3QxM/uOS
kwfAAamWFOvsX0Lbt7XwdZp3R+jg0Of1/0docYRmFxVmpUxTAExH/URaplpj6A/+tBUDYxsKVfLF
VS2oHCX/RMkAf110bx2wZudiOxaAwUztZgsZY7Purh8noAiPPVTyz8BfWoctOtKQGwQUlEmFXdt4
f0L8fTtZCeNdC4xxrv/iM/AaQX1mo4yNnSU7AkY9wwkQsGm/+HoQ/ZK5UMTTHFiSuRGf1CnLXG2Z
eI923u+QhDNLr1x3bTMJpBYcNqXNqDIxC8PbvmURI8X1jeERf1uF8AF6OwBnel0flEnEFy8Pqs6+
miH8znWv+dzrBTcso7b0PrVfV06aT7eXF9QjgPfUNERjl4kFzigvCOfbZh7BU8ATyvzmfXjRdjwm
fac9Xcwc8m7kL9P2BBytoyl9UVos5Hd5J/wbqy4dsRp11EEzV67Y3bYfsBN3hotRLGXzg7HK70PD
ApEz2CWqunILfleTPg37hTuoYNU+c/fTKpbc/JRY9Hhoo/2sh8LP8vvTvKO++L/Ah40WnpQy3iE5
yZCXx6voMzqBXgC6u7ZuWTN1cHQ5Av8jAabHqF4tjFHANC6cnNB66w+KeTPADNl0IbGXU5c18GMq
PmLVI2VVR30h1PQI5a8Ppzs8VM7obCehPM/jUCbSNso3fQbXWzeaTx8bYvivc3gQm3bLbTEeXBMj
FcTeg6C9RDPfw4Q0xB67V/WyFA2NDWP8bHeozgKLLoslD0YFxGICJ3snAAo9lHli8NAtgiTvpftN
wuGkIR7BslU1DNgE2euWdSzklsqD4b/6++V1iTHZpA9fz+GJoWMoeqVFNvgG5b68IpeogmbQeVAF
CBpEV3L4WHSf9C/v2JkRcGyk21D8l3DhaecVXd8fMzCBLvmQxEvYH0JolGz42dgLemdV/d3k6pvT
vuhwLPIWlfLch7vkH1QAET/2u402rtVFTxsf0jcin2dQuct08fz7d6SQtRleVQMf2LYYOLnZpcGP
eBbf7xS8e5i7NE/wZZm6gvBhX2yhlkE+TyEpq89wKL4DgdLS1jv19HqgElAKim3dU7B36z9ZNrGe
90maHQzi52R+87bbJF9FSG5k+Je3xczcaZ8arQRPO6Ma7nyulxFUm24sXf/hHmfZ7NT00Gf0uYVo
zaVQfHMQxMcQJshnzLhqYQCPTPCl5LQGOCjk4BIWWMnfSQTSqEcG21e5atPmWfl3xvdsX6GG4fla
P7SQm1lsMCsaZ727CuqJKfJlG8NBUJvU0AdoJhp5Rf6TesidYVhKgPyqwwY8zrJNQ9v4Ow7n0jsW
Llz8DKYzbLuMjAkVREAH+N+PtVb9M3iYwTJMzxJWuuAlWq7laSMSk+67mUkj+TRDi0LS6Xb3B0Vn
i9oW7eKWZJ/WoEMddYOM8g5LbD8C00ZNramnQJPoV8X3thZv90b4zT0EX84nO7YLjlXXA5LxmEto
uahWIiYDSN1Dg77+dB3vHCFuFuT8db72a9D9uXrlX5z+bOvGPFYZeUi/qntsoCUqd42vfMNRAg0t
n/mfWV06pGzNb5mm4eXEqh4+vdxbGvx25IPG5rx7B99/TwL5Fnt/3rkmluYblxB96PqSnJMUvMmf
iKwBHUG8k7MY0JjM7R1AgO9fN6ezix1v6dpBbINmID5Xzp2G36iW16NTa80BjMWHL2XRbO1ryuyr
lywzZVkP9BTAT92ixYfGROtZv6I6N/c+axU+tdcVu7DuuZIQ9kR8vU4jq6rw+af+PH3LNZ2bpWok
dp0CHrbmHCDhXY3V7iNX34ZH32MFcLVsRAcCnbpd7RrJn6rfC4Z7tnu/sSD09HblcjzX0JOxHjSZ
tedBXVX5gDsu8wujjmJb/OpEA3ueZhyE8sAv/xqZAJ54uVQ9ajA3tEDgMDK9rhhTxeDCo818nkwx
zyoHcQ1OnRmaLISPlbwz3BlxGqgLBxb+komz7vovAkQAWOuhywN3L8j1geBPvxmgSPjHpPQ+fj3o
lPE4XGEbu68ngnApGJ698Vad5aSpT6zM+W/aSmE8+cxo4t2Xtwfy0ZW7MfhEYCR8PqY/XDfdeWIY
LOzyLszLRaCKQC3JE7CBBtZ9qmpzV+8a+0BEH85TxIQWE3uWG5bNXRAzuUw/V7csjQJANBHe7PLj
ld/rM8csV5VZuCAS+6euaTP5+7b68ApziUiYTVXbAbtwm5oQWuGBlKMqzHivK0k7hcvG6RBkyCWk
nCRdEM8o/msSuFsaXZvilnfOjDfQ/J7qLdH1JrFNt4vZRGOSigRDAoMMfkCNiT9PHY+kSOWUEmQd
9ZcZ4Ai6oHwxbP+5bHZUhTzaNcDxlnU4sur1L2zjCOtBZAPWLu+7Mx5k7IhjTcldUyPksO8nqLWm
d9+ko/RPWJsAMhLrJBWpDuvdX4IKa7NQdbXy1lDaCTXOz83THbaZXp21MKz3bKS00pl1TA+9Gvps
LpZmYQ3wx2NRJWc5jmdBAxBpjVcR6gLTPymHgB41/qSHD1DUpsAAsG9ulbF6E/R9AZCbDgj8J6Fj
c5UoGLkL0KoqVEMOXxGtiz60zJen6PE8W6w3X9zr9GvkVXV12SPO8WG/aeZIqwIslkXVA4EGeZHE
xYk9uG9rW7dJehPBvdmAppJWetq9UkKyL9VOtXUsIxforx87rKdvG9C2/OpE/E0mE6qnrDi8gp5Q
z0GrpEV677B9ce38RCBxeqBIFeTHkMy35wT9pyFjr3EwamWhpzQImQtFl1Xjp8a8RmUnytme2cVP
RdnF6BqfE82PCxAdg4mrnRw0nCIuDK/w7suOUAfRQQ/o0bQ+ZQzkxdEld3JAk2vubwy+be5cWPCb
wZYJzX4Yla4+QGEjwNl27mnnVFlhsE9veOvodt3LxLoDXCZrLx0b61aOSHsQXfhDrLWWoYqd3wtl
g7IuawqfMv5siK4KD3Qe6OcEIzlnBfbNJe4pxcu62J8qHkQcDf8OIseZUI2cnkSCZoDs8PkJwPjT
/cxf4U/ECSxoPSNuZbQ84liETC2lWnJIWZkDCAe9issgubi/CD+0xB7gFv8PlmTKnWxyrLzL1lxI
ZyiZKhg+nxLn2X89s+EJa8OlNXIX7eGrXpwUl9m0nTkIdp7ObfomfF2v2KVc3k8lyvo1Ykv1tS2D
XNR9DCeIs6P35EzJagPLW1CVf9Nb7MGo6fgjCtLRaF3nfs3/GIUnWOLT8/sMtiQcKINw8+hDLHST
WYpJ+3fwCzg6E7kGycuCdMSKxDP2U1IHIrtmEiR4rTJfufQgD2LKG3ikv8LTbpg+8HIkdNP2mQOr
TehJg7uMbQiIDDE06vDewzebVbcZxJ7aj04pSq2i0mpffme0JBoGUCOma/Wp1oq3QGzWVj2MNIXa
pbxtbMig3cPgxYtAGFqxcQJ3g+5mR2T1c9IhflMLLMPxukBjDq6TwqAIitJIIasCVdouVZP1YFR7
J5AIRGDkc2BfIMCnBgjWX2CrZ5h3B8Mv13cXgJ+/kjVb+L2bOQsxj8VGJ2YUsWgdLrRQHnm3H/p6
F0+WgffC63FnrnVQK4AHSJGRj0Qhf9uHY5Hyfn+BdDFflC4sHNc/mNeIkOuMxQtQ01/ydwKoHpVY
DRI8JfytGUt2FeIbFCW9wmAY1iao81gfDraNtJqGiauZQutJkH7+KVJbHsDaGpEMzheU50tcLjkO
a9ujKR3JJ7wCDfhuiSrqQmxrf/hrXzc5Itde8nZAZhL+0MaJzc3RhegVNgiBPRbvFxvq0jCEo2SK
VYTZ6bkDLTDP7Ebs2oPHGA1/oYUfvvAUZ8pI9WSBOFuNoGPH9AzmBUCE/WQ6KhvYZaherZ0sfraw
cW8yUMUKGJs4MOE3/lciVXOL8VeQGxSuvfQw2adVBK1f1CAyzePdd71WcwPnaajZdp6YJNXSNj20
MnlZXVMrZmp3NpM40830ZNMCEy1LLg7JoFkDCvnSwciAfgpRb7TRQjYEdkG1BPHfFW39oH1RPr7V
+XfxjWBk9Z/Pbo8noxdoS/SNyiNHT4pEsKxMYaZunbBXG5fPXzLixplXB2KQz3Gm5+tcbF6zitCK
ENwwTeO/F+9MluZi2YutbUppWVx4SIMXlNsZ3P2UX7v49f5XSS1VPqTQPv3uXTL0LP9KIfbYjtgH
+FGVD7A7G1/oxIYqyYOpZA+gBaOmLuqLLikRthiqS60+pC31omm2nyvMWyKngBfZHOBn2YF9leC7
JLZVcLwRRrraoReakDPCQLQocMESw3iIDqXh7tXU/HL9EhO/pzJoLgj2SRZXs3Dksoqu8dx2I/4R
8W4ikfd97wL3aFKO+3m2EQYz6l6dwqRbZZ2lvIesBz5Zr4lO8IwtSo8L21NpLldEEryeOTkYmzco
itVchASoDdtIUXcmeaXzSYIX4mEr4cN/9DdDLmYZrz5sVVuwlK5AV+HzPOFycf7AOyi8qCY3jDEz
n336tBxJ9k6V+XxXSSeq+KFZszPbQhU6mtRRQB0cRzersw+SiNEfgiuH/QKHTJTiTKYBIOe13C42
a8a73OU3n7Vz6ZxDvzj+/GRzQOk7xERKqdE7n58q0D6NLs6q0yLzZsX8mCeZ5vDwcxOjCkYF7Cxl
RxvoJTCCFwvhsAAwLJfEGOV/HhlpIoemHP+cTYNmug9nqxrtXHkFxIbhHwKaB36hH6gt9lmzjX+Z
Fx7l+nMIM6I9QR3RveM8CrT69IdxjYSohwtbdLLer9iKmb6bYJd0xw92DGvPjSh57qxGOdz07Bzn
sq/PohfZzzzivo7DCTgosRxk6PgV1bwCasaxWbRgfriTySCg2ENukjTBo3OXWZGDYrKE3F5Oz1TT
mwHtzmSEjIGGAETLaCaNCseF15HNqkjNYbtiChZhi8ih8IAwCE6K6pj3FmYargtT//xfWSLrlvgw
r9RnomACWWXdGtc344nNnARoZpFPrZP+Vf9bScCx4qiqynfT0DA8P3QGO0+9Wu9N2qtQJrP6imUu
HZd9tsLM64VGwwCE/dB9BIngD1mZ7UBbfcLF1T1L6YYvKLp9y2SSfu9szImRBbD3hto/2KmDDdm7
+V6+EifLUHd+PedvN4dOVrw7z7Eknwe6nPElnBqGjY6BrR/Q2rD6TDdnnUmF6siKstKkyqeUMl+4
BEpO1chODbDM32xb658uFWkdSYov8GfcyEgVqN3xLJwkDaHa5IiyvbsfuUpJqERpOPqzcQjLXnlg
NuoFi7qkrPNFcHDumFe8TyB0ys0U7MBTbhKquOWFBqCl1q0GTvKWMOhWPZehgKxYgvNMRrSNwoqn
kcENs+WnSl3oryI5MicC8JGIsvsCWV1wZUoAYpKtai+duL+eShr4PxnqmsJginDndPU7uSoaSGJM
ZfWrpp8Kf19RrmmRKpjB+D1pYqgSEK1055E+WKX+5TYWwMm1d54ZHuPxQ8qtY/3HFpMavnnhl6ju
QgibYVUQOeZrR4jIk5GcLSXaQkP1pOLEDltVXWyIgCUrvBg4V3Z16r3UPqDW3Wul969aeRN2Q3Ox
geOMWD3venuhFZbtpY1gwWe7lccwNNDluQ2b6k+mLdiudY6/t0oDPXdrFwxbi2jwda5J6gu2NkfH
QOTXA95XjnTMaIOR6tVpeTdiFGjXmetV9yVqnvzVQxKT4MDYkQLk3UxwfiT6e/Bsfqe2DHs53laT
St/ER1pIqjFiaF417UO7Prqfrp1bL4TO9vlHmUn2dHDngp5sJ2U7pFfMCvtMeC32vhL2QK1kbFPK
zPKwd9Lj+8ZQ9bYX5px7YKZ4jTvdyZN4rxaZPOkEee9VXiQA+suKBmLVe2GxrDsON3qYmr3q1mrG
dsZwuWbj7iI+vTH/lSq2Szk8arpHcOibrNq4oBfDohgNsE7IPLYCs15eVjAjqyoT8EI/OVxNJYjJ
Wl4a4FuW8YYWKHS37+O4bdTiSnLjju1cEB2ICA1JNjgNBLerPMajZ4bs9HrS+ug++0oGlttj2Zm9
TjCUsuHrNb8OiM64aDM7sqTk5nxC7520pFV5edIRT9fGuYjNbLW+TdFi+q6u7BUKaxHXHy925Qam
7iQkelLYMelEdvV4YnCM56rzlxtU0ev+5JGgYlCvADpb6SUyJvMN5bTFKv41ZCBUc4ifazPA9rkp
d0JnjF2dVMO+55cvh+dsKbpGNWCiLQKTTtD5C6lzbewc0ToLN66FgweOMXd19kMRWFpB7q07x/AL
sizfHaHLT92PEjy8BnnnrTJws6u4jpRcniRuGGD2T1cUDDSRuj7HI91OyMabPozs2fOmGWJY3nf1
yJdYRcpPsbC+DvLtI+20OQ5mbcBZgPv4+UgUgAWPmT/DYlaCojj7XoiNK6vChDdIImFEhUxDN1mL
CIebnIMHql1dfrnFTKqNQstw0K+wUK8P+j12mW686TjaCrDDwi/6RQA7+0VgMGwSTEoliHMBm6dk
3xvjjO3TPaiZJRaWye2W2pTc7GxkLnpZbmYPh3SZHByDGzam3XCYxfQzfZXn8puZJLaPyZPMioxw
XltxnXD58ZbDzINPOe/5rQBXxhGzdxNf3/fTYohAZyNcCtDr+DLGATBSGmwMcuDKH0t7ZlN5hoTk
lsStI3hQvt18bnS8Z6rFA9TX9g+Oy3Rz6Jine8xqx+nR/zMv2i5/o5rwCHa2vkMp6UJXKJExYmvq
CKWfaN2dotaulGkz2VDEhrW66b7Sxsh2zC8b2w5b8OjR4DHOoLGJcC9tO+n5SDYd69Yu/O1X05k0
dz9Co302AU69cf+GO521eppfg6/qlT+kW21ZCloLDLn3RQMegwTPFsSBE9zFXPZoiS0L6bGlqVcS
D1EFCq6XQRSQHBIlArVxFaC3u82XBuNy6u+LfYucN9qBiW03sRd0lY1l9dbTICHFyjjghuy6u3F/
p92LUsd4ITP+B7INZBDhAZ6nodCdQBI7mIkNFBJjEv34dGgq6IWJtrBvBZ0YP+eSrejtsWyuHdt0
Wh3vm20658iryjJRjss+YjEkz8m4dvRjC3IFVNy7GftbdWvc/+FCgLOpMv1zyk8lV1jsnmMmzN68
f92JCAzk5fWhYmcnmSyCGYhC040BL0Kgr5UkthnJHIoE+Eq8A0pPpzekHaIFwerD33yOL66YhOuv
jnJbEMnOFP817pnIIaRq+ArDF7RvOMH6ntfUNwYLpIFaB6UFsdJ1BPpnyAelaetr8QzfuquMoWt6
XQ+qqONMp+Zx7b3UHlhzM7241xt6Jos0FNI+XHqqINYvLDhgpMeVuRj+cegwNLKhs9gir9jt0SnC
omuRF59v9rG+TU8V4kr99M0FR/uYyKl95YczAOzlzeH0JCr5B1Z1WVZh9tN8Hh/VIxQ3qYQyHvq6
3ljNKR5vxAyidiZZbCRRLoT863XPKnGnjD8g11Cem7YB9RIaVG/MnjI+yo/p1sdmuuXHQ1J7JFwy
N9LOHI9WZG+MxO4ml6Nlc9fgw1fX5C51op9M6YKxRQniIALCsirIP/a3rS7MPoZiSzZI5MSHKQle
qgWJKwM6HA0nLh457jMa3iGNyRHv80ZwLwoM4qNhSgdr5AnB8IjBLIQhONXzM2bdHaYgL6YRoxas
rpFBpme09DIgEWekJCtds8SyjCc0vEZCO0n9SXYKdIiPwO8m0NvtKyQlk13fKbGwt9P1xb1RZBCb
UfOaSbtOJK12Uk6VL2SRPWw2iy83r/uw/uuwUTKSXk0YrStCYorjeWnMsfP8OZtea5ZYoOvhKQQG
ANQ5iBNLk1Tkfhx5e5vNfV2fszObRiVyQGWW3nxidOopIJG5htGG0VGx1aeaSPuhC3vJt7VQDjCU
09knUH4CdgFibuHpGTaXY490GL9aO5HxoVRvJDC8lZgHrab2QaFGzUwFnj0NHysGOIoYFwFHXsJS
H2/X1pT3zm0YD1Y2EY5/wUQIC3ZCjnGkNW5SryVfUO6rrGjxBfEZk8+22RTzq0zGBZrKWC4hgY2D
3nrdDKZ0OvN5abQenVIyP9/GE56drBSlpdlmEEV50tlZLjnkBX+20nBDJHpDgMD55nEDGrtNt1IM
SpP13+IPwPKColzICHA6EXlfNV+NKRyDhZgfl4MaeYy0IktBwP9KPFWDE1Zkik7po5E7O1HaM0d6
LTpN6nQNnKYdS5c7JdQ4wZ4QlWScIanQo4r2grThL9E5/88ZySlQkx5/ah7+QE9US9yvjkuv6C4J
MHDyIs0Dwn0xiUjlrZ8orQjGXth/U6PzevVLUd1F3ayHfW7Aw+N1ywdC1LzuteGfID4Ppefm5quj
PGngcwEMqwoB+kMjE096D0zDwerTgpgc1CWY/tVkextgTkMEyvsBp1EygDZy3kJoGFQj4/Q4vMZ4
OFINcPqNgP7Trxy0ekyMUQ4+FOiEmkn0jCscylXRKsefJ+1gibBtm9YZEQkjgN3DSg9IPFvU9wjd
hyY5PfL3zGO4nC9pxOJH+FbGRy5yWBTlHSUjHNiW3drTbcquktP/wUlML+uE4zIaq8reeSc7FHQ2
a4hzc/u2MCPhXv2y+GuaCkExwODkoaPGrymB+UkONimfBhrrTA7fr1exRp15l+bo4xPfMeOq8+vt
IICqyFw+hBugCfu+2O4UKt5yv4w0FDsPusR1urihQ7w7h27/b9EUVJT1Cs4sPP0iX3GvvfX0l0iL
3iZsqLs+XHYXhqUezoTs7xX4abgK1IidLFQcBovnA3fUf5vc1Ge351L65UiREKPIcCGGpoZosSsh
qIT+njqR0W4BEM4bKZpm12WYrg3b+FQ6JsDeBXda5h1veeGttGo5A4u7ZUlTzP2zAU73AlNJpm6E
xKiFHTgsKBnhRJ6F1qYzGXtCRP/OrzQnFC4+srEreKGFg7FCx7Ig6U5zHrB9TWi/ane3t3MOpLQN
33A0RJyjitYZogukUKHHZYnbGlFQgjfKxA1jOlR++pg14NsmI7+eqwNfhTo6PPfqkMGDQJ0hO8h3
o/XUJOY1oCtkGwGM+1akIIKlJQE3GQxbzsILiEFmA31RTrQvDw4R+hRFfeRsU+IxPU/gUgC6kULR
vxuppr4opkjE61FFoLylthfkzp24OSY/ifqH0xjiwXxVOiNc/x5UNkjUKEwm3gu0BiKZUV7Wn7rp
1MA36JHR93avSo4C1O552QtPuPrpDCnTgQJvCN8RsqIuaPwFc/nO3rLHpH0OJGkx9MkCkQU4scWT
16B6qWpH95k+VkKYUW6RtlzwM569WvLPxMOG8v84E4auLhdDvgeSeytt7sUdrwLFL0CFZe89xy3/
7gDBeQY+yNplYOm3MnVyelISb8fdHbjKh/1Ct0HaaVRk8wVePshlbL4tiAHfezmKwYB9cVrpkOky
Vf37pTPh5/AIb//V9W2lAQUBjkwcLSelSYdEBdnxkq1bjT0eEmBhZfPi/Ik0IdLCH3EONa1SDCOD
m9qpqjZDM48+J9dDaoIHMBBM9BStuD17xCtuMpm718hYFGwli+AXZ/W0PqSyVdF8iyF5pqk6fvbe
nNzLaiIA0kso3ICnNezfxOEx1Wd17vBqMG6R0rSoOpo6NXHnFE2A1khg3fGnCrwb5jST2xo0mKYm
GPJ7H8pkEWNlwt7r6kOpHT7elaKWbydWNc1SgBi/Wvhs+lb7zmxZ0HjuixdVOYfTfkym2aYd0Vro
5UULZ7xFvpIkoa6dFCtRFqmz8GyJhQKNFIstN/2ZrgML80bumEkrHjpeZgiLaA2DBoaOeNoBGDNd
ciY08brAKRaaTkPwBna4O/AiFtLrtOcl76rTgEOUCviOiOS1CRdFQsyntBgCdDMFq/s+Mh+OPeNY
g57J/+tfjGhTQ8bg93e2RA7SQ+ItwS7hp5Vtrq5KPD5svtTBUODK7ntCNfdNaFBEXQUbX/Q50HRA
GfE8qT+W4HeH6f4a8jGpaq5/JoECjJYbW/yAZVFy+tyb1BjLfNFdZP0RXr9Yao1IESIs+XZbwxIh
nVXSvj7pKmFaMBxaumW8HHkDr8BarPpc5RtQrMIrMtQIFmWggID9dJt0IWxUkvBF606OjswiGXoU
BkFozC2Jd9MO04Ixr09wrJu6NxuMazeQbLnftiUtoMcIm8lLgNnMFYrydDhI+sJ2oGirWMKqIe/y
mTOZjFxTVlDDBatkzNxUOn4VfQiK/pVUTaBAUkhotftfrZk/4vVv4FABvNQTFf3L2DLnI1OWG2Oc
VGheXlFIdPcxLxciKgFXAcrqNx3+jfMJsCXCVqpNNgzB0HEk7Hem8wPEEh09+Xrj727eE3t7dgH7
NIvqGhAu155uCj0r/s1Sge7g4zWNPHaaVY2L84tKUsHzw/f0ex1FJxriFw/1dy+enLR8PrnuK9ve
hr4lYlOB5JSaA//Uv0gEDh3fvdERgpmi58mODCMH5oNPvmEmk3LMXuTziTwKJqxaaM8O/Mdql/6q
qnbUde1OtUHaTpFx8QQA8YL9tFntrmmAe2qA3yR1sdvMsrgIEc2eMK/f2T3pe2EB2cB7zyMPlEiT
h93dnp32MvadL9KOfpllbTyQ6kGBlccdOv0VkQ3fcloGKdEYnAVTjh41bEVAF3dh/mOG2drkBlJV
BtiW2Pnk4iu5yNqJ4oR+4DUp1MSmbdtbEc771XKxBKtk49lkYxa59KEMhXaj6hx9LdJbZioOf3Vr
Za0McbuV5C5QaB4juP0Oq+JrDYuQMUSEEyVs4OXFb9a1mleaMhJW37wfzdelHqMXaG73ikHcBWPZ
pVELcuIBQueAGBn44cJiyjbUcQCcO+B0405G5Nkh3XxtM5gcJFr+vM6X2fSMM01XVJxp9+tJLx7M
4q4iFtnV/wa8ZwA99FHuXX5X7NBhS8AGQZ5u+Y45cpViuVdEX9rq8xAZG2MVEpZjxCkCs1+oluPf
X0ld6AZuNdOjUdK3W11i2+5V5DzxxiZxMW3Hs28lXju6p0FVF5DeiB/JmfyL7tcenq2MwVI8LXwx
k+B8SuxSw+FkJ7LBLeTqf1v4AHPt9J2oh3yb2op9sUfo9V5eRd5QF7T0Csjma5GxRCFn4NXVpMRa
h3AjmhBA35jpnfp3luSjagXX+tMn+aRh8Ks6R7KjixwluD3ukuIljeoBWq+wGQm5UGhWk/gQ8G1A
h1W4Y4nWt5lfZ6LpJg7jdPu5YSEKgN3PglDjPZDxqV+rJ2lqk7KyVUswnqrI8MyYiETEhHK8Q7x7
J+evrYxIM2AFlMc9nDzGC3+rG+J/sCltGuAHBQ+SFVrK66Zfu4JsU+LTjRCpCooLboMU/QmSRayX
U9TC4LMwK3ER3ZjoWiiBPJk9Cx3H+OrrRFcJnoB3TR/WPIY4ILXe7rn5jBbaeXMX6A8MUdyIGtom
IDSsQm50L81C2vW2vVXmeJdquHSkGKwgi0OKOiH5ecwvVFY7rpvEvk0cxwDg/dTMjFwBqsf8af+h
HRmv2QznToNMPUZ009YJGbGv/HGICNgT0IrILHeP3V77lmiZ6euajliY2jd8N1l51hLOR+0ady2z
2bJ+Kw3tAcKO4PIhfk2AGyyWsW9JBAtRBpMLrlh6jFOgUc26AYyvyQY+qUv4g3J80HPWfhd1k+Mb
Zd/gBSJxFjtEpjJZ6aCr33bbrRVHiSnPLoZpqyMuyPvtZbxUBR4W7mbO21gB7ySvj7qS1x4/HXKT
dCsTasMZeRsUot5qI/pwGA54tTpr/5At14H9kMTO/rVlmBQlzWV5KZcN25bKkt2vhG4HyoP1aauf
XImN7yywwVaSFPwn1YUACfAb8PfGHVht4NHl/5CGblpZYPxP+qAGulL1mtKNKdBguelN51fWixD+
7IyYUps+vVVXsbmeeVXsszLC3rvcLdrecSQ8jq/ZdmaPnkbnOzXMgFpKpdS2XjyYI78/07EBwczw
pyLTUHhFQsIxDZbbkSH/t+wG2wzQ4qQRsORdmojv3RtZfz+b0MS6/dmNqbjbML9ScyZxlnnrsfAT
y1BCrwbXVINgp8UDWm1zeSSAENHigRYo834zypnB2KzNVMI5fiiqIzSlTD73sHA3ablXkDQUqVth
YyvnOqkcJIaywL8dE1+Za1wHV1wsvOooTeIMINuk2ryCIlURlUQAs144GZ6USb56caiUwZvFcFHs
QItk4vfLGD47IBebCOFzVxBa9aR9So5qaB0EwFHOystUpPTyFVZQUv3y0qMr+3lbo6pV+pof88Xy
2hy1EdANyAxA0fkqUJKaRKR+8ZXqiPUnOulYhWY39iN+3BHc14e/AFQoAPgc4Aw8NTWKuGhxvXd/
T067RsS0WZXPnstiTPmp8aLN2Qf6mnO9P2fho/8VwSD7JCkJQjezx8OrSHRiLLrly7ZSQiddWIhv
5ox3nmDURy5ismZPC2UxdtLnKPzUnTHY2eJRxZ8jTfC7qyf1Y/9ri3qB93TorAekgeL5H+4trt9L
68el4hV2ym0U23XmuhrI3amLVHM949nuL03gF4WCnqya/laMoS6lOZDaELLVk/Tll9wIUsfuoEPt
Nufigio0F0HpZLL+uF6Ll632Q4eFG3vGetLbbfHVxllNKFBF/R6tD0I2aH8h1Gg9wi/x8Kl/StZF
MSG0lmuJ7SiCC414xHUECTT+PMQTkxd8EWkPTKmFsGUAn79Tzvn8TN3q4uIGwE1FrrdU/8S86BvG
ym5y9IzzlsI4cTeqvvPRowJbHvVJnRoYiJMANuSc2S5wmtFuyjnMIaburkd3KjScNf+esXcxHHGV
zLhaLFgpqh07jKHkWi4JnCPgAONItu8x/ku7nvd8Pft1x1YkRcmI54Y0qw6tex99F8hGRiVRFbai
8BY/rDqpvn0eSTBrz/ZPYAxs9D4vURwj0jmJQbDt7bV9Fc6Ak3+M5d0A5cckUXZjZdHeBvmeCa3m
m7HcwauBsearPYnSgbPaNVCUHqEy4AUsOUPdbQlPsbcfftbn8kDXWl9bCNLhtQOccjqMcGhdyndG
9+/oL4Z5Mlp5kH/nNhCGLHCEtD6JcyW5Upx8oAoioxobIbqyAdX5y8D8GDcjbVMZQW2JnLejDDFi
hsl6F+rYgEAoASK6NOg66obujBg4/D+Kf4QOMhiEioNm16orbw2kzQhrM3GYch1BbVeaSvMAGBpo
UewQOu1a9ovqS4Dh9lWq6lPePpBLEOC48ZijDxSgH9A8mIDm2dPKvDxKtowJ92fTzCMnn3fkQM1R
5TDCWJOUOJGLirDJwyxVhdFU/qCaPz/BuA5Yw6p7Ajg3VIGU2z2k/Sz+sCHXJc03ZKK2eg8QEmCl
UVJoVXTsmSY7nrt8xNMaHmFm/Zjqfqs7SzLrueyuLQDlFFUwAj3IrUu6YWOPQn3eAh1yPLcIxKEM
/cFUfd8dxWGIoPy9JD5tq7eadCu9F4XE4WTAMR0lcfZ+6LQF8C65xq4pUqRDn7ZOiQ6QHl3FNGol
Kmilgayf0q/csoYLv0GnDe2GyY+WRBWUKlB8UI4CFfwKcmg52muKws9uzQhJAYH4ILbmvi08hTdt
UPthBil7ceFiCr+lPrZoDbs6a2aMmuJnlXLQsWR5iRuiNr4a0X+Yo+cMrux649clECAKsQhRu6j0
s8Xffe/dqrh9LiUzK2AzLvkyJcX9ox9+GN/M+wXlkrNXzOKkG1qCSuqZrUck+75EtV0dXRTdJgtA
xv1Ymsq61eXm17VQV1nrYyeMUTmjGtYguAW5tNw0KoK/hJNdGcggLlRjk+VSm21ChjUubKkXxdUD
ze4hQ6IAqcdl55WV363fYx36jzvFMU4In43zAWH6mcfR8/kj3WZ3Cnv4mHpogo3iJxQZ1Ksdr2gA
enAoD7WPgTwZCYn6nIvmdEc+VQq22Yqn3uOlYoCIK0DdNxrwZwmVCh7tOiFiiSQMXSXYr2XSL1Vf
/yc5vVDTzG1vsgOJtRTuoOvcvCZu1cOTQcnrMxpL09NmLQseVYy3wvAPeD4kakbUKi2nWgkrRKxY
G2FGHohK2A9iASTQqNEEvOEkYjP4n9vZ/YPOBBjo11yE1bcr7qxxWy58RGa0dBptjFC+OuKejNsm
lQ4XNxfqx/YGZW4tKOBuadmg15FbVNL0Ef9MYzp1w9eZ+jWLGXVbvawo7FThuQUXE2yAk8C/uV6I
K8EY++gOaSH+38M29gq2pjT+UIBK6yTIAcV91kYK7VAonAIPSEUz72rHvDcEAdeqp3o2Mi1jG5za
C80U51ZJoVtkH2kdvzcqdHgIGp09CALmSqBQ9LI8A1v6ujyrIMPE/gMlg4ciarbjqRCFmsftWV4p
cV0SLiWXDJoRjzKvR2sHOjw+F8c7mF1g2uCCOargmCANvsIuGS5yOfHWA1VxFBbIrqLB0nvhZtgW
Q3kJ2/j9EcPg5ySN+JeIM3dTuqKOS3TT5Fuvr1D16wDBQveZwL7unM0IfP2Au6EGO9TWhifYVzDZ
Ds4DOubF2bt44jAnfhL3Xsh1n5zmocd6zFeDrEDT1FQJtJCTqsktP6kepd1OzjmmT3EiOFRQ5zja
+6hJyqNYNAEPwLbU/YkfTHpNiU9K91z+lAi0l7n7bbhZSrZefe3nSSyY9yqkqBxiUNDettAy87fs
QmWr7dLJSI5PuJCKnagN7ATtGKOZr3kAlKTjG1w5t/8AkhquvlvUnsYAT9/RUnWKTtEkmBEKzowy
WyGsCUQbGnnvaI3X99VYg5peQIUyb7tyKRy4gAvmUndJArTE2ZcDXaq/ZJ3m+WISZTretMbAyuTP
UyCCOvSNEKPC7u2l/tXDnvlsWpHR2w2FsupWjniDKsPI/7LcR+IeHouI7260ZbLvK340Ttzo1Dge
sxZ8A9pNs3MyIgiFbdB/8ISbz6FjnxDUVOs1LwTOI4ZPJbdu62wpa9s65mnYCXLDBhjGze0HaBgE
KbF6ytTn0UfmeYICdJhdUNKkAzQ/nyqTXc4ZgeG2JrtYnkS843VNh2v6w40h1pHgg8hy6FuFA2Lh
NcLEmN4fdc1KrVKK24AL8gPHZ65BhF9V+FrrPqoWN9pvuU9Lo4gANk+Cnk7tl/c9imf6FF/+0Rnz
pzkmOsMgRnTCbqbCU6ICZcMMdWPEtIAaTDsgF03z8m2gYOSvOgziwLbV6hMAiOxM9BGuvjAN04dm
zp+wwV4+1Fy6o5CSYjC6SRqNLEWiK2exSOcirkm5hDZwnQ4v9p153dPD90yX/WpPG2yBfTtEMONf
jhV3xiZ2wWWTq2egYWthontNXHAfgslabrH4Bt50rGNPJdeyb14VSjX3KI1BG/UdV83mcdex2tD2
3ZijWUxBz7Yfd9OA8WJITAJG9UN/c4lQSpp0AjfrM3Of6EMskIsB/gjvipwVN4xSSwLtQPW3Rj+S
Q5F1wRP6fKkPW9GKd/j6L1+U6nigInV9eR9UXU2e8NC9zFq0VVJpOsmStDaORk2m303F80wf2+SG
Ic8yZ8nxCkkUOxUgdIjBTGXV5BTduh3qobnvusVwyH5HDy+stK1OS6uLGRu3DeZuOoSuxgAwfro0
o3i9NMQkLudfKzKkJANw3mts731CpEBsanty8KclU8usLMEjL0zatUD3IkCTvCFvp/6qxB/hsHO+
YX91cYA4gsgYg1wBH6OUY4W9p364VEgh98WATa0aDeM3jPXQcrveZqFbgufut+rj/G2iOyoSMXLh
nOjDqXNHO2ROc+4GkUS1rgaM1ujciCHQVmTJVsGHWsx7pRjJSmK00s3GoUAkkmQYgMyk2w4QkWvD
QqR36SYnQ4jRcmaRP20ATOLYt2dA14mZ4jbMtPByQVmWR23QVHHxn7dto7HMLdsyV9yNRTYDEYFC
ENDod2uHVnFjRW3EWWtNuFd3tYIc4wEW7FMqzID+FvjypKAay2so5odQe55hZ9xwh0kp1+815Zd1
Zu9Z7olyJ+rGiYH3wXopGAxLvqv0ngM4K/7nYu1vlvDNBdwQv22BpxbBPuQP4kYJXCQ+dlgQmu0u
M71ftmeyijMs1A7zPYdnKZ1NICjWlJraSfi8Dm2kPfiPwiFeRN2vFjH5mumXdQBo524O8NVbYWja
Zt7lpHSYk+sDNRabwOSCorEeH6+6Z1ZYtLTWyWtCZFdVlk3HiIToNkOMoNck+7RQ7OPT0BRzsmmT
Khj9wU/eW9xR8rEj0U5yqg60E9ajP9YOB2nba+bF1GKtP2pUmVSWFNaDm836C6RF44IcKquW/YfS
Ey71V2WlfG71VUAqmEOuc2LuCYgguCArrTwX07fmkB47wAcaFBkzx1xQASfeoWfq5nDoenEh2u5G
tBW80uMsh6ioOoUW43+dXoGHGBiyX7RUpndIogNzs8anO1D3AR4cyZG4o2AVJrEcCJstwqYC4Gmn
h8pT+yni0fOkrJ83pXj4dMz3FoJj0VJDwa5qthCa3dz/8A9jT0QzBW8YQqf7RmfZ8GSNnUTSRo5A
gTqxIdd3riLqSsR6h7p92y82hbpB+z26Xws9QIx2nwJMtwoGsBx5LFJV0XBJRrltBi1eXgfZbo/I
LFwvN434QL0VOYcHSSOZ921AZ9YFT6+YW+h2OUaTn+g38CHAv22h6VX29xVoYyaK/lT183Vm04X4
wB9B8m1lh7z7+o6iHDqiVSF0DaSmW0NKzix7RwJCTzlGYGttDJACl8ZuOu/kKSTMEkGxWZt4fh9j
iX+0gicMEpxhjhC6H/KZ9YclTOIandwLxl210zLfT64rhg4V/q6IrPkjrGhFra6rDQb6uYLVzNxy
5YPHa2FdN1kZDlZnrcpl/KTfbbIc4BvjJ4jYNyEYGTVFjCdiORBCW/FNxR+pBbUBIOf0GsCS5E1J
JPqfyW7yaQzL1Ug7e6I9hrmMSD3+C8dmgVvh0RJoCyEOz1+HYZgRxWLNiX0QXiI9m4tOKz6N387u
1cM/2ynVOggQ3UFHZj6QPFRkPbLeiuiTClu7wC3V70fbaxHnqJQF8MNuq68Xcg2WErjdRBucz7Hr
BkQF1qTxd2y0jZOXMr7KbqW8AeWL9s/ssy7tNrYLgEnKlQHs2ZgRZWob+06DvX3HydTw4MjD7gLr
yQCMw2V9leski6RnAnRg1xY4vSJInDpy5pRbrNFbiIF8BVSsSeKHdEoEwT41SzQ4dBy8t6vwI8Yi
HRiaLtoMTywh11NwQ+wmoTzICRPXgw1ZcQtKoohdzSlNbhSiRtNeotjjnirDD7p5mdUaWkFS6JY9
5wbPBX/wL+TfFxQpqcHWX3vWThAPTH9H/xkei1Do5T+b3iQT14ize072yUunpD5nXy4ZJtYRh9GM
/TXxGNWOBZmcO7X5Ok94kPmghgSFbX4OFwyyx+KmzM0gl/MYqFt+yDD5/uWl0Z6f1Ymlwc8D3L8I
gwZ42/b6nBmUJWUFt/zJy4Rv29b+MyoZzW6l+e2mk0Y5rsH++bXsU7Mn/Vth1TU8IVJBxOUnUViN
AxxfIpfR0/KEJqibAg5yVQ5VwMjzpcv6IhF5RzeP0QS/8ZW1/gAs7e4dWy56IXoTqNS+dkfCQbTc
9BJH9RNPxYpGbk9s/8hBlQyVL7zY3WjNbiS47XrXltBMjoJWi2CLfdma31eHgoyDLmDrOUKsBj6J
4vXZGDclLdqyqOF18gScZwqVOrECQWBAANhouWgZYam15J4HQhe3p0xjgIRs7i+0lfY9b7t27mX2
z0NI3S9Arnur0L5i4m+u49zLxDp/h05D+JKpKGKM5etXGVgrsggX5WwOgiE1eVLBIpJzXQXj0NCh
y7OKtowcwtvX5TrKzBQql5KrAvjr7HAoO+B1iDF+4bSpt+FmTJqSdpwZp6pWWgENSPgSLRaiIaTA
mA0wwJVj3+//gEEZU3R9+HIcDrZAiruRr16F1lVjBS6wqFHoWpx/xn2YybilERQOmfQp/EZ+6Mm5
w/tlZsG1zyDax7DJNJAoF4jTEfdqWPLs5rhGXjuYT+CtwbmWYuSbaQLQpnTuE/sz4jSjGwl3ztH2
8nQypei+0ROpFL1NQb9U+PipS0Tf6Hb3wtm7Jk1oT76fLuypi3ShA4kDdRoNNFTJrLP7999lcZ9X
HugO1c28dnKBxSZq725qBggY5/LocSLiTjYvEUCrG3Fxnuh3cNhB7IoKgFqsrBTbdRDc/esiLi25
zuInQ5MQIaJhrDkYOYMLsX4ef25KZ56Mjkx5zc4AoAfXwtntkOlD/cfwW1yTTjo6G+AqXVpQUfqW
NXR6z8lv0tXUm2X0Dq3xaotfpv38bYQyDI3Vv3RM5I79FmtdDUgQ+4pMHAUCjMpD6uUSS0/7LpHT
QvscUaJHwoaPFIyJQrFQia/Izga9SiCcCAcHrv7N0tqHQDYCtTjlYBJdbjXM4jAb/fQImf6WphUu
UUIo1zObz78v5n1rc9EWmFl5F3XhnjpoqLql8oW86X+Q2SRiPlFM/BSrhjbz0NxMSLaPqf7zPMza
WLcwrndZaSnVZTi5AFvncxYnoZZ/c3U3UDgNFvftjNPwP9fd1j973Vk9eZHyH/2lmzk0S8p1D008
MLIkiBQy8o+G/cLUCuNEOMvofAEyKF5ovlEOORTzcWQEJOssazTWX/LeP2bLaPr1ChynbeNOKZ8w
n8lBYp1C+LGf5uQjlcz02+7I75SpHesNIh/YKT7+IlzYi7Hf7/AYXYhGRwAs5APqBpo6C0AQPAH+
FisAVGWwr5RHLMfr98sbWxzKoWj+39fC2jGMGCN+qooXepN4jpVbs/zYTdNmNqCcJqo14Nu4vuUv
rbLhq3th+VyBM/HWSHDj/6H3WsJOYNfIDKcjav7kxQXlrzv/3acf6xUuOG7KxC38XzA3IhrF60/B
OgtTwDM3yildYBj+1dw7VQxVh29jx5ZJi3yKFxf/3MeJqXrFib7VJyGOqh34CpqOQtnm5Z1XFkoS
rPeiqtlAXVeJu6wMfbPRgU7LgRGDPBg1z18yk0334x73O97JcaWSyQyqJMTeUBa4YhpCsX9BW9Vd
8IMGvEtSbwTLd6vpRkKE+HkvjtIECZZrntAnOkSZcQzVDU8VjNfS4URbbsa5cD9XaajA1KSwqQyc
ylGDoVe3pYe234v4HNiczcqNnaVntHJeg6W4VlUTbguck0s7Z3sEBWdpiZ1UJnRrA7b7VM5v6ckQ
xJKnAzEzG9Wwhrle/LgoeO/S6RUGESuIfZmxBmkdsEHYg9KVaYhOJpe9FM5SUuiQmRSkoikDncxU
hqg0UYganIl/pvYnOQ4EWCFa+IF24M8JOY6QrpGC/WwwZ6SkCNxdNz4XJBusWrzJoxNEKAKPPaBr
eTkpC5GDiRMZIXOnP1VX8A/Q2I4QhcZ02vvdWdoi37AI+6QlEiBW06f+LoIetp1A8efSTA6C1D1a
fVAqWVgg3/AZlgvL8lHD6rJ6erjrs55ARxds8LEif34rZ/ogCZJm0ewnmMkdAsvY2YQcjojgrjO+
SaSWlEZhqd9sWdUIVtuVb8bDKvw9OJqyUMfWvM+OGG3hNtHiXU4GnFtGXizlTGvqvrnibR19yD5z
YV4z8eMbsmg8omhD9ACUp2/D+sbsXH456G32/Trjv8W65TwhPx+p21V5JTE3R5+n1kA83bqL0ZAF
mGA+YltZG8t760mHTFoKd6iznVjth1shH+GV6yXe8F9sKw1RsQURj36NI7h9HDf3N9tOaTGkKnaH
Sml6EAHtYcpC1tItwyHWWkh27tAEhF0hGhxl86cBaI5UWxnaVBB8+srizJVaC0uZW+EVle3LU8jR
7jKh8WFKLsxriE8XyWbFCyndUimwRjp0XLZGBOmAdxajRdvE5z65nPcQBxf4MGGrBNFvSJ/ZCN2I
KTCvQRmyciawk55x5ZGUwAKiwErVN3NuAc232RrTG80YOQzbwF5I3wu6QPao7CnZRaKesYM9y0HL
L/OTqdoWi7Dmws/s9Ub1nuPJwUpJKhAIa0VQETzREIAeRgwaL76aachZt+C5tVe5Tajcoq0lrlFD
XJH3AHkgpnfu+V6QJ6DuBCjKrAoub7GThgBF/qvgLiwVStLiyMAWA27hF/nVxtqnP2SfcWpwQUL7
w2VOKdGgJts0NThze4Bo+SG68Eqjh3qZ/Ay7kCGsoXBOW2PvAcJ8u0OPci6tbLCUaPbt6quvgzRO
Momak4S/Aj5fiRmNTKiBY2qyBBDA0BR4IUR3HlmM+gf/+c8i8DR94TTib/0xdHXqcpvV2PAXQxy5
pkvlshKauVPcXwXH8cfZzMJaLlQVLSgCLAqWzSZI/71ZbMrQIt02iuffoaSKkyLO4M1bWKzLHeiU
H+gkBEBcSduGD+DsbhwwEMRSeTlf4HuDFGZrZTAzRQA7DH4RdspyD+Wn+fROUYsjb3rhIka5vRqK
yfwvqQz3rYRvJKV9om+nlDjeb+pZiEwsqwHmbtsuHwKznuNWQ+0QhH3JQKf4FA74EAfewFi1Rt98
hb5gKJUWjOkSe21Q8wJvyEgGL+zhLu8KvWc67W3IgphoqXIM6nAYuTP0ylRDMgNflIb96ckRm/x4
bkFoxYhBBzIgj3L350ak1HUcWicSXj3dLggXC+hOJEyU6nE2mYo220lpDzX2mMcjcG4eyn+oTu7O
grg2rDTnRO8CGYhzmr5OMrJ5JB+OOz9LMVMvR3Tu6tW71AF+BjcWldkB6Xjr91Zr0Alh6B9hnTeU
s72ABtpmKpWdeXRWChcg1Ve2z9m8dxcV4rNOrN/1rfYDNkxfKK9/g0B/yLdJV8xoc4eCP5u4zzhq
Qco/BaLQ78k8sxtNSOAs0HyF3HGvg69uVWNTkxTO/hYmogQpdD/jdFZ21II00bGKYbrW5WmlTNBq
9RNXCDUf74iX84Dg9zoaGFZdquKUNEkOccP3unk3s7ACs52t7ravEo5oLOrctxb9rZiFUZxv0+Qc
Mdon8fqG525a1f9Byydu0HY0yNQ7fZVxXk8DF0EN0oy4I+31p+R+xaPIRcYayqd/QNuG6h2FMxEd
zwHkRZ5aF8NjgrOcPux6HHDqgIhCOzl3GCu/1J3OSHau3/7JQpK2SeyZjVA0vLmo4PhLFiohICrX
P7zLSuwyBP38QtJy3glv7Z1SP2QkCwI8SfFrvVO3zjkMkkOuzqKK9+j/QR5YdSmanvyASdezs6dG
tVRbB+mrOIDHhHXulyPsJKZIdvVe5fOxb06zYgJ7HLMBEjQhNnTcuZEt0BesDLrpvRETsRGN5Ykt
T7A/fHjf82lnX5g5WSaPJLUSM3CN+6H9EOGTVMDyxlvOy1gN0rNBHFOXafq6EdDyt45pq29fgw14
15v+WZjiThbMhFRbp7ACg7Oc8vMDIwX8ZyBcPiUtvFXfNpR4pbRe53pSCLbiEDT6ph8it/o9dOmH
mlE15nM+aZ0+XTrKVU5Z0JvkdHkhxUC8+1c4jvUylGThwvdPOaUBnb3qdLKrAVzn+pTlzIQFEXXo
A13KYEPt86HlJ1Dd1nJliuZwq6YGbfEuMT84yNelWV5BgFV7M26R81yFN125IMz3rfYRHWwAVeu0
cN7yACC7GoxolPpKyBaN0MIP2x5fdXRS/+Rrhu+PkR/0avVYYBWWuX2f7u8U/ZiqkBCKEXJVbtHC
QgAWSDHDqWQyT+kM5zo7ypz+cF5CRl/Z8ID6UnBqIdaoBRPa3vEWar72BnvwNPFnu2h9Hib7l70I
A4YvXDHdQP1qcjPwWkiug5MyvJ7Qhp3E1ZlDdlge4NM/kSdvUUcxIvOUbAVsqIZCf220D+k/+5Xb
QHRhVGI7+9HsG9/z+cw2kw18GDZ3TqIW2Q27HruoMqdG9Vb/eCZAI0yi3gdAE/Sec07xq6WfUYgh
9kwe//eIvCyFggDGwDVsLmrfDa8M6GlnU1ybkFhOZ/WCtCPubegNc61pT83ItpVFM7AiLLQdhqWH
Xw5Pu5sw9AG+ctOBK9qgS39YUdTKjH9tIbFmSaNL8H9+iJOjlcH8oL4Oo6wR6+3NFgjHmy9OAHST
BfPhwCsGcWF7G/bs3lgy/BnbwiEvaYiCRG0KpPN9uzHPIb9ACD4g/qlxQzjOupgeYJ5nLIDCkcpA
h7xIzWN1pMhbo90leGoSFk55TgETWMVXP4PF6nysGrdy3tdxfJP89GlLl+eoFWPblKc49ahq8UDa
OJWVEI2exq5mLRcEyfBwUvcNoKoAOXZ8VfAK/5PAuiuPe/LAJMjod9tYFJvcRLKisiJa0KoYfraD
Q9lyR75nR+0kmxYvDfdpcethB7RsR6OW0ucaJrACqLaI5//1KwI2eQ48q9LQSJRceL9exdrkUsnC
oPPBDNn8ZQYcuXCIExwFcliepPcX6C5EEvHCepBc/YdTKjdlKFyJOEd8lVyJDKUmQwxueu50i7UM
X7ydFLsJtwkmhliie1JALPaS3Rk72TMXMXSREq1VSdBMNpqrda77BqD/j7LmJodndtEnYaIfSWdr
h10kuXJv7lpRAkCC3c9C8uy07Wv6Yz1AbI8PPmO3g1a8e3FTb3IEBOX2OJCGY/rwYhaQnobhLkR0
MKIkdeDnaWjjxND2lA4I5MkS9XXnyOehIvxVj94RXVeZYIX5lNGJl1HHBncID1Sy4Iur7CTdQ6AP
7UhUtQECHBpReB3DrcTHXigjejgzAF4/YE7gyoeqmkG8aYkWg9xu/AJ/H37AS6SmhHJ6VmvtuK6S
/avOms7yfQwINUePL6ESLcrLe+Iv2UOqYfjrkAHmb1HDIvkOWVW+AMvyuDQVWifEW4kxXUJKu3CK
NRftKCtgTNm2gi5mJqrxQKTaw548DWyiniEGkodhxX9+SS8VchRCQNvgiwqJHSUI4xA/ZonHfqOd
XFcD2JqTvYrZqtAFhV+OkRlEHyhcqAbx2QkDUmY/V+bNm6GxpH01xM/QysD4enoczT6ykW3jp7ag
fQC2Cy7nePqnIWx4P3+mm0JupzAtcb7rVCm2vFVGyzMS4TgrIdtXixsEmw2Bsu2kMy7NwSxDhM74
5E7hzuubVvPYKtCo6ZsoONiIesz4X+LnWRGUN7FAOqTOk7wWJZ0rrDPl5+6xs+v01AhNax2wRDMC
8J6x7UbpxXxqnVtS/hkWA2dWsiuxg5oCk25ozphjIUWzgzr0c8HlFat7NrpiP4bRrqHI4B4uCQUf
2zOt7T4IKPFvedAPCjWvXIDiYwLgokZZwQZ09Xuxvf/o8bbRsZjYCLZgY6M1R3l4mRmZjhJ+1HjS
QxgFk6NyWEMdQKqcTjV0KbXT3wbjgpTi1S1TieGXZkgw5k2N33xQEKO71T0d/HXuumPZjd/thYmq
meQNlfp1UtvDI9y9/AblcW5ik+C6aeYXdDPlyTSo5X0UMbVCzVNhkI7Hu9JbV8i1u03dIGjlIu9Z
hh41PpSb5b5gL8Mv28WMp7UtK+AJIzQRn9gAQxgDtCbc0XPnhQud7yI4T7Brftneh70oPr3Rcf0Z
pOeDeN4JCIFGHH1OyDPxjxlXnVWzdqkK1ZJEdr2qdDQC/GJANMOYD4ZZNFHjv8mK2Gb/K4f0Dzgi
cU+3jxLNMf8vQa/BOAmhlKMWCD9QPL7NXFgFc/PyjMT7DjrjphQEprRgtrZFAciAtGohdcW/x0DH
2l+WfXuLVmN9j6XYconl1bOuUMfYeknmJNP6bFtlnUkbcqqmixZ9Hyq4anzbO+mBM6D+CKzqKLSK
iTWxyK9PvktN9Yojc2/yVLIv74Tg/ZFODvtRcLYgblSNqKZXkLxZ7iPE0rF9mBszQSl132jaDoj+
i5ZnTydtRuM/6hNBsG0YSkK7MSExwLjGBYolHikZYJ6DdXmYhx6iGEp6w7wEou7B5J/eARjWKM/I
mtsj3p/lTRTetWIGbeb06L+iflCyp2tuY5id2Yv/mT4ooAXWnpLYV7RQjhB2KPyz+FJHezjGSjEf
PJGMq+ylr8xLa+Z5PMuAj1YePoaPm3XxpKZp+4uFgxNVZu6ekONcEO67VJPRGhjZtJZ+r0Tn7w0v
kmUfGPE92qr2qWpnNhJ6OggA4btCZBLjJGEq+qoF7vWEp7higZ0dxrO72Hfnn6fVtWfKC4euC6TT
+6DRfveItOZsf0lqXwWKrinUzKttJdIF8TlDLP9TccvpqVH8euANGjSr411yi3UsZVrkikPfTk6i
LWAm8u1t2nye7VGfQ9Vh5aiyXfiyZNPsogk2sRRHKswOZStmwlaQ/WJzCcnr44O9FOhUtYQibkeR
Ko6HH4Em5Eeb6sZmoQ1QON8llOo9mMBmfJawAqij73bFvscGnoeSMsqQWRJT9W+6qbHdq0mg8CLI
kXSXA/LkCQ==
`protect end_protected

