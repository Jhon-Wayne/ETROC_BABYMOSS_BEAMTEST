

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oYYUZ0MeKqJUJoI7DJiuvSB+q5Ix+Iwj9N3EwG3d9aznfrZuw1+Fc2PVy4cVNiksbh9EhD023m7N
/1rZI7UBsA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BmgMGlUziZwp4Aeom40PM0gFb+Lk4HIg7NJ8Ke6/iR/nzJgqwxvBOYZHlsOO/Hp8XOgAeNb9Zd4o
mPFcvStSgKrLqxBJrTC4jOtTOOUVOGECik9X7RElVDiKeZuCTuuYfKks1rnTANMNKsXOPeJj6Svr
YyXA9D2NRP6YkUNuPRY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1jtnTjcMZBAylJ3gewlkrSdkM4rrC/SF7w+2Gpl8C9SK/D8Tzq+D0qrZVMnmX2MWMKbqqYu6bkIj
sy7Xox+kttnLUyhBRsrBNs6gr3T0xsxsJ7Gnyco/P3Bde80gstdJ+PNfjg9uJOXa0R4ym9WtfNGf
swawtPDRNO3XB4oPqX/YBORxc12Z2+Xzlc5kJQDf1WM1UoKUm0j7+JBzjmig2WrmokL853BM29jT
4Ht91JL1B2bOy9A+fEpZnVLxL5NzuQ9svrSJluHfL94vaMxePXlPq6InH4B+XQp0TAFlIitjElNz
4mBAF7U6zb9GPz8ite7f9+Ofg2sCbTc7qhRaHA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gQeqr96ZiBT2MmGHCpbhB9Ma/ONapmaS0FJH16GFlg7E/VRDUjqbqiiC9oovpVsOBnNDQZNmXNgv
dI/YoLxA/mPd3NXizDTj33SvvwJdHC+sPFJrC6pT5rNUHqY3WkLW4EktYj3xtwACazlM0R3H+N1W
ZL2jtTv4hCIZZw83DISHIwGMevxP0unAXWFpAlJTyOmzC5wsjnlwvjA6I18++KC1ECVIFCC+grSL
XEAA1xdZCU131f12m2UaGi1yGaQH3scoEe37TXsoGUkWCMAn3jD7PddNt1X5zhoSRxPsOfUDmtSO
kCNVtrnPznMY8kVS/SdMToJlnwH2sKbHJZ6YoQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aYbz66wynlNa4RYsWnE11uoqAUkMOGD1rK3oC0qHnHAmOdMhPdz4cV/CAQENwbN3ryQY7/k4qEBR
2l3bOqYxA0+CBRl+jt8CXXxWU8WE2qwf32lPVes4/pVAbKANmE02/Ysj4IR7MGLvUvtr934XOsBK
cCc/KqvEbWgnnzkEdl16nzyz9Je6iY7Ni836+/z9BA/OYPszoNI5lKgO/06ni9esrcL9aCuvKXjM
Vplsu70i86fjOGURYjM2YFmCk8Xng1M6ROF+0KD+TufNMvK1W5if6MPJr/BsB83OF/hzcDKyULpB
p2+Eliq8StuhC0n7jUXEo6ZGATEY2a8DWEYVhQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B8e2xR5DNyjb6SEEOPCOnfB9/yUC8O8izWpzVz5s4/hfcHkvr1SHS13gqMQDj1DN3uSpaoGxcSIv
a3uLHDL4nIDztAAEPOvl5rp/eCLKhGUauWJKGzgIaInIPCBXw0hsptiyzlIicQEO3rsxoS+LR4e9
ltN4asLfvR5i5+Aru5E=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o08P3wLx4KXr1Q02DiaLH2vPxf0H1jXIwF3rbwsiMxYgYGWIJGF4/mxUFC7J/WeIjcsQFoTUns3o
ZlNZWWRR36HJ1r2GmZoMunV8HAWjNjCUrk6RBWvB/4dYllizQVzRhb+3YUjmiSEMr4rkGsWsR9/t
W+i6luLQskwMDbMnn7puINFUehSDaOzDytgvFigNs9cj7haJi7XjPeMPUBa/JbbTJGFnxz8xzl03
55+BSHF5m9JHUn2eN7uDkExSgYolpcYI1EQnoCH8U6Zfcweg7A+n5SfklkTKUeWInYHoz9tHbIHA
y9aJwNoT7f6uxEt4GVf7oKjEfFlxUe/yajXHuw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 132672)
`protect data_block
ZDNsgBdDfmUioy/EdAAAAITFDXD8FZPyCGfM6polUQd9bZ1PCg900V6a0BLCTH9qk+zf63OqZ51v
iwgTeOOLLFhjjppTCHfRM1DhvA5BrC1WP0uZcUZUgoeQTLbl+gQ+AUelUTS5gMpwgYRPaNRxN1ae
AdSmBq+ewZLD5eVC/txMylBHn8Ko0c+FHMc0eilosaWoUiKJdDwVFf5vH5ageN8Uf6F1RBp0pLGL
VgtQtJzBL15okOj4cWMEnq+o9t0inXW06D2PjXuyxY13FJxKhwJ9xSSJlZ/u7Yaz3q2LrClXOM+P
oZ9027lKumW+J/8ZJrmQe72OxLqXfQMk7/PMU/3sbvqgodGO8LDjBzSzuwg8h36gx13NIOz09L0M
1J81Jtsgz/GrSlIoxahWy58YUiIT4ud3J4dmVwlIyCNI/h6m/x1DQb+TAnQJUDV+YEjMKdjNnlc0
zyuxj16CY/upIHb+1f8e+qQpLZj76hw8R5crB7bksedZe1Oj4AJWvhvdmIxKm0ksx6jRqqaIAic3
ldbLYutEfAqcoNg3RCfR8nEFCfPwY0iCR20HBnUAV45WUpneX5P9MiogmcqC/S2tsKroJFr5XbVe
QhJ3Nukh1Vgzew5qA622YloZ75//0XbIPEwozxgIV2J/5Fq2551Y0sFwep1nLFozi61UphbLfXc1
coT4zVEI8QowPGtoO3+pXap2qOcaX7Pn57iRgaXh7sHycSMoQps73GIIZWpJ2bZ30gFwuOQ6dsKB
NEdsUOacPv6PWcz5Ts9ReLrA/D6eloRaBeMi/YAMdrO5ljdq3ChxhXqGTETmGUrxe1xu42h2MzWZ
LVxhe3Xf8QYWkZLcgZM54HtO6w5ZKNQS5Mlnbtr340WBx9M7FjWiiWsW+0NxeJ4VF3Vgc2h6r8LJ
7Jg4zkl7ZCE73DMAhUZKDUDo8CAC6FmwAtAlngZhgshMCXBzrS6cB3t/vKlxSELpn54EexQNkhv7
Pnl6dcJaGYMOcBZDmerN5ZttUV0cpR50wzX61VUxyhVlmai0ykYSpD4C29bBe62ULvlSEQcdaDZA
KUlOgQqRL9yO/0ulMWhKyZJJGvfJRvXkeli7bU43Xlu1WubuSgEuWO5Ewd2gW6RTIcVRrVJrqEYU
ax5v6B6C04nD5UXdTfzodI73mf3OMtShlywOOzPRkEFg1nufpvSOnpgs7n9dJrN4A047EZdolMMq
DUFs8AATGUm5h4t/9KhkWMHxwm9UDN8JdnfDA7Mkk+SQwv9bAWGZrlpTHnGpTVcdd6AM05q+4iN2
RNxsdDC1iMyrn6cJ6Lpspk4XhyeBtCLP5PajFuy+OuR6KDsWmsO3owm7rw1ZIXeZwzxnRqf2Hwko
UM4TeiuiNtwYvXgXVRSi7ZZtMAfCVjIYBCDiISOLFTadn8J/xfv8f+Ssey/NvBSL7RMvydjM0pPt
yZsXSNBIGAaJjJ4fnZ9rW4/HOQrhf441ISxM/q6WNWv1GnYzlsE7/0txh9H58Il2AQjUaXDurUMA
lM8zXI9JcbJsNheeQ15UHleYKR7EjfvE+OXd4aIV2I5ymvW12teeZujWMQS3n27rwXc1XgzHM4gC
1yhDzwaOHqRvgRbxHvw2oIuwhFjv1c5oplNlBgOP1ESfQuYjzzaGUYNbqfiVAZ+4wBp3t2j+lJYV
IQ1EshiGyy/j5h54wxnOsz2PuGanjy9u0IS7wlwQJeghFQP2Bae0Fbc02LTRXhxIji+lEpCqNEfH
gXk7LYHEDwMwVNdhpQIXW2iBS7qUohZFUDRKxZY4MuzH0PhlJ2rPZDu/bnpO3ByRrs6KfV+eZ2dG
uWQNUcI+FvDy00RhqhysUKKCLnzn1W8uzZVsf9ha40yAwIi8XIN+t0vIzqoszSfYGfgB5G5x90T6
9Jw5d4LaB6nOaexpMtJYgoYM9M9+nnpZnhLVhetgMucDEIU6Ia9tf5zYYOlBfA9MKw0tRJh5YjUL
yIYGQrgDXq2si49Lg28YdJBkvQsMGwIdNKyDJvgF8Qk1E4amU1YIaGaUZuH+NEtbdVzdFRx9ZM5E
9uSn+9KmPfInEA4S2vju2gTI76nPytDHmeQcegC3TOGT6yw4hb9tHPUWn2URHk4fr6uV6TOp3oRZ
LKlGUaj3oP4u4MABsiC7fWWAE1/IvFPSD49Mw/1IipfdgX4TcPQ31KyaGrHax7aYtDe8tbJbrDzg
hq6n/sTitr4lA6jnzO9JIpvfEJuOnDyWXj5QSSrbtFUtO9BUWwT49ZkBhwkS3qFHhrPPB+N2X89t
4KgNC+aoQMrQBf2nrrT95jafe4261pcTaUsraF1PA1HO4xAiLtZbext0EkzOJnGIc6f0wv2DNEPQ
A0gDaP/wHf4QWs5/Nk1tv7AwmsUkhkFRkHoli8D2kh73/f6LSwrwZfaqivIne10XjzA5ZDEbOZB7
E6mmCJIL2N4hNTEzEXlg3tW30TXUvrLxsZYOQlJV0htrG9Pvx4BMr6H3vJL50EbNWPonysWEvIz6
vba4CvAgTsWjjeOg87SPsHiAzp52rKQS0d0QTVdXvpLSPvCdF89QUZPGer61URLv2LNb2yh+0mle
eQS8o6TYcf7Q9V6nBkLNHXSwDEin6nkI0AQixgUWKBAFPsNsq2GeyX7SLceBqdLWjo127GdcPW8t
qoIpN+wHPZMC3xWkw/d17B3hK9a0mj1/I13i2b+zjx8dHPWfpF3VTFOm99JYA8TV3tCjudQ27U90
bQvLOMU5MnwYKrZ/hX15H4kIMVAZyW4b6hPjCSrM4R7ykqBSUfF2iIjLbhU/oOZsEWdV2mvY2Ct9
2fIWgo/rKv2OCfO/B7eqI6+igC9g1JmxJGcEl+zN2mZlZJwJqGY5Nqx2IgbaDbCPCrLb8qjIpuyx
77TQOAOSsUQHKdg5qNJeYxgtVnI2tyGyTVR+5R9me2J6wJcgTBn9g/7heGQ82gVk4OZnMHUo6VSt
Yqpi3j6JxzHYfgXFFMtqd9DT//CqcHsMXKlsdaq/K5wxD4C0Xu+BdYpD1/oK4dNbA0UXFia1y9iW
Cjy7dXIHm8aZNbxChGE4vb98El1w2fWVhc4gVImIzAhMHffeGycnQ59Gr49XKFkZyouYmjXBLtq+
PKY5WMUeTPtuIzxC+eQT3X4EmBE9pA8AHle5ZrRl9UDhplLwGenCobROqiVGSoVzkz4BK38RtVXj
2THfyjvMbDSWoyZ313eG1+7vhAhHeFqVHBsHDQjqxRCWLBaBPm/ZpGtMkW6EugcB9b1zf4tnMPvy
FagKQmFw+Qvjt158bT59WPkv+zzolfPgLBjMgaEAfPjPscgyuUxxIkOqZgNigSFRu6YVyBR8Hk5F
OKkfTw7ES7u0KuoF0s6iwgLSA+qxz1jCRyEPtB6gj2SSBZmlaLbzsrHSQQZMQUsLvMqUaufU/Mhi
JTB37EAGNMXAZpIYBxzHHi8sLjpVDX+v/mEH3gyP5R362TAtmrKTlHnTA4mT3bgVCACZ6UD51i0i
soFhvI0U8cfszq5gbCMMDU/m1wsteRNqlB9yjs3E94XiA48YFtcRP7lLcxfI9Q9ULERDNrac+eva
4s3trdFD6g7Bplc5xVYub67Cm1Kw/vsvvZyCkOH1TOjBxSq/LBUNxAKJkT8coJx+dLh7Vho0tLDs
sSa/gUFESI5kWNJ37yU9h2hAH5b+OI/Ia/MTjBHJs7u/KG8dk1OgrqZHj8KW/a/1NfP+3b2IkVKT
B6QU4Uk+5HBt8yE3meaLVUNKPzDaW1Y3/k4952vjmadhImlhxtamYfNCw0FmBR1/xKa33f1mRf9d
yTEQ83NDMNrLcexc0OXh9MYX6dZiYoYczjZk1edfYNo9HG/tGefEVrjQRKvCfdQXieaCY1E8be4j
uGuYMGVvy6RBbzJZne7Ic9RpIGjEy+5Fxp9ZMTe4ZgeSqVD8lIH1GzrFcihqw2h2m8J+5yCXl7ky
nIQVRLGKmNlRjiUotyLf4vWsdpP38f9dF8BsRT2CPxB7b76WmdYe3COPqAsb32mLTQOy/myxoNHX
4l4uGN8T1OuW0awCn8WLHF8sqqSbVTYKyh8aLtSnvhNF4p3TchYu51R/Tf+PvkpqQjUUNHOw/xNX
EowHH0vrb41rdqOPGgYMa4rTMz1oEFE28KrQ+tdJpyUapt5STZvUbS1fW/kzZbGxfbvbsmLwxfMM
zsLc9L01h9eh/PvNUOftVo5x4Yy/O8EKkEJHahTLJge2jKDDH6iICndstrf05H2bz2vIZMyMPM/o
2o0d4NEF4FtpKlqT4QBDJYlJK55qQN6XXXZ+kO99DH3dtHMVq0cRYdk8zhaY7+uw3AA+sipWavdf
/S2mRlnaq4MBiensuWDE68Cez9CnjE4At1a5JHgSNaHrTpzvBqnsqnSWonBqrKfVSZNbAu3JmfZZ
me/yVnMh8rO5pe1iAGDyHp3jE4V2yBz/07tQ9dqT7so7BEG4G0h7M3aBEEV/yrfBdro8fRI8Gl/I
50fQZAyJN6u/8ZZM7acQd0f5NLYSHjBSUnFFoOALcaCSDVE/Se1Rv2fHRbyM35fxPdlU1LfBj9zv
0w0KuWZQHwGXOw3BrWbNWPVJxuh2fND9wpQU/swoHkyEBPkFTjVmquDW2VVWGwudPdSw6oEPr/xZ
enQh0Mk1ypmTwH6A5WWMAf14VIIPbpYK+kRg3KvwvjKS13R0YSerxhGy+qP7YkiVzxgBlb9d7wdf
hAvVtzaMlh/LtXQMCexfQ/UIAaIf9a+b7nLIwpwVkjnlpXhjPfy0Ud4pYIZjCv0aAAYhzKFgfmIf
YY8yIClcIoNkLYf/G2+7lKbNo7VBIFt1qBu8gdZOqKe6qZwysyufDD38iQnCe0YXCajb2/aVRie9
ys+HFL2U5NlTwMX/osGKZD4L6T1PtDXPl05pnUE+7OqOeYYmcVUPfL1A37NIEVA/nbT6WpcRjfiC
K5/93K0psnWmgG4tYVoYlonjoAgyPKOGmsP3Xy5IMkPEEQyQ7PI8FL14dEgN7js3ZAyBsx9OPJdD
dJr1dH/52IJE4/b4vdAHmLYGjh8a9UemvGNd054N+DNcvJmF88DaJHLyScGkPpeGWnhMTObRGzAM
+lh2gP5i/8I+J4gpkLzuQ5+C32jdr2wuRdOIjYqdGUNcXsgW0OI+i7IyT9xgKpEiWRUEH/j1y20P
PXr+Yav61dB5hjnUbD21ofV7hQiYbGs+LDupYM7BcihKOrPntSpICeU1WMN3eAy7ICmluC4nhnR0
SdfyUXdmZe+3cNPshYAMab8r3rrdiqyZlsduNO63pTTY0TuID3teB5RYA23ajXpeQsjoIz+8ttze
/sbzJNu7qEX5MSwH+qmXVDZXzVDn3KoPYNKQY6fnamMGOt0AFQKjU9RpSBKe8Zsmviwx4gqnG1vz
wRXIQUY0wx+OJ0lJNBzpI6U1SllO1ctwhATK7j7OIKmxYFO0nhMNvzjnaat5XXLwGqFVYQCLYRQ4
h80Fukve5x5iFj3PZcAqPEmB5RI96tP3OocsS1a2mAW/yapzzThC8jOz8XS8s1QXMvoV+KZB48sa
0EMlmJzsH/iYG7c5ZLB4Hfmxm+GOeotAdH8prNaK7OVsykoBCTCVW2fA8/Awi+tbij/gud2AXN5W
Cm+xxsTHGftWV4cRZyoC4DhQLv+ojsQvoUZAnE3BQDp7184IOWjNtZcT+5Pd6rpIU51w0OcLIlB0
Ma5rAGBV6PBaY6PJdccm+tBHZ1Wlz/6N6lgO5mjZQTRkjD52g8MGdxysCHQ9HviLoAGj7fgj/WpU
nB776/JEdyYiPf8B94rXR/fY+xXpICX1P+NPbS7xAMuoIM8VOcUUjce7icDF7WP+XvcWCSz/0TXw
FbDRgleyPZb9QB6RkmsjmEsLWS5kplEagAncQxzLnLjUdJn3yTv0bvxE3HCPQZIZDSr+cMJjzZfl
nfSKoJEkSKWo7P3BIB6dAyxo9Fcjjt94fm1GM8dXJ+OFhZSIGaaXJkwi4DXkqBLdxev6ukh48a17
IEysWmPzOH6gpRNQmKqQGxqe9UFCZsVcB7IrInDMKnNgqn8uhrgdWZ1eL5vX48DnCK3Bz5LwZVFO
FrycGSxYjL2PUpJP0Mx7YYZU4msIigqtCWp/3yCfsPzBEUhoXj2OtQvd+/I6vh8nnsy/+eMavD9O
8UlN8fR7FKVQDLyEgwTp0ZIpakOiHeW+80sk+fhpsBdL6aUxCFHz7SzlnqxYPd9MfZVnyBzBvATS
hqbs1lRnmSxpC4O+8XJ6Kdck/pMChWlQ4kk6hAfteTdhGiXfPCGAI2bVbcwK6Zmn4yhO/NGKebCt
S86uMs0fNrOvEjMewRofMOh5qKutuHF2EhJAjyWPGfwwB4cdFt0Q7SOzE66GGbLv4E5pTEuTVA03
RjN+RGwLi88LdFfxD/NtYQ1Q3/scZFX3V8w4l/fhfIF04nyds7Vp/NyVyQyLUncRyKJ/sHYF2ARq
U8JCHxqTtNKCcmx3BjRNGHO60B8xl62fwfp8gjKrw1Bxtu9JbzR6fABntHcImbFowarUg2GSFpjW
8/kJr7WKgxVvRRRU2S3ercWoBrX/4aN5oTnLVdTZBhf5jPiQJ3JY5djT28TKlUqWkTraPIHRPKSV
6dshfXju66EdJlvcWPWIa5BODrjTvvvGA/17iBeku7aPXwPZB1RNaxPuQcexMZk8o9MUPrpBGKa9
uiCFyDtd5BH79Ody90P6XqQ8WcXfhgWNcp34pjz0jjLIZaSlLUALZFnxFOdTaagHNV9sH6fNRtTl
KgD05nRLDUEa1R0TeC1Qd8MC8CuzIfOPyaszHISMaySl4iOp6hO1GcKSkWOEQzrchRrNRlrJH5GN
g0Xss/S/ARU/j0JvbNAOfysPTnmsXgZUuC3vs9YWtP0f7Fy3agoxmvNg6qECYwP4AWoEQpJVs12X
4kh7eP8XjVacPhou5FSgIt3WZ0FMHFllSUUlR8ESihVU5BVXG9eC4lsuVaCwExF3WhYPzD4PzPL7
s5aH5/B2m5ae+GsUtGb1ejEVs7cqeHOdSwrvTCY204k2zWewgV3jolO2ost9U6QABJRCoDt0RiUX
qYJt60wS9AZcKXmhr8MeFoXnpqfs9DnGP9JpIRkZ+5w3RhBWDIBa5Q9plJtnu/jNip9W/NgUzJHg
E+miA9FfV+1YX8kYJQ5D90hvcc/byas2TJeJX7T1ri+Ag0VkKL9ZwZEY3w5B/vdcNQrPg4GgMvnh
CMhh3nBpWsaW4NaghYMMfPc6Tlj4Ld8KfqfmymGvtOnHyJ1GLvD4z0XucoezL1H+Yc2/bm2qnisj
iQhJvR39vuslP5NT3fjZy1mpF2snsB0eZ1nNU+u/1Gygk5I619hf4eMCOolh/siUaP4foyGa/A3R
Pqwm0WPE45BTAI4u6FTvDFyvj9yDfDd/kn5mqKWbJio/24fwoMg46t42pyZ00FBbgAet+8UkN9h2
Ju42DP829JwAL6YaCYU0duDoPw/NN+94eIxuRsKQ4q/PoFY6+NeJ69EGqfba5zSzU52BIM9MUExY
TXLde7+tPRDX+1Npfa32bd20/Coe3W08eqDiKMlr7BOTY8ObsJ4c4y7QFtjGSpHi87epeEtmctuV
0yH0UBZPl9wnNiRAMcDBhcSXkSY2HMl3PBdbBs6FqVaFBUPL+nphmUQAL+mZkR5hmq/I/aAMMpa8
Fr4R5a87GcMnfa2tm9GaoFGYd+v9+M6HNztjZQCnjvv9pRecqc5bRtO7z/0tuofo4YZk8gm7g4nA
N0lxddH2EPPlNvHXF7ElE1syyYGzEQRJg5bhYO7aCnpLOrfZLlEmRnLA9+VYG6F55S202NAp7g0z
3etmIXm5loEn1pXE54FVFyw2OUUTErpJRotgNM/h9gfkydvuImMbyF3QD4b2peZcnaSTLKjviSD+
wChOo5Y6IlCLTlbpDqBVi72bj4md2czFzdBCr19SLsk+BH/AKLGWsT4eANJZQo50w9V9J/B8FHMI
zPl+AjUOy1EiOsd5tCaP4fSPqZWvG9Ml9L0KE94ldqQriJfOYu8zHaZlbCOrbxQELvFDUve3WkCC
dDK9GP3846ssCgRr4g5dUPi91+4agyoM1LvS5+vd72QVb94wjdc9CxpCGd+K3MXS3k6YQJ60+tcy
VA4E/fIlF2dGoKSQMT8nwTw+pwcnByg6zVHxtXsCzod9Ge5JTgtcG3p5quVWBVIYcxhEGe4Bvd2+
WmT8DPatfvvfiyk2rW6Ibc5FFFOwkf5obQKSaGavUV/IKLzFJie5PEkHCFlprLpanrTQ25N+QQs1
OhSZPbOiqiwJUFHAHwEMdWSvhKEQv9lh0m+KEysoNb29GgCn9KyBsZT6QlKOkwgmt+nuwXprWGlo
yy+C74h6NmyCj8vnolmBoYYt2OXRPYaLrBE4H0ShL7Q6PLVh6FeE9pyQsa8LlI0GXjJdZc09oWAm
cR6h2Lhvt1tI6Ng4CDCvDYeg4x1RkkM49CVcqghPg9JKa3ldCnfkxeEIJjAxq871MaKsipUYEZiv
aqBmVsaQ00obl/9+YLdZ5p8zHfuoX0bpVNTwEjdj49dANyJvnM92QcmKrL4RAN6TTO1fx8hAT6kz
IO9dy6amk/UdSDzQLDvhOZaBSW3nqyfp7sFzwPOuP9UfglIupDwJfBU7Wn1HmTBluhREnfmp0PLb
VJRbMaaam3LX6g3u562rqKAq7AVW8goNWl2ckvikQrpuyCRVpCrW7kDxppLpFKUavGZzi/iTyLlH
jfTJOgGcYfYrQc3LjECWwlcR06TflTALfrn+XTvlFJbqkK5VwtCqDTukl9KRCwkDXnE9sHV14Fvi
J9RppkoZ3gFRrjWa8422FPMbyIz2KDRRtEroV0nabrca53byGzAFLgUl0zHzxRayA2fEt7xVkSoE
SUBFeukLbUPCzI2Y2p3F5xF5ApKYzccrcEwMnmKToADQ7lvxSzTqjhp7aUuMd4hBU+xFQz0Bxbf8
b9o1wku5P6cGQelqL9o4Qfr4D14jQgb1JOTX/oJ1N7DPbd9Osqcwz+b3t4WlAY3Y0uJJVuXwQcdI
GVX7QWol3XyQz5z6WwoCdkLOTF2CCK4ysv+rwfyUzrB0SnNBcv+QuMjel2CfETnM4CcEfeCqjgzW
BaxP+3LZ7wPuH6dquoAbBQoS07kHmX1NIa+n9bvZCgFNafaShUzYzUCBM6ETXUt5rHZkTLqoJx+M
zExURqleJ5sjzaICz9Xg77rErYXswMqo6OCfjEVn1zJRl5kV7+wyK8shFwUazoysl+Jv2qF/I4Ee
qy86UbcIX9J5gzhHqTX6vwss5GpAkUvUt3jertY+hhiI91MiSPKA2Q7NlPH6edeGX17HwPqAU56e
3ImVkqcBTz5rVEFESp1BiV+9WaMQmhq+ogNha2okT22Sv8oP951gLCijSMxZIG3Xm80NgH+0Oz3g
WUJ2YWROp8cD/E/8jD+JApNSiZUdcGUhBoVROZXmnyY7RhI/ixmsSGV1aT5mSXrKWUAjQHeGkUFf
FxWUmTI00UKTFQUd3s4EMF+H+DWN/IEcfOU+O2a+TKb+S4Il8JAXQRkyeeVqM4/7i2tnFVntY+p6
7qaIEbk9nOpBqYPJLI7Hwkg/UP57tJe9QKjbERIpPkGw6e5lemkBsyudgrA7Acg6NR9fA3Biip5F
UaF3RMK3xO5jSRimEVMalmKCELBmBKrObxihwDH7pehhq0m0BpG+E9c7YSHTqIzJzHSfLoY89JwZ
wr4IZwubkJgMyvFm+lmRnUww4TE1jZlwCzRhadQ6AluS1RhSs6HhgvxVtQudMPd9GTFDxVeObdcn
vSlQZ4b1yveFy8xFyrmJ/j0e+O9Aiq3sRqONy8ecDUTsGk9lrdIabONaf4Q4dR8pE47A6pwP435j
6WWjwx4XThnVBj2MeChyWek29laKhYqMo1AeUEaWRSpRFMTNpp/nPQn1GkYPLBZ+gLp2Ie6WIY1q
Xgs7d6fAAH2iIzOXNQfN1HxszrFevKdMoJPxutjs9C/068TykhgmY8zKlHAKZL9SOBWwvFuOFQAs
nugkmRZxoXHeXa25K+yKcNZ3DtbKsHGyEqlf+uhX78smBjPpPbGjBhejjfhAnxPdvJUf7WULMS+I
PCpeD/n46uzjpDTxrd/TY3tB7s12bSM8HUur2Kh6gAXkGpwiL2b4oDlCiw39L119KUEHSqlFCGJ8
t5DIph2ee5GdYZJg9oZvhNaI5uzvITueoRXUVAmSuIsVHrtHeGkMQrWyHWqY//MA5SfXtvFoNqMY
pF8VwPrnBLBMWlhJCeGUyl8zimUZqk7ZzJ+cy6ylq4ZFsyKlnxMtlGLhu13BUErt9h5mEkJYkVWX
PY8M2dXr8RB9AUe/DQWegY4SxSHuSgfzZ7fluVa6eqXFi4XXzOv9D3e7S6ZC83Fw8ilqgy5Sf+Hk
SrEGQRdNpLRfFREaR1Qq3e3IjZWq3IWYu7IFctgmX9wDFn5GCqcOg3ffB9u5VTCj8G32EvcJpY94
LXQtb4h+Qomju3Q5gF3sTtQjaeUweIsRGEDSEB58ivWmzyVQz+SzsH0pUeMF3GfgPOf/5xF8fzCn
KSFtBlktluo0cE1E9y5OmylUx5MZwaX3NgIrA5HA/zpbGlh3OZdn6aL5QY8Q/zYVBowqJGgg6KjY
yVO1O9SQXmczYK03zophkd9EHB9Caj0vwuELiFq+E39rwRvlPEXOTTs0bhrRPMc/OstK6CXEP8mb
jljnDHqS9IbU3d82hkEdcjrDp4oSJtxH4pNb+lG42m4jBD3+o+oeo2u2yLkRUT/IU+BpLkv59ojV
0P28ITEHNP0dsUSH6o1DaH0qXr/NOjeyUrIOzxfyDL/j0o0G+PVWYyQKAjboQJTYOEVWhShIHN6b
FsRb9JusJFsGm/QM3Kgzlo0phQbkeTmI4nB3p9HBnBmj11X++wL0xSOkaErvwCRl0QjcnCfI5QgE
904apo8UQamLSdt528+MGevqAJlm5UqNeGULmVmg7cBR+P13w3PjoUH7K8XnUSLUCuNKIJgHGSUn
ZSV++RUsif3/vOM2BG1f3Q+4sbwEatix/RTvnMGgPnq2t/m+rG7sg+UMSAN8/y3m3yy7xfu0YFNb
kl4zJ3RywOz4IxH11Mu4zkHnef3cRHfyOBfPXldm8q7RwiTHruTb14MTSRtFJIXJwmOsCtEd263b
jZ86ndt7MwRdmSROnIxdoH+zwgieOB4h1hZzQ/Esm/xhR/Lt26s53qPy0L6WYSc9cm3cJtlkyyjw
m80u+ovdDtARX3wzi3ddqziEbp6QGCDKfHz5s8iXio+dVe8qJGtZbYfXOtHCwp4RhjDqBhetbDKB
ezcb6TXRfLWdG6AL3fJyANDxL3CNYW7wbMEbmbPdsIlmc87zn1rnFx+05JnU0r1yEF0mAZnYel2W
a2kaXL1Bj4D+sSkdf+NU04wrSaDiQbvFiouHsaInu9yR+9PMixCLl0z5OcdY9TzTLpS7iJ/9fxFw
/dtkoyg2IFNw+LF/HZosROnfqvR5RZVs/LdLLeeKCJlFjM8fEjpcCT4LfBfyAmD6nPo5Itn7lYeK
WQ6aWPQ9mZmfMJxZWVsmlaqI89Rnl5mPbhC4T/X2T+mobMAnZByFqbm1iGpw5UHsFpBIEVM16RmR
b1JOYcEP/AYHiBHBv3KX4Z5qyHa6EbzvSciL0xqG98IdQCO5zgAcCTs3gHZAfRDpPzE1+rLkFq16
vs/lVv5oWYSXoL3naAprPxW5q0h6XYk6ro0Jinn6mg6dpDllkeSuyWxdXcNsAfS7Js4yAhSdz9hA
NY4LFz8ET2lhw8CApATVTJ7Hqk6e+pea+VCXkKd2ITu1XDGB1n8gPp/uo7wnH8VzqPPfu7y3Wqy9
SoRxkVNI6Ysonb205eQ6pGwNwCXLaNMmWk85s9dXwdSklrcEpQk/wCU/2vz5qJPqZA/362dZKKp8
xmOLpw2z6HO6MPP1fT6lCjF3Qu/jmAME4ELMeJ7Cu03gQbgEfOV5PUMDfvquzAY1Zf+WujSmDzEC
PHNDh93mNEXaIUUg/jnEz847qXLMYzd9+XolwdiuKK+zcmL1aE192T8a91tJt9xp0IYoONrdIo4f
B/R/4Vgq/8LRgdALfhpv7RyOK08cRYrc/PHyZT7qJZ6jFl3NBRtkLhervQQa0gS2qmWXGu1f1f6O
GGRlQdhBvMWFSmSiEfs7WulbXZy/yS2MSCUZ3yscnc1uy8aoD/hpYfzxW56i8L1krQf46oeJADFn
xQyb6SRY68Tetlp6bhumD0ydOPBf/0ieRvKkm7e+y+pAcJ9603ld4g3sTgKhx7Gpm4zL0Tn6Obi7
W5kynWSrzuryKNCbclke/+osJdrI7F23ktnJUab3/d3r8ZVHV588GALeXwMb8fC+XI47ZXvJYy6M
cEDcTeXoqgda3UojjjgArywJsLgG/bZqxqdcDM3LU9aYLB7HgIzBYOoiySAIJ9F7tUE2VyI11UVB
cBZGjKoN/l0Cg9K4dEvvHiHmq5uflUQUA4y1fgvcUCg97ZAQjYIe5U8qhEUvSYxyiZxQ/KP+9tpZ
bAUSP11jSwF6FF+stNDAPvrHkyvkZfDaGMEuA+YYq7JtxpYumrJfVfQhHz6NyE7XBwRTVGWVXxv3
TesvGAK8+htjtHcKIXNuvhCCgOncPWVlkLZvmliUdssTVTu7C3mGnOAg+6dcznUqI9mhaZWVlkBc
adMNwJnEEaU82IhEyhEx7ZoeLf9gBFnSJWVerQScZgrUC7TlzcxD3SFo4W1q/QWVBFbHlwH1OZCI
1REZ4Brw96rNNXwFyZ9ra2bZKp5aRgAmIHZYKscXwguguTcQUDp1zDlFYQEPpvj8Pygc4X/vTjTK
Gl91GTb6yvp1lhgqK5F8Syfa5Y19cioRj2Q4GblUf2IKRCY8DzXyj8f2IF68AzX37yfVBptCTjKM
LOL5CB8pIQu+DdLHb9eVxhfiADPP3a5xOOY0bRZcROkne5sbRj2UNg2X7tXv+3qVJHE14nXASIEE
fGhfHtan71DTw6xZ0BGJwDlwf6j7yMm24NRoacUfUpCALa0i8THQWnn7IqwLYU/dIbC3M8CbYQrI
lnowqbqe5QamZ0W4LhRCKpraKaCC4sAayxSyNlEyPG0TQexoppuY64pj8KC+iE4dnfgE+mPvK+RJ
kYAAPyar/Uc/RzP7owr7sImdCnSnurBrA+ljUOw9e2NCPsrdQULWGdXgJ3fRMIkuZnKMc8nouEf3
RbRanWp0I4S3koPyGvRNfw+FmNG9bF/HLLa85HrswFJtVPMWBDOYqF7jf47Qcp1OWKAyQfiJF3H2
lsbw9hs8MMHYn6vNbvJq8ZEt9zgLkpPnoiNhWdMlwtyuRHZuWtAfFcodmoS6FmJHVu8boyJLBMwj
oTSJmCp9KaguzLVnvx/sDFDMDkQWDHQEhJx4I17I88WgHt+li3e5V/WW7NjNXis0Bozh3ugEF5Nb
gMd/GUsaZ5PhrCdmFIuWXwUcU0oA4hmhr/KV58EVbJeQswjMbQuxvtffItqzqN3J5bkKKjdgpJG8
zhchMt/5HBXjozYJ57GJ+UCsT91Z+OUJmmJ6+8jeQbRypl8mzDbv33qSmFdCvVYbMFnWtWMgJMVo
Pf33bDAo8s0nHbB7BIglwUqnZJJ0QhJqGqCkMJ2LXkBGqoXUvdvJ3YOKF7C9gKM73eQemiVsdrbB
xAbcRoH/3Hf5g8rkgD87p8Q649OOPzLLfIoGLqFEmpo71lUBoPx8zfGwcygbzhjU9piem/5q/1Lp
QXxKbOLLbDhtRjpxY30n+jxeONplnAmhGVRkiaTQC/6o2Ta4FMbFSPwTiOBUoxYZGKJzfjHJKLVQ
K51auk15GjVSo6IiruoKEaGGsjKCZx4sEX4jpHw1WkBdjcX/MSMkWyQA+DqjT0Q9C0xqXXb0isXF
F7BAGrlsB+/Kl2/EEIiTKuqf32m6VgqtuQAS3tTW9YFCGNYUIYf4+M13wM6rKHFEu1qBo//JvQya
DwU46nyeeO+KW0wVRVMwuAET+mv8NulnlCKbQGsCSpEFcqY/1tShzcpiKrwkjv2Bnr1AAa5idGJM
1IIKFQKXN3PVMubKMoVItDYiRZMPxzz8chSG/qL2E+Nc48NLoWsIMDvJ3U4gyUMCuqxkhQ7Ukhxd
VnCQH7evr9ZciDgy22hBkoFazcuPlcF3omAJ4f1yABBRdWay+fRr0lfhxXa6Oda8Yhl9vt7pcKKQ
TJIfLvE1wNboryRcoN3cZHraIJYnWskEdlKR3y8BZWz9IWn10XMEUH+2lkvJJ3jh18uvVtHvuRM/
Df3hBUnlvTd27xrT6AUC+tIA/Gvxvtg1M8mtL1uy4Nxjb/NSyNrck/S9dhJB49bn0Cz1JSiRKeA7
28KM0NlzyiBYMMFVxwEeRZ7UoZwsfLcTLnMGdr1BIza2cOaV300jzWtmw7H7m0w4KwekPTKuCM2c
YbJdLdNPdvDBFR90UMal6Yx114+naiP06byiuFL4DRlJg0wC3ViKHKTd1o4YvTfZrf575VwAI1Ps
7RfDxrLErWgvWKciA14h1HbA1m1PWgnL0y/zUuaeU+Trjfx4WlXE/KDWn52yo+uLO/p5z1iS+h2S
YhZIEkI+kMV5goYhctFVH3Ol1I4biyCIn8qKe4xrcc57ZKQS/TiUr1t6dZA+rtLfWjTTbfqMgSyU
gKUbNBaHpD7vEOhqCI6iInjocNjMzHB+JX1WGjNLcWgxSsuTrvI7cwyfEE18B7n+sOUeA8UiADBY
Gul3xgDah6pU+VWJclomdOAB+5XArB23KHnjam8OGf7R8DEkG9xfWpp+TwcdDKSnychQmK/an4dU
GTm7P+x+GTP89uJYHAlzZStd7Xx+hVhCz3mmNwuU2Wj2CSDbgIV9AUHgQ/RvP0rglA/oVYBsUTJK
WRIY+ysqgLGJv+rLY/fjYvLKKTnKUxgUX6s3rQ4Em1CTzzzcl4RX81Jwg12D3wDMcZ6Wn6rIgckP
qXhtgb1glFRm29dkH90QuuDDg9ySkUddTRGsjPSWUBt+GkY5eNziWsCp4OZxtLqVgehYoeLpANNp
3GtZYelutfHaUNQG4iU8MVsIybET3PExSqtNUdRUmpWFOiyFJ+pqPc3v5rYr/ZXL60dyrRNwTjoD
cVfhoZNyKPsUP8zcOOTX+wpWlrRgfrVt9nOp0fktOGa8fr8gA7iZsQKRfCJFMnhToisYHc/mCoM1
p+Uauh8Y9RXYEvdpVVMkXUD/oSIFJymwD2MCsw7iGUq6GZquplnnZf5nwlQ9aDmf7Wdkgt/X10pq
YON6BqKNDYe6FaEt3J3AA6FGuL45XdMrYxnEwjiiuaX4diy32PeFn6PED/Yjt3BALKQwm3JnscoE
hbWG0kYywsHTX8/gYyz/bl4QEpgw4hinafIri5m7obVXTs6TBgdkkszJxErZggBTkqIM6aKdMiGE
uqyd/JqhLKkwSKvoIasuI1Oa0xmuEX/WQqHiafal0ZV1Lg67zcHcrGhYQMu9FbzbV2pMLp+AJ1UZ
kE94Ug1narB+GY8i6dkWmwohTs67P41aXKX4IUposPNKUtfkmqOZkNQ2CAf094bCtF5rW09166YC
JYAeqOC4JzQF8zrkjxJlc6wGRmhSapdEF3+2uv+nF6/k+ZB+75y81px1JaLZ+QeV3dzb43V1uTr/
octGGnue7zfydNR7QV7FsR4aZPc9bBFdiVTxMsflX4JmbXjTDqqDSn2gu/H+TLZS5YnTfjhammh1
3dqsUDyBnL5QSaOW0aF2gsgCeUmxmFeQqPFJX4oWBJ4GU4vRxt/43VFZy2oKN/Y8LcK/8yOKBHL0
V/SFEKeuyuSprv2orpsPoDZTnX0b7FXeOYQHG4IUqUePUPoR2y6vpkxRdtE3bf+FskzT5UbGCcfJ
F8pCwj8NfGVW+qmAQ0ZdHZEagCGA28bCimbw6SB0pC9WzzXY0wUeIxWj0Qm5YRttzvnlR8qOOs1S
WUk1ee0MkFKPCNfNJrlVATHiJPTuEhMrwA+/9LNSlQbDuNJxe3KvXmMaveL+hdnSN1o+1G6gzWG0
ulh5BUzPst3eN7WnnVpoAqwuVQTV1yRpFYD59NBctZMtkWYiQGpZVLJFnFZJ9M2nC5pKhVOLKoxE
/ZcAHFf+489E7fDbz+nd7MqnrePRNBkCQnk0x4OWYbTzDiXwHchuKg40gE5i4gyrVPeSp2r2XhnV
1RV0EcbQhO5jBj+N1B+lv/WnbzHNzVd2fwJKygtx+R+q82mCdQkh6Og8T+gb2oVNQPjMY3nwHKDA
UYfaXU6J+fCwrPvogXhE/x5pa6b2FdRfWKCsZOaTDn1/YXlsulHX8r46H4SXrOluz1+aT8RinLkG
z01gzGl+cEAy9YqdgnQhk90PmFzQCb81yDsm/Dn9qOf66d9g4VAnqKoOMR2Q2UzhmoYAQFLFKmsc
NgufYrN2IDyfzdr+hLrRwkPgYYJzEHy2XvwO/F4IyqSU7wdoyWcxhetq+2chS+ld4tQqgNGQgLlo
tqqoym5IKS1UrG5hwSAHHUQHC44VV6eWAyI/dhANSe4d+f5SymPVdj+CVla3kLhHEaUs+Uy9u2yb
gSdbOLn9XS5+qWhmFKraRnyB9UvFYjbO0tjvskHh1D3uMcsiVGFFP4WUvhXk4GJXO2UD2O3lK7qH
gKntrzEfrPsDXabI98NabaKw0qcqNJ5r5gdwjgEryc50rcKZ5UK4zkV7yo1TqBbzF7hj3XvObzg4
XgbLSdJbq2SyvsFqNpxG5O49K5ykrZ+k6s+x/QXHvVNFXnyfiL1vJzAmwJoR2ZvAN/rjez+60dxk
KzoIbQ0RNm5XcsB5LfMt3D12MPdunGvFZyzCG1ukDM2q4+9aP69B0p7xDqXYtBxvIjt12Dm3Fn6y
pi62/vs810tzEhyXLSVpwSWP59PNYH98KXeviwHNKmzu1Jd/JSFj5KOhd/Q/2Sc32X3ofJBqUUPr
vO+PgTQ/BCv3q4bXPyQyw6KL6HqEJSQ3vu1DVMJ00mQxIV3AHK8WTwY1Xun4mwpv3LOKWdAiDId3
QlSEHB0L7Ur/GUbZ7TeAc4GgT+kPA7xBnLg7lg2P3cv0jhiZC0p3CLbrbcdk2bn2Pm10PmCRoDua
NyxySkXydVoQWMrMeGmwrUSY3Pe5AzHF4CtjkDpRWHGRNZpJF5ApPHPQmyel9gHNlSz/6yXsnLjc
es50eRsDq86E8FJGXXxQTgpU6/EHezeVusxfWm0APaopnI7xH6fcNm2EDMoACmdyaIS8Z25UmT1V
1Dbf039XBrf2gEA/E2ObR/NcjKAKC/q2X3Eg1b4Rb5ozpyxwZiT5403RagSIlPtXIAa4EkwLJlSK
jjXgAS0f7COgqsEkUe468GTJ130omEp2/QvuVTNYlH5stfqdQYUWz4p4g85kIkOJ1GYURjzS7dKo
Ex1jRv6cO061823B+gwr4pU5xC6eliJXgosVf/lZpSXqpPpwgDCyTf2ZWs3J0pwtHoEszX+7kLX8
jAp2ig4iq0kTgWkhDFMTfohKyK6gUTEGcGxeDD498CBMNcfF+nIJX1xqyAfHUI8ys1ayv5iXMpj2
UB7C0Y4/sOMobxvBZlMNZkEGwxUIzVsTP802venopElBUxsDCCAcuRJwdOf6Uy/+I6+scjNJJos4
FY6XvxwxMEt5nuTwZmjRz5PnlQ+Mc2DYxRwRaRuHj8Ryx4GmefSiqwjAU739mkJEz+tPp6c8qN3Y
B81nq1HEGU1XzhjkYmheNdHyLbwb5Jx79aLjCnChn2ULrXmVsn9z25B1cydORhpZEr7VZ/EEDgk5
ygOK/PGaeycmYcV++JyJjz4BED4TfzYz1De26qkaekofm/d6BqvHWLP245xSuH8YlKGfCHmM5nR0
Nxm+k75FtSzJGPGhRJ5SaAazXfdJoqkQvwJ9ws5s7BfKzLu8v0d0eCliNDI6bk1yPIVMZ/AkVhsi
TtV/1PGiplTgtPfDhb6OEHE7SMEfbcSXRBCZk07S+zGZ2CbJK4x0+XQLVwoKyK4VtYs/aXXtYfLu
mrSQWWgri7cyRY7Slf95Iwco5kHj722KIH29QaHw6N9KJv28npTnYrzO5H7HZltlryq8qWUXXiQ6
DTVqFkcWJ4XgImrNLvyWnmq/k3LaL6h0W3LAShFmlNxmLcU1yB+xstJPg6Sqsc3F0EDP1yQ86kZO
vs2jKrpxvsQPma1Twy3/CGMMPD/EDlRrbsOyRI3Ie1MFNaqoLxgdH95KVLafdok8v+XbvcEsZ+/s
B8G+4DjAbxfoOjWAayFfU/vef1pImXrcg9+6fTxU6IkX5nfdtyxD5NOunCioyqcai1EQbvpa8HZV
20OEhcbIHuiQtIVsxBc4us1nFqI4v6YzwsSIrHP+rwK55VxyiZzVs6YaVKMssaD15dISh9rkntD2
e01HVattTwr1IFQ4zbxPPEQ6PPp50Emt0/fu/Nz3e0e1A5BEqtimeaazooFn2l/aeLvQNDFj/kTl
Qp/zSlWlck2kJ2mwDDCqE6lkrCav70WC+jo37lFIw7TMEOTQA5Ig4XBgs0I0SVVdi5PeEVm08c95
8dK/hLsfdX1xjvcXTswmkx9XeSfUdlkIuyggQP+U+AoHR4KcpAAAhgPewYT3g+lmD5P6RLSqLyRL
Zocq3CXBZLB4uicM17oUAfoilt1ntLWK/wqbf9SG8oQfIq7VFak8FVNvBvdIWhnkeKeEpnjhmk1c
6pfsVCY0OgQ0OIoHwQs4a7fl1jykoWxIggjMDALHqkKqVk72Op7WOd2PCS/g91k95+VSlT0fYunA
RkJIt3XMuvGQQ73XKkjUT2Qjb1oTFpfAV2cI17Kg/7MzWopNhOVkfhAjZCX51wLBjGdff2ichGTZ
J3JnUOflaYfgnOdt4P/ZlTsymS+kOND8suB2AHj9WJMSZG5EmA3SkcBEtoaV6xYbQsqYRYltcYoX
/kr3XTxyOyoSKKdUCwNuhHTU1jcc0bW4BSR5n4Lm2bnulvplDPY/xuttGkjgj5g6reotq+bILnUJ
hYBwUmu3Jp1sz5KLS68nPt66ufn114Qn10AxOejCJ7I827Vx6xH/zrYjKNqUrNmGdwiEFZhs3SVD
B9efdsgk3aCJgnrkL+M/4KZqzeJVDnK4DU6kuIQ3yPo4L92IQznZN1hgxVdWOs3XVVLBHDMKfSLd
1tRg3Zmb8Kc9x0DPRIFP756W9t3dBkv1XhBpIgeR8dFhhMl0VWbpD0/7831yDQRCMwtIv5URNR/B
kfsy9znZKdKZjLrI/MOIjkoczbNVEMtK+sm/kSYTIYsWRnkdR6s6+tk0d2I/LUbHXiTo3eYxaSCF
FDIJvlsQDvubuM2hd7BsqEjNWQE6S4SrgU+9JNn2mE0huO+oBn8zFqgh29tq3vyY3oF4XikDtG8A
fXDf9+OjuyWV71tyl7jsS43maVjj+fMtjAD4Rw0ULhixNNXcK+I05q5fDMuXC0ER3g6lZWynFDym
vlgdNRFVVHDXXmalmh9XDcE4XxFWjlXJOmIiWPOGm5s2eYxIU8gR1LUuUABJ3AIB3iiW3RuPNUoi
bwyhjOZmVDItbS6gO9NSbjOM4v7zmwHoO0aarVkHl0TjOsbcEq0U+La953hTdgyDEVMkL9FMYU1P
gUSWkbEglT99orKsFCBxMPK7IbccsUt31EPhS5FdeFnjMWo/v+9l+vdktEz7/q2qD0Mayc+8RPA8
EFjtPbiDfig8kFZptZISzC9TCf06Kt53RsJEthkFB0zUrGVsWN1C1NcNHefLoOxGNZO1btTLlUVQ
1SaeI0Gg5tnXMK1SiMlIRsfmzgbf38H38N66VJJqn9Qpf6m1eMfxytdJ+6Aau82U+Bz4DYwc2yFE
BwRDWLM3vcfMPY9X0Cjj8rFCWGCQvONt+HJ5gKd5x4Cd544POQ7jfn7P5CA2AaqXlwYV4KZMP74E
ZBCgrTahDLbMLpN95OMVKq3HHj27C659IGGZxzwY9s/NKj9sQQMMPBaZBCDpzxHzQnibZdG2O9eu
nYVrJRGrWNBnMhJkVVscV85vMzYS0ilwDO14k8q8kYfhVcqxpAs8cfOfY4WhG3aU1CxO31em+l9S
lNZ032OPWE2pqNubslE9iovEzyiQUte/MU2FfI9jWpEcWfAZOwE7BhxxNswHZSRmvUsnk/Wi7irk
Wy856ne8X/2zkOXLiloVxr31UEbC/mSGJypYZxEMXOBrJTTZ315Lw30Joy5+aQh9CQTow6LH38GR
aXIBMIQeDRxJ/KZaJQChHav8FAgB7el1FeZ7/u2yp/1oY05JbHZVur6+GAjVwTTlElGG1C8IZLe9
4iUrBbHObO1wZmunVw3C+TNDUbOaFluwf/corw7bAVbJzkjEkA+s24ViAXmugVEk+2SxG3fzE2Ve
iYwYEBnjBVdFMfPojUUJv3SfDLn2P1Cw/70wmBYZCZRXeElQn472v+Odf27Q0NnlPGgw1V8GyE2n
WSROjwGIaxcgSIUKLf13TPB6Rtl5MirLryqNP9yof7KJ/sx8nXFYXYKTqAZbKm0ghDpqLomC7Mwv
Ea8GMES56XUaGSEyIveJxNwqJ0oO2hfDgule4vYqJfUZrc5NjnEe9cApJU1vmLzk3gE7iU4My/zH
iQff9KksjB27UuYL3QNkGmCOAbhHeXRR0IlVa+s3reFOS9+7TVPCZOYtfRbGGKUTh39Y4wXfWfK0
AzKp4gI1BB5X1bDnRXYWt5WP8xnU6YMmYT/2pKyfUOYJpYYiZ5s1483tsoAZzzbRTz4wTdmMo65A
NzdPhKlGVNtAEch7RQmuoTlV/Tu1IK/myYbJ03sTRazJdxb7GW6MXSPAt+nse1hV2kaVkoaNOn1t
4MvneC/FNBG7968karXUbPRjk8TZ0uTaqGq18YK5HRjpuj9V6vW1YO83+bWcEi/UKEPyOU2q25So
es35Fi0XGwpLsS/YB+LVRghY9o4l6YQ9YKQNHKHlhP2X3/k3X6jKV4zvWhcKqR9uyaIF3gzr8XL7
IkNXauT9Io6ATk8KQgtV4WAcoMwkgIPZCeyqFTc9P0kAwarFcjx9LNggJRovCYfMS4J+g0LJihID
PBfqQV1vuuugBl6ITYcSaLv6zv7Ad82eMm+NKDdKfoetjm4TOSM8lSiU0VIQCcerrADjO2Db0Kpr
LQI/a7/rbkZbSpC6hbZm1BYBvdpmFuGKNadFauW8ZgXwoq40NiNHZ8jg5TYzFq4tWf/71lq7l+g3
fntNwYMYyH9E6h451o7sGsuCPDIvefoqbD5iw8f4VLLm+tyaHPajxybSPvKPYVaPFjTJun0BIQrm
dpDIqn6//z7L0ylHTbd3b0cU/uW/4poWR/8UCJ7fzYk+VXkg600vjFUMDLcKdpMydpaEbKMtRlrd
ATgibdusGVEtE0O6STxw/6UJrD1WLjkbSSBtbLncAQeiLojfSVPegfTUiVezckY6V86EbtnRmDVH
L9OknjfWrPx64XVNx7ctOlqFqUJ+1ALCTguo+CeFn5BeKrsWzKyBUkIFFAg0CzEdyf0zd5rRg+iA
GtSEFYcYQG9MuNl2kvB33zlG+Iw/bHVYu4iRAkV6KJbKXkothBL38C7SKWrAM+hdZrNNPLXbQN6N
FD5yKElUuLFmPdOL/EQCZBM/RQSUVcg9zNhCrymt0gmYpR2jx/akBqct3nzV5Eu/IMljR4868BBa
0Dvy9GKd8zNKvUHxRnGdK4Nyh5yGxMsKj0wKeV7bZZjOCIP2reOC7EX71MeCI/pVETgSRbNNT9U5
C4D8HlT2AShh1iwu7AtneXKPRoipQjy8mpFy+Ur0yu43BL6JJMVoVaEl80rB1ZgcRYvyLhLSvpXg
dlMp+dxYmu7W7yPkU+RU9qkVxRqRkJz6dnf8oYrEq5hxe3eogJPb7ZFS3ZPrjB6CaHzR6W8erGM+
BePVLS9x7mFUmM6bMF/P79O2IZsUA6zVcFS8F1pk/28+5pJn0LzecP82vdMmfuykqHNb3fCs/cre
SdsBVRm6crT+x9ooBstjgEhLlAmEJdMu7+gg3nugn6p9g+xUaGlmeqh875fUG6zis/hQpa6YVyLM
fCdCAb6hWQ0NVWC+c7thPUVPIDniiOYyTQH7Chaq1AwX3hX7BVouVq19+pwSsnFAuZaYHYM/Mzdo
yMLQFpFnUcSegJXO3mJ2s5chmmt4mrzzHHCtDIhJF3Oq/wisnO81ZQvg4gCb1CMAciim0lOmlLEn
iJ7bQFbbiJC3HJ7IfP7x0fz5X1u9Eo+lSMRtDBR1k1UMHYTDrmabIYHj+5WIENt2b6JMcalHMJGB
zIzacYjW324MTOLGJtUCt0UXWF4ZEym+DsNTi/OTfEsHtryr1sP/WhOu7iznY6PdAAE6DRBbVPdi
n3uIqv/lSLei87HYjtSUe/3mBe5Ig+U7ylKgeB33xn5cGsmfkhVO8VHlMVJQ9Nn4oCizQpKsKx9b
vhSZgyoFTsYzDSOkEulRKCVX+vdw0jKHeUvRdkt6DRWiRo7N4BQlBq27jkZqWdKfF87YeaNHi4Tg
E8tF7CI3eod8V2ipfuXxTXOc7D7UAJKYuBfOZJ5NBqtdNYRcXiMoxuswVKUUhMJlcq5m7JPw0w8H
GoA5FzdM63wnFAfjwgPjGfIx4XdIEh5dcJgae30o24c6H8+HI96Zo3rwNDqzhxZCPiwqCEc5mLmZ
h7y9Iv/eS6so51fJa/me5J9OvpRm8Mjk35+yvUtbsYUZdebDghztc9lm7hFWdAzRngkhf8thsIUf
jKFOUZosb/j//hb1YL97Q54HhI23YXci6qbCxZzFVZwbmFYAzxH9F8Id5Nmu952ofisGeYNZ4VmR
RD4swdu0uJ16BYeTYQngIWLanmhAQdB4tk7hrhP56YGpISWPHocb9dNckDB4sDvsq/eHCP6rFCaz
LpCjCykVn6S46dPkDntY8EvHastzmocB2Hrk3m7VeOX9wGIcMxMSF3knKaX5Xl4kuLl3722bjDFp
R7UMHruwMI0IXGyHp6NuxhWwYGsgcop9cfqspCV2n5HYra9C71JvReMvN1Cs57HgrkpGbnVmse+I
NTgLLJa82R/ba5XiZKPnBQJVTMDEU1kvyR1s9hG8Dg45PkXwjWr4FI9zFK/IA0vKNGMvyUjqYRrk
1R1AldP/N7iSseuQbvTQc/LAty/EkSnpvYaoJcKpfLwIK7u1PuDJ2ZA9ZB5FCjUN1eSTpJk4cFIO
qJGgjrkkg8DnDA9DR9pij5sIbwNVRvN5ovP5g98J0tm5d4zXGmp3ZMoC4sfPLzGdJvAZgVEv/zqP
O2N8m4XwNQvWdxIa8SuNQzdyhwEed65gs5n5HUpVedz5JHK/n/OBxfdb+eXRgrEi0Vzt7znoNcgN
d+kv8oNUvuuC8dXQkpAsAW9yyZK9GpnUAKacXIM31uhrITUkgsxmoljthLcETP92N26uSiBXi54o
x+lnNStRQ+B7LjSEZaQrdIbFSuUoOOOj3aGJiB/tg6tSmp/KLI2vcGdXYWx2P9i3RdKy39YJttJF
AoRu3iciKE8OO3mRV9NLn/YLlhSVNXWDhRilY1PsrcnoaEWrGbXUU2aQU1d3GLtuaLJMzTD1CSVS
rwdaryELCTjZml1pG+u5bCcrqDDEgC/d4lsp3LxzYCvwTVXLNnnQXftfxGo9Ueo3tKPYa3g9IT09
AueEhUqfsrRn2IW0/yRkZMH2AA2B3H0e4BUhP4XQeuEx40NZC08FC2wLTXEEG8MD83IKoU7F/aUr
HXOaJYyjCj1a4PWIzxn91dmVO+0itke6/wlcWLaJlfItiiIvBbVMBgm17FYpTRV63BSHQvc2WYUR
wZ6ou6gaaqIepWfnBIlGULeaiJkMFGZVBhl0hjmn9vCK+JuwrLecDMvWmXPtE7JSyYIak8GAjAP0
6/6nLd/8e3LGYnmXRuPIwAzkAeeQ6xolQIdKMheXYCHucOchC96RIGZf2bwcIz+jafCi3jQc5v1L
DpCQXnSSqEUlA+lFlEO4gNBTQJoyZui+9eBoR0FN+Dbkncwkxyv9Fmtf3BHOxQO0T3bOfSHQaUFc
PUFlZ3zIZzShXVUv5G42+hIKViU8G2TzYcHGIcKj3YA/4ur0q4PJ7+5lY0jRB4AHeQf7VRP9eTVG
58WWyxf5LBtl++MRCa8kK/UTFh+MtVQgKO2FSbvuHdjkdiSlodg02G9N+spO/qWmnb0vj8SfTziZ
jIU7MqryDn3Bd7aIFr1mbLoej1f0xHB8hxfYiTbykRPeFGLdm9RO6AoGEE5WpW5uZX2YIdyLFLVy
rXgw+x939cAXLVe9UupiLEDSAN5ClcpJ8EVWcR/hI0alkjoj5r+GgDsXtbWHNgnhYElME+Ye41Qn
Pjbwaaesaqb0adrfii1jAeXRMqw6I8+h8UNSPh3FJLrL1p2MwlFG8M128T1MHcH6wzJkWA8WBbYm
ffPjRonyG/p8cArrsQk6UXdZ1XPpRoI5kRLUedCHHhdeOlUdAI5vXTvfVLxYpP2gYSMNnJ8zNZc4
B02eKcOLBqNRUYmLWJD/sUcJik/0uE034KcNvFmGEqvEOWaMCtfczM5sYH+SpmwNpK6qQrsBNBTh
joTS7SrhcX1jcUI6gR4KTTVjX7i6LdAcj0XXwuyX/4TtO33rs6WWVP13Ra1B+D/jPdkPwxs2kyZt
/dyA/Vyh4Gm5hwhpu+iH9AZER24nki8g7oh+kLspkObzLx8uOH7815wwNLjrk1mWTg8qPGRRXxre
o+CKWhbyqblCIu7rnyNZRVM5z8udUoGfWMpHpt1wfEZtHI27gK97s95gx2FmIORQeTthQajhc8nh
EJyrB2k3VXkbfWGIC+NpaG+roTmT6HCR3g+C0epaL4dI+67m9DXUF1N4CIQbW6klL9qmfOW5BBEY
VuEcOX+2mg2L5fyUJ9dyuNpcPwOA/asVMMvVef43sXx8NwvEItL1XP9ZLqYXVceZAZ1NxwBX8t66
srJoVGbTY2qvxsBuGkrhj+rPM6SeeAEHsNV4lRvsN+NulwRpCC7gVR7tUp4lt8Bl2mX1paXS5aRr
KHRuvf3inLP8wqphBDhkW80MP5R2OMhtAmShwvNFYEJLfdb5ymgbuilCpG6/6p+2oaL4AbCQ+SW6
CchBkz21RyHCHNRvC/+Sa08Zv1ZYxLmzhrDVIhqE4GY2R1Ye34J+zrkBPnSXzjfb4Bb2Hoqetptz
AULvAwkfIXutVJ3gIDU1hrwm+NOWX/c/dm4pbOGqh/KD9Hlkm96BM8yYKdlmkYHfC8gmishSBzvj
2FhskF5dNH1XsXKChvz9f3Uh0rUeIKJi4x6UwPinwKduYfWi+bsbYmN21UGV2gO8OeXwySmBGxBz
EQxMgpdduWSZemlWiuxleY9fq8h89iO2rkbhhMZRF8m0hP4xJbViLmQgJXAPB2CXP0/EZV/4E+Ap
tUmhZMZYTaVi0WfW5l3tvXqgp7GZUaUaPN/xE3xrHCumAqsKtscBzMWGJY0BfpAUWhER1UxOqNMJ
cQ7WxHV6CNawF/VFldWb5eOFNRuSi0EkZtEmM258cCJKbwpETjyYeKVufDMrQu/6VSW4TsEFtKib
6sTlHPmNDoJTnGNni9hMDGF71BTnI56qkabhBZPtF3qgCHM1BCphH7JLQOYXhr6CymLezQq3qEsb
jsdaiBE9T9wp890bWz/BMwp6c1UAAsMK+XiCEOb7UxWBCv7KyhD5N82PZa7WIfRS32QWnOEdwX8G
hDaIWIRFnKbP4KFt+2LcZZUdcI1Wue22eSnZSCjbzlc9AqcTlgIXpTyC6b1HFi6zkIuEmfJfz48i
CHTkajhhVpIPOZ1ZfQTWgnt69R7MN+5Jm7Q1LAcjCmOHMldey4rD3EmmiUqUvXHLLIPKiqrsCLRj
aIjFAuS+kNKM8kA+k/pIOR/HZaUqVZx/FcYzhbcdMkVjG8kJRieAS3M2Fvuuy3R/3bCus7cFoOYI
rZtOP8a7HIL8PdhAD2pmxOlFwWDNhkoO1A2Tp0u7pOCMR1DPF+QfvOGAJIVnf4Qmhg8wPwVfTIKv
lUsOSwsx9VN94yNLrN6N1UZwroBNbN3a4icXpYVM891pPWCGIjF8BpBN7H4I0O5cc7WH+fJxC3zZ
oAzMlTdHVklS9c/vFqPJLjmuwdPX9yIZ8Wb2P0g+u42f/UfNalbPwTq/wcuHNAORXYGkXYWsMZIx
iE1ARqHpRLRZ6G6VRdi05DwmyxrEJahx5CrKb+erpglPcAMJc6lh/gZ9r8OndbwJn1zVZDTwBMpy
dJSCKOR7191gxnLftF0y9AMWwRJBZh3k3zONghScJW3scx422CaJbHqyJSrLuxSDceh+3ALorbmH
lwQvbC2QBMWIAmwUCb3/6KdaHSagsyKMai+HCdUSLxmfFy2nrUw26PsyriHHE9k73NE9a1rsM7Ra
hrdMvnrNaszQ/5aLJSf17fk29dniFrHwx8CqyqOUIp/onfzM7gPU17xm5J6g9lA/TWKX/RyczCdF
hDdgxDSQE4NewfImIPYve863Oevx9jFgcGzGNIqBCfrluJV4fC77RHALVoTdVqmCEqgwbVQz6Cz0
ivSHzjnlKImszrj1/RJ+DoBp3wjUA6j+soKVxB5Bq03lLH0vP7A9rz4nOrCCxuWlwMVxvbhXqE5q
WI/5QnL0m1F9wOYk4+Rlv8nVHkFfi+THNsizht83lRUBWYpb4GbtArpacamIgWYCkZmLhh0V8v7f
/rpkU9z6X2JulFSu8VBR5foqidKjTUgP6r0cdNxSDIvNMQ7V3DFx5mwRw1GOs02DTFZGzs0xtoWA
aJopWoI6VwO23swupxEtQkH0F6ktTgZpC30zqbB59O84QWJW6zBTZv0pc0SzpdVjTD6v+0o8PD76
HYQHmzUNctBCV4AhyCqjV1fHLLEjpZHU112Odd+MZrskxu5mk5GLV8j3rnlENr/Uhska9e1ARyW6
nb9K6EhbAaiC34ZgYNh8PWu84iOp9wwzVkLYHgcxUrYF1098eYa3TdkBfPoa8oShT7MusaIypjwc
ztGqvV4yLKRy/z+ydkOhd1zS27pHsYyqR8TxOcDvk6NbL0Stjc9m1I3Bl3/Eb3KHb1c0iL14h8YA
gReIurfsxpbjSmAooYLHA46qnBwxJyOgY+yyHlznlxRflyhIIKAOXwW64+wdK0K+LkLPWiGw1IwJ
wr/K2v8eCTZK9AGnikbISoWmzZFiuJ5T7tzXdKw22sWODpzjXhbEOWW7lnNzYnE4SOy7oNpMz4lS
I6VDPdiLD25ImTNiTpGf9yaCEk2jQcQUig+BQLIJo2jp8Lc1ngtlhTUULpMipkf+MZ/llhvq4DKx
x52tA+tqgB/jXbBzvITt7E4A/NX9siVCDNdLVkrVtN+z5GvOuytIpXPwQKf5/kAJeooQqCwJRgpg
WqfqmHwvVBtaULsnImjspdI8u0wR6/iqfmygUdtkksWokPySi47nvDwjDMvVvh8gWraDkdf1m1w/
M5CAVpN8Hhtp0ENotOyiDay+fqfW7FE5WkZDEa4d/2yzcna923HJogMJB2dYjlIEhpmNuj++Aym9
b/DeUq8rleAAawpOiIB2jiL+UToXjkXJF0BwNlK3l1BhWbtJm9EX8Y4FauF9PdLsUAZHEbmmKmfI
63xwo63/bI7rnPJgbDouZjuG7HXRmickOTJQe9nocDV7oBPGk6pXn++w9RaJMc3rEuuX9KMLie1T
mBrXVFPqGqkU3hm68xS+dPhAucyRKJyEoP0AqsfW2z5K50YU+rIr/3hDFwSojCNUECILL0x3mo4j
/hH8kJFV5u3NtZ5LzJIucsRsu+iG9/hNv8on7EdPusIY4hYiJnPnFRwtoHW8N0HbCFYWpr6tpmS5
ZPv1jWqZfr9rsuM3yarhirA5dM0rOoIYUhm6TAJYwDiJIUPVGL/OMsWl4VjlN3r4DgTQreZdP3Eg
CgeA3KPitS+GjvIw0PWEGF0P0XMO5SqNVU8nCUzqKlj1NO/WmjX4Aqs76E7xNR5kS0ogC26Q6u0d
GA3vFG8JztrC09ZRyifh1RbU8bXLKWl7ZWq1lG2oxTA7Kt7sxokA36ZWxWVoQk4CWjQqu2bYH0LA
5tx7uG8wHRFHCmegbabSQkXqUkjBa2XthQmruwEaqp1C7VkKeb3O3+8mCZNLQ1Kvhg2Iyx4vIWqE
P7f3EyZQ0PyDrZrxHnAT0F3z6HNhB7ufKZ0tziXHIi+X2QweYWBXyxKTNvOU5RlGAnoelxG7Um65
kab/zkIVZZWS8oGTHTeR0FMMgowq1YfD3pGSKsLgfC8PW22Grt+d2YyB/YOiMRj8+duPVCSkJ1KI
CI5Ye50I94eQ2oXlqsHyaMRRy8jgL6RgMLE2DyzTRmDH/4TWyowyKI3HWsMKFNn3k+RZAWim+JqI
yNbNuG9z8Kv+qkZ/UMqDpguu+9diG4ZhuvRdU5JVBWPpxgWGC1ZOAgm4hiHxVGhTrcjtaKL7t6z4
N5nbaEyCG+RJzKxrqgbuZwlP5b1Wvocu5n517pYQPy/45CmvG8lZZ96w5v+aq/C4QRYF8EJsowef
87E4velKfk2kqbsrHW3rY0Pl7Obe2UfHxC2ILvfGNB+m3uUoUtVL1hYyURbCp5jVeojr7gWo2+J/
ySJVYhU+xneUj+Nv6Ek/2pfucfKY5CLrdJMzOiI1tazXyD622t7s7vFePNT6syDua8QW9CPw5/ko
h0Kg2sd82NhF5rPxPny6WnM+N8EvbRVH0ZIT1FzITzdawFQQA3S7AUjVjh9afRpfYQcCeVzyV1xu
aHyyMU+f5r70MF1v1gBZqccUm6cuAS+yfuRuFUe7bCjRD+x40s4/UZiUaxteCndnt1jZVJGEROHn
bqxa8Mi2J+CddBqIvx7wVyYxmZT0Y+rS5z4LwDtWQ/Mtw8oC0EhWLp5j9pRIf8ag+tWl2FlT1tCS
Fn7DbYk378IlAWv23AaFM+XOXs7W5TRglaFZcn92AGHPD0V0tECRFk0oYNKSS7M5twsCXIuTcX1x
B9nN9RaE0uu7zP3maet/k6AZT/5yklPSJXv+TMsArcpmGMg9fIX+cuKk1tijbXcFZ8mfM2WpfhN+
omZfH2l4Bg4NEmRFoU6R1A63aD8Y428Tem0gE9dZUaj3eHWUKpbn8Gm0r8r0wzRizAdSALATMYyG
XwXBExPe08A5x4XGruFSMePwOaMjt1foWzu0N+GHdtnVLosi7fxLCnL79Dcj9RukE5AJGLDggqzh
RTs5zn8I8di9kVwP3axqthixkBZAzzK8wPYVdjUBFD8fm+kJj4xj2nJAIKSDI92iREbnZADO3oMa
gFZpIEac/LA+n/7vIWnPxUUfcEMzDVbLdQsYRhnsiTqlNw57DRIyr6oVHVes35YNB4gyQL7n2DTJ
h3NJu3eI3XjrJ3eY5Caway4CYVUE+waz3Wet0f08V0nn2M0sdu7VWb6IJjgrCSuRkhnSq3TKWJ5s
SAMo21aAIiJpAdqFq7dvkXNI9Zil5bkVIb3MJ61IdSQtWPMb2iVk3uks5GG26VhcUlmxnP68hQpU
HDRY1M+Fuhnmob2/P+8m4NWyd3UmMgYdHP6yFEk74cXPrA1p3LNM6lz4QMeABX5EDFhp2TgyAbu2
Z2JCg3whACs6yza4Y3i9P9j5cZSi0KwAVU9jfAd9HiUmU//K8dIwOkMYf7q4Jmn2o+oJxOp+WCQe
StWblWeHZ4ExfXSSvBMpkPQBAw26ZCtxc/iuXZjp6CYa0JsdZCINdnRkGIJA01vXrNj7Rmu5WpUL
yCQiKV8Yvylj4w8EDe7ltcMgCLEkuxCtatcdBBp2KQrAFnzd8sAkpjITOo4oqx/nrJnJLknRDigF
l2UdPycaMOQJSdIGYdBzt43qGGbMAdUJQCOdFhKAKUsXYzUHez4HMQdrntBEUNzNaAJ4uNRKem1A
NwIxSsLhzFI1aI3sKLm2d5nSh7FkOa4e+h0WKGbUK+o/jzWGia18adjEMKzbXEAB7st1gf7FJxWJ
uI2pwyjyNzq8ZjoiqokCvpmjFcRBtSC2PLA1J+9zgbb/zPt6HkQfs/spE0ls5J3GPUTGc8PGlePT
N+72y8Ja9o6gtkT8ddAYRnW6VBLHKik0K9axx/81WELLaFLh8H9Hq+g1pEwHLfmACMcHVXHCy4zL
NjmJmWKUNKigshF+aca9aR+rBxtrHesAROVcj5bi9gizdQDi+JepyPeN20/blChQ9OsZ06zarP1O
zimTJHvsn9LYnJC5mDZc167adV/D8d5Anp1UkJq+TmxgzFuZwHqPgMH854W60LMRbvHGzJ5QXlqL
/v+KWkDAPMa5+wDM5hE4p/lLWwtLnOJgvxD2Lx8giylMSFODc4H0JSLpxjHhwwBMhWrX+WT7foWj
tiJvgps2/JXDduqz0UjDZEU0kuVpeSTXAkhVo76KkKlvIHqQW8mSka24muA5buaDaM+A0XzSm+Wk
gk2C/1OJXTA0OGAAGH5Z/BjZpWp4HizHRoZGaCzFVzhZkWkXud9l77qbkh+GsIlNeT5XZrOL0cJp
9rGl4/1CDu7/kkzhvvNgM6lTamat7SNKzlKNRt+d317vI+mU3hdPSY8KM3VK7DdX0E/c2J04Ce+L
Z5IwB9FsxyJJXD4fnkkqTdDC7TvTA4PuGQfwefcuoxRVHvaeKi9kF3P5nc3JiXJWfOji/ICmR7nf
nF2uHZpxLMXKc2bF/cmNFI5xG1IyLCnRWHX9lQD/CYpXGL5Ey2cZcur18mBeW77CzxDvFMjCovSW
2DaMKrYh9EwCi6K8tS3a6RhQNEEAnVnSCcEgN3w4soiayRv/LFIu44MRtHc0B2ZLK7GlVTWiKaEI
JsP/G3VnvfK/MHklrdg2dQJOq4aZcf40y1iMIhqbZRGvNzuFv6AtKpOghubmagP9BqxJte9JZgFB
IGKlETkSoqoMAEvEy/c7lxrmjyo8+QrhoXoMQT221cEQiAlpv8tWzElalSOPLO8KO2Zrw7qqG3iw
bW7+MNBgd8aRuv6+py/VyNMtLwP8FMYDrcEUlz1yJ2g+o54BCbLkqxhuYuyjfRqGWii3LUCMAQrp
NT+oqCxvx0nRz0cwjDseruirbT9ut4PLRIuVXl9TXX5jK0Dw64gSJPL57VfCuPmqlR/ljFY8g8W8
KcF9Untn8NL+fh2BTXe8vs0bouHC/QMJSVxtRoYVQS12O6AHx+osXA4HSjQEBNtaAJvq8RRtX6Jl
uhVo85EX1/6ISMyVy9bswQWZlm5AGnWcnDJozcMIkItlQ/O3Ows+17GC+m4ypxu/7vh4LCUQSF5I
u7TYIY80cmbBpBU++Areni90CRLhATGuX+JIyroWYk+eNiZgYAjE9DJm+6LbFEC69Sc7UCRVEaon
LRKSghdUp2oAD1ZP1410iiBL9+q+yNX/KR868W5j21OwwgKhf7SCm2Cco0pyCbHVTqGgZnebsBOC
YscD59He7CQuzWvtQcFak1HsdS9jtEmKfWZEfrBw22GWI1UL+fuglgWq5yRhmolPlFzJfWaCDWKH
Ury9qkLvHAh16ekThmE3nrdxOH7xqq9vvjc1kCGUOE716ar4pxD5QquLZUm+SOeGheP2bgCE0Xbu
EqIxhlNsoraUotlNjymj+zjKPF/DPK4iGcB+YPu27vjUVXvrG/Ei/zUxEwxlSuCoh5uJ6EfhK4TO
jkk1Z+2nBMx7V7DNUPRWZSYAR/WUVm5GHKDnueSDpwh08SVjcc3qTbVqzb9dPshpR0iyqEytG6+G
Zr8CrOFdtzTXxa8+pLTcZFsfcqg3+Y/CNhZbi8B6eklTgdkWz4UC9n9TvfNx9mR1bdluWCnpaOPU
aQ8pxdufTejwdhUbAzqsdmTDt660nao0/iw+5en/6JVecxdwXVcXqN9KAZJWeL6p9TjVlgFB21Uz
VlToZAGExLiVR6IG0LmC08lca6LGYpaarjYufoZkUP1/e2EB5d0TYPOTNlOULi39lqAlVXQSEo8d
eKcQ9/4LFPmeyV/VWSMzHPvbtZQzdfURPfkfpvOdJ3jx9q7SIDXLz6LKrVxS2gPUo3EAVLSM0dd5
2erzMfFwJhw2uVi+JELFbwg7ee5r60u1z6WwO8Oz9Wh83q/u4XcgYvD1PsofVAtkyGdTF/zdAHR1
nhmaBxFUMmPCeEiuiP7Yvemk3QnSDXQ5Tlzqi1lGSgel84J2Q7KQ+N/TXYBUwzyEBoxhoCwyYeRH
7dxgDmDYKqNmwwX1m9UpxC3PilqMpAKqc9ygghfBKhDXYiPv/Ie77vk/uTBMTg1kXe3VWIZEy45u
IZUiIhsjAz0YCHPICa35bEJeYgIPxBFm0Se2xqz1mG17j+4LIBP70PqliO8XPcmyvYir9qU1oN5S
CiCb6PZm8F4wtcbqoBBOMOpAZrVKAI+gsYv0DFnuAoG3JJfZ5CmxPcMT02S/HI/bdQbsebKv4/kw
OAabJuXu4TTHs/nLv547BmxtffrB7TX9AhID8YuNc5dc+16E0jo0b8hAWAZyv5TktO/bZJmG5zHi
T0gJyq/N/gCO+R/A3tC+gBQZcXR4wEiXZTZqp7ZWychvvonwPPRnZl8kRiRxCh4IVQkHYyLd+df8
/trjK7wsa/+pfbm4X5kXDGZ1vUBEj6UtBgihxI6KWjQ5YTFU6PraNTNkrRGlZir6OiHVT36OrRBD
KVNdHb+k7v9SJaGMsvA1WxQan4YR/uW+r7FOzrorNjJcZd7A4YQZx9l7i8Mo5yVr4n1kQna0AfZ3
jdPciz3LHsfC8jMP0qQv01Xk3FuVZZBZ6Xn+fogBuQrX7cAcsr4EpFhurakfN04imr+GI/l9/53C
IXhHFqD+Ri8gn3klPkoua4ciUTkLesUEpw+yJcmRm+nG/LXg5EPv8VWOqmlxQgEjHgxERJUcDO5c
McA9Qk1h/vPyak/1Lui2124PFrCki+ahUCcMrLOqb3onUPx/5bxar2ONHndmQJSEWwTuVIwRyrE1
MUkoaq1hlAT8/Y4g4XrTWGFg8mOi6vkU+V8I3dhRc90xj1nUjM1rcQ3LGSQv/M/CATfs3GDitYqi
uSjrOMQdQDPen1nwjzEDSXNDGrBf7NU/KVWcgw4HjaMRKqf6lYgG+Qhkt8Sz5JXK1mLkIPXj+xWq
NQ7nR5+ci7nP+tPOyiOsabgt4nTuAKs8g8l4q62DatuknLUSOrY0W12V91iyFgaS4oXcIKZKKzwN
VXyFAsum7K3ciMxjdTT4/LLeQDi25KSB36Xdh2iXHARKfQtwpaG5OdV+pL7m+IsWC4gY5VOyKKzX
AUGIDH8aAQ4zofRdJ/UIzByNayUqZZSFKa3XmYAkh6nIKXnH7InEakJG1sHiKIcv5OiqROuurCKj
d14yovqCTkgPnRONHRCTTuwaQi+pD2Cx3qslzTQrUasLsuLElv+5IArKB5Z4AcrRxnDXmIkctvcp
thmvI1NClhiodHNvtY/JFlErTFxV5OYM8Jxh8fTu/PAqtjaw2CfiVpURn/vzz6e5oBrN183vhFsA
5LPRChkNnuNVVO2Ixgh9jaKaIQKT0s9KMKChylEYkCyh854NxXHzVOCVijrWXdrEMhz1lcJYuQeD
2w9NSrT4zdCAUyN0lVKcevBpPxoKNLttuACWKjfFVKZ3luCeZfwXNTHWtSxRbpi1qqv7WjCxJIMp
sGjAiAA7avHd3z6sq77i7h2yH3oyQdJX2IJLMz9A81h5y8d2Zm5xMA/gwx6oah4FpsBR0fL7Lisx
6SPKlLFW4UY1LvNPhXPNfV0QbAF2DqsKU6f6h6kt85iTF9nsaVkU93ui3ItsPmZrVnTFhZcKpPNw
GEQTqqfyUoxJKXbsbmWn561rDdrdv5TCyAZbXgKMTC2Mdu9j/rrg8fLrcuX+SXTqz/Jt+3GpxHv8
6fS9qkWif4ONNYW1P4vAc36VjV3EFooeUH0XoPqCo50EtI3tBgeFGqeSntX/YPNLGYxXsWFNkRNh
XspgflV7apR/D2k9sLaSTVGFx8o/ycsTPK7bADZvEy2syMa91Y/zVk6LtmEnsLvUKXC8m07gFcai
lIWBelxg6S3tBvpjIRsVz6UlxkbVuv/s6OA1akgQxd/dtkgdzYvCz8JFAfxhZrcK8seKUnzKVKWC
GhYwdSwU8P29d8Xgffa235Kf6WRul9M0z2IJm8sQHLpPc50FrLys9XNJq3Qno3IzFmEi+Rjb5OrD
AbMv1Y/nYbED5KyRiesL4v3Dy67zQyTk0OOL9iy5wyTU0JkxblIWxrcJQpWj7TwhIECeVwgVoIkC
lc8sgXX6BOfvXrMWWJugRaqcLW9A8P1nOM2Jz6ybb+HvlGKvZSzn32HU8216r1qKYmTwKYyr9kXU
vUHzaambVdiPUSpXU4JzZ3MgbQUY4jgylubvPVLy5hbo0A7tXFvk1B+yckuGSYJrwcWpexa18GZz
WsmSwB86VuPZM2kU+RNv8Fet0r68TVW5/m4VEhl/wgpaSNoZBL9gCsn0xJSVBIdJc5PqyBn5e/1u
0HM4DLkWX8y1af7RLWYyHqKzk1eXYjRxoBzJ56Cg91pkMrtA8Y03VXX6kg64Bd/rbKAO/0PbflyX
d4VEoYmhgM01CYnmSVnsaE5A6Tqq5TrtCtembkZBgjGMXG97PM+ElOnjwpsAGQBXai1j++vcz6PI
jBbldM7ozVoX9chSTMQeIvNU4QgB+od6enZwyswZoXrNMt1gOSb5XPde4E4aBqk1VOaWzVkvca43
mocMzRXXq7h97o7/91NNmn2MnirG/4ju4K24rDWCZu4TXqUWQ4q8p4RKQSjneZlVAeDzYq74gmvr
aHaJaQMZvNflL1vbVBNksfzuCQiuvEJvcGMc2seTMyY5yDHSgqT1HwTDrMA0gJ6Asj78zWKM5VVY
ppwwQUfXU+aomtC77+a7EU68JNAth284S9j98WRDONTI90UFVuKz1VVX9brxMNVhGAxox9bY7Tgp
u0CgKTLHSN5rc1xE/aSsKerdsMpEiZ1kTG/Lp4OVyPu/D+B7Ph0XwO7ysXUCsvmDCtwirI2A5J7Y
iE8X6sRmyd01eMlw20/12+OejfTE3CuFlemVBgjLhXmJQvnL8sFqK45gAEqjJtJeG4UycuTQ2ruG
muedY54C5zaFu9tDTtcSeJkNW5bfrk6zGtfwrygj/JZcAB4Z1LFi/osrTt1lngkK0lEGThSPEKcv
fqnSO77iN02xgIfF2QEdH+xEJ3wkJBypnzNHMyk33rtePwjMdMnWZOyrCsSaiWCmYzQ8C/hqxyAh
YK0O9vGPIkpaNVt/hk2kWRSMZKd2roHwXTpJYN9T3eKWU5BFDIiPjtoYde6i9QEsZKDBDlSMwajk
8gxqFiv+6ZuMcl5dyxDVaebeZR9Q+V+jNN5U7F9fiHbPpvkddF5QBdiJI+smR+aVqBJskkiep/FU
RsttpaOIfPa9rpfXc6K0JSEQUjAS0UzO/l9D79m4rbOyIqeJfccZYmqOn40OT5gpHIduCBXlPsRC
JY1u1RRo+zLtu4Y7ec6lPDfaDOtyrXDPCb+W/7UTibKdecCHNAaXZz9l5Gv3ip3A4BLP+dN0M+iS
DEMeAI5f3eRCmJKCbXpENcnQlrsmMHAm4qHYQ3e/d2bUovrW5tLAmXBaM1nqxocQyXwNcq94OUjI
IhgdiknAGWQAT+E2ojGVyOPDmy+PfZX6EZVg7rVXr9s7jwzEXxjt2lD1SPauEFn6ezGp4lCsT+Rg
96QMjQrTzEqMIqUQdcjxbmi3hLsOlrBtCbMZ9HQ+JM8lEUlgDr2yRp8ASiWWoJqIWkBjQE1k5y66
64FMWRpqe8EhgucRVClg8xvyKjf4bcejd9v8JCBmWriNVQkRaTrnsrQeLzlIwqFZB6zwlTC13R3S
z9AWjZZJe33aaPhVGdrpysOHcAHzO3y3Js0n9/uIUjX12kiqJGD6AbEaGaneJYSTsMU2o2WRGc7z
tyQQIaCQRyWINywRz7+qHlBu8o9f8/GJdZOFV1ar7+vqo2qyIO4DhsWOfMj/Vga3z0BurA8/V1iq
PxTZl3QNsUGZnB25bpePaIETZpZb3k1DlgtMO5jL1okjsBtPFUZE0pxRNpty6sx5zPtgXcjL42SN
dHzmyD18KgtsifbSp5lEGVtXV+kXmXdcKXTWxuMboNi4/QUvCfBd/JoJq1fF3yRqoiXlVKWTlRNx
ZRCXPEjrnsUQ2ET8HSTf5IpDYvheTwx4A+4xWWaCTrSFGSbqYdVGnnBqOau+9kcAWkuDShZqHKmp
zMmSKedxHVmz8Gf4gmEwgz8SHHq0dL/92xsD80UPzDVYtxFoS8O16G2GbACnUflk5vSnt80O7oiC
je89XsgtDwddy1v+0jkVbqaYX2xBq5c7BCZNkcLcz2L05Jbbmo/Em706aOnBhhY5W1sSMpxn5q2i
PaY+/A1H+viI7ntLnYO7ONHvmw5Epx1ok7z90pivZ83yC5wMcaOh9leabDccsDSeNdnBnccmPMN7
XRRrOeYprzEN1bIdhaEXp/9zWjbrZCETtGKURqSJnHcO226Zq2osgXjfP3eZq34gpRdWtMMbBbK1
VISDrIHX/ky0W5HEF/aU5yHK8VthqG4Fk27yfOPBrZzRRhUCL+m0G9RKmtAZlnqrQR0vLZjDZpzL
v0grQ6PoiAI8irckLmp9SdQvCNhZ6VB+ruBnftVZzTkfdrHT0G/ZZTgukRDJtLGcsiIo/EtMVCVc
OmYqMDAgQHhMzt7OmtWSgFQ4bGBnaI0RCBIC/op4rhQFrOn5eK95Gn2KglcJC0EDszPhhvO07Qm0
VB1aOmop7pzeBbuvSlvTHSlJqNudEdXOToDej14Tj9kFh0gPkW3skHknk1R8RKhuCR1BXk+vnuAj
Rhwmoots9zJY7heNfK369khMkajJKfkwnituRcbLmPUMVZil5p5C9zzRN/jZE7fh67Z4Iz/Xbezv
hIlL4Gw9lTtI9g00EQ2OiALacftY/rChaX3Nmnec0Tr77S/Du+UMmINV5aWbpo2bn44MVYUfP2Tq
z+hdoeQo2xVqgw0s8yIOXl+xyhJv7sjVmAqvcZr4wdf2GM012rw4mN4YXYXzK5RDjh3ilvx0IAmg
RDekhb8aNO5+wr2/p7y7mmaVkczw2ryRbAumSiB/DOyLwaN2FAcw/amRDfZWUk+zahouKvcYoDUy
R0GAy46D+jmzaBcCoyltdbDj5hBP4oLsb4x2bsBUYbDQiUBhhXk93qkaLUhngYkNB4QvtBIefuQv
CZ9LX0F/Xn5R2dzuDzdbjebfuTp+tWJhWNzORCHNFpDiSpDTHMIknFe99/N3m7kNJOT21qBdtoDO
v6hdDtOJxjSZ2GW3CR4z1ivda7pBSwBn7L0L2iIEf7Ftflf6ianHmWZnF6e5j/gevGIlJvYkathu
aEpXeXMJwSSnq+a7rmffBYizC4/RM2aMxWfDtQXJqTWidaINeQHWrVhWIgfCtTpc4WT1I2sSuJB/
zDcyGpVj3hObm4QuMvyRKwBsB/6xVjOBVcaW19m5VoWoY4FkavrdIs3+yIZG5JhEGbA2spC/4NMH
83w+peV2wpe+5FQshnMepQiKIBN63ine9ZknKEItcVc1JIgLf26WS35ZTSrVtBia416zDd4Jlag+
XbiHa4X8jTzKZPmDffVQ0WlM95PTg9I+Mt+UwliKyqpdllgrA9rnRd1+UiwiUu7iJjbYrrMvDA+d
svzz29bBh7/WcLviWNt1P5t6wxj6OFyn9BtcS/rKO7rx1vhHUrovARltqR5jdmsV9Pa41c4NZ9Sh
7mR/HIkqlYLy+x6JOHJ4cfXwsodScQwWhZKlc7qJ97lOc4khvd3aCR3lZSBEv/FaZakQJEfE++jG
4n8QCHlFfimA5uVcuDPHQyNfC2K8G1HE7wQHkVpY5rriZoQeDajSjg4qnt8HAudY7qtuKwj2aCoX
ZcG4WYs0wmW0McUbRLky/7UAYdmj5Ar2PjG/15KLmTN8TnIdzxigtc1ururxHgujEPY3SVvWREAU
0RdvD5Rgb0vyLHeTcFpC/+0vH9U8X3bsChheX4jIugVI4qUZvhNGlZD857TiQsKLjw/y3H3kbY2V
lZ/PB6yIAHSOG48KkuDw94KCuhPYSppVkkght8wIBTeBfZ+r4R5LajjlXCkwdCcLUwgHDVOHAVwh
/tS78GujXLZ8nVQLjV6kJm8gUvoS1iyEIXRzJCRxsttzyFOXZQWpgo2vwxLDREE8RmOsUDAm3j7Z
/fgrjBz+KhoyuHjkY0l3Q3CP7dxdR8r82bRnvKRusrxbbS18kuAiOuiuL83gpt1C8Ya+aawiF+N2
vT4UMhvjLOSc3sPjSYM/Hx+KpZA+ZqLGlZxe4B0A2LeAj7LJNeow//eA2jqF49prGd42163xcr3X
MjrH0Fy898TrKIjNtwUOJcjLad0sPsrih1MRcSNXbr/d6PHfEvvX8915ekuGLyZom5Ga+6SeZL49
FCLUwFcCwmVoVbWokHJvQsh/SjOgFEsdCEsIa6+yJMakGOwcCepRglBSjM33BpdMKxW5j8vq2+6Y
6pcQmGsVgqmbkn6m/pmjB7tp5KhKfq9HA2Ed5LhXJ6imHVuWU5Ome/SzjgWF5JUe02cc55iDtjWN
+I/n0v8QjVHCjxKSKxLETKRidWNFC27DkQBk/q7tRnlXSCR5VjlB0sRIVsS3zbU/G58n5bxczBag
g0pe9/J2Y9u72eyiXJm20uzXsPjLNU4SjK2a9ZNBN3HzsXvXKpq++ivxLvFwpx3CyMWUQZ+keULG
+T1cwS5ATSqV1d52TA0JdXYiurbWzemc9jr5Xi73WTC7fMtFH3dIB0rRRxbAVBVjyCX9jHoErbWJ
bLjCtw3h2i+E1TXMXfIdCSU9kt3ujYzXtdMLpz/3fgNObtwSEQlsZKSc+cxOaw97E10RO3PAA4P3
lcRiWZn0KG3ar4kCWlsYn3shashsHyaYaROR7BIs2esztLgdgf8QbtR4bc27rGPVgjWesOS7cy2F
Xia/tXaOvWRJmIUUJpQ8d4GkAoNBHK7Pnvt6KNFAhUtb5hOM7alxIFAbM9UM8mhAdKSd0ov0HaeG
F9rl6LsOt9yVc5PqrwnsGi/dkfl7+H1oTR8vTFGIB6gjruY5eQ3edB/N2/RYkfFhdiMW6dxUJCR+
JTK/92hJh59Q85CtIioH3OVH/q87NL11iNhohg+9gE8TFMBXzbD9QgMT2KU4iq5Hadz0fQhOt5iN
EJZ3RhBCsZOHF2W6t0m/ERuDUlfWFmNmpddiYrnLO1o5lQizcFBS3YFyMWDD0mbbP2tEEt0nwd+Z
Sl/vLcfquK8D4ubEFKGNuyQdvsRZa+djCagSBq5FF1TKqJuBPNzFrJL9NX3qr9r57uQjmQJwvhMt
ljIRJ5iKY7EPvq63sM4OlGI4Jvs4VJrhLSFsO6q1A1B+I6AOTP2w8SacjUR7CuKRVYDgcT/Q8xys
Dhk4jzKCiyWmu457m+UhAEEPoYSSsKd5eK2mVyM/2jlGIxN0KJyvdHya92iGfGb9LZx8gPHdvb8Q
v9CI9vFt0he9NpnARWrEUBHuIy/I0C/mmr70D8DTcR+dYKbbbZuBXK3A0SfljOgCYeHjVP9XL04U
Gmy+rTVtTwEopSm1zuZzbAhIbvO58QQzmQYrXFI0GH58WspEgDsKJPnkO/KffV35FEfMDENOFzXo
VGEH2JBxS9yW/s4U7M7QEgckv1V86RM2jpTlArJEtrMNwO7GJBMuJfag5/VkBeCPHGeKu4b7MzSw
/OGUh4WrgifEjGA1nwx0wI/A2DtdIxQhv+aCv6ABRppv2GrXS1qcqzFRhwoj4Ps1NwAKWCiNGfy9
ijMhr7X/UXbtdW+n/skHt9k8gtLGpAGzHM5TLjqLlqzpYKQxARj1iD6DmtnK7EoYZZfXQYzovGA7
PMfiswlUMc3y2MYUQ/PwCMVKTO03b6bLLdL/YgRq5fBcux/qJlpgCFw7ZFuim9vncQY3XpeW/uwJ
Qp23+nNIcj/52RnIuYIsS9O7p2In0NcG2NmItWaRYh9eX2sLsBbH0jdzAUorvXgJEbbGnrMMA40t
5C2/vk20P9w9vIszLX/aOc5BOUo4VHCQGuYc8kvCKhX7WZkJujp8E9L3bscUq79daEceuI79eNWs
3Ed4qwv6bLsYzgdXqszbAFknV6Fyzra2q++lF/iZWhXMhcqYx1ITXinj3qiolJQqNXmliLAS9vy0
9Nn0s4Qq+0cy1jmUHc9rSHHnQ+D0ReN+2SHjWrxjtAA9zPpzisxrBiE9NH71wMT0rwUXnpDchuv9
ygmFty2PicEW5dUjobQ7qWyVaK8/u6R5op8j8Jl58PdmzozmPUYYotw80QIgBHMzxKl4usa7J92Q
7hHNh92HVrt+NSdnCPBsvtBqG54bltmCt/AhJ4S/qv2jG5H/QZqLMWYm8y72htFnn/fj2YwigDEX
1Zh3LO9vlNth8bepMy0Hx7JDTY0oE+9rmkONQE7ZnufIaVEfCYQVvq95+ftlPpqoNR+n261E9ng4
5bKiAK1PsWTLyjiDKQ2DcLraWLrpEIQTmNdLVsHOOMAYWr+K6huPPJevcjCF4SaBKnNe1rckvctR
qS/xZjer5/xnYVpc7/Rk75cKtsLgCeuu2TkgyCpUsMJtpAFK+Z7Yug8bLV9/ItDAJIapZhm+zP06
re2xkDoDuRt0NrSxu2IAlISu0OHX+sAA0OxdijG3A2MSEwh2v3GOT9Gsz78rgSGK7WQFqev6nQT8
Ze7flMEfvjGB7aOVlnOfArjQ0BPmO3xFJE8pCP9Wq4o2gVKJQ+Yb+pMJUGBIfZD/nxsRZxPzhR8f
sjOsV1N87STJto1toxSLZak6oV48aFNzJlLnmnFhsrmNalnwog+yPqHqT0/37cqOWRdAMhIZhIM/
LxZwPWIGhMcOAZeI6mIs0YyNhx1l0PcyC+hUU3cs7KGyry4HIqC/IqD+oDV2NmMQ50ZKttUvpLJ7
gtmIbFr2ooIXdK0NmYS3WoGTTtXsYB+GGQP/xtGsqR35a9SWSlbHXnfdt8zp6EiAHpgHZHimfbX1
txQBHsbD1/zYnxrKLpvV7yGeZ+gT7zPlonSZEAkf16EOYaoLTIpVwuIn5CGiUeG3e+kO2ob1NH5G
QkRBRiC6qFovjHOToMYBuHHWZXx+AtnoRBlqwE+Upn+cvaDoOtTADeE71Oyv5wkvQyaAasgbyhrQ
wYk2Y7nJKmySV1b912T7XkfYTcjZoMEbIpvj+jkxfNrGp/NRxqPulQriEvVcccLcEmMbP9DwNKSx
spF3ftnqZ9Vn2t9fpAcOxDKuN/9i/YGqGSmXYPN2yTDD5BhJQWiql638o0VAeC5KdyMDNd0zXWCw
bcOn6oVUF/REpqexxRAhz2f8XzEO0CLObNwcSG+y0o0iOLHY1oY6Rl9eMQADomQi29X9uRePOlxR
bvHze2GywLcvAcWupFQQIEU4yGFt0IVISxAUej9C5wCt0lYmf5JJoVMp89L0CyPoV1c4NYH77nZK
Csp9EvSWtTyVw8emSC/vII5+jlaJfDKjA1YX/ZX6MS4gwTgIqIZPSJWzrGB0MhEM9/Wsn5XjFf3t
3qvIWAl8kYkuv6MB0HMLtB3rQHm+JbbYoEumJ2oNKLLidDliqMNYFKNRLP8Ius0VdciKPxKXuSRF
sAbT4ILgjl1bg5y8rw/14A7NYkzO4spxaIfW+2rVWhGdCTnnrQnlK/G+D00C7a/cskdsKgVmBt24
KYyaXIlStUC8mowDkG9EJSB86RVAbQN9e5Ro5pT8GipxmCiTjQ7IOkvDoOXrdzoYjnyljnBesKRQ
HsFsSkNrO9k++NKeW/40pwXRtQG4gWbUTFSePJo9MOpDN0oYgscLY20bOHVzfuVXev3ULQ28KwSB
b5Is6OJR4HIljlUhM3hFZihDAzTlVcRcPOZcc+6JBN74lGGzQRfguIElXSD+t3l3fxbduFGbc2xD
ZNsiKl//z6wnHNO6P3bZkZEvLbkmx6cJ2yW2ahgV38xu6jdriss7aRxL7MS+4aK4QikkBxIFdxre
v8Y4YL5/dyIQFDhzRX0K/vpvyZ4yH5u0XqCacKctPKI6xPJGT+PL+Da3l8svcoIqj+gZsvHCePyS
xW2YJPO5LxdpVKZGCVhkFaBkYHRxi7kKdWIdCdwPOYZcfQQKR2OBzRQzJfcynRx25rj8EKSY+YjZ
7CviYwBh0yEPZWPCju+TlFg/W4Qe6Zj8dnFGPzbqkgbot1OnnzMtW7H5gmnfTSPBg1uTLlqTF9fp
l8hG3CaSh1drpzRbiSS6yeGCVDANoU4T65KBsqJrlKdheue+bSNnyOS6wFOyl426aQAvBh4+2XjV
xyyyrnWdQD44X5ENLETOF2Qmz/nrTFQlcNH6jFh3tWctN3P9GdRkFejQWp30XNSnqsSINmeBtxdJ
nLG7UAXFwAFA4K6LQKqprcJjFg6OzckBtq7KtgYTadq8Z1nz4f6VXMAmH0bZjkxwfAFBmPX/Vi8h
wGgKpxzqgQYvBX/+nrNOedBDQ/COoTyIW5ONZ+qzE0c7Uan9ADmS87fGlnbdCwC4iO0YVfcP133i
kb1olmjxF+RrTJZz38gGm4txwAYH1rV24tlY53dpphzaBze9+QfDWnoGNwkG/nmu457dsaflWwQo
b/vMQL359GSMN/9oIOemrupkcn+Vujm41o5Gfk7+wh2BSVOPoK8cnDiZmyeDOM/upzka6QYGJsB7
Rf9zbicCLAG0zNqDvGsrgEWf9zRBOFoQWCTeDMfa1FXUMWng5CVX48CHetzruMocO4YHGY7PrNSt
/9EhiDChHW3ZoW+yEXOawG8+OVHNnncyUwOEfjVbR9sFuK61zXfSW8EB0/SnAQuXQKmCB4uDzF5G
iJKjldU1H+yIR1BlI+I6LrcOyFDE9ADER4/aq7fKofSwLs+UG/oVJY1q+5KXQKoWXu7mdmnCEbzZ
hiZ+wHOp34poo6Opsfe3laWrHycX8uf3v+zXNegAzgw7/YXhxmLrTQdlBOFJHKGGtZE799/kEHlT
uRTA75dnuMn2nJ4DoQfKXNu7j13Mxkwaq7pbwwLrAwruqZweBBKAZNK2MhNOIml8zInuJuwP1aRR
9Ufx7VOTFFTt81zPSZKaNQrPzboQlTNwQWfx89oQreR3CT7ndI8TxbvRKBnxvvFIKlv23/PWaf98
URI9WwGYbj0qCl2/+7mZKeU6DB8ALhJTLuJpXD04kiH8dvOlxzqRYhGM2OLZpUX4GNVgnzVLHwQa
RKsv+FcwkJfWKpZKdHufitPe88C2D3r+TLy5l0Ta7yLzdS+4AyPyv/jayG7R11Oa0MUGnVEgEORI
LLPmBNR5pkyBGzxFepiwZ3w30UWZlGiERxI2VQPUV1fdh8Jifu/OOiZwXOma4splm6LWOE48e9ZM
TzGnXlET6n4PDxiT0SZXIpCjYvO8a6/4sG5Yg/kdj+Gr930XKc+YNqGzzk4eBqS2d5iKxN/wFfuQ
fiRC1Ti4wV80Ao+NQOrYJbngKTIn7SHsZpcDRgLSzc12Dl/GGKcyM7w20JIpegnAnGTt09fLIFma
4vM8zpYQzitosJskO1ySwllaNzh9yRxMN1K66EE3eHQU222Nzd4yyPpZyNLkbcqgzncooyNu10Qv
cJuzGNOB56He/QMVFNTUNkM4cm9vujxtcJQDqZTH6ZUBXRxciSWmvrLsddUULIkz6aLuLUk6Psu+
2HRoacsVmb3mqQiv9gsiMLwf9yOTWkVxTubXyk0spLe8Vna43ZCqc1azRFM+6IfuV1f9/v3VLu8T
b/Ov/lBjV7tPfTs9XSJUN2g4HeKgIKc7d8mGl0hqWeq9IR18Xo8tFYcumr8eAjP+mEzlWLlGFOOU
oT82z/wLvo0cJpRfoLOMLZmBC6dA7q7dc6xozYy//VG0+WMneo4oCnMThXHT55EjtJ3Lt240IG/q
vQZrijlk7LTG6I/L2ddQxxHIyXw5vNrnmgjSO9CuohQGh2OTdVxgWpPxSOPf4AwjrFJ/kSNwWZTc
JI32cjBKPwQd9cFFYu3W9uyDc5v327RHqAxb2lpuiwGjC2cnd4hNNjodXntiliKs4n4/uavwZmpU
dhc9jrpInUGJxZU5AhA4vx7StRy5+pE9iOUhGd3l1C4lObgA58A3iR66C+R3h+H+Nyd9+1SBoJW7
lextykSlYpKMBCigJgbECvasCftsLblSfQzwLBH13Snhtv4Gwmgd47/pErAk4+jSekl/JO6C/W22
NO7JAOQft7qtRpcMJjYTYyjuhx/O3bQSuwJ5sUSU8peBrO6PElIVc9Vf5rejv3t7retf5MO2TL0S
LT8aq0SR9PyBYVJdqdl9KbGXjFAgcRX3F/pqTMV7CGshfXsJ/xY1z9ARJZk5hcGw1CBWsGQmdUcR
1Y1yBvwi6R6jCH07ghLydLlH4KiPhDDGJpbFbRqSAO8f3Xo1AE88xvUyb2Rd4vyzscG+U2Nq3XFy
ikPrv0JCwLdhcJLm3hWfVK14IKQh1ZiauOuuDKuyli9ERUTt8GsP+AZdxKkRjtZg0YBkBwuSn+2m
Hk/0r1rR8uKuxJZHkhdB6zblXNzTQm+BcOJz0ovw7H0HtlAdffHQfOUnWJXOu9VYdPTPIA4c6Pck
AMdl8jKU9skdvjeMw3jr1GnrXMN59SIOAYAmMcGa4rss0RXHrJn7dTv34aaJKI7Ljx2Oj3IWBQyM
AYLA2Hf3L8YiZVeDyZxP45F/wc58n89O6dPLCLWNDya0l+fy5rlL3z5aFj0TvbBIM696zckCCZPO
gWCeRi1U9V4aWIwWj7y4tOrBL1kZfNC0zUJQUjpxxQvr2slXOgaBNGlpALgi0lDAV02eRY7y8olL
G4Z03pbZHrLaSJOtjRHf00/+IrSTcuac39C/MQGpPFvxjmAZ+bPzwyDznSxbAjWPCDYYP2u/mEvH
5JFXKgMizWVFDLF/cIyWrnDR/WOELhzR364puMVEXELKX1PdpaTMauJtCvSZq8qjQqHJbKBNhmdd
49MDMR/BFvqQkVwI7WDHJQHNTGVBToUngl4AI0RHoHb8nQIcfMC/dlgt0a5pt7coc9mGfuWLBBmT
eb2eRupmy9mOCeSiyTLVmmZFmBGiInpQM3y1QbSPbgo4fQJ0tgViL0h0RCkJ8eKNpwwHMLCjl1Uc
3GNCyyP8mTKHF3CQUmXFVov7F5nzOmB/vAcEH+k2utidJMNsTLHkTL5YDyf2uRR3RSUL2sSi980B
J2ewfZZtT0oVZmzDp2E9GOVimoX34f+VAXYQqs8s+mRbchAnZxz0csLkrtK8Cks0Uttg9NpuZhI0
iin1NMEnswtqGwm44zFMMlT4e33uF6WrihXi8sAjSRB9jp5OUQDx+vPwgHn3umC3zqTkn821rd8R
UBfbgp3IPKXAjtwASccyXJwWqj5n7ZInT1fGAipRX+kugdl8TkjmAxmRri+jmUCnxSC1fiHoY1W5
cuvCkU8qJ/aM5oA2j1dPuFkF/HVNwq2Xpc8egT7SUlse98g/WUnjlLi0gRxWJUHqkkEDpT6lsq/W
s6lY6MsEgFBBdvp0WoAXTGbGP+fh1HoHH5GIECw0XdepquZjO9HCMh+lmAEeABskxhYyIiW2PKpL
I2ofDSiteFK+RjyK2H94+hOaLzzax2dOVMSRh9AGYuZjpowA3ZTkD45DvLWHfDc6d5bgU7w17PhF
tKY0vem8Gbq/todAQijOCi+AugMuc/WBgcqH5UtVBNZHBbvfeC2XsUci3hJRHJUoxpw7oOyiut/A
vJhYXpNMtE01EswnlnZh+MGb1hU1xQF/lxf73NETBvsp8GdJ6sux1YQWGpsJST03ECizDpjOkvPd
rDHTeq8Dy4LE9153VCdlaEflo3nAJk9vsqiNaVyn/Wud2ERljeAIH9/dGoZzczIK2gdLs/V3IxIR
bqyVtmQo/kj/YQPFSgZSNU1zlAvRdU1x42tm8Cw0Y6BPRAqoDWonJuydpLQRrEVmrETPe9LKfYDq
j0nzys98JJT+0gvSyqsyNdmJjj80dJXl5pd8KaPxoTvdVCGikxI/wfSB6JpVROsbcdJUIC5HaXIZ
4VQ85QJGyu19vbPAWdMRPQcicX5L2KgeZwm2n3Dc4uPUS8PAyopbExx/4k+JCwFbR+FxhSVbTjip
tl4Itug9ZsudKDT5meziUCCKBgAgmb4apBncKrtbugaxuow7rddLNepB9QpTPlULbcKC0yJvINEz
8xOHi+O+NniWS6vf2TvK0pLPP6F4LhHtbX9KzGAetCgOEYlvxJVDHQQsa4ge1StHIjoI7YkUNpuH
6aSEP5hUZWqcyQ8ZgHt/Ff8p7DXGrEESzQ5ZdVq3SGMNbBKAHgP+rsxRHwFc+cM4xCov0EO+JvEl
l5KOoKKHuoKjikEVWCo6uyB5C5XjDLcmu6dYB7KftmbCbtqU5oNHSUpvVL6ggn0Zc43wJNQjOlVN
bs3NvomWsQ7CkHpgK5SIK7XSs/4A+z4z1f3h3pcXPF5wh+KQ847jG0S2S+eCw5ZUfq4RupEdkq3w
5A3pCd7hXroDq2GzmVnsyS98p9dyVT/O+JFpeewuRkLdzMQwh8sj2fdQn92yHJ9Aw4xpLw6uAb7H
+L1GADe2ur6I0aLAR73FBYmWlN6rbTx3gc1OKZZzTNjRQ/tz/WDBzGQleBfwe4aoEuosBF1omn31
zArIFET9/cJwXg7gEkVfohHlENgRqQMND0/NXgPdYcMUL8py8K0f+9ZmGHrn8yEzLgl46fElWbXx
oXHq1e8wQLbl2Rx0sb6qdRzXM/KqAxCt0WUSPAHsyf1iespvw8VwYcZ7GplNf5Df0Z01vj/JHxaI
NlwYnjHM/GtHy2j6lS+1nnQhgKhTj9HH0J5SS3nhyoItSRJHbyRRum2lKgC1T3au4TXOjZtaDuw8
ERtaT9hrDkiNnS25cUVspleMfWecozWR0OvOpR+UT+WmDRY+irg6uvdmWxbIbmraejdAi5ysYy6D
WAxe6u9dYJeYWYPVBsjVJXBF5pu7HZhUgKk0EkaQiA2iZVEOQ81eN/nbHGL6asW0cmbyPbXY10SC
00oMAmyJzMvVc45hAOsZ4GecRoLYzAZQnu0IxliH3H6IVu0+hvpgf9jkqMykXLDbqV4D3aOlQaLz
bMzdabjHItFNZZtQ8Wev9vMs1y/jXh7TtNgR1/cTCA47H157cnjQw7x5hsm/pzlgnYSnewOGDKpA
nrR71EUj2g3PzQuOsQAuA6LFEdI9xbyKd553G4LhH+WnEaISASgn5Riz31h1oJrPlqwnfgSiBwoe
UpPrUEC0NZMoCWnw5OgZn6CK82At5Ekiu7mbhr651Mne6woADQQqKlgSf1mXE5qkPB/nQsGOM2c+
JuzAEOABnwm4ufLs8TE7AUOKJbfLvuJpgyJ0Ap1DHkCSnaHR1UEwYVGUGYYTVKK97XGpcrPpG+8e
/MIkGakINr/83aMAESHv5jiv5+g2/rPM8SrScLh+QlQvRtVnyBd4DS2SQHbW9d/6VazxMJz7EoJr
SWQ68So+21vHxRXoAJfcudb38x25hSS3YXtIG1CXlgjrMBXyuYRBDoGk249/K4UZt9MeHzip/9Fq
DkHSNyxRT1hDn2eXnHZhRInqfeWv0yQ5Z9WJPwkRIRq61KrILUZJd2w0oZ4BWZFdwrXqnc5VZgCx
4vCUiyKIMRPHT7Ke3SmTYiEQ5OO7wlVUFpn8UK1vafWdTLICetcRcb2j2aLVcRFxwG6beQFF16w9
UnkYQM4tL51FmggKXQmK60hPkNHO6S8oQqkwhBv0hXQFiLi2WJ/5HlyBQ01+M2SL7D8UMhI5kLAn
mGk6Kutud/1osgOx9AeHAIIo32jSXnveQslMzzsKPlR0ME5480cTkQbeepuLQDlMS5Z+aKzLPXTS
Ta7eQfLkwHhpJzzNUa9OUcWzNZbpGsfgnezznRRaWvkI7xjrzO8CKfLV5IquxgGoBm+PqSWSnRnW
lpfGLb/pJ30XgPJrzhhwExmBAcTfNRnStWOKv2SE/EyNnpflFRY4kN3Z/O6/maf7fmcFtzJ90wVB
v/Qj3ItdHgU5e6bXAf7Eay/VcWK9ylqPHBZZBuXNp4HwNzlHD5r5p3yeDU+cJUB6hNF/mqbDE7+8
TL2phyvfEi/YnXqAzAyDTIi2qoA32vXycuezQaEJ2jQPmzhc/bl/nqJphy/2HxqF+MYZWWF4oez3
GiTlntvaCVvU748YGGBhZe+uSkS0Ca0mKgHCIs9TWTZ+hhIW5AJUUkoIFQX++d+MZ12xMBMk4Tg6
Y3oRkD8ROLpBfwEKkqZOA4dK9wwD0KiN0Aw86yLFrJPpbDYjyoEE2eZ7f541n1qVamb0QgSDPrMl
JwU7N0QAAt5l5Otqar1lO9Xx7KGN4F6OPwclZTHLPct52a1HmjgrbD2FPU3bJmiKJQZnkHiSVAzk
QkLp4J1nmom+jrHhYtzVLDe3uboQ7Uhpt/wy3uvS3/zv1Kozku2P+YfMssgqIYNTILGCjMftoiD+
NBes2bErivudkDQmEy/9OznI7h+3l0ChpdtL7J95lW0WwiwpB590QPfZfr8OP9M3Irv5HmY3ZHvU
TvNSK21R+U1J9bQfqQgTuz8GYFH+aLQo1ciw9+r92jJyyf4rGtM0vcAcpJquTAPNXmRg/eVaJuzT
9HpYtq+C5HDpka2h/nh+l1i6u172a3lDdZVbA97fUMkMBvXBhBi43WvUb0zu9kRUVMD0pn762kyF
Pd2Spyuxk+UU+3dtdg3VJSVJwxhnecyHCXOVm3GJb72Zij9ZM5QZdhKydj4UseR8Wwx82jzcgd6i
6XAybof/x5/ibpvqmgIPua0ep+yj7arnQ+KAa+FojgxWyptatHl2fFS7L44KNc8R64XFJ7W6Ib7N
mmNAgdMAgwtkfKI0ZYn+Kd6226+SmBof9gpA+bngFYlp54p/tSylKhnLpThsvjo1L6RtwaZTX6rh
ROLBeCnJIjmgLF6xX9lmiQ9PXDD0QJUqi10ovaCUGmcqKhPYb8b8i4pJpI3N5wLajEEOKt/BjOiL
fNSXYB64FwCLymH3oTGQyQphHq/Ctk/PH00ny6/gLUW2fL+RzBJwvWKOqvJ/no4drf0CbDZE5Qdu
+MBKfpOiPwby7hTLFU/XEOCXJqdHwZK975cmdJBatg0l8FCTpaFSPAQrkRY8VuKtKWBCpLADX9Ts
D3AA9ATvoREKDJV69+DyvKMLxFqM1mCzLIJgxDoahY6MDOu5u/RCv8tddl3M3l98UrvIsphzx7kG
7nNs7ryEXiGuot6g8T2oW+F/3dGo0TOpPfmsFhT7XZA+ZdY7ElhWrkY4+F07dtmicZNwpeftNPRJ
+jLUjjZ44GvRcTV/MqSpWC94rXr4A7Zk0CPkVu0ts8eQNNujMTBzfLNOrrHLF1smpZSeIinvylK0
8wFSdd8h2+20i+54RRYem+19+sQ4cSe5sgENgujZZdNaDV0ebFOX9G7QC5VIKu0wl2+AgYXpWS2z
WKWDH77K2+fwy56QufZokj4d4ArUDM02AsCo50db55D0a6xVya+pA567jiGuNx1c4MKii0sm6OjF
hVAujMP+HVbRg+rhJzHlCbegjGw1y5fcMQrc8+uq2SSs+u7LcxtrNGkjoVZAC05Q00hYEE4fg+u0
ycwOStVnpPjPVUWYbhrhKAHZZif4pHok3BGWW6ZGTXdV4eFcNsY4emmyUrNPr1COXQiw/wt58K22
TZiiDS5q4kpFlmU9ZSViQVaM02UMxEJEFlk8B8qy2nd+Zp9rOl8n8QBLXWiu1ql5vfPXD8I6Q1EY
oLwN5MLVdjF744S/9gInjS9BgsmZe+i101i9ysTZJ/wcn2/yAQwz0QRgLZh1XH0vW3pQhbibKNQV
3a7ZffVyCQu0mpClS4d2b17oqHU9EF52djbDA/dCW1ux2+d4lmTZMBpEt4ADzymCpIYO6ydb6Suq
G2Xi5FS6xYDzOeFCnziy4YSPbQagqM/PC203uKT+PKFwBxY3ZyYFjkPpgOZTOr0SpnaOw+daZnKv
HFgvXs8hsOxMiBfaMBix8huE0ln0p0AGN9zAg15bbkQvmOPq9NJ9MkXIbUkxWwQ3+gLq9e81xsv+
jnVxkFzAaIRUOLVOvQTXcNy445E08yXjflnppeAy5lqBtoac9SUmScA+DAdWSnJBj1XglKYvUv70
2UKVkgGMBG+0HmcGceCRWTNvXMraL1m+NDQYrDGXMMNz/fVWSQM99DgNJ9cYxQ0rSdVlmlt7j5fK
/nSNiR23ZsOzd5318o+vhs81conk6AJagL9WFC2oiZ3UgERg7IXiXl9Co3ZTwTHMTJeBUQ7HVgf8
RFnPE3dOUmdbJ6W+LFILXKKVhIn9lAhYG2v96McqWydkXchltzIdyH7JU0lUzqCKFoPkVFl+Ky7h
Z0Gh78WF++V25zcEvuaffiaoRJGQH7vTcBO7OMzmzfWNFFlAT1SmBgOuTI5lQXh2CfK3JSM+98xa
zyjv0YweXUhIGkX5AlkrNqQXORx1080rYbj0mFQJorprhY9LTUgebqfBX4LIwigoy0q103fbYVaF
K2YgUA0aVrh0dHmorbxXmGxr7rIMIR0RdQ62jHdq0i93Es3jNzXAXR2535grVLyJXxopRNpNafZu
IfH8uwrGTpyMAiZFo7/4+wZrgOkr//lXIOzm0OQCFkh9WXYPobA5LOf0Xzw9+tjWhncGcK80GYgJ
JtsGMEawXmTLt9HKHDIEJr9ZpfnePjYPRjBHbzq/pzDnsf9Ao5zMawPWpcms0ZYRyJBmHcriUXhv
zLaQ0cJAGIAWKE0iHn9oX9JfEDQ2qBMhWmEQL4KGOU4qNCX5MqhnND3dFN7qRbYlSV5oUk9VA96S
Vi5z3dgPqr67dYvKpPqeUKM7KgwdChUb0K1ZwTw/0yEWym/CQ9HO4Vx+sxafHm5yBeWlmYYDiV1Y
O/Oyk5/al+TCMsZv+INvktPnD6muqlpllrFavzOIScDcZT5gBHlPGvQSYKdjwxM54QslUBYskkxu
eqjJDSoNwXKhdOYApoiZqayu4C6vV7geRXN0ILJqiySKfeF93jXLfJnvgpILIvNYoRMotlMg3iUn
NVEXyStwqEqDaFaUNdezBfY+vpnDOomYPGL7GaIlQ2vaetQRuZyON5NbSrh7AUk9/z3exy0K0rV7
vauKUB49zsPNyaxED+zlNvabMDpa/aBhR6RN+d6XYLo09N26VuHcofESlrnk/x0f7fkdD9TYEfns
Cy2HfW8MStMw9eZM0yR00OekwXy+4s1FzEUh4tWLoofmH34fPNIPUcVEMJBtz30T5OrwxfuYE5CG
k3F0RYO7qSYNGLN+7/h4GGoX4WaMSavxb4i1T4BAunkIpygoDsAtlYxBm5cdbNZKfHSPhNA8s2eQ
Lu+IjUdzySFPHGPAFKjYhIl5QKypW+P8VNatSYbErCO56hNShtiFOZyo6HwPCE5y3h/bejf1IKoU
XjR0hhsQqCDzkrtWSYvKG98j28bucP4DTXLX1cfWYpSFhbASDZVC5wABbropdupBwH9uUz9tZu7M
HjKtp32abhrYHtPJygKq/9R2DnWgKg3CzIuvG8mDU0MsLydKEJSyCjyN2OIOYVt+OUEGi9HC2YeH
ULH+OZEeKXxg6r3RlHO0XrZpY+v21jSoF+HptLG9A7ljTe0a4EN8KX/7AP9xNqbOzaaHqem1IQYB
DO7nZZd8/yUbYnG1sBnjPZceRV069ZN0LSHj+XEfa3WpmGj6z2h/dXALpA9CPzwU0PunCnKMFAcl
jk6Cmt7LfJ3IrfAqnZ+FqIMKQZeY6m5l5wvDKXmkbSNejmaImpOTBzH7irZsXEeUpim2cZBNOMdV
mdtb/5jOKh64rlHQ+H25jOExrOJ+Abt/mP1hbzm0sVZjGpBsXbJvt8QFyXNasWcDVjQNwFWB5K5i
6ZzAVP+5xHrIUyJCcsjCkLocuVKp2Tj/lTAocJfPgrc/p90F5SfHmC9m4fV+dRCsACklX+AFMOqk
w7ochhuU9dZ2nD+HKtY188kA/uQjN/p51lKV83LEs7E/aTH8xtDN6CPBauexcD3U3cppmLjm+Urz
SbZ0Plenwgu97F2BIxkNdGvuYznMP+1+GyDXbL/x6Lp7b85dEUvOtT3sJs4tLViRQZFUl9teHPXX
8KjT+8N0K/kSH081+C6jSt4FyUxigtqGThtOlOe5Z/P7Yg+1/17i7TTf12uqSWP7e2PByMrJCYF8
Ws8Mt9hvOOekGHs7HjILeV9Mm44kpn5/upba0VatBuoomXlXhSJ48cJqhyj9uJ/7THWWc2yB4g1+
pU2H72cORms3h8l3jWDSshWN+1Bs/sOXxi7P6YpCxhSQnBcgmlgS23SWm6nnGxaLf531/q0/mYKV
yVTvEnCf9XReKKGZZ3mdFtv7q4clt7iC/dsraeleXVI2UUdqmZBsn1661dv1Ftjg5whjt7hc3v6n
UI34JjwnWcmk4l0Dxcndb1MyddM43alYfQZXdvBmwGLKZ01IoP1hHNNklteIBFE1Di5cq1SkQsal
BRLEuk5ho4F09BQ2OdTsrcrAvzvq8Cfcpx/PPQbv2RTLKkFcBvH4Wg+K61Purwh+QLX0Wr5sKPO9
Bt+lD70SKPs1sArizN8++xc858pKR7gjNTu/O+Bs9ul/fqBPbdmNHLmBqEBmM7+KeLHeC+prTfGz
UPaE+y4Q1HVY7U2HJcpCMaFbFY8Jq+3U7RHn0seutaW6gsXbk0Ynt9kPSJKU2Ibb+u9IgGg0zPZP
Hj7L3bPnOfnu+1+pszDVlEwmz45KxDIXqS51d+7FGmWxQn+dtLm8tIVliHpBvx43akX4G9H+l/lD
GSlEL6d4kl+u2/ZrfKwJR++xPXJ1U1DxPUV3fUl2tiqkvLncNRTrvLrjs6N3KFi5FzAM55u53w9E
zIhS6kdY9X3nBF/cds3F/YrggURRjRtWRXGVQzv14qiQJYyF+4FhERIdZS+/cRjWX9b05Q0bZtKJ
cnde08hkpV3Y2N7OTFPZ2EekVDs9ygZhatUal1otPJ3bhh9VZN62qQDNDXSHTCjgOpTgCY7qp7cc
TpgszNRWEqlfTXxMk+gLN7VSOfLlMUrdeUuPucSrihN9Ost1cK/SS8bnpg6CPBFffdfksebmdnss
+wteOFwSgELuLysRNzpSLFfDq2FUnnYb3xGxBWDcOJJXtRu0ACZ5PshTkZF71UXrNjlt/D0ViWqc
NsaL9oWAGFr3+decXitaraeUxCwo6WNfWBF8M0mRhh0twHF5ZNEgtc+8CcdgZtHOzslKMjKWMULy
9yYI7lhkwbGV148j+QvMbRIQo4KXnwzRMV03sCHhaxJB5h0IeTO/eC1+yOpGLfxkm0zcQB4Hrst3
IKvnxkLkj76wdTcGhKA3VjM9++GfeNCKm4g01B0mZc0EifSKKahakKBs70iRcOiKM+9bSR4q3UpH
gMO/ACChxOHTpOoaqG/EK/dohwJYcOiK1Toy/hr8rkdGFOMBsyXM/+tZSsEHjZtEAVkXpTcfTqCO
pnyuETuuIWIWzHeJgCZbfdA7L5brzhUOWx3pmk+TwhqR0JM2az+t5U1u43et0QpN3ylwmT49oSff
OYWq5A4Uf0xdCUe2QFfVOhCHKjJNZELmYnA9vP7C5mRyX5akimUK1ttyxpLjYdPBzhrJkMJBUAQ2
ITOX3njZYWUeADWd89DqN/exi/K+q4Lolg++9JiJc9WSLCasCj1bWUYVwkAVvGWF9k7wW+tDgt91
LV4Yjq13AnOnpHinuZ/gIcxEZxLktNVViL4zq1bM+tFH75co7QTRnINl+FspEq/fzLd8yJ/DRWsJ
bHaW8HQ6NcqiDGAXghUrLpbNisZr039yGc6B4QBlnwLMSSns0aRPlxkl7eayR3PoDbsfQ4l28g/v
EkHFUpwV2i1LBzmDhGA1TkNrlNUSNJTSuxH4BmFSCAS3fvH8N7Xtc6VmZJmLda4+RYKH4/a0etKo
++f406HMDpcLF6R2o5UTAh0/HiSU4Snjhg0ysfArhA8BAvZWJ23lNyado8t/HbT3B0anc3FLLkmr
Dvc3QQlId4rdq0f+0AWpwpgKL6UUQwztETM5OnHhfb9PeZIpV3NTpJOhXBftRMPfNooCrEYUr+6c
OCiy60CP0KMxEKg05lFuMlzwwxR2NqT3dCFTmJpCCUfm2do4IADBe4WwrWC4/rXovP08YHVUnoVL
JfY9DN6/rVTleeCHVKzE6acQ6/3JsJvISwZHhJuROQEuDRg7Q9fgSYf/orMrL2T/HnSXX4M04oGY
4kMpmsU/jSz5gAnYym5jSfpCp4eLba2+zw59a24VNrexC8n4WvcxIAU/dadzZHLqMPsiIFipV27f
GtkJNtILjyb3prm+f3z29nKuG5bjhYOvblX2aMXz3Ooq3w1btspfpd2+3Q5X0CRZhhe8Y2Prcwfv
lsJj9BfefzZUxMsQW7NCxUDJuxDsAyAP45KE4CjCkqJkIHkbfAbFtBWjgSg1wPElyOdr+iXrBjlX
nVPPyrjnxA2YZvfxswT+1D6HXjlqBL4U4JkTI1wusUlJpDA8eW3dRQnsRMyPHQHSiJhUvpVfInXz
ndGSSaNgXC+0hr/lSCZ6RovBvV4Lx3oH5BsWGlk/qm5uGTWHmGM3fDlwo2IVGrF9xAeX69p/j8Fv
8PB4vB9EajJ8ke1z8hvQSlzHPcbInGzwulgSpPE5uuF4bVyFG7wiFfp2D74Tx/Krg/NPIz8hGIzk
EmnyYWPBmL/C3OuyLgjn9yS5Wy6ciWRzeFUlI72g8NEGNjHuBgoiBwTS6dknn6Mx0fhrcwUNsyZ1
4kR+W847PTjjl88B3xItR2Ws2CpHJCDkHKjq922SJTpav6FF4VS+OgU77z1vdXi0Udoq9jaDoF6l
CaK9IP5J5xKpfSTMU7iwoxqEpeNAgSvWCBp0dbcKsNDel0+3zGTvi0Hl+Lr9rVxiImG6ei/TcRkN
GkQL/K+SBs0xCrLRLVUHB7hFsP1ZBuCPIAREKE0IvcW6hmcA1sNyhVadWUQmIRkNBTmjxc2uyiNG
BCzIHLf2402u3PKFrzd1max+tuA8h5gsr72huzMQV8v7jW8+S7jsMmG+n8VPySol3Qy+DTWEcOr6
GbYCZpjM+2S4EabeHJ8dJl/mYmTUWOF+aaL+HjASSzvUZ0TVI2HCIKSKc69rqqDLbfsMb/l/ybpo
8c9S3WRIH+yE2tBP9JFPadhhu23F8GkqHcuiN20YIwdZror+IYOvgNKfIQi1VY+aKBszWMvMbXjy
0Ek0nFsRr65UdD5kO/6oN7NcXI4KIWCP/AMeTFyTuJkxf182Sjxyqrw+qKXL5+4F0Qv1+RJeJaVR
ZRDttvrKLYdVgZUymvNqe7aoHWgPFgcZ/bYYs4HbOazFoNEmO0+uM5CX2myqHPh9WLuDNCM6L8YY
WGETIz/ngoQUOrMy90gd+Mye0YjF8Ljer/uCSziewklfvPpRlWxhp1o8sTsV7KxvSgRak5J6LPEk
O76jp3pxYkN7ZLq391c2Ic4YohtFar+fOZYP8Qg7wyoCKS+dLRlmoBMFHqfdwTeZ8sZvcTDPIRbF
/WTueY6dsE30NeEVHzHKnNLpkwdhJsFqrXd0O59Ed1m7fKsXvE6Tc9AJHXufpvbVURYdhOfiv9EC
fgMhMVPPJrVad4DqBzzq62C2+dYx4SJbH5jdcnW32av4kaSL/e4fyZXDRho7EPnCCQ2hg+yQgJkZ
PmMFdhUkP7pH8QJ0gC3KaKHHX6/vW3atUcnHT8w0i2IOG4XE91ptHRZshjRRMNr7G73mK0Hxooup
EfzaxEfQcNOGcyXndOuHoExoM9t+aQspzCq2ZUTOBIvR6puGG2H4rwCTWdHe0qP+ROhRiCl2z3x8
QtYPvuXMMxpjHvRSobee5DrAz/GaObhLd9VF0zbsdLS9v2gpoHbiKwSML07TBhMDFKLR5ydLSxfL
9PBSoFxmNjiL7nwa0f8ygmlA+Lz1mmB3OvX3LsOmAEgn0l6bAZll9jkfJdVix5e+xWdzm70lCzbw
3jnklicPTBdaLJuvQAO+klzWFKtyQr4T08vKGUXnwR0DCVPlwXjWX770RiBvHI2yTC/qQMuBsR9S
kKFz83XLN3aiC8ClmcdSkb80vJWN9p5TK5MwNVICYus1C2NBS/bWE/5GD+azAUSTI2Sx2XrYf+XL
URBbmhQpArOmSPuby6YW/UbR/1WfEc1C06pZmXuc530I07wre+M/vtX9KaZUuQ7Fiuv4IsI/Z+es
rKqRG3uOgIdr6ZZYWOf8w87cOIH5xVf37YVA9BtAR4S5Wdtchs8VebOfBVFvN8xjmZ6PIddSum52
q33PXCJtsyIMCcj9Ca+DUVr7avenPZ+dqrBpHMjk9IA16zPRsC2PF6bG9SEmUJthQXUtqIYD/55l
9eedTCu0/80SUm9+aXogyJd9KRu47JbtPuBl3F+oNul827a0yRmCf/ok4MXh1Bx+oXCOScI8lQ47
Seqxjp6T5i0wDn2O6hBes5sIzjZGvZ0klQKlObWnXAKfkrNSTN4pf/uagKAYzX1xr6n3TYiBxzTV
mDAkD/+pi1EApZBn39ievlDasjFzUMeigvWSu72hLiEryTIRFXDWU8xhjCBSAnUDlTozd5o4dz+c
TFO/vApOPvwX2xm4pcF9GClM67ZyTHcxZe1ZSb12Wh/ZmYF5uXfMtE7dDJ5i+kFrn07QtTcjeZc+
Tt1OQDTZCF/JsTMjbor6fVm2krUiAwrieGuBRWdqFDd8Z86NQZbG9ispcmfOAZuaduMf0OglNo1e
uUrsZ7c5INFfBTXCWvHXuC2hDwwvrCztsc57UVnUmtnOwK7dZ9nQub+qBAEtAxAt16USdpau4n34
YOQ4B0iyaJDwtsrs3YG4Ffsig+tIW7++Q47NnnKjPvuMc1wPOfLE2q5fPbqcQxmbne3FZV0Gzhy1
koqMCHICUaYKQwBNpiwxGFs2zfKtcKLbV24ikPQuo+mf/muVNNpg8mlBCgLzhYzd1RFYuEN7Yvin
0ALvg/Yyua47Zshn5Qc32VmXFUCBSa2ijRUIw1bYtmjCEu/5930+Qhy536pxauVdvGp8edAE/l88
moKh/Prs0dCvBm7SV4STBenH84P1B7czReG+bkAE2oZLlBpJyfJUYDniy8FEN4sjxiFppPE8iqJS
j0G06wXbLXgV84WPVVR47a2J48Vg1ZzDPjPPeD82wH/5Va075z1FtNV2XnKdsEc0NJtwHD+aR0+C
AXHnQ+XCMbM3s/x/qHlOrhEpmYeY9d4Hwcs9di5gvWRp1iGTxP6ODWoQVGf5/3LGd3Ivp7THGpe8
3k1Wge6dt63D2coDwOHjjoE1jJ8SLUR2xXR02HKfRweW/fzwd40Xrb3BEbN5j1MPN4uvIKVldLV7
QR7xRfMoTIXSYfIDSYT7b9BWevcIx/16jdUhSWg+syKtntFmeHK7U8sxjl5ufceccid7tCbUGKRW
XV/LTjcGbHXZWWBQRinyItmIp8HneRdcETcH2FO7zDJ0tiu17M+HmfgH0MUZPCQPvUG9LjFwOV2b
SrcGtlyVCg+01+qaICB72Iua0+rh+uyjWwsgRj2S4tvTzj1h2iBMnf77b1WmhnAO/Dl9T1+VM5Ah
0djZW74NTyb5e/94cUzQPSLzrCXsileq0nBifLVwJ0PZHQJ+EnMqF6ZyRrO+Y25o1lzDZXmz9cCB
jtuUojfWRLXEQpBvWLg0aLujyqk6GH5nRBpWZUwhJhzP712D6jZbF1zYCj4k8KoH0bUjCzRt7h/0
oifNRJ/risEi8qNnF0v67aksyELvjwfFYe0nIy0WKw81tL39PlF2Up/M8K4VtRmIwmniwkuYPt36
u70nN5iDTKuCchQPedjBaKUvANOtOoI21KFohEwoiIu79U5Yy3LwnFEAnCOsXDrSuF1zvfdSWIw2
ptwMbF2ILOpn9xeTjEnMfESG60d2JsGaKe2o45+gs+ujPK0/ywRwHmBX4iAExMJoYQ0Jr6OHnkV0
KRoI9G60NKMRcC8K3xom9vrsIR3hqshxqEet5Wdfb10pfvTjdMIhyD9JdlDbFs7UpLQtxiteNfyV
Su1zEb7JAqN3wsaAHvlxVo1ch7YAKz7ZRpcwrbMLkWbLpggjt3VqviZkd6n5cS4Boy1hQJ6zycuO
YUsdjD7vkOF9j/6hYXCctCZre7IiQvA1NYhoq4Zv9P1QgzwHsQMTLb9evZy+exOM1/JOvNxSiv8o
Gtgh3dqZgBf+k6BLQroL8p2riGYUSJJt8LU9waeU4dQBzzj/xszzbwzrdudbeCnuBcPRluPw7kJe
Jlgrh/sbRvQUrBZN2AbMQfJE4pdw6VbBmqoOVHlwMLPQSFpWrn5O6O+f1FVisA3l4EFXGMICVkXs
Kzc9x4/KRKrhVAaJjelO2LLbp0/VqklQFl5700Q0w8NEIxFpWtxteXgMb4MuVv8bY5fI1LwUAYCR
eINZ3bsv4lY+/mKUQnyJfbF+jaCRhwDXXEaAEq+q26FhYr6KNFFCzsdfBOCepu6BciAWWtPrEtTA
MkB0dVzYCWX8zU+NvdC8XZnUkQPFs68ddlhfAEzyo9Luo+rzSVNLD177bmbXz/NMzuyb9ym6g+fF
okLa8A1pGBHrv6/FnDMlPtHe/7TyB+/tWPBF707IGNBoW0i6sniEk324UgTOd0Eqo44dR133WOIi
63OWdddmoU164C+BeVb9v1qraxJ3HCVmObsdwEox906mNMRoAbSuF1JwjodwpWcdBH9PgDZCxY3D
KMPop205Xx6g4UXoB8GB7yxemV7Ss8gifBHhCoUeESs5jDWU8+ye157GlATfat7e6yDpqMtVOvmJ
SFw8oh3xB7nwjoEI/3aHje7RXiM1mEfuXCdQsdqIeJF9i1Wy4t4pRjLGizveKk+hyvixmkuIJ2Z4
towVt3IC6pY9Mprzb8B1lDwFOIZV7aJzXf0ACu1rDw3ox53/xNw7Oc/RnFXKvz+wXrK5crgagN0i
yuah5d7i5m4MnisKRA2FdWkqSnjclJInncqpgAVStB/ormt6DvteOTOBZgF1+Tq5ZOMa3EY7Kywm
gBM0W2iy9Cdrfp+teDD7CubOPFfUZ3ROTpWUEn+Wg7TLUjaGtmurRydv01n9CKV3J/ga5tbtk1ZQ
Qi1UWK1854+wUDCpuqTUhWq5CO0wTkYBW7eEtc6vMkOsLRkdXm0i6WB5+7qsA1nyQscVKzin7+8D
zOj+gWHNW7CMPy5QAaY8z9XJ1as/GSsSFZt2FUF56hoZhhqq3gYgywQtXDsXckHy3iSm+fhtQ0Oj
T1MZy7VaZ8kneL0d6HzlDDc1wrksfkIzrKZ3fUccq6yUmooRPTbMwM/aTCkL8rWNS0bg/5tEfqsj
73fSJ+PgoJgdZIDe5YYpubyWo3lMbS6aTtTt3k/uj9YrE9HxglO8a2hBFAR1ZuxPxwsdFpgEDy6+
NeTfKisNAOEKBpcJiHpAVimoulgfYNbVk5FfUDdE+Itdl0FBq2kFop1tSpsXaKXhLMUdgkk52tq0
JiyjKauYciJWddh6kWCiFr0w2Dw5j0Ae204RfmtQSp7YxRK3JwVQWqP5fZK1Lxs6RSeVUY59kJVC
ilnKrQ5m13nXjaHBmtqqeCGG1CYACQvwFy7WOQSwgci7VSNSlUM1MCZ2zb2CWgnh/AEqDIbRDiYF
pnEHdJ9B9qdBFfvBZq6Ko3/7BAeES9zLAp42PUs/vRnZ9/KHOGTeIbaZ5Qip2WaRMLNtf3ISKZdL
A53A023xfklnFCPQQ9uSBjYO0xpS3TLRjwfsSqZdzMMftIyXZyDVZtSqJquXWbAPlJg3XpLHKzRk
GYNLhAMkyKU0jSncmJduVMXmBtEH8qemcWghkUwBXoUFXshqBKnRpNKwF0NVRFw7g/P94Cw9Rg5o
kwQitM2gB/NILEth6Xi1ACGtlsAlVqoj7sAKXsFm/yiCZ0vb5uS+Y7auZzA4e20bkvlZ0ZcdGr7t
AM9Lpw6cqlO4u/vfJ68Zra86tklz0NnQbfVO82F/0/rwKrtt2XQz4fR9vGRtESyNNe04QUiGmazh
TB0Jj0T6+zl2QwBeM915KqITERtFXvB+4LEBWKsfCpt8/o0FUVUssPKhpOxqpX7i5f3EvFHQh58P
QLpQxK7327cSg5wutVdGzfYikfFG4wtknOji6guc02hXk9zrrPTISFeMpp57zkZi7PdMfyg1ZOu5
W6Pg4yF1VDa0t2g4RnmTUEzPzIf3mXrOAK7jQ25cYIfFlY29BvBRtmJZ/m+McAsPODaJh53cyJge
poGNWa6PNHVzVSW/Iub1b8J09fGsqpZvjrrHJkk5Y6fR91ksW1tBcBGNsntg5saterwYP+uR11fU
dfm0WzCn2DnQr54lzF9NsP8MnTrJhjC14PKyE1ZbwTpgY8q4ouZYLWujx+fXcXuwruHr/YYkbOUo
OovH4eCqacIvGNQMzBgCi4tX57hbnehflmcFNkLfN67Y5MaKgyuOf+FOKBX+xN3mkQnrp2dPIdtZ
SqvpHiNOyMG79lr9Lzuk3WUgEQ9PWvGq/H05SamSZ3Q++MIgVB4GZR1VHJVXje0bRi6dKVp+BAIa
+dh+0BMr89YrQIuKchPT5xoKuTKxSLpYtD2eR3Zo401ChOs1+C8Aj2vDNmgU+qko1L59RsPDAtZD
CpkINjsx2Mo/ewlFKhsXTMrxnaw/P6PDpg1vLrjrXY73Sk3FLavtHFe+mje/OcPLmn1XTXosNi+X
fprj0Z2gGsdlnaVb6mjs9iLqhKYkqCJ6eSGJd0zIrxdkob3QZfL1cHXIiuL9OQEKWZ6Kg9AbRMjY
UCtFDXqgIrg1/zd1eFCb+Poo7xvXefNI45QqReVrBNRwJ/B67XolEyRyxxGyg9qe5ZYNAF/XJUI9
g4xpnHKewL4vc19bE51uSGztP5jU/y8XOcqjKcNxENJzSDEgst5AxQ5KVFEHVc/Fbhh0mMK1aRDK
k2OI1eEVRQLRa0qP8mNWR4YY0tFXkmbwAITFl7eq2ZN6ggP1PEcN+s/d81l95bJfyBmgYgJ4p3Zt
s9NtAT8d3X3k4sHRPFCDr34q67amc4phC48TUe6reCS1Dcy2bBeeEgIbMID6E9fBf65zpaZtdrso
Hd7tV6Kkvwj0dlqk7tVG9BmzV7ly8NO5UMKauoJlkP6vz7LqS02SNeAmGh9eCPOBZgfMYChV7jEp
Hov9ciJ0ZR7mprC0WstIKSQiGzFR5ykGaGy+4Glf/mLrPWW6uvg4Zoo8LbZQmfDUQ1Kb0bRy3jZ4
HDh4lpKwARxgWpB88a0s7bkGPPJV1BQ702vCQytm4Vf+eWTT3XNpOMd7xKQagrlxcd7RSV2oJ5eu
Le/4TvaISYOHKZVOFALNpIudgyl2vaf2KyHlluqa34HpDHLVv6zhnvHj4fCNUEgk6X70lf8eAwKI
nFdleOFF0+zAbwIVRrIojdcLdksYXRiYsWBGEnFXJXZeOjPbEK21tLpNf8FbmHWoEGa74pY6BsdC
1BsipezoyTfUoI760Nph+Yzn3UevXv2QIjK5y36Ez6GZ4tVGh7awrQARw8DLSdnVB6vf3wlL/Dj0
b7pApEZh3vbQyxG6kKg7q51pOXZ3YBd5/wwzUCBCh4EdquqFOzYH5DRKOxmfOfQINOvsnmmJ8qRd
u/8PklbTZtdWFT89VvHQYJ0hR+9uYas3t6CL7ZRb8Rcu39a1l/tCCySjtTcf5i4vgJ5VUxG8n8JD
CMoFDwHeQy42d7dW7RBt6snBRAVQrYFTo3rQz2bD9q1L6Co8AEF6iUafobpq/HyoPeFmj51EfHR1
D/qE51ALknWvhbHYVLFBHqSo5Nv7HxaLw8oZokhfM0YzPPUnHMuQ/guWb3mvjZTr5A4TOXlrTVb0
5ETHPF2oGC3BiADu7DquXIgWg28NwHL6dqz9x5+subCmKwsWPszcq5FoG1vetaQUlF6Ef+JXFXqR
HY+VXHNYySldSepho9GC6StCC1MhNM6JWahmkgynW7EN8PWVScpg+jg55y1TRY3b1dgGo6BEfd2o
3zlEOxEo6qBiAD7OLveC0fKhOopXlXc5hzi1pTG5ttBsWRfA6LHRAgfRKT2dj1uJnkf5unbIcFP9
9OsoD2ZSggHRfIjbba6T04rFXaWVxn6vZfpPe38JXAg9vrWxchdgw0qVSICqPm+4yAukrjZmlif7
WxdEZnJGZqDCPtWDxHLeAuoNdmo0nYSKDh2d1rTqpdZwcjnt5QrJFY/9h5bncNTmQHCKL+a3hmMA
3ujKWkbXDomLgksEccYA+7sTmocl/jnLruKBqA/2p6sNPFF6WpwYonk/8Mgh+tbx7ZmtbQJolSHZ
6dV5H9GFhLGmv1ty+ibGUNCBSrTEjGf9K3Gf3R2sC3lMsxOtRyN8KIwvQkLQKgaX4MtrFW2wnEg3
oOsQIpNDNli6a+BXddwUImRa0PKstx8zzxcezHqt5JDP1CEL/MeRn5Vv02kFhwNCDhr5dSlj0MIF
X7CXkqjpnhWkMvlXWoBicQG3oeWDe104bE6z1UzvKFC92JXbarSK9rHpVZ0i+fbmjo2RW9lzdKZr
8sipM5nPCfp1Q41xYbrp56NHyXp6iGupmcyBcxl1s1eqF0r6P5hp0eAzjaaGlvAqycDq5aQjYkHV
apEYw03El1QJzhl7GHFJO+It888XlUQzCKlIkO/tnxIdzS49Bs46ip6D0lsiCvuEqE0ROE/hkksq
5U8/A/MI9vK7oTskg14xnTmfAX4ZdDJINK4hWaJLXUi9pDF9e4BXj7cCAPaGlLurRpDMbAratoba
sPhMacWzz3dG7h91hD+0v8dvlm4XBFal4X5Fwj1j1eHdX01RRd3d4/JHwLrg43Rn1P7vOy2BrEu1
Wn+9Gnzepe4oPgWHkC40TUbTyD3bKgouAWlvhrNHdbjkaoADpGzZ3Mxfd6q4xGEoNTzCbBXaeqWL
9WN1GM7D8Q5LN8FCd6MWs72lWuc1fYCPNxxG5VZc3E5h891RUPwRBIreG4OQZS9lYewfwNKigMOo
Fl8mbpBeI4NIuBi+Duyz/FQ7eJKPqa9BQniTMU8zNm6KmLu3tihevyvhHuoG63/j04v4rCUL6UWL
EupoxDHI0MwQm9ISNYjLHtXnUQrPccEJkezDIE4KSeyrjSK7YsK7CSHJO4Vg/D4+eUvhz5H8tZS5
K9S/rwNtGZmBbjLkyX4A8K6MibBzknobjql6TOLERsztaDsgWgI5AUurXgAlcfGcyGHoDpNTvfMh
5isqAKeIoCk6PetlN+vpyXDHHLJyQPCjqGSpuGWBJCOWWR7aCVlCj4GRfN3Auv/99rqdCGb2BZjG
ak18C98CHcYdezobv3OwbfrqBR+XjMfIDigHycXdbbYYiO5nLD1ruYsLIrAzaVp1xCM9ZJAKFoEM
EBa5sajx6xSGKxLJSdLRpnn91bWJ2iAuc8XY20nRdbRTe7Jl2xclkzz8hT9VDWqJ6X5f0nuC4zuu
P/uezU4YSrorNAmcN3jtfXI8VzASzx8uB22/5cLwHliPwiZLp9aCMvgM7W6aIARVN1ybpqKBccj6
qd8ls4uaIP2b08jcT/EirEY0sdWTJZL50AfM+1WOQMjH5s1G3ZwOxJKZoych+wRNP0K7cL4FkN5f
gfieKO4K60nsZN8QRYGzRCgT8U6GLFVVQlueBLZceXOOwifBlX/CUUydB+84vimRbtEnehIzF+Hl
WBRuiNwj3a9gherBJi8dgQu9gwZKywNDdq0xKg2BFXVDTQRE5brqQ/2X1m7lGMT9qwM45THUQr++
A2wFKaDLvNHDV8mYqjDg/xm4ueR4y+oEmcoAZgrl8/Hnja8mTRR0mCQY17FYcguvhuMY3NG8y5jG
tiP1H4PdDqVyjXUIyTaTeWWh7XQGGGW2u5QibenIOW2yYDkEkstxLGjDH1oL2o9L0OgNC2H7fi+I
pcGi8SM5SrGW+rZb3a03Mm+9v2Fy2unoMrZKOngTfOTiaWhbBPBs2QMYbyYYvXjIzNt1Me6/oh15
w1BLZ87WoDkufes+7QtZNmb8U/ga+cBwJvUdCWkMFRL/ioZMsxowMb64DLeqMI8ZDS+RqoY+7lPy
/3mlkl5eEETwQLBQP5Wf4/6YI2EyoVm6Nl86svVRLQ5odqsvh8BYE2gRgWY2AOiuyEnopwG8aAsg
AC8kU0JHEUkpxVE6jrwJ1e5e6ZLUoA8reY9urff7W2j4R9bm/7dvqWyBDhy9X3LlfhKSTSWLsZ6h
MkfYV1EjNULDUbYOPoO5lH+xpRc3fJbZEwg821u44fzXMdjoNwoVsKeGjTFytd9sdtGgpGYmiwZt
Ku8agyAhzXtvdnnaEo7iLHzj9ofIobpQUm/EwFmmZkVGL2MihZtd473M7fR401/kFrcxQ/99RRJ6
tufNX5umoscF8+p36IXfkp6WdWaRziWNK3obWEv3Rl5V5AnBns+Mn300vCcdKVPm4YoFpOTMPxQg
eTMnw6AL9l+t8mHOvli+ZbPN36q9bx3fvKipHDGcsjUCdjNAn5rFoeiAWgj2MXNmUivlfSYIjTz3
IQc/353JoYYlorCKfci/3BmSp315SITSkEQtRr2T5sKDpdSxyOi5syLnyWNcq33qHZ1wlDnaIgNi
gFOro5HSUlhjZqMvnRaAUSCf865SZ4DDLZWx9OOBiXd0r4T9aLgWW3qeCGQ/6iUwyuPJyMrTRy7Y
MpNCDXOVToeAHNCulbiXsc001z7j5bQHLk+qCLPvPnqsJqqD472Lhl3ct+Pvpv5UCSCvsbtgOAeF
mI0afeB+cLalw0cmw9cKAmQyyAWyYmED6Aqv7SO5WUBNvQ3A3E+Lj6RshHS23jjOY/FppM+fYB2W
BOWIDa0pUXVdnP9bzGwkaL8E/8XJ+LebEJfB9+3/aO54jYgU2+GiFczE3Yud5BZ1TBB+g59/SjM0
XJBAk5zXzArym1+aZ7MOA2kyXeNxm27E+/fBtCgpDVai/rPyWXApXHUeYbEUfX64HcAPOMbR1nK4
HD/nnDOGEAiYNRwiAgTNJv7dIbFwFRUQMF8yszj0Z91aLG2gJ6D11Lg70L969W8o8TvNjrUAT4uZ
0nTbf25sPXBChxupOwQbuhRW6wP6NxDMD1/criokcXx4Bfhv9DFSBDQ6kAgHJ371dQ31V+2/pqX5
xACGNXAfy9KQdE/gSlBbLkgwYBUUEfqsGluDGcdfln1LcRsFK9+U6f79uhLnAgttdcr2DHr3zu9r
jXv20xihmmIdUoPqlI/ihu1pzrKJJl2eeYvkv2dDRIpKUMqcxILUlkcc+Xkhe2M2smHobIVlTzCQ
PMU6roMNB9SaTnxNa7sDy5YUcgNspoeJjh/iJejiBrcDlxb4hUkUFz7lS1FWBz0BoomBphGC9c/s
qhtacMRioQQhnEdR2CNWLrhArS4/Q4dD5q+YSmI3zhMZqZMhiFr9wblF+MSxgqsI+0uIC5ArIwNG
tHHX5afUjkvL+49YC8Qe3d/mpR0TAh5ZztuRwYFWowvv4jYrmxE9Z54wh3SxMqGFtJI29/TvE6LW
sPvFzIAwR2vshQjs0mjygX1r6EZqeDJUXDaeG0PKQBMhZL9S44XRd0dSw3OPDA3/cFYAMnYrDLRi
i7rLd2oQgvuYzV3Ti0TM3grEB205wvpCb4zcgH6xLoHK4hOHN3ZOlUk/1naoq8xyM1iLdY7frI30
7Ucv1TGo3CZGIYiozHcWKcoIibAGR9vkknjdpCCCYqgyzCBiyWASS6RrT02yWLCW+4NTxp7IE8Mf
ZCiXPr+fe/ENrtU4pe5NLyQzrc6WFR/9TpiR5X+OgPcWcinVhW24ViX23y9bBqhRmzg4GjspGQrt
CaPKB0xyxk5jmKUrwdXXi5jIO06oNRRRjBQBbFjI9/mMrhaQeZXilqkZ/4EFOPtGrzJjUQ+zF2OT
4/KTDsQbmB1jzrofxKfr7wIWndfDXSgdZFnYbrpGFJQFjC7DzazaPAjfAp85DH7pUZCc5mJX9aV2
j+4akUTZwdWJCvlAGo8RlrtfyuaS1wfBE8g4hp6pUbrL5vG/e//DjAM7ED3jj7MH2hkwiaYcrLBC
4bX1Fwt9qfc7ZQHriHkmmZnDr8mjFiclhwk1NSkKwZNvda1ws/0wJjrTthfOtkAF3drOBP+ITvE3
lXQqa6ygSfnpyQBbiloPlW99kSONKeTe2zVWRLox807EEDE8ykPqXLkjo4VCb7y7VcpMrdFU6eHM
vTg7ITth7lRzwQXlblSt2LDNzymw1MuBGRSzuBwpvsj/wg+bRruKnqpszysECDo9IuHHIBbut8gz
8SZg0d/uKJ2hxQb05K2rR+IBft2hSfTc+6BCf0iR1nHPTDD73J40HfOR3rOQ1YY7KLZgreU1S5ly
TRzP7wuTpMHPhGIg5i7tjWkQTTipbU9F4mo5O7TYwnPQqVL190P5YnVmhNUN3sKvo8xpnG2j6Z27
WG48Dft30642MyiQjU6Krsel0Nt3lcMCofKLxoCr5iTU7dXqRsgDPjbPTjByy5BFEjtMaUaDOkWL
yKvwj9ba51YW+BLqi+I5mDrD0Rm4NGi1td9xHln+sj5HQJL4jR1aXt6PQ/vu93VFcvdfN/w3oRZA
IR73PxF/sOxjZU72yctNlUcRWf1lS7Rcyu2pj7ykhodkh2t980ePh4Cw0cl4JSFhLjV42wVuTUjI
MGKIOchHaeE4ntGyH/243RwiP86AWkgbBDrBTZcK0WjcjW16sazEhHRZjaRXsTxthdzBKgkmzweb
URukhJIfOkvT8b05NUYI3mCAcq8sGGN2TYNlFnsUiVpPSbtps1JTFCB4mJZetU1tkOovu+fRCIHm
k9CEGKU0qr5HD6QSQlRmmiPvh5udcC0tZlEkuaHriAZWaEo7gtTF1Of1v4QnB/XHBCaOVXPs+SSO
rnUxeLmxF5Wpio8/f0zBwSBhCcXszmnFrfrMEXbCYSaK3P5oYMfseBygqLPZtjMlV0TPrYG+Znbn
9idmSq5dPH6d56UjazOJdEKSpb4a0SdueBG51vZfDUzgGz/GmksNCjZW/rtPblvL3W7py2OGQ8js
b58jo/aDfpyZ2ybX+XkGA0cmHIbGjYf5hJKYVz6VBhwivfkKE5EgFa/CJNwVjCknvoMNIILTDezc
nirDTjbqKw68Tx820FVUcwmTi4nVR8td2sK4BeoZzIcPLn4ZjXeAy4Cny8ZR9p+WF0nmK7PCkw64
y3PPBW1DsjmNY+UgkvbMsWaNL8O0rD1a8/9RgI+DnRhjwJmpB+An0sbWlNj1d2ZVUowbHVhIlYYt
WLNMiFBrAeZC9g01WloRujJlAHtLhSOQ+P3DX0Nvifps1P3HmFxz8aKTUaqJecw68jrWMGRT38jV
to45cTqvX2VCBzp2AcZLSxXu/JY4zq62XqrD9Q341G8kPLH5wDXAbcwRqStbuf/kO65ExWfK+j30
LWovBK7YzMufOjp0wxIuzEMrc3ImfgNCV4Ci/h+y5Fcfa5qQ3CsgFp4SxLd2DOGx81UBQuf3AQ9S
BRIXYBtYoY+9nOGt2BDcXJKcVUK44+9+rQ2lgdzX8oRcaYJwA1Ii+DgvrlZD91DEXbqF/pYAMiGF
uIyrzcBJz9cLaGVynvrRf187l95c3zpi7eOUEE/k70UWFDhW5bsl0yRMx7mn3YbcHmMrG+8lFQYN
tNK6qPcY9kOqg6wInp6gggOkg3YWpRsPYzONqIU3vEdio89Q6F4XzG4eHE36uslTJx8AxcTl3V2u
kcUjF3s4Uj4wZZ1RJ8w1bZOBU0Bkml6fIg6XMvuoyaO1ui525Sw3/fsdepctiCw7a6Y8uXzgSQyF
iVeY61fRIPdCMdFbT/upWVthDT/uIhYTKOOr8TRWUQ2V11v9tc/Ssp/Ssh4/suoRq96WCFMll3fB
/vEz3isnv2J7wli9b3vPBI6vft9vhSbX83sS5E/sQLzwHD5uNr8+kG5ZT5hc1y2kDUijhI/Idtc9
frwU8XdTLM7sXi/qSJVID7l3pCVnGE+dseDASbEsptROrrT8v5tf7hkEzARDMsCllzpjbqTye+Lp
3JKJoFcq4Pm2O7MJqQa/OjgHYq2roAnpR0LoW1dk0Thkfq31Qvyy6iD9XCrdbwRWS4PFNjsnmb5p
KXutUfcJjL8E0pMDGSBdWHip1Q4vd4DYKM06ttP9Ifj2E0aaMjVES1ilRhfR+6WR2ijQ277EnLAB
d+bz1PYqV6EBWcksxhFvQic+LEBgG2Zq8i4/XblN674o6MK48B2B/43oCGCBcdJES10DB9mC626L
Rt6umXXms51IeFkvosCtiN9aJvUDFyhDMq8L/SkQt0He6/PHmHeVkPRzLrEw8azygmfK60WwrbTD
peXTundKlFo73Rd2cjURkPZFDnEf4mFnI+qjd4EdZzRRf/98OwMahdBMofu7Ke57VIg/56ssOvYG
BFFTZ5PGNS2ou0l2ViN/wMelgxlSPoLEhHPTI2TUtqBVCuDSn90W/DuKBhnq0TnegLKKJ6c+h/fo
oL0ENXVVeRfdM4s2w5mx04FQpQ/p2W1xK3AvggORf2Pu18mEPUKH9xRikPr8knQFFGvMTmmUVuDc
j5RuGTxPg310nP/n0i8OWaM71m4Eyr9Q+MBLtbOUXnlZlP9u6jDK5DppBHpVjmvj2Jo6kQDnXywD
3fnEU+cYuiEoE4E+bpJwG3qvz2vNdEYlrXvt794L9mtpqCGC6HWcORHOQdTE0UUPEGLbWioBgrJc
GhKvFfrBluxDTTyLTrPpOsh+rwWJnlZK7ydJCxivtmGgOwgz3Bf4B4hVWiALCKilG+K37e3fwjH5
EBKex0sF4f+L5xYgRRqXonVBSo4fSjNG7iKtKSgKs0DyHa0kgf1lchhm6AjNjYo7NriLxMW0m4BH
13HNnGg4wy++Zlr5Hou1D/UJvE4WzXeJgwkM74NombmrMg4mZidRXm4t0Bj9EIybFTO1I6kq7241
sbYUiokAWLy1IMPZOQ6C+8EFBF/z6bWL/9N6kLiELYiJuDNfqdQ07hvPLGELe9h/Z6ESSlWIH/rW
R8ySC63rz/D8aEi2WDxfK4D2xh6eBCIyv8EGmlJxlo9gbFte4UaeBZB9ORHecZBHahzSxKXocQmz
jxZcuSy2AZJwWViJfQC+kp6rw5yhPkgi5g5ZF5LlKIJhCGqWbFGjvs3+2UkkF4UTP/nPWgavTYpI
hNfd2TJLA2QGHuMvgC19HJ5dY8PbhplU9KnucllFKkTRX+rmnkRmOOzISdmJCIVqeNd5965bb8ko
dYeo8BaMJpCp85EShGjsFPMx7CtVBmKO1RXxrE0LfTyCVM+kvt7JQHHjVFjDi693nxc2QMYlM4TW
EFnYYOaEIuichWBK72Fi5FlzbQG1jVEUCeIIFOX+l7WyqrqB+TI2nasI9QZlRbb34kGY1o6Pi782
IkIxdgaTrkxLJb83LB4I0LmQ8xv+ILZb77bgDxD78hooIJ+TbW9OMJjjyXKhWfAdtNdM8Z7Btqol
/jspl1sGSfRM9aQLd9Gg+HdZEz143WK7ttgAEO8ZvAdATX+53HcyFccgX/bkOxH5cqnB0fHs5azd
09Gbc4cPZPThXieKc02Y1KjvpKg5B/1t0VafqonIlFRW058pNztx1Bdylsey2jQqk5aEfOnj7AmM
DZRGbN/VLjdy7+goQH4sYyeRwkuVU7g4ODFayrUPnbGuFV/r/BB2n+TYZoPtwoxEiANuQ2pbUAy3
eTBGHBueG472VW4qUiTfSmZ1hK5keG+jPq6PGDe3Y3UL3A5nLrIxVTixbjrQ6zOVgZch9kG+yO2A
8Z4npDRV1XBNfwOJqOdsfgv6U9lMrjRJttk5honjoXVqfJhQ0YFWPDQ4qtZYp5Uescn79oW0BEqh
gVRhvbe1ga5dP5iSm+ecPFVTIKigOXSJnOgb1WS1EtFpVhr/8s7erwaJP7aHYLlGteNoCYniu4OK
K8eY1sKBr+wZWSuXBpEL7eagXIQcwKDgVfWOPjm5TlPHZTvsMGGU1bxKbnXkmgHDGawyN2SOjzyk
CtVrbQPyFV08Ex2Yv4CmRAsEwaIEhBJJlASUSz03bmVaprdUhD34tOVkuSe3TE/aYU5RELscxv9X
GziPTw9uDCRP1Ds5I8tNZPIqZLMfyEyVgUnYiFitKGHpAgcG02iiUEilYd6iKgPiSsyiBrHpWyL5
J9CbYvISNEj2wbW+O1T0/CEGV3ehGC8nRlwDJ4x2ZBj0OTv1OfWvIsOZg2SVGVb1+JZY1b1stjNr
uSnRRTrWppUtyDAA0eoUCN/Z9ty7/Mj0Yn70RhhsLJZ18WJwEx3frU/2V9jJ62wmWKmb6NPh11Fr
1YjdzPwjKbsGDKVAk8f3DOgpwe4zvN2v+YkcqwLEnNzv3ne0MLqhWV9bFA6gCaLf+FjJXQg8nA/W
rcQB7p9rKZPNTzwMXHvVmLnvMdqO+1Ocz8KnmjrQ1VKEOx2byPkUkbGyprmhqvy5dAFwFVmbI0zw
hqn1gqW+kPkeZoNRCU7uRbql4OalWc06CSmyCgUhMP4epryh2CUkd6U1miYaI51Fy/aKAHZOwfaj
7HAoV7vUvXa6pGhFPl/7gkjqFljjOIHk2YR1HrsLjA2I1nZ84x6Obzy48GoVBRy5ptFu122syRod
CKit6nlX1sWTNzyHMp6ZCGLHUFPIzTbiucNfR29Uzm+MiXb9ddy10wogFZVevsouwKeg5HC9eRze
kFtkfvT6vk+313nxCplsiIuj9SLesj65wJv/3teGf1xRf4gRrEBPyWcGvqRLTzJY0oCQ95oP7J4A
Pmz9SFNtX80GW1JtqnH3EYL6RJdkrz7vQy7p8GknAVTq66gRGRfYAZoXfniJ+QuWk5BkSAoOr0WY
oicOYQTPK2l5JSsail16uEHkklSUAzUvFu/PtAhzZsc15/l/LE4w3eOt3vztvUX6KZLWUXaH1v8Y
Wd2/wvBBkhlya8LpF+3fQMrwAFmfQ4loSmVVT22MDf5uT8wdMs7civZIW+5hRXX0rgEf9DilKGu1
6N59WqNV6kzPVJCM1VjaMWBz4gvQdQe66eFXoOR78D0q2ItoDhrVBHzrUrdO1kB5YRCf6ftjsIbf
W5cl5dFISQdNyz0oP33V39OjqgqxvhfWoWYBuolMEqYgxDXITeEivk2Lr9uvEAHZfOhDPr5THf4K
iH2OtW8EWNkfpuvHzFnl/S/bVH9UKekUnehb+x6EYw4lDhY1zIfZLtFMJBrI0zK6oAdCGIfEQ5uW
hnawo0Q2Q6aK4/gN/xyOrWYza0IVzePBtJ2nnDoizlYoYS5is050v9bd1Da3Xwzs7SofqPCNLtnR
ZHVECWKQy4ZwjJB5S0HDsSQtbjTdBKDkEOxIfqhxAq/TKequkXflJwRU0bzK7TRXJMZcsaoieyTQ
9MLL7ykPzR7CIFhb4NDkcOACJpxmJTTqV283Vn9YdQ0qoJW6lBFNmYvaJmYXYrjbspSMsXLSeX+u
4ryG1NWOQiKG/hwy1vXi73lGe8wlo1nTa4A3f6mx34WKr/rGQGa9XU2R4LbSgcBnY58q0uj753o2
Xw4fXzfu0+r/gyg2iuXlCphof+y94q8w2U0qaeQIui7JMK/HJbD9PrdY5M2//zAQk3Wb38GRjqDo
3Z0gS0zYbxazASRM2M6pdiAe5K0r5l06F88lDlRG91776ZDqY5OYn4h069qhTeVI8kgmCIgNdpWO
6vMcwmLyShP8mp3bn4tDoy7V+j3lIW4ln/Yy1n+hH1rFKGDHE5S9NwswI39ABoNeLMr+DaUYlR8K
Lyyc2Blthf6mgi4tgyq386Nnoe1EFS51TYOuRpZ7oC75GZJ77F/BQXZGuh3fsyaNfhVDQHOskdz3
FOKPUBf5/Oz9xxg5z+ofeoe1/rSm3j0xaOgxMCaxmqYufcP4B7kYIIaVSSxTV7exaPp4pUmfAZqa
vkDdhh1GvaY1MoZMHfPhJKfSVpH22389/9qYUp3z6MMLgem7wm96YPJpw8x1ynksccz1YWXyZMe2
avLlGs50ASwls/3m6CzcQT+JjZxheLzHmRPB6/LC4OOSd9KYtLuHBfCI7JSLTNXwAzTEX2EH5YMJ
cb/V7YXcIgVJLqyg/cPpmWY/V36OukPV2TIS4hiXN4FF1SYU2ML4HQL9PUXRG05oA1annDaW1FFX
N/t8jyYno56c6NSRRh7ublcKhZa+srrQ5Z/Atu9zelVbq3wrQLlzYI1TjLMrJaWJOb/DPosS1oFT
ls4q5gi9nEkv8yk12f+L9P0RQ9h7f9rGrhLv3t5EYWii48J3qehypRwgKFiDgbcADNFfYnk7eQmS
vKt7r7+dWkl1QDlkEn24BikatBmYS2K41rH6WQInY3WoR/P+XXq7bYPQT8aBQGA8xPpeteFOnyXJ
1Jp46Kie5rtKXxRD1Mi4ZrU2rkq4bzRdsZZ5aneDyCwxo/w2sKSdL/hN6Vl5ITJ5mK8VCT166OhS
8LVFvRHtBqOzn+yLl+2gXF40Bd7V0iD6RcOwommChdFn6sW0XCDUhzmUP6VNwh+uRgGE+QX7ObF+
//JS9gBc+1jhhZxsLjW2jCBJmalPhEqqWBYrGvipDbZQsuwPbz8lmSE5MJKVREjVUuc/Meb30fOh
ZGRV5dBjB6EY7k1mQ1OPWA117heBGePDCI+y8NswDAQV8ZhOop//mpoO/i1ToUFjG3PlQy0Z3V8j
BRtBmQk6BX+TH2FU8ra7vAISs4/Hl8JUJoiyYs3W6X4td76jt89rJgHnnE9BmlljfW4gL9l8UH1x
DhD8Xp2OrQ7HyUO4WRP5eHv8ZrjdKg4ml99dmil5es0mvMfzlf/9n2HQXibXgvqfgrE/+ZlNj0aj
7ErwlFv9gQHGSPDKN2smI4jdpcee0N7iKqXD9tAJFeO/F0imcAh7sOnPhNrtEotiJsCXyIf58SmA
0PE3bR0t9dw4hiXyLkcz0xONbNXvgCVo+SHSFKcDlb2I5Jsda0kb2jBHwBOYxM/KufEFWxRrun1g
A75bnNYYBlS9uCkLqwDMetSHxGJnrZUq3Ye3UQ+yTdVvCGvoLqM4yK/wk9x+3QpWHGZiLLdF9Z2c
ZuDzA2UXn5kiGzy9eHPiWt9CVWmoRy+z3f6zAuM1L10q4Q8b11wSz7wJWcu/UgHoGnHIOtxxP5Oz
/9kqArhtoMW5HaaEiK8AIo6Wpv2aPM1wvNZtMkyQPRBoidB0+RhErSDFnmzxAVqy6gbXbkxco1of
3YAlkSuxt/bwpUh52NaKLNYViD/SP68cuzO+3UDQac4a8w1Q2VftA0HQOGlaxP16fZxsTeWiPOvn
o/1Xsa2JeYNsSivKOR9Qz1iF5pyUa4XvSvK1LmP8RiDIND9TA8Kp0S8bz55pmQN+vemimvr/a4h8
YI9WZnbhISoBsyeNgLoiU1IUF5ynHPxnLhVr3kuD2A1QK8TdqDMo+DYy73d6e19tTjengugm5c0k
nAZBh2z+XnT12rMv3d2y89YWb/sXV31sqXdNdvw+9/ySK7Ilbm02kBPAM7eXbinyXCncwQeD0l/Q
k2FYPynTP/MlknFYdSL/gvXhZBtlogugUsz6AxsuBcf23yMwpjjNK9TTLAS4Sr51F+NM9zoCqcOB
Iaga+oqRw4G1S2mtN3KSeqkVICFxpOVnlnHXU2GP5FRqUUj8XSA0ThKFRMmz8BWXnqxd/CawDTkb
I7K4cDRkiusMsSuUzqVBBVYaubi2zuQ35t8lJDP0T7H85dCpxOn5nY7gHeDFoSFP7ycULmD9IXkt
D+Peyvt35GFyrpgPLdtYYd5pLQu4LRTDuw20hXTquwGygZMKVAKMGdO5uD1V2ud/DeZIImU0ceUu
RpFWb4R/7D/VAd4n9lXu7tEys4DDHsTUSExX+/ysq4R3fRdLNsZNOSsm/t3WZAQDNjTunffL1nzs
GqX2x6Fhh1azkWzj2tieaJ4UyrM3HGXl8HvLBerLoz0f64AOWnp2EukpRNP6puzo/e7mOBlG/BKc
ofqW9cKjNrA1XVt3n8Pmv2Ao0GprVxBTealvoAhm79PxZ6xr4HLX6NgcYPIBqFSRzKBhPjx+VkAD
AjS01hIXV0vTcSuoUBanE0F5HVLoHIN8XSVQ59c8VXzH/kl0pZ1Azmh8YUFYFiEiy6Y5TZtFjBzh
iYftOdJXkguofXq3kWFLAyZC23LMXPW4JGI0HMklxIZVRflVxQIt+l+rcZ7ZSe/7pPIOqgSFdDM+
1Dwn9JwTVKKeR5dG5hSmBxMObrCTwCRWQKKDz53UXXRmWU3Bsdd/wgquxvLdPX87GIlCFKO18vbG
sE8Hc6Ohf6TrKdLgJKCf+xGY7NlQEYMcHXjtyjv5pOKu/D38tpKcAX/siRsAXzN5N9iICsG5HeHL
qvnemEhT7CXaZpJ8jLfWy01NlrGT0NUoFBbKGi91q9Qien26MAfT6WTNFJOIKI0LMXJJExtz4rXk
WCEeuNbH51vVey78tdYGJMs9AnGjM3SDYrmSvVfVo7mhKPJkE7MnQRMB9vRkrxqhwzU6WEONu0Yy
rWJ4atX/OXdwOxKU/YzAgmaoMDDQcK4dgyp0kWu9n1++q6ZbD8xNzfWSRX+J/nW9pKx+XyALnkgD
cfaqxkQbL/mmXdHE2eZeT0z7CJm4kyxfSMPqWpbI7JEQmVEAN1L8rvY6JNZ3b1Ha87viR6KVkQYx
DaoLtIM9i88O768AAQTOH6+la5LAD/B1HBK4Ndzh+HNKYRcd82XF/jnoWci38lQZvOzXWJzxoP53
6HUoFt4qXRUAJ9ss1ALVbuK1J4Aj4z+mPJPsKcOOF5mcNIbS1laIdgfapWc7Hl+taX6ClRd1DPpP
RELM+e32UilhhGp91LIDq5cT01NNKWIq07Edv1ic9t+/L+CDSgPLwPo7yY7PFdL22JUZGksHvFGN
VbgzO/oQR0Y7mtEwyGoPszRYbbfyBKQ8I35STXdIAoKqH3Vuql1bBdufebrC2Rkp/mMwDW70frlI
F3yDUZqcpBWMZ6eBFfl3rToFb9EFMmWQdCRz7FwB5jVX6zPs+u/2qrh7MK6Qq9CiJshAYBLVrtNI
i+CntuLoxlpzpuA3LrKSpkXz6WPaf/qXgHIFe5rPKbY6GYnwGvQFpU9G7SQzaFHxvNeHAVj+xFjY
SFEp9VGZySjr/MypbGkJqdpeMtIIOUoDdkTfD8XGqgpEP508GkrPvn62qV9exh14xRCJ+Kbj53xH
FkFO/aMwZ5lVr9Mf0JbKhd84yoMzDekP4GcWxJthotXReA8qhvIKrydzkrRRCKa/nHz6KC5THwCz
GciTRTLItFSmhCgRMFk7TVmtMynl2u71MFAH+U6g9seIEJ3susWY/K655e4kKdpMCUaMZDN5zLoK
lZMZM7rM6hofS4H9aQKXL6Cto1OrCFXobtNTqXVshMzXCGdm+BpkGQIFWwFL++27DXJAP4dlkrKO
7knP5YkLU/ZCdQIbKWJtFZo0GDZ3kN0d1ZDnMxkzcz97MLWaP1C++aJ9QNk/WiDKPgbm9m45JZA6
NAV30VbYiLvi+MyW7V9gfSq/qE/C3fgjBayRRqrRw42FICmnoeM9GxrvGuHqJukXo6X3t/xhi+kP
HBSQgOAAArmSS6GUeswqjFsvM2Il+Q+0VzdBbttFwwBfM1kcywb0cCHHEvjCgj36FIdnMiCMYadp
Gbe0EX5E9s2MxZv/5tBecA9xn/WLEOpexNdC41ka41GEXaUvKW4xESDc2TIwDgSH6wBoyNa63UeC
oYZeh2W+MiacF90c5GgkOVM42wA3zXJ83A9eLRhEssAx4H/PYtqhrJe9iYMNZgrEU8EuuwQXFtlk
mdOmYlaqG5IXQpjfHdyrbE6so0J8dQ6THEQ0LeGyxmtjCAzCYQUehHmqheOPtZgMitBeRPghvhrg
Lzf61M9/AsuPapbgRK/iXJ95IWQAgSGvkxy+4UmvgE1dcWbU8jLnKLH/z60zHZbAge2WS7dgJBFy
noAh7UkGSe1AHg9yEzuajVy2txPss/PC5RF+TmB+9XlL3Hjk/7Sc4ScKX7M0KpmCtWo7nvJSyjeG
UCRCDBNNBumTp1/cUtTMHvwc1ktiopUp8zaaIskO1SdicMySJi47MxTJyv9zJXjLnPZ3QtA9SUM/
zx5Ib/8WihcI7k1M4aR/0iX1Jzt7+14gxkTcbMMNuBiUD24R7U1Xfp4qizFOxBsJJcZ3/EFxOAM9
ZqN3Zy5naJHNBK2KmO891+IO/IH/5Ct37+K1s2LEdwIeJe2kVWBZpWVVVs7Hh0oc6R+Nlblu+AqR
j+9ayZ4Au3Ux9VNNsKWdCOdzU71gE8WioERCnarFnRbBQTHBU9XoKlS21h4rFtuA61vtIkCeB6a9
Gpr+0Z4KgJfQXcBP4nDDUlO4uydELMPpJtP6luQRHpTWMpNAt3CsEly6fqNr9f9O6dW2wvvBwgBc
5DLTBPCQuQFZf4MUzxqb/wC98M7lhOuBEDTTkRrohMwMqh+FFEE5Uo7IIajUmKgyWiIvllfo4xGX
Ry69POOZISnUM9PmEKkG/GtnA3Z0a+6V+iAK7w7PpCHVa9FU+6BbzLKoZdUYnyBRzPzD7Gj7a8YB
3gBLIVFifXyrVy4ErZV+IYZHLuXmo7D0qAZgTDsIawQCsdYujqIz9CVsLZqfGKOadhF9LH1EJkyK
Aahag5OXiP3U+WrT4n2EzXqbhL4iIscCrLSQJzLAtA+1zuddn8q7jf+PY6jHqcSg3PXBclU6Bcf2
vLUqkIJ8ZOEWlXZxAWVcayAiFbbUMUBT4GNSoQdi8cYlWdK14R1e20p/c8Dq/SNgsBOPqTZa3Bq7
uWGliXxL2yqm8+yw462Jbaxcv8ACmVa1NZESNl70vvVjze8Y5NlK1aXO3ToWL7iWj85swF+25Bfy
5Jm8oifrZEV/dIRbZKEQe3pFADMV2vjGllqxX9i1yi0ecV7W+IAlxZ/vM+2wbh+aMlkZ38sFTRDM
+b3Sey4PGq1VCf9lvWrRViexs8uQJ8UMjOfJ4Oi8HfW/FckDN2zW5oZ7l2dfRmFunCy6NLKDnucQ
kjTFoOXfT+En6Ha/XQFLOqXspZkV+W4dNobtD6d+4+3MfB54rEMqZW1z8z2F/CZ2ZOQw1Kr/dfOy
aGvr7FyRxnbHpm4VjzQrg+wlKrdDQtpDr80ugZ0wCGBVfIVtMRnJfbUiiH8BuXvEG4BgwiDEePm4
WtN16Gg0V7X4M1SPM9eL9y61+x36ltReyhzxNPkVrYXKDDWXQ2R4iySX+WU8qhsAGRTf9ATCizML
LJXYm6ENW7N5XA6Nle06qw+NKgqqEzgIe0c+SgGSdUITaSHKsuok1w4A4GFyU2i4zEXVGVNwtEzx
VXSlApt6kqVuUlXYB7ybMXExTAYFFuWjcmv3HtGTdZ3BAB9IBkbe/ocGu6O1igmLCuyDdfxfdBVL
6J/wOJSOvPpJqSoKsP/FMPhg41YHHuiSjD0VjCITviJkiHuKopHYL/MZK2K36TYkVTsEKvfsvF7j
tB6+xnjfmL8TSRwwTdgt9ww5dzP35zuCB6RevLtszpiL5G90rnd8l9mUF7WCPWMFHHIS/KoF7Zi7
uLC1k2kweIGdpT6Q+cz8sSd7CTFM29meiUp37r/mHH5UcooeaoDWVaUjxoOZaEybYu5qy4ZwyNVR
5WMEQJorfunvDFyY3bTJWGv/U2Gjn15+3h2N/YyWuQ84N7o5+vKh9QlHpTBIMec/GpDPklNTvcz1
6M4KyPylwA4D3/RUldAfIvnPjuP0oNZD67HO4fpOSG9QE0YC00QQbHw0iKzJzz77I+vU1VLv3hvQ
l+nh5LTxTuQZd74hvIDVrvGWmCn2xHkCitk570+CKmigoGhtrzY2Lw/fcWmKo2wwAyl0Ky2ecaLR
Fim4B1rTc7C2UgmcR1mCTXREG6fB5U7OVGxbSAWZy0Qra9bx5orYUKDRX5S4e+oVtnoGEU/4VKl3
OTK3ZOGHd4+o6HM3eL0vvQBzun9+FeoXeyedz/P5QSvVj4aLNQYfmegqc0V9lyvYfFf9VnA8lQYS
88vPp5/C03Az0kOSQ3l5xG6zD8AekDp09XI885x7NOiRYDUdVaUf200u54wWLdNr3LtDYqVzgBxH
wflp1iqzcp+JsckZEio39F6seVm8QKgPxwRoD73BZxlSrw/pbkoPUZIAAWO/upEKMhvS3UvMcV/S
ymQqiJfM2kunoEkAbxjy3LBilhHnun/yukr4pRB5uX8BHwMg2cWocxTJ9HwsEWIl6/MpAqQWDKRY
14esjvKqHJ9q/UEJHql9Eo884sixpSvxfQXn2tXb1IKGe1nmljl1QQrY8W81BDtL2M90IFUmvXv3
G/I/q0hCK/qEb1h5FrRlSahBbz9lDaUbaUCiwXegyUVEcjLPGFs14z1Y/VWjBkdf9WtWFfAPg+w9
6cgv0CWoX7HsX2ZB6JF5e/7YDXbFD4VQnzuNapEBjxRzE1mm+QTiKJ4S5z9UCtQXEzQwmFjnxmdu
0dobAGT2Rqfccs0MXOVdY8Ty5oBcYkquOfK1YuGaDb9mtwmbFNt6puusTbXvtKp0APWOG13pWP6B
Sqq/SlVd8rjgN3HGv4KzG7Km+cyo6+LmfvM9V04KwlKmZIBD2xtYFncDeza8EbfcJY9YRAZInpQA
4sFBCPmByo0gWNvI9ygORk2E40d2cnMqqWWhRTU/okGIZwr7D7UakxFxouPLKcDNA1MkkgYlu96I
LW7KV5aaK7HwPHFqKtdmrh0AFobaNM9Ba8zBIUOpnuCnWbO0mm/4CaRyNkPctpY6c5eu1a1JbppF
ca0w1shxxABactIChuXpA6InCoS2dKcymN+hwV0Ytx89DjOtxgsulrKENZ5yAb9ml/Mgyk4Q2uJ4
lrX5Z36qSFoP1fH4vbIatNIk+1EoIVspXS8dtKW+R/GUN+Cc0fIcgWbOWdaIXVb9cjVI11T4XUS0
rXjc8piT4cKVHVtYHYkyGZhSR5Dq1pQ91TbGFAyTA8doILm+yGe419ZZgWoY13RRWoTAvwWy2OmU
GMmPpxMpjKSRGkZRTE2NaEm0LQaMpSRH2rCwYfzqKR8S+kPPG093LgrZ73SGU7l3Zmvz81XFVkRL
ZaawO9W+n7e8GkoPmZy6E8Gq+BNOQWWBWxRd4bIGPIUvAe9KRK3jBmpMieLxy0jvVA09hYuI9aed
RNY448x2z1qhewxqABMKKQx2UfhfjNOMmMe2iHty6TIVhQ2QY/JcHChEzLfa3gVQfSTNfvnHX4DE
RR3T91pnbbdde/xU8OT6hWdoGSVZsg18PND5BS8fyCD2FLP8Ly8N9dGzuB0pnsurBsgHgBoDqTcZ
zrlgEKgnccb2b49xg+8W4oiXCkfyNUqOFVvcTTa3fO33ECQxbgXaXGOybXzYa1uxXCiQ0UNCWQ3t
fDV7zdrMX3Xo4l/Xqe9ZZxv85FyXACnF6qR7+gQfkfhztCnt9mff2dWxU0UozlSwQE5j+GlX5/kq
WmYVOGCNUTvzCRZRQvCIhoMrhRLAJBfW8wSycENZMvMReJ3ymjLRdiljk/hJvd1QScdeBAxKS9zp
5yO/D1fHgpCvMhloFyIRc071ZtFt2qJ14tNgslwaTOSdtXrke6EdbvKHv0rSvgGKF0DxSqDsXdfE
2fKRO8/KfY+nrLuiG+EWX0OkDoUDYA4jhvCCXM3b/fWXiBQGNy23Dz7BCTya1fNLMY7YgVLEtHwN
QV3XzDpGAPdCl5VS4PmMHsvp3DtO6fdEN8INiNyHhdgWEDBRhcRAPHNRCfhoIoo2fzIyGsWctiDS
IIcDkKeqQZmvF1iDRh0RPnvYYpG6KlCKNIVHE0gEjzmedk/8GViMc6otzUXxOA7fd1AsrihelYl7
VjaHs/sVogIr20L9xP3t41t5ueA0ImTa/NR8W0c+kwCQsIsdoZpuZ/izwTur6Ox3lhwEzw/isgNG
ZWNO2sSuvyahXhLz1Vt9Er0Iyc/vFvx6X1+ZbGI0bydNlmWpSmJ5rp2ATJiAzhwBDI4BVHIE0bse
Sw7lslQrmMdZpUVGk3qnpBnzO69xDPX6/xTpWz0OeBjSBOSCeEFVfwnUyt6WkMBVYjOIhNX3hYqj
XyoCoPPuS9IF6MzBzSJnGmLPbRBDwFtEUd8kaAiTL52C9hRRvgnTcoAcEd4j/D+kQhtWdTLkmf59
SDFV1oxs5GK6HhEhptMvTqpbF5HWuPbAcW/Cgcyz6pF8vuOWdjCcAHz0DcM52bPYV5j6FwHh+MhA
qju6AGlI/MiNX6U/2ADwZzdwsfsHiQHvc0+6Pe1oaEvBrk7imfP++Lc/sVtijsPVAsK7qYpv9juK
5zbDJLj0JA3k84qqedq/LxdEgYMDS36+GOpMeQ3FNzJp6W0bYCnKZjSsbxGCqVtoeb9zVSwXHIYj
Rsv7eXkzA+akFjeCxiPPQ4q9VbO1pkvUd33VTxnqQv0CYhApq0rQ3hBiuZJKcMbVJpCbPMRFAoic
3hJ2MIRPTAP02tv0ddtUwxDpLj2yZsLicNkhT90pNLG03vuUT3mhL7/jS8yWvm79IzQGP3ICeu01
HgFxaujlYIEGZEUMNdP9S7D4+EIanBb/B4cZ77XVqObkYS+T64+AbnVkKSnhvdnqFl4dhMpTnY+9
et7bL0XAvcJnvoe7q44gPeBgzclGt92C/uCbKEkVtS6Yvpbz/eXHDay9r9MNSPV20yPVRbRdRY+j
NO+0zOrlgeoIgsGqOj1OZCtewlBKTlg46Uhgmgtk9TS20bR7IaV7cEO95/r5X5vra2mfZds7yIbc
Q6jqu1xgCcCOMfHkZWSyba/HlFRzlNBmnHVfyTkwJhiI/8UsL+ynKGazbxO1OrPFjLz3Sm32lkjs
fkUsGbf8R77LPxWf8TRpoG/VOTdNMLw5vJiaCy+6PKn3B0VYDCiUo8qm5lzlBjNYQ9fZSdn/ucHn
GWuLz4Rw+BMkey4oMCTXL0yoViNSEyQ3HMN5NW+jbKtEfKrJZ+p2QNwOZ5OHa9fNJvVXzdKUH7Y3
FGYEsSCsBktraqZ79QtDC0fKpcIksdWDLJoF9mE0Bf9EzegaQJFvFyOrYTpDwuQEHMpMriC7+BE9
MI8XLiU8FZQXIf+C66Qw87tcgHeM4FU/E9j+Br4ev0MNvBUctQDEsZhM5M2YoycNENHNEK50giEr
B27jxfvIoDEGRg5pE4V/wxZt4N0YcOueb6tQUYaQKuV1+W6sj0LNPLaGq14AfKQyqAP/WLvztduz
uV0wKV80eScsiFV8NIXtMNm7zNHN+XzIGrV8QpxWPjFzK6d6AHpCtA5SuCFatjkERdoRwzAVxjSh
Vxoi8+81Byp6wf1MHGh1vMzzndrceX8MTdeQs6tPARqlU/LH78jG54RLqr41UdWL+hV7K78J3Tep
FFACK1pDk57fy1OMeWocneW8mlKo7+fgwDIU/0G1QUOSCRJm2yo3Wy1DPN/6NXcBN/dyvnt/X9iA
yX0K/rl0y4dmSaWgyQ1Vd35IeV5ahsUVHzeb4rUJ9gFLSqvMPsSpIbR4QboYRMBSYMsq3m1k2FrS
6QNwO3ZP8hS1RE7sely4/YUM8MBUcCuCubJN8mSBIK1f390akPYKMaWs1CrNu8DYs7jddLgADk/M
w7MyO0DItzHuD8lGCWOfyPI26fn/1oRex4MBPoypWAVSs2EXeHmzrJvOB0f1yo0hFKTENuzafwxQ
p3Nk/ZYT1UPWJ6zBrmuJrTYFFDaI7l7+QDfc8Qw55UmDokPeCep0MmwRKvDfP7pteg0D/WyQDOu9
6vOiOd0PBDNsQN016nAtyb+US2PE0LjxT/50TOrvBCa6V97kPBQZAWwJxV96T8BOC6Wv1zxrviRY
rsbgJjFhHfqpB7z2Z+ln+YdF2fobuANc5ovdRp9CA6bjcHROOp+DRejgLyeAq47SdbEWSeIDXRV9
uDDnMtH4mL18K6njXCWqBzj3oKjvxArZA4BaSGafAPqEBkT31VesEAxXJaxKTyhXz5X3syJtXnU/
FDDid3xjk/nOFOS+/+PIRnSn4K68wXTPeMZlE9RqN8x9iNyQARHVIylDoolhcNbGCSlICuFCJFwT
BsrRR9DsVDgYHgDdkeeonRaOXAWUwfRj7z4vZqOCKMkEa6nhqW+vwYHyZkMwYD3O+kfurYvHlzUv
t5vH2rh4+wMA34w3cLVBacJIYeuhbPF7TW9tVAQPIRQH8sELVId9TNOyCJBZ7Q3HT/l7R8gnMGJR
Z/g21zOvfTe/pfVwZfIi/tDnmqx2GqFFYH5hbabXnuuVkYnltrNmbmdwI0K57EvIJNJCpQcDp7nJ
naGidmf/ICS6VWfB+uCZoXllBfnia9mPQIuzULpHnaM/23ROgF9QG2DTjupyUVq8tGLrxL0/8i/6
/r0u0+eJuKGcJ8v1/gpOWl0B/+99FtVV/D3Fwlle6Xnj70PwlM7GP48zyld+9lAu+b8Uz6UkPN2c
L66PbfQUNcr49JMobqWnwcbGuYxH5DTgC/+PPIvNZ9bFF4UpIQXTTnwnrfvpIwVhN3RaArl9h3gF
lrfPPDsx2AZ4PidFJ6qmWdhhroDMTmcRFb/e2U2/tTARGiVuU3IYCcT76vFVT1dcikyw1WZJAqrb
zBRWZirgHDLPwbAOBJ6g+F39huJ5y69+2n5mBEd0kgVKYVrYmJjTLjfcm/IvOx8R3e2eL/X2GhRn
W3PJb9PkiJLRB2Cm3ltNj9b12PmUJbHfgs2gYW4/DmK9tJQjsLMmsCAv9dismDgn2KR0eYOmTXx6
InKYiBdjfjwiq2s3H/iq5tIIC7xhA8y3KYOy/llE4QvgcJpY4FP/8akPsnV5MsyBmaRPHJrzaKk9
B62+YEvt0coHzlZCwspRoRyCcvHBVw7nk8dxanczWyorHETLZB+ZWyLgWkjiPV0pRq5K/fiuEqdQ
CGOLZ2CTh+oVH2C4+VyZc5phHF+QTmVaY4LI1LkCogmEB89JqK9yRjbMrM/wzoO/rKlETAzp4yyw
V8An03VhXD1eenu/x/r20Hf2hi4zVKS27EoyN7ZjoGR5jK6NNAhC5t0WV+yS2GqCfC0ldj02xtQP
Q5zDsAcBxmkLohEr/AjVhB8uL2V67WaT+ltsJdUiYl1OyftkX5m4Oy8sp7ZpiA96OAdhqW4dzOGm
0J/fGLW2UGCkQqrBRAk3qymv/aWeD4HDlTu1O/GeTfYB1lTzH58sNxWz9LzvNcwgoIlRCqqHBEXA
circDqogiKaTAdcajmC83qmSi/aEqmnbyj1bCh+p+LbG88tQdA76/kzmFu8exsxPexnRXBIEsqpa
TBsuRxqFBbYKjtk99Yz2pkPFenI2XhSuQPlJdGPGUGn8Yu8lBsm1TDAyCJTzkESUx/+zlBHz2XrO
QioUQh4ArfQiok1TW2LmhLUqHQ+8xl/Pusqp7WDOti5c0U3rcgZa7LnyLvsthsMlagUvo10VSkf5
HtKBJq+bsMO2tYE4Lql63xosfv+mv5OaZZdgIMADttHwxP2Y2ti28NAXSNkpb2UhRjg+n1I4wg18
oB4wcvooo2H0T7Xbx/qiaRfkEmXJgyGkZgrDh3wldSH7ygETk/Ns4m5xnzlqu/J7kskUSvwBy9RU
Ntu3yiSM+RyMx5Sr1AkmrKHtwlWtSJntPqN9D/k3cNM7RRSbPuhWdMYfnYIDw7jalB3W8FuhyRez
zgBXvh5H0b4wnT0vMQSo6QP7Her5p6+boGlRILxBllZojLyzpRMxfdZ2U9AqzRoSlfVIl7092RFN
ek0scFDmIpsU7DripGpcDbYxdT3btSTkC0wkphsAbzCcwrU1HwGNQWX5LfstjsSnwg/hLw50F1h3
7bR14EFzf2Eci1lw3xHNv487vdXWYgHx/wKyWY1cjf/RrNUc1cVJ2DtoRl8+q4jpWNkPjb5TlAms
PByCg8EPwqCTmoDKF+24W6wYKwAmsTqs2L5/UUWYVp9VgzwwS2OhXLL825gSCTurNrGHX0+oXEOl
QMrMR0MWR8DcWfOlLYFCLMGcEgC6O4eGl/hozQc15laTv3j1PDxPJzK1thOvn+64/C0n7k+ZqTQL
eiII/OodHYRXiNOJDUtXhJMPNnD9rHQmRC6j7fnM741FkwOVHN7HkcDgaAu8TLx5R4uYggoHKYIt
jAzRpJgYXfy1y7F2NQPB5mEjgMe2BRO52T9MlJIHKv8NpOurfkGZtwGfuVDAY6c63cw5Ialz1oiQ
6xBtFEOd7+A4EclD9BGYHsLXcwjXG36dSSNOD//LkgnAjjXPvjHSCbydN5yNTTr+RfeTU+W03ljD
xPLM5VYqkHhbhLVjPjfX4UiNEOgRuz9k7lxvg6esJNpsXRE+7n3RnhRDorrw1tLWboljhqr6G2Wr
ppnSh5ZsVcp2jHGvmo8radaYAvEalugcG3rZuj76Zy0lA+Q+bct93WycYmyvDPZ7aIF7zSDoKgx2
eoZctvzRabZyHdDPcZ16OdYocCTa7/H+1/heXDUUaQHlvhjKmWdY+lJ/MlRKFMoTvaRylZ1R93ia
jNns4FqdIQuwhvabLRpRHUgA+b8AeJrDD+S1zFcK8FQR/7QMC5w7G2gF0cx2GByS2Zbdk0efWviR
MYITkheuQd4cpB0PsFgQe8H1DK8NV7lISz69rIrhQesGUvtj6QAQTzw+qK5k0GJlTrGzZ94amz5T
VnnpA59vdwyse2FRIQPPSqDeWRxW7Q4221byAS62g+bppOEihTXVtm0Gj3+sCXogOB7gUkKrsci+
8wreSs1x0bPmrUtItXnPIP5KG2/NSXCaZQRpUsL8IKYaorYEaHM9RuJHoeCZ5LyTdRiQxmQtSVvG
DcbHwccbbuJpzfFsyEnyIlXY4UvAdL0kW12LTC8z1JrC+Ry5GdKEakGBGdUffPYq490whPrYrA5O
KNa32VgRYA2uUrsykxBXScBF+R4hPYjS2+Ar70FmuzZJcHaeYuvxw8XldEtfsnO9RQYaBIX2R1lK
t1Eug7fX4LVbIzGsNtfMJzLV3H8JTJ8kMkiJ8Ssqy+IuDrQbbLfmq3aDGuo66JXBi4WfakTlukxm
OR6Xkkitvgyw/h5a28gTBMn2ft2rRrzMqska/5vf9tqu+14XFO/rtYGSB5SDIuFaoLp3M+MpLvbZ
vuZ9ov+n670Gsf4znUDnRi6Zn4FaUaIF+zlUcIKPYenSzzJUOjc+AP+2ndwmLglvlVA2OEVec5ni
Jo4umewH+ouFQk+P2r/2VoNpZw7abapPa4Z0wi8cSYOW/2xkoX2yxtE2BK6gzq7R8qwU750TPzf3
/O8RJelLx1I4w6785BF94+y7SjRadlW75R69ljhfIbdF5+xsNFKJ7b+pRivzXGg4oRQTLUIzRhow
bIlQZ0strvUIzy0Wm+gsVW499MWj6btS0swCWBCgbbHIVFCkIgxxKmDd7ewJVgBEJ3xYgDuS3/i5
xlGT4I8E8dqc5c/qscXSC4UKAr4h0zdaaQ/VysqdVrSZ9ShB1mtywnGwcJM+9c22iIhr+3yWbB5i
m+pVHVsDybZvrDsfdVFDWLldCMfTFAeDNmtMGqCN0YTDT0NUeSXcZo1CRnzSI3Sy/V58eDg4ysJl
Q+VrWNHQNBTmisXdMWXevCwzcht86Dk10TEsgffiZQZGGoU45V16RA7xHgQTNYhz1PMUthcKIeMm
Manqhs35O/ccFNRq6tfYulXy1PJZ+/ByKPXorFvX4FyA0Czy8kgMOQJNQXXebDBX66+G5+s3CN9d
trNNhgs3DiaeTvX4moGp7FbEaSQzmMZEl6x3FWvYBwXJ3Npew3N1qOW7JezRd9TTeiSnB+W5ipDT
EM70agYUPDKemKAJYsyO8b7uNiYtIQMThxFG8qJ6yUlpudM2k8cEBr4fovalj5tyeiKgIFwUvtpv
v1JQxhUK6UV8WwgkC5GAT/IobG42hwcAX/LWjGYETZ5tVzKb7+GchXhNxZEz2uIqElHyFswv5DBY
OWAGL/eyRKhEN8xuYxsAD84yl1DdMsieV5+xnck2AToDqCTO8cE1HmYoWKo58RomMlsLgzeMJGKx
Cd8+TpVPB7FoFF86xsu4OA/A9CARbzLucyOcz0ReHq/oLbNoatYJA3LfIS0/FqeasxJn94ZFCxBy
LwaEK79r1MdQlBp3BUZf+nxfLvPS5qPhwM/bz2YWohk8kNZLBldDxcYueBt93rgHkojKe44vZtoV
xyE9eZjfkkfFlnFsai+FxfiaKA6l+Cnu60jo+0Pfxyq8bLk39PIqfh/SnQXgvqzacuC8Vw/hQ3lU
I/grgeMalxdHBZb4KYNhEPLcqQy33UDC3GP2fujy8zzCUEE4IhfLBhaRVIO82QF5tjabaUcXyLEE
9jpcFBci5TtwEJ26XLEzG65WomDkipCeqNTwahV6sU/rojQbpHXZxfSp1rJS0WLLGeqYdXnBoVWi
5QVgMVQLgZJfzawrfPO4evguORBtm+PAQayWNNH12gC/AuPlrdcHszCtgX6bTCSig5QdjH9GUx9O
WJlDpa4LeXx+lNCcwryL3iahNVm42t6xY54ytTsy1UUBvoU/kxBYE5l5yozQ+476nmNmpWqMzMkO
MxzmmlASBLQyZmo4O2gQ8g7Z8GrYetKriusILS9YhFNdseS8W2z8kRYgKCEVJAvc2OJ1QlRuEt6J
0IRDL9a3Aq5NUbYxQQ4LT4n85+W+11wqydwtPVshgREvT1DK3V34+Mb/ARzuEFR5a1lSk45DmI0/
JQqxJzizzjs7Xfr8gAgFlCWMd5b+LpDDma3HDJuUW9AT6zmp9AfdLmC3DVbisU5DksptlOa/IIDT
Th9KFI0itEcUliWwjJvTd38mbbIPd3SKusyG2N9gg5jtIyQujIfms6Te/g5RQ15+JHeoUbaXTmPt
cZ+PT9O7gdWy3G8E+RarEfBhyZlSE1VuwUxIHrTfb5U5IN4yZHK+8nNrO/AGJBMZAavpymygn4Aw
wcm6rcxpUPIXSMryA5x+smeKZm0zXVOXxR4JOEVIXrGMM53wJOiCTMRSuAhSaFLntgv7Z7IUQM8k
5aT+okt2GB7Dlu2pNpiG15/uxieLbF0njZ+aFr4BsRRx0yXhSoCK9rOZ1xntdPrbSpQhNX2c27x/
1+s9NJkRMzK6uYKuA1Eh6K47FHG2FPfdWRsYRgfSkdNGK8KzRJDLNkycZSZ0cJJhb0yV9kZr9XbS
bpL6ID0gZDR9yAjY3/XBfASMrAnLEtPFtk/JNeTJ9WYolAdXgpeqYh1ODdyvysH9ExmxpGXvaYrg
Jchwa8GWlVe5yJTCHJKQfwT7ATByZNeqDhtdUcwyZAZ4WpbJN+Vi5izFkLc1GMmrNx8Kc+pGK5Y8
EyWCulwk4b7ZzXna21lQzUKo4klLzhV0gA8t+xQMXozQE7Xypn6lyviYzPimE9/D29s8lFiWrk9u
En1kK7TUlUOrbOWrDru4ei6EV/ST50ArTcuyWPfDkyCD72/kDbwypHgUZ0kOn052f8jVNci55Gc5
u+fQFuwMINmf+kqBxUTlfpV+Jj/XHNJYCGi2nSdh9TJy7g1dyrVxFmfFWTUNTR8H4WHEZIZgcrjc
LUwjMVLC4ADirNJ7kiC/2YENf3GVdEvcUsGT2hnQJaIlUXzhtJcC9ugui3AD+aJIYIWwkKe5dObK
aXxFXhtSLTd10OnbRfPgPrJevdMA/XasMXPJIxEyvPrl9US1RUVThBD4I9Y+QhvPjXnigW1r0kI0
UWFgDY/20pGQ/KqbzaMBw6EOrriPXMkegLqzM1coS+IBfHtdoXIyC+gmNWo7Yu25QVitjSwKlchg
G8O/bDGUXtARf7Gx6Wns27tEVTxrSY89SUJdb4/HoB64KxYqBZcz3G6zD26KdUIRecPN9qk+1KO/
YNDX6Tb49pTEVLeMsvfqtz0wSr4DRK9UPr6TWcrGg/+Q+9h3FwEmGYriNtU4wwgDvqcSaqaRvDmS
X02eI+lPRNSUrWHuqryKoZaGv2vUpsi6/eRq3jOmQJ+vxDgoc5Wb6SRCGVU6/OvzYMbNlXFsvr/J
RT1Wc0BCMk7AA6NMnfdPssQ1SE+1qDRYD9XsdzmuIL9v9WeLCSHcsi5qNfK1gd1aVGfGX14OAuqd
o9iMA30FjLAua8fZHh5q7tdRPl3IqsaMITcKuxV7f+3UO8AC5IoOE9b7uK5sUXfjjHnxbsvihOV2
NrJh0Wu+AWXkvj2OE/5mqifHQTyPtgddBpHkTFY/L6JkyguIWcCwgIzY7JR/X/A6c9pnJV2Fvb0o
jSKqXEGp3TpSFT/cNjtGfsJbZ0OjLXrX67Fm1riTumn5ExDZsupIpUBaI1Ke5h51ylFj7sqYQ6Lf
Pkd8uZBwZOrZwKGQkO9LuzyA3fisGXwiU1r+nyuUwxn36e4zk8nbcT5eeCQ79lY0XAGblB7/2SSt
LesJkN/QzqIAMM4NmYoDtZF4iWawZIjz6nLLnqZH7/e+hASeQEInWWGIogia7EED/FBtW+CM06wF
wv8uoQDET8N3scp5Jk4NAsy55ijty7d17v9jnAmztDRT9cBRD4+WnGeq7puHsA9V3Br10tP1xdrm
KqgbN+q/tuzUIc20Ez4n7B+THXHnWvU1TRF//d9AJmaO8K8DfLOm7KKHNYptAVTngk8m8khL64UT
6ZADfsOJB1QTX0eC8N3WQH/KOYh7dVQEJdLT1p5mVPOTK8ccn25Y+31ls4OdNNyeYuXmgr3nhr/X
tWT77TesNRjPRWIb7jUXJlpm8hJPkpT6GBFSNEBu6KeaUiQL3fK/3+KUdtUlWgOmz+MRV67Q3E5P
A8aldod5tZXEXXB+IMDBZFt6dUObI9r8f1zIw64YMjagqUCnlvsOo9SjAcgOm0iECx9OAlzO7fiK
JhC0QijGmOl9GBRqZAoxf7oWGRZ2IYzAuz/rfhziYr9NwzBq6XvrX9kfYX2NOhMM704iSEw04qGc
1GsG0pPiBnkcUVArq0isz6gKWwVsJIFRMZtz9KdhQ6l3zaRgxGerwcJb+ooFq/cEZ9LLpf0V27VT
Mo4ZN5sVET048zYKrapl0yg/hSKBukFAPmMnQzcXtv1jC+6CoYco3nQYX3wkrHPJBqVRO/rOAHhy
9on20qW63RgyboNpnGme6QOCytYlsZfJB/66Md66IM6CZforM2f0yymTdxjILOiWLekLAXz/QEBo
4Qigj+OIxbijWtlbRVMBEFm5K6uBGFNZg9Zv53P+D3/93L9WvFAXhJM/cFfN8/0M3WrR4RG5D2IX
C41m+SIG6vPrKOSioa9t60M8Tlb+DQmCPjDK2PkBfZ8xe6igRZRGVx0TG+ruATAEHjzhDo9B/M19
BsLSz+DIwq1b5j/IN4ejZviWtygRnh8jZGTG1gmuXsmdisE2EkC6mT+vBjT2PieKzcD/fOw2BaJ8
yOsakdYqrxkdckltgjlqsLCkQ1fNIXUhGay/fk5immC9JzKKCEldvx3wBLgXVvlfIpzo/SpqeihO
tT4dwFSNfzmvnEGMvjBX76QXN1YZrAD5vhy5ETJ763QwoKwc9JnsquLXGXyw03njhZk4cm0jNz6P
Dx2tWcrZQanC1s4CZei5K3JEB8auJdEVQahkP6YH/7EMNoIjqZVVTVdRs2bdVe5pZglx5WLd3Kso
kzcwmYfcfmzsI339WsTCh3qKfmoUk8oO4hekPTKQDvGnAB9d6P6fW6qi/mJtXMw8ZfPOObLGf+kS
DoijbBnD9oNI+3pjMCMT1YJfgzwkyeTXzA4bZNAFjyb3YY49wqamnryvyWFEHH7Mn1/PaDp9GmF1
3c+7WJepDX0kY/CODCt7H9WTlxHxoGYwMVMh1iQ1A8Ogp/C56e4r/+fbYC0R5f7GCNEjMFZiprxL
+qdloqQ+hmNc/KzymeHFH8JAmD0CuGAxHOiBje7R0jEjql2RAs2Lz+8yM4z9/xXQuWEwy9zSnFaO
/rhakFK7ncHJWeuN7+EyCG4I3tj0jBQZp78aw4FOD8XmSIyIWI0mH1qBcJ9XnPwziARTpg/oNbQF
rx2tIOcbdmVk2Rhyclz2KPeZsVBirbFQVpdVTs8/lNfNWpWZz/FBbwqK63h2V/uPtDJKdAf3Siyx
kb9Rtwc27hssdxj/iciGONp3KJHpzrpnKNPmt1t11gweF7RV2Wko6BO/YezQpW3V3ySJAs0Soveu
tWUnSXJsTwZCF+ajHkAI53qXL9d+PbOTEOfsOVT+Koqbup+uXX1XoMy8iyO37opUpUn5gWeRJKr4
hjWKip/NmD6QnzGgtfLjTQ9vX9+/WZnwrFkQr2LQMU/zBvViOvxFdlt6vcjAafEfDTg1GAM1pGo0
rkj81yB16BrPj8C1jLn8Dwa0EocHkTUwm81qQfhPDw83PGdD7GGQ42Dm3aUnr/OMHwHU/Gfpr1+n
cPLCVY5hHfTIMfkVkp6BcMY9sJwroFgt0I+Cirmcz9PiZF0GLZMc4FP4Uzlk4g7RdFHcIiMj2ARn
Yc4+mB6cUFCOEJm06SBbyR7FPBAIiWx3sNfksuap8vtGvCv1LaEpmpiwaou5uf4IDD3nrGpnUJkB
m6uBRAdMo3hlJ1E0ZqmMrEsLvUvsNbZtUMbLWOFk9L0D561DLXOV+dVBE6Vsxl+8RGOUUHmN3IiE
V9jOpTL+zecnt6pgkh7XdiALQ4Ss8U4mvsJHaxP25WDTrAqtC25dS0alnZeQ8F1CcHEiK0OC2nV8
/ngwxGTlVHnvGPutf5+e02mxc4+fyWu7GcF6e2B9l55lBzWwwa6+5adSGEjpOZ6NSDuImtFYg4GI
HNsmZD/ZOnz7jJslm6FBX5eQooA7P7Cq4q/8+h/0Zc9yZ3rgwZ/SEYXDhRZScjA2ndg+q9YilIB6
z9r7q3sSn2+qi/+u2ipl2yn0Tm8CScCRZ2O0Ql77OXkKs7f5hjwfy8mkqO7qElw2+u4fE3GvdE+V
hePQLzfr2afCRaByMRPE/j5ME9GinKf/Rd0Bxt5Am4Oi6nsGA1b6P4qlqB+bxAC295sczyFe5KLW
PM+19Krf+YrIzU2/1WVyfbUVDXMr0jQBVOu5GR3neYni3XDiODtU+P6QlT7VJ6kUNNS4LPnrqRpi
nMTTWnpx3tvzD0RjTAvxMSFk3fyz7TKfUKoznr/w2Q0VeHzH0J1rkmk2dL431A9AEri6a0AqUfxn
94uhf0e0pBFvrHAOBp2/NSWOyaY8RqgzfyAq9qnPZBrejMCBI0OWwRtM6iH7v2EMKvK3cdcuhTuT
rzOrdpXo3phkKy0V26rcL+aGsQLc2w9XUJJ/bdf7G0QIHVvOFcDA+N1qwM0hjP0E4D/zovQv616e
CC4o8dCbXO4y/J/MHkzj1YQOxhlLiM95CB9T9M5bgWNlXxfokoeyER9Ob3iqAM/iq60HFAQZzdmO
1ffMWTct5OkcYK7o6q8xrUI9gSYIzR9Mt9TxpWh+Try/IHSbbpzf3vp+v3I4l2/hUI+TKezBop1W
E0G48lljCwpaBSsTZ/gCPaULZCZTBv6ddHOSQZLRjyPMwUXL3Zz5p51p2NIjx6dmCg4455Ac9K7f
hrSt9gKDElQvtInqZXWps2hGs8hqwVQ/AJWKQbFszxvlYg1iCxrchUB+NfAGncpN9tNOa3HJHrKs
nebY3GN/HIAX//EgUMRf/0zAz8wdzJy7o9+iRLQpOFXZC5F2bDBcREKpuHCmhSuDRAbqCpac3OuH
skjvN7HmtopvYPe0QXyEL+Pt/Bc7+ELpxhp7GagWm0MFd7cKW5mk99Rt/qS81ibHzNyv4e+pD9v6
t2HxK3CdE4o5SXQ1iGtCC9BKAt2kDtFi54OQ0bFY6u02p1Ovib87r5KtBR9fCSWmiQDbo3e2iNjM
aWYa3xh2MiMu/as3+Qkm5e18Fgl50P27zrqpM587bhGr2kyUQKflspv4Q1gU4rXJgeML4+JWtGZX
Vz2lK2h8OMC/vzSQROr9yPFeTkKxIax3QqyYbjup6JnriYDYH6CAVKUqEPHqITmq0ZSpH9wcpsla
1N9g/nyqREbJ9UJ8G1v5knrJPMhUJvFCG7zNXDScOBn+d0glIrwa0E5BhdIfPNs9r0yiWw+PMEEi
wjm+N+snBKnJHsZEIEqjM3EuOW6Vqj/JPM4pLXF0/xf7rq0IaQn2gb29t+iSxytEvNGWae9n/28s
bqDeyq/qHcfDAJCLFYUa7Bhz6XOo+GZTKu7FnNnEl/6YqWg3urJCf036/w6puQymtvb1naX08WBq
1INlkYmN1WYiPCRfKkN/N5tX5dySuO/MjNte5CWW/y1h8IVYWTAWJeUZM5tZgr2sEUxIPyR+J1kS
kqbPMgT+qUOAG19qDHiPzE4DZSMAIxmjopb3mKmT9JSw0eTIGogYH4Gkpvcb+C+lAY74Jamn+WTx
SZckytuY4UbbdlJs2nuokASqe3LpFE3sbOIWU3yz0DeDRfCn2ZgUu8ouJv4mivYd2/CKN3913tLC
oCNIqXaG3xV1ryhgDNYu3Dgxrzpjgx5pQkxDVLqNY9JB/eL3kihJKWXoHqyPoAwGoYkmiYRFI3PQ
LQ1+z1mcNDmdrXE3Mv5olaeC0vJBZajoI6IrUjeMrLfvcXJU8kQOZR8sL0eYq4rATKM98V1ZTjT9
W4LBfb2Wy8vnhXUQpSO0XWZwcEB0Aqcb7ehovnnZHqnTRNlxuaG/Tsn4Y9oM4loCLvpDIBjrnGkr
jn522FdYg+7wJKnsYo2ifu/Z1QS737iPGONO6UTmftO7Uw5fCECLULrN6izKfp9Jnbj4KziYHq79
L9LJ5kls8cNDlf7AlCHEppYyqLfG5yxBdSUopn+G5o0Js9CUNafbujd80RH6YQjY+QLg2AFChma6
hTiISzBL5ButcaIPSn9oqjnm7IfMGSShsm8tTCTlhrHJcnE5wU0ehU9LQxOF1fV6DJSy1Xlqis7Z
WtN7hQnLZQbbngJOcq6OFVb/qULDy8qUAbjPzRsJeDe5FcxBE8UDt5AgDyBssjTUv/+MJAV7x6O3
gMAvJ+HwzsWbAfQKnypEtyLLG5pLUL7G3MpjnQIEpAIvIB+veeIWe33k1dSmXjB/egPtKQxXOcsM
B+DL65K70PoYpDmLR5fnPkMOpNVMYCcQ0pp+NEs6XRA+4NwBa1QBwaeWVjCvKp36pHVwaK4wRKwW
jo7oL6Yj3PhN+sKKKy9ovsunuNE4wDGI37UlXHh1xfkUY2sVaj5C8Cob2TtYVd8FqHt47AlRYGe6
4R8FqQfkyUxH3JZcnx7nRA2R0hHWirKC/dri1ffgvECkKQelUhIMLKVBEg0W/WcqWBC5vh7BFPGh
N9xNI25NUfL8xHDJWj3BdodIGBbsfIJq77D4JvC5DVCFlBue7O1NphRu6RzJjNcEEjKFFkVWnIaC
9tWdUTeE45pBSvLlj9xcIWFJ5ATyw8AV+vys1YJCsGsuMuLpECupLfKQSwwa6xrBNDUipfZCcsKF
ScAoCX5CvKIkmbV01JRKHYO2I+602OIx8TYo5SdyV+6lA9uXtxOeO9/5drFHIY6izkTVTbArrfdS
myQ0llQULKaL56lKifZ0sV3zptIcdAJmj54aXLpV6jmdhzok+hxcyO8r+AyDgsjHP8lbO5XrkhkY
VXKz+tV6Hi1+KoFg6boRXUGRLauXCKGndF2hLATItdsFayjXGXi1CESHYSzD0IUo5htIkUJz0Ndw
QFlVxnLCtU25aVfTjkht9RsjwYkwkas179/zSF6Lnjwelis3cBwgVtf1+j7BFwRDOdYqoXmmXHnx
J8MFfZ3gNsCLrXgnAPb6do/orjK8jKUqcORMUsK5GhDTO9XyoTLmwYNMAHGsILNbpp4/Rntk/or4
6cLbAw8Zh/g1wZcUPaYkKDPm46KDC88vqALpkL2ZL2LgHE7UpUZ2xDDwSYQEjSAZXwTdc5CqRA22
MRyq0Zy97w2C2sAfv2hAX7BrRXxafq+jbaEMQIBxB/ojs+ufzDxFuONhkjxlunN3+TxAOpclCUvs
8QgNt2CcC+JBDYd1AuniI1OMqRmGCxL1b2Rrr8sPuLOGNImmf8at92XXZQI6Yqk6Zd7IRWvew/bP
ssPP2O2zdVqTYoCUkgk1qgT+I6ZbrmjRjjvZa7AAXv9TpjQLvtDrStCD4rSyBUsU0afILkOowNeq
9Gazq+Z5RgAZlG4WWw90BkCRHMZgdZdsMb/TSr5nWcE+7javfpmkGCL/DbyZO1zsdxK2SBLSy8T3
x3/m6kG+R2bWeA8R3V8bZRgsakZ9aIHxQ6sGs0CjCEhsrXmRFkCxAsz3EwL2NTNEoJkYLnSuZlhI
ZEnTOJBahEO4HBi+vCKMSwVIMhS81A1a9Ft5Yo8GolVgO8tLwexk42GdieqpYgufWqUFw4o5rrqz
EmYusM34sXV5Re4knmCpCWvxxnORND2eCZoou4jhLc7dRicOPnpiRfSvE1/uhya1D/hfXNRN9jj4
KAMoInt8c9Cce2nM6ph1bmOg8WleMlBveOn0qRhRljADojOeuOkzDbW9ELP7sw/sffztI0Cm3WqB
RauZWv2mG+Zyd4rsc2GmxDU9v3Ya/TsJg+U4/FKriyEHFS7nWJ1D+r/l1tQhQHWiu8bH1JTirnWA
aGzBiQmX4Aesqvx2iEs9iTB6Dmd6vbJm8vbsMRzFMHij22bnl9VNPFso2ILi1XdIP4NJ+CDg1Ps4
vU16hDtTguu47ZdJQLa3YcsbHrps6c0RU5NMfmrt/3vMFlVqyQz+iNKnHBWdt4XoTJqobO3SRJkP
aZLUziRIdx1bSww8hdFyJhrshdKKWNVKw8wsD8iVre4oc+N2wyWNl7IWJT8vGp53rwNHL7Zxx2/C
9by+B9GzIBMx6z0iLKvA6hFSlObBTVR7AIjZReFNy9qTsmM/cGXu0yvlYamc9ixScvt2LTA4H2GL
ElPa+BFtruij/nhk71VoCyxfIN6AEIb2FcngMbmxIYxqlIU6dYwjSi/OigVxfxkb5erJPMr44U83
XY0J+svn4oyocG7wn4MZ2T1FkebmxGPsTkbYZv9bPWaejq5XHBmTr15YFhIcmQhZWPLryAOTqSOJ
qYFbfJY85WT3KP0UIIYi8WXyCWXduwTDNve5lDQHJVGZ887gcefIO24Mbtc8BHAy8SeXHyfynoJi
ud+nvXVIqpprhh293PKK7ixZR1CJzy/gpu0lPnWjLTgOpeb6p0+jmyJdQrSaFwtp0q5kihFun6Ra
XwgXNqexth8zCPAjJl+44BVyzg92i3dnkl4MSh/Ja0hMsn+3HZYaBboprN13m6UbRM4VPQWuZ2fs
TLXa69BK4airAsVMR2fF+Y2o0M3YLMvBUVApxP5ukytuN2NKgfMXfm29HAv4didxFnU+12Jp37GV
Yi+7cx66C3rdoIvmr+sRZCXUrHL0PD9LV1vEuPk5JZMPejSfTFhgPqcNCns5JWpfIOdtRSSgJIOA
04e/ZehDvDTFcdZdxk/qLHY4XYXQD/7PWUm2rgFkVVKKgKMR+CkEZE+x41FO/g87NlgMh4XsAc6z
Sa88fynfWWL8mIhHs6odnS24VPb5zq8A8jnHp0Pr540LGB9POe9RniJBwTxa6ZnL19v63DsQVfVL
F0iIXAPrwbyeYMrPeUqs6LgfITTtt6gayykwgrHAebskgladg0vmwISiQ075sj4oUxFkxekqMoU9
y39ToC2oFolVDxH657lf3/unYUcFODvdDhn8s3OJzN/u8k+IlteqiRu1FMZCEYkpzZTYR8kml4tT
DxmzfJFvAr2B+DfIumsM3smzQPzVdpiemeEDpZZOCIWrux1rFzRnID1U4+KodQrYPkgAVLOkbMYo
zDLg+zI0KcKncc6t6OYHBptY5FMcU9BLOTeWTjIZv1kiF8wOa24cy1SLfN01fsZAJEEshvxxpFes
jjThxVuGEFBw4ZVAFADUjIXzs7Q4vIR7Acz3jiYb8xmjhrVb6ZJiAngW4RRrP3jilj0LGZqfhAnY
4PVilfU58wxIlL98/S9hVY5xGREwvGiGVrpj4G4yDlaW83MouvyJPX2ifi59Rj3kuusKnEfYZ9Ne
1R5i/9hqg7scuZsKwQpdi1jbQ3QHtgEp7jwTwWxvNhuYn/as8zX6hArtsv+Rr3mwIKWoczUm2xR8
DizIjfDSOSi+bq9RsGLrchrttXrjOlUqSWDxNKHSFQ0P8Q+rDaNzcJixcfSymlvnnQgTtWJ5h5PH
0gd2QUErZFDNEcBtrpnA3GvkYqliPgT7N13LDi62yCL85yEYVvwBa+knNb23FlVrE72dncwBsLzU
y1vMN8ae3SxxZJ08zCt0N0WcO2y+BE8h+7yth9R8/nVzfM27bl6TljmClP/cf+iiGfFHuXt0qzei
/NSeVCrf7ju+iIf3XFuUxI7rif6c/VFXBdCcqLiJfyhLygGnPRK2xwqeq8CT4rlOLemoQVRNEhTP
tbdCKPzXOQ2WGNSfCQKibjlz8XOnV3X0L/6wUVCvuSW35ghMYDHQmC8ASDQmYhIgp5mgKHyUCGDd
2HYv1ScNBmJfy27guBHp8AI6y8LIECH/KSeQaiyRMqUSv6As1/VPIRDWTjDRJiw5AdmSu2o4G82w
GfdTaNgp82IPlOQgDYIxnkfE0xg9iABWAnUob+uzsq2wMfhPBem8thaISx0cpGDZatxvAeqzSdTO
VQdjauH3IhjAwLKjToTd9R43Worejlp5P6yMzsjYCIlv+Kz6KhJeVy3gtLVEaJiPqSy/39/kS+LK
m+YxlM0Mcnzqic9dlumV8Tnfi4tWOOQlGBAr0bJkA2W9rPXKWylPypM2WKEoz6hPoi2dB22eft+S
oxRvRcEC5wfMe4+87kqpELjY/OiemkNcq63U+qTTJhoq28cZWgLVmGkHZi9eTVo89YlJbKlcd03p
0Fwz411uaHPRp6Ot3S5X2eVJwaiJDrqLmB2fEK7UE+UKRJckp+5zaejGx+tD4kA1hEl6/P9oImtH
qHXTzFaqhzU/A9IsgC+3hyjuBcnZNYMg6zMjZA4EuFbBOye4Q1OX/ajaiodNcyjyD5RWwM7I687i
q0PwE6tWOsIWiBTzzBPT7L4n+oiadtBFlZAauc8+toqGuRwlpXPgTZGedU56F+QqjQimnDIkBkCC
RPnHaKpqFPB3382VdxgfhY45JoVejyJuAH7bt+M19IAGQn9fxrfy5SutUg2b5DewvwszIqICiUOK
yYjLO3oogfyIES2NK+l5709ERGOvCSaTWXrFEI85FNDQjRPUNcM8EoGTJuwMrH5lWMPic+3/+V70
5M1iGigNkyuuD/1UBOJ5mbP2XBUVfJFBPt+bE4OknFRG57Qd7/C/Bdl6/umG8W+YDoShLEfuUK8V
jb+tmOCoUderHjvjwAQj92yOsG6aKmT2mgKFbqMO4vCFcz+svvQwZXePj8oMH5gOUh2RFWDYhlar
dkkR1z4KS6zufPa0kQS4NNY0f+zJbACLv0oLaJjmxW7BGFAiFba+hyZ0MuD8n58c3gLoQgpFzwu8
vsIfIO9sJPMYqXZ14ucTJk4G9uh9rn9BOUh0tDimpOj9uaDG0mTc1vClj7CJgI02PX/1fIj4nRwY
yxpear4TcdLuko/RTXasfyWbckz/AiD/3M/T9QHD7KwgdzpsQZe2svnF9mxSeYko0Mk9804avD6y
TJy8usyLPk0+xVdaV/h0RZ1LW5DQJDToDTDaSYhYQW8aa8LnGYu0Bxl+kHb5nXo2/sKg19b6Pf0r
ImD/bvJYbJEfhSYMihhYLdn+EPvz8iQQkhJxRw2DjcHuak1Hb690ynEc7WEc1zw+Dd/6zD9HVE+T
Kr3Gli6mDYdA0SwOGqKYrfgCLIe6LaVNbS4b4U+OEa08iAfXj4jFpTXjEwa62BcihffE5WPHY3DU
o5mHG/3mtDdFujccx95KnoEbJkxB/SgHDqLBofDYpTjPJNv0dpYox7Lu/huHk5Nfck+CTp0Ghbj7
3M5ODctX5F4JZuIcbeij+GuqFbWE9S7zPdZW2x7dmModQ2T3/6M8kk8SAIMkq5CUreaM2o1PJ6KQ
HJTH7aWobp6bf7ULVbmOUNL3mdCXknRumdu+ObdQW43a0lHkUTlv6sg8oZH+Oo8oLLCyCG4tWc1i
HOGKh8P6gPtgz/TkL9ey4L7LhIa6TUhMBYZ96aw13JFks5eu7S/i/8Gm3CkaM4yz3+EODD8A98FV
O6eBtjGZSB6qsRvJP989AdIo6CQNjDgIbpChrq9Guxr/6kffLePzfypPyTntIhaVmr3+Fmjmlah+
1Vy341xp5YdkU48UufMUeOSpSSjwoykFSFLu1A0g3n5F/8vqW7HY0xMZBDbvvRDQTffIqmO1irAZ
CpaBqzzJb2GATMuOOAyWIZNUVOaCONJtO+e/R0p9FZkR+dZH4IE8MCgW0vzAb1Km+ltbtAyDUlKE
NCiJ6UDS+HoxoUwvotH0rk9tney7fkeW1ZzGY1X5cLMk416xOjmxdlNcNmmOE5YtKQeotwOlXZio
mEjYegS40ubpsi4vQEMNT5ngOtbEg5kAJel/5inxuwqkquQuhjRX8SQrGuOXL/iTsyjKFLzDjW5C
9NHJX5xKrP36M66MHD2fMfm9XBbqlz61NI3nij5LFXK3Ar+MdxXY0PaNb0cz9f7HdWR2Mn0mzsC0
8SSwztu7nEI4wSeqbWP1FdddmYtIj8VkXI6BW2n4C32OrNcSa7Gnj8mOJzv6VAocMgYVhY/UkgRs
Rzepnf4lJQhVtWXEtD7dvSnpZxshVzdTw4GjCn0plgsWXDw5DJcfQcdevVGXvhcGHTvTodU1c/+F
cipOoIm9MVTswaR8ev2JvFCX99kZb9yYqYTICG+uU9NN7dbceVuOIyacL5oXyiT14G35RU9i9xsM
lbQ8cclHg19jBIyMzVbjFgmR9TCxJNqPhyYNhlzrYFk9HHbhfmIFouGOd9CqrPgHpL+lZ4o71v48
HOxETXOPAWPyePnPBAxk/PJrZjc1tRNAgxujdNQquzY/S4HuKkBeUrOgtvSV/ODf3UAqSZjgAD3f
YGYnwyqGA3uYVEoAG8V5cKko4CT1F7lelQnb+8MaPCGgwL6UEdliySTwipOFGtDfTQsQK3JdII+8
n/D0tk1/J4NYttV/Ta6tCN0hZlC7QPlWdjaN3QjE1iwoQryUThdNzupQHRJfEnwtqw5xJcNSOeeX
//vUqV9RIIuxxLNzN7/Lr78kTxwWwpeGcujQEl3sFblXLnSwzMhJGROKKnq1kD/swfz/8HHdZ/Gt
5Q8g06Yr7hqottsoPg0/oc7fc5wL8nlyKzG/DTHrVhgoVXBzHomI0ZTS+6XSsRlcwEQzSIiIxZcf
nyuXcf/gVWwxX+YC20j6QWcA3xz2YQHLst5JNpxjYEDbf74QOiCtZHpnQzwX/KmWvXjCKDmqyI20
vqzeZ5MlswngG3sQiqz+fpxwDSAhF9m6HLaIs+AAkw+4jG25J8BrYg38cdM8MKqa819dAq0Ps1T5
E4jEBG7DWHsvK6Anx9Yh1u4/UNVtaTqBtjmVX/ohdWCL8o7GpkcS8ehSy1Rrpx+bFY0vRZ2Qk69w
qikw2k9CjJdWc5e0N+z0Qrti0j8ILjP3JkMmWjBl36s26kCUtLdFaSZMSVYaGzp1ffJf7xupgHmt
WXy7efuewTQd4DHnrysg95aCkGcN7ewS+Ca+DZvepWqBeHXFU7GEzAZPkrts2t77AMPycl/F0R6p
VoKf6pTDYnXUWY7LmYUqkgwH5/xm7WhVegQv5PzTNWzBdaGNmNDthSyxZKbjkpNPzHv+jeXGwesz
47bSYy4yD5mB7WZVTTRBwp2wRsa2s7XryyiTCTcZPg1pKkuJoAhT7eHHtxizWmGyH6D7kKLvU/74
WCqWsvMW1IyrBcQHzKp0hOG4npW0jDXevEb0VnNFYH3xmQbMA62L2a9PNouBGGGZ3Mdcf7JdGIsw
Hy+czULcQM5j5XbORN46MnsN46lyLP6JyXjlav7aCnrXrkr/t3KaIqv8qNuXwRL8u7h6aaDeqPV/
DT3BrxSjtTHnYmXldq2eDSEkYfpNL67e9s0zSol7S/ctSzUCkW7J+N7AUTOkbaoJFp5p9dK7S5cZ
4gsD6hT7dagEWgDa0cvAd7RcRXEUEcqSkMVw5QDn86ULt73WPrfsoyuPcVn0uGoIn4LetidLDY2P
KhbGU4M7KZdl9cUEa4pf0m41EQ2MQTYPzRVwZe35IjRmmMHoKw591X0XZFGfix+F2MJz8ABjvj2t
dejDwn6bd3780KOVsLCTl9eyMzwneL/Tk7ziikAv8YIg9fmjp5VKSPrEFfc9uB6WHaLm2MLy+VgP
JSFejiWr+JY3wIK2ssyLdX6569ZVNtwD9Qgy61NF6zrNkisF/1lu83wAV2CMzE0oOHXgMaI/frhd
8sSeubhvXW3c0Wdtt5s9TsKt8Arkh3zYjFZu9WfSdfNKSeFdDlFmr/oA7YK+CIoj64TvcuEngSMj
1q29Hek85Y3k+JFtI1aaus6vqCtb24duS2pY8NSZFcE6FBZbdn5/fWKS+72qDO/Xm1JNkNBjaXJ8
gTbOo6AmcObVQykudkhmf1SxyNy5OfawNAhjzMpa8xoGPZ5QqcRg27u4uyM0iEbfdanily7uaUKR
a8g88aqjrb9egOSGGPUIIsT58sjOzE8Rf6Wen7M+Xmq+KLDEFSip/5qqfDIf4SRIwQE0BdfWzPkf
jvn5+QpYx7v0zkA45H4ibX0aVJ9eHjyiDtyw3ZLzRpy8YO3h0Moz5Vy97ONFIe5OC7eJ4+HvE1ME
sytGXwGzM897moL5pdjjpGac7DiX2/ctde8vjKCtKU9R1x7t9IybdAbJufFPM5e4mglTIYQhOwSQ
3Aijwbi7MHMZou4hAXwoMzz1tKBoGpUaqvqKufqmjcoW0igoB+pIUuXbUK3DSfgn/Bkw4zy+SR5E
h2i1S8QFKD231fQjO8TYlzrf2VtaP8kkNnYu0LimFrp0s4nR44GFINbVE4Rt4t3FfPS9mZPgvV/3
eJmIh8czXrjBZMxpzi+XpngJn1TXycApcz1Im9LtVet88Jcaqi+lQXc8JuPSdg92mZmMVPEV3ZNu
0Jr93wdtD/upMsgjR7dbjlril7Nu06wcSCORkA7sczfDLQ9IXCgdtJ7WrNS7jLyhUlncMzCO+uq8
RRQlzgp19iy3B3rMhjJt0yJ/4jJ26uItuTTgNuk32dyeyCa5i8YjAskx0mZgnwHyzsPbUqWgvYcE
cMTx7b73tNlvx5CeOScyrAGqpOMGS4ZFlK7vj6r9Nozg7Lu824HFVuq+7a3q43Mi4ArCOKWsEJhU
kdQ+HHg/ntXcwz/JEQoMBxtfkcMeWNywgJ7QWxfIo5B2ep/dwRuK/gfpMNf2pweSPSlgZGClz+KL
vRHWjgTqqz9HIhidfP+ex97HBcVpUpq7aQ1jV1RfrTCSPurr4YKUGdJxSrxGYC68yi2VnLvmEyeg
9lpW4Qj0fcXLZU9XA9kDgtT5Hx79GlBG/9DhQ0dfZhgGUSstjy193yXaZNpD5QZpOhQRzro6YgBD
KpH8i1Zwu1C3Efw53LF+FRZZrB+dqWPlrS/2d7D1ShPFVW0rM7Cb2tkdT1xBi4QM05opYw4GXfiM
MNwmHA1iy6FhTVBBWXy/VWdMOKd9FUB+zPXEP1kJZOr7TFtC0jHOXjNRn/z09lqdZyu2w77yhxj5
qB0y3ilA3CAEPZBZs2NbpoBvbDtKs+ksozm3OXjHUy+dt0wj7ogVLZAJzsIAPMXVaOYO0XasOjb+
sxOCC1KQbkMzJdb8Zh3FOerXKvPbUnlxuWMRvM3k+f21qPSy6xktZKLb69huQbPXt5b4g/Ytlm1P
ODE9QGzZ6/Mds5mUonvV1DPcF80GyzCVUunrnfRh+1jTx9d3tYzhwseZTQtA98s7XfUUUmzjcpJG
8zDEPQygvpNlZg42jjwhJQuIjJpi1cRbtUA8xFoI2JTZqPkURXfpKt/4VM9b0aUGk3EiE5zQhPsX
SqN2oS9K0HkXjWdW/ougytrldnIexKl8ivkiAIONef28gK6GN4aAm2gh4mpk255U/Uox4aFa9z4C
l/fZ6s6TbUtVdVi5qtWYN6S0gHhh4HSre7aFPuLCsoCYfaGNLUWiMMT4eRNWOhRYdbUEwHCL57nH
yABbq5i2sUSm2gAaME8UYc5Q2iE3XZCfdKbj9EYUuZVqQ679wSEasdavF0t72MJhRfeE8NNoyYT2
G3Vunrm5MCmoSbEGzWOZaR/dXQrvB4ORnpQ85ZvWSj9/znU8dEnR87NNcBjpJxpObmDBzd+xRX7R
2AmLQJkYrg9+6vc+qNIJtm8FZuh6YawK6BGbyIhGPFPVyDIEUudndLO938btG2rGXCHwPO8QqkDi
iCI+GnKgkBI/VAIUP3G1MJfIV1nAOWk86+z40E7wEi//9wAbuv24vKmleEJ0q/jxxjUfrwp6lgks
4veg7GoNgsTbxT9ahfrp+VobF289SJFt7SMcBL2k6hIJLFN9imA31kZxSutM5SnUQBomhQP/lbtz
8XvF5ETSM5oXSOOTvWhwZkIIDK+fYXL9fmLCwC5u+SWQBlcFhTa4q/L7lb5sLE0qTDpXSJNsi8Be
unGbz0wUKRgLplaEjby75yPyaeKG+EyNrm9lSz17LIorUlY5S3dpoS/c1U0xxfl2tGQtaC6IOsuG
hGHKvYMH4RTp7nUB/uIQUsYxHTvwzheTSFXMbDQjkwOIFyyeVPrRkGgpusSyJuAihOaQFUmJecFL
fuIQx8qFGkMzDAYBdaUftMRIyj7RWIpcaGPHbf7erNK7RUq8GMv+wUGeto1jt9EPrfHLO3ZC5RCg
5O702chD9H884i7VEBrgcHF51AOJ4covSIaK/AZRZXJDSR5Hjt/A91CQa3SdbkVl1DEOTZTQDttg
/JtHdGtqwzInnz/CK6NqCRWRQAHRrHUPmKyPcWxXjW2ZtM03+zXW2ytt0UPQ0GvKL8lTfunr322s
qhw4gR4siEjg9ATlCfvYtzFM1SkBTqxLl/rAncPc/Vzaf3tLRIQmsoDv0iDUI8Vbsb1izW7tDoW2
l4WwMGs+liNygKmovBFSBgoep9YAYDIM7XNV6gFEfuBgDIs7u79tHsDNNbL8CLut9M8+PVO3O08/
dRtHy+bh3DM+9q5mdyN42s7RQlFtzPrZQ6qcyw2Xkej1Q5r8g3n8H1gk+KF7qf+PB4OzswipD5Hs
tkdImoZUEOsHiUNrQqv/JyRt2gxFJY5TMCwzwNAxjHNeJQzMdSNnL/FQyLHsi2WFrI81W6XG8uwC
/PNG9q4jqoccD/8IUp9Ir+Cdx4oMJfpDAQfIrlscMejIsBlrX4bjFylQD9WAxe0u/YO/8bDEvU+L
pQUTEC6BIXE5ynIS+p4vdP1NLNOizAI5sO89YZzvn4s6UP7CbQE2FFepwmk13UbNEmTG4xjbZVkZ
npy3xqssvfM6+ezdn3I6nwULNAJMJdt5/nImmvLc/INXQ8klMCE9KVZMKhhbwwuBqo1iyStx82KD
Ha+/jANiVcRRLNGKIzl/1o07uQ8jcD3lhCSrWiRe5XDYeibGTPkelAJmfQWZ/tT10EkXQFXePDUX
yL5BQx6qS5g7J2uA960vB5agO9dUv/89AQx+I+548iCvqEZH+3hxToNw5gI3EmFhYsewvEi0Levx
cylNgrDp4RSBFIELnbhyeMT0L9eWMxRMwpYsWckUnTfiOkr5mIb7Vyg451dThPtVBoHn7P+wZKLZ
k6LH/6qYT3/BxaGPHghv2DIXUc5oN4KFdgW8fYvrqYlsVANbartQKdYNYsx46rCREXMprIt5cxoj
fnxnoPzC9utY922xeKr9ikwTuX1qIt2ke5d+IgC6+Nfn6/LJNKxKuwvYWG1Afgbq2Xr9t4LYJO/u
vnsYZy7f2rUzQS4NwWfpGeMCp6YIUfd2UmCtCTXfYzskC0sd8eOd7gnUU+P4cmQyZB4cNA/AzU9K
SEIzBl2qgpOh8b5QbROzs7SjulD0deXtmGbBesCNqcO71GN6M1I0yCHZjMpm074cGM4Zt2Jz+C0z
R+vVTO6evAeE+CflriNM2OUOCGvwtnDzdiemTR1xKtxRaWONrSN9ra7CVBG5O887QY9Hc7Ap+IXH
dDESRdjFwqmQj4p4UtTLTnbOz+XeuTJHG4q6liUOcN5yBUV4AajrOrX7HcrL2+xtohUI+aKIb84r
R5YQoTpaYCFaRfYjM4Qjs9N4fE75sEo+O5OlHI2+32SRYoOhp1fOLh5vwMsJbsxutjt0y0jkGCJq
VrLpYYg97/YxMHPv5WellAvh7FZRBO6bvvGraPmHnwExKyuQZaWFBiMToZ3MpKOfNbDVQcmdeU4f
xGU8j9iDQfU1zD88Pa1T8wEOiy9Y/WjnqqLoPf4LWme33F6MzkWV8XTMgK4Q9ZvgCkrQh7W1wFTF
Garr0GscJRmpXeZgvcHkw8IoQ8lO9GfmnlIlK663fHzka8wRUmxmX/hlsD/FzYGp5urbsDRHNO4N
DMb3zfXb6PWQ0y8Kni0l3+A4nq0T7vGh821nS0d8LWv0wj+1pQQy+FmB8dXrfU+5TJMtQauzrmAS
nnxe6yTSbHMDY7w7KWbdtUqRzRHBuctU4ZNpjSFbcpaxvnHJyUEqpUKcOHFqKaz+akOC9tr47TA5
ckpXL1cfi0gggpOnAfPiC31T4vIl7GUMjTS2AvUOdYt2NHEV4pyvfzyxqTc7RIHnVkkzDF5j0rNA
rsOYuneiy5xILGn0LaWUcW+4vCJsAQoZ0SvjKzznwqPsDyVl/YsLRudcGRslVVgb7nymX1TVrJ1T
41Z7V0NOWQpVF0ALce0VCEj1xlZrHw4g/KQDY3Gtw5MkV0nLmiCbTL1L44c3Zz7Fi2N2DPMMLrTQ
VShDSuVlYcgs+72LcnyMQQVxlBQOWyBKH8B8668EtZ3xXjSih/IvIXJ6xUJYXkuiQ7qR2NdPX9e1
0aqkS9AaLLcrLtaLVHmiS1ugIFNJcD4KXojs9EDoe0hDSi3jNLSFeQlSE3221yPv8nDPuBcg234D
wT7A//MYJrGtRLUAnELqVNRw6I3DNNWKKs00VC4f92RBzIF9s8rBfChnX1lBkQaXjurJzd1R6iJ4
EAk0dvkE3k6pMTybliVPm7RSHFjHpRYJrwjV17M5dFrNdTqjJAXdR1Ai9k/EKUwXwy9YW2QFRWLe
J1/evdJIOmIDHJiwDKra+xznH7AanppEKU4nP8u5CWXSKWGXyMd5W3koO3EV+0aP02QIibhGRKxa
hlHvyaQYKkQBfI8JBnl4J4sQ65b/v0NYFYAiuljB1a4CEFD89OKQklIynMQfdCTB4/4czY+x2/1v
l2xrxzpQKB/ZfcSZZuozCBENA9bBjJr98N29tPDWWgaBZtgbIuXFL7fhqy38l2zuDrQZ2yQazfG8
A/j+IPMYO0WSNCoWyB9N9+ntcSrf0N2fbeH3CNwHPGUqRJKJjQunrksyGUGLn+rMZoENaZaCMTQY
cSVyjztulYTVSXanZBub9BTDi7tnqxcZXHiQOtacm+M4VEoQHMKLPpZv/qB0EEn6Q9YQ0Krv2t5B
DwmZF3sF/LTNmSqWv22GoW9Hsn+9BxzMUv++jH6Mk6EQbZYcol2ZsVx14CaOUAtXoo/UbhOfX7uD
oIDvfpRpyxcYzgN/CW0ceNLYmanbC+cpMEUp8w0CYMQt8Uj2Ukq4aLlAcHsrLQwysqyi+nbYpGjs
L4inqnvFT1bl0wu4Rqhozu84XCzycSvGjQtwGo59VgaTz+fCUapqjBgRz6K5azCuVCsgSqQ3GmJI
ZyAJMHG1VB+IeQMX8MRLfpQu2TU6Z6vMWboXyb+tG0RAOJcKHa6v4skXbQEuqMDYn+bOi2PpiOWE
Ier7w4ib/UCCpjV+p5jfxpqVPYYWdt1FihVr2vXQB7V5V9OAMpUXU4JJ5NHiaFHcpD2hv8QsO3MY
dksuR9RNBJATD5Se1jJstt3xJ5tWiqsTPA3M1ouzJDsAqzIqKSwLUiY3sbso6rP2/ZUwQYuyOq2f
BTcmZXT+x4l6KlYQRxBMDJ2VSe6NaU7G8CD7xpFY353DoivXfwH9dyruXTFFQb9QN5uQbarYNyO2
GrnkuGWNX+Ip35BkDpSvuv3gT8DK5X7thXmwp8g495phzyXL2T6L/jO3nqttqbNxQ3knab1rH0Ht
yBHKkpPNvC6XPgMB0NyzTJVNxeUBoFIi45kCmY0sN/XLrehfGB5l58h2V5SMxTbixSjlTA3owaLy
zlxuwsoLPvKq0mPP3kIuGtMoXaprC8jDNNk96umTOMrsWgxN0SzVhvjrw+Iv3vymLo7DERlcgTb+
k5OzJABpIyBIF1BdTTCmHa6TEy6uonVw0I9a5CEKEgx5l7x2RFQonvLhRRpWkKZAcpRwNbGP/tAU
ekSQCp1xssbvuu8MHxagLXUB6R1FAFfkG4rUBcjIIf5AS7k4U0s6PD1GBGv716On95bxUZdDQIIr
1OlYbKg80FBSfP5ufpwb+pEbyAvPnRYMfCkHd1lbM+d+DSpQW94pMPL9AgO6wPzeABLECgOW4xSD
Kx2VpV7bAJEuE35mwXAfCn+jGG3JTnbjQIf5Mjfuk7QQCx5y5GYFM7EtXpOEzUFORci5PiJgUDAW
bzyALTaAZOmLnbhbsuqrwO0qwc3B4Q+FRSmlnjwuC9GslZ/iIeIUutN52S/I0IikSrxTpPvo5Zaf
T7XKp58I2OF0Ta7yQMzfKLhkZMGfXClIJdxxiEo7AuFvXHQD+8E0Xd0grx3Urblb4+Dzrdqkx57B
BWWpH/cKFSvJTg3CDKcaI5UgriadUVGn813DvJ3dgWhKXMY1M0+GDsWbcaT5E/jgZFsnKO+taYZT
8bPQukyUD2jtvF8VMHdGsqFa7sJPeqtvkR7Xbks/PEmFmqfckvAurUFjGQCYSIXDjHvS/m+Fqqhd
/d+Pc3Z3koU7UBBUQLUIlkv+vZm/J3vPudRpMUJ7tSMgknWyD5MigVquaKhhURVpSQr10QNz05pd
KBH4RThdBA40DyUtevjRF1NBeZ4qmjDo7F3B0SRaQIPcM1mJjqwfuv0GlR3zSlEYAYJ3QcGNgW2p
6D4UfZqdByx+jFSaKTvATovxw2TY4eNtVkvkv351LMpbNxt02Ld27zEbqFADoL+syN2gqtYoQOn5
6MsfryVIZ9bgOVA21vpDamvHW1SK2p1XPZpwsvw+V8lEebas2JNM48N7J54E3sgqaMpms1rTA3ew
l2SRZ8vq6taSjdZPlDRRsfMYZIrBkYDf0P++9rxlVSQ6KeC5C+TG5MvwkArDY8WUwFMNN/XiJqx7
JPXL2aLXr8cZpdE8mpLNuBiY3nPYQn6PeWkuozQ3wRmfeu2nVlYJMfML+S+A1YWLcKU+OlEBQLWw
9fIxwi6P0EFOGcPCqj+PemBnrI994s5RuzsTBS4zdiA7uVcyHTr96dvwST8noZtIqL7esOKsIomO
5AOFsmvxGPb8bJfbL1EAFhLGG5YWcNa8COyXrDZlqYyuWpddjiPmIaD+6YF0a/sXO2DK8ndvnZMt
uVHkeTPCyqGs+6u0w4PyAaYONooDKIRxMYU5JtQtEFsUgBKhPYEyOYXcFJcjrVhS5XxWeYj9X0oz
m3lqdCNf1pEVXExRzq3mJIxMeexqNKNi/znse/uVjN46RhgkvqBV5Hr31kGUrBjsHs0UPLQMqJAa
pkocVU8sdLtPu/e9tq0kcYpjn0f83E9f+pJLMiAs4tKIZHRsX+NjbX10UYoQ2ABa9/OJRgYUyIt/
HfI/OfszJ0tMyavZZ/M1rKJ/SZosaZnAulxCNIDEBHkaOHyYgbQ0h+JLSwMRIoKQm8TuT/BmT4F0
u0S/vgkIQ7F3Y48qcJy2veAB8UI8DuQA77JcAzzMC3KNcNVcwtNqaEtarVgGwyUSCaj+oztt2JhD
V4NURDLAn8UGMWSqiv3NTUXboBCA4P9oLgKhnpMFvA21b1DGGOLCmFXTfSNojm5Z99Yr4NgdtuIk
nqb3rWV8ed7HgpyYE/zl6vdMxmCHIiUYDtlPKTY2I9bZZVxHsaqtEsWuKg0Bn5TSukzvTcaPKdAP
LtoJI1hTnTmuKcCtnFF7Qsv92Qwsw9PIw+9HACbhQqk9fNws9M2jaVjGvOqixdphIrcVC6lx50Lq
Oc8GM4SfAZ7LWt08BYf3THpmqmuXnRbizUPv9+k3fdOSj3bJAro+NaQOihzmQXFDPTMhPsIYl1IC
IalZp9/sf+gSjXfwfaO2DcqtFA03eW5QSOE9YtfWSi+ZIseoyTtz/6GURB9GNtO6n+LXfyjbZEDg
Q2TxPmqEkptY/x7cQlnr0n+ra+jhHUG1Kk2aOG488P8mkPtfl5DjfG4R3C8ljXz3EmL5g+sA2KSb
amA7PhcY7o1JRi4Q4BvbG4231tmliCXd/Rn6vLQD7zh+ZhKYkMzN6/3MxcCFareHQiX/nqVQ7JtI
xz7HGX8hKKkPoOGXANTpJfRcYPVXLtF+soV0YkmguaSlKM9PLXtkeWpR9ofK9oqJgOm5QosYfWB/
0QvJnucjqY27NK6ZbB5ellGBVU+NZ1z08RU0ypXiuZyU1sGOYJ/TtpGvRGdGMd88G9Avn2gFl7xU
nWK3GYbOT/XMXJV8W5d5QIEpf9S4387bQLeGk1V2jRCyrfaV2U6klm9eCKGE2R6ntG8iNYvQALN2
Bj67r1FjsObhmp4a/mTKcYPAp8yhjoDZfHOCUOMPP/P8RiVWdBC9yOtVAmAI6NeqEejlT7DbCqoR
bHTZ4XQMvJ/boLuoPklrVlUWUbfXOE5njkpeS4Tb315L3Tl6BfOk85SkvqcCOjWC3D7tkFeXaZQ5
7SKWIP3U2qKm6C9lQtufIzSrI16YZPUWbgdCCx90p267gTqDMQJ6cSTzcCjQOUOXxm4QMUNMvRYJ
3fcq9gJHvXd3vet0AdvBphw6OgznpHSllf/3ZvtauFbhq0hf3dFUvN38CiseCO1OavJfm7K46DSO
MiEqs3vq/9Wxf+Ju6DaC5Pi2M9VRl913O2ApA/Q2CbvR1HGQZ0JvZNSH6kBsrw01N31TpaQ9vh+T
l4mpcbGTdGjvZadsYEcNxQatlrsjkcrH4y1S7qPi49RcSd8MyvsSFWFzdunbbL/Curhefjo7P1BS
6cu2UUn3J9g7nwkMQ2lnLFWEB4AglpV4WE/wE3DRBV8XegBeSR++UhlAuLpS93eM+TfD8e/cef8y
Lp9vWzVNADc6ttq9Qq3FlRvFI3X4i7YRMn7Ri2Szv0z4M7wt/YttMzUNRJLZDTE5q4kfQvdwhrSj
VK3HcEie319d6B0NVZry4pd2+w3oAADpO7q9VciL5Wfinb4wVctsQhPABYcLrBdpicS4WvpzbsJt
jdMPAEGLODaWfYxvx8Xkm9emNiXD3M0uIY8HnV3GT+EIztMw5oYzBA1P5dsCNMfDIpRs74A5Liz9
lS8XQDrCT/R4QYPHi+cX/W8P6nPuUlRDys6WoyqooUHxNwm1X0K970IrYQZrIl+ukepDVG8oT0NI
RnA9sYSaoFAfJyuq8i3BaI3dt12lKTJPCwd4VB08pqc8Tgn8FSDFXrKL8CyUOpxFixt9LUhTYrkA
Gybl44ulGLmjpZzUvAHqyxc0BEQwd26DYGxft5D7oAV6uMhGEkqOqjKz4Vb8WKxYed2898yxHPEP
T5ECEEuHK/PTe67OEUZvEgZZWT3sXgMSB8dYenGgEvWyRSr84m1lopKgqFuekmDSy79sNEsqsgdy
KO/UOhMWFRjtFlXWLQniJATJaCaZdRfr+DWdwTAqWiN8aHKBldOoHa77ODlS3wX6Sei0NHLiiJvk
SFiHQkuKIXTMcZBM/+6Pw55nuVf5WP1g9K+7qjXG7WbSLr1uiP4R6R7QIg972+4xbW4BLhKKRkwD
hVdhxECSp+uUuSXJxNH11m2M6Gaa61G2XKooOP7akSRymBI9vz5N5pxXeZUwdzA+w3T14BWhr17Z
WUYyjR7TFqZhsLtbUctCJF48ija1SY8EGG1tBjbjNAy6/BkLCrfPFSUw5XQ2i4hRd820Hx+qNK+/
FEwP4In6zLBzr2bMtWvEm+KKWhGli0XHtX3c2zAPaXZ/rHiFgd10rMCMmXJJ3WJHVM50mr8X3uqx
NNF6g5XsRQAwtuT3dMYsA35TOAKZq025qmxMF6cAYwhoWJGbm5ZBKaGYj5aNRqzx5Ok7koucqEKx
gSGdnonu3EKfYRZtvBHbi2m+VIRcqHJYofaGbqSbv705/865JEvzuFXbNo9XevzZ9q557p82mPFb
RGHU1sgnGB260iVRh7CA4MTtMS+qmfyNg1ENGXRb8Jqfkpr4nT3+LIKcGygjtma+0hkf/lZGdgTr
n1KHpZa04sc1IT0HyUzlNG64CToodI7+kl4PisL+2WNidV0EVn1m3IWt7yisuN5SN+Ck641nfRQh
JYJavhq9DExtuIk50NC93R0na2plAG+pEm0+MhYXKi9nyspmS8xOwwAaEqR1eemvdr8a5wtBKQf2
IvtxiFb7Q1/bAASS5wkePpZ1tpd8072K+IuNkr5DuCsvs18qiCagxGwrWIWNxlIaP1NMKuygZQx2
gjnPD5Wi+m/9LdYcetP7AHbA7SuxJPhQmzzHdH+bpTJPxBYFyz65exuvOzUFeXS5mBcV+aWe2iuW
BoQDimIlRIAYhgIVgR+bAsTD/DzPM7n4wHTkOs5fKvOteFg+gTMaIqOqZeB6cCj0vaSPgI6i8cuv
nNBk6Nx1yECYckgwkVXcVQmpNrmlalr5ac+NpyMc/IEjlhx9jFl1SLZxghzQe2J5tKFuO/F+exJW
d/zD7Xng7f9TgzjCK6F2LGVk6jQ0dLZKdq1MP3KIKwPKDISy/bVuic4Kz3QPXTVIyLg7UV4YSdhD
xE1mjev/3lwJAPkM/z7f2YNSeTVfdiPTdda4qxGf0/UkJ4irq+yxMHIPJgortyeOOcDUVSJldKlL
SAKuNuR8I2VgeUHnmnr5ThiJqaFCAFv+5b/ylNl378MA01ibGiGC8kafkvMWE/QD0kVPvNktUhZ8
7ozNPpr6WYZZ7im0TbnKlsX0kOIwz8eAvX09EGWZ1F9siyVwwZ878FsBnXFGDFgPKLEJLXi6lTlQ
Y7DYPo7riWNebUVes2XOW16IWEs2ImBPmFkC37Uey/r5ddE54UKQBpO+M2kOATNJrjvGW5pUiY05
aFc9sLqFbHiVpp7EuSlUq0WN3WISjKqGjH281zjJ8Udew69VRJ3aY07UdQNPwKjEJP6RW9a9wu1t
yqmaqYmqyYChn2DTFlZQ+Sk0p8N/airClen4+npmrUoOsWmnCDIZUERkB9A+mKhf48Rgo803rDqx
jq7rClIKIqO6awcvBpcT3lmiNPrMM8nXmsIx1j9D41A32f9BaQR+KI7mIlLUupwKyjWPmW4LVqoQ
d/Cxc+vmXb2uFnJtRZCK1LWoLfodX9gH5FNaW73ar1oOTQjOEnZs3vYPfacFsXmpnCRfKMV3NDr9
QTKT+ajeixHsysS9MHTl/vfdkl+HYusPy3SjECS4h6MYvPjUhGoL3VAkl/xaprOfFqRyLMyTWkvm
RHElu5PMgH5uVVRvNyQMBcUf1OyJEc9clvBBlN+FIFKRH9Hbffaw4Of/0Ku6JxMat4yTnPWJvhaj
IcEQ/IjfxZ3PusF8+5uLMdEo10zDqpSPVcQ2Zu7z/9lvR1b4Wup89VEiTX48wN6qbU3kzv37gGqc
zu4Kj6naSGuYvq0LIMgNkqVAsuJLpjeyNb3Np6C1bmGtrtdBSFY+MBuoO38+9OAKOjX1qK/ij+2O
WvwqwmvkYsY21YeZQhs1LhudgG+V1b9EEuGiovkuc3WOkl/ydmFeNbg5I50M4tBxIONhnq2+vZAd
J7fSRPCV+p/2bEX6T7vhZ8dElqPhRry3EBV1gWBYYG8Gl/fYhYIlgzxPPnRsxJVmvrKr6o0ptKcU
InTRxhZ40Kev+RaYkZCmAfVl8TG6olrbcwRKRI4JjndzxNwlhuG/a54vGCQ5D7rfJPtQA+llPFoR
+IQx6GZCxbkB4DhyYECQ3Ki55gpGRuLJEFYQk3unwxGZqjy+a87MTRMVENT0V53eR8ti/8QX/YIZ
Es82Adc6EH0n6k6373adXLjwmT+19RlvacBOypjNCVx/Zi12J9aRNjl8WHG8T3v9ZCwln5qpfEQE
m0RLeIL0FAB83lIjCDSNMW5eDdEHgpC5pw6SsATrSgkGFcUQFWMR1NsrlW0teil6fnM6maByVupt
uXii0i95KJ1Q+NFZ3yoTi0/sD9BNAYSIA6n/pjyjLXevOnkTm4Pwn95Gv6KY1TwLvGa6AzFFpys1
Z/3Q32NX0Z+9bNn+xS9kFpKJlAl6LfO3LKENrEwN0E2HFYNbI7uepiwSG6WAZKeSMNsdTylpgxLl
imTjFaP8QbEg+fzdK+xr4+277Qcid8sgkYbEtZNnnlkYohtYO9Q9mf+dd8pDmSffPnz3PeC/sXhp
Ckkn5w0SqkdNAwU5m/f0aOvcRWwy4X+fjUW03ySlJyIlv8ZrHtOXhl/Xp/uOwtDq2M/htGmidext
+Gu/pxIgx/fLr6JqS9Kmtpdc4RDg7OEUCX3jVX+V32pOsw8ko6uMQAxuJGbOTT/6Zz6pYAhOMKQ3
9wSIxJy9wPIfO9MWkvENJV8mMPjTnLed/b/T8/RCUuSj2EDUC/lh/DzO0v8zLD/iqRDqSYs0QH6K
210etlr6HejPGTNxs4LK6G1qoElu41f+lmCTpE7w+kSrSP5rXUtw03lsVVCBADBc37N4LcDay6p1
YVKUqGGwXypZlOLoTezTF/cyNjFD9/GPpE1x1Q2iaHVR2Be3/DDfJZifhkHY7EW4pF/k5RTuT3dC
lfrBKZLmKAbSnsDKsaz/oGZ83GWHVPR+WzuZo3ZeQlmwuEshVf1NVgSW/Tgud6qNjMvmqzf5vSAC
U+s6qpG+fdJ4ObDV4E7Yx48usuqlpncT0oCFs4poH3ZMwDMQAy4bbhlmLX+AONA2u9xvFXgAKdsj
YXLwoEyLF9MhNJ2pT5dZRnzIYnZNLkcyFNTaVUPaXQnrGQVf/4OjdoyIGaYEB+lgcpbL5MAtPk+X
ZoDDjlJWkWslSsiaY4HUox397YMTD1bnCnCsTYxAKmfxuphBG65a8nCLlmJqINsMUlkEp0H96X9P
SYl+Q63b8k29cGSaf1J3v7aQMBXjOeFaC6OErnjBN3RN0n9al5xhIp7lrSIAVO5i6kbnbWeW9W1D
DEnInIQw1Dk5KDIpWTmlPTBzNDEjvdgqafO9x84GtFav0fsO6MCaz+3I6FXa+EsUJcrQsqZxo0vY
phekXGgN/bXbdNyf3H2rAPkNnuBQpnwtH4q5q+OUtaBuwd5TVxSwEFuX9wWKiBSMaR+dqkvb/vNK
GvS10yQmD23MXWMFBdxY6dfFBmMR0Slh6EPqtKvEtfxftZOIjQoB65p3RYZdQRTns2dd3uyyH4tn
kWxzyALHTDlV3QHDsOPkbBkOutwSFBMUq8F0cTG2dNklLjOQzjULZo+ztYYgqCnvUQhHDMO4Zy5M
WMJAZXS7GF8kjuRlx2XquxJqeE0+3xXmbmaYjDziytZNKQrwRMsWZZzOf7AUaFEZcYB5rDvFGC/f
gqzY/V1wW2wW2K+WSUEdCUqB14GlhtFvsdd8fYJrVwgItsOlD8JqfLjp4f/4qaEFNORgUhwu0mOy
86WVLzzgdKAvW0llSvhvEgRPZPN29wVAVpsvHB2ASvSbyOeNyR5vivw6dbsVwhGqNNIkEhWmDWb0
VgpfWQiLVkt3L5/i17al6AN14S2hnjdeVPdiHbXe0wej7VF7LcXqPBr73K//r//trErQHbgSMRBt
HW5xtTxkRi6hbz3rN78Kcip8JIPiTUuLSDnDagPyqhejdBF/atWkQjKJEUq8vx4UNotUj02ancbP
7+e46CH+6L0+7DmY7pYsU76OMcGxqnUQ+vOMtauEFFycevOGbotR6gkixYdYz452nCoZrnnYBkeb
cVakRUAlZCx6t1IvixDSHGuB+QThCRu/yVEGjYD57mfKglf3UE1bQYkPORSkSJsY3MeIrznl9pYf
V3MbKOBqvBxu2EY6t4dgsytnhpYuDtpHUOOAFmEtKUYV+h4PK7y2O6eTD2krbdcVwY1VMi8abShW
Q0yIdF/IAnjY+600T+9+4xQa7Nf79F080QJO/3255iOgcCzbzuel8bziTqignEsIW0nopsExxyf/
BxPY/0q/erlUwM+sX1Z+XSGqERHmXTMnqofmaIJSfJw+IdPx68a5p8oi5fKvlPBNLQjgCUnp6bFY
5S5noQ0VsBAhBE+yGCMrlJfsOQuPAFQ6sKFdzI7PiVspVTwqzdYA7Zcx/+9hStfsvyN7XevwGMI1
7l9udrZfgsltolhys4DR/R5Fz19G679DgEaZcnsVNo7M8tXX7nh3vqqBNXuyl802e0Y5I8pz8qEc
ECxmzP8guqxEx2iE8JHukYe7dyj5q4gWcmGLbdo81UFf8DzwU1sMpxkYNDl+CfOJ1LJV5PA/31VY
+tTupPyaC/3KVFoV7kLTbfsvcWL1YXd/nsShB9V30Q81igpQVFn5k9SfKXptTElC1DJzsvIJnryl
J51lk2kvOC+k02kG2KMGEzRU470igrdLjR2sKsJ7zq/atUZ+vRjJhOFSTC1uHnGUxjY1uuYWBi9+
ZHZol5LNT+Y5CDy4dGxgSqUzWcr1kVBhyArPtiVZcCuAVX7egOu1sDL+Kyy6khLLFgHJljRisjwm
uDS6GfsSLtyGZYpdaXdpepTyZjcPw978cSfiXhDjPgKIlhtuJiD9HM5nOnJlqgYkgHZsWSyQKlgA
XRf7MF4zXIFF+SidxY6K5LJejUsldIwgPqRBldSbNbaRmGEtUHiIqL+2waedZrnhdHiAHfBehN/g
aBiRHWu3mdnU95XrQBKxY8VhAupGv5TgevL9UPui88Cy9IXu1KS2usfAbV/2jgf/59VvLsrRKNEa
90DEOOpe2Rmd2gsbW4sgucmYOx4WNipQOOfMhC2dWHzjmtJV1bBxVPbPeqtRfq8CrBTnIIf1bTxG
x7gT/ZP/jXUUdlfT1j/XyUVTmRx/nk+kv/jfylp19l2SL7qFlb32RvpI332mztoypM7Ld4pimeMU
cRWCzI4yCR+iv3ZOmaTwdqtBnXYgET4GxBcQmtgNC3aIt2cKgbhDPiTDr6HxNXPgwft5YQrnT8So
xEzjLTfFzWumZKxEhHoMJMICUf06Q9duMktg4gvkH7GfxD9obDfnYU96AB8D0N9wRXgCE7O9u27i
QM/DtyO93y0VW+FuWhlZ3r9h+Ii1hyiIZ303vBUDeUvd5aFKWrEFjNuNgWSpCNhEnLA+jHi0tqWY
WgkaRwu6rj1z9JLBRn59fMTR5XplDSCrS14t7w/jOurQ68eJaxI5ivSRWNDrPn0x5sU2npJild9y
kvWziHpPDEi37zC1hm2kuGDPbqgKxtrsYtU5sPdIg3D+i34bWd1k2hPPKQ7FSF0qE1cioI+SLnkQ
PKnWI8L4iHOlgGmZqxNGwhDE6TGC7LIW/cv1O6KdBMZ5LFLhn0oIcZsw5K/ksSeCir0tHzuKfYz0
onx/wqpoZ8i0DO7YqghaV1BztzrCWMjKD/vSV7r1vsMsCmZlyBFCCALGp2LEdZ7GE1AYrLPvyYpl
Iqzqy+8DoITxeRO6kgz33qac+1lVIDXosJiiLak0Mx9xziAWsW4NlV7itl9Q1MkipCT0hnaQoDC8
fRszHPATxvcjzC+hqbcDCfCGBkne8zZ5X/mKJngxLooy5x4ciU6Q9mgMQ7mjzk8vK6iQM31/hX6q
jiUmaQDDKiA/WWO8dvFi7xHSJ7tINeB/KNWR9/jJrRx/MHSAqzq7ZDxWoYdQlYXYgpPyAbR5lyPh
Bq3g8+gSSPTCynvjkcyXWpXkTr8n7aJ4f13NjzSWyu+5frzRgTwjP4l8+cO4Wr6t7e0kVXCJ7WIJ
Oh+ZHXwpvJtq5Am+Pm20SLSCv/streLZ/490JcLw6A9uzwkQrcdetiAf4U6jYUet6qjM9i+fAfXH
8E5cltGkgX2qhFbcxWeF2N+7K4RNoNy+7ReEweLh4ESUZ0rYg14Wz7lwvuoEWYPUIgDYWfJ4sDRg
Iv9mIKk2EZxSqRsNFZs++hPxy6AnuWMFds7VWpdPU2JqWu3+yIe3li6e8M7y07Ds9mm9/shDq8Vi
ggq5LPEm5agcxIWRgEARYOGBxLj+MJfkEYlffZvK7BUGScjcyqpNd7eRqLNy70rjr5f2LdVbBI7m
SH6ZSiSlNjV8fy9B/aAmLIkVAtGaThZ1Fy8Fu2X+ucqBKLgwWY7FBdzQ4UVUYBYGuX6gxmDN67OT
cjeCVhGptUMyK8KQMMP/uVCe9O0Z1r3kNV32P8q/RwE8uEUldQPAY2U659L0z6MrPdeeMjvWxMLx
FCquvM/+8oEJyZ6V1EchWs7CmBv/WQHl68WJSXY7og+ep4qV4H/P3AhESLgndemtueQ6XKsWf8lB
pq1v0YHZlhEl/0l9gG+J4oBB4HrqFq7TVNJvpi08svwijv1uTe8ldVeDO/hTB/QTLcjSOQv5h69/
G+WoGdIQmqE+k9x51YJksr55J29vopRF+RLRQrXijYxwnQmEAmYYIiRBgE3Vjo+pmU0uJlD0SsmR
jSUz2WeCiyFriOLGpja151YydztPC/8mzfQWSMGnIY29k2oEtLz6/zfBqkDaFrTuaxVu8g0Lggiz
CJ4xjecSkJElRv2V/JvvIq5hZkf3uSlGcQowIX6D1yixGsKatP4dd9jJleKLs3t8WDgQk9R49A7a
8ZZy/Frr0i4VKE3DBd83EX7AQaSvckt7gQ+Tr6JX+cfFLbznJVQ5uI8yebSLx/NL54yuN449oiog
1LmomR410PZOFP8FD3E35Rsbd47eWF74FmoOLgpscHUIrdZt+NMfbe9sjHu8OdnNQN6W+soxFUaB
Gy2mSMmAn9LTMHhtRp0UBf78LpTsWonCw7kVUBDWhgHlM4wzCTEdgOlHt7/1utt25AFKwv/JiWlH
KAaxXHYjtjJ//ctLdId562ZNh9t8+3fMgTgjbozi0RCVbG4Kl9j1fCjEqrAro4yFbhpuaSilRtc2
+woG8fEjSYikOR3nTxIW2yF8z/ZI8mOXgLNmRCoddOYdppOIehaUeh8DCe+E+pi3mhb9h3InXyad
+HRARYYyvW9rLMqGHNQe6PGDjzqGH+wZtjaQp3uLei5bQQzZUOipY+ktcd607CuFs7ltY3e/2sqZ
QQtI914OEPSe4eGE0EOt6WYo5QWtRe8fF6Eskzm8JgNcMQWmbiXyoJGRXxM8INbxCUNaRJ8GlLOR
QKVUk5K0FQFoUT5waVS7pnom7w5yieHHbyVxk3998C/hGF21EOKeo6SquNbfyMxnFZ3Fqr2AYDHW
yxR5IQshkljxvFV18V1x3Sjz8hNgQ+aqFdQZ5qG02KRBO+0s+kje502pARYPvLubshFFeChjpdNt
MAtnnNirlEtPXQOs4kdsX+VVcDKoipP+1HF4yigNxsmaTGldYosN7vZjq9/xa0WhnUitFog96/yh
/THZzn2B+pxazPkGDZMHEgFQKTiyob4uMLML6De1I8mJOjyfbHlOcvkpXww+mkaNuoH/yMmjAPOW
s1S5rt647DO9FMfVS17ONbwh9km0pamEWnp0AfHNK+Ty6xWJO2qnE79ef08NZT+APAlBEadgrZoq
0djja2UkZIRRqs2xAYG1HUQXFT2ZIpWXEP1erN5Xn8eRyQfKAXug4pgoTvxsA6VIFm7rZFjwdqur
VKHn4xR7tC0clITQvLvNkPNEmxjRWWLdd4tvNBbO0ah1CYbMp+tco+5g/rlBa5qsEi07hXeXUDyo
VkA8HPYazMVhKQ7Xm8/elOAnbDXIsHg25B32/z+r9KghuY2gPBieMTQXPf/GPgz6poBpZ+pWOBn4
KMRDVeDXgbZI3+82UN+xBAMQVm1KwEj5DC9sL7xmHVKCb233PaEsp2T4hAeC5sZDmCOy5zeqbeIh
TJXOlTYZ7lBH4hOEVrgGodWj9Lh2KzpnbMgccIcdcGMWrwV2CQD33tf8Fq+qFAmQay5D7xqNaDEN
2ZjBTJPo5+1TPmzd2t1mTg6eehetzOMe4bwLABc19IZa5g6zhPSy0MvfTpbuBeynP18ydh389lIw
3yW/0FclDo70OglesDnXLagHt3COfAJsvgf1oPWgwCPeM5NZjbxVpMvX8aMIzlWU1O2y7ZpzlcSI
Luh4jTstPE6IqaZaqAclq9JVNcM3k0AApGMCWSGYB1AIASFBKxuD7rrUPS+kFJily8AxhfVSChu5
KdCwKUXdW6l3PJPh9bqCHH0HaEuJOR746FNnuzb/jR9kiW/pAtGgXvhMRVDb4BaO0U+xNYSRFwhk
aafcKr9RFf19mwsqDpe4OLkg8ltpGHVNElKNK1IlxK9i7EiGYhCwtMR7uqDvHJp75rQzUjbucEc1
18soyYYJ+RZeskyPn6RLsAgpnvZlGFbywvv50tPBeQ2qv9/CD7n3v7IVtDrOdLVtZxJm7bNlm9ML
Q7wx3nJVNF+LtAl31+2ASEye5/S+gZwUxvN4eLrMOT7RQKqYigd7AkY5ehXtwEy2zWiP70DKBSfx
0ZPRr93w5ek/EYbsI0oTcsVp0xaw845qoqKz2EBjjD1El97oW6ipvfvEUxhKuMy60tWUtlXd0y0+
RV2RX9VAMBPQ6H9ZdabiQ3j6dGVGbS1Llg3kpj/S4R7bSt8OTpPQiuU4olcNG3fbkA5kUrP6H1bF
NSPhV7xhsoecvEPWvqvcb2liMgVhLJK1BOJqJ4yrK8i2SNPGHjdmtCJ+POC8wy3anYMbdU4kmmTH
0s0Cxzds6hGC7QiDcoaE1ydK5UZSGK33idBcGeTnQN6MbCspwluFcYL80vZPi5U49B/kgXfMXb/H
o+zUaUvCo89mxR6PBhp+7DhTlwhlKG/nTE666KjfiM5kbQ8zIwDK933fm8ekETV1Q4zzsMvCW0jf
EewuadS+R09AwTsCwK7msNk1z9z9H3cuEUr5VlTdjC6DG//DON2Zk3ZRpzV+OMIzxKfd+GjSyAi1
gCE4fpqbSzuO5CTLVSKdmT+MZdTu+vnsY0W9pu2DRMUXowGf/jyGvUoN5JRxBAox7sGDcPI/KeGq
mp9Vm2iPiBeKWf5Icykn2oLztr+K8pKtYdxMeEwVKHcIp35rXcf21LbiFA3xJOH5SpsWF4PYEWMA
4zgW/Qg+ZIZPbeJ6q9vRLllj66RIJqzdBmIANLFnfvE8x2uAu+k5tGRw4dMOu6IL98JJAXHsZXqN
uakdOBhaDgJV4gNM8WZCXTZSnI7ohKd4MFedTRhVu82XTymo0/IfUwnffsTSw25AQTls7ITvPpYv
HPCOu4v+Sclih9nS+rVNO1lDSs/nHxWlPIcVsmARupflXPzPxRI0rHSfkOmnu/c/W3bZTCe0wDA/
2OWV49vI+upWdBDJhA2bjmZiwvUn+nIojAFe4H1r8+Xts3a7MfekGLTgQt44lzJHv2MFxOONy0dM
lEDsNIQ0n+zKu+zAvaCgWm5uUplgmyNcIj9as6e8hsLUYi2ApQotFP3uEbJ3k9L4m4p6sMhPSy5G
ABkgXaSsdJiQU1lJauJFIeSFlVH3Cxb0sW9nfklsHKd7QkPfgjB+Ww1E5wcOfTqClSO8yHPoovRz
w+AlLu3hRbtKXpC2TEKLSb+fmkEir4X3jolXovXTGa/2n92Dczy0ZRttS+Q5Xs1zntTTJxF1CTir
7M13qIw7QkqJdPmyd8coXhLmphR6EbkpjhygOo10NWJtH1bGcfV9FtJ0SS0SjB/40oy7ZEB2NmV6
KgeiY8HsEGFR4RKgB/KJhYEG8AbdS3FauzYql7j+vd+3dBS8BQblUppw58+MdspnnUJerhbN5l9Z
1xZWhIFqH/FPzSR8AaGMMDWjVJjftEQLCvHx4MmgATxw1KsqMWVmRr9unOy8/1xZd6vmqV8I3ciA
fHGGTh4LMOmYe5W7lRwTb90bkSZty/1solcI/OK5NNBMj9TQjJBc2Xp0223xGkAjGMv4giJxGjIH
wSbDzU+HVyPDyE5i/Fa0Qo2U+7ynLRjeorMtp4wsaJ0CzTWyyfWEeMHateMP9Us9r5uNThNJsSuJ
WL66S7LA+bniqD6Lu1H3o14etBpHhv5LrrqUvgorWUMg0vu/Cdq+/VZq8kIw4V0ZVItK8FkFV5Ds
ugGU2q+fzaBGvjlZtVYKmTQVWEJGqq6LWj22ZueyciPov3ZE9awiokrKI1/qnLmrTE8r+7V0k4Gf
fnRHm2BeH6f0j38QpkFXKDJMNkR3c/W1ECvPPQH2EOwoX1GSHiKApdxeLRAd39k19yQOY5keAIU/
ZThy0i7qtHM5im8QeaoPl56QcaBzDmtZlvM6lBG3EK2Y3mUO50i+x6gEuffRZA62uFTK9ILn1Uru
nX3b14M9XV4+zn8dqm8jsayeBFypyHJI0eNLg4M9MRymPF+kiIWsqwUV0HijMOsFMaIVaUDpEhnW
v97trMA92S0VedgnqYND0GptWuzj2aB6IEYHU3WZTWViX8hikpDBVlEn9VoohRPRFr35VFdy9WUe
8ajqLUEDDjJT6NzMrCh6HmvyDvDWrHB13ABVPV0Q/5FQqWtzHbzjePLLeIHPRl4syKeCJ1Ypqqxf
Ftma+YIei+f1JdvAt6k+QqYMWQ2SbqNgrWqA8JasHjxXWCdkQ4RKz8PoE0Uzs7CJIcjecoH20Vyp
cgyW3QVaHaAraUHd6vrsg7cM5qi3KOczf4tRCr+bDj8G5U/PckLJKaDO6jAGslQvpfDamH08fnBc
zY+katgEBc7fRyJsfpPOlmkhywMkq0VvzrvHWKBWdUYe8thq4y2x35LltrvFpUKImpL6/pXjOMxH
/xYtqSgQPGBMmSVKCf/6BIpNPAGBT9foZ6EGaVZiavfk7SswCizeUezLu9n4zROH5jiV1FcqgzNZ
6dyMjfE+DAmKQqo8yyxkPPArTdqYS4ii5eNkqqUBkyBl/ayXTvtT/hwilU8yVVZPnqQq3YaDEWuI
vu+Wv7wO9Vl99QfQv+bG59mQpNMbGtrksrKc86tmjcKIo0HYm6TVqAFExq6o2INj3JKKn/hU5en4
hrSoRKxwKhetJCmBvhtCbju6Ysfz7mBICNbZHihujd6SDkWaDtERe+862YvvxJTLcy+gyS5joHv/
YFOHFmR2jwZCqjEA/73Z1Y9Hs8yghN89oSCGaT0aNEAbRq1xKx3FKWIWDIDqwnnbHstaaJt0dbn3
rxXW7l5xsK9GNweWj6sVY4TdOLQ6C0vSMQ8xDuhVuq13/MI6Ye/M0gYWTBQhBNRBnwhzrlazApeN
se2pnDr1EntMT1gRkew4zr5GxhQ+Z+caIAdXh7w9jiYDRphlvG0E96ifPIqLw9JsALpP9Rbo84dm
K03JrpXe6DgLA1jG5Q109FIVcvkkbE9VZdA2kgHNh6Q4EUjB0t7ohl0pynScNX7e7yRCS77QkBaW
6IvqXG/8vUF+Z2ikf4pY36xioMzpDI4wXjJd115MYbXLOXP5nkhWfVBEM4ufkDHb2vPAeV1hoWx2
yssNWRvADs5HJAtljmsx/11BYgGi6xLFJ97wNOMrZA1jnfsUzKYwzL+yvJqwdGX2b4o1EsETHyr/
8a4sJUHc/9Sl2/1bIS3WshAeTDd87576C4pjI77nM9nAYuw22mOkRXVqTBaC70iAxjoO64v+0cJz
jtCh9RnRzX2P2hc3v0DtieKA9RkrtWyYrM9EWeaVk7VNAwIjNSrmBIu795TQhOhB3DWy9h/pNDY1
YfdkvAtwIQxN7z+pl8PTM7kGsfxAdwKeOQ25VEP2P1cxUOuNOOwA0vDIbZhQ2kieNmz5ljfoWSjl
AouSxuiVq51wvoQEJIbmvqGsYZfHQoC/tZMQ+73giJoXwitVCz+PK40/pCL3dalx3tFLdKHmCjgp
1fg9Nzl60IWsx+Xc0sk7guQo9HkWyLgMVbUjzjftSea02tGCpV9Kcs3uHPzobIqxZrmlHAqcLbd2
bRPfqNFownB+q01Arhe4TAorcnhOxjJtUhQTuA0qIHG6wcivkNCU7pbkSSZcpwmtJIjqLhh5EuAG
TV+1RrvbHgbT+0BARZlAb+3eEWa7kWwIRZfiZ517vUpivDczoMBeDM05YsJgPZlpaDfQIzrErQpc
XFKSpBuGvMUz+db6NOEq/7Dnr0cNv3K9uE5JF49CeV2aWUxh5sneOLvAFa60c03lh5BErccPYVTp
zJ5sLgAXMZgqL/Zt4xLj+9Qn0u9oPfdtPaFb0dmYoSNi9iM0HhBrcny8uGTX96vznyu3Xx3loSMC
OxShfslDgrifW/CcgzUWV6pBVKg0awyIvTfyTj8Rkss+5lrh/k3ltISdLeHfMwCJMNie8p1M6Gps
Fk07Egj+jJs5ggLNFEcKl1VLukmoa3EYaovluBEPCKmS0QcOU0BJFO/8+w0rPorT6dHVrAHVa7mh
jHxW16zM7IpeqAzHfHyaRWqShtIm70HhrZimnJIvYLdtGqsoKsMDqaMfW8EKn3ogtD45L2MFf0U+
KLjA2IW9ivTQ5fYz1TplM2mJUrbQN+hYpKPEKC2u03UysNzeOwMGpdyGdl8UImW9NYOuu29lwGzM
ZJwYCLdxBq70OPbZ4HChnHkZKC4fvYEBXFIAnVd277hwNDBwvlBebfO7Ah7EbJkqoMq88IZSaDgi
9bbpZPuJ4mFaribxvCBtRrqElcrv6hdNnMty9o+sH5qhIY0+LwPeTEI2cFATuhVW97Gh5wjBv5GJ
1LCQwvUOgOakraTXStvZJAx3ykJNlYaTPyLGyqYagqDrHmIzYYtlg0R41US++F84oQmTaBld9tsF
hfReO7mcX43J4OUhRVQadf60nSH1ptkSTFfYu4rzmPZVk+h6rfcc7u6fiMYQ2ZqXDTazjmPMnvSR
Cpz/mCnu2ITrv+Xc9v1VM0IlgKpqGHJ5/E88pBv3Il2KokghPNMopVnsjoIROztRzPYJneObbNZM
En3LhteNY4Fh7AEnSa6rMcGFMCZrpRLcl+pI5cVqWYZhXLAWnhlBAivgY6gfCy4vNHDZKTjQM+CU
MWjBTxJUBlAcQnldwcHuSXXS00btPyR4rlxXnhKtKc+gPaI2B4tq/hTo/lnpyYAaBzDtmLxkuIu5
2jfOZItBlFGeRyerARcPPrShX075rXNNo/JkCjj7dncsDMQx7JUms3/IYOOJg26DtsmeaXflLBGl
2OGYYbObu76SfEfJffex8i4OglCjxoHRBjbKJpTLB/nAma08RJGO417kWi8Eq+VZtwJSXW8wR+LV
HfghYXg/HQew30kFhspd57sIsG14FOYZ78ujZqqVi/GBkrrnr3nvnU16ACbtrLo+6EzP/Il6bRgk
VWHQ4coXzmMYioPpEunIoSiylRSlHv0t2TWYyi9tU/wcXwulmi5SrO4P1ISSkBUPBB5mk2ju2dhQ
RZYOmE0Rb3uAgfJMehB9Rbj7DuEH/qOAOnv0XeCiB8DxllKz1xvSYNbPxzTqxvmAtpJXtySONkB1
pHmI/Oix7N32i3RE23Ta3TSDzxdLaeYcgJN29Md92I9mX4doWzTCPVxwa9SkAbz3CEESOw2dnrU8
n6BWlmqkF7vkOxZtgTyKq7jPBK/EzcBS/B/N8RnrQwwDmHyKppt0isOzpblKa/3jvuouPo/Gk3Fv
oICacY8ywNAa4nJeTXqRHf53FhXcZb4yXwCoid+sciIcGouWJMmQgLcn1/xfne1ZfRXjzUGpDDl3
23SO0EFumfIPv8rc+BWMmiXpqZzI+dc1h0Ifsr3pHsJOMAR6b9x3LRnVZ2IUdMfiG2c+n02hb+vM
fRhytsMVGxShi+YedpqAJVnHOftHeMA6ioz5eWBy+OVONEfAozM39XxtOLJ8CNE23EBiVF4uwOWY
oUpkSo/H6pK2JuGmy0fd9ILvfVs4FlOXZM7CxNYKHIe4BTZCRM6TJXIhcDjcoatlUV96B0GqQ4mS
QUGAmPJ8Pi8oUBz9+eNLKNfhJ5S1Wd01AZLQc1aCUDCAwTJ2PB2a0m0evyKixke9TGxDCBLabjuE
LOTt1hOPy3J7oU+hDHpaSPUIyNql/OwKgZNvNnYsLqkRSp/rrtuA83WvEdWGcoqdH2tgqBRoqukG
yr38DHJTKLUyrB2AOsdi0D79MJWl6lJEA2tiX4HOZQ0QVKqGlYcfVzDVw5nwCzz0tyE61FssVt2F
RF3WNSZL4nzkF35VAWZn55O7zqy553zKPkOa6Rzc1nCmTWs4ilUZn94Yln2r18/bNrbMi70CRaZM
ItVy755p9RUhQChMq9cjQpTnyu+NqHzP58ALIvRwBT7/MA1x2GByHd2s5KppEEckcrO6uhaZmMNO
xlMXAeiuClFytvlUQ9iE8QdruqP+1u/Z1XM81s5tz1uFPf0oBTa50jzPOibT42P7s7nmEvV5SLTe
mWfv8iQuYjWcpu7eQyrlXXaiOG7fF4mmdUzU3sQnZDO2S0xylLomuGpQrHpK4KzY0kznkeFC3kuI
1i3TVDcEGvyJpQA9HIvDdcq7h5fWUGbWyEuKF8279QnUyK21W84o20nN+jevU7ckoxAYsmIjJU4Z
fbixWkJZI9koIXyCZ3w0aGFFzkOG6KfKu8eZp/Aye8KNnD7dTh+yz51yIGHkOl4b6USLQjmK1/3N
fO2gNPa6ZG8EShjMbEknNRBqTej97u7FidWYhBKvAgpkabp1agYMG+tccUKdC4xtRLS0B1DfRq7S
48HNcs0lzg8RPuQUAOu420D/PrtctgRAWdG68CbUs2hJpl1VHjETKZ1+1887BYRR2P+j7BO2X6+u
t4AztAxnyemVal+TMbl/GOYWDPuAhaCqOnp32pkELFYrsrqadA3tKbI+Zz+stzxzsmmmDCoH+NV5
7UlK5aooCGawtq9j9IeZKaWfyauKAnw29NsLJ9ODDL5YW/33qkrGeH7SAoqS+sJPBAfe8UgClTFU
buT/OtogL7VHaTl8jPoqRFLkUtAwr02NuX9+5G5qhG+bkpGtJHE61jF+xSKB/0+3ZY01UqTkJg1H
srXPhNU6H9v/mv8HRdownlGzRB5JLZY/oJtxiBcL/fOsKg/ywUNOuZ972bIJN8yjiChVP03iHYjf
qbrURM0BHMOeN77GEpa6J/AS/iNV33JbuebFXDbIAHzd8sopqPlvgBs1ldxT+6u8gtsYSytVsXPY
kBDRgp1AevSD+MG0u8tXwG63pqDVnW5+XjwL/MKHtkBwxgzLJGS0CEWWbz6v+L1yAQ1XTP8Vgh3l
x+mYf/YQQQvgywGRvFLak0Jrks88GLJpb4O+l09U9DZ44cfftZCvf4qG4tb7D4S811SifjaZ6kPU
H86fHVmipdI1tBnjzPPDPIJa9HURul7dHIXikihcjEZUFDT909AgQrC1fLgfDzXE34kn9YDJ2e1u
u6hXIjU+LlGBHPoayOt8bAcO0++yhDN8Pw/KPQ/VFYc6WOBGp7w+NiEho53SPT+hDnHr7nhjx6mZ
ubBa6jmmonWT1ar9tUZ327zvKOdtimKrouWI5MStR0LSYeidO/9Wo2LQD5keGn5s0/8imSukmA0O
1zMwAPImr72a6b7RHZjgWxJV+yybRZ7US8/wEL2AY+FQk1oUbLey1rvld7jrwFcTQ4ySR1SB+6Rd
gMePKKZWOd+oq2aJq0NcYLN661/IHmiCovGlavozDtXdDc6ix7yXVZktOZvmzFSBzBuw+IRl1oZ4
J71pYMTUG9FWYSrVcDykPNidpLyc6GkisDhXyCgznhyJ6owAsrXufeld+mtWblpDPkulzMb+rI0U
u+qThP75uKTNum56OdtXpBNmikFbvjddHRfZH46zAaIclJX4IFimsWRuYWc2oIyDlHDfD4bmmLoK
EIgBpJILksVVXnNtBsYsSE263K7jr3MmqjvdAC58yeh7LbPMCVx3DdQiROBKRXYym/6Q/LhVlUBI
2RXWzdXqPJqz+jbsHJJqL3URhxbPeX0sCbkX7jsCPcwaEw1w0KrElCBl9fvsJxniT+4OmeM8ThZ7
ufncaFs0sYp+FvrMNIZSIa/K9TXwZNwRdQSIUcS/XecmK2KaUGGuSlxBZG5kGDOJ6n2C5Iu+iC5N
gzNcY6KrwG1bh/OAOTEdoV5hs/Z6vgFslem4PSl0652Snlivqtwwa/FEOkESL5sw3VAovR/ghirQ
9rpQ0sNTkn1mmidaf17hoO/bJ1s9FJgLXc6A6XGDLYTEyCPguVjydCtl9s/WxqhLExtF9EP7i4hx
nN2ax17YqbELPzb9sq7hSNyXUIAFNyPgoNSWlJWr5gJXMVBlztZ9ba6kh0puP0JsTg0Ej/Sv40h1
bQvpbIfg9synpPE918V2Vu+nGxeoi2NWkpknDBWfmD3M5Ldn49f6mFVKVpChGBwHlsoPSJiWvxbB
cJ/bheXzLP+pTRHfLOvlJHpzJlLE5b+aSNw+Np8HqxVceuvMkCnZ1RCRbNQp4iCo/EbXXBKJR1fL
i87fM8F5Y72lzSqjg1gPgMQbWvHi/jUVcVvrdXCucXV6jmckJIehXmyfQhf9/tdAklX9F5fp6/Pn
KT92OadUURV+OB8VNwvTJyrAhnt7UUnh/d8Y3hJQhKjQoN02dWUOOKBT91yFUpaBeO3pBQRLoGlR
NnqWsNWcR8J2pev/44Onakc5SCITyT0Sy1bcu3DZ7qqBxPAVUnCkGyzNwuHsCju2RBn1RKDkpjHE
470Cxyrw5Ka/kmkM/L6/fSdDV1XCVfK5bAFd/IJ79gnh042CVoVwEi6HZVTwWWyaYFLCv+f2c/Do
6m36vC1fhQvaJsXTbyfC0l4PC0suAH9XZuWWQSU6Bli0h12PGO4lwOir3DgdSMzql7jOZnA9kEp5
3VQo0YMsLD5VAwNLmXvuXO+Q/oA9XenPAaup8ncFNN7717tO/6eO/NB2tT1RMwn7l59bY8veQKdb
zK3/yFxN9JtV/ugeI5m/W6Q7QVxk2J5wpsM4dOBnEMCdNhxLJfFqD0pQes/gYlItZEvF9PNc6t7+
1xP5VHdA1Xc1nMjRCQfjo6k/O41e2mecCufARSwYmZ+YVHBCAVXnv3pGY5guhtV0Qj3PNSCG4ZWL
DwwKblz4DY2VzErVJEVLWCL2RmCODFXNL8SRXlVrA+v1mEzdWNZ1uWRPixldE6KrXArK/aR4kHRv
bJcrLaOWrLnYwFLW5nHI+lOm9F+3ZlBmAM1H4N8bxLNvDL8UkOrZV0OjV93a9tlsp4LdPCpvPBZB
ZOMEgRTPNWEQOQZlUI8ltbgf63zVRB65vhdoRIND22tiCrSnBHfTDwYxKgHMpaqZZNgl4ZNM4Dse
8m/1D5ux2v/UPkV9J/sIflRYjX44qnPHCGWbu738fwcT90O3V4wfpvVSoVGAGKo41sdCp2XbAZ5+
Ex4hAfwAg/pWs19YbXlj5im4lsO/ySz+XXpWwsy/HFXILXY53nNL+M+xeW5i3SUVT8kSy5oBD1NC
8xP4jV8M2WOZ7lJ0D/BCnV35nHGa39WCoYzWutI5z2zX8YX7itl0ppbkf9466HViaRLu9vD+VCQ2
L24NKxyxNEKlJdfyLy2NCnsREQk1EfF49jJd7RlgkvIeSk/sDeh3tTUPIhOIrqUhWuPyGzf/XIq+
b1lW+gec2bHoYhSK/ZLhpsRnOnYWDiTio228ceywaYzFj3nS8CGPRlWHQsaQWL5TJJQldxBuAy/T
Y3MiUiZNeUuru0cPcHXQXwS9IpEmY0VVszbSJ+xHZEvz8Gti2I5wBV0qthSjGcpuFMhsESB8Babu
MfoNkPkmXWejQxzdCz3Do2xNz6gZUiK/s4miV4apNOzMCa0yzryhrRHcif9Uw0o1b50iAAH7hAKT
r9qqWsCzqeEhY0KCOkHdsT/qlJKgY8auqom51nIBbuEqZzKN3tb0hBR2Rr5FFKpNOmmyd73m/WGJ
RT93aD7ym4nFrIWXzEEfo5thR58k8DFzFcHn1g7pEqhlXUrGnHoiXUmrKDM2lf07CpQIYB0J0kV7
W4GEnOLg4MoqzG1PtVUgTZGF6aa+CZ8rNr4RvlatlBXMXU+PXjivPN0lZZEbv1oBET+DzgrlgzB8
mVdDaNHVvqKDRYUBXOh4OkqTab8IlG1NRg0m743yX8d83LYO6RXGWmANbANRz7D1OP6a0hAuHO7C
Ub5aJYwvJxLTqhzOr2nlKqCmJvJ1JdVC9hs1FeLpF/B8DUWT22jJjvL907pnKLeZi6Wn1j8Sh2hE
4a4wvx1z+MuhROZoeMTAaQ4zdGBFAyLEclqJcJoZopZf7ajLYtxM3j/xUXOo3jXXQv2gQduCRDPT
6/QTZ6+gmE11CuZ6PidlWcPWZCOFz9SWM2MbLGOC0siBgCNmc79A3neVylWyyOxVwjcDm6AfiPi+
6wnDj2fsfO0UGU8Arw58wsxKtY6bL+Xs5kv65Qeufq0izExaYDAiwV04cpGeU/LuaFwxsOmamKP4
a2+KTdfj76R4TaPIP2hlETKB0UZzFQAKx0eiZeE6JJPvPzywCtl8uYSs5ZhM6wdZlnsL0Saqbzz3
7aWgtp6qpu7uK5dJEyKTZFcVCGDuOSfDvEVvX1B4xpLXYlO4AEGQ4hwvL8XPvhaVkEpVUuhx0qen
gGE4wgeLlxYXMrIud9HuweLVCr10TxWgRKENV/vMk8R/V62h0tNKtzy2cBfQ0GPDIg+qTS5JA972
aHuzVDT1OdGCAUahg4OdtHnIf6JGnUFPEOUEwwKO1LRz+Pb/s2h0enQmpOib8rXS+dOs3TL6e39A
TSI9uoSo+oVnoRUq2zib1XbwtTiVXhhKZGACjDOp7ua569CSNXOEWTZtuh5xL+wX91wWNxnt8MQI
1vdiZta+9B7qShXgwcnWbY0dVMX91cu1+oXX22AHpBYPXAt2lG+yl7aa1VdjhT6vceqOPXqV0skM
xI1V0VvIMiLqHe4u3ctJtfsEyzOoi08HgcXCaOyqiMSYnncCyYo076XyBASzr/cYRpbKyNv2p+Jz
PcNyUQMIWlpwQKvRKMzxkJtRmFKhhPnp66Yl3oex5TucKg7xpwjWlrM52tDjOq7J465qJiozcfXm
X9NGyl7+Mn7jRQqJHVZlG9Mj2ToC17qAXRiJW4bGgEj5hGHSl1p/k1Ty5n2bZEeXmegVv1D+lnEf
e6kkk+PCchEviW+7jlyJ+UviQmrk/GMEN/lIsUvKJU2iCp5zlx8jsffTfzwBv+z5xHxZcbQCOLK5
t+S3Uwb3A+P+7Mkq2Y6Ruj+0Tgbxd/Dlr7YOfmQx9afD+bRqG9bff6VXmfK1x13e7OMXjLBT+o8J
G/AMxIDr5fD6SrzpPq0+2r7E6UDb3r1GS/bUAdpccg9e/Ihxj/AS6sIuDsxFFjiNRvjYhtaE5xkB
8gBFUkMBn0SFs5PJXTFI+QSJEjprnNvssHLQH3ygE2+DPnOTAK59hlX6dfKTKcufpAyM6R/T7HNv
lJ64Uov36vaYouRj/BZSdeMYz7a3mgK1f4Bv3BDHQEA1eeLwW3fNfNsfdghs24BExRjaJU7SdSN9
XwWAEstCkrwkurZ5Ea30uoTHv9xk/TBfZX7SP5NLHKQGtxN6a28HhhnK2FxJRHg0dsiuAwWyXnJG
oW8UOqEQX5D5MYGAWH5WCFAgVuUDSkOTderOi5aS9GbgTaeEcr1hDocAiP9rkqeIXN//lTxdouxk
kRtbWt0I1KeHHfcNU4pG2kbUdvOgh4wy64V/BH/8jIsoFDgP28EURWvisAwbHqwcIs85eZqRy1iR
6cUlsHAS50h/YztVuGVOk2YfW2hrbV495BWccs2/P2payms6and3Bgzj3Z5R1IkusUjEYDB+o9ia
oaRjpWKI+QCK6nY07q6Pd2lMAHrl4hwuTC1u93ZAbYddUYHeEGgYJwwtATZ7BR3GT/5rScxYmWBT
0Q4QpwKWcjIwF1jJPbobnpGtSvav5/ttHuehn5J24iQRb5RtwexleDakLQUP3tWDGWciEC20VQFV
i6NjYIk9sViplbjjdL6cwZP9K5Gn2PxHmiuBefGpqFJJKggjtYjCfXdvQu0lMbQE1ilb3wLFpdTS
CVXKchRZ/7xKTXc7tNelSwawYLZXR3b5mcvW3qzoZLGXyOMlvNUdO9KTjEV3lORiUrVDXTq2v1sV
Gi57ZKNAAZP5P+WPlqo/B99qScdKIdwTaOU72Il1q0w71fF8tbvH4JnrvZPg7bpcZkmb3hbxJY+O
G9b8qUhFrJaJk4ocSlSrwbif4u39DrDBH1RPV60aQQF+KPLHfT3fSaSnBxGVLKesB3W5G0pa8lLu
cVm1mSR/BoxwNZUUpr847xAgsb17KFw/YigFSyKTSh/nmfQ2GBV72R/0tIU9ejTsby9AZ3+QKojR
C5Ei5N+mAETQUllrbCt0Qn5a7cyYdeSt3SrMo+5QCxLLIyeKaqp1JR1E3urujHborfU5DUNi8JK/
yb8kkbcImEBxga0Ot01kSN29LRDVLCDUHeT80apKuBFDJT1rtpvhmd/idCnnrgyAgmj72l4vxVnk
Va8hHtjo2jA+50bvHCGK+LPNU+5ru3tX9lphwI1CPbnP/EJp7iSPAYAgLmMQfNXTVFQiG1WiYwsu
1B/C8+WV/oRvS0w9q3tRctkkZaIQSyMemTtbYXvnqWdwdw1+5Qg5eI5MW1CkwAVhHoV2F6jFM4WZ
1Wbugg5cyH7kmLiDLMvenZrKINuZf1vMgQIQN6g/ytNZ8EMrCLxNZL+vaoamxNk68HlNBv9xOO5Q
aGbok24EGJaezuuRwdTjeV3tG1pOaX0QHibzwWA1orLrkkK0a329BEF8IPJt1PtsL6WW+hBZn1Qz
6qWbrqysoIRQ+1CPoMqSrmou1NEVO5XQK9lZCQdZrb+i+bbzVDk4636yTn6pgoiHcpsbUviamNBV
DComiS1nIT3vvFas+ySsV9kvZ4y/WEhAWqvyLSThwKk5hBHHwM4n+sio03610B0Z6cCZUfEOh1Nb
xzfUMpuoeMuutpzCGdQTjMg6EWT02K6bBH5EYT42mQJVaPLGzlcneVf92kMBnsTPHqY66LgypOM9
p89+mMXIFgTiyTaTAOCNG09IVC35Tr9I4rVkKMEgZQeVnv7aa4Aur3fx83iN20EEgwiTbjrERsg4
ROVCRiH3seWM2aRTCEFMRVGTRuA1SxYTawOBhsO/TpOyNrCpPCcCT5mTqC8Fc0XTy6UpkzwFDgpW
Smcd+7WKSeDduTyLmYLtGTIUHV7BS3Y9djPVwFPOCjWX6jKtELM29Zi1lm7puniHU0aZzJu9yMhu
fug1M0CMk9MCfCo8akb2ttLuZmtgo3FcmAbEpflJl2bgb3hT8x9l6rFIB/Uh6Rbb+psa/EqYTJJn
AXNMSjDOr0NrVK+6D1NVUKlPfqLSnzUz+RpG3wd01oD9HG4cLyLIWUH81YaEmiVno/Ss3pEzjiss
YHTWuymhZK/VpWMlb4/UA8iAidAmQnaKXZr/nd0IXk9TfzZADSYMz947eGTV3o4cJqmBIKODUI5F
nAGt5QTB7TmhIM5191AcebiVMHjepnkwJ4CJKFimG/TVbq5n/ePReOt1QgMeEMyByQ1QDEtxY2fT
08Y4O5p1AkRJP4eKhWBlr3hEpgvksq6d33wK2HaX/zQO/XoQM51BHRYyq7CkhdAvYjuDgi+a0tks
HX6QedDaKUcTUi0VGO4GqYGEJfS9dyhdr5mfWcx435nHhmnZMCefpdZAzlxlivgbV92vAbbKbE2J
dGmXd2N52XfYo/M66fxy2/RglVPeWV3f759LDCcUAsXQUFmshIZYoBKoUL5K81RzKzgPEZ/wB12u
taGu66Zh+KnD8s5RoSyOwEZ4ju9kYXjQZlEJ7V4IxZFnAqj2WtaL9EzWPqM227JYoJxr9o7uMpak
pXBUUBKtY90zwrUypmlAL73RNVqUPJnqCVwh6sExMdmyvtgcsBEWo+n2CbhSjmVmP0LvwBIlg+S+
az7D7aTdiZTDLB/NBfsPayujmLLV9/71O3PbG/52cgI2hKwJFzKDnWxCXoZJTnZtd/SG0S1YaqrT
E0y8cnAdBCVTHABW0FXhdRTyD7gh+h6VkFeDY18WyI5NJ4xf4F5XoMHvPKaEe/5iAAeIPOacmTQY
3bucaIYpPHTURMkW7wd30saYmXyEAe64hDjrx7U32SIPWkCAp6ORh6fTytfN3DtOcUAOx/6DdCwG
kWiONkQsGq6hMwxvN3wZhLCW1ZC6Abzs+2YlrYyq89VSqzhQLwyicHrdONZpLhGDTU9jNfCzTVRr
6K0yY7pF7hcVcDFB8PHuna/mkkw7xlrf9O+7huPE3vAWv9aF+dHqaTCu59wAEhDP/k5wowsvK7pM
JZNWjSNlvsXkwfojCEaG745Yp7/3t3hbCdYKyN39E2eDygSE9gRQKSf9gzcYx55JiCVCrgoT1YGd
JJyzlpt9n8cbwphTpJ3/C5wcyu1w6OCr+Ndi5/PmQej4y9332u1iTOBaBTPrViAnO/7qDqmtjAEq
+xwuan0TTdb6Z7Rg8YMuLoMDFFYUDdXWfSr87crmrgEuKVcnH+Z1J10YBgP+pipuJ/XOony4YqyJ
MWHcapBxPyL0OT9RURa5BjaRCFmjJARmP9Xwimy+zycvIaQctnLG/DcveL32Bs3W6oaoJfqZLPEa
DsRnGb7VOmyicPoa/loGJMjsbqvi2HBBpK/Z+KEYYBpMlGzdnJTByp+ofkPazUFANiGx8diOAINA
iDQZ533OuEBYpeXOhQ2SQBoyz+p/XphLjeI7E3WKaO4pEz4ZheNQ6YaTPBLLQh1zE8Xcz6bk7dwD
skKQrkf7cfo5579ufSq5xulk4qBchFEFPP65NcKlqtUh0t1RyPAA303GugNMngdhIfCJYclgrpMa
NWJq5/UZz605T3yDOhvnrsmDTxUMXggErZkAXIfSj1ROYY8k427vIxTEGbta8Sm+9SR45RWGa2f+
25rRpUJ3Flsi529s99IPqwSVy01pN3tPdtPRJyI4dVFP0L2osEFvlgGFrW/nvkxBZgTxZgK7woPZ
xl9JeOiChwNn6KZsDOtznxgkgBhoyNU2G3cM2+OdNfKJgQAsJAqij9Np7KTtiwsWa6w3HJFatAMt
aXwi2E1lR9Jn14oo1gT/9Afr9y4Bbt4H6ESoTrKpwA+OIdceHWKKxQZkTSEYtbua/x6Fe5z6x6Go
hDzY0lMFx988WJ7WJiZBlcJCd1xLMY0DRESnGa2Y1Ex2g9rb2VyPEw2EGg9t54cYiE8IAOgSreza
XIPBpShxZG0EFwe2L1z3tlCrvb1ztnfBOEyWWgPZGBP+WdpQoNUUM8GkIof7CEneC95M6QDHViH+
ezsG2ttwk5AJ9BHT+hsNTT28gGEiGmfIgGfGXWYRmDIP92ldAA82m6Rj2EB18n2ZkiGZ64kq7CuF
qiHjbIsiC3CnKrLxAmYCJFP2pwdhpJPU9/jCU5SnL8MTXSv0GTlWMKZZ/rcHmPMDNJ68ThALVPhR
kqjMd2ZOAfnngKz3J/aoH9jJ1SaiDG+5wRbW9WW269fSo0Cjn79GNdTTbUoRVClP41wzGffXcGow
5x0vggT7pT5sBbLffwDRc4zHR8sy4deSjHBMt2AMEb2hysp9xUbNy0JenEKpyc7sQ4XCrgpWLskt
ynJ7RKZWBqq7cORqLbTs/srOeBOBmH073ufyvno7Eg4BEjWm6xT/K1QCgYVTXJvXi/eG3znuFFWs
kdCOz/mEK6/APAWBqkQQvCiC2FkHTcNBD/3qrED3SgtqERm0WNWflDs1YjSHXkI3teFx/0RTHgcW
tuXlb2ozyUsv686Ur2H2BVv2fKiJaUYaTtoMPCfl1Me2zyXzfGxtcLhK6oPl8trnPG0jGOvUiMR+
5QWEz126YHrKjF7oSus3qWPM2JrBcBjCHGNuPXcGk9l+50n0ii3zs1EwCgDsY5yhSdPugIzfHFxa
PHB9t9iMkFsV9VDaGji+NTWTzAKrmfDbnJH7kKT0K74PH89dPT84fesaL01C9uNUm4BwxifWA1Yc
cKPypdSIN/47zmuyrxfPDHuHqx3q8oW3eyIvx/A4YMMkafIsNq4ra4aHlguNtEqHCvx62kWJl+LX
jUfo+Q7kzj7BQ0ntZnD3wrISHs47gyr9T3NhNIhyluRps451+F2kHeEp7wL76KEu/SvoIxlyQEtX
fY42otJqdirOBXn4uLaQetfY4g0rlbHEJkr3BtNY4RwFv2iGGAuCCx9/JrwMP5XXyRM/0DGZeu68
R9C1yFARZqqpcQB7djfIYuwBIVgqh88S1N4xPqsIXFb7s0PF/P1zkNpucJn7ji+YMIQ7ZgDTtgGk
b+OfanNXhZz9nu86ltffkpJDOuFCS/CMGv7eqDtuCWJbSmXX9kxw/mvSuKddON5zgmJ4br4RwfmQ
pdseAtIPgCzjzwIM53Gvfy68zHOrMzLRmPJzQmwfZ7b71FfECjSQ+fY3KuJdLqwDQWDro1l8gbqQ
q8l42Bt73vxq5bFIDgubjF0vi0fKAMMV5EXgKEqNeUT7DihHg+plL3a8PB0kEBwvNkfatBFwpnBd
igc+jKseVoz5YbYLLKuZ+k7g3Wdq9tZSDwPXdhJI1ppJK9L6PO3x5j48Xp9IKSeKQuXvTl3FmNXK
TKbp1JJvBwEHNy5+gb6mOE5zVyCcyhDQVrXjujw0auqZ3ABl9Zo8JZLTJ350dQijmkjwtinh4l+u
/SGFAFKxKauR47ZN5quMql/S+PpGKvgBRE7jv+rwqe894rNPo307dtDnrZi/lUp8KLml2MFd5M7V
v6F3JjigW3QdxtQP7unA7HlVy+QRpVB11YIhUDXEMeyZOYvI9jppNkkKRenp/RMVlX5bEdRdjERH
wMjNvTbbJxJp1tMC6m6Z/3MiyjNisXM6GeiPWmixZveQWcxPsIDy0pCvegi/uephbI5uWrkRB7Sf
C4Nv66gJh0SRAz0q0G8WSBx1LoI9Ckig9Q1M8Jj+neynQ+AmJ5PGisERKpYSQRObkzxhWuwQZWnv
OjSGi5JQlduovjJCQnGRFZ2ctkXVlFSbXJWzZnX91seGZx3RB2zQZatpXtFc5Vry7M7digZcf4RB
fcfv0htgGViLZwLaurIidF0Y/lEXL6/3bPg2tvKjeZGW9+a7k8UKaG8Y4R+zaJE5nWI4CvWtMe3W
eJYjnyjUJguLiQ0PtRsU6IEuasFxJ3aWbzYscqfwy/1T9zW3z4Ll0nUAYQrpDh4pAvshwNGCPk1O
WhHVKN/PZEXPYEijPYR1jOCD9NMtlwjhHSRPFRUWtcNhDcZB7pDu/njXstFLXrO3Vw1lSUkp1skH
SBYRyMBjmBxVUOmww1Z8PF0HVbo7izlLKaWBeFJBrwtyHfLqWjzt+16BVemrabvRoEfzS8MSNpof
WE6fpq/vSyqy8iqpsssNCW19FcMIjP2/5StRWK8CMrvjfDq0hnlqEKO2aZ1qAssbx/kafxOLjQ0O
U+Bkjk08Hksad/2Qch1FGUmps6EsxwufsmBshmtBChSz3uDgJW6AbvuJwRFBCOLHWLqPx0c2WghG
aSWdeLz1A2o9b4BM16AAYMoOmjNsol64mUt8F/X7Au6q5SLKOVP4T+PrmujnSZXdbEuN1JFwbyCQ
g1LnZHGfshIsVjlATR1uQOlFRSHFDaRwJhv/g3NkITD1vBOxoQVA8a3zNcQZw2HE1+mp+n1gXkvA
AQ5vtdU5XTukYZKddhuCGdrZROxnVf6codmfMU96QXB5Wwh/AkSodr4wmtn9gNm6fUaG/Qf26dCg
9aefapiP62dtyLdv3WwoWmihyMg2CcntevvGaUG74HuiUX8IdjOBNun33G7uFjZqX5WqVjxD/U/O
ETRTab+QnZEsFyOyxMwdNWu2V5G8PxOpXRPjfH6+oR4F+TCDOZAwcjnTP+tXE6HkBNdLjSRBtV3m
V2bHYf2pm8UnWGg/jQMjNQtHjHqyHX/jiHpgdvh2DLWj/gUyuR+E05TF1iJdU+MyL/3u52QL62FQ
zcfSFqrKaF9aPygetxqyPURh3PmyCK/upweav9iF++wmBJgGmBo2RnA9seJn2qlEdONB91HCpyaK
eXAlTqh70GdWmYjpS2aaorGo789cxMQLy36ATZb8Wabci+77XvEZfgIguqNfHegO9nvb3Gx1+4ac
J8QmCZwWLjehbXXHVMD7GE70Xenn+TijrP5PrcJvDiadhcx+RFa0lN4rX008ypy0PUThs34sEX8+
xkFCKw1g35nGiy7noCX9PA3jTmkURquty/07wMMrriqFOs56S7vQ8/jyBGGv5xxEDcCdVKn0OBzi
4uQNx35HhwA7k9LWhg8zxV1x9xK0vkJmU2vkH+jde82X4Q8Cfd00l/LKduDfX+xiSb8RiT2iPagg
WywzNpmEgMCNJM2Ohhk0+69TQtFKHjhJQIAbg3cDyaW0WWosEDjS4SL8u/FyTR49jwxI9bI809+0
1EjD3qV2/D76pqX55qbeiK8NhX57jJIvSu6xnX0WcWpv1enaODfSGnB8EOTrRTySKqj6uCbDOOjb
SXU5qwpMT6jNZzGY+VAbEQ3NQzs8Ge2QkdQ0aCQUJ+1uLxWg+GWKFdtcXg3wAAyl9tXZRxmKVeAE
Tg2VA/fC1VqJ0danYX/QKKVgAgK5WwRTRvDCTD4Fll0R/NLc/hzqj5NfsJ2amlC/cbyvVwL35rZ7
M/CuR9E8fZv/x8ey5wmApDTWvWzlio0BaA1i+GGnIrC19l6S7bA0nv2gUA1R21Q3Ua/z1lqsoqAG
JnJ3uV8ZjBc8cjnStXVtTgbbfoEV1Edam5QGbO/PeH/OoXnW/EGSyuI/FC+ka5MCvNnsG4emNpZv
jWlagyRRgZNeI/WCGxIaZEvlpPWSqKBx6tWsybxXW/3vrkXngbNwuluUoncUXefv4Zl67HYdn3HW
ri9E70bxfBh14yIugKLjWClqYl9ikNTdwL3b1N0nU6/eZqxG/fMHw7kEC7aFh4e/aPZDUluW02iW
WlH7UdNWYeUDfhuIMieGkpg7z884ANEuLzd7SOFxCjAXTEVkFLSN21aMdyZ+2MeSX4CqZYWi+elq
HciJYXJlwrMyIocOb3wg5s0W9oQXtIZPteiFEOSyfrpkErIrDKki2oJrIpG0x6sf6xb/E6uICNAx
PadUnVM/Gi5QKLYgmVD/DW1n71MhTZJ79s96Y3iNvSObWvpDJmksqrdvKuttSJ2raScZtKRi3aZ9
FXl+YaGrvw+PnIgQNEQqMtzgZ71DoaXUZVDysXYct9YoyAQ++bw9tkTLeTUT298FnqdNoKw5RL30
gaoksmeXUNnx9ZY0utD2Nfbh+Wke+49t3Is0fxB78Gqm3vrhtfMvqorZ5Ly1aEhxHkogwlW64GYm
xaoCuTgxEkh0pmp74wDjqtkwE082FYrtkpzFy8PSzcyNDIMT99ND/xv+pjtV9nP62UDYYRVPxIWz
s2XDS8sVBbNVXRFU2Too30ZPfclfS9hSA8UrieHZR6eg8SnIDwb+1jMTz39V4RPcuPC/uVHFaO2X
fJcnJYcHTUZW5MLzSYkvc4MCvptSbGmrGaGWTi4fk/GKLgJQBeF2hXJruc1AcmQU0yCPf8Kgf+9J
cwRvLrok8mFcqFnSKu4/6NXj5KqN+bNDp7GLXClwzaF91Qys8bVtkYOdyhSwFejoh0IPPKx86tGq
IrLW0A0DvGzRWrvzjPP9svuz8l52BjOWzrfI4igUe9B8Wzl2FE3g6JIEINEadJsKmzJ+OQsqvP//
UZIsbMEpl+rtOD1vxNhfZTLyV0N6fJYjtRGi32ckxRmQdIKlnOemfrU9b0WiS4/zxwv1Oa1Dg8Ij
0AQQ0YQrCRopxvFlmK+Q6PYN2mG3TE9cDetgN0JWnPDv3Ub8zWPdevkF0hXn7x8TW+6PBJAma/UB
dest9l0RSPoyjNeSkboOAG/HtZYreUG70uL4qwgWqOisBTwYow5L9SQZ4stdpXMHuoX2wIB9irf2
OH2mUc3yUe/NOdLCvoW1Nfy+VuTFjNhNkbB/eyYJODQ55djEqrxLKJnWxma/g4WV6BSUY2x47EYn
3NbI4x6eFiXWprZxMhgjoVzAS6wHLOJBfuSfROx7gVYqjNIKVio+eiRtecGSCJcUUXBteiUp8xRo
pqLQ0dI0ogfmlsZ6aagfSYpuovciFk1QvBrcB28jyPbgWcGW734jRZPB+2Lc1exujWrJYeFyi71b
h1xXWVLfJuModM1HsziQhXOUp3RskKSODbzPCZHrpXDeL+dJHgfDhXqmSlgR9yo6GlTcQIKIAByf
6yRKkwBdqG/YW5dIT03oSmdo7kfASu39qZRy0ANc1ucXLauT78RUylB0fCJUMbbx07y5rfba4Kb4
/UZ0vq3ULYrCdtDFFRXyIbPvVwZRNpKBkJ4jdhq77xa2mPUSqz8HZu+ro0lpOpqUqm7WYyZ2UUX/
HMOTxgsA6szjlJGiP6u3u8aOUp7rfDLRAUViLkK3cWd++hEv8Z9hsxeDkmjvm4FwHQVWyfNpD9Fe
1UX5sp8tQdp5zrhv3TRxG5txyzkb34pyt2b9Aq+Qt5ciAF0UeeGFjTg3mp4gGOWDlbUE+EsaNdiP
r+Uqqz8UcYmmck7zuwvocW4ucjttAQU3rLEMFpCnJMx8ZR+FhZmguyjWPYM59KO9qC03mFalJLso
BxZgldwCIkisyRvoFuIEXChj4F+ExxZMPbXzIjrGwVdo8lVfA2Q8Xz0GONHHFXcMsP9l1NfLqLoP
45+/p6pEF9fommQpotLffyPnogqfARHiWiPD899/vUlK3m1BLjtI+8WzEz2PcRwVoMhM62LUOC/k
nC0BA5m+50RGIcL0v0FIzaZ2tByS8yY6wCQ3ttNOvWZ3HvgpkrNQYGh5PB5TGLX0xqL7WjhISdak
5OdWWxZjLQ2/he2IpnoYGmsKvSE802FT6QagEHNg4TAkgvwezvnTwHm4B3O7O59WpIsCRqZaJhS5
+8Ez1YNOaeeydGa2icdGOKgEa7Mq2j1BYsCil7pDANIf0+BwwLYd5ObdmHZDJQoInA7zMpVJT+Ok
wDoP8WagGiUfE4Wi+R/fm2LDqAUc3olmFAXQ4OBm0P8FI/Iwb1tf8PDZmacE7RWkmlKFx+pQHY3j
qRwKB8QDUYtPsChzv7z+InOeLliXX6mBnADJjIOqoiOHCt1YKorQL4Cm7wnRLZb4FMgAv4TV+xGP
+0EpSGbdr1MlcA7xnCg+nJS3MLtV2A9EDLdKe2hgCDsHHP3GZCBq+HhcWSr6AmbSg/PS2dfNTxU/
ZRadyb53F2IftMNidwAJ7+Bv4/6PYc4aPamK+cGLPGZ3EmxytnDUtjmxO8jQ0PjJRLg7M96jaxmS
/y7OWEltgKSmn3dWPBCwBiDpJLNIogwqurqPAB3GC+c64INi7uERqV6haIUOftOOpC8eCdLg4m3M
PTkxzPAGAUQa3w1go7v3SXGcvagfEX9+DvmSjrqLsec0bh/zoCa4F2j0EcTXeBpyA6EomYeDIEZz
tAZfk6AbdG731a/qUtRC/4GYyA2aMse3xxrw5dEctbW6AFNrrvDjHQdFuE8KIttOXvVzFWa7X/fK
reQfYydX3zj3+TlfqhDMQ8kUwEGbxoeHUYtvM5NWMaFh4Q/3ZYtyDm9nEvU1HppqQYRF23SptymG
Q3cePMkDRUg2QYzaGZb7pyOMqInGYys6Mm+tMeSkxcbLIxZS1MG1jFCqiXWgWPf0W02M5lp7RIwN
4s7da4XhJpzscnolkKjCb+J+dXt2HYxxAVdrZnyueqFr/kLmUqV5qVasIa3TUheoiNvO6NfKbSJg
tj+QAcahtV11p9Biom5mIinPxkrpW59k+gISk+u5nvYkTHLdsjPlgpgBnK618OxD9ItZsKJ03crx
dpguOUPmRmOs2DlXbvEM1IAEDtxMH85ppoegL6VP0pUeIQDNmvZ8g/GXA3MTd8a3W5GAU3ZjtejO
lye2mG9rBb/gKypdwI2YYHI3b2PIEb5S5FiWXhzJ9s94juroyEj3ZZs3b4LGXTVkqMpwI0/DhdSz
LvLoqDd7nD5eka1iGbRERGsOevvup5xmlvrwl1aEPGd0Hwx4yrLqeONnaejCAiryC/rtmkowRbwM
LxTi8I7sXJdyIBN+EA05XnHL7mgGNBqFv3A5Ultx1dylVbvuYM5j0GCdOS10qa2E49A4dsUzHguq
qNc1qVuO0ap32Kygu7frgpmCAV0uTx+NH0YPz/AUBY25Dqpk8r1k7dQKOKNcOAcb6N7xUT5SaM/Z
G76+4o1JbnQmJ5pC7kFS+ZbYcD4WtjDG9vmf+XLR8i6Oawy0rWRZ6wySg+Qk1xrsh5DzNRIqg63N
MOLy/h/9C4SGqJpFSZfRQiFqnCdQ1As5HxFXfdJ3Zc66awK3ibCBDu+cYBRMKcf3YxQm44b04lSC
nEBwH1BvVz4Zgopz39wCRCQp+sposViOMyeA5AkYHKBy3OXMGxufKW+w7Jjjgu1C/i7d9wdkfN7v
pdeIlAPtty6M8tJR5Hz/rn9fy4siXLp8PdQvD0CwqUPtQajQg37hR5Ah33RPSdXeb1b67/R/NOoO
LJ8tKMoPdDbp9sfneL7wBi3691AyTvNonE4ync7lH19ylprZggvXfn8oGYgGGb+1BKNcnKcVx9o5
k3EL77EVUKo1yOOYklyQPD7FwThcrMb1lVS40YcXAkpTSvvyM4ikDleVIoyGtnRqpSw4NZ7bdSzD
GjorG60ohaLYBWhGnR1b125ZC5lwUSwQU3J4fWn4QDAo70mZAiExBsIGnVXpCLtN2NpF+6LLsn87
ZnyV8cMU6hWhqUCD6HV6jsQpMj0VxrcxcUvUEsqe0yyU01pjDKgxYgqCjXhWTusxlQo4NqZwANWO
nmiVSqmXDNvlDWu+hBppwTb5UkvWSgGRFF1xU2mAIlu24Ua3JykAvmeiiPMEVVo379K5rhO1DKvG
yhUQ3puqiuhlfzXbn+RcwNvtJ/gp6VF9qXsLMqWKmjacOjSCpy6J97LaqMIMS0ouq9qcJLl5u/v8
FK9uFkQGexmM9P40w/xRydRpPedvzOHBavf72BwwJYer0t0/qBQcAXOwgMtL3+vnT+NXmlwV+rye
kMOZOU7Xwxv4CcKbIXofKlKV2qjJIBJbcawy813ee6M74aP6XAOZ6fk5ybv9T8etUTlfA5DtHVJa
BRq80tYnCJ0GsLI07QmAehMXHq05pxM0UPieXRu/udzJGTLpK++pLI1FbL3R7+H5DR4IfF3Abz7h
TMT9uxuv9CDO3zFxDLUQdUlTvZxK0yZ78WNXdGTHLsY8qubXC1t1zRfHOet19e+rJoU/dJkwPKaM
+lwgAneVWsMURngCLXC4M7QhAmoSzk4sQagEZ3UezW7OjhMwGsVQk8W7rcaUczwQ/KSErQfhE3W7
Kk4CZFudPoSfBm9L0kQEg+6aOKybr9Fa+TUGshuhPwUz0zI73q3svm8bIq0QfkL3p8Z1sQkniTlv
02K7C0bALTgyzv8DFvHp+TtemPubEzhY+VqU/L4lV4HR8NA1YsDYIgn3yGP3YRoCdgh03qWGKGiM
18UveVlqOoqsR4hV68HiVMWUzVPpqyb2vj2HLWmLnYZusk0SSWDUcXuXeqdvUrPk/VpYJj0lLzVA
r96TlvrOuLJEBHKivR1aAcsH3UTdHP/eHdPoEFcUiiULlFMI1LwOSd/3vz+dvLT7Xpgc0B2jntot
x2VpwYdgKQ3IfRwqGTMfNXU9OnM5Dqu0K+fPhZ4EJ9GJ3unJCwyUZKbXeooeAmMmIl+BEj/Hb3up
PWJFNBCNwlRSFuJkaQhhagzfwS29lS2IwabYPRGjWKG1yqzSepS06qpHYE6MsA3AWSixpqlNzzuN
0DKpWdx/T9NCd1WExAh0wjmLeyJ9+GsBfDg4nhRkOvVMsgIt3/8G4TItrzO9vBvRC9EVUXolFuFC
ALj5wcLNw585PcLn7DrH9VFjXL1m20SwnPqyhVIYPxQPHdgRUrQYvs/051ICcTTCcQqc2Ocv9/jl
R65Ixg1EsEt7/FoRPQMQ2MLMaOeVXISkLTW1jG7szLddOsUjRhCU7bHEsmbZOhPhBep/w3yVRs7C
xdjU5v7krbHzCk9uTIc7kUZqxQQa8yzB3SD8GWXn0jX3iS/hYMwaFm0NFnmq+mceGzWB19mpmIjL
YbCTKSN91ptP/ZiQOar4IStJs7g6qw5uKSOCGRfknpidlhnmasHDl4fov6uBH/83rN+53s28tjsO
tAFtHwCjWtQ5LGdmTPNuC7zdA0tmFvTBg3M1BGr8hZe5Ktwm7hLRr91cMWWcCGPqR/3R2HtT+Cvp
f7FXQj3EnBv40yuV6qkWopMSOTQB/qflhdmfjzDxgH7xm2XW5z4VA9oFrvPiVdEhx0wqeQqGBQhV
x6rUbSWv99pEyCchfN1PBhGMFKGMZnVaUtAg9jTUfUgc+3AibasuVnKmishiiqhUPkD40a2Rg9b3
OhYkw8QcYO8XZOdcTxtrL3WQdfg5ssX3B8GrSGRFP/sVq891Jt06350LtxdgvOy3lSHu6rHovrH0
TGaG6iTjfECGf0bj8566TZLOEb70KLOVo0MQduOn5Igx8h634QmAqk10XVqlBcYISsFrrLF93z71
b/kBESBDCr4H88gwNhyfdmu+Bgx/ISO5sHhyvdTmf2uuar/3yfPXyxLQUMkW/TEGOGnbYzk+TVYV
Q+GJw4IaGgiRgae716u8dDRV5sC2X5Z3+P2gFt1IFLWAHi1OfwUvnGfx8nA4XFhvP3Za7eUrZj89
xhDbZgoo5iMpX6ela/GO6aWReBYZ2ou53qitg4HsLdlVyCIylZYZlQES4U6+mXYbn42OONPZW/Uh
Yh1eAcwjvW2HBG6XQ1bpSCarg9RtiYB01JlXIctEENVCuUH6UnaTzjJ1BIGw5XTB2JiMJt1ebfmZ
W66dccE3x5Yo0nriupIDp4rqtRsAkdXAUA7hzECeScklKsNbkwYyGk0WlursIyZXvNK+nNBjatsW
YyakxgULC1ky1gnH8LGxXn1xmv2XVx/sRXVr5C4f+ijZVsVkcjHYQKc/37CMI3FywpcV1chi90xK
mtgN61Ele53LRGJ4go07RGhyOefOtUNivvjeKPevCko/jc/C7zG5TZNFmPkoI7w79Z0vJYyVuzgz
Ktge1tfoNkBBV5pMATt2yf8WKo4ziKTOxwOKiKZjhYilDtlZuBvimrXlM2l1HpeKZYsyscoiMc6j
Y6XPW4PHayl9yVFVvTSH+OMTlchOhMPfq0HoyoC76gwZbL+6mAO8zDkOyHqV8QpzzyxNBQcLDbhA
UgBIU8DoTPOnwqad0x/lCUy9XAeYGMLOK2RaOiO/YdUWideE0WoOdiRn8KB6e+tLIWwWdxH4muz4
CKFTgXauo43zzgs6HSMvQgvasiJofqyPhsohPuhKGpfpBDQVEDQ6RHrWK1oiZliiGVQOrbNuzLOe
NpL5yTmST0i8jOH035/IZGyBTVeXx6SYR5ZLBQwv1/KRiHNTtzcwrDk7DRNx9bWzWK8nVmO6uMDk
yAYnq1RWpdVejLr0StcSTlEwJDIkBexfQeRSjHUo8fIDFzlOajjFGxw2NixbxPJonWhYxKELIR3k
u5FTvAQTadQ5SMH/WYBKJQsfVXot1C/C7QEq4pQ9y6MwoquUDh3Zv8t0UsZanxq5eDNO5ywHIKho
jR8tvNT58dlFmxVXnjk4SKrSH/ZxrWBq5EAFC35CURzzLBuISM/gdulI4WEDwQNLxXeF7lQ6FPaB
mjGG/6a2sgBVyCWyO3WMkEEmqVBPXhxeqkOBHzFASKc88R7VcFUaRpKjjE16OvkIyN9J8L8Sy38B
ju5KGRhZHHaivhVFRzLQ1PrqQp3uyuI1E7W2iXST7fIqmfiS8rlPoelz4h7IFIfA9/ayoZEgbnzr
wbRvgKfU/P+bRDmLXkt2nY/l1TR6mozuTLvNa5PwMuDiTABFNi3iJzffDMePmA/T46wPLrhm9gFe
ShiO3cH32rTTRyxB3JYkakIOgldg3JJtrvnqHMjMlgtxvekuF/xt8dUSSebi7MIS+em+26ytSTF9
Jq3YuX2CaIZ0h1AmqJhASHEldTzePXONbHkkEUOk/G9kvUUDWcfuaKuQHCr4Ca1Abb3rNUCpw4tk
wB+oaDvAPkAeAI3E9I1XMY0TmqQde1Jk6P2ch7mlYshW8HhW7IWhZKO81Y5EWIj0ai80IjBi3oLK
4x2x+Ac5h96jcnG0lJ6e9WacI0s6xYrlnR4ETVYclbaQh29w5f6Hfmqe1GXVFeDok/He6WLRXUbg
j+sQhtPDE5TShSzT3nmPA4v1gYHG9ffR3bNBpXART2HqMf1C0raOrHVKGrHZFG1f1QdBSGqJ/qyJ
hOZnkyR5RJqlVFsMC7cq1vTopExzqQvJB8j8vAX6Z2V3YHpkudZ0/NAqBWPcOg4WsPULW8eHurBx
/CUGbTKGflZCK4IXvAN32IKvVEoig7ig4R5LgKT9Jr67cD2BwWFkL+la85UJaOrumNd5eMbLPw6p
utqYglvJP2VK1Q6ifpZIJBa3f99biLN3X3qXSh6Kpj/Q5tIwwmIhlMPT8GhYzE1C4LhVR+KF9BQ5
DfWNI5pPRtmtekkPq84JOShRXZjnB3e8uaiSzGKl93rpi/zXlIde+Q3IcUJEiK3DU3CdXwRJF0E4
GaHPlyfQxZyjiJvWdCkaoBRAaXGzauvVpWbPZSEqrJGKcLr////ZB8N93pscXdxKSZHJq20nfvcd
+FdqGg3CaxJxigRgjQfAb72YtL97RwqsE/KXY/itGR8u2kmQHYRMy0bYeysXPUzqhgvy8n2Efqnm
T3pa5UK4EfIyejjd6PaXcbZAJ/lk5Vb5uwvgk0LHXOHPvK/QGONBteVFpDVNxxJnn5HlZyJdeKhO
rpoH/a1kCeIJwpIlCirmQlBhrqg9MMi1OsFyos9y+426Greh9LDTR/wv2PKcfRXuJuqKLO6gYEF4
/j0cb4FLaeouuIx8ay0WAlxdRZG6ZErDpiQeohzIzKbLa6q3+TPFM/k1ShwrclivUDv2432rP7wL
z18hgLUp6jYKrlNjND80Z9KrjHVcIUDIaC8y+D008d5vPEIircZhJxkecpRVwbQ43/M7C5Vf9fKL
pCX0oGRyTQ7VHm05+DL5qsEOqWlca0MSGieCcIxpxvMTrFCBLz7L4XCc8iETB5mxjDEc5RNdCPHr
UUBTIDYajij7/ocrYYS4UJJfBKLehnPdukAENJDqZrk4409mIYHH7LyKN0LJMTHcGtZnu/cklFe0
Q6mchdxajlGjBAUCbLNWlgs8Xrkzl2QIhKN1+NdudDpn0cVEMCn19Z4ib6ypnZOCYcHOzVrMxlkA
C014TdThWgt8e1Guk1IlFzFrLYOibz1KsYKrlHfNwLjoyr/PCnxpqlhUiyRVlbq8KaP1XD8D95KE
0S0Vo2UVOthPLb3+25lLNb1WfYJFMXeJf86ZKsSV3efVNwXwnbdaksP0PHNPPRWOi+iU19rWexGL
mr1deTBEKOZsqBcxxiS1n/vQc49e21eO+VR6PClk65jplVGZkBIuTQsdEU5acLzvLgxHhjmgxuY4
kNqpA+fUPFAjCp9cxc13eR2g5eKmsZyjs8Chjg+zNkpMoMid92UWBKE+3KVzFSjigPJBM0deQ8xR
gaWUuPjcIFGSPsd8K876Im0RxeC0EMFwyGGXbm85BqkaoBbTCtK/mF39SjJS15zUUSDAmJOjk2jH
MBtmkeVlq50wedGmepbLa1e/N+Mjy5USQjcRCVUSEwNRIMRhHBk/24d+9huJm1MemZXti6FSakjD
5hX+yu6j8oJdeMNrXraNjhjGxOUBu2tWlXwdM829V8G703tzJDrhWtyKoqwKsZXuSPcJ2kGzK9G1
i32cg4PG4gBw2p+2eolR1G+p5i6Hi5NHtJr0aovyITSIG5/vqG4L9R5I56DZJrFqHnKLUQXG79O3
WagQGDKwPwyUFzYT7N9dPqSqLcPqxX7Dhfz4mES/JNWTZ2/G7HuYyInH8E5HD5hP5wq8SLyE8ulF
K3PBFYqFum2DXyMOCO32cK3C2qJUVgqH5rAPPKEN5XxLbylTFyGfsCt0o8azN+4PnpNHfOf841Nl
wQA4pQ25YmZV0gic8oLAlz0tafzro5goC9G0B09wK/yYH2WE3a4EJ5q5aV4vcjv0XICgTD+GkAZJ
6Mr1goRFCmnDm3/o6YtSb7kOZoGvTl+VIyIOpGwQpyLFK7EmHQZEhlp2fU5trPl0XRVo5l1pXmMM
AiPxftYjnVhfQAILXCBWJFArcQo/fYBX9/o1IhFRyow2jUJw1g8dg4GzFT7gqyWAVmYZbTLySRU/
peV1tAuiTrjJNwNNeKncSFQr+KDg1XbWXCY0yMZYNnei89ei6Ymq3TqEkw/pSTlNp69nRMgO2bLf
glGNqxXP+SMIN0BT0vrJq3xjn8QgpEAzBqKU8rhzW+GPgShQSqidyiFtE43IHUM2ftlr7QZSBTfS
6BhZ5JJ89cWuBPYuELh2sSqzDf51z3T5z09aQOY5yjlk6nPfeCFRyqBr1c/snik5XIlNupsPqMwS
TB3I//0mMtMsBmOcKyDeKyK8Crh/acQv4tJZMSyyg25F4ASQniQYZsOdtQA0zgYCNNrxXYy/CDzR
tA2u2Vc9hzIpod3itVgFZ8GPHrjx28HbpopRBlJs7FshkN65svVZZmyIVB12oZEVQtWmSssPnJLR
ddVxtFdLw8uIxpXO/1F5MZHBORTdMOSzVmeZsUBmsWrrDL4uTq4tZnQDRHH+xv3RyQiewb99jpNR
cMsM7Xctp18i3SRjMubzO/2SN1pTSeTFsCgdBGcaBsVePEh80wXUAfYPmHD9l3zyhtpgGxc8miN6
LrnaV4R2kTfDdOW4g+RQe9W9XLMPEYJ+Ji3n4+NrbXirMp/iVaE7cBmteS+IidJ2ScLhcZisMfAh
F0fAAqJfRbP6MEKxso+KtESXRbQgF02Y+kbNd/0XTTMTKpc/r7ROB8P9uRMhEAnJ6i45SfjMuDOe
uHJUJzMlrl/JUVpVA+SR2rAzZV/6UB+LlW/WlwHhmQaqTbK90wpSnej4Y7Kk9it6QZR6kJeaCXcF
s10SX7q+PfvfrRPpBWdnF2yRAec4LY/XbTP9+t9HtrWWLQ4BhevdYb81OBNXtPKGCI9jLChmCVuL
E1M54gqbSlK6vdTdw9kJLBiQkX/k64EmeruLOtdUhdc5LcO+FUx/f5RKp0jSjIhNMIfAdIwGFAVm
xa6HxETilAt/bV3jhMi967gGhfnNmGONaHm3RbbZBLVWEdn94NgqrOrKv9kvjLXhZf1KDMbGbJ/b
tSeJ9ey6roMeBoTJEB9EwX2Cuvv/h2KNYjolBBYx+8NxUAT8L3/NrMUsKjYaT6ahhn310vyKHoAY
IXWo/qvVl5fzkUFjl/XZAxmpeWn4RwPC+hqIqgsqXH6Quuc4J54BZ4Rg0/SztmdVQM1UwVmmjpLe
f+F2RL897M6+kjVqO6XVV790kDkpqwsOV7uqr7wDfi4puJ7BuaGDMvKi9cyuhaG7w95yk90IwnfW
6OUWwDTEgEjOnZDo++hjK7gHwk6kTIA+O4L3oKDGSozr70cobjGqC6dT+L1OAFchLSPNO7g7y9bc
2su+d/WmIA4Bk8bC4XVIKtyOT7fWaQks9nCfa3dIscrzE2QutogihnOx8WxS/6RHXrnhG/tb0Qqf
h71a9eY1XZRPj+SHsaxWUhGNz2MDpkC1GaffCJVZspCej9UkodI3IvVwoK5vkiDDyzTu4ZWCkZfK
/7/muCnNLi6g/Mor602qxOt7WmNm4G+9mhv4G7kTaVwQJUUopPh50ZropnkZVNYfmpAlvLqii7lN
MTBSop+Uaf6c57mKe89/6pMwjlFkVFR0RHW9PygScH9AREGmmGMCv18lA8mFUDPOs56QSgp3lXoX
TGp8bb+v9aPym5S/goFPN+HYa9c4GINAIFct+al5xTCM1iegyVwnAAiyY7n1YTkPfbD/fGl503Ie
uokWW2LZNfOe1caNMO69ErgGfcpcBpU7LDsbtmVNkB2VCLTitKOBx8zCQkiZJRRRTa36Yv6ONp27
64gw/GFsH0STJW0qaMYDThlzGTL/RY8l17MrAYhYAYobBvwxwyob3ld5HoJCP2E+IDi2G1urAvp2
hEcjyqEDaB4Q8UDoao0zUVIQaKHWD020xpqn18OziCPK8O2wkLb0UgG6MktrZ1RKRSn6WPuzQ1E3
gJTF4zUsrIwji9/Tn6UN6MLdSoLS02oaQ+uRIfwKfmE1TvlwZJq7Tl1O+KFIy89XWv/QdWE9VOm5
4FoXN4So32o2PvJ/NFvQ33bNgFqgex755CERAR5kaNuRBrUTdyDtvTUhPlzWNZMtvzQ7c3FPaimG
cgUEr3DJJs5Tb2vtsxZqTchZVciIcvWEuncNDZPJU2LZGD9oZ2TY4jBnC6CZipX/rKJRd+ONXSVD
JEtDEqH1ZlhAwRHfiNKrpNZC1lZIhnBbvJu0KmQ6z8+6cFDRrEyV1Vhdg4Tgor4lpyt+yRn6M/Pl
/RSV4orWCDIDpZEJk6wigF1bYiTiVbsL+VY2XCE/F4KS5LL2Wtlruh3mVoVPQcrnlecdg02KlSfm
vOmklD3fEzCmX6/ax5T+1LUS3IFwvyZPZqjI8Luuh1O33Ea+CU3BS6N0wFZYT8LLjioFIwB2V5Fp
BbR6fWrinmKvl3whXdZSmxCnfUwv65kbfAC/kGcGMNuU+dJoCvxwcJGk55LGemlzYdtKlP5b8hL1
z8dx8KXjvNuQjMRQTqVamtqOobVXRJY7vy4VTBsHjC+SMtlSXUfsQLYb3bq9Z6Z+5RsfjzgbGa8S
NUbAaVKld8rBVBpporlAnmP0z3kxHfCKslM7rPvWN3RbOg3pXEti6laZK2HlEKc9l4sTMc8TW9wL
Vetel1KtzN+BO37bTdpVWgA42HXxDgtO4bD2S/gCeQ6uVFddTiRRb13p+fQ3hlTJYs+sljnvtJT0
KKFXhTfdSX2Y3VnTq2feVE6Vdb3FN50L2C/iPfPNTAKKd5FKYiQ+AIw9mDElDdObnmx2blbaMS9U
UA31gUjvpSzWFGtDlxGuVODSVls0R8jynXh04OrsLVgC5iXvcD6JBUC3sTXNAj5p7byRk7xvF9uj
xevXDSSkkF+laIkRWJ/Bu9+RkP3x8DyjV5DWmcZUMA3kHYOo6Uxl3DAxHqgu+wm+RbfVOWCUlGW3
32HSImGW7pW76hzF369hegAw2ntYKBFm6Do+hhqwvRDTx87AggvJEbXBoVsLbTAOvobVRfXFmHeR
ifG4wzubtwKwIS/5u8DQfWZEn6Ce7vZ7RbR3E2hCURkZi2YJbWitdSIt+SxDcO0ynxP7LdczyZmv
bZv0p6VVmyTBYyy4PI23DHGKxTq4pAVCXjW+cdb7ye0wXnQDIrJRKnL43h1F2YEhlPk5x2rGsl1S
UvcYjrBCb8Uun89PPbdU7RMOlYxCER2FBrdVIKCBclfimVzkQScTVyOTz66avzt5GtcL8J3ZmV4e
cEUzipPJZv6ckkXKqInSU04qZCn4TPy+cWEzF4sUtK5vOxg0gP/Ob0z9m27QdSFy3caCGghPGsCo
H1cyUk95IPhEsg92uat2d2bnyPIW7xxYK0AhvWClWbRbRoiOXJ9RJL9dVxREYsop2BQM6zRSYG1E
SrjV21vZUaLIUIzQrg/iql2Tp6z7dMIJqNbVDcIizbkVm+SlaoMJcP0oLGp4EFRmvcAqVoVCkZlr
Orb2YUdo3ngwYbGxso0IVPDtq4oAwz9qhw/eMl4D34ka/o5TDubfe8pYWRJJ/b0St9h+zsN8bUH1
Q4HiSFuIHcmrWTPzLJWMfGgTTcycmr+uA/mSufQ1btTgZdb6qUZJcDw5V2EKxR/FbwRPSFozXjQ4
miNL3/NTkGpMX6ILjCb85kxA+0lXfH8FdGo7MjFv+LYJFJ+F3G5l6WbNkarwB8eGJiThMOxiTc4m
4Koili7axWDlWIylH6hJeNHZe5v1EwNVVlzNzATJYf8kD80PdUdXEhBceYO4qjU2xe+klo+O0f4c
a5cXsyvKUu7Qt2hpDScSgnu5ArHpigXPAKdkQgVQWeS8u9rHSIuBYFqR1e19jerMFaHpmSzWfkIt
wF4pQeEZr4BA3l2SLaO5a06n9j884VAFBvxHKaWmia5BjFUc+NH3MKVqh/sCqu/ub/BJp3Gfk265
+/V6yoMMS4tsBvI/kGGlqWOPM07luyLjLEKIurlYRD3RBQEUCclsG7dJnwKULp7094RC9SX/Vq+I
aVGv4UqgR3EBbHh2ErWJ48lAWzRY58bjwRnUdlb6dvqtJQ2BIcrHkqYXv8fWvGVsOZIwrjS9Qcl8
J5sqzz/3Lzye1TgxO1fSBm4brjGEq15NyYSFX5uEft0Fi3kymf+kXAH1+MoYCEjJsW+WkWeBlPvu
BXt+/W1Kg0aN+JSk7XLjwvco3142C0KYoanjF8cmi5kDp8vldyk6iroEwCLghm17z3n3kH1rIqlw
AhK0dVz1nvBEci6I/gxBtpozXrATNSByiLCV6V08jfrmNoUN9hIY7xEqXNaViNADHogIHNnDNpRj
eMhDYYXT8vOY6J2Z345VpjqkNoR7x1xmEwl/KTwpGttczsX9+Om+xhVebDkteQwxpOsunvnwZLBY
fdsytRDvXWsQ84HFz6pVDl5HkZHsCFjEj0Y+E1BZ2isz6M3dInhiUjUk7mVtSwenkKlOe7T2mrkv
uQ+n9xqXzHUWsvjT8jM3fBrrLiAfYvNWdYTRb0wN78dZUWVS2mFwUTofTQd1MgNZnqvC85fm8YpZ
TyHXOv70F0hPv48aP/PrTeL6nlyN/RqaHhAmm7n7ihD/rlUj28aol3/bYakBFDw5vgExgTWbZ6bT
NfmO8YCQymOLrsYCCymiUc7WwFriH7U83zzxL/CT5Lpl3C5tW4GnHhctn4Q5V49x48Pf7VEDpCgV
zmGUw15DwJrq1XMqw13NZbAjoHjvoZHGA+TtAkZ6MA76SXkxMk+Ihj2oZIDrcMud1UJKJxk3zDRS
bGd9am+XHXU9L6LMxDwhkUXJDkJbfllqnPsgxYUyzmLElryLa1sUhw0gZozOv9KLG74YX3rJHDqd
+olswJVvE1URt16cxM1F+KA3feTzQqgb39EObaVbc4oDKgh754fiuefUFNJzBXRVEyIHf+rZI/wQ
yHemIOzIkgstV+BMXbdaqxyEMZS7R6eIIhGS5I73ZOQ8/MA26YeMNmhiDdO/2zUGfaHqv19Ygqii
C9ChqGyP1v9YSrvHJtNfcgAoO1HXYh8j55rsJBcFp/ENoyWsL5dEE4n/95G4H/hPF2o0p1lYvSFj
yRYCyVGZP7jH6ZU4vIzBLdNke2VJVyp3h1hRbB2iGB5PCEbLAI4k/Ei5wStrHBVA7jvnkERkc8Nc
GUU5lkR3mHUfHjh8OyZhUBNfX6uhjgy6CW5cDxNJIj+9R+ybVbp+CPjvC57Z4Bpiv3+ZJFpg+Zkk
xz2vpSYmrE0n9FL8xgx7eiC0uOMqjQvy6a0KZNvHRbsFZJ4D+Z10tjJ2T2Zot9Y1JqBGfNaPui3R
yRXvdmxXINbCkPe/Gt5a3SpnnYPzEM9P30ZBHf/+O2x4eNQkluM2oIqeknPJY492P7A8BOPZEVjP
hTEevZmss5zDmIuOryHPC1CNUvmiC3nEMVx3WEw0QUNhUr/Qw48wa/kc2UGlZ7T7BFrO0e14Op+f
y8IO55lDon/ysC4u6vDvcT+lLDnPFJ4JHzYf97/3k9SFQXnJXyWlAlf8YVzNk7cGW3mV1A2f0r2D
603RIV7KG9gEM14uaSV3HqJY0Z5r/glODl3rDfdws3RG54JBR7bMSnGYkCvFU4yWBf6SQw1gHO72
zbjiAv5Vtpr+n6Xvx336vyEi/53UjeQrjofiegO/9emNZhABPjh+/3dFpqUXxDLQTmN2EPzkhx2e
KhiC5olSr2DRti9x/cwaQiLUg4kToua9zOvuGmiXksNUg23kzKMAJ3LpIsOP9xE8mw+KELnxXyjB
1QSyg6MBegJF0BCEZx7whzXyuTMPn9je0MhOGYzULvB8TnIHzzNwCV1mvrVU1P7ReD5WLy9XOaQW
HpSaBxnaMag0ocWl2IV9iO/rRtoi1/gE9e9g1MA+k7SBWq4tCJR9KpdsMwAemyREb0I9QHsNbawo
0f3sJgZkpwaRsElx71ICdrCyEXZioXusmmAqdu0W3Z08AXtgn2TFx2VDvD9ZXMt0dsxqCqF9Nfq+
LZzXob+KikQSXL1yKmXMnrYmDaGwdHnXaoL/WhCi+88l4vuNju5XG5ka+/C5lS2tGGRujyJ3m02P
/NmUeFSmiabColEAqHAAxhXSoc+e0VQyflt6xZXRs9UfO7W3zVjL2FYWFShKO65/ir52zvQplJs2
Dl9oDUeCeTbbSLdelh9qnVtZ4rD+o7E1+MSYiDTW55GS24qlmM8TzkCjd9t3sFiZN+5qCuY1PdkM
t9auiBw0R+W2dIbXa0CnwmkUHo0x/WRUGQJ8KM8hpMBKBl/OfjQ2H1T0uBD5hq8FMBA5pYJRLnIw
hPzZ5BPi3IDdVEOn91tbz+dktSKcfUePsG0Xl4AqW6DhXHrPY0DL8+KgIlUHQtA1x/qyFsw0Jy5P
bV2VzircaNp5W/KQn317nUfpyBTzyPiqllYFc9LfuyqQsndJ8Dh+NvfiKWyQ4xT9747+GPKP8EPr
FRGWIYUpsjCu1eRe2B2yID078FLHq7bqQeQaQOiYWPWQpj1RPeErvMOETTYuZbl2NFLxz+4JizbB
26lLdEYLqBiaZHWcuU/IzcU3dS4QTv7Kiq95i4hYW4bscQF52qyuDihufVCaaBwzGZ+evtX8n1Q1
x3Yx8jFKS19aX94NY4bVDV2S8DCITodmHY8Fy6cDCvni8M4+58VIvKqSc8wzkuUrao6wFvwXjofS
AScfYIEoF5Q+MpL6f3wLuOMRbFmiIF5eqJQnSd+MpLxgDfpTFb6MjZ1MAEfZjqjtjIooYgN4gTC+
7IPL/+acl7RnsT3BWm9fEwuruO4wRim+XcbRM57PnEY54m0NpsnICANkFPhu5M7wmPbdzoq8h1wk
H07dpuRDKKlHqD+0/gWDYzcEJj9zyM7FZpYUB2LAEl7W5QdOLhRGKXdfCCviQ0VVo96cir5LwDzk
ia0jEYKzHbwVHjQvZHWeA5DRm6iExKlToKH8dCtse9835m60f0FBu57NA0EF+/MGnVOhwKEwO54Y
HLPDQmbyuZrZSd6mH3iGQXODquKrOY3gkZBWNsUzgi7shdT9xzV9l7lrFF5pU4HjCi+f4LixPNmc
CXr1uxr1QtoUXDmGP+cfwGHlWz6i2EbyIv9q6w1iKQ0pQqD0GHH1Tu3ORtvwAAur+C7HA4QQskBS
vtOVFJTO7zdNbckyuRA81jrXYPCb8l0Utc4x91kdFyl58Fs95tDlByYnGIQhz5cvqvkUVybgmLZy
foYpNHjNehTSlRfhqDqHJsoOEmO7nl44C5ZnNXwGqpfXEQ3+gUsQMRLu7Xl16SaCShaB52H3FQqr
IMZKyVuTmyB3w4o+SjK8wVdzkAEeyuuvoVDC+x+FQePJ10GRRWIcohoLVVftDjrcalMNL2ZqqP+M
Jgw9tzA6dzAqYT7mYkY0uG0dku+IdZpSV0NCSH6eWMd7lfHz8SsI8sUrYLP9H8nDIMTVng9hppUh
pTgKNEbOc9tl3qzi9mAhiq5fXKyR5IyDlZO7jR6PZc8Ut/LofNBt/5Ku5AkdC1ivN2dLpUcn2Wf/
SR7BgX4l/JoCWuFeoKQhKRs5+yj9LV9qHij/4yCK3uENV2jzI5igKNJf0Lr0Dvtf5hZspfPCVX3Z
QL/gGDpZsPswTiRbd6ZpvkpO/zrSktYnP+tvz5gJHK7G8+Tmv7k+4x9wqMgx8ZIJzfZRXu1HTKOS
FfM4vpIQD0SCmiIfkZ4pyOrQ9PxGDg7mPbNNImUjL+UPV6/g6RaNKRLVZXXZ4bg2jPNAd7mih8iG
WfE0NtcU6H3+efphe3IkqrjKiJepI0yJbI5LVrDHi11olfpjGhTx2IFnfnOrrtuJP0YvFqxvtZrp
FNmBVBmoN7SF7z6WI1SLCigj4TechUf9Qgr1nEkXwzpoL8BO2078tUOkuZNcJ7N5FRmQrwMAPYve
w2/Fli3/vhdqZswCdg0WtfGrLi8u/n7byaSNcjVX3JHVZRsO3eZ2GL7wrNPOgT/TQoTxSPnwUU12
dedi98Jgo1hrlR2oOzWJXI6b06ZzV5pK6ZCI2KTKMgwHDKfSxVw+bCYbh5i79URCzagOWG++OrAD
rHEp2XqbJak9NVy4SvbSlmz6ctIMO+VKknQI29UZiNo/+Q8vlsZdgh5m0VHWA+Rj8w050cdtwQgW
B4IgBoLFGuqyYMZboAcTeQUeI+/00MUmIF5ZFQYwy8j3scp2GsCqF+DAhPKyC9uAtwwSiujAuwYU
xzN6xePbD4ScRHoOf/J94vhGVGFDt3MKnAZ+abigiR9CoitWILD4fAa1olMGGyXOoN2r1PBTuqtv
bwBjpcpXpfv+YJ7VpXGq76iJiW6YvLXWPkxyrPbq1sX5CDaXVH50FUeheFSjPrw/HJ+i99rPjfhH
MxURBA8BklCgThyxssxWolHUdLCkDsvNwJ7XfAP3IrivKGnHA39ibNPrwcRvDBJZq7LFyVzVJc26
xnzPx/qFcFWAAUwbqhm9ZrO62T44wYso3yX2wTI7BY1vwSyI1F1QYURojHi46cof/LjODYckgFiJ
KZ/Pi1FOv4WQzAOl1rSR3vz477bTplXxLZDUcLiN7sPPg0lTIy/ZMrS6Bw8yBTv8mTwVeMxzrKBf
EEplaLpzK4NQPrynMw0+hRhAjc/SxDYRHmjPMU6jOjNoBy5xLSn+TpF/AaAmZ2cGiEiBek9KQN3C
6eaNOb51I9q3xwpQjGDUDy0mET25zLlOQZ7RSxWMHfQ55o53XvJjKU4QEfHlM49QrLTKgu3RznAI
C+jSmGKt6Sk60DI8i3Py+ZXSEvlnFZ4fyESoBYfewqEff8IMRahT4X8wEEh6dFVNb8uW1d2iOIeJ
skV5KaHGFCLiCvflhaySGA69M/1Pz2/zI68gfxIKjUfWiD2Vw9g4bhV/XOojBOuzcDgnOiwh6/Pd
gYrl6kKjtEaGZ97NeBXTzHN163ch25i85wPeNHGQokl9+PIHVOAcABDiOjtIOYoY8gYVdW8Kjh1o
zqwarA5s2aUndi0e3uXqYcq5bYJp5j6ZYkR6GtjM8Va9pH+4263AsR++RyZ6dOslYz3p8p63FiMn
URgTqIjGpOlgITeaUbgJbMsZn1TQ7foZdVjUXaMwlGjbeTdWn94OfImt/6xcMqIDWoB46oGtQNzb
wR4OZFn4zjxXB4+C7cuK4b/ewPA7zWjM42iW2QhnT2wxZVgcC7Lse2b4aKV/Qlezm0Y+9a/33zln
c4sS3kiCUw0Kl3WybXCBL4jgCF/mgyYrsfLxgXQ32gzLnbMQmZD2mdTLdl/pbrKKlMAJDDBbAiQn
3H8jSe1REDwG1eRtAyMmoCijAoi6WoTnhz79VHGumBtG22ezJhD4WAK/8miPU90nR/1aP9KmaV7n
HW4dCUSyC2zPzPffzHWapw+cda6OoIMIkZK6C3yjY7O90LeHnUhgUw1YN9YxIZDcYIxPo6w6hmMW
jylJ53omA0g5n1USLRlI/uvcjlVAkLdhx0UB1AjbrbQ7iYeTcr1sQvC3N/3JPLwfBVsnmhPF6+kS
pBou6z/H4Il/tvqoA3a/6o/ULVDdGv75G1ai2M967ZjOZrURHCLnqHQAjg0Yd9zyZWxnurcl1ciO
IpHDmsvaXpanTUfRM4vfqt+32pg74knapVhIhe8SDvrnPIdM2Utv8KWjL1l2aCHfbc290euWB3vv
w/L3Y9SYzcvpE8G3mWFKwsNnU0dfovVsiByagTfH1laenyiYrw6LXKdR+P+pOIMocLZ70mO/yOe5
hR03xLiYOMjvMTAP7+cEIVQIC44AuGq54M9Zb1V9IGh7c0sG/c1TLkAOHqqQhwD5a7XZ0Ds9N6IG
vygaNheoDDzDNVoi1g2mj2itfGOYANdY1pnotFb6DbBNs1mKJSRw2vw4A9vJ+vGkMatGGf1jbTKR
lybV1i7Y7bGAQIaAfpaEA1ehQksjyyacYsZjRYZqdrvwQaU87dZjzvad3Mv01tGdsSFoUJniiDik
BgCTxti0lzevl8XCxN4yMSoh0RaXw3lvIa2375wpupQmf4KQrBLD0mEcuHJZpbvIupoo9RThc0xm
89KWkddkCD9UNuTlPkTh06Wk/pgXZVI9vFPe0WcHJ1KMkSq3Ati4n+qvVl2ypy/e37QvBx+B+KS7
vUDZXqiFnNTb1t7Jd8XCQ+9V750ypa1oFpTD2ue9YPn4I7ZCW7AkYdbmpYpbCJQPW+LNfP5ibwyr
cUyasdL7Pbiwo3z94VP9oY2W9yGPmbg+gujwZn+1WUiCc/4EzvXQJSDYI1igokrpAYUJQiM9ZfAH
eS+ZfKf5IslnzAV3b45XXQMVXsFIdaiojok5rXrYNA2Gixawk+hJtu72sY6bZ4XegmG3UKqtFa6j
7tYr01pVCxh3aSF3NC1e0+FmwhYuIgWcANX6QVmy/4SPoU4TKZcn1t/DdjuCEm+I9MOwG5CflEzc
oCfoWAp78M/Qz9wOMchjlZZ6EJYzQ4VtfGwSep/ysIdZooKVgtQSt9EAWtxft3vPkGSMpY0Cb+wC
CgqDk7qHsRVjybyFxI2RF5rqYrxNfwwJlYJyLKZfaU3p9PuFmLLljRDLV9fHuWSb7RzbUYbv7B3E
6BnIlJZ1aL6nxqhD5Imn1hJ9rnyqjFtnDGpKqYrceP1+JhbxjCCLfQibiVOAD7zULwYXUIfWBLcq
QqOhZdmCbUG9nV9xvml4eROUkz9BcvJKthvDVGcGecjxFJZuQKCPDAVfdrmaO8xF2Y3jUnbfHwK/
u0Upp8nVri1vOsC30VGkw2ojoQXzhepIGVxxqcsHtalE+9DnvBGo4SpS47JDpXtyRicAQT8z+yYO
qnYq89ZBRnLPAeNsD/7DFtYwEHLLpbvDPSneVoEo1BVGEZqBRGEr7suqyC0/3BdymKWkSiXx0Lm4
GeY30kIB0P5UqltVKqZ8ZqAPWpEpg40xvO9bBb4RDEh+OBYYPQhaYv/iUuuQ/ciAk8y9Lp8CIqyL
93eXcwrVLMlv71skggyrhr6ThHbrH+hH5oionbrmOBAQy3sAvvJUVPpNNlD4UsT7WKGu725nndF+
hhE1UZ8s7FpBK5oo2kfVjOkmvkk9J3eCsIHaS1J1NBSFZt3Fj+a7zfpfTaVm5Biopo13SqXIzBZ3
HeOk4FucrnQ+OQgVFPAHoe9f0FK3TEHXyMn3ikxGYXxBpS04kv39VDzxu8YsWmBYMmOt7Igr4iD7
tzA+EfvztUr+LhWCYbfi97F5fwfoj89XFBLvafJ20XQAs+L7l0Xzt1P3YOMBptEmzTY2lldeN8GG
Ofm2gDCE8l/GjPERCPWvvxyaTkyUMHERIXkImwBOXufasla05WfhaC3dYZiSLFSQA4ODcF02sFc2
qe+aPchfeRUdQL7B/wyG4JsE+RT45jqjFsJRGuQGI21OAPKms9KkF/UszPcswmuEvwu0ugFXk9yR
/o7X9Dgs/k0zUIyOM2vg2JxdYgmJ5JpaCznS5rj5suQA0NC9swZOdNPsQi4K/ffHhPu3t4Z+Wy/H
Dyb6bw5DuLDdzUNtB5EU00sKZHm7ZTl2tKaQymq5gClAeOk2S7ORqDfcnfSXlPeNBon1rToIkHRv
TLhrR76aZiKh1dVJYDiLnv0v3FAN0MVq4UUIPhM/Un/aIaB3nEuk550NTbwoOy230Sk+nhupOTq+
KVEcud1SabWqR2IksjGvxcXxXHN4/FYfVNceh+fl/Mj+wPVGaenmj7FMpaa98WelDIJjJv2DmNsH
oN9/dKELG8C9vVffwObJKrmMBm/EPstmAFNcj0fwzsJ6RI0VhEUvKoLk68wwfZY9iX2wvZEQADzq
KgFfPZA9Dd9MP5Lv/mLfkdQZHlFDBn8z2B4X55wLdZfWyFaksKnNy9Ysk4EZnp8DzXp6phOGXTPl
gBtpK3KsbvZn2QDn0po8gUm5BSkwmaj4yNpgwN18WuZpTmzZTRdWJzGUZhhX2Wl95nYeoGi+ROjW
dCMQNMS3Lj4EFBKaJAv/Rp8OaJU7OX1tg7Fh45Tct7eBOD7VcprSD1m2PzJgA1INxyXNX+xYJvKL
7D9s7jEqppve4pnsY37cxkjrHbDmS4c3R5z/o1VDKlb/qH4Q+giYUf6fFMxpKNN6tXGRxbj2/yaT
sGf9Fd9NYpibCHxAzrumn3Au5pYAh8zzVHI2WpzV3KhOwG+ATn41DmHr5yqRxMtmH8qLn2GI3Tdh
7jZqK9fS73F7a9uZB6GQrr08O+JUGY8TUGg7llxB2DBoq8U/k0LFsZT2C5Y+uHESo1bvZACVf7/F
w4THnSeQQoTse6neC6yYBfacz5tIldrTykYK/XwZGi+VsE9pOOBECdVAAyvOC2Vwsq+LA7ZtdLiP
pzw6VrLDIptD5K1z8h2o2oBuZCgnmHwZOkRXbN+8Af/Ac63Q4IwLDgQFRX+DIGChpopFXlesiE3w
d++t1/LA7bT4pfdm2OH5LMq5rAOYU5qucCOO5XSWWTfTpF87mhqhyiK+HtSgIXS0ppFc+6BAqTt5
ryR6isHjT8m65iqaWdCWPVwZPUbO5E/uDP5Gf6Ai7W0BNbDl3TeUApJ2arVIpomlY8u5+m0ibpyq
EGfjpgHhNX1TSspzQS5rfVd9yzy6CAG1e0+WlJ5wNl2Nn7x3xKG7PnAUUVS8JOOexQ/aNaYepX3a
VooodGoRBAwiF0rrjZghMBRuPnYNiIewjswdKxPhX2IisEp13il6fSHpGlmGPc77zCpC8Ifb57jL
3PA+n+MkhDfffVvWTdrrqmLl4B2TWs663lidDDxebJu0Cxw/qr7cJW0Zmu43sn69imkVoccvQuEs
mfZ9Dfe+iQYAYZvMnLja70DR6nk5d16Zd9K284T4+373oLMrVwJLXHhg0X+I7zB7fatLnFO+lNYM
Qrh1rOgyjqEHHktzWc1nIGaWH3xDNul7AnuVfEUsN3NQBMP7h9pGbcsI1F1ZiCrzmbWugjtn3a88
8jCcxd1elfteuKz9Zv69xwBVNJZAP+A9dPJgDeuVdh5Alfb+w9qVH/zcn+IprDoMiddAuHJbcrfZ
iz8aUHxMnOYR73GWLNRAnL3Zqhh6B3jUH0rHccx49pO3mp7Y9NgqjKLvxFqZpetxPM6s+QSjO7Eb
+PGSQ4J1SHY8QVZ7cKqIJKOfzJGXtVOhyKXvjg5Y/RkgekGJA2TR0KBpalRBkRcGxVxNvYZSnlYU
bKIZUMzCQJfoOz3qXjNTqp3I3gOysK/rBSHV4XmMtiJY1L6B0PE1F9KKYMx4+YQkSSrGYGfZtRpy
whJ0+SzO4OJUmkk2qcO+GMjsMC32gDkR5Irw7jvcJWEWQ4zECdyndPTCtjsk/kJ6OVKnxR1NCdju
AlbchkZfjQCtZ8ffdYu9dVhIQgyCD2vo9An6xzbyQjJH7bGhE4vwHAsI9h6/pv2eQPCaRbN/fGOh
DSJSOuxKOePvAG4N53iAVIbIJRfOzefiwOZ07wyxBXTbPSaRl0wt0+cjI5g8UAcaxPVV8+9JYNbB
S8l+Cur79EqWQDxpbWSZL2P/WTMBllIm7toDV0x1fECeRN1f0CkZOyfhVr4x+6Q/v9CCgSL2BylR
MMQiLTbP55o0o3hfYWOa8MrX5QjA1jyuABEDklJll2+uWJlxox+xQTYvhCy+mMWO6W5z9ppiWFY1
pt4+ralU6JGBCgAacc6yKICHuwITm3XyyufygO3PWVV+7ez6c2je7XlreVlddtcUdV27ICNIkdmX
cjUGkgjjmupSz+LfeT6z2x/sBnEdJTf6Nb2rb8TRhfsjnV58y9aDCmwGBysIgdkrXfrGh8vMRjg9
S452QihUy+9L3QjYBCPplRLxke48KlZsVjRz18WGwRzLvdUs+O2PN09EcpTBSifdx2B4XZYTKKkF
G8FO8pp4dald73sg1KKcZ3Ks4hw9uMLnlGQ6KJZX3cofNQ+YNdeyVkV3/eVZZw1yN1E05131bNw0
z0ipYD/XOrjcLJCt+gkdEohpuZG1zhuF6KOCxDCNzgRpYdKkvAoZa9X2i7kJWN5HGP0+p0dgkpbr
SscE7CwPfCdpUCvhx88Qz/MV/ISJIejJUH/hLzxcgVi6Y9k9PCjh6dOdkGcNUlja/QVCfCjwGZ2E
uVkr5ZtnLsaMARrqYEEmHs+dzcwYoMhhkqzuwkFt8s7cfvAZTruGe4WdKEYe0c360TTmmlmt/qPq
T50c67qSkHHHbsveEKkz+x6dv1yyos1KgpeG4p2vxxzsqkbLuiJnqY2juCbGIdP+qJHHHC3HI5++
ED8t7hZmjus0vpgtulkJfEI4ENf5koNhjVvMtAZwnMIMRQ0CK0WDjPu8ZxhRVLkt06aye4nEFw2k
H1p7p8/CjVeQIRIlggQJdZF+b/OS/47YIQKhbPpmpo9HgkFz0W2ukFmn+/XxtaFdxapaZfUrPh+A
C2Wmr5Nri/WnDk+Wgfy59nxlpAIz5ne7QnI5KQd5hI5gm9RP1ex4G1/h89yuZVF6LkONOANp3Xfa
IfXKk1oJX1h6dFd0ZtQoJ/kuxhezjWY2+YdUTvd/ELkLP365v3U0ertzh2R60+4niLHmQWTReJ9k
m9X2uUmbT2LNw04FE1HHeotW8VyvOJv3PAGJ3P5mPcYzheyOcRnExQ44313pkQB4Atu2mqPM6QRN
1J+BIgLStpu2saeO67fJQKobnIT77sRAn+Ae+CjS2CiPsfB3tqQE656SD1pCyimmgCLbMIFGGTGm
HJooVJaGLVMOPWk/0puo5L1+eFlCgLUBjC69YR48UwTRwr/7xj8tTQpNVi4v3QxZLeS4s+LprFu0
8vGkIJZ4yh7P3cvBCrAJz157lppGRf185LyVpfCtBS4k+mwALn/ukxPPGF+LVkggzuVwBl2ZzOBh
wMYQvowffTgViWhhFu+cuiomvS+Ylp5QPxVH9q6dsUSs2AEEqv9b88roSY6xv51EM75iCx6e8YG3
2/+sBr5NbNAMwW040h03hSWDD1OYK64XEwmJlw2WHtba5DxwIvCXU1V7PBai9BDmYnKgcCAy04Vd
buzvdpg8oS4XV6Dh3O/iCZq/0oAw//c4aQsNY90EvSFvkWb8fhXX8kixxIv4XurH0K2Hkl9rz8/B
fAFzcItnqVv+nn/h+n4Q9iqK55JbIH6q0it3oL6WUh0fmjTVgd3j+CmzLgDIEpymC1yLmL0A/ehp
wZF2xwpz7zvFej/IxIbvxiNUm4YNEPQtvSC9v8QCuajLYlV/BTp5XoKgc1x5Ngn+Kxlg25uktgh3
vjhZz0yBcjdVfp2TBjQfqTLiteT545MIp488YT+w3xthRGjBhiglH01QDpGXxYliC71f6l0CvMyh
I3oC4jXbKw5/4lfNIwzlvvSbOYbGY1Z6PNFced53Id0qTvEZErJiA6zzV5ETKt+egeMxlKf5S074
LbXcdIEAkZK/m22WgjH1KQ3J+wpWoDstJfl5iD9vY25hGRwNFrPfcrPmqsW+1N9dVTw+BlToU3Gi
bGXY74A6jwYh5a2XUINnTs0245jQdgqWR7dm1upmGplbTJjTo/6isSUzcvTeub1eskmZFp5vns4c
a8EYQyqkowzSUlwRyxGadyp/jsbyAuGquZJN1+hhx2ISnb10mw9CQr13ikxtKzwajtlxY/xzSP7b
5RZePRsqsn9lnDPpgkHbRhetxzj8Ho354yGOoxBr0Vp2r9KoYgXd1X6qTukgq1+Rb9hFV9FcdSyW
4xRgph+0EN8nOUbmWq+cZcMaRduMgy5hkuW31ieSzFDIPXqxukEGrtL926rMkjtgYLW/D1JFVcOt
bBZYdv0HF6xq7HtHpYO6QTwrqug9kjXbNOuGU6AliiaqWbY4ykhx/opY4UMCH9AKJY3+OCtFq3fG
82kRbelpMaSnPymJMRaKdP1ppjFpx7q0YElJ2xwsG+PCvXd2rNgnSP12cUWgIE7LT1H4nW9gA/IF
yJza2L5ubz/N+noZvQG9Y1gY2//O3d/ReWg9sZG68ZCG6UCi4xmtianHWkj4HhSBKZvhKe7pMHwA
BiDJsG5ZRh2y3l+16iEfx1WHzQU/NZHZtcZ6O5fcXSKZLkGFUjF8QyOVQqbT33K0jw/P/IZUVfB/
kke5hz7Cr9EhNQLvL0MzxdrYT4UMgzZ9JOkzBLjNN3pIelU1h955/b7uIFUDMU6UQfyX8HKprFQu
d2MLqzF7B2RWGhbvh1tSoiLtifMa6WGF7A1gO1Yww5zw3hugKYHarC5bI5x/HjeDVbnGu1YJjv5Y
Hd7rHblW5tHWtJgS2iewKnTzixLTlHUPUojkKflTCKYFNAXvCCKU8lMW4BVCNI1vr2sW5kdf5xhA
TCsDNrsYXQ0agem2R2tzA70RqP9b6192C8kk/YSVvju7Sq4EYGL2yyy1tDjdbzq1hv0lWm6b2kKA
4tXDiXkIUX9yBv/wvvtAKUYOXK0OdeiMUDJJN1GRdwRaERZ7i+NKHyH0aEmRvsVI52UT8kGcfGnY
pA3EJ+T8I8vEFGf0vIfS74WTjvQTDDQf72rVJvB0F7WcVHLpzdOSl+Z93ZYltIGNPSQz74GJYkwr
+p6wyPpeGt8A0H6cjCzutHduyJ9cz176iOmC625PkaMWE55jujuJxu6tn4s6SWhKVlZcT0nJMRLI
D2O4f7dpxKDCRPH+hxQHKS/OoP9q4WAuk15D4aGcXE30k36iMy23/zsIjravHu3wpDyE7oJ3D7Wr
1mTzSmbu2ZKLnWsG4cEBbALKvmgo/zWUOIrvY+eOIAsbS1h1pGiy13Hy9uS4612k3IgmkaYhxMew
cU1+2FILSn/xjutid4iGS+wMFl1y6K/PlmOB2SOkALj7rSTIg9oe9rix2+8Fj9J3xQ1tu+aXFf3T
eVHphSmaBLXYgYxTEBjAAyC2pyjLP9mOXIn+n57DwQBbdVxIEbHr+82aRk8CNCrgGxYX3rqLYLWF
3L0duFl0s/zMtIebdUaP3feqkB6rtrPoOaO/YdUuKSu0B0QtjckF5hrWIiRMqFsOxXJynb9gGcqW
9wIrAT1Cf76XgCxkrntXEGx75lEqbtwX+EUx/IWkNo7PlHd/RXHJjxqQAUxgqqVLHIH7LLPFm2xy
K+SAZny79/DQmCytotXXDpFXcnhfUm+WR+JFXppZTNCGirEE4azyIYT/d78OM3g8j74jmvs80sJD
zfpUYtoI+1iOQe3q/h07iWnzJYtBifgHXB/1I91jVtKTNh33Yxyj4ukUWd4bP64rR8DVrs7xfE8A
seMsXJGbuC1Pu5dCh2Nkneif6Q4PtxgkGJJCAdIePRwsTxqgAAWoLiKXTlX7waLzj8J9rKHZuDow
3+f1BkBv3K9tgfoXX3inSh3tU2KrMDfk+jqtq9x8pb69ceym5yZ5rcWATBxtA5LvKRGMBeZvP4/R
0agb60Rc7nIG2gLa+teCsGrbVdFnRZN5M8f13yODuNywq8yLQJY08z02dioua1PJO2AvM2JbHI8W
sd2P4pkHIyjKhzsAUfTj/k+W65okyuPfx6Qev6yTqs8xiQW1Q3iw8d3tT/Ns9JG/TCJKACEmpvK4
ILugVP1spHHveAb4damj4LSw2Vl0O/W/jRzqshgyj3Pvj/LXoa9Vzf9kJYjLm4N9dvPv8G31NOm3
HG9oqhylyMe+r41raph663an27WfPdZL1lp9LG8fCgqB11EV533jhQmrWYXEpvXC0+8F96flYQ1E
jjmKGijc4PXFsR18hOXehwxUrVRukfqfgYviOsrB09V4ruVFELxfK5QVfckzZ1AQitKf/7HvlNjY
QNFCeomA1SDOmvYzffDs6FENWcQzegjf4UNl49lmvrYYFiFbKQStrx9kCYkX7PNHK9faRJULIQ6J
BcIomIH4hmKqbI3YaGYE7bob5legk0HxJ/6jT+Va/1LeYcDr84G5jS4JFFgawE1JlK761dowFlrf
ioAR6K8NOOkKy/YM1F1kL7EpQL9kRuIFN15eaw9h3anWHA10GsI7SJUImAuICDxLtOiBSpE9B8yB
mZffVA1y1KSYTr+QL8RGzZZNBckFIKkPY6ammLvuAKW+v6fTi/bf2TxNMh8gAfSqQ8bBo+tffx2S
SGV5iRTpQ/7csU9O7POiedVcM5QJqQHNTf168nMuCtHW2nLnVdA1JXPrfrHt7LaS1DEgKOB6a1Jn
rzWKYH0JMafvcbYK7NM2KiyzuWK3b/okUMW7wvGIj6UBpFBQ7OBQy7y3EN0ZEdJvW3LoOCYRY+AU
YGfZke69AFic9QiWnwB5OHOKJbuvdzztj8j+X2T+006gDFFMWqHEMJsGFIAjD90fW4i/BJ0kb4RB
biMrJdroqiZc3dR6oping2O4JIVYMzH0eI69AeHQrLLzYqCldNUX/zsMWxRt8FLTotHOv/jElOaO
LFSBGpVI+HI3BT44s3HNrcvtTsybJYfsVljJ0A6t29LTie2HKpKU+ER3odgV2Y2QKl32K8T3hxyV
qr+E4POa4C/kcTLVN/GozCagzMvPCG412fmy58yDxjiQ6m68xokEWDd3nFq6djv5rGFq03dNBMAO
XSkRTIBbjRUk8DF+2X8iXMR5FZfTGXSpK+L7qW/BaIjV6tLOEAwz3tUPO/eQatjfqnUkRxi48MSy
JkP6qE5NNs7I0n7PmJnlSfmTqM+fO7icw1vqZS3dguxHj5/4EQSWVtnpMX85MmCBePzYVvTE54RN
bcr/3lcJ/I/z74RB+4CRaETBcGZdgyfM+iZ7VcW6jBKVHG2gDq+KjmGZl0VnvWy/Z8TOCXBjmwmQ
Qg6Wo+ifVOTdISm8WQYzzANPpKtNIxDSAl32Nq9dUKuBRPwW3NiH2HLqAs8BZEISWTyuoHWjjmsF
7nXdqQ9X8VjEeu9JMymQjIKBhFUfJPkbV+oNEmzVsrnok0TCk+/9eIcoI4uZg/yrieVWVTQx6Q37
OyT5UNkPLIQ1mjWOgd7KaY1XHl3uLHDdtLtj9gOiuAtpj+McoqhF/05Ur5b7ZsxorRFcOhqIugD9
hDfaXWc7xN70d/5vvaj3aI0Ms+OkPUSw6GtwJx16kaT1HTuvznvN6+clKkVqQ9XGv8kscu5fedtQ
G/gNqYbKXLWQXdBAYFJ6FC1uySeLYgGFoJMqy50T4jh8lqYaOnzI5i059wrjuzGRkZxY5zhShgAw
DlcU+jlLWUg55S7sAT0rsh9k9m2dRKQRHwDelIs772tL7CKGKen7ufSvfW3vPaBF/66RkQf0xxKs
QX4QuYnH9Bu/9bMe6WkMYGu4FfklZ6tYKlhHS1vm132lblbvcExWCDDRkroaatsUfdswtdeYRLAC
p8sljVYYB/P5O13Gr4k1zXFFf51jmPxaedaPf+oAnrFGYMkw2GJMxKMoOFuJXtsZ68XGdAJRtf+k
9KvhMN6AiXuHXrSUWcJdLu80z2CwTZ3EVAF8AiUUG6V9rLqZNk2sfHFHl514QYXPD9LEx7WZzqqq
/iL5YXOvpVtFcz8AIsJKDcB+wuM6VaQqCFuZTDnxtYKRsqT0QxU2whkXRbEmJcTdR4zagjXtdTwE
9ATr6O5VkQUSSpQsO8hjodpPHJcK26u1prbSvM5R0LHcH05mb6IKi5oA8aZtF9CMVec5LzBlI5PH
phKTd0694Yvgcn//vLrXW9SBF0ecNYyWtIWeEIpsYeKP/q2Hzf8NgQUMOddf8Eud9p1gZe8i+ub6
2RDd27t3tNJ6KRd4xV0Qy+2djOtSVDiNEQ/rCL0bOaD7GydgfQ7S2WQxPwjsClewjaJMsTxHcjn3
x4QKFaBVqhgV3p5tLfr1niqqMxOfkybwFpqMUAQzG1PRzF2XN62JzP4IOkARUqc5T/5b1hwZtyY7
E/v2uEjtkYEXzG8XPcDmER73B6m6IiVhqdyH41/PlgBpPkE9q0ViXv8OBqqToK+tvIPRFP/jSdxD
lAljfRntXq1H6ZeCsRjr4ZSkDkbfu9ceknoOHTAlshBp3gmMgPIQJAn0tYB1ICdB3aRwFVqb3y2m
8iIrNrP4HvZlGHlX8N0STtHC2a+jt+Gg7G/c9QMSGTECyBeWj8+DKt88SSVdvMhNzzbh+pbvfk7t
MC5AZDkfo30U7x0Tc6h04z6XJhn1u3rSc8ra2VarM0FWVBPkK18CXacBgjPU3cNZA5iW3sACKbeQ
UAhXPC9RZ75aU47t2nX3Wm1N/hg8BHX3/E4HiLYAvclCFODHz0ybS1DNQa0ksfBL2ae3q3kh//69
C/KTLTzMlHmOwEiidqoUIMbp3zUXqyWwk0r3Ro/ouMyj9C55AjrvN1YcVI3eI6vxkAWrbjzMJsli
G3afYhitKvfsC9XKOJQ3UNMmhb3oSKENLe6SMNQ0qAN6aSeXfNBSK6ZZ8M3zXBXNYmfaxLGen9rc
+a7/TaU+phDoEUWZ4VvLAO0H9SX3eja5L960Ol3SMuxO9KPLt3LNtQOpGTX6Ql5aYVyxjvoROuU9
JFaU02tDy3zwebdIuE6CG3YI7kz8pmmlZqSl6HPO3My6Ao5sLbFfEMjr9t+NQmNU4euXffg7NtUD
uIzb0SG8aHmTH9bI8EmxU40mfeg7mEJwLkSZL3E+cSyQfcfLNJK6icuIbO5B3TmCnwBkRMuUKozZ
rUKKyike8zQjK9xNVEnfBk3fuvNOFQ+jMfowy8l9VfAnZyPGFeht+GHWWC1TQkFpTG814Oqx5G/x
teYDw+KPnrYA95ghnJ8r4JjjWG0Z8DnYAUGck53yia1S5pOZZdaW+A0F7nJyzF5cojDn8V1NBk2F
aPrwHhuTYBb5d837cblHhU0pum87SIrMba/PqBUUmgHoGEJ182MQflzoEuy/S4AjgIIsq/S2I9wl
vxEL5RxukDoBF7sIJo8QzkhkzjN22WpqNdR1F0MUTHt3cnKm9GL93bGa5ikV0hhoknrLjzXSwSw8
2O/xO9NZItEnlkxwOLhtbFisFSX4555PVi4lZkyrIhIMSAyuVjFjT5iNknl+exAMEJP8Ge97dUZt
d+/zdsDb6yi8VLpqc8k5r6dxBif1sScEsY6T2qFRty1i0hTjkrmUbld3lKj74sURvYDp8y4Z1mE4
fo+ZQzBjtzks0aeqUpw94DqKkdWDuqTM1sMeHJ8sxGrFq/RDFBdlDgphsrsAdoPA61IIGR4mOL6B
0lFC6QjyC9V3SCRscNQVwVMTg23nC7lgPqTZQpOi6AdZggcQFYaOfue89+ZWCgZFtJHJrmtfB2iB
6qZV/QfSUnTgodqM+ZyYCR4SJmWVEzR1GgQo/M1FP+qmzxYHep0el+5IV8Rs04K/Mf6boPmvwDBi
3D+IQwYtdK7q8d9SmieFQBbLw60min6+5K8Og93NqgiaW5xF1jshRFgb8uUHXTYaXfmQSRKUK0pE
HsY6puK6FLV6RqKE1KUII8oD/4bObG5l7zmEuPi9wwoRkiORGRGyC6IH3ZzrY/065dqNQFZuq5OJ
eRIhX63UNCtkcx+Qh0RfQRy3P4iJ/8CqghozWNZd1CmAwHuyWrcTnqVr91pC8y5dEaHfB2RaGClR
f2DwyKLw4yUQuoMxNqyFRvwtRwODrybgdaX4gkP9QWS3n1T2BwiCGP8lgh+WZ0EPYSgAWYObiVdb
pWLck+FGbKKKZuL4BnV7uihwreeOW+n0cL6jlQraGn5TBZoxwR2jDnehUuziQdzhHFmus3ocPRWH
3G2zV7jGKNQ+OPEwfWQeltayB8BpmpFisbIzLfkG9aLu9W4g8b5Ge1pZpfAPw0qg0bkcuGTIPEmb
osJoFGZEGMSoBQUEafARt/FSMmmLnpy9A5yAW8bE8T1muTmmrNok8IcemrOdddLkqZa/PMau6aPA
hxfi0FmiTFt2sW+V+XgBFvJ/JggeqsHy04Z6cP0dy1qdYCHL4j2YoqmkCJxaqDANomnE2xMPU0/W
moqQMUSwUDClme1OXWUG98PR4/N72m6xWJ1EATKF+hnIFEMwpmTlmhG3k5zOyinIiKbwEXRwmiQQ
Q8fH5DWJmmjUzkjF283EzyL2D+1gS/FX3SZKuXkm+PEq/HFCqu66NN8R6rnnD1OXv+idy4GJCI6R
TFphESIwRQTAvpwpsokhjO58uUkSlTgHl9C/ckukdPo08w9zcG5+vQ+8J4nKeYq0z1EYLc7Hajnc
LI+8MdJy0BzyVNh7F977mn9UOGnl1RQ58CMZ0v+V7ppwNC7DoS4s3Jpmg7wrnaL781kqBjsP4Yfv
4viOt7uLDQfoqHZua2CMpWodiWw1NYQNo3nW4BR23vdoMprJhY2TR91NPq4O9Q7fpFyF5KGikdXF
toFG1BYP5hEe+wOHcsr9vSXuonOszXcq41nvrxjygqj7WFSOSL7Z8SVCSW3W2gBX4CjcfBxVJ1Ck
9r9/cXMqbPouSVlwhlwXoI1QVNyslPzfTXgsdNc/gYVlxyAu9ICRZnAOUA59D8YJshRhwJoYyYfy
A9GJ9tTWKXsVnbcFXg4GQBwhXdK3ZW2+p1BaoLkTO8oYPYOTK8ypwHaKg67ZOiaY6KOfGHH6WztJ
xQkf5sfj0ZSwVaGE6Ym4Ro8sSvcJB1MI4W4+casjxzV6cdaLeFDi34uMf/Whxq5ZkIhsGW5Vf1bH
UAdoQPPzTKOcuQ8jpJun22lrtTnTvZ8p2PYiOMUG45Yuq8SN1T3KwG3edURmXiAmV3lhPDSgShWj
OiwFcG329AeUj2DuI5i7Uz1QZKjL64WUGSaJNGl9Vq1qrry3gazoCyh8uRxge7WNM6GpR2dKZ8qX
0H+dtxRSEWjpTAQz1ZfYcY2MnloSbfEjicHaQLHeouh3aq5UL/P2n5x1ypHZLMEs+snZGHwENN3W
us+ZRiySpRzbMQg5XQvm1NAw8WSDSQl6mTosYPU9iJ+D9mrpmsANREyViWOpBPRmpy94Ra8qSGPj
Rtt6XPWxSXQvG4s1pktXoU6EjsJCOQqImp6ycV5G9fFoxvSj02itREjKqH0AvyfkaTaGZHPd73mE
CR8Cs63ho9ChiiVybt2qTEmqCR4VXamx4IpvLKTszWEYjT8TKo2TfcHtoUFOXqHwwbtmOFCnBFjb
sGE7JdTBPcfiHkuQ+6Ee1oRp0WXKiwWF/I/+7FTh0RnxIIFL/F7s0V1wRRVbI74NjJwLq2CySKDp
IB32IwWfKaLugRW+XbQhd/86EomQXmG1upZmmMbqxfjgdiP40uPWghmRRceGjLlaOiiL9LonMile
0tDNKCI2Zjk+ifwTgNQhgN47g20jq1O8tfq/JrvjMo0kzcIcyw/YJvWlFN/IYDs5PuTZGNaTuqdT
iE331fgLjdpvpzExBJ7bKM5y/6xPofa5sVLkU5hp0zA2Sh79CX+Y8FkDIzIeUHFVTzJaVPec2Q9X
RWnRyKZ3Sk0ti83RJWXjKLx5PfEfTyw3ITmsqLO0A6dfrZZLlyYC4sXRu4nQRIxEA8F2XB0Uz7+i
HMD1sYeeqUXprs59xBQxQ46WW47wDb9A68bB+2t3unJd4uA4xTCqMU7wDdL1RvUQOr8YVzQ2jxEr
Wg1LAj25FyXLpZ/ncAZU85OvaCzQptipdvpk1VwOW6pt3GJ/Y7Fj22r0xbW45qq/p8KDCWi7+axa
kYYMcMVk8PhFEPWk9WAijrSI/bukZFkrNwA9nFeK1NEtzp8bCrQYoJHgd83bRpx1cgP+mvWl+Ylf
jfPtSUzHO9caCuAuOYTsFIW7mg2yD4v/M99ALrPmZF2iCN9MZA2Jtyuj+qgpFAFNNvsTOOYWH6t1
3x3Zg1nRnBmEEft0V1G833zBqLC34HtNrp5rdZeGzIca0GCPOyYXbNCMn+/au4vFZyDg9/1L0ZZJ
xrNayWH02CqCvz3cLfX1Lk8T9odBW/TUHc0lkSgH1V239ButuFrp8xfooXJLit9g3QZdGqPIynaM
kNZqT35l+7hhqH+7Is1N5uERt7pj6ImX2vn2NJrRzlVwLpRFkwHPKecCohU0Ly+AQ491DGdtCEIB
0mTCFkzOp6PGMZBEfpdvfN7wopij3YNcKX5XWhUupzKoOQwiz3DQu4Yu2MUcxe2Txsj7Kf9+TyJz
5aHstorCR18qoJLXr1VlmGHN/DxHcZq8FPcBRayyODgHEjZkfQln83dhuBFBcdC2NZXWlA4ywYF0
0VwcGbjPVPzkqRb5f1hp2dj98rR+LshT+XxWIBLfBO77wslmkJI5HtwpaBsjbLtsgeUlaNpuDR2Z
vzqEpZ28wqqUYsBeDDBsi7AHgGaF7T918z+YAWlPHNVL4DHuRVFE9bgar6oI17PomEFM6POeenLe
XcU91ULs2tJmJZgESHBiEpcRJPavKrvt2GGKuDW8odsAMHHdgMNNXTsqiLiVB/fwDlBHeHQ2nbOn
LwASdH6SETB1jZY6HY+/CJkr56GULE6u0aQlRRgsNsNBfKhUNFMIP/XpFVwMXfEZ4hwtJNGtU3uR
FsgigC3Azj/JvO+6Sy6Ph5zvaq0zyrVP0Cs1VoMe29wMFJv/oikY2HzSfZoO7U3EHcF8xpFAVZRl
Y63P35DVi/2Cylk8JHnebyouKjRV3aGCJhk31OrZiTDukNCbG06F6HKWVCx/2Vl8Ln2hizPPFVUA
OiG7dzHhgInihy2hA7An+Af1v0WepUOeOhJE+BiSlXaodSA5LOl7xqendw+GL1aN2moIQ2QnO48E
dV9komLtJc07pPoIOZLTYtO5CZb9aBOoqJ6jTdIdxoJlKvYIOpBz5+3TiaKAsmmjuCo1hVo7EEZ1
/BkhTS9BlSWveSy6H5dgJFEqHHH1Mk+aExb5LBtivV3fyLGI7z+Nle9UdsUFyxkfa+dH59WRAksB
gK/pMZ/hKxKyKuj1HZQT0WexOIqbwvRlTirE7CzIB6dF9ejVvoOQUCBJ+OOrkiCdrv5XV4w3CF5S
t4Eku2PRMkcViJOfRPi3GCijlS9I7vQZ6NH7qBA2SOZ41L9hQVS7pTULX3SgoNRez+CyDuwayPvH
8pRQhb6T6AcOiynWsm6y6Jhmso7eJGMUUhNPyWqVsCd1OhPgSRYvRDbRj8pz1mSx5TcX8HFl4EWX
jSxnym8zh4FbhHLVjIACDZqBmENdH+HxVuB+RtC7BQz4yYj/SQOuypZT63+Z5yA2y9qNr2lJTzIl
/1CcWw4mp/sN+ZZZ2+ZRB2eJXJ//TjACdiFJgL6ljkC3uviD7hoU5VlHuWV8uC/Omci4aH3B3g5R
aSlisU4gDLcYab3OIjarXXXOD6pfKgicxsgHw3AD8hjOD4K782kHM3mL5NMyKXyLoNhanjtrveUf
/ooaoOZI/gxIWGwYmVTrEggX9whxXVWd9dvWLtCyGxPtnIPjKvAtOOUKN7Y+W4Aom8TKbu4QrWIa
BSufLOiF9eh5cHauomCe1SJNHWhQ0MEtcb7mubWpOmimsUIFg46aJku5Dhv2g5u8PoNg+XRKp42s
5c4xePlfe4WvEidxrKnUZbuF9qHoESWvo1OMQ8SKk2D9+SZPd0WIJYyxQcJMc2lQcxNaCwVwI//R
Ik2tUHKt29z15DPO6SEXSFJCFj+9jToizy5qpYr3wxC82uCtohS5d8gPdnPbweo8U4HqdUrfLMF4
KqBj+F+lw+ueMWp8YC7wH+CKdSUigSRBdOosQzX0Unf7aRD6k4L4ibuNvKANJDcKN7fOvTDlR4wa
ppkZdtd0Rm6RfQ9UBfzyme1mVCY/9/P0xKNLywTx9zRnKcZhqBHvae/p4aVo7xoqzEbboW51bsS/
c5fONYo9v8sQiKwq287XcxpaCKW8ESpdfwvbraPfXez04dyqNQkYXAkfuxAlRqvFZr6DnrL9a063
I+g27+RwfMuZZPrkM+g8qyrwIK0lj0LyLnwrF7Z6taHa+Nt1X3o0CGc//MohYdcNwnxhuC2I4USz
piaoEufbRQQ9PRlMiVOn84Uz39rxg+jIACNIINljjSYnJf+beKl6x6zxOazaB7w+4HEeuBRV+rZW
gfybHKsGVnK/Nbgn7Lx1l07zdpS0txvCojTIc0UzPd5IfbzOSvSXzNoaRlllpiuO6W36ar0QMjTP
Ft98mvVI1AdfBlEJFBzahN9PQoALlOWLekbClyufP8Hsg5E4Hr7vFUCf9oCwkuUTA+DrQvc/UxHL
5J4Ic4/qCSqoSGosvxxkGgYpkyks1Ym02+drDnqodcP5Nq43vwecFVXdzCvkTaas34l3jxOTKZa+
qVCMRVS0mDxeoQsXYrx+5MLgMHThCzwMd4FpW1kbYxz6YVCx20FE24yLFnCyHWHR7JCpqaEeMQyW
98DMDQYbxAl1U/GEsOr+EgUysRxoLjxYb5rZIZuuvcMg8aVT9tzkRo8Xjm0XqHaj7IcpO9J2T5OA
9Q+7mt6eE7f9CJLKUo+Qd6xJkCrlxyKcRaIjjWXn0UvbkmR1hABYjyxS09KdMIg1GTYksLtFnoCv
KNWO5evhZ329WiUvUtRE35e5wBg+6iOBAGFoh+WYyZbqZOiaDEKF+Mlwzm6Lhqm1pOFtLfv/hGis
JFw+BNgFteuvsLklK4dD7gBIgBDbd1DBmVtnoKIZZtHcJSvc6lzF1Diu5h3Xgr7K/y3QK7voiPEA
EnOvg5TVEmNCTvDfkKwyzXvLkXe5hfdjxbSDXQT4wz75+5446lZH4yx8NEVVxjCH5w6ozgEMZ0JP
WqV+FJunzcGqq+QrTL1WhldscY31HQDlRGnDHRbVe/irTlq5AJr30R5uRKILqENoVNlyCLpfisTE
k+0p98rRwaEooSCZzfDLFgc12vD2Ev5F/ABaGTte6mATqKgBpQarJXk8l2xki8ZJ1aAsojlPc/yI
l9w+eAJeApVD9qjc8K+fn3eANdYssb2SlCMQ1ft7BsoD7B8iQxPQyHb3+XxqksCv3WS4rr3ii1Vt
lLtXgwpNWk7BoCEh/SW1a6dIXRz7EKFwXEywDeJNvAjEtU29RPm3LhNlS2rDTmN2Pw5bK+rB0eIQ
xS6q4zzS7eONZL+b3YYY5Cr92HIgSRJoBogP5/NgsK/FxWTdwcygW19gdBireXy4Ftxdqv0N6eRp
/l7MkKCwjqWU1ItBCMBFJ06l7MK4Y/ZTP9IZpzqErqntHG10kNEpsfUZ2JnlkLktGeOiY3qzVC2q
iIwFo9T/lVcd5qIY+OuZ3HNyy4npeXZpmpwUlG/uod8HbdXzF3NRN95vn8oS0Zm09UXZup6gYrMN
e9/UG0C8RhP6Eh5m4B52St2ON3n7sgtkiUqHW1pFKYkjMK+lhRGB53bmNKVbQtCpyzOEYX3nucUZ
0PFRwZW43K9w6o6K5Nw1u17b4i2TvbZq1o3wg2DBHmMJa0EPNc67lLWUk6ug0pIiBfQLtZL7UUb0
8Pc/iu6SQATGqjIHmmIWqb3ojnQpZnSP7FBYvL0K18q8qOMTGtfCC2V4TW2iITrQhHKBWdvKBwFb
cek3MuSuDKoxPduzspy4lOs2TGnABLZ+USwttQJLhUWckOfalS25F6gfys50KqmGuaG+6ylIvvQ0
2hipwNs4ackpsD7uQyIgmRvz2RU2yKeVddQYOGfhWvYweC8wQajhWACcvfD7NUKCm9FpnTx+G6Ad
V+03ptmuFZvpNQTP6ND/6+2x9vHOJu/+IEM3xwfOPq98uzDHSmSHdG/GgxZm9E/dQuatKM0oiHzs
UJaU2ljHTN+um6Z4i/WZUuHqkR322D1FlavzuxJ6vw5zsaLFgs1OqJCmRVZOjCJmfuZqppZpI1x2
dwf1QDHTYqk/tpfV1QcBisofXyzdjrkWYelkRtz/n9x8qE3EQaxLkwezRiBhreheF3cm+BogN0ho
ynQ5yyQgsX3FipxM4c5DER4CFDtVvVNE/GJuJSVTeAZV10OHDfOJUJhi7fnjijukHI1TFc8qYiqF
OSWbrqCmoxSgJLxCQWoUnlZ8xx8LZYKiGq6xiZeUTFqnIfBESlNpkDmv/nzr15gO/IC7rCNQoO1E
VzIZxiu3KLA1oljbkTizEXsHPAVTpfiSYpY3MaDEzU/6CSMPH9mBVK6VzzeBG/+yhhNmEf0NGm4/
d1XcawbepiqjDONHDcD7Zx1ZlY6Y8IQwl9JchGsGmgsYy8tPcU6b7KDguWfGb0hxcnTKpEtKM2Jj
eiVC2TQL4qgJtcCYm6yUQFkTtukUrGfinPREpIUrfgviulyAiePJIrAPxfsM+4EVdRa2v078ahA7
UGH/zPXCE1e1ocHExRXrNfjFAYbwD/huElBxrFDSvcgg2n2ybt5KH2TqtfOmU74CQSSDg97jhhl5
jjrmFX2cp0/P5idRWLxYIQOhN0z4iyND74WqT2R2+s/ZR70Gm4/5ie0wQI+xLhqw+Mi1srhS83pt
WUIEKX32psd1U13ApsTt2nbWUk1ogRwsPdL1k1Ib6EZcq5MdoW0AuOqFO/CJQWl4tF1bcJ4ZwXPF
wYP3Pi6rPOOe6BwBJIZUCRspN5lYrS++F+b5tL9xmoFJVXxhAQDbQ0UALql9mmnNmFXfmD9VbAmR
Q/cv5cmzJIr0S8Ffio6y5YR4yxzBBzUFriVHdexG129P8byW9MbbBoR5f4PV4PcEpOzh/W0/ZyUm
Ef/o4IL8jGr7SfRN+DZ8Pu/A7LdPiFvpO4al4u1dtHtZcmCG02PHaCkDXRMJ7C1EeXSnYBhcd9WI
C/A98sdzVkKpbUb+FfA3ry6jLyGyAtrOQJ1oVaD1CfDJD0TI6mx9CWeJf9sljJJQOhgSytoePCsd
Wf6MSi7rtAg1hkPSfa9bCbO6MqVvYI7oeDXEvWe22S9tlwabc93U5KBvyYpgQ5E9v/Wfbnbr5kb/
hwUN2ByGj2+k3NcjTKenhjgH1+rFB2J+8XN8Y8XvYURcnnjIiRQ+fPGAvSq9IkCEKKkA9sPsPapM
JGnfUyTc10b35X4DOBfkWW8MjXscRLQ5eyYC/UPwyBQ8fqA6bRvhByeBolbEMhQ1WuRMy0Yg+r0/
YJkNBB8yBpRmHszy9cUQgmbrhknZatuj+Z+rwp2kjEFZ9M069Bu2/TRh55iYL/fa46NEZxaoq5/b
COJzNGkw8fa4KS1fCF8IbXUbhgQ+vXHy9pk4+FMDFmYiSZ0g1SoccTWtU9kYqY2TviGhrsk+72x2
WHcJ72aKncMzA9NTR5marvWjw4L+863NNc7/AVTsWmX2Xh8+9bN7Tny4oclCCe9FuLI9HZdni5oY
gEmGfH+lN7pJLU/FEeTSB4Twl36+0tolXMwN2qYsw0PdKrFWKgFpxpPG3ifKR6zxL8WbTrSEkpK3
FnNtAZ0AYXsC6jxLAvg9lWSPa9ALIG+n1767eRTUIQbm8M5Ds4atVId7WM2ghwsvR5/w4r1Mwv54
8x0cHuW8xdQpnEEzW3q7oapT6QWG5JW94ERNWXsrZtEEjir0aBcPMQ0cc3Jo7Om5CPuXSXexKsde
X05ChyXF/QkQ4+gTehx84/yz0CPAbGYxIVKTzrJ1u6GsYbqvirR0qp/0YqgfV6LU7g71IHV31DxW
XD896199A1EVgXe2x/avHvbABLnhN+nprJ2JO0KDUJ2XZItp3H4P0F7ECSsBzetymWrIyxETdM9+
4aGO80rpyJ8KUBuFy4NZ2Hl1sMyu07p6so/ekcbqsnHpPCpLWgIh1Ga0FYWQuwEqLgsb/ubmVB1u
I8iKnhfaFG5rI1fM7L0nvRcZwoWaJq8BvUhEQs2aSk/7tk8wD4+HvkOluGgOsJW9fLkcHabfkp+E
9pDuo6P0BMnKZxRq2K4klRiHdevasrDEO2KUz4MR5P//zLUr7zRxA5dL63rW1UbK9fK6jcBQxt7V
5cFRXk/SiCsUEmIZ6Fl+1XFj3msBD0PNqs46F4f4j7EyevWwS2CVa+JnwpuE9ExDqjuwOHLg8/Pn
xUvSL+0z1JVeWggA1XLBJXCRregIWhh8lcLuhCz5Ths0mev8fjxd/Sh58Jq22lk170e0PFH59JzH
QTuJgo+QHDxlMTtYgs4Mx7Ayaml4h0npepV/XcZL9MHxCG5KzJno+jTwIkYMsqbHTbkdvkNwtAvM
QeeJh8UyEKL3ynbcNKZv14HLPX02iuQU9VjGyuTNs4kLqQ7az6+9nweOHJSULLk7dXatk/ZH9tVO
b0YGEA4ch0ynSNx+xZle/yUzLTVwCM6/0a3/cbIrKjGkta5zuoEzSSaqCAB5JikqdGxlSVQMfGE8
S4vO9HZ9YcpKFrM8IdsX7jdoQA3OlZr09yxwdbFHLFXc+UNDG87p8CJh1ADZO7FKEPbtKtLc31HB
JHP4WAIy65Cu2OnGlZ+qwbOzKyi8hd5pSE9NTK0hjWFJtqBtndDgUR3jIPDC7xTXtyXxBepQLwkw
GZo2eIaXFKHSt6X/AIKlt7A4PYa72//AvaM7IFOP5XrEbB3rHIuH//gO13HjK1bC0bZ74fcFfGgb
wPlPjFa8U8kLFAXq0doBZ9QavR2bNFco5QXKKoTfNR4TLANf/YJDxySavb+LedA83yaE+642f08u
5em5cyCw1mif77qrC6hx6l72NEPo5LcP/j9AWpSDgHDQezxNXtTlCk8FOmjzfvuO9Wu3CR9ROnk0
k156W53ljsHYPdKi3+yQurNr7nRyYG4U8vv1uMFmqGN4I3w0iA8RSUSgfPm+tjAq4VaVHbd5fuWY
4+jYMiAnVyVE7POjpyDk5onlTnwxiX1HKCwh8VjVkC9dwGrC8MJd1rEduqJ7Auyzv+aerb9ZBbM/
UVuQPELRTIlOVKA86B4n6MOPWT3DT6K2BJemqHcjvHldb2FRGGg1zco6Iu6L+1WJO+p7ypoVZrck
5s8geK65+BClTBtUoc/7juT+dVihGMmgPTzxCf3s64d2jUcjzwU7QIVTEPh8R66DH/GzozkcQwq9
nu0Zru5UNLrLFn2ozA/4qGo9jI5f41Z1+REd27B1B9M/hg3228Pczdnup5hMXYvpFQqVLL7JFnoV
/wxfCoS+wjaRJQoqc/Zxe1i5neLNaER1qkdrKhQKwCnK
`protect end_protected

