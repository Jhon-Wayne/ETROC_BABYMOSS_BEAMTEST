

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cQDd3XIPPlgRDhqULvYHvwCty2ZrVwzfefmANvx1dZIylIMC/SlAcj88wfYJOEUSOPC1U3p3rRJH
cF/G+RPdfg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hcwXqOGXIKp1yMXglvtwKNDD2csTguI/218BbAfP1Qe5YaY7t7J14bh3PN4/sY8v5SUfs5PPhYYF
AVoQ7+Y8KyIAkFOjVjl8Q3cizlaMAyaX6UCc4wmflvCCOjy7mkT0VJKPELyiFH5OE1gTiKu4NfqY
cLpas2QiSAVn/xZw83g=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JJiSVarYWytdLFzHp3wkrD5+jxEb6zxCxwIxMuHES7X4vO/81ppoMZmSB67P59pBX5Chyu0EswKT
bCRha6XDZljqkcBWrrqj3cLRE57UCaEr1RVpDNBMw7hjNrwCb9eTELEwb3X0mZPKBqVrRNroBMN5
Mb9o7SPJ2GKhIDEDF5Q=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
x9rjekK3vn0E248BFQkRU8rm2REs1XV6NiMfscimCVnt3moe1QOgVJzTLPCcPYvThLcZJXwVyFUX
J1k2lVxuHKaC3FNNToKLX7girUcVANbS6jS2AjaAfdpYmQXF6epSjXy+KOWM7AfrGv2r7XNIcV6T
P4He3ZDDIABlWanBaDiVD6NYtB9SspFXaifjJ2faT9Et8gWmYJogYQ4BjXl960BUcxWS5faBudWm
MidcfsfVFpzH5bJ9L+thBkdIh/P3Rjr9ssCSzEagp+1l0DsZGX583KqMaKiaZiIsR+KyQ8Hrld0H
vh5k+kh3k9z7ewkJNwM0LCpa2Y0qGSJOxIauzg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bMGW+/GNxe7XIGxZQsPwYg9NhBUySelE4d3DawPwcsMkcAefxMJ1JdlslSvSp+VjxIobQhkauqfs
plGQEEjRkhr+3m8iz7uiwT6s+TtBZQ509t+m12KAHsziCshi0m7JEPgqnpkYUxS5ZbKQCRgudms0
J1TIIpIIdBJiHjiJWPFKhl2FSk46olekE0MQ/LvS36IE6UC8sP+H2MLZpAxpzqHuZ9TNFvVcyr9C
pc7viw1i7pElJF0USsLWRjDFrkLdXdznJwKPhjmDvq2WWhH0UZss4B7FZEDrUrjB/HO8EjVy2Hj1
fpw3eQ84VC/StEBHWhh2/ovbE1xsoAsXeBE8Tw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pp8HZNaXt/evJqKzoiOa8A1cmkUh/1mQf/2Vkpam3N+hCoX7wAAqGU/zZVMPYP16RpMjeC5zeSin
YvUeVcdgv5x+e+joKUcjexTi2LwQorDqPIl0bCwYx4LccUexnWG6I9/pSM85Q6QNP03F3dTfZ+nY
q8I48HLVTNxhG5xD9+JTBp8D7rjXe9TJGi+hVikOsYhuY2PrwtvuAWhuicAfJnsIE23LJrp0i1cL
6oyVsfKsx+68L6qOWniySUGZ5yDe5zDF3WoQ1oHIZl8/tfnTJcGPsIRyeo3fpk/6/w5zWnz1pHuZ
HvGPaU9zIF3KNoE/3qKTDNhAcVbvP4+ohJfKxw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4784)
`protect data_block
IysePaxxzJCAR6tJ0yqBu/bIdBPqhFsRIW96g6DHhlwwT26leLJchAAMgqwqDonYb73lVfBJjsXl
di/q8LW6Nhh8rHzj5gwsH2BQg5TfcUcydNbcXI87BbFy95EKnz06bL43Ws6VnYBiw2vNMIN8Xc/3
HYB74NKx5p5s00arPpJHmN0BTqGeW+ExT1L7kpTvfHpQ8xjfKTf1dvxMe4rrm3KuVhlP9S5x1hZN
6ImeUR7eqJziQRoukS1Uts9WPKUjcnh9lRfjfLBOZYEW4QyYKsixrK4bzFqfSuZ60HAitAf44VZj
2ZlMCsQxMO2RSR6O1Cm4r1S6qUZI9i0mrlJLsvLuF4K8N592xu4zg9ZR7a6j9Ifm8BUYISLiF59Z
hD1HDrwy91SD1sH89sy+KogwD1AxVNbSIVVnUWB9oBpetRka7RlNsLF0eIfc7MLPZezUa41lPyJ/
QmzcW3SApH9OyTVNfXeVn1v7Ac6E3ndiBt09JNbhbnW8yT1NDJhGXsp2MdPRK0WTqIEc054ec4Ga
X412PedhoOh8x+jYb3+Jyao1Ltc6RfnCVmLQoFK+BmFhkFYbn0tg8TjBpzE9TrY8fmkBqSJO+V5N
uPHs+kBayNZ/86MB0iw6CoqtsRQH880jUDdGT5+NGi9+uJEpTetIhoFAToe23R9Li2CxQ/F1Ut9b
6YafxfZismmme7H+XnDTIAincFAqwCEHuwSzQw03fS5LHveIq921dP4Wun0KiJBd6/WDvxJmbdm2
agcQNb3aD9f57JIxn97rzB9+2YPeFhjXCLUjm2UxdVpBXMMl9OvBVXeFzCsA1pQ79ZrkPSLg3wO6
OsS3W5wgoIJklSB9xhF3fOLEoNYu0lj8XKxK6MaGaJmXNn2HtVkS0zf/LYnW5fu5jllWIx4MwW3F
w/0jnxDWvwduXVuS6bYzXt7V/fnMdPt2yUoU2jTs6GBKZmtdZ3UMdTRocJNjH5durlobD/5S45UB
LWn/UwzWrhd/o/4eCf1mM++NxdkUpiOz3Ox+UAVlvMtZCouGh2nkqay9LNl1DErOKODFdB44/8I+
xNbN+4HMvB3a+bQ86ou2aWO4/UGz/0NdMTMUolrtsjmn2olQWuDsLXXrkK2sLnzdVf8Pel+9QXNk
geU01nE/evd2HIG3bmkxDt0AJRIRHmKmqFiI+MKdMglIeylMq/8dXbuZxbLNhqHzxtiTtkgjrIkM
erh9JKRZbG8qDrYMmSg8+VkumpVMg5tRc1gtwLgcymGkCgv+nqoXO96nRKOeAu7dwbcpuflgC08v
vRWnXAtnmU8+GO+zwR1s21mjWd5rg9hGfutbFfP1YnRgd5cqF0ERMaNP7Z49vSlVRfxMkSPVcrsX
uCrvH2RFs3ORNMRjN2k6t9yz2bfU6ySM9Gx37HgpGYwK5+bpZkuECHNMmJLV78ML4hFjZ6HuGZS+
KHyHpz3DpI76vnVieTrc02+wr7PfFNdp6pKccvaxnmuB/PukZmBUovs43jOz/jcXdVXMdvU2C3it
8k1rS5A6qyQia+zxxcu/VDelW8Dia9FdAI0KgmwpZ5dVFlzVoPazrSDUvPmQRTNkAV0hXTuLrH1D
tTTHTgeuXDQME9ObpIEKIn4msq+K/iURfinmmXRbOGePh1yh+F9qclh3O572OALvbxXWEuTiaHCA
U83kK9aoki19SJdbPzF/7GC7K9JvROFo0ICRKYfLLVHtmn9s115+87K3rEus8Lfa0+4pmdoBU15F
uJO+G+L52wykDrc3JfadJlfQl/BM/brcwbXQDr3wHBEocVD11W6SgjPejM2AU5uW5XXOlDfQTkW+
ZVk9pLVWgordNlzsBUo4sl1lFIatk7a/h3KbDrFtRoM7T8m6I1eDtYPRtN8bjrbgpAtXWbV3a15C
xAfpzYYfz/2CmkHVJTXnBvAn5MY3zxpUQbCBptG2GWwamjiIvvzFRFgSPV/hppYHANfO/eVLSPfE
414IVbl9bFSeIYMlpYyjtDTgLCz0s1Xe9Prd8NL3kZ3L3Beehoo8WZyEJK9o1YAUkBEPvqaeV0XT
Vuk7diYDE7XeOS58ud0j4phVWhUJJ6Y/coGgjnZewxECbz67Ohm16Bw0RJkWExZVErz5Z35elCzM
9f08A0AXZV/gJO/ScXSMHrmBx797VMp2wPOiJcEgH9MX3RxiooG2Lf8/JXDgpOwpmV+j4Yhs4Svf
wZDyOUQqyQrgvwid5zm5RGcqjCAVD2xkITx2WQP2TPzgytaGMIKUNJ/adVEUPxw1hVCP/3BxkALX
yl1UpUZpdwSNXAV5qH6SNIGvr1YgAB8goaCPlTxLSvbNLkDPXzPcB7fQFyLc/chKiG0R73Tqk7Tc
PNcZOZIl2nOAb4bjef7wspdzW/e+CiqWo6mqb7vnNSVK3LLuoipfovFEQbzAFrIlRoOsge+xuQbr
cy0SZyuP0weagWZzQYmzTO4FfONZuCiXoS/02A+WlMYCFz4iKobG4DUiQsPFmCbNKXE6IvG5H95H
oAVOR+j1xNna4kET9FN69Hg79O4skSc94wbXctEqsaRoU4vDx7XXurbSsB61wFXsMiK4iKwkMHZI
lRwbKhVZdcRKDgbeWYkbRWU2WPyHjrj60Rsf7Tm/eskrrRVaygM8CqF0lpyjAEvurk1Sc3UD8JxO
ROOkghVutI5SqhlX83ka6Q3cyiK6r36leACaIstMzLaM7Uvh/iDIn0URiFcNhwArJ/la8xJ/Q/O0
3F5fxFV31p5jE7VDFtsqnyinpyQStCqSXexct+hozpWRqeKqN6zLsSAuRMTH5Fsc4/8ZNf2HnNG5
yxstTz6yBbFoN8+LYA3fg2wYdtyzouIOJ5NhjhFletROVi8+bhKX4eiERKkMURZ96GRvG0mqIPWB
WlOg9eFeJ3hbqtJ3CG3zV6/+dTs3mOtneDlwtHE6PL8Vy722joheY70nvyS5Phq1oTYCCm50SRdd
xFxAPXhUpJS76rqV7mYj0rTsw2ZR/Byz9ZB9uBXUFEyw2+KWA53w4Ek0kQ3pIioo9HYV9meLwnIv
PgE3yfIfk7qeDttrkKeUp8GgbQtji66EGot0kdoxTCH6/hLBN3S2eQJnhceP2s82Me/3If9RpDar
wKien/0KUI6DPgrTwB5/CwMvu/OPCU29f04GKtjR/MhT9miBzVE+PC23SbZfdM8TOZ8R96eeRcUV
9vSamVhhJINmtIyIOLhaiJIu6/i6sjUtZSTAiaXkmWqg29aXgVVI5uQv5myO2JROSI4wFo+06pyn
bNkEUd0hi/95uLXiU2kcDwFs8WL83kKXwKOmlaBN40awT2jZFa9SsPls9x3SxX1QrLkm46TaJDuc
MnF4ZnAatSCvEP2bn6EwxF1X2DrDS4gVupOW5+XPQ0gIYCKD7xzzO/6TtZqSZ5/rYVqQhDmoyhme
BsEIgL1D8ana7PPK1r0Yyg7ExgmktgL5RynKBLYCq35dVfQFUQx/ioenm1ycEkzdDcqz1QcaoKOq
KCrgVfd47FdjhQ6COJnY/Ke6sNYc5X5HiMv+NLDq/X9GyyUIoazDCWDSa3mpIByDZD1Ir5nQS0q/
IFsdlVPOurSSEIVM6nkWvv+T4E0TqFQpCCrjdMko/ZSdpEnGKRVAh4ijd571U44mwJSs5iQPBfQG
IkS8RG7YuqENNR0wzU4lAmhIKB3MSL8lXpQ3nfWRInf101XqVmlYOzm+4kG1b45uZnS6zTC8Lltc
AtdYPBXCzxUPQG+hpN9ofpEwiW6lHnU3Vxdd2JvsoAJWS1HR1Gf2YmhdP6L64XGJRcpU15fanxsw
DClhFZOP9La8cgQBzFS+13zOUVrTL9mPdHM2lsSYWdCf4dAz/M+hXp6z0hpPOwym9BrAh7bXceV5
MtSvLWI4uFq3J0oO2WbXm5UwRRfZ7e2xycjrcTc0Bzj62jG8pFIiT08cjizkd7SPeydONQj9PFqm
pjLxaE7DAsiWHdY3eAu1EXmbvasp11aRWGrZ3oi26wLWQZGkCPk80xucVfsogIHgH7dCPHOZkb2j
73OLJsI8K9h/aTriP68EbZ8jxOAad+gZmEVS3fHBO3tUWxQToxlOM5Qxb2zsnC560/h1Rwzl25+L
gnE42O6+cY6YhwONDUDodl3oV9E3uPjTTYCjEkvEB2PAActW75bX/d+0EACsZyKoRwQ6r54OpLX+
bQBlqnER2hFNNTLhF0/W1J4sUlqly1FvyE4isH1Jm7yZBHUEvY1nS4nca0WTyLcnXJB9wDrGvdu+
DWsJDkAE+XTLEdlvWhZVl7hdNLqMB/wnuUSegqLtWFzpTeCgENLDp0w1S5zbHyB79uKjdj9r347A
9Mp+EFrmcfKd46cmrx48NsxHk3lYX0zEE6/vrvR1MCUKId4IXvqViUj/EMm+Ts0pq0jo+HxpgZOI
IOEMA8jELfQAFRiwZWhpnd0htLqladTtbBKtGr7Xj1HwahZkFOt+pp6NyraOkfNM2imHPpdU5w0e
38XYtUB1mybVy/Miij9ceyeubXahOSFb0cw1CQAWid+JUwwWRmcpD+gc0blQCv2cqm3/KtzDp/Ty
UzFx+65BZBxLQyn8JN3w+iRydRyT8lYth/BATP3gr/M+kwRWFe1shnPQew0yFu0XBWNbvTXy+Cgh
XpF9ot9HYpkHso3z9zP7YJhDy7iR28Hv7gRph6p8Gp0HBaaPvhvAiFWqwje+k11+pho5NKAQMAT8
WI8rYZ7ZmyDfvs9ebJk/CswGNnc/xlKMLmH5fP6YphysTm7JxHVOVSQFpxul1YNIgEnrYIPTRcv2
W8SNiTEkGjnl0g1jDMBa47Nf/vYHZAn2f6NZV6zVNKDKwFHzBmTUhNuvrmdFKgg8DUuaVZA3BPsd
iiQUtrlrFWr7Vdkm/ACIaGQZ74ImBlvpIgAl7kBmg7mLr7Qi/dDxPuQCM9G0C3Hr3/Rulimi/zi7
FJRX02cgF7auF624U0Z+gIREo6ySufdUaFkdjMLQsMzLG8Nf9jNgfvP+iCz/rw9/Hx7Fh4QyRmxq
2F84cryvC2d5doSs41nyzmdkP6m70isrGrxvJraBrrTcr/KXoiVMRVWMYec+X/0vn+pcMFVHS/Sx
R3kV2jgETcpF43R84glhfWUYLJg9fUJNmk7zeNbndNkIkw6Sm63+CXZxl58C4sKnJCriZo2wLSCs
4j0DWVm49e5l9vth5nEqFL8C1jfXd9TDSyDxVQDQhhdhOoVq1mgQAabTYSO4reNe9tBeuRt2cvpq
Nv/LcowXsoUy4BrZCXEiLGhQe2W01/r3YulDZCyjrIQyv76fPthsuJoLROZeanblgkI8YNSR1lpZ
W7NrPjKTq/Btz0EOAdRgezimhWkhYrO+dGT1G5hWD7F14mgl4MATU69GG15euV3zgXwdCFX7uBkr
X5TiU1P5WSHOTpEjqXSbCM3n4+SVZou/4rprCBgPStvtRS/NRgVcL76vyXV6EZfJBJjSlgVghXLA
v+8By2kOOUDIfJ9ba4zBaF0Qpf9iZBlv6UFk3uIcAFSh+tiU797NrEbolKS2Jd1x8WTfh+gnkwIJ
Jjbz5IHjvzDYnDCLkr9j50NEOLJMY6v4CBIQNIfrx7QI4XgJnNlSYb5q2bTp2da6CTMOXMWqr3rX
kwHstcnxT8rxkZcNNRtspHHMXfoawUc7WYSJrGKxHKZ0cYoTet1r5C4ltWJlmgGj+A30A+/j1pD4
95aENudov8ueflsWMM6B/t0vVZuOo3QGD/sbBqq6WTS+E+xgwiliBTLwUP7+Tx1Nf9ghXLgATgmQ
tqPXL16l7xEYAzT58I30SpUPAKupmc22MXTEry0Ul+5AuS8clYuX9Ilas3Ir8kFNV3x9f4jrFkQc
7cqJEBJdSlziOnfgBg1qdo6d01b6cl2lbkx1bh9UpTU5EWpARWBzm5L/E0KKJS8yh19jThP2+ilh
V4xIPLgUNeGFRy9NfCQcj+nqq1GzpJoVdW2IAh6JoMdlN68Pa+4oXcSiw56kEPRWZCrPfoHPQWIx
iet5TWAkOcFQQh2nttUoI/N/IOn4GJJFGD2IrX72rQl2TepL3gk4vdwibHRx22gypyWOnUjkbL3i
HOYP3hfVo8XS0TCskihC/xEcoPcUD81uWGI2tL6AYcMjIfOP2wnSf50XLAo7YwFJXcq8dxNtbTdJ
xPh6afkQaSdtryV5dwKS+o45QmllyCJ4jtlFWtiwDP7hNPJ2TD6w8Onxt1725CRSmGq/kW3SVg+I
QOHxxBEczAu5mXDYPxfI7FeMTEqruQhdlt48RMMUa7v9mCIzT7I1KKgD6Cae0Nwv8ecVjHPvRUNL
szI1+WlG3WiBW3UJXlZA9PV41/PpEWXEw3UW9yP0ij+EVNh02kpbZ2FnsLKJVkQ2HC9x58U=
`protect end_protected

