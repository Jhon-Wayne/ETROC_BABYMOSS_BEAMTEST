

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dtD3GNErsQQckBQO5gsI3QX6KEV5E7ts5EyKqLUcTl1nwscBhbrWkPvqYWMRydPjnBTBoa9evUwI
eW27Fq+haQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oFqCFRLETxY+F99DAnFXOEG0LNv8AH/BR3YZ6PVXco8GYLMMd9KV6vIm5+C+Vn5HY+mO8D+YQphM
iT6ggoff3RcuaQWL9i3ZjDl1GBRsEk0uLTUs9Kqo/a2mHug66MVP4F57SXjq5TzXcKSiCGzszvr4
UvcN0RMZ9JMmnhPbL88=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dUuCsN7w2Ia7j7Q0zaUBQsXxD8yReQ64sMeg0RFnfoygLxvK7nNNhyyZ5VM7b2BhPDex3Y1+/HUI
RdTBcuNkIHefWDCgutTO9TVEdfBY0xOiy4OGbsX/OPTDnAl0LFJ+EeKTP2u1KI+sPxuNMOr6ZAUE
xOxk04Yfz4CZB6x2gMQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xhN6lxizkULPoPRd+P+1Jgxd43aCEBEjYwquDYSQqwPtbmDQoUYoUVKq7Ucgv1UXB7oXSEDiOK5k
UiRNNR4/JdOEYKKFMdbk+2DdFKIt8zvOj6Vy084Z/twNrqcJnvzNIyLxBEsfbYcGK9Nu4QmNiP5j
ewWJ6sf98qt5NqMv30tVy+RX+v8wrK7L63yG3hqyL9j4Q+n9lfxzSTQQIGHS+SYp0NN/+K2/PJT0
uIubVtrxnl2QUS31aKTOVDtqsjeAaGsM0OZVNqDXuWer80fVF7Q8zBgYfEIrXXV/13MSal+q5q4v
wJJfhAhOrW7m+6EFwKbcAXNla3LO2uO5AuXj9w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
riDHupA7EDOiidnqinxH1xY1/c3WAySU7Hh9YnDukuwyIlGMRngvANBJFw+wbARkxNJ5Mop3eBX5
iC9q+75362b91X9QGjDpZjxLCuVZis3zLqDK52AY2Rly6BKO5HoKAmvXIUEYzzWRMNi1b4qsQZR2
vH3GMNcnvFUhGmXsxSKsG1Ypb7JZqfuDSsjRlBY8VRvCq1BidT2PBx0omBFnNJb1jqKV1rgDVQfK
IDms3jRfQKzBFQYQ74G38cWYQHO1b1rDZirv5v+iB+z0ozneNUYQG7v0rP2uDNG1uiPCFKlDisFR
ncYcLkKyw9dVdzITaPdZHnG3mUAmDedAbKkzhQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
E3BMI5Y0R9sdenj86S41gekYAgvOsWUAwBPXMQM2N9bjHn3fHL196RqOaI2vL0OROC/MuGIrq9Xv
vUmCL/boBG9zWccOsrwfp4FijlBojaTmrgC2ziJ+2BzXT43evs+NNB9UbTLUKpx/JTajjMvPa1Lb
Fn3HjiraVE1jWaIccJRsLmB+e9+GuqFZ2tyIsmgCO6Qhp9zUTAWQNT9hX0+OCLU+BjTug+KgDkAt
gbIHzAKcRjh6LG24DQm3ZxQ6cc9XJYXyrx/MxQ0bLVIzih7+IWUHEAXXgVtxO3knw0LSKMNDPn/j
iQ8C2+790TlGBlZ12ewscMR4vwYGvY5t3HPBVA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504720)
`protect data_block
LpJgHFc87AXPRV+CnKKKzsVq4XPuHvo1zq85xFfELtVC/oDgmF8xY9aLXyZPdc87hiXz5IeLcGgM
MW9cK3HELV42AU+5ZWTztP6UlqzvOLEQXObGm3TxxdgGe/CVOUbDsF0DvpeRVvntvGovH/CctSI0
ai1B1bYs2RcOHR2SekYRmVdEGnWHantXxOl16sZgDSjmbuOJPZ2/82hw4v51C2t43fV4KchHqr80
XXjut1ypXUheNx3/yaWDrfEbt+wfI9aFfq2eORbQk7HvxMLg3BAQNbpg7ScSducv6sat6Z8eap+v
UjvmhVSkOKRyqTaOkJPrvhqMTNGSksLG1TT2CFHa9uUC8F8IAcw7brfF3OPyOlUCbRkUFXP/ETx3
JkLS0IJl11p+L4rQfA3VK8HdPfN9KOSnlsnqx7je25baSIvB9LjkaJQjkpJc9ONvc4HA4ZYTg6VD
Jwov/52pZcYkfyLpvpmTZT5AQaZ8YRdKebIvTj06m8AKA6gg5ki7YPD1JEf1lxRtJ+m8sjrsxRRo
/3V4b36rup4PFEXpXSIcN8F08i+iFMF8Jb12Nz9fNfQ1RMYFf8cMLB3vm2hBNAuBCtNucC8m/dU+
NJMtM7BjDYRtcWZ+ITEMrVLmxhKXJMWXmLNxlkEd0Fl7YMXVek0tP2lAMupaf+EfMD3dYNCGmUp7
V1uPX5WtcAWYCx3W1IJ0v3L93kLROhyyv8ZnoxkZuXb0/hol1F91cAao8HJwRrRXe/ISgsJrR9PZ
v2muliylJ2gUeymdOETB9iFSIlmPhWHWYfT2BJpcrAdcmJmqYUP4Mn46C17YV2b1HaVuxBy9SVTn
x1TF0pkNHgQ/aBGGaq+x6PUw5Og9oFrBjZbI4U/v+KaDC6NtK8VQi++Xc9pWP+iZFicDH7NiiQgH
HeJ+YQp0Ur4MooWm278OjtxSe1BrnYpEwClsDBe4EM0PgD1PGdot4nqoQVfZv5ByJkU1iGtIbGTT
qo1FF/Ju+9vfC3XspQb4rpVAWab1IDiTwCQGukda5lZsq2WZE6bIsXG8EL6d4Xq9GRzn8oyPaYRG
zPSCqvJ3SFYDZTLsQuBDM0ijl9YBdl2Vs2FYV3xcNHxaCMPt27CbsY3Mb9UmB1VoFPqW54urc4Hr
G9slW0pL4xzzfZ9AaBFmM4hXBiFx5dDBYbPEus+trwYPO0gzz4JdRelAngzmDNKeOrIoWTaArI5G
VspSBSFRW6dw+Yr75KnUdBQfpjZmnaOiNhBbT3ExNygasjLIP1oVYRP5UKbspp7UcrwBtFumABFI
b3R3Jljm6H/008muvPejgqTSJcVv26DoJNCsosjFRbuCfadIaKiQXUcqJUzc3s013OuIb9XB8pbs
fo0oaoLwDKHOtzxOVngVje9cENmCo9914YVg4M2cr5Skxcnu3dS6F6Y2JAMWR/DRDR2Q+4mqDETG
lIgSTqDpNhWUSxxQ43mzDmBF6l9OPyna4vNBWykPYNjKW3lq1VmBoi70iT5hTDvkXmeSzrqq6p1l
vBS7HTaf6LRcxGF0uSHOpwu3dGFY5p+yVdNX3i2aK/z2++mERYWEUZtkIj9d/7KLb8DBEBGiS7FJ
P4DAssgB5U/kUeHJ5z+jZtIQnIF5pWYG98Gn2l7XzSOti8ultW5H8m/p2FPQ/0xjZBF76pbyE6QE
YZRKDhNiQTxxsf3jlXvTF3MkmCZ8njbkdwTuAHFAWH7ByNwEHWjuNC3VI65CcuRi5UAYeH/YYrHA
y3Pj/6cQyKFCHzEbvgclzXVgtR4G62Vr77eJFd/HyvGRneg3U1zXON8mA6gYVfK7+v39CBVSEY1K
iWNu8IyjI3EdrjX88PjpegGfOJYuo6tbgnGt4ZtZVTK8JXyG4SxUJ718l1tQZO3laC2469iQfQDK
6g4vdlPI4LTAhNjZU5kkEGDldxMnG8lLgHuSBscln8o5q1xBpfYAhS4ns/Z3mWPvikP3juP2/Zlc
1AuSu7MD1yCikZfZu1ykH1KA+cfZ4llOIWUaZZTxYUHOW4ImULQeM0oE5dxE+a2crd/kGNuztTlM
LXrJQcUwh1iDaTCaEwkJEFJXpVUGlMsvO1uJD2F70vJKXifxWM/AxhU9y7pVeVU2v0R8rvi/YALs
mA+//tQ2UhLV2TfnsB2V8Jp76TMbtw83W5tUwTMZCHHxottaVF8Ty/wS39AdFIo6wi6S8xNGJiA3
dylWpONNlzJj956E66vxTBaGQ4Z7qnos8vRlDZRI2u9s1VdXfs6bjlp/U/bE1he3vZaHGyAZXcy9
DiPWYJ+TTfkNYGs2uwyUOaQoEyoP12iGMg6PzNmiicsyGLiOkHHGa/bBYoNO4g9IlLbYFeIIcwk8
awaqt0dd+Hx3u30qn5p0VhvVgy1poAuZ79QnE3be88aeqrAJ3uQpbGAlqwaI+YMil6vaghm00Vsx
f/4FgMwcacbtMyC+QQqSPJfoiniPV/aZnW8oUqePOQ93Ox/ytK5BbCfsLc9lC8yHsqPRwanWBF2T
lQ1c+qUVgA/6Y39YmA5eWqfYx0PqY2ObLFTVl/okQ8hf8UJoO2x2uOo5nPKcDNEuTbxMHVDeFh1m
+p+w5o4jp2bahjnjedN2DH2tDsuTWXzWSjrNIyOZ5prZVwcS/LUEK8uGT7UrMxyfoK6xP+9aAkpk
vhxFzMHKlKUwtHl+WmtzYwD/+XbKzIv7a8A8+Y6W/r1xd8IZBHNEN/8KmiJz1xADEhuG6ehAjeeO
3wqNgaSpc9hhbBYL5n7ojhcrD0qbCJlsXH/RajF9WyzpyzbIkAW0RsQADJNisztQCc76QX3Q2JQP
UnWCYqTo/ZeBIkxB7/FwMeMzc9lBUBVKo4ohj+n8ARM8hW0RxKZWdqPBv7O44N1WSLXcPfY6wezb
iMv5IF3JSCkMJcr7ABlkV1e1ItYES+9aYeZbZNCP8huAdz8Jyf4wujAwFGBMllV9KskhgI4q9G+U
M7EzQD//u3/yAAPQem1UGuYT8lhdQYxbStkul9MTaWN/M31MabSJp3x+zUPdhtT2pB0/PKHvzU6r
Z2WSBDTFb2WsIEsPAxJvorMQKZDnG8/SsPVdf7CU+zCXcNrVvwcSygSEK9gpYoEH0EvRY8LdqpcP
Af6rej+LQV7HhoLnABxCW5taBauEaN2paOEdQ8lBsN811e/NZlqObxc9melXXb8PI6TUGzz1YWq1
itTErjDrxEc1EPgzGQhq0DPueVfCHk04zSIq8axHARLJ+IswC0ucitCwbADGg/PmRvQvHW0zVylU
DWqOv/2+FpDasMf+KRgcBT63H0C3Z+MoO70sf9FIiZI9uOhMGTWJwxYhsdodYAAvi0Z/PxXQG/ym
KKZIO1oOnpzpn5+3jt3qSiuLqZ5OIHYtDsEpFwjA4HsYvwUcCX3aIFK4+PzU3mXzETx8/ABvVWil
XZqz9TZ3D3tF6rkyggvmePm422+3WWm7iewVHrNkrT2V5gyw1tUJ29zGwJ/4ZE4nMeeDDugjYwLh
MuMGKoNKNdeRykRyLqhpc15NpkVuIMqIIcilaed1072H8cizpSu+zTHZUg4NKZF8yN2X7SJH9N0d
U24tpmc2HcH+GDe/XV9fW1Qx3ha7OO4U3UarlsjdIhWW5v9FYmGlqUDjUFI/jRf1SXZVqcfJBi86
fP4zZPGOB144mZmgk9vuagz63SeQTEwYBKLkb1uCn4Ezrzf1hS7UtUEIuxxKNJjLzwubQaR9hBbH
oEikqowLKfJ4Mz1hTMDlp/9SfhrE7zDOQW3mpu7nw0sY6F7m303t8SCTSOn1K6FiU2k0o+268msy
WxwkQEHR+IqmKJY4jjjTmU+RcgDTRk8GhVFEH8DfXj41nF33XpDjAraFstqFtb6/dHh0of3N+8wH
DxQUSnFh9fpJTPhclRwHSLNfIkQt5SOvga8bjWQDkwmFG5gOCds4UgdRNltFPHCG9nJM4K0pz+kj
HFwOeZreJnowyr7IQ5zlwySZ2LuU/tLm1V4zrws3hCsNb1AMTEGO2qKbEDJTqMinDmFb1VfVaGzg
g1HrRZS7PZyD3pA1F37PsitDz9aadPPMYNbVIzs4YL3yPAilB1PM9gCjkk7RKaRUJBX6iuOJpj+z
GCoYn3jouWt8So4LCjvGDhpQwrh1VzpNZPYatAEuqOa3Rx+zY1gqGPkPL3YVs6kvKHmOZE/nRHoQ
sZ/6S6KXCO5MvQURmHIbjSPkSw1PMZnVBv7oo7EFlS7/SNa1HcNVUSW1ZDdR+6HNrnkgqfSqY/an
cE85o9LaL0muF3LrGKJ7XRJwtca2q0YKIjbpqldHOlCZrmqq678lBNPHqOxgRof5DNZYSDbdzuJb
SBUFLMcORFaAyVwhu6ZmqJi78ByDlhmach9dx33CgCb0XSmdbD3Yig+JIZF3X9Rptu+T0uCFw4sb
z+9sUrEqbrExmqn67XEBWX8lwB5GhdBSmoyouxEyFk1Xy041tVBHdMA96gl/e/PGZxT0v76kE+kb
mQ9nm/XSrvhjGrME7tqSN9XQLhPQSjMXhMXWNPtChvPfEx87EkCPfH/syhGLkbYc6UBg6mhBr36y
3HIgnEtmxsHp4o74B9WfCmHN0DXNSZWROP9MVtdpIV5MVIZgMfsyp/UBbvcWSMfX9TyA+TyUQuVK
Q1KTF7mIzaAOMSof1qWCK9k6ezDsOjJfzFbL4tg2eZUEdH3tmOCxj3lB1x2OBTLvRs6+bMs+bfzY
UTgKAxF+7QkJjwrDI2lODDHsR226fSEKW/HDn1dSmQGPGzTQHmKwq/CEetQpZoGmHMtLqSI1x1Vg
3o0BkQhbyZo8OLweXehKtG0yJMigfw2ILJnSj+t5L1cP9sjgawiOm7Y7E+aQcWhGyX4wB7i1Gcjy
gmqgZ8z34BNLBsvTJhXCkLEBz02lBPrk69NYZURGBjrRBayHChvBXgJrjD1bnBsfx+ATGdE7pkmz
enPN4nQVdin4T4wR2so9KFUT3sGolMJANOlBahAg7cb2xw1MbGPx3bATn7CiRHhV4ghkuXM4hx2b
YG3shURCNxdQXUjt0Rb3zvCYbfygl16IHBTVYZH1bn/M+mAH29HA3MgbV8k6Lk0V9067gELSLd4P
Va7bs1qKt0ZkiKioF5MdQWOvMHQxLmIc44mhEkDde1Dj2rKtxg8hr1REjhq6cnSwBEcnxyARnZ7L
5D42EC5ttlYOJdjH+mGry1SdYzI3BcSl/VJ1tZJmlxRJf6zqvp2tOxQVxr3NuS4oG9x00qbKZyAB
QRxcLX/kE/gYcShq/9HRtNJI8EKVZJ7/A2RXs77TO+zKm10kHcncQX4Ai5LZ39q+itNyDzYG8FNd
SIdxFuk26rXn3cvVEbSKikrnYUrtBw8meTTrSE2Zr9SZE0+dL+kr0+/ql0hc/0pD7QZ9HlxajB8S
ndaQsYBse1y8giAnvW9WRE4U6L6KqeSVkBeffutLl8g6ZsstRYVp+HxUEu6BvjS6Aqs6fzWqLuVS
JBaTpnNRv1BC7Qc2xL6sX0w7Bcknr1dmFlZQ9sAzEuSnTX7pMRO1Hrjb6qaDu2+7h7PW+4Tb2sD/
CZiajdHgwFZihcNqHseVcvRs7KcTK4OX57OUv6YO9ogUDVgw+lbTxvs7o8WnqV5goJtFiATTuuB3
mk+DTsv2QgZn96Xt64tY5CmDLvUpe/mu9j/eF5CdInUYwlUv98DZtTxwvSBdPeJfyCMwk2dcMuHR
u0UskZ6kgfEmbdhPjIyaawn0zXnUdlIfYyRPS+XtpAB4RT2IFEn7bdWi6dZXaGX5II4AG1y/fbrP
Tan4raWXbvvSLXTSgxiDcrifeFt5JIvcdnufD6/A+UkugUlLo3BMGvpFaag3xhhrO24gKglBPGgW
HTQ7dS/fuETgR6HGA6Cf/WjfJ8A3w6FEsuIH/95iid7TddUuBICI6expn+jf8z9A7rXNTiLeMaml
V5UFNen2vFvKO+gFlCTEFXBBIEZUhNBR2xC/8D3R66nthWXuaYEBOGksbovSB3+yx6nMgnDn23FH
NnfAGmwPMNnEi0nsbRcgnUZEFUXGUrxpa6fbd7oXHmfHe7pHFXvrOa4+3SJObP6vExhn6FRh2l1e
vvseweiiH8J/hWTuXJ5XY8sB14Pqrqd7zRpAm1G11w3fst/yDuJMOs1E1giTZAHHtQ6DrdIkqG9n
NRf26fKpwwzLMY/jfvDz1pDEdBeiinftH2FgJaNGChyApER8kHYKFu/WAsKOwuKNnn9+J+tKyGb0
k7Bd/yo6c1/uwtATe/6KHtMtKPHFvahwxH70Fgc0aFUCZkauKXajCXu0dzN6fj77C2bTzsnAABMk
yfh+AFBmn03RxPmB/i7cxB6bc+BPhjfPqjQenhwB+qjy3T5E2dLyno4Dj0H0rvYIRLePy5HADmlj
G2uFGK09jbHHdkjMD7mER/swMiOOj2Fl5bcsGB21sw1MHkBZ22YnInSi1YGG3GNXXL/Mcm+CO64t
RDMdoKqfXCgibWVZr6ePX8vKWibnYFuV6R1Uc2AFwxgIPBfDZp2CChRq7lIrzBu1frlWlAfPdrE1
TfVNEnrjUo+kxhcwE9BPW6zeaMg8KnQ1/otb5T4HHHSIfga1jLoYL/kzfVAHUbqEzJylNfjhadMW
TXFvtFgHjUB9J9Eqv15mlOGhiXIO6LZ3j/xKuetsm9YAVHDFQ/mTmytoP61wB8GXp4Cn0HWaJU29
dlRozjssECCIff8fIcUJGO/BKahSo7ppiTY37aVnDvROMyrrstVJSz3dUOzQgv1VCw5o2ipIO7j8
P60PcW1R8rc0f/if5LCYZdDkDaarqrC0ht3CAsnXHkYBY/eObradQ5ZaZjSbI5VOwtQJxNGI/9VM
JEkF8Ua2QT/aIBI/MaMJm1HX+bBm5Z6CL76mMICaVQHGx99piRpqiK0EM0q8F9SwSBR4uUjzEKp6
Y854LPP36V8lflI3d1El4WSzPtt0GI1m72JUqoist5lz3oSR3O5Op+RxENiFwn6lc0x+rXvTpNkr
rnZjmTww7MxJge6pODvM3RUaKk+4aEIvYioRk35mWe6sBsFc19KHwC6A2O+sDrXOUJGQQqXrZFWK
CimwwMcS/8c1i5OPFoNgYAWmM08ViLwlN2KSaeXjgndTqgegcYAySRukvmlG7ROeHNvk/GI5C9Q2
WOGhrC9VNqzyn9U4V/DxeScOBrkinSwBiB23kCcwF+3Ersx2/jpSKqNaeYZ5ge8FaFtdSIFakQ1P
t8+YDTL5ASpO3wWZUppGVL0NW6LkUr6oAgOIzWYK+lkeqWyDWiIlbsGDinCz9juGIC5Nyvz62z/U
gQIu+kJ/IK36MZTTr5zkITLiNB5ed/B/AI9ca8Bh/sTOmpUylE852ZucZ6ng7qpYPuwumGj3E5O0
Otat+rvygb+u1Xp4Q7XIEVsWI1LjTxLjtGYKVHWhQs/DNA+pfs6Al5tsMLRMXiL0ViByRZrmU9Hq
VSAjrsWCpVVVOn75Vt9wAjJhvw0r1rS47B1t8kV9MECdDKXuA8l6gbzOTOp8pJEtXbdP/c8kAhtd
hj7OF92AQtz8Lns5gyFtke249RZGLJlkmGN1nPo9VHWJDwN4TYMxc0NpvtjNhTxivJE8ECe4h29d
Kjy5HNwUlNgpRqvZT687Gw97deryes8hvnEbQzmM22FAdvkG6YqN1L5kZZf3K6GmJfLD22p4jYlY
b6i/tWaRCRXrpGB9seAsSl1BC/4gpsomeJ5JO2D8nUEXABQQMhYvkFxrI8YsciXZuJYh3AOLaiZ3
ffZuWYRoBbig/sQ2ZeWDKOvan4c3/0LwN8OgqRhcIL4J8KyPV9wPBpB2Bbkc2TZSaFiWiCDOQVB+
oK55AILK+CsQIhP5MdrWOipCWlhHDgADEV34nb6rJO7M0GMu6Kzu8SjMnwW0Pj5RpVUfCM8H4P4H
K4VbMUW79Z7DYFhweWM2HMCQrazC+RdLNXYCJ8kPpnPCmPhtROFlA0yvYrE0hkgfGWmfgJvA59FF
IG+n6gqy9iZ6jeXnfK0UUSLpggznmAe79BHRjLinbL3gCCbkvZ4L9OC5UiWx8pDPQ52udFZfM7Ac
IPCWEiN2Z7T/gCOy2hapbZUnEDbMwjOTytGYDS7mVxF4khmDKtKEgbBIJWinvAFXEMfy5RCg9uuO
47EEQuUciItm5/O74CVODDrdc5e++ePRfdvt8p/Rlp6s6x3IX8BP3lbytPU5B7RCJfQfNuUIoEK1
dwxlRgD7BfFP9k9ikNnL/kumuYhHMirF1x0DCL06iRnYEF/8lwRV57kZrc53ZH4l2BlgM2mkJAzB
1xwrqpkV2ACyD4SQsqzbaSvfD+gBwUSCtTPyhgVuPeGiqU2zw7idDhNTGeM4D2qAie8exQOrL+/1
uCWX3GtxjuFcZXfoH5WzYVT2JeKzUwOr5WFNKXeawmlpveboNx6tUpb9djuI+FPjYrbZtw5I05Di
iTtFi7b92p2pAPuj+Sk/iq+B9sZe+pMqbxIHykABvrWUqmk08Qf6X22AbsQHjz9yic1irDhlNP9X
MBp0hRSvNclFzaZPmXaJezYeW/ES8ZQUIjOGuKO7BpDfwIdFIJCRVEN9yMHIk0J6rLMP2lUqjnYx
DQKPKXGCSulfsgMD2g3mB+rxkkpNXiwBb6QFkDr4tvKY95jaiyBxHERvoN2TNaSFJoeYkn270Ac8
ipVdNnaP8hNQEUlJHPUHazF0UoeF+WkaX27x8dpKB5YSMnzPXIEpM/2B+R9eUV2OS+T6nd1SV1Cm
tNS0ZhFjzkVk3nU2XTv7pGDT02LEbY84k3XqUpyUUdEZclrpqhT4DONImHpUuBu/GvisYU723URJ
PSDsZII4DoV4R790jOgWzBZHqJdn+PE+ENar/dZlrvLPkCiDqdnS2OshbW9m20pElC6I7+y6bB6Z
Q2pVoppMC1CjFaHcnVZhYvqRGAmcrqz+a8vIXpDGZcXWGXPdQnw7wIW2cn6GcN2ZpAbEG4T/9zmU
A5IrnTes35eEs/2jjkuarz67vaONWQDxrXbT0rWwmGYio/3RpKjH/Dr44clsRrqmTM4VRt+OVAxg
TiF8DmA7xtU0oZ01XC0T4XydJxx+ANKBCezddvDEVV/PC5nvqWVIvQ33YZaBGhxYcQ9PNkAwPb0F
xx1d/Zw4EuT495oqPexmSi99HGXpiR+k6dzfhnV9Rp31eK7KvLj3hwlflL5EHzkJIm+0KrODwt/z
/i4Nv06ZsnLx1ivkGpCTIgs7vKNtQyy17MgiVtj3F0iFf/V6M/9dsKH9NQ5erUyDvArys8HUsdoA
rqgH8O1ihOfMyEf9Chh0fawS+Aubn5Zlx3Z6yCHC6wz+KtsbjrZAlLzy86bBK1I3AWSPldUYJzVo
/GnzOPKz8yEPBZOaArlYwLljRkzC6JX++SbO9UIFiNIVRRPoYpkgWkokQVk6AEe+4vWfZctGbmh3
PrcfiOy9nI1X71+84dDgkNAAjR+FXnvzDmE9XZHk/HY5IqaF6G44klVMcOEmSElnfPI+/JmDo8IK
AMBQzfEXyNzZGWL4JH5frim7M1phrt7gzjyQ9iBjxQW8Ju5dbUyh8U7VfV36gIuhX79xCopivdCu
d3Cvj8xALdv0H0UKB5kkyFhyswms5lWrZNp6jeWBAv+OOiZQIR1rdFLRJ+x5IboVTY0otYnS4697
4sEb4Iy8J559i9IdEBB8WZTKfDYsjOzAImlI4v1w3Ubyr7YE0ioj2w3eM/CJObilaJiO7QOxNhYV
fibyVdERpX3BUIyJXpIqJTi+z6HbFdadc2c6PJxvkGr/JHiVuMNi5J+o/d3cWzeXL7lwXu2HDFPM
TNOxdBoyi59zAwY0ERg/+oSA8p0mvxzheElzAuuRl2OGOuvugctWVfgkXY7SBGaX2NGuPaWLmgwj
PS1/zeiFopayuSKQP16La0TL60HDCgrC0EZSbd4HtQHw9+SX9PusDdqlBSM4uRGD0WzbOy/jV5Gp
HP2WYuPjUGATpwlmuE7iof3IJRSsl4mhhW3hiGheF/iwmuo1bSw0O+Tb8wWpzswKvwjEuwuUWQh+
Q1RAOM7nlmGhU0LigiGW6locuVzt7D4QbsDAuaGESDrlachyz0XkVsEtCbkq2x0Quy6PBdt/ieaT
67hvLwhKtk3nn1Me/9PQCziiiF44IGoT7bcerM6NdbqNxkuLmON1I0QGS10ctgxfFgoAvKUPH857
+1AS/N/fvyRzGK07JHHiW7v6+iVyg6MLbf8W+XYgB8ZuuzdCbQgmpD+Tc3jV0K3du3GOlRPDAtA4
qf/6TLuIc8t+MnJIrQrx6Kd3oSg6ZG/PgLXjmUq84h69qhpA/YMA07X0hC7qy+FahbgDHvSjI4Rb
NON6h4ENdYG6VpRHOdRDrT3F7VCq0xGLuqk+LdfR+K5Gt/e2QSfIsqeeawRWhYJVJgm3UQ23/IWZ
FkOV4+BGYMdoJ0io5cIx8LqgoF7+du7oPs8EKHJmLIV1+2zCCF5w7wAroDC5/d25kEK0q4nSHthR
11QcwKEYH5sopCB3laX9x/d5uefdwQK7px5vuA5d9ptpAps26Vohvi2bXPkjvtnvIaoH+RVmwjOO
d/43l8LYlgIvsMXVGi+2dk6ebkIC9UdTaEjD3q28fgefu4xFzc6Jokdj2dpnxnArQ7k/Zy4kRK+g
d1uucl5fQIBd5/ULI641uPELvDc5UMY8IQ7lxdovQXFtg9T1VhuHAbRwcNPqVEdjZGjwBaJSdUu5
To+dq1Y3CzLdSVvdvrvvzJhGtQZiLTlQKwnlASxx4BzQtPH8Lixm1mLDz9VbHsHUp1Zj2yE11Aa4
fFuZ1C/PweOTw7OyKtT5P3qCDt1qwLcIyND1lYqFmKXIO+QQBrJTjvegeAzt+tl+Z8DfBj3e4bj9
hEQT2tL468nylFHEy1l3Ke6QkaPlp69nvqJVnBGGVJqWKmMHC2O0WA/bxPOccJGhdzZ65jv8WDC/
Tsu8qfvI66kRvFerSePRvxBbit4e2LMProblvcRMU2rym97a9Vwtd4LuX/UBNIKKv3PMeflf91/n
h/NKzCOTPxoqYNdYqpEhFKdZMx3Ta1rxuY0EjDqemuSTZxISiC1CiAeAZE1kNxPmVHbJWM9sadXz
LGTWYqWXX++8TvEOHopIPzw0LWK8qMrWuSw/ZyhLRdXhvz4T7g0W/7g+BrZqTPKIyQ/EYpiCp5FI
swk4SBlKWOvyScCyV18/LxGumXm3cYaQlHG1hvaBo8ii79xK7Q9sow7DegYqDGb09CUEuX5xqijS
I8ijY91g39lxRK/c9Zt3i2KXt6T9abFRMED4stVmrT6AlGN0Qu4uFhoYCcjEZirD1m+ocd+50wlg
+5z/JSTCn9PbO/i2+rcs4fyjCXH/DpFJ5S0TeTEROSJIJsiXlsFvixI7AqZ4xfXtjeQ2Oo7tKWFJ
uy2D47HSnVh4ET5Ih6wTZGykY3cz3L8vX41OCfKh+g+WPVOZLTWngZjZpFj8oPOz0DkxJYQ1urfZ
JHcNpup/S4hTT6quPMWJOFNMyc+mqfw/dBB2cclSkSE+YYMhRgk58sezLmNk5JaIQqVyUBcuEXlE
K2I+Ebo8BBS702wz1hoMrPfX4MlvTuYRy0UksKF9f4oWpReO945KW+qxZMOqGFhSxXRDNJGJbDXA
j2lwVJBK0Spyp7YY5CI1ffa+a8W9hl4DHbZudSgNsjMC7ItV+L4eFzwJFyzoxi9ycn+7hNUJyyBi
HXaLQafyFLvmaxeuLyd8uFKev6PmA9hJNRsytFIkqXXuIkngtEmrOwAgF6bgUxTmiANVm02vTQzV
QPRSnKwCxkMxA1Ik0HGlxbaqNAYFv93kq0ACMuh04tlyjuQ6gkPEQb7mjCvHSWQy3kCdXWFY1hNb
HYqd12YtYWbXKwmPyX/TskJuD71v53fon/xVgXSeJLgjOI2klWYtAHdbiIOJWJbHkur8cYotDve6
FVIq4jiuSvh0J4rsFC1Bk//HboJZzWzocYxWVMphrPj2YNZUElTBpUpFbqIR4WUB1uxxn1SOPuMh
8BPtmhQg8V3C9t1XZ+xjwLOFVPdfTWWq5O58ua9zxfuat7QfD/13HfalxO+dcOj7tZzNXO/neaXO
uvUMJSHQ/slGqSiPMi6WTVoqjl16ddo4q8A/ym35UCtxsqXoxneVWp08/wgMxi8nQhAspR+8SNvA
Itasp/Vrots73ygeoHAgJ12LWLtGOX7gY1+lh3AwMSCfHTr78unjU+cde4UDaTkMTJB5DnFduYf6
Z/taYnPj/G3OyBAKa87qMpj34tQcT/BllTLQkvKQj0zgih0NfG42LWqMXEDH93jFOrV7cDKtJza/
NvI1oKtiXjDqJgvVYa98d2bnTXmGpV63vsv+22TRyNXXGDR/KzsSVc62QRIY8o3c72XYu8ghH2pu
YIxMJx+vUiAibGkaNz6Hdq4LmixRwF3NJaBlNWxgLFKXCWW9+14FHHktjNeD7a1pNBPbXJ9N+p4D
F488UOfDQrar2qEspcex5vKoK2etrLbX5hR5ZBeIqMpcXI/YbMGPvOfiTJ9hBSq6QK4+Uy6z8StT
f5AanE+pAplJO8VjsvLg0GJIQDffILBo2cAFs2rwb83ELMbbRQqOdVbSf1EtvVRb4pSsbjgQFu/Y
IlSkn6KKlYISfPM1IUTPwqGJ6iYhGIgpBZ1TNHgC+6FIzBBw4DWo8XRlxOnGzDYi6XH3RRVfMgE9
yHOoz2vGApzlQZ8RwuCNOfb+PeQrfxHCEw9r41hj7tDefnc97uxqmsVQrclTmgNtKx0ydmixcl2O
gQXUhHadDkGWavCf0M1db0hgTu+z6T28LQTtjcSBQ4tCZ/jTpQEC2VfxY4Dz3DttQhZm3rgeznS+
ZpWf6d0QVGOozUYiODsYv9UKwmh5c3EoUplKxYmPAgvQ4lKimz+iUZXLSVdD9HMpqiAZf9So8/Mg
W49q6WMY1jO5ImrP6uUXLB6Nhg8csmbLlAEbE7TENxgl1XoZEUy/6d0c9yxAUnzTwnhD3y5NLdlE
unPQsxADexGqe79NCGjlwIq4qWEmIdQf8CuuNYAFCQaomm8A/OM5TY12z/eOmzvaDJlcZY5FHOGF
JbTASW6GUIFWKIRi1Xa5TqMJSrvYgbC/XuMQ/hnObKWETU+m9BYywAY2U5gA3ehcy9siXZgq4h02
ouMy+6BTEhCym37RB7Uukolfo0avqm6aDdb5GqTAD4bd1f0B7FhLTveusKgo7BrhQtyxfJrHm+7l
f6gJO28vU83irkpNbbVZ4TnqQvAd90in+6G3b9sjAzjjvlR5Th5D1XbpzNAnQCw/0jyVaR0qS3B/
gobeJcnZaLuzH+WSW199bl29pzEkRS4jkBSHHLQG8JK4Sn07fZSsn3GVlMB1F+qZsa+Cro7tcpXq
founiuax0TBdbJi+xuM1PZVMJFbbYjUfKqJFuMP6mlLeGn31FO85Rw+Kp8lTLdGcMzMLikT5/tCE
ralfjeLHvXcMlTXYyNGb46a4Lx5jmDuGB2Iizk51F/D40c2ItTAELHDjrlWwGkttYhlKA/2HJlrN
6fjBnHbe+3Rs155pd5832stfesG14+LH6VBJND11LUcgco+vY7oOWs/CvyPhbc84hxmFnOlIgm5W
UH7mey0vBTVKB1W1simqVVMxEq0zVGWp/yD4V84Yn2Qf/ryY5KZwrW48gXYBr58oFBKhSWhoukkk
34FQhbnIJghjkIOKegXP1kOVOiFC2lHu5nKKMAk+MFP88x2EfvOMKtGWS8l0WeYjvb/6gsenk5KZ
vDf7xCCGUpq+p2p+XBJMIdMZqzcTFoMNgckjWpSdcBmdr3YrdGEIHTQ3O7keLkWB6j/BCoIXhOlD
/oVoxR0Pe95YUlxtUhBhxfKE2Udr+x+TXUNyOWeFAvr8rWosjGp7dRQ2CBdAsxavmea+wLIlpR5A
alGxIL/tljfGK5cHzww9QjcZcLhrt6WTEptxa6009gYf3R7fhu16C/LsFF2MzKVNlYP6QrEQ1add
HN4jH+INURH+A7vzk6Br7ND5wBYzdUJ55Rd7tJXrpnTkDBqtPYjgx/o/FdeUr1HjiEOsyRsz0tdK
Aw3iBXn81dVLWXoZcf4kgIfyRUj8Do6mQEAxth/Ht5XTNWQwqqGSkAwxhK+WPD23EEYtkxNW7iyu
+teYzNJ/bh83ohJ7/Lpith5a9ac3cQ1PFIUowEvobgd9p7fr6vgcqw+khzPZPGZCEecis645vbgX
AttIpZB73GHid1bPg3pryVDe+hJV48SvjZQMdi8Oi+vHiDr95JW3U2GQMe9g9v1syMZt+E9ZFXPV
97gI9y6H+LcM2nmNrZTbKVsaxYi8AzrD8Zb0VXP0nGMhaycNMeahyfyXC9Jc2NX0bITmIaPaPIxv
9yGPenIjtS/YDDvaATyTBvjCPJoYsjQMFug0AyMFXBTHwn8HdfLWrtX+1y5FpA3WXGS0/Rzn7i4P
XfiiuX+fxMLMGxsQ5DNiNIa2dgBlbWcdQQfoEM2/BWFNqyD9TNMNJn2fXCYZmuHuHRKlxLp3yLyQ
TgsSkhtqQxNdJ2u9q+K2mGRzNSrjrr0WhvHLdnOP135aq5xGaKOiZ25MLXbcRCQJ6saMDKQVXMkp
1ZR1HqHv/32KnqTEkIPPAqWWFTAQPcEF0LSsesAOuf/AKtJdbnL2hwjADpaFL+9Qf+VlbNXv+fkK
xDf5T26DpXcZTTeQnTJh7BMXFddXq+R4zofNXPTUAq4P8jPnzcQz7spdguw/65ejRH/XZQjXk9Ny
lFhAy7/fUiklxvEGkdo0vJQdXvGkWD2vEYQ3kTNT3vZzNU3xpWmeRM+oJOKUiM5MxWvaR6pl0LyJ
J/wg2y/vfpx6EFbwbrAj7Fr3h2FJmA3pWeve/B8KqrOiV5vv0g/d58jTnDsgNirJZ1Y2lyHQGfMQ
btjQ5FU/rgSd7rrix9GUNkoEc0CrGT6YatTIHc6J3dYeTnTC+ftUpsuYE2eTAWyC/3hS+NMAx2kR
CmYrWFn8Da7NEnT3XDFKmxrjtyLJeDQDPIeCMzhsKVgT69ctRRr/S+VdF8Dpa/vczZc3/HRWxfYB
WeB65H2FUF2STuP6vxbAySyphNuPTCTA1qvzHuL6MSIre5noxUMYujQ8lep8y2sDDcHX6/hMrUP5
SpaCk12hYV04rXC3aBT+Bqoh/rsE4P8mVIUpBLGMopxbkaFWNdy/qbWZHKr8LrBP9j8FhvPkpT+M
m/PZXMdRU6xM1OBs7lCE1jTR7wj9gEq5JjntXxzUDgqEge0ObYLyZgkEs8EhzFmwm4PjnUEEyM6Q
ES+QYTg/E4R9qBgUjhMj5wUtydwGXa0aP9QFwQlGvTedfuyfYCBSjSU+GtL3wcNLodf4PtQ6r2SQ
9yzY18PoZ4AQcZnLVUh9HKkZ/Ye0hQsSyBEkWFDAg6U73Ew5NI+Yriu+h9L0IJUnYuXLjXguIbh4
Z2mN+hCW33eIn+80BeSWt5Z9l1A9kuPF1Q5DK3nxZhnPe4q6imwnFJDLUEe7QB+dRhIFtzzUeB+6
FiWXrj6WgaBgl2XZxZxSn+/4nJlkGvDsz2+ynYc7G4oYqFVPoOqXqt4xrxhGcwmYoYU98HN96BdK
JS9bdhnEYyNZ7SO4/aKsRqW2NYerPOvgY3H136FNW6OSAwHq+3F6xQnk4LVTkuscLYP2Oz3GJN+O
t1xlRUIe/C3MzV2a86wNayXtcIc+wYOKOfTY2XnXUwSS2qHGE35Jcwymd1UIGTCrkrIDi+RYdHR5
8A4navIy9s9B5iG+QLbVhLPOa0W9iTqyMUip7mlYpNaFIMWHiTDWVKy9Xw84e+jxYi39fLB00NA2
VU9S5FQh4TftWiLkS1+ypoBFW3+sdNvyCJDp+l1z7ft3TUq/W2DcqvZ6SNOhvjP+MO1AlXgQWdHm
oqhWYLFyvNnz2UyrcoNUfnOLs19Kb8/bEBHXyUYoBx1C9mfSjNCZ0mywM4eZO+f0o+XgC6jB2Nje
QpxoBbZr16sdNpLeUoYsrOfT7suuD0geU2aoOfu3G/Z8ervZwMbopg4+dVEtb+h9Po5Q9DOHwCFO
s+MdHkEshcUcLGsnoFS2waaDRuP0MUxcTO7hjvdg6W8Y2yitnMZyUANpnOhy4ddU4MJpghppqD1J
X7PAYMjkpXQ+MGDfvppwOL1907BZxBliP5C2oXBYJpT9E4eKs9AJr6m7cv9T8HHOYnsepty8pLPS
uoblH9bOkbz8HI39je58082QKNLmF0sMIwXfR6tQ0l4U72x/KTKpfIZiDRWoVRr6Z61Qdp29ksW7
m3hxYFuqz2hO3GECyH8/s3iP1g7XYNGPTwbBMmgZZXaUT/rMydyKk2hazJRuCB+YUqsl+vxOc81G
nDkG04KPnbxIm6Z2lLp3UFOxezVFBtvnZi+8QBDsCyfXIjw/jstMxo7tl+5k/zwBro407r1rFDIM
r7W0vSmsNekRmL+ZFA92Bra4mvkh9erkoCD9cevPQhjCNd5tWEreEOyjFk7KPOhnJUkYvtQvkll3
kMsMDnp6zg+NFT/8AcXhNuwUd8qW9FbvZR6/U8+NsCfVPOFEhtAB2reMgPQ3UnUMI/xp1FXhYS5b
nDl/KiV6qE0oyGOkQ6W3r+UBdE2e5zZdB7+7iS+LVzER8UN3YubQHNjnMKksnCjTeIY/RxghaE6C
gfCr7lV9/P8207L17/QBjWnlJsriJ9jhikio8PIFFB19I/HleKrgfEsZ5RKofLuoUL/15+C4spl9
sr0KStH5+S1chyrsu/hSkoxAPLYRJOpMTW33yLVyzOgyZBGlYwXYc8GbwNVSGmJC3HX+7tByf/YB
iRtd06Mz/RbB6LZ5AYio7mhLsRuZa5T+uGC08K/kW/x9CiyamZIUMxumhLGJ4goCRVyYFtLnheBW
XrHLsOtmTkgtaS3WotUT9CmatoVmEtQMYgRL8tH8Gg1hZ0yobimC9Tq/MGSpHLkxwyfOtO9b2wdS
x0p0Qe8wRIHV5UxUqiutyD00d7K5YrHgBkzuQR4lELQKzMlfw/saLeylmwHkqZ6MN9vVeQkKVUex
oKgg2e1JGg62dwUJbLuUdC/vECt22ehicTqz8wF/Xl99xATrelq8TA4xENNsuInLpwfkHzAfYjE9
SIjYrfTy6BUmpN6smUqH//1fn93v9FIFeiSRBnxa/yGf3NkHu93NGLy9VMHIqSd/ZkjwHGJ/3HOB
G1HW/nqbh/hHKXD5PTsIXQSWkOasBVknSsjUGjGyMmVloo0zYjvJYMFISdrzcWHmhMkMJV6xlQ7J
RHUE/Ph9O1IsOfeYki7YnOqpgECqg5pOPuyoneEgAvpMyS8MLWASeSS/Oxrzy4uQi/QH/ZXkl9M+
SBokzNq96BCobXhNPjiICuYDf0ZYl4dy7Cp705sVn9/ExlNsagrUbniFdgMwic5DHqbulUKn+imI
IrbrpQcgbm19hskAgET1D+p1YgvVuYFRTsa0ARL7KAsQ5hclbCqdP6zNdx/uWC8UPdtogunwEDXI
6kTinDd9J1yVGY3jO0119UN5NzNGUGhH5dJAvJkd5Mo8zM9Y3o5DfIeIlwdJMjUR04dByZR4LDnv
9/OgWcBE0AZwUCoA2DMDdu2S2/9qE/ym7+sUJBfYhoqSU4x0qqR5xY8g9+5O0Jq5vv4k5BD/OYI9
qmjKACPjpOw0hf8TlzHUNFH9U+ybDkns7w5bxL7qSJ+UYvAgtyed8/yebmU3ZQ/8/q5Nu0KPb8xK
Ey5t82+CMv8v/DfTPH6+fG9lROxPm389uoj51gq2paCqchLPvb5sigEh3ONhF+xr4pEi6mkGetK+
U0fdBD7mvgF0bhG7/Ow1N128zK4cPISvTun77CMGonCh8YCO+MNYlF1up79bSDwZJa9gvoTZKzaK
wDnh+zeUoNR5wwdg+0rl7qY9dkay5sXJu9z7wHsvrAcudwZ0UdnbIdNQzRba+wZDfwmJHz9QCyrg
/4ZRDR3do/AAgyYhgI4FT3FCOhp4KJiCz4NsYSCHA+I0lmCdXMkReF6KNEhNpoCLjX881r7U6SKy
MH/vbWYdMiUXTAO19J/VAS5tS9iz7LrFZreGXAeUXnGTV0LIL21ER8HLgeU2b9YTSSOgCvJlBFCX
yBSwVXKuM3LWTlEl0uz20T+a47/c4x6N0Xvl54mmuesvKjvbMq/DFNjA2ZrZ2rvGngzux2vQY0q1
fQKqi0ESYCqau1WSB51Z6hAjfaBV25vBXFLDEQlleH2PQYoG06NI04eHWRT7Xle4czUfsptwsryD
b61Rgboe4hnRcdZ+fagXzz0oEr1qKYdYQWqTan6oJQNq5SFeBQZ62/SqjY885ZfTOQK6XzggrA/6
2rN8IyvupGoHRU64guh9aYYNcD+ED3rwhujKwVMjfD9VYhUszlRcYFd/5h47EKVuC+hTGvGuZWXo
Uzyp0rs+EkbkwKdjlWoAVRExA+5n+8fNudZ+irwrQ23gV7hAGNFzvNG5FCCMoy00ZtGBDhDrduWM
0NFNuMOoO5HntVqGv9vGOot0bcaH3Oqj0xsQvWbo06xRtIxneYf1+V15dI8vkSTFwSReTcpzKhkB
kKI5r2KHDh7KIcMlcHPQWzlilkwpc9ckVLvYpm3oRyqWGAxFC9Ge2dAl4kiCVsuB60h+4yfvFzaq
lSy2Fs239PTL+3cV49FGa9BWvGu42VOteUIKuMbggCLCcE0YCet/MUFybar5yBr5AFhQn8Fmuml0
FTYO0INTf9rvChn42vY78PUTkmYbjEO4sZZp0mRAcg18AAevgr2pcbiic5eAmzdPeX7Mvw9lKY0T
s7P+EgnVsHrgHg1PkRBfd29UXB3ClcQl3QUERD2wVZELyEe8QrJh0KXLNi6mbKGPtQLf/XB6gQ4y
rMIlVUIlK1Inw7Xu8OuP7wjSIFkgmGCD/+YvnCkKhOkxnPgBxLflZUsbvQIe846E68+Iog06K7kf
wh+rTohYBEe/AuQcnPfz8+6n74PmWacR/tNQc6qTUE5pPjARridrkMbrDW7PE8xhK/GdhLdhlwsg
iYQWHE+M0K75L6pPH4EzFCJssCsN2sqMvrLahL+NCYB37NIjjIcnHLPIw+acoVFTtcXXgf8/H/by
9h3uudieFin30vGvDe2zlC9jP8eoGd/Gyj+SkV7y7k+nTRIx11lmey7OiTF8PC85+fDLqyDRZv6N
dAQ2veqQMPhhIc46dyNbFX2ed67XOmVrssIEw1CcoRcaHVCZpnbrl3xEQYsnAw1gpRBpowihwGoY
QsBUAbG882WcIs+b66tviU4Sgzgc3of4AAFIhwnirQ5hgTngtuZdsKl+KZhz3Rg9KrXt3JdPREpc
VnGotEyntIb7/5cCZSlAu46rg5m6ABtr48pMq1ZOfaPdvIZlXUwx5q4eWr2IRxxRQupA9Zkn1N84
BFRE2Ue7guqJI3EcuVnPbu0tyWZhFvkw1pDd1m466dfzUDrLXlP0GnHTfTQwHPXIkAM8y39lqHDZ
7f+3FjCDRg7rXbxPQom1Ej4eiNEFMTckUhs9Ry2c+pzRFBkA4FBXkgj+6p6BwrQJOnSPeYYPJWoE
pcnJc1IhCU4K5b18a2MSzkgOnCPeNR4YrObNAutN4FuI+9/pGYUZsW3JNDyk3YzIrudhqyktMNHN
a42uWwdLfkxJVac52mOXgRg2D9Ad6TvTKnQkJKMGMpQZiDW0+iQ+o5KmNg7EYlONm8WQPQni57U4
o6YkOsFEi1jjdBv3DkY8LgIO/ku0JcJDnrpMUwvvDfjhEfcvuBMDW0t/nnHtf7nw8EnSQnFm7pTN
RWa1qlTzL5f4D5+LJmUm9mHckeSdwLsnEK4OCynhcBAJvHUcQ6qZwtVydSK4Ai+qj5RCUA2oHbTj
GfN6Qe7Ve4aE3vamR5PI+OXUd3etwhM7/p8qdqBrUDAEnwpyVWTMfasW8T1gXB3aRCMlRNu5telo
0ctvykrazt6fcRdsuHf2371m9pu1XqIAjsQVhKUEcGyuzUlTysjmGyNKCf495st9YvC+vxddG9oK
7OV+gADUxxK9hSRpskNqnajYJYnk52AMRT6jfPf19G3mnzUFBScWYs0DCzjNIX/F7j04NOTHxw/k
S9UT0KjtPYh2VwRZgmbJ6eaVstrHD4YSx3MwYiwkCLRgXQ/3vE9v19TqfjH9zTn5O+O02ZcrNbec
rmVzSPJaX7NdP+TLdJzEqvefc6m0cIl4cqrhPRL/0X4n9ljFxtId/zvTUstkPXb4Ok5AeoKrFNiD
ir4m9c2HO0P4WhviSWScZ2qbw2ubejxBrdtgjhIp15uWZam801hXIzjgs54o1tF79vgP1PmCKlA0
5rONoHnebrU1vaq0jQ/50kmI25Q1+aYxZIt1ere80qq+aaTPftGz8ryXAEJE16hQeUewc4eeeDTG
QrcO3s3cZtyEfL0XGNtaziLB6S/GwWva0OnTlwU/rX3dSs2D8f+4hgPni8fGE+hHu2IjRCJtouyR
4Cy2qCkwgJuCKCjIVzazxnvnPvF3XXQ+2mjYG73mjsjPcwuZhJMDDMKQhwwcyg1uqRPPwI3kg7X3
Kaz03jJ0ryNmbqaP/cpBDdn4UeElSPTrRlBZMO0gPw0KgfjltEjADwDVrcXgy3AESbIjdpgkcDRn
VKr1cBt5it1JHYr6BoLAfLABOXmw+hSasQtLbeX/NHn5L/roosgJacP2zz2wN0UmH2HRFRC4ciFa
5aqDVgFYH1P/9/c8vaurXY9J6/Kt2ZUJ/Zt58zY8oc8H4Zw9NrJmIAjbuWTyh+DtZOiyk9xI0Kmf
EiZ26EIflLP+k8r3JGIrWcqKBFpKkRh4z3Y8OfhSKtAsyBiQCovaea4pJjBGDVuXSXxefXUxl9Lu
uxyyMrGovSkQnGH/xA4gInksH6FjS9j/7TTP8WoTO3lppMfrMtQu1ZZ/cBwPm2nmWXOn8+j73LS0
v+T7Q+k4vRtyEr66ecHYHZT3t4ZoqE+gfpnNds7u8qriPVGGF19frOgNwtlM02Z5wT+mDGrQMieF
nUHWbE7KFpGwWunmj93pyBZtWHVo2zt0iOSRSOe4H/GiXrPdV/H9c22o10k7hkcGv90Ciq0dxkdc
E+cDPVVku+SD0Rf9ysJcGeCFr/j/tu5kJOZ6f62cjweFhrzlqcC5n2Wi0cYteA7+BYEkCqBq+Cyn
Lm1BHf3aNWp5vdASgauQZA5hGHL2OBr9cEFhefLI30kO15Wqh0AOHA2ZBjyyy/X+2f8No2BRY0w5
MKNLDQF6BGnlqjR7N2nJ437/8Ilg+KdXrjmF6PmbvviyODyc9+rTHDM8FF9n7Dp99zXDN1oOogci
LGRtrHQC57G0O8zb9hckdXLRZ9H4oXEdJw/3129L0fjwRsK3EjIfmDYVprL/ji0HDZUpm+MJtNrT
Yneh8UTiNaGA4AJzwXht2/X20n+LDraTAsGlWoCcih0yu3iCsqFzxfFkKTY4BH8qxQI1EiOeBvyW
vz777IZ1IzGBEDjB+10JCQDi+VaveKdP0LRZfDNhg9mKHAMj3HxbVTrKxUjrcCjcg99Lmt+LVb4G
QredhsCbol6OpEIlL0s3JSnWHs4wRqJ3jsRUsI2iB8nWcahMvIrCAU6s/uBmvlUKCMGiUSh6TztE
pO4DGCnqlQPtSciOT7bS5RyCjboYUjdVeYfe1D+TKM5zpl9kSEJsw1cv4ykUd8hffNEsJS5lcQER
IfZjNiMWFQA8/ReSVl4E1kqkHKHOhQKb3Ib/Jn/g4ypnC94ZEruZ4Ls/iFDJCX9Ix39V3NNbfBnU
ZMckBaydHIzdmcEx7ggxrdvKp81/yYMT9zB6PJc/kd/JjuVeNIDuPOKhzbxOzwJrCV4cO9/0+hWg
73Fe+4ktqOu8fzujduRCRMDi9w3AbihvsHIILL3xyQJ0Hiw3JHiZwxNMEB4Iv0HkKdaZcrijPKSh
UAT7Zo/AZA4LOLE6td6TjV4OYdf9nyH6FGw9JMbaD0SFQKrE30WHKr8AlqKCLTrbwRwoKIejKiGH
wEBa3OkqGowsq+GfA2YxJEMKM2W1ZpGq8/HLU2STNNOshRnUu2c+T5yv9HX1ckZc59WB8Lc4Dh7W
ogyvCpwJtsyUuyon9bHk3wjRSTwlcn1bdsIBrVe4f9yN61XNHQbbefNa8GWw52CS93Vh8+teN1fP
M5TvnIm4yOrTNKQwzHfCirnBRfZNsU7LQjZIicyyiFUQhWgnQ/cvIK2YhL23R/57idXiE4auhlz0
Y01K7oLwHaq5mcNY3Al6xyyiigRqF3q4MxTzYWChqyv1GyqcMhzh42UcHQPuKVGOwJ/Ecwgx683u
DbcZylqE8SPqCKxg6p8erdDLYRi3K7ElNwLZ8O1vNsqjQCifBF9y58TEq2DWOOP3epduFrhi38++
jRz27zvIbrbeopGuX+4uPxfIoAIHwSgrssEgPHth1NdZy4zYKwEij0S8Jrs5UqgZcM3dR3ttKune
OR9Dve/fPS3tedC0Cy/dhsPU12auLuN2Z2aZz5W++UrJVEXWZL3DBCqpU7wvK8xEPjXO9GlabQn3
2nT69X4rxGJWHagPC4KeRFFaohxQFysxDF/FHHG6niw2jb23gZjn5xIFa1DWHLzGEumpeh3aSpwL
/z5OHw6Of/+pTJtBYDgFaNda9nLXUQyHE4R/tJhJxv0MHP7D/fFR8EZuHjs5vblVb18QPPvfhGPU
tEUDPRTzmPjCVy9CKcLh6LbU2uq4praW0VcE2DOJs/Ye4yb7o/sxkoKfAPjZkcjU3vxeybWESZUp
2m54gSokDwrbQK0FcM+nnjRi/cbcJZEWOZw2vLoE7EZ+X4OIA4Np7QqoMwR4BfE1GoYpMTlqdVgb
rBRsKROu3eFPS6tQ8fMSEPiDlrVMYtnOxSy91SrGRbLTEcG7j62LNYsVzGCZwj8FtJoQPc8zDuW6
QVs3JXyMEiTUBi1GZzO0/1h9Ob4GUnubb66rscpFizpRDUkNoKfvPp+j5awQXf9TBn26FeDy7sD+
8wN+giwdc8dXb3uz85/ZObKzuczY45PkT7RNx/gk+t4d1dtp0Xw7TTEgg12XxpQ20fq+8FrZ60i5
43+YnemPsEo6rZ10cL4G9+m82SXryTff/IzeUZ26yidpoGNHFoR9d017smUXTsOTY2Lwp+WzP7Vc
tK7t50mmWpwwfgGrhTuINVTCg8pqTZsmtn9s8GL3KExBuah9BfA9m0+vHERzaQQg/56ymwv7x0X6
Xf6tHZiCtLcTKsR+5EiNy25Tmq2tb8tmt6YfbEvSXLX1WTD3RW5vXhhsu3bw58wIaolC5PrBZCkD
2Q4axTILJx+wjUJ+/FR18VlNVAPQhycy9IlHytq3UeJG6lIU4RoZkM6yJRtNWIanYJxX7hnnZCG7
C/fhv7+pFsbsbixDMRTktAzOCipSVsoekP65aYVKenzGSfBpUn27GdjwMB6p++hkV6wc01AOP651
NLaK3pEGgTwtfALwvA2BWPWC4eCFlYXdjbdcHDDwRjmu9ppboHu9745L+6mRfs1nQZt92J8rlmHd
9RpE+z3OxcN2rxk1DbktUq63MMVsN6kHv1OB1wj1PgMD9T+SuwCdV7ci+8TcP3vk8O9NR8ALNcE8
buRvyqeWPrkm2aGX5DrOne946qsqhS3vJjgrzPgciTOiaMYRsxLdQhF77wU7sVtkDtuTA6X4JUpI
1z0dyPDAEM9b+6PvjfzpvDA2hcR/QppbXCXXEkSZWAZJ8TLu7rGxzAdoWHsfjun/4jl0orl3CF+9
rU4lTumd/ThLET/OGha38r/wutHn1hKdVuVWI1gs8uc9pbFESKCiKXEhrESNlzjSRVCw8NOUMmin
sTiMym+j6x6p9UiRoy/oe7FGyuOlC9WDEZtYCUS+QRjtQP5sSNzDwZuYfh7jqsvadxWzdGTRPSYJ
fWmu33Pe/sv0hX/H9LZy96CbObv4x5I7JacZLZbrgZAGjsj9g3JZA0VTgfaco6lzhbiPWFjUqVFM
/oLdtSAZNf1oVxnqNGsAeixLBJKuj9c7CHCTmKSftnlLu6gZvDFBZTcubgODBKUHzXjKZ+Dw3FZH
4tx61wgrHIYopyN3kgah3ahGekwodaOVSzChAABIFyvnWTKQ93D/sg5SW8vPnu94hv3FJ1QgSEf4
MtUFnRIJb39D8Ab+XRXhQVmobrSkUvesdTJXyxjmsPtQBXBWJZVhzqKAfzdK3kVbmj1QmIKQ2kvD
dHcJ4ntVKSXm6t9xQheyri/vDjWKwhJAfJtG4E+ExWas/Po95VdWpoXukaRyW/ak6AJB1r+fiXyO
j9PNUtbc9hzL3LKGb3bSVqeCiYBy0v6BTyrgOK8+4uAU9IgqEAPkg3KDpyiiwYL+ok7bkximHPL6
tRRrohe2Kkf9ATUTxzkwDTWm2JXIM9bmV3DsHElcoGGgGzUPiBu6HSd8qUqVaZi4ijbA4m/phEg8
GZCHPqQKm57boxxS2sIIkHHYW4LqkJ9zCKe1R5r8e/HFHDrAJ2P77jq96aakeYGCLuJYaqvt7gyd
37Knj26bwsXBYKQmQMqoqpmtQsvE4Q2ptxuLB07vf0RaRclUCPg5szbB+K6HqcWshMQc5xC5G1Cq
HBWplKdAE6dntvXfHNBJoXSh1bvTQnhfff64We5EUzyk53IbBZHnOEDY1kg6mg/LXUuCczl3V2om
fCvgzRrnr/Rkz9QipP0/zUCy3U2MkjhMrGsmR9+AsWXdr4FanNGq3y29inOOMlCFS5JQbf8CY1JH
ezOi3NkosI3uvZEW2+paYOrBBQs/ZnudC1E6/ZUToqKXyK4LYAdG+9sZN7iqEOk01Y8awOEfOYbV
GwE94RU79Ht2jsrysoJjDH0xah6e6//NNsByW5htYTVtHWDNsdN3Lsu5+Kt13qPcPtZmhuVuh0ZY
1CqTuDUU6YXxQKyjifWoOK35CNFKQq3bPVnqDRSiDY2N7AWWUsYCKCuWLldhmLa3UDTQfDAuNRLv
wQ94wq0hZg2KkT7l3u7lrjZitDGELe6Fpw7kNv/XTNW0n84jNVeuEoH4e5zp6KOSzGGErWN/6NAW
XWK+0Gy3l391SbixjcQBm99NzvrHKzY/1cn3qCUKE06AnRW7WMUxZLj9al0aU/5fRb+yl4i+Mo2y
kLiZIALBd3jFMjH/bmCgpB1QOb3BIS3Ih+Gk9O8wl5qjftn6BCoQ+9H5NRyX4XGFwavB2IUMcf8/
vEJ5/DpSc2bAmPrB5erYSKKqxi6bnw8ydCdUJfkSQetVthHtn++2tmnC48M3je3t5yhPPe4SPIOm
YG31t7queoKzicfyPeypgIKMOTKeQ9oEH4lxn/HaFrICmovlZqMcnx5UuAOYFZtyBvU6C8xigXQH
7snqxRBNO+UzNAN/SavdndJdl6LBewqN3ezNJB9VqTVpvg+PB52lEUCTGmtv1mqBioXzOVdak5GZ
wa3vycsr/IT2ZNWAIUHqADqq/zwdEYN8/2wvgTjJAdlfvAt9oU+ieypfjPlZuty9BvF2GuTzBRmV
hWI5UqKqgkLvvFa5TfchGIVm3cqQ3EbVvjHmeMVyuIhgv97DegVABNNnRkqAiz7QIDVMIf8vgY6p
qBFqA50/jRVb+1jM8mwwrDctvavUkOYm8g4WHsiXhdbrWkuD/W2nd7cEz6DYZkCXdPgOul7Tjnno
+naffyxfEC5OrAghcOql9n0DnVhKqdZzucWoZmlwD+/jQ7K64MZ7SU/fzQiJcQ3qbAu079YhqXqC
aRi2XvgukCXfxV4y2F6TLG1OxjabSnTRWmrH1V2qYc7Ay4JxjMV94EVMO3jNGoFTc7CWfcFpKbO4
fsNvnOGQOSdVhc+bDdAvzaxNvRmEUPGO/1s5pA96fABl4Zn9/fTk6WMXS4j4iFlbTDkwLM1NbIbT
eVyFYextSPNiZ04GGvbPT/5Rm8Lma9JQC/TN81GUsfhpJa24Pxb3sCZsbzKwgMZMvxp289HDIpK4
Qm2UUc8OYJHtVTbwsFUE7sCdDpshItLywmwd7wylX05QSVhV5SYTyAism8jEBT3PCnrM//sGELoJ
rCTe6+oB6iUSL0lYrWaJL8VD/vDHRwStZBHbEyIeUWp1NnodppdP6BJxwbKJCYS60/3ALLs6GNtR
Yq1IDUevwzB4Y5/jupRWvQHkE/weL9/AYZXx36XOXhLmkNuVQUxm/TTzYD4vQlk9LtNFmfaQvsBe
YK+DQLjvwP4qD4tV8a+7t13p3GwqyJwJNB0ZQ1BCzVGouQSBXRJ9CjLtvIhOVK3LWsf+whAsBW4v
KKpn7kUX1E55eKsoJcp+X9vVSqImFuZw6865YZPQk0l3T0D752xEicb253kj6+rSed/oyTrN2RvX
ERa4P6Qacsb6SBTS8jcOfDFhQeamwnEl5e9jopcVeNrQPc2vjeiOvphCHUk7FaRSmo3fQLJRsUw3
8eNQoCSevYwdan/et90qkCzqPJK63lDT0VSAaIZtVlXeR9xbvIkMApoLA2tzHaDh0hZc3Zx6Jnga
J0GTLtRd5/E8tRxhGy5vnI8kUud+SBY+eZk6f7h2CH7Th1d28mE8OVhO5Em49TPCjMy+Yj7JkbTn
i8H6YqY+GPGMXGUXTRSl6HX99MAPdwhUQLPLIQ7ItdpNd5bMj+6tlDfJpFjA/FH+LeyvAaOCZzoO
ChT+k4i7UHXMTZohsKp5duUJii4hoGB+LiBcF20y6QlspGmUZ67D/yl5Gnlmn4UPC3Ca4iXwCdAP
vrbrRfyobjEQivo75DenJADLkAsCKNr+PILU0fmIynA7O6+NXGdU3qcZUVczTxv7mmtld+9X50Zw
BEgLcyhqa284qNaRuDOTBFxV2xzR7Mfo2ob69z1chIqfJ0GEw4bXtyDG7nZL3qAZkZxiJtkamoYB
kmKsAw8xtGjmp0JlMh7ZCzm/4M2oJDODB61yUc3UrHt+yoxpi4P7vreqUxuiI9gCOHFRcwIiFZjU
HKoo399nt50i5lJxva9zicx4ZSkaFOXPzrpHQs7pwGB6+euQfD2ZBEvSxVbDkjyCIXnGZniIf0jh
/uifD9nC6EizltYzMUg+WgyIVIxb9ITHjZw4WdregI3/1Q7gQSLnrqcigjpKa9Le5dcZnlwXnhjt
gjqaH7mA7+9jsYkfyx+xb0GME01Ox7UNleX3GGV64sYDNdukV3q2Ietu5z2JgGpTL80F/G7Gif2R
TVMXxUlw6y6euSxlJ/tDM8SqtKwyGUDhwGnvh0ijWct6ZxSmP3LUzdluU1RuQwc+9sttjZOxdDaL
PR0xEWqzHBBARojLsCFMpD+dtuBOlwXBxfzsqfVcht0ImgKdhG4mFv4BrrKScTnQMpfUygEljvy+
8ZNteK3Q2IMm1ididfTrqm3zF5cILUkZMnwnb6Zdtoxba8SGpFdMI37D+m5W0aaVJjjGyaTh6DZo
Ssmud/Cdvx91ELfA9WcJM8R40FZI98mg8u2aFhMBePpioMRwwHyOX6TCTqmzHj8H8Km66EIHTJX2
PjdHJYciBg6Z0Y+9acog8N8bYTTlq9xNclb7vzhzqpGC6crp6XjmRcd9SsaF3yloyZL4baWY2asQ
I0KkjvPA3TkV58r+KqiBSy4pxfEl3POHuuM+sA830SvsUJtKuqeQX7ckIoWIQkj2lTsrJrhJSp1K
mZOXTHsb8BrDQWl8lQh/iN4oLjc39bbBBdUmgDRLdx8+hYoQeLX3i7KkCjbMRAzAOJ7NEMAmYbrH
fKFy4N/bIozSWGLtQ/4aamc2uwx0RcwV4HDwWtYzovlXv5wTyHaoxf2mvAM37o/0l1eYlem36qJl
mQQ8FEofPVtmfK0bM4NPA+8pWTPM9kYNnBQh9kLHRaxW8Zu0j1koROp4bnuQdKcevpHtUNr1N4IY
4Nm7Y1snm3Et1MtXf4/XVE2Z+GsToMcBzOQKK/cqd9ZZUSkeZepCo53bdpTeQe8FjhenKjIfLXcA
JrSYahtxuCLCnGp28wjJ1fKvjB6ri9e+pabsFoz7j01qTrzFzubnksb2ZTLGUZxYA5XmbK0VASk9
MhO7TS2kenprMH3V6qQ1AVod2VanTyLzarZfOpD6lJDhFqLj8YSK+eXxXeOL7JpnOix0TAW+W8nZ
yStOccmW7niTaC4o9mj7OFBylShkDVecfD1HXktQiLtHMQk7H65SwWgyHbTFUZLsOzT5nP7x3UzD
HPaKOpx/cjOSZnU8lslSDVsi8Jxk7c71DQwEO2UiKe+tl8SRJpzMFCAu9Z8P0b321JRGhiyHCiu7
7v0QXfjNn2YryU8cfeK/eEstLnjY/xTgjsUqo7luQH9AqRuJLgrx8NTFjzcMkOEGt9HG1nscPWct
iph+bQflxsfKd3y3pPjBPjkLdCPuNsdCs+AehR8LdwVVUQF6o9LBTmgaxgYjfHZ3jQahz7GztzGh
w0RNIVfNf0h5J+h0F73RQK58WXPHNF84PzrZU/wVv/HL+mBUE1DBtSmaG2FRhh8ME1S6UvbrCmvy
5HboFwISvIuOMnfkc/HEOdEI4tvUWTdDId/QYeEWB6gE+Zt07ffRGE0FPbv9gigp83XxOpYjiU8/
1NAtHTeEgviZij3KvLHd3hJz7+0nwJQGetv5SlIh+ARJYvMLceON2yxImlS2fvJ5l/fYd+j6laj4
dbOgbrxq/Qm7JfahSw/8aamDWkcBNdkUlhyEtxOyakHvLKhM6SH+zRFXrGoABzxwKP0HzoAyRBm1
L3FpHomSuUu+RTP+kZEkeRKlWtQs4jeGA4MKP4SU+czzHtpScN3fiyvxBE30K0AJ2oGejZdMIK8z
CuyhcDm1KHlQSn2r9yBUttw+Wn07KMVZBdHO0kkln5ef5VquREKD9wtiM33Y1VTgV5Jvx4/Z0f0h
FkKniLuvachK1TNDXY6MnSpj0A1wqno49cmKqjxlvoskKYnMvjU6mITZf9IR9YhOIsyMUCTGFdxV
XFFzvsgIvyeOlpM9LoeTfMQhqOtw3PqrACXl3znb/DpLJfp7IEsCCriQyjMawfpY/cVobx8tDy97
g5yHgZvM+j3ds2F8cVxVbNFVFX3ey9TQJvMH5sfOp54rvbX+hsuv0fheukWqXytg/tmdZRqjyFjt
o13f88oOZzyqHbfsBdKsr1K4zn6qv1+MEW+D5DwR405Hllgaca8ktieA8dUNjzSYf3gU7D6H14lD
VIUOvF9bKEj4oSfHs0sn/LFO6b6yPgrRksvHbfGVqeAXCK8g9q7SK63l/R1mBc05K7jhyndmadYE
+smFAm5h64I6J6KnxXeBkkVDr1KdZzOP/m96l6a6X8AxsKQLzfqdN4x3GCwb3VLJaJj5GVYF9BMZ
hZtcbNsGLnlrKDJ9CfSd8BMmAhqruGAgJgyWjJ2/cwSFt5CjBKRey1L1Qttx4/nW3vfFqDL7yNR4
/pWZitf5leM4SQPW0ZQVwQbJhQAkqg6QVrXjrjZqsOSrFwhZgaOrivrxnl2C+KJdDoMYHTTQ8NkN
kaudj8ToPNDW3M2qBeCvJQHV+aZO931TQYdj5WW6J4k4A3A+TypVNpjFvcsepoI27EJlKR+RRd5Q
+UVmzp7mR5g4MORJpdnND+9/hKXn9DaOSEoZlQzKQMwZoBihfj51fqopmzZ8JDubNf3XW0nJvd5V
uwftpd/N1kQ9thtaDLF1jpRwLEgV35EdxFizgCj0ZTbr7BZYNP5laZymhNY6/Izf6g1UxOCq6oDc
FJrb7U4eph+eoyFGY5vNSP4Svmf1qtRFB562HX+eFxblG2FvgRB/i8ZWnIeK/ExOMQHcVxm6XIM+
jt3w+RKFHz9myMTWz7xkdTY1cbDMUdtfhSEJ+5AC6PWhIRYxE1pT6S+Zsz3XP2e3BRjgZJteOeU9
8+ilYOqjEhEf5VVPPWhjb6s26OGsmIOKLfdw4XnqTRYQtMwVn7HzJxJwvxpciVty/g90zF3RtsDl
9Hi97F1tctADSz/H5VchxRS5fVUtLdGT+WMf/+79zVT0J4U48uKi3wsuY5q9+aB3pDrK/z1EnZ/1
9B3OcI736wp4VpVcQb6yNqu76mly5SeZUAzJMjjubAYLusJQ77HH55Kq++rYNKd2e+4I2aKdh4sp
Liz8Twu3Zk+XNN0AUwV1/Ut7tDSRcAGAj5V1qYwVurO7NjNbYNExLGVSbwyBNzB9adpsfKlEezIj
gOTv+jEThlaQiYnyqd9Y92bYMmeFYDO4GvdGGO5t1C+3IliUIChDqc5ZIfhhFiB497F1eMQ1Ew+k
pSv5pnRh4sADEOI0K+cb2tXgZ0nYx/DyRgUoHwQntPAMJhlkj/AyqsVMIyzyrpVOJb07ZRohhICV
QiHSjitJzeMAcqUXLve2Tb6ik2bcJN/nYnVZaokyzoWxAK/FMmD2f6398sL3ws69lG8H5VNdtPpJ
HsegQDCgws6JdNR3Kkv7eE2qgYUsx4tkbtS7/JP3tYRYaDS+8fo6cFgFZ2328TZWLdh8J8yPe4BO
L6ayD0wFcHwfq81JG+85R9m9+9MtjsqsrxuSHLcQxUUIaUXT0rHL7csSYkv7LCKhl0vPcyQYVOph
vAcdoL3nLeLRWLrTHTndAOtGF6o7qTw5vUT7DSnmgaza1k+BZCe2jJtu5d8ZqjJ1G4kbd8XYq0Rj
902rnZR9TbG8KMaUXIiHLSSyinvmJC6soly4Vp235IWQHzdi9PkcOu86qfmtQOZQ/EHY61+HP/Ig
E+HYMwwE+hJtZ+XYRC+xdGRhkoVjx+Bdj6+51CYw0+i5w+Czhdp/RQeDFP1QFMVjGy4zgePW3G6p
iEBKSgIuwYCtVR6qUynNp/9VrA+1UroxIKKkHg+HnAnmfe0B7AutxD6kZSzWJ7VomvJzMGwyPEZ3
WQExHxvuEchTGDolEHuOYNrkU6tZOmq96xYDk4NXoI5AIBExSrXBozzynCD6+VLFq0+gCAlHxYlR
pW9rGJqgVPsFjvZE5qEb1qpFvclONOH7JS7hDcg8G6/XA2j4TYFQ3izQaySxKsGsyPp0ogRa9p5b
bPV9Q+3X93/9YgkZ1YdMe5GZ8zB9NsAq4KRQJLBplHmfrOL+OegjwozLCb3E1P1qnXWkT/geIUlP
71aWi1ssBXpI/cLguNH32zxBmPb9VjFyBd1tl4+9Bd1dxya5SpgAH5FsMIWJYN8W0R3taQZWwJaA
ed5dJ3o20ZXnu3Ibzdy2p36ol98r3g0vL3rizAy3St3ky6wUUKNfdP8asBxBV/lxwkJof+TZ+lfj
d/7qtGrNvkCCix/bjzyUOF5vxbzronAA5pDBtoNBFAZcJKMw9lGMd6zEeF2cwjrwCNDNYovPBwn6
BzeQJjOFdyxxJq0GG0rIk+O2KyqQ99HiYqovzANgIoMYr/17NMtlbKPw9Ch7RK88Axjoa2JLtnMc
y2HnCWJNXtXDnE9oyIFQDSQNRMwu4M2op9EGBJ2ovEd4KJcrOe61Og5W9Jnj1Lk5Ge//DJ7Z/QRX
jiM1lZ/g7+8WGE1w6ejiQCupUkTbLmFsYmuq1ZkJ+CS/WJyOXNo7v8jA2PE+bN29LlW7ixCIqw+z
+enNw1TrQUx8ARPt7IBXjSmYmj7jQMzbvNqOSjs0niWoVBhZqTjEM+qH3tcD3CVw07XBBkgNQ48x
P/P7+ISZuO2bvKCLgrenoaIImtKAriUcg9ZEaYOr4e3OvO/u1zSDb0HU06/WBUXflKJfQxyQf5uL
/cVpVqRqNWdK02ajgi8zlCF2fsDLn4ZVDsm1FfNBdS0Nr3loac9m3/SoH9d0ZDd5zesXGyXx5EpH
mNymORXcanGqmjG9GZRiiYe5SLTzkgLFFYhhk826IIk5WOIot/qhXPaPEAABylWbwr4K4s+xXCaT
47JfoWvgr8BjT9ABSUEMvcaqZbCTAnDJayqp8JKD8Eo2U8WcCFP6GwIbzyJd4A6AUYMnyMPsGjGy
JO5mdvyhyfN3TIbqgaWSbp43PW5xywn7BplppBZrjiwZRjlfiSXwp7Bb4dZ/FYEgqQ3+PgcDPqPt
2j3OMm19yl/nAExzxFaMCj90LfMQ8PNlSDH2Eyg4yDeXbKlr8Osi1u0zMpAw2YTbRc0QJ8xskb/i
vZgu9vt0VMIkh8tfNhTbgeVzUyE+cd+bUcyHhaRlfhMG6i7rxkfdqySJxmmT5mOCWd5OnNPsH26+
7605/j+ffRntrWRsMUO+wpeOyL2++Oa6yMSZJFptregYL3AyypDHKZt5K+up1l4hXNbQya6ZB1t7
swFb/PIIqXc/TKYmOwnRsZcQDB0c6/IWQg95ft6uIsQVLnxPGxSdt3oZe6N0LzEB7Bh5MX6/Bg05
sx5LLzTP5F6Wowi4Rlxqfu114T7xR145hZr2OTAL15yS3TrL/74mzY8+DnaUCKJhunmLVqZZpcYo
O9M3FoctuV7Th2/ZlxUxpYhUG2+U79vJch+CQkCoWRfDG51G36a59U6a9mhZmtX6SKSnia4T7zuj
Q6Hmo4qD7lBwHh/8tpXkpYJBTDguxcjZRzV8mRDUggOnmV5q3ENYRGIC+fRnaxy+6Iy9k17Y7f9V
is/8VUW6AAI5c/+UIUpb7UeIbg1iyN2DNZrJmzhbUrsvwAyuu5QnweJrKmptlVwFCezFyEuwaBz0
vCgNDwbHdtJSe4hf5Z6pY7F3vd9vakXxO2nI4E+dxD+4np3U5Yb5E0+luqmFM8S7c2rjuXaJZ5Zd
zKcotIjnYY2tW9V8SDQsSv/MOHceNqjfPPKnZLg8E2th1FKmPOwjrjX3GwiGFTXJQBPSyisCNu9U
XpESKz5EbyGZ7U3xI6+8jDzxCZBCcoCcOjcMk+OZZbEl6S5c9A3oAea0LvtDvt2p3ixZI8N6DRcC
Tlh0+x6WvLu65TUMOJX3P2y2y+HbIKxaxe6LEPzAUlMvZ6JRRCn9zM6BkOiRaJdI9vsAV/MZ0qMf
pxKUcyU8bExLDiSt5R8wP9CqCP13l9xF9G4EfZ8w3c1E8dKyUv5uAk9COvKS07Kh3qaAqHoSPF5S
5kHXDzrHYFLvbFko5h5BBJR/J4NxTrFdAcEel3k/VUVBtHJ89wSZcLv1K5mDKjsCaQza3UcSPPJ+
wi5fZ3w8DQY1HrboII/oJTZW3hsWGtI6K9b/zHQHGbUV+8Wo2KjxrKtLM+IyWCoajIMxQ+aWc8aR
f0GP7KxagEJZmIGsK1ivPXtHPnWP6zrrt4gSEh6E2ENlVr65z9p1TopHk1XJY1gNsmJc1FSX5cOK
hAhhc4TCHcpj38j3py/DcpCyyE1MXx7IKiqNmbVTPmFynhjZu9Gog8cKzGMsnGQpL5m+kktw3yWK
IQG5GCBL2Fdy6TGs8viKrwBPnGpMCJiEqLeZBdt/sgtdT187ow7hd1x3qReoudTsMy98o/gYq9m0
j+P5PPhkZ6z8u3+AX++BtamyMN1eo56dZrL2X3FJmqDpFv87JbjoTSyazY7bWSDw+BbUbqaCdKaD
1VyN/Ey0P4C0cbVrXTyRwWzcaxgo9ykJYsHvCdrXNV4qiIwf8/w1T5I/LOGehuJphOBiC1GUWvz/
SGgOwPhtamQghcwm2dOQYzPRaxGxnK0yFd1OfXLGsJHEEJt20KqdzolP+tGI8xBLvlu9wcgbINEd
GECEKaPTWXdJtwV4FOb5TeXUENstCgcpIQLSXc7NGzD+bV9WQxsfluYxNLVD/+wKzpgRQtaMbK3H
mxGQzE/rSGqkJktarfMtNl15MXqwP5GXQrWup5/CUUFgBNYzfwYsH9DOkNnZ4FVOLI6TB+aAxkSw
VLD1e6YwekbUWMDnqkNwUu60u0qZo5xQ62JeEQ7ZQ9iW8PZil13ik6hEZmtBCNtJsPc9rwdb+dQN
0Bp0SaBnRJvysOZNo22xeFZcjT61Dvjnn4AmGLWm2Ih4Pqc/tUNZ+qvJROnWNMeyHHn+TUw0Y2Bu
7BQ5n3roU5qZIRy1iWvtvPMXFr1T2E9/SbL2d4SecABXzy8VbPJRvC1grlLOpsqybjh2oamOL5/2
1BpKO/NMfw5qxwAiialbnKI9Z14TST73ierDHe63xBBLAyAGWjHpbrTE52YfAUOk+jUTDzwrmXpN
vIOPQSSydG21R304CrkXrPvmj3cNJm4ooLCBW8cqXDJNJu+cB/lz/esWDreMWv5KDDV4ZIGUzSam
guswAQq2VdKQAfa9Rpq1utGpoMeVsLSbzphcSbB3fhpMOvvbf7YlukaScXyFMjN9tHwEHm1nR9Q0
eVmTCdTrXPkVbbVlyMXJbl5ypzsauY1hTP/OFb4H64dwxs9qND9/MPS0gN0Mjutl8ECR0s/wgVt6
9LhaIThG0/nlDc37iHEMIGkCKt75GuLIuNBWMI1CQYaFUlUMmFyQczqQRH0VfryDe1i3mZcfAFHP
sKT5vS89nlQ4hu9/8ti2FZysO9pcld7VRvkjR7r7ADuPuCsb91OO75F9HIkql+td+1RcYu0nuB1F
6F0/zuHHAikL6Na1hrgj7iwNPouY95M0CLz4ZbXMmXUwhVV8fi59J0f3hbNFvrep8bWw8sefEzNB
SuFQ1uMGY6Dl+P/THLjgcZm2qYAAAjiSDh6IuarJ6RicPkYJE4V900nvn9RmOa/rrCx79utR1xEJ
xIJToppiMVEhvB+hBDnAqxYllBzsniOCzEolKUyzKA1F/S2vD9hP1SctzaXR9GXIGVUN5cU191pt
HVPviNqKQFq0bcHFfyowcVjNszTXx3LXBtZy7jq+D9j8UFy308UI34QcTaE55HQ6rqxpNQifjob/
0zqdpByrhLRDBKBJm5BoqdOaL0ztJrpd+eByvKI/+ncpd8ms1rggbLNMOABiA0gfG5zh+yeAkzz+
pYPfTWZIpAa5h/y87Izq2DzDGP+Zu9hfQs7gbf9GPlbTyR3FJzP2jH8aod0erkgDShh3AaFPXO/3
fTwc+RfKuOu1pSle/Ep+kndDmlGQxEUySjUzRZI/oPBkYk6cPjBBR/glrLyFhLDEwci8zOV96cf1
Zx5JNGb/9FKevpOWsaQPgKewvSq03Q3kfVujhC2mm7nDjgZk6vdWA1jQ4fmAsrI8dx3ujGAU9G5L
57W8ztHdMbqo8L1+RNHnG4KNAypAiGerIgUrIOyTkXisecV5DpRAuxb6ZkHZ/FWilvCaKiudA13f
9g73PZbHroMXnYUq5ziUgwMqYZmndOxQmIoIzTHky+bc2IBP7TcfRhzfp8PFET/e5SQg2XQGP9SF
DDF0ssnjdub4m4YAEJFmq+ZeTOJ1eRTieP/I+dZOho025kmvJk87K9coQ3H7bCQ9r1hK63GyVkmb
s9XbiaAkP+8VoXKBr360uhahPwj/idnBtZVXTb8TgKuJs3hTHdEOd+LVuxCCBTmcPXz4FslOITFC
2X2TxE0Tts6JElLZB0umeqjSvGs4CadRF8rbLcJrRGhKdcnP5+rLmsxR3Kywnppm6hjvcewpUQ4U
UmRPKKrmdhV5rsFIUo5tso2cLjN2uYXPNm8bJIHXP0iSqD/GTVCjTFMSFqy4QE/MWGONJdsjeaPx
K2LStAiecgUdHUcPplf4TpGmXIhh1pD1zLI3HfL29VWezXEGNwCpkxwxGOsaAgw1AVmR94kPoN6G
Ea+xoXB2jqfn3L3pG2HvgVyChFCF44JvkDIddBkAptr7ExGM0XhANQqFXjffY+SAq8x0batZneqG
ojqquXg6LY8AGIs4HXM1IljtzfVLh4BYfI664WM8bUAmN9nUTLbW4f+amlB41UDKKS0kQxwTuqkS
2Tm9g6XRt3/+DPMKd7cOPyt81dZGGhdmFzJ4taP4SIXhTDelSt99E4VJSLPjVYCqSIRmVb5WmZWI
+5uO5A6Mcxlz5tFT2XsRZmY8DauabUbZbAGncx3bDVo40MqZjPB5UY78RFWm3J6Ma/lo76MaT4Mk
LKnj89H9OQG4lxJYuPeDn1lfhyP0R0BQ5ajVpjCl0J3w8WcSYLEYIGNY+SjOSyvKOCRHkbUi3k3d
eAzTRiU9EOgDwtZLlswBBpFYd64odbN2XjfwedUgzRTeAAAgitfAccGwvYMHzrVq8BkZ3lD0kj6x
SpHXn0wUG5TuAOhb2jSpuz8l3B+PzZI8lD2Dd2w2CANHF64EzsvmTzId34nGk2cRqyOuVVsd2usx
3+vlzzqKl3x7ioJNwHJRH3N0qATF578nrTzGg3lq3JHphUW9c6h+EjObLFlE3soqiNCXae0pghVz
AN+7nzGxmdJyW3kAvlW/g/8uNtRybZDuhFuG9CBpAn1tJqy2kFzIXaA7w3Zsq16+RKSSn5pFlG5u
ahz+C279CjADdXuED3X8oodMm+XICLu+ZgMeRTfLB+r69AqOy+u5wSVEhUoqpBppqnznzZCfCaPH
izSW4HV/YoA54TJLl/WSTosjw3a6PL1Khpw8Zuld05T57Z2ZvZwU7SCmgh8wo43gTS1m1YA5+GMR
+W81N7MfOEAM5kOfL3XPQm8Y9aeDhrgL+r1UMcwlWmf2YJqzLkWbtHgHNFUVAOen1kYgRwG4AXTE
nlhE/1rmzckVRxCfbXXiAP5pHVsKqskTnhXkLsAkegGxSqxyp6ejL1WDXr54naPgz1PveAV5xJPO
XDuuMBwRB4RLqQ6+NJIR10OhOgZSdJzh68gRRMXsuHnNj7Pjy1a6iyShbufYJsMnIhW8j2q2FFj/
Ai/O36vadfbD2NvPkrspRZiLxEsJRptOFXwOI0zukSo2Yby/fpOBO5CAiQoIDLjLBk/XAJaPpJXp
lBhoFWi6/injNLbsRlzJAQRlvuLdxJHgbu5syCFxuINofWFb0bdFdqWwntH7A/tqVQJ+zgRXRJQq
P7HnApC5TPVE9BmMEksWx3F/1c+v94lm94I7WriA4wwoOWuRK0Hhi7nJ2SI9mHUiowe6SzU4m/OF
c28q0QyVXn9matIe6lhQE4vidH7freL39ZBhSmNaKp4In0y7vQG4XUYcSXtbXcnYx1IyYNLwmQAg
7DkcjWxztugr41yJCsf/SLPXMUF8j3bxw7zw9OneprjEsIx4unD0EpPEyU9SrbOWMb43YNy4/ciA
cJXQG+ty3kBL4gN2IR7C/M3HQcmi4K/HvrnBewnAcKUsmBoItbc89qc2cOu43Q+s72z8fk0AhNeg
uVfZsU7cAl/W0mJpuhJ7qad18bDqSQwf39EiUWw2tfpkJpiZgf1UyXcK/AeOceHJyf6RMoMPhtFw
Zl0V/TxbKMSFUUL/1mML0/wcc+uhD97vdbErX53sLPotPsSQSS1j2Ha+w33u6xXnHNWHF5NdCeEX
QnDqJkrw+1vD/DDzmHXPLe1rmIsvm7zjqiAsDnrSHnU4NPg1w65yjdNUiBwa4oTx7vbdc9YKMf0R
S3R/x4lMjLIpc4ahZny+WfH7RMYDMACblN0sB1kjTuKz7yn9s57mvgmKgO/TstM20qtzLrhd9vb8
mDnRYTmj35VFJZUqSXCB0ugFivPKZYwtwXkwfo5eSDlvO52wu1BsD80PV0VPAgmgB7nwF2cGzY90
KmsFP0J7GYDfV07gnOCtQLKv52zGb3R+hEgzYEgIq0h8ZzhAlp07xqV1LsXAD/ZmhAPylZnQTsoo
XtCkcwfyKgmocO1kQOylXWYyhDlj65J9apKxCHE9pl+oK/HASRADJACQjba2ECZ4N31GUmin1MU/
yTMTjZej2OZ1Ef66zpi4ZaAZjN6pEfHJvDWiJshq6fOgCgJmaafN8WV0g2/+RunkcuBboXr8JHBS
IIuuXk2PQO8GpJONsvPOrjtnCBSB9K0uvC6yxBT8FmVFzxetnH4oAIsnKwh4OXYv4XjJx81218P7
VtH9beEUL8gd2BiaPw9odltujwsysZzDGF8tzArZTXmNgumpH3cZfwruYtzz+VrnVbKCx1SlP4Fo
basZ2NtZZvydzJPULCl318Pzz1LM+pGDhVx4W7XjVhCsWYE8d3q4Bb1j1j4Ns0OvZgWLgdMf1+18
KBOo38vx0dg/6+IIqL5633GLIJmc/1Cya2+ANvLWtm6OcwSTnspZf2usgtu9jabQwni8F0s2TOsF
U+VLHH/wsyWK6iZsHb5DobJ1EhC7Dv43lBGiyUDSCGwcTo6sgcGamnY+JQqsc9lYxK/1lbd3xgM3
5KAPNRol89n0XD6dzviF25hac+d9ezBlT0W2QGDUZITtdKI+Hw3Oa3YA91Qx5OITFIFYD483REv1
jSHyuNh5tZuQdc6qu0BCQdeU4FnYHqiWwuuo2zEmDo/Tlyv76JzSH9ezTJEqv6lXH5Udsq3bVG5c
HPSNDR0BWqU1yJ5Pl5rNuEJ2c2iGJ38mypZD0DtxcmPZnWnI1wQubQds1hs2otxA9RaLL/J3X3Z8
vs4i6aKM677s/SMVehfOj0uTc98xvT67tHbdiaI4TNnVdq8rFiqguW4P+LOG1WiE4vQ2zLfbZLqM
pAIqQmPnbWeE8Y+9m/CeNRGille1112PTiR+Fp3kWoNyH3ogD7SstPE55zfhJtqBhcvW1NKy/r+6
4NNAcIADHa5KQRBeU3AwtOZ5LgxyPyXXZrmuUTz1iUS98T1FzyGvOGHacYhhnxwYmJdHZ1SrLXAw
pcBw+BVjA1sTu9mlc7OjIZzWSqvkMSUKhxCaV/yUxU9jEqwiNv3XPq/SYvsar793zER1z4YszCzv
Ia/rfqqKSQZnkEboZt9jZQHQBsgnMjF/J1xNfMcigF8OOU3G8HpKSyZpgI3qb5PKKdyofpxRQa8B
DynFrJ53IC9ka3ENAwvAIiOKMVEHfvBGFssCPN3IomCcoWLdmLQvztM/V67e8gEic8frqNBk2Ol9
sBHDz/E+PnKlCsiPB5fZEgIanZhAZnQWQvjnPQluelBedZzWMnIK3674QW5J6ghK7dKSiyomspQL
CLPedNUc8L7RcRQ5GoO69kNDMPPosigF29FmSmYPH+1l2V823GkgaehAsHni5tZ2BMaCvGH5U9aJ
8jGDdtuuZaxNZ7A5Eco31Ss0Mi94VfVDxO30EQvUet4kSXdMiRapUZXSTEU+JaPClqZ/8MEGsJtk
vn7Q0w3f9yD9DRojd6hafFOdOzqGvynPFHPWF/Q+5TVrzkHw9/ySfGwwWhHfvsf8eG0pIu4YJnSA
qCUeH/CBcSP/QtH64soX9Ytx/WLoFulragM8zrp/XWv21hn78DEfhO7PhQhiSh6leCgniwZCgc4f
QBsif6qCYdgdk31GCVh+gywXUWFn7XW5lkdlIK6dre6D8p+2kdfPX2oHDoe5gSGq1eMcyAESDId6
MCmAcr1z9zyaK2Vz2gbmalbj0UojXZp2zkiRkAJXQAtKLtGqj2ZUKmsfeS3zNeQ+ODbl3i5u83Q7
GJiZmuGP2SCUW1PlzpVyh8AsG5gFeW4B8/cESzS7TfJpKLKg1EkCxIk50hgUguK3kNDXhSadLk9e
8pVZ8C/aLB2kbqNk0ZDsJ8jg2eqwKXJWMcsP1YoKdKNwTj462aL0/l958HzPZhVnpIkaOwcrulIQ
RF0fAcuweeG8YQBH/S4Pst8wQOnsINaN71YcLOOM9o5oTq40Qv51gkbWmXI6Y4lMdPrt+NLWS2T/
ANoALte4bLNzeS5L8igXaQXKB5PGW/+SwISbXnvdjbBARto73QzKzv9ihS8spa09mmQFdCqseJok
lrRJ6WYG0emFz8Sh1SdRgmQDSADoynEtC9e7qIyNbCaAFbsMhktfE/ysFKFV+jPO24ulS1T6Cy0h
G8kELwEgjkuHqOAG3o9j3XW6IG1ATLnS3sKlV3cZHX9MpPXZDMbP2D0FfFnCdTJZ1nMr0Crm/m6b
nGAvkTWAxk+nhbmFwd17z92n7cd2UVbDoHpIF2RDHVMkaWbcLZWPa35jmYrTXbWBce6OOJz2hWpv
gVUgpJw9czqXWP2BMskAPJ5lIk2Cgh8TO+rY137kQjWp5NLRk1kq1lPYA03HkNmKRaITqiTWI7uc
caoOjy7VK5sroxuzr+/nCh20qNgJPw124vYPL52QUZ2HEbj27T0qRsh8GbgI8FW44NSSkoY32x0O
d7sqJwlHLiLsLlouN6K1IeBM2fxmb3IArWCXrL4nr64h7WmKwxysoj9xg1bMtLt4i/DOlHjskgcY
QPsO/d9mq3wrOoZBM4iQ9lsp2yJnufoQ/nPTUuf+WNRcvTuWNWwQVrM1kCAiis/9IWvClhRohUiQ
m8oUmLrQ3pFof041mNbHzsJBano13vecMDaNBG/0YETirIJZWnFajJRdc7yF2S4WAZVjhSJRbsDV
QyepFxTfEBH41Ek6c7AhrttoqsxrXMe9V71j+M5w7+r0z3bi2+KHnjz8PE4mXzTW+VBFr60QrT+C
e0ldL0JnL1UtCg9hNe/mkhZN2L7fw+6+WCPMrHg63SNaO3Ge7O7e2KJuPrhiP8SzZarIGL4cUJkr
ldCqs0hDGxtTi7WudeTlKsVpj5FIfxA6XqEk40KowABHGkMoO8DIG8cOKLr6Nrov2cnTdWQn4AVE
yDCMlnKxLmd/LbdsUXyOY73G3Qds582+aZoEr0jbSm1CNL3VG0PULol2sVAetKAsd0FYC+MEKjf2
SWUlJoSojmETwOnMzGqBIALGtRUw43Yi2ZI/Ogc1quQ9Bky1cOmenQO+cPYAEq6sDBB6KZKuz7cS
h+Y1gdlHqoMinvneQAgLOFkHJfGZFGXS4DvIvPiQ09DhFvCJdRrZuASc+DhM1KlppD+qaYseetct
wcLI4QP4BTnVbbhmlYHEN+xYKAtH1ZDuINUjdfLC5BJ+LFcOq4O9cbLEuFV8fliA8bv4XRMsb2EH
X/ggONUOpx/mHGRpex36yyZsoi2JeJB61ts7nndMhiMxAQWG/LatvvSzPyc0av3ActI4gcrmE0Mj
EXRUxWsmJaCDHcCq82ZV5TyKvzUHGovxnvY5aE8r37EIOK+fTdAU7+5jQuuJo27rkEtYXBVCYKRb
q84BOEPJcXT2vq0EJyFkhhFrtgsoP8B+Bjn+Q4G+7v4r+JtocBX8Mcxg5G8LhbVlNsAdwXFtiG6D
m+xINFYLX/ZBf1Bi16smSOnZwQrW6OSwtKA+9qxMp3qjUtHTGxVKw94QNFNHuE34EWWUGqhyzI0Q
XRvVnSmR3W4Neopn1UoBoWLg8v0fOeFTnRszARDHeX7sVOFuRSfXHfd5Vnc8O7qJxHFRtHcTj27p
iz8SBckbVzqGIun+cAVxvkTN37mkVysD2lwRFLifWD/ZYx8RUKNpcnNyQD3yMnkcJ9wnwP9k3Kfd
H2eSrlJ+jgeaYRUzliqZfT3GQsvH7Lvj2sZRAceqTHuhRac5ZskP6S7PGbRr6fyitqbMKLLM10eC
FX15uguiRfKOKbSLQyaTq5aA6bYFAyduCxCxsxnRrg9seoOtvDH6idHNViCWqNwsBHZb9xSpf2kf
rLddKIcsV3u0TCgtqcOtPfswmFg9M+mjCvaaWzNWgvsz9MvVkV9yvbJtV9lSKMb6PCILRG7HOJkn
uCnyOxtVnIcl76LsiAcLM4EQhqP6Sq/TZp3wULO6njHxS8qSgP012CK1Hx39z3lR9atVbI3wwKDE
rHHvBXvKi2uE6pBjERtRLww5mG/ex3lEei4lIK38k/PFGeRBU5EjGhvR99YajD6uQBEQ7UNw+7nE
ZCm6paT8aEWsUbtHrMDDOMAKmAOp8flllHViQXgJd/zaQt1k3XkuM3Ppi13RdpOpKWpI6LAzXNTv
AEZ3T0oqWlp3G32jg8E4GuVfZ84tYwZbwKBNjWDMRUOE15a3CNAvYTrJA0ZByXoJ0gs50eoF0Gn3
hXspB8wKlw9yqZtrqnvP/A0My8kkFMpxpiRsz7IrMmNEwU6ZArIeGcrPxeTSaosNJbt99TdRixTz
o4a/1KfVVlWDhp+sZHvMi6QEyzuQ7wqS+CIWJFJ7ZeygEaJ301EoB+wITBpNBwwe8XqFe5M98cM1
e8zDj4l/vnpUBkVunR00nuoORhovGKwfNN0FbxzkTYClfVEqHaxERpc7/fpZA1nqNXo1k1QG2XKZ
Lbxm0n+/B6KRAHy/DgXqRr5ZqF7eda0ShrBtYBA3SI+PFddNXvnjok7fgxoLREhok4NQDMhQTi+A
OR9KHLI+6BH7fzBTtQh8KnDcfkBReoGUWWHZrdHVJVJ7aGnTB1wZIm/eWfrBSbOb6Aa6KyQ/p1mS
KG3gMhdtXaDZEO7DtYHVtXLcOQL3W4AlpbbBYdVjWVDHx8dYG1Sg3sLIhof9lPxHzUhK7dmRokJy
MaPZ1Pm2gazFEmKPi/+idQAx2Z4bO/3uoJ4qmLkmvvWyr3B4PUEc4injYk+S89LLJubAjozN1DdD
MPNVADiyBjmVYh153KpJ4FsgzxFsigVaEHPawJQpcOBuDs3WoC7NzRZLRf2SK2NYfuHzMCcv0PUo
IWHga2jJN9OhcMz1Vx0TdE4sltNksO7frdIov0Iv6XIz2oj+UFP4tbNiULoLCJ54QtLiuH8aIOPj
AQFd19s/0DQf+KdN47IKF8679wtUuKPveKPfqorvyKFPRCgA9cWzH7sYnCdVyuX8SeWXKgH8KQsu
fuZwSfSv9EmJ2V8p7hFgRmvbGIscTsjz1dD3Op6NEyFjENxhfo5dPHnghcyTQFSAqIdO3q6ovC51
dtApXp7eI2aXWZZZtN72SldOWmARBWslU0i5lDKYDr7BaAG5E9VwbfK04Bbsz2bcG6ho/AXbqwvW
ueVwPWfnBMKvrSuEqmK8zqWJZeSx9q7IqrMYyT87//+4vwJ9FSPGMczzJFm2T0qktQESSQsvQ6e+
Z4p8/Wa+upC2TnXorfG1mEoYxZ5P51F3fP/gVImC7lX/7pGmALTGmGwnRxG+2DKPpZeG70hs3mbG
sscjXxsWJztmNsx1mskGtsPUeBaCmR/f4HxYE5NK50xczsVZjpN//6VeJHFe1uLhpeocuLlM1Pv4
xwFHQdaoAT2RYf4jQTMIK0yWntCaZAPbQDiwYbvYy/6MuyHXLk+nbyLzTIMUBKktbU08IZAJFE93
cB3+n1FjL/zeJ6k0SxFRUN1MXEq18m11eQyQ+DLaNRPBPVsatL/AtwKm+1ERHVCIiCiFpO4irAT3
BcGW0x3Dz4ObFZ7Mb8ADE7z4Zo+fIBInLSVftyE+/O7WGutE0kEAmcNZg0KRjEG0iXAm4dF7SerP
5orfOmniWg8LFE+ZffnhXuyFN3BXraRg9dvTKPyYCsf2aUIZTXpwcJn3uJdjhSeo00XakNsO6T4C
8uHDYo9VPrPktEk4VoXHU0rth3FRg2eOpPneS8aBgZhjXhFTqQDejrYBHAlAGtjaMGbyLdwludo6
hDAD5xG79pSuAMi0rRVQLP5BLNR5GNnk1BaMQVVY8Ql5buhh9LRzQipCUfo7X9OymDyeUF7LmQlk
deBK5WQ2C/HhNJQy875QzxpbrBOc6kFmd9Hy1y0WWi7ahs3uhs+H1mgytIjGul1lJRAWJARMual+
8k7vT6z63ryajHzEpScaKlPnWL+GG4WKVeRrcXpLfwXs7bEujFj1QLetoxKx5p1PCmLa4RZZPO0c
RRl6MtH5vCD1sY7sMzKi2oKe7Ks3YktTgHwtVJXPxX2hcvlJdh1zv2yR1JY1N+rgjaGl2d/bijTC
zH3vWUItNq2iAjBJcaJqq028KcyH6VCC4e+QU9Lgvh5Ag5taNHvLKj4JEyO0mfIWlGNSWeSigH4h
go1AWsx+ttzhJeFddPmxwGUNoBvhdq6rYxxcW9ui/+57sr/E8sB0EYIKTfjamcyGWl4TMrernNHP
3koJU4CTM7fvXaa0m8TTSsmhyt/T1LqaZouj9SUPABWLcD5jEdm8ifXQjI2684CcmKrVZYQyCFIF
M5t9+Eq1YzvRgME8rnRF8QHnxojh+vMxz4NFnmT0uKm6H8ZRBiq7ULMa3Ku8phLdubqtR88OhXQA
bxp5H8v0glP3yCcEDi5ZjMbwQxnqgROkFGzwQ8XdaOcIiFQpRiucGMqc30vmWWxdVo6KDP+JKNoU
AvLdpSqttETj/7ACwJxC+cAwWGZWDRz+mBHjmkQW9LlrE53LESzRGOeqcREOxA9cQTMgqv6u9n1i
vVK06Y0wM9ZfkUQEm4Eu20FFKzHIR/r3b9HtMaQdf9vxcCJwVA6Ych4H8g0OaD3cyPXfwNXqh8m7
M5NOK+xgU64CqLxIxM39kiclClCJGuu/TaRpnvhv9tE6N8rvS+w0PpFbA+QD1+C4SPf8fUH1vrvW
Om0PsjyObbKfx0BeambcCR7puzr4/0PPc/NZRhrDA6XBf9iChND5f4spBSDor7soHJQYnX/tzNgg
FtwT360ejLDZBXmAFBp1Kk+O7r+emocubZWq3SAUTzU+h7ulnu4LAuQlfvqIcfa6T+KA/UCBG4Ee
nQRd5v0ul7hvE+weoXBoYI5Nrna8+/7yybtfYmUDd+AUddIBWe1geutjCSfvx6eNYLH+pwsZLoOk
KVgl+WkacOa/ir1/x0y0z4wjVC4fwU4BA57ummhardOjcKFFKNrUq2xq7KstR4dATp8C12pAWqaY
8alPwf6r7nm6l44/6lfYlq8ZQtHOfQqpnFwLaJh/gvObE+XjNTWvXcCuzDX1DkYi0qf2asFFzMYr
xHW+EVg9D4K6apVeXeSBPyx7KGV4akT46u0Yr/+SxxqcWTvkvpBP5qlssVZEQt8l+pa4Rkjrk3dK
XxsQxoPvJPHnrMGdaoGvuJ7Q6KqnEqUUAzbeZdD5y3XSzwIO0zOe6mlR+UUe69wk6acA582j0617
ZOSVLF4K7TSJ4s2FhAoptgWodKipKH+WLVm1zUxxpvjUZ3Rd7nFOFPxpM2xEV1YITH7oOPBDi+1Y
rztQKR5gdUmdVrZ/UBnC97jX+LGKBge9RaKZYympuO1ArI4okpPNZUAePUh0hxDhenzVl91De7hy
HASDOBGoWpj8ro86HhPMgbWuwQmttOD1IUwK0XlWhcESP43uJ9FSCO3LHT5+AVL7D9WgjunUdJx3
mM0r58SXEiw3U1DZy8idF1q9CcqHt836rA+LASetOSzRr2n2Py7rU9PqRfafGGULJcsYWdiDnzsn
dAm0IqoFMvaLG7DDOc3kRFWbZU/ScHL0BAZ1oQZ7uW+OF5MSEftH0s/u29U+jjB4xFXPKnB7vEG9
3L8DCPSpuAVeRG7ihv5I1nyWFUYT59r/XaJ6mW4i945WvTe2L0Z4rb2BhY084LbQ8AWx1rpFVjAc
LoN9TCRAfoYYVmzN1KopuJyxpZbrd5pl0jRdgCk7lNdPxpDQK8tr4A6KYRN4aSDo7OgCy8HBKl4j
in0wbm+31WkDpaNi9raV+yHmdRGIWawDo9nIGTPp//VwTpgSVVvAxdK0Q3aSRDNj9Mme8O2Q+9mi
uo4dK2bO3aF2hGNLkbWJ7wb/Fj/NyD5a0yU/q9E3VDFuhmpf2xvszJ/OasMeYo7q4gNz6Ua6xyJB
ZsLJrGaf+rTs+9fEtvEBjAaixjVlHL3NwE+kRtyAVMiiF2F5HQ/cywruAg6UeP6EhU0rjEl15Oqc
g97WPSUpdrzAD95h5zKC0hkY/CcibrAw1g4Uu3IMdDZzUt43dQ/oeoUUSYkfsQbhfL3ii9zCu+TN
AnMYs1SujsUYeT2E9VIcG9GuzsQ/2aFlnfgJkUxOezPrFzDOob3T693SFQCU/P/O1a5CFbUqn8pG
HYioy6ALlaBDW+aTAt2JMMntjIWXV9ZREgPMpUWvT3zKFYqIUUv88YkzBSnnc/0xHr0l+KErF3OO
VK0Xtk7Oxu6u5oxSv/G9XdskjE2NiOBbEcMBtmKgMy3JfIennk5dBMd7DMH7hddMHb7x5fVW/thA
CHXY2kbpaaFQyX2V9Mc7TciAvu+2H0dW+2KUfXNz+E65g2snHaxOt9zEC9+B4YDY0DhUAbsbyDVG
xpKwN60hGQx3peaTLASVi5Xu94vBuES605kV/kpSpFcFEsLCrF6RNpYV3vQIa3BIXQi33yOJpxmd
M7Yei9srPLQWBU16M+8crh3wU5V1RMgB0RSANGjKt97ZF4rIToZx7IzIOmd+n6tbdNOCGA5GUVSd
snEi84a6uHTpo42BbyLLQU1sRTea/Z3fZkRQKG3yfh3j1OMY4ld/e3dVdv8up4NBR2iG21IqhADK
t8xuBDKSSomzsLY4/1EOZvl7pSN/6Zt8aN4NqkgP7zsnKHtIeNGxEAGGza+D50rtgj7E062cgx1J
De8HooRzLJxCuC6kpWiSgLOqrk7crRu+1FceOCg6Dj7PdV8xprqAXEVNrP4oNyhvEzHyLIv6GWl8
ulYk6+alcWX5JqZQypSZgdCJa+ylYAZFhzPL1za41yZ5aDevTlWiF6T+48CmO/qfnQ/VL16Z0tkD
B9uK9WTv+HSliOeLkSo48vzz0cgHiUKIC1r8Sxspgdldufcom0l7W46ugFt43MW/hGG60jcEh4Hb
qOqzHjw5m4az0iKgwQj8Dclp2ut7M+Kbtnem1HHWFu3y48DL7MaWOxEXPS905X7LKe5QvJACP21q
yA5oEeh+QpyBwyJBzXxJDdVdmAnC2qTtJS30wxqCqKPgVZNg3nHbTri/+cHJT6uecAUG94INgCXL
RG/rgmNnogPqzGC6jzLXNh+Q9HFk9uGRWe9Tsc+d672wrDTs9BwmgIL+WWpEtfzUNWE27rNPzZ4F
Asr+2PLrPlZLxGrSYicuQgM1QatSBupZ8IHv9eARUIDNxHff8MAH+TcUxy3kKpITnPmRe6JCazd8
R0bBelvazhaSluLM0CcxMGhwv2iaCOEBpUgMGxIofYUYn8n6h4gNzXhqf0ZMxK/Ve29yGHsB0/Hc
RC3SN4GT9mrG0POSMK/Ke05GLuynfvKZWIOJxvfI3ZBiYFsJ/Bl3TT7hSlew5pTQVlYQ4fIrMFgI
rrlTa4rUBC/8+jc/EkjGwaKifyqBL6BUOx201NYPD1EzkC7/zrJTEvhsm2K9g/KX4h5bjz+rp597
eIbvl07Qwzh8mxWu/G/FdHSGxBbMuTLtLjaA9t5WoFmFjlzHigrutenOfzMujNRkKDq9NTFnPjpI
hQ7dzHDYqlS0e4iIQpCdmc8wxSv5ZFKXVMn9MYSqfpra2AxeeruktVTGznQ6eY5eoJPae20oMQ3u
/BMzaYSoMKOjPaz/UskYXwdNwJZOV/pOjBek65o2z2FprvI5PTW0XSY84sgpfCBO69L43eCDRJ0c
6wAuFaZObK3NsS2mtEZb0kzeE9SX/HJreB+ulU8z3HyVGI3beuXfFEcq7WkIVSf5Wl7E86DYUc8X
0tfAiV/VmiTU5K7sdpEFdpNeJDUC+9/pMFellUEjctNO8DyBWI2ip8Z/sMRO1U42IPN84O5bR8im
C3v64sXv2FvjKDGA7Dt2zAr9ZRpHG4Ae2jOcUE/ok9IiJj8chNqLBni835Q3qq2D3JlI9PAa5PT6
0G5aRbUicelQZtYY45gu8pbZHKmkmYZRZGrWcoEyOVsGIJy7BHYmGgeloAY+SPrDpsh5bjIrztJL
8lm9sSh5XinG6e0c2FI+FYMlwruC5eTgK3izrdZbTuMGCQz7PZ+iht/vl6l9/OgzO9SeLuq/5g9t
Ha+sBK4DsMHwHEyNzVMs7nx1gpe6XVRGYIhTUXQm2L6uc7oXas88STzaU/7Djk8HLz4s+NfKQbqn
pgchNNQ2MmYmP/7aH+WgqLaq+PLxFhddXaAF4BaWni7Wg+jdfLheioNH5UxGWmVtNQ5n0d0vs4LP
OeUcfx2dmr1MWx5crKY1zUPPIb+l4R2JGusQlTnRBRkEtJS2SOEt1OGmt+jQ8kmEXlv7liMDgnPO
EHnSa8t6vEpeVzR/NLa6aL4iLGHIdVBWuODEKueNkSQZeNJ1rn8fam02w9duZQhG+BTXDEO5VVKa
HZvfHBNaTUTSM+lGNWJcPCQ8Um4Tk1hY50SUsnPruQdXa1VMIfG+wmyAFRFoytDVA7XBUBIzlIKm
3ce1Q3PeHUz0YO6OE8qBUwbm4KCGKSY6tHdhMgqLYRQOzemIu3w4VQT9MpCxaOqonEhAU0/xrOXZ
OCVPUHcJJ1oGsYFZQpj918mMtVglZFO+rbVxRQnJgZLf+7Z+aE0li+7ojGsVY68y588T3Vv5N95g
dRWJB+ro+JxOKyu94sHORmmnnyZpnlerRiJaGUKZNHY39F1EvQCfyHGfYM986P17I8/gBIMD+WQI
Otz1tP4pIkH+ifBve52bWiOyL1v+2O7NlueYgG6B4hRmOQ3gtUVk8Pd1JtVwjODKeRHcFhsUWkbM
olCqJy8/hr0OrihkObpVUBHK8xg730iacJ4j3qn+ayJ8zot2j4lfr8KHSwy9MQQyygHO4y+Q2ijy
3Aks0C/yrvuM0pnXzKTxZFCVdPSqnouoK0rSlV+Yb2HbNDfItJS8MxygO+0oDIsi1RZiXIfONZEk
ppCL8q9IkktqV8qLvFq+ul48LtlalxSjp1J8OB5B3mRvew79PSsVwCwWtskNWNKZsJ8m2S/T6lKF
QcMwimN1V+yLLF72wf4pWSiTMla76iPnKUk1DxsBkKPaSpK8tnoBtim2gSQNencL3e15SZoyQDXr
D4R8Ptr5MPsn2dhFr/I6fLxYJ2Db4jvUO0+bsQ6GtCgIpV+WnYp+VMV/vTeFdhZcl0Gq4Af2jt2B
RAr7w0cxrxpOoBng4aY4K+l2kFoz5YAyBG1/VVwY+dZszdu1drelkPmb+meO6dTJyUivNizYthWX
14Uvm8VILctzLNmOnn0qYdlL8w9wjsxtSi/5/wpgVB/flNd2WzY/GyrgCc+Hgj4A7iT5n2FNziQq
bi5F5h8hnWUckYLyJl9BIpkU34suAGu2M8HoS94XjJs6MGBaKyZxwe7+ZLdlKWkDQIuIGK8kIDH1
5D/HfdJcIrglpXQDKP1kO6ps8UsZglm9Y7w3ADGPdxmves1it/x86sB4rmOUTnCKX3UJDxDcIEJ5
gvsZ72bOAeIQIqOv5gUN6SlB5ycRSVJa+F+OVxavgZmS2qTjcnq5Gy40uYMM8WpI3q2ggkCzNR38
3Tb9sX3C24o+SC1/BrddKxOp7OwGqKtDNhicuP4WBMiLRdNAOQrkwNDNDwL7G6WxpnvFCZJA6qH1
1V/EGBb81Kb/ahahsfp3iXzkoDl02Cod/jeLwABzaXEB2wjFgIEEIapt8/ED9rlg8uMxHs/U3HYu
XRHXZFqJra7f6moUKdtXgDTHJnRam+6Pu3VAILpCEbnEO5+T6Y4QRyHFkr9HO425rfaeQAaehQbn
yNeaiv1NfgGv+Kkug9pJHY1CDr/jflQ4tTzGdolXWuPX+ipipFMzxD6pHf9oOLA6aL8LbU2W7PET
45d5xctlNLkmGkwqYLxNzjOHfuaIdEUgqyl2Vg2BMeurBuPeeFR+RjwPFW+xnrsJmsG/ahoCAVa/
n7mUNRhE1jg+3wV3KLoDhkvkUkvQizePmZ15Mte3tFChaUMEweom071RBW8RIoQFZSqfD7s325tA
S2KeO5k2XZkQFeYQ5NsPLMktCY7UclCdaeCV7lsAIEZvxIynL1oUehQHixRFLciw6cL9OjVfldeo
9s4K5niuxKTDdRogotbm4OCtzCpbUTsaCdrEAlBAGkTib94Qi5yQfRoWCa2/qt3sjCUJUPC9+tpo
QNMoahykO+CUMiFndzHCNGqF9Fyf2V2ml5EFGTyynU1t6zzisAXKAJehJg+J715oGXDG7nY6+72M
sUkB2Ubbf/HpDxhUpRQ32HFUuBC17nsY3Ywdq5nvpPkqy7tfqEdFwBO8uiV7zTFi75D0Myq7EzOV
lDUkUztwxljoTfb4AC4dKoqNgAmwgwWNVJsAWCGsC9fSFRCp+5mzClSldM9ZPybR/BErDHi9GrKT
2eUrgYCM/Og9DoEuzAMcM6ivAwXD7HSgDGPNpzOGKsD27r0hNtXVK1uWHYXjFhnQFW/AgaqMEcOF
fvAeNYiPiVTn9gJC5NcUO5ckqXUpOLfwuM6Gxd4NPCmllH70siHWCzV6Q182GK45Oe0i06wAKh19
rQ0F4GBXmTdCPvC+LHDfW7EMuYkYzrGrqyG+jkwD7nJUpFWFG2/4Y/6NroCwDb1LjuQJFWiGoCyL
dxGXDzq+1Ff2ZfpotJ8AqyNOrnb/i7UsgQVmPDVvbUj89+bvN+prfc/CG6FBrDScwOZ4HJwFHj/D
vrfx05pL0vobTlTvx7EBFtDLUHoGKqIaQWENz7hec1qYUe/1IQidxcnw3O6owiQsMJz3JeRgN2Sc
0jZxhsf9RPlU/3QCFZs0Ks51SE/0dlN54OCE3NebHGkv+KYglCynaGPqas7acK7DdDhTXRT3iiIL
7w9n44bdTI3oBpvN42KzoP7Dht+ZpiGKAhEsNH91jOK8X5JHtA2qWsJ2Q38kej5xwfE0anOBWBN8
pGTs45j9g2u0wcyy9yMd2uAtrx+ckzoQ+k+Gavhb1/AO1lvuM7xmpmLo28uPLE0JmypvLCA3a9lc
QJA6ElUcIe1mtg+MakNUq/l4sVch5o34UX4+kfzogTAS1ofM4be0TZ5gSE9cRWtrevqR4TPKuu7R
s0FhXwF5LEjWLwJQtpzBxtxLdlVwNDaGPN2B47St/083dm9DEpvh1VIwHWvejT8whGEd+KpM3ivw
lJnR0LiU+P2bN+pkkkqfJbUZcgT95G2rEOsIVMJhUlT+Drm6JeZSyg/WyMI2xu8h2YUZ0b2UswKX
EEceaGBQ4ysZaWJSNbTTOT2CVRGyDmnh8McYPRcWXhfDnukVBWdPcxzSQqnMz1jjHqpxcRMy6hoQ
JIkQA8AKrEv28MB5XYvwAzKq0HaAjgSWp7avUpUwFb/2/OQbkhsq/chGCGVqksqgEHTE8nn23P6P
PgnVbjI9sg0UjoqfYCM5ZXEx42tqSq7MixWIE6pLNqt0V5g7/1+IEhwR8HIt6MlqzPKtdAVGORsf
2SJsKk0PEDvMLSyX6nfCxAHGt4g0eOBRBmg3QF6NdNPA/8yE8zeo8BVZe6Lh6Xbk0wdjejGFWz5F
RsERZPMjbcSi9culAiEdqCHb97GKfvGZtB6MBQ7TxjbqTo874qNuFcFkDjhbuXcAeNkzQkEI9aGz
3LG5LhFUT8LR4fIWXhy+3+eijSnTs06JVEZ9aH5pYMkmNoxIvhE8q7DWIGpn2IBbOYe9CWMsw6dg
lBLpM2B/TygVQzFmaPTrSjynF7oH9cOYpbnNP3zskcqwrv2aAM33uywhokP/STdiC2DnK/Z3owx8
1Ulwnu315arEIqqzWGpSL693Q4MHvJ6IHlJVanfMcQFEqqWmStnJFo+jsSl/DNJpdoSSjD5ssexu
kVTMmbjorqCBNiEypYnsg8Ts9krA3vJwcaog97qOIlM2tO2J8/ue+YNL0Ucof8GBT+GDnF6nUUR1
vQ8mzYKzIB6lJJzOuFxm/OUsGJyMfRy4MILZRH/ARoTSFZYIDH4Pa9DNrZ/9bQ5qlyoDTOtRNiuw
ZEQKNJ5bO3uAd9H0ogbpryaZbNcYyYlehTJSgo+jVsdY7q+0X/4key248XEKlpG28F2NRqHf+RZ4
qRFmTfIck8e0AxowUm5GGjxh1WCQKXEXlcjCjawJEew5kwCxG+2uwOTiRzZFYoYNHhSABjMR5dMM
ZX/qIAqwxsUVmj2uOqZWjoxTuEjLjC2iF4FYWuuB0d/GVU7246oZt+7BcYF251uBrRJ7Hjtduu8v
4U/mflup3b/KeXhZBl21Y0iSxsm/aZxTAEMmj22WfBWmR1hbaSUg8aSCMuZYJQZSCQJX3MhPoz3C
Ga38HXMcluPDJ05yBmSwcM8S2FwHV3fIHtzjd8swu+wYM9QVtMOjH3vEvA3P3pcTKqzcZb4+b9dO
xgfQsJ7/7CYkCsBhGRT0Fi7xEk1uU8jyh+G3T9PAE4+vYEqCAwrPpnpED6MzUdzG23Udxv0S6kiu
sPS50OJFS00eBmkNU09rxtNJh4gDQfU8PmgXCf5HtHjWOAegwITM4XN93/fbl0E6YPRsRMaDXt/2
+s4hBgmgYBLyfFJryKRr0CAtR0h8Pkyo4CzzZ8VpYpum7QNOWE8Nrb2bYB7iiIuV5imOerQ97h+h
xHB5b5w+Bzm4kLjZDNm1e1Lj2kFqKQYF4rwOkmyESeSUEmdnxofQbNx8/ZdQEB/xadRUlzNeswz7
2sWbyLyeu+kpHTYiI5LYV3gyoOe1dXJvzbNCl7tirwiKNOVC6nyw4iYb6ylS6nb+Xc51NQZKpkXU
pDeoUgrz/BM/9aAuOGixxrrSwb+4qJlfQWfakG6B2QRZW4d9L6Mv9S0CWehmfzZ/JdjF87N97mW/
uuHUF6arCQM5cvqx++H6Wr/2xv9b4bg+kXwOfdDFdV7crNNnawzMvf6gZ5Rj2xUyCUsHx5RfT/Pt
urBtSVlSAVefCVC1PEuFK9CLrAu76+oT7EVbG23rcDcPs4Pw91cF2LGlMG+oWGgC38XomY9Ojd9h
gOHsFBEayajnIFYUXwdxPDGjBZbidj8tZfl3E3nlPDwEc1dqKqVMQrSjT4vO1xwsP4l32XSLTto1
uxBSIevGNbBeLESGAlukqTHcZJsHGSYpjR54raKbEN8JqKOAF2iALuZrQ10ZiEjjyQ1SEJL0E+U6
V7uva5CBm/LKVmffO/MKI8033pU3Cg67njaF94qrDj7pINgsVJZQ9xwsOqMCkgjCCMbomVDJcDD8
ykkqbRC+ZcWlspMre+yIQLOz0PW1x7UB48k1wzm6hJrKEdkmM6Q0PIw14R24nUC1IaJcblI0BYuN
H/hdfyaGwHFrAWCehvn8xxbN67gcdYYW/W2s1iG/C0unRwKm4GWKhQycw1HEi/kNVDnRxW2oZ0UY
RLiIQ4cqt+uvjgK3vj5Wz0bmSVCJ6fxxyvjCjF2nVXYbf4F1C66ZMfP7/0k/fdPt3gIfJ/kjqrLN
wx0hhN8DCS+JGictYzxr4yCuJPFLtv+uw2+Pt+lSp3KdscETKwcov8MOHlwG8Iun669vdfaVqDTH
HyNdOx2VZPZ3V/daygfhVA0O//zM4FMCCtTzJMLswXgkTjViS2AtjJrswwoeTJyRF7DMHrFKGoGe
bfW1Tpw4Kflg90CBPq0LUfvXmhz72yRsnl5SUXoiJj1TT10UxgrTZvnb86Bs0VvksswqDlsgCG29
z3Ba1XTZDjg9W1G89zWUeod33OYDNwe+BVd6mag8uPcHE7roVoKIOLvS1Vj5WILvDRRgCErUydxc
5xTD10Ft9zaW20Qs7W5jpzDn7H2Wdpp1VJ8xj57QUsh2FgbZID/dEvZp4PpQ54T4uPh615nKpzRp
dCkfAJmjMw45bgaLFP9vfPnQzdO9/n4TX7slYolKas0Sxg8/CAQVvmtsOVnjnVdCkfN8uvXGDpJ3
VmS/xdW95lsqzjPjQRaApz+UIU8TIDIHT7oRof2rigjdAWV2E1uwWhukizgsQzivs1HYXF16MbIZ
P25xQTpQx1NRU5LMzHgHfxVq9rIzn5yKxFhHxUo3xpYx8YbGwhGWUs91GRhL01A6xUvyZz02OgSe
s3knxp0oys/6AF5Wg+Jjcho9AQevczv3t8RboTRExMz3+7UqBrrzfW9XNyMUH2/wOaryAgON4Egk
4bHidigN2iewWRI8XX3NEIAzEKFWpYPHWskndYqQtFhLP3VDWK057OwnEQ/46EOk6Q5x6lX6Tx8E
D3pnUBIeF/uLsttKor/O/9M7BGgWMEzUfqEIbtqexxFa4DwqM0zT/+wiJTWXWzTcF0kHAhJle+/r
tHKt6EhRcum0+Kzcy1WrgnP9okARIkogYpZuC9UbDTXR6x6ECxXWtwJ4ANeugmWimVUf9FQZ7YPi
QAITJmP0tWxUcrFNvToBT8R28vgbYI/6QWvK6S6D0/uADT5ZwdI6jP5VUmaTqlLkWj9eZ57eFOE/
JhwaVVnlxLyORRkYmufWZDcP2XeQB2HVbCEaHKXjWPz9jMizy9jD641W43YD7pBfbchgmQCXffbl
obsTDngXab2mda1qQrS4W1REL7Jii6mPDwDlKhh6IGoWsGoD/XYaazhTw/LMn5dsCElvOZpRYMRb
lrAqn6Lr18Ga62h5+g8cgBr85dGecXzF33vTSP9n4o3JvcaEW5gSmiGAx6dX538/MSE05NY45SNZ
10vs5mPSekcLRRjCyYrp/YmszL3l7Q5zbnGnSYcPgeNzcjHbsgAGf3ko2V40OgjHz3egxslREOF3
J7NK7vgsEHkE+cMc3RhV9p55VZ9QuRPnyRHerIsxUD611iQsNDrZ2QCejcVYk4g7s5k/VZBKovWX
vHB7GHW05JqAnl6GO7xwqyGjbVE1k3aPGy/AWqF6t9qQz5EN87RS0zEyNk3sXNxMgGeGF5938rGl
wYCxS4JTLQNx4uVZbQT0rjtsXu8Wo2BDSOhcP1c4+aEoeFlGulG18DNH/xeyw7+XPTTl/mc4nXWU
bsVyhZpnXW1P1kO5VfBn04tGLMsJBKZlY5EjQixeKkPtlUdhiM87Ujt9rsgm7oAaivbW7EDUCahN
o4XmbvOyCIynrUXt1+mMQ4m9HlusIBPbDpaU/aUGbfYMl2FWdvy1vw4TmJkYej9vsIs9W2n01gQa
3am2jljcOXY1aHkRGvn9i01WLJwysJDhOQDWNo3JnzBYtr+pXWKMgo7vp9GsB6HytGAukuM4geee
AI18tUPC/uZswjrXU8hakOShG4S87UfsI5jY1ESpz4lMcQw869PmQj7Pj2Oys/gLBEKT+RqcUv/e
0bWFXChjIaHbk77uqawE4XjgXItu/5vT7F447sFWs43I9Dq6FHB8G3PLGFpHXSLdc0fntJbxqRGL
DLUCkgV37PJo2ClHy4tdBzEpTFD5QXs41e90Ss+bUfIHS+Sm3d2UmZvVcf8QGX7KYVC1C0oRNXUk
/ZOdWxE3xSAeyit5bHkRPHHAMlXTpP6oHvixp5YRBRsfKAMwIY8w7SmBKowkf6/X7ZqioSVHSxtR
14TXe3Q8HVBTZchnRCCr6rsKxK7fZTXpI0a4GX2E76JpjXKZzpWIr6JePNZ+7+75GhM4A7vE6ISS
DXt8MN426g8l1CQTBfBRPYdZka7i55fOrm5oy/Pz/Mlp6XqSCqpzkoCObP2FUii1spvKSC57HIB9
ZkulsCr3HOVbaSBLmzuva8Jzza6ikd2tNijta5/WJRdyDU08zNghfeFQF+7ICiX/084X6xQ5Hzhn
Jxbpb3hQ8ZKWdXpMvkeqSLKumFgbqeuhFY8iVnZK2/4aoPq9XMg/aBXhMlB3jyGspAdOuLEpGvFJ
ZlxJPDUVbNjxrG/4CH9gIrAOzd+d4jqUcfk7A/c1tLg8l9KJFwL3MCwI/hniy/eT6J+OI0flWPOn
JpPyWfb9YAAl9wuUpVEnLdLrKto+EX1HxU9ia0qt5TKxhCdUTb7Ts7ycp3ZIjxpvkBQJyAuknKhZ
0EIfkVNNPPsa6sGh0BTp/rVhEQE9Jsgz7v7wSOFkmYGfbpcGnYmJQaNXH+31FfCmylWWnIVMURO/
pt5vm8c4kL4+Xaurhk48592R15oH/lY1ybwhjCAbFR+M7jGtSaFCXrN/bb64YshFvN+YH8TaksOf
j69FhKCfZhMQtUOePv7QwVuFhOA+paHl0ioSSlCD70cAiymnRh5ePeB3gn3E0k2QTFZXzaNwHY3K
vNqs6ecTVCUjbuFVrCcsAXQjtIFO+HH/8Q8x5v94IjopUZI76FzbXhD5wR+kSO+P0qtl6C6QcseG
5gSvb2cSlxIEmKIc8tfa1uOejqZDI7C65qkXV1s+56UUBUNDGsBG2X7alt8dLeRpwxGO6KlUrCQM
YZHCo6d3Hfx16Sbmw8yK6X6I2swT7INqgHW8kCzaAnc4sfegwoJF0rK38z8zzA1RAaTtUCKxfOD+
Isq3g4gvRsrzQ9lAhBMEnGhhWJReP3zJxtgX6VOpvthLOG4hDSjHi3UtbEicxPqCMxOoXO/PpuNU
dVlhXpS0JDxBFWUl0knCiGgWbOoVxE6sqakLCCa7snmFVpxocKcpMx9FgvwRkVxfXVQnJXUd9QXz
zkiHoLNbk7oEZWuh3Sy8T1W+uBSlRll0LmfGIUImq7rQURGXF6OpFIJYjV1BpGIioSDk6dxIvBb0
vB90rEcieK9AW+18tmFjnj2KTYniauFpqNmJAzUs7Gm5npOtP9K9Ou5e7S5xt56K6wbof1UIaMAD
vI/ktv8BxbxBjox+1k8HReSLcut/cohPSUaypwZ3maMtlvBedkPgmdW1gb4Sd5aWZYYuU6OgtinK
4PrOsrif2/Kg9ZVexAGvAfE6Hjumnf2jRjpkW41diLRhM4Nod7ZcKsN7j29Pmn7FelUIdypalo9V
QQWZnKtnJhVvlhWy5+k2Txum+D4n0PNMHsDTNf6aTi9OFQg4elb5oTa5vQ8V3ZqelF4jBNEFU3kW
S0q7+UXEMnPyFiOS7lHQCud8n8UnyZgOPFCX8xdye2EnuOncgKcr9Sw8mInuXo0BltyHAvrdBEBv
6A/UtDZBf5+qS1Lu3/heQZRrDPkdXaOQO8Nd4CwFltxFWnoLDuHRSzImg8JJA/i4YLcCNvSGWct0
hZ0gkae4t5EXWOa/2hQ9GzLkvsg1IFwnh1VvYqBRk3Asov/LfDSgmKU6ilLHKn7e8TTi6B6CdizS
HrkydpkoUyo+NHoMOhznW/uwPYTz6uU3mUmpHUGlZvxMfF2aIUJZ9XwTjnyz5ptkwhR1gPVanEdl
7dgVasw4nGl7UjBdgWDrmTtnaIndK8GAOLrKwVXa6Gh6i7zkN8h2L5dVOULFtwOrqflg+pCWYIEO
tAAlGRHzYcUgVpOq0oT0p7vA0U5u30zMEIuT5vIej3eQar9EW9zwWllbbqLpygiULhJY4rXpEl3v
FdMD/SM/foMQQnluN14wwVTu1t3c402UZ0ztrsItl18U+oKuncTpeXe1KNxjPI8+PcrvQ3wE34yn
1YSks7PA+AG8TBWf/uulKIZNON//DrgRSdbX0g6fpF/T1LapPlNGQq46yBHxUYA8NX2a4fFjrCuA
RulkAU67jTQqmJH/Nvl8fMklVImYo4QzZDXGpmfAu82tYSxXkmcEdrggIQIztDVdjXP7YqsN7Pxs
W5QjbEdncbNbXyB+NvUY4Xdv/qDAbLnnx9JBIJnNdEXwOZ093cGDr1vHJIG+E01UaWrWZGtFcyl2
nU7w4FsHtuOH/9yMpxtXA7RcXujllNlT9/fP9rWORBMEZQC7FXtoC3DfGhBY9QQJo8/UXnFpDCYu
/PB0nHn3QY0G0M/ozvJZqeiPS0vcehOVpKihH41aIKJKDPN+4nJ3BU0joN7nv5QJs8rt/Hd9eXgr
9ZfytJZpFCvftWUkvPApE4VSZYXacCqbxP8Wt6hLGFhDjhLCcgKtyXsUUPHaQGqTtGoKpBURXYs7
XTDOKSkVqQs5tMJ6KQzV7blo8FgEtxKFgHyIr3LXRplMOGwqd79gLlqUrYEjonGNa59wBKwSCdWK
lyynCddKn1UfJz7bXTaftmgzAWISUXYOWTHq/wsymPgUkyh48NZKWoUIjoMhy1vuYFXd5J8m93fD
0IiTQDwOaEU7OkpXepsj2hmEvWIKl53uLzDnmmdhutNcRm6nVdYenseHagQyF0D/qAcCKeKK2HVW
jCxCEENMrNUY7Ppzhs8iZ3TH2at3G2LXjCVDpGgUg0p0BDE08vntfD2IOUv+XRRj6LsMZj8c/pcn
3vUw0A9RnD/gR5ij2VY5t5AADE2LExQOaUVSe/JaZ8Uqnfjmh1dF/PHXTDMwKcivhJlXD4v7tm6X
M/MXSVWBAnQj0K666qEEryWwOf8ffGrFmqJTpYsjNSUbi8UeOePfyKthvCGavrelV2xnS2PmVSpQ
nXj0fPuJsYbGK+/Nt5t3ONO3iMhhz4UKUpOy0lKRZTfbyoRDhP2FWYQ8vxQ2Sac9EzVqVdfKLsDA
CFdheu+aYBZUtvZkyJs2pPgQ8+NBiEYwirTc1TlqDv3I9SO/m27FRD3w0w/s+IkC9NkTwUU4ADqI
P0vCR2inp0Zvf0FAdWIqTPfoOg0K3c6AKhyYJbbF8dD+Nu6iVl1EITwGH3yUKkO4AMpW9KZ+ZW9n
swd236B8yIbYswdQXvChxCmk8MPUClqPTYgBs7KxgDQdNNvz4zqqdmcRm9/GkKOR7TWF0mLomUuB
un/4Ax3+FuzmTJhhsSAg2ikEYJeH7kZ83dLCDO8T/aZoJPi/uv2rFFqk3MpEtg8twS3GFbu9X0gV
8E2Fdm7rgyAKH4cUJr4/DrBlXdi+SkGT/IPGvi9Uoml0b6QC6dp/Wkcu51xV4ulv6Gg50flTUV1v
c1swyK8ozhbhNVmke1pPOd1CZxcxslOCWcnv5UpAa+Laf16b2sreul40OxryiyOgVIFq8/qec8fW
GcMSkCJXuwT+t0qdSayqHlI13WjHSKdPmLTWGW2pOKyF5dxF6pRY4Fpp0wWrl+2cQ7NQupr+esIf
KVyj2bMEDbP+/i7jZY5vZTirbEhV0Q+GIxiB6Q5dF97EULB4rw2rzfQpzLPOA2cUG7NGfQQ/0HlS
323RMdUiUynQFf7cqcBHn78tx7UlU9op9UXG5OeS8XAJx39eAEClcbVQRRTgr2GN0H4jaEp6DADo
Xv2ZckP5LEHmzZ7iP3eknCGiC19I+fi2mMwCjyLnT9GpdfySa9A82Zxx4+U4Z6vG9wEVZkw3Od0W
B4hawBDhFKG9y45YQM3jW0yl3xZnPdM2p0hP4yz42ivfhv4TMzlci7Bmy/yG4BHpEnzqlN5jIATE
/YlbFfR34XfuJI6VUlNiHhgP9SBsuKPgmvm99NBE7mnlfOyCmoPbjYu0Feq1IJi0aZUL33KUj3N3
mD+iIk6YlMWqboPBm+lHJ7bkI8fZk/7hExU0yM7o0fl8+uC684zYIhQFhSqxay6wLPOU7dd2envO
s0ylNp10OpmAO3UglJWVh0qbbdPPxIYVETcpbOZr9L6Zvc9qFKRrF0U1KZDypYYDD4hZwdLXlaEj
jEsLYXM1Fc00KHgnmo1cQwMRgVdx0TCIApibu5Nf0/ExCLTqd1txNNaumgt20HIBO6oVd1CZGy7T
e/HF//JKHUMH3vyWAZvLPM6hC4gB4FOs4XiJAKIfy9mS1Z5DMMhxYGf5l6EQGkAC/4iUpZXSSqor
yV16OJXNUlmcPqZCs6TZDjUb7jmIjT/t3jEF6dXD6gTfd8RiokL18FhsQDVBjvVpwW9mLkOuyYAJ
qYuZfba8ENug0IESEFM2NcdzDdTrgb+5qWXqmBlczYIgA7F0ZfWBt2AFZIDX3Xcc4WdXP9NPVYkc
sovdMl6Lca7R2csLNTDkw0LyJctIXiF+FWXcmA9ivgRfHoQ4Y1/fjd9vyx+Lsi8XNTAB3ha0kudE
w+R+bzDDZ0WFQ6nCeGPsw8UzH1kX/uLSdJoVD/WYe4dmDwhqZD960jUAul7/zpoRWOKyUdcTquFk
FUjcx+S9da09u/0rZcebkw1Yn7i84eQpXxylrCJJUtBr+FJZNmRY/dxD9Hixu/BAiriVQ8ieJhFk
n+LU4xVt7P0ncfiV/HhBhQKhCas1aQFOU5/A77FnOEH6M6ktv+YJ9/AJ9dyjSJXXFlPS6snnMR25
fJewYKvLsOU8SFAYz9udpdUp/Lxau47Gl7gcz4Z84kMwSqpgVEtC6adMSiaxGZoMLp/Q/O/Va8Fa
zSMks+ocl9Lw5252le7MehUmb1K1Q1vv+xNjg8TPygP4WQl48rn4j0/ZdurrLqIs3YAEif8MTOE2
Nv2mXxGsHK3tKu7LijmUk2K67wNE9sUzx3TS/sJ7kzfOYyMctrQVHJnaw5slY6xD3tzU4V1CYqYF
lZj+6BbGpbtTxSZF2JktKy4GTUm1evVxaLQEcSOezsnN++dnfDnAJny0L3IyOoqNxVT/SJZVIaWA
T7X38/Xo4On4Cm4WSgXtvoniy2ykkIMkM0/5KUb61G/2PMjCbL+lVkAZKiegTfxM692co+B2pjaS
rnv/QvCALF9q5BCuCwaWNu+xG9eTyFFoxU04u7M0LWI+Rz16C5OkaUNwvQ1T2Z7HgCO0I8Q0yovt
w024BQSqBOIY3MUJyAK5M97fDW50VGlpgCRDyd9FQRuG5rzHus6/ZZCgT+LrBjvF7gokg7aWg56H
g2Db1/j5W1q851+0x0hEVfSQJz2tRWXK4fz0GdsGBnpSdGG47oysYmNE6m4mrx9CNEVrsA44m+zX
YNWIuUTrcaBaIZeqw7zGdUVn8181tY0yGcqu/LD7O2cxTII4jjFDs/C4/H2+NJVFwsAIVJtbM5ht
k0aOYZGm8uXTMmlb5v9L65SoCY1BVWaWzflMrT9paPCj5Wec2bKZZ78kc5Rsvy4Kqp36pmLhH5Xw
W8Fw9P5QTuFguzq4FDMOmS/NKvjddoQDKwlgIwRzwsRzDnVR0EsvXjyTYztcKs9boEn9oElr5Omy
Y+VGitsBRiO0l/qudzvNubMncPS6spCKASy3p8N+sgl0PC0DZzaAYtrtKxSGsPjNxfZ/TeukjKpb
NyLiQyf039h3WM3m6zuYb/kZqcbPYoMp+ael0ljbpS5tjjR+sTFmk3htJ+mcnS8QYRJWKro/vN7j
gFEFZoK2ueW0T5XoMgNOlY6d3Z4zZ9XNp5/co2myk+IAW0m0GsT2660uXIhH5jDFfvthxa8boLch
dEJ62RpNirICtZ001MaHUFmXxZdpNf6K/7DuYxUowEndo2hKgsWOiflXMDH1Tywn0W5yuRsThp78
2rIoDPExdbrP0Dh52TK8HQIvKT38dcETiqOQovcCn8z4jigikrImoPYbVadoRPQxJFyKMxwobll6
wk6sV90W2cJPdAnr0dOItZdOzuljh4jh3FxmivpSj+Rp1H8Ge37QytjCzD9wYITPb+4HNC48r8A9
yNRftUsNKIlQ75Q/JzEzSBIuL7JLuWsaQlR2xlj+SRLXZzicleIOO8O+FhELPhpRCskt9Oz6vtAB
DF5t41RQzg/w9aSeESBwMnfEY2M2p/seeJn5MydUnvd9G4tLeGouYnrDSHiFYX8L3XApF2VOtmvq
xq93/WhvJXMO7KeY2/MEuI2Jo1o0hkaLDjM/oRnJHSk6OExrc175gWEVaZHB8OnpHrE6XuJ/C8rA
OtcxAZeFOmrV5V7i4iixqkQSDhf+w0KT4B4WYJjYmrlgLfDQF6JS2o027LS2VctOudgGcTt7z+Ch
DOu8sTcULJsyldLj2xYHvIQ/7IzIPQnkCdPR/+hSHu9NZFSEhxXBddrW8XMFBl5VYKEmGGghlLR8
Sc0lbcMNwnGgUSa/rQLG95zO4Wo6Dl/wGgfzFDP8iSXwp6YJ9Vt0twTAH+kWmNsDSEGdK0Oy+T7x
dMqGaWlvPN8THWzxfZ9NXFS/m4URpPW+Mquv4s74e3fNUSdYtjWzcCwhgPYvgAx9KAHftt5/bywt
TqzHY7jTLBQufB3+crdgXxvInlC3ktyeSrZqirp8HG0qNgulBtba39RRJkS/JPYfrohFq8Pt0iNH
FG3vNE82PyqmbpkMaOb4xLBgzSvtGEENS8ENWGGnX/RNaefq1M7HfDw2oZpmlD/ie1D86fp4oqA2
6wNqyzoAckr5RsK7UHyCYz+0bGLkcBTSCaKkS+/mdbihjtHwOkkDa+CsNnrjtHJ/DNr1/dxj8Vum
bikv39/IeEzljUEQcpL9kb0DwlgRumsNUqxtyJ2yfeGMEKhmfQ+bwf/MsH3Wyy46kq8+Tu3x6nVe
xqMF2hvEC7v4ZFv3woIxTD8puOSkdg9Dibgi32TO3Bu3DBzlFTh/F2ca049D/KKqK6b3cRhvUPGs
JL+vAQpoU6hzOe1kzYMXO74sputcIhyeBH2qMmweqLalVcZgcdRWE88DZzAM2YQ+UnliHxN6vacY
P8NDpIeEWZIIm1IIiKWFNiMgLN9ZyaLM+maTV03hLNAlackWlsHDqgSxVBAm6EzbYbskgs/InC+y
Ymi/0CbNM1KP/DKBUcMZVnFIVoQjJnglo8Z7jxzeZ95+m5oFl8lpG2EAL2zz8GJvyDql6fOBb6As
vDJT2uBC3NlVYQc9koawEqa522b8vuwCEY/vfCYXAH0T6PkC+T3avMSfECn5kk542g6vtLpptpSc
vs/VL1WyD+LNa33vmkGUoQ85qYo62hcD3O9uqKZY+24dFu+h2D6ewIXJ7BnCY796bLV5dlqVeTQU
sgbqSIurCzBgfWQDEWb3w03xki9XqVZGFa+7mdHL5h+iaUryp0o7jlmvEDOybWoZp2qTUB6ulVGp
GsJCm+5Tzvd+ajVU2a8AgKy6kGiDK7zwRI3U2Jkwsrxe0aWY+e0/iRR8IiYRULyCrRJXJWOZHMMO
KhhKTjzcDtlj1w2NguYW9P2I9n5x+Eq54ARVRJ0yXd/ptv7D9MkBa3IndwtmdKLfe4yeNcrJlnQt
lxprDZuIvy2PJKGwiJAEpAqPe/+AjQORQD9vHkVgZKsT1ShmQ4mF8TpZvlOE6m33Jk3XLTvN13pb
a1HdWBJeQvvlsnbaK0Om5lTCNJs+Vq4NJ17nuhta1hah0MHiTO1/H6LnElw2YHlgaORX1Ivp2PM/
iUNqiU7GzQCACuYa98EF6EZR5fTJ8xDZEiCctB8GaOuRj3r09B+Ki2UttDtJv+1i+a9pdVqxa10a
zh3vG5j71uwboS6df2xP/boYHLAi890pCEbOjK2d6E2jLm+8iZRgWgCMfZaecP6xM7w4y9aPLCjz
1o3OzTn6RWzkA21fAwFInZvek66KQuCCoDxag+u3ikkBruqslOOMHo5E0OTc2lThKmQaALRTQ567
aXxcq9p1gKI/jfJ36ZiHs1LimwdoXMjWbmtIsBzhIQIZ6WR0qtR6MabY5rsXyz1Jztqew/f4YtTC
CoGLCA03C4xE7gu35dLiSBu1mi8J8eJfthC4D5BlLtG2oZhjbhuJKlA33VneupgOknVI5SBU4W0m
gvo5rxMf2SRJjJJsAelHD/lShyIQWF/r0jNKoHG7Rixiaj3DHfgo8JQOcq1ylTqQ5eQ6NBkoA4OT
VWL5ri9i7WmL5+TwQ7aTBH0ZryObOpHDIZ+/Qpwq0/ouCbfoCexKSBtBCUuLePjV2gQcdtvOMG9l
dOy4V8cbIkv/r5ABX6QDA1ss8IfDWtMVkR8hDWeXscMj4uGoawJEN7fDoBNeF1kDzc4FSPXE4zGE
T6Cw9PQCcGWaoYOpH3u4EIWfHM7LwURue2LsCdVOtLTp+Ri3Lr3OnTfLy3xWd/2rxkgNdH07m07h
N7cyXs7uV3+mOhDlp4lsQRXskYBpKz769Wnb3YllhNJUuqAzAuPHHwMQiQvfPQnRtD2E1rgGWws8
+9rJ/oDblYtW85Iz29xpnmz8z7ncolLLC32wAQ/QnfEcTDOqmQVxvtxQmfP/3JXtE3HkdDtEooM6
H4DeMO58gFJR629mbdo2Sd+7puVnBY42EoN7vr0sfnh+8P5KaQgIoOenEakvcX3kS5dL3u1tLZeV
viLLObQAggpAR+BQGtXuVkHrBkdiIRDpOSKnaxSzJUXYdE3IT8BmS085XRsGUCCgKAqm5+pLPQx7
p+drMkmcRz2U3pDq1uyM5fELrPULyVkUjT925p3of9kU4aUzFSZix6/1vkc9mHgJCgZTeYBe1YEs
CGRcTPJVVDYHoMQTVUbExYQbToUXZToS5NSoQc8Uf/c37S19W9fhJ3mwZviaEL7xRRGvCSno/BZL
qp/h1EOQ6rxS3l6WES9QdSqTDRBqgLcfQhp2Jqq6Td7fY5ZWtGmqKuFOkL/YBb6SeQcQjmua7zCE
rc2u1tMpvldvzw8m9oxa9UlW5l2OKPiYOY03zF7dB46ryT58W/SHZKCXDxnzxRG8YrrOH/IBahbm
SYiAyk6CWj+T/TTjX82cRUzjGeR6ePTsJq/AlkthGJNAvvLN1NWpzb0gfE2VY1bq4CRCcdmY/zFf
gR5VKMQsMsIAnNGMfMbu4ihu0uYTQwS4FRZ3yHaC9OwRG63U3cQzHnrq6BzhcKYihSA05Ga1haXJ
hX3C33rSCW+M9qVF++7St3ckzyGkfWuJjMV1PvcHyvX6F8/KI6OfBYMD0WCo6YszCw3aPbXCFWzw
FItGKKV3U5NrIbnN0sK1/BUQrskO23EYvPJfJg9aSRLGgm3m/3ED+w3PVlEh1QkWfYxO0m85gNme
UhTCGzyJcnShMoLFnTwjrHgyJWH4XPxc4yj/KA2CWR06KR0QGMRX13Y1Yt1WaeDIDxfOTmDZ7sVo
KIE26/Ik4H7aX+PEx2NFYYoAntkpm1uk6t1CfqZCVNS1ofRw9AAI3jkzavOVMmhIrpIafgUA7rPg
LB2ZtiBw4MDenR5yy+thhjkInGUAofWivBTAI1871yiD+CdxfiK9eyZV8JPnjsQUD4FJ4mDWydOg
gkzb5JoOhFFyA8L+Lo5JjO+WVlcadanVtlLGIgFyY4GOpXdOaCCz118qtLHHGgSlWSOgUeLJrElF
Bqve0eDY3eZoYOJcj2ZMgD8kdy1/gRDClBVJTGznlMBGMZj5Dllr3/IjLKkFgnZVsPHULSJW6Bsg
55ZgdFU1H9RwNc50HHyoGw6D1SrcRfNf6L3TPu21xb0FmnTb44P4aeKwWJo0/tHHyMsf4YJcoGUs
A9+EgqXS2SE9UnJ6C9zN5FE/LUTTbLSdZ1lniZrIv/ZIq+Qysks9/x3jQ76NG0QDWbAS3Zt882uK
t4f8WOI+5RMyuI2fXYM1QD6I5AkeVe5yhJUmAP9aKcngEuA33rpbWvtgy+SQ5H5lX4XpeqGd6yq5
QCJwBZTWDCbL6wy2nALyv8AAQSiH37H+3EUavPhwlZnvL+Tg+QntHxBr8xW5tZpLt0/dPwBAx6oM
4kuXGHb3jW5qMSGK0F8b/c73GUpyxiPmPpozUZFEekZUlNsh3tAMz0jFOi9SLr5eoAQacg8qKmez
vc/HxOVSKuS2LCqkThwU+9BHihkpyRXjmecImeiJC6ABaGNoiVcZZ3TSMiPp9SMBk3kQZ0qmUZ7S
+YIdKSMaQ36Xo2R11g2HaS0zQQeoGUo2kkJFHBDtYLw0NTqVFRTfYR3PDvIYh7AokBMZG444CWLp
fo2Jvvd06nhg7ix2mLiyT4ozvQHlma3e4o7IUbw7OHUvrEwierb01nVNnJ5QRx/95xwsAMXesoPs
x62AOnDe/85xSl8KWCLUkrVI+gZq4Va0Iqi3f1QSFi2JcbU02B3i/NQEdhLSaTzG6rl7qg91SXiu
+2gMWQZzIenhAGg7KkWbivFLS/Qhgu9pZ//6Rmm8kt77vuyI2XqAGzFZr/qLHP+Unke534B9ddjS
miVE6Q4iUOsKrE57Da/fgTGD9WziZRBPNOR8XS4zMpCs1kitQdiYfKcNZ8fSnBAbPUOgMXGZx/Q3
sMxUS2fL4xw3BV1Zbe8m0job2vDZyuSnIGse/bPZ8qMvs8RfMs5KbFzOnVbyu6UK8w2AkOay36aR
SvpRz40qtwqQ3L/lAcH2Or7yhpY5pYvTqiqXIYDoOEJRuwP/7JzdWdbxSsVIEldyN53Ih9rMgUBO
x3KdfnXyrw1ah8WYTB4WczZMReSyy5DEVkNC+4G4KE0bsdPIYv/WwndiAFVhdCe/LYeIB4n/JqQu
f6fuuRKFaAG27HfuIwTLKy4KY7dJkNSICECcUbE3FwCcgS8A+IfNHgLmIbIF9xX6+LSdMqOlHz1L
bcy+N244lY73gmOaj+w5IkZSyxhIVX3cQCiVlfTC7PkCZGm3j1MpAF+6ctlUwglqJlluijRJOkA3
2lIb+mMQnpBA6K0LvQWLuHf0aNAxURml8m0MvkeLJdbXB6Bldkmyg/1oIaD1GSYGCU3E+pbTJtCX
TyXA7Mc3lIWpVqpoUi+/S8MpbCB9+oeMDGcb0XxyIDcFi7pSJkws9BcZsNH+LreYcKogeuSgOxSb
brOefVPgYYHzhCnps7AutIt9uQtoeqhcMOwYkodTJHOgymkpKPq91GfvfiwOu9gaZ1O97xQVtG6n
ecAaZyY29Dcsa60WQ3tvpHS4jTVLSn5KSYlZlZJcW92aajdoLyU6Lj7J8yihNLGOm1p2+4nlSPQi
NjE57INZLK9K9/HiPvWvaDr061p9bzhwrLWFsxbOK8thyH+gacl+l2RF2NnQWiMYxBWn/+PGZ8rA
6zWBOyDLjQ2T+CkOwla/DFo5+mKZyQgoP+zFclbKImAeZcCkI2atwxfSgERo8o6XJVbEW30o0SCN
4kc77/BH01EUTPhopyQySfps5Q8aWz7ajlUgaWNm0WLg/ZilZoJRh++17ZUXOmkZ/fA2XjRdUUGa
1LcoZf7/TH+GIvmBc5Sr8PSiFNYzZhEmgC3LUo5DEK+5y3j5p0axSkEabsEKRKH43BzbZy4TZzeC
e97+vIKqi3+F5LsxjZCefBrG1LWr53UIshsGkBgju5LmEaHcM88RC3pE08ZR/gAnqOr+1vGLRf6j
dnZTtC0/aE1auDx6f6gib9hELaU930u3ml4EchgTZwax0NOVK+z7ZAnTHxMVLvfUxkTeqgtfbq/c
8Zj2gm3m3Tl2lyrlBwUOjdAnduqEfJLtAmPvZdcYbgDMrnLobMNnPlsIouMr1sb9omwXgh2am0tw
BCqveS1L/cHu1jEAQ1kmn6AzZOqlknki+xv5IhbJi2zzE/H8ia+LgbbG0FkiJyc/jrs1i+lvEyNw
ug7d4caX+BrwBqBJreqO8T78uZJ4VYVN3aO1QaPTO1L665WkWEmKKs/w+x5CZbzVA6WROq4Hzu/L
llIwe8boau7i4TS+XOhj5aaZdFzkGrXgHoeqSVE3LUSqx9rO802MRIP+jD4FqhKmJUkxekTs5JmF
QckglrXZnGBlCcahVm/WX6MIEVzs0hMVXGEYRwaHJBS96P8dIkIJ+FRGLsD5ZnDAWCY6K+U0Tuvx
BqG5MFt9jT1Pgp0B6Yw3FyT5v8EuIwKLbhRhr8v5D49yYYVckiZ+fRoAdYocDSp3ES5/Ed9n5lvi
vbZ9YxhNQnmVdVTiENaUlF79Q/IF29APVQ/3GEkjdkEh7Vv4XR9AyK0KcQCP0oIlSpRz/zwq3bq6
2hFHTXBQ1PbP4G0ZHmQwOvtnfCms84foVsUxu44P0+GhrJ4yUFDtvNC7HO9z+AEqmcO/Mktwl2Sw
ocfABJzEjzWwmzObmc2d8Yl21HFzkicpRBtKaFO6bxNfis9MXhsdC2NnAOw29sSAFu2/yvr0BMs1
A/ikJMu6MXnJodKHsu1OnBymvwFPoN3uu7sVIO8Mat4VD8sljjajAVWO+rcqvxI7lcCVacMbDMmj
9/YaEbIgnA1O6mspeff6xu7znJTFTHjlxE75wnTHC9KfBimlQ1727+KsCeczSK6hJ/EX0jVBpIoY
37+mdQIZaOWUCU53LpuFH/kfpWmeahHpm7v1ITMyB993nt8A4CqBSC8cWoYh7LEmOxH5aFmf89Ma
WOFOzdfGj/pl46uiIIdBWwu4vr4wM2qXjq0U3/vSEgV+vnJThjfQYRlcXXN6gteMHCG7cOQdvaAK
lLT3CWPhvBeY0RMNh6rgu2mIK00XDiPuoN9jE7kGio2mqXfZCO8wonnWPyqCy6a7jLtdN32/RpnV
mxcYsw+NOcTsS9DY+ZnF36G97K/7jDccvJkI0TIrT5e8lJmdLlTgQnEAi6WlBfUy2bQ47ExQ7Or+
t5tS1LhIk0Gb+Sk8IPRX9wd12H9ELFSv8SWp3VjRK3q0D6WmNPcJfZw1/xDiWB7/79bHr4gkthn8
9AhGbIMCkmVJBBZ1an9w7yKKZcPOmYAnqM1g2p/BLmyU/sZWOx5QNIScppfV0Qwgci25Ni0IK48a
zKox5WUvFpywQXsbRw3ehIZNAt+W++7XK0sXhoPR8h/MzjsI2g6DnI4j2q28HAIUdBFik6l/XcLo
BC8Tct3FzRF0+OazxpVhPKS0sXm3E1v3VeNLhr6Q+kw3AzvqU1Mx6df4b8AdPBEWMlSEyN/Fo860
QIQWrIGFU6DBo5Y//mlvMlgNqHf8xwmhAFCApXNKDCIQrZUoZTb+A+Ob181QN0T0UN84RZlBEKoR
UGQQHlLzog0KN5XVhXWBvRHu1BuId1m21CRfLEVKwVwCjOydBpBTVv9Y2GrH2CTbAGRST0n0Ryn2
wNDQFzQ+z1HX3W1kLndRt4189CKoPOX2r+NI5QeOlgasilHT2aLrS+thRvIDfndhw9x9puQ87e4/
merQlDMilXdqwX30lXVyr0gQmCPsWodNJEcffJpRmF2SNPU1p8Skq1Wlr2TomdR4uXjVBCX/jGHI
hh9IZYDP1GBjUMPjlqFNhQ3omb4CQGgEGWfWGh6MpvKJ1SX5pWoXyjEwb5/iNlh8qOB4JTC3QmK2
P1+xTzOpHeJ2zfZRRODtlLEKdpa53D/1cS9hcAWn6CFcq5O+ddAzTeRH5U5B1BZpYGMeBQbqb1uU
ARK11PZd6uf0VDt8qhjxFRjs40JFVSNUCNL1615L0opi55SGk/eumtajYJLNgTqlmaMhrN4GB8GK
05EybxvqElaLrd7FERh35xRQMbpKloEtzamdqlsXaazwX8sGX7sTW7KlVVc8xrMxZbqVL1LAgSYk
vnfwSF4lgIf1q4GGPq1EwPFJeNH4rZkCIPoQSHyp8zsUCZ1gAxDjJW55ZBdLEvqwDVOw6bFwc6tE
oCNNFvVBkrW64uYTb82NeGHRA6Dj8vIxrIN+a6X+O3nUv66AQAZu2mHOoXgS+fvRUna6HUMc0yF/
eAXVAgRFsDZklMKZ4OGt4YawUxURfEr24keaSFPhfwdkwEjfHGvWsI9o1HZ9u4veIsPAVzBhZLNp
ixeYz18RhVKSZ9XaPqGkHlNogm4kLSIRIQhP9SePyDsI/rtmCKeZjxDq2oFCqoD0/MBC6nVAxhDd
alvuXophSk1CQ/OCqVyyRvJRauV3f6uvzxQ7sej539ijbJSKqOOygtSGNtBjwS3IelJQSDvz1FIZ
KpBeWIHcW1x0TrYtvr6U3WeLPNm5I2ZoC5JVu1HK4Vnr42IqHj0/pzpppXeq7GMAgzXPBIMx2Xg+
OuKB2Js4EfWUzABz0zg897p2bZjfposHZ3+a+qBq8Jd2xbnTyTX5I1Evw7+tYhjBLVOZ7G8m7O5q
OmAw/11VjtNLBjb5f2PvfB7LbrIHS2FFHDbUD0+8uZ/yPOqD8NRvgSVaOel55woLyOzXBFQJYPmR
g68HyHf+tj8mm9YaB0+WlH1AU+4wz6WYNSYZKw8pak3R8KxmdbAO1zEDkv4pF+PGgvy4I3a94F7I
KdizvLi8VFHATmOLOmxHeTw1D/eYVTJAHighzl9HwU8F192280FOYzIk5qDs3/5vEsOUmMU6D2BX
Ech4m7eo8wFjGoePK4kyW+cDzWSk3J28AopXOkBi0ZS5iTCWZ/GwFPZ+4cnQN2UG77zhpqA8gR7/
MHWQVynQuDq0TH3/9Rs3dAUEMbjO4d1ZpZ003W7iyrkj+jfBaQJEQ7dq4CxoiDCoFCAhDKhWu0Pw
fiHUB5IKKbryXYs3TVHYcoYTqjia4M2odbofKN3momX+7pLoKjDnka0OFHdkm0EI05EbTDKqu7oc
WcY3YFdT3jRs8icKtFr7nzW8f3XQmsXnxQE+q3SkoZ7mr9lH2J/5YyzCWY9jOJtv+hnz2Yuz9Oyt
oo3Pqbzd8bzatFXeGF+1aezNIR/s9877c8YgT5Lky6nBzcM1x4V8QcGaoh7oedKJWMWwYoaj3yGk
BDIueBPYeIg4YvK63FIfmQ9EEuBzpF+FTI4LatmcyRk7CEQX1QQKoi4khDeDAg3luQjFeVgGdL0b
NuH3aN0YYtGTiPV5V41RYHvF2lRYxtVHUFtAxQijmUZogR8V2mGWMSCcM8/ZkSX0bJf3IDdKs6Ji
jVyomwf0OYdmRpaCrs8oyUDOwT6LE74h3FYzg/ho/lZBWe/0y2xs5S5GgZElW2i0PhAGopWWTn5H
9K1DSWIAvzfxFCdu19DfX9T6WJJsk51F1Swy+dsK7UNtAkuFIMbR7u2Eq0OAKjH2k1BvVN8soaWJ
UKm+tcTPuqWNV7P6FtV7FNi+0+TsoMfCDDtN4b87fcArtyIDd3ReTywPS5sn96l4yOZDq/oN8EPV
fUp5GQyUyLtR2ZiQUlNtRK5vnt3NwsxE4FDGK+HPck5g3K64mvbIxjKNGGxd8vSYUGs4Qeb/7wFi
Li1OiOxWzYcvN4THLOdF9mjcNscGoeaQQJUnUZCBc/TESUdiGccKVFM5HfVYZdtiIyU7MRy/N+aV
4oA3245m3K+B6LBU4uUbtvxa/OwRiffoCwKfRxnCfu9avIK9In93RSfDz3hoMcB17ykrslnuB+vO
TFmFwgRQSNvrynNnTbFczmx57Z74TioaZsaMhrhKf+bPNOHUgW1MDZ0l06Y4nIbLltRm6dNrU48d
YWVX/Bq4O/+1/aNj/1LqTpffiDdAQFjrxVg8m2EkkJYdG0wiIxStVdczHCehzjH4/tN8AQr6ldMT
lQYE4hjX22TAYcOnC9gTEP/MbvRI5+ERDjDRU278J+CzBLtA7Fr2F0t2rGDK+R5FjE71tAZ1jwTL
UFqN225g/U0tUqs4s9S4hheCtNjQkafGel8mL2xQdi9MpxlxwPylRnNN/4vO8JOn0jh7YV99i3P3
IDJSTgCvcdnVQ1XzrqHZz1RALNBxhUjUb/75YdUjU9cDekLRu+KYS/+aZGN77iyCIGyak2lHQbxY
sgmh0iTSjQnguzuaUGZei8LwLilyHDXl8uvAo46++Sky4+jP3+25VPb6GfC2uf+YFg/AxI8eAswY
2nu3r2vWzvSnIeBQ2FeEzj5U7gIy4FWRBs5mpachKK3qtC4jYfEBdRnW4digOOEYz3b44FtPAijA
xaV7Nuafk+fj7Ap2Goq4ElBkq0IyFajQ7Iyfyuvl4050L1PsRHKEepNlVQLT8Z4ZxHCI65TFLn41
wnKLHEepDCYft2jV2zjgJCiNmTw6x+/LEyGoQSYNYlqc7hvUqtr0KCN4q8TuS4GmrXYS3EpPfw9u
pkHDDXrEQM0PL3U4OhhyuGN7+BruKaGGeE0jE1T8DpyV/a8anxnqVYC6wV4I6rRCWj3J28k1JOB0
aM3KdMFUYF8TFvFjx1KJyruPHDTc+jz3Uil09Pge84ZYWvJCN2uRxdmTSMOZi7Fhl1vBc1kXui1m
MYdu/5Lz3owuMAKa86iuVhy7KdBVGnulbfXOhhxe2A1Ocf/tUCtm0SYYLx7gzkY8eRzDdWmxGjy/
frdcVShEdUvxmCQICoEn7Brpsgvnsu489qqoCcw1qTQkJyhBAn+Sa+VJrijkyKWZmcVHn60cZgNd
+k/pD/IDsUD+MYSK2LGDe6exEOjd2TsdovikA9r5MynVkLjH+qpO2ja4WWVwxyYTQR8SZIALsP/6
59Aljfmdlqf8arTM5j+afZE7vJJn8w02df1pmVIsdyQwqp6YH2NcY2mZjJkETm3AK1blfZfp668B
IeUHY71R9r9g5k+utkXRdfDvNtqhfKCw4pR/uKO+rYhrLGpY/wGPD0dRf1zMYFif1hraqBAkwtn0
qCrvxaSmvwEHbS/tzEGwvxiScXYR8yiZt5WYTphvQZGouMmZImvQ+/l8WHkvMyc5yt5FXk1OmjU4
gnCkPOctZt1hbVCKRGfTMfQ0Ds40YVMQK4fdfN39QMer2H/b6c8zjIZmpFNxWqQ13qiS2enAZhXo
ipJ6tjEjU19AmtSMuaIF4pKdrI0EJMm0DMOrJF4Yx089u6aqNU+2J/MGF/Fw98HozsnIHwPYASvh
31744f7ATRuEGcvYE66w7zzMOdhj8RT0Za+pzq0Hia6qwjEUgoqEr0WVSImsR2mzAh4q0AxNU91k
OcJgEFIeSOC2xRBvMRFkoda7Vf+vOE1A+cnm7Jjq5BCguh09rUYuIUCiicSOhR/brYUEcs1SXrLd
GE/VnXe8eyOZb5reAobmO/DffLzwFfCeWTVgHpS52SrqYvixOZLM0bGb3V/PqJx5S1sfhdrezfMb
gw8mkJODXueKo/b/MAcrrs5bRNuNemxeYAowjfSpusxVOLomQkHih/X7ug6Ar152s6Oo7+kcT6/u
nRoC6JUDNODOJ2UNIh+kr4ffkadSsiRUQyaa1ydUZ+h7dMNpPZzERInhN0OKSNWuR50vtKnmIAMu
MYfkKQHk85GFwnQdfP2mjqEAbs8luzqxw3SLx5rdkAqH4rj4nBDx6jwSSr3uPkk6Lk44jfUA0PV6
Yda+fC8NUQ8CdIb26xF0xXTxL1H/kArx0rI2Q7YV2sOZ1tI6gWJD3GwiX5/q7iaoWyT9Bis0KhOG
FYToK/p3GadUxjNtFlk45AqpkZ/zvhHvLcWKfzxJHcIHP0PK1yi9xchmLdxkxQEl4x0IuRiFhAKC
5dCZTUEJTUVoGth77hQwZtzewgaAbmx9WzAURy18RQmS8yonSgrS19Vr15XZCirsmN/14yCKDc/i
URZklTeSPMWSmIQk3/Hj4RROyewE9Rs42aIpqxbPvliWrOwj2Y10U18UgJWe4d/iX27DiGPdLzmJ
vjBOg82FHy4aUPf6Nlq630+UdqoEVvB9EyHeABIDP8QZwO5/gLXiYzWYJX7GuFLebTS9GxwPIlsC
xNdYea/jGy6s+9fnWOng6OdWDKEx5Ky1Mgq+tqnh7HX4Bg8+SJlc/tO8/RCqMwtJL7KmzoXGTIV6
GzGjYh6DOKipItn9sn9JdWJMVIaOsoNtKgHnIXEYGvqUPZCHuCVoBZJOOSCQl6QB1TbBwGSwM7pf
6cf/xbg9K0aVnmUzDhWcPpMp1IduC5EGK4u2uhU1bYx590VSh9teo+06Xg9U2XQ9BZskjtMhoWeY
/0FOwA+u6U8CakDLg2ubiQS3khSHt9vLHze4zhCRnTZJnQC1Ln29ERHxs38E++xPnPmGn8DMGfSG
pnQ8sdkDvq0CKUXOREj3W3Y3ENOQzQKQl8uwXqZHPkl1ZBUd7fV/uDOQwGbqmqsGamlcxlgDWU6l
4E286R5yX+74znAciWABVuPSvRx4FiDEjkQ1icYdpUuwNXv7mkTbC9qQoQM3PiZJkT3qp1Jomwe3
HQwgG7ZrsZA8CR0tNaqdbv/hWUZ54+tisPnKF8y5maao/py2cwylt2dcH2cJgXFPZQetjfa3qxcH
qC1PdC1szcir/HzrqTYpFqA0kDj3aS/sVTjt8Ey/JAx8ZAx6Q2UChbfT8ghMlVkmsmq9xoOiM9lA
ZWf2uvxECHVYtcak27qoOdOvvQt5eBdNBexCstR9VM0xEGUj4TxhUa8eAY4B8n+hxlAnPEEKkwZE
ILM3leBCCfe7Gtrxpm0kY+87rD3jp/bVnjIqti3CWwL5zV0L8CIsLnG7Idn7Pt20ttrshg2DQKnr
aJwplooOI1TBjrGX8aSgaXMTa34GWYKdlEaI6298UFcOt5+J3momjDWS9sbE17TF/lZWgj1G+vWU
dSlsxZqhi+qAsr9/Ftpt85+CDWk/ggLKsvneL0gbIO1e8aT9RXOCzs8WQQ/2Zv+Xa0ZtTkCU5d4Z
OPAOyQp1bRBD4isuQkIaAnlGGSA9PRzE3E3UdTrLKQ6VUdjUUULZiwwQvSMV/JhKGVTzznaoR5H4
8j3+XrcoQa6VUlNmYXegEvfP/VkP4xZUpkPT61zd7ABYIl+M/V8Q96dt1ahAKYq3SLcTc6Usw7B+
ihmImsbUHCixCEtQxCFYpgc92PM1YfQuxjq+TLAPra/6F46fXEF1y+rTfB/HEbwwtOyvFMfnFpuR
/NPusAvynY5HT+5YJyGbvOhKRFaCGt4DHxqw/lv4BZEbWqK5rgj8i1XJTNh4NYMJ7Oft2Tzoun6+
mYAxXezK2vIVGLrpR5k301HSl9mTVWs2u9KSVBDGxFf3UxV8wnQJWi1UJSvdmFLEBtQsy8G39Pxy
3h1kntcPk6/9rwkNSxZ5IuMUBKpFelnrCNWEd310km2rki7Sd3lru1DPYllEGuZ0Wq75MAU22g+H
YxMJDE1sIFb/04bx4x1Wb5RfuM8maZtjW3iFTtLoC+aVXsAJMuFmkwWDvNDirmchOeg9fP4kKdy1
t1w3Wu8sDfP6TvxJEMQ999nC+aZ8El568ZSuk8ydVBC5zGT/nkyH5qq7zTex7isCbdqnn3as3/Ek
kZSEvZuIyB5lP+iKi7A77eSNuQ5r2S6rNBEnbfP1bUhQxrupTbw0FECzWi9/kppcsBqI7z9AmDDa
2qRpeyH27Eoqf+OlzKMYuvSpVQ6tmgAV7JwEOjURrbmusaZupiwbN5Y8huN3KPTDF9s119PWGKwh
W4Q+ircpvcBWvM/gew94QOlPesSHuGFKrr8NBdIB6bxuFSrzH+1Mjvol7TUbuIHJtd3sU2g2xOmG
ISogCPMkLxswZ0sY9LfB2fxDZJ3UKyq5RapUVQk/tAwOWmbcwkzzP5YHqlKb4ueSOJ4FV9YGwRmH
/LmCEFtXF68v7bEFQo4OnqLnFHMUxCAfCvSbyRRd7t4F/LHZgrH5z0estV3/1yo23IRBzfHJCUkG
7Sc7RVlHeVARoJGtH8eK02Qq7gNIBzy4PbQyx5ewSCiC/BWBNZ42eXYkpcY7mlzsfJR9yAD7xRBX
pyuoOv/30TBFvpMZ/sAEMTrZzq9sFKdCgBmqScGpQHrhrLC7WLLTFHtArCec1oZXijpZEdGwFlxa
avrMdYPPOIthwzuBNAtO4pKS2yzgMDrTtl5MlRl1EvT67QtLK2mTEBkuNqoH78siOq08q2146csI
LNigwS3QdTesKpV1FN4fBPUDZaDmTQunfIWoo4YBZ848neX8oWG8yFKcf+15kmmjuaGOFjyzNFjG
o1w1xI8PUoDyWAGf9PmKt301LuQ80mvV3gJlO6MqvslsBXNNR1Cy/pfopk9eiGaHQTMHLbXC2BhW
pOo6+v3l29k1rZ9BbkTV+E7N7leD8rkBW8vJ7ZI9ZWJdn2eo2DGQveVloxGqDfKvILjfvr6IYYOz
mDyfmCzs/cLKC1tq96AvQnVQPYFupnWyCEf8N/uXeuJTqd3oH0JyHXFT2WB2yjvIBp3ENPqIXVVN
lS06QXaCuJal/MEcyfgIlMYQZU4L1g02c7EkgKSn4benGYdqDT4T+EoP12vLVG9ZgdXBFcvW3UF0
DoXI5ybNwW48ILkOPdKqhhMz5sRW+5q7N0O0c7yXakpI+ZFBFf1l3iRMbkHAPhWEN76tu4ADrgHr
H1W8+kbBlthuGBFYu8M+AtvFHMEqa+NQ83czlMnXC5U6MVvIdUJYCXVRc9lzktATygynk9nn0tYO
7du+b796zvibl+MKTv4EuhHV92NIOG9HfsozCH2U29p/YsbJk/GSe0syS4kFwJTudKWMfOZ+X0TQ
kiA5ktf2o6XUpKnQ0LVMoovzwzsTlQIzKectdFvTFCTAyrR1wAEVWKwlEP5y9xQcFjErM8Kh/8UJ
y+1kUO6ahd1zL7tcQObwBI3fYbqFaelxutU9rf8lupnPeeet4cZntV+qomARR5NobkXHwxNAszuL
A3bf7FybpNPqJqgtiSYs4I+qmDJGK3NyY7wnUkEbea88kCdSS85jppgBklWre7rEOhTLXIhwqJCF
fnm9XqDLEC+jhvN4I8j3Qe2rIo6c7FWe51YizJmNITSjIyFv2pOYqzX0CdDcRnfZXG+xgbAkfEUZ
cNEiZhBzHzO/yBMnLLFKgM78e6ZbnRxYp9CSCCZI/BVwD9v1S4BGPCfrvATFZ80CicCFcxb7g7sG
s3WQpX2VmHeS7VTY90KqRxGkyvmIfNakzvIj0ohLCf3zcgunV8qR2YgDTHhrwy8YIQb6lkBBW0ZG
oqQcp+8CC1eetj0vOJ+Gvka/nqom0LEXbTF6j6jH6bwXz8N7doZJKFs13NK76U1/ZgNElqb9vpJI
p7BhL7voToyN5dG5J3XEmUxmuKhcVxhkg+o79Myj2miJzc0L5SY/CLyNvap0PlPH+jqKOlKeXHWF
adLXG2L38E5gSFdheJHQJoUVlcI6mp5GYVUQX2/aHeV0gjjS1fOLuOKrNUNop3So5u6wjJxrmMv9
JDdxLXudRBWBnJRAyoO3wEbzj3iukqc96DeXUnFDHGRy4VAPqym5WTM2kUKZ3zqSw1t4NEc4Eols
CyNv96UO2sbbzVsVgZzaxfTIRcP14oFCVsLGkraeohplpery+bXwr8v+YVPDjcs0q5+iPre0G6Wl
zAJEBFlgnNpKSMbqnuBHv8ftNyMzphOOFAXLvauGFRRTxZCswxvUeYW2SbloC7oUPzWQFK2Ln3WL
Dx7pgCKnRMjEZ4v4W0zDxTaRFhYgJT03j07rFnV53fuG69QNNYkLE2nqkBA+2xjVODhShLy+lKUF
jTlP0lf76w3DpfQ55mjKbsVVSsW9HboqXBt7tV4xUvM6mYu7osiSqA88a8WWsxcrdtCE3q+EcN0w
OlUtXk2b6jCztTehEGqnzn/isM5Vi4GevBDhsWi7sS1xn209DtkZzVIJCmvNNRlZcsnZR04fYFoG
g3JzFlzjjBf8JMuBXtfogUW6pbFbmECFYfkbdCX85mgu/efYoGrq72F/RhW0g2X8Kv+QPqpms8dY
34xORy6XQMwGur3kRlQ3YgRlnMiyXHIUTRemR7JewZhls2jxXV7YjZ41k9+mg7LRXI5bIPbLfe8i
NxMOCLGJdQmFbHT75QWNu+khin9xXsxspYsrwKDjnmprHNH1Tj3oDZX8EWTFhCFVbqYpHohLI2qh
wkcPcGTKSudxebTa0E7XT2jFxYBthPVNU8LbKda7PC+NKx2TqD3/uY6HISBJJN8PlJx7u8ngqZga
qMollSnwPtuxURtCVvMgN58Vx5t3QIGOg5F/6nKxu+QaId3XzkHVqX9QHcEkLTON07aUM7/JTacp
IEqT7+dlwfdd7ySXoG553rTf9hDVJQG/CyhHTNGBQDmxhjesJ2sAnkWVNRsGZ+Q9anCry6qgc7AT
3uDWMWCj1HQ+ui1T+bMrB6ZcUWxK/pRV3gl9xG2CAQWmPGZrGuiU1G4ZUOY8kB9OP8m4SBESt6ih
Qzp6rC0icbpysvbzWkzsjg719zvxsn3drf1UXAqwELqhD+bkQMqbwuqiLIBBZtSdhQqGTugepJCi
HKOlKciApwYsOqqFPU4PAkZet9ElRTBTFOLOU4yPM1F6tW1BD3IH0Xc9UZl8jOIjzZXvTpkaFHfd
tocjQU7itmHem3uaRj2wYHhWsjfRKWATZvBdnBEC9Zij4F8Fum7hDG4rdTSiXmppSXnsg2bUthZ3
I+bj3AHeuUh2pEtKqdlgF4e+hGUmeUGsa1GFZwoEZQ+NapOl22uN9Wi1tJRt+Z//51fUg2celKL5
PKxFb7hiT0PiKhyFcGZbVkRnc9odENFvsiQ2TNv4dWwEYJkZU7pYLLocHF6TNYnMm5hjGEgg3xVg
DmKvw5hxn4hWn6ea27ImHeLjO/uYUjfOYedWC0iaH4HitI3ZJlInVBcDAKebzG7/GPtUBCCSVSz8
ntEeTKKIsvyPMBv3dWr3p4vnV5Z/i7UJErqKO/PEOvLVZdxtox7ZGldTMWJMUF8Zjb5zLH4PuK8b
XmVFiUdqT9+Nopuu5AHcmJ15u9tdgGyk7t7YKbPiyEa+uz2xGej/1usKsMCnCunhEFASmJh2O92S
kGPl3Kn4Fwo3Qkl3uAvjN4xFV0GEhuPedu9bQ41md6MlCAM1r5/Md8K9lIb0HD1a2qTmW+rfKydy
bfIZTy3KG6xdSrWlADgztrjFvkQemOQkDBpNjOqWb0uM84ajQOY5NxClrfZfk8NpOVgBCbVoWf8I
zribTJFBUUkl98NCQY76AcvMU861rape4m4reLtR2+GQRLP0kpoK6W21MMDKcpIYydgQpds82nJR
h0JbF2V2y2kaWOA9DeIrOs0Hhz1vAVtrpK0chqfXvhHeP4bdLs3Pzx75OAFdsl9CBUbnl+OjbuvS
lvmmkG2CwkKZLEN332EDgZclrI9sJ9pQI0di2Js8G2yCdBaUZlQ7Va1RqkWffHVfDNr5LbhxIruy
iZjHEBpZVGZloMjfZbJhDv4FB0n5BaAC/2k/hO7F8CxLgCIRCTjqC1H53QdDy+nskaTE8hBArs5s
S282W5s8S5pn3Gn5IZsMZD3iE7qvggLE0zVdR0wlNXwTHtZym2KrNyE59ArCgsKJh6ARkSFZoU/6
D4VrIQyZQkSNAl9BXU91a0PZenzHKMgGcXorOWjxkDk7u/KB7xmFpje3ksH/yi+2D2l0ZW+ZR8pd
2csc2x/WNfjkm8mKja7ALQvH+ml4ZOe7KaEVcEvIpmVwmDQIitS+sC1z4VX2yD9IyIrUwXyiQ035
SGjabcginkKbzvPAN4r1WzG0EW4kVnNFePOLe1O9QiXurmUTZrGpaKS1Y/sXhfjnjcZPw0Mn2ASS
AQ81nLJsLCXd/fn2VkOlN05jQETZUdEgMbCAcAonmCFIK81fWvkeP9oKhGXTM5ssSo4NG+LzJp8h
SH0j5CD0spaA0zzCZdVOBjd7Hjs9f0R+rH0/KAPwLukOHPYfa6RRZuH7/lnGxwtmTLxTlpVjErsC
iq7Uofa8QICqgkEJE74264zobpcPTsbNF1/QqOk4fRQJsZ5gios1VUwB6VmEh4YR+WX039E33ID7
BJF96kFsuh6tVs6Nb7KFApQDEMrfO9Q6gJasLFPDP06jiu8SVwxuHd3rY99pq7XfU5kZQq/AIrVH
dVG18fOs6fNFtdr+tQuOFwS8OnWDfG/80ixjoVPZYRUe32bnre8ZCjTkzVObkGOcfekGs9ffwpO6
iFoET4NcdvG+bjd6fFGBzwgtgdJxp2qandIh3HbGb57Pgd212TFlvheEKXoyfxZBnYYNK/A/eVSP
zRNrG6lBv7K13RztIYA3t8rUSoZU7iOod38/Y3qvOuj7MsUNT0cQ1wkjKJY1DM+/yyw1vQd6vNOp
0CJ1xbrDfSshdWANKVdpRkx7pVtqihgZYyXKcLzQ3tY5G385v04tTutEBCEDPg6lrfQmWKyEshkr
QGHiGzmVcrDqT+WuREkQ3jsIba6Z7HBc5gb2P6p+nfWY10BiKIMQbdqV5Tik96PFy//eKI/YKwPS
R0xCBsia0TbNb8B0UErMQ0MNQwmWs5bLbgGCnLv7HcqoJTwltcOIGXB0nxPjg/UnptEaBXLG9cjl
FuyWKCmklAvx7EOFYq2fmjz8mGYC+cnG5Yi9qwtJsQJ/IQTZweiZQ5X8bulmdz9GMTbZ+3huF+3c
BPcZgOQW633JsavlIxevvK5KiINA6ADhCM2RMndtrcfLiyD9ZRfDQ2m48sNs24AKkOuJSDg0E4n9
q8M+MvQ+NONDmbVLiHHD+iqL7w1HJl0QziJx4kBZzTU6M4jSFzr/IUxUxhkX/EZsiYQu9tjxSubN
OkB5JiQpyAdBwCO/dYXsieG+B3Tpzh78YHUpRqOdaVGkf6AItxh/2OLqqj1992kKQv5cQdFZosrp
B62nDXZs/VfTn8XVZkwHf6HRtGxI86ZKgHIVhE9NOxMHNLduDahJ3De7bBNBOv/3n2PCCgGL+g4i
eyqdOWAIv8W72Pr2iuT7AR1gJ5iuKEc7e+AIgh7E7HLvznyJJw5MA3vybMFcTEfQ22I+HiWbo1nY
yKL4MsKXo97ZSa4Eu0YQqsCUJGjQpXwPDV6HXUWGt4tpU/EHORzywkxGmzenCYbd/EsFYOXHlkCF
/PuSZrcXSpNmhhFy9/Wjeb7EKKYku5xtRmdtxwkvN1Lnh54VFmXYt70rIgHwmLqs3ifFGPSJeyIi
dnml1Ss/00M+8YnbP6I7dpE04TVBwbFnQS5OsWnLj28c6BYv1ag4TCTFliqhS/iDqNoN1LTxsLu+
L/q6MW4Jv7rcLteQhnHPo4qNPJtqAmrsT4QkQQzgbxjUwK/EIhxT2Jjpd0Y3FLeWGzDRYJ3Yzahi
LZbwmXlYjV6W7I345OIEiwd1d4qv+EyGV03gQMnp8nkzdx2N0MXwk3n7l7SrbxbWofnY/Lo4uwFZ
z4QJONqa1hK6IfnmULro+NzkwMoOBEAH7+8cDYvNQiBb4YHMJ5P5HIN79ce6LSij9nX26dVJA9MR
pSjmONapeUSkEZmvqiZk19iM6XH+stRh/fFwPKlSTdBD6k9+wMLAobzAjYuYjagCLcRI5/4j2bYz
xiZCbkfUuMb7PupQGzsa1nrEl7td7S2UUQNX8XY3tKD5RZpo6wOj9l3xyQtAaGRj5ZF9xs5kM6p3
2SCwv2JHBhsGsWl0xGxgGPl6RgUFt42BCseZy9YakdPqrFKe2SagnVdGUw1wA1jrO/7qp5r4gKnz
2KIP1Qqngw8i+2x3nWLxdTRdD9vuqLiwPAI3SyrLkuK0piWEKYPZM4VfQuEZeBx82K8GOJVI8Iyg
NW1v27YyFdmhujyxb2qHFCLqoAOqaRAhBGbOr24YUBSGFKsuQWzaJ26Vo61PPvASP4UzWwqEKgrg
NHsgawYxE1UrvCWKcPlEe9zxlW/7oJlDnsy09btdIrm4DxrXpqUT3+c13yWd0KleaH+CLjzfAWRF
MInIiUR9HOCkKxuXWEu8a4zFnJwQ5Vv9qqiiop8CANPB3vBgeYqjs2Cw5bp+HJf6CwgkghWqLpFv
Bf8kLPIO0hbK/o1QSEaTPSLqLoDe0MzXCZ0uraHcr4Zn+ZiaODIiQ88reQv/Rx0O+EcVnXQCYoBP
sC23yyQRqvS39ZDD8+Ax30/7QwzZ9adLX38dsSpiMhTRM5phF9cyE+AZKZOQNZPhIjist7nHNBa2
rQqGGluN0o9+bkWFDDS3AE6HZdOOr7kbWxyUBUrwcrP+Ce94YRW18kIVkB6wiVfkux0H1GXkERFQ
XCoBLzV1gKQN2QCobwU1PItHPdIWtslygAfBl3b/TuFd0OVjvTbWYtmHbXL/u/Ovf5yQS5zByb15
8XnlaT7C/B1ZYzWxw61I5KT9DrrgowjEuS4bvk4nlYH8kqRIB/F57LNzkjTOVevnOAdJf2jt6nsH
m4L2jYZ1k/5j1/t3KoMxAD5SFCi93CPqCumARrB0pZfnDplodCzGk5j1PBH/B4eAI2ICqbZ8dliK
u80RJSwWo9RlNnyHn0tIL9Rd2LEuvnTWUOpQvOfBTm4OYbJdJ99SJP9eC4PJAzpYqWBLIshqSrfV
HiBoQU8Y7cs34HAB18wx3DwW2jG/WYqCR57GPO9KbNVm3PSk1LCw5cgmwK4Z4mrf09e+HYl+lzUq
+JJUISVxGVP1rTCYbtnwTwqwLLsi0S8qwOAT1l1jAqfkGR4h7BFEz0GopaaFKwbCoO889PPfzpNT
9dhGPUmeKyNZkoqZzidl5qd49Uyvy0FMZFcP8PD6KAnTmrceaoKgTgB04MbCjb+QXvF+T9K8wASB
JlFd1kpqz6/E36YEzgzLJeGl7hFD1dwHWjyrwaxWwBPhS4PDbWUiE0gikUdgt0Ksloye6DyL0x57
8juNyyPcgQe262EblFGj4f5PT5kUr2pV7hgmDE+Z/lnn4X/7I8pnd3IyUUwkcgtRcXX1ThPKrvmF
433Qvc+ZBIRNSVE80ZxmnaHkuzZ3wRGWBITFUV80hW+HMzHyDPX4bP9qyiB8GuwwZ5rtUTeaHMjd
dayJHj/lV8GbE3nYHZkPrzPO1WklEgGBRyAjHToB3qbynto5CghRFL3yn/sGe4tXpnrDaEYtq5qi
QD3LuD0lM+mqxyNix7P5I//FL1hZsp9sJgejMxqqvfgxIGOrZM80t76HtbrSMLZvWBe7ahtDNjio
4h+fkDVoI/FjIafmXGRkfwmTaOPvnG/Pzkk2UV6TR25e82wmzOjBnPHoG4IlmfrDnpsAgFHSaLOp
mZYEn6R96Q+i+POYr+0PeaEyj93dEgEE7+UsRqjNuWbfdZ3YXB9ch/mTOLnpdqpdznIywi0xVHTp
jbyR/zW8LXS1x2oQ81MP3x6aOD/wuKq3B76Xm4+MuhgJ0qkwdMX1H/3QeP4rIw4C1rLHkBKfnlMZ
xQo2bam7fe70G85rZDbOjUUifm/C8cIEvjpsJ6pEbxpAKsQDhcfVv+DL7XF8y0+WeF59V497lXqF
KXAosm2RsgOv9IE/GEilqNFm/Y7MV8m1Ovk4APNhpbLLvKlggpEAzHTnOzpyCqAH3uqyfE/x7HXf
5pFMHaLD5V/Vkc/l6VZYE/6nyMhCS1xFIKRc/EUh45N/Nl/pMyNjArq/3ZJCKJ8ymkawvr3TAmPz
7rym1YqXYbmqev77xv0S/KFElGnjjqKpWVcOKYG1MndVBJPOV2FwVHzsbJyvBwdGO36XEbSTgSDh
+pW0Q+MPJRZM2b5goVo/9pzjhLELSEbGB56reoI5maaZOWQ4FkTnXGw2YUaZ29lZLBgi5e8yl481
HujfxHMs2Hu3Jxz7C0NSp8BleP9kjOtVZaUpXy0H86+D9qWNgSOit9KOemBOPs/fBxqneTwgYpbn
B4Y9vnLCdfqE7lFs3KUAzkizQ29WWRZhcAKV0uq+4onom4zURSfGp43TRUBVLARiiqcbH2ykZrFN
RbhXV+HAURld8EuJ3MHt+IP3S1G6ogvbCJ7S8khWJHTfVVlGvn0E8/G5dkpXH3/7Km9pzM1fSP3T
Zto/hMHOtsL5rCdNJIJhO9/KkMKHqKkBWd2kfiFfSdrvxbTPqIBWhAiVjZIMIVc5+VwU575XVAY5
Gu8SqU0ryjAkkLJZ1MwQJQdQFjQ18u5NHwQWlccnkAJrKl5fedBnmyXByWrlw440wyraJn1El3CC
QsYd514wpD3U4oeKwiPDEGquAUqYVvBqOR3p0mRT5i94FHobiAj8p/66uIFrP/BTWtACeXp0ZFRC
+Gd3z4mFLj0cI8QPwqbs8rfcrmw6M97bamaIYmKFsLS7PI7dFppQs5XH5X5JSSiNtWt/Bitwsuv/
5BtOj8dFP3P31T0Tm56WSRF5oywjxW1O2d4kCsR/ZeSKgx2zlAfc+qEqt5ch6i0FoNYQsYwBDZSA
lmz5ttZbDG283enLpK87NOezcsNpzgxSLq2I0HabpSuxHuErgGcy4rSewqOG+WRC0pITZ0JJQwas
jd5fKgm/SX1lwJVHdCB4NYJ6ogruf2VF6woZYN0x5Q3WptCA+gaSgpKdtG3WNnHw0fPKhWiC4IkK
9cKNIP+c5PVQWX/ygpWEHMrYcJBIUA98leDG382XowW+PhvFcuqZrLVGwbdAu6uquwkEanbRsgay
1zFlq9IV/AdQZxnRmaXGHObWrHx6wWq8Qmy1hct3szvzMzRmPuEJtIL+6tQBdK+DxEWPI9osZFbB
Zy9onR4JaUbFZwBaFMOEKM5YnQ2SE9QRZNxpPwPImDVzO3UUwbCDOmMTGJuV9XkOnIEw6ATHhj+3
VEwG+7o7CUlbAGEa8p/tBZMRmCjc1i5UF6QsK0Nnj366/IgIEl7xOt1RrFb7zr67CMjmBa8i9wG8
M+0HGB1aDo9g2DQU8E4JbsFUrvmAPzLocSCWc7jHzALnm3n0i1tfU/44zF2LOqPvhgJEqZFsLVTR
xcubCl75o3E3GBvvDZOmoy1ocfzSZKNdonOFxWe4zBoNmbcZdwaGzGnidqZv+MHRRaIkO8oKDzOZ
B25OnImYqHMR5GKc0V7ATsxE66MA9o+DT8+muAm9ECmmQaCiAwrubHFKzU7TuaFHxpxgz2bkxvwh
X1RVrxkpyOPOm3UyZ0s78JHXo4ZOmgLzkR69jGLb/fuio4IBSOAIIWrZLc/5ZS0vXLA1kbIhLGCh
724yW1feJeBk2fbB7cHatyjW5SZZhd2ETfCM81T8Uwonebhi+7yvN91bxfdACVUXRi1oK3hHfGLf
vCLwLjHdvWkTK4ZSBthkme6Ft/hyTx5LYhgk74dyygNj5EgpPihGNJtjQ0uFYXB6hb4Eas6Ho7J1
aYOA2ddL8ZhBnJ3LXYt2Yw0ZA+ldtbdH/CbzJX8VOhsoxANhcMF2MPafZLK5g0siamWvEMI4rCqE
QTFMD/vpg7PhLCAITCRmFaAk+eQrU08uYigJn7IY5/MqlPiaKtQliNdyM0CBzubWoP9g0Oet5bQP
8xNIea+gOrLnsJVJErLlnjxuqJd90Boi9MRDCu2pwsmXjhGQmy9jKr7j7Nuq7L1uSREFVg7oRe57
+PdqMvDN7G6YNwrDqgKYWaH4JURkY1qvZFBJBlSIjKtHtMjH1ciDhBNve+cjfU1ny4YrSbFVCxy1
XwXhOrrQ+hxYwEkBxbl93tMpzf6rzPjqbu4XGy33Ln5dhFGKm9jmTvCEst14mhQanSwFB6zyPdOR
W1NsRP3pkgKodFaNebeAJiXkezvPouYOpPuEL5PCGMUyNRZHm5EN1+EvhN4Mtt5sY4RXVFxxDCbE
c4KEyfEUKs0Troi4WsqULh+v0nGsoQg7sX5rN75EAh3KzKqMxD2+y2dae/UY6ezNdl6ghPONvCBl
inXLgI2Dx2/C4wsJVLS0U5pU1kSnDN1yvVT2qmM741t/hPu64iKZUOdHAIXSPGnyJeFiLWpF8xSe
DJd2eT62ShTd+o/o5sQ3lJ+lh5Revbq7b6IN7Fh8mOY1SxgUncXsvCjwsWy1NNQKSbMDIHJDt2sW
KI5YXQ5DdsqXy2KqyNxxQOYAwGwK15Y98O7sbD6MwF2HJ8K9cDNTDti1Q9IbhWp83hfdoHoiKnGg
f77otQ+ODPwlguGJndn/4z2nxI9ZKR2Ds9/UWKy6XFcuDgTE/pc8pqxf+ROqGnlYP9kgyc0KGeOe
JqmWil0gif3y1mMvfwn0ONWK/Io2VBENsg/YVdAT804p3t2haTwpmFlGwmhKvWVxldwiSDkvwVWU
1vLB5CIlVhDqVlAd2OaODZFOO8wooboplr7UilcTp5luQSfJT9PzV6hILxyFUkGaH5+obBO38cHo
B81VDEzKBmC3Kz2mWM36HXkSVSISJ51ieMyjw6Tp0CuwtLiFFqpyQRGj0PQ89ELuHq1OxqySuHyw
EdSr+uWZd6SRLp57ECvGNFY81jy+ZY2/2qxtLDFeBZ87R6sZUdp9nUI+vp8i+qB9x5kIn3N9sQFy
C4kjf7ai67IJ43TwfBZUHuz/kn1Hj+rIChACofo8L3dSxngkwTnbz/+ITJEDTMYzIDwAV0GmgjF6
X8ft7pk3Fgwl+AZPavvW72iwgeBikdX98EK1zrSL2ric43yV1Jq/Vi5UakHTmzzn54bafvAHbd9I
FDyx5XYvK0jsQJN5DZj4VD5A7xuQJDRjIPnyDMlaTcWMkOlheRVO4cInfbt1tTP1Jpsa/W9BQ1Sd
YeocFzRuQtJvQVVvRk+W6HCyNY66BGzV7aCOr24qGbOOZgqLaD1bOZNOyIz39xepBzvacIObwgZe
cmb0aEAWB0XxT1k+PACb2aH+4fXM7bzbmu+DvqkXAAqTp2z1yb1LqBEQdaE0aywAr91XCqc/TUCH
acJt5K5GGCOYCnSeDcgL4dVROVFUEXvU8TQmKcSqFYSvKtBEdMIAqiEzfC34j0af58ca66VJsbhv
+t+8iScvhygZIs0d+1UkFdQjfqvwt6fMkrapQ6n2r6FL+NRM9yXBdBvplbNC2ZjcVAACmMAWArtT
4E9Aga82oxKuYwWUdmsp7QDbkGh97Hts0GEzDbVhx43jWFn5dSGLyDeb54rAMsieiU477G6cu0W2
LWxpngABg0pQ+zWlrO0dqU+0FgAtjpchK57IY/IGv97iNrUcmo9U9MQR8GX6hJv5EtO1AEHAxPcL
SOwTaIpPpLWtNx8I9lh7ZpylMmHx82e10PfmFsRDnvs0gKMCTkS2ABO5JdWmzX3lmz4TmSmGOAAS
ynd5B92JHmXxW9uPnOo7Zp3mIJHhZHNBgwJuOHlH2q3bhcm6CIR8FrI/KozqKs2Ca/xIGWWrqmrn
KuiwgRPtHb82KMq40azt7jpVqSx5mycHnuT21/yz9hSvYKxzAcjUjrEjjCXCIIEODoj/kTnczSb+
nnzplDnmfsJ42mUuVMTcmfLuFex6IidbhZXt8srQFFfnA5wdDnCqFdyOgNrJLm2Ga0YPcfa8zIAv
nI5Yq6r3uDGrTrZrOoNNUYmaMZ6inQFv2QbBzCpWUMhpdL1vjzmEa5ei+SC4kfndeQfOVjW9cByl
8fYn5KDj4PMk8iUx7JJJns56qP8sv1C4T96DI3CNWMq8hfl6RHi7J+I7y8+YOBtMvNoNSLWjQFOK
YdqgxMMT7ehJ6rPzzFpIg0us4r6eJmdkH0JDLRdRY5BkRuKTDOmcUMWg3ExIpbcff0zsXtRilPlo
yUbK9v1zdVO7FSnMryMZ6yJLZuWszxbYjofqo5xx146JSSwC6AFNaMLsJtZlp2VFuTf95/vRsNdH
oOlh+nEskJnN7aXYKD99esJA/Q9DxXsGg+yRvhH/hd2ilhsr4PT9dXpKyvQ2638ZVmIPffL9dvde
3himyikgpYov6LNI+VDxoz2EaljSVqrW+DAEKYl9jv3C+Fzgkz1Eg9eqAaXmtQkrPdgWpY02sFXi
83+OTHreAnOYx1gsmWEiKL4voU/zCI07FltH1Y9GWp9BNGRA7l8p6O2ggMK+JKldvPRsy3TYHLJp
SmGh569rLkcHShJAJSHaJHwDrKJg9+xewQdDew3ZKusHxVEjsBHe5eA74s2NdSMHZEWNeQQmlff0
WsTvBIO5KH/Z8Kr6AuIhCYmahKtqSHgyQpPDKfGjGyE7Fkm/53LeV2jH3Vnq5Q9aQHTuGPL1WE5G
J42f5e9KxNImXQIh8iqP6oRqVJit4SnIcGyCHX68x2EHNEKmZmx2W8Ep/CcbtPj+buIHMixwOj5i
wRjMPnmebxl5ZSbmaztEpXKGMVPebAmcPhiHQDXWzSWTcZ2LdCPELUkIpvvfEo0mG2czkaEblPRb
vzi0Pgp/GRqKEMKpvohRzgk8mw6GV1RRrRZnYVilIm7nXB6eDrfxvcAFAYcNHxrnSQSTgyi59cwO
xbLsKF29CpEvPb2xLxTkhfQsYVBmpBbYTzdufKD8pFcQs2uJ6NM+t3eqf143BfG6aN5586tKLVEL
y05YjxxuhbNkBDYpNbVRcD3Den2yZqMDN3Y0vkyLFX8S9Y5JlybA7Sann20xRqQi9JU8o1V0zZvA
N84QHBi/2nJt8CeHrNiXXcADih2s/TAPL82pZrOTE1NZ8viBYiqDLdtyjNSp6txkw+hVQqIAsSvD
M+2z+6O8rIp4RThFwQNGZgLekWZqcn/o6r4UMPTP5+lA8A8LknFI3EEU4kRp1haOavLeiw2U8CXc
1bfiSVkBin1KrtqVPCgUQhL+yxYQpCEtaJItNjdsZHprkb7jw+otpWYACcJdKomqeepcKhEjYLBR
2T9eQt0YccdgOdZpsfAMkN9q8BBSV17zjlGTysbMFN5GhMI47cLK0JUN1cZJkfoDcfqS1rHNx4C+
tbpeOMIZ3f21HRkGBKnA/NJweKsh1n7hfORaNJfoYBlwPh8tJHklkg9+HC4ziBGrhNXL2/MvgKHq
v9Puye2TrIZqgYilNaCRtReL7FepGM27L2MFj8I0G5vPsOZ/6GqVXjOafV3V6LOlU+fNBmVN0NOT
O99SBYD9vrxQKNDs9OtaCJsggGmTSVGwtYB1BgCCHR7aOppdVCKi+3AfsJHQhKXRMcBNn/jMkcAX
p+U096+FEen2xecL8rFAWKNCzhWoRYVlKfi1XquJB34/GOzLc/0JjfSiJnO5ZVTm+Xjam6f6gSHM
w6eypTjLbZs/ag1mxN9z7QJVTNTEWrQ8zelv8Uf5bM30vv/E/cnIWlvwoWsVdia3n/vTKrGDDcOa
JQI5p+mBoJvrcaJP1Q0S4kqXtDkV08Flu0aldRRU2eoCcs6Th3hQJVRAe0pXdumqrORT3EVJ4WBY
Bn/fEhjR5PrFbe8Sw8+pUuAJxJLi6fHr40uDGH5cbmemq9gqF+LPh1rfGZ9Q7dzm1endEcjFCBmc
dSYZSLse1P7BvPGUaP+gvRCtVkmur/KVyLenHDfabXWtCSmqxbQAs4LtqTfsBH7R3jEobUKyLfi3
b2Xxsw0Hb9NxQ9ccnDG9NDeLzd3Y+nR/aSTFXiJqLC1ZUAqUf0emQ4TD1VPv7bj1yyZucYZQ2GaA
oBkYhXYkLUkMO2b4sNKhK8k03TcA9ASl00puSr8Z4nIk5tIs5IKvztwgqzt5hfdHqSKHURbl0RBl
vJl5Zsjt10I5QUpta38BmplZ591CE7c8epcJXkLC8F3D8tTs/QVTpG3dA3wMld+gAQz9Z9pcc3Tq
oE/1Wi5j1a9lyleE3T556ZfyZw4n6X2yc+xHdc9iCW4CiR6KBTbkaRWNqwEY05dzMks5A6QROSxj
IT1Pui/IWpp70oJV5pncz7p5yjYQLdbmPaY2q7INVkLS/v/G1yeshda7IBcMfjlYqCNthId+LVaC
JLqCe2sTc/VF6fuju8uuBcxwDQR2BnDsOnhjzly8lVIyGJi6ZthL2L0OGtDaLglxyV/MYXpqH7I+
wgPYOaCY26lP1Uj+K5qoPkVpysgLryzH159XAUj3bvp932/ItkxnNwlO45H/U7Ps23VAX2iZEiow
t8AlkwbIz3/3HGjPWCe8/8BkWWJYGoY01Lf6xHZNw3UX9CSuvC4e7IV4bXPCmSt5SmVLBsnQhWub
ptpE17iUDA29Sw05o3+LhZb6QX80MTj7Dkzs3Z8WrKkjyBgcTHz6Bo4QgEmfBjVwyVz1CtAYVFdk
1SuDy1MA4bunq2ZOierL5eh97RnhnAZZkjLAlaEZp1dn3dyaWrlr+E98280YaOpBn5J2d7Vxdg/2
XyRL3wmlG1sk84JAfyDAN1AoSPLzItwEMKypI1WRxIRuhf1kT4YgzEa0k9oRcHaeBQPkMwyZtRGH
BCLZVwZ9aJwVvINWsInoAwgUocogAUY/6NvaH9wL++H4FCO+DbL0HGaALzDzvf/osnP0nWtETPLx
+peKO6MYbqqKQKGzqU/DTzch6wWCtp6wtW3hyt86BYvJQ26Al9/y5dAU/GbGvEhtweqWAFGMQwv1
3hMXRObP8RbS2K2Aj0iCgDetAA5e+xxYC4FXhbSrEov4eEBV6THQWDuSMn33zy+/JyK3mcYKBo/L
PKE5rwIpzAnxtqV0Aqm3jIs8maUy9cHV9jBBzvxVsOOcgfdK5Ph5grlWYyg11CtBG+pRw9JID3W1
d87+EfxHLO/m8FZ+kNRP3urmDFYddZSdkW+9M1wdhHSSQaPBo7r8YSuAfDUQgv8eEhRBuOvPVQdC
EgJ8dWcwsSzdUfSbNy9nL+0WuTxKiGJwIIQY4TfldPA2j5fM7FV1VGCueZ83NmRcSG0wvuU3hvN1
Grb02kQXvKgJdgB3gtKZ7rtR4BzkUYTt8YlWlNo+C9V6eXD1tKTYEU3rNFrJ6Dm3QZKWSBsed+cI
javug7K6VDJn0tnPbotS5HehIp4PmUWx+mRrwjjRdAjV1wbzN2QIoNNsvGpV1bGsxBWYYGr72eoW
f9uGU9qJ7uBytnKOyk8RkxHzq9AtzHN7Vn4+nrhrPo9RgyTY4RlDZFHmCDm3j2rwu+JobJxS03Sl
S+tesxUAxQ2iOiLZAM87s8zAjzeOSeJPDlRvPX3eGCh9Qhl71BDB+2RWs5ijvGPiN9NcypGeFUcz
VXHRfjMYyJAleX9JY08kvhXPzQyoa7AXlLcYfOZUebqF8+02f2Y9YlQRkgilhSoZxkMrF7ghCBz+
rJp77i+ELSJVm8xcmsn5BrlUXgxJr5OvKeyFHWRs7lhTZKfXOILWYHDezuh8/KTEMdnMkEKInKjQ
rE2ViBoDkTumbQrvTzTL/QkeNRvYZdF0waAPjozQChjmiBOMb9z1TLgOQfkdjLmp5lyMqI54Qgnv
x+EP6i3kMZaWnImWtd8smHzyHXsRsboCf3t1gvcKG4bwYJ76YhzZrjowe9RbvpPJ1woCZ4Bu0J/P
w3BHIi8KNj2TRR9ST/YoxkXO6dIn0ZDhAlatMS9z8iIFy/eIB8j/mm+lUXNrCnJzYJW9/MYXXPZ+
BN2PSLgF7X5izOwtWxtJGLPtTx1Q/ZUbjjBVCRSxp4C8BToR7Ti8eHUDPQJWvWiNXai/1LevpSJw
T5VTvh4KAIL3MBl2V/mP4K8oalQ6gpujRmJa5C60fj7VjbjJeKPSen4bGFRQe62Lflr/leTE10vs
+0HduNGD/3GNdrMrhnWZkSP5l8+2fbb6P8fNJjI5S7UH11rQX66oMjwx7AnXjij8tBAWWR8NWG/n
EXRxN4U2LfUEEDV3AOui80QyoKN9YQOzz7Lo/A8oK0OWk8PJw2BE9UoZGAoHCx/wcs2WA0+BrYJT
TLNITOU8YiiC7P5uj5FCncCYBTjiutz+qfOhV0BhncL3oRVx2ezrDrv/wMp7YlKcR8ThAwhWBTK2
1iFqZsMOj5JJUXWhz2LQGBj4Pz7JLrYUhMv4Yzc11TOQqkhpzd21zj08icPLF4MfVabnWXkXCpBf
BxBDSYcz4Oz4TNxisw8oxMPQwGdUaDGi42S3Qusym55qT68Iy9Kg/jXVIRgciUiFQZLk+GfB1bum
dNp3WYetSGZ640yjUwAtXZqaxyPfRST08JowraxKbwWBCh2SGXu4t5dOETq93dYVKoHksbo6RbTZ
EVuDTskaVKgSrSuGxYzA96ZsYDFsiXtbNuTsRPgEyohgoVegqEwlQgh/uDeu51hEantalK3f/i1e
0C+GwFfgfM8k9KbJmt2PBZjtWLChEorm/x+vgQZahAolmDr9oDlXCW8YQB++ZfEzZCkEe9mDfYLn
RpJlOJcbkxcLLFliLbnI+PjRmVZ3axoEdAMSER0TW1AaQs7Bz+8sjDbkfAsaBav8JtpJLYJUgWfA
Uc9ctaCpA2mMrk4rGfpHjwk1ULTDhrAzr4hKqe4afVwOSefZyj+cF2S63uPt7LTsM+ogDp06mebe
mWhRGPmidorKIosqlX/RO+yA09NNQkxrvi1Ghnonb5qqXbrxImuEBn16jI5b/V1k8ga8WuJztrKb
eZbMqe8C3vAoBbFzKNHbTKjueyE8ozTCIAhQna1OO7VlP5U32nov3xzrWI2fQPLW7YGOk4VTBdwO
pm6g3Zs0KoPmvp3ki52dNuxYhh5i5d7D+TwDEizE7wrlcvd1QCCCY6zC2DdSe1OHZ5Q/EJBiajX5
j4eIubBhm95pD8Db8qxldrz6EWJQFWVxTGb+ZAG0clDSZMJBJe7GnFn7BtXs/ONrEfF1wTLoKy1a
JYKPmDl1ZTLoyrbVWJvvRVg1AzKe9eW3ZOqitEfMkXiolkOdnMCoLemwjdTr0maofuSgLi3wfBTH
T2hHKd8spGsJ9U65Fa0EMEKABCPf+5sv6Bpy1cAy09ueOLqyENrBzf4sBo1VZqHoEVZU4LG5DCNv
Ih5JAow39UMq5m4KhD+ziTA19/cWPaU0kO85MOp7RvoXTmQWmDB/r/PpccUvoR8sDgbyY0flrrbE
yo3itaN/nwJh9BWKs0+6+00Yj1dOAcCuR6NHu8piZc08WmaIfpaJnx42ooXBZTUE1SrSdeWg31OL
DJcVvsvGxIvSl7bKcoJczUPJ7+qkYmK23YX2XlBqLCklG7y8LJ61AIcSD6vWQGm4MgWFvArDNgdk
0xCTocANmo1DmUYcjyA9Y7yJ446ZQtA8psDn1LzdgXQ2wYuyFL/mhSODl3CWNTsx0Y6gczYvKMVC
0fORCBGW5GQUSPMMHHEDJ7qqKwyfHCf+nCWqy8UPWQsjDj7o5avJn8ax8hkiKO1sQHeaRMnAG+XC
ZSBZBCfVrRY6B/h0OCdSFLRyb34+bUeYRKLbXRq7VBGRfHOO3vF+pr6jYX/3TjE2y7Plp9Javnf4
kxYvcqOhhlH11+wo5UJj6P+8pQws1eN8RODvzxY+a/MP6kwt7HxZN96ldmh4zX5WqhMCRDmkFThU
RzNoiUcMvyibGZx8wB3fjSm3Pac98PI+ft2G4M2antaFh7NdWa3/s+zKRxsDuGVfZHY+TnjAll1w
XPmAV8G8UPMyRhQ5B5Qw6mx2MLXvMg2lZFhFTOHUMSlHyqz/MdIYjp0UBHUv0IxVfX8WnEKP3pFB
ymrT5wb01KSVWz5WhAABFNimMRqSUxXfa4vDnWWOL0+cEOXV199G9TWbR0FYOlEf8OICjEuBqUoh
ZEIEW0b37HjbbU/eSZKfo+ssEsDbzh4JC+Fc+7rPAid5MuIAqvOaJA5wwztkjbOtAGm8jSsqsoCN
c80gc3hYwJ1ALnak9LA7eoSH4vTKhO9EnII+ZmZNIKVcmlgvlYlsfwDAEFNnnABtc9RJsiyM/M4W
ZrAq+dUY8tsNDpCvrIrhQcyKZxSzYiSFAQoDF44cIlMLvb7hR3NkzCP5Hn4VsmCtyQ++sMrVqV//
4s69KNcldnb56CVjtKVh/rnKcRwG7LScowaP8QoOSB9yQ57y7UqnAal9vI8hk2n0e9F8sA1jhxq1
IITMW3yTi1CFYdG23o6LKMXL3tzB8Qvt/fNNzrFZ64MIjfdeUp2PoXFjqweZGDM3zMTpk72Ujhvf
p7d3FXJSJkf81Uo77suq9Z5hMqeX6Uk1iN5LpYpzQyRlXVAAZ1mDc3XNIueb2odSTLkAa7r7gTZ2
Pg5UYonMm/V4yhZzixsmG7P6KQxdTl7FIiMtRUm5Vi/o1ly7JqVjAwNbvIi+TgIgCxe3ssruEoi+
mvSzIXg+Aa1ahD+m+KNIWkqbQFqwRl7GbBVvRIsglKzp1J7IzgjOUtX030Jy0puk9rw1G3GZNJ/g
2mkapefXNvRAeJDMO0XZn3IzsaPo5DWu3WRJ7OFbKSwTLulQABPRgFjs3Pv1pFwH6M4NkgP9r/2y
t7VO71LCyVnQ9421ME3ihzC2l8rK0NWFvOAQUYmKwS1QUXOHlX0tv/drfsCjIieSeKQBlxOxd9Dk
5/K2/FyexPU+cfScTKMgRBPCOaKYFgljtRGy7uVrY7kx4vWwywK1pmRp5iJU3iZqPgGQnFJUgoNL
6gN6zFurHZVjITtut/p3eZMVLI1VOtDL81DWhb8qjKqqQvi2wLnikymvUUkbbUfQ4p5dADsNqprz
0EdHrSRir3snIJi7gEDD0KNgP34wGzypMpKp4u6oV5LmwgCWwsLhiIMjRKaK5Vl+kCUbwo5xTPf6
HzPac0Z1pmuJyQaAsiTi2lmouApNstzNv7tT7iwkANSxxYo645yOy2oke+UVIsJmJUyYxgsMkWIS
jrkDJfX2i5yh4E4NNMckQruV2O37HMDvYr72EyQw1N47vB/VsZQveqGmjjM3DhHoh50ARp5xQ4iG
MZ+f3bh8dGe1fLKCjo0XEH0xhGxz0bk3XMF9pWm9YFrfb+H5yep0POGXcXvYyz2Dl47VtGEBzu5i
tY3esip8Zt5JPyKtcD24CHplrkZBBn6qekJNP2t/AV71/7qOHuui9RFH7VHf4yxPyI6Qmie3rsJb
kwCQvlcwcIFLLFN6RCzeeQdxjahD/NDvIxqOIMD2ne05o2dKRd81LfWRgT57mvbnthqyQHqYAo4r
I2jWl9fLN9sL00vNjon3Qh7+2+vPlYuHwj1rF+DxhO0J8xIlw/DidZAzPv7NDfWA2NmjzzxVG1bq
h2nxISDqXAeKjHTXFlzxQPqGPOiJy9rZIRVBu+J8lSWHOK4EAhdPUciJIe2cC38a7xuCV0yRNfwu
kq1V0BztLV/67NpJomT016WUdBg/oaRplL67hcS9BUSyNqUiKaGTZahOkfX/RBwR1G29Gt0b36nI
BVkH3ND7wE0Uqdri6TBfKqkTftKxdWaKfPUJEdtHwEaBUp6gBfTxayZjBGngL0mYfDpWQqewBP7x
9ymJBz4qjzk8y9k/5QWjoccEbbRyKpiLQA1uex77YvL/MwhEjs75Woe4wBhPJpK03OCWapbGfW1S
cHfHJMoLCmU11EzO/fDoqb/+uEAeJYhJ2JrrTybZT9h41zScY7JlcF6WITlkSl3DAzhiNpkrXt0x
ydDlMt8goy86k7DSeKjNfYNkEW92+QzwrafabdKO/aDDoOagBE3pZe8IAoHGqAIi6rZ2ZdLT2SM6
JnanMCOZLhmGb9rrFwGkLMMNI2YBx3CE9QbFz71nJVyoNSRy9rXLReq7D+rKtQorMlU9AeJeyG1D
cWnjWKnj9ljh9RivzpGTxytaHI893K24TntbPXpND8vHFzwmnZql98ehGFzGGYbcvOCMdecQRdYa
1rubv5vDlbNn4wDmkI2SoU9I14av8u6TROeqYVLF3fxsVgpvNmBWGdbzWcD7e3WEYwMlOFcyE0pL
/6CGYUJ/PPcug83MjrFRKS1p8RAT2vnraSbCocny+bop5HH0l97Y0baufs7wGjJ3WbD76bdJa/Mr
Zg19OprMMTOnFfgWrc9cDlhpzLTkjbHLEoqUOuBlY1FQodVebGOOy6yxnwa7jawPfYJAiuyIc7L7
aBTOM74Ea6geKihEhHD6J52OamA6rNwvO0uSYYvWW6+au+7NT/WM19QeKIWC5OPNXafLpWt888oI
GAne47uFE3xArHOPDecr85nWXmYtVwtSiDd537yOkX3kWKgse0EZSG7i3PtjgNChoXjNQSts52Pf
9MnXFhzrdzidMGQ0oWyfbJ3ly+OkHD8efrBa/n2iZ8wsiv9RpoFBGql2um1ixddXDQQyHzP1cTCV
RdqR4mOfFSm5zeEDBoRRwO/0h7lBDtZx0vxM0TjHEJJZ8nKFL1iG8pIDIMia3BOIVoDdx5ksYCek
qiecj8p/0h9ab5JgPm9Y2o5OLJbtCF2vtl3dqNgdTlRjs4BrjkS1f3mzWySp1d2SCG+/r6khWPha
VTWkq+STg5nM68MdTC/K5V/Jz1f/b9F8Trw/v5+77u04eEA4aOd/Uc7PxAGiQTXp3IixzUCiQnuS
UfgG/pVQ+KQFLjStdfVG5tRvvmcMh6OtPGCkTREVR4VSMEvaTt2oJZDMpl6sGdw1KKBzUBNtQy+M
W5SS6sCeLsepRDjT9T8X/o+zYz/l+fmWp25azbg/WKiXuWX8alwfxUxXRGZZhFBfSzb1tLIS8Bj3
keNxaFcKQMe2mP2oEaU4Nkg86uvLxeEaxYkaHEJsyzgxjrathBx4LR3YNIU6NyRsPb42MM9MEscl
wodr9pe0JskrC8nAyE/2LztdwgVFDfUXxxPh/7v9DY2aAc4SUntmqJpgd9oQ9Knc0DmDsw4jBmcb
s0X/xhqWPmkw9DkMM/SgI+rlBqzQ1oCws5HF2yS3BCJ6ulCOP2ms3csmfFOYoA9RodueePQU8zg6
kZUVHFWZCoVZ2WLleyyI8NrT3GBq3xn5MoBlyuLFqWeaCQMXNBhWIbjhhYVqquccvi1P8Ohev9Op
RnYs1WrOAYqQ3guM+t4c0XFFPXHK13Id2OdajIqY6J3xfdNjQOUPqNRhlfUcuQ/e9GNVi+8xRZGr
QHxQY6rWEcXTOpR4UTn16STseDV1kz46qlH7sc/QtrdDj96Y1GnEyU0YNOSkHZ9zyozZo6h0u45o
zlMNCa17tNVSESrEQ80b69JGsbXdco1r9AbV3X6Es1W6gFiHumtv0KAHQlG2fyrPHxq6+e4D3HBX
nDuJNUFpGHsKZXQSKRPsV3V5tcSnI0RyD87zG0xK9CG28PV607c6HB8oi1lwCxeavf2PbdRFYdaG
kBIZjGlok1MTPnVSTpQoQ0jzxJ9h5T5DRi7Lgbf6dBWvDQawIj7QJ/R2wSKM4WGwC8mHzYFL7Kj+
1+Vp/GKFQR/7hNeXsUJHBaxilF56orFmE861XJB1YV3BWCn6HmPujQwuLEWZhFRfNyth3QaZCo8F
aWBceg9xs36azlUf93yzOKXtCtY/mIQIGbvJ6dR5Po9QZTNmdwfAzVFhfhRMvWLi3HPgvUGbngLa
UvyQSfVXxWHglwZYnoT2yzlQgZ4nmIpY6mtrqx7wEG40lUTNZRYggvNqLpIBgUzxX5Cs+k2kPp4Q
TVSc9gkd525cTg5bBJqhx+35yHD9BGJgax7qyz25+ZN9bwqcRdhXsqaavuy6SfVEi4w3OfEyE3Z6
2kc3ao91NoimtZdIFZsPlUy3Z3k3GhM5P/XH4tw5zPToetwOL/Vo5Knk5L3jN465/u/JFUpgCqtQ
8uchmeuMt3ethDce78JHleQCPmKtqWwMICFPRsEFTO5g/2CDVyB94Xib7Ogpqr+DGgs4imcI0xOT
wXYLTek/z7yWEEFWTLF22PYvQ4ktpS6wEcCyMiPHKkLbJQPPD7FnC9owtMSyrm+3fAXDhP+ZexiP
XEJu0LBA8nXzfhfLmBtMkSw6i+AtJ155u6w5G96+AFWtRUgXHaTCrJQoN/Tu5cF8uM/znMXv1kXz
mDU1r6C+fy7O4R/zNsemX1pyKZayfuijkrD28lKdFY4Tnl2lPeei1upzyiAq3ApqHEIPA38JVQT1
GUW7JJtnTwdb+WEFGHqhJ3f+y1QRcM22RN9mrPvDF8VknqvrhlZCsX65SgwvDigbdlCZbvy9MOT5
l2/oCWMbEY3Tfcbg5HjwASY2ENqX4uWN5yLzeQuXCQAYQq8mfSvXjRhF0VcbGJrpFcgeZngg2RTE
UWoCeiNNNlD2PjpqYipacfcXFHWbFtkLgMwb2s5n8N0idABKf4Ev4JXqAhQpRCy7QphDq/ZqKaRX
qPH9C6hjCn5OmwidkowXNkux3uGFIqG9UjmRoOnpjpesZvDyjNoLAo2MaHpCLwEXFKxZZiN8ebXx
2D50PRzza7t3m+ftFiQRLaOwJgDUGELoFGXh2IY00yUsw0Yh/+4gUICpsLaHTgxbJnXan87lwsYL
/XATmbg6dnCb12Dm3Fwpbqj2B2s2BbyBFlrOI8hg/3C0esdDBcvJ5vdXX/F6W8YTkr29tb5wQrEj
mSYlprbESlgDbxbYLwO2zHK9AewJ+T6AsEyPXReYs68166D4wpVHj/sirHh2bSJ6B3zR5vsEt9V0
NOua317fMLZaSzwV8WJnJkeourNzm9aADg2xcX8QWWO6kt7NysW2B/xkQfIiqaIrHiCQyW6w56ZB
KutAcu/z+BdebWLS/NLeHlMVqjBSjaoZBMFGkq+DdPwQyT6/U8qi3Ooob9nt8GKznhlafRZQHd6w
lAWRWvwED0qU/SANp0sVfxEQJgjtVuqm13csdFNJJpIyp66nUjSKogZANK1yB75sH1yCn8ikmaYu
Qk8mygVHWHi55E4PopKT/t8BF0HIomR4vMC04XBeGwC43vGiaQXo7LznCmfqQObwxIT27nNHMIqp
+MqRGY/NB/e1+cTOUK5lGJ236vvKWpoqN+Gyty89EsApPL0UH0dATQhg2gw0TYBiAOny9jlWZyoj
7usROBXDGmmHZSL6O/CKkmjaMg2KxxCOkSKl2NTh0GYFmJwDlHLzGc6YlwPQpIvpO2pEAXhDJ0VE
zXuBUVR/qsyoWxhR9NtGqAPGQqtO5izFacEDxYXc7KKj3G4CD1wnPx0S7ylHQP48iNlHQTDKy/6O
IU5K0YIdUZyeclD/XLX1wyQ5rNUfIg/7thkaja3niWLJZAeIm0nrbZg87Q5fvyFKafljvEBv6Vs+
ZSjHlgmvzai0Osd9c+CTrL6MPsFmVs44shtDeev4iz8b4SyZq/tvAX4RX9NSyIzxCpO9Pckchshp
YZq+h3e1Ly8E55pmdhl63HvfDx56AP0zkNdHvffq2dbj+IsZlgq994zhzTOYjWeD7BB2CBfMzZvD
je9I3Y0DU/HExnzOqWKR9GovO9mvceWyHCLcbkyWMg3M1aFViyEADua+XGa3F8TnFFRzoi728rAb
3OSOu6iY0vSrrPW2xzTrTG7fjXkTjG5Tclw0sn05Hv7rIoLad7DYnhJd+mYZqe5wp4M2losoSoCX
q4AXs8bXrikrF/94U26AncQfpprHvcztBbiGdOydJMnuhnZXE8u6oewfsWDqteoZRfZCuJZulCmZ
CK4ovlUf2oU25CbT8S+lW4Sdo0A8k9VM6e8DTLcA8D4HA4sa9uoIbaGy4co0OLMk3ozFd6uoc9iP
iklKlfWfeK1Kwjpg2odRoFYMeRkUBVFGKgQOt3GdFd7mvQ9gS8ozMNQBL87zP74+0+GUTPw0aC9b
0/6WpdvjtGRx+5jAiXxyrre1AwPnV7ALm1vWLIuAzkP2rZFBCSRBmqEUPaaT1+ZbfFVhpMii4vMw
sPSNBvcglRc0v6uchqXepi5fXNsKKXJNwc89SeHpeDCZUJ+USME73RpeOqEjUkUMcl3NaareyjUn
ClvH5tTvtz6VciH4GKklzj2zNqgKJemZG1em3q71GYsQpHsytW04U3Q+YGLOmuykIA9Vxtk3Rgfv
Sw7PCYQBavRneJNej9K3wj7dnyxc/wVfNX0G6Gk86HUP13rEEEiJVMpMeJtyqZx/YZXRC2gj3a4o
GTeFARty9F0V+WTsvuDqGNV05LsDS8Gl5b9XOQut+cNOMIIOK0PXcmsICMCzxf7nQrPA6M1ce4K7
1P5H6MvlWTIM9becYyt3/7gb8UvwVIlp9cBIkkDt2o/i7H+8j/8J3EE2mptyO4ThTnCJENn22V7c
7PPhR80OBSsMFFq0aau+wdXmVtI3JjB1/s19tFMEzbQD1Z3CuA0FwUtyzDBJmf7Y6wEpvl4rV3yY
JMkrZemt3JBj73XH8Kx99PXP+wwZ67c4R0BllLc+7nc0W4DQZBEBfd7zWo/ktKytADT6cz62mgtA
whSKbJ31Ie+KIosIuTl4BN5NRz9ZXby24+VaAEu9Q9IIfzz6SIh0sF3TqeUWYtQVtCyd65MYTBPM
LCg80unZv97NvYy7v3EacVeXsPb3Y994h2hlCKwciTSktc91qPpyqdGKKUYlOT13yZGZgREOtOkl
3BlTMWFRaaYki6WFGvqquuCMCBhVQxQYriLSHFIVngM0s1D0U4BTOgknMlDWcBves0gKdpkf9gwX
17XEXux5v4l8EkzcV5Vmky9Bu+jFQGBBs6qWJ5cTcBDGjmb4tB//XCNA5+gdhoHv24ZaKrRMu3tt
/hLV6i27J+5X1tyssrY6AshxlrVDZmecP7Ng42R3vk64/eLyHIupVczGWItwYrFzAr2dsoCNn1iM
P0h+5zcRZSPyNWCHCHh1pMIK3wcQqKnXjidwXaBDufZLKZ2t9ueGNIYC7CeOWNFfIPLKWEqGlFUS
FmLYx0elwJEzl9RuXIlOtOjYRyqeDgVeOFChtPIACPOhQ+OhTP4WPH4NJmBR+KY3Ys5EM5NwcCzr
DzUT1co6ILg6B2YVAifrvaeHWSy+Krungui+n+RPEibtaWmQN1Fb5UaBLAefnE14t02dMnZyLpDn
b/lBP6O6ZX3NONdDH5Rojau/lIte1FO5BtcoRmS7p0S0uThfxVB6zMPp97BiObYnzu36jyMv4Xqe
jrktvoeesCXSiXNgj8jB4bk/Xfi5bzvOyTWu3uvt3cy8anml+FsjqNxp2SecEM+uhNesWcgQespr
2u8tsWCbeq+xkdDC1pmfV7aMg07kqivxftPyjqPlh6jPKIZToEtxNZtA+va9TOezPZgorEICpdJi
oKwjlaq5WJQLM7ePBThxfaTciFxTP894PM36REAAhTfgTtWK3uz16cJzDP5DozIRVepKvdimAopt
lgDZVWpIh7RytZcH18bvIhUG457r1cRGcR/SK2SKCBN2/MABqnTX64FxTo7lnaTUH05XXmgDTLOp
010pHi9/lTCfTGq6++UcVEMRtV7ZvsMds6v00PptcnvgfvKW7ZC/LPDuiOBluuwHBhPUbLEPsWik
ZZPA9fYBwEGPSCNnPu/vSLOrxtPKbr6czNov+TeN30K9sPLQOVsePxrBMh+4AwZJ6Cli7eKPpFb7
ukJJme0Bbpt8CCUsOwBnNJVoTQjQ/gdbkPnpyE+Kk1PMt7gH2iGwuH8J9aptiwzfCXMS9sfV240X
iAc32X/uRNOy0io9tWw0cGuBLaBpC8GBqQFUAHOsqzW9MO1atA2mh6uGaUjOdVyBqrsQJa1YIYrI
Eq03hQHvLZHZJFabwvbiydc5j6lasYBCtJUwpEqM5cIZnGlwxezVd59qyDz5FOnYWegqzMk/rOiZ
mprDort7jbjkQJhkYD+K/IYPBejZ9lehDi/uR/WSOJR7BeNBPRDtUFlbn6Cfu6heTWlMYr7kV4b3
tASxvRn0uqOesfMYyIpykAoKucT86t4WYvLgRNseRHQSLS8t4knnbotit9RaGYGFBaMDk5fQQm8Q
z4VERzLcfkm9h6tiKt3LrcLqNnQ7CxZpkZd0AP9aoaoEhqWvE/cHOM7t6iN9+QeLCvmTO5iwDbuP
MzleyQVM/AVftfZoK2QGIdrMSAIVHx5qqLAUMMRXI6AAVwFPOJf0pKdHn2H7JTX+dhjz5A5lwD6C
DoUDY7wuVnRb0SgNEghyYZxR1H0hy3qvdBSKfc7RUG4FdedZOxXpFJGX93l2rL7Ad7d4vHzbesGa
/gnqJ6HHL/eXOzAlsyC/en9S6vJoFaCPOS4sLAGCQIkrVfr9RZKYbX53QsKuVf9Ws5L54WWOCDWU
jEXQHS9tp9Ha4kzH5ZqkdIqJWbOI29n2EHtsOJo6iTfN6khj0sTy4zNH4Lb2rB4vUKb7OaItpbnQ
rwSOJHV5ssxtRMp8aQk1JjFqVL31WjarlurZexl+pDST2BmrYuQLwOJdu9bHzM49XYAOX8+WyyeF
gcgZJrdWxiA/C8EimRXkLShR8PSoVd+eLUOCf3Z9n7q5WfEoUskNxxM1P1+vfaEPNlteqoWd8r9x
G0yOcE4LxgaHVK7dRpVxSYfFV1cC91/rQ/H3XPtnN4H6kZ4RfGxuMTOr9+fGjseftuvB10J0BOtT
rUrxoJLzudjS26JHD5wps6DPXAxZTgzFWr8kBF5eDemCpJ243MESK06jWDfijTGqZGXhzJipSx8V
yWeRhvp5K8dNbiqCS2xNMN4jim5Gl+lLhX+B32kAH9/526CAQBN+6LVUgZzck4BU4xZ2hFqzydIo
Y8WpJNikl1Jxk61qIonfff4fFLfQccCUgniJX5JaeiQFU/aN1Rn+S1lBAEKWu85e1VXALjDlARI0
8YTFWXUxZZC6et4oye8zNex9ezB1TglWUToR8OSUf6J/lDvevxfCeMVVWOUfXUepyRnOwQBtO1cr
6GsKYWXYZSS6qYmaPNpZh8TBxV5hHqTBYYPL/gvs5IyIUf+5BS7lEbF37XpX/VkmN8u+a+SH52dO
a1qAWpEBIAI3dZW9CMQJer5MFM2QLto0JpGFbWhU8HObLmX9gNeKuWzam9vFMU2+t10U/KxXkHkd
jkGLjQZA0uXp3uOcsq7z2+sPLLyV1pRtLgcNuuAygLo3POgTb7WEekaGa4yNm45LwtUdi3Ff+al/
G/AQAR3cvrm8T4ImVIJvlaHTxWjyR46+dr2KG/oXTwG0mmIfdWPG7fvOKNRQWpo0XmCqaUiLU92f
q2WjPIeOeCUfM7SS4tdK7CNUNOhaCndqgeTVdZojJc6x9hCyx1v9rqFTi6eHNeymbDzD0LlYZZq+
vkmoPdlYpgkuRBLtcwSt6RksWMbLB7jbc22RywZKirfbE5pMf4/hYQzACTf7n91UdTqTxHmFDZ5o
8kYKg9eLcptkdAB5XUWfmc3K6cwbOgnf/w765e47KzA2KSBjehJwDaAY6u2F5KCpgD4LIhawkrMr
55Dx3HOAGmZt4AF/9BekBu3mK4OgVsluWIMNXz6oDqpQM1fE4DeUB/2sahD9NciygsXby4WKbZRe
QO6CpmdNgJ+ERypI1UDk4f0vTo4gEW9KQ2Yjej8lpLWUVAKY4fJHfIGH3kX7BMJ1j4JO0BmgYux2
SpqoOIWaUVjhMovyh6xGi9+jmiIzpztCzNBf8P3gX12hoLQAh1G8Urqj1l4zMCjYye9bMsUEeONL
SMLG48U+2trZ/6j+q9JMuyHPFdUTKlgx3/QVCSR2G/Wvkj66xV9Yxz5s/Z1uLtr2ag0d4q4ngL8P
Ar8W3tscELwyQR+xxRpVOrErVmpyNOsq5YK0z4wlZXcJtLOoGgQjfqNk+/Y5L5/Gt07rkkTo+Dwp
YCLeHURfapZqqGWHuITUw1Chj0XztfGcJM1ZmxuI/7nXNbq9mRB4KIcnATHqwan265+VW3OpTZjJ
LAkwmp+UP9GMjDt45lC8j54j6ngzccVo+5Txc3f/QX7e359XZZo9ravzF3XEhjBtWd9ueNGY2/Wf
bKqkmpVCzK11nMCTirxoUlayZg6y2JBWNHYZZxNixpUp+XWO1r4YUaqWlvHeeQyUM6WJe5dpyKu+
t7lwsrq0qJ3Oz0gHlNwNLD6P7zcI93SqFfpDlny/0nxUJ59+tPYglY4nbGEti2JhTAdYO2wHHeG0
tXuBOTMQBM+Bo1KkldTd2DVuYFLgHfz5wLA2OLhhJl+hV4+14gMSQi/xvSZ2zHA/sZSmEtIuNG4a
pmCzQ+t6B15HonYfAzorCbXLvbpSF9ISlz2PLdBs3cmRaas/Xb2KC8fVpxU7rN5qy/LIUStgdsCm
hRkwMNVU6+4r8P0JreKaVVqiYN03QKl12zWpCIvmk9O57EoDiwmN0uUe46B/AMY/7AqRDu6rlaMs
PFXDN/RGwHL5IKS3/UEvS5vW9q4z+IGXlXbosPUtcxN6JC4hReE2LYsjXuFFtv0joMpqZR6G1pFY
OrDv796kqbkGiXaXo/7zh2k/BxaFqtbHh/YMLsG9PzofRKChZeuXQw0SQhcUsA2pvr6//6S13qcc
BvGQ5CZmq/6k6ErVT+YZIPHAIodIGa9g1Nwo+vSiZn4JjoKqt3cIdFhmNQ1mjju7Od7wjk+wjeN0
Hft0kf991PKHipZUxEQWnH5zR0FzyXRnLnpNW129WqKTvQLWA76sgpnXEFE873UscxwY6w3RrVKz
jRdPAFilADIoeWB7ai9fRsMKtJ3LXIdN+B664IopFKQ1b3QbItSnNOivU85WoqDS0f/aCNGbSEYv
qAN5aLxhqNhOmmqJomUSLf8ZuLpBu0jPAhVTQPZGTaXwytOT0aMgB1srYJP4Y91UJvnV2U5dRMWs
onan4AAEqKUiKecwbszV1cqcAEE6+ixh6pJA1RSaapE7nkGlA42dadPlHCFnKx45vIN6IZmk+6g+
LWDu++Cy8d7t5mp9Mpuj6rGjKLPgkwoGItXbrDQ7NnEZYax7hwAakBMNmcAuNk7xHbQ922tCdMqQ
gd28srz7YylBymiQJLXkTQsIPJoq8hRDMEDyrfiZTBO58jMSIWtu9ic969oQUM5RFDz6R/JhARVS
LnJmDj5lalMAYOvyJ4xgncBnN+BBSDAKC87aAereLgBTKAfqQLlkKvdoXF/aUzHQ6nf1uYLT/sBR
UGJE4mUHbZ8Hdbb+u9chHtx9QLRyVIRhcs/SskpV2Bxn5l8OAJTuz9B0DA1CFC0Y5nEks/oaZ77y
WDvfhKO76pbP2aj91XUlDBjBmVKHCjF12b1Qsezbg3lP8rqNUEYWvl/kVntXQucOpuGVKRXio2w1
9ssOeLITmF1CX3//c++Sb+/Zbod9z1wEyHrkDOYugblQBvBFuK2y9KwnQLQrvbKIGgdIufDv0G1w
aSYkYcUlHSYgWAOGjAjssP7MTCNDEqP/u2Kz97i5T89RiVZH5dC+P/GwnqbVlKmH3ebdsLLfE6u/
kOVre6XlKXzALPJaCQ5BFjZimas+uGGuUPUBzVZs/YJobWaM27K7cuBi7irYjjORm2CuNW2rb9Od
/t2tWPz6CsZog40tAVMJEF6VHz/6TpKkOYqqPa4G7DhNHzNgXC9OAejfptZaOF0HfnTtZ7wY/av5
PtBTRNu9hDBaaS9PCUF6KF8xAwb7BgTY4jlviJ0jadmgzBHIWulHhwEu49rzxbYnVJY5lTPGCmJb
viPqnia4uMcxEhu8aEMWN4mYnycC93NouYZbaoi2Puc8PvMjtx8HY26LeowIuTEI1YnZk5rrK7O0
+V5hb9PXoI/2+WuXQD3bKR8j9TOIQQCDk5UpZDENbEYORkqhrgrJp3kWoioB1vwxRg1J9OSACrF7
4OHd5BzByfHUtKlK+chH8nkX9pexWMym7wpOm0CAbj6+LSw19+DFnKYo2lpX2JE4kIjIonvn20Jh
qFBordVelvrrqJoryJyUOcWsdH5Y2zo8O2zjfJEqPQ2q/EhXndoHGJ7BhtHLrJo55RTa5Y7VfUe5
IhAyWpLlNHuqb8RPLRSWeutNC+m6OJ4u90tnrp7U9l7g7dgW7jrH+ixUwMhl67RcV8viFPKaLRmM
C6Azg9kUQ+47tyGQzCzJ0jVRCqwvQF2E6Dmry6oZyWMm2+pLnlw2Xvo0nxbZkQnV2J/etAl9DmUi
sOTQ/OSY4S2+GfzjJVg3nz7RJcVhpVS4VmXQxl3FofklaaR2Cx64wXzggTflxxdS21nAHgOt9CaY
KI5BUAZvtUBF7gKspm0JnZitsgctUYy62CCqcAPL1ro0uWHIhyrUmmVq/Te9bwvrbAW5dqb/yStH
593VMDuk1z1BoIO4PS6Ko+uVh6AjTh2C2vkdQ9df4ejxIFYWANHpJlBb5SuMlK7Y2wB76ywsNUFL
BG6jeaWrzmGj14lgk8byL0EtBVXVO3kXTsVqCtyuN5GH+sllTogS07pHzVSdHJRgA8BTYQ4HwCn9
kJFK4w2hSzv3ZypI52kRYbJ2ldbrQBYuZaE0qGfUEQvYMXGyH8oMXSgMlZwbB4Rx5gqdyL2m1Xej
6UCITXRMnOlHBCSZePioAVgUsNrTJzr6VFFxZLtAh5hEKLG8YDE9y8nFMXQELFZeYVlwGOS4Wzc6
gvAgI2z4PZyVAsgVLBAswZtnmkaHQSlnkfcz4m1QJPEAz44htsRveneQd5Mq/FqDKog+aQasdui9
4N9cI9s0FKrl8EmNbBC7vH8/Rn8eHr8nAK3L2YTVHBsyY4/Qf4xQmLQ1deiRJBNUaWU+D/xuhxGw
uDVJs5iB9hO/dTDgm7oyJUitHMJdkyWIOCPG+KR2w7ZU/ChNdiBKtMpJNPyC6peb3BivsMqe1d2a
O39R/WzPTQdA6dBsRbmTRb8VOQaOizP3GXh6VAIeXPOKph6ms0w1ciEQ53JtgegytQdl9to0d7fG
uWaly+ibtMhO5DVzgUbsXm1f5iZF17jGBlPgcx6fbddF+CkgAflIE35X2hjfHVISo0AtFB+Tpd2P
JVomw8vY7i3D48elIDA77pPbMrQm/evjEUovW9ecImSSU8XKNC7JRyQWQajXNrXJF3GsepSJaOmM
0naJo3bBSUBhcu20Npm08m3LAmkzdCg8/0QBgpZ0IOmmugfkHI4aGL+WnjNOPpscZNgzy0iD2/En
URfuXZA69Db4Euf5zXVsaqRh70ReFOx8bUWg2v14LQNp/Yp+RyXZiCGgVDrQdO5i4+vugO7zE5+F
hyjEApPIc1nNJoNpfZa1bqaP6qI82JE6DShm2fLoxPsysrb/0WWTLQc6hDAiO8FZgvEnsDKkF3xN
sCoCUFtU72j8fj/HioPygACJiu1fIExUU/5Yp6IefHbTbEuyAI2BhzDlQP04xtT1s8zykmaIAoWH
bN/SlX+lvsHVJ7vS/bAJj4Y4uKz8+9jO+SM/foW5k68jA/zHOBZWw0eANDmn/WKExC3sLxh40Vy6
mYPWBa+bU0s0RA9ZC8YhB1eK11lS9c5ItSoGZWj2jRBb+aYOoen9RBe6ICvN7ysq1UDIAdqv3wbf
TJLLFKKzqmTM+R/2Ujz6/05foEkbNWJNKPVCFWGxDzxrbJoLeIUAwV9/n/BFccl+tVKxww6do4ca
SKUKtCI3GYjOiWiHzBkI0NM/H3ky9isZ1+hFR26iEOjH4Dq0C6DFdA/c3k2HvZdXU9LgXfLJF0rj
PCD2+1gNmaKzwBzPAd20dFKS/eyhaJxpDnOXrhgDJkRjNvyUcwFPvnaMmW8Xvl3x3IikQj1LBEJu
agAHfvX35qyf675jTkfAjxF/TN4AvsY/1MEgDV7rRDuQypQWCuzFf3rG5PU87CAuj19X5yIkEXxp
bgZKZTl+k94NvLTE+Zcnst7/I/W13xB0alEquERMUzmTkpGktme6pXRJPcOXxx8NDltIE2BaSAuG
hd3591oWVV0MIkxIOTh10wv8NePVYgUZIN6QHpYO/h4SMJCe3Q0GubOF2Wj4OctgCuxdBSmBKTAX
udv5Auv29okNaADn0qI7eyx8EjWYTa9WT2/P6xw2/eUj+RoR8sI1XF8wKID2pHnoXjO8TznoqPbz
79YzsZF+F+ErHM5MYJzImPund7p4N7b7b4UnHp+7JO/FDGSh9m2kFwp07h9aviOiNHAvxnhYczlM
nduAuRxWrA0xiQoemIHZ2QAsHufWZ0CSqI5bDwfoGZSuSpyf64B3dMmjZCIMTn2T17Pl+hY8eBtf
X0i0j5W8uMKG5JtJgzC4z+cYcRr1//nix8CtPS9D1iwDJjQql1foKS8BM4xCu4jCmtzCtZfGXDhy
dLGKHiyDPgsL3eEFiyVqRXMqdOuQ9JRMwxCosHr+aJMbQ2Mkbhg3jLtJ1XUpdfC4Due4ZGBz+FwL
77paXYlDbQcmmefWQ6D9QOdhOv3WIN4V01OZ2pqgDX9x2y2bUkkdnBZLIjb047BCL64sTkdYXGsD
Zeq3Ub3NLcxawiuYhgE890Cw3g4IopK82xV/9UbVw5BVbgojSCiyYs6kzi/+fB4CEaVlwQzd6Kxn
meRB1JwYTEQLqr4SxBCQF18nz7b4a3T7WlNwZnmYgM6qj0mBWyhHLVZjmjLHYiOZ0stfWH2mclPr
3DOGzWrdG33tiBoVHblRWD0ZAla5CiKYc4SUuFkOHdFUOeeLbXUVupnUhi29AsPvOvDzvwhgQmX0
So8e+b/sEUSTw63RRt8EtNa5CHYeXA9+d+La6CUAICV4NmFhH7/rRTQgCf6rVgcocodc4T0h1rpz
gyxWTIwU1L7ogmOgpmD01owIe23rDBqy3YmMBMF2655vTKbJIAx1fdpD4EaZJhZ4udJvzxsda2eq
dMyBTkJe/gO2iAil8Ui3I65lma8u1KiOmPgK9kJ6yqGkxyYk1VAtj9dA0Sf8B9h8zJ/ER+E1xou1
SayyB8HeSOpwImFqLCAKsGUPacBtCo4zlbeQxbUMlqju6yWVz+pVLwitEITOf8sSAt30lKyNpZNs
uPrRLNi8sFPG/x2IXDFoMe/2ACt1Km/eVicXwqZaoSmNrMPxlRgqxx7Wuqk5i85YSlPEIcIZXWUm
7e2vmIHY5O+19C8HKRlHWwjN/Xejw83DDb1fC1+wkCirruwU/wz2Bs+W3rIA9xQ6dtX1ZJjNiGm9
L8TxkpxenvKkffbcQ4PTqt7NWHiFzyNdFmqj0K/TA7e2vY1fsbcZmMx6+ZQSZ5a28TLywHFpB/aT
WhI113RgshLdbiuSrdigUsFizwwamWctGQZmgsvj2wJ7HNr+uZY9K7gX8YryJA4USvaZBjPXQqcp
JJMN45idzcnkLjdpSkQuUATrcWIxjNiD/gFjcE4K5tms6PExq7PDjcIUz2nmgL53n4dZRTbX+4R1
+5Jx8im+/FupCO3Ii19C9vgGqKw/+GXa+gOi2IwxC+LDmdipfro9jszDurR5WVZlHbOIU0dRvZPR
OiD68nVjtJpgZl4BkPFk/QmsT8McYJ0uEGFElsTcpg/Qe0wDrEwFozoNp40Iici4Qj7KM8eqEskE
hJKx0mM2ePMDC7nTAe4kcQ5RtiWEcy2oKtQJOQ9Qd6nU910idyQpFD4KITRuKSyTywnXr8dNmt40
DNsRD6s8Scs7HQgBYyZ024Ka3JAhXqF+45emtxsd8ZHddog2XUvIG+MuHM8by2jTTAw/vJMl74jZ
Gsunc5FmXiiqnN+GX6KNClVuZ92WyajchMS8QKAoMer+k7b9J6esJ5CC+9H/sziXkfCDhW2zD1Le
mgB9rVUU6nBxYLQ4JIuR+pA+52WMM0JA6RTR1VHrI4rfCQDx6bwRRu9HDeWUWxHfXDtGBza7jK3f
CsT5BSiezNsjjlA6WX3YS+K4JZtmSsJ5Lsyd+++gdClUn6QVZqPPdDREsBOS/NqlXOSlGMuc8DJa
oOLPExD2pAqTIc4FZghuf1enFpwKkpj2WRcvkPOP15acnJv4wR7TDVxdTEI2id1fM0M0+82pl25u
xeW1YT9l75XSWFzZnw+B9/5RrQFqtR9XPr4hgstP1x1XSL1vX8YhmbOKoDMg4c+rK9U2dweRW712
GTvG9U+bzW/31NLt8jogPZ6m6O/n1OpnBuGSNYXtvNdgiMCj7as1lWEE9mGTDC0uvfSVnEPLUyjc
S3qd/5h/143ngHMH/4iT9zf1vD6r3T3k53I4Vbz5DT4enJluSIKv6cIiXKSGOm4hmlXCOTriyqVe
EwZlSOz8AmU8lpx6a69MNbnqr4ybNk41Eq4TOQ/iZkbj9QBWQd4eDWPH5kCZ2TiKUt1U2Hodosum
tJJstW/jvj+Tp2/gqtvIpa09DDwdNuack6UfHU00Xeo8NdlubHdqnCiWxQ0hJDubTxiAlg5+gW0l
2U2DScQsn3068eyukSjQ9FMFuFi19xb7Dezr9jPouR2viuQBwJroyNtg1GBxISZdSKG3VCptSFzL
rjuZBjV9vhNX4rv5VZVL0QtNJl7UttA5syu5Wc9jh/4O51aq5azUNX2imch0xrhalPRuQEeYSYsy
Fn4Bq3XlLNsfSy4rZnBHwCmnUk0wgstlMtrVbgRy8GpAXN/zQ79ZaHB80+l8i3QeuOFR6tK4Y4IZ
HHeuxxmg7PG3tqzX+vEWNW05ckW/xuMVs0wKlas5lwfo9R53gtXxEAGBmHai/4WqeY4xnV+NlMnp
UfXYkfJMXwa8Xrqhx+xVycYDbEc4/DSkb0z5d2Wge5x1UPj9PQLsica1NiJ8WFEHcVJ7n2lS7ici
tDePcNREdvaS172F3QDeJn09b8F5L5VjtzlYwtirNSwiahU03TW3wm1TEnpVP1PfE/gPretR5Bki
uLRBXP58cU4QfClplS3VJb2xipjB30ce3XOecixZv7CSVN0URxr4XsZhriHwBfYO2NGWzWuJQn2v
OE/GWhT/DKtgjpE+5rD7Tu36zcrBc136lCsZ0WRXnfNy9/sveVm+J+STxbgPyklhrPZlSpr9Qmuw
1qMH6zEFAPWfh2vtRZ6eKWPRkKiSQHDGuMU+W/xWsEW0QsdJ0UUKE7PjGK2Y+AmJ5CMHwloiNSzf
koriWp9p5wnhYdqXfOQIF0gGPPaZTTLwVtfwi1s6AYNkJilBXZqzrxNprfu+ZSJkCZHPVFiMM0r2
cSW1KqqV94g0O8ZxwABgeLJyZeYVmZWtoTcofL299HnXvWzp5i0Xtnz2wnHMggfQVG2/KXVMBDXN
Ar1g7XSm2ZYWomTn1CDtVWw3JgebGPzm9T6JtTB2e1yqm1DkN4rYe4CQRbm3dMGRZB/i+/qMNk5l
hRVj6ytAN4iGnHRwzbjwqJkePPe7uebMXiUclOnSWVbn0fSx37OliIi3/Gk5y0zmaTpX6s/WyRC0
UP/+RR4mAUVhbBdvs1Ap/GZkQ6UKcf03ZAYtQVMbNCp/4bfqBfm6TkOuC4xQT2cj0+eTIrTWqdcf
9Oqz8iBbIVaLCb2VdMrF4fCRkU2HJUwLjEdjJVgW0Z0GEo8FWhDyCJ1kwFfEowna9DqCSUUtQ51N
Ywl+4AZZFQxao/zwlAvFjNdWEcckywOxzvcLh23qedpObsgVit7RhmAuLadWGd9Qqhbx1FaI5Y+I
5ZurkEbkXIU++zX924+IPdq1vB6EPdGqxbCfICvqO1Em/WQPJi1AWedVFgG+M+w7oetz33Wso8HK
D15+Z/i3DBLesbc2sB2SdQW8TSEXOqZZbtstJIiX+p0XfDF5h1yRBq8fmCjGkeXC5B2x+JPoy/PH
7+BJvgupyY73CdW4E+QuRedZcEXPmcdk+/ZtWdSf1xPS3OPfkns0QUhHt6SKUQ+chV9Mzc9pasRx
NJs8wTE5nQOorl6rfOVVWKMsUTcROH/KwjMVy0D9OFvdrszyyifAiSgB+CA/+44vFGAIwkBtHOw/
kS3UbZspGZ+1wVKBPnA8hH460fYaa0cGZ28HMvTa5+Cvb0xct1eOCNRkNaKES4NTrdMopRhPehf9
auakcDYfaol83ep+nQSDH7q7uZcaIpnhWzzNQEJs757NUzNWZrwujj8vngMpt1V65NtrVzYoYMfP
+kgIqkNsE3pQdcP/E/nw4EgHwgLVlae6eXAJidgZ+5z4LUl+qlq2cRYv3rlgDyr5MZ+QQ1nxrkNM
BKxEw2WVNgm/+zFAU+QtJmC4TQ6Ebxqepru4kkQfD9h7yCmTw/wOuomhnk5XkfifH4nlOMBunEMF
KtEvcjoQl/QlIRNM9GQ9SI4tzmqN8/kdPkqjafwvYjObVYLKQDcQMyKYVq/0GbcvnSsxBfM3Cq7T
CnY0b/MlyzXqaoBFU8UN2ia6kgNMOuRJLZrDlIEKGvrUS0nKu5Hs8MnvSVVOH1Kyq/RP3NiQGDyv
SIqxLxGIUjlrvaC6FmoRLfaRjN3bI7L8jr5vTa+IGTKJTxsAoqLoXC20UFtEELUTi3zrby/U8kWG
6kq9/vcHyOvIsj9fyxE1959vFPdyHXVVOeQsktQz5S1zqJt7x1Qw/J92TGAnio0PqkG8xzvC5WzT
zGFq9yUrSUDLIDUnsDIKlMZta/vepEHsZTRcc+oh4X/brgrQ7o+DADWMIucTV18w1TDH4VRGEqVB
1rA4ZgrTtJ1NwA32STb57RfpRoiqLMkHWI+KCmcJTpoUCTmeeTvF5mN986Mr6fDafZuqu6+xiajY
N8REmhYvGaq7YidiBIPDmBMYkOTfNoP02BWC1RbkuZp9/KTCu1NKSP35wzb6dwb/i4poo0P8INV0
mjPeXN8Hz3uaB2qeKFWpRY/tuwbMyjtHBnOpcwTUXbhtQL0zG1anDPU3woZTZSNBxrNnNZ4+A9fL
e888sU5SdUK+f0xct9DnS0sDC2KZo+pj1U4jP98hlo8bxVHnXsz+AGMNGY9ZAflbcRDafvC7v+m/
GzEOy/R2eFDq4UsBLHP3NQiCHLJNsfAQMQxQhcECmmwXN/9LZpgScwtAajCVsO2wxaow3KFqucgy
rOMZKMCkED1EZc/SpTa9IQros/C0eMvnxm5P2VwoSg3kykuNPbLQdaEJ40/pPCoJZhm7Wuhcg0eM
3S7N8fx+Fvlymbs1DXqmIxHEyJHQnEnKiet6upy0exkQGntxM1VQx8qY1l9E3g/CIKdihbQkKn2g
61/YLL4tmGd34TuSvi9FGEpNrlP1gHKHEhgJKMWUidWM7dsJvAyp6+yR40HQGVzxap4OW9uBPIRR
scnYwgxI7fTR2o/7HkRfAGUpvQxkxBRb6ODBb0rEJGlxeZSj3SmS2jWVBK6vXS8aCEFxcSzVvSkS
ztstb7a01BKk2bt3dQpYyuBWV9eqffH387Eo7TKzxakGf+Qam3e30E2l5cMsmBhSI9BBJm8HcJ6E
yjbWusca92XZxkgWGrqR4rM+wuLcKUDwtKs8DoLP2EQ3vqOxrSLvostdKAHLSIU6m19VjbkHXe8f
qNBwuIQN558NYJxhqhiyFuOpHYogp8vLKh12I30CIx4dLzpm8cxvXOe255Wf7tWbelljiAB4Q4jN
roXcCP6X+ZIsycUYDqkTkf+QAYPFrK/Z9itPEhAdkh8MVDODwRjeimIjYsQ8iSC5a7+VrXGKbqeY
/+AsLsPgRzbZFhA4wVJbNJd8OjChlANoCfLBc3dgMZmRy22uT+iwJAgIKlbKM2bjHLce1X4KA9IK
qmN1J666Y7cJMHG+zH2e+2ypt3xbJULnGHG36xMyT1EVxvWRzjVvBC5yboOSuSu8iVX0eaDdOhhS
rtkXVJBCETosVJ1wTw9P0pXXOR4CFQ68ODngBV9Rop9L9Z/tL9H/UVcVrVQJZPMGj8Akzam25sPQ
6HsxDZlCmKoGJcp9c9CJnV4GhLLI1cW5baBhfu+eXohr80mQCjbV+xecvqQJbGqv29M35sQS4B73
/rq36Dyt7pFfRM/qRV3Wq0hTSkQtwYxH+9S10Qr8TO4qhBhHfePG7r5WeUI0KHTtWD2mz/q5hAfo
0XYoRoLdf8e7Y7gkOHIBmwBkTl5DJQ1ChFcMQZd5pOrlZ4mPjkoGqq31uFpwSz52uwgvsWAjR7zv
DhMGxJxRKE6B6Kv7a2gAzXLhg2BSKXkZPFddpSWc6EcfFsP91HLxyZvQV5+BC+Yh6MHezTn88HUi
01tf6xRGG6lGm8DTko7dR6EBkFps4Cr0y1+O3y9O2TdOxySLoDy9579KDz013BfG2CtbHsgddoFA
nCzGoX5bYdl8hArAyts30O8sqcNjaiy5Gvr2qzCDHttBmUTWdx2dGHRtJoc55aNlSZHTi3GzJWIA
ai1PXJeekspDA9Ai6Pa2psV4UJn3BldBM5O+TvNSut+xLmgcls8TaOXooyqxsNzCzWELnMENQluY
q9+Z1qpzH7rO4HpbvP+xmS8ucVJsITWc+1ZjpFonsYMse9V5a8H5aumzj+DaZuzBTKCocZ4wL4dS
e10LpgkBM3vaYphHi9BwCOqmAMhC/xa4CDAvxfCsSf5gXlSCViW+URsSJ0cc/XK7AEpR4LjgyAeW
EKYkcAuGXIvGegthJW6A8nSrW8reKCOWmLep49VANLQIeSbaZE40WVZJPUtLhhtiIB/ZKcKRBh29
lZZ2OQoGlWrfk3BlwV453mkOD+jAfMFYrnplf+c7Gka4EIB4yVwa7/W0UAX8JLNzJs9qugG0b3wW
+fr0uhby+ybl31ZYRbZvU504BKC/eTPjhLfRqb93w+xQ5/MFV0JOQ6BgasuYLJ9kOAZpCSQzrtLO
+3AIl59CdWvAr83NyR09XgAavFd1/U6aYtl2R5/3ur2JtlfEovUN78+UWgh9pyiUH8ZzAP3w/Xtd
NMu+Z/tixKaxUUexn0ZYYHIxd4r5iRd301KjyQ8hxLGat/zyGHAJW58JCtVasPfljYqvfyeMZU7k
3MVLx6w989cscRGbbiYwrPnkMVg7z0DI8CW6ApLOqPUumyjahdLqtcVyKi3ifKwT+BULN4fIIYr2
Bm/i3EAJNC69h0qCME9MaiqcgQB6vws0Ur0PYdqgFuSyYng8o16TB2PCvHYy4S1OhGb92BBoiDPW
sYRxXtok85qV1Fd+rpXKHGQks1c0W+KVT3XX1G3mrOnOjqQAxuf7XQPFEjGIKXySfA1L5srMzpkF
mWXj+zGzD3HMzi3YKRxY5JQfPDkABYFpZkhDufGadi9buBlpRDnjKIP0lcGOYnJm9UhJWuYXsh+X
6ppLKcWKzcDefFhzt2DNVqnpNM4VvDVLi3qw49QuH+VHpqO9aWyzcVv0cvTEEcXxXChOcyI7Pnx5
sD16LIdBTcpoJWg100nOzc82l9+00JfVmMy1b4UpTP+iB5zVJm951pVLizkHauEeAm2Ov1RL1w8g
bzDJah3etioer/jtvwq4qwPmCKKJaMDX37aLwI/6eNfRC9XWMhysu21H8Mg+H6I1OyvwkJBU6l4a
QUabDP82Li8zYCi1u1zfzRNsRImMqDqE/7/Dj69SXc7n6E56DNBo3wgeBOMOWUtMrlov5tRxF+yT
yfj0Q3HwN/Z2EiFbGREYZF9wJn5K6Tk+jr8F/fSoWysL9bOE9LfVyCRiv3xJok5XI6U8TQd+pPyX
9uhFrDnB1QFh7VgDhvV8GzCdL/TKRw9J+8JBkScuacMRcn+/X8+kDEFKSmUu1ILYUwpQobLWXIe5
5dlhDLyRPA2lOZu4rQdAK4kyoC7XkZBqoaDWhaWyF+m8KMoGMqDuuVup6UfMkhIzTxIF+vA5KVnN
U9+wQSmJQ4IANMyHzdeg6JNijaDqku3RqGiQO8Xv0JCAW5+drYW2klQr5tnN/nhMh0uKRyseH2wr
zzzqLFj9dESduGcO4ewmm696ze76p4YV5uMCwrTImn5S4Yeau6HRZjFihn/smNmWBWlMef+xbg9R
zdz7tB0vAZkKkKcXOXlMcwwQEpDuvk5INe+CluJAJTI+8XPmfMSXMq1D29IMRFYNkUIYViro6Yso
VjwAEvC+gF7niK/2vQ9Mr1cpagRPvYNGPj4yUYT8q1jbqO/ZmbbTTyKxE1R0os98/cy1GURhF5gW
anUsjSfr6J/Bl39MG8D0+wj5ZF2uXdT6noSyY8cvI0zSZR69wB6ajx0n99Rjr1L7oyBaAqBDHHjh
ckHqa4nEq1rW/PIEBVEQrQnKpRo+PqHWAW1IWcBSNvAUtvXgTJd1wpKPSUamtep+jakPd1J0u6sm
G4bD9k9yRLCBvpM/8sko2Aa1thx8++VyQf07ow2tybo3QrKNiqCfTkadC+Kl1JLmZ+hsggFnzfz/
t+nM+7YNedtg9PdF+W8sFAeR5sfBtyWqRaspNnEH0CTVhmE3OdUq/2GH4laMyD8KjeSc5+abOMVY
NNt9xCBgXcbB51TeczpW40bjalGEqVUJrhTRqE0WIAqgNjdZCAkBFyAekhRY0JR+uFr/2LxcrXiy
bQEcRSOt1qrerxPdaUdOySecpT02BYG0MlpAgQQT71ejuBgxD3gQBgZOv5Onv+CigoZnTRJYGg45
P7dXkqUT5t1vp4WzVYI9MHV/CXZFc2zpKSmL+BG3/pK+qZ9QEAc8Uu+m91hq2Xpmsyt+X+Qai42q
TwKfjaxZ6B0NFse/ufR7uQKLK8EI7WRdCBjq5nm7KBvlf3e3gjz8xc7cFxGyp9QsYmwbuplt24hA
mwgt9+sRe8XXAJKiaFNRqsc9XMpfEge0TbC3QkRYOtFj1MM9ocDfOIsfNXKzE6eHsRyO/2htdejR
LhjaTQUsB2K4HrfjTk7cyL3xm0thFXIDZb3C9POodA79aYPh9b7Pj7nR7N7y2bqXo98tes/Xay+X
3u+wefypJdiLdnFa1XoHNHrezIVVQ3UqJzf4/gBTyeanPTDDEDROQ0bmiciuR7D0VZuXhisJ5/OB
GESSnVJLaqzpuwMe6epslpFDYQY0l1S4tnMOxftgPDv1RvBqYmOejo2F/5SaAQcHn5B/UY/wn1XU
ws22Lj4SMGH4jz94/ybXzDOpJttcrA9fKdmXa589lyq+fkBWJRx9ZNKwnfBqxi0rAP4dkY66Go3Q
9ChmiSFtu6x8gx4ND3lP2mk60bTJ0Rcju788EWFyNpK/Z2oRzZkJ8/g32Re4ZjSG19LAFXPFu4IS
SyNmCdSOt5P+okL0I/bUpI8u9nXHB1arIsSmSNG5lRS3l3FABNwVngKT5Hl2r1Y7vln58jI5IxF6
uM5shbg1sTQRNVSva/pOjuVC2bYvPYqNZXemTa041AyOeMnAto7X74GFjOfFA+pBwX/IzIHaLZ0d
8WjshXtK6M1d3cYj1Ow/mBEVHHKBpyleQ8zAHONdlTLMYxNM/HI6gCcK7YjcdfGhR9oUX4JIxGI4
xPyVPgqlJfmQIP+La7TTcG9+muEeSL7MR9EIOQgxSGeylOZA6b6VZfMWn3h5EBDrnP2vqfrJq1X+
VlbitILQQ9kP2JNjwLsPpsO+/JW5KdF0Ukv9TRsKVe/qxKCmzYY8oHlQ2bN7rwMSMgL+FkHGhP5G
Kt1hRsMkGeu/Eh5JOXTDYp3HhMbnqpCNiQSY8DDr/KdEm5FIDybDAoN0ceQjiYRK6/F40cigwaPy
0GtsPqvUafgqgDbRuJ7l6z8WlQ+ZTSmIAI7my1nnEgzhfgCyGf8gf7Bt948z16mvpIaXrYUL/Q8k
2ngud78IVVknVAhVpj+bXE8qhqyfKLHLF0vrq9AxWCDKCI0dxTezVIB12Gyg7Wmrw4pyPC+OhgAH
xzGLZ/Z7FsXMTPSVnTKN4y0ONFkhW6Bk/r12kUw5Tbm2RZV9Ag7WTOYFCyCw90UVpilJ5vIEnDGq
A3owN/viG71jjTcfYiSe5Bfg7BnJEjCjv93iSh0VmX8OdYcpFwIF5w+ho9NhPliCz9jbvFKauvyo
PhfhQP9eylbNo/YOjm+9/Lhec4wMad3oi/E6YfXzj70GbYs/BFCGSum5Qt0N3PsSpjge9t/I92Ba
SVML9fkNCTLhUjCR0NTEY9spDPJmehtLOOouzN1FNSG3YoQSfG2vFwtzGKcXAz1Ng4bTVJbnbHed
MKaYef//H1QCwa5ok1i+zHZQR9iOSgO5F+moRxwdjJKeL2gqopSRtN3I8zZSzjLKRuUoSgV6fcJe
1F2MoPwq3+hnyiwB+3HDv3BFat+0hnHovz8Bw7ulCQjfZtD20gGrbyUBmxdeZ967LzslQ5pMtdeq
TEn05djiXniBNB4x3lUgQjkdAgaksjkXE0fXiuctch3wEvOwNGRiInkW4x/nm5bJT8EgHVNgkuKL
9yrVEXJsrViNklUf8iSTGJSyv7MmEKb5rB1V0tFLNga2tZuvA9FeRgY4iGn0MpwMJZ6BLBbgBexD
oN74brztTFmH4IjJhTcbzWFxykyM0SE/85i0FI8gwmtj+Tz2AfUkbebsT5hOa900HIr7zpQu+Exv
U3frnAX8jbAQaa64GNj3yhUT5zbTyDipMDpSbuVf1CULiAqAKwGiFB+Di8ds3hCM7JIjr9z9TOgg
o3FDLlrV1z9CHpbcilpT8A0Qae3aj1fLLUze5f15WZgpJf5VkOvLb77UQdcw9H5cVaOyXeTachDy
ooT7uMvFMBjua3jvDfmKZuqcvEdMKF6ursW2Bfef4UAD51COExDh5GGC/QbaC94p3eHodM2v1J1k
UORZM1487KZkBAYruBRJieKmw+eOgOZHY7oDErnOvSNPtwIwTL7YEINST9pSQl2h4zV/pBlGVeI2
P1BFW2B/Ba4VnEsHTws+ofCHtSnHOriSsELhzTiFFt6LZGwe2TTUmByUqemKqCtm2KJ1QfRfOxRb
TksVgqx9r80IVNILHk7Dp+FlpVeiUr/fvAAoM1iZWU7WiqKhJ73xlAZN0wmoN+RT7TME+0mT76Wp
balo0t1/77HbET9X/wmDepJtG22Te65aZpFHiWgFhFvLhzqLfNN8jH2ILdgPAZew2oYX4h6N9ozg
1jl/SzOU0BVrS3NBx+B2TUaf5hbfXf3xnzAGotqBEmQVynGVadvn28NDLxrwp2HPhCUXDODvwlsy
hbTzQpTLLN5CAXQk0RHWbbFTI2IkvJwMGeCIIhRhyVTSWNeTtlfVrqJ+l4aP2woVkOAqX5AL2L5y
zD9uqXYAfPKuYhCtF7luDRGeeCu0x27vcqXtgqyrisIBP6iHtPwsNzPhWAWsbagyaaX5MpPATk1h
Qn1/jeSFn7Kkfx79rOEaKfI8tg6s85s1+XUBAOj50KD40Y6Aeo4DBkXKaxiE97lQX2SX9cVUDBCg
fm716rU6w20sxp8ZgOODSlzFbCaklwXfPMZMPoU2bq4I23kC5P5YlGg3wncEgwBLdZOVMOJj5Gkh
/eyOmZcg2teI/OXwQ7MQfCnffCu1SoJzIQNJNXPfo9sPchahcu56qTZCyhu9h9vuLGeW2oYF2gA4
2BPSnfH7igP2xeD88o86mUo+4UFnrsJrpYIFcJee0iMXapIhmPYe/QWbyXKTvzZbBH6o2xt/Wv9u
WUnjnvsjwsxAYASd5Knsj8HP19niUcYCxcKMMRLVrH25sONFtsyFrp/NsWMD7pogZo4dFphVt77i
7LpNv8MQxFrf8XKxxrbpxKPzq67rnXqHHD8MeqQVZbDTJj+1rJ8QCHlfH+Mb0R20X/qDl4YEvTDP
/0vQnbep8q02lGlA9qmyRtnOy8UvbG+pRouGhpxPW5TQOZOhg6T+hv8YVgRHkV8U76jLYSaoejpi
YsDKbXbM7Y6RtWvKyTS6kVzkaDKuGBUgbFoMPvqG1VhBbhDPZikyfxx4gh7KTwGmii+A95ITDfEK
EuI+fRkwZpkcVQYT81mtSUj0BUmuUu8pXnPRrWNlZ1FSVqEqQ5P3ScJyjwE6etaYYQunqHppNxEh
N15fT716J97SW0V97oyg5nEia5mfxfmKStgl+c1CLdCRHo6Ny8nuzTnofw0s5azzGzLRSHgRQ5Xh
Mwz+4uhTsJFZNxYroOBnLJfBekdwxMG+kfuBMqfoAZEk6tNSMnB5qvi1pg4GWUTxuKS/Ipdj/bcu
CkCZzgx14UeY+zpREGQ+Uohp9NTjALTvQloZMDT1XiQ8vzLE4ZFhh31gzmCa4WqeejP5O4/qPybn
JqcbS6LRjBnpXCizLC0LtrMK+vxqROh2lBcnE14/0YyH2ZomazOSh87A8iMnpr+ZydFwVYRL8sIu
kl6d9LcpDKZBW/mrTDKoLIdh7V252BiifS8asaq4z6EaEjk6rutYhMxlarXDkKTZzHM6gFO//ZC1
VwjMvkmGul1UhP4JJTJlw/4w7NT60TOR9TilBq0Rs0YkxnM+61D5yncgRBXBszsCxXQcwh1E/G2w
uML88mLRg6AHS8tvAU6cegKkpxfSeBJJkRr5qd6Vg3TGr3JxyZTFPhgaeUSqRWBCLbtlOQbKhSJN
V5OXOkQSXnMFKzq4CDT2BNPGN2LsOm+HtuVed/Gl8LjALtsogK/iLsJexMk+7yepHzy4Gi6U6+jB
nTI+96ZiJCUxcqE4YjGLd7/Go/sYDSlusVkWubWD9avHtRDyeH+fg+UETzTENM6ZLsljVjae71yC
DNUPAmdAevypZ9/leoKpQFoCHcoguu5rqLoRcB6W9S77FdDawjjTcMNVFHKO0y9wBzmeY/y+o6za
5YiIW4Bxgop2PrqYi/kwSMStaY23oavwSGgjKVCixqmf6xx4GpjQb7I+Nw3t8liFj3aVa232u6oy
18rUVgOBT4cSuIVUn29ZQ5fEwgjcktT/MJeBR8AbEbZLcIU+IjzFTp6YDlr87ArTmTtCgB+r5SYE
x+8XKrdHW8sjnKnHJi0HCOIEGrmICosje53hF8x//S/rm9sRrjCUTNLEx+Jy3ue7ngu3/ej88xD7
p42PvpKzacA8jVju/+JAwqVG1JrK/djpRYJGjbc5gZK3p0KTITTshiEHt8Oq/AdCgXpgZZRkH1AZ
tDgwYo52u4Y/moRNFWTRC2/hl3cM9JM6adSPLFyNgOE+FYEHOIIN2UAfuVA+VrLbGdmSh2CrBpvR
CMZ6Zji43wBubxwJTzuo4NeO+PNTdg+3NvOvJkkjiHjIjEMEergopzcQ8cfgreLlzmI9ybwsyl/1
yuFLRcnMKmXGEPq7urNV/UBEW53NF2j/cHi9Kq3Bw/Z0/PmIjrNZwqMO4ZZdgTH7DebfhmSAVyYy
n0+azA+uGjjS558edDoT5lqrHxTHP0tY7IhCxrtyn5q2tnS16oqFaRjTKycmDildasrb95m5yKkZ
5tYBPYbo3XCGXrV7C2OVRW3HE7fMiIGaloiyHYB1JoYZ+1wxe23IjBTRrDI4jeRjcfV2tD4jad17
RP1InTATIC5qx6QRv/eM5pDobw4yrD4wLEyg77VrL9L9+djDzBV73qA9gN+e5Eni21TAqWmNuzME
+MQw3g3x8wljF5dXbqV7lOpe8c0AI4Lf4n2ucvjztcTiF3LxvajFgEl3E0bu2AdGzGKa9MoK9jBn
qEmq3/z2ArmCE9BnuMOvc9Jhlo1x3anrTEt/Wi8utjIPwmmwd284dkMrQV+5gaULygQFcR9Szr78
I4n/cFbXuXGv9rGbgvHr1mt6iN7QD1sqc5UJu0n7zLqOy9tot/BSvvWdnCX/w4VZ1FB8xwVufjSz
CrRGVsNfc7Hkvt3Q6oNbcc3YwYVCR9XMFSzhsdyWP47m62A8W+48W4ewIngXA7yGSukxg4zHPBOG
2A5wjIxvlR3ZP9GQ8C4EiCbih4cVZIt4kdueAha2B6/Ee7kDR8kKSsOAAsE5yD30cj4zehc1JDSH
V7pLwD1FDY/2cTF/Nc2/b1v8aNxdKDVl93qvaXpb32karfrw11B1WzqCUFSpxVbfNFrwRLPZ8FXt
xl/NHGcDPvY6YaDoP4Y5lHj7zbzmXJgT1yKlnVRqX5Kk+VuM0cB+RgTnotP6X3m7l9YqG7X7opGu
Jovc1ph8to2vPx7uqMePlbM19l4mtsbRmohoQZ75jVgl2rGspyBqC8w7gCf8q5WSLdhmLh2lO8MH
lRhZs9Y7xsQmmRVPVUB3qX3nkBHLuXdSyr+0Nd61gTPF8e5pxIni4tFvMsSU/2jN5ExNUe7NaeUt
WiwDg6/Bn39sy55XOM9y2BOO32zMdYiBJtY89UWGAxQrOvkIg7Yr4DOi6wXSdHaLwtHLhda3Cs57
Sj9VACqUDdSDwt4VQl8dqYd/WBHKGlMPaGudQ3UUdO4VqlcgQND4Pea+sZkv5JrQU64W6NapWiIY
nWiDFzopNkCeYeP54oIDPWN4z7t1A+qF8BARqfOOud14V1fRlWIrrK4KGkFJKeB59DIeGQ8KtVp3
FhkL6FTK385py2uUth1UgkTy3fwfRc9/3/o6vpPH/Pj9SdI8MMtU5KwKxanUR7FHX0fafIYgiSLj
vK6Teyrc+jxz7zHRRs6/CRlEf2NBC/22VA/TMOrCrkl51b1KbwLm76p7aC4e+azZjsVcirmjMlKl
ycQ10l42+Q3yzb5pT8NoMZgJll6U3S4fmMjfZ5MiDLPq9fBBOvGhbHUueT4ot3aVnj6ypjjX1rOH
gjigvy+If1YjbMT4OlkQaQ94s6YoMPfl5Dahisiscedr9VIcHEcGTiP5sN+7cc/0bKtwwcG9y3w2
ojD+737xSPrsc0hU+qD2gawYT/uEnaMawlUXRNQOTXiLsWGuDv9NnUWUrUp7et0SkkywP0EOLnmM
ZSC2pYKj1KCtQEgUiloUzQoXZgsMiEmZ2YWGy/tn+IVk0AlJwgL0sc6274B5IK3pjsBkHTDi5oDB
tjyVzPaGnywncZQU9wsvqnKhy8yuYodnwwRDpcYM7VfZaz2JJbtWG/CID+pytiUVLSLANEsxHwxM
KwGYGM9RYHpEJrP5aTE1h4LUy6AeCsUvdd2zaUyaxEAGP4tttTVNM/+GJ2OC4C2mg+Nr986RfL6W
5f2V8NwdhsVFqgcFuZ+g/yiaDIOFjYWdizTfUI/JNUYCL7gBso8LIlirZYDUEfws7su3TdjhwBNd
BPVrEgD87gwLA5NFjux+9VsWCg8EJnbUB2mayngpMdtk0ZwxY4XOSl7oOjKQYfcgrH0eFN1K6kbd
PRi7TTHZFjI+FaVU8mt737h6ZSx5z3Jdhfcwz0FUSHxTRimlzU3lXqr9DviRB8KSy8PqJRfXRjuK
JeTS++6UyM94/V7WtQNp6BBxY6wZ8ielXvA3h3JQZq8pQeuk0dMNAhOSsLrV7yzlBneA+TYDgWRH
M5n3jrV+7OmQcTbxf20Nou2rU1uGzX93kv9A9VEosXPLG7dcphzP7LkgBfi6x4vNiyCCDwERtPuS
DH7W4m0VIfUVLEH1tX1wBV0l5NvXg0Y0I7gxJHrTi/27Wr7A+w5ia+AzGYf9+AGe962PiPPUxQZN
aXa+PhwncR1jCa1LW6QdNIincUgFzjZQnwCuajsc6KSTeuKOmCLU+qBlBoS6lYtaY/fwCo53fseX
gPv0Qq/eBg7698AxVZx/zoPuFOtgvlIAITACGRkuzpkwJz5CD4Zd9f4isynXS0epbWnW6s4qtvnY
/Gf/eKCIrRkVfErWZ8esWx78Mr+MIUzsdvMdJPT1q7CwIrBrd5IbE9G5fBp8ypBISzIIr85PqGsS
w7zoxd11272QqyqLA5Pwn6V/W5ZcET3WSh9gI7DWZb/ijvOJL6aka6HIlZXDdnwst6maSot6PqEO
00WCoo+IOd0XzJmo0syVmBfAEOsYSaooUXBWavrnvxGjZedU57XWYTWyO8rvRM0BYRlPci0kXp42
cQtZmaiGDcorvoyvlIZsHG91Qirtr/2xsd5AbuW24deY6I2KsL3a7daD8CLi2id5qpMnNcE5I1Y7
O9wi3CKvG5uHlBtgjLfFJwPbVj4zBX/P/Lf3BTWzFirAzGa4q11oPka1sqFa2s1gnURDHeGZFVN7
mSPUJIKTDf9Vh2K86n8NJo249ZR0XUEltkL57xDUUAMi8QsduuJUbzqhSHlOHtteIbonx/8tY1Gn
+k1o8fCfEsg0VTAT6mvNkBE3yXnFg/Ktng7+wlUJjgx4rA4pv5uVvS4jwOgTP1pPNvaRvCyugXDA
An1SDkMNL+za8undu61HaoxFRTAg0W2pUrnpQ4aC4WR/y8slpAijgnzcxZHbJLW8/goeyGAuNn/N
k4V22tCqMcIistoUqzq2JmOiKUNcHcqmvmB7WdtaoeuLRb6+c9+vGSwjrrposQtq+2UPZ1T5wlZr
Seq3A3cWHzvD2DbVSsVqBAfdZBsqc0GfTLELb7xAuprpvz+JWIhMG9M4qdQTGwN+0lRk91XrHWvV
AuNQVO0Ton+RHyjgM7Wyl2NTozG0k5laDDtUlVWQ3Vo0YFWnIvxqmcSl7vpFpzFeKq9acPzFCYl3
mQuHnNJAREh1sYni/iYfxUL0gD/s1aMUej7j+eXzCG9QhPHmRxILGJeINn5nGcwcBdsWAieE6iI/
URJbLin1/YpWI7tZO734XG3KDvQ/0bRX8bGoyC34N8q5QUhEUQk0eTnM+cQfNa6I5amjkqmCJtay
eiopI+Cp4zpwPP7cEonq9i/U26YckanUY7AoAGEnpyDyS4tXbJZian8KyMEJPgx3jEK46CG/9tbY
Z5PAFw8+kXI2NKoZnHF2TwGORRpU7dibFYiya6Rbc8gc7iY3z+VAr6DNxQIinLCRFr7GW+jOZZV+
Da7wXz7xsHoefTM/O6Z+YvLIPStIN3IfDiL8Qz6gTakR9Vw2bpPhk9ZLwqnVzOssGksKh3NU+YRQ
8+zU568HfcqMRN5FQjDglgxCYBSooA2UGGm2jF/P9w9m0Cq0k8y3WflWj01CM8SFkF/QUcwVeM5n
lZLXhrqrU6Sclrnq1Egi9pmLic6htO+s3TyF+QfKR7myyTDve2FL41QAYIZhv4OPA5xLZJjPnDbY
+Bmzgyp1g5SImwDwgppMJR7fRF7XaUN8s8y3HBtrSpM6lQzhQqBJQJw7B3J3pHPTzLZEE4Mb6UAw
LmGuVyBJvwGkt3FxTcjI8gjyAqNavO/rGqYw7oA1R4sZaFRKNG9M1kIsulxIoyZ6kvRFtQ0eq0Am
5235Bdhu3C071O/XURPZDCAz8ZkHJzFm1f9kgBJSeYBf3McHJUdbu5BKcy4u6VS0MKNnpTuxB/I1
uQJ7gJnrgYlFFL5AS+EU0XEPWCc0cV+cqVZlx9uHry74qFRrAIV+cl7bUse1we5fWmqxkvcb5QiZ
0RD6c8aOd3FCbdlDNWg2QeZAL3K/XcUSavC+I7r2WW/6gsNuEBtwZ9Z6SN35hdh2MmqCTSAhwLhH
epoFwqjULmRgs7zHi7qBdqmyti6CxBO0NAqsRw2zYs4OzQNGQtbd1NwWdoY8GTAP+fDeNt5PJtKn
489g3hyviCtu2E0GGnXTuy85PVbSLADHHD0Q/iSiYTtjqksEe5TIM13oI9UW542jpfoJcwZ4r+K3
WlyXT2H7X2eCFK1EAU+kbUKXax6rrmgppUTvktiLr8yRV+dEgppv6zPpF+QdWAMAxyl/t1WdcpIh
zmvE/MDp5oYw48RfFGT6sD1slEGRWLkqj1R4zv4PQluBjqUcz+6lW9Mn8AcMITXqyuS4EKBsoKAo
YpQP9LkNlwrMFHe6tappgzJFKcKGCOY/SzpIs4YGzMKrUMVPGsU5PeJpNrWe4WuMJqy/NtWZvXaO
VDUQ0GjhDLTuAEwRKz+8v5GUXpo3AFPs6lgYue3D5boCHB91W1TGCZp+R1KQuvBOmBaRlFlKXsUQ
+4bvu5bMAeUWw4Gk88f5Yhul5FLaRb0sweAmh4UC3LghMYCZ8pvTY1+tZ+PoUyeDa5jk0QA4Bsgm
/8TQVLyg5OeimMu1/DhFTWxkhPTwUVG7Ntk7yEPXj1AUauwHmp+RAyAfbE6QKMUtQvwICBB5pB7j
3jamfV7Af5YOEjfGqwELsE1rJLoZstqzMWpXwtm4c0PukyqsRsfDOS6nB0f4HbLQOhAcr4+gXarW
O2nUxyCV2ooDGTVzerB189uuogu10fCtXVkj6hxCgx5HOAY3uFvHv4FOgCUYLUKOy3bN7E6C7gP+
wjWk/SmQyAU1iJA+yCG5BJZ5jKDJ2D8EQEb8R8UH8dAzKP6SSAzEuiFOxKIjqfEoyuK/nSHhkaqf
lipYYtEtSmSi8nGpn+A/Y9H0QyKUvNcdWnql2eWBLSo2VeRdsF1hqNhEvK2M6QJHS0W/l2Vj43zw
LEagKlwGHR8gM5NkVaaJvJSfenNAK5/MvJ41wLjJddzEbfnVTNleakilM2UM/cyjxcQot5kniuQe
Z243+bPU6OYvj8KPUm2mRQbNae+wRzsv4Cre6hiPTE8MtskyipXaa3Li9e2QegCsGEqhWbpXaVzi
cu51jLfyO/x3BnV6ADOOcW5TqI5kfTU+mo4rmYP8G0OciQV9B3UBAuEaXJp65FUONVOXePbBki4g
wzG1yTaG3o3Uys8XNLlQKutzWWBYbW6B1mmw/yb85n77DFu4pKLP62GrGe1ZvVfDuQUAMTGlTnXA
jTaxH2zRQ4s1Ux4OB//G5e60Z7mcrW7ZslM2HEKoc106GG80ob1YrJEf1L28WItzWUubQq1ScV96
x8qJRGrYfPs0+TUqa6p69LD1X5nDumziJU2Lo13ZqECd0UsK0Fn4VDdg7h30TbmufdwsgsJxKh5t
H07C96iKBuHx0Zh7nc7Qimdi0475ZQlrFWQUWYYIbBXGrQq1Nr2Y+huNhv0Pp8+jEfvfo4jMlP28
noK13/hFTJtTUSrwXlMPFTrTxd54UU2ssR7AetPoCkUmwkdfl+eE9ji1a71jupkKJi7Aod8QCWLf
1VuVID5HfU2FgMCOwG57kCRto7k9kSN87Ax4yQ+Vym6SLyXZ0Q1KCtGbvmET7L8uzhUcHTsYxRfA
RSbcTKGGp37YIGzpUeBsWgi0seEvFZ9qNS48pruNrk2t87vG5yiKqqYE0cvw/bZMXOrMN7rneHod
Wn4xLv4vGXsBNY+16Zfep4KC+If61TgNDtilEYD0uJZ7bHvv0JcA7Zwuyzzk+/13kTnqN3owutb0
4B8C/AyKPob1cz/d2ug/ox5/AjP+JE8ipb4gAo2bzNTiKa6kezIfoRvHQADtThktbi6gq0b0rxQF
Mcl5zwfG5LgyKwecRSOs/DeWFhJ15f2kOWgEPBKZ+MHpU+I/Phpi3ceHDAz8nBnYjTg9MTfuAfdq
Cs/zCKYmOv8j3xlMaQ++YSz+EaJyHS4kAQW1/9GgIULwZc09p/AVwtUYKouJV3kHp74DIk/3WIrj
028L3Ag96+7MTqw939iB9zBLzzkyFRyi6MuTmVmhyvdBRlSxQiw6q2pocGzDwNn7AsoN53C46w2h
Vsz+QrpJMAJFfPy6p1rwf4uq8Frz2kO/6gPiVFth9cwGXW1A+hPftgGCrnreFBkHPPeBOtE4CdqU
ag92dMXibjOyXYwYSZoFwb2PNs++RosVkvvfUl6690f83MGQb9JffZhrAEGK1n9mSaus9M3c8Tz0
WWU3piJbnZcaJ8JEuCX5AZCbqAyM4oo2FrjAH/NfOu0zwJ6pZzHyIuGctAd+8qFkuofC4fgV5u61
K/pX90ldE2mtBGaJxewxivcvbd9RJEsPptB/Q3pgl9zOPI3AR4ErJmigbk0mWMgfFFLBW3zVXGH8
hq46iZyCur+GT6V3JwWM/IOKFAsP1/+s4CvhEQDFbRvmfZqEbUqJoIoYG24vHhXl//zH8uzf7l1h
GZpwShvBh3UQ8xHh+IvDv024jemQysrLTyxCPqR+u52mpzA67wAzedebR+OwM5Rogp7xCBm5cLxX
uyyF20/znMQap5uzXiY4kxx/zSIkTbDKPcz/0MwFEkKcBX9o2YUYrTjOu2zJ8FQpdWSWqoK2R+8V
QvSfk6JZxE4caVvMg+7qKdY78TIgMnnsWNOO/+Zzb6h/+Sw2sD4XjtqeVrTKaEryjAt1EtwSUPed
YgtvMAs1WFxFnyhRhFBkmP8PBvyIusOeGtcooxEgcKYmjJKoRnG2QsHUS2m75dKndrojFDa6+OfY
99GPgUP120hwOOJcIMhwxcwejLCGikF5/EFKN5xFfa9esPXvZar5A/awB2d6HKJdmzuJMkqkLoYa
IJWniaz20YfeP0EURVfvKAHJJh+EKgJJN59qpAwpILJimnWq4qMRklUnrh3RAKFl3y/pXhnutL+C
Z15OM4hXWVFab/tCRyvQfWuYelAHA7Ci43D0uR2R1Hm6cGH8vCfFrdvRGG1/4L7ilfJ0wU87mNk0
979ppVGkqkAmadzw3eATGdMIHIwvO4RwWWSN0kAMUO4S6QHDiVAxOJQH1B+TThL3l0nv/7WNOwQm
iQTE3hMWjB/KNT1betavhdRG2w1ifl+NC/LPlJhOQ0UrjHxwvVQITkM85lo99fBEfZ9LLFY5geN5
dhbbkU9tRL23LFXqoOENWBmYHPOYUiILL1uHyFsTdPoeetaAebYHwM+xRPuEG9s/cNW+AVvKr9oO
9FQeCpsSIAJpmxN6FXR1KcV6ORX83thLArO/Bq6NM3feymQypvv0q+dNbajzCVgPnFU6SEKxZ9mk
do5L/shULCnr1r6WNbf21ZJSBmIn/0TnVLhm3lvdOVc6RMI9tBh76xTOEWwLc2+U2kyitUmS1d8d
g3T/gzGN8u7ZIxcn1PGr93l09XASHVT/4hLjCKGHDZ+T1qu9HIYW6ygpWdN76GitBEVElv3g9Q5h
ER4eQoEzXN4OnjlUkhEp1y+Qgkyk83bskkKLfmMmM2Bqo9MHL1ws4F41Dy386QDpR9V3ypC329Bz
z1tEY7kDQy/oJeTpePHMAVx/xe76KE5lQYAEzzEkxWNN6nytu1x8ST6CJrdLLiJ2fw5trV69CYSM
29xrSDKN9sTJrtieUaM0oyUOInYC2dIMNCGgSsq1IY+0+4mEdNRd6W18NsoOJZp/G6u0obGNFkoU
iXEjgBL1HRaapLtY+4VhmPUq+0lpx72/evH33Z64wjtrmqEMxlhPvcCWaE8wZRZC95exK+0d7f8e
LhlhzCLHAUFTGqIuEnFbq1aC+/WG/2COv0AzAHU0Sd1RxNQBe+iEIk2oTmKNdxb0LnXBJ1sdHtnl
aLOfGc95DpHKLCutxfM6zeHCqEU1g+e3/rcHAXaT8NM32nuavsbp6SiIPIlWleAuAxdYjg0bfB4e
1y2QyM3ZeNv2rUMnOofMLrloQxl5eIZnzOXWmW6Jc+ez1jZkUs2Q7x+rq8YrdoC6nCupUuT+EjUk
BM3/QoIdr9b7gu8nGKPdRRf2BYHgIwwlriymPyV37u82XNX7CLsNFoEwx802jPLrTzaqddXTemcG
5uJfzpee/qEWMzzIZDU2U5XQ5qJom6lo0dDXk5GnhyPmrPGy+IP02Cc6Q4BLgXVG4lRi46Jn8vjU
SFR/7c/UWSuXDjwmJm3eZuybrkWfB/e1ilOMKY5Ybj4I8IocSujfukH29RAXZRRQYvGC6Hwbs/pE
QLTr+53mmD9G7Pq3vAUzngf9gjheJHsCtjZh4qBu0r1/FGCPdUZRZ9RySZIQYHCfGPOTTywATYm6
lcwP5/xGaoeBsgWo2wECdDu/MnmazxMwy4299+w9kiFRH54ib894G7AR4LWuPdvegrCdNSXE4kXq
x68XIhLrfbZ/TQVDKCY+Jx/wQ3CKczDxe5aqcL01Ycr3vN0U4nQHlSmzSBpvIFBWHAIpMYKXXxp8
GcKHluG2QVpH5kX0USda0RL+2tRrDQ+AoAEUdewrhhXFnAIYPd+4H02KKj96lb6BgnBxOXTaoMJ3
JnIY5v0nVtMI8vA6AamE2HN8bcHIbI0oxteQcKPgeRRf7EamIsG1ChcOuwwcz2+nQtz64wzaJHex
y2T3EHo2D8x/HKruEkBBr+MCiHyIJcU4o7bOGVF+PN3lE7+Ru4Zwc+GsIBPCobZQYIMKMRKspBpH
12dlVjDRYVqvhpNsx/x3usMDrnk0KgeQEFmhle4q9mHSZ4VUbsSWAqzl4nkfFLKCg/B704d+WZuf
DtcRa5jTpANQiiRh1FhIfIsWicjwsIw2YOIrxFnM11bKfCmyCMeG0k80tI+Qee4yiNAhApbiFwbd
v2otlNj9jYjAelXQZxdd+h8KNau09id1zacPR7CI43zAzBKdAbbJDZ+f1vUYMGslYjHuaj8fVtb3
noU81wB/+yEwZj2WMqjB1tvs1Le4tA5O6z7u1RHmHP3TJnoIYAsQ9YPn2JVLYYS/E489bzvdx6J6
V57Mrc+brVbRQC23PvYSqk3Tt1XaISTag3yrB15/nGfIztnrVyUu6MGySsSlGAx5re93NwJjIs42
f3Xbf6cYqbgq41WrQ8+8XX6cnOEc107Q0nxG6LFHCk6Kw+RwA5DdjLfc9yS8JknU33h/3nLtNuFK
FEGnUnWFBFWAaItfcCvfK0kw40Te5tXLNrLJ29dTnQSBelSUrskoUudE2ZhKI7aY+giXguu7Q+sr
4Z2F4IVFv3l0Wx2BgIOVTKEB49rGRDCN8D7g/xVUc9E7TeTGKmUv4b3zK1tpDOz3J4p41HAZVOUI
eQ/9o7G9I5Ie25nwwdyiwd9nsi+S/W49kVLnz1XJdCxp/jEYl97NZwgGoWTVl4du9GqIaK5292ly
ayj8d9O0AN3A5i7/F5rg4nHw6PekzeyPjxohmaQroUsp/ICHNOeFgc06pHmKbEnYDEqjQeDhA4pe
1dMRB0Z870kqV99Kn8jj0UV0+dhkJk9AK/Q129RdYT9S9Fk03CB4yRDAxZ2+gFf3lBkjTp5mUTMT
90LX1+J3RcR7AHV0sCdPc0foPhJXXgZYonbIaYcOWd0w2J6PgUp1htzE2R2kNxlXlOKEhx/xx/Vz
2JjSggm8GlqHTlotGXZnZqRbDfo0tTikwYF4p1XQM+VDW2NrrSSXiqdJM4UeTH/2UMpKkGwsmFLF
5ymmvbzytHQ9wPuARn5/7FHDxjV+Or/SliQSDKMMbeMmEVqI7QV/tz34zmb+aIy8Un8oylIAl2Sn
H/5TbJOIGlRBpR9QxapveI2PRVUHDRQvYOYnYfntK9P24sy5T2DIqPSD+TKbz+EVP21c7iXbBAyB
PUSwKIpHPf1au2hc+DIs1WOsCbZhZj82DJ4T87+uzTBi6gduQz3eQ5YGCWI/Ooy4z37G2NmnAYAL
+IpfBVN+DDA9Yge6k6cefa+BKI3F1N2kJUBysuxORYlXbrdgsL5JJiOP1/4CIFGtMcxUjGTEQU6p
aRRcEvPXbY5TfNbn9VC28VbS1c625bUxDStze+uK55aYfkvrgbTo8JD3/gAHAKXiXFB/ap6+ph3y
5wrmnWqT9NEyBQoKVbOIcMWrvOwJPxpyfo9FDmetLeeiIDvDEYn7Yamv41u0NeaYkAz+ZiVCTcZe
iDigf2g8XeafjwffVDniWwcFhn4N1i3XbhvxqS6mBXaZgkPgaMYrX772Grc54Ifbbzdq2ijqMnIq
2uZbNqywibaQTJShnkTbC7QGlRDUT4kWX0h64mfS/kKAjnnSmP/ptUVN10fjlb3M64GBgKjID/8s
drTD2oZZtbwojju1Fc9PpH6+nt4+XqEvgTW/BnonWgByKa4o2vm14IZAJtUXLaQHymktbK/fbwg9
/0EOPWt3NkiKSwpufPsCSb1j2qNkfnUuez5pLzL5WPv6Xhb+me4YfBEJqAApnG79z4K4rKrTHAWb
sYAFJfg3tE1XeuswvZTVsUBPWB6jqTRBFOulvAfKxPl1BODd84opOFpkHo4uqD4OfzJcVdbplqSS
WcPLYdeB5julCT0Y6oxJ+Oc6FV7GxS53gvAbGpgg6gVf+gVWZW9A+xK2Y81v36axGK30q2iv4QdD
XlppHQmCvMR0yYIjiNS24pfVNHH0/ma8b7u62gC7KNFKDhbmbPoiMou9nP6/DMa3+6AiJVQwn/sc
oGsD9OETd7DfEQPWm1MePAWEsEXs643mJUB3DFhLP3REBcIQoI4Zc/kZp3Zz07+jmTD2V5B0iBy6
TCTMcJxwyXquxDR9qlMg0V/eFJIaB5LT1zV5Bs2DWkztdP63kFdy68CpUrxP2sh3/QcgjkGwZV+t
QqOrRgXugIB1pRSnL98FEOxh5R8SeZ0JSTidj8LIrOSsdpxfe2Rv0K12VAwgrSJ3YQfaPE52lt4K
A3blEMV5ZWiLFnBHMYFTMuaa2MwRj1FPoMelzS4Hnfq3KUcuFM598sB0MABj6bifh76u+t9yZlqm
VYUeGDdKAF7I2AVqnTptuh8fvGACv22TbWHXJwg+xDC2hea6GM0idUslN/M/vztq1xRAdYycQDEY
fsmYUm+bwdPhm0c8FJzaOQ9hdc7mkgJDAx54+fcLje0wdjXqn3+j+LWJjxIR5H5gZSoIIW4T+GTt
EHyszkmdtLYmVpoSdj45fIuqcP+R4Zx9yf+BUXH4t4sRxQaQCO1mo/SFC+WsDMAw6kFcrzJpehV5
ZvhO8AqGV8eCelZ8uxfwD62C3xp9tVhUS1kVB6ZWy6lRjIeNUbxtRR7qE4T9XOpBkuxzt0tfaAvc
ucLnP5uVACz80vuZAtyG3e9Ymmhea3JoC9qQ9F+m9/VdfbptFRYjKYMsPToBS2kt2d8H+e6DoyTz
Tvztx5kYsaKARp8n/tRJ+QdX0kpgoWpI1uFhQgw7D0nAsWy0O0Ejl8i4N4DbyE1Dgp0HMKU9ffBy
hRA7I0YelWiJlehaiqicxRfIsZFRRN68zvZh/rMmHoufqPJhF2EC6sTO2sjmliYcxGWpiYIh0wsF
MxLsvNPXp+TwWVXJ2Rc6PRE7IniSKNIwaJy4F4PROIkTT5+0IVO1ItwlpJcCh2JWInamnnVF7CNS
kXNFRL3Z9zXL2mV2TUr4SgYtT6fZJ9870ZsqvW6PobIXBnpoB3Ady5g/j72ozqSSB7CFWgDqDVLY
YkUXpJxSPmzWO81c5LZ4vO6Z2IEtlEVFRl+zRoD0YbqH0ge5vJVyi5iAPFRR8Q+ksEMA5DDkKhxf
8s1YZDRL0Ox+VZm9PPM3xTK18frG3loI45wo74gR/8rjNl3r0YoxTJOj3R8s+oA0I1aJlYsFnexj
RBDNL/jj9O16RFoLwRD48OFlqJyAkjZALQVz7eLHC2N8XNoUI1fJtXZUyNPKYMEIdDDGkahKDKnC
7E8dwZsGwKUTCwBB+/DTGzGyYjGo6FKVvQrar0OpYoF+nTgxmgEjTRctV1gkSlb/WsDcN1f+Yc3W
zE44v8icmMsC0uFWWSgMJ3RbwtyhKa/f4guKIKBXba50zV83jALwSmFay1eHM/SCq66a4MdlZ0Wl
7yHiMvAD+5meVm8zXyNblYq+FC5Q4+v3prQhOQFqTEdgBqfIyZ0nne1Z7MmPF1+qFp1VL+psa0L8
FLjHkDsFi3vaGIzmZIHEIXHcsyuM3sfBbOfr3Ted9hfnx/yZ77OVLLaVh1sDgj0qU/TnOt0mO1Jn
jr2nrE+ohiFGpoyILc2bG6J0Yx9zuseeeF7Ysp0Go7vvr+umB9A39rgSUOxUBgoJtujw2KQGlVvC
JPpsIMfWDj0aipBwTjVCtfopgGI7gVWgovY09tsg4/ZGddEosWd9q9lQ2BCzrctUVTbz0UQO/gEB
jR2N9oB/cItcRBfTuyE+71zbXieZqj0CbjB0Z286U3im8Zd+wPSsJ/+UKyNEsVAlsjUvDeRYSfBV
fYr7beRQO2Lbn4gIUz237tF5ttrMC4s6aHUyKqj5k2iIRgGkc102qQDBxcchNdnC+Do9L8kf8ZwL
Em3Y/p0nnEAf4hknIeHtOeppC80p00WN7pMcnWnIiwIoUo3VBOVJfnjBNOqMEWM4hilOA7uBNUma
gizrK2OktDm6p2SiFeN45ULF7IKaEXFi66QkBy1a2817q2u0J4AVbR7CKUemm34DtI1FOs9V+bn6
4qKX9+tbRzI5LHF7y0v51YUrfxV4eU8UTOCpLq0QPzjh/bNHDBjEoweacam8Ard2XsMijUJhLIsd
7rW5w0DqBahSBRqNIQUvueCfoz5pJPpelcbZe+vinrp4w51m7z5pfihu6zqXW0JbiSKgMNr9L7Jx
1wl4iwCvu6ayBBx4CjQJQOlt4PZdtA4uQ5MDWEN3yXIc3XSYGx5mt2vZ1KzgXd2SezkKljTxvTV1
xuA6DaOcThs7YKWE/cuDeI5LCvHhWJdhTRgt4fEv/7xMU2MD31zoYZWZ8bKwHeShZXfdiXpcQOgr
FU+d0yD1J3PEdvqBajDtlTSzM6G3dghIHbhZK+Tq/d019wZnmsQYvIfy0ZtvTyFg6n8u/aSuzyBA
ugIhlCcnEHCiNrDI/B6H6zJMptx2042ELfV0/aN9gAN3W24LaDQQJXZ9dli/jz9YX5MQwI8wRGUa
0U9y3zZ913yANdsAxpyYKs5EGRHPwb5QIUbyJ84VmBgJWuUZ/NniyvxLorPGviGXSHVisi94Ks2U
RuL1vQc7p8/Kgt4MF0a9VirVJshQfGfMt3eHxJTlSy4hlL29ChHgE2ZD04tevdVUWDa5ADfWG/Pc
wawSy6fjZEBl+30CecniT0WH+REwJ5Uv0mQJimd/4dADd7wXjGYnj937MzhGBmi/cu7P6SVDy/vc
XBZiXsx3Qz08Xn8djeBwt2/je0FeB/GK85nOI490qID3ocvZt/mWOtDhTcqBLdPRHoGqlRbgn2ka
tOSj+PSbQClZTTqtfHLFw83/7uG1J4XvafswMlt9KNVYqrGIsACy5zJ7aykSan/PWofta9H8k0ji
ShgkeIstnKStmYIY6gh/zJOyFBRaju7ssh3LoPh6DH3DEdqHaaCrTWGJ+IKqcqSWgn3EJNnSUBI3
x4L4533NrZMcdAFPFuIlFZzC2T77m0gCkXD0UZcOlmxbvHOk/gf2fv94w/s8fwGUBcve7b+QTxzA
/xT9SGe26PpbdHToNOWx/6brXSfGAwFJA7bIP+iuAmvfLforj00FkNsoldM0qnF+EcAtBAC7rkma
JB+aT5pOxF834DIQIHuRiX11+o8X/FDRB+iWHL/YQEPGlWOBuwvfwN2vZqchvzHTfJQUNTWSyRs8
AgzTYXPiSwIzZce6G10hSQOmnmF9c/RKWamlGe95ISPs840BR6WcpFvbwfQSC9xsqHGbIvwGEiDL
CEN53w+4TBhRehJT4eZ5TSNBucmE142JuljB2oGk6U8XyPwCva0Xj78D9ddiZRX3NmvuC0PT3qhx
brg1d5y9kzHOq/0IDEQcg07vNDRPVn2ck13dzOMhf2IWoD5COPq5ud421Px4Apx6XIzcokuwW8X+
RtpU/2J8GCWJDzC0uUhQ5+PyQKfi5ZPbcxObZVwU85N9IBgm6JJF9W+BY4exOfH7qOWK4yRQKfi0
YHQNt/8gvqhQZkWoVx8tfD/KlwmBlpWtsBrJ35gq0zhGlHNv/n2QQ8Mmf5yv+xH6v7rXHDoX1BVp
ECJzjYwUn0Mz9LDfiTO2mpBHS2zmgLTFG+FAiq7O1flRkxdCWf96ogJ/JDIilYPQEXE7M3UC+Cu2
ZXKd+CfL3FU0WaCYZMjV1r0e8E5c9ynzUwhG02lD6PhwaMkf9HBu1e9gR3FLpwOvlcgV+Ix1R9bs
hDdv/eIT8XhgsOcRsdaC8ZJ/Z7EBRDKEbwMiggHh+QWxNF3TCjKDyeyqBIO1bipwf7WDIHI8YqgI
d1sVmnzmQHofzAL7t7bEuZx5MvssRWx9MGfgUXy5VqEuvCc8tSldbEl9MFfx4rvLEyQBoLwi+7Oq
9cf8lxgG1amLcGH2J0K65FRb5XaYsN3ufjkiDAOvdeipfk8V0Crjcwc94sZfdwcih1fZMCvFPS4e
MOt58B//oSA+E5u+Fzo6tdoxkKiZRRsWtIHIkGh2a2dI1SrO9J7CUH6zAm3Ib/Nd7ky4RkCCnBkI
thaSkQuhTOUUDfz6F/ZZH0N1Vu8agdjmKpmZ3DxmQ7g6TxpsF7msDpSviJJ8RB772FGkuTBaXy+R
i8+r6KzV4qg3BIUm7JHga8wTINBWrPganuhX6xJIba8gjoT7LUb32AdxHf5kWQ0ru4iuMmpeswUY
3KtDM1OfibsHE+whSewkGdyyJmfL4r9lAD1Ru0tF0DdcC5sz1j2MEzYFWHBi/Mo6cDrrhJbC8vK6
J76b3SVInU3E+JPnvJalKfprX3uTXIELdHslMpkP/lLugCIuWTzBSNH7G9XLDQg3LXogXG9CTx2d
eDzyJF7rvkamLjwGwcYF9oFLllHUZU8MCiUZ1pSwjSJDsin1Js7kL7iPYSwEM5EZnDYMOAPaDffh
BYYVo4ZHGwWQ1B07M9ZVz+b0U2j21knpklYq5cOmUw2nE61/xD7g7uX071M5c1RwZrSaZRVEd7iS
q8OVkhz0EDAxfwpIU5TllQZLTbXo0CAR9iXVhuolXM/BcovWYXJqrWbRopX9ocO99FGqHTOVA5F4
7iZlPL12SF4WYQ2f+wxaz68oEJqwIK4Z3m6muq27f9lj2HzgsAjCEMo8qh9Q61lNDzdPn4hwykFw
OxmMIzR7x+CzOfejTZMcHC4Fg2zEM3Ov0wlU1g2PO7bgZRPhVKWQ4cn1E+123cYQ6xOva521V8jp
tTMLeePDA2eaEDB4V9Ka3+apU+gwI/q2cXlt1ik7oDilrPsWJaABgFPqft0R7jfL/QD9DNyE09IQ
y+L9Qo1BIJ6UZ5tQOrtO06i0B6mTL+BDvD64YGDO5mBM2Q+QQtLcBHi3iwmmnMTi1QjjGtAtcJti
1J8pPfz8ui3h2B61NnQySQ2HQBwfpCdQbI5mWzTUkzWaBUtc07Yah/EXyl/jDtL4ms+MhWmEeSEo
t3XWMKUEGwWmkrzdRCezJwGPUIVjKUeTam7/CZZqZB/8UL3HwG6sTe41LWukHudSYdR3goFdPDh2
+IfIAVEEKQGWVthv4AIxi5EnU+nfciERDESBWZuj7+pa7VWuIAnAtXBrkk4aNYgaDT1FsGkavIw1
Wd5l8GZBtoOh0gCoxoSdFfOvjG+BSBGDMrHF7Nas6BKQbqgINrY6CMSpjmB4Ga6CTd/rdU0MYvLw
MnsgmZQKosvMAmcEe833cqEz89kOK2f6QBq9K4U82+qgzuqawOUvRT6lv1WIF8P8O0bwY7CxXn6k
vpmX/LwYQ83N/cqzXNUJCe7TEE65LpuO8T/drIwhU1mGi2AvVwWTfdUZLSBG+wBNhs7oJ4ZDjxip
KiS0lymu3YZ9duTY1oZ4fIjpnAU4ECuNlOWewaw93G3X1xwE2WCk9gVpaD52c4s0mplX8StlMPpS
3ra6xRV35Mvu2MGup946GbxvaTVonpUCj5pCJRPwOfV0So9sa82TE8OnUT7AdE092aPNa/nHF3T3
gMdsdVXGHPJbYRFUbm0/VFukO87GAR41Z9XS78Y8fZHkWuOKS25ZFKCa3SWIpeJN6Chc+AGJI6qO
m3e40VMAAns5XNWmJpomji7G8hhELkWn84DKjLVTYBbhYDyMcJETtiDkwRbKHT3vDU9p4khT4ZVV
Cpc2fKSjsGJuec1MN7st7MXV6g2h2ERxcd/rXEyagL6wtSPBJwfYi944Tt5M4h2PCHqjImeuaTxA
Il/u8DILI1nUPLvB+n3TZott31cPsdUhEZLBmXYIU8GLbLyKrdP0Xp7m7mkFn0a5G36fm48Ttftf
oBTrnZFcYFkvU+IBPTAoyg/eWn/Ma4Rt9Jm7UL4eL7tTzFeXXQ0AYLCOO++bAYsRr5KnaOf2fA33
Q/q+51dFX39REEuodPuBylPfZx/dSZ5qVYZGZw+6D0leRZY1FB8zPIwSa1xOOKNPqfPCHrZVQdka
BNbhxJCfXOTamYcfn3WDiVm5AY0/iYLTKxT2yGuFQNi6r9Q07i47RZT874eAnGbEhiPIDIbj/7V/
iucLMSYL3mVBSuQMUOF4UPHFB6gwt5nAKtgeYZ0qv5zQwED63Bdj8+5rwFqz+5YEi2yzb2aH16Ob
uZoZCEDruNkFKapkCCHMRzn/0cMI4HhoS6VAUvMz5cOzz+WwGNRnID9lNz83k4vfy9smVFM3ZYkG
WDGf7Gl1ZKWj8iEuJPuS4Cg6LlJRnQOA/KxFwk8cDT02eLsecA2OFDoD2hUZyvJ6+AcCLqnSj2qF
cw+u7EICycrUhgIYUa4py16gc4s73TLZ+g4otIo5VDD1tlAwAMmzGxmNlAaOeBdIwIplfc9+X/6G
t9QTeOi7UKp+rAtVWCnAzFj5j2l5Piz5a2pmSuPny6fPIxPIHjVR2kXQKn+hlgJNVFFR5IuEjLhf
5aYvAS63p8usNdbkXYyUmKoIZ7XVrKtdXOuPF2fxmtN9rscGlYa4Xk6xGqpNLPDTSpY+jb/o/B0Y
CszNZSyxu/E6Swl54++QqI+NY+eEEPx+u3bJ5BGqucMFUdMh18EMS4VTKivqfk4YKLxVG4jW08xA
kuc7tVvY80rib3Luxbyo2G/E4Gy3eIJBnTkbs+55gx+uJ3tikOKQ2OaOvD3Rzf2niZQkkdBEcPB6
S9brn6HvRJF0NS5q8lTb3+DiH4Z1Yok83Mw9XH9UxjH7tceVaqlK0iYkH1/iBmy6+slhkJySkCzE
9MILbLQtV36d41ii/CPvAZrvT6UojIJAKccGJ1jJzoWbUm2hIH4+0GIS/IgL/5HvjQZ7PS00D1Ps
f68C1Uq0pJJjAvo1nyoRe00rNC4fwoZ0fdvxZXnRMTooBI/X45nA/ymgD581VTvY1wZ1JzWRLaFK
1g5TWskQgmwnUsKJ4gChBaMq1zYMwcq6uU+my5ekatukc0OfbvEinKzbBsXDJ0k9WPxcXCItsr3s
bV/QzZPx/5d/l19I4UCm4ykMtFld6roZ79pO/AF6+fSJeUKfhpE+TFVHqokqyvwg0KuAKLxjuHxe
InqSYAZuFqOsTtIQLis8xukCFIfHGq/R4a1SJHE4R0g1CL+JYuGH7WY3w09zHgUuaSCGl5D2MKvt
rDHunYnHWf8JlTsaHUKzl5G7A/yWokb3dxxya+2Y4Ehe7i87yqDr0BJ2YfDfydWlFghlrWSCiI37
UVQt7I2AIblbm/6V4xidUkJaKJlZknetyhdQ38RLTWs8dEbDrEIqEQonyjT+0Tf3jZVkyzBjPq6U
3dIr9gVa9d3U4UJ0e0pmk4G8T6M4hCA5QjFCv8uGb0rEt3Gh2+pme8czkjLPTTkFlrBN9M5hPQRI
MUofKj5vqQpc1qg5hbhi9xNWb0v4uGJZcSBOHgHSFg+P6WTR99lQWrGGELwBH3EtHnU5rW7p18H6
tpI3IweuxBJ5p2umizutD5nCqX/hBh49mWQhXaM4JyVMAQmTb6r03bVFWOVxuXyKA0lStQm0+LOg
d0K3/sF8XLlZwHRKTSGy5dh3hipU6tZ6UUS1KEfOsTvhzR5ET3scLSd0+rk/rTIhBRWxghV5hCIG
jAGnvML7RQ3IFn5zdbfN96CETNfEVAkpwPE8vwwdESBrzE7fMsVYWbpsW9QDS7+8LvNduvKAKQAQ
swmLTeP2ig9W8covPBZ2XibqLsjdXVvCnPJPLtzrDubZFjh0kY1z9IHZup4gXZ5ac4kaLXNeEvLu
a3t8xeUPxJgiKbtVZ9Ul8cC9Zn1wZlU8LrLTnGx4MjoX7ilqUx1VtiqEc3Bk7p2Ydx/IFcB861oa
i/0LYQBU7rtSOYf691SUVRlRbSw9mflpn+PLxGHEXbNtaUf7DRRv3/g+GPMj+nGTj+v9G0PSqZUr
tJP+UNEkyarVKxg6KyrJ4EGIuva5x8FhbxNjuJC3ft2DstsfVkR75W8atgD0A+ObQLVBalmdMZ9r
iHxL+0SUOj8tITif7JCNjsGYplEwsjG6ffS+ygqkCvDQ/eBnLUbB4aDlX3VArdWUd2UIvlqbsHF2
F6KXtIvwQsEMYRRks2/aEcMe4FUzlPWEsw08ze0cY4CSZAYI0jcynAeaVxjB8ALKI5tUyjpCydGS
bC9IQpw4+VOqBIsdemgfhp501pFcvhJRChMyDxFRvLifBkeYD0hn6s2cl1H1PK1Pbx9Cv4aBFNJl
fPznvJ/5CrfYc3FdFzoB/lkKVwzlcZUaB5l3u00xAQrh8EnSqO/JXLMQzkGqoZfcyx1eJn0xrG4f
cYOoYkY7BB55ZZwFKHUCz/l5Wc1VM3ikwaRFXZZwK3x1efSPBgiPMSgi1RmFPAE2Vbhfg4kjTRvw
fLhOZB+rH1qbh57HIxbkYp72n9XIrpnavSr4QUnRBrqOEALK/zZn2naZ7anvvVvp1kqN1jALNDmg
PBsWqhOmMdS6Q3ZuYyrT+uPXHJQp1XP08p9B0vE+S00woCsdz5ZcpxTyZ0oBNlBK7hIB/etx92J+
ow/TDm+H1puWL1F/xX1haQWBzfOcR+r9bgkH5VBtGcSVuwbi9Amjmx4VDoALupVQvK+X/dmhrxju
7rsJEfXtkpdA8V61FwGCfi17Ih9SXuQOLUGQGNwqUk4SpRhKDFBVj79xcDynst4WKEH9FzR/+k7Z
3K8jjEVxfQbdg085agEMbMlazfPAJ+mKRuqm+CGBtPC3n9hkXMUFcIG6z5H8aZrYCR95ukzqgf4t
y774ZaJvwfSVCcBIJgQN8HIv9QDhqOVMO2xl3/q+SlNI/WDlObbzEjDWT8DwPBV82MyJVbBgyqNv
DIjvOGcfFuuXyi17/wkeQ4rO0LBL0M/4ULaNYzFy4/rgxXnEhWvNj+dR/dOqSgJzYpbXZ/8KznRB
8WLjdnisBG02OGPNt4RDknQp6V49CXDXd+RQ65WPWWbZN8xQ2Ev/nBTVbk2GUqQ7XXs2oBIHhvVT
TmVXu87BSRMRQmnUPrZc0Xvi3uinZfD8cPl/HdRM+QiVxX3ppos30hJ0upaeP1vkGy1D4PKWwhXM
hjBebWy7YYX84v3jimVLRuuZu0xNqCPWokTJYmfKR7g5UbGBmp2xADjuwbBTVURLAkBBS5ScJUqT
2Vb4P9S6nOMGSiEiweR+EA2aUVnM5EXtMW+jHLdP02aYtmMZNvG34Wf2vtzz+Kp7fycu6y9Tw/71
8yHvzDJCQJKGgwYcN4UbxnvZp04M/XCEubyfDkmbElI7nW4wJiAt5v6+T7PPALMpPt4smFmXhh7i
v/TLH5B32eK1kvL0ZysPaQYhQkr+u0Z7jNueRFcuGfu2t9Sujfq0vnZricidAc+bzbsr4N55cxBI
2FvC6XSE4zwEmOranZyFGDjCcY4fRvpO/V0vGvFFg0FRhnKlTz7dp0nK+05xsOfAlcEw/N7xwH7W
x5s6KTdzEm+KDVALT1uyO9KD0N8FpLuY3bD/vvrBtdJqaU/gk4tGhVEvQilvhvBu/s2zV+s3xDZm
IHkCutEkrn7kyReAGIfpqr9+x4J67J+Q1SSiJ9voeJO+0V6GnAAu+R6xnqJuX0MRJ/UoD0xIGi+Z
+j2cahvnTRMX+XTEiPEsbAiaiZtGVJcdulkz7rvz/rZhfNIMpWfLVOZtOc74iLU8O13dgJ6u+R6p
2vAYJYSkXoIn09i5gWiopoxbORXF0FfSXHve0b+lZcwIAOsZBy5UDtHcwu+odVrvd5Mjxn/2ICcI
fe83gfrL1O6fHQncED1oD3WcfiuM6TtAsBvSoA6781fIihByTbt1CtQmZXh2VTc/rBrnzLhJZtOH
K7Jbkq9apaZGLBrFGxJVpbB0w+SMae0WqenkvxqbVkYAAvFRRA3/I4NKUMJYKqAobHaMoz8c8lyz
PoODm/ky3xd2UHUukzaEHPfHm67sOmopOEGj6ofHt+zdNCVTFEbFxscd7Fgex8HztkafH4aUW008
58gxvHa0q8eWaIzwGCnBzIJIzyDa+Jbc481XieSnujVhfuTiHGOdbGkXuhz3TDqp2/jKqW8Tf90q
SHPvvCMam6VLr5YDmB6TM9e7+thIOHyBHngtW4AlLOdG57a8v7aIWP74Yqz+X04cpnuQ4qaJ+Edt
U2o1CMC4uUZd6Z2Rww0WWLfgPkI8Bo5bzEILanYlr4fIaFxbwMXcUFITLojD8NvxgVv4JC50/2y/
uXNP9FXIYxKxHU8crNribfjUo7l8hJPLUGrSCxY6n56FIuciCj+w1cwKCxovpPELUzQE/A1USJnL
Wm1VL/bQWa681TaHU1L7thIXgHoNZ4id74h6ieOt8eAxPggR6AguFoHDZFBJtctXCu74jIdlV4wy
kRb1n1p6givj1b+kwYxQDFMJTVhto0RDs3GBMYThOvkb887CEVKLobqTJJK7Ao3GLafrpyKWUHO0
eKZ18EK5igACLUv/0YdiM79ytvL06MceICWWmilKtTxnK9R20tjD0BSce0Yw8+6DB1h92LDmRenG
8Tg8qBkkYrsaRcxHUF6hQNHjhCTMOl3SXJqALn/0IjuRNOYqpT7nGgWWGi3BYCPofNyR8s3m+rM3
whcjUKW1r0O5LTZQWXIF/M1uDM3umF5wfdnX2bANY0QtYbfQLfoyNieASDVTKv0mNOlVJlbqc9OQ
GFdIVuYXZjSIenLNFLe2nB1FWzPifTafyIe12F2FFUj66IyIZuF7sgVI71/OC02p+oeIiOP55Xa6
tCroM7MFyhdBD7g3hZl43NQ1/rmqlgmr2/byONyj1na7qsDdqD7NaEpR/fZ9pLSvy7AU9yuDWAlG
/Axro7VLgCjz9SbW8S4QNg6Jl2x6xF2902KU11qjM8bMymwhaXFF30cBOJrr7e1qpTUIjkF2IF+Q
HM0PoDt5RKahzivG9nkyk1q8n6PmH2Q7xkbcohOb0Q0eC42ikrAorr0ClQypZl+mdrJeM3AMzer1
ujQER959HseOPDQLNjJTo2J1yAnc7gCyic44HQpSh4rR/wIo/2jP6r61UHdIPq9uyjytgNlHIwqD
WqZxKjVc3kNCIRpoiBl0Xi7eXkPpvBD1wn8zvP3wsDiNn1Ea8MfuuDQv8x59Rhs+tok8If15cuj0
SrlHRMXrzVDLPgflyNBdPtcqwWKVEks6nt4HIpfVi05CLNxF6KDmg4JMvWVtsSOOW/EtlKGcotKw
waxb3ECk6T5it8Jusmk4jzlPOtW3RlrThrn4owvI01FPKYNU7RO3meXtYldDuF41e1KutCq4DpzA
s8zyln3NjsMI3o39iQAB6OohoaJAhGal2lY49UPMwE2ZOE4Gy/s6UhWAJH+alGf74tADBOQ6dlJ/
5WjSwIOLK3EV2tnqBtm1lT5Znv9uzttmOvdewmVTzpMsYMtxTRU4F9/TmYusty33sDuuA9d9mjM/
JRLPYwfrKmpXolEnpfI5Ft57Gye6WJQewHUHK5cMFKEoflBG+mj8qeKeGr+Q5bbOqkKm5sm5Iqbf
bDt2AUgWmmFCEH5JD/15oOkHofdKX/RtnQkWc63CENeEVjkWhV5Kyj41XkOGV1uhMpPHRhOUpHEk
ExqQa77cQylWNxUrLnnCDVFeUr2o+yiYHxbhletOFXYFMhjHvYFkBWXkR55rVMi6iu7yHYPV8cWu
NpzwqueNswQ50qujeMPcH8cL8M3f5nall8NQ8S0/UyxfZ+VFl7Ito4CrP3HOyPh9OrdVzU/1AoL5
/427UpKFOMP03BrNmeRC7zq/3Vwr5q0BIbyEqjZ64sgKYhQHtB4hJSGAxcjNO6igp3/hBgd3mVQp
7TdyaT4tND0EnBEFBB70djEWZ0F8yVatVXBI2LWmQuxMerH6vK2HKvBOV/EtG76EmnN/LqRfVqjn
AHBmSJIM4OlzJF8D8jA5PQh2kQ9cmi6W0l5bl2j7xcE3r1+v7/2BSf24jgZHYe9w6E+8tbe/bF2J
NEDvKqcC9BDFYYFjah6rbz7/jxGmr8du/ftg7yprG7wS5jthHAuIswOfzeOz/zB2WztniPD6rF/t
bjfIK0mtpwgOMk7oYXVad+kbckGDnrkbAc9ABjSx7AjxHrGkYXlCD4chdjxZlGdutuNzvZdQFxVj
OVi7HaS0Ai2JgMq5RjMXIiShHuwba4pWP+kx0Klku7CLg53F6sLFGOsVJWgusvLh1ezA1u0d1oyo
CzK/waTdn6X+q36MowaPOz0ztnfeh/DnV+1hcQVH0/oNh/15cqC8S4qVU7c5nLbQ9WOFBRNPRF/P
6SlO0qZE0B1UxDF/wXDzm87DPTSqzAegQIDoELh+M9lZ0etN8nCgN+qE40Hh0s1hAb21Y8IVLFcr
9FF4sBQXA8v9HZKU7IulEPUc4k8H/nInti9BguC5jFmiHyrhAkI3cNMst9kyZrLKUPUwurcslAY0
J83fi9lZDL+/oVh/DD3Uj0eVaNkZ6OZAxTxuPR0QY7Ehh8wKCsck8BcbaxeU7trRy4f+orG2QW3O
KUEa57CtJyS7cyExwm+gD7ntd0I+5fxUMAX2xr6zFEQSAplfxaRinNRDbnuevl1/SS1/WYlrjifh
S+g95Eic3zJLq8I86y20Nvzw8GpcNnvj2qeAI4JVY7Fhab7z2K01V6+MDZPZ4Xyw0anggJFKkpat
kXuq6SujRLTFYN4+naoeNNOuw7ZyytI+susngT/i5e2TnK3POWXKmltYavLErSj3nZjMa4OGhiIY
Q11gINmdg4Rk9NFfxPQi79fHL3aJJoXJn8xVMYe/DFgLhCtR3LylWnvEs7a1gwraZLrzjMozFFPL
dQwzUH2dztTb7Nyp8TKp2hh50fjrkwGJRF8s485ppZlB1XFwxGCh9hg8l5NlcW5Qy6MuVATjZomi
uoKKq0TWcm0K1YL5qlJeQBTWOedHnQp4polzbKXSlqMQM17nA1ojn2ZUrS41qbKvusr6bcrhjdht
tICy82ugO4G6U1oP/RaAkyC8abwidPXnf9P+6fRlIG4Z1Z8CVNFA4G6yA/0HgHCXWQ0K7o6FxAff
U8XvWqo1t/tI2Dz8MakcMBHLEi6htunChpuh/+0to+TUgbO4ZveIUFlLUUM4QElq7rqDIHwH35k3
IUzo3P2/LKBR/3JC8FuNrUrhMvo3YLwmjm9E8ruIm4YFRKo9uW7EhsT7bwgARbkCYfU07FPiCFf6
jHAcJJTWOXoun018cQ5ceYar3IyZOT7R1fS+CHa20mn+PorPYqjJOoAa9s3HZ7gVIY7OxOdF0mTz
qw45jVjXWpKReFVJVrAb7jzSdxQasVy3ul0F8CZa0neey30A+6KWExGjtrHxbGOuh7A5y83OIUpi
kyGEforqk/SqV0Bsl7LUVk3zuxtuCnhwUaYjE0MyNeiZ6rBD135IVcbrAI+tQdcs0/fZPyRvz6vb
+GiBzxHXuM3A8QChGi2ZeCP+mJ8XC7E1/d0W7T3ooz+Ynr5MFbKaahgTyk2WaW/NmqgWxAxXgjJQ
2NMa+oBIQxZ6AwvmLqYCMEw4q0bev14JsWMuGkTL09F1hp5xU293EyykGHrgV9gt8J4EstpCsDeg
XUPKrT5f7TSupKxxjxtVTQKWmxDPWBUO/gk061lg4pMSie3x2HUUeDezFEtxA8jtD6mLbqk+puVJ
HZZsqCODLSKfm+10TakBWkD936WG72Bs2jLj2uyoBbYftOQR9PlMJynn9e0cEoxWwfX1kEBKNVIj
5Q5OhBO9maisWSyTTlgrQnr2tHnIcA0BKiME6Lc6fuka+v3p1SZs/QqKXrftxr3Zx1+hB8zum1M3
qjNccbutCRpv99dofgBsWELwUqfYSm3jHL7dGYsUMiPJXcQyWpE2LJHfHyYr4HNGBap0PwCQDPIO
ieOt41rvqENn+HZRofb5fYTX0pbdIpLuF6OreX4xHlYCBJGUEvrxj36rp5tEZlxWjf+XffIgU14v
MOK63SEdgN88CbxEt6sZc+RJDROnf2tD6LAzuSW4S/fVpI3tEcAaRVC6dryC6XMBBowCU81Wz9Hh
NXuOGmFG/TJmr/+hOed80dhSiHiBM5w2OLuuf0NpLJNTSy9FYeF7Rzu1cR70kj7+F322XVhu+nrJ
cFOmahl4RDQxfz4y0d18yEgTT8DqR6bB4ePnnvrxKTSndcx1bySN2tUvvnKACE0ZTciOOsnUc7uQ
oQI/R+0Q+FH2FnsTfrIwsHL3zqNgDJbqUCt80/FpbScPUEoF2Vn6M4r6NWtyPdLC8oKtWo1bovWt
OcSd7epG3i1icw7KlEcaz4fCHIw2P6kJpdGRaCN2Af+IpgMzbp6Q0jMSwFFUxWNmHDoOTEh8nEnF
9R3WmoDAoQurC/fANFFoa8NjESfwOgtfLL3dG8E+3/ntjdePAt27m/b6Wrl6fmjcQPun9bW9wCyq
xGlQz++dP+w4CsHbSi+0rtGZdQxqeHuCUMOOlGIkMyP7hL+so2UGMb+EqW+iVTR9c78FFFO0yJnm
2lcZNuY4076ruOfbX6joTsbaDTMNGOcPgCl6F4ghRrjG/E5ffI5M4ldyKT1rU0ZNVLHycO12vkZI
IixP7eyKQMzhK5K5sBX8qDDfPwLurLbGdqW7FU6iVtVEA/tahvpdiKVbnuE7IowM20FFdY3WIy/4
sBz747Fs7ptgKA+/UCmX3El+VFMtftx/q0wT7CXBYOCGR6v878idFdrztgz8dtW3L9DvQkX5Bw07
LPQpXYVSeA355/74nCo0atXoEOSyragMf09V2QMaiA9kCJ4pA41cK7rSDS85P57piguF3PbtpRpN
s7IIvU58XjRjOJB9m9QRjGvm/sCUZ9fqVP42jeCBC9Ram+wGuJMotjOcWdfK1v3tbzNax4/J0Yw9
CuPfumsFuAjLktHWbxREv4R7DvAy61Z2V6EQVfdyOL5j655aqp9DoQoFc8kTnalybivBALj/Zr4y
sztCN4UQDY56jKY46AhOfaf5/LCY+c4LDfNv2BDhThi2gUi3xMQMMA2ISTDXLl0uLGNji15MHGWg
vejtibHXI9lIbGhfFjtCfEpi/MUCBEE205IbdVINBM8ABFZ1NHGAow0KUY9xslowmmxdRbdYLQrG
4Efo7b3Rrz8tYdzYgHyYQeYL7w4qC1twMCgXGDgvSj3Zo4bHeDVD2Vj3TL8gzPd1XLHzgoif3q8W
745aiOhI/Ir6Z+1cgFAIMNVoCyLIOCN95lYy7t5IeTdlfiRP+8KH0tb+dYUvkc8e66wmNJh2Cc0m
YflwvRKjC2wYPgu7bLIzUrPE6+a+v6V8t2L3yP2X9ewQJG1rTStkZon8EF99UpKPDlFmEyDKE53f
amUzNTQ11bCHw6boDIMdC50s6ea0Ewyn6is6iYtzYnq5kLCizV9a1jkW4kSXdMfqCv2EFq2XMf3c
WSItUkfpMlkrlszZqfikc7LDoLAiros3UfMmGa57VZXaWMom31YrbdpDbEnNQv87i4R85H/if2bl
+NFgHBpCiGUtsPUvL2RBSGO4cTB/I9czfxGLuX+3H0hxPJyBt1/9EQ279cM9HDaCoJAMD80m7lgZ
9u87KwfH8Q1yGjfIppKfzsWq1Ax5GFQMZNiW+Yvm6kSZIO8xmsL4D/Yd5NumUGCD8h4eJYm0jH/h
0XB8T+Fe6Zlw3Ac7J/HGvbZzNpclS9qo5W+cx/QQNvGamrcsDfK/6mg5c7RoWo5Z+T6ANDSWnX/6
ujN8dtWCZJ1rxOCZURdl4R8lzg48TW0punthA3H73kCocfbSJu/XlXBvK+u6qqX1NnRdPzt6Njmm
kFwU3hR/xk1Tn/nWan/HCGxVl2mpDogz9cqFd02/Eg1tXejF28BsI7hlwR7MLtMiebZkYQLusrF9
clyaUEYlVypTYHNL26CwlwmD0UdqoAZ8y9rwIMFQceuldvAAE38jCjvquQfBtKh0HQ0PnQIK2qS6
HUvBbMDqyx8tI5h2nh1NOvabTjz/5JS8Irc0fUFxW3HzAvvGe8QhmF4PLD0TYa8kc9SuZrm1JmIi
Y1Ac+ib5rL+Xzf1VhhHeIRNC33Szni6E2N8h7BcM/CbS1s4jhHxYDpjC0XowySPSgMaFh/7Yk254
zLf0zhDb66uH9ju2d/2jgIJhPIP4ZJ4jVt+F2ibhYLtg33TXUlxohHWFDeicfoF5UrYCXwgOWtfC
kJrMuZG9EJW9Nawl7iwLW9AwkREsXYJzdNKl55yjaDrdi9sFZ3/TQkS+BkeSfPM1JzmR6oSEMQja
o7PiRiU5DW4GexrHsg2ObQabtluv6Ryhiy8iMg5PVok0YXrHSb33tnV/ZUtE5K4u9KpNDtDkHY0g
fF06cHMpaJkqQBbw4wuxfavEqiRx51NAI2KEvgk9TxG1SzM3/L598dSsCZlr6WxxJX6srvtScW98
b9Hs6JXPEip+ZRRePrchovVi2GLmRmHQkx87TzAXTDauy+f9+Grf/l0chz8SvnW4W1vDUIOnjhjp
sq0qxEuVxu/zaYXf4kqUmbnHW1iF0+F/iip9ez0RqNr9rAtd2DoQ43eFEEI+zOSRHGlFQg3Y7lae
6p2XGOAuWCmzOhEfOGYorB/El9dbzbRFidxhLAc+pvQaFG0kioFz9Sc8ChCD+sI9ILGHua3+2gPa
Ukhm6GVm6Jkf7Qw76IHoFHCq7nkDZUDMwruVRwwSaldKmmCJDUZu2KwFzKoB6cETlR9s2qA22yF1
V6UzfEtuUl/mD8trh+i71+HKRQqb4iECakzKB7Rqjxs5nvSBoXc+WbDkGYn8+fWnDaViDBiFzehi
BwoWRo+MSPlhk4MWFDiQL2+7T32KOEYRnqOeIJQHHhlgSGAdVoMZp7uCyaXQnlO7gsttGY0VtG/S
4tOBSD2UMYiHa6binwQf3sDuYuqTxfrGiFbeqmAoMCkDFim1HblQmKXqPpZmPiSJJydXJ5tlraew
mn8/CBWlpEr7jxMQbjqU7gIJpMKmiIWpMVNUnyHIl7IpjyBViVJ1wrzUmihcJn/JZT8lpQp32S6G
r0o5UmZMY8FTTKFZQypCUqRryVmmwAhk+kC7MeTT9mgdjxw71/8BWp+irUZD7qiPsDZyMAyrokIi
CdttApLp6SbloxN0o4eflCrTunVyYSfFSJY3mmvPZ8OtF/3OlesA8jwvwcWkggf8B6iXTnDQXzy8
NYewG/sKg3NbcERSNRyRQDFnX+taiAQoOlXvw53eyl6oMVcadnNGadGvbqmdWkp5BkIVHdtrzdeG
Nq9k4b7KJQ+OQ90WTF5dfsv5tI0hYnMOdXQKK1sGplYZbohYuIxkY+4/5PQlCj8EbyVZ+wlZpFga
S4tAo0RDxDh64SWh8kb0ZgNblFR7TyIWBEXHGClA7gXJKnkcqpW7B9BrwKDuZgAc1fTfLV1RNGSQ
QFWs32Ldt66PNhziVMLYe4IMCexgI8j3+r8xY6rOFgQRTdgoSO3/SRbr8Uz2ToGfGOK+OpLV7jwW
52qxjAvXS1sx5LKjRPSq8F2Mv3W/nifCCy20NP5QQtauvOlT2BUbF5qso2TlcH+WPRsbbGoFwzdN
hPrwPc7i6DACMnTsiJsNZmNPX9MqetMAuFwNLdvzk1EmK0nVHZZBLtteTELLu/cZKEMASRyaMY6V
jbbBYUpY2DLDW7zzPr4pD7BlHn+vZXm2GmIaWZU0A9DwtIe4EUBUjPXOs3PXecJKSlfRyAqUKDfO
EH5KNGhcV0XG2fL2Xyc/2WjjT4FPLmoetCeUD3C6ITmQOIf/lx2TThoRLFkNlg2rv3YJc4QCO4Rd
3/DbqOUu33rvMQorLsaYrrTbUjQsy4lnCjPmb1TsmLUnHiQkna8NnAVrfoapeiiJQAe3iug2lEUG
ICslThZuj5eydbFsdPZ8+79ML7GuBb8aw5a2RPrlGXGFtyblf886Tg/54uBySyvwMdQp0JKHk/GK
F+ROtRrycJXK21x2siGDSBvNjwt22oeWfASssMVLOHPe1pmwWms8YFOytI2xJ85EdSqRRvHR2cZX
8OBixt2FmC6K+39cUJ9rwB8mCVvogWGTG4/nbmO6GeGRQIVhUTDurXpGiotclNj2mRRSth6G8cBG
mypufvpOlofJbebXGzDyPAF3gT5uz0olnj3HcdJdcXsJUbhyHo+7DXmgw6iF1ucqAcDS3AffuVv0
dKmEGJgPRsIDcDR1UN2FMOUJ8BH9dompn1Hn7WswVNzNCEwSkNKAh+yv8rwCWM2QwmHzh0PYhDWb
rCoUHZNBpqYVpzSWVOzrV6XjqkSeyohglabcku02THEYk79tM5+rDRYX0ZxdvQ5x+8qwDxWTA13G
KpqrWja7xLKm3sv5i6AUjMoO4j/kpev7pJ3ZRDItLrbCG77nao+zkUtaD1bIeBkRnjPKDFUY6bsU
5KNucoBqfXcL01G++fNCRfDc00GTXW+uF53NSxAANdyqEVia6/zflFOQYncCpD5Xngif25L2Mwuj
rrmb9JiLxc5w6A8wEwHUpAwVBhzXFAamTFvcpZwWQB4YXtz1FRy1fqcIDZbXR9jWfNz5fFV2Gffn
9+3nE4XxYEVweYfxmXqk0dRi+LbRfRhF0XpSndOOHz7VRpDEdapxlZ8hTgLcCN9yVEIYOTD5lbwg
nsTjobtfXXDVUd9qHZhciUR3Cy0/61d45hvXDWHsFKE4PAdjsVrohqE4muDjgYsxQIMAIvro90Pn
6mVhBrB82WMilgXZOhZojRssDhwp52wzGZfEm+biF8H3eZpkmn7UERVF7RRS4zc2JTyN3DWHPYJg
kfM7jKVIZmd4l+ZUhhngO0UtnOFi0gACxURPK33xncKi/1f9VSBFBaCz2a7Y/Vv8pvkzu803LgDv
kjZRAG23nfVIfqiDGpH4HZQC8Pj2WnAPc62x1d4buPcGDhUzsxJYl4hAHhA4gwu0nPnD1YHKazch
p6cK6eiu15RCxPv4fXVCGTAv7ZYes2u5o/aAyy5LAce1a9aoHDJD/zpFEvJ7qOm0NBVOQT3eHAXX
HuBan9NV0NAFaxTraZKm5Az9CwMuGXfvq4KTM6P9RpBi+Ci9DmBm5lhGDkPCP583fpE5IzsmWIcV
AX1bJhhBXu1e5zsgOX1Tm1Ae/CVBYk25qK+6HWHVUzPMVXGhBADbfjEEfSMQHH9v+1q+4UN0NcuV
koppziocH8JnKeF6g2vQyxPB+dfH0fhBWvMeSIvOrpjOVSOg9C8O9Lgpr6Gd010GwioC3nEg3wVG
YVcTjPVgawQSkJRDbyOVPxiE7ro2Fu6cIZX+PEHAIDpc4RbSAlb9NHCwPJ9pJpTUKfD4kiIFbdhu
uhaf61bg+g4Qxpvx2UAcrcm/IVPeh+6iBJLPRS/Q3XZsWtVYUxbBYXCc96NsqHWrtgLqKcTGBzoW
eLVRqpbB0fbynOgdOo+ajsGAPvjZyx1mweKx89N2vZ58nkkMmgBJdXC+2DePVxbEO9DZhs2ZVXxr
vFaE9F0jbQ80FBCfV3KlSedlE1jevONc08sgwxe1TsrMj13wZoxuR3J1z3sUayZbcxCpreHYJJBC
c+k+B656yyHnEJu02qO1tuS3TYwjZwIOvBDI3/WVwlVxCKYDp2XMxb6PLfJRADEJFZbxkdNSITjK
SNwmleF8mLqhh7Q56QoTlqaexqlj7abDJDEm80O4Ng+yaWzhdavBamOA8bWpOkzpiwKoUDYsjHJQ
s/HOZz+tysQeN5Z9boq8Z8+5JHGl3Wyt3Lm6fGLI9XW1W6mhkHA5J0RCSSgCCrXiWaeB9WwDU8go
DB4rWIGtVJLl8Qd/0Fb/Wb+gJT25w23qCeB2/KgWQcsAHs12uKZ9m6pVG+nn+9OCIf5v+HFWwVXq
nxYr2iTG2suHw0amTestaGc3Z0hDzoSe0cbLw5x0eHGrEiWrC4K1/++HzQs7AfAILkNqEkqz/Kn8
czPR9xY4kKJaZEgrVW8cJMtAvzfuCBy35hwUSvMllaP/t4ISgc62JPkn9OwbpoqwYHEnHW3pJUV+
BsYXRiuNecl+jxjPvI04p78XHQiWGZP1F0gC2UoEsG7ESmkosI+OeitFUGCMbRpgkBZ/PX536wkk
pTXl/aXX6iokSmZlWYgdnPpgjHu1nuC/TXO94+vGPEcUGyzcKo93hgnbtAEZf3nyS0vw5MAvHwxs
coTOFbGlfStbweTEGY1wseaDfMz2Gy+39OZtM4aUJgfCN7F3e0/OWxtU8KErTHwhuV76ETuEg8z3
LypXGNCRtNJXx/MnFkZO581X92WHPl+t84BMVfClr3o8i3IVPO18Tmg5gouWfdsJE+7CBC1YzXIl
cerEeLjYSk6ctdp649720TYW1nQBHu+DIX64Qh54wzbheEKV1VkQOLBfoCiP3jpuEOo7H39+GCPE
WMB1C/y+JhOBkMc6ScrDA/pGRtuOn0/8aREdb3T2ru5VWDdMLAYGTJa4Nfnkk7Ofw3fBoT5ixbRF
fcLQMj7qi2mPVp3mBmafU3mOQD+3T5Bhmaow2Gq3MdPX1P7IFDvhzSjc3SB5pY6MKOtlYtorQJ4u
w/sRmVulj3vfpGSvaBHvhpodoVOBfTmm7tG6o/tXA/KmbR7S/Zi6uuJwA35xY6oOUpq2vLo0bzKv
l58pIoLCZi8rjjTkMwToH6rF0ugYOFT9cnLgm4NCBpiqSiT1YhBp/JMLM9zeyHOH5xJBD/4d22ll
rPJvmK9tKCPO8nq9GgiKCW6LimEIITJiLm9FmFfKDNMRkBTLp31jIjlfPbqJjIDr2xMLkvADfHIC
9WDMvmq69GrN1PMqM1xTvEWtpCrofMkQ/Poxiontlgors7cjeFyj0v6kdfrXMeRtJQjQxGD7L66D
FdFM6SNHYnh9jLwwcTZmJrAVq6BhDTBPwVPZtpWxr/dhMKHxnegmWg3cYU9/gFirij0+pPqeOR7n
0f0k2QNqVCKcAqdqJGQRVvIgAArgPL4Wat+g6BTKJ7L4WoC3/wafAjnlmyEfNGdBV606270gOb9P
N0vY0YxZYWNjvLSZzQZyzGrWs3dZpFkaw0iDriAljzBa2ViNIt5bXbnUw8at33ujNctx1/pksr2m
Vj+7/xXxYwaw2HVjpmSydRc7oajYy2rgVMvmvwdVFYapwrE1rxfU3uCqThD9HzQjvj6VQNCjcFUd
0jCGvIiFixciKr9LZ5ZzfyNPNqUXVMqv99gAEpMseawNBr0+ciARrQFSbDt+Ia7nLMhieLujKiKK
cqEBUJNf5Mnb+Y/Bk4we1NXZK9IBA3sf/bGxW8+hxFK1gDGoTqHbxGwgeKptQvr0D16rDLTfSlE6
bmS6CbXECiMLMFLRFWfYE9b8UOQymLBy7C2nw7Utc1D/lKEeXMbnUtk9ORWmmD2RTS0b3AOZsD14
6eYTLSc1PKcQHZNzbEZuIQLBGTdJV/9cwiDsy1RCEkR9OfxyoOt7/RdAwz4Bu0kwVj3Yt/81/ulL
s+Cz1nyM/E+dsMdsDjX1DT1oaXvUZw0gNVIvtmguSgjjK37OH4BWF1DCCLnLC2YGSeUzZMPtMgCZ
Gg5itmFye0C0SB9SCFbASK25KGQXIsZxt725K3zRqpKLlPdIVJD8XsjNtiN/b0yUbARtYkcYIP7E
uc+ulQXNp0rO36R8H9dabshrvtR8zlv8ybZg4y3Y/x5up0x25TXxewCE/I5BBAn9iH1Htc39ab5b
zuZ1+GRmljezpFvSgjjiDLt52VwkUrnF0V9PJ38ol3Lt2yigismddhrJOXbYb78/k1vkhXEMaSxG
E0HAw08s0asUo5yt+rZ93o+CYTKZPMDDvL0IYrrgZax2nfGOFCyFf0KiOuq1AUxGDtmn+vnjNBJp
UHKEByzT9CFy00kisfDTujTUuGC6rJaGrYKyfVUhsmRR8mj89ZZ9l/MVdzDq7ilKmutIzGyI9zjU
CywSFfu8kyzh+jVXIjoRMq6Co1rMGnOUxw55uCbMqFkiHRy3h7G3XKxIlVyGkDjB/8viEjk2sK5U
iq2aqtOWH/2NxTA4cYyXEuCfTYxIqxQb67BK9r4Lb1osHrUGsjZj7j2jTsmf9eGJeOTgyxNR3YVO
6MFv+OqEgpRhZfUUPluhha0BijPNFEhGsPg8j5ckTWTAkTETBbeam2QD8ICtSjAo9S3aYh8k0qyX
5mJ/6dqrhPPCI63dO/jK8Puyvrk73vNzp6KBuzvPwk4i0AOetkeujjSlv1VBP7BKd4PxS9sJLhD3
Rwgu3ftHdnuPYv+0vuhwz6P3NFlYQMcciZ5SGZOUkaoRA9nsvZuUvZ2JCM+15/o3spFWKEQCDibg
r4KnD6sy84dQxTEBpXYsAMm3uScPhqMUmChVCceTdwc3Xv/wyGOQw4dzt6GmYhep6uAXTlou+HIw
soClsn3mJFLt64lwC2xDW7qQ4e9Uzcn2anqx1HfAWnR18esHODRviHebn9JSRIE1C+ZqrKs1Js0w
kbNJr3qxLrc6WSVYSJq6PgB64PdgJuIvbkdXvcU9WFKDVwjkpyFVjSFmLNd9TeUYfF2/+VC6vCQn
nwIPBzDfxh35KZ4ffvAvKgsrsOYIfowhZTorUC+a8U6UmuaoW6vSu61aYg3SDdx52y8+elhDEE9n
WTahNi1xa5B+63VS3p+qbq4Kc2Aku+mn4s4H18wftlL/r6wxPk+glMF6o6sHM/EYUtLNqWYXy7FZ
q1Rqz8d1hKdzhTrly8wsjm5Abh1UzmK1VuSuq7YI1HC2cIjbFeYKlpi8UlKo29JfDS52T4W4sdEd
fQ0Lxtcp3ScKpUCev6bO+S4xNrTS1xZ4W8pld68nPM3u6Bhf7Qce8UGci5LL90kC2eGPs71mGPlE
0hV25zoDxcRGCwFDTTiL/iKzuxdtagPFr1VWYR0ROaBvdGCBA4hs92e3tgAljXxIqzi+bUi86I8A
+8u37l9NoIkULbqmEY08QePe/p2C+8BaModuBvFsomvkFanH5vi4cYEGmJu17DU1ubunSM+hoCSB
21TJB2A5/hscH/iTRzpKEV/HGORrXRQkttw19xSzN0C50vTtWd+ZXfsA3mIwCl4Q2WbsP1sHbl88
du6S1zYcB+RluaJXM87mhhRvY8qANcw8AJ2+7Dij4EL+bdlwBLQ0+ATaQW0Dljhaoi1D7O4z7y3m
RChKm+ywZWDq71AaJmudckoEOrM+3DcINpuCBQHPHAhwMWOTAJCC2fx9ALzMLlgLpxSEAtrHpV/N
/txrGmgfmSJ1AL4sCPKGxrbcc47pM8A9EMVClaHVIuFI6OxnOuskCFU7kkkqTKu+gXLnT/2TuJnw
i7Li4WLfEr5PILEi/Xx3dn50+i0Cmj0nAAhtIy/A5T35aatAGJdQxW7b6lHHIYkr3tRGOzKgQbax
bBdmVjxrWos8XeAMQEBT0TAQfLo3C5DKvY63l2QLVOj3UD5ayMKcpsVjX87w1aVBtVBkM09ySW8p
Mt93bLMzTeCb8Ftwyv/IEjGDEE13xPfVwUu9x0Jq2TVL+BNqms/tAE+cwA5avhDpyySqWJ9q9pXJ
kE2xTWDbwRDV4kmu4nXZv4B7haxxAxGA8Cb4fNDNHLM4iWmrcJm0copj5cXl6KoEq08SPyl3bLcY
PfD1x8nrwkiVlvlILfAD5QMyl3JVmKI/3nFg8h5tc83lRd+sdQhZHu7CAMm/g5SaRW4uxwy0YpK4
1NsdlZhbANxd9NfJqFIMayHhlQmV0nh6UzVXlpG+uVn6XqV1LhZgFPobV9qemqVulFQ4bi3138UN
+XTevudlNf6wKZLpofBrStDTkOROfHdu8Y7mjnbBRaSOxNaS55owRilLyIr9kIfiVkwBiPXiBgZl
nsiCmuXPF630FLsbp8iwB46GqCGu1GY4sOCKSE9BWasefFWmoiZMb0S6aDIeWEfn2+gnc0YzYlqy
3+0P3KRsIa1l7z6RiKGvkR9nUwqwOLrmrPiYrFucqyEnGMiZTnf15wFUOEKbTw8Y421LVjWlcYNx
Pa4JzEBI2t7f9QBR21lQY5j5ULOKvuq+QWNaNjwp1k3zYhKvaO+n9gDQg9uVyf2QZcnnaAH7VuEw
GkMc4t3setvtmLvfx72H4mPRXWkVwlmRYUUvQ4Kt2sXRKfQSM+ECEEsb7+pmO5QtwhkOEziPGsVC
dbLCXRgXcym1OdWTT6wOJJ90/0OCqwYIxNii4SD3YX6DrCfAyjij4gfT5DiH1Uf/Fwh6+paLwcB9
J9Pa8a80n0j9o8A6MM8V14YMdAWYiKTvIRDhJUuOrXElUWAHStLYYNoOrk/wAX5NAN1lm08S99Dj
ALO/ZDoLWCJXpJxwyEUuIeLRxHdZuIe2PbNQhWx7eS/ZBSg7jcNavlxA4qkcMhBV5vJkaChRQoGU
zn7rVGmLHMOvbNI/8z0U6ZEfeUwCw5DjuXM5TPRtCavl15MDMx429LfwLWdctYiE2Aau6zvhQ+z7
7dNGzJiTb87xqIjXHIqNHGJ5uvxuF37OmLKdzrpDoQissLIJFo1j36OTc3p480Q+3cALIAsMGi9P
vDGbdzePW/aizGsYRrYy1PQEwzLjY/glq82HmLnsO1yUBHAPa6EDjFG72CLkf59Gfb1Y2fyi11im
sRCu9WILzVr+numUv5G7CbTguTpYSeRlsFUy7nHkMGi+06HNfyoEE+wuQv/gTCuUPjSUqJ3Wpvr1
4/7swyiGKp5OVUjhlFNt+gi8RvcUcH7+jHK/xgW1f4xnBmT/b7vz6iwpVd8sAA7e2wYBo1YDs+XO
02WH4xU46CzSGw0D92Vtle2KWJoMpb/xOtTINmV17bMZqHahpApJayyta/2ArMt4eoolGZBd9bUC
CIIR+oO7NGqaLWzGXElsodgFNRchF1OOS1IHtnXFfxSqs3fsBYagVZORTlUc/1ZgBNJsrThvaj2Q
h+FOf+yr18RL8KNytA84JrTdLiVKKm2rTL+dFFFml3LPKkSiFCZG6jLSNAFCEQW0pHyMAfMAZ7x+
cVjszYWWw4BeiTBPJUBxIfcX46//sVig54krVhdQp2P8upUXs25pkMyk66yDLsKBPt1fpR7XAUku
1a78NgAlqHXkRxd49Xhn7duHGQce96TbXKZhegnG1bz4yhrbm9JrJPB5PjeT+gDQR2r2WqqQtpie
fQEUg0TLzlDOR4Kax/pAbDrkVrY1hLedwjXRaRStm8aC4G5Axc5f6SOi6u8RBmJObJp0lBDjJPVw
D5hnsQKiz07c/lVpYeOSGVgak6vs9lrLLMSjeFIrEFWJeiJyDf9pzc1haXSZH2at4h0OgqP3nV5q
+HmW4ZH+RCafCljakJbu+rpthas+3xeIrTL46MfU6Vi3CeFwGkCbu0JZtFHojUy2TwGjGojFScmG
sJhYlQy2JnUNlRXQ/dLXyNdoSxHujf/IDVEuoa01u35B9nRhEDHjBxYEYC4dA+o92zE1Wm5zZZMU
bnIXQ+Kxn8I06i0x6kPLx3qRs2m2kg9o06OFbtFXrsXb8qVYGlFWXYscQFsrqxGD+qqWX5DUFgIA
F+T2Hw4y4F3jO9pG9fkPjC690HMLam0W0Sh3tqP9l5AtowW6lIyxV/7+148yz3lvklCSR6aco2Vj
7QUmZE0aXeB0swah6HO9cr61fjcTEsTncHRUuEPJnhxE8M27O+YQnUnNtqTmu84v3Wixts5tdF4w
WhoZ2fDGr++YWffKd0Yx2tvuwN7XCNSyFm/2BmtrA3MUeMHoipB8Q4AS2q3aI0NxNbIhK4irH3aN
F3S7uxnvBknZU8KZnKmSuSep/nSQuzhnJu5yqUDz5zEfdDN2oyE42ceFCZXoFAQnYQWy+KI7noqa
xgF2TKW8dvZK5E9ac0fUAuXUOf1zrKxRuQ/YqOTLWT6tnfUt+2fA7UrU1MKcOCwvD4Zdm9zdYqzY
78Dpg00utMgag5tLzdCeFgVe1vBTyIOzKMiTDGJxy9x4sNcD/dxNS7ENziPTOJcpvSTXNKVCYk4M
0ZfVsmJHox+e6gazuJyM+9fgDbPgvtDNMVnrg10PtEmgosWDH+opqgNu/NCpLpi8eTYdbg3ICbEQ
Kq9Sb6bAFncX8JinOV/NVYYb90jWmshyXR5Mgngye5kDbP3dGD5mdOgWJFLreNiKgYCGAH9gPb4P
z221ZxUQgbncQaPwj6ONyi5v0lgc1Mbb1gPFaOhG/CHI4AFYHYnMNULe0n5NkXUUoJcAvVQQkct6
RiyBoAkfLPUfJ0N6GFZ58kTrm5OPqSiPCTlycK6CDv3AXEa7I7IklASKJPRsLLV5m5flLbQj/tC9
pk8BNfoHVmygAxOjNnYPn8Glz/FKNeg46DPD4lbNORcldTu8dL2pSip58m4oZlXsy64zk5fzqoR6
idaA+whLerycH0hNu3fX9H8vYhdUZNR2uvXSL1Y0HTvSUdH2DeK9nxzYJteTOjshFBMsC9EQ4eHo
mw2PPG7j3a1M5CD6ofpywk6Pcf/F/tOpj2XOe06jBMTSZnWi6ZBxoOES06RczzHSqzFFHpx8Sy7W
bXdzct5oQskRJkLqwgT3Is7QTcC652D6yLDuEd8P64DtcHlD5EhSyBMZiocMz3iEiae5ZZjbmEjg
fj7eL7DtAqZr6Un8IYbzV9858XB9RtvEAtJQ1oOmZ3cX5g/mgcGIIuhXdH2OJRJrJaEhu4IJdru2
sBfxtS2oWhUciZDSi76CiaL9YUWE5jj/VjFT9AbHWXSnwEj4HBh2hYZnYskUuTmWhY47vRqSRl3x
dgHBQ/RjSeNdLaIoE0k6rlR6t9rv0qMzVO8VPRlpcjeQYJAWLno8VrpOOzruUUCfpx8A9RbjAmgp
YU2cZZ0FCPeiFbvjbjlKPoZ+QJc4q/mpWqUJjl5GIHEsd+x37KnE3zPTnHXdey6QlFr2tdR0FwyW
tb1ZDgijjXyViRHBOWkJkTSMKcpaGLbcaFzVFjrEjmaoJpMZbRpa5JkZx2odTXTJaOg7Ls/t+kfu
sm+lEJgWvVRjW/bCLU1LrYX9l3NrFJP2Eju/16BTcb87jQCBtbOmgkFnggT08PU9aUA5p2DzQtdp
c5JL99O8biMmxDiGwehXwLtRLrhCH34HTIqvsUpW95sE6HqSDr09ooEIXT+/oczY3mbEB2bFPGGX
nuP+0tzoZpNwJAPZGhY+2QoHEf902z1xvMT8qr/o1e0CtX0RwqUtT+AjaJhyrX0mMAC5fGDlA2Ye
W+8kVkoreuYuPzUMpGP7TXj2NYplPy18Fu2J83GRbiX0Q4wnYMc01k+zmxT5kFHmq3N/gPp4d+aL
q3w4NPlH2YC6wAvAJIC2ckUyqAAy6fKhgmJ6Yoxl34EwumldUaTmiYu/O1x1Xn+q1/FPqOm2z4yQ
+//VkKCGP/fCNklHI7kufzERg5mhGZZ0stLLWckG2omCVy+RpjLmiGRKjp5SbA1BRE85aiCbTMOt
RQsPLpOR+LQtSuaCBA4uXTQ7pvsUIle/s0yIFJnWSui+ZXQd4TrKkkWxZcFWEu3sWcOs0lvT73/f
T3vWJbiUnpLhBWz17PAAXheQ3nzZYMI1bYY4sRIDPCEcczI2ETnqYqSVcQZXZtCsR2ADZUA921IE
sOWTKZDgqtTpY2RMFSn+0BTJ+Dg967drMVglNsGIuRKLFJAD/GA/+LjcnjKFhoxyRjzCVsF8H3H/
X3Mj8pLQkjaOZCpg0Tm4WGMILXnZ0fuQ9ocPyhDQMIRr1MhukFgbxAKfSi/6mRUcT5uFGLy05rAP
VpQsXNH+ySKpeKA7Ifdt5DBH63MRFk3L2nlgJTpyDMj60w1ZofAgOlu/byoQsvENrYwvjBkNnwW6
LiwxtCUD5guTa6NiIw+PTTlAr8NY18jDYRE9z2gL5d6pCp7OQkKa9vuVx7woNjuM+I0EdzhNBSld
9vv6hFaYNaVlHcoSN37fgkLRqh4kXrFEg2u0uUCCeoWc8H3t1fmCOtWE1dYZEP0S8IMMulhsCAUW
i97dTsgFeTwYfhZE6uaJrPhoqxbCruq4GeW4IPrJpHyve6hqHJ8MVGLsB4mTe2MH/tWrlJM4ulCI
Z+vtrslZKGgoe+LF6w6TBP2TGALyHhu7iqbxONDqz0J17jzxZKbHjjmy+CQIPpAEYXYislRTLcai
yLWeQo5PlazueL+BqfrRr6M4GbCQw9mJcOASRzen9zeS3AOHIPzQbg4b2gWsTS3rJjwBCGcjbmCC
VepniTZzo6xfDgeyP4aSwt8f1uHiPHB1wltYx3HU//8SmAxmBadxTsuUjsoDtX2r1KThS+DaiHVB
UF2unQksS1ESuEhTLBWNQTUtk2DqLm9YkXZkaxdkY1Pc0jH4DyNz47fHOWB9xPfBCk2AFN1cM8HG
m4KOXRdP0m4M8L8MABGJ7f4dvNeDxmZYjNCv5nMpLmhwqlUIxYC/VRDF/o6Y9m78vaRk0OgVS0fF
ACOgj3gaWj1Vd67671fxtsRHRyIE9VZKXxq5MADlcbyzEkAEzpHZB1Di0gYDR558tgiR7sqcubJz
BZgp1FlIPzYPzuHiS7ildQQSp2PMMiCWRbxpmg1UL0MTWfszel4lM/sj/Xy759hCrle05/xDH6O8
ufmtfdbkzxoTKRpxysoEV/gxiMqwRAsbUi26MbQbf8NPvzvdYTyS7LesKrO6Zo8z1xjZ4uWENpbR
hOmXj7jE+b3xzkXMFqeJvxB57CkWWhS8AOtRLN5Kxe1XJj/MlfNZfNGTe41nOeXS+17UQNDWVl0I
3gzVzUsL1BOOZp3xGEqb+dcFugM0+FB9j3Id9EVYnAzbpnOv+XqMV88KBYy4gsAR556QqKBrQOtW
qn/xirumN5/SPkeLWtWee0XFMf3lxTnn7XBz0iMGRRVYmvyrbJ5xgutdKMMANGJuLvWylpPBbihx
XfTCuEHnlwtz62SlNn6oaCUesWTpSYBI2w/hrdX9LwOuIz6xhWeWRe0Ai66CndbVpkFcXzzj3Lm0
lQGc5L+OiUl7CniAXPMTi2MQ+L2p5dDh5fnHvBYOgye8AasGZUSakgqSH6DLl0c92LjxKYAiKtz3
dOkO01K0r+9UpaqggQcdEk6XVlQ/WrAIYrcU8y3F5Fbpfu/fX1hAgpTGIIyMtcbGjhTL5qw0o8zR
z/wj+KGFslCq2/wdJpTuXZqKx14sTpLlqea9vkwSlgisWtthc5WIeEwTm1F3GVs+Xg/tKvcRQbfQ
uy7htQTXVyF6vEoy51AJDAfY23g3zFEKlqYnvKf1Ks1mgOBtJ+oJLwiPiFY1gjcPyKoEChqNcfke
fo8AEfsLD0Blke8VRUhA8DpObNBD8a0cVlXloFbqGcaP8N5SaEF0hE4+2jyyXzgZKs0NneKnM9Tj
ZOXr8WcBD04XYL+qGkrP5OaUox66kZagnDzYXU/Ha12dkcNTcC8fJ5fbDS/j910ePnIVI3q3U8xC
0ZNAiZImIzMpL+3KyJ65PPop2bImrHR58cDCkmYK/JxB+2v1DTmiM7p+329/F3wH0FNZ4DjeRI/N
8xJPhJRrXAxMgLnmiq3kpjeS5nSXrNLo4AgvTDbjqfmLGAUQn2DBFGiJhblBcu6ekvKOCTj9qb4L
VQ/it8/FEIZlXe+tLgzei7qI8ZUUc6qr+BNW3x9v8m+Ixh7UeLcQE+rrfH4dvCdzANaI+kQfIAZi
1afEe6UMl3YS6KrekMI1AzzXJna22Fd7TVr4IfTPW3A5ts5ZsBCeurtBHTRlVkBSHOBzP5tp3hyI
kkgHiBdtjBWEVJ18bDs1vrmn3JEN87va0O5wtekCQu0PjHCfyZuSFh1X8sHbtHS8mq8w0+dx2BxJ
T6zSjq0gozk1lWNSIqbQ3BZIKC34b0Aulc/ofdyqsmr7RMbVBMpZYV8aTDz2Ojs5MiAHmBdQOlDM
tCowtYkUf6h9Iay0iQNP9EM00bO1P6aausAXQbFQeqkeqN9Y3dlhop8eY+a61mH2tol+bZV9n0oz
9hmFE8RQ1Z7nEpf83O718AsVjCX4EvohCNBCumr1Fa/u3AOFW+ADyXAkZddUVrXW+mZWYOsSHqH6
z9hpp08G3i2atWfzHjAlM6dOc87Fo6UQFSRlE56yYKCQ5v2H6CY9Jo+F6MyEKHBd7jIG5f3SkaMe
lPEe55Ejgtn9exYj/EpwoVEZWDYg9u/R6swX6IbaamM8179uner7oN64JJMEu70NZc99MKvtsl8z
dXEuTmqQEI/JqDmoHgW0BSiELAP2fizj7Ndkmfc7SG1LrVK4rSg9HVq+pzXKp7N6OTiJtkwjffjX
FmOM6POb2+PMcsI+6x04hLVDBpYv6nZ3h0d3UwnqNDHPUm28i9+XXIEvXwwxn9hyKSF878kB0e5k
4ZakS9IYm1waH8AIeGPcK+n3xwM3kFB3QIo5Dh6bxV0lpp5ZtmiOMp7BLfUhMDoD1AAAaNcpilSn
4Um3Z79kjj1rFuGecNJt/u/HIFyoogcyszwe+4kolU5HY+yOfvjUihXoWSoBqbWI1XauI5rjvL61
PTR6EN3kA8AB+gHTegGoGOFqvHoTtUJMz/JGuVEkQGb7rwozPtq407hocmnEfW6C9P9WxMyAtftq
aWdwCcNtmEfWxxKGlZwS/IRmgjRnJfKcdwN3YKR/h9QpmU23dRn6AnoyNrp72yjocTJQyDjClauT
pqhU9gKnsIz9UAhJze56miGZJ7uzg+NpNkKI7uh5x0E0bVuIlA32MAHG/x3O6bAZIVbPGzQwWyES
6/v8CcdSd8tI76O6C4Kz2I3w3Z038bJRUNXx3jEgQrGVICz/45wL+yaG30uxfECnqDl3HA7jyLDT
iqBwUXGkWLF9HnrIPbOiahOVLYXM3wCHuTlDYmG1aS2RjU0pRIB9TuoMLviz8empPgKCyi1+I4Mx
TR/xQhPVYYjxq8+9QcK7Ozvwr//V90dLZXsTUiIpl4l9acR8s5poblIWWl8IxEcDJs/BFAtZtYIN
8GQ90v/tXkHz57SzZ2wMproVqr5YBZiYr357tAjKk4l8EitPxxcWqlUBvXqUrOaOwEeR6J4uuRgg
zi9LW8QGmggYYN6OUX9M2NW5kg3/5mwNhslhEhrce+zP93fwJWqK1XrZAcHcHfUtkEIZPkNRsnK6
InicYlepXOS8Xh3n24xgAFEZGiiEbSL7FLg1OvvTV6V71i7Hnur5VXqiOcyR4E8oadtyRhxB1D26
KJUvmdb+1aoDtS6oqQWZoivffRrYJbu6DWdS0L7oD/yUXw28K8IX7u3jMAT0f8oEsAucLc1Ki5Zy
cW7GijbPH7796RxbkZq6ueb4ed6Ab+3cIJ9LGCR1xmAFyTMfFSjmf2DjCl4dy4ObeLVm9OmKpZ9M
nJ2MmCvzvtH5GAK+izzdswf2NgRl3GNZ+ZWhM8H24f5SrOeKoG5YLxLxXLcbdUu6Q2nY+Zxywm36
wlVy81rFeuUmbuObG7oNtqOK5TezfND63iH9dBtrFL0VK9Gfv4BzK4Unv8SUXBvmtzwjUIHGmFj0
/7sHppA/1ymESDx3mwim3VZol/J3aHoS7DOzMaRKErMOvER+8QGdeAiwteKy7rPoDKRarBC/K+7o
AjkJJR4IfYcAX5Z3hu+hVXaKYAZGbsqfuK6uzYE0R2aZRR5zEQXx8/ABGw0zsGSUdo4+3ZOJFjUm
ButvekIjlez0jh/tcMUYFSA3pJ7O9cHGk/LV0pYucYh7HdzX2Yj7+GCBoUerIaDCXeiQT4+blIy+
EhReUFheMm5ABz2rV08tp2WTzkhfpJ983NhdenOtQC1pr+xPKzPALkhafkQhtzrZ+xhl0z89kfjl
65PGEFILERsloxmQKasaViIN4nC8OUsSNneLLu0PYXlc4yaqSahrjJTvFpSK88PU5lXAYnkKK/ig
kvtYgGcmJMrSBgZKuvUme5ZYBwDqk2M4EU+Jn+exSP8N4TeOhUrVGVO2AZtJ2qXQUrg7Po8CdSFP
CAar1emVaWeO+eJBmtkQc3TjhELhwT5Y4pZQdHl7YC4wbBrLCXKoPnfs0lBtq8cKVHZv2diVECVv
aERSzE4ckp3Jnjef43RTh3t/R3ociX7GbWzb70V9+4it29EsN3acN6ZJrSo+8worIs8DNTvkkPwu
KetdxAjxLmsOIGDIfZclnmWrL0CBhaAmljRGH4wXLwN0EoNiTLkDIecSk91U7RP7p+97+4GwWl4J
jEYz1etpBFzRowQEpP2ZUa8msoth+ZH5FDTC2zYp69PtH1Z1bVIynjpvzrTfTrOSW/ekJll6eaFU
EL8HMR9zsC9s1ecB/NKgS3ZlodF+Sb4REked9a+UqKanaoU+3FZurijvtZELPl6YarL5ahrtE8Zz
NDHPKy2V0q+wCiomun2eNbnm2Euha9SWGvAKnVTdBa4SnvQAC6A9FNSAdV4rbZeN6qnsBtPmgSE6
wdDB4n+ygDczuUv424gJO4YS3yTl/QgvtanMOoabCa8YkTxvtebhj5TMNHfwcM7UbT/TfuOm1ZpE
nnAIxN5Me8wnXiRxNhR+JLmziEL6z/zbh0GLHZt9eT4d8WyDXfO5e9o61qBG+Y5k3ulSnqq8q8V+
gy2BbrnBS4u+YYe2oz/ZQAbt2zjv2ZWxl1u6byI/DDypZuUzZ3ohlJwxH7DI2KdgSlsmieT0CHTX
SG7KV5eZWJkZvr67pQDi/nNrrhXzxO2RRem7rckEtp9q/Izr3jBoIzAcXIO6nKpBVN1DY+HIwt2Q
RT8MsqT9aydC9K374BlRoPKP0+rsKYVB+waJHOWH2UyKGKykkf39tU7URLZntHw7RKNlK4vKOt6s
t6RDqH6Iu2nKHH+XaGZQNK2HlC6U/N6G9ePdB/UieEifmX9puF8OMjbW3VBCAHXMzkuzcttwreof
vwKZyaQjOHzbeeaZKB+lG35ytsbHkj7vv7x8yO0oWjpRopF9Vw3ASuCtyLzKjmBPD3F1FtTIQ/ps
W3W92w54iwdsJZ13NwYs3ZiH8FTG1SjIVmw8m9FS6f/DeRVr+GCDApbqaYJ2+v/rHUAegw2Gnrmn
zTo0RPs2LhKZ39IYC+KYoOSpw9S/qzSBLl9myk+SzPxXhEvkQjX1YwPwxP4+gRUG/OlTf4EEJW+B
oyUdnuZnAh+prxmt4xrxa1DmL0Ed+P4IrHTgqWLgX5Se6Jk/+r4ZRcCiQLEDOtDW2Vp4ToG7C59d
sKraSc5ttrNldAzuq/UJcXqZy0LI00qnGgqZyXXyiCOfjPAmlvjgWj1cx6HrbreIby9eISER/opx
KnxxfsWAvgWKew2F4ZNm/ATYXmR6nELGEzX4xIQ3A4MLnzmpenQKMs5fVs1CNaqqvMU0z54B0UGS
+B7neG07xojV5G1OGrCXEghgUc+Xkvj6rxip5iJxQ0HNMseOYchIQiANhJ/d8RL0R3Df/OCin/Ay
JcXQn6lJgAkMhx9SK0/dhr/XgL5Aqq1LorpxU+oer7VhU8KNQc/FYZs9ZfunsP5eSKcYJVx5rqGI
PrJzTiSrRseIIEfaoOJVLxWmi5ivmMoNakppDKOdkhKGRhop8568gO5yxyUVtoINj2IQrzYSSose
lLAWgyuvTXAQCiHN0eXJrhjbGSxx/+SgMNmnCqTHfhZM8ZjsSopzaQzcHz7g/Db+TMoX8e2AeQBH
dcTHU0MRP4G1mndECpFWZYjj1ulT4YBkyrPw/IGJfTX8cX4kU61MIi5hdbcrmbSqbgkN49iiWfIp
bKpgsLQWzrqRomI6RO+zxdQlnSH24uLL2kJnAjUfsQ21EFvdBK49c7PVq0PU5El10jOjmYgvV6yG
CAT5rRl4P8/nWuV9DhmcxkLDwRRYr0rrCRPmCNkNq06lk6UOJuQah1+DnC4nQssLRN1MaDSD1jwO
JqNaJkZK+7xXhIwApDPduMH76boF70Lbk7OtuEK3rWSe4uMs4OEbH50cRs/O8uxniGUyeMmXAdyH
YrWvS5B+Nqcr7Inv/Ll53+QfRYbNTYnVf0TLtQpdIyeoyKvKXS8Kwp9aBQl2kPGulE2dix0Qk0u7
v0hkF4S8UMaDaUNfuvxcd8kc4Y0+6hrrYSuIkOMYOIlapkwMLlF2jMrqa2UpoGHrNTcCkO+iI8gF
gPIbYFqbRyqCecQUf5U3lzLO0BoYuKw/lDFvI7ShpCFLXzGtHueKBBsEIIUMOiUeA42H6eJ+9kcX
dhlUhrRdag6L5M1pLAkBYfqI/J6R0xlIfFnDod0+J9ig4OqjoYdpCnPsSjqfhUR0W1HSbHr7IJJA
Ycb8q4y38grTpFDTJFoJ1JLTXhR7tX6fH3aTJJcu5E+F8E46A9jDVx6rmyXjxU/Pg+I8zpE4cTt7
hCSKL+7IdgNGVUXxOKwOAix+G56N5uBL6W3/5y0AL0d8gTsX68RneHgVJDZVySmZAxCUtl1tyjQJ
QqED+j8GEH8vWRw9oDwv+M1QTj9+IilNB4Rk04HrCAp//kyy4UzLjmVSBOC6zSIf2u1NjtpFNfLg
bnUmJHELIENUW9m7zkn259+pyKiV3UbuZ4xSznMY0dULXesDCfb0FcOCJZEySbJICJVq528k5IdX
sVykgK4mT+13m7d9StAoVi/V3RW2V/IHeLGhZo2LCEEtNrMgjh0TiBDhlS/yK93Fj688wzlFD/va
7rBCVdPACkKx6FEcQtMTGzl1qkpNsIr8PEjxiZSHA3G54gei5w+AftaVLx+GALCOsxJKAuV5LHkM
gUWYCFgV9+R+rI2P1UKRqHsJLQgkj5e8SuKDYQT68VVm9cHiiZrbPA99/nNCDgi7LgAlCjBdi1MV
PcAQ99WKt1MmHYsVQsdNBDVghl8mmGJ+GafNU4mzHARd8q4zz7F5ZYdSiPfCCq3ozFlhf+7J5KHN
GjMP32B7QSQNu0WZE5Cxsx426UetrWGPBtzqjP2CM5Zgr+Ux0IPhnBDsbvICPiBBa0jbW7VnKZM3
RBRlYnQWeP1tzBF9q/NmKEJ1shTOYhUEHJj/+EEfpWF18IkhsJnM2BeA9PBZb0LZtXlME3ituXGR
5tKjB8fW50S2FRiml69H7jbmF2mFMmF2I+NossFotdTK1Cdc3ko4dY8bo42545174nYYG2DedbKD
ZPh5L6Toh15umkUMAJMGURkLLnRZBWhHpoG2TxueaOzQGaI+c7Fd/8eujNtS7gfOfgj3RvHi79uf
ITGpdn1AdHIKk1KePptcYSpggvOd/oOdOvTdV3L0sQWUqePmjwC4mQ494s6pPE2LAqAPdCZHTFRr
dqJ1Gl+XdL1qssxItmFPTGKBc2ATNeIrT3dtjcVpzTjO50+W3XBpbkm+xpL/6Rl/WAWVd0I/XyOs
hWA8xywg6cvPbH5o9bTu+BjJlcLNslwPAlH97RhQImUqffrzgLtspcmRDlnZ+rz576bhEQrnNgtf
r/LlSgAUett1+eEK+R8gKahZZxQUKlqiNUmNxfj9E6UbYJE6svwY3cRnS0eGrS/6YyGj7HjqN+XG
UGJW7dgOG1N1KDh3hSrQ9WJKLNlKhv44MXnNO2/Ah+TajgUQ3f/GFSrvuBxi+C6CPJ0A+vtbv2ZN
RoT1/Pqo3JpL8kvLkprXXUCv1e6LqM5GkERTydMsV6GCbTcZh4a2qiA7gqDusnWe+PY8NAhkXvHs
zXAIDPg3vaXiJbkGtG6U/zPcX2h5/lFdKKcw7kOguz0FxoX1VPkTGPPDoGJGMjhsLq7TTSj83rFv
KB6towQhmPOrCHJobMN7Dc0xpr32S79V/rRJfj/OfwIr5OKLRQD1eCdrHjKDIcarX7D2MdzEqneR
P1xds84hzmzZ6SLMzuj3digU9LbVzuKcPDsO4KVT1T+KKmS7u2NL9P4yiQMdO7wyQ2cbXxUZFbqh
mGm1s1/uupUmRfpfw7Xej9cft91j7V9NW9T156W2Tt0LhHUqjoXlBqySI+Zj/qS93ydoX9dq+Pcn
MJfD3M7b+583j9Gp5sJZJW+g+MpBvMDXYJhr8yaBkMuytuJjJ/zszr0Xk2Jh+e6e6QtGj9zUn9d1
jvZ9UdlO0ZGvGNSERVskao7Cu3G4CCTsn37GMb0eDxzWLHYh1lkSHAeoCebANK8pfoe0gt3lQihh
0CixyIf49IpBqm4y+HX9Gco1R256sUaklO1EKTPjyiXiz/eV7k6WyGgCtrIgea7HiG3yUl6SAnwW
vHfjD0SiLWStrJ1wwXkp3IJXoik2QSVMh06clVGKwkSVo5hn6ggOtAiw3SkbjkQYlvPit2t/1g3H
xK33Dl8puHcrb5feIJiDR8m1uDSEQVRQ6MWOoVVBLIhQbYbS94AtIfAAHaJLqqt76nxRRiuqstV8
eGf26bJpiKfoh+SHRwxuworWygb9uocWe6VY8YGWt/URB7pWOhVQJWhUwp25HsQQ3mtljMZdw+AN
/TI/vi/7aYCpgFEZ2gGgRKfdB8+4bzPNKK8BvP3F6qo7NROy9ncUvL/uhYKgzLBn1OcQSazT31to
AKLvye0ld7x4wN+VnuHTTn3XA8YnF6AZ6gplCtaI1ZK/Ds1B+qO+CAKSUq/OqJkKFxr0xcbgxDCJ
u5IkMqJ5/eyJXrH0FPYQa7WLQ1VHHqEd2GJvZCjsa3jHjc1O2r5vrthsXIujw2T5F9LigTLZO34q
5aV4PPyT3v6e393I9ub5MHFZamc619OGQ5LBFpJ9EnjqE7wbwbk65qi5QXa0mTZiXBeJklUrwdZU
1bDOT4s5W+HTDuOB39NCdxW1or5ZoHXBfElMTIWiL8lxgjSTLlEk8ml08qMq5hfB2NTYpzCQeOrX
9tOlrTGW7C0QwjdqCMwBk2gtW0cQpj3vCpKZeQncm4qpaO1NxQ+jpL557ix0hSFo/ltAZQJeMohP
UKUTxEX4Nja4ad+TiylKGRp+EHSxH/p+RT9ewSGlzdYFLOZS8OlZnTB1k6o4nsr2Ma+Aw1u9Mx5F
W6iD9AcuMx9V39V7BtSbrOT3n/WJwzBOnsWTlTh67e7NRHLXsvWgZgCfHpUYNdDwlm+MZ3zMQioX
H0MNJyXYR3l/Cu9FwVeRU1mwjFl9OaqIcV1TjVZVvByxbJkl5Rru76EpWnDibTMoqzjg3n36wCwW
OucPafhZV8MeIgaUGUVD6JiG01GbRZA+UVjYSH/6I9Aomeg3FpAnvr9MWryhX2iJJs6XiiF2/Yi4
ekfiP2K4X5c1N0RhTSismyzF/XXxrvuF0M6hhH3zuVscbXR+0AgNA76rcRoUPlhqruHkGyCZRbF4
f2cr95nv0F9ve89gUQGYR4I8I0mXM/r/sVYf4YvEwiB/p6max3V+Fs2sLblUvUNYPKvYkkZsS//b
gdSUHmhE6bOYTYHfZiLqnq/snWs0QIFQBZjEzbch0/ZRMUtNK08IqtJ8ETzb8PEwuidw97YUFjpg
fO4Vs6O66axK6dcMGa8DNTmXl1j1ollYWUDHeqD4NIPBjVKaj6UInY5TMHnnFDqd+DIskDaQ/IQW
t4F/Mej2ANTPGX2ZNJaBY7adoaOP2ILjpN0cRUm3+A7jjeIhA/5iWih372ylrdH+DCkK3/uZJgOu
jBgSOXbl9sSWoXl3VYwnVzQZ1f6Qhqtg9Fd8spZgqlUmqfLitwU32cLD5WY0UFIhlT8HnGJsYw9K
tV8ioWceQMJOQktpwX+C2NAeuuFh+8w3wBMx7TUKJqveH+OpKXDK0QOxBsVpjYDghK3uVBF4U7vR
v3jv5nYYKM2EslXtHqU3q6LrlTHyKBgUg+XZ3mwK7WHky70RjARnmK9Qp+XYyx1WTtArLQGNd13R
fgbXLHwkEDXhVMaESWMO9wfkn+S3nDJCDrCE9BzbWmCn/rUBw71nc2mqRAZtS6IaSQQ+idNbBD70
MclJzTdR/MuShltnXDLamKVMv1ZjDbWMwVvGdl7n4521vyvPCaDKB4IgR+8PmBEmWdQIg/lxLw/t
QQDfuS6g4kAnAo4Ww3s89AJ5qQP78bUDN1DVo8HC3/mfJC8ezQQ6U6cCg8KJDPTH74muarHSXh11
/LKVCd5ZOAh5m0nlhLvixZFOInP8mOuX6wrpKAf9r9GGYXGu9sRQRAyiFqRvphbNPqwb1uW/FDwZ
RTE1AC1opUYXL38hCVV9Z0tAgFU4+yDRU/5vC74iHFFu9eg3vtP7WwMp1rA6WOx3arHk60YAPe+V
oMDOSovYTo3FH4hNMIV0hZcGWQMNO1vMMFtw8fo4NkunAavuw0NYr3PORD3soX4FT25aQAfCVYh6
X8Bsj1C8EdRxDg18CSHSMOpTR4q7V2SL9kB1TJqIwnxiTIgLElYMLIPO/fC+eT7myh5sidwe3Ym3
zHetWX2wk66b0kFT6OnTTdMReXJG2RCSORSKe1hzQGi9nXi+KDBGyWoT/WtzOUtDgNy3Xzr7nT+S
oX6wR00W3L5sjVXr4lSnu5ReZPhfNGT1zGombOf1O262J5YUQJMuwzCPwyaK8N/e3VCX5fpkwh+X
CCfYqWhBnc5MjKTVSjWmxXxIb2sWDQ3cLMQ3D4J+BMd+wCkf9dj0Qs4LRAkY/e+yfHz42WBCq5Gb
sREX+e66Db5qc2QeCxaLjVHFxgDRhFzsHHVgYrq7fBF3SoOFfq2Lf9ln0Lpj+v+NCRC1jWZ+ASu8
XX1tmsdiQtAHNnKeI/rzNtphT80VHgcifB90FiUJYDdg1Xu03YwGWixsK4WpLJohz0FltmFJ8VWk
M13Enkt1BT0YG9sQPCeqMPEkvMOSJQ6Uo3oN67UDEXkmAPvxjlSbT8ztOhEUUETUQlD/Sx5kHUSL
h81uejxcUT59YBNphVzvCJu6fl2xR8qw3l/cDjgclW2ir1FQ0rRsldGbHABNRaV+yVXMyGyEDIZb
9GzRmhBMDNg2cwCP+eN9Ce2JoW3wny9f+WWgKZMbtjmGlJ4apQzRRWSFK91kc7x1XDSX2v9AEzzm
EGPYbDN9+1WvUAllW1jsGktRijgbE9LgK9550K4ZtbIqr1qwkSNp+phMA3ZwbOKH2Rp+S8Bgehht
JjGfVeZj413u6wlaUV+gLhNhRWNiD6Ek+Lym7t9eHqD79qY/9EhkpZG+pv+Z/0oX2TcQXois3zfp
DQgy1l0ugwTG29Wg0kTHFVz4MERD/ACs2akts/o8GDLf3/CZX7JuQhSP9lUaiOAcyaiOW7HDSljd
qleUEyxHpXAj4tJy4NQ7hLFTtyj2jKDyACHFX7BiZOFDSoeeOEtext4LozEVPvbYFLoWgdukKi2+
OpNwbH7rKaSfdLSOjOJ8px0TCmuM8AgmEDU8KSnpMBm5azPiS/XYg5DpCGGkJMDE7+3jM99ZIsll
wm40jfcAcZ2rscDKUNgkK0rkn5Buo6Sk2KWLXslWm9KregpQWeQ9E1RNjQ21Va8MXQoV0sorsXmP
Qy6LAIY0tNo0P+HGLCC056S/OZxHozJS+rE1lNjKtO+vzQiuJfr1Fax738XnS0uE5U8QC1RjH2O4
2/ORG1j2jylfO5wuJRZHK+LY8jasqW0BodWm4yZnDtGltrIK+cggz6YZbvOEOCsbzWrAJyCg2/gb
4orbPby01dd6wmem01N8JeuIK0aSWLerFZsBYespeOJLV+A4SrWMlqLbhzeswQyYIW/J2jePApZ1
lspjXyidi2ZDBwJbwttTZ+OF2IUA9OBNPhZA0djFtAxcp/bqonHgCuq2+4UEzvnugcwwjcbU/M2s
upHbkEaQ+nO6qUdmRivEFfg/t93wz5383+dMzyzLSw6e1JFW0M0P6J4w+zFcOmuxMsNbUEQYlfRQ
vt7vZTYMnY78PyZfdhyLDhlPcT5AEP+5m6pfQ4Ugv+XRAdvt+Xq2M9MSBOfdne+hCsS6NaWZf1rS
11+B2NuKlZKE9Kz1Wke+FMglpYj2Au1EPVsh3783tjEzf6h1J0YIzKkbUsPWHv7LT+sNExbNR8e+
e3Uf1Zyf3FAp5a0Pt//XQA6NDv3pTAvRw0Tzegrdi6BIr/95lzO0BufjRtKWN4FMSenJyOvqYNXe
+4xYXST17Ciarne/Dv8j/6ojlF2VDtFlUpSM3fJEvRVvR+vJiLuDpTJjgOGQnNBVZoezCKYfiYD3
lKie44jeWg/wzOxcC3fKyQjbbC3ksCRIM6zP6HBJV+FPXnWeK1lc1Q/3MCkyNEMOEr4wfHdiTuFJ
BuHn52dSO8n2WMnRyRWxYFOnslWF+sDTTTe8chlV85H6HpMR93ixeSbr/NJGbDnLQhcJ29sDJb6g
XHfM7FmMKiOJs0ZbglVUL2TtiAtW7YvNf8tqNp6E0GIEHTtFoPv9FgktVfBgomFroTi8d0YD++Am
IKmQdL56wa0Hktmv8QI7XK36NY06xUhKOuTibMGThmx+UCnXYCRDlVVoaeAlQp643z46GXJZjcfK
k8LnpRseUA/INx861jWp0FLKMoh/gRhfKkLMUdZdZtt/7CWveg5SweoRzecw6EV9TIkaSbvfY4lD
GCMLKXW9fVZ54qNrnCk8AmkvOkbPXFySDvFRcRd41hlyfta9NrKTobZLFk+Ayd5yA3tgJrh8RJMT
EKJsgtQRJinMSSnx+CI4HAsyfUJZVqokD9SPh+GM5UQ0X2esouIS6rM1drLm4y6yXF6Iqg8lL/Yt
H6ii57OcfPQiu+loTEt92VSg4eYRDCHGg+xbSNef97wMpyEdW2dNCLanbKze5YhjiGh8IhuXGBKD
ni+9iAWNBbHw+FAgPacxczKZb7WdKfBOBxDLCGHYi2uFymp4m4SQiBeW5yB5NLjvY1cIDoX8ft7x
LxCMoofPxVH9HFWaWnsr8G+J+DPz/ON5odDmex4bfbNVLpvyXc1yHIdvkFQO72oGYSoIcfuiZKZ2
Qd1n43wfqNgJsPngJGx9DdPa70+Oop4I0ifr87BRFXvaLwIonyr00mTWfyD9K+CKRXAQaK5ydFfq
dpdZTa+mygFx5dEKCP8kuVKmkUw92Fidxtltdiz9V6tbGZsxMUUIBsy8Dpe5kQpofx7Tk6MI9fML
wbbUVuQcGoMVMZEWRkhCnyWW7PG5Ctic17j3XSfQB65lAyx14TEkwXvgzNvyYDTxH2ezKejG2tKZ
NTFwM4iMs1UZnWIhIpfnTHNf/4fq0SoAsvWPGEo//IAIeWKO2qi2bCw4pwfVDFkSiA2A6zCi+Fxx
q4wk9Zl2XuUc63ybA7OpZq/QhdU5fPVybR/p0jQgq4Ua4hixsRtx92e54nrw5nIc1UWIMkjnGDML
1mes9cr8fAwSjBHxv2Cjma/klZJH/UxdPoPFJ+rq+4DiwV6BY6/C/Eij7vB047IbWf6B13x/2CQt
JapfJzjKbUw3+s+76+YvdpIUslrudJLMZ9XuIl656OGzhNEw2spHKoT1T8I2wLGghe3Ja6YIDA6q
VdM+noegPIxIpuIlDQjJcq4Nm/rfWg+b2UGxu3yGUfjtnMKRsC5PPwEwnH/T/+ncIuRzsFv22VaO
ItezUL3pCppN6G6LvC5F/Ljz4qde+fe7W1y5Ox8gSsG9WBha8efz41H0mBqKqbD4BKdz59ccA3D5
xRc9HfuymPKGuJBc9++YCmwj7FjwvUw90GQvqWu6BAcsVkz/nDBa3w5hH759c2285W3ncMg3uk0p
Igkk1PWN3MLlN/sCAh05Wpw2lxUWVbenFvB+NpoAOxHogmsRKd0Vc/L8IhWn0LvyqyUeM8NhNRpa
wSkZzTHRh+VPSm1HtNqJLJOL3ABlxVH/UUMP8Aw5Qremk9wQQLQQMhwge02M9FN33VUBI381jSMX
lACf/CtHn718BCF/R1hbPg2QQEAiu7ZKPAcmN2a+xuK27URf/tXoG7IElW+HYRo7KCi625LZfQuI
oJKJANB9P9Ph0aDTtQ02SSnKO1AAhUP3sdYRW3aQotNQYsI+24Sn5DLV+VPQONau+4wqR6ZMW+Uf
XbV/KiVSxaIhZNx1JyLiz1yrXwYjf8PMJhy2IG7bkX9mYSe74MYWUyvgFFcK1hJeYHhRy3Qmxg35
gVeWEyaH8iAUUX4pu36R6FMA6XXQiz1OfdA2xLr+oDmS05F8bW9kujCAJy/T+19uIp0ypqotXsOl
WvhphGC2v25IczRMRPjZIbMGSax/CoXr1Z2Al9o3cIdI/NwnDTDXKVueC7dW8D/xPjAG3yIVIU55
bGEWBdwvLk3EUEMvBAL+6xY5OkFH5ZxMFUFr0k7Nko8w4lKKnq0CQrnyiPmtBI1qemgTF1QDgzPM
VkPnt98bAh/YFgxKE1PNmCr4I0moFn1SL49firp9IFIqFJuaz2Ivi5RYhv33F2G5mhW6C7xe098q
BPDNhBHHQkR8VuBQX007Ue+S/pAPszn0ydMzwWS9+4QVBQPiZnl7k/ijoSlImxfy/31nHEAGm9MK
2Qm+CRfuv2QtctEWD6kwhrFFL2LjA3jiqqK8HmfWSRbj8RNh8LnhcFmSTNdT1yvPUU59EUWj4tBP
jUIj9A2/raKeBe7yiFnViC7qUGAui0cWhUyeCkiX5mpBGBqOkg/udP9Bxp7q6E1A+ljLIJ/5OU6d
sEOIZUJPLmiWzRNLRYsMn8zQlIbPzxYaZYMtO8ArgKh/20CgEch0BhASH1YnzPbeXDMeVlw4znFm
TTfxB4lh14LyeDnzPO9Z1tQWvYU6beF+E+5PSU23OoWQxMHsG/9C8ZKw4OP3GV6sqvjaKeKSyxXO
aXJ79F6dkMn1QiF5dlumWlfsJCYsKtACcOsrqXBOk+kdqrd6Xub6ymjo9rMZ2veTlEV5x1QOt9UF
9d0eNZrqOTvVr3GYiKUD5pO8uSMAI+KopCoIHWHCaaJN2ObGT2HfWiInWn9EIMBYy0QPeRiaqJmB
MjZa2Iv2DbtU+UQZT6XUNUKco/+rJlTs98wcgoLb55o+L+WSsJGrN2C1fb8ISezHapITycKMETtS
y2NxddLXMEr3nZjqwQdKGXSRIA1ldsKzfMjYXo08DPHvINq2y0ciAEh/FHqWqK0R/mkNvlu7WAvM
AZm3aEFZo5RKEvsBoRfF2ufHpBE0Lyab9LPEAM2SNHheHAcSY+3WrHNq6ifF3u+uyswGxkUKGGhK
4ftjCA0L0EoPqw0+1e433R8zqsObbcpCWtmhO57wyCbShnrssnOpne8uHisiynalRmeaWfAVvsPz
nk+LLihSuADAVn4GOjF2fEtvDJ3OyeyeUSdvpeXE4C3C6bbcJbKroCbmr2ixeFmJS8IHq3toW8bG
Gt4Hb0XM8kWHWBfp1C+ISCq8km5LONHpRQkQprGDiEZIhFMGjEktUycCmZ6yKUvQa3MUCkCq8rgG
S2ntTN/rggnFGltwU6ERxaJEAe+NLHvpry9aRdytx9uAyH/KN1uuT642FI1+2gg1oSJxHv03o9Lw
wUth3G0H8cuAU6IMczQoucHkZKfMmVj2mEchBHeVej8pxmfjZOWTYAO84qxFH8DhJsAsPVeXT9vT
ti9Lx11N9yPB5BDxXM1zhL0KtJpa2rtli0Gz225bjYlQOIMSUm//ZrlrQwdbXgCOY6J8Ksc6P9Op
/MRV5o6mzImY4J9dkcsnd6XYfrw/QethugzuSnWczRs7jFYKCQ1cJSvzYf9gem4+ndilRO93+FmW
AXxyaAN1Eb4qH2S5pu/NfHKuwENqkIBmWLanOF5GDzdmw9mE9fRDspeaTa6I0DYpjGCZkfwTfi+7
q582RWaTphNfuzxe6tU7PFMBfm2yscNcY+hYB5XsuGRhxsSkH4itR0tycxgSpOBMjf80WcIC3sr8
KakGUA7oyD+jKLJDME+8b+u6zfW4P8uKFe5fuInyDCiG92iZ1jZNoDEuxcGm2BEDBWdVc3WNMhYE
ShOOFmUgodbl84+pVrhfLFselEsWK5qbAoTJI1fuO/AurT8rHod2zr4xEOi2JOy19xBlCec3kgCk
JDzKx0//PmGDUr7hP0p7xDpvkMXi/IpLU0QTFem9eQhVSVyhVsqI1FGDDqDAcIMxuKL7xQeW4/bK
FTjyC4vmVIYafs1iRDlVP8edMlMQdsj4MrZudGu5iIqFuDMq7dfkVBuSPuJcwZXJnI7arBLcKEmM
RL+Mq+eEFtG/xb0ieFlvwuDsMySrsLeNgF91uycXQOfqDi+fLJDsOTvJQe4lcAYrZNl5GcOC58nB
5FswUyDdN6oexAxZ7TziHWlk/FBeccqvUMLZGX2uab7zTfscFq/0ByCJzN6wObGhO0EYBlLBZWiU
a349AnYn+/2MD5xHuZRWw/nUXpUftT7Rbp9syzrn4NqFx6EdTp2wiv+AWg2ZBsJ4P+CO4wNlGwHZ
FYnuDq36u9OM8Gy6O1ovS3zgSWUtg6VdpwYnLTkwXADd1M8UNS//5qmVZYXGDlwu8OZnT3oCGqDQ
RT1gP5ePGg6K41GiUhIlknNOqjk3nLJUVfoBOWJcWKq+6VXTwhLiEmf0ZGqK1ar6DauoiCiUjcyN
o/OXEWjS16DD943Y788AAzEv4sbS6coOcx+fG0oYNZaL+xSxWORo8sWlcoLlc1Uqg6kxfc661d9i
d+RjDrEMMRo+5u5PkYnxApD1dQ4M6YiEnXlsw3CaZUffhWBKRBm+yjBgvcZW7u4s6hV6PA9UUfba
EdNgGnHK6KybAfi7gJA+xufdEZSE6uDhhg7bX3RNZkoclaj+R5x8pog/cOb6gVt8WoiCmMY0Xjj8
+OUnLeA47mDTJT/puVxe67+/C2MIL66ToW9tEg/AKC7aKldUyCzJUgRqoI+JF46NJVqjB0RaYzub
fC0rkcESVIIemwWZorc3lEXrxyWEilSF0ygw2+OlMYS3HMLVeb8ojedsei1YvGm3EYOZtWgKSYOu
rKQczW1KYaVhSUEdOsvgALJnou7Qb2kZhgDq6M9A/wTxORNQ9sC0Z1avKcQ0uWW8qX1XEYqjWunl
CWBcXjXFx5+L/kFrwKo5d1lw98anahSDsnHAtqdGiCgby1chIbb5nhAUcc5R3GcfyUpMm6hhE+cH
xH3tIZh02INM8ph4+DLtBYgxA72XWDWzK8TKNtD3M5EC+HmLbG1AZ6Q84mTli+kQLODXuyVo8Zfg
9e2NNGXAwTVioF0edEXe7d595K7tfaocSpZ0zuyOLeT4xSwVD9iYOLMZ6VsLouJWUZfNrtVNUq9G
ZE6wgn0AqBtWef0rfIK7NYg5X0JSADFX8qk053QUnYht6rTyiComlNXqNC5IuBZN9wAg+62/z/0y
4Dmvw4muPkC8CBbJZs3YedJ+IQzSmlZB95I8o6YUmyJNCpnBNHADvjok4xTS+xi4QuTFY+98sxt8
8rVgpxm8BKknWClLY1ikhAtnDk/brbwF9risbJGnAHAapu2yOsF35ps/r3bjrbxqJwUAnAlw0cTE
tLVDKzSG1QUzvT28xCZ7RdGNl42btuWu4RdxtvZ0T1n3IWKJot/XRYkZP5DY9TeUiYhsoFkmBrtD
kA7XTP69zH2wQQBfxg6raMXSh65HTgDacT6zx3ZCcnkjc/fZgzmUsP7Zgr5j7JY5+zGe4mDq1JeF
P+4rBtFI8QvquffdeFkVf2jWwjcsN+oVFAExTrxp6xvnAQLIxp8VXZF3hxLZ2B+GX+eg6mWyfKyP
3X0AAAuxVjYq+2NBhWt1h8M+X6pA/Ma1ZVJuyuhLgBM5upqgfwfk8h3Q2AvoakrPjVphdyojgQQD
tWN3CQV8TJMQEXdhGXCqSTnpIsLYwryH7mF4DUDvbkskKZClZJdARhiPwP4fQni4Q/fa8WndHaKK
cgJiIVwMGKQb3rYyNddry1cc2S9C78/kWyktE5EnqT7Fi75RHP/IuMPMYx6u1LIAFjYma2QjESqk
cCgiXv7hVgTd0MCKXdxxtvzMWrh5+4ji0xfQmb91gAcbAK2JA+0TPSOvaxwZtrQtVZMKYP0NkvM/
Sla+HrcVpnbFv+Tag7va0cHSfM6kpOur7FzLIxl/phNzb/Eka9xL7lAYybC+VYyNNS8vSZ4GZv3V
mB2fZh8KGwbHFHMKd/Qb2EV6Bvq/uS2SZAuYti1QAZx0ZgJ/n8VZqLrUP34bpllwVMKLKxxJUvEM
+3nabs6VePJMVqoK/j0sCc9d8N4I57G6KEcPH88EpVAgIJEwgeAvnOdM9FPLJEeh1sMZ0NWvNN16
jcX9cftwWGlfb0udT5W2KjQf+VZnaIlTq3iuuvIqCeUW2YNBroxbJUdrQS1EmpC1jy5j7VhqL4iM
Eh9dBXnd0p1YZz2+v5f29Tr7JsB60uiQL0ej/uR4GGTx0RT6duQkXQMb3f4mEwu3qvQtxgRevT8I
ZkZqU+G6EInLHBvD9XCLVpPiGSmE4fOkHSOCbgC6mGTI/YZBUOuc5tblAaz7avpgFZZ6x5Gu06cy
NYhtIf99CE48JK1BkNlk6d1jHZBT+DNhKuSV6Fs/ISwVIyFy/UwHLQVZR5oIy/L4NQiF2ff4vrC5
jUUMHL/RfOQf0O34mBo70NfJOgAv8eDyxjmD9RGdnGryKC16WeyDOnyFlmyeOKvCDpCgM8gv/uGa
CFlH8dXO0X0xXHn5lc71V2WxB/OBj/OrMLtCUkMqv5cf/0/I8Nn1tzXk5GfZwIldvLfA4oVJcaOr
u4BVxruTXByAPZghcauUsVRxVILJL4Ve7B+x5mUy2rC64/sww6bto8ROoXglQL1dA/5oiQotPuXF
xTjLoOjeoihgAPhYKagI+79ll9pgjD8lVeRtve/eOm7PAN/XYpsKZDdQCb/JtnxrbMQuazkmc+WN
FuK4u04FZHqvRvXugtjmBjbERzqv5dt544oHU77ci1+uaXB4q0SYWTNlsetBlp5yCt/KptAHnMzf
GR8nIgqAWetQYiwNlKuH8USlaL/jsdk0potzJDJVfUUvfSHvnWVqYGdTdC4AY6H51TA+heOOoH9C
v0FeGg/DMGV7dIbOCjquyrzgIaWxRDhSljqdUc0v0RP9Z/76Fn07F2Is+p5UX9XgG1hhWFFhoNEv
/kB1XewlT72RhS6T2kULLNse2UOsTX96VOEsy83bB9dzKLjicLY/+Wb060mP0OwLNyajmiDaz2i1
HAUM8YTR86EFGroRXaTLKGEBAODwcvsqeo77sZ44Nqu6Pw1d1iMxDsiGfHwJTldwUieDHMNuUv/s
cNel0S8z10YcjhYXsRvlGSk/3zU9feBordicsGIOwRapQB69RfBYUyVvHtfnFxe89lSSdQV7xU+X
xMeBiJ3ErxD9liTb6fyM2CKNys0mxMY/70I/aSDypZ6XYvhgGk3g5xh9+7SO1K4czIq+jbWSKh5f
mNEzo/Af7NOg5wz9EMJF8NhCQ2Ekz446+5S4pvpk32cxQ1EG5nhoKvFZxs4uVE/EDMvtBt1uShKQ
3IYTus1MwhMccjx0nS/necg/mdvNLhii+iYPW43MksGxZANy/rd7SNoQzFHh9S6QZB19gVwtR8w7
qIC1dEXl/z1SD8cfi7LpZeyu/4bIGWYaPX+YdRLjedxN2/CzwOnMaAPZXxthMATTScV2X4G9C2hm
00NqSFQJNtRh6ng3vdR6XWZSczmrVlSPjZUU9GxyK454AlcLb3wJWUAmfdVewvkJtD21mLC7CbO5
XX+RXAdlCpkq0RnBbqF3IXSbUsNRI0PC/Y4UL9hbTZpXa+9cIqTPAKBX375TaRTyCXfAPoTNL1VR
tvZePdLUP7P9q2cJJahRNN3qgYS5gd3s3MkU77gjKEEtRce4eDrZe/NXP1Bhsw/vxAcqSV0mbs+S
cJxI0dGpNnO1rj0uxsSa8EGwKFCmt1+tBGggr7GSF3UX7cw5OxIpOUnsyuX+GlcaMwLhfCPuJn7j
QFECQtwiEj1JpR7ckGFLr5jMrmbJYTJE1xQaUxw7SFTPbr2qldH4AX+fNXqQmiBCxPe4UAw5nKgW
KZWJgItYoY3uGXn4G2+pNfus3E+mSXSzNziA2AOnD+CsONL1N/Ok0CecMGLeja3cwen8f0DRbOrC
aifKuENFfbt0IoHH/NBYuJzdH2x/Fc2YG1EfgktuKvSs8NxKIQRsmt0KJPksuAYCtLXacoeFVTzN
5tvK4dOHvAxKYjZJqdlymaGwT8BuhUIJxRrNggmrWIBzc0S2eIFGAPGFMOsL7kbxeeMmRikFmKsw
S0K/vAT+8F7xUWkA7Z3Njgwxohe1LhA/0QmPFe4mky89aBEttg/Uow6VFDUktPnTMiOkv32ONndt
k+XoMwrY9vz+EfmDm0uNWNtmaoqa6pkpRyziw/7ZXNoY411jxWttZvv2EqvhXjHtlgpSGBXFKphI
mnBsvHUSg0zW9Bo8zAihHRoBXhJDRr1u4hH2gvg45Q23BVInFdrRemHaxwYcCfvo5deX3QJuHVaD
Xhx4KPRvMSg5xEgvCh8hNuAuKT9BMKLQYRkLPgKTVI3l3DIMwA6oWTz5DVe8kAJTziL0r8tQ1Tr4
c+TrSVsxhxHK32Q5oRcfQQbviZITXDefu9SmLfvhWtapihphsQcWuC144MaSI1xGkw+4iArxiLvE
UUVi+fB4lpH2EvsY7xSv5/XM953OEKUmFkl9glyliyC8vYfM0b1V4h5HE/lXRKE4xp2Tyqb+r+RP
fBzmf0WhuDO5rwHP8VGJ2RszOtKWgn5ETKuPiaMfK9Kbdn62mZVQ5pOpIQlTToq55HqcWo+1WAl4
0ixjfxS1BW58C2lO0gtlAmBfBxyhGnNmCM3eKwSAh/MwMOemjx8dPsyGX4f+uPChpj3FCC3HiLSl
ju8HjKxpiKDHcYaL1XvcA24XSmtZcC7Syc3cNA6yXv7Lkh4AWtM8cJhwMFW4pZ/4ppxYOSgrh+fc
Y9vCgLJ7lVAoR2HTnfAe4ykAy6g1wHYTdexhrVbtCWzj48xweTq5QFLUzo7/FMgtt2eICLoF2Bu7
nVrxrumCdsn3vajLD5emxSW2f3UdZcTnnxJjJZc4GyIbLa9la67HtZfyJqcUNS2YN9DXPV0BhFNF
wRTfCqsNf3kDDANpxt7EiUp3yX21MpSjXffTXlYJuD58Qs/An2YRM9PtS13uNLFPH98hzpZ+/64Q
4mgyMsfDFIiGbX0v3SfQ/m41Q1Dbbl89ybSW3AZSonJ+tX+KdsFEtpDTqTj2/ofWmqaQQcX9Bb/a
MbBYfPOAHI54mTeZxWj8EmbaBJ8jbTLCUfRA5LFw2BBsfjB4eQ9KZQxlqQTBFCbc4+7M7G+G8jPn
6ukVCO2IbVUkT5snvdwUsqSzboDynQ4f6RkfI6DoN3MVNOBrSgfhwurlveSdl1ruGjY4+T0fhrTc
VI5fv5kbmIR15pKFD6dG6csS2AgTf5O6b13I3n4O+b5arMGXwzcH/7p2nEKkrPi2ebfG+GmTfwkH
84/EpKfB9kQUv7ohUluqU7VgwOWPNUzEWYdx4HRL2Fe/W0h8Xss5mkx2XGXu6rwEyr2oBoSQEdlp
XA6YsLRRUEADLJPgVNXIUjTdGvzSQ5bL+WlFmv3wXxXhdiiZPojuPg5WFCKS101x1GqoqN/xWqoT
LwB+et0LG4wb1cAXshEosEX+qjMXDlxbsRus3pZVv2SI6V7Y4g2rvx/tQ5MOsP+r2qMH51rsgKzD
/HR5fDq86Xt/pOjJJor4dK3XiASu/l77wV9BwMXRI9rqFkekpJTSKrD4XuG+yIAnzr83WqL3teDj
Ig3cVffEow8XeK7bHQaKUTXe9wWfFY4tnB8G58GoW5aTedqYcvRbXSChw8dKz3+roR2jlfP559WH
Yd0PuavEhHTy5DmBT6+suHnDFqhKQRBMNWLD6ao1waJgSm3uMkad35KonqfNjw0nL456lZ6lWED5
oXl8E3ZjDSTtANbeNGXJHgG26zHnNT90daNJjJrWytm0uP5IojusgN1SaPoLKr5DCJqcdCkUCnE0
/ZcHMjEj6Gqe/037gLNUguzJe10lXY9oSV4N1VIocuKkZ+SJ4w6ndja9chqTqUtz0f8B2LzuTXBK
xc+TEe4AjshsfDX7OQKNiAaR6RAEpoLCS2UhY1pCC4BEQtvkv7Zsn2fVacH/T9ApbE1U8GC/Eb9Y
f8V+GhBq+0ZSlMoG50i51OYOt9wLoNJZkYzEDuHa4rhWwFHX/Lrdp3617Z6434pKs9pJFX5qTBD7
onqNmWlTS9arZnPLh4xtDutfZk9r8xTMC5MuXSk2gLojnKB8JbTCX3ehVtZD43V/+mAf6nIisL1x
srQHSUw1pWfVFjL4uQS/Ofp/IxRYlxMRbsVM6vrKqfaNdO5EsGgEh3vm81dIqRaztOs28LfVtzp4
/Xa+ahMrmhLs8d/lki8oDkKnGtq3++nFeTTSvVGWoBBJxrrCjVylqfkM3hi9ky14rXEX+5pzGYO9
qTEHllc5+IBsLpRP8A+GgPbfaQ/A5IVICAh5DQSmRpmvyl8A26a+kqrJXI8YjH+JYAwnEzBSVFbc
RRuWhV9CQlXwcGqPwDj0TBc63UG0KrtVVIk0rKZyBQwJPjZC4HUEmEwCU+wTBO/SpEmRXLXPMvIj
t3OQz8ICoL087DIPM4MZliGUDHpvpvxAmrs8IId0e5zLfJUaTdl2uVRWnBxlOeZ33VcdlQ33YZeX
oPojdRG8ySimOmwLluAsQcMlX3aArLAZXcUe7dibwTKqHITIg7/uyQ2kiffUKQx6poM4IRgJWWLM
shp75VjiOR8qdCQsIOh3J4+X/5F9hErmCrQBRVcbqJiW9beGFMd+sF10sGzZIA4fzV7WIMZ/Cfvz
dVyg0EMbH0qBp7bXEnMu7J1xHWKQZBNqOQcsPgAgHbQE97PHOZJOHw+xLb9Truh9jZoT4qV/LO90
yA8dpLaa8cbswqKJxeUqOnHaJBigWaLvN92gFc6hFx6LWRqOMMhFvcwJa/fuyAQiOxwlyVAOAyTP
mGNg0DTCocM6VrJ2hkhguukT2dt+87gxNW6D2XAOpDqXnR7ORP7Rz3A+taS6vrP82BvvbICEmzud
clo0BuHoezx0CgzxGa+93xHR8MjtMsEsuXFHIrp+EgnFJPeu8TN8gwV1a5m8O1Nf45ef7YgKIZCV
6SFAeIjF7tlCSSVZZtunUwJDrw1mzMFoVnBvZ8UBpD1uDdM06ihGMcaRi1RLCxHW8gE3F2aaA3nr
MOdv+jbgwfBjFPABC31lnORlF90TZWwAbNu9dD4bjLrnU+ifHeHXWLuX2qlE5AixZLO19l7fA98s
gJnsSGjVHi2/FV+wSBZuCuu0lWAoQbJih3B+GuIjL5fUE7effd1piUr8iivyXXRj7WXqW54dPuMA
HMUX9mk69a7uQoQ7Y56+6fcDRHEsCc1nn1KpoC610LZZED6YzP3eS3D3GS+lDOElYYwRVFD3oMQD
d78VkmwjILEEDil737BuIbZZW7Nviq0cy4o7po8wbI14+OuS+xhhpOd/xxRfXACIRQT2XB6dT72P
dunG5NgW5iz96T3KeyG7Gv8mA9oMZpIWx0zv9R46IJZPUwsb0m1NXYY6OsIFfJqUGurA3tsemAo1
Y5rnlDb20IFJtwfNWVDK/L/btU5lJhpkC4ghGoDPmJltR/DEUxKQq6SeSptoASHBfKTk+ceVaVCO
SRIQyynGVtlVSy4k3dMwzH6K/AAet7zI/U453NLtNQVZyiM9NwWliSdfPCu76iXwiWwQ91KOUV2M
JS6IgsirZhDphV6IBkVArHVcqeTaPQq7nVECVruV8wJKoT/a3hC2Lv2g/sWWnwCtn+rAiRNeGy08
Aj73j9xrVGRX0BmPiEEv18X8+xDS9dntVOlVUzvPyAID+RbNf5hCCSeQg3w26DCdwomZjfuL/eKM
lwXzBpXVq4spVTrzCC+J24uYRIzOEvJl6dXdClXFQN5d2+OOCQtpIRd8wL0cQCKyGjczMizaBPPh
3PgTZyHej7jYyZXzZx0PcFG19LczDqszpFmuXtjk/75fWpyDzBdP5s4EIUdufDdTTh9daor7LCBk
CwNW047o5W7ozLcGdECmioQhIIIiAVJQTQERlzb2Zh6qjxrqPXQraTCw+oDL9SrS2Rtb5R0Iouhs
e85IDbw0QiWChNhLM3eIByylLLOvAtayOevDDoh3rZIlBwSd8d9KTrYJSsJwfd4P+bRa9XpDVSB+
+uF+FF5MJq4GcnX6po3BSERJRLxhOy3ndEuh9/2B9pxmuhiD1aqrSCkko5NEehI1twvx0909VwYZ
uTjIlLLWYJ9i+3FCL6TG4BBN1HzigEOASAP7x5vVG4VHZnBB/DDjlpXcSYGrCyOSZxt/RPVjzw2s
TmU2QRdSfsKK6j6fjpGnwJXhj3DIXJLEzuQB/+VcT2VOY9yq04P3rSEkz9npshGOIutkGIWq+6it
Slk/RF1NF5rPTD6whnlP8ZULTIK+HL8ebOdyM8xcocLoNnKqF+OKr0m8B3Hf0n7scPwLwqGB33cN
bOctdAX6YrcYrgBy15/efO+RF4tetE8ZbP5xv6y407fLWPbnNuouNRHw/ZejxDD40yVOcpq/4Vof
/fcnLL13MWwq7ImSpwLXtBw4Qe8YEs7C/hgKUUZ5tb4bUfayy4oT6O4UfaeJ2650zU99pDjx3Sr5
2M/O6FVeheX9cDgn/RfXSjfog/uYwM9HOHB4N8V5CgubqSXlu/3QDpUccX8YiLfyyvKNxziLPWiJ
ppoYWaTMqfoL3d6q/OZ+Iw48DL3k9dCIwI6YO5Dcig0HQcttEcA7UhY9rNwZY7W/tYRygtCwcOFP
RR6UG7TpD9l25FlPQWVa+gYJZ4uRDq+ACPWxwxK7NWFrhNbBtfW9Fo4K2aEIbItHVQd0c7XFxB+L
J5eODGp/p7Qfs5pYL11Hm/I5jIfXZGYRRkkO9jed+6tk4Xv67IvyO+oGmMN8rjCqNmX87DL7D4Rx
eP/kxZPwj8WTGK6t34R9yqdTqkVlJ39WOqBqeD9Wq8w5MzZXA1zSTz4rZKqE3kMLZwh54s85dHoK
xwy+ERDbl098fQAX9l6x0Wkz/IMMIwVJs3RxHQ9BlhVuwIuRgNhYa1dh48YBCILmOUdJ4+VggHsn
eFWtaYsn7CBb64r45JdA10eblnvPtthkxFN612l5QzZ/3fN4Vps4dShTfDjq/l29xh3nt9cblT4i
PWv0X76IFsu8/0HoIvaZoYBP7t1507gUcr/DBkRMQ0jYBijmKcPIU6MnjdZlU5hTvlEx51KRcqnv
QhunOpsrEhjZBsbrpoJH6YZ8Tg59uEJKFEPJENUuFNc1ZJlJgJC74GUvmySo+UVOlR0sJa94sArv
uPsvVBKyfe4GxQw+DQEr6c87Ndp11ZOs94Qg1oz9X42BU8x09LEl9khr6+tFOO7UWsMapuwvFTzj
0e1aDaJI1cPz+XFWScvapEtcRT0k6CSDhisbjFdN74Ty7Gufhae5rQRnR+iiBWqwLYWcic1Zjmj4
f19x3+oF+OEbcOWkQpytazYLcvNexxvTGoRfNizPVS3acBjNLrkkKXcdtqtq2I4MqLUcP92R/HH2
y67axJZ8rQQugi7n8ennLJCfbuxrnAKQRunnboNKhnXMa4h1LLvLN4chn76N78crEY5ZBtZSvzYV
DScRBnO5pS7ZYnvMDaANTFe2gy7vWkTX/7OvOu+xfu4lX7B9Zixnes+cF9A9bhDAI5O5xLS2LaPZ
EXwXJ3M7yNRsIs4vIG7J01x3oMSeNx1T3ypyvDqRcYqihbaXD82SUcRlyywjqSKu5XcTnbuSWEPg
6Gf0lbaXD0z/0A1zzWBbYpSuqEMA+B/Gxr6dgTHlP68g+A1vsJtOFTXQ8TCRCifl7RtnQIxe0tnj
kwy7lW7vWvqVdy4l7TkjA7vJWGs+ZAH0PFDxBx5+mWK19BeaXgFXMXqWrfvcqEQuhlezsj6bnm1Q
0T1zFQbX5Qr7Ahg6F/7r01llCqNd2uWTB5UHPNB5N7z9UxNgV213ImysFCUENgK5rvd0xK6eVDyb
cC6Er9yoFcHcq2UXwn4kRXuyCtrjzNkbRTP4Y3R7gLkMmqku8sL7AO0J1muXWz9LxuYkrCIKx0Ea
2mtYRfSAq6WQravzkn7rfUhllfjiSkU0tPhnujO5Fcm4lRUuwjPlzTF6DFgDIXUk0Hs09XpclXfe
0Rx/iExX0gw/eLlNxGZCZbP5fO+h6zgTWV5Ei/5bUEgs69ZEOcoo+7Rxp/oUosqewyGiZadJb24n
NE3Adr/tpc0Ilr+vu2Lj8+jqZZbIaxDXSiIYAoGSpixlQBBc7HL3N/bfTbuz9EsQdkQ6bpnsD960
wc9kLbrUZEtz26+2sC/rluXpWPuOA8ALxc2AiPtD9ogoA5LBxVfDZqQgop9WN4XM92ZFOh+dy624
shBKLPGNZjRdqrCajqVuvykq3C9afDWf8CWDeqfVITYFfuq1fVWBGOUGuzVpjUlACLNhI7mAAJmG
cHP9zxW7zvbfucRjKW9ly4B8V6TrXwTmcpcH2agnIvTEMR5HKfPXv9+YA+hWBLUlblIScqTg/uM6
xP81o4f2IFGy69AYr7MLpEyzhAnzkmYoB95TCQvOHBeT4+R65s0XBeoSy+wHitscRFPrld2RNJSN
c7/4qDLavNO1CH3sqUOKuKAJnCL9RAWYpnqX/QQ3Bhf6+Wb5x1OjGy1iFpKZqZ8g0NZyzYDtPTUg
SWdyAyOVxraVHUkQgeD6OC8JeSCzUXcmBvaGLciR0j2LrkaLbWLEbnJ8dif6qgic0b/qIHmTR0P1
T+BsDu5Xdch+Hn6cX3kZs5OQ10dGB8GnkY092D8GsmqA4U8kflpgZGjjWu/NkpQra2gNd649SLRd
hK57Df7q5HoCtmuou3u0QhntB4z3l34ZQNzfmhGVBvTPoblL5SO/FSxF7gKGxE4N8RmBdP2A8BNQ
RCI2vdGMM/uGNdc2bLbJ6Dw3rULW6ZHx7agKaviANzE4oUeyi2/bmkMHKqC7rCZTj2wtxZdwT7R6
M2YoK7SXch0JTjFkHmiwSMxc1U1uX6feTXz4XijHhW4uSw4dGnztVTMD6Unpdg7Tg5KTV0ns8v/U
8On0xdl5qTYGaAZ2Z5sHCVnpHjasIpgYkmpMH6JLpXDpyQEinW8L39RA3uCp/0Oo7Bce0eyaexRD
6zFFqnXzOKT+EBccCnospDfgMcwiV7NZgsNPL445I2qtEoHMXuXEF1D6SHP88j4H4ixcfO5h3w8d
maA+Yn6rIN9ICPcGjStexs/sJbCsoAfdR+q82pxAMoX/gSWg4nKY1rg9iGDiNSXNwaIEvYKW3+6W
k6lN3w/6QeAarQRG5gIAOTC8rOvKnwQ3/2eUvhz0VU5cBVM6Ng0ASnejmuRfMKZr9GThnU5u9rrk
zcaY+8bF3yRnS1x5yA4EIpzzRkwhY9s23WF228dbvmzavvux6dds5qktJCAhS20tFPs9B39Wm+S0
m4f6ClbhDDZplrrcVSJMFS3Y3/mn4GKkQ7S3keTkl48PosPsMWlVFbkDBo95wgrXaM5hRO2MzV8J
97kb+S0sbiBnJL4Gp2xIwuxM2S10D/5yPTDzxqUCP2A388x/po86s97hVk0dzFLUdlcW8BM4jH1V
olUhAA3kXZcPdVDhr3PMIOd42cFbnqm3iphI06CTBtHDsc/yYEtgVJEeq9JwhsT+6v5B+Q+YXpmL
Dz96X/mp6YKWd6c0aOxs8mxPw4B2GjKTeTDm1qolBbZFUoYv97n4erc3ZmwFZHsGiauJrsNkDKvp
wnJeBX1P/OIucxf3J57VvLZ3Z9m29B7Q1SB7Vd0J194SCdc9FZupiux1EnTUaxN/BDgYE+nDXqRv
bwWC8cmMhAZnk7hGRM4Y3SQL7Oy4XbsOfqs9z9MnUTWJVDKAp9uVZMrW1YmknNAqZ+bYAXP70v50
tY1CtlrlDPIFl1VsEv7LcfVmiuFa73cS2wNDqZRigOV8Iv4iqHxbl9nKmGsWjmLXmWgJBH7Y4B2Q
PDK8YZOFz/sBiWiw9+3TGXt30wSIFUUv6huX38S1eCSVOGZ5upVIdIlKZLMXR62mHM2K8wu5oASD
v6dGEn0ALfC6cKcxgcYjLREJgeDPMK7MLVnG7m3hnZoke+ePiRLYkWwhNVOTnW7iG68XrfSiqJmp
qAyOeTfgZVxZZqw44Grsh2Qm9mqjLiT0/k4/YAV03xSod+G+YYD1vv/OizeOxtAazNwht/Rhlp9k
atwqO3yrgHRgJDLlGzkGUZTuwQs+KQaO6CyT0mwVuJcTMMLa5f5IweXoGAvfZLd1nRLUqXP4jTYP
OHLGlFZseY7DfccnQFQEdq4HlhtGWRgBDd4x4u4nJHyhoTebB45u6h6oybPAPomqni844tarSH2U
Di4fsdPAQJk4CatnCrOJdGt+ojjD6yJGnCwZYHS5Qphj0ojP4RyLP6LzQQyHu51bygbFjHktguJT
0sRwbNL+968E+AcEnH3G5XGk9uMWYSBVzRuVRNSbnkNX6mL8sE8CrbG3TGopVPWF7CwqjadY7egi
V019vhAMnaRB4clQhENpdqZytap+8dkDtBuuKeuY2jAm0VLjZj+2yLxorvUhQL5r7Upmo4wHO56P
QNngeKSwFpK0dY1IWuR7D0ajbXrhkvZRGF8AIgRsmDDtu3QW4AKi0qfz493KZu4hdbOgdj/Ee/9x
/cBElw7FXBwWG5jNrE4tHM/0Hitc5KhKLsaBeqyu4m1lS9wx9/pnH1U7lvI9cJYsNsHzaaAAA3kG
7dzmHZjYlb3RmPf3Zddhitshy8KWB4ST78eUqxxiJCCbWnPqZdPnvQxZzTWRE4S0DPwqCGint4ID
BXa3ZvKFLJOLUeSWmlqKf8HQY5a4nkQR0aPCJMNMoczqM85Z5/MSx9j7iOWReDOp7ZBDCMFVV9MK
PngonPwBxwBBTN8Z3dvlks8GhmH4yi4nLsNtw2iyDlwS0hFTE7chrDKjvMRKIrErzvAw2bGl0gZT
gbvM13npqnjEssd8PpDEta2/sIWrZghaJaXRtbZo9uaKh44z3oPq3xV1ckl6XGmceIytySSxfb48
cApimiR9f4/J5a8gkMhFCNOHN3Tqr7UYAAvcVJngRPng/GWmvdCMPTavagLCo+nbC+QLoiyMaB36
6Rn15C9ZVlxeudOKgl1my4zsciv+d17a8wsL65W8OzT+1ypHAJqzuv6piWUbMR/iWQlc1pw502La
4rE0QQRTca2o1hRlB5OQO1h31jKXdRu7CuM55B8aJNrckymXs1WhS6l1RY1a5Q3MxG0EFdaKtQz4
qdS8eqzvHshBlTwSc24l68j9kI4d0o7jyvJD521IclUynC0L17fOhYGq1K5gLMDYiMOkGX37t35I
Vxi79ZsL9ccSNXyHs6KY3Sidabl1o7/jho6RnN78i4K13TmcpjHZ2ZAXDYBUbvddYc/O8cZqk8VI
8UfsEHt919vFKu/cIjn12ISa6xUELzZinyecuOhmQAzcuEmbag3aWjsdCpzGDsD9n1mLQdyBtmBo
0+TswXeVf3Zq/pHimXEqyS6KudXkzuTrPOP9EFW9aEsEaH+OsNl66UhjSHwpKy5ad9ahXMruBTHg
pzRxS5/nnm2QmVsGrLDZu0RovsEpnIxJgNT2V9hKrSuRXb569z7ik9KNO+R+jgP1A9kaBWG/cGvh
nSPLHkU4J7NIvXWCMadf+WvFM+xr6zuN/YCO7GEdLQIfapWEaMPZaVSkXCaUtIBAesDgyTEl13Ft
UcvjMK0258EHQ57p4VdMYb1MFEKDLCxC0lKNWTsuAUCRyXKqcuUHEqcDdTlPkg3+7dNbc63c3+H/
J0bow8NaPW1SyC2D/bk+9Hf4QupwkRZycQZlrVRl0av2rQaQNtp5OzP77Ir08n2dkXfU3svsISEt
yU8B/S4t6MgVwZIPkWMq/N5EztdAe0bXymtMNfZXL9FHPP/Ij64+QxU+eyBBd2Px4WEejsT+ojRS
LOCbYk3PwDKI0IOZwiOJEYaII5m9yx1Pf2dbow0S9Z9J8m2qIO8IZqY6aWrzA6JzBBKXl0SNm7kJ
+xnGppSgEXyr47CoY2vmigmwoTXDcULrZmYyJj7FF33TH96OFJv4FyCC625Xjc2XuvEOJqr5eSSu
L7nEg7TR9SnHwpa6HFfIYZqiT9d9Pe8JeaLbQUs0/q/OJShUGlqnVGI0EHD2HQdYg9xupr4e/kzG
78quV1ErF81kjw+Z/FF76IIXveZA5VRUPEPf2rhvXzVDVl0gQMYQIW0Z6iqZnV1QtKsb9iOEV7Q2
Ub81KzoldchFlTuanHzE0tJKg+fHW+Kksh9Z7JDnrqBBd9rHsPmSvSM67pHLHBBec12VP/aYtafn
XLmBkNLLOq9pn9laGm9ciU5FcNCy9gGpd1l4S3A/xul/pzkpYjlJyCAj+sLymsvWcQUV+2OIo5Cl
SVLCF6qmajiaJ3VQFpRoFtjaEjlcpuMCeKVAUlzNb7dLAK7XOt+Q62zui396BB9FKprH5yiFlO7z
99mROLYup9qHrBv7eOlXTzDSq1pSOfZiu4y4o/hKHYRQuza70PjVpp820Rl/E5y/bjQIxgDI5S/g
xSY0MACkFw1Y6AFGsDaPNKNBdQrt+6dj68iZsjLTGAtivHXwpHb9AnaDs7SYcLK9/k389Hj4OLDL
8ipuazcHwAQCVCpYgyE+6PhhmWqQKnk0sc8/ZvcLGqVWzxJDOU4xgmngFwlDdHcHf5TZgkDyuXct
byNHaaV1Ip0gqoue1OpjSQl6xEQFW4/MbBHndE60BXyXtmaIYwt44Eei4NLkVUejPfUvWHmKTO9p
uwj8MMv8QmAKGj45Bw2Y6d9Wgoj9If0Am4Cq4GKKopv+zik24iRJ5+p23mxU+/DyyZVKVsJ8ePu9
toSYllcEsZqm4kCZKyGC1D35fWwfoYghONcWJa6w207mVZtMUJvtHF8DHsjH8i22/6UhJt1rvmfa
60Vs1TFOyOBxsJlYqXx+FSaWRvlsxfjOzrhmlhSAiAGLe/x/Qj93/0SqMDiwPykUMGHpmUO+/w1J
8Y3Eh5GMYNxU+PRHjcRtlXo5jjWhL9GYxO37KmyGvTknyfdcOelkTk7hM+Qx58RhYwQKXfBiitCL
cjlR8+xcrDc/yVpm8r7u/lBff5VLuQZl23p4H41II9LaL6NfThSdfLtrlcF+b0ESE2xd7aB7ChQI
uKHi82tjja9gdztLiLTiGdLaPstwT6jqTf1VDgXwYnsG435LZ4wP/lsg6SAP5ccc3NKBi5vZj9OF
FaQ7CHZpTrO7dJwAU3GW20BiGO6pdTa0rry537TvXuNmDy4bUMktV+XIcUgWW0kdcAN7RtOk5FYl
Cwj27KxJw4DZeiLx9Vc4jxR/q5g97GcyF00v1zLoVMMO+ui8QHZdexQecEBg+PLc/AIkCgyg2IMu
JA0b+T5KRcB85szqyCLJs2v2d612RMVhN2b8x/O0d6OtPguO2ji9G6HpS7wJheiEBL45rNYPUDOd
F8B0WVdA3j1MOA5Xkd8irb7TkcZnpm6hchp4ad6pv+Gzr032Ht4dRY3c9R8/xucqNOHctxMvMjls
Uw9FriUnAbt0DmkM6eaEpqxpUnrtX6T+p6jwEorNlXx8ZOf+Two+qVyMuRdjVEo9k+9GaouapNXW
HQe4nDmGIPidrtpQxdjsKNVz1yY+ksL73T3Jo9k5Up6X7TMr5zNocCyKuchg6MHl0IYCClNHGl4Q
56QwJIg6VIMigl39GLQUDXvDheBpIViIHcOIGZ28zi6D/btN9w64gprKWfp1/azoeeCIIIay2lxs
VXJz+dOcg21pZ6On+WEMvvE9gNVt+5AjQ2/3XrUhABNTEwC/Tv5UGB+nYiU/E18iY9eOv5Vg4Hl4
YYDssGkor1oEnE5hIwJFOQcbjAfvrVIHyQZBnoMNlZ/7kQP5gLDPp0+QyPHK8ecCUevFiGckv4RA
XASj+OyJ/fUTDyLs9wQZN41RZix4/1KRxYrLS0MiXYguIeC5x26ucWorVxv2WMaXtzWjz5JvcL8s
uZGhgnDWtrwCHlp7rjA2xkQhhIz7bUJATWUGovGhX5zTf8zZwJehXEHk9lFEWbTMtRpfRkG8IYNn
rR8WY0kUI2+VUT5wyE7KIM9LkIPRk01m/tXbR5T41zqrOMsMZ4HBz/cdt6n1n1eI8Q/yLJpb24lO
9RY/X5JyorT3r9MDzMvcIKIGwJhpYaIGutJ76EejYZsqxjxnUXpCtnUZyECIAQgWMWZHPdZpBFPd
2Ix12emHEoKu37gvAMTMrDMz29+C9q8QaSCrrzrwLH17hFvhHCdF8i4OEfXc+dkgEHt5azaYDN2u
QsuY4LpqmLdLjtdLdYeNu2YwC7W1BIZm0F/KEOCSzNcMG/XYmr8RxqKxKBjGj++KpXxYH86pc88H
S4YKIdTmSrzbiGQy/X+SIKuMIcpvamhxFb0vomTYWTkFT60HCdG/bOWKqNMtLsHk7IgiBKK6IfJZ
Rby8iEIxrQCbibvxS3+cIUXaJezZ+iX8lk+5X6H+iTPBdHwL5zn0FYTr3RS8ui+47JVuufuEfg4O
kQ58ILDEJTtqJ6PqEx/7sO0v74T8HMWIp+Fn4d0H16bcg3JE3Dc59vXYudikqMBJAXqaIJXERui2
pAF49+5HLO2PZ2z2rHbYdttz1/+sZTER9A6i95LK4AsALqyAQE8Bl7qU1L0JTAnVjS5xhIYPEQ6F
GNBuJrzJ6+Ih6a+Dyg5dJKNvjdszngYmT/1H3uZHba8ywf7j0zzGJFwDPQh8+dn7V/nJvizkr1Mq
7U3eo3vkpoY1YlmAB/mFuLKC9x4mm1866YXWZn2Y5tLBJuPQ6EsbXi7EVWEsXkmXDBlGit4G8dhB
3PTqmjbim5pMcc5P9byF/LERrHYtjiIKzcnW7bYgJf93iXpOPVj3chX0cltCg96FCpdr4zEv6saw
337Wkd3oq9R50p5L06stJvXcZ2Y+Rqe2LxlthSbV7Y8tbIlnPn1Lh2vNyNmkv/6XYR6HZ8UN0xI8
9mnpWpbXHFMVVH/L3nzGL2NvSRnKQqKLukdpSkUAC+PZMeko/0KXI5sns9ewL3IVfBVGb/aTScTQ
qbYVqaKeZiR34QPx6MHLo0ke7VQAOVQ0EWRsuUnnvG7y6XD8Aq9j3tUkmH0bOIXdrx0hr8rfSSU6
H3SWIiaREIK1ulOAeDCnIjrfWZxUyU6Nv/t/07O5EfgLwVeR0uJ/aNIAEKnpBuLRld+AKTJ7KuDy
SQ09Ov1loSVkHtaxORXip+cp5izx1Cx8jlzrDwIyJvMN6F0dOGUNkM9ECCXlgytZs3ZRdIEzDgt3
w31JT8qn2uQVKjwzgQryGcgbejRM9aK/HXQASZg17e5L0bYQ4Xfjl0krlPRya3nvSzZDhmSFxlWh
A5/QvHw3WuVKsDFQSHZ22I2hq1QqGGhRAHKwdah81ChL5pjiTx2C3dJGBx2LOUj3Jmre2XjJfMq4
ZrHTwwn9EiuvorQT9Bb4V1gqI0PXxxn3/dygvpMY3vhgb/vVWZdYpHJtvcTyRrRfcWwB/20sCZVN
nbCym/axoCqOBdilVWL8xp+j7i5D6oEu7wk7Tg1gnJd+ZhFSBM4Asrz6ST3Gc8VpcsE7E86PfImJ
ii2zhYPqn4Z17k757luVUbpbfS7e/DIgCOya6Kuiac4PlJMz7NB0GitCXwKvcRnrY1y6U9UFqpJA
u7j9sHfILN0jdIAaQYiM6mrTc0V2Io3FbOXcTX9V+CytU5JZrsPGjgvym06r/2oAv+tR6S9nOkL0
Pdr9O3R3LHhtnKXmg3HmeO/IG1HrWtk6Tn1wp1yaXjFSWXV9wTa0IlsUvuBCof9uukJSVFpxNe9N
PAS4/OuJnLgpqk3hXKZC8ycoiMT9GJ/4lhTjw4YjWo+d9V1VkET+vxv0IK/JUTo1orWVA3D4rKJI
rY/dkUgB4F4kiYT4M25jhRxhrA80H03IddNR1CknUIOaTzaR9Kt/jZeSIPpPAnUhucgfZzulMEs4
0LDPm/jx48TSBy7u5MMAjFsjJd1maLhW7P6fyMIRONjCTJjbTu9QRZxcbZvRPRp9ZOA8PZ+Q9nDZ
LDiN4084ElHSbCBri7LmULexs9tumoQ8pHYFkUtCXt2HSvtDDgJQVBcbGb/ANMBoxq7zRFUFU1Mj
soZzDGdz4JhZBU/+SZfdiI6nI5nIRErLkwV4Z2juxytFGyLNAjwtO4sUtpuqBorVCu7ier1DnzSZ
CvwN04gBt5M4J8b0XUjgIuF/2P3xBQRfY+ENIKa/TnovJt4d+HAbWKyORlsF4w2Y82FRMf68Qlbl
SwJyT+cBy/ZATrs3KMwG1jpE+i6jgpAbXhZuQjGh2vilzYEs+47Q6glg5QqiThfiZDXUF/pyVMCd
y3miSqHfXurZjO6mhMyP7x+4jU/zSNJdCAZIezmwagtfDI0g7wQVcvYCRYkAaPLcWAZk4o1zMS2n
/XVPF4WfUUU9B01rxkk3bzX4jwzf9qg1kO8+ApApNg9Wdzp95a3kkGPr5DVEF7PHHeMk+D/i8nQY
4eCRSz0i1A6AL8o874j1XP85fKyuWHmN+ouNjseYAuKzRXWKbd0sY1AXGPfGK9eGwaIO/IiiNWMq
wdZH2xMSG7oBVzjJ7/+NsFH1BBlwcvLGa/M3L9mXoHyJIYxxDXgJSheDotHcJ+2/SAcMmtnlzIlo
6yfFtLGKuM2XMQ5gKVikb8/pyE4G2iXS9teGwd7pvs/9v3lKngYEb2BoLfAF7jaRiImFO5MpGrW+
E3yhqU1ikcNev1pPWxJOinaSDMTvCxVzblB8RoqrCW2NnixBhs/rzTSIMXnb2HCltNT6616zAWUi
HPjPgBU0xlNNU3DdYzBcBiA6YGPyeBo/K5Uh3e0reQTPYxDrawGbSGv+Os/Wg3z9hD4fpWXs3e5t
CVtuCVOyrOHcE6+feTV37Af1TBZ8b893QKmB1K0c274C2ruKLAxzds84bl6CAKAWeuYjfZguBmTx
8pKdPXywrxeFcalaOh5mf7+XrdyoPFi9j6B2VP/yJl7CMEpPkCyLTmolkXUlw1QPqouYPIQ2oLFQ
4iUQOMnhVv+1kva2lqxKcUtZh31QT6BD7fyWZ7PoFJ+Nx2SjA6wuCLhkhOTQuzjcoPxSwRwecfyK
Vb+4TqWx4yGVY7XWJpVNHaOsD7Lp4LPZyTmURmnLQsX4cbWp1/NHR9vEs5A/UA78pP1lf7QAWi0L
yXO6NzlYDQIfcpO3vVPt3oUilS6aDX9x5QBNNIhXDxlNucdW+Y766Dm5oJLvxwFvpdBHVFDTmQJy
t73EbmdRuNqMHoHuUJwh2fWGsdPJfwRZJuBV6F5uxDFIP5yOozM8c/8Ix61mgVn8Lbpzx+c/YzOK
ufzUrXsbUY3JhnExv8LZNTDJZa9AVsWJGlpxiAqgq5s3ESSIDdNR6wiQyySLeFOSSdrIYaSHfm5X
bv/wR6IGC5mxALZfLcqtxhwyJsHeYq+zE0qkzzgNppB8ww0MeWY6sLHEWhIqcawIupzabtlHVLeg
lQLPu3uzEZ5/rSrKAMm9KfwmJHWKnOGpj6XlqeQzbXO60k+ha97wq8TFFgRpGL0VzCMvAuARbSE6
tn+ErP/nEJmWwyNuJkUvqpd51l4PSHwxCoDMdv4NfTSyTiRECA0hLk9aA7UQIwEjo0C9ub8efVsZ
xkm5kHNS/FTypOsnUxc1hz8CQy+xPsKOt1C1K9rJ1AOUIkJWEzh3Y+r+f/lRV9oEwMc6SNYIjo+J
5Bgiu/9lE3DgQ09voOoOEbkVesZ7/W2OHXrtK+L61WDbbCmDYbFRyfnah4tcti1LMxGIh4NwN2A9
Xz/6vHwEvm4cU8x3pyKdP8Hw4n8/JhTWPnmm2dGBzDmGR0/7H3Dz1QFX3+taLRbheBnVeC9UJaHW
JHMTeb7/mSb0SaSJDk3KvfozUdCFm5i7HlwdgKwmlSoJQs7ZEcowPLe0RxA//Q0HrRYKAVGuTu3h
mHdYmoiWns8ig4XISRhUqeRJ7XfXlT42QzWvlrssxz7v13RBKL5m7VIoLBOEAwSfwEYvC1vkc/DZ
kb9JguN5K8pW72tqfFrFDtJiQB4LH9/ukd2Tu0bKTtCSlTYRU6taoywvjfmce3facvV2MtO9+boX
Ba038efTlTOEP23pmmRbCU0Ke0PlBDgQe6vbVsx2ppQ9tYnpA6xTgXBUBuW4OFVjV2AIpJ18TOqM
q1AG47fBZJLdgrPD8qJBC0rVA6c4hBgf8CAdN1MNGiWcwvA9mSwyE5VSxrPayZgZOpN/Ap9ZoI21
C/pq2D5OXzY+BNkoCtQwH7ODWaA3GwVYqapjFs4VFeCzYcZaI0x6wDnJ3e6BPxS+5n3xvkCPrIFc
nuvGIJGjkUu5mzcH0gOegon5LIpz2c9t0enM4nn+dDglMpzhS/hg0MNzFwASmiDEbDGGEHraT7Z7
+ldjm48VpI3xS7Y96GeVGfYMSiH8slSyCGMJExZAuubBj6TfMrdVLnE6QZ7KCTpn8IM1Pp9+ZcYR
1LNSMT5Z5hBQpEHu4mjqQFbS38jyzmuXHK017y+GiwqMd8csxOnZqxkgLiBHPUzT28nxuebwTeV7
ONSZ3YposiHS1LgEa83iwTYYxIDztm4xhdMLHU4APNhAoLvDgbBL9gK3kNwyOOGOTmwZnyo9W4sF
Nos1csyQcp14gCBsQRppGrTC/sq4CHUJImh/GtrvrGxTaxxu+FktQpHxvQ6eOXBtHwqjERj6oKEd
C5Ollt7pG632Ps4snvXGCCFBYI5u55I5clcskj9Fd6pK0ZPmioI7kaanaZOSIcecfxiVM7hB9s4T
TKCgMFaVCUsYZzmCOwBt0pNov+D4XaNVGtJI0UN/fUusfd5GchhbFfmxz+1pWj0FO/d9qAaXmyLS
PMjNzM5KRD+CZ0Lv2spa8SSMCE09UsJ2Pxs/qR2kHUC5CAbvCxkuqHLJHDn75B0dL9XmdjnODL2/
aIAM/kS4LM66BCU+2fl4huklCTekuFN9QVF9ifoPzvGvCy5UQ3ighKSM5JT92hUY4ThFhwHhtR1n
hgk70RhcvNeZLxZlpVR+WXOz3NX685ddXKFxPrKyZBCM7EVAgehzDNCgujdtPOYzpUm3rPnwWjrr
7LaAVsRHlgmdUP1dP/4Kot7TfqN5voVUc5xh49kkz85QOPPfdBnQgXenDdO5kZ3gupmIoMXI3ulb
GZSkWbvWKqXzBInamvedPrvlNp0ylBldY0yTgMHrkdaTjbjVvVcNlGY7RV0+VuAEuEaLUx+BUPR4
+eIQzKuzwKAB9Yf20+kI25TAMkLF6nkyFij/1Hzb1UcCs30U8ti+tvGFk5LowQonByVEuAYQBDZm
/HRy1v7WYriEPd7c0P9kQj3nXklCbJwxkU0+dxBKGUEVSzuaoGpOagTRgH1zPWbXA9R0j+ysGOa4
socwYYWrrOz2dJ+wGGV8wgHwNO2ZrtSohqk2xXc9Kr/6mxEDZHxCn35ZFss8lW9fiFIrnZ3hOvnK
S99XJ+29JQjsozoXiPzT5Ey5EK1G4c4OrW9Z9bzBwVnLF5uuHFS6ju6SOYLpNfj26E3l5aXStksV
y3uacEt2B52JwD4sPRMIbcYSK2f0f1x+9pbfnwp3f1qytKvQg0oTTbD6yDWJSoeHsUFR65vcO360
cgZ+w/lRuwtHvrizkJQl01PMBWWPB7yCZCq7nwYCRn/Y+fMhQN23qxBusq+h4qtKDATJ98PYXsYm
3qbmZM6qg6/mPg5n6MVsKPETiIM21PEyOd6ZAxdMsL85Nu0eJM6ZDfg5p8WcJWI66nn1pjHqEZRa
rvAwFbqmdFVQavIEqGtpAiQQC4VwJ5BFFzzpp/NjgUGfN2oZAD35b/D5zlM1R7w9jihw73wE//x3
KgJOE+sFL/sDbYkicnBnn//+od2xyVV2ADzxqEChGnbN7/eY9TahbuMan/gx+BVLDardkMo6O3+j
AZ3O4w93GcXTw39UZFLcDHYMdCr1GYuvhqpmlC+nqImqd611ZVYpApIv7YW1n9WqXOuKS7syjs7F
jofWQzzsych18gM4i2xEyrEeH0FrvoLstWMbeYvGpNW0GTjJ7Z6A3TEyH2yWHTJ5kGAdd8D6T2Ub
oTccHjmJ9j4PKeQYVRhsvuGEflI7G7B05vDpShxbMD5vyVBRvGolHJ2EX+4iKMYwx+0wr/zkGaqM
3UDRRgiX/SKQZyQZ38EGMpNoP1NV8l/5kqAKpI90d3vbH7S1ODWDIdL/IwH0hW0dxz7Mcs3KO7ZD
xdtOyaRljlFGqzkBjazJ/f7nDUIm3TFXZAusAOoMfwCL3rIMspjpmqRvMXy2xHsRiK1Uv05bIuFh
nUBxqgJ5KjVsVrpTLEcGxzzwUdRaL1IUa5GzLx9P/GhPb8RhZJxCLwiNaL5tGaSVj7i7VfKmKaKo
uXVDbnu5NhK2zQfV/qchPSbllZuVklq/tWErpM9GSnmI3l/NxKA/QsUrlAXr+SPuzDroLwUMWdd+
+WgBdZX0+syjKE9+ZLSQbM1uJhXXKSqBm0+8XTBU1jA/NMSs7S0CUm1lIEp0rgpKn8NNdEEME3jc
ez4d/+JtelEz/DsHUIlRpoH/RNGKZCEHkr7nmk+AHtVWpnVwEs/qeou+Dgllq2nkqGcK65zyVEpr
jJd2UJ2qJNhDPHp1iIh5KmfQ+gO0y9T9UaYcLNFpxHfrnC7M7HI/dJ0fPYzGJoDxNU9dDBmJuur3
Y1K3Dqvt2tTwYGjDTYx5EjykJKrKbF4gxsmxf+LJjrhq6kxc+nNZC1dwq9QQeo09mhuQlfYS+9ib
FwLQ7VAW6kBOyUEgvYHoG6BMRDzo7Y1JEyOR83ZyLn1yC0+WU2BY+O/QbEz0U7BVFB+zvAqkUDmp
H0A2KYYE/AwpoW/roxaPaLJ55NpYQ89xk1Bl2/UYCwa8Yqr4BEIR7Ojvs0/AsIbRBOcl+dYqoygn
Fbt6Ke1byO36VpsC9qaapn2gzariURexIvlPe+xTBVrP5hvrNAwEFcCi63k8UZSK59wNG43tgzIs
cr/aXCF4s38whZ3jEahhXmQXQ1OfuGj2HTORPrtI9Xs7ag4Lwh+HwIZZUl1ZNh9JLnPPr5Gg/OEb
S8Ug/iJ7u6DQVy85Cb0Z0AiVhAyBhjjFCGq3aT6SvWfyPHnBaS3/QRhDmTXwytp888DlBZapzz7r
w7GDgJqsGru/AUA+nq08uS+5IRwXwHZQLz2iagXil0JVm9+70whZs5cD4k0kxuIU759Qav13w6WZ
mMdaydHbpO/QEJu/vrIf3MFjaMQeXEv/bt5XEHGHET9eO7pEYKKpyW8RuDtMJvEcSr3iiw060gof
WB0AInjEL1Vl8o/vGDs9BZidAcoSKWPj3Gi4V13+PkwuSCCCuOatnY5Vj3vlUxmuZcxV5uL2JWBm
qMZAqmp/DV/vJoUaQtZ2iCjy4SIQrEFtvK8B27gkPRTdt49OVYngQFfgcDf+FeZplRXkpx5KjAFu
CIwXJKNeBcQFs3iwYsst6aSK/eLsfXuW46iayTedV27W8qn3r4OSYIwrYqLIQrD9rnMx427SEZC9
Q3hYIJz8XV0I0LUx/wx4QkJFHwDRtihi9jk8qO+YEGykL+S3Ky0fWXpbS3SKwK/l/UPhhnTIRjth
RUPMzDa6o+FEO08YGlMtr0ngOsnhBOKi69xLeU8tqJL+zk9eXht0AT19Mf7QzSgRjg10nnOLMLBp
THiwpepFj0CpXIiL5ddduR2WBOvtCzNfAE0Fk0ehwOi71UN9pOryp2L5gQ7umzpCw5hrI655XG3H
NE5DkZhi8EO0bXQAc686QScGVJ+prVUrLn2KScaSZwzSD9f+08Msv2WkfGPyxvhrerHyOR3inlyl
0B2KaTcPcksxGgMo0HaqiJrUMu1NcnXogSlxgkRZVEsch5AXuijgPPmDXvfHYx4AfIThnAqdXSBy
ixxfvfWYFQ7bPl/t99Igk31682Q+kBxRzr/59/wjTwdrWccgJJEvYewuQW7KQuMnuwiwMt9EQOO7
8PspWA86/kQT1ZvQ75Q91yFbs+hRpsFDFU5ski/1Bi+TjLErW0YekJA4AwO+GVqUW8ZFGlC0DFpP
Y+A6Rb/8or+ElYLDqh55ll+VUwuwf7SfSn+Rm7p9ImTRvzrylqMHUX/AT6XlNCUcV1SaMSar8h8v
jXE3zpdS5mU1LwyuHproCuGIfxP6OqRXbMmYuJCOuyjkOlzMXPu2M+gMk3x5xBEooMkSRBX+jZ0n
PPM6X2D68KZOCzAGxQj2zd9uVfIqEeSLRCwi2P3k9ziDYGzRpOMxWdgJwhVCmZsZPFyqY9yDRgaM
1rixJxjrWNWZofEwqFmyT6rN4r8klOFWmrwY2zPa6I8gKt8SJr3uwV5SmHcJHKoaBWHiCa7hEqzL
jKDwx8Mqx39JOI11Rs5yPL4yX7OMfTKmcmUDkyeqJpWIvY25hP2I2sr0L9VWiYRJa53XaEF8yZnV
nxTPbly+p9qctqeu0BCjhgZA7jcnlXCZauE1bHe01yMEJhjdD2aNVKJFu4uuKB+KHN6rvao+TYhE
12b7J/FPJIYT6qQ/7McpCMa9AE3LUYkrj+pbyRr4X87Up93fB3QhK7cHTQ6ua/EFH030VRP+x5+9
b2jOO4n4NXQfCINpzeJ8EA7Kyyu8ZB8pHZglcx+ux2kC8wYKgQsau6qyaHihYZgM3MG7SZKu2Fqm
2DJm/mykPpVjTg1VSLOH285UHGAB8bFn6pFxFz76OniHmjfWE4xWlBks+Juf0yxddRLnauVRwqe/
mIRVJAC3bGZCw+RiIFEozXujJIpFeAuwf9Pdew4gRb4QJoBxIyBEbxV3JzGyaRfOC72FFver8Q8M
tdlzSTdVPyyjcNX1lsgdZMb31vzSME3SiRNNebzl+lTGRunVW6fHYz9w5YELf2otiMvMFuY9OMl2
8cCVRt+hSdwGfy1f0Jk66lGlT2qtJGPDEpFIVW2eJR+ZXG1q3dB8hx0pGBw3dl29VZ963Dhyvprs
oFeXEChOUt8tJKsEP8/5fVTf6tJ/yH4XQ3Z71iDg6HR3IsU2TxV7UhpVKO2Jx9ay1zwUzS8tp2uI
Mtgmpo25RaOoPJrtGhPDRn8Eq0uAPu7h/iX4RpuQ5STmd7ULoFUGB6a0BncL+gstfA9D7tj0cvgu
GiWYZOMHKJ/o37bfgkwnftYtZMsM6Nb2DUnCZDgN4yi3RKhzDGjPNgddJykc5yh+CsGpgWDkJcHN
DTFQt9s/yhGijejqnKhktozE6/SnT1fehWfUPEGOYs9NkPJb/9LVVpsJZYMR/K5alKe8skf2f8cz
Lk+xHDi7xYY7YCjHvCm54ou278aPKgYK7DhKWv9M9qz2HCr1MvDQy/qzuw5EkFmeh+XWuhI43loz
OXyTrNySOvgTD390gq+nODv4OCIuEa3C1Q51LTMS+uLOhRbspsoMr/7Zo8yen/yRUoY+m8tZvKf3
/jOh4mVTxrufBj3MBihn2J7tSKMIXNgXBywfs95Tan8mqkbXn+mR7gexNPaIi1mF9S0Y4HkswNWG
XZjiX25TInQNPjT5rFNYEju5o4G5eOLQd4uyDTMSnb5N2O7rbhGvgKrq74MCdJzB8G63CclTpq2M
1+QwzvOmOvkjBWYIG+hibsIlxlF/BMw3Ic+hKJgHxy4r0P474N+ilziDUgV2xgfpNa/KmMVs1gk+
W/cj7uwKFuxtGy7DJUcxQxTzjOuoyElJKbeh4jfBW+avjdAax0sDmQ3DhJB9fVYGYtf3ewHFa6c9
DfT4HiM6K4bBTkjnpn6jIwui5dJ05Ziw//RoXKzjpZPpW1hAjeNalC8NSSmLeuAfXqbvRjghQGnG
9bqduXInuZADXc2yuWQpMwq+5NmsICN4HUvmGZSCbhjSGCDGNgBTiEZ0QWGYJaF62qzzvuMy5F3f
Vyp9DVnSadPrq5w+RNUIkPDXR1hiaEOF3ZjF65vFLCbF0Sgw5CGUnCnzZR07A0Ld352Ej1h77sF8
AlXnondCDnXxpEFGzAsuNSBHBQo8EXs0OODGKNPG+NcrH9J1dMODtT8zjUph4ZI3G/GBBbU0d8SU
ZuoeT6nUXH3FLqHaUAJu7c1LDhcrKUwIYaPQ70W86tzyGKMrPq9z2xYnXre+Ri2znuNDZq2tXAYf
mYu5AnLW1SQJ1UdGSObkg3YeJ39l0IaJLd956k8nXorVA2SDedQvIYtmV6XpjBn46AoRIMvcZLjc
TWRDU278/2Ikf4KsCTQJs8o8/AqfFuLKAQrMIz05nMqNsZ08bkxeRADzj6WTc3h6/az6u9hzqcEe
4AnJMMI0Z8BkZQ+n2jSmtdUbWX8DkXcK49gVuyZlxehmFgEEzRnvcJcWlqSgoREV31RCXGq8JOvh
O2j02JkNh6FIwxXPNLjR3eVASSBE7rf67p5XeywnZOmby2fK+Q66/tGMuw4pC4XtTxuVZBNuXOhi
YcGfRW1ByfLWwoWrvcl5p7GKNeXy1JJNRp4p2BkuS+XP1xeL5pizv/IHNvH2CEsqMps8SsUSVeYe
dg1MbO+qXwrM6uxYseyjVz52Mt3rdg7XpYbzva8MwlvSDRhgqghwSxFC8UJX9mMO5eE934Ae7kC4
lliWjHuUl1sSwhsBsgxVJo+ARSlCs+S2kctSAm6PzkxDkmIUdt5aHr8D2eK4keFhgOxqeKBT52ON
Lz/qYdrPtKPsbWvi/bUwE4hLzqZU9PPVGFuOY8CdhJPMQDHpMWUpBsMMF3SBwUsIZXQDg3TlVl9Y
9T5xo9KnXter1LP4B2oxBsjLv6+jGU2DBsK3h/In4uqROQqrmqnJQ0RoQytOcu/V+KPmEpDtwwkj
RBBVTPe7dLZjC8bYAPoqOTYYtqOxMCMu5nAABq+xUiCUa0dgBmmbbp4hXhVZjttjkUcI711x0lDG
+cwcTIPiMfMJGXGXF/XnRFzuFqoObck9YRuyN7xYpArPBfLiPhhAiYoBW9aMKVIofnLeMqyBLwNW
0NyAu+pUPz6ky7ctNM6u6Zivhzq/FkiT214DMzNEfHHp3yR6vdUrgeZ5CVjCmZcyZQ9CLwSxmPyO
RbPYWMIhs4ghb9aWVK0fO800f7v6kTpobqc58DRy0yoQnoseoYG8gJonaXlrscJFW4TI9dSwFTtK
MHNUhEKns+bhZnh02CgBWu/YsazYnoVIdJ7E7wK6Y7vyfeiAHbTyc5cufFFEn3lI1V+OS/A3f/ke
Cr2KENkf7RP8vlcFtumTyVqwj/4YmR3E4HEnPtzP93Nq37wDh5Y3tOFg6Pq0Dlybhw1PkMyTEvEf
/6HCSIEDDyRhrreZt3JtLemqqTzanf/s3K5g5UcKAwcgEUi13WpI5Y4C/sM/kHrtYjW59NgFct9O
82aljYGianGy83d3VbSWYaT/gl7OL2BtpprekRj5dYAhpZ/mop4Z/onNi1GXXCtOhxMbwAs2TPzq
e8S5ZrHI5uL7pM1Wupj0Knm56SWZ4oz9beOO9IrMYR0be44RrWe2IUY5zFFoX5E5qdDdg4LEbyhu
ZqV+Ni/d2Ce632RXbwNW3KkNHDzdypqeVvqecIwv/0FItvb5sJwQS9hQgeJCOxBCS7QUInrTOSav
oi1KtpTGZNrwSdl/mnZzLFxUTCZXQns4y1XQzefkrg6ogLr653wPEz4DQ4s258W+gu0siaRNNxzB
OciVmkJ+3zZXmG4uYqDIKUMHZmafP03aFF734InaeviJFVIbKZM0jxsAwTXlPmPj/NiiRJGxfAkW
ptJS+v0yCEoQKKwF3vlaVnlBlYmh3JfUSTEc9RE8IZ0XuVfO+95xq/AtLfRsbvlRPsuRaIAYaR3p
iNErRnvPNs5+JWH+vHTbN7yUxcpqIOCL8RQp8FdjkSqCHMQyOhoMgpQlXDnhAOMXpB7P+XudBCGH
ucdR43MUMvZ4k6mvg3PrPjBacDSoAjx4SuxnjD6VCKAYmuZa5QlpW0QxkLWrddxKWMqC6D5UGGcd
7thWvBu7CnmHFKncJT+AYBXOURBRVFTVw8xYMorS44oiS6sSWa0kGP8/QqcRyMvrSs0Bp8zZwDiu
Oj369+0dtdPtpCWNK6Vm3vrlQXN5z+RqHFhrXW+yX3PGIOdgzp1ImtmXkFULqC5th67cpjzVERF3
UKzaV4nmJSo7H6ye+dWJSDQdl/Rg3sonDbNnz0LkTOU9m2RdyCDI0qJ0nBqeKGMa/vGz02TiEo7T
NU6SlWrFhZsvK+5uAWUav/ua9guwXz/RMgbOaAE8egB8aUuUMPaCMxJalJf6W7LFT/XGQzskwzBY
35G71ZBPz+qtL75FUy3IxM1FnUN1C3S30dweZEwDWjVHu0TZQ6amBO2pn+5kHiaJ3L7bMwiODHb1
avi2wFpcYgolLpBoO92cKTgOZqISK6RLYNenLp6SgbP7lLXncuAzUi0BXKRjR/pYJLomkWpq+y5f
OOhNdgUKyPFVnkuKJHks/vDgvPgCQz/vyi5BvDY+pSQmFYwZuxMzNf5Bd1VH+/ZBWb4ei34af3pc
s8PDabaVKZFBi86L4/4d5FWNZcUFWL/GmHFqhnzPbr42Ae2pQoLOlkaPRLiInFdA6PLO0k8AFC88
aUlAkr2DT3kldr71gPRLNKJXnt46rl8PNG9o6q23pq771dSGrlvgkiumpODZ+RZRl8CZ/hJiP/W8
+wFLgfOglwno5hAMl12lWvph+JlCMq2KjHeX5+Mz4HIpOTFCDBzWzO8ZPu0e47cXHF2ysHxUZ+nm
aXs6uJ4UPaV3X9zKQd0vJrg2F8S6UzviD9MXFjgxPSY8GndIWrID9F4w6upkyyVR/LGemQrRZv7s
h0AgDLx5sb+MvMZUtALbSmdk3aqmR2vI4gepCc27OoxSZeLi9VeJMeIBe07MD5AhhJBrijCrv7ct
4aMvQOp/oK+MAaREWI5BFRlU8l4ZLxH9PdmmJNjJEFUpKy3za8pW2okH6GHTAL0gG9CuujdHslRp
n9XtNpD1a53S3SyWixx0GzxCb7+7QQNY5EZFRO7p3wRNVSZDVBgk+PKry0D9aogror+NbarPLf9W
noSA86kO8tLyyf2V8fZFJ5/VRZKfj077wNsxD+h67MyadhnpBqUmf20aQ4BzEJeb6hNZ5WPav7AO
ljWmgVo4FhKYzEQ/YrTtBj9lLACDmW2k3r5eSCaZbmNa+AH16tcwqY7Iw2Y6rK9bR3A/fREZjM+e
FPzVTFojib11F70i7F1tmrcmLeM2v9J26ViYrnxRheSdQCV7GPoqPdxwEAD3Dqud3Vu/RldZfhjE
e3aUuOeAWpU+ZCNYFbBQBahgYpKskO6mY/yWY4EdKpC5DkstJSJXrfJ5vyRQuZfQTo2UFgse4MM6
fAxtdhBsv4liuudSYnPVPcdSw1C7Fb6oxdpqQ/veG5xPWjjsUNqFKlgH9itn+CGgnu6YimE23PgU
wEsVySSpQfwBI6MFIWrnV1SxdSq3i/VWWEFWwAk9fMRFQjx/M9cQy8coAAQZnCH9+pdKsIrPjNjF
hXUCqyUMt6odslQ98wHc6V7Qj1avl+b2A6SGd5n9hg0SQ6190+Ld12i0q+OF01mHqAPRCB3hBKN2
0N7RrRUtf+xuLLr/7gzrJDKmXlS7YeaGs5VYVqZEDO6rZwG08cB2UuZOIgsPycVTE+2QyZ91buHC
gq/0k7rGTwXa6zhEVKeCJINSead9uQ//ypJh3CGIYtg7zNrig24XrSPC6jaEU5w3633iXKuC/DPQ
qTDwqEkcZJoGndBbpE0ON6Ct+eKrAC5hI1zZbufrPs4cW1PqiOXkkx40LmFvZkyIjdWM6Fe5Iph/
p6pJHbi0j5VzoG4Hr62W0BwhYk15lUUzLRdJRK13TEWyNCZ5c6BIJuCF4vrakhOzTI7yU59cGO+u
BXA9cx8TCO6vtbH/XrOvhhTQ/0hmQTfe5vhtnW/HIOVOrbW3TB24KzbrngDBgM6CcQjw3P76IQP7
G/FSSczSww1Gx+6P4wWpOeY/hocBBjmvAVcdc4dZU+PA/GS7zocjayxLEtmMTCZbNliBOPxDbCug
09Vt+IY5DLbR7VYzw7afIodNSJZ0FO4NDMjExf6vibBaPnXfpXYFkRlFNoJTRMmd8VFPdPYJQ8UO
lCYDxOr4V24WwB53BJcgfHBoElj2/Uh5qBIYwcyUPjEZi3+gk1cLG37eyBCU7qdRcfYxsTb5p51s
mCy2yI7QSKI5+/UasmBPKNISLwBU2rr3ZvxYsSvfweEbx1mIYfJszxpFkUZM7aCqpgtb903POQnz
CX/PJ7eDUxv6Rk3eFu9U8CcGi6er2qPaKJ2u+c/kWOUKakdFyrvXu3oJ2pNpcd1kBV+sulabnVNZ
ai7rEGYR28j9SvAepLtqRl/dzmSDT29smdQjrnN8O4Op81pk6DOL+w4bt/IwqY73heBvUaNDFPrN
antpjvBgcVh9X08cTN0q/e/zGUYz9Ud0f/qJvnIeb+m34ajlygag1XksWixt+Im4GhodvDLZNo+x
ilBpFtTzGqZ1mEEphwxhJzWGklnVeSvDoulJhpOt+0D19uhNGVidOvoQVsSZJm+OaLHmCSaSHfTC
xJ8cSltpOYvNKbs6qffdMyH0xTyn7T3kNR78aydNCCQj5Dw1lba8YYOsIplGtVKp6fgMctx8g7qo
bkNRP9Ek+n2gRJosYiahiI2nTVVudK8p2KnWewOeGAY2kt9tAnvV6VWIG7ds+E2xIqhEkQ+bdXcV
u5XFG0ELfgtbuRjFeaZh5ULE6BAfTA979WgEHKHMAM0bNIlrDk86zpTnE/qyceWqdwhIHzWiP7nW
hGSWly3mDKdJ5ffMAqJnBx2i5OYtw5XHMZKcLD/gh5LTsq0ZFGqs5OEjHCdb+Cd1obgZAUJzGHeu
ubpz1knrQt6C21TtGm85rqI9F/NStfje1OrZkjt9W7QDlMvCDhQU7JPWwGPqg0NyzPT0rnVDitH4
2N+EfqIEtdT8hCXxAh2tkAVmbtbBVhuyGktT2FBVL+DAqWUcCZkaE43sU18NK+TAxNtFrTGCWsL4
vpkce4CIeAZnRINHdMrYAgXvFq7yQxLoskldplPL/hiKM4x2EvghjYlrM23Qa6vAJGM9n4SzAkC4
TIuCkSAGjU3HlIj1AEpEyqeN7HZZEWTgXOdFz9F7fUjZ08fVug8IPt/RS0zT8x0Lu27lwcG1BKb2
vlIzfh71eePbMTv1nvqacBBPVEP/IoSTdjcSBRNNU6nbEjOD3yJHYNAEHFdgjtbuwfrnpSccVNVn
/V7bIHoSijV9rkcAAxGbojpkMwxwstIrL8vf2wZdJ9Gh0L6e4ucax/Cd2Pu+qsT1JjE0IcM7hIT+
mQyMdzR92nbirCtJIEx8lrLnOsc25OJtJnjfIv7NPM3B1ToRuDDNmy9OrU7PLmNcfmpcbIRUO94+
L+nev6GI84ioJy/2Y6OQF3xrMDuz7vFLlr4GMEOaqfZcaWKJW67SWdxxwSCYXF+NzG4cDwcscanN
ClkGy3pvSKPYFQhRrq7uEz/oapGOv3rC/BRFHKf2WrfSccLv/9fPh+TVxbNg0YXObWEIn+fKlPJ4
AFLeb8Swzux9g9Bur4Yq7IXtDeOf1326Yzi+fWRM1TiKljZ7l0jOBN4I/WJtP7umyi0arLmFNNgT
LJOlRCW6Mo682dQPJJwPtr19B76bPF8qhZLz1c3hVQoWzLUtQnyg7Z5QGeDIgPbQk/itzTTm6BhH
ekwwZP9plP/kCD4LAtGTQ/TsX9xozVYBXoBDSlnym24Rarpz/r4+gfY5LlRFU9VJ2lEZUz43Jbrb
9eWPU7eHm2KyIX1TY04RbI2DKMf3NBLFxR2oGBliDAEnUD8b941EUQkJ4aECy7u7Q/HiQ2bhhGkw
MsUjgvMZnA6Q5amYP5/bKGw9hHnblS0R9T6hbvMFDzSKWSNjhd1glMPyCRUoUPTnVRWHvj3faL96
9mtO590LyEgoQcgQZhTTtcGGyCzLmtoGcn1u0Y0nWssv2HGXtA6qKYS+nQ8wy6D5XDTm8Lozy83d
Mpi/hc38zdG2Ee+AGCMs4C4SSRk462veuq0gfVvIzTm+t3pOUjnWVXVPYMz0T1np84NWrmTMTAm6
ZmiPFgj4UJIJ8YGBR8AEAfm9lF8WW4IKWM4Zm/5VSIyJH9b1jz7MPK7GpaQ83UBU5nU6fkh4I7eb
9gzYc6wrj9BSFYtCg+vsISwoXaTGJNKiN9OGvI9pygS66yg9te/dGrXzrQd2p2ziRL17lbNWjf+9
Aw9dSfgvID+EP+83T3nHdux0ESIjtBvdtXnlP5aiksoo/4hLy6cGe03Q6qCfE2j1ca8lqaVdEpFY
FItZfqfwsNn6eZHjwkUdCJk3hdrj0vSFj5RTc3rTSsng4f9ycPIoGgf04jn6cXVstfeiCmX+kSgu
2PPRnh0gsNuz8yKEgPpGiggGc3D4VYUHm+zo0H65L/hDXCFYsaxGwSgW91Pbwxf5+T9OWkLpV135
qcq7ywFqKbHlgY9/N8SJ7UBsXVdNKttyCiDovmrY82co415owDeMGaSaDs++1/1en29zALioX6dU
CpYBYly1jzQwWsqKT/RVZDocO+HT0b0RJtiJs8OQ2UsVVfUOnL2+uGMnwTuy0PwSHcL1VV8LhrSZ
JwOAjcXFtiqqcVXR5zhRCCSXlmvjE9o7W2sA8BSYoNZkb6J8s3PCT6RkC901UDih0AD8pcx8wKyY
WqMPtpc9f9kYVHgOY2Gw8Bns4N9zYqUATrcnOPf+b5hX4Yd5aBSV2QgtcatXq0v/6+F8zdlbJzVH
l/kAXhefjP3lJtPYbJlaO+FX0wiZDIInu+0mRBjpLs9SPXeYJbNTYnZO1ObI/mkHYF08yJhMbt43
nkHq6V7+83YmEliDsQClpjUzkwnjKB7bMLZuT/SORfLgqUS+/U6rJfegUkL6yVlzKc3nlHh4e9Gc
NgOcOYCgbq64nX11x7otSFXwYgIz809IFwKIlD0kWnpr/pJCvukSeIu1m8QECy02BBV0LGaUrJS3
d5P0c+r9qhUpfqvXGBsZm1QEhLy5YCkjDtdirkdq96Oi9y6d9wFhBOWQNC1xE+Gx0Vmq9NkelM5/
WU6c4TbjvUDGkwVM6XQxj1DVh7j6JcDTSLTHTxDxlHv+RUSgYGT+z9Zbn3YNafbCtSz33bSg9v6j
YxyjXsTUSeRQbc5XF38h9MaOm36fYdLB5Vk6vP20MOG5iJc34eHcivP2Fj0swZ7nAiwQa12wsfln
HCkOBzqiSDChMWjm6+W3/CGudTkIic0fvfiue9yQiBTGjlvIxRHiVRhSR6oj8A4gwLpivRIi2LAL
SzbiarOmM1NaXEXGWnYs9+8rUuPSLyGHeIHGnLtSejvRa0Vyaw3ebWF0nzYeiHtWG8rGErgslCmH
nd1rqQntAZ1JgjBrJ9d872a8josn0KL39zxqe5N22nKe3E9hNbcIKGtpabZ1lGmcx8kvMOXRze5J
vrz1W/1Fb2syx9wr5WdllYdRxQ9DNpNYOUmu/i6mUE9OAJiX1eeNP1svbntQWILTu/sw5NUGjVss
UbYTu9LpIeE1d8REGKDoy7jsIL4xVp6GFrefiIjp5A36x0J9A6H+AjxjJPZt7RMu9R0eDdCIciQx
cw4v7Ickg6OWzU4EDKd2m3PbcRcyX828egPbgZn0kjP/gO3ZqgQsV+UeVY1ExN5Ox3bTwhUJbLlL
cKgHTiHV+clK5lq3y+iYidvwPfEoWUStSfYz3I0qATDyUsV7iicxmMZbPTgUqVkhdOREfhOtmXfV
W733PTTafEzY+ZN3xb9CUyLQHWb7ENoDmQ/8Jh60nir9bq00guIbWChwt7NnfMX8B0X2TUOfJ6xA
IVwGOwWF/L+wBuNzH7eWstNLK/6tacuiQdC0oVIaUuxtv7cW/h+XAIf7vCIyNXxkcZtrLrgHWe2f
Siy5La269REW6cmaB/I6JEmWQlLrAr61RbJuYj5vSloqK74kH1WbBPpwEgIgjPbCOBCwkd15vIE2
ST8Nz3iuVg74IsgyNRxXXdW1z9nnt7sr1NRTfZjvmuY6rFb8vr2xXWY8Pdvs4qvwEwECllOdaUmG
+XmKdol7vMmwXJ56tQzsX/NcUIU0UGKuo87snBPTQVAmiY76KH6fTu6SUkCSSwjylEwZH/8N9DpN
go7Ci8A4EMWqZu/ALOFEvnduD+zguZz9PLe3TDbWxdTam2JaEOcJFvJihpb07K3cdNjH37X5FpRz
l3esMkaT3T538h+1yePdhcy01NcywIhbnwE9tHAhSjrbu9gUxg8ZXI0GOcKJQezwFNvYD41DOZ0h
R0iNpEhHDVJ0YNKeO3AX4pWjhjhJq2VUH8htR2eyJdze5M4mzkb9UHaMOYl5TGYONxmnz7sjnXGa
gozCrHCTqN3vk7gHUKm6k9S40mHuMYVNo5wPDTFasQ+vLn02xzhp6ddkarl1Rb6hNjlwL7Q36SlV
FY6iU9/iuj0WUMMmdjIeVvzdwwf2wZV4xxONZD9ZfI6VTDOGABBVNtmIO4yYfwLVuGdYkEAaM8Em
Snx1HRjE7uDagB+WnPlpf+2h6Mq6csKY0lc/2OgTCQWiXhMUUBnpvyZbkxLOyMaLLAFVQRrqAJ2W
N8bF+vYQ76mh2lpdS1kViq0393CzHd89nJx64MAJSGwt4JP8bmLgX/hcgTeK6vo2MGmyKDVM9Chl
NEBi6lU/zsDddJJWF07djv2+e8hDY2koaGkAG5sx0WtGhBQsAVmi8d6legr0cl2p52HWpl+/PjXN
YVWu0/MGYRmtLqbnIAtWBvOxEgG+AEL/apwacGssCkZmzMDTyvih3xZAsqF7QGmAbisLmNiB3lAW
mruCViESSf3MYiWLLKnUGvUVFsltd7Y3D4zF5CJZFbzw6IUh/2l6cW3+1mNBIE61/7O38Mm8ilB9
8Fs+tJsCmg4Jb/bfIbKBM+O/Z2Z4xf9yYBvma73L9OpxBCZNlaA6d65A47vpnjKPBDiB9qt4jvfX
eE0xVzahgq+yeKeeKB5X4UouJyUsr5Hh/MR67NZ0Yy6s5syAMqVtbbLQ22ntkZOpGsC/BfXkoUX8
aTEem/LNGockt/MRfkW1Ev1yrIxWUnI1iLqZ6Fojs9RS4cd0XiJyQEGyB4IO4Et5RREivDSR2uAS
tn/fXCS7zgXjKlOq6D4Ha9n9uOFRYZV/tJsXboUnWGoyXPt0fKFiCBY12Lzb1ggwoDQW+CB0b8cd
NvyvRuKgi9QeKFf02wbe4yCheL8UwDD1b/mtn+WIO5sUlp/6Mp/abm+dilsPtLLdmT1dBU2oLbvi
TkbOnhRq7ZeZs9wGyBQZFGWBpOkAmgm84c9CmdeAZttHQrkKq1eZgABwtHg0zxArQ+BKL5wBrlfe
WbUtGDp9CTa5GoJ/B9FXRW2G4ujPw+CKKFARpW+VOkbrUNFUrRabx2eXMUTQF/CE9Bz1qwvYWNE9
FE+lcUV93KfJ5XYzQum1XbRhaKohSSwo6EP+sGdqHSIRzQGvEK8sIs3LgJzrE0d7oMHtcVuxXUG/
7euF41OMVE0EWhOCEKgMcr1SaCAuDJy4ftMOyT6aUKE+VMV4b5FyGJ99B6H9AN0ej4DDgMZq8rWd
SdadzQSrn91ExwR16tluMQrU5aIMLRh+Va5sQJuKMeBWiWBmt33e9r0MGxlwILCbUj8kyINtN6iI
DitW2rO0+x4Zy3jQ+Pwk/XXEWwMdmlJTQM/57g7hEmXmbTuHS99/Elm9Sb4Zb/qWNyYrPiJfWu1i
2qolJiFStKHWc09kinEDQSqW3r0bdJTMHJgP6mu1InN+37dmcoFNeGVDzn07LWCRTlRWsaLjoA9q
8twBHbw1ZwQ3NOD6flbewgxh/gSluRQipm1m1gB/d7Z1rEfqs/+Z8r70Ns+3fH/DnGtgB5JxmByI
kj1psNQVuKzhUZ4wTu8C4BSxnie/wLn3249XUhi/OCq7WBE1rTqzqOhan8vpyxPObEAVK/0nBNCh
0k85T6Im2v7U7kiXEWqz0rneI5MG4MSZgTPjn5NSiwTr0Unpjzkz/9jIyd4uRyaIYsDHxOBtCyqa
pVlgg1r9luimHT75bP1gq3lPVES1zreaXwMLUF/6MWJt6kBPujmXMb1r7fOfVIqwmrIgRZWeyKTk
kwultqZgo273cqqEQ3GvGH9Wxj0wClAh3M3T/MCS+P6hq3Sk6hDaENoavqFeoiEesatL+VXqx6qc
9+XSO7OfnPVB195I6A2+1VK58YsHSLnYTplG0P8CdFHIdoQEi6Zthw/IJCAzh/khN0lJ3+bwTdQI
V+C7p8IUJfbXwon+G+aGXvqwAj9m/e9vFPKtqRkyCoEdSSdyx3ys3Suc35OELUQah3svq/MSRuvr
4Gk0ZfjsurczS0xZxQyvYUPyUAsSF4sj4Xa2bbjrMKPvy7kslwP9ZzvAe5KRvmyS13Y1yvx0vnpo
+wsVZDj8JtwjZBHv0caHHybRmKfaxVrFTpgil/djVNxXT85Tpi2cDbVSDs9UovDmM8J2LUL8GpKG
/+2vZah5csmLuse8uu4TWk7DYA6YE6cFPZxFPFyUjSYEurxnvYQV2gH/O8gvcHKwRof/vz5ApfnI
MzAl5GlZUwaaggVkD6pX63m00kN1uqhOJlaCk7XCVaT0SWOm6yOZ1WiRLzLZDmFOx1SOUMZK6Kjy
XjlN44nkyiWlGEH30ZkLDdKkXjjVNAW5MMk1m1XTZyXqU4bixCPHt0D26zarpaQkACwioHmWEpG3
cPWqY2FLRQf6xPs6z++hDz5pyREjLgZmUD4VA/k1EA6Cq2KLb1pW7xsvHOL8LoUMWQHkIIc07EuF
oBvejTzg7lboQZAp+T7xYlcssrfKk/OLXqcP5xmf96p6ZVxl8U5HN4Hc20/eflAvBcoFdmZVGHDT
G773S/zt/KojgNJjdA6EkkajuFaobFKFy7t/tsgjapAWtn4H/sQR/9tNDK0se3V13Qh44Q62GYAf
7MImI8HPoGMNwLrUu0QtHPrG2NXC/RTpzs8H4K4MNlKQFhgxRp/s8gAZB68CjESl/cjw5Z++a9jA
8jXDi/ebndwiFGc7nT+jNMBoJKS6gb/55C3IMGwSr7YJF5ZAqsA8D8SbFr+HSgNfuAGhTUff/ohJ
xnqLQqVDC/3uIRTLT0BoPRWady/i3tiBubgeGCjeBuyToKVy5LJFnuAedy/hP4E+kDJT+4PXNnGx
QY9w+c2agH3hhGzp9tfylJW6i2nHFNEohtYLxZnNzzx8duP4GK9Ev2PWpkdSYsJc3sX3nK9V3nkN
IFteVFczyzegv4JScsphhAs/CZSJg6RxRpmALuN/NBYhOOUnJsxHTIFfLRviNwOjzuS019LOznzG
M/JdKg41GsnpaZvo4P/7wC6w5oyBZBxB/IUImrfFvJEwCMLLTOiQckW4aSKXCY3gQtr0v8fOkuMF
E4H3UXciNcMP6hP0CwqsMg0Sbd7qLKD4volaVAhH5+EsMVddrFNhJJOxBcryW7cA0D+t7Llas5L7
Ps2oeMHXnPfQIFVtdfw2gO3WMu34AcWMi+MFwIEqA6hD/XAwYUkKFyVSZyCHklaFNF4qatXN75R6
0ta56wH59wNZy0ak3+aUpnfNYkU53vQbqBNaiJBI5TaYGk/Y0rNYip/DDQQbKWZCdLyYr9P9HZYC
7i7UScXFdF6lVhi0Gzpr56DIxSp6ibUh6wIvbu8qyHphEIg/OJxCxM/apHmJKkfb72eGe1Kwd3r+
c64myZW+ihw6T9wmhdTcj+/c9jzYEQbvS7sTVz1YDZlNLS8scR7+Xjhg4j7n+Cv/S7u3BDYjWviq
nUkb3fGhyRe2oYYGcnCxDxSiwLwYyhhbN5/5Hnrnqx0Axjvh6LG7aRnpQ7UuDLfiuYo18hQG9llG
5cU40Fbzrr4YhvpPhVmx+gcgUZOo8G5RX+/walMcY/amxU24qbBdQhKKf7+j0sLCKPwt2sbkzkWq
PBAK4VYXzuDzwiYxIqsb6fxel7vMpMlL+6+JIgU7WpPHJxTUlQQJJ/ORYw+xnhJIHsiiHnbjPhRO
Ju7EGea3DCaF8H4fGaf0Ckn9ETHWQSMyPg76cHflq6qWhoXF0Reqng0viaoGgYijQV3KUNAxEZ+H
XR53QuFinZO5gJcs1IEdN+ChWcWnERZOjP23vh2S7TEOZHSAQqXEDqEVYYmIhNdgwDTtEgAVY5zB
i39uztPZPq37+tljS8JrhskDTU0lGg1VMKHG18uB2uoaDQ9cuZm+xtXbjg8klJtkPXcf7XV2dTHy
fnddiTuIUyXQwnbVcFQ8SidaNCKlqkIEfaPYFzUmRgS0lrsOQuDFdraZyCM/GGH2ZDYHhMCk2FQn
sdkfvZPHLPSYt3uDNy+3TjGXrSxUMjxbniZvCw5ipZN/M8WOFJSgxlcBox+cA6XQP2I53/3Zinm1
DSG1HpMbtSNHePgqupE29sa+KXuAiY5Hpdbc9lk0+RR/g+y82Ixz71cLQ7/IcBD8EN+RxWOUNnWh
ikjnntd+lIjE01cdOwZta9ETb6c02ILhX76GhVOFk3kuaBPjVJRQcMRfcvhNGqJ093EgaKCBLx/J
JtpU2KzLNiFPK38jUfTCtAipD6yOSOA+EcYpo3NtHRp6IDM9oOpY69fNCiILy8CfdGUtWSe3Txmm
7KnyVLfG07Qnpc666CcBNqFGsQ9ClS69a/oetr56XA3j7rX2RzrxmHqAZhWEld6p1zuXxiXNZPCU
CHzhqE7kGqO5azuOSMUoYPRYLaKNp6FAmaoEZnCBglng38OExHLVsiQhekbTnNFZg5Qzkt6MLVGX
Ns4SRqgUVX9WJNVOANFbkXVzdJoVEJftERK2CYyaU+4nbldkbGaWzKQ6kL9UxnKWITZ6SdUHbp6q
aMY1hPyUSPVxz42msZNT5A1rHJIoFHRREEu3avgfJueG2wtbWiZn3tZzL0tpFPnplzXQugpCLSKC
f4+rwwtJhsgrCwxl5mulieePDBMamcd3llExJv71nh1LkVuqqcX/PiDJBG3rZa+wWEiyRQiEyBg7
lkit858cd/aySGk9PLL3CHwfDuuC/pOsuzbvqlC3A/eJEcaNv3zCg9AaRYtHwvOW0fDa6y6xNvFq
b9/+oY3YurhFPolBq0/pADUQkp7jXp8DY8bONvPAvJMsjzjPV/2+4g3ltuodxtLeZqfO4VVEolQ9
O7vjRkaVlmYuQ44hxLnxJcpMnkpqnrmodRjHrYW7MrIILuR2qcf0LKDdRsdQ2mznlIEFqV8bPNPR
Kq9PrY/6/vuAxFClY38Uxh1/4y3DxxBYaVSrKD8MR2SQwqiYWika22xwMZ9iAHI6BKNI3rfzKXA9
mpVcKHSJu5PqnoqW8ylAxJMJ/Hlb2MORn/CZ6TP99qeK8SwoW7ffkol5k9BQSF1Gj060MDnM5+qF
+eyqmadAy5qeLNwXvHO4mmM4MuSuf1dUsEmp0uCbW20pUGI02PVOESAy53Jsvm9Jp4v3cNGA1Inz
ez3g4r9bjUVer3ak+ZrduDmL+qCm6SKbwl5K+t2t4rqdzPHelXUFE05iNsc5F44jGG+lVkx6aHMJ
LAMvd8AevWKc5AXogjpTRjBYhGH8DBsQCgIICoQi9fR7ujusEZYRnmfBusacUiwwtnPtre1mnTUq
4JlR5e7FyNS+10Xt6uBHvodWoBUMpj2kMy7Jk7RtClUcIvtfEqIbdeAgIl9pcRymq/fvslHWnPny
H0nIHdFWDftaJhxzNzwKgXZdaewR0w463xLEdugid1PSdfcWxRqg6yBxBFJuL7yLCxKr0wPrPVNI
HQCT9RIgfZAGyseqS8N+xBPdm4pZORgRCpVue42anVUhIzlf+ETwLKudqUERXPt6V3z/xRQPPvpH
LmEoyxLEoyeW2O6gxFUnsaByAPWRxBUzz2nwSmDnmUT8Di9lzN8Tg0TGrDC7Q/46mwOluVMcIznD
D+7N27rXHeDi2YqHUggMF+TCQ0Y7GaKi/rDl7Hv83tQiuP1QO7Vn8CFXaD1XrRUImIBdD+8+hZjS
6ZUSazsExz776N1EaVx69bhw+uMQJETGETio3sq1XKNHugIDjeAvXimqOVNVHAC7Pqpt3x382PxH
bBAF6QotgFRxYTrIIX4wn/LePa9cuxgIq2AQRr0HVb9CNWBR6aTgliDonIwgkNd8+j9jjAQU6LXX
YJnSzZbmU/axCNF541cVQcqQG8KtTYmUm+s54q5NYFK3KTsAgr0gURyEq4XdoYHY5guC5UioEkdp
EwbzXXhCtJlXQe7oi3sjY/t23un/VdNTIr+wrutvZVm1xIeGp3yfmc852op/KVMvCqjDIVwVpENg
wS7tXMSIXcri5Mp6r5+nbNPzI8k9UAImm0yO8n50RAAzJzjg9ddgzuUwd0++qJr6zCjB2NPynpmN
Zn8+kM0vOUPouMfkIyq5LILdFnZtMs9etlBTLHvQm/om1Oxwgs1RL0uME7wWTEmq8jeuqZ7vLmTD
23BKlMY/KXL+wRI46WQIudNBDnR+ouMUDhdokd7xKFA1ihidlwd2a9gY0MCSfQ8hJHHWoIXe4GJz
ntaoFxOA7e0m/hPeJQedrEpiwNlgcl7bZaikRzgtO7mbKR6j1ziIlofyN5McMuxBI5PZS+tNcWLm
z8a12Z3+bgioJ5s9RCUe48Wnz58PpdSe5f5C/sNbuI6fOsKYK8I9cOLdeXvg4+WS05S/9nFZrv/k
OfYWglG4aQN3wZfydFDrv4dNDmEDRIO6Fl3uxp4pERQvZQuw2waYc1M45+W4q2R96E92dKf2J16o
3Smnh7uddaCyLa5Plr0tUiwC1n3hQnY35znqSp2IjePzP0p7jtoKJiv2qEF2NN2BEMi7Apeb5d3x
F2rdGNpeygZO1ArnoaLMW92lIO4FID4SEzVoRuLq1qwHG0kYMWCAAoFcfpHu/CSqSFziT4oMfznh
AvXi8im3xHCZ05p0EK3iXEf9qyCPOwE/2fBu2f6SDftU9lQYqZj4zlv23GDvzYJlPgpQsMYmtcH8
mgRVh++k2wKK8+xR7ePLGLvlIqMBoFOHbg5l52ITIAZC+FOE2dVxxlszejldFzxfZivZIpPAXqP4
qGV/p2I9Z9rtNrA4UZP9V7ZAyC//OKOTyHTvwBfM13OAtsYXcPAaoqQaOylZocc6hqW1vBZVoKkT
/CvOySpR3nyaqqflHmOnh4/AQeVK8sxEEhwin9r4fAPyFgSQ6ZPTHALmsz9EE4HqDB5xf+cn8+33
WrlPhYw7koTjVZUkqOZfLMUYLaFS+Jji/5Ym3h3IDlTnf+P8Gd2iqLfdb/TzIs1aN0pFdk6My4/a
/xEOFMFoCMezwqvWXODTsSPm50yzpIFfyDAuUvYOXUVcszqlyGiqVUNK/s//evIKY4xdviyPc8DA
sUZFSy+Dmd5xYnPrI4KUgFrJ3orLy2kcfgh3A4rtT94cLGUTSEVYk8tWCESH991H0a6yueKreJg3
4EG8es3GNUGlrW/qp8LdkTFKAiXrVvy2Lg1+f1NpsoaK8QncWZtjw84KIVhDdbYC5YvrWz17JXV+
DXuNyt1fwSGmcCi3EaGx5cVu6/f2E+lTgJHw4cihLN8hAeXOqg3d/5ohVZoBqF/03qQV/1k/jv6k
6eXJlzCg4Pkv5QM9+S765HWEeKu2PG663WkK+9lqY9mTI3VOUq7V+4w13yQdi8qNXo/rhstz5IPK
uf/Kyn8aYobp1Xl3ChNrM2O9upM8rnPwfXd3qi/+JihxHFZ8L+uMUOM4NWvio/1whYux/saQC8j8
1gz93UoMQYNP5Cnj6ldlmdHWfdlWNT3zrl5pbd/boUvQUO4mdiydR7kOvBGolHWTvN0jjc3FOJIl
sjR7sooMULu8lyjqExqaQ59LV4Bw+9jOvhoJlx0DbRrIK3zFaUbKts5pWqHA0sRS10wEq2JIgNZ4
rY/FAxdn2kvp+l0VrLkUu2St2Dsmf1v3U5aCkpW3b6iETE+2Wmu4t3JFYlnE2mo6hvjYe/z+tb7O
a1Vqw8wHxkbqz2U8AJDGLvVmd5H2fpqjctAQi0krFXXzsPgWun0oGfh/bO5R6d2eE1qGHsrOWW2H
mYdQizd7hOoR9/xvhJeMv2/R4eAMOXvRCa9uRj0pxCMWBV+YDuXG/BZr3YUrjJ6rnx6awmPBiIjl
vE/zhYFzE66MgmDo5inNzCmkTw2zxa3czTTNMq+gUhqlSwOu7ipNtL+DT+8GowlYqQ+mRd6YjUfE
79kWQtFkamMItKWGjZ20eBOoEAAj9qbS33lJ2csYe0mnQfOUWvhHGv/iaKnHRJgMjvGPRrcdQYO3
rjvoYHpR1gzCOCaTS5VeTpVqa3NSZs7hHorw30sxv42FDxF/b7SoBsJjbN0xOfz6ePPw3L40WTMs
U5RoAq7GSRJhmOzGufyxMtAlKn5ZZYzFlwECSNP5I1FBQ6iDSY4MgjMhWc1Syd/uLk6cjC7ZRUCz
pEWoQDkOtsuVW5IGm6QuEsjVHdEPY66qMvuHaj7tyPPVui/RHlRzdQlLMapwwUzuuxVxvqY2jef8
NWsvRm69Gq1mS9ueA1ttzQcxIyx5ciO1gpZNw1gGKGZc3uXlyowkkVNkgfEhp0s1XFWNhypm2Px8
pOMyPq9iMlGAVAK/3PRQOo/7AZwc6xyKx4wbu7zDCQqqDsSyl8sUtTW+PfARu/9BAjjvGivlU/ZT
hhES3hZH6SoA+yTcu/um20k1b1KnarTwbZos62VCrM20qW3E3yLVcO9t0YbJfUukOurj8azlRoVJ
Si4XjysRPaPpGhZCTFxf7UwEeUK8jKoZNbspTOi82HDna6echxuaw+83V7QSqgS/aFL1SYU02Jqy
/KpLy2hnVjf0ehCLR5dupW3OTT/VdhbkS5W0QBQKHqpVNl09unES2fAVrKkvaO9vCbzhRb7dySt3
jlRHnGAg5L5KuFfIvm0BnEnFJsg8l94wH1EV2uVo79BZj9GEE4l0s1QiL0FzcMgOjFTX6/OMqlzY
hcdf/D6AlWxLPTXMrtw5nErFYduQkBvTv1waiNc+qS+BvazWKCUOkwPXqnMSjnTHPcOGFrY8zkx2
U0HErdexsFnZaZHT7DWSWNWFTPjJx4ihNy1oYZNHoZLXqHhBJOqE9aEpk4w+aSWr5UAmUtCjzYU2
d7xDy0GqeunKnmx49P7cdKRrLQyiwXThiBSHxXNeBZedKd+A3n0GGGQnlyuI3YIlLxxmxkdtnPW9
Yv3Bdg06HMDthi9s+0eqQc4zAMKJrIw9neinLxw05c+U9CAH3OCBJGrN6FgurE32CbUYe8WJ2udt
0iJONI1l/mzBec2qBouezcNMd3hlhP55H08sLUhSRCFkiV37rgliN3iWCliT8x/5SCFXK/cjK6bT
XgCrMoPpS9LJFfvjpxL4ujWb+ryPV/QVAVQnxY3IafKDRHNRBECVwzHZBojpLT929ncxGv3QnR0y
Osyatu2DKbKhAL2xPE4QoJ/BEqmYnK7d05FTiugb497jEXgk/6gy1RTeu1ABFjFCBHFNSmy2e/Hh
BLl2tD5jFmj30wpasCUwE5mGS2DQudEikJVP+YRBmr9WRMkdgv2CzZcUB0l3BC4VIpZiTAdHbAW6
05/83lnggLSEAEUIBKG46sAzjguvJFxKm8K8SRT8zdNMe7OgwXo8neENi12YUCJs5JfMNrQ9LORk
imuh5prbiJ1TDVflWWZKwBvJmzGYEJsZWuwZHcrLKcn4SZ+5YxJmSYubI89jZneO0IqdWI10pJmD
4yN33Bl6IyoxJrjLb/4N6K9NPLjrmQY5uJjk2VlCb1W0re2tKuGUuw3F6eJetTRoH/z9G0gSdVrm
fEvDVWtfFSgHDg1CBjwwsRtovhwOiwjaOWXPn6JsyDK9dHkaihGUM5cqikZxQXE32yu9jtTbwn9q
hAqFm/4mKAEnp1IZSPyKPftASU8nLQQc5CuaTiaN61jgzKzMFnfN+TQ+MduYHCGm6ZVn2gHwME1a
rDRWwyt0flcsmcL95xd+jYYSk22s0qgbtkaVngmDDAEKTaVoN6TPVNKX9a6yoR5UjTEmoqkT0DBE
+i/m7sq1ITKMP42zqXER5GUn2YtinKj6uzFJz6KNxCyYBbkqxuzhSRrxj9CHjHTmxT1tlAXeUJBH
y//TxaAWPwRGgGuVo6yaBcLTFKJLoQZcV20l5LpZg+BIn9r2aA03ezCJh1zgQAQyNVeCvpOUEYpK
Tu8qLg3LMK9Dh7jbhtjhX9S8U41gDcFBJcU8qcE6lN8v4+j24ms6pkaNBw3nAaZRV7v+YFNqhHHx
pQqTvbYBrs9GEegRQwHEIE8piurVNtcPGtpZu3jGzRabSDQwmRrSQZ1aQ8kodRZGwHWJi6aI7yQQ
YF/ugo3rToKL9O0+2jgfcrhEs/1t3U71w8P+Lea0oiAuuV5IippEfElvbH6SXmIU2PqYDFSxQrsN
ziJAQQoQxzPhaJiPXpZ9V2u1RwunOnXKlp2kXAM9sEoy/YMNqi1GvkQi5M4ZS+YPX56EKpnhr2hk
ZE/8W+/qvs81/8XAXYJpsugz+xb9Lu6g0erWzZIc6VRh4XFPBwMshdrZhApr2CbF0SLcU6VY+AQf
gSFI6WbsHgQ1t+yb86tOccpIDfCva8ye8Xeq96AfdLP2d9AsWsQoebWBANwokjFdW3PTJzoku9b1
G3Qkk8vZbc7QbRzTzT3UipqBPo0+zIav33BG90AD8AGffRNVrSvaEvTFNfMDfuUyRrYs/Nc8K+TP
vBGA0NcZGa1po27/zE0xfXJTX8IF8KGIoE+kbbbubP0mvAQkZAOnUnDx8/ZjWLEeeXmRD/A3earC
Oed5NfxrE+7HABo4XXeOp3iNlsWmPXwY3NQvGa//ccBouh4Kec1JjNyq8nwBsF/uJSCpOVEV/xB5
Qe9nCrgK58cELYkyc4dnrfjTJhjTPLtF+Lwh/5cLPWXts45JEyJGT/Ie8cckpLhai4bUVbWMHBvM
fOkkOOdMHROL86On2pjBtE6xHZpvfo49tO+niZHrkKi1QetYPYFH919MC8dY23T+7bYdHhAkctaY
r9oWCjvHPwEXEavzBdRYmLSj6MyWh1yxf8f5mQ4oeRXA4w5NpcW6dHjYwfT+yT7SpufZ43IkdMtz
VfeRRDDpcO0aYkfN3o5pcMERAxKjAILw0kVcRzz2TMK8DINCh2DnCraX3wnvsyls1oHTMeSyPJp9
j+Z9oUwDdzU4ieBTzbz/Gfo7s2UmpWtlU6OKy+Av8/O6Rz22+Oomyw+8lbcZWWFI0AZbRTXns5QA
79eNhFVNVJMoJF9SAEJDepAnSZw2QKHkQJkqJ2Av41jU6qCaUkjF2mJ3n0eY2F1kVO8671XW3+nE
JOgEskyC7Ff5i18L0CqB77oiFoJP3BQ8BwLZSfBY5rLAl4Ndbkms+v+Q49ezfw9LJ0oL5zTeTYu1
lpEeS87KNEMzE5ymG3TRIES/f2SqrIYGkvJq6Wo0FzkvJjqxzd4/zlRkzDrN06w4eg5tUJRgO1i+
2T0f/dtU40Us7RsuUgJMCbP9a3Wixz/blX8RciHm+GEvB8SNPPEh7IqQ/kmc9fEtfwGch6u31V/P
j74cjaLOvcF2Ov9gYt8uVPvFWddI/8+UHw9tnwk7c1asMAbA+IYBcPvbA6wIizkVkBEfzQClcm5s
5f/uYnrwTfkmidGr24VRjFITcw8lB7pT7dCqSkCiXqYQSoqe2r2yEspLM1JHO2jX0MVC3XKHbNoU
sdpQ1i/mhXYaMyavu27Tkrl3Kso0/22hSzsNr3r3o4aVGhFkNMW6ItbkMdbyuhG3KbjTb64qya9m
25irVX+kCp6mNNKPVVWiq3aNsrE3XylHQ0YnnWMW5ncUqqDmhrCSkf9q8I4DgOJg8KCcbnUgiy+c
H9MwH0BC0R6pBU4gUKLErWhVEw5g4xa9k1r4p8rVjdqP2PJTZVUTYHJ7DqMRUFayUgjIPzc9h700
fYStY93sVgWbHM+kVceFSemK6+PgIv4WtwvRml321dk3jBjrlqAmGxm+67JY0d+GdAsTUPzrQwDe
Ghu6MyAs67mIPcvlGNdwX0gFKVLqgLWLHscOaUHwpqvJfl8GvuF0C9oGsar4sQPoDPRdNzT/553m
MqVqdGZQDV6H82VyvR+FrAmkIKvle4Zsu9lcncTbCkhnTANUcb8DA93nlz4Uho36BT/jvQPFStts
4BDLFqqNMGwYnjXiUw5hoRY9Pb9eq7W2SJYdpW3V0ir2XAJuDlGR29uGhh7nuYQfd4e2iQt2NWoZ
ZccisQKrSVwU6kXRgwQtcHV+SUKVzYUDLAl4txJTGAJFxngjbHP0IcAObH38hx/u4574oVMbRpw9
e+UAyk/SNPEa/pW87WX7yjc3eOHEvnP18fnskCgI/amRSp08jDp6m5cJj1KtNq8Cpux0ec/FF+PL
+eBcWHbCl/nJtVRrZo6x8iwZWOAmiFKTK4FgVNczO73yrm38FnEf36UiJxiTZW3in+jCQNhj5CJw
ysCg7wl1ItE2ABHBFX/xSRcCpr8ePlurjNGpDPrbE12svfHtGDxd2wYhUaJ8qch/OU//0jc3HtTy
H0lFjvSDA+Zz7tp66uyX7fKwvfHQUE4rsynrN0XozwdwabCJpj0eLWV12f5VkEbZMQXC3kO4JGqm
muC5DJD7bP9LcwNoK+ewrU8U5LUJGugVt1WlRKZ22KIV3xE3vur0aN/KluHtAIQb3o3K7ADHCj/W
sdEUTqx3CZg63F27+FHa7IpBkspkQj3Q82thdM43CMfg+WViUUOLXUgodSGasa1uoVV2JU+nDLjj
hUxfLf67Nk8VyGQwRMZdDgitiYAa/ecS5xd6j6vZ/AvSaZQBKlyPVQb09f5TUFhHNpvFsrOoe/vD
PcPCfCxa5bR3WM6fWQaZsns+BYaoox6z8048qofc2SStaahOWUq+ya+VXIK5aNLyEQfi4/+eMMN2
V9HEC1RI45sr+n01DREd7FqKP4NLMNa+6GQ4yOQlrQcHXsMrRGrK3yxmt5liSpRlAabpYhHhbL2v
2uPiiK+uVD7yJaw+uGcD9kSAg6Q3Ai56gYJ5STur8+/LWkK9r6ZX03qsj5AC9xlGXeaV9x7+V1mi
BUPgPivBMYyGI2e8AEogYaiRqog5YxHw4bxdVbGaylM55lZH8ZqW4XRHSs1zlwiJ5BE9aZC/0r1v
lcslPOt/jVRYAC+QMBca3+pwqR9io3d0VZob8SBfQpkWb8YODPhYrsvGnSN+JK00c5VS+rY5FxLz
zHUHNPhgAxXT+AeBRJImgkJQvntxomfnn72mXZfMc9s0oCpE2Ilh4/ufBGHMS1+YBmnK7eYyiSh9
MeiTNGJRj87CF0JMfYmoCmi/dmqqrFTxeVE7XUMh2XxggpLmtub+En6AqZcXtCXhGjs8QpfesVtI
eAXOU1wVhcPlXSp+j0GJcpRdedLor/vJSvVdaoys/JPqYC2r8Xl6D2qmDMAEezjePtqLdnAHqlG5
G7/++kVWzSlbCXY2LCIdUDjXWYzI/p9hdAbTGRtg2L4HCW+0wfDh3YE+9q7GwQW6M0tw76QNBQkR
sgg1LOwxsedCHBs+YlZ/ovidr/lHhVSS9mAzXRa/T4GCwoYmzttc+7MS9MDz/D+j/v/ertxWrPvp
2UcueIVtlsgSkVuZ7sOqN3gB2t5uINjb0aYKAk4IXYb1m9n9bTjwVMG4XWbjjh9cTmCeZQ+vZ9VS
4SLahgpr4ENqmLTQSbUZEHR5D/eDxLwFXIJAUVGK2FD8YhqaqXzm6UTd5rtkRcsQ+2FbqURzLQQY
e+vcdZ8WUBZ2JPdJcraTFcRWvfcYJLx6WjvbJmfU12RllHsXOdcc7QZ4MJzlzK/f1l8rJ6Y8IemE
Tb8TVF5/T+a3m1ZaY3GstpVNMPHyo8pon9L4Bd8LeOm5iMvrcsIhbqNpAh5ceLkAE2f1xQLRgI4x
k1t96Anwv2HQk/+e/+8E21Lr5uantFc9Gk9PBRzXbKEbfFLxd1S2QnCvJrRNcpk6Jzpxn2LZC9ll
VpPjuevvwipzDrapu713YvXk+9BuVYKiqbdLLscJsraXJbqFBoQZKshAbVsFHsLc3FyR/LDya/zf
3PrJL5oABwabw8k/GAAAFSHXRJlIGANhWd0uRzY651QEZVNLIxYnkw2M/YfRqhkC9ezF51bCzdBJ
6oka1TQZ7o8jkwrXGGjKwN+Mf5TfdPelYU1L4RNRQYlnw5ASnTGz5lGIrcHzXG4TrlX2392a4RJA
MDdOBV+U8IoUCHaLUBFqaLfTe+9/jAFcsvuCjhEaKlnRXtx+Gu12SSoNyuxfO7pM5EqYgF0Lxgxl
y1M0q0qTIhS07AVyKv6uxG3ASkRNGcyl7G4XXHJO59Qfn004S51Sck2Y7LS8KnS7HVNYTbKAf1Wr
xl4NXvSR+pTx/m3vHtgohFwcuzyaU9yNTvPb8UUWJrsqCicJIwm94XOnqPsZISQgtesTLS2tRVdK
9ELwFONNfddAD7tFffe/RFME6kqW64uDjj5XXd04x0nXHupfh7uUn5xXh2Ma2x8Pcf+/seJzGMSs
TZlMIWV0GJu75jFnPIhfJe7lUGORlZaNu0SUttZx5O8ZoB+CXvr/pUGMxKPrdH8hRjWoFnl6GPuG
nTeAF2hD3UqXZqX2llbpxOGW+xVXfetRbxlwJfSaLIjlTHrU5x/IGPj+p7MQF1fe00qFOJbvH3la
ZFx36R72dSKN3tTuG73NLpgTZ1HVGgsvPpK7F5I4F/S7ENo858nAguO4IAtTe2/jGbCZyLHwhA39
eXUQZ2Q2lHQY1lgEJ94o2CeEsBbx9uLkP8ZF6F5zLXMaHvQMWFQ29WxBQ+UigrEAsf2vqKv0l30k
QH0fTvW8p1s71JzTPdLLOD0i/pVmmcJcHyegNGvx2vNgpINtVBiAjU18ZQz5SOFVswP/gatoAj5T
5untQgYagKG5FoN7fxTXRED1uoZXaSijcI6NlTu5qbmcKMWGqIc8TZ8sGLf20J3FlHRKHUi+1daQ
mzO8dgC9hL5O9ktbcaV8rvnXHWEDJuLF+UbMsd9X+h7SOHiZo8pWq/OM1/TglA7oq2UJIbOYFaU5
5UZvsShCNkl3kSaV3OOeajXEaDB9duJz//wJRde2mFPDa1/fYAav9BQUIDpFrzqUY89+Eg8r/O01
bmiNGajlL+M400V6aE/vvKe+j24zklM5FaZYSLvhsnu7LVSCDRpBNzVdfFrhxfqAqPfRvw+FDZKP
x9bNt+Gaekk4Lyrr1Pnu7+tEFhwcTmIOkNG0vefFpvkfiL98mg1g21B4vRqt1GUtyN7VpHq+SHuq
LEu3z+SjKo/jMGH+0u/fQ97EWoEiQHU4vlm8K5AB6KY571yxWtCygoQgJe2sbYDRBcTXpgm9FcNY
NvCHZIug+ik0leAv+nSU5jqrkx5HmkbQUr/OpxasdyfRvtLnc5p06s8OIMr2SryrhvhlLuKoZUKq
xciXcrlP0d4hKHuI6efAG7ZzKTX3qXeYz3LQpwiRQt057L0mSNOLhN3gVGHgNnmIvLUSJb86xEDE
mTg+fDQ25H74M72hzjdvl/9nydgsnf9MJh6aXsdGMgU8qIC4x0GG8XeZgT/65DQFzIyRtZf8YF9z
16gzG2QuiBIUv6hMUXyDERzVbfsus02MMqUfPgPuZX4Kdr1xCVGgzzvuxfsOFRcwd124bBy+/V+6
2XhZiaQu57fe193vRDKusN8cWbIm8yH2mplQV/MZh4B62MFrO1oQbUIOVmtbwXCftpI5kBrRhe6w
wd/SGN9dl+f7J2S0EgqjbLPgIhbgeQSTvzQ2dmnUYu3zDiXkKGla4mySTpTZgUNSQvCCzGk1OsPY
xsZOPkPAAP3k0UVMFmXOFvA3CM144DWram86ibpWGRPFKqJwRcaz6eF1H4Q5N3laR5X4MSJulXhM
oCYykAOgkSw9xQzwy7nh3rcsTLyWp8EOQe2taWFPcUWMJcVP2UkCYrDtorzRm/HVELNGtQIjy+1j
RixSbtjJTB15sWOEum2JbOlbqYDdIGdTfUKnrX/K0/IcJKyxB9RLBLxvyAVSxoYREOdqh+RyPeKO
Mhb4X4ii1Cd1x8nVkKhqvThf/05SR0By0p9lhZxFpkL7laGuX6C8mU///jl67oNLix/hHNskgQqT
gmO0w0Oykr8ZVSy+tX4gzHOWDAaZxoFlK+ovL4bYV9A2lBsl3KPMVSUK/jCxel3hSF+zXS36apCr
nhG7DDzK4eVJqSR9Wj/q90/Z1bKgQW0Eq69qtqa2eRjStoZPi62RmMiyaALfNaYA0S5Tzso8p3gq
++Ehce9aY0e7+ES74/V3N4ibpNmlMCk4OXpS5medqwnN6DbSYfxAgoPmFYrwYH4b9kC5FU8R8KOf
/oQQ4zxR0FE8kMnFv+ymu/J+w0n0c62RfwaiRyFfAX+RDzZ+ifyho/vvb0+tE/f58zT9osoKrvmF
Zd+LYMLcB5vsjD/hqVo6MeCyXxdJbcjw/n7v6LE+zvXZHQ2xabhYv05tp6aVlS99C9JJLiM+9+2z
DKr+0pCqwJt4jjBlXXy0diooGXjoobjvyQRj3XZXWggaCxA2uZ//TevZXjjMQz1UWFelV7CYu7E9
gv1n/Yi/lKjzChJc4DODH6TKCMk2i773WjbOqx9V/PPmnV17p8LGERdMJmUK4lcqzf/GqHwHVhAr
KWvQ5gkSTwCyP9OLbdaLDnE/tTAo9vWMCefb761YVvOJQ+7oAXszprwE1aj2nT/kTX5QRvOvUuSe
1PBGjESPMmuYrczVifR9iQUu0Hty0rp5bbWmNsAQdv3N6Bk1kKgNp47pyu5WKNMR5FFDWsYPKiOj
EblkX4l5MquPLg5pvIsvOKID00kBd4Q3MdxzpfwbuSBIc2DcxVNTtRTngys9rTq29DaXNyyFtz4+
TJlXRRhArmdpxj18Y1rlT5KBoNt4pDwgt1oGMTMom+pCgB+pSoSZFPOX3wOSoGake/5VwAc3vy8d
agI7nCn5osxzGeQTw+AzVKhWOnQVQMfHeVfr7vwMYIbGy0DS6wlSwGhNACLKKh3KEP9QftD7kvks
fP5H8SbUI69s7SoWnVuWvRk3jhyWBpZHE7bPL6O79YK5LpeZyXiYj8cWbK0mXQMrE/tOCnmX/Ldl
FsJiUfJbWp6oCLe42SOTocmqohvOxDhCjRcupp65FDTTTRmlACtITl2K1wSNLJJRfhWO+nXRfGNU
Qf8jCVxpMS4vgAVU4SavkvozuqWL+SAIp7RjnMv/9iFoTLen2qTYIrLNumQ6q3xEbNWYAxW9aPly
jM/mTYCoPiafOoxk0WGm9pIFV3cYyoPmlHOtrhdLcloxfuwezcuM0xtBdn+7lSqHN4sFKDOl+jwB
7hgebp7PVCYnXR6Q+3GCDgKyW0wonrM7UsyUymVyeahfJjo2nmC0q0GABHBo612rkDxiFlvFBS+0
xnhHDxNFt8rlPtuTFIsD1Aned39PE4gdxO/jjCq6Gtl0A4PGR08OBB7BN8c1h0CPoyxu1BDQosW4
in9D9ifPtV5Py71fTjwHXRMdiNf0IrJG8pIUcoEeAZ1HAv8REIX6AQ6R7zbeCfuEqSil8tSNcj7v
bQeOWZ0SBPZ5YhEaH9kECmkwUfrHHqWJ8FeftYHiAlCkG/DPbjsEMCu94zOTtE4dNXV53Z+0IkB9
8GYUnZig98P8G6ZpJ443rgMMGo37I8LKolz2GY/d9fxkmhQzcxyG9JOcvCaB/uxMAXPnLTsep+AP
NXUHAe/4Z1MJxTlEC5wm+si4G4yXiAtjk918WBlFI6GEPiICJD1JHt+bIO0/lhHm05Ckeosv5L/B
/AWHAxg/k2IkDsdW2n1OHxj5iLv/2Ksa9RlcPc/TJOHBpt3mKLmYwWWOQHApDvRsmbo/TuYvomxF
67vrlMEAaNtJQjVm8rHbqL6yUXTK38WStDbilwPolnA7/d1F8izm/pmooDun5EJ/EKBPbQkfVSto
Ge9rDJ/3VMk+a9hzhYKpWbWOWyuBUZAVx+MRvc2fpSNqvLlSOksc8ydBhQXjPRqN/a0dGzJBWi62
d4qowZYpzonXkxposNlhz5Nt5buzz/WIksavKeAcsbJ1W2wipXBa92ciGyfQ16NsHewetcMqBsDi
bgPsUQHFy6ReLfhN/NwEAsrq/3YxrSlMldINhAJGcsetK83ZA3p74DeHVziEbnb6CrCxO+rDZ1Lj
HfYRbCmCDa90WS0ql8kbQVcJcAIBYi5aeRxNmB7ydF8QYdQqFsma6HFELSEhS1prA23VmS/1JJqj
pT+yjTOkrTCIgxqB/ebgNz5wdnl5CkVynUCbE8WmctkgU7odlBmoyswms2sMUiGDDyfwuUDXZ02Q
AiU7MtYxQM4b5qUMAzIH+EVwG1TbBTHU99xYqkRH0vp5jJXd7HIV1L04gkUznKLm8z0aQGCJrVLV
/MPPsbg9+TsMJdiBhiwZOhC5mqD7bsadFp0Fb4FuV9JOcXf4z6ZK4xTbRFTo3HUOOeMCZLhl54NK
6nZN4YePgH4Cc2Ny1OgfEXyi3bpkg3ULa0v4eECtSdIPb0LVX2qT+tonBlw1VgqF0mZoibu+xtOU
IRHaTZ/G2kCSeLvST1g98bJtF6M0SOyCBbW7iXjeQ5EePIaJFiEk6Vc/KpcMl9CDZUOEYFsoZp1z
SA3J6cRKXSE73GV0dHPA/XPx0icFfC1DBCnkxb1sQZZ9MgZtghHq+HfXicAgvexqIwOSGOA5MCxs
A7p0ZeyB+vabisDmZjcJaU60tZl6TP7C6kek2x/FjSG/JWx2k92Ou3szjZiQKbFz/BkDG3YOn2Ax
dWuhD2ggZthxgFoeEgrG6gKaCFploUYuibePxL1Whe239W54yImz9+FuPZTuaEiSla8S84PUGCKq
q549YsOnTV3qa4G2mI83X6X+ttixap/jtI3baVJ6Xm/dYiMsulKrGaz8isDMLjugKzO/fLNB20cP
aRO+I1ooWHjaCYJfgtOe6KtrRF8vc9mat7DlPauokgZlJqqj96wrOcnx46vqhf/IYJAbgM5OoWsK
tYL7+iu8meb+L7FcJUMhiaFkW6InSaUdhdlZn0ggejdEY9n4fddEhzRl2dGZVYFwVnilW7L1PGhE
TyrrGvOaQOLCbH1dmFOy2NaQHbViTudMdkZ5hq3PVR35C/RPcJNdC9ylR8B/IAg/Hpl/GLMcFZ7f
/4Zl6Pw490k4xHRefu46mFegJOquPa4NuU3CcTllwBUtr0EgZFp39TgmcxhpkIxf/dQI2+01xxEc
5jZeqbDRFn4h7SEMb4XzDitYrbbOAkmr3KcwbA2WjS2sP0rfGgFqPaeV1TJ1YasL0N/8tU32InKv
WFj5HJTlqIK/PpVs0aalAyqh+ozo5GQ2oGWZs9o/YTh9GgPIb3s1XEIrMK5UfWTvRUkngrI28V2Z
Ma6Eh9w8KGUdNifPZxxnSUUGJDqg5+XvPi77fD/909GIG/P9P+W02Zd12Kj8YXTC7LRfyMQzFrV1
dosBwlkxisT/5fJyAnlwfyMtTjr5tHS0WFYX2EVopnIpEHWz7HrSoEpX4KXmfCqOtMJdKqdRYmcf
F5wPgCxft2v3Sw5NRzfijKmjtsWeXg+keReRkBkFJ+3gGo9EA4FXqDQt3uoXVCcBowCiDDqezPsp
2c3mVwuKg1HSF/JtHPkfIW4x0zML8VAnbA8x0rrX0b+7zjFmMECs6nk3koSZo6chcL3lPAeRXgU6
C1TyCMFH3JyZwWdQ+Cta5VcRupqX38WNgq6jQBUSA1ZXroiLq2IxzvOiqk+3QTUnEg+xZpoUMRPu
8r9QsBHeL8kSNd/KWZy4EBZc27LiSThRUzCPfqjfyAQZs7aDY1aRYpIuO9d2L6QBkmgGW5dE4bUW
W/n1543NSS+HUfbIvQM4BsyDj96nL7LgRr7FtoUP7oNViwrqTsr+d1kM034YZIKVy0CCbV94WVwq
thSEEVo506g/MYLwuU8XyfVILGckHv5SzpfY23Z7Z9nbyYi/ai9P1OGNf1CaydcrwnSElytIN+1A
3vElXiexYpb9/lbPMnwBxGSjXx0NDbk30/AT1Mpm6tkvb3z3cj6lp4Zv4uLOnNsBnnpEN7cEwDWD
aiSYbqLADrIRHXQ+PSX3qsUf2eU0yWqb2LLmVhkiixTkhePI4zIdMu3wgII/OxauceHMpzN465Ro
k/owGeXcS0/BsLwZnpnnznOaOFt0fC1Yj2oEj5vKxY2mUh+5FQXlS06sJpYBgBUAgvhh04orSpNn
ojdxSkJsdr7yTJe+gnYa0tK7h+DFIiPExO3sAz4rS6Gp8cuAx+eWPBqv7MaIOrPf9/kBh2oCs9pZ
A9L7oh9jyMzfFg59gzwW8g07rdCZPa1qqRQ3wtijo1mamZAPFz1QpRtGXjMfoVavrzmEx5Fw+fki
okDXloNVWkPOYS4NwYZHlrfdzU1ac8GIev5aDDV0BLxtvFDZBnz88jlXhQ1d2J3MBXSB8RqodW5N
W7JsGQS4YuOkzdryInCkm670pvdweQCdALKglSUQadIPcjVH8bcWFGV1l/tbFec/dd7279oZiIt5
lqXLS8oNBWnTcCZBKnmoQP21vNGZVxun19ExpYIuES1UwDzd3kzvkKvG2GDS+iXyjdQ3elLnC5hY
j+Ws1GrTAyL3KlgDdzksjEl//QI3/qu5yOfkI9h8M8LCmYcGH3w5m9S2Ln1V0BjKEW3Hvd3eG2NF
68nVcgNyoBg8uWwta6y+a49WXvYaDObWp3ZL3xOacAsvMSGxz/0ANJTfgRnLsN3HTTm5hfF9DEox
poXFF6lkZM+bveF1mujTermjWAAsI8XeJw+Ojjh9ykJUwBbHu8zUE75WF4Qgx8EhKjZU9IA7IREt
/J22WX/+/KUWFTyhDXLBdQ182cTlOvRZIR/lsZ02DnRjz+7mUP8RhV6zgx4cz23aXoQxLkshY8OM
SekX909AZ8QtveKPxkKHrkE34NEsBA1BBbOU6OOEVC51B7VyLpkZPpg0x5wsXXAcvNalvDeku6BQ
CcNjOXHqfPeeJpc+Jh++O2c+E8dPT6wpEzo3M7JWZP0T2OEnkcmfVvBeO0fxP5zFGGrd9Q49Eh3E
JhVoBDhyCDX41nLd1YfzVS1L6HPDPjGoeYZBsAyvvkt6OYY9z/YR9ZoG/rRC+H4tPuM8eSPhuG69
5obVa9cr8gXBFATaBr6OQQ4KX7YW7LeRtxwzP2QhdUFACz7A/tq7f0ySp4vKeuxb6pf5hpsy6ueF
9bpPGe/T+Disg6H1ZejfmFYmZM+rQLmCuxPuCJRyB4assUvhOlncZ0Nc+lACERfCdK9JokZKF9px
vwsiTI4XekhmncKdz6ieCDpZxN91RK901gQAjCODIJH0dcEuwTBmEMyVknIY2QONzmVi+bUfv/Vt
qmG47hAOR63rh8gZNB+kpbejsM06Ylf0KjnT6vdDQCxlc3NOEmem2pi4j/nLiJVw4NxT0+0vajQn
IhUrW7clZC38Mmner/bMVBUyzMdfZVSarXS0EaID0kpZID7NNpjcx0sRWDKLy+g2peUxGPkWaQkw
XKQQY2RFxnBNGBpfCU7A/5DGSFD4Qlh5TBnyQXIA1qpcPOky9KFFa5aJ0/wXohJVUgkfTbYueyfv
Mc33PrhN6Q8EXj1LS7vXHLQaKZD+CaMklKx1TfI+BHEXayYhG1T3++IMGIqeGJoJd2loUi0Upgxa
RjwYyUbNrIB2ZMqWnYlvI5alSY9HOVbIgOVeexLrpBiL3LdFBu9ljhJ1EGbIGAEtlkQZD54lJMk0
gGG1VaxuEEh/bdFI2bcDvGdiTyiD9p1GEdQ0DeZcqg20jSfKecB35OlSTumhhSMQqhujw2icsS0A
cu6TNCXBcJ0IxpAwyVc7sNFgLzHMcfiQBmSKDWbUw81ZiRXdqr70vrTye1cxXunjAWc7vFPkLbG3
cySjSSAKfF3+SLYYm2tOOexnf9zAYeeSGJhUBfl1bOV0BXXm3tnsXBn9tCSZVMZO/HRuc7V0lvYg
oWxmQfGIG8DvrMZV09wq4ceJq93Mw9Et/+GFwrMSDiWuzSq05bR5Y1Ni5L4iOM/4clU4kGbdnlGo
gZgcpd+rs7+2n6stT28SaSaETD+ncb6XIrCtH8dnhW0krGDZ329w9YbVyOI5FGCVdLbIcdyKlYL8
r8Ki+9gSU5a+Dw/mNg0OceE62lq1wl/KdL3e21Gzm5nam+gjEGLSMiGkVRjIyFoRRRKhNUEr6cdI
va1KYOBpepkw/mnSQgFPRmi9TRnu3EP6hUzZeb9DKDzM5Cr1485iABnqDsH3fLDmFDpqgNWBBnpn
y9i/MvSKky9nAVczVjdHvWBP9pJ9inlfIg6hG8pZi1I0VrYZLjnuAyX5Hd1kAAaxnaVoF47YvgIh
GpL2nw5J100DuV227XKZ5jTBPA372ERqW3baBr/CBIkbRwA7xsbnB8jcprjUaAFJGn3tuu4UG2LC
Ly0koeB81xLzevPvytw6wvM2XWrs2pGDuUFSw9g0zBztejmA2IVws0YVD2R8vi4cZInRQS7O1s9r
4j6r0OPlbO6sPqCTyLD6GQ7HZCqNUDhXH/SHby+CisGxQ9l/HAUaITW+lPDJGnqYczAl/hRU5GZc
X2eHWAYu/ApmL7D6sk4crEnyMLGB1A8gwoej8AatLf4a3l5I5Gne6PUJ3xZL4PlkztX7pgVCD1NH
oC4a8dvkoevZMZsjTj9J+LX5rekK67BG29EkHPqCQI5GR0bwMxa0dgpJqNHYMKLgTUZGs/2LEMFp
j0OgNLk8cFTjNteL5CHLF/4wvGTMGCq6M9l/9vykmUwNDnSRe4xHG+Mz9CI1xiWBgo89/dt+G1Qy
sEFgKVsNt+tG91QOLn50gOk7Hs9GqXLfXkMY4B9mjPlyEQO55W6q8eZzKgZIrfPGoGgr6aCgYlIw
NdTybP5TPhcIMrlRBgs+7c18QP5VTqYQ4gErcr3dmbaGSl4mblDILaeSKtQBWhoqqm2CcqFYE7bz
hcwyF6jfm95zQbw9ofVTyGRVcrF5gAybS2Kx0kgo+rW3TrqrLz4ahUO47qWacHZthez39+EnjQmu
FCwz6kuMikM0uKc+hnlZ4i14zh8FvesLxOGZpz6tpmyZh1gIXv6L5gwLAHZ/gVya7zWUaelgKt8X
ctyZxAtX8m9GOrwDtVfraroWbmd+q88dmZzMurCcMzc8+vTIFX4WvLlx5+7kIlkyll8/OPxiP34N
yrFY3pjGikwNjHIPGLtTFrSxPQ/7BGqMd7wP9OdeH+tevh2h5u2Kd6S/nt0SPQkiQAaa6MZUNk3X
bpS0hEYwCMISA8uTeYhOm1cz6gA4b7yJxeBwoR4HBPVkJ4IX/dQKKOcBGJpe8+lXnyD/HERB32je
t2omcr4GgFyh8f/8IQZXAdmnffDBc957qW1ApWsX6UXLfeA7bioYDwWetdoGNTpe/WYbXYbL3XXV
cU3EoUV5P01TBqeagmoZqDeaNUryh+eS9xMuQxpSs0q9LgXhyRIDt2tp0wpVi7YwE0eLsmyVNYVn
ixItGqtzGU21VsvUTJ6dXBZoVEnRY9JgTpI1imXW0+DW7hCoefxCFPYE/3Syz1+8Xw9IL/Q82bAg
vL0r4iOSOLBvPpHAdqQGFnKjCR6rDZ6vvSepiU78l3I04eN5MG5AG1LjA4kUVGk3CQ6lozszRN5c
E04yJSa1G89b1Mmz6YtQnYxYcq+lAML1asNuBw3QfjyeGh/tR7B0jD2FCB7upXjsskZuwi0UXWqq
EXDctdFUO65OwvBcS2CUbLvrQMUBAXRZi5fQ7YxgXf6fsvvErrgZkiAT0X1j93f1wEMDF986gmOH
j4TxDAUL3AFbVjAPdqBIPbfSIxSZZ0qZq/wNQcZsSjFss1Tj37HpEvN5GFQrItl7/6r9qWvtupJo
FCS1144R13RzsxytlIRByzMEQYQlIUnaAOqiT4AF9z1A6MlzN/kkS/Ddaj8y7F5HeyJm6Mm0y/Rj
hzdpikov2SiEb5dIoREeKJ6RA4q6Whlhdw2XlfiRglFqhtJZl09ERLuYa0mVEtENvrJ7RIU6fFvz
Mxf4FU/IDWtEOputibHasrEGdY1rqNarXJgToEVRVd/YPzkhTWirgIcLUGwXDX3A7Dw2pmqWGADJ
V0Tb5MedATz3iSgcHvuY9foYic6alUcjBHpexaWkBt9SAU99TZ85jxs8f0yDQR9M4O8TDPeoj7xt
w+aIy4/Tp30ocTqO6aWrFjicNgLpq7m57tiMvh6TjtJdhIt9gRtXCxeUtsZVifY27nltqFTBvpfl
FQR7MlNjp4uGDBrFoYBCJXo4TE9tPeWp77h60Hd0dpUZD+PcJQQ7MaZhcsXte244ahT9t+Ef+yxx
3GBqIukaiRD/2D4y67jzE1V4hbKKBIl7O3qFAPZGd9pxHmf2Wf3wY7ndXEs/1hcklz2AiKuYMmQI
Hdp0bjyIhb4JYNHQUIwRIoK6L5KingbyPeHamPNmeLW25a8ZM2BTQFAZGb9xwP/qaxXQzRWOei7g
hRXfFz4LS7yBdVWU6JkOjtmBAJxvgn7UGhSQIkvs+HB7PcAedxUhSUFzbPHHaee1hvri6qLflu5Y
fu/x/Iik2nqDsiKEra7aVEBsEDkBQYjBdawjKe6O5mFU/yvmBtFYO63P9gWhNlB8Dk/CoMKwA/zl
EsomNfoRP4fVz0bD3s/0K6HWjbRW5BBy2p5EgbU8jJx3JeBifTOVhQCWoyohgm7WfkD0jjNHjek6
cWXoRMpZjS3Pe69LkPfIApP/CpBkfMFtwwlVyyO1kDY2rZlaui6U0/PvBynEQtQLK0SzrdQkxCFu
4TyanQClMuhJ5sWoDdmT6emJZAV4sb4jPy/zypiUOKZzwRjevkfegtxuEPvgbC6VLq6sMn12Cx9e
BoTsXfwNCKsaKXJIHq1ba7qnTxhl0cef6DeyplxZ3ZMd7pADtLNwVIOSgESaVoAvWh9ZRHrt1EDD
cb7xoyNfPqkcMnyKHs9PJfMRhHJBa5Q9Eo8Jtuz4LhJ2+s1pveES62bKn6bC4MPx2s73Hl92WtHx
+U4iO7kTHkK6wBmORnYJhXX5fPj4+l33azHQxq9h+sw6Dh9uDZDF29w7fX6Fm9y8ZKyM2woxGuDK
TDCxI/kJghATqm8N1QSJQsN/hw2jjPyxTB/JAmHDsKhpuH6khie3bhpg4SlxIi3j+yKxUF6yk03Z
hFo2R4Q4QApgLNpQCD0nalANTMQ8RjbZZNsx8NR1yjFiFrME4CMR4gaua1TZBCGXolIFXbCBK9Yk
oDiy27E2wMgam9fFMtxhllL5F1zoNYhx9J51lL4UOPAAxiwTWmKO5EzDvLqgwQJg0RcYR9WIgoz7
4Z84dJhLokU4MuiqoL2qp+MMfy6/PC6NCkKAy0p6qIGYIW/oXWtJ6N2ga1mRyEoCWTAveznOdb0B
jlBRKsLtRKwd0mfuAFioNZIpTR6fXK/owMxURSxawfDmiAu9DeDs7MwLGiVDodr9Gwv/UmduxIoM
EOwRq/zQDbFa4Osb/mPO6pG38RH9XT4CHLstovEIFGTbkoKKBDxPPpQeUDv64Rcr/uI12LCZzJlt
EmYWpLU2mjBAgqP9fCw7trXkEnWstkQSqLSLjk7rzKu1d3aHf2XBKWWEwG+4EoBbuzbRN5K7uUO9
Yvqxd48QX7fOTg6OiyQCauJI2SXl2exw2YwF1DJHl4UncBZu5lUNfIns9XBK8OpP+W3IQ9XEZsr4
/7yC6unrgh9YUVN3RXd0zQDCTkcKqXBsp7T5WZzoy2nLV3UidvC495AdTyK9Ld0TDx/Phn0snauP
WdJdZoXNgBsiY4cRqzwmB3I4sG5x1l1vbonB+APde8LdUWKHGapxcx4517wO9D9So58024oIh13a
HVuSHBuDCtx5sDq6fn1oSSxRGsRSutgJneU5glYUFd5Hxjk+4ogfSJQRG3BSmnQ4Kz4BMjDf7UZz
T0l9YXoVks+B0QWU3gmse8PBEsqOXwL/AOJ5yBKSdlGH6NF+qSsMi+DkGYtFafgsjH3lH9j40J56
ZAl1qaQ9wWLBaDhKTR/JtpsNfrOpMrR5U3H56eVCSrXfAjW8YuQmfgsFiEp7c9kgztI234F5WPdz
FhiRPJnroDjU1ikgJpjC5myezKuGFxmJbsSAESqQgUR0CkC8wOFyddexSKZCyYSL9X3X1v0gHeuk
KLEef3oDfnOXh9GQnT8CiEYUAlZ764faR6hPiP9wSTDZ6igI2AMp7mEBze5roo8OYFh4lvj28n02
qZywibS+l2fM8J2rH51GpEzHu9R76O6IMvOoTZ6cLWmjjm57ayMu+aoE0fSmFxjCM6oiRdIWcYvi
tg6E2Osk6XsLpEiLfz1GQdKnDDYJG6Q0h62GE23aKuE6qi7vBEFiRPAX8S7uOAPDCBZFIFCXdCBT
2DQqM+6jnx3sY4o8OoTW7jpbECMcjfe/1Spx7WetGPypbg/68LB+DWYgJtBJFa+fdgclGZnlbdk9
IJGzZvR6+D7jmIATKp0cyR1pCsqfiUGVbSnw8VvapHcsgZS+oshJuqOGtLtiNMrLm97lMhQ895i2
/d4/fkmfbeTyxjgp0xsUMd6BizC+SIAsqm5R3cTNEAAS+mSzhrueS8L8rZGlYNZlKDgQtEMNowjm
g30SJSnhptBRnhAPuGlOMN37BlUyfkmMFL931amhhWI7yIjHMacXmijajOyPBdkpnma17HYFY/hQ
lXfYY4SptGZAXsvSEEA9RkNTj1xOpwuJRJrz3Op1KvJRpArPKuzuyx7UcyNkbMcTXizgffbOGlrC
uVHkG52nijZW7YB0UFX2O5qKlEac/zlNQYjtuyCEa0Mds6lJXWfucme+ZiKUeZ6mu0CaQq+Kf+Eh
uqtINlr7yAqhHfGEqPtZHPaBSMPRa///F9mb1k8IVGycjUaN8mnn6Ysy6NGkB7G1va2OtPQABQPk
H94yZML/yu6VTSTd96zvrvaXbr7SP25IdZKKYqepsNwupk+RCYvCZBlGf0CM3/REtdLf71aaZJfv
HQZhvDTu+bDKe4hnQ+jWCN0NTdMJtyNZimZA6sxtuNs8JctCWhuj3CqjooVgOGtgrXI6AsUBzvLb
xWsJZOoeZchamedPT+3eIWYIT3I09vf+RgV83yNqhbnr5mVx8slL30sIKLlsC9WsLbs5P+Cyo5kp
UoqWMcwrAtOBvlQXGD2LJ+XpB5yr36VKHIN1iwyKiBBZJhYrDqTBLA0fyeAbhSMZOneFhThxiAOP
8La+m7Rbe0QDiQ7A/IixcpJ7VbTJ3Mo1gqZR7jBqaSUtlrXXiAAvlMiXy2j/i1FVVJe6tIzRZkLw
lThXP9sOou6eZOc4kLnu8accVtI1AcRDRKuI9tV+XMr+QkWSvuQSUx5V4L935jDAZ9X/jaehmfjV
7znAxuZ1XEgUIdT0bRVb+Cb+hoXtulBipCIqBrU/fMEoHLlF0dBIpnQ/Hfl7855m8kXtQhOcO2PG
IlayBQWSSrgVCjK6v7rszqNe90mT1y1qDM99x8/0RsOIQsc2Wv9xCYd0qr1zIMy3CrAcoxahl2Q+
WrFfFHFoZb/E1qnifQFrl6X/8HYB9byUtkp3wEW0LUDjkb9qcZmsSoQKyAOKBoT7zXrv5jSNJ7I3
4ifdfJx0uU1q+fq7dIvp6UuN9fXzjI4RD3vUxldabIjXh/uk+y3I7LxBmJbfOEvlvKfwj3Fry/BG
nUd45FWsvUPeJTUmCGjrkQ4rli5xHecBTTgnLHjeXfFfFoZOmsipE9JXPk32SOZqsTVNmAQAOYLp
yA0L0p32G/qvbaPGuFXp1kbAd99vlb6z8i3b8863XAzTfNR32bIs75aEdfRx0bz9Aar1Ol59CIHD
G8gEPlOuH30rPbmBHttjxCMKXNhUmzqgIuWzI2ZfmvWc5uAxn19/bG6WoaONm3opdABB5P892Hu9
n2ooOJbbQ5MePNvwCNzFDW4Nv5PJIvQ7D7lzagJv3fEtzPIm0ZzZXzYjMuBalfu57QNkPUAuPWg1
lpYNmdB+8vpw7T3OPt5f5lCRxOYPcUTfpgRBWM1LjkwA1G27cEZZ6Ux7DPaK51s59/mBNwbyI1Jd
QwsVnk105oDmGs6VEMqj5KdpbA3/3+7cPFS3iC3JDA/K1ezjzT2V0My7ynplqCQ/zN/HLBUGzw43
fl/i7kb/qKikQiPXkLHA49MphVG2kWfpzO7X+pFIC2Vfbfu/Kz5p5C+tZbNhqSh1Gh7hENVyYbfY
lfQLUf7h9SHABmpHfufMy5KLqJNTymREKt02DBtm528WXQRXq7M0mHyr2qmROjeG0SiAzh6iwlxE
6oCME0ji4aeuSdJgi3yZMXwd0egAp3g7SUK+qGIZndPLErSPUvcPc9SYV7xbyWPu/6faXP2Tt4cF
irf47Kn7nI9p9L6CUMNwkdcIudRYDx4f+Oqv5LZuGLfT9deBijDKTTlDWZaIaoI1cfJQSyyDc3ay
AnzJVzVkcPNQf7u2KWdJeEo1GzYvvgSuPtDQXqh47d1JjOo7RXeegdgLS2YQ51n8H96rlSC1ef0e
y4pK5fQVhHoz2ussopMNta23s9Tk2w/oLWyHiLodWeanX4bPcx9R6f0esmnE15rRL8ULQ1GJGjR5
SPMHorFCZk3SdSN7J0XMM1noeCfUXTI1p+wyAAGZjRsMHZIHAQ5zeWf0B9RXQ5kY0b9ZFzocz6tS
0NPTh5CZdYzRMECqyZBTs7QhElVSeerpZLjDTwPVqD5RfsTYiDW2E/+xa182d4Pq4PfXpwlC2VzA
r9dBJ7W+IXQCKgjRkukaekKCMUXV+p4jZpGXl21Wj2tYLBnTYotGFEGdM081CIQTvqn2n+RXiw+4
jcJwOV5RWFDkCuCI8tgEeJePjZOkZmali24gQRJYrKu1scraYuc0wBhOcnZ5RUAFlqYByMwVTRwH
96LbJxXABkBm4SVtWvw8JkH0ZwO9u36cvHzc55jKfeYSzhf6fCWt6fxvXnlPz3A7wwvqxpPBlpN8
xcDCiWg6WRN7OfNJK9YAzOmRWVofKQMCUsuYuEY/AI5ZpFM81etXcEvM2mUrv0onw3gEYhSjsWRT
17cn+/0AVD9p2JSzSpeXMpGXDNTjRbjCgcDz2STjVJWYfKykTmgOstxDBlTzhLN2Nr1ZV8LYRbNO
Jy5oUTuzZDx7mMMvhaEGkj6OIA5+R/vA4gIEOIWaO6yoZjDT2ZbVJSlmQV8OThBDJ7xB8jIidXjm
pCQH3saKXmulQnOk9Nk4478GulAlGh5H0DyJUKkRrPCIBtKCvWh5+HBXq63SSFRvxzE3Ph95XjIy
5Hrr9aElgQ+R2CBizgh2HX5E4ele0iPECv+xm2wVgf1JuUBYZsMasJf43UKnLfbkP8wH0Xo8SsDb
XP3diR9wItAULqwy9IzuDWQaYXW+Z/5XnAx7AexNzU7DkoxSnrbe4uWVgIImUvkveyRiD1roGplY
4+aFB14zrJ/lXs9hqSEUB0GnY4lIc/oQIsA9dNNebqb89hkNdzdVZpdXB1nqaWsLhoHzfZ7AHRRJ
52GZayDwT3PcsC8tGRG64vRS7ITBwNmMe5xP9Hiy/T6XtEFkK7scSQfzhi+3dEE4rRwfXG8w4HxU
73nffSSyOutIHrumysEy1hXkUvxH2RGNFAN/EvNjMYqeRyiXXwxP00d7gSYZR97Ku0WYIPIU1jtM
AGqO/SOrfs3Z4sjFqSNNrkqzh3DlHi7pUfa7NAwY16FJrEbW35uzUTGhqfozGu/1azewO+GwZG5m
WotJEjl3grOhIj9ndhmTHzvx4zI/XHZnioPpoUJNwAJnakLOaIqN3v7eCf0qD0ZQp1HIoTAXrR9q
qbfal5t4SlIExqBK6tk0v3BtqWq7POSjNGFmP2nBNgSwK8YRFvF5+ed7CzRiSwvi6z6C2jrF7KBU
Ca0DG0Hf8IyJgf+9CEzMqz8lhAPpS/kNaj8saWRs1f46g55mt+YRAhVAbRMGrHzzysit2JvjcH0x
pQJ4B2aCsG9o2qpONioK49z0h/vDQDYwCa2tEM1T8Ybd+ormeU+t3lJ1JDnaDMHJcRYBJbbfs0al
gGUAzH59wgx9suMxIEq5alULvLxM3+sBtcW0ab2rJ58i9HOGdBTAsChXcn/mNhI6jJo4KLU4jAmL
moWXQA7TUEYOeiutI18vmZovf5geGizd2t2mRJkm9+dBujv9LCCPtOQ88o5LJTax2e8Odx6zq3YV
AYlf/BPl5LggpYGFwy3Y/5zYu+9iYfXffeaXd6Gy2l24RFal7Syw6MLTilh67oM5Oh/GC0DMAOQ4
0rVCuKYknB+8jen5ieY13Y4i9l0JhTIRva5F92EEB+CEA16L8/kmu97umn1uaidcvvsD7jK1r0Im
UEucNM4mvf5xQIoeTdh0RWHMw737IhQ2j318G6dvgCtHaWKT6TQMWug8aVzZ9n4UFARIxhUdBuDg
/it93dX+AsKaGVVPDjTXBFN2ZWA8yDUMpvZziqqo6RoOkk+JItp2WC+BOqOONguiSFAXL4S77xNJ
t+10PaPHTnsju6QXhJhrPgT1DWEG88VzhupeONDRKO8uZSy6yJqQeMTT+bIBLbzByWpOtdyr0A1L
ji5WHg0OlDvjBsKk1HpDZwFmVlSYHvMbq+O+LZG0VbUS5B51CXft3lYB1KyVwgJHMSKF+922J7aj
9WPI+gGEP8AcDmDlDGzD88m3zEIJuRyyKbjPksNQVwJ7vCY42myz/LndnJDH+K5xrCRHHV4IuoFm
t8sI6CEQnJXJ9JUI0955dbzQLZ0t8tpViaLtf3g00K7kjVvJCcj8Mtqi+/hWuYLsK0XQyRJ0tdBy
86C7JbVBfhS5swepm0qYN2ppx2ix+BcpurBV8FiOGg9MEGapZ4b0epcXE5Tyn3GrBCXCDuXPTTZ8
LT65QLwHD1X2aPAotlLVyozoDQVYzVfQZMh36eInSGisXANDKe+xSfHE5r3VFNFxk8V4ewVc5VKn
jstQSvnjxt1hvkG2d+m7bh5wFhLYmLD8kBy536d6zs3r56pdwKzoc9f5sXAsf8/zc5ObH0+4cCVx
H222fb+Uve3kOPP+Ojd5j1xjzFQq4H3F0q2sGlgIF0+lSBuELOUDPMqmzmL/PHKfFXiDZilwYY8a
fM1HNdR43F4TXSTuA1PQE8hik7bMnmo6x6HVHBT5thVctZN+WpdHbEmYr7lSUHqoNi4+kRFkBIEL
YUycM8MbVj2vBFdJpVWf5Mnp4McGpmfyLIMtcEr6mePW9ozImivEoQLSQOu/PvpnA70JQmXQW+xy
jVXnEPFjpum4Ak0AKsyC0t1bHBKdtPFzVpuiF5VwHsD3UYwr+/UxKCcLGh3o70gzIY4jeN3hK7Vr
BSViGY0PK99PCQugeCLRzTX7fYhYYc/IkPsPqGyvwr7ExEtXuzgad2sVopDCah7kpoi0r6M7BeTY
bJiW6n4wL1cLwu5a9QsqbNu0VlBdRwrRk8BmELRQA2bIwRJV2AqamRyfLoMGoPbp7WJu2TzgTEgE
teYjvcHn9z+436UMnB7ThHlcV1L8E06RteZkKXHZ+YwObQ+rtQIhAmZsyPOcYANHgR9ZCTCdi2ta
ij23lR/kZtMV25d3iDXyU1sTdtSX+ATv2xmM1whaqgv37edbv/R57qJu7v65fmWXlLX3fVYl7zav
ZC0kD0nJ91Wult3UTeL195uDiPn3/5EarGLMDbcb46WiN7rnxE1xwi3TTHGwp4zgWZVDnMIRiXXf
sAPhKdygotQQM51yS5uwk+0r2QLrZoN/2gXAj4HD1EBN1WLD3afHQn1AR3UoU1g/2cC5qbhLo1FN
D2RRsOSgUB83unrjyr+rK4CGuRu9S5zs1PhsBIrF5MtJHCFB2NKzqW+kB6ableu/h/2l6jY/GZhv
NchFVrickXBMF35htmSaVqAYIuIFNlbNT6FtFL8m1ytNgun1w2Ulla6Breh1Oltl1JLTT5YE6J+k
zpYKZW2cEKgwDLQoDj0bXdFSvPwsSic5oXj2u5vq0zVeWlTBr/27EExoKRf7wqVXDO1tsTJifcqJ
5rFT8/5MwGYtyj9kBlY1/maE9HBWy1ALFEW97QzfxxeOsx4EyIWv1586A0yoqwfh8o0GSTY9UoQ3
eiu8AMCowtAmlDzb6jiBqg5jy3H7cbm9258eI/zLug4urzj9FAdGHaEbWc3UPDfdcxhGhFi0GdMj
37/dQNVRSQah9ZpmeZZWXyiL/m0+vDhmq+3+rV6LZYGLNvkJ03XAML/u/9Cv1eyCy97Bp8XDS7gL
S8g0SgjdtezeRG+hQTlP+yxzhqBMaEP74urRIZKh+Sb53jHFhKm72EOJgQR813r2ep/X3A0i2ZG4
sByHgEIcigpJbDrNXFV0K/L6CuktQX7sZt8OadjZWB6Bm+ubZPmLDP5DZBXkSSmZYAub93i0Vi7d
gpiKfXonVu0RbfA65b8gqu7eQ6o9N4it4FkTIpU+2G+IH9lUDbky3WQg2eEqg0KjAZ1ho0EY3uZT
IVrRMMQhfEYFHo3Cxcn0NEY4xOJbIZvJdGUKYIn/fGsDL49ro4HUTi1K3SBFykryLWg7a7+SQsDU
fZTNsOVuwXU6sRIB6gAezeO9KmCXjHEQ9H+i0DuTskkNktNDR5mTfEXBtA37UXkzihvTuujKjl8P
HXCCRw7Bp0rTL8ZvlS80VzvsIEuMYbAd7xotljP6ncgJuSgrk7LwTGJ8Lmgc7pL9JUv5UsiKRmrT
5FbBRScGLKFxJYoH5Z2JMtzwaBvODgqkPnB5uB2GfNh94iQoWLVVOivpuuQvaxmBKdKT6ygy4pNo
hVntuw/6UP/cTAkctGbCEUPT5A1SsISYi5YsDnH5oNxxC6qwaLk4Q/iE20w/mtN1ZdJIdWwnmCLh
NEOc2gTNT4ZNkFV0If777dxhEIO0Z9aVugj53F2ZIscLKpXJjsxDgMTYTKW3WOS6bRlOcrKNhUnr
H8CMD9BEK9uPPGZcJx+2nvl8yNq3KmKthKBMGhxNDRds/Xrviq4ZldsTKsBGE2XeggjPTVfN32iX
yCQ3hwmcpzJlcmWst51FFXb77s0VBJjdLPPNxNkMDLIVvzSQoMRiIoQX5RoySu+kATQyweVBKonC
rqO1IpBPqQEo4to5mey1XqW0G2zADZr1X9fxGvjIhiFPnAUqmCsjIVOb9EuQKDpJ79Vj63+aFH0O
WUtRHeJPaIh/zs0c+vvpwPA0iEgqV9QgyTPZg6wfg/Lud8EcA2nhCMdmNrk+8KU2bb68mbwhi7P3
R5FmSN3D048i54CkemDRbDqNgGiccNHY+Bf1oak0GrpiSsndbazFpuVJ7NHBbSKyd+9QOJetERhS
NownUVE/F3c0qjQhdMgz5UC5TOPWQdeAB/ZcsZJUfD/BQzk3jz1x31FsrNF8SCnMOYirD3NPjIek
G2bZpGcvtJ1Y6NPS835L1ZLvirYMg8L8PXPS8aAFVLJyPQbm7uvdN9vOHyyTEYUgHQy56br/3cS5
K9JwvFL1X13B6ToQU6nDhjzcfKH/ahk1bcxdaJj1U+ylKsoW64GOgCSEh8g9BbMd4ldJRneHNC9u
6Caw+KDZiqIT34Fo99jaEVBcmD/DwXFHQlmbz2a40QtFRutS/rnVdxQqiZqrA376B6bZpep8plBw
Z2uumebiPAfu6mfevId2lPlHcV4USzoiM7dM5QOODHay2LiFWoy4lRUmE6kTTIVzZjDeqi6IZwyd
M3ZIpZSKpKrYx5XNNdZQ1j/yr6qsjP68pT97xd4hLkyzjNjEQdU2lwLxO1Jkaj0BrhooyNbr4Egk
TK5P2DwvYQ90kGerLZEJqU6oemfYHhz1p9ejefHxNZLBW/S7Nd9Rd2LZdXR8Ua4J6BCDiXp6VoOO
/xYNeicMfQmEySK5CqevvFnSj0FhPrC7/6S89VOJxGrHGPwiJZjn0dpOCp27tjtORQPippwQrt3K
HZ4yZZKczVXmzbek6KGMcQ8eHQJ3QeM1Qlsq917RAxmN9cq2ur2MgstD5A035FDMyg0sjHcTIwta
EDWPSGd8LiYoLKPjfo6PWxDlc1k8TOZeLE4/05zpxaGVORVpxNjTXoBMbjIS5IWcGj+f6HGtUwqn
TjaVZ3tnkjXjX1h3xSwuIQoknus5XUqsux5XUvmFQQVph73hR7eKeDZOc7n2eckIbVlZV598ZPHD
1zgTOyG+wIXNylILBoRZfYb3oXsE2mNJWXvnCxga7leYn2LafPoSf4NXxLY12gbswmiOhbSDyN2M
0krgXzfOziPCgB4zxywrGglgLkrP+FngjN/Vxw6vsffwTYI7n/YH3pnym1ixIJMdJD7SRm5QkbIa
cLO5hsHRwPFRJ+v5GK2GGjoYbhev96d2k+ryUuXSwImUb5pUJGlgorTVVJwJ3qm0QKF05HinJvQt
SCNG2XlhuDkaZI+LgXIeWrXtxgP5UjlXvlZgN2Uv94unYjpBQiUcFLFYYgSYd/oWXNnuuy5J8fzx
T8QBzVlWiRbE9OYmnRxesRypoRaWVKVs8mrf57JSIfeBCmHcQXMmd9v0k2mOwCtZwLQHpL34u2Uo
YuXic58AkVe1anZLvjbG5ghup4uVCEXu1VwVwif915VGC6WPLdwK/tIzdj0eLdnifaHk15ycooHL
3UlOv8QXW6mPoNhHBiykCZ26eDJ6LGBK751WixzujK8qqH+oaynVth51i+iwlWqCY6l64kV+3Ab4
j16kAxe7JZNuX6b7veZrUisUJLmwzym2K9V3t+OA41WIEhDEEZQhVOeu+lxT7O2CwLY+hLSsqEkK
Q+TWrS8sPy0VQHD4LF8RWGveW4eJrr9pP+ab2OrtYS/U3d39NpuqMjLw416tXv8cRzD3UR3nPYNe
eWoehzgpAT2m/Msw4kX8mJCS3e4BidpA9Xg6ZOG2AOFbJUknYZPZN+1cT08azCas+1TULeGWfRUC
j6UxABIRCFP4Ry228aa36m84C8z9yHw5KpgLp0EDW0KnZDQ64VmD44I4pvZ+mef+nRwyjrhaYd/0
8gHWUNzBfD95Z+Qp9/kykEt1LzuVL/Dg++xjNcxvBz8iw4gxQY3nWzcHgO5fbxnjOGkmhRmQHEJ4
oTUxatAu5+zn5GRccZzdIkBCdQxbOAAo3+ewjQ6K/ahSKUXiugDq856gXTS4MNwngN/HI1gVAwt/
WVNI/D29xoSFpjsnsA2Uhk7V6JgRPlkSZ8DtdfcKLkE0r3C9gUOs4Se3rDPn0wi8oKCTx+PIjdAz
WVQKFAXvcdpajOatEMObewO5qId37B98TzILOqjbh/sGj24m/QIYZrThSgfpaaVw48V/tatMMO7m
oxJcT8VX2Ju0mWhs/binSe85g9c/VfR9anrrZQ4et+dv9W8JSevGc2MQDgIsZJcavfmNWIvkXzuY
B4le/xMyEjKQfeJE9rUSi4hrMZ6AUQZAw/phNXKEvpxMSA8bpl5se5k0hmauWeXKw2HqhUS9ffKY
8wuMNPAlCxD0P701jZCMDdsRwfSolJg373eICJNi8OVyx3hltVNB9Zq8Ya7RvPzlyiv+qxPYZGOp
21O+Rtk1mnSa3eP3mcHAlZ98b2gMk7p4ZxeIj0HPilLq4iQ8kxeXrYXRdMleTD8UjrGXXP6aoOPl
fsfVHy3hTo55vHQtc0Nirlb+JiGB2yic8ptGFyWYSGlBMqkcVegNOvRLU7MGcYqLgM86Wn/OT5zS
yXo8GgL7W4yIPrUxZfJh7uj2qZpPO7JJdRcv6Wglj4Uqd1iFK51Jew0CE4zYiPIFR4BKj6X67oT4
KYdTCICMBt5h/hNaqNK7wxgi5vFvMTy3XBcZHYlEoxjlBj2i8dtDB5morJy7OGt3vDDPs43/CTSK
FN5KjFWQRVHTInAd7GMCjgx1zY3gq3ge7o09WEDjNN7FZZ7QahvI6QApzYAGKUfZZb915CKSvATw
72ITec5O4Heo8EIsUun7Zi6w82/kgRhniukYS4E3GEl/9W7wA40b/fF/gFUipBlyl1jtPOMrEwzX
8+Z3EQ5oqckwjirwAAsnNjTFerpJ7HYWdlZR+YiJmFI7mSZUX0i2zX+DxjftVAWryIG31ZAyy09z
e/i+F2IxItxBbX9K/WmW2O6LHR0WTVybVREfxgcj2R9kjoDn9wVbw2G1sFpajDosv4HFIapA+WTu
luEVmXuAHphVJXwwYCwzzaXeloL29rbcYkDGuzD5bqrdqAKxEz+Tl393bPPO3MGJCVQP1v4sjHMm
1yO8XUO6Gq0StItJf6RcabnGxqabSozBowTL0F1NkaIcRqSbNwdYCUccFl7lJqU7kn9Qy8Tq3U3J
bUA12BYL+PEzdYT3P2V6/sRemc3NOTjukTV5QsP5MYJGxZa/qLXxMjRAUscgSJ14skZx5QC9TNZ1
Ehn146w7VlXYRbYd04YrERWo9XSlZgk2pQh1k9HlbGfb79apMcTrPoZCnWgS4+A/JpzE/yd0GYHv
alFxJM5c/zWIdsrMKZUSHLJklXUjA70/N+NSu+yctqdYo0arIa0A4a5UYYck9z5PnAqjAxfbXl+r
MLm/uU5JiQlJ51GrKOkeyrIbFiKTdykwUrjX5e9qK2l5Hm/KDcQJmZcuFf0z81obey66/h7bU8O7
Bn4F6xZX6iUSVINNywEf4B4CKLWtbHOXCdpLUGflhGb3iFNzOJI3ci8PmXeF7z6ytVtSMbM0cp+k
W153nrUKsNOEGKJB7FNflE/RZHyZIAttlzT3OHFd8Vl5CFHjm0ynTjfyZ1a8lJhxZwdvLZj7uLR1
nxAT0A52XSTlqP4SMdE10+wDXKwcz1GTrgtUqGDyPLcIiCQntCLUlkfi1tvRmcVSnwTibwSxaqch
8VBrW79IlTXn1OE+qGvwsICKCgS2362GyijcElLpK6KMAoK0rMPmYiYYjZGUIuJ2S1pWezKasf6L
mtvpKOXAiDIM1u3yExK5JaBhnA1mv/Zmv6MTrMOnXE5LBHHu2HDlrUrgCdd1qXx9hUQ78wN4W86j
dy7+o/fINPuHSwl6nNK9UXJ3GcwgRSxbvCU2Idv0AZRCwy2NIv+2WgF5uFpN6v0Lzr0aLE4rY54M
bmi7Vvd0HSLkd8z03RTJBbpXEBZmT/kySEy3ZQM6VbpzXC//thblojbw0g7L2yUjVEdBM4Bdfao6
1Dp7qznaubrfAbOev+zXCfb1B6oIUPvuQI+j1eBLfLPCI7Nh8N6ZDgnsrl9tdxxU8wCbUxzpANPa
kUe9rLh0Z83pnwmowd5vo5iBoYT6gTudVwFb+L8xy9tsFdOFmzDuE9T6i0EkzREqK6j6fkxAiiKt
+Im0DReJJgcqiYeY0KYSs81Iqkk1KM9eUCjgqGtOj3+CcPz8CWO2rjctbjRzCi4IdBcrZ8awweiC
2nw7/OdvYW/LhoKBUU0xDXUf2jntWZ9lVnl+pNyZnn+w3+Z2l0kjv3Dd9mrXIO71OSm1MiClgB9j
CFmm78ZUtF0FYoxJNApMi5mNOmGBp2j0O0rbEKtJ80qE+oMutmjDv5mVCqqpVPdXZTuHay6P5VZN
Iy7MPpl8Sus4WfFBkmqORLK8uJ9yQVq+81gMN4ijz2YxAg/nXrgvb1GeDkbQz3naUJUMFP3fYYGR
H/t4UtqjI5XMnkjgFmWZYTop4rFWxJyv8AAeCAsz03EvzC7tRDH6kjQ0Sb9TDmGaFVPV+Z7BHZN9
9EBB5I4BtSJXh1JS+PXV7eSgGp/ttD/KI/d4LbktfRBp6ydI6wEo2dNEJN7M7WNxw74k17kRLNmo
TSkgvURWjww5gYOUvUI1j7UbXpjSikBvPUZbGDBef7O6T2+Ijkm/05wvwGhUUlQsH6uL0HS1naeW
imklxnMQldCGfRWhXV2GC59PkEO0KoNRk4CVrLM2t/dWEyri3/fTXpsAtuWVM0EENYf//MWiN0Ch
k4rLF/NuhmLz72PDChUmhTfKi4ax30N+zqw5CqvbdwyPVaTY+Ar032ER9eboiNmGgK5hJmmu5h0+
GX9RpBr/0Em74CNWakrQADJnNFaf4KSIcy0IZ7RjPYksZ6dlTAEWb3svhJMddAGE6qkO8dFpKtHg
NhiFYMNYRI8FoZbCgH9J9rc56J8YWInWN1hW4c5kTWFMtwqpgOLmxS5OanDwsTtzhyiOU4YZm6Ov
vmxiOmnC7UPGxxC5TPXkGvHZUMLd3nv6Q+inCZmk1Vo5koFmYyXO//6qycPc/6DX5Xg286WdVnF9
WAtv0ZY3GNBMlLELWN1Gn/orDAwm9TNcT9Zyv17tnXxidQpkvWU+WJlAXXF/XJZpGx/SrDrqHppD
nFWjPpcsO60wohTXdyp8FRW600i5blHs4bnGEujY4snPU32jD0lbSIE4A1gOP3Qxx6eguGugx29M
kjbVVhBcV7TikZQscCLVwI+1xHE7dlhyu1in74mG/LJ+qq52u1wYNiH+3maOD6RmMUwhBG3ciyOI
HDFvbDXneZN8X0y8om1Yg7cdop+bq9eutAe0BuhXo813PjaEvaT2geVpPxyUmjalY7dR6Q06qUqn
B+nBWdx4RAxeYOhEiFa3VwIqKPaIZDlsrMb2Cq6SOjhcGPMCXKoCz7FDyJQCYn7i+/oSrsQdZKwh
OxH5mrtT63xMZNUPdYf07esd21X8owsMrRRSZsw8ajjN31qYkx2zj3L0+9nL/6U/P7SsZDityOvI
/RwyFGWHttH8oQkHB2QKAzllMCIqb2uHv5xsRYgDMIq07qcTybxn0KTMJ7w3hxErM9u04bQ18yCt
QMlgh4T56yHY8kXDXbjdKqJequDFqUa+RJwy7E8om3N25OFJm/cPvnfEQ55c/n/wJsQZvvOSYgcb
k4Wu4uah/QF3sa78CdwsJzmYmxG9OHDG4/UBu9eqmqS3lJNqzew6Nq/5OqQK4DwUDB6t4mR4hcq7
wXiK6+ku4A74MW2dONUlJ5pJTeMtKX9VHULknnKfelxtp3GXkeStR9bXtsWUSm+LuMJCQAlwy1Rc
RdFlV3xwRLUvcJ49fsUPGO9y2C+ZOyWDWwvce5xbprV+KLvNj9ruftTCYr12No1+mrEmFkAwGc9u
7JU7x1B3Rxy7/HK5J0G10mZ4jcMoC6sfFYJsHctcay0SeMlPL04KZ0Ck4CBqkD3QFrmIwZjlCWKA
pwOUVl7DCkEas9JVXl2RKyGnz+1lukVoMpqNfTj90zm752gZV1ckgswjntyUibCTcJECuTGufFkf
LbBdhkLp24EUs7Oo6MqScaTxKqkJlgzaAslxDf70T6r2Xyr0juHJG4XeOjuQvYvXG5/rOLr/T69h
zEHXNEsqqFbvMJ1QeTTIzC3vslmt5CdmMwrs7G19f1l4aFnCA4jahmJ13LtnOmYNYdmho1owVj60
UzBVb5p5gfve0GnSojEaO39EDTj8y3fgG7VoxxiNg2EuDofo3VnoKoOoOtH/kRREhn9skB9fwNKy
1tsKs7wA2pfnKEt0c/FB4EbtMenKrxK6L4n+1oaMpc4IZoWolIVCyjLNEXIWcPzZMm6T0FxpFu6X
1QHUL3b5AbcuCePqUlduMera9B/4vr+b6LPlcNYOmcp7SdwTuVG8X4CFUZ6ovr3BrRplJYwDsoa0
Zw7NgyoA6JbZNUu4MDzrO2np6iRuEEZHmn/T3MTpC8BI7TCGekLajDaIuDdX8RJHk1My/w503jCb
U8H0TATrH1JpfORQFJjLba3Ie3uOff+7LkzrG8yhKuFJPVfF19KgsTiLr5k68RqAHYZznGaTBLq/
ISkZAKurnMNSpusdi7tWsbp+E+MeBZI0gNfIgPrl6B4oJdMH5NIQ+RGqqnoBtpsLXYBUfmzKCuLN
Hhi+rAd0sbFOw5lYlIja3gvMzcMGvhMqwBPqk2c1jUwpZl2KJ3URc+vt1QCYyrNR7oGE/CwVJMVw
1GQpN/4Aa3DH6K5e8EvCMOHQBvgiJnkpUnE6Vj5cqDLhWOQcYo2mxS32nLX5FqJPyZmeJY6tURLX
yRA0Zgmc7PwLLrPOcIAWHHFNhj0H4Cv9SSS87IlPDcFXAfJB24Alhh4XM8vEXYTLLDPpfFKGiVFH
xX9A6ilsX0ZlGQfJIpPmavuzLRtAeXoEOnzPYiMYbc27kvnRRYeXSornu7yVhNtY/19Q44AdknJJ
2Dshd6/cpDggL27XNRKiuDCe8G4MnTT87usKnV/eQaofmliLibAxPQZHYDlN7QEonBSKedu25QHN
y/nlMe14zDXUdl6WcamCTfnLuLKCAUA5wKFARF4XRfe7Jgaj9tfJsEp24SnctPkwI4ln6yKxTEoV
trF0dWMfaWabh5uLlSUpT80DYczFB8fI1h7D3eXI5PxagxtX6TTT2OL540ZnAYPBwwyYx9R+eNtM
7jS4aDk4/dSegRl+1tIYbC6wn/JKP/wWdi8XM4f1rW5SELBhA3PhD0EvaYgm8neMrmkr+v7sQL75
21qToq9v1nM5h/M7sIc8YeSX0RCQBYbDWsfTt7E3JgpqnwPcRdZqLWLjHWD78jQc1QW0EAfOnkqf
RCcCKn9daXde+AKkvMjovON4Wt3ePnjozrJ9Off67J5oiyHFTiIVNTNdtfVAl71QB+ClnYAb3vJd
oYx5F+YodH1t8oYZy2zN2oM8uVRhhx6xpAlYWRbqVEHJM1OMceUzMgsBjmf7uV4X1raaHloOV3ys
umfp0Mg8jVJg4b+AzC/vH+PtRhLAwltGUArh4ZtiVU8sz+jUmpFcvpJ9qzCOjhDuc4jbQs8FMdKl
v1idtfDW4LhHlBjAAswnHNBXh6Rub+AIBvJr+O/N67bWuyRP+vWRY3gwNgWasBDSl7shOuOxDB0S
dXeh1BQpSQkXCykzDgYQ3Yj8jlfH0end1dY8qnzVdqaSTTMOdRvAX5JXevQo5ToxBKARWOEC1uk6
6ffAcuSRzdEDJmtL+UC0QHfjv9Qz0meFvavcjptnVbYorUOjKzVfEFMWrovD1xnPaLspmHnJ2omh
NmsS3BGQB+oR8DGonPsDad0mk2Tw/l8KbRhjGgD0TJXLnXUuy2sXirnVux/W67XKMBGcjMtBW1Pp
/dhfauKScDgXkllMKFam4Jc//vVX+sLBgtRqkEY7y3dxfiwbE3LHscRlRfYw4zZmA0rDm+PYFD3r
uec4qAytYdGAxDsrAHpqnAmOqyVtrD9KtG/dEO4r/VI+uOy7f3SpR2mE/luUmKiBQIHdZLAjvA0f
X/V0e126YNah/uNXE9fgfBE4K9hg6guW8xRg6+l2Xlsk0RCk8THu6ALj+MTE1X26o0UIZcBPd45m
zF6lSa+m0OS+AVjXqR9DVVpZW8vFOTiV/+1arUWQUM+II4Xxkf9HNKKKNgDS7vT04tdLDqjKSQz/
CSK9/6O/E7LHhgeBxL8ATE85IhVDheD33IT/bAXeByRfUNM8zPrezZpXFc8mPwQAucH2jXgCU2M5
JhGCA1lSTMVYRagOlQuDKt1qyKW30Ue4wEXnWxN0P0jpT2ndDdi1mri+ubHe1VqCveCyd0kbwbQh
4FyF+3YZ1E/8xSuXHqQqYdosc+bAP1Ep7+6kQEzxthHMSl7GSL54PqPgeeBCTjOSTrKKTu9w0fZf
h48+DfV0uIjOpWVwIbLiB4DZcRV44qKcKXZ3Ihesq1FIKOcSEeDLNwwEQMtfrB0jnDOSdOCba79E
NSz3PIxBvHR/iNEz2mlFPU5A164fHXdXs4zQ9cJllf+OZx1Ze9K49nKjiOnP5/LGmu6xyxwQ1d7a
+n3HoCE+A8HbVS5DPSV7P0Wig97pkVWhHH+EO/2kjlafVh5kMzLTcTo9b9g9gJg+0GTQc9QdlGpN
fMdI+VX08FajeiyGkN2Y6rSf8ivHR50IQ+FgKaIR04eMcSxCSRm0CX1purFKgzjwCuRLmCHCh6AZ
keJ5o5zFe15eFZZye5FeQgt0QPmYr8pU5VTzoH1TMnaEkCwXBXQfdRVCvKGyE4Ys2+4TkA3+U4j2
SVGII1mVdrX8u/nLM7gAivOAQTRXcSiNklnBKp57Do6hh//ZziD2D3TjcH6myIFo7sbMS3WVmBwF
+xl0w8kThhfs8rs5NNXS9lBNRsqRC6I+uiDapyiSlmBhKBhW3SmrCtoVSzUCN8kTKzc5c0lwOWvp
nI9y46A3hQ6L9gZChb72dzWuKHTddC+Fb7VlxipCXs/bef1ElDYoYALFRAjg/Od2rrCZkmB7a+GJ
Pm8nCeWfVmg4LsB56/ZJyR68n0qEutBZyoJbppGYisCxVwns1ObqKSakCEhFWjvTOtw1xZRV6Mrj
bnncdIOLx79d31jv4qMMD76ev5xFNU/5j4pNo81/QQzTDeRgg9XFkPOdRpxg1WDlgr4rECCxfcJ5
mSz0zOga8tS2nsym4nvdt2Eedm16KpyYe4fDS9VanX4gXWJ91kavp5WV5S5tv2p0WTp+Ntn+ZySL
hekragBjBNJHTxRUhA2l988nZL/47hD5xNJtW4zz25KDWOUAiMlGFC1pFdapWQsy6kOOgmVCBx3K
B7RTsFO9tmNcE4YWddtmpMRSgsXNiKaUIy2qcuKiIO3sGv9H/xmH5LtW4F8Kz6i5qA9IKt2cUyF1
bJ09VhP9lthKTp8dTpgQ+w1RWoWSB3wp4X4iXaErJfyFkpPWZsUQVKkpklZssOI2Zl7+4OntY7wn
6GNWEb+ZQ8dHWNk7hRnTeSvgfH4SG3ZrLD8L/OJL/zlZpqHSMNdOm3exxC6I5RQw7zhQ1gvwMTRW
kOG9+BNLUOuGJtAB3CIZbphl37aOyilU9//sxFEIwZ4vKyAhuXaXdWHm0tAm1EgcIHGKldVKbML1
zxmbzaQ9m3ehtKD81JocitTqf2sjF80oOa6e3MlVyf7G1d1TKxxjiVeXI1lH1fioi7v07Et6SWXP
8qZhCPzhCpaMe2e5w6Pn1C4t0VpW3Hv85kLePQsYM/gZDkDmgoJ0ZaN9K/Y8mPouQmCd36KLKjXq
YcGDm7SeZV5lXJCE7626m6Y1+HT6C7W/GPPsRN6AzYsTvaUSRmfxgnP8zRhbgV6fZHEQkGTouhfi
g2sNo5egI7LEUL87f1kcACGMJyA+u9HmNqNaxf00W4NHiPeGeCqhuuTX+zCcBYAPFt5BMOMasFxB
X/LEV+U7/ek/BeittumpM0FTDp9SRr//b1ZPgLaYicmfXu8fEkFdLeakO+xjaUJ64syWMSOBFmrk
lqt1pI6Zv4B0CE69sC2maAV3ZUvG3o4n3e5QxreXBU9BBSDTxTC81WfEkLtU13+2Ggwir98F2wLI
38yQx2ezVpN5DHyMxEN7fgWSLQElstX4B3gvRqNOGnSvEH6jWl2jAg8JNO3dsOfb37WRI0N5U6r0
RVKKBc557VQVMpbFvWbAAPx3KF5ZruiocBE+5xzhPsiFzyVHtr2YtKtKU3vDHCeKoN6gGCfMMFsB
7x5eEMUjXfc2wk2lRhOr9LZYCCZxtSO7jyESKfSh4nkwq87lX9zIer5huzRipNCYomJEU2sBd2bM
6pbXkrEvQkszck2QrKefMTE86qyDhuoGvSJQMPnWxghVg7kgBWbci5G46HzII4WWXexcJ3rYkrAw
9ygI+FhEV2qlADz+oWIRfyG63xEYiZLMF8TbW2krCrU1pHUB26S8TBat1DrE6Art+ws/4rXDJtUQ
UZnzjBioGuRpAwDQDLmv8XzPWsU3JtS2WAsbNET8a76y6tfXDukBEDI1DUazyhvxJztQQsl7J7fY
RO+Dy/ER+hJ2t5LWSYYQWMF8F0gnodqEBnU8W0e/rJvpeF5t0eMRj6iH+hPN/h80bOS4NFeOHeuy
Z9/yyYy5ynjOdAQVaUR78wK/XMH4a4FHlgJjnpaGR8AYRj4KENVJrwCIrblMVKCo7Sg8q2CLiLdp
HbmYaFEaFHf1t1qW7gxeXMxEGfVRjkddZLtexfP0eUSOXMLi205CazbbgxLAb4xvLVYp4a+KZfnW
Y/QOMWS9rtcypi5s+Bzy61vZVYBqqhK7Vgw7Yjr1VGj8eH4RDWvonhfTLjLcOmM9kKI7MTxwic7k
9TGu+Xq4gZDjQc5OW9gXe2OZ2WQzIqwgw5Y8sufTkq53hwg/n+HuLVpKkXtVAgks5vaIErmWpGXa
9sVibDPIsskMtj97pgOb2nij6DYebc59DmAVA3CfMWW9ZkaVQ/5ClWE8BmZf5QOeP7eXZrbBLKXj
JKirmK0887R6vGSSbn58bSEa+hSoxbqNBhdmN13RssNX32Cbds+JJ40+1Isuuyvb9evzBg9FAQhu
jCQ6W59OhgfrJVRgAxO6LHu8oMVTM7bLYFRxaw13Hq/IunmgKnhoQz6SlfKmo2z84w11hvqeNS+O
TV0K0ubD0YQY+w+JCmtIf0ztwEMFKSxxtRTWALQ63MM+pP8JLtQkIBGE2Sz8uhcAZOZIh9+iv78W
+tORdzEJ5K0Y77/uDTHa/q/N+bVRuLZPYtWzTBzthMQtJ5QhTlNIFcHtB+dMNR8f+0jSndB6nWk3
FtAq9/G0KyKKVNhiW0PVHy1yvn8yjk/J8o/0s28p3WXvMi2ldDWp9PpBM+PkiG9fx8tJmYrN11Q+
tQfR/dpdBaQf2j3CN9r/hXH5SD586gfCQAiyMFES5EgLtp30tu8kviC9ERLdtKqrbNxBK3uLbwcQ
gAI5LeHsnhnKLSE6UzxXGeTy4+PaZq5X3EpG3oVM7xfABAh3prRapuJT5QNGhojHzAia29x0JTF4
ab/SBPuN+07mALOAX0is1rT6xKmqsCHWc5b1dcD79FZ5qs2YteKDxXhUPaui1YEmNB7xTdbTLqtS
NY6F+gREIO41GG17OpuzZfKNaUx2q0SMCFIssv04do+sy7kLhbCT9wXedDq1UrQwQs3QtRzSSgO7
xcyZzcg4mnI4NJMgLt/qtsimoEZsN/MGu6JJw7McJZ7B6QKqlEo/q8c9/RK6oqSgkq0sj2nWZRzk
qud5xYEdcU3+hXtaD0Jt+HPH+BHY9g70J+GWOdtPBVZfx4JszlUNQnl00XAdGmHoLS8F2KotB98r
0cbKz9iWbahvt+kfkpImzAbU6XPcRsU3rJ6HJwBupOVbnprlVeD2zVCjgwgvq5HDyqtPJGWGoMGa
alx/B7Pj8A1vyiLExUBn8+nl5z5jml0yNsaJ+cTsK9r0VrH/PaHqgVGzef9ZCZKk8F5hIGiivYD7
bISU1RMutbnHVDdMEXP2Uo83TwmVF3KVtRrEdRZgQf4ksCpJE7sQuuSP31kIVN1fkXlcwmgsm5DN
t7XruP2GGMjTUC+dkJIvkJNngdUcXEUrgpoJpWuxDyLrpotzx36gWgRl7U9NUurpHVRq9o0UflON
NryF7vAGkQqcjGOqQeHw4Gmz4HpKyQHFXfoQ5HXKH21PGa1Cm/bJ4sV90w/0mqWcubUBWXX4UzGL
7QbJiKBYxNcV+IrbXKDQnRajK7lBm1nfx/4NFOi4axMpJOib6qsy+0oNoehYQZZqshZ7yHn/Hnjz
Gd6Tv/pfy8qKrY43raKKs/BlhnI5Y82YLCxxZMCUf288F1wlznpNsg8VYJQvWs+2IfE7SGw+Y2Yb
WEOJJEmQpOW6EWn5oA0C8JnKRFgDaUlAv2pPYpAHJmQYDBAmZuAjjiD3407G8rQtGoNbex+HHLk5
+WJUT4VCXXZMHnWSkMFP7O3A/dFTupzpij9kvu0msVPMq4RpAqSOuiHD0e5/SXjA/c4lsTYGGHIJ
9WlpMmAiwjlQAwKkxr2gQiCZxLcqeVDobb3O/OmrDSyYMNNWj5pbNN7yS4SJeSukk3DpnE+pgwPB
NEWjsw7EXE9VjqJHysUPnQ5W4xFIWLDAsXjTFzoWawhBripKtrKbIFrRNgDg8NAPkPOvw4gOFboM
CFvO5gWHFTzUCEmvmEmhNHVjCzkZBD8sOEHyst2R6SemV1L9TqgaBhjOU/M+Vbsi9qWcfWwPh5aZ
EHdZh4ZtY+gfqt/ezNRwFAnAb/7oqbzdWQ5U86rPVUvJUSMc0AMlA6jcXZIntZonXCbLW452NZDh
Q1LSN3PUmdDKGJeJcgq9OJ2+MnJ7QwbFbZtZd9j4SD7QWBBQyfVPJFgI1IneEwDDAXXpQ8KrVdjX
cfLIBP3xKbuWKXW92tpOI10bPD4h99MaHJRRwqfULit8UySm7mtQK6srsQgryytIlWbNmLvLbgxp
PKuYpf7+37K1tQXhjFqqW2yqCauSZeaMnBp6THXC4koYq3j+Qj4mWedw0Djl5FVV/VwJRMqWxtsZ
h0Jh2tmdHllN/19iogQkkLpUSkz4U03AzZPw7PwMWOUg2qYIBfvOOswE9dilkdvUAmZC/p8VcFAd
wI5vZU0lxHUBCQkQeqR8FtncLCBabP1unnK49BxVkt6xC0RtGMGI52qvAvtI9TgxOpTfGoV+FS75
ND32WL+adQmRK724A6NvkbmUzFfF0LtWRdmUSA4jStoz8lRAgjXNKDkHbDaI2UimrH8dz6zylgLq
SIcN0LvyeLQmmZ/JeoXnc7wyARdTQjTc+w9shDAGcSFMCrajbzWq8al3/74K6lHhXQLbRa0s/KFR
ovEkfBglqSUcS2Zok8hzErDGBSt+L0noUOC2LaxtSOiatAZhsUOadQoaZL4AcAr00FM7UD/5If3A
K1qqunoCjTewbD+Ryk2+Sz1ev8e45NbIxn/ssWuguxHvweVUR8z2zsaiVV/WtpxzyUC95Ji6Uxd/
CbbyktSFndBDxsLcnlMTZjs8O5WI5hsxWwe6jrlyr3Qq3HXcqu3NNvJH12NNEWiroj32QhGtFFBT
pQKysV9+5VsgqCvrans72hz88Idqg/daQHSIC3sTsA33nqEFGQpIOyZDvZIpfCSI6Nqr1CTMhF0G
FAWbtN6agEp74KiTyisb0PJG7M6c6Ye58fsT8QIGDYuYb+1OsE4K4aANP4nt2nRBuySjnqKUVwc7
v7FQdHa3SeZOGstO6+9Gi7A2vxnr/ccpeKY8ehELeql2aPgugi79YIuf20UKDEgelDVwStVOTTEC
lPcBDLBqaG96QrAigbyvLgGYvoAqmOSF77Rq3ARKNB5ktIaWxPFvQ3QKbthgVyzFzqj/rVG/VWYN
jICDnzwPPQ2lZCZdl9bfnG7qr31T0s6ynS0B/Wttg0XtEm+Nw7eY7Q1RTaeDjeZFrRfcaNwYYVYM
QMrx1ZSI9fQ3k0rpPRO1aKtvLRCI1bwhe/+yu+5MpSMcPaOkaCPknbeT50wuJtcS4eg6JFXkaAWp
WeoAFoKcJ+6QD9nG5cO/hVKBgskcSwxtQiPCFSxlAG6PXwHG6SVyKZSt+GPYKwBBchNBB66Mvr40
wXIZJUFm65aLo+EKWsbXEOKkspcRfMu5w9VSvb22/YTFNF8Rd5EF1bstdDzsLuELKeDSLueDftCh
xwXwU2RNjKKzGPGZyWKjwNLABd/FR3x3A0pfR5y25ptZp4BX4mAxs4o7htHVEyW+Ja/kgIzbOjjc
yOUiLRh51HviBdPEcyix7joJp76jgIZKkXArRrB2janSxtZuO9nCIqmvfu7xpISCawiSjLG06ICj
NiPiNe1lTL4YeMdyUZxMnxXigLVlqQ/HiASb15/dI2Ygg+U6Ri2iCxF25aIv+wzRcddR/eqZzom3
Z4wR8YJLlcnsLlMHJ3XEZ88VmRqyidZ19O+jCacfmiZq8Iyb1fo7tm6iYrskbzNFRYWgbDyf+fz/
Z3SutD7MaM72CE47FRwlI4P9kgpWs+A/y9k09bY7MixSObxhzH3325//pF7MAIy1qHeFIlKldSiy
BGC9XpALJ84eBdGjXDyRSEeOHDXxNGw2xlW1caC83P3ZIkAZz3rmslRYlJj/BTOOx/XSOEFmKI++
TtmuyCj4sJRIcDnSUhv8DRLLl3GrSgZ7t7aN9IpHI4b4/DhaDaGrbrdRowmVTNLnF4mpXJZGrJ0R
GmzxZFgFECfCZz1m4ebjXMTOpgJ+0rRe7Zex3MmrLGjx2H1MaH2fiivG5cosz4i5zeLyh8joZ7I8
zziwgdSTe8kNwFZU5F4wT9GxrZiQNYYIbIelhgWDjIxtQQyUrtcxtv/vS3AdEENBuAwbr8AyS1oI
MhpzJSlPqiMHAWMxN4dR0qkTfHZKc+3ZnWxtskiHuwMbFOTe1nvHtZI7gHe/UeLBVpmsai3CYy/1
jvYRB0gVDgr+MkGCT7RfyZNlV5wt7y33QVVVWZSHUJHk6T8Tm+AUiZO9dogoJ3OfGdd9tTZvjl0a
S/SBLlNtOdJpCqTj40ExsHEuwyHhH7FYx9Bc1YjykPec7hivBaCKvthBOq2OhwdzOqsyH7Tsq/Dz
jU9J2MG772TwDhoh91F3d2CwvHPrx2Au6GH7qQr0Vdt/lP9w1wgVU0k2C6L3Li0dXdnyFU9WnQFj
xtU3/5mkmLcBrUY+PZFcSFDuo/WYQRX65L0FUdg8MzW+aoaolNYAxpCysYyR0xh5oe4Mp0Oj5JP6
2bZBKiHc6Cs7HuQPOJmVk4D853mblMlcjufZaV79/fZyUvnMsXEMZTVJCctiZWGSGj8i7exBeJUx
L7kre9tE8Il5ylBlqon10oEmVNl6ttCDluW//1rGmjqZEZn3Owf2zxpOY77AcugTaTtNlvtKwWsD
jC9UASw3anz06aUjX2cL9q3Z55RsIVkIWdLIcSdO05CuApokVkg93gyin75h3moH8K0KHmbkmkji
4r3f+Ky0OSqTXinmZzwuUoOyUrgyUlQDpow+BAO58ziLM57xBb1ny0rHiatoS30TKUSqDFDFuF9j
Ehv03qFStSkIbMW3lATT0qz4Qa9OUfWqWrjUBgU+C/g4kJHdyFhIvxPYVXcR0YFxNg2winqYm3J/
YqarTajJg8IeWRyW3c8+G4P6h0Vu/7eT80+zypukrWiR4BBX/wGkklhd1kzH3d9IXXhy0LIrjljt
+Gd5KVcWBixvVItAWs/0zbRbaDRCkKgsqOjkugXPmNn8WXTVJ5u3iJ9V3kDuIlP2Qufb0aXWfu+g
2jbllLr/eII3VICSR3p9Vt5f7ImmdlOKZ3SQCK246L3yOUHK5xOvJbZWV9a432rat9uhrKNoed9+
NBtYOMAuTgQqhFSIuJUbKJWlY/wGvrYbkuGLtKPXLMYVTxMQGnnAlTDfGw1hnD0MhO4G2WUnrZ+D
ABNlfT11SQo2uesAIZFONrM3lOQ8t2edI7E/V7TqOb37ySaQrdmow4j4MqwTfwLThiDmtgA2AqCF
QnJAbTMbfOxGfMTTuPbs/IIa4cJDC9fojWybRO3WFlC/zqkJVJpMe8eTr0Eok0Os9mEtLP22gLbs
FlVJxRoKkzqIvGWwloxCF22Do87VeEA6qbbCr8H/xcJIv7Bb5H9ewK+dTD/ZARG7nZrXaXwYaU69
OAR0OeLeSXeTs0qtTdmO1/ga8+3WomBb8NoWtiwbeNZj9u/6RPXvjY1GUN+CuMPwhVcTxqsnmS0/
gQunI+O7WXlF+nMi3zX03ipw0Dvo2BMc2aH4WdqkifP0i/gCcWaBFRyNoTlQypO2GSqfNq8J1oag
DRFwR2rzwlnMCtETVLzTTIdRbx7yhfq7NEq/Fi4/6hD00oMZ3FCXKLjXXWqWdPxi4rFVk8neCdJ/
QUQXv3/A8nyYXN7aEu+4Ll3qPDP72K/UHAN5a4IhFgMVyFbdH3Wa891WJr0XkwYdjUcdKRkO7xmk
1usEEpNw9QCYEplN3QJ2MTk2ypoc+MBu1B704J1EHQVzwG1WTvTWEZXvuQIxNhCpzxELyLfTmFFj
Anb0MaZRUC6DB1Z9uSBORYuZu/QCZYtdiRoVeClOYH99qKl+J4PBJLwXTL5JeEfHFrEX5Ov5/W5s
aqGY/2urpEdVlWRrqJBF15EtemE94u1BwyHLOioyAuq3ebbXqSZX7XwRZf9KfYltTr5cxfJclzNB
p3x75omqBJ8GqWYSFMJmaoOnxfOox8GITS2BqxdMA+ckB/38Xc4JAFwpdQSebiI7UzVlAM2mjlrv
jWygElJdmpl6xG8VC4f+9MEJJy5Mv3HO16n4LaSBIqrrpZBYWMJquz0DycU5NKuAKx+WyT3ztnA/
QWcSL3RNDqVwpLTlPYGW1fh9aV4Q6mgSvE1T/rU6i4uiGVjzRG1dtHUhI8nppCZQdVzXY7BwAV6G
ZK0BM3ALmWdJmAOnFhUYIXnb9ZJir3edM0l7D+VMERBVaxBEBPE/vA28dN7RfUExtY/oNGtAOYtl
cBpXdlIBoL1Oi3nC+CEGMFut87KxRWQ3pfL7hD4UjM1ftv971wbbuc3WD2JqvhkZU3f+5RSUK+EQ
lW3MalN1L+0cVzCHLzaw5GS4uPfYZSUMDtWfyKYSvaq3MhBr950K8vwhYuLPiuvas/hZxQi3+idP
uKFh1XdYfNJhh21bPY/H1BJJLA20HlHYnJ1PiGRsu+g4hv/RIqdvxhDcPA70/H/a7sSHKePqeA5q
CBEj8lfD4ywnxkmEv8gKwCG9GbgT9ztNqbqtdWk2JbM/0JqEBqJioi4lJQpuxi1XoABTDfc3HOIq
Sr9FjbYUa+6gmI+4kLdEjAIv0ZTnaBTG0lj5UAjiUyoZNCC8ntQT0/cNr4orXQKo5ingYeo0eWUw
mwUZrcEr8ERYz0rv8mNZes9Vo0mEjf1hCk9uLmcu30AE0htP/an4eU/hHPH5LkzFgzByFaN7hTyI
n5taX3Pd2ic9pOjWbkNjkvtXk9e3gzI84PhtO38vgxXcYwRlPr3zQwETQgE1nixuFjt3KUnKf2So
4uN5tlMp8nCzS84CmCC22Z0EoGnJRQMzfGIcVeJrA5hBCIx6j8M172tu5ugkHR9zcI36kNW33B8Q
AcGZWLaialUOhnG1148GXO2EPpHfJP8LZLyDvl3PdjzxJuBrRaub5PQS/kTWcQfbK6Ak5VT4sfEH
8Yt6Hlf08xoDapIb/ai9v7sI2slaX9PUdHxGiWDkXSlq1pZ94f8TQzs1QNbR+6yIlMCAqHjhSO1R
9rO7qPQSsWTm7trgveNk1JLR9N6kxXot4EV1cyMF+wB/s6zo+zK/StRmdekoC6R/nEZTW2bfCIJM
Dx1tYkOe000J9RL5d07zm3yukcx0/tXjlY9KBrKy5JUhSNUR/bD2arhp6d5OnJTiXSNM9aM/FMwD
Ew5BRLkY9qUC5yjJVxO6McF1cQZNVIJTDyXW2YXkqvbudeuQcZKGFCO/tyfjiTCxWe4+/HZBzo8E
5a7fgxS53y+5tjIf3mFGfyS7BVqTRxfcAQ30Y4SEx0g50OsM8PqVUnUnzSA6/37VCRz7naBw21QW
3Fzosvx+1xGOlKxrXLWepxPiEVq5YuhluFcDQFbl2NXTn8BzFO2llK5NhBsK6q+sf5dEoaxhFKbM
wBmMPfS0BFzVTN5+32FDZuJkauGIkL2vI3dnBRFkmZCeNRj8GcZzOjVjD4pDWCFNK73AQWWz99t2
WeDvRsgDSAkGzYF2Az6DspcJXRYGfcPP942DmbtnsvgqiDvenrXyxt9eGFSQiFnBRHfHzo41pq9D
/xyoW9TC++iId19Yfe5rkoDEpAGnz1vVbi0k2o07Ivx8uAS0aKiUuM6B++oITNWWCjO7j2UulvuP
2kVs7e44fQh0dnDEC60FXN2CXQPqkJ05K5ZWXW3dzQdE/qP71E5fqtRupuntwb2iH3s5uMLb2zxf
dqqyLypNmBPYsRdVbprQV8PxX9MxrGxr52oJmvUxI8cJFN+chGINStCp5snIMB5TZgrbJQzDfVcJ
f/KuFfedW2qdOv1OlZlEHqZRfhC3O8zasgZQaz93Bokdiyph1CtnhogC2WzUFT24tYlb6je05Erz
kru0h3YIWPkISiMUC8s8mAivCsbZaqu6zEtu0HzgFtia4Sp9Phrrua1nB8yjcBY8lVq5juwASEji
UBa2vMSTlWOBh2EAFcLaQ39Z1H7bwX/+ROFSC/c3NWVEgjFqN9RG1QQjQCfiXQoJ31VLyMSrADh7
5v34AtNLjv809eeDi0coSCMA4Dpcl/T9ICmj6EwlvxbkGKL8kgltyeS1MamjZWk440fwoMzEZ9iz
HsvrNUpmuH8pgX2nAlwbqxKstqCUzvPX4yzsNoIx8moI0/+4jSiGsgp6x16mFEvFJP6/MKB1d9PW
zqDYqe7jDSoyKPNClduETBVYN4c61CKy+gcjfu9hU+4z14yNcGfCNIFCZX9TMUDQDFweKVCJ/YLg
BreQMQZrt5N9FZdRNrXYudfY5FsFrW3Yozj8N6gtjkrwilz/a3Wt0F51NkJrK3yzFwk7KN6jl0W5
FN6IQiy5wPzV8HLjLq/afGQziAaWQbDBJ2859goOB5XL1CgQTp6JhYAKwntisZt4nukXh2Tmecef
KSDoLBEEmGZqrCQPNCUupYBVs18b7Nc1HE4ywZfGLblp1lzdIZihmi0pBEGaR9cGFN0RBq74Ugcg
4uRcC6ybnmAnn0ZXU7642yfKh0xpSmc+2eQzx24jiDe0Oz7ampY2bhrjEkbBFZQW+XjVn+jS2af9
sQYuaWza7//72qDL7jz6f1rU2IGtsoZy001Vuottxp8s0X0qtMun1vw9DvM7A9groTS20mc718bg
3At/wk5cBKGkEtitAb4LDBJPEvI4UyeVGgatMBB3nz+HLGEbKPa/oNrOwp6qTaQ9MkM8zSA5rotI
JiuGi2Lq4QIR2I9afOLjEX5zlZsQthMwDtfOzPFZVdXJk3Vy5Fza8QA5G51shOVDshKqZLGrvBVM
ol9LqSkmpa1fOn+V4acMiWH+6PfJnK9UQ8VoAoi3bzbmZKT77HCIBzvct9WLqrVTqoXnzI+gTosl
RrogcMMC2Pu7iOqZ0cNy9fj2/QBllGu4y2YjgcyjgcfmKYG5N0LAx+wcOgSM3kKyH2kGzSCNjDYj
GHMtCdyNQ9JUCKLhWnwIyneVBpGGTkf64RrW3LK3mB53Ue9hQDa9eNkxAyOdT0rqTeWykYtoUFWU
XFPCquMf5QvolJDmKUAGE1QVxwdGPpHfrFbunOkmCmkYojfiB0+JJagSNPBBdS8TZb6Wrvwex/nS
fqifZP14Z0E+HpTrcA62O2c+JlPsKr1TmzNqKiEuSVfMosiMRJHHBpOsC3BmGpobXZ4eevdezwxm
JWFxf45fmQDJ78+jUS5mTRxTrLyAVxc01X9QM+dkLUXjZC0eVy44WsAi1JUrPxUF3CdTzfOg95yZ
mxdd/LmwNPClK27lKKTuUNtLlG2tVYJBFfRycyqgzNfBuMQuFObb3QLRA/F1a/wBQDu3pGhaHeMH
kMwvUfIUvtwKiSwybghCc9zgKBNFXTRdERAttNaTofVqyMla9i9FyZgNC3rjfLSX6He2Ou2axHtG
6XN5heg6FbI331fNJ9/mkAgYo5S264h++9hSm6w/H26KHPEtmWKrRGmxChHb9PJoK/LXBHiDJwjj
xzkKDtppAoObgKVWa4yBedA8n4R9tgH8t6M0De1qMU648ADYUgp7lBG/I6kvMm9qL4k+ZxrzeBa6
sqs2bC2gJaWQB1LHz778Vo8iKEZv4sfjt/GR5Y7rhF4fIfCYnrkOVja6abzs+BLuZURTQpb6vU0g
15ACHXAvgxaOg2ORbqBlz/0Yv0zKSNKbUaJSjT2uZpzCX2rc+N37ln3WMFE8gqmnrtnqWdlp3u1Q
oG5UlCMwPV0hbhuDXCRN8Mw8MVc6NCOt2qUkdhFmdgsPx18D+TxZknN7U2F+5K23Z3S6/SHX1abA
yjJqPgNQmQCxyVnoSkhen760mm/v4SKFgBSROMWTXNF9HfDtj4SZDyYiRCaqgmTcQzFyZ6hfKs2G
9BP4QwjM682qw49h5Qmu7NkN8yuO8Th3CkzobFX5vaKRQmeCeXVIL9eh3pxxkt+QP1xT9yATjwzI
XIoajOlJMr0vxaFHvCBFh009ws53YoFeJfjrAsC+1TsXbs5omJ25KTrt7f+5+O1fDK2ubffvdw6s
IdQpaJLFG8SrAYRxgDb34VtJsScyagCN9u9uC2ySesgp3dwxpjRihzduAJC58Elfkz51jawoG1Ry
eD7Bf1OWPNKG4J13RSHKWhdg8UOHHqCAntMVhxoxaAfw17Uf/JbrsDidAkQSYqgjO9v0U9g49ToV
Y5xC4kyhvlqGx1Df0W9i4uaiurz5ZsoXVW2BEWAIbDn9PaBNwDoX1eukTEY7NjMur/bGXlPk+PkX
PgLuPS6izlNfcK6QKqcJ5yM8aBAxnIIq7e5eHaPXx9hkoVwwChGIC+9UbPRmzqaK5FQuLL3Mr97H
fAjt3MkbazDxKPQZ6wRch5YRfF5pebMp+zADT2kDiiFLMJo9gFZpa9gnWtMBMrXZat3rdzS1L/bB
7/4Ymv9CPY0tPe9EfaGra13eJq36DdjYyZQOaTKJYY9OwrrnQnqh7NZwbchDG7rp/ybskBKSketK
aZcXt/vDzWhHmg76QClH2ZCcUhIFcCd2RC1iH21zre717wJKWKUmILwkjdl3/Ytjzj6U0HqsIkJF
xXde3yfa6kiDanjPOpqaSDbrF9jo7FtRE+wczEwkptU9/CXtKOv/koz3YrUgo5Ot+obqLCT9KKvS
zLC0Nf1QJMWyTz/tOa2VGwT9De8jVKNbjccu7H6jOuqhcr9xfjgV2gSOLznkcEhAxkQIponZjwx1
yJAiCZlF/NAhEGV6Ld3kd1PmtxSk21T8Zf5EoGerv70ZP3cp8HsQDfrCK+vJnAJKy9W0TjoqiUZJ
O6JwFNc4nAqoRfXPtpRDI79vhK3WstVExwHoKbfIJKjfGUr+h3F7lYhyIQKXebDkiR8QRvE/guaJ
VQDrkkKd4MPYZpWtsgljBcad4uAiBwaMHk0IREsQ4f3/YsQE6SnhLdpJdDXXnYIK5PAJnqc97N0g
Dwv6xvc/ILRdHXdiztDkO0P8kdgviLGU+0MpIa2Cdu8Au9kWcapAZXgHf2d3u9rehrpibhx5KaoT
5sC6UZ8boGKGvC3gLoSwsG4pu33LApqdUbrgKMQIFvP03rpjOtGwVfSPVIZBNKtLHwiGrVacybMG
o4HtQ9s6YPZPi7OwZESDSrPlz0uabvS6jrt8Y+D2f4MwpsTM/Ct9LgexqOLgawI7aUY0U0YS2zLf
OIWvNDq8cjGTHYB+RjNewf6at885xBXkAOPX2JWHM91m6z5mX+pZEUHf4hLIff57Leuv6UklShtt
oLnhf+gH0xBFGtQ8D7hgoQ7UAZvt8wqPkrtO4RrmoZxRMidzZIzXuQw+itDdUxNDeA/s7lw989H/
vD+DrCXcTsfCTeua9FEiurJM7BSTElFcs7DE5AakNkrStO0FRUsmGLiNI1b1SimIzocirxJio+aE
uULOcS47W6vEP3XGEES7TgH+pG7DEh8UDfGk9bioYw7cjl7c3zoWn7qz3km0S02q90+SAIHx91J1
IackbyvdCz9ejRWOfNvegY5HLXJedqkftOjaQ6qCGimHTRfu461NCpbWYj40YSghUkATv9KnFlx/
orpgR7TckcY2201r4BKIeVKPCHN6/qvzj2+SnFh73BLTUNS22vkEN6QQiQY2ayb3t9JBT+dQpgMy
f4dDq6BX3TF4aCM/CyjHli/B1dbUnV8A8kDBA05ITKKtiUaYraU17AdOX4cTSiUMlsiqibWYlggL
Gvr1B1Lrzkc00IVMHE8OmwwWGo+N2jdAQIjRy5oRlNqt3uMjx4S+tFcqsmrnE8SJh2f4Aem+DM+V
l3pcC2Xuq7Xs3hkoCMZpx2d8U7lZgf+duxSLxkHSS/mzIfTfvy3NAeo8Ro+AJWZbaVgf99PJoX7V
FGc42/nNnLvtg9RaBL9OQ6soxbgKKBU2glXI1ALFlVPrvXTJLH4poRPOd2uhn7JJHAzNOLfFoosm
rQBD5DjGttz5Yb+iRaizB+RSJD0CIePVtBwOBluGoeOhe6KFqOTNBaLjVJzSuXwZ5JpGqFppNcm/
/+qw4GdnTTFIoRr8H/msRoYEGcXgSyRXbZGaHyzhR55TATU2EV+fel6QL3yA2RigheeZ2Wg+OzXX
0kzPvxP1Hij/4sd0d5L1ObBBZdeAO6Tt+tAxUOAu5SIdSVcsmhwwBUCafUaRNwdZaHikmQSMqo82
oaGnwUluALsZqZm1+1k3pu015bdSitewh4GNjZL63OPt9JWohip5Dd1K2LbdauGCSC6ySM90O0Ep
2ArgB422SJJ+av5HgPjA2vERXZOoXJ4cuqWKgIvKHRwsQdvJw9f/iBxCHqukpBGDo7X4BwkmlK+3
X9J+5qqqzdcg3bCiH7AAWtdgV76K55LAFI/XuAKnvCBihUThamXNg4bcMaX8Ux5+dHuMyccppN6A
HUZUo/gnrJMUd2uPX9pITkzwkrL1jJpPO4hian5JFDZPQVEqqnjkCh0W0zfuFLCbDApTg2lRRzY7
/F8MzWxOhjBm1VbI6eySytkzETpOc9wsBNnusV9r6Dy3QAfgPtl0VvS+3jgsAMW0vXxvwUhrmFAX
7eatNSPb2qH4pTDbu57mLNgosZ4nEJerabaN707znBl6Ws9Ad1KkLS9vWzMsGPVkeb68U5p5Ke3A
+oS0iJvI1Vq9xg4jlVrWfbbP3VvsdcWG7Nd0abPhjrsOAynboQSfjD/4+kb+V3/cBqZMUBJO9lyr
AoOrco1P9LxcjHz/Ze4YJsLxwPlid1YZ/6mlG1y/HMvBpDx3uTN5tiN4d8+g7KndoFcfBkvqXcfd
IqM6uas243NSLAyv3QIZ7bkV/IkNYWZ4O0sxP4Yjv/MLh5RjC1nSg7lPsxcW+0G/mgcRjuWyEngb
XdYRXxSkEx+C4M0Fkn1IT7d3gi8r0thvpaEcjjrCaVj55D8vaAYg//winVxeYhldcT7weA2wm8a3
eLFdwQDfiRtB6+jds1C0/43SWNxRIKujW7voE2h4diZg6Ss3KHu+kkmlGRnRc7w/WPyehyePRQRu
DAOXi43ehtrw1RYBqGAikof0zVB5KzNPyR3nCBgRH87jyum4eOKas89URJPDfWqTB8/VstppvAAq
EAJEBcCLmtQUiVq7AXRyMqbtXH7thSaGA+2OLuvYP4sWb7H7dsQ7UNRWTSKDScHfcxC6p5y7821y
0PazJIX37F0/oU0RiFJzSNxhCcovJzU00d4w0u+BKF79pftFI2OhO5dL7mFTCklKi6iAOSbC0EA9
olDJasse/JjsktLv5aumwHjRBImnaCL3x5n9Ladb1el/xpfwIkGLp/pNjANUjXbS9pcCdv902q1h
FSA/kiuvgMl6FaTrt52I6N81FMDxKYySp9deOglfsQuVjIimI1pNe+IXjhCH5V0DgHazviggUwaM
jhVu5ZYOXBk3gQm+Rr9Qhqvs0wUG8Vv8X9LeobvsRzd03RUntd+BaWPVHyPF/EElsG+e0De4wtar
IYnAB85fv5o3Zn8XYg6Zb7cnccnrsELna4Fh4Y3gVpl2JW5v+njwb13fzXFfHJUUzbcYEAhHk53F
yo5DkzZmPHm4OS1n8MoD8DY/XvlgFsT50O6qK6RgjNog3KG0bwDPSouIfh2oYs9tQ9uy6tsKKooW
nxCBfwVvv6stujFyrT7H6mMNDrCMiMqynwPBoKV8ffXcNVZk1OTh+fN+2Gs30dbnvnTOJbKvZB8d
3Qvf5uvBcws5kak/KhsBoPdRo3upNPVMf4OM0pRmOJUBq65mCwKyzuE52EPsf3/bXvxOAzAGlovO
na8fJdwo2I1Dx7so4jQHzKhZGYdG2hDX3D4XFUku0mCMSvpwfkb40Rr/kEEHOI4ElAG3mrDez8Nt
N6eIHIJYM1jMsLyi0MdvesHOaO8uDiRlOC+fqfQE/6OPZ6skckWPRNP89YRi73NAyxICgEwAvYr6
q6WXON6NhvmD3j5RSKhMARwi787HoTnynecvyDRYUUVQ86IWo4AW8OYOck6MHQ3mKX8v5TcIicFU
4QReQaZa30dXjylwdgq3lvMh9y3olkv7vB37PLsm0c2cROh1WfMN6suuUQFmshk+XxFvUwPdaFAP
WyeI8sq0x8YXc8bsaXrPRMn2qK4OX8nSOk/s9spMyn99KGE2idz7WE9NnzwM6OcqvywfwFG9JNfM
QuAwsXaaAQVGD5NGGzGr+khCyBh8Slqe4aRNvF1sCgcmIL4/nDfrqanpGqiJTeCcVXKgVIxWBnCD
rQZHhqTie1ZsHKt0SjNV4nipQG9/WBAqOFSGKGsRJpkKr3hTiGtKEDXdv2XZ/KTTgGGSHIjcoRHq
0eLsEOwekTmY2QC0svluCdX0KlN0HE5UWbKJ2+LINHKeE4P6/cmdLcHt7jcnp+Un75Wmm0qhZ7lg
KJI9CqjMqWDFCWPfmn/FxAUFwznTCbsKdgwgESQ1VENhqr9OAWvDYzBdkqec3ntDZ20ffhyYI+O4
sXDFRz/QOWs/EMoe5T3TJD6lwzM79c35IZDrl+h4+W5jNh3m8e06W9h/W3LpEBicK1s8mlu1EhIZ
ryrYEYx4FG2szKnITWpVvCnyz32w+tB2deNQqg2Nlc/8gqww38fldVaT2AhAloLB2nH0iyJ2ttGe
M+yDACtBnFDjbnrZl4Xyy8bb17CR6no2i8z1Xt9oUty2mNxhPuP+luFy74Q0y6siOM/6aBEK6HrC
8Y8ofrDK8sMx7b8odeWFZn2S2hExkizhgriN1rsR7vC6/GE2UBApW+Uf+PTFy3PFdHkix5rHoRWi
gG3t3XXeChPCdoq+ESt2EPkOvwtDg0AHLjXJqZBHw72tI/EhR4VlCDYxPTw1olXKJ9xr5IvzJc7e
k9Vpm9jR4knrVEk6Vq1EgvI/oBM5hklw1aunXVk4xTsKFHjUg+IriMbjUGsiZYdsH28D4Q5f0si/
O3Ejn6O4Qi358a39lxprUikURgqQpFId+uXWQrAYQ3OplanOQPrN0llAh/7f5bvIoQlTW1ZLOdrY
Mg/VvdajrG8yud+0OL/g7FmtBnAuCz09n6ix8CBNjgXw6kfW0Y3tvo7FQNHNZOmBaMsvz4tRx5l1
L+cFoOZ7d14vg1hIJyy8t1887knzq+WCrEOgLUSFQOpJ8jBEMK5xenuLZBm/bjceVEp3I5T65l9t
eF/nmhJH58yNkQJ9YR1jX2X6Z9Rl7h8mXFoDWmEMyBgLgo4Rcvwf4kJeBcOEJbhaZYs/766cwV2J
Rg9FfHkTHf0LKQwc3YdI5X6v083Pt3rYd/3VY9GSCTb3mb+AjhVm7wQcp5vErx4DvBYijTvrLBBJ
8+PHcqbp98orTdfdupETXkauA3R8ONR5C2/TCnQAgO1MHmWq+NbERidGiZrlaa1mq/fTbRglzlH4
iOIAehgWop2s8Y3JV8toPSkGO93+5foNtDrqTAoq0RMW4TQpktK819zP0n3JCl0NwbpdrAsScrnx
+DcEUwrmqpAG1pi/TNwW/EQzzxuhcQZr6A8z6LvFSeEmB5CWFCMxsjx9KwpiameB44KR5VMRMOJT
lFrdbM3VhAmCxg7YhLJsaUaayeTDLK9QElV7kCGJH5IkilF41HrvQj8her9bE5Apb4y7VGg1MaVy
5HGLX3CEtVp8UvpjeNRszKRNSWFHQ4XPNiS1/qqv8IEcGYa6ukTayRHZplke+EmA4GkwVz+RTG/D
g/RnprpLXz/o9NZeA6rc/E5xn9L7qZhphudOU+mY+4AUSQUYeZLubfjrQncgGphWSbPUCHhGpTbG
C3Z+Vj6BVBSF2Q0L9eHPAv8d26o2BSBmPRJp/YDSGaEYnZut6qmJ1Y7CLy+XT0Jepm5Trdu0ed2v
iJvdLXO7YtHUPqDJ82u84CK7bXlOlpZYIWSsu1Ucl0RcCyIG4qV/i2AxkJGaWyyFC2TeQGPOmiH8
Jb9wWPoCgUFVHpHJdrBTpXhtuvl0bAmg3X2pWzHw1oWLIuhzcPCRd1DMj+d7ShGGxcEme70jWrFw
hCZ4NC30bv+S3GVw1EnO6P8rMGl0kLPDwMP3uLHB2iOz47amF4qakMRTWtqwvutBd/bDYMEe9BNq
Q4TWCFIeuDFTwL9LsiVvNIkESPo/GHI0ZgbeDlqr/7IB0vZvSNXwzESrt1NhFYrUBlLrX2meyw4V
cLWXj59sM0kUbkRnfYfzfBtTCDajBljlqPH7J9iVQu9J0wNx++K3ggJvmAt4bBoYzBVB1a1+ejSh
7N3yOqQkdgzbyv01X/t+ObNy+gNMVXL+hj27ompvUtAoTQbh1+1oWzev0Fe2eWgmxfMovqlGH+hp
jR+tboHm1EVGcrIEmWI7E+kGgQxj6jzM3RWtcPLdRAE4+JNR012RLe43Uas9qt353bNnTAO0g0nJ
5RQLb/KDV8gqlh8J4OZa9vrt+RPGDjbrFy9fpDM6MMliW3d6C5x6Q0uiNzTrsF1k3VRsUaj+XVp/
sSvJbZc1WYDozsUkch8gniSeYPmiv6WAmsMN4R5JQoGnGfwdL/jCrdclYBxZqIB7bx7QvCcXwbkm
MttRGyjS927MKU1vdXgTZh07Fr7abcXSB8diFseo0evtcNeOJsxZnv/z342fddY3KYoc1vZwogBD
ErER6NerwRwoKc6S0nEr8Wd++yDr8HmjaEXr3hB5///JgTshZjlmrkW7O1ZsaX4c5tIG2e/kWWKD
5eS4z0tZNR17cBg/FLIV861RskD5J0BdYSrWhWgxrMFLtzYdP8HX9d5+HLnf0sgYX8f75mG+Y7ok
6Jw+NEdpZtKIDSTW/R/m1OT+8SD2BDWOw/QqGp6td369LGhisklMGytgqUDYq1RRAw1YCYRBMe+U
GwXr3ZuLOVD0y+ZXwbXYk6odHUlpyfR/cuTjIIsGXqOsZWKyIW2qaoQ5TY6O6qdNSRZvfjP7jnAn
Y3iCLUzz0aQvLuLdYE1lTF7m9JvMph0TuhVhbVYyVK8uU8PKF8VRMXfF9p257RDuPxND6zHh43al
2M/pMUOHtBk4uDf9MjrklnMeHzqzqEXeKKSSGntQrijtsNTD0dlHR7Ebrwyi8oay4WaCiaiKlps6
Rj0IxfR5V4AG9NxS3JWdXIBahkl/hy8SuQAmg2dcZoaPU67sPBZRGOzU8n4AZ8846Rxeq7xX/ngi
7V0zD1ANXyQwZYfJmAyJ40sY3pgfN8bjd9aISvM7zZTlYzQdWJQQik8GW/9x1PDF7kxQwjNwT0V5
U/xnbEqUtx47zlMux0Y1JOaDWm8GbpLPwzem5+0689f9dBcGYFJfUFZbyGR85W/wm6P2Gt/47war
zyCoLdUBLwpLs/6moGs66nkVz8PxHiEa4AoebqkrzWW4eBgQ9WmWxJ9AEKiRaBesLV0ppL+vUzcb
sQE3OPyBK0nk7/pnBMo0CpA+4GuvK/Z5DhNzl4wkPgCB+kaK+ufB9TQd1HU6/5J4OAN3PyefNx3q
c4p3ux+VErhHfscKDAvem/dRVXuvAmKLuI/2dsO9yCNkLARJTv+3Z07tmevbDfHZSqHVwJ8VZz8O
Jm4lSHC8hM2c0vjdk/uyfZ52ohtW5R21Q6Uqx+XEpsBk6z8286qDuxyzM78K5TMoric+wzbq9csY
fWc5U42F63JC4xF1pwcbVZeooJ+3TN3z4iimbCr54kzBfXSDNdeOBZAnr1p/XIWrM/oVmjIcHdDU
N33Yl6p2yprYVhogcOSxI65qjq9oK2Tt3vVJC2DT6N/uYxtSj9KYSrcw6Ewmc9YVjur3amIqf4AJ
s9vKBLMcx2PT0rvm7p22Md+COmodSCtHAkpbPTR1W5Z4iXS4FUtSF9U4hKr33Kkihwtbt4yX1w5E
W4GatNxsl7e+GwA+akmLUDAa0YXKGIaUTJ58/O7w+VbznCfQCRbJiLGjCO2wRJs5FrtfILl1y7TK
xk6YsXENxVpQSDtp+ZSWHjRCCRhH9HKqruOa78hUp3hpxKnf44mwDpiMvzXzDOFugge9e2t2VcQF
ldKEw1vkicX+NUI5pR29SRPY4yCCHycx0Imhw894H7cUbMDUOIexuLLVMC4mgpcg9vAFS23mYclm
kz+hxsoIC7CXTIy9nLlj7DXkOLrPKWL8JEKJfcaJCidWfi//auZGa4kMTK88v1tiNoq5xlD8wBPU
new0cwHB3Lg2Mi/D+Z1C0sptszYHFIjBmYYjxR6tT8jC+mJi8h1hi5oPi8P6Evmn29CHF88tLCvm
bRoSqIRcYKRS5j7CCtAt+r/m2bRxR9U5cy1buxyA70igXUchfYeZ40PAQMN+P2X76lu3NemYFmCa
EeUxZISoiryedEo7ST1bwT/+UZXg4sglGRxNhNw2NE32Bu2j5iOFThp5xegnUolsW17KfZZXL3UK
ugXdXpmw1sb13TPdKI6qc/2K0bvk35RnI2USCrXLwrLNHDNExuMm2QZr1NpJX90fkmR+VkU6o/X+
nB0P0mtgYyjixNTmdzTmeC01ozKhQj4MiROHFatSeSYGtawMW7yVSPH7GUKPjwhII97d2CJOZkK/
+d9n5nHQpBLF+MTj0DUAMd6ufHpSr5BLevEIG/+riZvjDL1PWJjSQgdRg7Q9KPwMRYNHE2s+Qo29
lGEU8VxSTbmB//NveUGRKHZE2Wwk0MZ57qelV5LFwYzpYHnQABHWvKz+AVhVw2HW8083pOMBvo+L
y5YbtAmPjgIH3wi1iPCBaJZ63RKUMKqLFRePPnOfi0A6KqJLLqY53lcIWvoC70l6bnQOzNcWCvtM
ue2+lmZWAZOExgEnGMgg2/A6oU/TEMrEcPy1v1/+xOZLeRYOH1KQ79zh282iDRHaofPSXYg5T6DD
i3bhUh8LWdKNydPIjnWtD6RGxXk4rN/quU9oTjMCYHGK0Nj8jOp1dxW6pYX8pYBBWlsoTu7Q88yr
GeCN4MkGAJc8L7kkGwqonwtN7RiNgkzwbz9EKYc6rGoBZYW5JDtMq99cPpCIVAOzXdyxWK0CRa0Z
Q83ZeOftICEBrER0LCOpuuR1MmCBHDhMsCsNAHT2/jvwRtMRBtqab0iaAbWpiXi0HxfaPJ31vg5n
aG+LEHpTmwYFuTu+Xs6EPFt+KcVuOIo7hH2vxktVrgKjEJTadEOLSpDK3jdQA1E09aTVKFEVQfkI
YaPvw+MSKXB7nWjfbI4s+OZDNJrD3fkkC/BaK/acp47IP8J0JIq72Fl0LBTCWeZq60H780gAmEJW
iz2dAEj0uRhjamHDAtO/7he4Inmlz7sbpEBlhSF3kTgLfjDRZERztGl7RkiAsMdbg7gYc1iVidBV
3UJkUWYSox5GAs7bnhVb8+JkhGEr9Ki1S4OBzsdm5I4kjdFya1IsVLnQF3nPs5mYFbsPQOpLGpuq
WO90d6nP7+Vb37Zg65O8dzOo98qq0MWDgyz4/ZGJcdBo7LuQtJz+xralNLw6ONQC/FQZeQgVDjmg
3/PXq2lStiN+RwD+g2seujVB89Hy+se/53rL+ZAnQVnSvomw48KZDiGrYytqA3axeFFkzHd4pIp8
bT/qaZrVDEiC5QVyaaMhG4RmvAiGHn2nnFkqBOGMV0hzrXAOMHnCvR6Sg+CG743fHwk5SxH2iitI
l0CsZYRgMTbjy0H8lzM+AMmTjWeMyBh1qvWmHAy4UXyYtqbr54L87fONbEzDRtDF2yRAzjBbQM+x
tUJ3rrCvO0rjX7mjIEeVV7496tEzX+//TEWJy8FSaueB+evSHENRyeOumFNnZlURyfj815UsS9SX
Ra63PYnkVuu9xPpKexJdkZwofXuGLYO8UaAJ2w/Xwa/cIKHpInMjy1/qaEFv9ULBnDNQxEZnU4hQ
M5CoZXpE8ess7eaV2vzrmpvt3pvEDAzm0KahmsRKOShz28UNQFKoLLDEeUPPIg/pm1PLgHB1XhJA
sLCXLVdDx96YA/L1rJLLZIOwrV81PRNqStdrrjdDNQmZPpmk62j+GtrhCuo4obgo7yZ2PRgzI8xh
cwmBLmq5z4QvfBb1CIHUODXq/W7AGt6nxUZtqqyHutTfWiY9JVYRnCOPCoDLefCB9dMeznJubKXs
PtCmSc8IYxVOR2tkpIKKopXUFR8yHzqSWcgO/KIKxsbRfAkPSwVgnZDCC2wyRs3HMdo27a9+rscd
0iojbbtwVuTxh7nJACFMt2cBIweguDCc67qTZCtYn+n+kv+UYAYhKzxx5ME0QIyczgsFbG9aebfG
znNQU0fNdI2cA8wTBzhD62uaCHlWI9Vu4Lr6mpweZB3UBZhTv8gfEMrQoDuGNVDf8Ht0tnSqrZKS
VS7PmWxM4Oo6eR4QxV5YBg9J83HHeTSH7vyYeo5xmxS0orVT/FDQjsnXeQENbAb6PllHrDf4FHA7
zXdxnAbBfdZT6g1Y5EB1Rzi8k4UDs7IAFGIstbuO7c5xNIJqc+SzlSUR8Y2Gzg/Wn6/gkdQSRJzO
6P+Tyod4ic+5kBXmpsMDs9Z30HclO/SOpjIJ98ZM0V1bJkSJ6LUbI8c21qpyMPCNLberGO7xrfJr
VmyHbaMJK1mfiaV4Cpx5Wm4B5F35+unrzpthiUo+kl8I8DHGulhvUnXKriPzcyjiaxIxEEF9Hm9l
cx4I2rt9UTPIvi3NyKawvisvcn7N96Z+b15+LKIC9IdO+x5lOBxygu4B2Ewqy+dnkO+kneyHv5Sh
ELHLDGZD1V1Qub30ygpQia8yzG6miQ/wxKcHo8ybZ1JfbNX64yr86eFYj44tz87qyFXKnaTBq2cZ
I04yFVsKqU88NQf39Orwguatf3aRSN7PyLbBM9XMA5xzACJ321ogyYzK+8JOizI/KiLkc2JMXuvr
EWq42c/ivcsUplaCbtBwbf8iJIYjt6VKE0HuBrh1OdfT3Bm8NN9ey71SGa4tVaB6XImfjVg7RN8+
Vr/572IfjC0uy1E4/zeRiD3E+369DLLRONY99KRwt9i5Q5hNgg2mPcLbWjIbhtzTJmM8jqVuaqX8
IIK+Ln7XySmK8nbIJT/HeqeEtpsck1TytNfRKyXJ1aBH/TOunnKgbuFC4JCPbsGa/qGLLPvaVOME
gG+13BoeGnFx6HZNBy6UVK6yo9eqBcyYar6ls2hfLG6bzO+iYxc3Bpap970HcHegXchTxyp9QrYk
2AZ5ILweZURARSSuvN4Hf9RZ3+QlNimZ61Mafx38uIbYM9MMMSdMBnH1PEQYhZ/zKZgKq+RbdpuJ
OO46/PvBKNYk2zkkfwO0BiLBNgwy4B/2v0vQEzyUtYk8+dellrNNs6AxuFRFNQGKADX0luYmx/ao
/sNgBOuUruyIR2q4k/509JC7BgAbqRW3nU25iiUp1mAn33A8Jpy4fxp9uIeK+4wsUBGI9QpJUaTw
T1eYPQybp2GmdRpvmVZ7EAIkbGx7ccBrdKTQlZmeUOaWWuR8rQTP7Lgp0x3IdTTSLujTh+VVfAuo
qXLlhQbWturntl3sy1PLgki0Kl2c3mXTqOv2vwaev3boPaws4eauAd/MseQhDlAL7G8bsDP72/wJ
dayfgRbLatQf2VvzEpega0i49djMgdIkOyUOIINhhRiDcIyIUB8kfmkuTPlYB0eXkW09M5LZs6of
/f5/qe/9Aubjt7xVCp3MYqeIoa8A3BvFc82vFE63rJ+WtEazDW2vONlZPJSQ30855j+xPtfIVW25
ho/PmK1cT/qTyu95OMZb8dcNFbz+c74YDVoK38Jf9cUeznnJuECTfND5Fi00JqwCHZjyGlrV5XFE
sJyfnzZm5RferZ/6EOcGuhw0lMI6N040fzvNZw+K7dTEukkDTiPyYH1kksXzFkPGm2DW6A8seAnT
ea5s7F8GbHtiWH6NLvfh4BbskiF1n2zsMWO+jVnVMuPTWnFicb46R4TWz1t56U0mkBt1UcDDb96g
+9XZtRO/xNZx09rBsuXaXSJqCnw5RyU2wqyV9Km2Om7uwYPLt5bovdRS/b7q4G0d2cEf37CE73DL
Us6KaDn13JKrmzq+ePiCcBTgDmO86V8ZuzHhNcP+BS4F0yJZF8VxieeoIiOrN7Hksf6l/PRRudy7
aqTWmcQicmqH1utY5+uCaK26iUg7aliMnUQrvZsKdXVBVgEZugGWlYkHiSSkQQId9Aqq/tE+WZ6v
INSgwZJxhzMPMt4mptYFrGAv67nXqOe4kuiBI02MSRIAfAE5n/KeiKIKm0d+jrvoS/63cikhPmCD
rCZmRSIQFwQ96/uM0cUnjiqJtClm7b5MP591RStOokSAY9LHkvwX8OMYww3aEXuRxFNkDBu1tt1G
f8828QZEhkP07cQOLRCOv/o2Gq4Wb0XM/QPFpM5f+bT/ZEnQPmnvs2HWOxRAAp2+KJob1D56aBVV
dMUzcLDvXboZjTP3RCUOT+fGPBzj1iqLcpP03CV2LJpLM1WieT8b02NRt24OhC6X8T71FSOf3I0g
Pyjz/BmxY3Jr56EfPssfF02B7URWviQbjVg/MrQGdI12uaBXF6cPeB/2GXBxQg2kTyhasNyPZ1j1
Xjud1hj3VFQ5yR89xHfnjyRxLPBgH4vVZ4XXJ3TQc5SFub1fA/CdiWfPczMGin2FjDM25W32OgQa
CBRgKzlqvYuJfvTKfbphG4up+PPToyOvgiTmepUogMrtQlEePV65qxV9rvN4gSwxy4XLTbMPcuwu
3EQHzpLAFv8YD/KtZALcb3FTuDGhv7FSXtEeizDFqcH1R1omA1g4JUVv/d3UYNQp0/2JkwXfyaNU
JE+whfVhSl+xalTEleXq3OvdnjO0kOFkUO6M1jtI+igt4JMhbizoZn1vAxP7vwx0nUr8le+j5asu
c8/efcwazwuHleye6Ch823QWAXT7/swjij6VrzCKOjn7RWydmMh+RwospQIvCGF5sJwQO9BIrZav
s3z/GJ55zsc26kXa9C+wHmB9QzHSmD4uTTL8FTYUCyJ20FTe3dm00zoW4ZJVhVP4+hyMO7xrZwqT
qHoGfg67sbvNAstzSQD/bie/QaI/QW4YFFIbiG6N9iozM9EI/y6b7s0HRbGV2pOKizWg+PwdZP2I
gy+7p//Tu29XPlRon08COBR9IPyrxYo1Lm7RFlPKvCUB5DADZTM7lPhy/dRAsA781a1CaKF3n0H4
UAv/jew0Zk2F2o6V2KgOWlvqpb+glbLcB0K3mQoZTPJ/KZTlAT0cUKc3soyy2zc/dJoSgDMTMjgt
dg/7Oza4VzFLjcjv1cqU2P3ReWpOSxfnF6IZgciXOU2UvEeNQx94ESgtcTqLFEoLgDji4BZSHsNp
7xK+KlkUX91Impaje+DZLYOc0YB4iUXe8VtOBuEw3/IIsa+WkpcBt7xI8gM8cdQsZFvHV2Nl9h5z
pfVUKvOo6eLlBiaK/Nzn32PPior2P8ch3MQzDWZYMKjwLbAw5HtXwc4rELZg/c3Rym3/OQXdb8yO
tewFQZ6PrM2YJ7POcL3pSb9EaArJa83ahup0g9YiFl4/DQNDqpwH+Q8A00Wu7Lpjs22+zMVz1Ggz
UxXXGF+atyJHjZ/PxNpObe8S16KyB75i+e6hJrmolmQzakYyYIfoB62qU6r0gH/20X7f/2mKknNx
BrDwPYxEu+jESgZ6qIWEepdDyewXuDSHgSyXT4LBITMlnkasZsxQvMCg4oTk7Yz11jS1Fa7Y+mNy
q9RENAtAvixMh6R4aVkaMXlgVvk2teI4GW/inTLMaF5xdGUscI72py1LSngXEquu6C+udgawGMF1
KQAP3W3T+BjLbjZ6erLq50ybTpeXP3SjPu0SjlgXqZfk4+s1FDmjwrQeDZ64oL4hCxTQZgU+b/QX
wmEtnwLkVEW7qKr8K4PVzCdXOWHOpYzLfBRkRHSSTD5viUwpX1fO0WcqByAy/5/5GHks5PjYknvB
DWSRWLmB1JNrVN/Xp1LWpw8EOcvgsMPIp5sPTnQEBCiPo3HgzoPIQ45gyqbcWA+oKzAvYUaQa2ZB
0FLsxEXoY8KJrnb1eRrSnFz5bYMMRfCB2iX/UV/JVA/I59hL43fzSLn8vxpmVemUDkaG9SUOLPpm
HV590OX0HVTtP16SMEuvzR44DM2HndDiKbqnzUNcBWuYucK+l4JmkFVzqLh2T+0p3gZ5GefDP1C/
vf+sG6f89AkjGcLRwWsg7+YqY3cxI4vT+iuSynAcYApSaasYfo3EIV4tuLzQ604TsMg92XpkgBHR
B/ac8NfqM7yHSdyU68dSe6a715mpZKJ5p1eloc3FAr3xg5m7HGp+SkGQcgnoAF/VEo4A7RwpYIze
gjNnqTL3wK4moqCAXErAxWW6XcCecsFgZf/RuuwBNyKI2h7fx5aQxEkIMH4OqzLJncO6TBGuQC0f
K2WWwqfXUnfi3zhWBKiS819HPO35cilxM/7JHl5Qi4wy8FXFmu6hlVZYrXvtsidlTRMYtulnUYi1
F/RkSn2xM2KYhImjfgtrctE1FSYffHXGmhmtRVsVSYX3W3nB1pCkPum12xlVtgpfswLKaWbJuMy1
E66W2Gdygtt0+uMULcoDw61JIcCWvzJlWfNZppOejB185ah5IfU420JMPi78xq4kadhBcfkQgdPg
sfQqTCflOWQGBwu9Z8UMEPFRa1IdN2+tkmanzrUqAe/On5ZBGlFzqyK32PakKnvXWpg0/PXMTQyq
fP7AmOeOwpsVTCO4/R8zvSCkkzgZbKsek4VwDEEbd/2uyFrNiGDunELXNyZZGnJGP2SpWSBUxN7q
JdhCduugOyqid2IyzmMCBf7PlPjUopHYXPXSNde3egTCeL1N6/oetKyE/zhChM0g6sta4I5RgxVp
eW6HQ/gqh8dPJqCri2awwtiSrNSTMZF5qD9DvNFNdibv4sThLCxIDiJEPk+8pQULK0CvqjcDq0g3
fw6YsRu7grTrNzjuwShm5qJi8CwfX65CGoQQIJLNnDglPTkLVf3LJvHVIDkC3p0L6fnRtJi6I8NV
swZtNouEFPIXFC4u/mOQvZBrcZD2vsQgpefeUn9HtFOIrouCjJEwj+A7YaWb5UehnUEk29gEPPgg
WiAMUkSxaw68BBvhgsN7Dw0wB1OnMDDS7mnR60WsWtxIq3eLoccTnN2VXVLhyQOF/W0RdD7Pnlnc
g+I0/++M4zhQK0/sbrKJZN6m56oLnhMRRAunY7kdfPFh5dd03HDvsiIZVLEmMfwpE6SSH4apPr7E
Jzlf1BmCoyb2QuE2gmwgOClpFG1Ty+zknpAPTdczizPksQDs3/Hz5R3IQ3KW5JsMqkhPI6odOT4L
BeEgELjtTjeUuqEvjXTV5Oiq+beEbYnKNWUKt7Q5cSu7iw/hqkOcgBWBMrw2T/IG8tEm7OniOKFw
s3bjMUXbkdYxDEEMExTAV5cLsuqpR3fhofxJ1SV6o0I77Xyc4Rpk/Ey43rTsOu0ei1BfuODiCpO/
zj0knVbz+icHpHxQ8MV0VKGP0IJ6o1KEMVEo3jkueTJslSWZVxKEpEI1RP3MypYKLCi0RjqJCGiR
ZQNUJofz6HVGr4n0Ucw5lgXkYgfLVIV6TrASsD3VIH5SQj6SqmdbHZ59Vt3xH1pWbe56Awrw+ZT6
kaB0pRZblwc3q2v66YQauFgJslGQW84BRIYvw/U/CZ+x9dOskqnjEM8LlTYva1vpxEHgmGydBwPA
KZj4tpZeojjTuLrf1jvAIWBmp/F7onIU16xOJwDq2GDzzK8VBjmRecEmWJGqYl52Bu6S/+7T1ybt
/KpaS1wp4RQ5qOWNcMIEcHwFZ4XubIds9fu5w4Kg4EhZiStW6HxXnXwLDt9nEL3dbiITPqerkvCX
lPFh60RNAdyf1PS24xy2hFa57u8VKjijfJIqSLnKEd8ga2ZEkyQ+lQoZw9+I3Dv/3RSfHBwE8F7Q
m37K8of47sAe04QnrvOYYBsf/otYICLHuztXL8foYzGVdStU7x5tKunxx3Kc1afEXCrGtcwgl0BU
tAP0v+Rr3UU0KjGCIx490WuAnWiTiRM4WRz424AbeqelhCw2wqd2zIsZ4XOqoovoOIZ8UVRn2zIE
zDgz8V6itF4kL0y+iwjyM6Fa97uxJUhG+r70Dl6hNkdJgWxmSCRuS2WXbuAyYNvwgCT4mLaV8a6O
PtoiIZuNEy/w/lk1iFrk6LEjwgMeuLj++v57fHzsYK7uUIkO4JwSVaPqD5JvHGkeyQMS7ZfG7/qG
Mp1JALIQGQF6/zrxJKoepgZHmrFMRR6q2m6skOqh0/ftAeOnw38szWHRbIHHMKeRasg2IuFOmcj2
iO0H5jUqzf0V1P1ZesMnw05V22fkntZ0Hba5zkV6HS72V5x6bKBYrF6T+1gzRHuf4V6gQ5uQ5khC
zo4inrZxsIfRyPZsQpoWjfbXtLCYb/HLvVwf4rD5gRSksIn/SExFXHLYi7Wj7tbqLTo/k9B2rFZM
MlKYvoL2nSlGppnNnT/s/b8Pjgk3W5cNmfXW3sOGy9iIPLm6uXYR9gg43gSI9S8jm5iyofXepXCh
7oij0PMEuTMZxEJnBO26N8oEJzA4gxQfi9ewtel822f/+fdJOZEU5ilgoWbbNvbnJ9iCSrDl+FwB
H90tu9UQ0r564nA5Ot95Mya6/NY2eFJwGZSikCb2VLiuvRnAq9iyEyx+W1cM5pDoZNavB3nW0K7S
lPFwKHFtvRIwRbRrZbbdtU9IHN94O3jLRrW7f35uZHLo/HOyB+xUgKKQBmmsrWplRYv1rtmuN7Jv
2dYVn5rDU8zJuwlq76IesflPunsv2+euNaB5ZnOCWrCekAgqGKM+muFwaVX+OkTpVVw2r/wuirZN
ewWZ22rXGlTGF2cVBKQbA9Bi3NNfBkAAI+HrHVHLvnKxJNoBN+W/PS7l/1AJyLdW/mak5PTz94ah
F7AhCb/8Rag7SMEjGp0vNXcwdj0sp+wt8BDg0NsmF0nk+jgSn/gKGZO+iZFEqOQMRFJewQMJKqxn
xW2UdZRU+2nXBdGa5yUJrks4Xd+awEcCzs9BaXzq6WcaVs3BGGltHKORjhq8/nzJzCViTQOnBDtJ
3ELlwMv1OD6AOQ2FmZmF4yEJoN1mbly9UMis1UxchiBlzH3XmSe306l9R/pnMpqpapoBgW08K/Nv
sZ779G/LrAs8qsvBewe/8VOAYaCHO3YtOmUvnbtsWPfADTpz6MHB2DGYr0MiQhST6lpaM7WOOOAT
fqS0vUWMHfOrFCKH/xQipjUkOZdjaz7M58b6kqy8G5C4QWvsYvAjZ02OrFxLLq4JKr/vvb7ZBbmj
790b1R/8+Kiqk0UtO4OwQqbGJlOAU427wc8ykC8g0/Ep/06B/U6ubKqDXCTujZTvDCXF2/oN6PuN
XMu1I5cmBM6gF9tIaujIYaDWlHgkXtGvICUjnf19PHWFwp0dCQsq1oNdXljhQi37Ff0PxkCGp9Ol
Ea0qiqX+VoXH8uQmwB+BO811M4A9+81UJPwYNBRed26MfMRIvJGpR1fX+6KKFOHXvCykNITlH7U0
2B05LMXPdKLoBGP+gUPZCwNxS0lSX3uUx9tDtfClHMdM8Pt7w0ZUJuui8yjFLrL/C7mnFT+0s2hG
L5NTwFrMMWELr8OdJq3X6Yvz7pE6fAhvLbKqV1J2vXc2JowtseAwHear35Q5rlYqGRXc5rHc3273
ikXagfXkqNfOizmciyA2jslO8gAZokIkRMjooQJgTPmgOk1YS9GhiLwfrbQzSqEt5Huz5NE03Q1V
4ogIv92cSSvhpWoG3YD7l2Jj5zKrDfGcnHO65o6TcmSrPaniHJVma2UlQu+568BDQ+povh4W70+i
eo6ZPQ9Zo65qWByS0Z3HT75XPMeC6VNIS8QOxmEmtQ/Dt6GbvUlcz1q+TkQBg6ZpGQlwsNE3N3M/
ViVVPHbS1eQyP5VP3vJ63YDIbUFgoozpbGbBf87Dvtgrz9esX1X5V5BhXEakGYWL9SQuebIPwVk0
M+bIFhIFj+mjH1rFWDzTrximKIy3+BO3ep17sz85HCLuemNTz5WwwGfrMkRqrUSdVBomOPNpKYZr
qmrYohHGAr8uA2ej0JOu3PJHSWVFlPhwz8qMahVwY0/piM83Mz1ArAOYPoYabXZQaXLA/dvZ4Jqn
d+oluyvENzLrV7YUZSd/xDbLtB9baCdo8OPWDKkMqKII+WHE9ybAdBj4XCH9ErBWpXNmR42m4StF
Xl+p0eawf9XqlM8kvuXPziu8vMJVv+pB3HOQKecKJDqFoLy81FmA3T/yUtQFfkyL/CXyUz0MUw7R
x9U2w2X0n/B0xvqBTUUMOPuR4UjLltkhM/GygLjYQru3bbuKRB081vPQ04xtfTRny6gKiGq9FXu3
AKOYnm4E3fr0RdIeJjjKLL1QapwlPiecR5gQ6z7Z/4BqCHhXvbjgFYRqb4NYfoo2Cd/T6Tlygp2k
i4akFlqjMgLgPGlmFRdQmSHYNkdSfRV3pNcszqtz+DN7g7xSLYqWHgHqEmuz90yAkQDG6ynRHJ7V
He7Tp8+fbsq2Rw+ySH7TOW8HxFIuiYEucGUlt39CTpotbsH174HKvwp8ocyOPRyBZVyfk8be/Oy3
TdYge2Q3vWoW8ibZ2thWU0lkC21o/GZM7IB+n9dv0JUOevZUfGxVWAi0aRGwz3ArvLcPgVgQEgU7
qBKL3I+ogOXRSmK+/lsOrNp60KxlFTkcyNPPk6gLqkCfLr9MHJckM9nm0xeheJDW9xXrHjAlrpi+
xduSwWLillFudCUNSgsV1QGqNo2giEizDTMM6CbRksFqXss5Dt/YoF8+2L1RoNI5xRGbEYAknf4M
cQuM3yYIt5CgogWaII2VqtQzr/fOG9YTkR6QGagT4deBQeoEjzEXJIW3ghbFCBC4KBD/1qyREhxv
MN1u5dWL5b9KfagvRgZyhNZqmdclGtaxZik27EMNjURMXdju05p2G/Fgl2KTtvNt1OeuVKJG9V5I
kMZ4b4RnyBZbTabhMcpVcI7Gubkl7H79zyaomUTqWSU5kY2MFFdEAact8x2i/1YKGctk7XuLT4cJ
P5z58bdByqcRIQfcWbJGzwmQGm1KSSvIz23v9EdQVZGtix5DXhWxZqsQKZbzbtwtC0wVg9rbq1GE
qLdHewLVsnZUBZIxM9P8OrKarXCZ1XoiLFBwMtfxX0aloZ+Ktl46IT8b9smzTOagMfXxjR8e5FUY
sCrxZ6Q86Y3D+ImAD+rXZWEkrOjbrMSPCIv5gS4YbmqF344SIUdP2lw8kfkWMz9fXvYEeMZNlCoy
1yXEMR05Fdn7rO1FnALovpn1RRlEIuV/4gFZEmn228fAiBL0bLEVugDgTnmicE8VyPOikmSVpC/N
TDRZPUXgD7mSAMRzDHTtR9knr+U3QhESpF96KB4mx0wF3g47eT9C0Z0ES6kauNAcU2vJO203nmQ2
7CMjECYkbGj1DCkR1eCDNtVbi/ORM2RntpYi6Hnuxd7t4na5JJufxnUIz1GgLuHT33vDA3siDvSe
9F4LRtESqEUYbMjVzHONlZ7NAdPqKploslX3tHqf97lKjg+erCENFEinbbv8iNPm0KM4JPijwh34
OyBb16VwXwFLbbThqz7zuiYUtTWzO7lO6MHq7u1C6DhIQc9QTFo4Wfr/skErWYHllBh1cI29mZEL
BPvrqx7YWbsNHa5Fypn/dzR1VPk3D7OnwHke6EWBRK+y9tt0/RMCsP0xgbCFRAn/efy3rdS0A8S+
qE+mg1QGz6d67aBgykg05s4hxV4KEjGNTOV6g5P0WjCKehfx6MQdCm6fRiGUcnpfVPxmqIn4ct+A
A3G80TkfawQENxFoLX1hPB2eDc9g+4t//MFdQcH8Ci2vs4KzxUJDEH/Dqz5B/Fx8xDyit2+FcwVM
Fy4Ot5g2WovpCQaH3zC8zBKfb5KuhL4h/LCV98vwAzX4DMrIX3sCmgUv5cJ0+ZKduVySs8X2En1c
Hk93Yonxf7BiktrzLYVqP+Qx8CWHv+4uVQ3Myj+Lf3s3U2KmL90KBJaG+v0uJWHGzZF+zlYLh74k
/Zee6eGMoLRiXxaYhBEIe8tsNetNhsuG6y1arXuCVP9OFgnXlhOOs7CUamVcVhhV/D/U9Gtqzus2
eVQ2dYyP6NcsVk/o1EP28S3AjFHmVFJgxZtiKP4XJ4gd5pR+Po5PA+kEupRFjL1QCwfE9SGjKbrK
8Q71F4eXBvOwmzE7f++GF0as1rzigjNdlgt8I1TsznROKVuuIf/r+mBj6c0kRDQPE3sETJjNI7d7
I8/namncVfg+sgaoxayTsynwyWO+1KhpYKFnpEvOvDuAnjhH/mZv5T+jd3s2NUQPF2FjzgYEPTjZ
ACDPwa6/kpM0V+pVRlkRlJGW7t+cR/zogMBAc1oowS1wXvODWhTs0wj+9Pm4YyY7u5vkclbXUeg/
ZPpLlqZooPe0CAKfq69u/EEM/tvEVHa757DnDISA69wATMaKItbf1mj/7RfcN6PAtHtMm2TnZdz5
GqkJuozDWOEnfo7wvry5dQsaRFyKSccd2FmSQF/TkMhjq2//Ps9TS/gOwq8t90MEVkJfHoH4U7tt
qG5fiXhbSgm6+mQcpHC708NMcncPd7zzVcKl15RA6bnit5oxaVs8ZiwzyUoRqwivuWsfyOMXAKxa
bu0PHI4RddNQt2SPe2bYQEuSoQEY7Q5fp+0HNi/l4TINsGIwhwgfMrplCjFJxyOJrBHecbvQC67J
lcsGN65fFYnHRyisSNcxa3a9cSgr7iYd3HOYen8irUM/YjqQvEjXnMmf64m2QDJQiDC+DlLw+f32
hPAcEg6p/PpANIEEcTK0d4FO3Pglku4AyxVwciF6oYkA9PtoHPkRWLMO2hZtrnfFogxQF1JWrK74
zvk7UmW62M6A3Lie2TarLhznfbc9MQ5LQcw1DV1n0PJ6zdoFNbS2PlUCdGODKW15JyK5SBVCnkwp
ri/x0mzszOF9n9fOTC4+3Y8ZdDXwJpGw1TQcP4Jem5IVNuginzC/yZniXlLl1YqbcqYGS7uWBHlO
bk7BDDJwodXmUTFj2EB9es7D2uwhe5H8cEoVNBc07UlLsU+bnBoFfZ4vD7bNuDUxT3BiFWQVaiZH
lpjIfjWneRXEG3pcnxv9Hi1p0o92Ip1TRYjGj1siLkjkCy4pd+crcygT73PWTj7i7cx/eXC50Zkn
upn4bpLJ45r6ijpP3AMWNDkvM+e6tSedXsnWMag1ST+pwsAfgXCtLHE/pVxNN09d4c/hBHlA0N/V
wKnfbVHw6KwEkcSg5GqWSuCJK3HG380ZXiCl7cxhaBO0LmYAeb86vtIncET8h2VSgvbzB0CHnhAV
gtfAZtHoF/F1Jw0n4l1/6clwq8YevINNE0/i83eSCvpcnB+hgsGhrImyOlT0qy/AFdb9HATbIh5O
yFw1HTY22Cfvg8qlnr8TvrIwfSEM9yOpvQ5OSDPKWKOlxLXMcMU+7sn4SGu6mE+Xrz+pa8AMQku2
xtzqAVSHMo0HbI64XN0gl/8UcDx4ClkF9gzlhfx/EbnoBet5aMKnCzSTAr8NFD9uJJ0uDuFV4Tkm
DgwLQCZjwHsUCFSH5f8/vyu+CKD8xh/Fpg++udvqFJsOh82Xe/XFY+dHLfWhfT/MuI4koExRbzSy
U0W0FdfAmRq67BFc7UpoiwutJP69IF/+d1PChcNNijnEpWuD0ypVR8KXKXbovb4xL3waUmKVuJ+G
CxO10510j5vpcUGRM/XxhqyllqgmDWyKD/PxsdHf2gNYtnuu/1zB0vjlk2aqu4PLMNw8u2L8C6wm
5uOa2AHf84K4sTkSU/QLWtxTAUSfa/Z1jSTtKpsiDg/LGbMxh2GETnCKX8k2ayGd8TernZgY9yRr
KadxCqQtcIaZsBQvp/XzDBqLcLB8zdq46XoAowm4iWle+phHEQ+lwUgWlKVsMru6OyUgZ4o/5F8T
llG3NUR/Uee4jhQCM0cAAI3sUCx09JppkXBGo08EKKAW8fT98lzUWC8jQUjmgAjLlbfT5crpcQvG
Y+vLkh7T28y2JQflVyvmccwGVB1EYnrMuwhT/chLGPzKynFGJkCZvfIAwzSDKHGqC/RRN9DPPjn8
cckGcYeSWxGl+Kzy7s2sktyvOF4cn7uWxNaPnOnD1NMA/9Jnq/m8dOnlyptPRWN6Yguc0CBru0K8
1umrsugXzMR5+xfyiXWg7kK55YjIBTZtw7vy8OWnCKB6J5c+ed0+/uuKFa94BsyFk/cwiF1cRFul
z1JNO75/HhXjsQkEsS+8sXcZcvoaZOUIhT8LbSgjXcVVVyMZlEgXTIGk4v9aZU485k7e3yXkvORW
diVa8DGfpfsRJgqdG+9qwW3vzXief7c4ZAId1jdaAdo6qVIQsbrnuu9ihcNc8PzcGRFOuEQVF+7F
ehwkuGNx//zz8NzjElNR1TP3+nZVH9Lt62eogsFYeTGY2GWJQknYZ910B7h+LDX3oMrXnEHCnDEH
zNcU7h7B86+BwCNZoO3pvGJ5V/LLYVfV0vF2zIfFvRUShQZORSMu8KdAXy/Q8wdJSZUfM9Or6k/x
5NZ48Nw2FVdGXg8vpoYCjrkJfV+b+FWWMU3f9xqG7nRfEiN6TSNeBiMx5iSHSaIbK4aLcRrGiUOA
7nxch6M8mtnMQTJvnP8d2q6PYz2SAu4BDkvyk/pJ8leV9phrAxLYSM78gmKRbVgS2HsxMdLdnfpc
EAT+vAoFFWGT7TyZdXKaTafeEiWLqBytaktbJMbMhCKhHqMXUvQVMXoDYmb4S2caWRiga49dtiX8
sYuaAe2bC6RyBC7GI2hL37FIX4NbWnGh9O/TPCxBYqUkSMKgDZ0Oa6LQu6uija5rljML7pTjiGaB
UggPthgHsxhW6UGB5lZo2hnvmPVbS7A6OIUs9bbehCSnWilpxag8aLH9n/ZMEYbdq7gQiXal+O2H
8eId2w8eHcOw2FlMFhQRAPlwWWPKPGL6TcV89lY+2TG3eWHqcn2sjnl9n7ZFQHuAUJToYHxzA4lv
wjE+r5cg2SeKq8Vv2EZsttnwqk790gQAvM7TBvHaNU9nGZyjwYhW7STws3yU0uQYE/DqtL1h+eVR
6OlzwR077geOC0ydRdD4Atnc9shMMhPBTJh5ZOD7atWg89r7zXdrdqvfmx6FSUYbLYdCwVpz95o4
nGZFx9Ol7Be6vnqVLdmFFz6ZvgzLpPl5plXDS69HllsQWgscX0vtvtpNooRQpbYFQ4kXi0QK3umT
h6p5OoKzm5Ben7udX1gW8tl5NVt9oIC9JE24jOFvyy1f+SVPIBlkMTcqVdQRSh7+2git1h9Slp7a
SP7gz+ppYUvTxqz3sr6rdqU6PfSAFpC/6QszzbKr8NvdJS4c/M/I8B6CUYRH5Ak5r58xGHZb7RHe
ronlouYC8WxjHAjbjecXw1okgMBriNLmHppxO5h6wp0PZQTonqi50//sXqfQS0Y627rCHNjK3It7
SxOrgx1mHtS3tjpGxLY9aqY2Qp6ulu08Z5wdK39ZG610UnR2yAYFN0hdoCkayymlqASAkl5tgKGD
jdyM7CHv1IZsBRh/yxYcJdKa0S21HJe2k2WcjJAfs+8EwXQksVtCBcXQ0FznlTsLmi99e+4FXBdf
ACRerYwNwzSs4gEzoTiLtSWFwkezlDmQiFrW6eyvVie+twbP+2dRwHbZb3fBPfETEAKYc9BVJcF9
j+42r4CV2Vz/dubs3kauuVOasnUQI3A1YxnaJ0CAR6lIQ7zfckYsc1hHQ+9eurZmyyUBraep5a1A
KWTxN7TO1Txjxzm+kAURSgnm30sKA6KX9yM6v2VSc8zzn4V4/jbqQLYtAKnwuUvu8CA+dgBao03v
Otn65PwEDOxcInnm5QUjFw4gKaXvojsJdk9YLg7hpG/RAn6R5XDiAwy11lPMr5t30jSxsVLew+iL
4RKe/DWV0qrNawsqY1Yfzgo4lJK4kuxwPiXpdMuBM6o5YQKddm3GHGLOo0V9U62yYJCgG1ELP5bi
eSNuduBqYukOPII4BpICRC0T6CprJN5k8gz/UjRrXfRriNnE9W6+GLuKcIryVrFHn/W0ZyHldEyi
5ys0P2FtQdLMkZBZbatAtwduJ59/FGtgVZQVNRnHGS+KUviCnERqri2eqGwi3LICfNQiwWEsh4Ur
qvnqqNGljbIfnX0Y8sRPWMEopRluiHQtAutTSWg+DDDe0hm0eAH8GwS7mtxM1hcnnpIdEWW6SvLD
xQudH/0oWQUXCSzpg7oGzopsTzRBTeFDWG4mf6OGDYJ7mXGpc2PIQepu9kMCBOqd+nbfX1QyRUln
GdZm0xhS84qcvDClHs/PUs4Tjj6cNbzDMUpGFmRB+5tvTodXpsbQHURi9vrBMy7zuS+haygQDnYQ
kvNiqickfc3P7BFLwiEJ7Mst5qgsU29hylFwx1qlQzb2ODBrGoAudr7XLB6nSUXXeCNZa3eK2A7E
u7wRzJ5TLhmM2Dg4ojTsFB01C7b6B+RO+2s+hYZxrQrbPNgbxctBigVpYpac2K3EwNFmP+DbEucE
DfpSUTBbKn3HVw5yi11QX3+ioMGDZeQJHnMYRxR86Eq+56GSnEeMh/D8KiChpeCukSIJsZzaYyun
vqQgd219cMP0EEHF8WSonJgHHP9EtIAQvG8qYev8YtBF07N2lwASv8qUTGxYsoO6apODbgv1lpW3
GRQgwxC4he1dAvf6aYUaQPFgLDTbOLs2ZfSXvc2FAYFUdfmIcH3F65FhSqK+qbt7eVBcu6NIlF3V
C4prE9r07BS/ACNUR+u1xQqZarsiSr3pvuAHfiT9qoSjtc45CtIN1WGzrCAtf2XeGDWcRA6bGgtb
hsxGBBvFwOs+M3to6beQOUO41ErCDgefrN+E9SLxpKPMdPcqZiUMboZbURqfEle1OjAGtJcZ+KSm
ZT7dXjCT8sMpqYobZPp6T5JXgfKP6AdfXdAirALYa7hbm3mm493wTbXLl1BQZ9JixoXhvDEnMelv
eW/NmzASre34yEgdLq7DIog5DPNj2AP8xewjTasl+B2CDHMrIP7BOiUEpqbXPXo6dyyeMNiT70mQ
TwawXNPwPj6uu7Mn/XQrIFm2k+d/Ftrt1ko642BF/krSndDmfEW9+ohyv85zy3Gu811szuV6R+zs
QN8/M/WkxCZFjmWBghHWKYzRTA2BOglpIDVPLeY3BgP8631nNYo4BCUyZ/yGGYcAanuExPumqFTh
gV9833TofqpY6fo+VV4KRbpBCnhSVC99tV8itJlAAyy5hjWaq4u1uWwLW9FhKKFrRqFd4b8sIqSX
6sKGILxXkvc/fwq34XlwlW4b2jybNBTKcOqvI0dUM5cnJOHjtMTJk99/e8lipjIdJV97t7ThAQHc
TJt3hbpPurN/MmIDKF63yeoSeEFflsPevrv33kKKAPNgW2egVt/4lv3atz2vZ66ypMvxQe6peLJi
5ySP+sKafasSE3Yx/SpOG8WxstSz6kazNUQ5Gy2bDidhy+3hSs0dgsbYJOUZzCAwAo1bgyVg+Iw0
ZsYnlN8s+wESrl3ISGUEW67wWMh7xHzQ8ihIAr2ZHcxMIjw4Hzpk/ub/J0UY55UNxxhXNICDc4vC
rG0NK+ZYJ73ioHXmfPYn5mzSP5OKL7qawI6eNOupZAj7GOqcuOIFup4OsWYv66x1sZNv9cSMRNaP
WBa/mETHrsPZ3BjwpwIsri4SYCVNHDeVn7Q/c9oKR5BKnbWUUkt47+B6Kz0/9cnAi+hTiFIU7jao
5qvklJc8xq+eto2cQ2QP9qe30BptBJyYDBvME0XvzyYMtV+gNJ9RkLtOwRgEu57aRThmksCOa3AI
ocIk3tYvf9AhLur6gj3aEmtb8vWXN3IDykf43Z2yB951c9MbJBa4ARanCCbiKOeRRCkS7c+WqVlt
dvrfjQ55ovxqE/TQfN76ZwmAwEiwsJ5Di+OY/9DBYMPkAyn1aU0QMIKT5q+jKTP2ArvhXF305yyf
qcpte9Y89vPIuzQPA8XDDjhuGdYd1ratLYQbvx+8+njtDloIOyJ7c01fRE+C4Bhxgmfu2qBTZ0Nx
t/v3idqUo+0J5/KzxksEfTETe3cDQTzQLgQ7lt9NXITYcPCZUE5qBjbTxxdDqfuNjcwEj6qfb3j7
hxHR26IHdpjcSJQ+si3udmuTtVblmkApo0BZ0kloSpQbUqWuOSzFEUEE6q3uRKDr4nEB7QGt1jJD
NwKWqAEZgVXRmdzB4J0Q/uFzFHQKfuoEtDvG2Q3U2ptu6VIIqk9qZnGNJrZrzRdXFau/VT8y5XZa
SNGccFSxQZwdUxmyxEtftPW2Ep5gBHic1e93Mmn39ep3m01tR13C6jMRD3AUOTPOJEIDRMz+TN0h
XOn/Swb65Qjuu7rvStEXnpnRymetDnd/vZ2LXTx5Za66LiGHAZfH7LpZeAumXvzav1yluL/FuVUp
Kq7H6YFKI0vC9pah0uI0W6N+nZXHcsxhSneiVjepf9W4N927ZWZ46+1H8q5jkNYEFALA+Bi0eh2X
Su/neQGXQps4TpPH/9yEO6ajST9cf62ASkhyu0UFyl2Eq74KrNTjUIKgN/YOKHFNAqojLwjvpWkd
SAvmyrtTXDeaxLBIIxdHDbQwEjlDjit3af5aBgHryifYGthTnGd5oHfUo0KPj/+lDmgXJb8Olhvb
VvM9e727gHh2fPGUuX0KcZwMi4fEX9Lx7CbMLFvMmO3vXB42hybyOjdHaDE4FyeTDBvFkjNVRjEI
9hiE9j8Cd9UzdzotiRXXe4tBkBRwWoluxr29nQwXn8vUXKsHZPZicLfd6DkeHyJcjQ5uL4DFUbHM
a0adw4yVnbNUwRXDKrB7E5uWheCBiKhEWNcGEviD0hVrca2tNB8jkoT7Mjk0jurLAAFU1SFTTBwT
VNrPUEMEdWTJUFoCMa65fiZHNx2vNbfJ/RY5JoJRUYlZ8yiDVx+0RYMfml6RAmpVGwb7uM30UxBc
m+YpP39TEt9qldlEFFHYz28ssCDfk764r2QQeT6CxjorT6dJEBZkys3jYwGRGQs8NaAhqSimKz5d
W5JkDB2VW496goOweto5Fxt28xzCm9QDUwqMRk8Hc1LW99n3jjuCtfs6/TODHWgbhzWZWnTuyT8r
5B890Y+V763hiRBbB5q9ACdL5rF/b1pKbME2j7Bg3oYh2KpUk/VwBkzK5n0jutDGxtJtW7lP3gSX
KaLtr/DnGV3F5XNmKCpGLECMiphAnjNYBlHkO1GpPjRNvpvAcGdbYZNFfnYiQqR2vnRzqzzGFhKx
rNyKdJRY6hkMJ93rCn3/gywlNIbvPDOH/JRB0CLj114GGCm0Xh2A8xeyBhZfyqVXW9kdaNg7WIgz
KRpLnQz8ovNleqSTMRAuhWKqFp8aWtUa13MFcEWHtQ6UIgr2FgPbvsXPqUwKRkok54hgYNu98syw
RmHcRzclOMhCXUu1bxi1hlHHCQ3NiNmwXT7x62p4oYkvRo8OBtWV7obRuLWtx//kTQ04ub02YQGe
A7Py55QmjxJuv+kdTtBxrBnEURs4e/+LDMEmNjORRxpymmnViRqbdGg/7o2BTsvj168OjDBNYOto
Ss+odf4Q8/6DNZYtrtfNeH7oWYygyGJrX/bI7ZvMGtcu4WbQvbqngg2z+spGAhxNb2MUQctvm54i
FfSoZKv63kWNv0hCFFQYzUKESXb9EpE6NzD/ia3MSz61CoAB75rTSEjfEAj4X1DvG5il5dQUQpwy
+jrfYbalByhZgQiIbH/5F3qlVkEjeXVxSZaQFDfhGOwELjiSGNKQ6dCG4j57ZttDohsfhCLj3i+a
v+pcThL9cEpaAlaq2P0OzxUoCRgictNOOyhcVa9hwJnCYj1ok1T9EkrHervsDsfv+Uj3OTWgin1i
tB9Fk6S9GZPZz7koOqW/VjQASxWRByMffljGZNO7Ean8QgNTUmFYiqin4qm6Ak8XZNusNhBZ6fev
N/oy/qUb5TD11A2t9gRZsphZag3PGEIiEMJl4LrKlapkIjrgAs/2K/6XP3TXdnw+9hx6gC5FaPfS
hZli3KInR6ef41dWbnsWuD6TyJSZR2Fp3jh8ZSmmhPPsIpqzZQMT2lIAyo4arcMmEF9yT5qgXDsk
hjkB8ar3G/s/yUiGHk2svO3ik30yqHaPaOnveHqNha+YLqrMlqpvJGnu77ItPtxCTJwEEufKMexY
QOBxQbGpxEggvfNGL/mhseI2lsZaqFeulMkibf5b0POpp2UdADr8SfP9bNt+53lxpYAG8FFPnGWt
k8xnPoi7Kj5C8+s+whbJ9bpBVDDmqnFEzLI4SZRou1k65xc+BoAf0vR+2STBdJMIyxyAmIYzEaTO
TIP3G21yrYBHcgJLHdGXiomVefsJiS1u2KghP3cgVvJUu4pdL/otc9hmsz17XFi27Gv3Cdc7lx0g
Ec4GJleRrdHFkegXJM2YjmftPuDm500eTAz8oEXheILvz9pnGuE/BUmoFKBc8WUfXNdf7QdZAo+O
wtbJnemb+gYtCC66EOW+CTX9hdlKGG3WMDc0Wsgk9DSF30+eRtVxz+f+xTa2elWl1rqw38w3rFGr
pFg/plE+11WUtA6UqWKm0KSWJQOTm4WnATbqhiDf9YUNbcfwZQxyu19rU3/susNoEFYWlhQhxmvD
Uqi0s+LVvdS3UB97BVErgHxFJPhIWSw/Zio+qTosx8eLiBDcp2OkVM2Pw+hYYbyDO+1nqj9V4iLP
vsQ9hAS/9QDRV52Mb6SQZ5LYPDvHvMpl4U2DndrPqwdZGjgDxBGjos6ZFOutsQjzAVu06u4E36KE
iKMtGY5XE7zDOoeaX5DJFaFBIYEOqsrSbw/ojn/sJQqw6JGsyRpHLm9b+ApMxh6rQKSmkBF4TUVs
PPulbaVYQxwgB8kUpeSqBl3GfWAD4TBJQBR3maWtUQWYWvVrsiPnixSWH3HORGqRGP5cKUg/4IeP
ZE9K4UXV7d/rozVsBrtGJV4PRsXKaWCvMXiQZF/2IlzV54lBFznoEe/tb8dMEjvX7i6w1PCYMhix
z8HprMH3hGQTPJkbCsXvZCd3tninzJ2HyRghiZPETjCcnMsEirM4Dhs9mHqCMfUtzpu6hZ5eQwkQ
EYMJltWCQSaeLM8nuA9WkmN+G6qhwScoU6L/NDjWpV0QyIYAuz2YuvT06xh+szpkepq3vDgn49xU
h2VROFrfjsNztKmiv5g6RJo/C38PntfjTA0g3yUfvbVlrU9QMgP31ZdXkt/r7QBnUtQpEPMncAFj
Oj8k9Rv7jnuHAGqud2mAFwepEqR3kwim2XCLxRNrMPJYAqBozX16Jy+Vh1ARwq3ggX8SBjMhhX+L
Lj6QXXSmObqgBRQvmTLt049GFmg1uigxnPrRZE2WiwZ244EUX5DEx7iHJAcM9KAN9tEsr8hyp99k
CL/AUKmfuR9O4UGrJk2YIuih4pzuZHmvucbEOrK+Zi5874zM+6dFhXiF4GFcUhsHxxhZwHVwghiz
lVs1k/izxqHX2l61N/4GdxNWAU19ZMWryWARNFWUXcKmzEUU1OXiPdGm7hj30Ct0D06E5k5iuwLb
h7oAst/xrq5SNiuFB8Z0JoTLheMAaKrhftsqJY+V2VFgbmrc53i/a1TspDbXzWut2eA7bdlKoa/U
+S0VT98v0VvmSGm4iByngetveYF/PdvVEFuvTnEiQHbBNZC+aXIPiSL3n1EGJQ8EARzzQPQEiMHG
OFAQttbE7yeFR9igU3IhwfKoG2Dwux7OJ7wC+Msb9FpG9rapsL6m/rdJkCLS86VHK2fipuXVrKLp
G8Mo3cCcakMQCgZ5sYjUHPjv/1DwDub6XZRsTnY5vq1izpL30Exs1snhMdN7498CJhf9ZWThpyzi
rKKs0yfdILPxAzXlUGLUkr0c2/Dk+VPAENGiGFEKx7EO2L6OdYoSdyOteYiCwJDruqIoh4sI//zd
+gF/rpYmi1lsbARQT7vYFzSUUd2LA8nHI3Mcae7qwVGEtHk76kvj9ievRIz2JDvLtJzFXbSDUuvI
6HUKEZbPxfMb0uDoH3uZCtjpwYVDiwy8aJ3doOJ/XJFqgdqx5S5TTmOFGRRwJL5NpiIwvTIK3JdQ
8I7vHK2HMr3GieB2J5uNCS7JGDzR+qlaP0CpIXCEpsvH6N4h5G6Fb43PB3wjakne9CqNzckQGBzP
Zn8AMzoa0S9gj5VZpQx66rSIo6F6TYiWJmSH9xkNKE44s3WDV+ZCYWmdmwq0oYSvEny2yMH+SUeb
0nXW9V05xFyCQfKz5RHjtFo/gTuNeS0fGYvICvxTLDYsm0jzbr7ipeB0lTLUKNFF1470YQCYIu/I
VmTPEWFbK8RiXiawQK/wFoa2/e8bOh3bD5+iUpxh7wWfBUxzCT8gAx+ZQ/YHYA9Sf+oPN4HGRWU0
KV86bsVXAqmtKjXISeUvwKKb8FUyBYcFniQ3PApfyGIx360Bz8jayhse+k0vyVN9oH/+IhnNZMIz
im2wDk301YzpvA/jDryUqT/gbhY/yba6k8ru4vtI/2XNXI1NxgtUFe+OrEoMr9bErLEOS0eKENK9
0NT4MGGMfQ8Nb29skSn4w6FCZrR36LPyU/2mz+QL5rcRIkNKIx4O4bEzYylcF1LVnNSU+TjV4IPj
N5UTrLrK5SvX9u1UJDJLGJqtj1qn6EUz91ZcwkOJXp1wAufOO9Kh3q34FoavZ2ojmwNbHo3plcHM
dZVNmz/Zl/gAyyZxKwMgs36bSkCGf2xDlEfWrMZ2eeG3karpHNot5qKeQZ+sj1Ou/p2EnqZhfW2l
U9JfQiE5rBpCmVJKFS8ROIst7bebPODtOU+RCBsYBVriPbLPXtYMBig1BbuxhKOUYrn5mNLsD3Eh
XGNBPFzv1oDBvKys1fzHlFXJM7Bcxkv3czWgA1jan+xPqRi2Lov7w2UHAH6BbFHAFDQa3TFLoESq
H2yxGJl1RDnyud1Ye4AS3eoQtMMgkRLbkOiWsYVI7J1kxPe5NPAPk5fRcDN+SBJUGf3d/h5r8TWd
v5z5pvQGXUDM3MulR/ZBKjGEyivhk1Vf5hBTtF1FLRdbzsH4Bv4RRBF2+cEFY283k3USIlvFyUyq
vRJ8JBHDnmOwa1KvGczlcioZ5cTQFK2XrcWCRditZ1DWBfc17W7xh7I9Ytft0593c8miAORiOPg6
3Y5NdOLAJNaW++l1Svi1qWBrquRYRUeS1TsvS0O8azvVf7lBMBGqkKI3cqdYNe1YaI8lO5Z815Vc
0mnf0GBDJ5WVO+6dsLkkCPciEZdclk9jG6H6+GM5bgGdo3yJDFaJeZpcpSsAQig/7IW812xlBd/0
V9vrqNQJvDzqQV3A4NayL4EPU4tFrm5jMfpO04caMsUqXIMCtktXDhkSi4MR14OS5D7xP3cOj/po
R4oFDvuQZMaaKuNPDH2LsXa0X9jWZcCaeQJXB29xEVDtW6GZaNTTH1Gx2kfXRx7HvgVGXO1KFefc
aWdh0WDxM2EEbA3446m98gMOuv+RphQCF20bjpDo+pZwjIeACAI/yjZ71jgeNhm9CWtjznR8UXHV
RpXpdFMa37Jmrt8ogFBbEKz5NB6tFmZKFslqZEiNKXGBL8OVfi1RIbv/uUdN++ImXftlLOwKtscu
p/BUv1nBIYk6LUPCqHcLItuD8yvVIcAHkIXkIPCacrDOgjHLR3Vn0VgJ0BrJOVJCNbArlfqJVOsH
MAjfz2bH+KCrXGWb9OTFZL0zzYZwxKuBbmqXalL4BVhamEdUzdx3XukdU5IVmSCHZJVQarnX9R7T
bw8iLz4PZIdsCAD9edn1Xblmnzxm9C0rHNuWitZXcT5iAE54rgo8Z24KMH0DQXS3es/x63u4mz+D
RD7343doLoFdrMLe7myMr1CbmuJvlufYBEmCe/5sUAS/aeuHKlMt2jMb2hyDS1El4NKe2LI6UCUw
b6Yv6ZuZ7l+kEf7kcMFqzmb62f1YrW7FH0Ar2q+BvOkvrmqmZ2GiJRz3wI0fjR28PAWiJMnSA4ek
Eun8htXGiRbnYVYJhnmBtW22TRDZ9TAmhj+hxLargPeNpj2xWiidlUjLcq3VwFmN8xVFTQfQvTeO
EvfF5Zv6kAME9R0BkrAGIDqBThzB3wIAPhhBx4xZpXv0obOSUr65Ij6hiybcgJE4V+AdPp88LqO9
AObNU86fAgHgDjWrO3L0Hqff+AiTaAB2d29AgxoZehFDfkQZRd/osXY/uLpAZCk6ehaNm3JCzKv4
G65PmtFF+Cp8QdbqQl2PQo3GnTA7GfhsLEt/SxIetkzOOxXzImAuRskdq9ugLBEHzgiEaLNOXaOJ
eA25p7AeiNhIRbUJ7BW+vYDE/P2+KxYI69DxK6bzNkUIhO1GpjPRoyEC0zNk9Bk0plobFqyGmNp7
BM/Y+PHNPIG+GWeg+94J7quzdlSlmOeNDHae+DzxfL12UKxePdT7Pkha3x3eIYIyWi7xQN6uLyd9
cJD+Gh7mV+Y2jf67bDlWNuYkGySlfCPSMXYNnFCV7e9U13tsi2iw1p5k5urb6C9GGI+OVWhiTg8i
6esj1lz0J0rrqsy3X+OxqFHrdZvGSZKFqI/wv4AFLTI3C70FvLMvkF1J6d7+giT5iy4/wE+zsvR1
GAkosUBQUO3pZ/ocapo6hyICPzkAgUP4JBRRgGAhtEcO1oqgkYMSGq/Bh2ihdQTNWp04EIAm+ljv
iPC7c3Hy4QfInfOrtpUdz8N6HV+kj33tf0Js5Lw5KWrRecs1CqwfU4NThlTr4yS0LkN2CNgIlDZk
xkUrjXcnu7wQBOlpTkA0W0lZR4L14OI2qAUyxBY55dWZFuEWnk8BKE9C/G3j8mt7UXYoo/WFw61n
ZZfgKsTz7P6sIkpfxbO0dYJrCcfl1ErI3X5l8hPpftKRlIDCukL2YQ9z8aak58Q+LC4Qnu2oCb8v
JSQ5cujDSORzMuB0aPl1ZRItqB6p2If3F2bC0ghSBGVPwvrekZJXilNsMvdsZ9hIPTqCPCTvVleF
+5s+47J8mQjUNovxypSma6+5pReUrjHKBDNNJ2Rrotvq9+MOdj+SDwEArfAiFCrEFFdM003tM4Fs
6GL3Gn25bO8VFmeAxFifRqNWYvwXU+o57iw5DZ+uPy7qbyGGU13+oVTVZIacV1LnxL5YbSpwdQlZ
+jzG5eukAGt4eykAQ5QbA7L9MaN1tKkrB21cbXjpY/d8dZ7XvTl4jLG5ghoRLNgCaZI2/zH5wZD8
B0WiYFnb/2wiymUy4W3OHsvacDbgO6W32p48pvc0YpUtmzSaKltKD22PlmiJYjJLveC3r67vNVXm
M3bYajf7NFCQghq4SFvAkRSIUUck0TupSC27MnAfvwPPrL0yrQOXnnMFNqHo5rNhgDgeDj1mOj3B
peUSFLQRG550zfZvlX2BmDRZtOK7tAP3Lfpn4rdZORvbG4xOl6VKrZq0nxA4xhDubOtUwh8WREIh
lQ9ulW/nQOF9HYl9nM3TBUtqfAnmT9o5NP/uN3xJzAda+cWJqu9Y/8Xht6UFUMObWCGg/euabpfo
O4c4/ldGkUdhPsYsM0yNNGfjahr/9lUiulmG/iQWuIMEVtA15PeDdr8KOsIeDkMGcooLdIrap/h2
iOfs5x4jIzT0EkByF2EX/9qZTt4sP2BCLMGog6ObEX6dTv5wJNYzCmPTTdbSm1XxUPYUnwntJ95l
tx5RarxnnKtSR+8qI8+tHX9mMRaRtIIaNJ176KJNpefQkMnxNXaUs5NB9v+bpr5vH837krxxL0U9
FoFA86rO3QPFRy3Tob4VWbxRYeHBGkutWN5K+QV/s23TcLDlE4+jXzqXpB1ZRIbv/U42rqx1yNwR
u1DCFq0DEgYr4WUXZojg+VgTxD52ndxQnLCVhrldzp/de1hTU9Fc9fhZ7P7dYRoqW9F2+sgcSTIm
AfqSC/VAFeeUabkMpY4VMvBeajncDzsIcVLGqb6dWbSGASmZzBuqoqHI5a1pdvmqr8f9SkmcA2Br
ceU56xVxaIMWTx7f1cT9fiK4ud8bjeo+f9BYsoWs+JhIV8wFtX4/rHbTrdmTlwqaMcH8DyFkOu1n
9le+sq9yxYZ6MGERa5+4AEMzi0LSmSqqkFDNlfkX2x/uo5oWII5slI6sXElDKFKSKxl/PSOn8W/Q
I5InZn/5dABF+XlD6s5l/escJGZ6bEh77oeTnhWWE+OU3gqx9cgQbYZLhDQNXsdXpWLF93v/bL3S
jIeGQebeIApWGkNkJLYJqmW/wGr/NyoTBmZb3LXiJfpCOeMeCnKQTRwdbQhzR3tXj6honGFw9Fv5
17xl7cK4nLQYzGJOg7RYJj/Vt4W5z17TqxgmhnraAG5a8VmjIb6GpluJJkcADHp1d7YPXmbQRbLv
N1XmdhaAbbO4LC2PgD3+OEuFTB8yrefKmywdCjGS92fGp9L5CzHY8K2HB0ulHviw9MK+O7t3QYLY
oPvME79l75L6DeRhMpFMKRmGAulUu/Z9kx2XaY0R2FdSQYSST3uQL0KM4+cZaP9Ld5VBElJsBSHa
WDHUAf0kHF+/PCgUyl76TSnHcNGH7LTUT1/mvUtdUrymrScDwUED3EDrKIeP/KqNteqsqfGRLh0M
/rHsFWLwvFST9Ec3RaeUrcVycz0Xh00QXeJW3L4fewiSC2wl+TCPcXiZCdE0GSI0RNkiLaMtkMaW
PWMnw0tiswpivtHnTzgwxZEsxWmYBzmBQheXJhJTPGl+8DhTSY9USV36RI+6TMfyDslegJpesxHu
g8q2xuG8w0CQMOoK0IMi8++YnwGXpTeRlDNWLbOQ+fDEnL9YItzIgfuHcnZkHGGN7KUsgEDxpCRv
SdMfqEefcew4bcmoyi2wnBtQBo66iBtjf3SiN/W0xjmweOUI/i3a7nexkzbROFf7e0H87OeOpgnN
HTpuGhBcPbmoBvkPgBFH7xB7x1LfJdFfaCGqCzxqdeOeQINE1kKi+2+06Cz/j7hadR7Gg+Lwi8qo
yV3tjHV+ErTYSHxvGfjlm1N5NhdM3IYNA3/FGkqJlUi7snS1UfeBmRuhsnMHbD8hB3KsIRtZQLWm
GHaZm7b3KpmH0jFHkpyWdp62C03VzaXw3UkIxHxTmBFNen/9mMKzpsDsxg2KFO6gsLeWTWdFTIp2
kEoMRqVuCnDhpjTxKATnKwhaPhul6tArFIU0VXOOC3JNL5eT6r9Wr95o89zWFZo3u1p/ChIUrrWh
c+/ZOG70PG979iiS7j9xBqAYP3C5img+wr0LQUwkOFxIo4o5+XWfoN3oOKAj6FxboHi3ki1VMqon
sc9pEXdrjL5STKGQQ/BDCZITmm9B8+xJotZwgnMS+fMphxPRlbEKzvKlwv8K7T2Q8XiTMsIYzcoy
gun1Ju4nX10VOuTf/8YeConrGvOBaOaswmkoe7S59CzBS5YeTynQryTSCOyIa2JjNnnT3Ls98uwR
05lf76urtmJ1BBmTajzvLH0JB2vH6B3fal8z5wNTa4qlCG1GGFUcL+BR+CMLg+7fgADCXOLBpye1
Av4n4uHfnidLw+gyJ1QwIfMgQ95I9pHpo+hS2/Vae+O1xTMc2PIuxdqquiUwD3t6RbZo1yeF8EP2
qPwQf9QPDYDs25lQcSMN28v61xD+VEac5RYqvykSAs+NNrit+xXbG52C6p5BIsoaNl5v2wFxF4/J
7ZfydKhQk5VZ5LnNe+hdqs7HDAEmBDPfwzHgn3/k8cz5N+74kRHVxIhxQ/MHxs227lpV9oB21dTz
aGV4SVaqiB89OpI5Z2DxOamkYZS+NIzGV3CV+ezjL88ogJIvq3/8UcG4bGWP0u9mvJCi+0RbOVRG
CSY5m/AljDgiQVn+tTL+gIQsJgY8F9O4sRlBnuLflpAofCRUDVdhfDlqw3IeCL4gxwx/OUsAVPEN
diZFz54diwFSKPabLoPqmq749kuYa8vt0zc5t0ZU28YtikJkSh/qARuTDbo2mrAi5FWsff8DM8w+
UO0KvDm/g5M5nnpsULOOTTWm3LgzplrSck5ZdhfODY2sc3tuEfIL3vofNafx5xpZ+VrZZ7epDH3Y
taotTVOuKlQh8js1DdhbK7pLa+hswJ9PX4J1yK+2NohbtiVZYIV5g68/v2H5gLn/kQ4IESM58U1l
BtPXaILz5B5i8zvygIhdLE6oFr4T4dwEVWWhctkaA39RNUlcWdOIiWomBMfpEoXOkKbPVpvTaSKx
oDu9kf6+JAFofJ1XKW71PvoRDDj1eW+yjelvXbgkL95jCe0SEzu37QdaPwZgBHVJK4PF0NvcgvxZ
un1SaCXrfMFTV0yNvOoAfEw8ufD9sDfO9rCXoHJZnL5b5rrBCF235TyqVXXJ61xVQIPQsdc7VXs5
v5SKO/4Kv15L1bIachCq5wNze+CBGWhJGiEaBZ/giacK+UAxiHl30EQQ63967A4FyKmmFyFibZc2
PCgKlLGQD2X5DGWY8VPWEq796VNRVd6EVUzK8zVYPUo+cRTz57y6ScFcRuAKQbQxWrkj2eZoeHWN
HZPYXTqZmi5S25V5e/NwwE2C9N9s6TuICYWXAGR88EjNWzj1l3Vcp5pM7ExkQtycj7E6Cyghbp7I
VVo6cbEVRg55G7Ort9Uq8Iclfa4M8wBY02LFvLDWOyqhnLQ9ZRujqo37cVCFhSVLOL9xdAhOhLJ5
JXPJ741O0xgWt/EdDCy/WUigPGykR8o++1cOEY7djRbXS4iiivZ+Xq/l+03vXG9Huai+AaPaHpt4
9ic4nHXuxxHEro1ruN4fIdAKnBb88zCZ+sYgg8CWK5cIEiQAV0ZJKxE5wldiQEPPS5pfoRDI6Pl3
2e4HwINnZP/7wv3jMrVqZj7BMlCj2Yo3ALYzeyKIza9HLZ3fe3+ERZeGqKtMh6S7+ZLd/rfBT1qX
pFHqPXnlVWmPgOTlMiHwCIAKyyQ66WP86HVzbVNFM7HNg5c9UbLU5HfpfELzgyedZRqkf6Muy7kZ
Mks8q9xDImlGA8D1HQpGJ5CtvFShSHEkaF6DoMpP2/xX3i7lm7t7qHKk6zpqsu8KP3WE1FIO7svB
fUhokyxQboZZWjPhWqO6JFxxjky8eSrKCf+wJy7m0zUOXeKSXMRo/l/JvXF60NTgKHmsDsSnJREZ
hHFKXKZDFPbvidryH2dCHEQd1FcD1oelNArk0l6+H84B/s/ymvWdnU8tcw5CEo1Jdp0m9RjNcNJA
KsLkPDFHESSxzr1rowVqdnugSQNqHx8i33HFoPvXEQB3WowD26YNjyXYGLtKq5fKM3TvVSe6VSeA
pmpLlFtVZFh6k+BbMm0Ui3dxIRW1wB7wryomasBXHFOuNWtbE6nFnTuESAFW+3IyU00K1n+QYFo9
7m3WsIA1bv79ANGFIpw3ZnmoAh/105GTltR3jIwYW4/GVqQtapg8EtAJa9RhrE6tYltPqihD17nu
DRKEp+O2m/1aVXaakz3547vnJM8hvdE+y9FC+QEvyTdZCH/7CKeMJbMg/mvat3H3EnEDYaXypua1
NbQ8Syc6jrZ25rJJbnpn3gqY/55MfJuehMhUJbj2gaHw911pLR/vN4mcv4qA/gPZHHn2VwYKFXDM
M8ysOSgTJhSusef4GMxdZpivi6VgjuRu+eJx9FXA7d/U5W57eXjXIRt7i+vh+eFgNNlzPkdliY+H
ngAKdXzfSGc8V9EXoIcNiswNyCwvZE2/euAvxPFplklLuXwGstR4rqbI9OXWKkjxujDYHpHYBnd+
nwtEVkGZfAgFybrnxtg5eHIoYArqnRbfdC6q7Cs2V2W4PZpLMvYBHeG3Z+TLdlGwrYMFSnOSqytb
/1n5fSArAh4dd+fkIREEmodCd1+yZD1aYF5Qx645VEOdRczbEPaKZnWQswdcjjivZh+NjiRMoLwp
B+CgAVlwoYlMglWQ5aC2P3FbwBRz9/UqQn3l6w5GHj8sR2+M6Lf86BMpxAJ/uEyv87aiL65TuYHx
uFviI7svQzjQpWFS3ZN0BN3ZxA6JccmPSberHcfxzDKx5XVJLVqxQfh7BGwVJn4PxvKMBqnxhc9G
wiMqRWLpPqilLMFFGCEZtnDTl624hfcdIEAzFPBVMWIuPOTedOVAGigN9WxTS/ImytKks96Pdo4f
wFXobI2BDHGBfwtBbyRh7jolmyEbJJhd0f6ysF4j81Xivlm0aUPJ/ziLWnv21vn9O4MDSQjl7msQ
ypJ7dwu7SXvw9ScHUkfnXC3cKyJK48INBO6U8UflzCnuL5Qwzz1S+NGXkhNAD/hSiS/KMw2OcdSM
s1ORsUgWp76iN0bae84MeH4mjosiiNyKoABV1DXCAOFdtovN9sm8ZhUiB/CwmI8FZvQSakjbk6F+
BtxdIT+BKmjfhx8t0mp7EI8ZSscOCD21BgENR7qYhLx0VYEf8DmQ+PBhe5yY7lsy5REf8jz7zsC7
sFYAXVcBMk/035alZWYiOJWs4Vnq2q1eDo/YpIPTfXOp+HEnYOPx6p8dj67+c7jBaV0txAnKNs1T
g1kVHdugJ2WoEf3q7BJeqBb6Ti01wKgVYfVQ8H//xUBEffhB6OH3jgvx3mjYUs3VYTw5MRwZRF2p
IgLpBQ9FSe7YNjulCTzkB3xGg1rf5b06xybsX28h0y85+FYfnI08jM4vkGgz//df1NerAhy3IQNY
U44NLVom2Pn7HQAR0iigPTFk60OODRYFLzy4pphWXBRfD4q4V5v/E1chMGHfYUlOaz0lc4g7+W6V
aZVmqwYcofOnJZHCOL74u1rkbop+uQDUpXXTkcmrYpMS7+JAdPGEz+B9VN53f1lHFzfKypO0jjaU
Vs28cY5ZNcRHzU620/ZT/PwXZUDo4z2QXYMF5gg68Y4+2713JKD2xNevz999CFTR/9cMcbcSeLjP
pTzAJml9h1tPIUFa1zg4EkgCzBd5+Dp/4MylyqZnXhvCbApjzjUV5QQpkYEoe2vP+IlYXQNfYfqf
K3avVcSZI5yYwaW2aJg/gxHCha1/ly2gPPlhUqGYnKjaxS8m6EQuunBfGUdBiAwgMtvtkdWiTo4L
mjSA3fOKMSRKr22BfGxdJ9vL8IcafmaQPjwWZZ8hgh5jZFemyCd9hvyToyTOz5vo27OwKMe7KOvE
iGo8v5Jnpwti6tiq9wseGON7zbjM5SaoLhoPAoja8Bz4zog+tt8d9l520yPJ+0QUdc0F3I8OBkXr
MlEPp3WTxT9qrfS13bkrQi89QVnZ92C6IlrPEDj2sG+KL2THHukjeilRsT0qNaqMIWpBgYIt+9vJ
RCwXUnxRpbgtTaZoRrW8uYx7//Bdfmr9tCIV9sFD8al+qwfcVumokUOYjhTk0uIk05SsrfpswuzE
hC9qkwejBMCcpGQLcLJrOZUCZMYZOdscaJz043bsMvvWbeo6eLKGgfqLBvXFLe78E0WBPFnwC/3E
Ij1bnnLM0nbP1MxPIWtaNc6GbC3uiLIaGxqfKOMj3wQAJqid0+N4eeDfzzi4TzP7DoUdhrnbuna5
SQL4Ve5iImXCXlV6U03mdpAZ1xpzL0ATCXd/c7RqVhQzHl7YiDJH1E+I05IBegEzsggtM0K1+VU+
hMBxjP/yzu6+awfbeqDG4PEghFr+ebgBqfb/d3TX1WJrSMUSUDn0Tu6GTzRGBXTW6Se+7uNG2/i5
NZqCFhMZ233fLZkzxPN00PJ4dOLN3HpAZkFk77eq4aiecNDtSLHc1Rwnz4ZMADH0XTgo1v9OvNi0
hrAxukGIbb/lXbIzghxy49QhJRQDggBvFNVaer7Sgio81Fkz/XcxtApZvMXhMvMboJjbPo9swjHd
CpZJAUjo31+Q/G8gfU6BL7mL+jha1hYWwJkU0B2gmFeH992Yd8F/fu8ZgRuKhpA/aAHBMpFx3sDl
sC31OgZ/jWTZ7y3U1QPj+Tm1pDk1Id6+AS5yWjyE/JRkDBSIcOD7Zy2CATZUEIjXOSc/KpNhAZWT
BekVK98Bv/7EpXO2WslE0mj8a5yrtsbhQQQA6JFoAy6GAyKhDhsowxJ3bfIz9xIbx1RwhuDYlVPN
+PIkbdPZEjfMTyT9XTkPtZXy/rA2kzObvfloVkvFh0NGRCBpfYIy177xGXxHbfVI6q153BlX4qhZ
Z31ZgAG3aELAhzFl1ZQPLWz2wPLNslAHyOZzLFygbypDHwmPIBCfHeTsTceW+aEV3/Wgf4Yvy0Lb
a4UP3LZDiKgdV3USuLNcg4TtMoCwbp4GUIRQiBisWaAhIE+zUc9VU4lzuueTRt71+bf9vlXmRoJ+
wsGCwAKWzoN9H++JURHNVYm0qqI99At8rQu5NkyJK/7mmCaHnVebwbekLPP+WoA3SXPTlYNOlG9w
6Fl/og/17h8WdmZLp33FgqGcPULxNHG/aX/viS5yBNdKSZsIc+77XZ7k+VFJAVHAaAPKSK7mq71s
eKlFm+6kxUkAaIFicAoiqIZimgAd276t+T2rzf5V3w/QroiNuRR6xFpDojZ/EPas8sjEx6ft5AuG
slJ8Any4xB33yTJZsB6Q3CNoQ/uv0do+b0SquDH9nGMNhvIRKB3Cw5VVioKLl/BUmoYISUPVDfd9
5fcp3HWNZB6AWZLetHPbOZF9i+60qiK4TnKq+RiQYIEmqyPhtekfq0hAJj2Q0vSkZp39g88HvbYK
N6ZvurjOV4VA5JGtqtwhdsTcmWvUz52KRYSKtGhu/4Nw7CV/QbOH7Zznwa+954WDA7/gCeewBLiz
NWimEilMMxK37plDSL6wuryVqL40OSq/+aKCW5JBBVaf8HzMKghWY8TllvlUQEe558qzMhiagLJV
pfRBxcLXD8iAhKSL16U/KWXFVLPJ8BnDfCBle5pnNSvbXaUfWy29V3+BOZR+DlyVjAybuAHf9V/X
9jX9YO6lisS2fu+numKIYv4W3YorEc6QffLCymSpa6qwT99wjmnoeDX6nxVvdiemKaSV+9aBkRsv
ozEogOKjkgg3rIYMJI1QbrG2m/xU5g8bTkplZYU0V4GVkDnFywQ/R81RZg5Sc5/vlYxsn+Cn7hvx
K33Ht+bobvazWJEgN/IiEgl8KtX+LVQcwA58KJx1I+zBxnUBbUngxJpibYa9Wx8iZUeszcLWOBnb
T/YTcA85huUIvnqsyPx4G2QIAEhjl3GUyXKPTXZ1dNcCg78rSjgH6X2WkWSE7tFPpBoXAtQ8shc4
iNQWZDWc9LFnX2qc+bYFEMG7IccFawnAZCdXa+V8f5RIUTvFtJNPaJrzrgeAzRWn2j5SjBwhya6v
tde+EWXnnU93CNu0NB4N2enSVs7spqEXUFX9BA55JD+N9vfUdPSDAoibqeM3V09cepZyOOIMMC2/
3a7Bsmqr0V0iu4K6DLpnVkbxQZq08eFncvVmyYwAlYd0jVTb56KF9iiKz3/S6gw59atnPr+P68AM
cDvWEgs/cOA7leaYdaG0U0y3b9tNf1/Wo39IZ0PCFYY3awSYSD0IGaXX4qZ2GyfG7gE5deqbk3qP
aRCO1VYNiogsdAMNhrbAINOkUSl0XMyffqTYeiDRiqVmY9bXwvSYy1ZAwEsIGVtBbLD2s8rlsNDc
VbCCw5iX91Qy34XKmYgvUYkpk8ldS51rDdGH9GgjzD9zTqP6NJJK4orpC9e35qUxvywHbyzwBeQA
SORUHhVArvzAzpV3E3HPIs8tj3dqat78wQNwNt6P8qemy4H8E2QAcedjA5XO/zIvmbAHSY064sQZ
PnXumasX7jZECv2xB4fs8szJHb9IGp9DVTQ1Dq3j0eBicjtw3w08NgXBdDvpAG4hRBaavUW9Vt8H
WG59EiwAyX9VvXVOXvvYvKcZh7EeSWDteXuUEhgRvgtOyWH1CMRrTr303qjt9n3Hz0nNJjQ0gkDb
deF7uXV9AYF/x4j62MdF5gVYL+IeLzan7U6PxIPPXCcl+JEStLelynEcihB/9ZBXWcmtwOc4aM22
27nmqLk+GggUGKTBCu9mtqxMTfW1i/5hrmS2agLAreVobIHqUdMHe8tqWk3jtn6wniZ9epC0snwp
jOTTt2gduYlEgybLrJS+BPuHRhnwLsA6WqfIFUE7k/yWvjWsreaA6JImgcVUYjdqicOlf1lq/pKO
KCt0h+32UtlJwavfZsm0Kx1iDEVPeJsuD9Dg8Nn80063nBXj5mdihDPwNsCRUdz4LUJAozvFtwDt
vLATQAPkuolLFPUnIdRBJXnPaPINVvKGR1oxgByb41MbnnIS0pslDS+pgWKTCl/UWDBP9pKmrtm4
8BqJ1pp7qCiZ+N89/1IhMlyvMcGsCdRGF3OjhWb/oWp6lh+9zkxxfvExLOgL+RQQ11Q9Y21jJplO
iv4cNAXVp/X8NAdlUSkycg2qbj4KugjLBjxxCfsvUZnkQuhCAwNfIN7ghOae7tMgprYL/o+P9u6e
wZP8Msv5Yn1rScELN7st6GFFFH443NbJRbLGD4GsjFYwEF4PdsAmAovO1NGaq9Qnh9Y+98pspCdw
A1fdEa1bdGsgbYozWKNVZepJFW7sVNgHOihgDt9ZuTsNdCTW7RhopN0LjYPxbDIj99eZln7paDTM
1Ny0iU5AqWqzzIn9wN4NrZi5ftZsguVVEO+Be9798CCDDfHVipTuXqVcnqOIhjFkv/MUq2tu9/QR
nZZSPT9DUxLoHgRrMpOCvIO5/JqXCMOORva02vKoic45KMlJf1A8KG02gjDuUZ/rVl881GZ2PQ67
wzuXyXxV/vn0jscdfyzdmvSU+6HGfLqgnSsiSDwItAJVmIaVxN2dK3tV2CWBjmfqfw3/VHt0FIVf
oHq3S3KTva/0wAyptg/+77eVgxZvr4FYc8Fe5V3KEfs+HKbT9WlILuS5zYKeDLcu6sLm8PLTyG0e
FgwylQQm1g7zCsD+Z9qZCVtiL8tC4qq/CZz2TP6nJ08dxCTAGxIvOBpgBORBlDYEFiSgTfmd4BP6
INxIEKOGK1/zEfTw7RP5VZr3GRgU0Q1tQ7yTsPdRHXGVq/mpqO+v7cvJLxzbS0twlJpEBZe0quPR
zWoG/Yv/Rq5kYRAKN4/i6D3qlN/qyNn8WVx4PsVbjq0Owg8R7N6VhBxoFID0DUp8FDTiDPvZbxA6
jT9PnxZ6dNeFHA9f5LEzMrlx7iHXjiyjfDeT/juLzIsvLZlGk7IDL03m5jC/BlFWXeHv2tiKba7G
fwlOGuGaLKmHAsNyplXvSXUjYGufskmQQOHPlWoT/XTG/FgCs+Sx/YRxb1NdaQ7qmZpOG8oNzYMx
vmq1+Us14v2pRMR+Yh/yBUWbdthFedNyf1lTVcMgKLDs3woRNs304EIYdKZcPFjWTEHzQstMOlQT
d6Lbb9QOMqsxZ7QZSR8sUi34NEqbxAsNWkknid8e47et007SyiuB0Jlr5kEfW0T4b0rIu1aXHgDv
eskMN06MPAS3odGeVGizGn2Ajm9anHdZUhBfmE1HBvDMPr0Gr2YX569QUuJw8gmE2Mk2DfBYPM+Y
FqcrSquDsFz8ulG/W1xeH1I635DfNNt7aXeDff423zl/zDLGzm53/qXu8DBFbccTVhyVvriY++Kr
XkTqp0387GcuiP3Bnecf1+kPRxt7brofu73bjy1fVY+ZtspsdVbGUIHwBos1E8ys5wHBGAAxH6qR
hU04CmN3yu3QJyhqs6UL8mQa6eSn5LLm369YAF+RD3u6rYWiD+FhwvaoSMKXPgRRA4XfTF00lrZz
19U+dxXHv1chhUVUKKK1dwkqyE4XNMcjoEseu4lqP9nThhMtNd2EVPtMLSrOZ+D5hCJMhJ9RA4q8
qYdZv0gtLfcKd+FJyWJXPP2zOCn1pRQG9tEzuct2j2Ct5nwulYaaqJ8onhoNqsKaLNP+qIHI/LBx
If3iggg9Avi/E32rGbbIT2FB2XF+OvuIqvnwexCuxLnVJv2oudPDJxZMuKmz1zOM5rvsFfeto+Vs
5lxkwaYdar4kk7gc+mbkktvZsZ27HaEXL2aNK8KnhI7LSPFwfTz03qHAXqYJkT4Q7R2xBOPFwzq4
XVUzdMOKr5cZsFYpLfFaSM9QlSpxUuGWY3ONEU3GN1J0SK0wYGstOgq0D8vJV9j25dN1IE7pR7vF
njbf2FRo7AxdcfNJnvYh6avZqv4u1MwZko8A3GEhG4tNwY/Kk/Yx84Y/JiEIi3pXq0ajahsmsACh
hIRG6y2/WM8xY12sqRPIi05AVekbll8ZeBCIpU9Soo24CF78v8xOh1a7MbcS3yY/Tlxv+/ccH21R
QyJm4gDxzIQgJGxvElrheJyAgy5X2gTONKwq87HpbxpeDBWeyIHZ63DLRecys536BXe78s/ZykHq
3zY+nHSMuSp5ZZDwBBDdcxuyBdYySJrVYoY5Ffd8OB91H+zRsHGHxYEqdWGtlgTj1Q0eEK/5KqWM
4LufG1dw3WzdMYxERiHyX5KkPZ16SEz73RK9eOm4mFE4oEJ1/MKHpgWkxcQ06ftLu51sP+CzgJfd
KPThIlGCwu/IEa8KH6/8gEtTO64j/UJivr5ABV4JvLwapAZr9sxUWcTM5cdrFW5Y4+wLfc8h4f9P
Iar9K5OtW1WRDTHefcRI6FrYsrfJ2/nTTuFnT/VIf7FDCNb/Z/ahT3xhzkmOOjCYzqO9dWkK49Em
PGvkm+xZG1vop97xhPrIWzA4F7IP7NCpEhPk3BwCGwUQ7Ce5Y/pV5ubtrw/Q5+AncxEsfhxWTHH/
BgGJGzj/RvLooA7554yHMOeia+dbP0K6kFlq3kE29VLf8qBwgICZ2y/CtWnFm5qYGPUU0QnjaKro
KCD+KEAMGIrII+XKzvAUmQcEcs1rdu9UmDrZ9R9IZCB6Fg7bE/6OhfztgswEmFM4hJMF/Ombmb3S
YNjKyCSu/hjn+EkSNvEhhfjLg8RZDNISYSdb6BKUaeQxIWkp6wg7puuOi1BOCo4ykSMuXffoBi6Q
Pl2U86BJTeh6/XPSd8LqZX+3V3xyiYn1AnHOhpNV+9vRcKjFrxKBho44LNQhQbYjVBzBnEJMyOuN
bk1ZIr9SmvPSQUIpA+W082qsxTuNFM7pEQqpmHUxfiIP7hJbcxI2nxhLNY/SWDYErxTk5vN3xjCb
Lf+LG1+HHXBuQwhj/7t3iSl6f81PBgIGbnQh0nhMPoy1nJqPxUrBWxN796RC13XBQmNWmdGTiAhW
BAJCWpI48v9SEDvxJ8asXAyqvw2VtGCzktYer7QleWZ54VscOHD6A1F4X9fMFMJIxw6StFNyN0my
d14nHGrA4V64mUz6aKZIhNc77cxwztQED5VtdPQ8DcSf8V9hEgqbcIzLrsx00Gbq6C2blw8m0Fqu
Ql7f42GgwT4XDdmposUOx1+4BEito9VNMP2jizpET/zjtug73+CenAkOY5j+R0xnc3Msv1vsxX1j
vb9bUnRv4SoY2zNCUeTFyZ2HlhvUwCOejGwaOACWAR4CGxXMpe8pEi4A99oeeMJv6YaQAnkGdXYK
qpxrVHGLzpHnr7vw78kqfXh6f5gryKZbDsQshQWIXMzDQVtj0r4E2S2zPz8wkN9y9YlPrtJxVHnd
l1lYg1zAVhEfdnikDncZxS9L62Vu2rIbL4qQEysEe7ghO+plbeuVjLkt3kLFAndRmx5HGccWbKKH
SSMDqu8TfAaXCXv/k29XsoRHg//lXFU7ZEsdSKRM3E3ZT5KC2ZoZ2WZWanXqwc+2bw6OSExIT4Pj
qTuosiO1cpkxUsy3EUSghEqc+mpfPCTyejSEHY3lefEDT7YPgnvxbylKOT+XkgKWJMgVHFS4l971
NyEppCwPF1MAek7fQ5KVfkTEbbGTLAIQHGeV0p5fljCfr3PLxW5vw6aD8cRuyvJyF0YwHdaEelgx
j61YJA93KTiV+BCXEK3b7a4LYZWMXwNXHjuPmIYvYBDaebU0z4SN+qP0R6S2cR64QVBLLR5VF0nj
V20ZYCFNdV/e0fqN/IMzJGvwiAiRJoya4Q9ASu7YSgUyDa+SWK+noivN6yi9IXNrFOIzI3oygKm9
kiHthrIOLi5vgvtPLPLRR53mjzhCZy2PIVF+Yrbmi7YdyG8TsBeZc8iKTYmbsycBdhRD/5h5I1py
7OKHfqDaj5MZEpjeQZFXAy+J3tY5coJksAjhgEvH/Gx9WYmUIZQIitrVheF/wulrlvrh7tlgfxXF
caAmF2zImN99IUD/PQa9g9vmo1CtPGrbxH+IYZuAQ2wnt9eelu2Lj5oluWvauGtGvsqt1qiH+uf+
lMUrOBpwRR9wGyddLRwjVonX0vcvmSi3onS0orYC9u5q6Gj62F20WhWGvs1O/1l2CvgoXiOrorAy
FpE5nEn5A2yJPRosXfIV49ZVYBhuT+FokbYj0Y7WHmqfwYB3Jg9HSsaZI5mxOnY0PTxe4w1kQHve
eZVDrM5/nA0yF06hgcU33xwqg7rXJSufC4KeUJ0DGbbsgnCgHtaeg4EFESOz8A1HC12FIQAzy39t
Shqk67M0XEqjEG0+T79aGng8IPMP0ZTyglOuFW4WdbADsmw7dc/cP0NImw0rrc3UzUDQ24xYpqjA
h629wdSTz5WV66vgAPM2J16CnjgAINIBBgU876JgS+VTHrPcCP4ClqBAdWXE9gKAzHIhIYfInkot
gRbyDhAeIDAIpcJiDjoGxqAvJMVZau3MJMmaPTViUqihzrKjYBwgF56XuzrLWQduDpXCQSERBn0z
aA0bA0M95W/hiCNZ3iFxaB0v3BP+vWpC6cndIafWrz+VmWJbP8ekSdBB9OmmhApIM5XLGeynqnxU
6gneBcbiaLYWt0g//RDe5DJA2wcvi4H7x+eFkaEsgh5NUg/SozLDpiuDGCyF5g5ERvO2//pQLxtA
17dm5iKuArulT1rFOyEEIcJb8BjL9mIKXauK4jjzine9XgiKmq/C5tJDHQY6fv4JebLRhgWXrrLh
LWUPJKw3KIEnjII4AkQUV2xYbjM6mzUEwOXZ1NOymduquPhpcUjPS7usPvaD2/wkgllIqwhH2OMp
nJLrGCaDxGa5+kAFdjSSSCfsgOS+RHn1U6uYc6KUBilLwMtDwOv6O4cNbzRvnb4tso6AmsQ0lggn
kxL0BfkXDHnYsdyV78s/h5otwtHL9YJMGsUWKvXWGlrYYlAADr2njr2igOlZmkgOHyfRR8/M++BU
Tk0K+g8Hj5Me9tAJ7n2Io+db8DmUpOMoAHyBN9QgG7pwLsXA7aYIv6l94VeziFXIaFkwwFNWWVFT
nBbsJPeubJ4VZKC3QzSKPX9OFTF1BtUw02qDQYUc3ZqbuoYQlxpYTedyIpF+jSl/kape/FC3U8iR
yACLVupCmZYEoxpfeEAGARxXvtuPRaqJXWTdPgni8N9odLKyOjsv76WWGTNwcG5ByjpRUQNXmR9k
FbmbFzrjscTpujCcyK/2gUbQDK4B5hd80iDzTL82oIy8iiTr/Z/zvW6TyJNQO15c7aLDUaAEnYvq
7CikgDs6aZL0Q55j6ImST1KYcP2byJyJEvYYgP4+6sU2vWRp809pINXWp3r9UC6YdHSj3+Flk7Hm
aZVwzp3QUdDDuAkzwZxNaMAcpGQzz/G7cvuFzGOQAsyHNEqpPOOjyKrObpEDCKOTMLFsRxynBcrq
nOuv6CCogLc5WtWUL0Pm2Y/XWoNwHaeb4JFIVNkgBiM1hG7WUljhaU4fy6ICjEL6NHqw5GitKMMd
G2m/9N82TFXfauHWsPUWNAvMt6wi/dr9rijmupHgVAwofJHN3T+cf0OqXs6dUqe3TRxaMwun3Qdu
EEQNrlhyQZeVqi42pSNJWqPkY+HjyN2rh3ntzPafPPpXrONea25C4Qrpxd/jqEG6cESRz3Fc3IBA
FZjUky6PpBhs3ymanySBxTa+8Ok4j3pUSC1CPEh6q5Idu9DoLLmBBELON34SIlRRmziNXN1T9Sx7
FZUtce+xBzfmqShePlRIh1SdN8+oO/H57BFBQiZlxXtjLWsxiriqUY+gInlbM6JdwGCGfNqjg8If
BG7xG0T3gJx67TWiykym6PQLY/6K9QBb0Y2hd1Qe70o/0VEj6xHMSRLtg5yNp93cuHa3i+u3y/O2
nlSW0o49hxrIo2+nIH/x8ru1UQkFUJ/dWcghAkWhhCzm+wPpeaYlDuZ1OWTaE3qOZGsktm7cLIF8
u2y3bz0rUggS/T+Gzs2GUvUtKHdP6k18KFGqN7xg2av08Lha9TgqIo/S79XKRJShdxURM0OXJwuq
fx1dJvusvZJN1bdiQDSsRRt6q5y7oOHQjxLSkFcv2e6XnrTJdMKjRimoFa6cCBlCGU8Rvf6G6JMW
RlrqqBDlTyazAPtn1ydl7LvbeoZaSVInY74cbGhfaWBO4EjWHeX+7LH8iewe+dnGVaZGE9dhl7Wo
wfqxUFaOOMDKnFUayUVFznAvSpkCkuzCL33YeweJXAAV3dbAMZnu7JJEu26YP7PcqNa/UQPrZ26j
nTOIkMI3ox7/7ik/DVBYsjDMn4epG8F2kMQ7tI8vpZsidUYjWWp/vzIu2+ziNy9hOJ/nfJL4mnWW
+DCBxYWB1RJzuWufnsmUZnGiqh1gLWBCZS8MRjFaI4D4uocvnzttMujSY8YJDyRyT1FG9LFBAcWN
Qpcb55hP8FgE8xjCxLY1hVCidTg6MVjW08QGfSfWxvkYK83LEVkqkUpOpFtDHckutpdNdebwgbVR
0BETgYCtUvRUJzcdoaOOcfn7a7psIgx+Qx6WMbcxRM8hZ5bex3omAAbBQrqKO6CJPdeEQhDLNhrc
pEPMvixwe6dRJPHJelVGVrTHIKf7yw2tQwmmCqt11pBpzWWD1wSWmv19/qOt/+q9y3wZH4pcGJie
b6JK+mIwFpObJwLJuGaFwVKcjk0f0QWDydjLPojAPALwAH3zExS4O6fKZG6oPkBOX5A+3fnbBkdE
VlsdNvzs0WsJbbgAuc9bAGqy2wKIXXHRBekHniPrqf33I6n2u6oYchLmZ02tSUbKlYO5yv5n05sG
sEcfpy1rX/ZOzoc8w6hfX/QOvIHKVWeb4+LdBHA/TIkTQVoLvAERBDTT745CeoOnPCRJePIVDVra
wSlIEtiapwJK2TY8iR/nvlPT6WvC6a2IYUZJfXXvr7NI7d31/DtU+70zraOMo4fgMcBjZFTKz3TZ
4BDNt/jYBrHJAnJDKyDoCuQPidjPCkD/rTopMm2g7fE1ma6vy5WrCyZqbyruPLuzpCjGrNdLLfZb
UwSIsOmfITTtVjzFV4OPRHT37pdMRFqEzeuDg0zFU9tR2xTd2tGvqnP8K1K6ZOhgr7MwFYelX8V0
8EmJLO9fgmIdt1QGWCXPv11PSB3u9C+zWUpJXDWgPKTiiXd0UyypcAIX/ylXdlniFVJsmj3xHd08
PSHTcKK1sZoosydipCiQUdJEJ7YOHJbOEwpGGjfQLNLg9fp4p5Nzx11Y2lg/lWuYnouw3kOjIpy6
kSgIJmU77J7BVXM81jiZ4B2IP4xT4DQmozFibfQcfw10ZzrOvzp2ggwjvKcIlf0BoNePeHS0H1yI
6/Yl8VquLhZtfrEqQmUwvX3UfHdZkpKcnOcB4pUWaqYsNNQrL87pjJvZtQ6hiVfjGa81sl+O4K5S
f0fd8RdLLZ1n4LS0Dqq9rLIoIR9lqmAoi6Js0uto0BsRK3EOAx3GI+Y8gkwfgExhWFOnUExDuCDO
1Ry4cVrENWmUnbpBV3DDLX806GiSXT0MOWn/uGFVIOI7SaKTh26Yu+9GVSCe7Z2oT/FZsCclt+s+
T5NfJGaEcng/5RFiG+4Ijxb4UZYXzfVLjvkNwRBOlPNC/sE1u0mzKNxGwTyTOac4NwNJ41XyEYVy
7G2qSWm3R+Isa+PmrmsLWYsHtHE63S064zAQM1M1/SUwyF58+ViIE/nOg716Rqz3Vg8LQxs6M16M
IxiM33LOjyVF3AnF/NAjhcBtx2yZMZOk9CzP30U2KrqgtpTZdzpVRR9iOTR0tiEAhG+sueh9T+/q
QDcmirzuQE0J9dR7tLZhlyclO40PtAdpcqnP4CAlWpiaDO4z+Dq1ohn+rmLOlZYZtWgBgW1VesnL
cC5+SDwPQYFWL7nBTf2+SDEamdacNiiXaPsrQ/coOZQKA9X8xPXRAgo7INXriVhe/ILXeUGLrQVz
J62VtQAC53srXQovLEauW4QtQs15UGXjWKmIWrPhPVz8Wy6iIEn1K2EZEGnngh8Y29TDq3wwNRa6
Aypn9o1SpnRjOC7UR6nrgrxz42MqNRUB5psCZR/x1ePA/t9nBvyvp+rtV0Cev62qG0bU+iQivRn3
T8d0DZ6QQ947BOnwyIMM5gCmgBE9qn7DhX6yOxPGULr72PALyWr1KBVGEjzviR30bof0JG3Gzt2n
oqPrWfMw7z4WK0opktJSaR7f1UX7Yk8Losfp2AHKAMVYWOEzIJLDzlUmx0N8rkM8P5N2Tk+P7E0q
9fz9fL25ouO+5cFuSxWL7DiIViia63VglzdPA2fLQC3n+iRmOkBeNOmABqHmyBd5QfBWD6qtttfO
02hHH6TSuwYL9ujgif5oGBfTFxQVjFYr2FHMHcU8z47b4S+c6oLJvAelPBCdmNUMDrxY6s3E4hqo
/r21j0/uzsYs/FD6DIQhggrmgAwQVa7ysWLg+EzRkPTutBG0oiMr4AzKfVNa2maBwAjI8hd851d8
FOI5hzYpwx0ba8RK79tlWG5B+z65tesH6knxre0uES4ArRAyan2CtugDY67xhV2UGpscT8egHDf2
ph4v7MA7i8PD2cku311porZ6L6JmHnR3Z00IKVh/Msl2Y2dxk0AfukS7g0BXo87jJMKBbgV3Cgx8
gLaHE/DK+NA4MGdAkNUhM9Tzks0emyeKaQz8G6HG5M/Ff9G5mPr0UnVKCYbMLo3dWPsmKWQbgv+2
75IoI/MKmtGD07SclbooW6Zh4hACASGhIcfZXOAvx/8s0TPBAoC2iMBuyKW56ntVYtRZuAeFQVMp
xyL6X2aJquOAiZZyUtOQmR+9+znqsGEZfhHJfARUDuTQrFvoAK2YvdYckI8+9nUSzAj7oCw3MDX1
GGjFqb1CpFkcSbSNMrAYU6BB5jbhsrfQyuKM1Y7Ov4ftp/Fwg/jz+sMNMLGqraz+trXPdT+xMXqC
ZbGEkxTOfzuloJqKqdpqDH64NmTGNDUqsWQ7IQhCoEm0a3VZLZMz/i1eM7i54mHmJcfa6CWz489o
HMwlHX4dANlzkOtXVb5bVKYYKP4CsIYdTQLnHrMqVKegdBS12+XgkvmQRw+iW1+xl6aKVmEdG4MW
kopa9CDE7yIuwiZqFQg9SOjlPj230osiDXW8xX5KVq4z6k+bpw+dkZ2Rk+SyWalMccTvJbm/CG/L
0nFjBH3bHv1TIpqDhB/x8GTnpNMknQ8yaA4TjzchrDyr9BUSIJ59QY+sTlDiuGtWQDUyXF1kwnmn
dO/jmSyrbZJ37kGbInVU8Icg/03d+x5lhthqkPNiV9MkzgsC9XR398e85k1zcnssr6doq/M/Exs/
pYygHXmAu2tKuY9fesRaQLl2ZuUtloyP0ERVHIISALRsS/cmu7czswPOg8fiMDvY/fMVQnyx77wL
jG4lIWdnCWQJXLlciJCfywge7HzdRo3Z43qtaOmP6FRd6/IsyqaEaUlwhEi4+JRvt8yyJLRdGCUB
VpvVLvlnkzzqeNDLb+MSYcQ0WOSPDYtcLnDKpMJqnyNGbAwE1+S7AzSnAdmHRK2P2aQ4DBuCI6Za
rYPYRQZgBd7Ajz+xbsJ2AygUPa1nT6c33poeb5cbUtxW4ecQR0X97xDekRAcE3j1s0P+SfBChCkI
v6VloIt10XEcA0b6Nu67YaAhO+NPM5tKGXNBK/eR+jOLYZI62kHwt8VzimEWUVdV1Y//uuwfCXiM
tD6p6eksjOCJoEJgOPWzZYT+/Zr50vrCsApc7df4ODIYB/AyL0IhGyYuxlns1sID2qu9O5j3nKi/
mSGPdhW9mciUAsaeFZshSlkVkz0JlL6B3Exy6aOt/bD2BBBUzIf+GJJR+cGG5jCDH/LsEgiNGyuq
HGq1m/9KKFqg4HEcD9dxbkjY7oCZzauGN3msXPDItbMexug6k9SbhIMzRHKM/HLniGOjM+Ky0c+Z
PRLMrsTsd3nNC42BKFTT10+KAIHX2vXKkpzKd6FVZ6A1KIlab7SqCPmydDBQHz4mxwQqHhGUDmjH
4Mr1bPYhb+7I1CHhZFmDpFJjGuwJcONE2FxrXAQtz+mkxAQGlOOyE3/ltmnAXsaG2jlRAKBpvDRj
fcKjVBEtvpb/kqg/H4liTsIdef8BkbpCSCCXu2MLta/sTOpmi9lH8aGI6lZYVjqRDhb7SiW7Ke3s
l9oWpUK8aCehXyCT2ndvLxBgZLvrwH4Pta7veJnhy+r1SogsexKHCm+Je9Zxzo6/NXdLIqd7TJI6
VS7rKY1WHTS77oVg/hA1k5BM/mnrxoa/xacIbUBn9Q6PkQujjsJScBDsT8D7lKSt+X9oPCJ/8owd
Tv90IeB5lwJ7kz7S+eFo37wTMoVQel7Y8W3Mp1++h9x5baARCKOvLRpIN1Jfk3DlcFMkxT9kSKCY
eVnMErgbOjRzg/i+G/q5e4a81bpOvCcGXoscwDQyNJqPr/ob8QulxjgElHIGK25r6mhhPv5DdGAL
0FEzPK/airktapdUBvrTm7eH8mtMHHFsd5lk8Gs8Lo+pzP1c/y8N72XOixlYYyKPuyWxsyYkNZ95
W82lFl5IFLP04xG2HJRhloNcOpkjILWRxK+MoCPYua6fWcqPru49up6lYyel4tUG5W3r/Vhjid6s
MFvWN1uSwguTc8KFM1aI3hdE/1U+SVD6fkuncskdvsdU3k41RmQVABX9i/X+9d+JK1LK96mTsNmz
csQuMk8FCSVV3SQ341Cm9SjXO0PlYdCmsvJpa7ncZbrjIW0kxKNneknVnICOWJq/cJK0GJi5zoq8
EiQjJGfCPxzim5g7yR92Fv+hlkVjYS3PBkLnmClKMv+FVqiwcxr+TrDkhaa9YSEU0A+SZjaPtvpo
b2Uns/pVLhyI9R7Zq29O8fj/XtNhHo8xPczKowpCSfHJmFzyZHpmORA/cwM4jF/3jsPWI+tD6/yA
evldvIBcRxoI10o/35jDWkf0fCKt/FWtCSPfqaCCxNjGJwzqytWS0DIpDkPQAk6a1Jn+ZNwhMHfZ
yOzrTXMVEWo8/mP5LE7Z2oJ5vVDj9P8mBA1ScnLlbVIApSoLrI0u2kSAXSzKCD0oxdpgZI4TzSsK
0Saou9BnNIK42vK7PL0t1rdzrC1/9ca6+sq+IBeC3fRI2+anTHDG9pfrI+2O89HCPAreEdIMJ5tZ
hkF/E/meR18JoTTww6eIYnMOGzGnvRHPX4UzqYaktzBt3wXSXp7IVFuQewFJCoCjzW3TZBjTtzC8
7W8RDmF2WF6v5Q0+CaXjytOSh+HHBopLpFtIJPD3U+h+gdUCHeCmT1TxhjtkdBFENiYSZqHxuQm+
dYj3qGu0nzvHoVl9zt98ll16UMnPzUZegP2g/+anGYC8sbKD5uSbYh1I8zh4X0zlqOt5iT7o7Ijc
+73uLK/acTUP6sJupzwsIrXuwmC9q9kmY8kfh66J3waK2ry5bpfT5KWMmU7dwhyW3N6utOx59EPN
C6SBLNUrzMRvR3qIeh9sYG/3MooyM1ajofKzLt0hj2rqUps4WquTukBBj6x38J57HcXwa+QoGXXi
quTpdHPMKW8Ha+9rzoCWQTkGGup0BLmhCx6YLDzgVLKvTKHgFSE2D+wtBZvzHIe2KqXw1uboILO+
qC1+m6IDQC3Nau/8A3zMHJg9oKKw73TICI0Bj64/zkDsV0KL8FevYdxWc5it/E0iXqZBJ83Jbhpk
5b/gLckvkDv1dRHo29slNOkyWNauASX/lRSSO9dplBfcbDcc9+gDhWPxAvHoRigewsw1yqCXRs2x
L6QV2/cxtiVic4n9CLsLXJdi25KF12WHlAtpKeNlytUgSCiM6S7sZSUcESiK/dakajBUtslAEQCw
lImCVdTZVuXf0umi+4ziPZEqW4A9OZIm2/HOuwxPnao/Wz6sE1bY3HvdhgVRTxbbTHj+yQclQ9rx
Vv+TmqdUVKUlFD4599xSrxmT3f0y2OqOea+eQoSu9VhlLnZZSo750k+mSs/2v2VWvR6adHVMqLha
SGFHGq1CKdEj7sygQq8dKx9MRRzZQ8A9cHWQpyxoSL18W2OXaORH3VDc9mnpspmVMii1sEqS01eu
Tm8dmvqLMDj7kN3WQopqN7vypuoaNo9fd4iXksr77EUJ3pem4k1QAA6HI1KMaEKxPjUYa8GSpGUa
4fAoSY8mIQAmkJBs7S/9ijx9b6UTQkK77myf9imMzYfcsfZ5foJWTCZLH63Bu7A3Wc6HXM5uuWYN
EXU+TCPGmT+BVH/AXSEgrr3oPogPvvlutFyfh6S/hOLA0+g8BO34w/joyrqHOWkexWeCE4PdiZcA
t2H+B3RYgsVS3pZBNZn+6CZu0C1zmEGmEvMCjYhOp2684dMYra7wYG3Fkh7JzHY1K6YqzD2WYdF3
BN3D4nsv3tBRyfxKjvNTEgrJEH0UpMYp51AxSUCcW4BbnXiRPHc4QYoFMr9n9QkOAM0nUyrsAQc9
eEX7D6ZuuWvvJglyRp+LwgJ/Flzt176o+7/kmIaosPWYExQm0Z/kooYsfSfH2+QFBK+3AfKisMrk
TWZ5PrYrHPza0cCIdc0AkY7Wt991eKzwEjhE/PcJpp4ixSayrlc+r+1D0tdbNivkAjqNn/OtWf/Y
2MnFt/juS03MnIdtM9JHHi1TYi6oCyyJyiIJavtFpk2n7Mol+GygZkq/tc/XiHnaT6nejQWUQ0j0
WDtombPN5lwi7wMSpXh5hMon+k1DpBthGUrqRrQgS2YwCrfKUfKyfSqXMSG0QarTu7b6JwAhcoox
Rhf3nG0/fQR4NcHZ1kiM8ODmEEmrp7HqpZ6pIo5Oeo9ZqkPCU7IvkShc6c1C2x1hoS0rmCQqkyoG
gY4kf4JAQT7N/ssbMii+YuYvoXSb3v4eRmuw7WirXfiZ7D0PjLxMqFO988DBr9lto9SLINKyfDs4
Uv/vwiOKfYJaZ1xP8V6yWd9LgCOQ58jdhfOXDPX1AyMvZxv/7XmNdQUai52x9ujl4ip8wDzqgyo2
PkEoB54zWx3+PHp8nvgIvP38dNPkG5vTnvXla3mZza3oyF8JzYm0lrr5iiMuFLTFGlDk4Swwadrm
rq6SnhUzHCM28aaOBSGidDvXWIe3mkZxqU1ssurkD1uN9xO6elJZS96/j6Dc31chBcKqjNtgRgfT
tSsAaVpd7gSqDf2zAME5P8BKAtAb1//UH6i9P4DzsaQ9gl2m86ns9thZGT/eW6QPg2oDZpLOLUWH
T/jI7UE/4MUurcCB58FdaQ+bGYWtOVGY4Sk0fKwhIgVY22mfQODQNn8r8NGqeViBh9E7T4IpFPOY
8K/rDsmACWT3/9NniDQY72KP9fxgqjg9I9B4nrJfora9TeNqFLPtsdWuIG1ZLXvvsMTJWwnI6HQR
vXiWSDdPPEX8i82wJ2KinYzC9MZBay3m1t2VJud68Qnd0uV/GIKrhXP+QzXfoZifHrzp3P1ftrCe
f0ZtBH/0cv2pJUg3VV5iPICq++dsD0fiLqTep6WJzrllU/llVBxJtEwyRqXOjmxN3lihIfFHw2PP
DFsZ5L4B5IKqFyFkK9FOcOzIKbyPyud7jm8wCYQcvcqJB2BwVtdgFqzX/fqFehsprTPEmilqSep2
ngGnwku8h6HqWeCWMw/NKm6U4ck7nwPCEtPg7EKA07EzeF/Nd8bRxy6li2ZCLDzvoPIBN1NFJIxu
K3H16R0DRWUPn0zv41GVJ/nFIp53jX7iOL0oWjpMH15ZoRnrf3iVUvwOIsZHUJJ3a+mfCCFNNFZ8
XoE0+iNA+kbSM3pSFyIJfP8olhHGH7hszIe8qK+VWBDRlI8CDV+aIQyZ2CIqjs8VDPnWaHChruiA
T77MSuaJoSoxDVrduCMKOsfLzMvVWm1uafNX+6RDj/m7mC69gr/piC8XnHNp3EVXC5/D4jCz0BuP
FHvykpWYw22xYSPDh2XklnN9Tymhq64D/56sBUlrjUEbZ+i5pB75l3SPj0iW1nj+oBfLNZwnR26S
/htsmP63iPFyZmAKQkXV4IHkborZ+ivNrOd5ZQzLDfJ0KD7LIs1OetjGJtgVbGdHkYoG3wSkoaRz
ELkw5YrUfXN2XE+Y35he0JZnVksnJmCajeFMA6u7jd2+O5TS0twbSB4YDonXFzNhFqwVy9prfZTC
sICWVhGoHWp9z9UfXqqhqCVYY9ssS6H70LI2jF7VzpukIUJv6JgnImqZ+39snpAB1DRDwMsQSSE5
LyRl09UwUMpkyV4v1egMcJJW7zX4s7Lb7Pd55UsJUyJ5mQJxLnmG6M2DoJxP4X+5V5Xz9saf3JPC
k83FeBYeTqkirEhNGu9zTWRR8F4x0C0yyWdEWA4H7WBE6UrpqZvqkqCvn2Q4F8jnWw8GnQbJTEHf
awDym/f8hQV35RbBgD/PQxET7vO9aki7RVHLOceDtV042gEOYnH5+ZEg+iiaCLuOOMc42cU7id7a
atZZD8lQRFDm/uXp3yLn4lntzK99XMbRdF7+dHM/TSA+xxAImoBMk2T8Y6ZINGr4tjlcoCe483bB
Q5j76ZoqpAtmWnAmFyWREprlfKgz1zgc0yVCkKjJkvZFpbRQLGLdo7JCaWIxibxOb1Kiz3IJj4Te
6UHE+8r8kF3bvPOYjDNlfGm8IoPcPm1R9UVcmcntztVPOeECfqdw8FqKiBU0olr7Oq7JV+OVXi8K
5V+qkPkSzFGZflUlJgFX459BxRCxsMW9WnUiv0WmI3gBFYfFqS9PhVVwgYH1RYfv/8XBvVVdBOzd
l+wNINAqvmQKwBTgyVd/N0suwXymY4wUE7Bu0QA/pRoAvRvwRwOzaxxKvcB9kuzfAJzgnx2ZsYzP
5OOn9cdNBW8q0UwcsAZ7KQluPIF7Jco1X0AfquYWR0mEazWKodjKfu6tDtmZD6FrTRIrw0fuDIAw
ZKpnR2pEoaln4f5bYrUGWee08jWLYYWeOlUDFcWZF8AQl2lLa76bhpjaw7vNu1OxT6yQ+NMGU1A5
JZpm30HL5gI7f5DQ35nvKAUKDy//a+mf1TFDyEQCZNo+rNZd3Z0j8Hd6GLyuikJLOQy3JeMsIKU2
xwWYRJnQ/rQO+4L7YmB+0SNOC+Gd+lcxatQkGBKaiodJYX98QwWpW93T7oLM9voHcZJhwy+bmYOS
5uo1z8U9TJ5WZWKxNOfDNHwKQaNHoRORSGJdTyT0SA84L544722UvgE5VFppdI6ZEPfmHz6nwiI4
NM33hUFTYtcQmWUt9hNsrSjaiH4/BrfGC0ONgzxh6v9eO2HnRtzsOvAWNdChDMyzn/PT711zT7Xi
43oVWcUhYcHEygWYR7jV85JPMWAoN2evoLOzxC8kJTadJUx4zo16T2QzayruKmrOOHyl4G7E795X
nr2OEiZe7CH9quT2sVnClRBh+wbBzsOGz1EGA30qTsz2x80GhQWbj2ISdgmvB0nZa19jn8y+SsKq
AezRjdnr2Qn7/S6ySxX8Sw8kxcRiedvmorgErBJHwTMQUTHfz3lBXDUZ+OgY9S3nSGHeXv5IJSLo
sQzSsYROk5BRhGjtpZzwOknPh9q4kXXmOCNifn/42JuppICXGP9/hPWHVaDoEsPKVZmekUza3oFW
VilpGZLuILWVkNdRXSkHJC4g5FWczSro00K7lP+yoz0YIrLgOCRAr4KA4B1ybKGFebjgTE288eEF
3akGswnb/S0lsiIgul0xaWZvXBVQVmrdWnGCNtugIx5TGVG5DcBGH/XEkiN5PUwMzgESMqJ68p6E
cFqgOt7YwltpGBadUZD863uN5RmzwCr9C+NiloefHGUyhx8Dp1u0YdhAFaJKZcsjHvoidD3IHlJ0
CX9qkBaPiRDQ+Jx2AvOELLU5qd6hIS4JeioMD1T85n22f1Go9/0cEVQ0j84kZwZPB9sqEOYtsb1u
7bmuFsAV5iQxNdj1kbfnFZkA4GMvF1CjgTmNY63eDw+5l6w18igX2UuST/mh3M9RQuw5vze9+m+G
jl33tT7/dwCpnfBOX+5z8tW5i4adPgF1bQULAgNMsnPkbz/9Bg6NhmxG97lsK41NSw8pqEtJUKC0
2YVDF62G4EzFq9fCB3Qj0AGzrYRj6PgD3Z/jv7KQTlmN3OO3mgZlMo7oLPRgiOa//ZMwfHjSi/L+
uHA9TtcMx0sTTTuVRbnOwyuoTDZPc7Y0pJsHnFYYQKXEngVoyk/y/VUCD1ijTcfNxO/kHkjMCjWH
vcHdYLDzgDtKtW5Tp/52NskI0mUU5DPpcZ/dmcAf1MfM6wINYsnwd3UPiFL5FnmsfjODSsGyYcZG
NwNvfnoaQK6pTlFOz8jIea36t/+y80n43pQo6kNtCObQ99KEOGBG0z1SFYbw4/YreHFeoGAk2hPV
3ZtX7rJ2v3Fmp9sDfnyyQ1mU+2QGU91OnS6hNKyPlGx+kdTIfC0F5OrMiy9ppLLtCljgGtzifFTw
gzcJuNQ+IZ6+uiN4gnJJ18M7pRA5WS+5fGtZ7br6VOLRlu8njpMek9Q5vafPhlRY+v/BMmDc4Q5H
qn51z9lNHuwYFaeAca6tViyK9tGG3ckHhD7zrRsIEXT0x1D8TK0OdIMF9sjE++JSZeo4JXJbHHlo
IGz6Zo+YqdRRW2lC4VuZ08mXFCdDHcx6ed1iO0a3T+ERGG5YR4bJDWtt19SlLCXLhBmYitEo0c+M
Uozq9OQRQzg6PzBz2/Obnxm4uaeDjT3Xf/SEIBYVMv0xglEqpM5eUfvBn0iCNwgsE/BnN4KhUaEd
LEbEKwQO9OR9z+o4QFncYaecIkffOpADgn1Y0oDprdNPQxdIjJGxryGAjJ85B30VirAKDutlW4zq
4lwRQ/KZ4w5pDeyfF1ldGC2zHDRB3I11CgHfVu5sH6dK16CJpwUTgLsV/zxuIOUDhg81ZWUuFO7o
NOpePIB+KWMXZlzOT5aozXd5W3Utpew9Gwf30lTLLIvESQ6smqwSRUQqTEjE5gBKBh0pEkE6eGmi
tcDT2SjecRC4vYOn0uSNHLwKkivrJ8FzN9poTxOHQurdipMXutXTGtxDcqM5XwaLqlgWE+xcxMW9
n+kP5FCjlxDYS4k7H6W80Jm2YFaZh9fCVjuCGDJtf6EU0FwzLuJvN6b3Hm2KidzM5FYG1+I0zL4h
0yRvuFUjLkHcuwbdH+eUsEOG9hPPpQzaFF4U/L2ITQulAabooHPvfhdTO1CZYQjIfuefXvcurBor
mfJH9qgKe3RBGcuF/VLdsAvcp2mOCwHXB2SONTqqIk8WiX0iBdEy1QLSlbYJd7ZZll9aUzRVHB+p
3suB3+g73YUKIw++3nRmNjvIooRDP1jWuAqej9ypbVs9BQTScM4Wlal0KU6s0WvFZr914IidnH/+
qgpgg0u/h9DuhxmM086pz6NKgJxyJ49wIo6Pr8I/2WEO5xs19kc05nnwJrV1yc05ChIqPS2k1EQl
bca7bwZLu+I4mgdxhpH9e2tyUSwGbomp3PZ4xBGMU1T36eR83YVbGW1KM1Gbzs3isysTlCao3jOB
IF3VoyWDrSqf6ifmBEyerVZlfgJpBRWAZBy0/hCMwHV1H6seIF6OvVc0x2PbxagwM9D6kVq3qKwQ
5/3n5owAHsYGqWd7qXfjOiiRYOsjpmVDRhhO8aVkH6MzP7NMa8uxdf7DNIn+PgzL1oJUFtiFTpTT
c4XdnKN7zsTTl51tH+pU/4cKEjvf0o044zd0V/fdcYpN9JS1LkfV1rwqpeH+FjZDE/WPBsAbtfyp
16LuPc/VBAUHhRFJe+2qTsO6HursE2a7yFTzjo2iFazP6MiO5bw2kLtekFRe+3yR7PnwjlLwdg7N
/vVGQQBTP3/Mbe88gv2NNYToC5ToK6+QN2uuDIgcI4/wdfJe4neowEr9mN6/BHLjKDDQcEGBFe8w
zYyjDsRbIwoV2VdvjFPwoCrl/xwHiDg7pfcxPget1kMp5qD2U7XBnNGs09FVUBb1bcl2CrdswIBB
rtl10PwAwZ+/EA4UFJbwWw1dCPyxlYi+wifObnHY6SAv6b6qWZU+yBw21SafH1et4z/Ox8o7FyyL
l4d/qJUsIpxrru/TFHQEKdTT/vp3G021asWFuGAyncKI8xl1IpUDA1YGjD3o76Upt5MtlSLHtztg
UdJHQggZAOjJxhiO6/5pIwf4/vO0odWIokT6GkBu/tH9fj8mcvv6iRR2Qo1jvkhx5Mrtws9b7+vD
aP+9fZyFcgJDVIIqiZ1Y6Z+HC8ufmMk5k0+Zs22k8/jH6PHyjBhK1CmJnsWbwHEFnoR2w71VQzaf
OtUp6+u+hD/Z4Q6f0g7m+86JTQB75qvkk0pV9kmt/f+tFNdjMH1yeUYE4L3e0YjbDB2DKZAdxq8R
VsjoM6uauzTd7j/znTSJu/SMPk7pXF5e/UsDgvQVPKwJFc67IsMiqDsrT26XwVd3QrPB1ijIVEoS
y4bLACz+wn+GWb2acgCdo5SfWQkZgtHQCPVC4l/TfsERpFtGcESZpqSDLYgtXJY582G3+lqkvmS1
7bM6zW8bx3U24ixEdJz5GtrCUTmoMz8K0RulJiMrr7erqsEYFRYmkMDOluDDnvcOY52fhNHWvJWs
zwuMki6i1qzLxUn6w/IrqJJds/CM3W1erS3UGJt2UTmX4bW8ZI4Xiv78u7ujjBTJOVvjYtw5rO1b
l+gKnta4xIA0VxeN8TksyvN3/weux8qeckjNYOSO0iRyrFyzXL81AivMltgC43hLcPIWLb9QdxWb
aySKjVulel91n47twd0AYV5yZUt9rGQTR9vUdSvQcJV7pzq/F+nIus2gbdv5xxITOMDkL4aOF3yD
m1NZxDS59JeNvJjIMH6z/6EohCi7zD+eDeu1/c6Hued2YX/+OcXdHSycEijwm5GKEVdq6qE89U2P
Ym6i1ih48cPAqrtK1TGLsIaMcp4w7r2z1Kj+FHLH7lX2FJsbhInXxvm7UFK1CWn6U5FeZkFbOCL0
zeeRqtSZ4bnipQqRI0p2PXkbLQnRWUpYwn5CXlSaIzf6ySLNLdCqfz6LZo2iFuAn3One5CpIGcZc
/OwYv8X0ZTLQLObd4WwfeANjBsFHp4YThRpmNpvoR9hKpEDnu2js5RxzgnRZtDDSh3JjXsRdBuLb
jKsu5u2sOe4q5HAoBvprLfY/kw14bT8I2JSOeniZ6w+cKRkg6c6S4VKSsqB2VTBwZkQHYmaxeKij
QAc8ftuqDQKXYYrrtYB5U8qFNcTPr7PLgvzMXvOIOuqdtf3y4+mGOmsLNZ7335U/tnaYzH8rcjyd
I4rtHgDX2jepNGRiF5XrIhvffDN7M1rUOiChCFG9+qMp9Y+y13oQSib3LvAWpj5921Cgx+sKLFe5
dJUqliP7iA/zQ/UEG5JbpcIRy/MZfVAgkJxlRSveHEZJMhHRtCjmU1vPfHZ2oOAoOo9OWx3pYVDt
Ejxf24TUu1sJLj8sBJ69Y4tx2JwKb1v1Xk8EJaFjRN3U2Ifz+h40Zd7+qTI83P1Gn2bSqZUC3IiF
3SDJlnW1md1TUUDrCqecZ2QkD08Hb13EvkmZ7DN+4D4o4cNrn3owNYNKB0JM/o4MpKKr3f1LSlDf
Fke06DzeldJurMRo4XWb2Z2lbL9p5Cv8XFEork8N44cYvA+pW4spGZmUgxnXvHUguBdWN3MW3Zah
DBJOcj9DfLOayn1VW0f6SaEMS4EwvQzIUdowHx3d6Ovo8G88iXhssVSEKjHrLkNdGLnvt1CGVjuz
A0pf5GyDFUaWtgCK8XsJOhZl3foyN7HGwwqkJ2A2pKE/ct5aTc+X2bno5MwTX4c94VOdmo/nEWlp
aRR5jd8d7TNaLbTny0SWwHzj7EyT4pzKlD18wmXBnO0wXCkJOWsYK9EWY1Yahe0CedSdYAv6VxYB
PENkczaxCRzKCQi8P2snGe8C9/FjVSkyaAxUahlzu3A+ndPK3iNe2Pj5Rf7oFucMRcY5r3+nYUIr
GYJiw69yIXO8dEezahmd6PO4mJdqPrGStn5QamRHAO/NuaI4uUChy3/A2Xs2iVc9tUTE/SrCnypO
uKkJe4Mz++pSbMbzVXYI+moQ39s43jcm/8HR5PseFqPlyTbIhKwU+K3UfJvQypfdGM/jz+t9MgLs
3ZT6RDyIB2EHnTcPBP3OwXMjDNYD+GugMdvu5Ghoe6ezGcpZAFqXSI+EmJsz0zWxmar2mi3Xf9Zx
fAShgmfeps59z3cJPRgQw1gSkkFMAoRIZ+t1IDMKha5zw54kWGI7OpUuAZ0xLBcMe4OLwcPnnnms
iqlUzAGOd83qd/StITvzsJXiM+gwE9TYuHC9KOSyekUU7APMSwmwFy/nOXJb43MmOFy7PianPSwn
sF4zaphOtbd3FAj+/vjX+JgAffZ4+eWFCGbxShRk1M1qqhnP9TbdUMEsQ9ot0JwfzB2vUQ8XZe7R
cmaauvwLslD6ksBEMk/gDTL0A4QydL8G8QeNKgeEdTjfVjDNrd7GzK0l00m53V9YH0MH0c8UPYrr
JFZSSZdqyvbUXgviIYfuWobrH0qNEZtVKlDaxP5uOCCtETYAjpM8hFxmeAKPUNxQGmE+nThTLG0Q
a62QLfPro8C/GgWeP/AxhTCYv8s8Fy3aC3Oqw6s5t/H7So8Ol0FP9Q863Wx8QTCaUnNzCbyYOJSV
4l23DhAwNMM31+QNe4kj0e6M1xxGIUjVxjD448QUnzX7zqknFC9eR7wWP9sZehSPWGOTTcfAdM0j
NNiEGdtNDhoj+3X6vd5rMwlo8qPN/6ndBBHMxB2QJyTIHMkLelLSmvGdccxfavfX7cMdr8rTlYLo
DZWjz6yR851xzlrT1yPiBypK+BSrstcu75iMJzV5oYzR1oFWBYIkKbj5nCMUa/vzWJ4xAyNeApfd
sySRDa02W7puuEXEPVevqyNGsSlWA8ZpVW/FJc0zypcyk/2DtEe5WygZK3lRG/tCDE3guTsiw7a0
U7TeMvHUWaaHc6CMPinZMQJg4TizPig3R1ACRE65SzP3g9GE7C7tV0FQoiSMVkGfH5DW3WqAjg+P
Vt6yJWQLFYG0Cnf9UndlQKUmr/1iVzczz/4wG1tE9j/Dax/uoWg0KIy/fpdgyxchlKLHj9q7bBEE
/gfWeMCNs3xdiGY8xFTz58fB263ZdfI7AddQk/6j4iVxJy70un/Fo+Qxts5W7haY8cFXSYP8sB1/
u0Tlo+Be0aBPtEN/l1FaPlBhon05i73EzZ3q6aO2OXtRIYLkAdqAHvmXyzgkKCk4prbUJCCHDfpC
kN9Xr0vF5IG38Et0k89PebMaht7iWeSeTUFj81Cr8ifrlvJBV8Vc9ZPotbLSgqu9/p/GE5+zzZHn
Nvfo7yq4LONTHPctpHdaf2rJ8coKDCNFsUqScg4Km/4XHagHYFs/LqYXKfath9hj00DduvBjVwci
DALXdvKOb0oBI+VC3KTjGwX8ALDSLwcWIQUMMU+CVufl2yTeaTmf34CDhWfWb3wtPodQU8Ojg5qJ
EF8u6276Ze7pGqHtTfSi3GLKYJ8Rn0jXyparJbQJsS3kuKtEe0kuagBlLxTEU9k+q1JPCM7z/YbX
s/G1Cj2/xhkP8/Gpe3CKex2IAx71Lh2Z9C4KOmP26Q9V/DfLfj9d0c/vNpmuAt0bU/uJGW/BMp14
f5pb5AZ5sIOAPbBCmFkc/w4r6/H5VQwS5omOa/i3dLwF9AxjBAQMf2OH2KeyC8GTQUmjTTQDBWPe
ZnP0fKoty8VqJJKuvePJ8GSfwzgpINYjGAtWwHD9E0eOxq34HKsTfWZLJS9/rTTbDr6OWRPh498+
7jn384FxSTJTrHIR8/aegEiKCUD9Opc9fVUSAXT6ZBazsQu69VvxYSaFizlTRXxZSba68CwbUJNq
hzUuK0Ea/xcIns0bO4oTISKgoOUynMENz0dYnw0ZCMvgwTt6rTHNjvWvcdndkYWzk4ny8rf/mgSG
pU9mdV1mzaTIj+VxpKM6HjkjcwGzv13Bw2qNFOVjlcu3YTc7iVFBAcjGyAc0jh1jOy2+xEc+42CX
xXyDj+6fV1DZc7Xc8mb7DV8/2ZWXLsXPNpI9RQgDFFWOR8GWAGb12XSeWktF0jRu7PkH9Vio9uli
PrSzZqXU5vqYBgrP55K1heXOGOUVBIg/tpTeuDG06vh/xx9uS8Mp7U1oVVOmc7/3fEiDWn+YF6Ft
cJlK991ElbOWlYXLke2a+GUGqxJKA88jG9R/APKi3GzWwoum4Kpz/eVHXD0qJpZIhtB9NdGSr52m
w5+mzFfnOYBCAoevgJxtFWNLt/pF+5VCHsI2vURE1ATZnuwbw/SJqH+ClSuIh3h9LoolvdufDOdZ
wUXyKhJ2tekvjU/+AwmT3bjA3Q4JpHNDpP2t6LWI519ehVMm6HACEE1BMPUNqJcAjkRnG42Myq+1
jYajshBwIzz+2IG5BqClAWUmBC30rXPO6XNPdnGXYUQIN0c3XJGjt6/dpcRSDrBh+4nuQIKTy1AS
HfS6tEuSkigFeBYBAmlYNo79Jip6htTo9E5Nq0pKLCEsdV1foBo0mn6Pw2KTNNeaH3BL7DCpQ5FT
9nd0I8mC7ke0Fsdv8byiqqdxrChTpdVsRKk31KBT7RGJEatMTkOwU1bIbd3+xGFtiX83Jzi7r/Ld
rnKF2erKfi2CgH0o1wG8RBdsObgvv24NOoAchyV1oaOVCaAxZDhqWaH1w57nOP/fgtV63o0gDIYg
eqSAf/4/m7J9wjHo1+WQDZP0rOd2KtKxKTXvvuW7H7ZHKRbmWyf4ryn1S8krKfSnkuhUk4QJqqDi
004IT94jhDecTwb3k2wdJfLFPZjJG8wEFBvgQBTOINdJaTZfAddUZt5P4BJ8sU7pR2VvFqgmMZD9
3yLPdFGUp5Ve3J/B8OIaKw5A8WfD4e/L6X2y1cvL2KdLq8q24PYEsqmB7STBER5sCAek0eCB0HtS
jUzlZ1ZXkCEM35W5rGlgvKrYervDfKwGJKNGym2Um3CQOXcBB7R3jiZUv+2dTN6QdOGEfasRHdWa
Zj8wJPkXsKgCMU+APPclxCDWqS4QjpBKSL30R0Qg1SAruxPwGgFkEzJzwZpAstTm2N/qFn7PXCu1
ONQxYquzRIhkUt835PQah9wQ3HoubrKtTshTvS28WC7DKwRQS+mZBaYDd8tB18uYwvVQ/QKAJcUz
dw6pogjYHm+0jGVazL9d4iH/3h8CaDvVc9k0ddRHd0N9D/rndnM2CZ6h30rn6xtnjYiAUyvVeGAc
8hbBZ8vTXFjTTEZne/FUKcXsufJilYHQS8bFnEw+85JUXDfSxwjIQYQfmbhvUBC6LB1irUjiYvcX
RXanJuAsxxyHiEhTjrskq46y4YmB+Zyx2IWEOyK3iltQnDuqg/8atQxFbMmdaogtdymfY8gmd8d+
BxPq9EHrTjm1cLdSYbTFDTPVJfRM0GXtnSWyuLz3mu+SdsCstUZUJCjY/5g76tgVhCnAeYcM5lDe
kwEiLmfCKSgcCO6awEgUL9DI+6S61QQCWTByugqgkI6VvAyUSGdhgOxgR1eeo6JZleJ4GTWcUtrt
0RJWgFacvwQ3buvzXzRc0GERAlU6GeuB9xIkMPx90RIfLy2jZFK4dq1uGhN9eudmliMoRa6T8c0I
jLuYC2m0rGjV/ogb2qO9+h0KsGlSEv0ElE2xrFyumuvygJuMfzdxRsf1jKh11Qz/PxSCDUXsFZgi
VtEBYcWvkNRntOixnyY+x2XJSh0llspuNm62ILU4GoSHMBPxS2qO2kor2FVQSeoWjxWQZ0pjlsgS
GI8a7W5SSr0xIdbYUaD/SQEmpH2CVBoUoJMWv9CgYMSeBJgNYmNrWH8x8GpLosQKRP+JdvMFFmIN
2yKZ+UifW0+TPKlfrbClz2LZjJJWyrxnjPzV7OV7h0YZARs7lo4Q5voPXwUEGHV0TkIBs1IQ57qT
GosTLHdlDWYhEr96Wxs1k5/L3F1IHG23O4bvMnRmzmduOAg14YZXumqDLhhOziCDCt3w3XsT5V7D
yjH7sR6u+g9SzSfUJowPvFuy1cAZ2g2Sv0xqco3AjlY5lm1qVOBRVQg9TdNIp6wzoHTbv8qsYAdh
rRGNi+V/2fHHlFjl/02xdcJdGwhMLj+8uqQWGKvaVsyUXgyP58fYZAI2lvYbShj3wI6Uyvqsuwmq
QBSPBs26QjdvDu0b7CHIdRTvsmu3zxf3v1qUbO8KsONkGb+VtowAp7379pbj4TbkHOa6cJR4QlQq
hgKmw0ErYQaK+O2wvLNH4OSQkhr0C1StehMboXxm2qWSnxT+4RPunSeay1I7aoBwHBBi5GEAE/fw
tNSTbNHrX4X1MpAn7CdJZ4i8bgMfgfE/30lhNugjkAe4DOZhFf+XFF21qFPYdbkce2VJvVddc7aH
5GuSvA8psqC+meJOimNw5++80uuIgvczVFpYgMxo6n6C6wmttgsu8P0oppPznwf/FXMVnYTYODba
B3jaAi9iBXS+p9qJ7TrAxSNpteExQ35qSE7FwFtuYo8aTwGcC+HF9hUWkBPSHOOgjpm0AM5kV9s6
i9mcqhny/M4jaSu0o1sVodNGA32dMj9Yqt6RSV2GmK0e1VR/ZHO0VCxgXncKknAY2ydxOrveXZNc
og/63BW/FgKjtuPEtOxCTx2E/lEDV8rp6aRmNy8XWSyh5YmlvoVKQyxkxrjFi4xK3ui9y7rCj0I4
JloSC/XSMCbhPmnh45b3Onh/hUOoq0hXq6/cBduMLv/wuwH3p//vyIK3tJBowz917ywGCm+cExzW
StS2gDP/oM50ErjmaimdvzJn0eXsexTLFxPAFBikztInaKztpBH65TRJtIirhSiHhckliqhdgA6Z
nGC2E2tBwttD7RIjEFgkSukdsikxOdSAIDQYcf1c2BWj/S5hKwV1j1EcDw0uqViMg8MwOYlAPOeO
DRHxJQRa0dTgXyFBBy1RYp1ObDr9HiOZIsx5+MPiTyfLOxavlPVPzZfWebiuJWb7B+agjTZoBxSb
bjzyt9dyqQF+XHmYTbljeaqxnNFQGm8QqytBh19sjThqifxczjw8RiPx09RHzZZgqVrvU5n24jl5
aGDS/iul25gQt0gSxmeXJuiT8nhAomMb/biWV/NPijnUvnT4K8q78OozZQa2g++Kmy0RbCkReOfP
O0LQ7tuX5Qvgcg+iS2TsCv4RNzyLpQzWvFK+KvymSGsgd+2yMqLWLulkvx6ER2iBA0FgI3XtKVWg
VLmE1B5hgQl+VoVWWsRfPi7WZDnC1Z8HyjSzF35UN98tDmkdAb0wiMgPCPkSyXwQ7AUykljH08rb
hbBXa69OKYZRcpWKV9Wacigco3Y3IGAEZ/JvDTQCfra9tfeQiEZ+0FM6a9I7Tuz4QtQAn/FJlefz
nqWJUzqmMBHOvvZj1DKf4+ZMzGLjbFpujzSxIjm/UPPc3qRUbK9WWevJsM/ZjTtipDe70xzW5zNo
17vVXfpNhVhtp3gc9khtMBZ0iS6OpxlSqLPT7OY4ELbY8jUNO2T9TFCYgGLe3vs13eYwGTkQFHxz
R+BBT4aKe+YSYiOp7lpOpdyFhO7C4bVVCjueX1BHJHUyJwlk30Vb62Ra6pJo2N0U5bA7ry2HsJWX
k+s7eSdAKCH56+L+g4yIGu8ncosSwXSgGJdauCJQc58aDwfeuJIXEY89NDUYCB6wa431yeJ/Kb/G
ktFGkcFaPC06ahGgte7lbwE80KVQtsGlpTFf6izZn7UPPlc6cvmsYvCMA71W7QXgExj3KSLZ7pxR
YOGQfpW3B+wwtCYcBeoVOEQjcNhVQ2goKRT290U7f7Fe3ojx4wL7d2iFJD/FY1vKc/tMXMDuiglM
FBK9wQXeA3D0iEV/J6NMW6VqpGGSVPs9CVHnL1wguO85g5Sx+GFCRjILwmhJxTIPJap4mZL69P1O
5gKVx0WTuJz7XlpQu6v6BK/1DFoSAfd0qu2lxtjWtamCgIbWsSSodsqTTlZv68f7RUgS7ME5u3HZ
/uOnNPgFkjGz2B8szOEAN1gqwXDitnCsZKVx5T0Vq/aCRb14XqP/ruKKNuObaWeHFEvKhXGyr9vE
UG7DMUfUrfwVEhEYzA2X3oz6roOOmXK5ZP5G9sqPkIFMX7KPP+36f2Mpiw2QLpDg6PXRtJfAcki1
XiSRkW2rzWKHPUbynIYDvEKjTfHtdNbY2yro9jzozyFB74CHvuRAJiddovtADNXAFh3s+YlLuxaa
tJ/+ZdUiGwmkJyp/CKeswX2wsfsx87zERrSsme2aH0bHbClCICw4Kl92qkQvQUEAWAGT3RClr8kS
I+spvhmAyiXP2DFM+kyoo6a6X37RxIlsEs3xpfc7gKNKRtUWQFG+Jw+gQMrWphTNkqLXgurZh5s/
RLZ8qHFgDoKqDzZiEIdxrV31q6KmMNqSXQcCmwUODOKKNCyZKPcnUIgluh+e35uWGkkV7TCyBg0B
YUGQfarBXa4jOm8pvVJhRrL+yC3of3XmQR5b39MMt+d2Lu/hKTbpaNcxdI5/rGh+J2oSlwNmu4aK
nSDLgUl2I88GOTCLWL403GhCswTCWf6DwyCPB9vm34gf9BAOM/btv4yrJKKQaWbfhKKpMUhyMVUm
IOhiAur3PyPP8KyAhRUQS68/zamFkLdNkIT1OV5AhOvyTqWRMwwsbsbABk68XbVfYrLbxDhZoLaM
k4/ZLkAV89QEL/7DKSwOr7GMH8W221ZqPWdD5UjzXqF35i09zJ31LmPXAquaepGUXmp1rP9SBWrs
BsIGOWBdKQ3XdBLR+eVqN46mFf9gcHGptjcm80/mlEFwkSBAoI1l9o4IG8p3GodMSr+wzyhj+OWU
GK0rsVu15o58RGFZ5Vr/V8/91UKMyseiWnCZhyvui1P9NllaTWSc3XOXktoC59C+iNayDjpDPEJ5
ZPGeTRAIaQr1PoDYq4bk75LKLSRc4UUT5GJBuF1nwYNJG2NXUih3mFX1Gp7vhjeK/Z1hk0na02qY
ov5g0/k39OqnDr7fmb4DsYW+a6BAR/puuttCe6ZvD8H13vVD3Oa6D/dPnA2meUyaAB/wZya4B/0u
6UTmQPHzThVs+8UMwErnCESEpu0CLN4RyUh8ZX9UE2XT9sVJo18Shd1sozWm2aMlfxv4wZ+0FoWD
08Gk+tdDhzdswH4yBjz0JvONwO6gjjSWp9eB1xVP5xOic9EGWGdonNQJXTLpKYQcZgmEvkxoalIl
G3cAWSNS526HsUEheDDBXtaCh1IaH0ouG4vSn81wWtDFSxvhZx7P8gTMliQoTpaOH7NbRLZf4Qmj
AaKB8LK9usGnOJoOq5BeLnN6DbGiY4FfW53h7WLvEv3hcVfiJgH7PYkUGnqxDDkiHclRjSTDQZqL
sSB7OfD70KWC7mbsi3jv3OeSgyb0rpAFlCrgnrtvf/9lOWcIjOjwUB3vmJwlpNKM2jyTbuPB7TDB
kfOV9q6vf7l68mun9ILHV7b148ZerOAlfVUXIiBlc7fX/xCwpv5SXcu8wQGEcPMpD16ngaT3yEpA
a/ThPxl4JU6HdqinkrP4CGV1zrX93bQzg7mI9APIpms3WzoQvOad5GP32s3UMTt7u5mrXTTE16nK
Y+GCGh870AqFLle4i3qk7IR7JeILZ1H0FB8P0sRl31Gybv5QahRlwgIwhVld836iB4U1bGPMKAMX
CcapgbpW6tom2rgudC/oiTpiyH36byqzRq770cUJqvJrTUoB6F2ovomUUplyJGP9Yi9vzjkTA29i
n3b/w+p4nmHE25g+SzU7QbsaPbPzasWGli7GhHChgQpIVpTiNN90o9fHpDSflbc0C+d1k6moZpg9
BM5lQGwcjkGtOkA8OViaQV2UICkdJLtRe8nMH4tVihSXvyjld2w0ePCVn9sg4TB1OOlCzkU0Q3df
vyu5we8skv6FEczYOW0y8biMBGnJQjAORejakfgUSW+wjHRzqg2E/SwNDeX03rijQLxpSEkEhQyw
fet4ICaq9aiwKG5mupSdgvofnO2paaNeMo1ejcQbfyEuxkhR/A1q2Yl9i9Mk4eA0ED3Auut4IA7o
tdMH7BQiqXN10+U8gWK4qmgFimP9o/XK19Wb/33irqIFWvzZM7UG49ljw1KKrS/jEeYQXNNvdYs0
VP1D5ML3GGWd9uKeDKIE+6dr9sOyuvGG5pM2/BmOomUuLoaUkI6qdwSTIJfOTHRcfzgzsNTqi5zK
NYMzwdHzJcBywgDWK8DXivAfP9KJN68iZCA84jd15R6SNYbdmjQ/JWTF0/37fN+PXarRCETC2tTy
XHFED1P5XgJ/ZCSzQj9E0rrPLpjtm6Wtvrc9R7lPVUukjHMYx5BfkFyfi7N0Xpy6BjnAV6GfYx8t
VptYNw3YBZ4kJ7jhhls1ntdll1L4XbJld6ANBC/q9tw3YOSnNAHWKtYd7eI+cZbEglUO5Cmw99sQ
tlRkJV1wgDZ87ScCKDbU0UIHHLFAgt/Sf6W3mxJ93A7bkZta7tmAgrba2dQnNAcFsXN5dhkYHHqY
otJO27Su3yb/JzDRR83veZkG+zu6/P31de4s1INh82FEBbkLl/nKTaYecdYjXcgjaAhpVbR7aGMI
j45ZOaencArPEn8rS9sczzvjWJoH+f3JzmH2krIQB0isiFlhC1SHV6Ero3F1qz1NHymqLaq8Xl2I
IM537gthz3cTJDypNJt2GDfxVZWP8snr7ZR9v9UOQ0hm+1EwskrpoowbSY/HOz5RDMfvbYR/I+od
V7XJoXhKQHg/hWOecTZW5FzY7VBsQ4uLpiDh0Z/Ehs+XN3+uJH+Ku9o/9b5dTIsQHCa2cRd5pvlM
BDTEBQZBdWyrgBxT+RTEbeCMFT2PpdTqP0KqNhvJwsWsOKNAI62q2I3+E4CLZAjAMVq8Szl61WqI
9HIEZ2VZoXBtHzZF/MwrCGNeObq1eXD0zlS85Yci4+wI5yaWwmrd75eXnJv+tFr/mSzOoafcUdWb
1Fp69MVbFdrEvZ6/dHpD5DWw3atecUNEpsVKeBsrXCzmOO+G3DC2EqpvKP/cu3dYbOYjDQWhG0d5
KeBAYGkj8UNxy96dfP1C8d8umz8MCyDuQFabbyda99ZYUokG0+vhoYACWu0G+6vbW46Lwgou7CgZ
ZgUZvyzwa8KxOumx1dNxuVYr9nn6ch1WB6XoYoNYuqY8R16lCbV25XiELtSYiGkE1x7M6l3Mcpbr
orhGkMlEyAzZEOUgjs5Iqr9O5+/GEAB2FSFbpfeGdAgd90yidXeSHnFnY03GDo1COOZHNDeAbQx1
7HzH/x2NUFNy6r8Ce2Tzgdyor/o30udrHpVSAX/PUZuxCJxctB3RAV7+Y6Y/AUJlKmZHX+Dk6ss2
ypM795RDW08UYTZod+3sYNqdZCmwTKbmzwFU6B9VKZWehOkAiR0eb1nYtCfR/titemDZsx4QOCrS
Wb5xCFzsL472TcmYY4KPJJxhHsHyCl3abQtWOXuREkzt8bz8P8KbwBCgM1KybMR6t0ECFUNwvFSK
VPuwW/OinFVm/7kSfIW0toZjgb+u35EXWUg/16o30w3JH5Yo9VXYP9OVoItLOIqugzOE9vOcBYrI
M2J0zmPOrI79tbswFDcGGu7LDKG+xQRRGYxhNLekWlHWwIM5mmf+02pGc370zlDQHFQosQu33yh2
6RhWTIEer3XkMnlcR/z0QPvhqBevHf2y9KfZMmjA71JvUGNTN7xkTRXuN7voI4GDwaigmOwIG7xk
IBHmaH/j2ng5qQJzBxuL3a57l+RspP5020j74cx7hjccG8o/6RivJCiDCUfEtjJGI7YpZMSAAVFZ
cvQY7GP6C41t7AdUxkAZyaHO8KF91jfeiGO5jil0Bo2Bo4p9lOn5qOaDWyoFYwCT0ZIWGwu1QzSg
kL3EICzoG46Q0rrWQchXSzjb7zFLkXYnr6fZEOdq+U+RWIFpAlcA2nq5qSXdw610dfTOawNSHQpJ
vhIkErOAN+6IG312MKOmj/g/jIaOP/XYnCFw/qgXB0HJo4zQ2JGB20uD5gguMD333+YFPW+elgqx
iFJwrq53BqaOqHz6aAERb5oR/6ZX1jT4aWXFrN3AFroNQpdMUWtkWtJaGXEnEtclaioei6V0SwWY
9EQpkMwqsqiYjAA679Y1FfHfgn7DDMSMEYV7ROBDXniCtpTp8bjG+cdx0MghkpPooheThuuT3YEY
6c/qXSSFf5zf0iJaZSTqJSLXaVDmSjubT3FC79zxlHfNWPCEZnz3FbqNoCdK+ok7PfLV41khSHSc
CtGb5gsaubctLUHOB1BguCpnr4Zo3Vfeh8iUWd3lhy/eBdAS5bqJIwLcK2XSmGVOFrM+qzdSSveV
h63R8CKyEnHVfktKMUk+GwUzly/doGlQOLSHpKlumRgj2EC9UUBbh5hq5PM6eEBq86OtYzxouF4W
8jQ5Jca6DYkRHQLQ6Qe5kVpP1FJ/wkktbm9ziBti9Fp2gfgSv/UdVu6wJXQrXfWTOSgEZTMP6ngU
5ANF2W5tj7L/U8Mi2dkwoJL8KnmWMed8QUirs8vvZyhYMhxKASHZ7zf4VXo9PO9roAPH72M7mZhd
VBEIxpADVOiHJQ0vczRwonrGroXgEZRmcnQ8j+CvtfM4zambOClMqNHFALwmDQWa4XAPwLWwY8fS
hZDeKw+fqA3bsagnrfGgc+eqvgO+CDuDOYNfJQgjAsxUKlBg9WsZQ9Ke9y+Q+GQwDA9hGaXnIn81
segkaL7hlM2vYoFTabEXcqR6rRCpDWncNvUzkOs3UoCld43WjF2b+cL41EyVW89jBSiup9CEbji5
9kEiH9LXhUPi4AWCqvbhLwa8l89TUkLLQo7Z7erBxocdwRYaM3EfayQ5uVd6jYSO8o1Q6uKTvCsn
aITWPRjRAcgVLuTn/Ll06pCo2e6mEBoHtH8wCjwjseyiftXFGe1ZAAcPtz/y1as5PAtZ6VdW6K6f
BTKOzc8dJDNKba25uhdxF84+8qE00KxGlxm5Ah0ShbGLgt210GSINcgWrnrfBm4r8a4vFDlQTqrE
iTDsLzy5boO/MPwK4/KQdx9WqT6HfaDoPXwT+4AFhC1WcQ9UIkFxnNyTIhnijiA91rDPO9JMYkT6
ZWFV7fTPi42XBeKkUqfCAI+Jmy2mQY3fMNp7F715+lr66wiswoGSEvrOGIDFFIHmJlrPJdGi15v7
KiTCcRf6iBaw7/hL4t/NgqdMVmrrW15dzdHz6j7w6rbORg5FYRmJcWc0F/lG2DMRDQL6F2uZTjPt
INSmJZXd68w+ITuTxSmT14v6gn3LMTDuQlgoqgfiOI+ijmYzuw98RS272N/ozD5EkwbCwHm6PkjI
Htjc5YkHsnFzgZrDs4DU1lFYBCAMt1ZDHDa+wxTxjwfMIFoerqh8ArTNOFErl/uTwaSjerwf3VEV
tYRdp4yG7FZu0sTT92f6WGOfkA1bfv1Qp+F4cB/2PwCnGmT5nREJ116A+bHJZ06EspK1MjP9Aon1
RhwsPzGlrhZOo+rsy7VtwikaQoUjlUIkRVQMcybq0uad+YnFTNWaf/ruDCLALfVWrJOeTsmBCktR
ksFnrKevCsG6B8OdeGfNYGMGO3pW7dI11DYPOz7dv7SvO3ftJg57ZlF2xggFZRB9MVe6TX30MV27
/wuuWHpKfNVGbDGFrkidxfXXZNR9sXxGXH4Qry8XeeUXMg6CmqARCyMbwNKLe2X7+Bu0XIo+8dZm
RMFgWpZlyec2bw5op+sABsSGrHLUL1oTQINBeq1pecoQa03xQ+0FAdjiXWmw3g+xjDogh117Rhbi
+ntejmye9ypmSp31GUi91t783MPT0mcdkH8cMxxm2xChApFH+ZWR6QqT6x8UmGGD2cP5j7NNfM9P
OymERuqCHcn3P62dtx6cuQpGZD99L6AfCOMrw9mxeDJDSkKWeuv7BStqx7V7RYVymyKnPqGYfwDa
q+oUHK5gLPlC5kiTZP059M60WYcejfWt/OS4VW52D2tcyMZYHgkMnB0ea8llycVNzmlJVmnhlAM5
8WsFatZxV25oOWhUV5SWvI2qc5FJS4oYrkM1hP75w5z673xlI1aIZFXtnbXNi//aBtm5US3BWI4N
Ti1ASAn6iqJAGZ+Tdw3KAPFnkcBkb6mYoCVVDrJ+HhARtfUszl++d47QKSTuoa9Q05QFNoF/KF9k
wXHE1zfdKV54ERi7UOwfzRwOi3i1PkYrPMmW2JsGk6tYiLankdEtPy1k/qyTyrKxhOsLK1i6jwmy
9iYSNG10XPxaDcmwLvo4RTwwGtu4vfIDAWNtUtqC9TDh5U4I93SagIawJgIrWS+ZvTogB/6Lc1wA
d+BfuhOIu+etZ8fDtbkfVqWiTo9jfGW7aVupMkr4mHp8SncIu06taMOlK/V+sc00/36pq4eFi2cU
PRkeJ0ci5x7biEQgL1hGSVrjEijT9D16Jzy3HbN2nC/TiwZ5tmAMXlD6UPebKx/fFuhCkEf6GD9I
T8+IQGsB3IInmwPbjdy/fwTVm4fdJcRW47U3heyBatdDBs9DpTJ22VRs+ytKL7McsnAmepDjIUvE
r1KpByNKEN4dWG2PUAPjFuU1mLzOGLjBsBBmXK80enp3PZS5uoc7p3xGpEOQCRL6dW/LbZqai6ri
x0K2tMZ1DUIlB/dx5gW16vIxpio5JOxdIaOm+oCJB4chHFHnV/pDFceWFC+1ynnWeZzGS+co4TDB
TftG7L0PfcvVs7ZGA7KVdS7eqfo96IDNUjDRktj5IDm21k5f8NJjFpz0I/L7FR82uPMjVTUft10A
WG4TB1HS7u4Yu1DyhSwIltdJlsBTF95uaMRMFPJcsl/2Rjtc1cpLQbP3qn2LrZqDxIyuQFPf+aBQ
9IWJxrEMLPx8kFy2uLrCOzQFX03kp6QD/c8xbFenFsKUfudTlgRlyGYItT2y0tkZrhONuVzraAPU
Ka0vorTgl3kKboKWH1kpAimP3T/4Rrm+wFk4KFcHNYwRsBDFa7wcfZ08F8GKOj1HqyMrlDjyHICl
lZIfOSoFy3oTYt8GiqRBhrDNCn9CPBHtCMNT8z7hxGYEjm66tdL3pED4ppNotFAZrAdoEB+gG4dD
iKkNLQXSuYu0J9EEUJYCD8fbkwTugOaC02ECQjhJnXcmLHqvi8WQZL8NKybHDiIXtHDaAgdIscBi
NfCU7wO3+Xv7+EpeycxDmqQFneUKyTYKQ8t1OtxuurTQP7p5v50YxmTEJQP1bJcrS/t34Hg0Ykf5
j0PD1MPk9RoQU+ZTOMpXy2RYEoeLMIgLPIo/R8GXA77YW1uOyYghZdMzy5QhN1hGIyd2zFY0xqik
iJ5uCfQWroh4WU7e+pVjZkcjHCsVJgXHtsDXNVwV9jrhZj1L0PAEYSn7rzZYfWSIn3vBLkXTTMQB
YCGtfbDATa1IxyhOrETRZnnpEN5Az7kbB3dxLPsw62WydrsaGYpyZi7Wa5BjG5h3PR3sn7fv+wDl
3aZag5gL6zD3pK9Wo95NVp2rli3IBVRkYdd9SuwTMG64Q5hZwXVbiRenoMp6NsRMwRiAAXVD59UE
jmpkD+YCDU5t1UaVHVSvKwgHOUY6WzMAc/mixcq2d77xSxdAwx33VW3nng0586aSBfCNoDHlA4pe
UJrEmaJxKEeeGDAFVsMFq86vdDyuOdQmum4hyuki9KcynQen6vuKy6wJzw3fKUXf4NrW34Hz+B2u
/wG4yyAyMLKLcdQ7cr9u9YWXfe5nCNPj0U8vW9YTARlMKgFOJqSq1bJuizP9Vqh3E3qPRt1/+9d7
33CmbKxYtqdqK3I55RWIy3WtjKRsZG03MxqN7kFoztwcuRSirmHx14dwsLueQneYjxrzrkgdS4uq
SrxgpXc1r+YI8Bxfaricv7cwFMGxt2IDzD9Zx1nQBiyW4DovpmQaO1svJQ1qye0AxZvrnrujV9ZT
RUhdvgYRmpHCLsf1Gl866iTebvBPV3fXrDBX6Zt+81n/wSTOTvdlwzBMwXX/WpBTEATk1BiaOm5F
I1y+8WG7vnB1s3uL0O91jyURMCj623AGwC4+eYaalFt5PXsODEp8CXcfwUwbKUpMJSyaXcXAi1wU
Zu08wVbwD1gwJGN/Yaj3yLTxg5UINzd/zHfl5SrHLQ4FLE7LjiVzDo4xg/+zNMk/lZZp2dzpe1y9
wQ2rMFiLuGjxVH+8FzCj+7nkQFzpAwQ5siCUUuuHwfdhr99aprrXegp5tVKDlC1cmhVANDx5GYSZ
EtbjR6Yrg5uXsKg7+v6/b4qj/LMwxe5l4pYHnNvSFDu2Cm/nD3vtEzlZfXQBn8L4nF7Ilcyrh+Q5
o6ZP2mE8C6Szzcm4z0p+EhPR5km7TXejvFkR/RZ+Q+oBmlVRnmSdPyKcBBV1xuY7Eela5ZT5hXlj
vWlOfG0wu3skHcEMRYIBBfmqzgc7eqoRk7J+s4O1rbnD8+kMKe4BlDwfiNJQj1HFM84W4Aw9IHh7
M5OhRfGfcqcLNhuK7rjXQbv8pf2yP4n8TT7pSKM9dYHrbyHcS1ibF7IUnaO2oQbUkF6Ga68jix+h
IOq66LyKKogfEeP66K4ey1qfcAreTh3q+uOpW5+cT91D4QGp1Jqq6UzQSAC1RwuVmIBzmLy7Iujy
bQkNXYAfdHc7sek5k55CekUF8Qk3oE1XYoG74Gdd4H4kEFgib7Qb4Q5mer6QZw2WMw3YOVSsROCu
R1bxR6TC6qFFFxbb2xIKwUYpMSGsLqu1G/hwQa3mkQ+6PhF7WbBMtxPcfgwfjpkjCM2dwDFQmnGt
X8tADOXUzJbpJT2tu78h1u/xzJsG5Eh1HYAQjzkUwpu2AsoLjgoWNBngUcj2nr1O2G+mfpRFNu8D
2EDUk+Pa02chiYfCyAdgffndAmzN45JHGBysNyS2wdS3bmSmr/Wxtf2ZTtOqyl8ayndzgTtWH3s+
rm2/MB07ItQx5zxYj3Gum62eEQWPvCxSGpDlR5QX4ZowiA/ce2H5F52Ks+fl1nlylsIzG7IFlTeL
h66L3TWXI+ucZsYBFWPQ3rUv4C/74C6oQ+yy0enn0Wl08dqIJqTfq+TfLvIXy5wS9rtuIP1B9hHD
CR0REaQVh6i13fAKKz5KANH1Ai15AsP/7iQjq6UyZTPn8l/6iAkcFbHCNFteXkxCUvXEqbgNh0PV
DzPX4V+4d1VfhXWOU9oQNZN03s/wuM56OQJmsIMAblXhmKLLButmDkv9SrXU9tHVHRBJdxCHx5YC
PmiMOc3zsKY7Y9FmRf+HulSK42CGvm31N8lMQvm972nce+mdaGntg56xhAxz+H5NTfYrKmeqfNrw
cgr/fdSajJrVGrZGLJD+NiI7y0Y5NlE9BxAkOdqQ0TlbXtzF7byNc4CoArurwQP44siwv8UKm8Xt
xcVvUf74CMgw2izDVprOyp2Y5zvFgA/fZVupxpL5fkG2Sl/n1LZf+OSHrtABcvwGk6GwVdXdacZx
a9ztcwVNk3Pq+10gmK4LFe4EmRRQGLrsGPIRLUkVB9n+p0tEU/+NK5d+UDkEMsPiIR9ZJ7CdWC3J
dx7x9GHiLHEdvBZwyaegvGB44L1q5BCf46E5PJaB5jgPqmAYfEqRfrYPyN5HUG9xRLoJWGDpm48a
gAq+bBJy5z5XQKZPslAKhd3YGRpk10PhsMvksiILUrBRTVHk62otiNQCyq4+ZM0jTpc5Tcqj1qtm
IIixHhgQDiG+/jVjArkvymwqXaHwusyN6B8F7+D00RT/uekXpgS3aA7/v77xUTbfdnRUtTq+zgDI
pL4yK30npBq7OSvbBFODryIiAYNlFm5X09CCno8yYxe1Ku9T8OLeWNId9VY1BZIztnkDcJQjB6LN
Kz3NhMs6DvLcBq3YqDV7EHcnTH7uHZ4f3b0wWpy7CYog79d4kAklAw6QtBRxLnjzqg0xUniLsTqF
j7x9s6XShBmi2jkjWtPF1saEOaKMLiPNDaVboePjNfOseIKxO+rrwW+M4jQ9WzeELzz4tu2sGhSw
X0m3cTEdk7AUrEajzC6FHv5pcBkwsNA9F+dr97Pg9y2PNH/Gu6ss9wdqtDPHsU2OwaZ++nuUfaFP
x7V3aBQVtUAq3cqkQGCSy/K3xUoJxLSR5u+JDf8y8kU94tUa2VlKKhnNqSd/dImbB0iITzpcSAi/
AvodeYNtMZfgYj8Tyf+ZU2wMgFh4SsTyVWDLY3+kFT2xUJBk81a5d1KZgWcbn0TnplnWTPTMaKYF
bp1ImY9J+m+deUtV+iiiGdyIj5X3kEjpWI01HLRaa++zZqvCpoespfjym7PUkOmbazemYDdARNSF
yZ9QECBlS0H3Q2kZeDPj4orr1lf8YRFD+rGyIPyvbjkqFV3dbGd0oOGFXG3ZqVkpITTyk2/OmPnc
i6xsat0XZuzLelTfb0/7ep8PsybEEdSRwzpZobateS9MZRCEqE2l7JfzJpYOaIeTbHO98RjFRK/5
hxYFihVCOb4cRnOqKNl2kJfo2J4z8OTLXwOIiFeYX7h0E8lBzL/uLv+dOIS1VRcDKFRXh8JJgz5T
YOop33MvnDCfmupsjHzDhTemVrGhVu20NyftdBcJz1qozjnRBvjAf7pLXdc+SrVT0b5njvsMlm2w
qBf/kRigYnYEyvlKv4S92rOMsMP2HmceEhZp6JW/rXibsb/v0Ynjsico/VjE1tIlIRt6d0o+0quB
6IFcpbsO5HclEfb6PjBMUlRbyQrUZx387BY0ON+7HbuVsPptQGicsGYHirChxC8YoQveguzYcTBe
VIeG/iy/gO8E5ML3wRhhpQbaWExzW5eLmA3uoOYoDfYbrAMHgl44MuMEvYeboMCVH1hfIcBZA3oa
PJUV+ulEzOcti6FY+zNqiZB18k1fJmyCaZ5Lk7Lj3wqCBCSbirY2fqLSU2KAZJUhsbgdPA5ryvLK
Oske8n6mKLrdchPzpmXW3TWNbu1R9+IrcbLtfjfP4rY3n11aXR6cwyEnbIBAn6vH5I7lPose6O5r
jDDEDmmmMbiVOsA9pE5Mqgw/6SGNKdvu6HI4hhwwjssXvUIlJ2ad+PXBqfnaEfJ7iZurD5Nbn+fx
w5pe9jowHIhppoY6MPECbzK7eTY1qRFB0qlAhr0EZs9gbbRSH49KjOmJ7v+3MaSFWcEtl4bcGI4R
+fAZNRaceHokXNfvPjafuzRXwfMk7NMDmodzu8VssOxKPAb0NaGy1Uozp4rSHDcr1MxcMT7U85A0
8XJRVtRa4PI2NevfmNa2jPiA6l47/t34oQP9GR5P9NhaRR9QkzjZ+RAM3lcXFYR7+mvVcVX6mjGp
RWvadW5Yjk0qaWg3g44z5ImKBMNM+JLyMkFodbVUR53+ZRA/KX1Gtar3opeI3UOs/L8BL3lvSeaz
qqf1WWlhl8bDiOCDZMNn2Sh82wu0NPCMJljD3XfSiyk+vPTcDEvNn+81TuIi0/wj4NiHbixDuJYC
3t9FxqVvZzpyEVFc4KwwwjFJRh4CDehJxGxKHb5GlSQN5FDYUIA58rMkeJHlsVUUBAcJXgMBqYge
KRhMaFX6ezlEquAKyo+l/gYe09vul/CyhRuxirKgbnTKh5xApvyNr8nUz3+pxgm2ymsrkjwBe1kp
Gp4pmtvVB0dbFTSKAVQA/6Uzk8J14HcitV+FEsil5RhOiruCLgWUtLEL3oGfEMTGPNPmZtTAuL1R
lCNSmBH6K5bWQyGKDwSTMspVcCw3Wp5Mt0Zhfs7XKDw2MJ3I3OJkbYPmIXyb+HLC9OUlzPyvd0lK
JOj2XGrUpTJRxK37pmrntXVuhiGU5pVIw2AbKZQOtNodIJRhcE2TFg620HObBu41p1Nh/w/W0I0j
y13ubleXbjjgllurgUZ/XYBs9dxh1FW4BEczdGJn6Yid4aY7YwXL55kIymItM4i1R54t3v8ctoYw
58N5aiESo1PDC/KsiZq2PMuPnAVUxASwWKly/GkKpNf1FCA8zEJeTDQaoD50P3UfkHxCaCEnjOeo
LoMzfZ7vS29SMjJtOAgqhmnll9HLkaYSZ7KpKfFEbYomHPgZ7WpNrJiVdbTOaBPrhc4uYJLMjlPs
mw82Dll9/W474FEPj4tqSp0nK5D/lNAcyp9uumbQZKkHYFPUXd1NDN888cw75R1HPCAaxUljv4L0
nMZUWWF2ni97alddsyK7J0BiseuV8D3QD7kCG96LHzHOzlW5ByVw5dceaJQ+FDUgcO2zzXwrQTOj
VjMJ3o9DzhGeO6ieEZnMp/Ut6Pat5819p9lnpUGJCcgu7W73JVhJ+wvkQ0EP8c3Nh7ppqKOf8pOQ
Lq1oaD3w/XDyKzuhbHG+nEeC3SbjhT0KQMBYVxESajIwF9YqtZAYcRSUkDxnfwUa21zVvVn/sZit
GpUli0zl289w9j9nzGIFlqCU6TYDpjpGf49MrRdc9ZVmmByyu5vd1Mab9UO3YFcPR3BznhtoAwYA
+CI2XVHjCb4aMhdQJv2GHpQiE2A7mcYywaNyqPohpXjVp1WfC7nUdhALS9/PRBfLn2XdpQ8seLK1
BACzB82W3FEpp9kHXBr7LO0fnJlTzJE8EdA0YhJv/H3wQjLp1YzZPU/xD725sbhq/czo8x2S73Kb
+35Js2wYYHmGGEuE8LQBPWTHr2Uz288STP++7JtSORkYAPyiMK0xhghM1rL72VkA6N3lA82LxQDv
rf3BUxLsQ2/uEzmcpYRDyi+ZpiSzo0UaMmTtek5hVxa5nTOASXK9FwJG0Gu8IAo8BoJ7HFptnK1T
eSXhzZiKhGsMzFLozXI6kGPBugJUaIP2aBYBqNu1h8SbEllkGHWv5AOXhFT54pL1iJLFHtQBZeVn
fMlPutN7Ig6Z5Z2563Luvgg0SU9q79tDZRnHhv80fABPpRKSv2CiYyDrbzmTG4ZTOpXdQpJS/DsS
JSG1xDIVJgMe+k02GCVpZEd2a6ctqGFqkmtd9kqIaKajCmc/9SIFkTqpl7TaDjif8YZa0vS0yzpB
t3u93mzyuIhhiCje/RwyZNNaPcp3xCeIjx9Db6SDGaFIcaocSKsEBS4x7n//f4JkNX1ZqhApsZW4
hecqlU1SDyT6KpkrZJEK6MJrFwwk5kAQzTQyl067vZias76ozAqxwA+TI+u09ATwJBUzPVysBPjh
tJ3+KF4kRUJMO81X3M3uwDgBl6oaNSKrbkq/+irfDnrEoD6uC5QArs45xB+cbILxpYRpMwInzjZF
8Ysj1qgLhY8obc8+9voA44k1nNHETgdLry1xE3BzJ2E/VJdZHDbjCik9NOgMm6qzHoAnHn+c2DPD
RgSHF+tlikXUCF8tc0aA24hDOje5qaIsLgNtnawh5DvLJN+knIfPSTJ4GiXBh6jWas+sD0Yw4GXF
gr39psHybPbflcENCIn5LOMc73QLWHmjmFdK6Sl1lmHbSBpUhDiqaj51DZDxdH4zOGEIp2wyVQZq
w39ID+PJRDviTMeoaykPH9RNW3hQfYR/Hj/HZ6vnJWdXF70fCMSwdZSYYekZjA8XtgoGqz37q4hJ
QDYuZbOy1PZLy/z6jQ5M5fyjNzMgu6rJOYULykYxxaK9R1XOOfpKmrFqcStLQ/jZXwFIL2lWjq2J
trbg6YISuwq5ZpGzs1ENT5TruA4MpApedblTQdWwiWEkCr9mMpnBl9MczvAxszsZGJJA8FyWnhSM
e85NwO5qVBDY7H5C9WAdNBhVgbGNinJEeXkddu/kkpInNPjqDePrlOeeSTtCz7iuybmQEoWg+fSs
lvQ7I59sM8EhIdbzPY06kgJPwIpN9WUw2ux5jFf3pFmeGJUnUw+35/eoLNRpD4BxsPuSMT/mn//z
Gg+ne1aFhvPAgyAhWoRVPBjNcrwZ7Aiu6gcfsLlz0mzfvt9nSc4bJYSX07TeSLpKG7/lO1FiAsD3
mtwqVQV629kSP7r5eqyC088pkw/9fIzD3zpTiVZ/34ASGIfIiPEv82M3O/tR6bqMaSJv3xS0Ue9p
VdC5Xw4+jBE+vjjpiHE76Ob/SZYI1cTT8S6UoqGvIyrpX8sNU/hHSn1lCzFpHJUbN+01hMd7rXU7
EmlpnoahjMz3gxCkbur2gSQgIAdBgdEBM0tV44M58tz8mhQJkvTk9QoA0LNazcRluvAOTJUXDyMR
l7wB0YAahWIL2QQFvKx02uKpa7fNSRQzw2OPI3AVxBufODI6rPyDLt6VkwDhcKG1elkZo26VGb4Z
HBjhDxeAWiTY1ugoiQl1VGXMx6AgIRqLVC4IUL3gZ3NhMu5+bosVv8etVbcnm06Y/f4dd3wkUqmC
uaDtsVMX7eK0FocFkRRKIBzhzrUqnGgyM4WK30jfDIVGP0Ti/EpHN6prZOWt7QBL0iMArpc60qJz
5AvxnfTQm9MFc7jW+xr4XXfMIdfeqKIz+7p5nW+ZjfxS7/trtqHYErC9xIF0mtt58BlxmTtrAneV
CSM5uxPZFEOY+iumY9enpQWfPMkwZlcgijHjw+ySEfS7FRH9AvL63dLe97fDnbHNhH3mn1LO9Nhi
hHavmZ1NIVTOTdNuavRb+85MvppKR0RD14yEdnvYl6+iT/jvowD2gX0cZWVZd7hIcbEAx1b1Ktc0
Rf/tXMK6/IZxB6k6hMjTaa78qiCWP1+jf2YwLFSt+k/Vv0IvnGpsZBU12VSz8EJbzkm5hzVh4v5E
m9MGaFQbDCAbkCF9G1GRdkgpYOizyouQyZPVP6nEKrNdiZ7O/Zng4H33rQU8NYtdyDgG3fXdI3Q0
aq7cYwJ3LvKQ3zeeZ+WE32i/XbuoOTCg7mjF3sbk6M5WdWbhsKLdc3zcNvyyvnd0w+z17VnccX/T
cC/lBZOFMIqO8Eq4lM5oN7BakOixDbDXJ0m3dZnnDcn07Ys2juss97u1lGTndmQD5Z352h2+nfBy
arQhdSZ+AHHaw5VZNnhknr55h5IbqPgA1txZJuuekfnv6WoLpkj9RYOYHS2qYh4DkO86RfbJw7cC
5IzleZwkGaOfj83Ks+qMGtUDK3ecMO/di10u7OC0Ktz6plco07Ny6zf7hUJPdh551DzpAJgi5Ox7
kgJurAK2UaBfVThbmqaKQ+FRqFd+3QpJ6/NLYeEtAKaZooqJ4fmdQdTxTe1oCWT+W+fQpE/foXqj
j+tvr0jiKVA/frh8ueMWrth3VS4WWrsPzIm7FljRXxEFFkLlm/I8bnc6i2XvzLvytS7na9+gZnDs
LlliTAIfPZlSQxJFGrMyd5U/aS4gsoxODg8s31Rf+QeMWBfPRgexiMfMhIJPgCzgrU5ApDmm3lr6
kyReeP5uIeIv4UU0P2OSJsnUB+c/9g+/rX9O5tGLKUOgf97QT7SaoXjzo8CGVvudrTDqTlWcv7Wv
EdQ87pAmdKkMF5Ab71PDKex7t2wMvO0sXM/xrKuNoOLemU+ueS+wAdv45kZgkiNvdW5FDO9+gnMU
ZAoUiMz5qF1DxMfCeU+RFAmJ3TmcgYVMqohDlSSIcr9+f+lGKjklW1zZUr3bv+94ulXafog3n4dW
J49kGFWgbMv5sU3461YRLRXZlpcAbhiOuVwk3BNh5Obef33Bw0iU59koh/4wHyRXGVsWm4gS9e+L
R02+untV1BPebCeNNPXFf352lZbutoOHj9DSOnzLjXa+cDOegr5dAOhR/VZzh+CHXunfEXKZaw2L
T5YxfzaQfIGGKZ5/sjeZj4hPJb9P3CkcbNsCQgu/hcdgFIQenUqpaMYDW8732s3qpXVnDnfv8jFF
X30fW5CeYKqJtcvmdWUF1xm7ZyvVUTI5jauUP4TQIdjWOxNHEEHT8N+Xd3d6o8eJRUXv1ZrKN8/t
hMikzHeNIWlpwCEj2+r4FHUQ/3e2h8HpqC0HZXjCikzmr1aDPxXNe6uMM03ku5MSTSCuvvmUM+eS
TPblRZABDBh6PcS2fbX8oOjE+xt6u4n1GxZqGXN5tSYKpFb90K0HEFqzG20ENSIORMGamCKbFOgV
noNXsAaFfaGMemKEXVI8qh5emxv3Pr3d6NLz0v7FcVNJtGSA3K/dyqDii1O7J6AF6JFddBl5jON1
oxHxel9Kq1CejsUZQgDs8CwL23bGdMqESH0DFc0/6RPCKjx4wScbYfiC20I32mfaGcYnXzcN0QWZ
tnoeI4kX7vkhZr2v3WEFfceCuRTlMKid3s+g7rMSgFjmWKWRi7KKVA/Qf12DkkqmpI7Ll8oMK2F0
HkmD0cHWEjs+KejFEcXaj2gCrQWVJqqVjPMpsxn/tIEKxurI4EZes598gfBElTXDlS7Oz7wr3h+1
5hq+Tqjwu+7V2CHaOfa7Vy5xDaUiA4MB2zxgjxfRXbmZqRK7WW5VGdrzc4Cm3//5EHyWKsQHKuzq
mIhjDg+5MOwCCKnV9UiMlta5CXzqcmo4jyVhz0lUoe8s09cd4HG672IiduJqKhojPhLCBc4uIKdf
/1RYQiVfuiUMiiDUTcdHT66hZPftJgrK0EtFatennOBKw+vZQL66N259x9HN7FBT0nhNVnh8pb4c
3OU3j/+3YrqGRA+vp9Y6C3XmoUvqfq2V38jPN77uuTYEzO4Ce19x8NYEnIgDUF4mv2fczP5q1gqC
khaRaWxaSfCf4r90c17BoIPZNhLDxVPs/5Yon0p6BiF0p1MpNnkRoV6fhvvDadLVimdMuRkHGPd/
VU7B02MCwgdSipu1UuGpSv/uKzRG3Mdfy4jf+Mdkh3zdFMTto+wed/Zrgl/ng+F3ZL85IKI9azfn
kEjrSPx4R+zZM/zZVG6jZY5NpKZe0XUFiIFipk34NCmnBaOV7BiOGskQdAbDUPx4T1jYjVebfhQh
M4Fo5NHB5cbKPyKXAPLhERCXIYtOMRA08i6oyI9b2S9IY6RevSuU3IOOl9wa7Kd9bQwtvZMzFTVb
KqF6LCdmboV7lOT3sQoMi4DuM6evaEgItVJDafKa7WWXyRBaxK2HvdDKnqEV/R3y6LrUXioMfH5k
hgENwalFMz896+uf0Qvg5eFGMrSrgJNDe/N2cfKfa3bIpm+3pOh7v8fEdvC4IIGQJ40pYB6HrdKS
BL9T8hVeBX7a+i9ICFz/3q6wDeJMWqKAT3spvLTPx5fwU9tBFEE67V+z7pdoPxHBo8BrzzmF2Z0S
UGwqJw7NKwm0kn01C6jZ0nG2nbSTdQKYt6OUFmQh5yabFikbbmDbgN2+0gjhOm1mZzok2naEuWgN
kab0grhDVYy2McLqm50eRAL8o+azNGWxPMuvuthS6eiDLZB/3GBKeqlBddUpSW4oMUd7Ntz8evGS
y9NlP4btnF2XZ2YGntf1HrJ6lQJJNO/UNYC+KBzrhHEIFmHlJWRh5u2BJPRxl+XslWJshndKfVOa
nYYGHlha3DPyxI4EFOxFxH468QRcDHdRNcnvCLUDHOwN/tuBOsctV0oOfUJ0K5lbEKph7Z5vfZKc
eMuaPMKxnujTEHR/F2DJeR9gdAq+KGYpx3jLJbFZc5k9VKrfdEVmgQPZ2OdoZmN4sqTkEQRp2hsV
i7XglOdRkM/fJ4U8Vjl/GkrbGIND3RjK9o73YYneL5XCEBW6TQkDWtUStKR9GOmQLo4DWkiEOF5u
IXv3j5bEOETHCjoNHMmeR5NKTsqLdPSYI8mSCdTMy+c6EfenJmTYcJLrhYLK2qOOIM+NQefCMsFY
v4fOtq0310oxN05C4uiPJZsZBkHdlIeMen8zaUIKOpM4QX+jofSmC7RtOYkZIt3KvmJ5qYPcLvim
1/sWI7HVanoanwg0Y80ZHYriEWSCV7uVQvHO3wdEz3GuLPB0XZWTsUiTWxYyZNKW8pchEQlNrtwZ
iBHWryr4FUOU46q+1Ud4xIELT0vAN1+grxfCSPZSyhnHpMfWRcTGSwW5f7/9YI450JiLEFZyp+Vt
wHSUYjK4cClrbrngMFz3AiXI5FfNXb3SdNmnTYt8WRLopngHC3piEzk8wiWcMmirkMerlZBHcGod
2IE8YWKyR//hUXHY9gD9n6rmShs1KVFVwhz/zpE3lNVX1vOqIuZfqkux77u/u+ZwPkLS+8uFllyh
S0kaUUI9GAdy02UW/clrokJmR4RcZLD/etjpA6TjkCpCy0OSFJ0GDsnPsuP3jbnb+q6zUpWw9PYx
MMdNfN74Hcpapk+8/x280XjonLVLIccMVW+SRmPgW0zEEoOaobL7h8AmdTLXHxBgU/tITbB/dwmc
oQUeEWkNMThEvPTymOTB2BqUhh3xpZeoscAmhgIa8orEAVunPEJGqStJszMxa753JwatC2U5OAvc
E4O2QpVkfZ2Z85B3apXEOAUOUhhv5wM4vZxGe9rqihpUauxn7jN4eBtm6t743SLn+XRFxSv7jWH+
Xd/Sj2o4P9anzKbJf6p5Nubpm4DNC3wO3vIjVAgVIPfWzxv044xeG0idsQnNQ23jeyaS90E35zcs
vnPfZHE3IqHdXDdLYGf9/XOJxB3VXQ/fBOvUoSEx1SUn1YQjLN7Z22HdD7QqT+E2nsZcgvG1zkOR
kbgfyS/sJrapeKOkZEe+OS+k9JtBy95BEmdpm8b/hSGW/zATFCQjpSKikDeXGAcZ951Pzfo0CSAd
QmwkTxkRoieYdOHEzTgMbpNwM0BYxoa0z2fKUvfVJrUk7MeRLnl3CaXyK011th4Rpv+LxJVm70Ty
sea4E6OePbF2ZYRdb8sVb9JahH2CkpFXm9AeeZW26NfmOuYxzJZkn4ZbTFlWPsOTWFyh1+8kZOtQ
SX5qCLGHxDPWajMIcE87pb1dMAHbOOXesKXm6iekGh4GnKx49ij4KXjyCz2SzGRX2s1kA3VglAZv
0vNedf5XVm7UAIOsxpqFU1ZtH0zX3W8Cj9zzyhIfdaeojmCIjMuaNx5xaHfNVXYsv12XHvLWpavQ
n3sP226m+Mfilzsnd9yZ2xQ3/S9Efjy7P+ZxVv7/Dq1/t+kAFpzcBsKFQmT9KTmQ23lvVnN+BKek
ivZ4R8n5DRbrkj1PliLV6pO/qFNXz/u+1SyDZcQJpvlm+xJy8DlhhFKgBUPMIShduvTZE7OedlY8
vwdastmebhGSUGAKsVdCJieBO1c2T1ySVInymFzLcj9jAGmMFjeiUb724DhGRdjKlK5XJfrSnEZB
1mOMwAgsDDvzXT5uCt6Gh7XrLJQTzl2TXytLvbdN/mKq4o7sj2Gxmdv6oVPvuEFPs3xx89FBqkTP
tGQabqpBOOpLPQNZui1mL/1jxRaWD2iU1oT5DJfFHVGoo7rclmYv32cVXqE9xN90XYSvFzmqe9q5
FYADwepxxItstEvFZQBE5JuD2nRxKpGG2At945p+l2m6w+wO3pfEwg6BRTEuawviWG8qdhQFqTmq
5F+JlHBKFZNdU8l5yx0evtMtr8Oge7Xu4vSW+FeSAu6ggU/8uJlo4TRj2PkBqNcvVpSifjLWwkaW
AoR3jQWjdNy80eZlFHx7hCpn6zxutr9Fxt3oeskgKmiZDmq0mP3wwPxPbZ5/kFCHOFukoMwF3o3d
fMRvB/OSgMw6oLpHZ19lWcvh6NHlLzgCx7kwnSjsW853dLIh0nrqacH5RKfLN3xE0r9pYpfL7+F9
ChQBM51aJoW2Dn886hWuCRIMXXZ1sMHuMBLnwc7maF76P/C/lTJg5DtH7u5RFGcuC6drFLG2WTVo
v4+NZaSTAcGZYmqjfzZP9Xt6OrtwsINFyInKw4bXsiOYGJxCo5n1KKNP5VKsjMamGazDLjFd9Ill
CXS3kuEinUMoKMfflmuvwMYvq/We3reqVtfn9kdTIgsygO64Dcb9JtKDVUT8IKJlWtzRQ2FZQwmN
PmSvs0v1aoLkDKxfCWjTa774CByRpGx4VkiiS34ubr94MlQfUOfBJYKhwxfGuWCvnY6sIfRjSxoo
BCQBS56wUeVIfpzS169mVMRdacuFb7dcZPnHcE0qb2lGegB31BU80Zep5iIkcg2gd6TfIWjbpVhZ
RKFz/1UFg+p6Xh8x8x4jpzWG1PM3R+7UblBHspkG8K8NOwkMr8kQgfmwHKU6oxD913o54wj020ko
Jr0GaFn42yWxqzq71rSLEZC/CcKFWg7mGF5gsC8uF/RMcs/fpML+g++J0OCMz3xklk1tGKkv1vQ3
kE74sw+VnRo1PxYgZJfuvUQ7KBa33RrZU+b0sx2GkxrC11uYVcW++XY1lhY/ll7UniVVFdy7F8PP
uwcxUjqgAKGbiHnwDVp9jq/SxZjdLLmOBPKE5h8EkBesrBmOXqjyoJwTBDiJz0yCbVf2FDzsxQS1
Xm/CeAjDEoC+quBoN8CGVokZs3BE9q8AViIgn7FyiVk43GnqKwUan6Be2zSTPySxdBPJK7DUkyTo
owiA/6Ow1fQIQV/NLv3Bx95CtQyCaXNgtsm4+uWGoDZo4vRssPT1l1SecMy4ZYyqxdqjYnOtI/Vx
JD15MF7ro+Z40Y4OnmxV+mvM3dBu/h73hDQ/cFtw4DqyMJV0btlbfw3Zllzki5sAg6iUF4RfFSZI
pBWUJ2ku+UBR2UolvO/q5T+Ydm52ok2PuxNk4ekG4YGKQxRtKgn+XtyvuyxusiLLO8IPAiEF21ZY
+r+aAEb1EKkAYJtrJEESuLSV635I6lcTvFFfkyFAWZ5bbgpe1ZB8lpOlqIjAuyLt+nlpA2nuejk8
5nCyn+gAaOaV1FKWqTvrkvvhsd1yRmPYf5SlPgPov26eNrSv1JJa8oqwOK5iyoAXsLowUCUPXgfE
kDvU4aKVA5lSmadC/GuGBp4bfehL0JYGeqEZezft76H7oMlN6GRJqoiGVPa4msQ9GGnlzOjre723
Vr/lN4SpD5znuentsQmYXtFvX4I2PNzOCMxUQGIVRyGQyttQCt440q19F8VUs4Ohxm+n49ObjCAj
1PN8xm/yspY2IW4gDjFuJfJJckYiok8IcTU5eXXImscxoJ2mslvN65iWnkVneaVV250b7QBfTh0X
BRDl9J2GS83PtIrH2L58U+kd9FDfBpEWXaCZSUBu0GbVflLJ3/lff55Sw/zyz3jDQdN7rbZOzNTp
4k65W9bm1arWTKDcnvSlYcahqFiAFsgSA2kv/8RmPai9Ad2PfsjbiPjvMYLwZAzyumycQgKgX/Xk
Aw0v8/Mr4mrE8Qs+XDH1V6M8BZxAjGQvTNUKr3gzv7iVRE86U3ttUfTgzTv0g6r8RkS+fC3LPSD3
u+Y8zN8O5QhD8YKGp5wf0r6NEvWxr0+FIlPh16VgEkcfDN1tbnauiGq8BFTdzTJybp/usUpVvMYH
LmxQzf5EQLIWgPqhulUsILk3knCqQAwOPzEOdLyDdVQBf60i3z0LKhtRI34FiaW4Nsmo4DNwwC4/
dqzdUh88zJd4AI3DQPh6gN2OhwcNzMLY+AZ/+RMDx6H592vf8WpDefA5AUATDLiM7/JAg0XR5Rkh
pbQyeDAwUxSx7so/RFB9B3kwVCC/zHTUFrjldtgwsghcjn1kWtoBBkZ8rB4GY+KunewPijWXcH1v
/DL9wBYdoBMjsOPFkb+GeTsu6uVJwlrK3H1Sg1Wyz3GJmc5y+gOoA3krlicHjrLUA1VYTGXoG1IK
a/v4iGISewzE1AujV91YdSIbMGd+Dh5KG6FL0Ek7rei0FjM2g94UxrlUkn4s63BM8yFYY/viB0Ct
KrTZgmVmp1yKsAGJmSwBkPLR5qOBVIigCSPtBsbA+nKvlhtxjUeGrUo7x7qV7BFWDkvJ3XhUE07W
kjHdeHgDqDuZpvwh/JhGydzH1yZZNoZoFV2qIAoQWz7BaFkLXVXta6U9nmrK3S+82QrXBsrfMYwM
i12rDvsZOcyIbj31EEvxdWTHhFAeSJvTxeXJaKfepr0xZFJqaEU2B5/6JBMcOPWld0c0tv1rJaE9
LrRcWP0Y6CUKrWgUwb+J4gSQi1RSo53Le6PLSZAwHZkEfl4Vy5UIPi5f+FUkv+9E82t3clNLbhJm
tQAjaEYguq07BngqBKy2aZExxIb9p8cw5aAdFruwBplKscgmo/AgLUGWYUeEQo5yqkernc2ayxws
1fFWJ/hCHqaREDfr6MWEcMUcn4XFbvSFHwOsf8oDOvACAPXAGtFFE6rrVShSSx+Ovoe9RBGGVkvn
bYxCn9HyZcPU8rs4lU1KPyXQEBOSKCcP2ONm0xouvBkac2cJdvaTXNqCOZZQuM1jnD9eD2q9aZTh
yxbgVaBCxxcWsBm1M9qBM5ymCgpx2DDpDctrHjdibvF7FGQnbvep1C8r5eycqAR9BeND0Fs01oDG
PAxHCpyMx4uE4GbwNsxe1G2NWWVgaxfTLp7dDSGJKPDA+fytlkI662JIxtazpjKgCIuIhnwRBXK0
CydHMTDSdJHcmj4BgjSlV/Sk2WSI4Vpj8jso5Qkqgd3tYFvs43yQ4vJjQ+j5BU5+4nJpekw1G4IT
/qmqltMXmjTrhK8cX57HX61NJv6wJVnAmlfpI2LZ3EJ3dwidkDgKWxFpgLblD0rdct8Wa+Q2ZFy9
gHugy55zdpawqRUOFBZamw1Dn9SXG0O47N5Z5YZ6fCEuihcftA3VLhGe1amKvAA7+A9ZrPS7G4dG
w6Cwrl77F4isHBfV711EXOMBLyu4AlM0HJOmTK7y/W65RzxH0LotrvZXG9uAXXGi8/IFtf5xktKA
IIt7Fd3ulYrYVoE1n4ZD+3sW28pN9rGgWRhwOpjPDCZ76dLzh6XOumFxHhkKlgLGMr3OBToPgzlm
GHmXODVHr1LnpJOS8GD21trzUrhiVExuH31Fu9gWHMLmYD9qgw8aAhxf1E5MZ7WlLZq+FkDW/lXI
9jm8qOVx84G50cUjBG8il4fqiJWB2xQKi00w27dRulVin7nrVJv2LnVAIzXNU8PpQR9FgAAjhhEI
WJD+igWJKZ6Y9fxa0L6QNuGEDMxsC3ZLk4ukL0d9w/FRpYXiwMkhvUifFeSTM0Me8PXBUEPMoFgS
Yz7+C4rQDRQ6WV3kzx3qfI8+uoUf+4Qys8/C3QrkF8/exuvZdyrri1s1MNjWXyeTgIoLLSiyLwu5
QpJsi3rprV+y3C74P1UULEGlfxxchVH8ZgoOwA33RRQscGFnUgORryQkZcjhNUlp8uLeZ7jNZgoZ
NdZsO0lhrNpAscCd9d0h7PMWlMwBVVOuFei10nMlv0vRHNgg7FhdiwnD4wDXJT/QiRvB+9hE9Z+W
b7cgDLA6+xJrgzvETeTr8aWC9W72k0Iz+jT5n30B0UMGfqLsZaWd/TJIR6Ado6bwkUTWDq1r854d
45twsRethlqzDh+N1Cth0137Bw5Hr3/nECX2CwwNJKELQDiftMgOo3ktkvGs30GjtRmqu97fOYOD
L2LEtIapKhPm+1P2n93HPzfeRT4AC1H166OUVxLDzBorz9OZoEX1fAzyj+RgSNZXye2d5pA528Dq
jU2gUKMy40pCTPxmTvuSgRMw4Qrla191SH9FN2jFzeFshymkPrVvoolP1fczh/9a406bpOldwl7P
42zM/aqovT0GLpkm+HefI65e0ixyZJ4m8U8HrhNoZS2EN1w+QUB5Wf/aRmSj/3L+WCa4srHNc0Ci
zKccKT4EbvTUBmXo0gNL4YS433Uo7G1bpflRru5uW2YGrNLU/QleG6O8gDydTgNUCwBnt5mW6KFV
gdQ7XGIMfAGervNWe7wjdhWt8VcBePsCF3M12heVsG8LJCyrvR2wVaBi7ZpJzKf/RK+5CHVo1FGI
Myo/df7q3klUaWtuJCR0q3fC1xQJZxr9bbaZNMt2xksmkLAF0tBqGB4eeA1s+N/PibuW/Tb7erdh
bhAewcCSBZpS2jRFirnatNUgkjIW0cms6FS/tRxMtnt2l0t8i6qbGx8AY+CliCHmt8upOoJB7ZL7
wQuFV3yYuXKWtS4C6PHa64siz9E7CJILurVCneDj3aFqdvsy23tNn/3civA5Jy6rkSqg5cYeY+Cd
exJt9kRCpKVCY5LSnNG6EC1H4QQclmBrJ0hWN2L0h+170+8dGS1GR9XgVD8UzOyCs4vciydZoI0A
XJzLJD3RIGj8EjqLB0OO2uLt0HOKufxBhvfbBUIR95vMqiq3FlSmcVSKfM77SIARq5yNYlUBVE5M
ZVA5A6/f8tqTFsMInPIsjIPQLpAeAYTGYZayH4+5M+FnOS4aClfnKuOA3IyCmFy6chTgMZ87LKpb
nqaZAxsJpvnxkC0Gv6T10o9zm9qZTPILxIraOphrCHHi0B08qPFGNK5ptM9NhSAAC9WQbvGsf5ZI
JK7w3Yk5mURvDHOKZxuO9u1MC1zpxXPBNFMMxKRRPWpauJl9pfV98S7a1xPb6Dw+Rxh+WCpaKVn7
5XLnKfMLXAGZHruYr003mblpJw1ludcSwqV5O8JtDvIkW3eqlTkbAwA1MRn0pGDhr/T/c0Rq2F8j
gKkDcIp1q2kfuvhtm7i9zK2PLAgIyOMksjd82hcreLy4cVbmcdZaSEJa4Z1yKOvE8YqE4R6fDd35
FKz3uSGATju5D9WzZcDazXKxJZzOmoa6SldWNP38LCkZ6i8h+K2C0YgtdxF4CP5k9Ux+dUDY7BX1
4e1WxWmGW3o8aZsuZwozOUoqAKy1yWNb9Z5FtT6AS4CUWHGwrGKHa+l6Qw/36ZayaMmCkT6VYvuL
PwElYoj3iUddhOil2TMLBf43Ti3UyQ1p36NLSwo6VoOrwBPV7wQBFh+vA5LfSBUnfkKJILKGxal1
dsZfWNHZcTw8Bn7HXwzeY5MSNwXU/9/Ybt6lmTDkznzfuAwhp50gVUXyGpds50A1xFTDTSvTcURH
zKuy3Rwy1mRFd3+RKhK98gGYDdIqy1mU4BJnYEV73QTG7gdANXP6BlMMqWLJLqL29Sy/N7UzW5A7
h2wQa2VfvQ5KOH+pGvzW8SOd5VFMaodCXE7dL38WnKY4VKTBoaXa8eY6mlfuzgodcGbjP2kj4wT/
iam+NEeeufKRbxeR3vPrfCv0aWjhsFEiGaF1E6IYvO3vc2IlvgH+b+5qs0uxX2afO4aMjdAgdJM1
n8a8tnFEYIDkO5xc2SM3VXiK1JM2SurTeI44z22WZG1FxqzsbhWK4Bd267AWGI3/GD6t/G0LEbV8
wzU/qNMSBBTN24eeThLkXecaHIYCGotb7EHHiOg5j/xnu1bT/oJ9BaSrhczbUQ3Xh6hDxC+ueOwb
gwmlkEpbeJULtXyGIoys9IEVLE9V0sIY1bak8ZfMM8F/RmDWng8sTZA88b8yEizrGCD8tSZhXQo9
3i1BQu/7k+DMQhwGiHU66O1sOHxY8jZZHEQ5WIH43UvstQOVKqDB9w2BRMxTyCkTrSaLSenfwWUN
sNduIJZIF7z1Xl1Gf5bY4rgt8WYwLw1MdqIrNSiY4aMI0kyWgtabyKe1NWE3dTazL+8QfYDb1vE/
+zRTGTKAPJtUCLMrZ+edFWsz+oC9MgXUTRmTjbWDzNeffQkjiWIDRemHsThjBwW+0uLZoRyH0d2f
w1YWXlrQ9Ckjr4nXRKYLFFK0aKoPxkfMGFcFj6m3pR8wynhWuv9Qk0WKJaGYp5VTiHnNwHQnXg+w
o6NKMYTjxjBmQccujy0Qr/gyvAh92uzfi8Oq4rSuhXlakZ0uf8o1/1wVUyT2TkqkA9gt27yLe64s
/R76fN/GT5VaFSuAoI99z6+txP1Rvdker5BGejnfxXY0zYtd/fs/FHtX068CKXd9CspcIggM6kRq
88hVEa/ojXrnU5Bg1Q+J05nqZSAxQA+XtaE4oSGJ43zq+v1k1CjyfVMAZKX+VymdvfuTYNejh5Ls
D9xqsjdhgr/FBitTDCwsUL7p0zxO3Xq5KXJfO6JqznxZJAcvLOF5VmR6dWQqMuKJ/3pHycj8cZZW
V+c6DHdZffYd1kznwigsJx2DDkVarRpJF2AFOW4DR+rfLnMlQH8ny81zZ9iEaS/d3mtv8a9LcdLS
3HZ6GOxvVvB3bAKQG9f4bWGZSRvzd8j4AxMzWW5lYt6i8HQYEE61St77u2ZUmDEMULSVzgPI6HJX
uezMTr9frqvSER4bKmygpQ03+yVE/nVjdU+pFEwkQPIS1KHPvg71SP3NASNs9WbWggnrLoePvEny
Sdm2To+3wihsRiL+U8cUKZek1JimoYCj6JMJbXdaQ1bj0RCwyMquxGPBdG8aTcA2QCgyqBNY1puu
F791xYmjnuR7bgFZFcawg8JSZivgQD3aLpD3Mb4SKtEoBhLuhY4zc+fb/8NxQuGPdpQmpHyiFm/F
2ligGt4yaVOY7bG7Vj4ePuislETYrH6hkeHl83UJtonEi+kReeb/u0z3OkAe+C06g9eeNlfdSiA2
sT1KDt1J5NeLNq0+M8wMH6XVI4d6ztCxaa+vxOUmFImNE2xR8enUsGcMAmy0mFVlbXNkMdSPDVOB
iKx3ENxfkD4iBWMfAmxwHc0r8b4F/2Hd28dIXV0qyhq6w41fq3jpzF/q4d7A/K9zzJ4hZe0rGULY
qMy2arteW5izBVmZ8vhVxfBBZQrRAxq0Tf1YndxsLiEGYWMqoL2wf5OGMND51Rd/2EaEwGLmULw9
UDM8ammVTfWzXdo5zgSasNOhUPXaO7+xcD+ssHrR9OyBrd3gZkIty67RiOYOms6hlFHG+NPmhVMx
8pVIfHLa+iJ6J55+sVUTdNFroWfXWt3qH3m1r4zOZe+kzA4Ye53nZQVas6FmU98oFmerSVwVq0oY
K+ItcvqKjzm4RF91XGSeBWUVpf2e+cLUW3bj+uk+JBxv4x5xcjhWxANQV96VVixXj71egU2yzRmQ
kzH1Gk0GbGKOxeKOwhcCnakCVktGSwnmwPJURtMcSilUjTizBznYxy6zCTDQHfb8eX9he7wcv+Fn
pZ0CE+o8sPGtn8RPfpdei+/lAHbPTYXnTd8Vvutp2rduY1tOtdfcV7Ya3qu11eavV9XRnzu2KCKM
2X5uPqOKLABQ6zgPHrByDXotinHjKAmTHaWCT0Gwz2rEfoHtLPNF+OGq9LHSda5qFqtTMK0rZTBY
BShHv8i8S8nA51X9bDsxA505EfhXskZ7MImAUF5gPqWI0p9WSmYkSlkRuyahE7fJ4LzIkfeSp5yr
1HdP+R8+K9ZaGw2YyjjAEJK/LZIU2Ibu7PE933ibpHZ5gcXQMMCWD4HTW750ogSS+zX5SFQqJk3R
I8nIma+XJKq6tZv+MSf8J3qe4cp70Ay5/55xZmsqJ8qkA2l0lEp31wjeLtXg7NfBcCbU5jl4RiEf
wuOjkSf+IbrNJtRKi4fY09zmJYqQuSIwkyF1IUXRAUx5am7cpM2vFecp9Dru//fmwHLZKyZcnsYw
RmuGHCgOl5LB3hrDbNLvCWATxp6Q9QuSCsfle7uTWGZinFMkA7Qke7Q2x6ar1r3bl3Zn+t4CSArg
Ri1kVmyBxIyPmtzhgpGNH9a2bAgR8ggoGDT0SDG0LdI/2pTkqMVsPQv34Oi8688bd+ijPJUtvGc6
Wbk4AWApD2f5o7Vq89ArejiK9bzwwvX3olUwmvIFIp1DcslVvaWWpnNrYIJpzbJQ3mrymW+68Knl
8pklCcxkP+gQLMtAX5nLl10CJ4jrOno90ipuuOjboNRYRe7ciG7CkWbupx60tPLEJ1BQukD4FrA6
6n+l8Xlbv7TthSXQw7XXqoH7DrBbzPaYU72LJEKtb//mstN8MqeZiBrei/JL5zF9KPZoUFipGYk9
FuAnMqZRJ2jYLVA1KmigcId2Mm3zPdOA822ecTvHQXGJyzQxxOcLrTTzYtJ6Y8BA2HspywOf5xOp
HcDPugZACS86k+L1av039uKonOAXPJSc7HlGES3/TpQ53ZyaBrdukHK78KdMx9DMTDvbaeJjg5CZ
tEPI2rLiP7ec2Ti7eCcAJB24FlYQCDtAwbPE/MH7XpcBrfR4tjBiwtCE4jfQSjKvn6pHBMHm4rFh
Cz1vdosVQvt2Z3+W19Kku+WIiUZ434TTR8Osi20qEwX/Wy9D7VS6h1ew8itp6eWwz9eFZSvT2INg
T0meob0UeZFviTaFZkJM5v0okjYVnC2BTmkoyF9RbgQPdhEG2lCzfKQZjtZ39soD8BPYv8KTMRkh
4ulgLROqNyhkYQ/TcC1HAhP9qqYHFyw9Sb5dsSwzlrTecdMCp0LRxd2lwgy0xxVOh+BRFVWFCpGO
iTnByZxdbsDhHZLTK356vrcVvefxoTvRR1vuoemAzzwfyy2TdpZ/P/9xAQ2O1T55hvvnQXrRpjFH
rJnq2c1QxsPJtRWFJVg2w9vkdMWx/gdzwkXV6E0K7H5tFE4fJjCUdJzM14kvQ7jrCM6Rgg0yvj1R
SoqEqfvby2JpoLCl86tQwQx8CRyHHIcTnjhW+prOKLyQsJ0TbnzW0DNkXAxWBB8+/h0Rpy3kXy/d
pjw7RNYO6u66wDOI6oqKRjNb2d9TbLdAWmm4JBH0860vB1LQR4viXFN6p000WVwdeO3F+H3H/WRR
A8GVYMvZZQzLOrGSpdHPRe43vYo6D6kPIu9QbxI+5B50BSKu6ONmuUkqme7kMK9QfYBYs263d1ZN
0/GobCeEPrzxbR2Z5UcHeff1dXgG0VIHaCGczyd1fW5k7IEbab46GWjGiaAyBsnUzJuSCaSTXmnU
1Xs2NUE83F1cJwpCi8frZzrhqOyf2KE062iQQ52NsOfXV1a40acIbCZ6YjlRRWGKyU6Wa/P1JQ/v
neZ88z6wNtlfJ9Jq05GYIAhq/MmvzyiU3hI9dDA64WBb8QmN1FXnqrDBbKHlj9fMdS49dm2Nh0Rd
vZPnFgNBj2bk/vzaSbQfX1tundWqBAm2DoMV9vWAXkJPOaGpUk0tEFOQForWeh0oYJsGZYrEebkZ
r9QLRibXOCGs8VtDAJ//lOwqevBoexWpUnYQ3vokeVTc2Dp1VO6kS+xGf29xtm4JotE6rHuG3Maf
4qadL18evYpjoMEkuPkibqviRIeza0jAH3ZWE9LvKWnyurzfcXTKDiQG3ji/5vcu90l8ctrxopuv
snmaobZ2eeF+ec7TNKHIYI+RQd9wXlsX3qi4OE7gADUsgmR8vUSSK5hbBrwf6yRp8jCs4xsQBMZt
o3jJ6Dal83b/SH0VjVqNvXBswRK/CxETDJhyYOevaIStEWTIznoI7mi/fa7sCuVFsf/CQagt/8DN
DjBULifPgw5nqKm4xs4wnic38ew9/g3hzXvMmFk8yGojSHYvNvWEBnA7RJh7bHb3jhScQqq+mubb
HDroiU0VsMdOKWPZJW2mRLI8nlY8hWISU48iImUIIV1Teh0c1BK/kTF+JkmhjAfveeFwS2yTiAEf
aubFUQT9r2M/tf9uAVActbTiaprksu4DPVhUd5AIuZ/ZdnHNh4oGK/FU9KZNWa0ZKXnvl0QzqgGh
o9C+6mJ7pGSA8nP5z4QIjESQ+iFueTxPcl2MDr6LVubQxHmkxFrSjn5Z+7fa3voKewx7AD4DBi7+
H7IDuUnKuB14DAh8iVfHCu+MQjwot+egezS7TJgd4ej+rw7eJQum8Ud3Bsm+Myon6Zgsyn2S4Dmn
annB+5CPo7cwvpWat4PtC1/v0U80niKuh5fZl6P3uf6+xIBkB5PQeowkmi3TtiW5CS0fX1mplZmo
LTOAbNg99p0eJqDrbzC1JFmd59/EBRCe2mKwIKh3vkEI1prP//y6tgbEtSL8HrJzz7szdlCFBhcl
aA/b68lKm4km1bfmKRcUXE85i12Yke0wKe61BNABuO0xYJqFUYSdDRBbm6BC1uhDEQWTvcM7hF5q
gbpY+Pui4/7tr22rKr3/GWjjZrlbv0E8u4NaKn2bTYzRI4reGMdzG3YZ/VxQ2G+nbUqZX4Ua9Iwc
xIIxUSwISw4Gu+VbVjg4sZdg5E0QKzORoe1pHwEyWbJibxgvj4Fm+S8/4ZEHDjVgchxrkgNWKUpi
t3/lz0BeqGLZgjJVJ7LFoKz1Jz/aUpGPCbFs67Dm3N3sqPXXybVYBqflz/m4ulPjBXxoMaiKxcI3
aA5pCYyjb5zMBnShLo7Kp1hZlWMhEj3OyKNhIpAemMvGSIgybBZW57KN4rDZX43vn+kipYZTvGFH
0EtKHVbNfRXfnDzVxY+/cMx0RIm58LwcNQP9nG+TO3IYM6/+54oOuHO5sAN4nKXUB9X9V0YUS1Ix
HmA5vX68uY2suRltUoL9Nbx0B9cotktSr9qgp6x9SyXnrCG+E4jl+hrmGxasq/3SBvxpMDN+alJH
cb0qCT4J9n5paU8MJpa2IwC6oM4sZgQaJTHp3AzLmvx30FphsEo5Zt5Yj5NtrUAJpfpz4dcMzOwm
e7sW4J2S0kSBcRCnT9p5Y0LQYaAfU4SymzUrxwY4gvbInNlWwokgkzxvOpimCkRx38HguEUys4ko
c70WjnmNLTY0IRWNPC3LUSf4JcwMBZommUCdj8NXCxDRhO27xqLGdhB4KUFfCRoW+9hPInlHid9b
l4c79vv1a1Wf6rIypqvChgg1My5WLoQM2E60eDnnhz4+kckm8UqlcF+HFl+LTl5v507jBPCCY6YS
w6XNdStp5veZ9l4ZwR1oj9jAFhYF26gfycywFSUtSjb9onZjcwGHkg1meQkGV/HZR3oxZuu6tw+5
x3IpoBm8LdO1b+5huQPatO+KY4P2AXcBLVjvFAIUrhdFd3vxeEYThVN4L88xk2hBd09FvcBfPHxz
i8h68Upy4trmgGn9AELatuG1ZCbDTm511via8DIsqGndCLfIAljzdrmSnMzELaRzcY/wRkJPgn8R
l40kqtOCeOxy3mMrSYCML7vIVnb/PoHtrwtVR4MzDj2hndgezXOmjkVjGamXc5nBebpOEoGaOv7D
/YxI0x/JZyJKqArx9MOER82FiLAN1Jhc1eA2HoOkNd/adXVqG443UNBG1ow6y7dqf2jgydW6nRlE
bobKxvmtRGwe8FMLAVR+8Ba8tY6EhuhAIYlMPCW0A02vlM7mb7xHaG4kbq2NhjbEvMuArqH6Q5+h
1t8xwB1pZjjnRJTpwqrHU/EmpcztJ2HehOKOklsOzx73UnCQBzEz0R/4KHToOv1coKM0iXiYG9sv
SGYu+I/uJh/R22IZXJlfUkJYJjgV9ciCgzzyCVrCs6C26IxFI6TG5uzEtYo2mQEec9hAR3zs7CST
hyo21NzRXJhoECYC1j/O5yUjdFJb8sEnW/ZOJgpvB1zasBlAnUvqemGRyrlYq+IF6OBnGgHh0+r7
w8nh2VVUQKLOaUh7QHSgdL+OZOs6R7woVv79Z2knhP9oHGdtfkhW2tj9ozXIsevl4cY9FjPC3tij
b9nYHAsiNVfSFpoUIBxdloFvAIGJHpw6E13rR8i0QlS8KbocFbH75jCqaNUvl1CgbxY69Yhvt7eJ
SfcIEP1XsiXZmJ2BHmOcr8uQj1UI0Q95bFB3CHoKFmLNxSLe5jjITn+NfDUletxlkBdM/qrZb64t
YkXH3PUuqf963Icm8SBZWQRvp1bCSyTCfAZkx/fhKgAVkoYJmMsKvyf4e/98rG8ZfSoUbZG22un2
9q5O3WFpgOXV9OOeYfBm0Vj4vtdSkTU3/es4lbrnKv9dMTqWBEe0naZO71ZLR5gR+reg4Zev7VdJ
672fA+ACY0f3Y/KXK31aMKlvBL0fuY/94xZCQIBMa23pFX0L8o10kfChDmKUG3ZGwvu5yzNqGlvP
7Dwr5pzwxPDE3GzYz0COK7ihehfb5o9WkyomUIElOtOBdSbPhWs7/7uftcV+6EUBvDitCwDDAtV8
P64aWx3rhDKnSn19o6IEmVQgePl4TzVE8wIYLLsaHEK4r+yrmy2gHf/7dxBwsTahhemqr9GK1UYn
Ygc6wv5/NzdHfmV4yWlAA1MtUeK1UYLO1WGhg6YU8V8gHLATxFCNh8Kq7S7iY1y/Lu5kyqafvCKt
Y5afAUCW6+wuipAnwRuKceKPmSyJeYqWZAB5eG4o62GGdzx9POs/u/i8pWc+BUd2u7w7PAhpzElB
tVj/DtVtPTt3vimKE4x16YMAlnbQ6GLg0H65HpBMjEXDswx299M4VZsJDG4pHnmwPPmIrTraKfpn
A+marU0Q/BDY9mtet2P6OyQXL75CqAqB6aJPxgXdutZqoa7slHBbZS4ArJpFiyYQkr7lk+cEKw13
9WvXHi/8HbnMGDcr0VJ9QwCrN0+yAYBSOq/HR4RziQJlxQ3E3R5iOTLqeB0vm7WONMhBrG4EFLRd
QX2ZTFyYU2ylFHOyaycm8Df1nlNmQUqmA4gpA5XfgnF16JGSWvtSln4SGLPrrEg8tTDpUHEViAJm
dZHvBFq/7yFwWb8AO3o+09ltPn/MtizP6p6Tjl5i8UzfOUMmAmIyLiP0++ab/fSd6P+ACY52K8aB
uFWkN9ebdB48POVtLsq6rHG6l/SuL9qrzzK5qQNcRTmpSOFh9dqWR4tVCoiQ9d7VVNyZ+L9c7aBv
lSizhNm+Py3N9jVA3uhjVUMLT4Xf0IMC03/gyUCyeakLp/iAefHPW8GB1URt+TGcoWx6wmkxYsid
hn1dGynONVd5D331qxJlP9BdSQydSCqlsQgWaM1oYXBx/zWT7ztH74IXKGavQtoFakwusGbmPs8G
VZ/yOYGN55NBFiqGX+Ou08/BQUr2/TBQNshLH5Dc33gCxMR+M6BNa7gk5Lwe2lqw0/YsxDfwhQpr
oX1PDaq/30dVOGleiX5+qhc+3wcAoZVwPMSgHo1ApcRzFveQvS6Pu0S7TBQVL7gX+MRPg/dxioC4
+MBUwvSWMAXTwL0kCJpO2T2LGQwXsScviVf6p7ep5BP+riii15LTdDwTf+1Qd6feneFm/DjUqujB
7/oBWxKAWwivG2bS17lU6fGWwcb3mWV94S7YC7hPLcBC43+qPab7odYDWsXTDXvZGGr8fQ1aWF1p
bBHVR2f4oNJ+mN+Ld6Mx4WOBp31fJFpa18j0aupmn0HQIawhTLRrrqhb1BGmD1g0e97pARMZKY1L
RaqGj3mc6q9FnnxqP/Jq2zCPHMdJkPMKutLiYb/TDZ1Y5XptklRfHTsjqJhEd9qfBZq3nGILQo80
oBm957SJ8rP5TVlN07hZ1risdDttjRR8IONsB6ryIeRyb1pp9/2wvSTX5c9mn/YP8I2NivHo5VvH
XdHkNf0hh/ZolNfQVgHIggQ+bzdwrvYX4PdDOtp9Pa9un/p92I65WdfeKgtrKTNeuGn3Reu3+0uC
Pk7qTlLy0TiMt89TS1xjA8MeDaRp6EALTcHw33r08lLszkOfa1g9dH1RH2yF8jXflmAUUSzhQNbu
ZeIYuOQEatIFi5myH8UcHm3D2x/fHQ9XejMC6F8TQe26ZzYPEZBM+E4LpU4qhfNuhYzE5x7GpDiV
EFG9AxlLI9hthPh289iVyR2Numay3LeV82y56QcfvUNo3ciJQAqkyPFmGozl9v/4pDqSN1bmFRgn
HauVz2Ie4u5HlURoOD8KdOujU5W65uWe9J3tlBS5EdkhB+K9NGq04Ymi4+EmamQp06nC4KEnH8HP
rZlzui7155au+TXfjuYh26PZ5MO0We3RLV7Rr+LfhmNfBx1llWxRCZho2JUGEBuzVzmj8fYzg210
krcJ36/XPWbGnwGwiwcZjJwLl1io3tDS0RCxa0NZWURz69UXH97msDM+/eQVCjKt5m1MW87c5pE2
QMzS2Wj9fNbBX5wD1/23EVWWkGO8n3QMZV387dYnGwTSgKWA4qZ9+gD4S6SzWQK3mHZd3crnVYKw
glMTvjpQiLwPacxGcAtODU2l1WV7m7HYieibMoVzF6NZCOfQlC9mmYmTRtDYbc/t1IPk3Ngjluh1
sSXToRpc4Od0jJMJMeQAZ9ARfZjrsrBkUuApkzfKT1l5HCbg1K1R32HXDtIqtPwLYPVJ4UyP/47+
VvlaqNYU01fvrVucOkjykxBLh/Q0D4v7QlzRbxj9iLlDipCga+gDMb9MErxRr4TVCI/YImtMLiG0
VhMIp+mDWbdue8iECEQ0GgsVC8LY7tz6lglEScWCUguUs3UACFL0+gCf9yqyzeYo6zv1Iq+a4Cij
xv/B1AxLiRzAZKSF65OMBuZSnrZ1cN3bcdhV7DRyCMM/vOnaKpST41yeaZSJ122Fjk4rp1x0gAzZ
LLSFu/+kDLcBmrgHXxkzTaWgidhZivko22VJvzl3OSzaDARLcGSY+hBE0BcfY/DZNF/Ug6bcN7L1
exFFMo2rkWHreDfx4tLDONmVQNJKyXkPA23iZO7dtMDcrTzZun2Q7OyLDWIsePNHVHm8zj1oVltA
KefcFSg0klnyDXjx5poweOQcPgmSH35G/98j/cMwgyG3MbSIqDgIm8Iy+TXSPKFobTu2MdDWB4w5
OHNwoBijgvjZGjatiBg3vbNCXPDd/k311JDMxk+QItw3Zkz/2cA7BFHnZgez8kS3jN0qYK57JzvF
fZNobVso32HIW7ruUAhoWYrkpDkrFxoRBKhD3Us3UTylyR4yve2qtYoG+ZYpjbt1zb8ofVRQe9hA
gFEsI2fYD0/yTs+tbc5004nndeVenuxlOi/CmjDFdowATYDf4mPRTPcOqKpQFKFUGLc9jWyVIwXm
/X2WnYLiRC8V2U1d7HgHaKA+M5NkTLGkUIIY9bfZ5oz9WkbbO26kM/+UMonjmFnNRnl4fxuHUcg3
o1zM17H6ou08kQAmXjTa9GDRIrutKOa67b2YSjJKaIM/r5kHX8LswfDj2yXwv80UeG2Lv9KhFcCX
E9JUUpdmsEmzbf5RAACin4bqoQ8BpW0Z7K1q3yZOzUmS9986Xp3PGPikm+5Y9WqPeqq/kwPOxpvQ
I67Liii67PcmzxTo6BeAe1Xcq0+ISJ4wo0vOdq6UTLbgrBcCphT1TOuEsV/WhFf4/QzGMWrwKKsP
CT8n67zLzbFMO0ktzVi3NSZHx7ioejCS9alDG6D8GjwfcA/vwbjqq6Aaqz3bHxc95g7f7ObkVniT
f7mhW/+MUa+7zEkHedHMiYDhb21m/5iTxLd2tXHsg9+1wNYuhKWtIKG6kIjz3XCr+yCeCGqmPPxa
TNitK4VHHjYkd/whvaqp6AD7utSJwySI4yXg5w8JMriR18jbBdPniHrcNTWwx9DOlvkVcbYJQeaH
QWoGzfv4GIOW6mJEH59zq4g+6cbTNd82Vh9V9dcfMKIKCAvJpYIumwH8jbXwZhUILgHsFEBQ9Zne
g4OT5tRBaEfSjx5rtcuR5mN88BEMCkbmFfGkz/mVmVog4MZdup0sFOApDG+x5kolFMbJclRR6654
By2IxfrLGdBXQmqoWTKyxkEk3TM7gshI4wMUXkktyCxYcrig/P08KXetQSg7N1UyH6pzQBFDU50r
M5IqreBTRZBh/vndA2hSohEjQRG9CGyiUq7rDUBuOkqZS2lnSu6EUoPBmK8+JuA1/k3QgqEmeNsM
vOgV4bzJ05NImrb2RxXiBgVT/rq9IgOy8sF8DidZlhmesasgdFPX7iofmLm60jYpnYoGWYPzJ/bq
4jjEsyrRlMkt5dmsM6xod0JTH0nAbD6UduvBIsfCqN7+a8ISbyKyFwr95nQlBsIf1twnvUhGUExz
2fB3tENJ7z/mF4bKDNoe+ydvzHUDGxU/YAllYiK1GBEHU+WjCtBm0Hi9yjPQU+Ytho4zICOUZTh6
suWp6H30Ecgz8qTW09ttqvH/XVl/ogFC1OIhiZwGlTaVbxHv4vMd7rBhhHKo8Oix0y6f3iMXhqus
Ob3NVJHtL0UcYfeBFrYVAk/3mQ6eT3SebFDDchOxudAyH8HsneowohT9nO+El/YwC5xPefAFzQf2
2RaAPt8lDqrQy7kSVpRoCkKHBnjoFvn6xaR1Py23vyyKgYdGrjg/IcANrYTRt9x6NaKNNmxpYAZA
LkX1MCj2pWSU0gWDr69GEDWAGqXTGQR0fR4Ef3c8c2YNdrjkFVhHs9g5DVkj85d4hnAXWr481DI4
mEe8zK/WTCXCOjcbE8b8wLI4BxXjWwcub7hxwCq5HgNkSUan51XcHypCsiliIbiB90YYLu38xCgW
4ww3W7HH4Mcyhkz7XbcE26ir2TzIo0/+pk+V4P6xgKLS6sR9zM6/Vsae6sh5Ez+PnXSPcL1CUw9i
5EocWg0H7EtEfPlD4QzGde1ar+ulezcTNJKKhoCazIoERDcJX2j1TivwO/VtAB4mDy1hIG8e0b3m
1y5vaH3S3HM6OL8jrdO396lcwRDzOaCiIUHHFZbiPXA3PcI/tIX7dDlpn9Qy5hQS6OELuKIm+sFA
9H4v2rgmDQA1WLmoecsK7T+42Fw2PwKZEcYI71JzMsgqNwKYLG47x9Mfb2ut/ZHz4OGYj9HWX42J
Nm7zQOY9F49kbEwZYVnlqm9TQTyOCm+9DCbZUD/mhZ3euI4IgnNctKEdLhjGrBrh5DMueZLfKggH
fa08cZQti4SjXWI+uIipiuqZXO9ExJSXpLRUrsSWd/BLeJGm4lBnXBz0eOTDzMAS2mnrMy3H1e+j
fWyKdL8BI3/j0w8EQ5+ZUUx72omKeRNDIyUxHPPzBZ17+xAbDl1gz40TtzHWv74wPWhCGxK1gqEh
skNxzv3UukAnvK2PuQQEJQ/eyR0z6A4XqI8AttBSfnc4kG0F0UlCKNSSf2L/t8fkjEQWLY2cdFp+
je1q+v5WC9gBo7saF4uB+FbwdSecGssHSprZVsRmI69uSdmsKJodrHoEIE3QkI4xA/q/UAWZvIrd
+QXPieGxkVzzz5+o7dZPWzhm7gSimQ1LWMN8xwvG8I0vuhtzWduFHE+DrymvdyVwi+PHNhvC5EPO
VJgLLMwM7cQAVVVvp0jkN6VKbF2R55X4QMpuOPHg4MGnu8uUkezUozjyLBdJR7XnuQWZdCIp0ppD
JNIS8H8zTW9h39HQ9jL48jxncOPYqpm5rLCmngrzh1tFgltFsGF5Folz7qTNXB7ifCcxbMUHloxa
a3ZPqnOgd/dl1zNpFhR4R6JPqUSdx81+zKh9HvhFMvuBGO1xpdTr8/5h61jWcTkETkHwzMmgjRVu
7p0lK+dp5YRgURs4qyYODDAI/TYMro8cY6PBmz3fjWz2EXhfJsaq6BW8O+CB0Y+wmXrjBUh7hr1B
CdAQu34uon1InDLf6yL8pC/kpPQ9ujP0ZLoKYZDh3Qb5rYSJmewE/Z5sJOvZVFjNQFcwZXGz9rVE
z2zx/9sFhGIMI8YxkQjHcj+/WpV2Wi/fii5rpZ/mpnlYndNLLah1m3Mid/K64SHUzcEWlC25w4Ey
ikdmxIx8vXzxGyFm0p71gK6DPYntBz3UwhmDDTCcqFcScivk73tfwZZwryDQ23y5r7QfN5PMimKh
5k8k7uYQhv4pfioFOOzzASa+zeinsJkPYG5UKdhFdy2cLJuDcxps0LEJAdm32fyZgqoAE4S5PZwc
fnvQ0tRotWgnZh6X/+eEAwfMVT8gEF1EVwjHCKZkuoq7TSaIEHnkVK4ciqGyJ1B88eMdxbIbvUio
DkPXyqy7+qZzXd8fhonYaCvmlZmiZAwn6xVg3PfIFxSpZXuJpRSUc8J2/3oTy3hAz6G6nvN1dNeB
BcATdPVnPcBRP3PFuPOC35e1JWPpTk1DzD4iY3qnAypO+p4W2cpDqWLdJ/U+5iyitEP8P5EaaKyf
GuEVnWud1VQlH+DKotH3h3myVJr9R8tUEzP1tHe0OUffLoalBbLO20uVJrv+hoXE904w3vkHLRL4
64pu5hXPjUpeXGnLnAmXsnuNg5MwEO+CBYL8W2sJEeajxQPeA8JCSwjTJCShxgBiOQfWW7VR8gou
Zj+8TR15I95aZXgECCW7lOGYzkpiibRQP/Zv5hNBwNIUUwENcm2UCfSq/kvGwQSVsPZldeY8DCZw
oovUvHbaut7IKwsy66u/Pu7daofjH9gMKJ4pWya06yn7jlpOB9jSas7nMMhDGFfE5dsWMlxOxJ01
nIdVk6kRFD8wgy5Vd+TjjSbXBqAI0ZUBvTtJnVYqtkj2Mj1ERrZSFiYPxmhE8m1rO+qvNa4AKaMf
L8+DKV40tB9AzPU3nuwCpunxSGZfoWe+R6kAB5sFzSKQQ5ZOdPYPdntNbZYBcNTpzwDu1OHIaaVf
S6h7DGiLdpgRFqpowbZX9wZ1yusVPXVXIoAmuRSJsQn6iOIHLDxYS0TKronxR6glUArdKvSKcNUC
Xy3IB8yQVBF4RIJjO0E0z+QZnTtODXg884j6d2vtT3KikHK206HkaLRJeQYb4NGowUmylcI9GRJk
iSJNEl6gPXPTWWMmRoD4icy6NeA7rdpoFOwlhJKNqaKCnJUrzRCTKpU9KlFFmI649gED61byeBzw
sqC7bOF2z0zqLYYJUX9yRgeoBvJ49eYKhUHz8/0eTU8q4HrhB/OW2ZlehJsacFf3hfr09Ve3ldcG
w4Yi0J0wWsKmPrBUbajs+lGVVhD0NAemee9EG4xntGjCUkw64nsZ1pU4kU9H51MDxOp5kbAQC03r
xOZaNKAwtHnWpOGMXyci2wA+P64X1FP0wIAVtreWGzdj/rYnMC5yAVYeJ8+4tJYUEamZ3P4yBnLt
jwM1fo77cqRiF7R3JfGK0KoIgn+x0Xd1WXcnTmIFy8/aHgx5CntkCtxcnYEdRsJJ9KSt5JQ41Hhg
2HPWBonrS/RhIHHYsbrJcPm+0aUDY56QnzrbBcjHY/K22uCleVrxXNKo6AC8pFhd5ZDv8tUqkzKx
fXPeWvrbS2DhOrCQr9c8+Zl0UA93yOMV9iI9mRzjqCaSflhkBiqZeUlHob8VL2VjQSDNTPQ+MYMF
CSoTrP/la4x2FA8fFVO4A5LE5VmUtnlnpVvaKLMFfGamle+BFRk9jBPPg1ngqUTsUlTpnstyH8LE
AF0MmXYCdrpnue1gu+taQaKR9jPpf4mOvGMydPEny4ZswEU0uAIAh6z2tqx9KapYZdvqWRcZmEbh
rd2ZLWxTivbIhdZxYZd8cbQHWKAVkWz+Tbuj6gGNXNVbYpMm+JMleNi50DJFDBbLoGlqOrXASU1e
kP208/ygNEojnulVLCy3u6PZHXR335NbH4JJOxwJVZvY6J4i4MiS2YVK437PO+2Mk6vlKTD2FY5s
8W1qD3XOlvLoYltGox3l917nuY4fMWJD6TmX1QSB02VIk6oopZFOw7PPPGvxLDo0lUf31YxnTA/l
PgO0mTb5cEpu/BUPvQPNKITJLgfiThUg3NGT59bkZymOniUjcmhIXMJjG4oug+ODpQxR3gOh9K+G
Uh1Q1hAg8NKufqWEBrfu1fdA1zDL8t5yrdzr59Bj00glZWuDD31UUyMPxONB8UdcYVOOEgcmUDvn
G/A1fVnQpBhvg6xduSMZnO854EzE6Gx+jlMvCHdt2dxcsfQc7o3Fhn/iaSS6OUJM6WjKw1twSR0G
ygJ1+GXjaeDWUJc3I1/AqOBUo03BRa06ZTjNSLwHEZw5GTZPSHVwCclFgb4u4iMOebTWS+K1vl/V
03aDuEljvTDAjXumZ32J18+vE2Y0oamrOHgEdNEDX5XfSU2TZtkF0Z+sZQGIt7cR5H55rMmK+/oe
u3+9fcK+prZnPCpcst/9F2dsgLcNTJat0wWIjbMLpDoNyRXbajX6UEIawYuSZdmrFNcleBg6N0aG
0QK6QHkjS4mzkKso9Mbl06EiNUyr83oduGdMhO2b3ERazatkf9cgeC+WTrN9PXaYYVEqeKTOUAsR
3P8ESZkAWaZPEqmYk/NlZ7/v4YzEdBSTmD+WgfB05tlPuD12ziniZGMIqSgQt2dfiVpJvqIt0Md0
bDPBNrQ0tn92gYGcPex73rEWHqqhippD2aSjtM9KQ5gzRJi+htBqslOs8nnqqMDyen9/JfXbG/uf
yubJoea0uaagpDwysUqDJvypm3BE6VdXK3MinbDOiFUiLTXojwYuUICuzAlTKK06Kr6G2p0PKhNu
MUx9eZwexl4bHn7CHgC1JckxPgVPfEb/lqe265eSPP069mJUeWdhcnHm0H6k9+r6IykFn0kzusT3
62nHBCzV5+Zbe7G63lCk5rlw5cqJukFPM5PUm9ODEMNs8LCo6AlqRua5q3D43wK7ZcW0XJn3NkUM
V8z5QbLqbMWugzVlRFLOZK/IRYNQCPnuiTZvCnmNe0MXtrPF8mmnD4EHCOl0AeONhlEMgmv1Okbi
WBkK/0LPqYHLmGmuNSdYvl/M8RDG+Us3e1C60OrETuPpDryVyXFBHmzHZYQ9LUOYhT8OW3SHf0j4
6nW2XjFQZMo/cSE+UWvUkSAH2buc9EcorkdMKwhZ6W+gEGzaAR2shgnp22ZsS/TQEHwAbtEZBduX
X0WasSXLch4cgt4lUewdpjwIjPBQpps0EMMZM27R041KFHrsIbNF4EJuMXAcaIXxffDNfVzCKc2i
hqMezt+u0IfC8VGc/xUicXv6aCJsyb/TDgEghZLu6ncvDnuAQBQzV/PduojxlL9B+XrmZlokWvC0
RT0tNzdK4u72Ekwyjgd37paBLjxGT3PjoB2FMevFNouMv4mB9XDiSukvLR9+XYwUs9Y5gpoI4Rvr
4l0YJz9Iel9tDEg24HvBZIBEmzZ226/vISGV/EVgAEd25f0EVNMSrjS1iN3mUtHhQ7TgoULzvwbP
vIhLhicThxm0SL1Dpdq7RKKDlS7ACC9P0dEQNBSoNSEVPzR9PQlviqbcSm2KMYgeDkUpYqjuAzeO
619oETvhD4PgYlzDQuTQOu5yvQ+eRFj8VpURNBGHLUYC0qNRLScH7hTh7PviydDanWgz6VsDSx1c
xLw6VguXihasDIYYQBzoCkA5pIcvYzfEqWgPe+BwoTP1TsXTQMzbKwXqMOvTo74Fy0lNynljPOi2
dfThgqHKQTwWH21Or6LxJx7OlN/H38x31JeNubMQ5EUABOprhU1613pajBG7D/3N85ARU+1wu7FS
6uu2kDZ9nMyzvxvSBWbYk74FFq1W+NFGERB6ulxplQ4FjSUtssWgiJEoooe41c9+qx3SgBfQWMBy
iGFFUr9VP6ERn+OO0KwVHOqaNrjHUJBbE4MaDQApi6eRyMhuQ5sHgnInjpQf84JujBGexnEn0uUv
Z1YK9fMURBGrqd2Ta1gTgRmyGwOflMipXwjwYaHPAEwy3Pn7712LTGinw8Uqm48HXBS/LmG866kb
8cnKfu16DVmUkk9yl6EZkQpkVe6QuHisnJJuFndnB8omRev+4yjNLudDNbr9J8U7rwbUiSjSoNRE
/EY+gniP5jAJh36AOhokP3pkfKZcN7HMnCSPG38cxZcDMhbi1Ja3+hsGwEptQeQOsDst6re9PYJE
/NkU8A5aazoS8sw+sNtYy+w6w6SJj84uIj0ZormIp/aYhjuPQYh+XecajINwpZNvUeNHVI1Ayd0L
pXMTCuVMXSOr9zUZMaCm7rrLw8bgaIRBVWD6DvRsYjYq/AaDi0f2vb0BZcpi9+ExY/HX6LL0pjrT
W4tGgfvkAtDmDSGsIuMU/Yn/XmdjuYQB67RzfG379qCvFGp5BhRGvdk7F2gEoZ/JNdPyPJXkA4TE
Q2Qz0Faw2xWSYuL1yQ7LwRA5UzIoInjLRIXGu35BKkf3l8bQtXS4jokS1X4vO4Q3sc3F6G8vU9Ho
va0uMQSm19/suxYEezYNb7W9gz6DuQx/qlWaGOT7CS2MK6JMn1Jmj1SB0H5CHk0+g6npOPVYr+KF
VQWCDBi6xFvCnGh7Xc7nXKl1ivSlDWVlY5jlDe7SntBrTxvKvAYgTBQlrdI3m1r5VU6vFqnhC1yg
twGaH55hSwRMADbGJeucS3uJbnbPbNBl4CegCDxcXPHo6bIhmCvCZjb4YXevyD1ICd0PpBc6/aQ0
ND++4UAgVkgfS/PNWHZRhez1IZHvSiXEBCtHKs0WTcSDxhcXomIKmUsGiLOEzKmCshd21ur0qmkR
ffLLjBSlZncKi7izOvsiIhUyQwpdKdbsxo3kpFlBEExyLmNRi/j1OHoIqgLzyyPdq2vt8CtpFbuQ
CXYM19I47tEsD9e32Wemb1vbwjH39CnEQDbQssiKDhX9WrowT+MVELyQFskUpxn+iwTd8R5xaNlf
9xPsv78tZUkN42V5dNmCwqoi6KKI7b1LS/ItDOTyHuO6NusHLQSGvpuMKQyAkGZV24nOx2jVEFhZ
m0zPklPFgUQzuBY78423jUlRCTIieYRwOO860qXkr50wHFCZw5iGhQHBmnFYf/3ZgIZ5ipz6JbEl
3oyC7jqoggtYaFKJ/tjGle6Rfg5JAvM4AMSU8DRntYmI1oabBi+drjQlcetIX1jdvmIwLsyHkvjt
XcdyMfawsHsgxVHxg8nE9J2N+DEw7/EfBAAqF+M3pjuN5i2YcbodMqMJb/pmnWhvxnYSMTG9/qSE
dxcvtfnC/MEKdWWfI2zOC+tkGwc6s72KXfUQrGlM/hQ7TPHo2JFzcoeOXe8umE+YtL/wzTlFIJCa
YW/fnXZy/MpdJbHu2ieKG52oWQZ5UPBO5i93JRv77Y0iFZ3d37CSemnxNQ98Y750Y/h2nhmKXSm9
GBJOzV1oavQb/vtxEfZhKFxzwHOgMZ3f0YGZSTsZDqt3vum/LLMvJ8ww2tCeIkmLSSCxn1tJiNbJ
GWgg05sNCzDitQjaukOq5n1mVIPJ9zfMBkJTQdTcmsVrcv+7bUvsszyeuPbgea+2krZ3TFPe5JQG
ieRrz2xfwTwhMtNqkAITkZzeqOPiB0O5ku1eKhJJWt50F3jLJAFeORNrdDjKvBWwJX+nYvQ1lLDm
1yggcVQw2T0vnc96KpqVQ5nyycytz9cedLkCbUk1sGw3XM9JkBxfxRMC4dGnlYo+obYs6OnQjtx/
tm+Ygil3nGG0m3FQTUQWcMr5F1fzmqWz5hMJMFL83CJqvbAY/be0a79dTR+GL9e5uuyTDlUYcqx2
gT8fntEEjgIFVUc5qEMzoUyH2TDhLlmlo+rT65twCPzpcT5hfVEpknXTmPGFZaYxlKI8lY+x3Eb7
l3htUDQAVXmlvCGJEoed9qSt5GXu565/lYmfQ2fx2fQ+upT9x/5lYSzUX+Osakem26fH3QD++7l8
ENMuzIcxKKo/YPx1YP+KeGkh0QgF9HDI1CSaYus1nTWm7axu7VpXLDcUIjtmHTEKRNiSWA36z7ji
eM7+9gJxjnYDCPPVDFWHtOhY5jaY1vMjCrln9GPkz3UUCRIZZqr80kvFj2MEov6O2ivIfqQ10bGl
1pZnsdjObhidZcvLNhppzP/6euPaqyBPekLse5oT0TvsKFvLPmaAiuOv6HFknlw3iPu1H/bD2Y1Q
p93m/kEPwpN81OBWhIc+RjJ6zSjOx7GkRv9bPNwmvKU0uqVKFjruN7T1rZzAMigAMKLdmQgZl/vD
dwNatg9cXyG7uV01TNWddMMJJfgLcuwA8Psr4KyifSYX6ATByv1wBqRXTV8i1jZxNewbHXho/+VX
HJSnCzYwEWkYgovDif5hu8sCBSKe/11NOsMOKGVS8Pm528WIyDD6B1hmzBhDdp7R125pGNMiyHRY
Zah4ckRIj1xCrtNbz9zIUbJVR3zgM+v6cKCG96C5PJ0JBE4k7VEK9Qr7xbwRy3/sw2o0Vs2/Fbto
SPBxCtqkaOaqY8q/FYpWvCxiWfInH7XXKVF/ARtxxHernpP0OdfsyEz+idhjZjA3I7cV99C1H3AP
eITPAymax2+8NBQRuwZxa+3oTXfsTbf38I0LN2MPqO2vObQXJf3nJhFRuQbBtBHNkL/n3zNTLpC+
qpEo0zgbjf6GPHm4WSqaPFEyYWMFSOu64ycgoSAqNZWXGQ0h+Ts/4i1L4xq9ba6LvTTzbprmHmI0
bhwMF3sXOKyNB3MPAz3nCfgqOALJg7BxW0fDgxtf+uVr/oPQxgPRuxIUQWqrDVA3ivvulO3JfI3L
dA0F/fGA/QZe1/Ox8EQ5S5rpD96KSoVTopt/4fsrTpFSIHVNCdBTJ8V1x/bFP0PSTA2cOjSHgwCF
q5QCCCR8eTN+i7UDNf3elsvE1waIHrtQJiyt7hgZJ5FvONplAoh0kvqD3wrB+ftL+wLFHl3uqpIK
NlTWPdBuuf0MchGVhxiQhpRvNMCA2ko/dk7XhnEnmoZ3FjeQALv3jGkozBXjfXyKYhmIKIAchPEF
YlxdguNz4euloyMMff6AhwEEhmWes1aBRn31FCaFpjd5Vd92Ci6HuSJn6QdtqM0dqPVZj46ywVem
qw14adnBaxKD2nu+zvnq8gxHf3vvCrg+qpnRKqPfv4/lAE762ohKFfLfhKR+7g7SUUUXg8j30+Z5
hx9EJnbRRx+1FlFqkpxw8FSBof3YreRhU32j376D52TLUNxFTHHs9a1tpyMZQOGS8e57um34WnAA
WSDFH2L4Y0wXSwCYa1MrlfB9Z54BS+s6mYbZmYWpN+yce4nduMVFjIURUZ5V9BvOpxII+2YBX/9U
RcHLCYKSIrDeDk+3PypnvQ61RCPE4/jUc2WrKG5ANKwcE+6LIr2OWoPWZxTY7R6Iq0ozr0Ga5Mq4
Bg/NIzfx7LabwwlaMo8QyHo1NCG/6iACvnlmOWAjFIpY5PZaP/i2CgXG4dUaxu+l+S8VNRQBkvRM
ZUlf5Yak6JA2/g5IGpWOm/wV/gUxJJ3nHCE8R3qbUKv+pcWH5JBg0rj4DrDI4/9glkrSdnpBe0w4
7oSu/iII3X4wKEkebskUjh8BNXmXhNxVF7ycnEKh2yzo3TanU5O4918cA5gY138oc99sS5xvB4wp
ViFYead4F5kLWpH8Oa5PSwQf53NEyKZJt8vCCZEk3nkYkGosGNpeHkWTxPKOcu3DO/uDffaDlwzA
iVCi0q/3DOxpqSrZwzNPI6IvWy+3HOYa09JDWz7Z+bYMcBVlUBpULmMh6uRyCZQr4ZCdi6WoljsO
2pe3g3G6G4IVwOR2KYCpuJwDEOI3ctgq8zKtS8eDfQl5T/WwSV+rGmdb4cWiRfMOGvbKRYMZRYB4
mbwQvK2Nbjv635ir/DoLB9MF8kBUHFInhzvThz1afGoH/IRa99HJYRe282lwC6aSGv/RzmGIdcZm
GjB/oWDkc1SyHsi++WoEe9/yqyp6/bvtfQnBo1V3V5LCWfAuy/qDxFZ9410xh4uYX7gnU7CLbgsn
0JdNpOPMsMMNag47zSzDlPG/rc5kdDkAfssYj9/RBZjOC95sj53ReEZV/3yyn+qzFlby+yDf2Bwb
gZbycKD4xm0f9IJ5zP31Z0Z1QZ0gjhTkyv1t1xLPJfaMs9LMoIy5C/6jornL/AkSKu0/ZATSToK4
JUrEXULBc812t0dVWSZnplZepwMiU7hDRPcEvB5e1FNU4QEfh/92lzpLWVpa5+QIQFWgfUywcQs1
ab0sxF3kAmJRjl73OeaM9OO618KCLX+YfGqgkQcyWaWuF1kj6TSuW3msvhMFTOss0YBNCx7UYss3
jmY97IRrfxbAedDraaVZr0JoD9cBWrCMfgVrq+L8V4lZfJcbuacxyWjzO7Su969PYCxYYzJxzcBa
h6ZGSF06Ba7X67o9iwuP1udioPMdyhqeR+8P/0eqyv1ToEXPorLe6m74pWNnRNWuGxET7j27Wnd6
88P+V/Jloeh1t3HS+afAv/VxUaIAopplrFg7nemoxi9scSEkqQbbhGkADDPG7VoG6ANgDseU3w5d
yipVD3xAD6yLVlqjPZ+tmbz8/hCRt27081OunLhvwpO0SSvbq5TkGWL2mzLtmXUnELG2tlym6HBI
QiQquVyMIzcC+ueKJ+RJyopxyzKB2BtuTRAEV/4yeFbRdjJnmiokdv3Zl8bhvhJ62Qro32FUlOmk
wNvntQ75ZFOl0d9tqjQocM7f9s+rwmHKUjGF4FlBK82cCdvdQWWgLtEq6ORa022dWw68NWAJs9XY
Jqv4/hilt9wnZJvmZqejKPsc4Sm7+prWnvXjAsJ7Qnt8QZtklxf9Za50mZUmVMmn4kiz4UKyYIII
X62VtCVY2bNbfh+TdOmMJ9Auyrt+CKLn4WmmiNdQYk/9IEM/H86jCEqKS26iAQ/wD9z2m7YaW/TT
/mCpthgFLTeP+mGGCDbweY/rE3gs1UbLhwK3wL06g/BCWmLag1agwTSvn93wuJ+SESUShZY+4kvL
ymg2gBfO+91byekFT0xGAH9ARf9Gh7IEPZ9KAqA3ckZVT/Mi1cMshCsn7qHPBQf5WGEsMgOi7dux
pzLyM2ZF8rUzgKkqkrhgPOS5MqKdWeY0/OaUlpjFy4DgloP0GxV7hgp1P7bYUkA/cjhGF67xUoEe
GpjYEPwVu5wvkvcZlTVEngmFnmMh2uwrLpyIImjxF+8Z1M0hXupoU1m6Kxgq4359hr6qxGdcUItu
K8Zy8R61sd4lLJlD3koV5IqInaeOnYk5DW+R/acV3miyBGFrH741+wAGGJrcORafty8WhP5xtm8L
uxWWX6r7i1UI9BQjoFmnJc6YflXRNwlf7wZsTuEnfI98L5KmTZE4RWVbQyXQsHNC/IuxOLoakjTZ
LpgVptnyZyq15Je2QIms3KrHMW+XZXd0UepmpqoAVG7tAqu+G5eIn8smIi+bLxGCdxd59L3IaxH9
R2Fh//bvlr4n3eE6aN7UgQDde5YypkFSZ0aGT6T4qH1zzuaBOY3maCYrEsT2ntJaRb8WqFuspGV0
61FTzfL7rtBMN0N7LDCka23QdbW3N4sUGUNnX7S2RaAmeo4HfQLpGTDZBa5lAGPgRcYoZAOqD/TU
LR02RhaYBhVtJOAb4wbT5ZsYoeCBf275I6vRdz/GmEPCiUyTdxlxJhpuTNwJynizvSrjz/URAHOF
KltCDW4AMohC5eMBknxXhV8pb02Un7Q+vqBEeaiPxgJMDNkAjc4yON3CobUWkwze9JpfIB6kmUlh
wygfGbQXFYp5I7lWg2UGSFnNZjAMcuG7NZ9c4aAkuLC7p4W9CHfAR1+gd/Tjj6TEEYS5BJrNysi4
yhGypAkM1pzz0XTrtLP0A4J9LlYRJ394GF1ZXGQinq8sBrl6oCj4VCdwiM9FN910dXhspuMIxNi7
VzGIqGNBQ4JNOGqlQEdgXSe0M6p5rMe2ivB/VkNeYJQmAGm+IyItUYHREIBSDlTnRgShiHrtk0KT
tbExls30qJjllCbKKmM4EPyYkt8gU0rRq+MdxsLviXydwx12uUpScSa/XM1PMs75OAztT1btou7y
RkM0zU6TJlsOj9qKCEcEOiGBMe7TBMbrylCO2uSsdshhaGUMYV9cVv3lO+d+fK+zcqWgIQr8kdQt
fX7w2FqyUMiZLWwDJ20RSnagMwedluxe4x5WYq9ZtEgoJrWNyRpoi8VXuR47M4pPMswOTixmBbBz
0zb9LmOCJrYATbgILqsD4EBnsQMprJSd58IrHnyiYCNqqFUeRX1RT3qKibY83GOKJCrXPRoyKrNX
yedRaiuW7/l709mj9q1TCEKc3+W5xaZWg3QeSJZnagVprcobZsua9oF8KRrgqmUL8sWyyFUdJ/fc
FGtQNqZzJTRqoj+YtaDiVgPc/2ZDqJsoXnEB4Sbf+Rv348vw7igrqLw3qNMLa0qRwPYZ1Pa9wotP
XKfmqdexYJ2PjrOpnLGjLoA+shzfQO3qCoM0dACjRbggZIdQpY5hSJNFucG2PEsYhM52i6bu7c88
6Hz3vIUmgNgKaKvMFT2ytztyioSRmy/G3ZHFZhXSIwk0YrZpSeymSaEUZ6L59cf6DerpiK21JsX1
kNAqOh/H61EqOgGnkbS6shrt9+EL/iE5nuMqwdgx8YWsOi3zbC4s4f65igETsclehXUstFIt/jBG
j687C4P4zVApBzI3lE/5xFxzGTS3Z6Ba0XLSQhlQqCZ7VwZglTf8S4UXNwfAWWd0k3jibbgT/wsh
ikeRx2/Dho8QMUWeH1XGTw5yYKnRdLkhepplbnXu3zcQd4zHVrTgjlSQ3vKRRcN+OMsOr+IPiSrl
PfYYgmZ8/RhtZU8pNiZQ1NQOX0e51aHJ94JpQNjqBpXJZbyilCJ+jLuO9mKSsH6jqIGaSQurWxPj
NIHZUvbCGzT7jv6wPomTS1SQrwfstH5neUmWY/aik77SHQX81pdaVJMfmOJdwsJWLay5Z8SRSxTc
zNssJGnjbFaUQaxhDeR3dO4ooxWQu0lARnKbtfGVTqX35azOFIEcgABN0I72hmau5omfpd2AJvkK
3JP1BlKUQG7Q7XbJkwvTklgJh5ZTHZEE4/92LoQ6VDoHPtrZdvAKBpEbtfyXUi8SyR9Kkd/qNQvv
xWrrcqD5vVQXRGweEhiC2u6kTDRPW5/DXHPmU7rUGKu+jb94kQy+pVg0EhjHXWrzshXpQ7r87OIq
SGVCUXIxpPT2vZJd2Z/Yn8GmoIEDHd0r1n684nU+rIWd/uviDhBuvGAIy5HHY4w79NKQHClCv0Th
sPZTzqGLrM9bhROd7Pb3IsTdasMHIvZR/zXeJn1tDhLg5q1FkxbSaFF7PUDhtYc+uQw3EUUWOxgw
Vb96A5eE8wqNs4EFDA2Byeqpw/S0S2Jdmb7LKoTzwjkRMz+DWTZ4l1SRv11YuCSolo6asnR8kjNR
C6hFe5bo7C6hq4Xjp2i7TCcGV5vAej+59kK3ZjUj0WqnTvmQK5zKMrU5+ilaUu85zVKaiIyvL8UM
QUwGafBxbxJ0rxTIUVQdfsMgNhOIgM8Vax+rrBnVsMBrHtgEqMOR1ZmFsqgQv0u5un5XNh6A9ZjL
zus+YjazeBN5GYPmokCqIuGByvUOHz7tjvhFUzRGkIbRY4UlnibPkHQOCWaMjF0iuU/aOY1mTmwZ
9XNkI1w8x4kco0M/ll7hFI8aHiZWusoGNB0Rjh7ZFGxkHRsZXYog1SKo01YGhDUuh+sc1QuQGpzY
UPu/iGVPGhJJMOfovEtMY4OkSfRkn1EO0e/rPNnX1/nab6w8+bjy0y8YV36W1J9jx+6i78C+LgrE
SqUF2CbZauqedzMV5yG4hWmI4gie86718zw3BG2h/mXK9pIjNdR2xW5EunpIJ4q0fXPXwElJygvg
Vs5ymPsXBsTDO0zQ3eLbicyg+tcgPe/lXFTXQn7sPguyjeSiFHYlk2GfJH596XfcSn5R0CQRU1+q
YPmbJrXDrp8s480ZEB8xnBgUO0s6a+HxHqvZGYu7eIyKmmoWo7SC/OEDnQUHbaBSg4jZHbhAfekP
FlbWVebbJGDx7T0XV1GIQqu47U0fIZFDPR+cAFTssu0SQp4MMECy3C6PNW6TJHnYiKBeXDaFj/6B
6h/ZY/HtacXdjXEqJnTl2D3j4l9OA8MRbbyzcUchd9H9uIwPfjMShQgL1p+oqJ5iQsEb/p22D4Cn
Fr6pvAcr+26Lksp8T53heIrftjleKuQ8cEAhlNa6z8Zn9PR3bod2CXoNyQx1i+vCDiXFNbjMxuuJ
YBy0wlIJU+fJC2aydVB0/3pcPFcXaEBi+QDDX/ZjKTeYMz4bFdFLZUw3O2OqH6EEXhNC5VCj0TEb
k2Ep4q2kMzigy7TNm95xRHdHKrrBno5ZDgHKpb/ShBwoDRHgiWAAzen7l6XHJ5LhLcXcK3EfsUFK
S6R2JCz8gBYf3B6AnuzCfoloJr8Yig8fcsMEZWE0gNJ0fcSPaIoZVJT0MT7EiveRH7BGEjBWb+k1
/OtU2V0aAxu/O/drxs1xU8RAYr/kMnZH2a50F+zqPTPMKgBBSBb6NHwqJ2J8XwpwWSKOP6x8roF5
2BkzZp5QpqCxS3JKs8JF9CBrSoecSMgX+by5k/ItuoQ+Wf57fOOi+BLsVnHP/3bWh2JQZKl/jRTK
gTsNhLchWD8xMt1hwIgVtbQMX2riOddZvO13A3+r1uO2+P2ej7jyiQaEk7VGUTjQhqOBchDc4w42
2eKwvDBkUZo7nIt5KsxSwEsgRaNZ7R4dDDRms/xLCIDmzUWDP7bzexgwjsBufvgL5Y+FFHFnV70r
gGwRCZFABFZkPdNCdHxunyzwyLGoPQNIl/Siha7ubjzXE+jvEbWdpMGKlvIuuRDo0NLKzIwYgs1f
+nvY82yw66n6DfC5aMCSKpEesII77mC+DmwWQuHnjQq3Uyo/jtEjmzH2iBRIPJCLFRME9vxlzdth
LN3tGpSiZe6r691b8sWkTxQTHPulCZ1SyVc0uXyNS7OzpN8WKqUcASFcCYch0U3txs8G/7bRIKco
ppU3UfQTdhn3RYcoY1d7NwIe93N4QtzKY/EqWFzeE2GtDmFqC6nK6hXd135HOOz6fKX6WJyAdG9b
evSweq+IGjwZ7QkaQKhydd+BWxeEL39gpGfppaVk9Ma2DJ+Lx/Oeo+xWPtHKuy3uvlvBLgjL4JIb
N65EhemUCm7f2PjolWcgHEzaj8YILYcsO21Za9B0b6Abuyjk0QvYD90lTMSMxSXuxNhyIHXwB3bK
lHe7bChIDPrWxwgn36hVkTGCRcQTp2Y43d0tQn2A9kN0lK03UpVjjttcrYPFqxIexnWZWDNz1mwE
rtPowXcpK3CsETI3FzRT5/JOXFjxgIqnYPKLGYxPloC2IjrYI6IoaNzoJ8IqX3GMGhNAk4aiJT8X
AeREegcpZndLIO3Hbo+P4VDANftN3Kgh9tYhFQWIVE4MsF/qiomS/6ArO3jT3rVwmpbCTwXTc7GK
K8OkPf78NAiVz902vkIgJN1XDDRlbRJsFSQNCjAkBZbeSqTzYH0hWerQzn+7uJJNE9C72GBf7mTF
pAF2R5DrBg0iDMNy3kGgxOj4/Y8bfc54ey2vyTMbgPcGfwGp3ON6WhZ7YUoqHkMzm7W2sug8WWjm
EHh/Rj84626j4L6xVJbu1dnhSAcqZupcR+14SBFNXA3qav+AqYU7Y5U6mLbAZiTBgm4UXCOUnAr6
/Z6CHf8q7vx1KhQL485oHLWt3SlMM8OuipDM0IcegeDcg9ZI6BT1dh9UOLcycX/UnPor9KpZ2qVo
5/qsGanhOphIWN5vxeVrp3TFkLTX0WkwZWpzFdwhtSh6emqUFt6MybVtqeRrBa9AuO9QFPWhmYS+
+8V5ESq/LQIfbaJ32EHmBF8FjyX8B8JXzDri9dyaPhbY9rpulH+3TtC7uoolU8UiatWXQd6NgkeZ
Vv0oO3vqeWKNUpgE7VhJP41UbSvmLiGndCFDxIQwwmck8hfpFICl3VxgZGJe6IQnP2SFHNBo6065
VBGoMDZms7KOSCJthb4aect1sXBBuy45/4iDPdYa7rNf1kxy4tas13SVP+/LKdQjlj5IrMzqTPZq
PWKzgKTk/1zmQFL+fOVH1tFZCdE+iXNwRUukTVVSHDoRrX11+qe7kxo9G2TrIG2VU0xLc0k/643c
Kb3GeHDmJVRjnVoVHhG8V6j89fGXETI6fQcCbbvSkhn4kQSCEwDiguOVoIKDv+/jd+UkxcA3FjuR
fmko+pyny7jirxSZySKS0PN8qN54KJeFF+sluFzupa2QDVSl2ZoUtI8ZUMXRZSI+OfvsrBTavgpl
1aTGant71RmMfbzwcSUAznFMLeF0ythTSNQc0BA3YsFAMAUHCs03/8yXa6D1uOX3xtNH195dmGXr
t7tCJGCJ4wxrzXGfWvpsb688U9h3ZGim/MVWRJIxoSV1XLCaxYX9Gq+aCn5EA6iTCSbvBMGxdQb7
LQr4I2WXloEaF5YJX5ks0GsCBqbC8fYsscemHaUWJPKP2lBy8coJJFC7zylZlLWJiOSsJXDb9eJa
SZQNpHotXCq2X8ZQB5Fl6JfM0G/m1K4isQChrdTsGVdZEbw0b6ZtM2R/V4iY1X+8a/Su6L+1XVwJ
OEm43dBJZLo0ji3fM2x0Ip1EPqXoYNAF3CLoI1W1ZyMRd2aXPNbiZ5gvTlH0bisiojUpN2xZzTla
uukqiRe+DnyRVxdjq3QMntZuKqUTooPYcCfs3+Fr62hXJagCA9rpWkv1vDqW95bwi0/bt8amgVtq
69TsACKZ+pKuLrZNq9L4kLB7zfI/r1ixw0qab/Gl6/MYcSkbxWAngBTXjUmYQToyy4gIthWruJyr
V7u5yOBHdqFpj2WJks9D6XKLFAwfxAHqGAYCbsxwp+shRExezYyYdCVju+Oo0HBlX+tiZXEv9L4M
90ZJN93JSKWSp8QwWaMonrX/sfHmdrKhYv+HrvPzvFQBHjmZSde4UJNO0sTljK3wr6W/mHlHyWHg
9yWNOWYh/xnZRsFwcXJrWo60mRyBnbEY4ppOnpS7zaryLPinkx++m1cR1jS9O7vd/ehB5njcq/mS
aDnE0sfu7QuZpH+7wqwAF/MgoMTn9N5bA6uYbu2L6WzSfuQsWdbVvhgUkReeEImfKrny7WS9DaGx
shJCRWjZctyEz9AfXN2k+oXV1h1kv3hO/+FxUrqfq7ph/uiQvHF/K+YXVqhCDd7jGakNpJ03Whr0
VVHv2caC22K3vCgWkkixUhHSSy8kuqIneF7eltTJWvVWDNgyCa7bzTh5rlQdkuHOC52yyXLiaFUB
LM7LKDwgyCWJ8qbRRYDqdMSmM4HZFTEvrYGVW8CyHVJAE/fh3zm4NfOu4FhsxH2LPsaODsGdTVmv
2tYAsObP5ugAW9UdyA/GtAxV9Sid8uOzYZE2noi7VNgzYUGxMvYufD4Jbka3mKUqFHYCe3fdUfKD
Pl3NK5RwYjZ3hOhPtFbI/sdKp/wfQyT0N9T4MJp/qkyIKngYgFrru4lDz/QK0Gk6AwDom87pZ3eh
kwre45N3M1WgRjcc3qj8tN45piplvvCAFRuj3T3t/hfa8n8ZWLXwXeBsw+YLaRF/CnE7WxqfrJhT
e9IePi2EV3UJIdDxy1qMhSgXXHuhFYw76JSFFScOWXNNkbVcBJVQvkOPwXxCbqelfLk9xeH6AefD
P3akZHtEd9znAWNqPl1jaaHjyOui0ifcoz5QImK9HFlfpCrtbYrSgcvMeFkN98LO8LSQ+UTbswt9
foc+miAgDxV0Usc1+Lhe/apKywUzuFc/CNUrsTW7VfzZ/zkkYRLArRjkmFNXBNLdymZbBGaQ1hn3
Vb2w3N/8V0l9It6rpB8+nqRBTMlVKekCd44dCpHSbcIOHjlNKI3cjB9dK0rJTX+LYsswFyZ63WVb
8keZaz3n0aJrKuKKEliXjql+VcGhcgRLsBFBnbqDnxH6MpNAbHdNrdCyEur/rM0sRVd6PV3sGixv
CD5x5aANvdAUI/JtYznd08uPYVeFCgVhb6xD6gljMbrXmsitGq1O4pZYw/Hr3YeQJ4Em1TLlpGcx
wCNAZZNVk7pLhNQmW9XSpQvZwaWJYwPwgD12AS0PY4S/ZZSWM8Gkb1qBdBNhZ7wsnY5hi9v+EX4x
8//qkF2OUOYhedRmNaIJ1NMV5i5hwijZgjEhHV6lP971PbcuipkCcggP0Rj/nO0Qk8ukxMcm1CmT
FehdgzmRIVe1bMTH9JdpxzHH8IZAiPfD+h/DUllDLeVTEZ0FbcZdpoiSC3gh6TMeA33p7pvaMc77
tk6oXO3Zbyj0SzdXdrByRCeFVyGYSAqmpNVavoxzO2DHpOuF2zqbBkIIJXsg0gIXRyof6ZOzMKAi
xbaexmtOFB+0iT7sXH+lSx5s6m8S3dzVYTd0ZNfW4EwYi3qvRB0oAnJ/BPdATQLp84P/7+nK0zZs
2s+gTgeyaS/foGuHKJkAwBrfFa/DB+TQjRlYKm5alvzJ+VZEKSc6LE3uu9ftJu5/fkAWR6+RyNeC
UwmEhHPCrD41CxodxFkNWdBMsTyYi+2OIq9RqVqj8qQX5b47TwzIH0kbqYUltmicnIjdn2ROuHN3
C3/YmIrD0DGcgxyB0s8ZeFh6qOFPGyI6WbAKM1PBlvGfz7IbEyWzjwS+rUlKA++fOYqNEJ5Ut/VM
rOev1jL1IhfpxOc5tN0ulJ8R4f9N616aeveytFZglw4CwdJ6kQyucbY7fzGq1Xt8azXjzwufZIMT
MHy32u3w1M6aK++gCinx5ZzANTf7aKIzKRg2xwh8TtaanChtxHuJy4N//j/gWoQdAB5+NLEgWsKs
SSN4aoEvuhlKZAR+s4ZJVnNtE2pIqvcxxjLcYzBAIwfIka7VGR4It/rnhoy2Ijdwt4Lh5CfSLUNO
7sxDWpThxDpl5NPK3oTQZbleHt7K3LZtFgQxIIjr8AsiWFSc/UdSNfNhF3MoymN59/QXCD9CMWDI
oe8MDI2xfF1U5oTtFRPSN1WQWidsskBErWCWbvfYrnCd9SllcYpJDffnJv/RK2cJIVP2G+OJMUAD
mzoRQZSVW3j7n6GmM/+yr+EHloTs3+VaKwVuYcYDnvWVoSnnKgK5IVT47FHHXt1G+MU5NN4hp9tx
cj+2qqSMzITNShor2TuazxZeft3z9699BkgsIWzadm2UnwtrGd43wu/m56b1XuViReUIxDJ6e+ro
T1nOiI2PPR+9F/ke0UwIg1L7oiupbnSp+OHpjLkK5ozs08qBIHDex8jyNzJJWc+n3I0P2hPJBOIa
dyBKLmIojTfP57inbl8P7bOtJpBb5ZH1/AXgMJO/Hqs3405HD1Oy4BCWog4lgrEgFchYdbsaHC/X
erYoUEZok8V5WQuyeSjeAAF6Iv7YV/G8XbICyXOHb9Wuap/UoBKPBvj3Ossz2t+9WZj2FAayF5oL
6SZjq8gioM9r50A7us62Z7Dmfr1buNFXBHtGsHMV9Mk+mFGbVeEwBCw3inemFaP7CYka4n94E9Zl
3aQS2wTGPgmopRjpRIabtb5i1f+sVIv8OeZMVMhkIuuYoCSPVPyr87DJrx+Lvvfz7z6/VrowuRLG
5DbgDZj+oB9yiouEGl5Ed7jxWbOQaLyX2fiTXaDeZcLc5JutFp4pNox0HlfWvOGW8Jpna0q4GeiB
kzlcW79UkHtd43X/Gwi3JWyLoXu1M/evmSRQijp0OkDav2LrM6+TXaTR7jkxJAutPOqOcmnR/OHz
SGri6GdmNHdsbzHJ0yuHVfo0w1eRV3iBc8otC3OPttK6KH56VK6wX+Gb8uNDHC0h+wMnxnP1G6zE
hV8okEGjQj4R0BB2sB1+BzuDOc4AM9eimAqx8ORRD9xA9JLwp92tbTNEAjpH8rIsYj0xMWPM4Kug
oq8exegLSNAJWnXcdTKTfYMfObIf0jeO5AE18mFnJckMVrmstLm8LNibP27Xvd1oNb0XT2xzLpcJ
t2+G6oxkCg2dqnk5vPbu4KA2WQfb8BKcvnzIWncbwwznFAuxNI/pfVup/Wg3nvsSZWt9botdaoHe
9NsTGkFMO74XFANrCVnGcazXP2v+Lbihb97+K3tM87g9+VKTt0VAuSd5hTY6TU/2shBHbQMQC+oc
9Rd5WeKqr5Sfwm7zNFa/U3KiCRu7U19MqjWw7sZMVTwy3lzTzUuSOHreMJAHqEUQB5jLPVK+v2lt
5xu4JJYGBUA24vfWTz25R/5QbRvNZ8p6hudlYbHCW2x9sHyH2WVccrXSh5Hh9Ng+aCul4XJSeC7y
vXTmdCPK0RPdQI7qAg8taN2ZlRCLmrM2sDMzn3vqf+bfpvS81vDFGyHAHGaacXVsdyXqsTMnZ4o8
d599dECR8HmY4RfDNwevKSm4UkDuv4BbJPJxFwvBb3yUz/wFTapdXtOIViY4VVIJcPAuTmu2ajNW
GXWZ8H9+QPJwHF/tNrg672/ZOelBPI8q8G7v4jIueiW0+ezD9gi2SKOt3Fah01Pk6bBVcjLewbom
+n4HAA71vjOT7x+IAYZX8+tpDUZ8FiSIR1FlRZHVJ7rZQCWi4xEVYUgvBEL4AqvN4g+0IUP7K88p
1OunDFJilGV51vo30KmJbBMeFyHRcg+Shdq5N4cWznmqeKFgyqST6nkfAniRgeflPO4UGdtX1ryw
IddtN6paSMEKKgu5/oGphQrpE5C+oBvIzqipjD4eCGyJCUC9XIQX72ZvYPz4IWGFtw0J+Fa57KME
zioGgIxeBZOTR4lx7FVWCLJgPEdbNEGuqs1ZgrRWQ9Fn8HmypUitxSinbjfQf89h3waPoVWD/N2o
FQfAJky3Pb9ugFqHBn5HEn5qYO3ReHcDU8eWI1jJXOYSyNkWgbQpGRuDNgd/WEiQ8g4On0KybZz1
RT8gr4NzUb0WVifHvzzFsRqXw+VKEn/I0nJ8HIRRIQpuoGXPNBSa4g2aqT6oI9XH5mC09fCLGHT0
YQAxsCmuwEcHuxr6zPh2dGKaQ5zulfTUGt3vmlWdl8xXqSb19yXzvI8KdCQEHRGIfC907cu4LQfP
2UQxXssghzDSsg7WE3v3YAR1cH7BmM1SpRJD9+mNmKzFrfpi1omuAvHgQkTToje6YZFrGt8zLAKn
1/I+Ieg7zn0ntflIwexrDvcMOX1G4fL4AgPihOp+CuAGb6R7D+vWiXk3Nm+YPMWcn+7dLHG1CLtH
NBEQVKZnS7AY8XK2VH81HwhuEfldZ8meYEQHlCV7uppN3IssvcR8ikwfAGc/tlXwvp71tsJZ4NHB
jlEUtbf6uY2UzEjGxn/OUMWFfwotJw45GJX+r8SRNQo9TybAHP9/a2TzENTiV9UCdblYpsYgGTwU
FEwSJfJbLZI/3D/cd+/Msih50sCIgf1fPyeOlX5KX4Hvvl7HC9UsNh2uRPDbwH6RDeVFRwojO27J
Vw5A2zZz3yLBE7Ht7npEQxIUEOZU2idIfz66VMrG0eW/zkSbdTUrBTKgH14SFoWoI0SuY1rConm0
EWFQhfzuahX6GemqDqmlEFC+ebHyDAYSvMEcyffGigW62S5jK+eeKwSYGs8ZltQdRKV4t7fiN5hx
7b6csC0vFIbskwS5rPcQZSbFHQGXGymU3VgPWx/kkaetMNOjM+4CPnhHGPTKjlWOFO1nFGlvjvB2
e8cyIuHbD6n2LIKjynlhEylW4nt8uaqKbKJuCD6ub1O7SOlGU3ixSrfnAuidLKVVjZW0VkPaMZER
fpVCChdBsK+qgWmdlWrbInLXmuQ2AeDkM3/nV7EeDuLA172OFqTkQHQ0m7EbaET0dL+l4JGr3/jN
GQ33aWS/J8UuQDgfwAKHFD7EngkWL+qeonVhVBiWDf+qD/VXD31Dx4hBNNEZ4XT0Zu+tulWIht6H
+Qso8BnTB2xEJXc8JQdr4kpIAKsEn+0W+iO8utaxMeSMAHbdxEl7eEcK1HV1T5M6Iwf12VYCYgfA
sGXfByYTxZQ09UdtBr/XHoYtmuKdhHG7x0YwdbjEZo4mht8uf5JTIVzTftyfljY/Y0SZ5huG5OZD
dZ7+9v5BQxX1hXSRyVITlMS1VKGleQuG3/nKbonb51aipmhIC8uw+B2ScQLogX+QtjQEd4W3DaOV
SxoReiPVKW49rtcWgUDIpELY5tnimcu+Jws74Z0qnP74bgk+htCwiEztHi7ZjUNtNxunYT790+jC
Xo2079ehL8hXrMqcnZTjQjCUTVahg1NFe/9Uh78zCNuzKN9KQJa9mBA9PdO9faDIuMsVAIbw36sK
sJi2vQ1tyXUSDzyvzIJVH3KtPJJnGdoi5A071rP8aJguYhG1u2Ar62VKcuTI0aXVbLpocGyGXPSg
940zuOA79YvQhNN0n6oxsmBWGcbSn4UIhxFFTAK7M5UJeJ9p1R+pkk9g9h1uJe6lgznwlp4RGN6F
FD2y8H3gscgjHKwIBwmwR+q4TDaJnStQwxMCty9zmxYTilGuk8Wxf2x8JpyB5avM0YdCmknxUtL+
TMcEPrtUZnukX71w2VzRlIVVuijt99hF7ub5AMLxwyITCRVuzxue8/pwYYazcR5NXB2bQmcPdubb
utBWIEF3ZjePWSSSC0aFFjb3KNgh3xzPDGRqXLBgGFttC/dyLLvNhvGhB+kpI6tMaCwXUYmb2qYi
Xt3fHqrSQZbd9ewUfERcmwywlTicj8JiH/Pbrz/Yebv6vnBQS4I7ZpZNR3JEaegRIcGSySrNvqpD
Y7s5clW8LzaTs5e9oWqIep2AqW8GDl+pHABCM3dMyb+fMSuPqAFN9jGDDn74XVeaQXtGZEMdyBYk
267cgtoEjOhA3HUSSDr7CdR7WCPBMukUEQ1NU4Dkx6yGK+9alWNyfoNe6vZ6WVFfxkXHZZrqll7N
ZbpCltBMey0UwfoDk75yKHiaQJ3BW/6H/axzwBYsbQOzYAe+10bpf0wdtfcUMdgSXsHeP43DXBNQ
rh6xlMFixzCNN9efr7MBjOPTIfudaPfgIRjzJD8zIMD9cz4jZ7kqAPeNv5tqMiuivkZGsdAVVf/P
ZmDcZ16BgdKj/f2lFdWGmcwEu/OSaIMBqpa8LdZefnmr/nlwKJGm888iILgvvgSoD7K2j3krUByz
ZCo0pKercmDhKT2TS5eqQIq+D5g/nVYjmJP/o96gNeU/4h7GUwpcy2IiuRJDBYyp+Pz87bvPhIYr
d+EyySjkm7FPun3i/i84PQJpfwwaAolFRUWybnRDbqIohJzsUSFryQusu4kuveEpaqlaRMj3d+cc
iV9JrjjcFn83VQScJrJ/You88NeK8hpurmDS0qK2xoN+JHUVHks0zwG7+3YzKDIZGR+GyAflnpiq
Prt8tvYJepvP5QJ0sZxcUN5wCxmlGux90SEuJwegGrUFoPddHWpmHiWcLWKEe6U3yfIpp4LY9vPR
Xhxn1LNZ2cSuorxpiaGacm5huvh3WPndMdu0QubZAO8GEyLLmDKmxBVD1Oqjq1mvZot3tsK0TaiV
OQQZI2MBQM8jnJ+JSx5h7kEKy3trszgDvdsKJAHLF9uo9vjjRGpBzARiL0B/ZMWj5A8cvkFRYjaz
a6Xs2za1Y0dKxDFAmEkZ/ZXMsrYhKpP0ntzr2jW6hHiH/vJnA3VPCE1UXGrGstaP6EfhkYeMBI5Z
bg3WT4YYZU1cEYgfnlkKjGAD+WyRoSzhAUtAuESrmEmRTsaTErRWQ6aFTLst+B4TG1NZaHuPnrVK
NbzGuH4qD6B48uVOwnBdBPGeLrJnEOoXuzc2TMbjBL65oP4LC0nvpK5XoALeTJpfB0Cei4F44Kl0
l5OavDeh71kXhf6i9oOzm4iZfKWcDSIeY5eRk3T9pMRbvbRvc6/Yg0q5/Hc7MUBpJpm0Fjuaf+o6
nQx6k+cXes16yAQPuhVHS/sDWHS3PsSqeMqfoFqLLNWNNyw8jTym/g1CxZVdULcEEYMuk2BAPKIF
Gr0Xw+1/aWRTRbWI9dizmBeozYEgNTSU0sDDOKnNH0Q/dVqw83Bzk9QXI3XOzDJ9B9/UppGgC2hN
cXkUGCYShXRQVmMPab0l+VCtsdFPJi0sVronAsn9Rz8rQwA5mDEgwhRgLcTAReFnZ8/gF88nY9hb
6jp8xEJNLe4b0UiEzLwN8GH8NFOJhVyMN0zzREB9dvqzsaXZKzJyj/i10VwXZsTFWmIIrCnWUgua
1meuAG85E3lQUplQkzyyVKZ+9LsneKUFrhPpBcupAYHpi3tAPWI4vXbaxyST80Pk/g0Aniig8LiC
C6NFXRvt0JhWXlHR+JvYsBYGj6KTRM3/Y1hcBXdfClNfhzRQYbEqMJmh/VTo42n1cerofzi27OD1
xLbQQq6+ejDujbyeWDbUin1F/AFeup1cOERzwGIZSMgd8f/wsaFKjC8fwvPfDQ+FH2ktWFeKv7Gq
iT+VxuSCsrpav5mwci6xrEHXHXOxRBYv+6gdHI8sfeKhIW+Teco382D0SSA+eK9hEac7TfUkHYdh
WBmitrqu0qidqMI1ie1f9BpFWDFykOhitpBsLOX5Degl3IvwVKAeA1weVfzVp8zuumPR9ONcjmlA
3W7A8MetOKUYBJLcqy2/SBluJXe+7K7tpsIOq3oD5c4RRuylan9IkYWdO+U657es918k0BE4Azz0
eZSw1qkUG94kLTDAPUp4FpvNnmQyp7ltt3bIRfSQyyjxkFCCVR22tpok3J0wY8HakMv/Ah2nRaMQ
jbBeihCvFZTGnIdb2ElrbcmFP1qBlm2ywDTcPBR+EhBVwMUsHTazuMDOKbi+Y7Ba0PHFX/Z53c6e
a4ujPrpHsC/z2gEaappxsvDuUemevjMlAgefsPZQV4WP8m6pxVTS+WFHtgUURIOv1joUEc29LwR0
3wKABSjmWJHAU4JfB+AFfKfy1yIKO01YhkObJxQ/7vkZQUl3J/riajwGyZDb4LRN96/t5+YnS6fE
CtHXSfKsZmkUq0ucey6yBqKBHrG9VXgASH4kO7v9zBNttyUW1hC02IwZkxF4+xvCKs1m1GaM1uSP
PIBL/AMNFhmuxJF0AzmDBO/W0R1buHin+chJIbhbLzKO5nZA3CWcrexerPngS1z71sSa2VFEu9Zl
IVh1ZRsIpZyQB/ZndzA3C534dB2n8kKaAoZVbj/AVLhDuHa2aghdtabOEdR9P78mfpXfT3dSJTnq
ZtQ2e28tXtrNaGBhvitijWnRNnW9pgyY2uk4B3L6l4Llv17imQix8uwWALXpbU9uU+6QrMrp0NUq
LMIRdwPz3zT8Cx9Q37Kl/81OD6m7ktdakommze4OTbZkK6RLKQm2ttuLxabgzzizeYDPmcSG4BkY
KFvSuFPLgh18fZIKOFqGJtSi3HuEPU2Hjz25ySJy3a61foBsySHLZ7wHv4IBRSZUoA72OezI3PDT
AaN/4V/KYuxbJCIiqKNF7IroWYVLrCS0R7k79m25NQ7/yOAZ4nzP6SyObUH9v58YaZ7hWeKC4+3y
a986PIcH0H414Kshyne6Zp2wNVfcB1XVBQpvCkzpyj5qywJuII1W1Q3VmWSRNtc+xKs1yWnS2s+P
lNqvCBPZsmr6onpVoYAVGxL/yo/b3AOR6TRyFG9c++uswNxn5w10Pv/hJ/35exLtCab8PKUETnsE
O7t4U70tHdihUeU/svcyQWku++3265fajB9O0AumRZhe62Lu8gByJyniwX4retsVMKO9cCH5csnM
nz0bjheoOWreVV5ILqO+eMtb7CdXenBlWMIv7UYEVVITbmf0uUwmWSeFm0oSC36/XfVm52rqvItT
sKwY/4JT/lCGblXson03L+VZrx3Xt+dISy5BfwKfhIJajVCvqKqaCePaSBH1D3mCxj2Bn4K29Ejy
ZAwUv2Lg1l4P53MNndc71GEn8ddbDxp18825GPMC3AoAGN7psQPQJEYfovmYvsVZ62EP+GKr4aQI
PzxFXNZu2k2/ihzdBwd5QFh+YRdCww3Hhsqd4TlBTHRlvDOUcAwL24Ha6gSQ3emVkbsI/30EKnpT
Kuemi4JSEvUqA2CSuADdy76YaveFKVDEuQ/ZK9qFAcHZQMcte9jkH7dqQ5+UhFBMmSUwyDj+8afb
KA/+m29GhuUwgy/GCXt0s0mmWTKBt0QG1oCTUiT7g24xc/ENLrzaoQDPlHSDoecTkQopgLwSxs7+
MLG9x7g8I9V5VP/k2k2VT+jnwKLAPTGLfzndtOc+3Kx3joqoKXulz6h2cOwpPfR08KgzAPHHIUOY
UQ9IOambjhVAq82CmjlH7W3PWWw4O38V8LpZ4My6L2DcU1753weDsNODeEMTVQ6+7rpFlRGwpzUF
SHBLZY2WbnSSaG8kW4ZdjFpgDVWtJGvRgM4rBa6Xxe4yyQJypxJhWg2M4KyRGEzwxvNFmoJnEppU
5QNCpQ3PNoLiqg3LYsMf6P0Y3U5FePk4YoxvBmL/3jU6UnJPMmdSppXhM48V3C+wI5iy7pqnD+pm
SKaUZN6OGZq0WbMlxrObcnecMWFePt7wKKTgalT+dPGNFVs2QSx+kaW52Cjc+oQPQtDKauSGvCa/
jkJ457CilclkTm1VyUyQn1XfbOK5LDUkyI2uCB8A/965OVv3ueYW9EXxVSgfwSKqCFjQpE81i2MU
kt/PyyXFlbI2uqQ7tLdl/GTLfa0RAZ9rfWJOZB1lN7YXDI33hwmt1/LZVd9lkCcDcXctCf9CRcAT
6R/Tb7cecFFnn8O2eCpR4JU9dTvNoGjYZWwAcdiuKQ4nj0zEiaGPjwtynwIQ9JVt5GC88odgLWqh
mS/psbE96p4ZJJjLpTAAnyvujFYIdl+dXViXrTbzGBMu3/710T7xaZ9QKSfswHa3k3i9DLxrECMQ
WMBjc/0ofXCjZSr2196IUmsDMMGxnMt5v1R9VS5AAHVjH24VJEd1UkE2FeP6QzZAJuyT3ceD8G5A
ygY3hg5s5BnDyeGlum4QTezMDaQGuiW4ZCef/Pk1F1Anh+oKNHWfIytNGA9sCgWD31lq7b5A8Bzg
NlUm69W5ebe2mIu0qzNgd3pf3wSVZ5vygfJss74W6EGX7shj/9MYK5Ime403nDxI7RidQ9V8+sjB
axdHGQ+XiOUI3S74nqyg08XNMU8Ekfdd0EezmbxOMA0TZVQsTYmoY45VVhYmqD7KgH6Aa/yfqFI3
UB4GmATT0/Uss3QN0w1SMckDOLC8MSlxCOf//M7GlsBQlqSdoNBlJk/dth9qq0svh+1j8OdFeAiV
jWwAGIMNrbNvx3SSL8bWt3ErSu8XbLRkXZRO5+zQu2tDLYjWZkmsq23Y3DmhwCc99oZ4eqm7ijr3
dOGo+1ZfwaEpDLgm16hh7lgb+iWSbfKOuy4iaQYxhtNVOWo0yE7R06BI5qQYPPa6isGE58BsKqvc
b6zfLlePf+KKXnCEGVxY03B7sHAmKjgP+lUBBDgfgspNjoRSG/jjl+Az9bD8R6og5mpZXJ0nMzem
fORxzFKCtI4L/XZiksnw9XjEvJTealw6XfgYBWG8Ti4tnaoc/Bw1HOROUuD0c2l7rA8mpAhPnt6L
5MbY/Zr4QmamPlPQzVEHncwmOAs9oiq9OD4FFRVuwJ77/hNn3pGIIZTpGTJcpbYdu6mnvgUIc9B1
asxJclC+AB8gME0FAs7PyazgMLaZsu2aKPw93E+u6akDeeL5Dz5JcF7wAW8UEMSvkNaRmT54uhzN
tUruLWj2L3yXE92zFtxe0cSX6Tt+vR1epgCaVkkLb7bBAdVbE4R7zDN3WhaSRr9dlleT1grn38SS
qdq9PncydsxFmvxPjaVRpHvh912qpnMwkfCsSUzd+dw4WbsHnzs2WIZEy5TiMGjnVdnDPT0OfkwP
gO2Izh+27r864Uuc5PBn96UWmSg9bnHyhq4dM/nQHy671mBUXJhMo5N8+s5oGf7INjgcyHKtAvHq
TXv7xcqtDhzBaReCbv0go2CrzKBhMEl7GpFtQ5f5dc3Ki5ElS1BU1DKWs/qyr91C96C6fwkanMBg
b9bKs9ETu6j1vSW7u2300Jjm++6p1viy7q+XDCEhNsYQHafQbzXyN1iZB+BxApSGjT0UXldIANB1
pZzkjDCvKXAv5QywL7BXxw5cpayoYdYZVhtkj0WpM8RHIPbv00nfHtuScNgCIex6Tc+4GfLhnsCZ
Pgrm4Nbu3hQtOhUbKGxfPiPbWIarjE1HZo3Z5fB47ZSPI0r6mEkHm5KISzCcU4qDqEg/5FLBI+tF
DFItKnCYn/w5eE8bZZzpPaWBPWPvJmj5zWn2gjFUcKTTBQjFSPauEVzgB6/W5YSWlBnKVR65ZO8I
nDMZ9Paf5PNsACL/iZ98G3tViv6J5bN44vPF2K7oFv3CuULvtnYKJUIKiLcSAQSplQf/jv45Z1uB
4ZePMyHb8kU2ks5piFWmEzt/mkKrqdKia+jiq1fHPsJOPTmV2wPqSJIYcWh2F3IaXULEiDFCYYdr
qH8OWItIkcIolerCtbJ+TVag69V5vuo+1/3eAPt/CBOXSyTMh/IQ1uMnTjsRDEk9WSQRsf4Fzcbl
IMVmnssqddzauHSOIp7se/afVlb+c+dIAqitBR4ul61Pfzb5LamU4Yrp+HRGqPZbJa8qQnWxM2q4
hbntCRMZ8jDyPOTSmMn8LRRbdBeNDjY7LrVE16ikF+xpiezoPpPSql1PWoe05hL+9YEvyh9levKg
lD6YHCpR2qS9OtP8uv1vrXf25jQba/PLvIK+ucEcuqFc7qc0GzfG0N+/EaHFmiU9Kzs6J7Lnlo85
m0epmf+ooc2pSAeEes/c5sD8ZrhUzqTXD/CHF81vYKm+omcSwGPGKeP7Lp+l2kh2tjTgi67dRE9i
UjEGStgi/5FUfrojv15XYhDx8Ofh6WYWjnyQ/d7mEFrXuZfJsqMxHTUlNt63wF44ppz+fUaiLiW3
BTop7cyJsx51twgB8mppt5sY6ZRFM889jiT/eFXJRErH8o0C1Jkfk0A6MamrXvGXwdTOzPJhGnrC
aCFmAfdGai7uj13FmPu0yCrPEAMYCGrB25zicAID39y1QLLsQ6l6HWrBvkqVwv7+qbb6s4VztYll
sUxdDlZSXoewJ+VH4OcIJDhd9gm2GpoCUxyx1vkY6elnhVBk+5FQ8QFR9i+byjl3NTNq4AGRKad5
YI/qO96GnQ4ktNlNUF9SyqsBY3b8mq24w+xD7Zd0mlNtPZQJJ4t/prd5KQVmkcXwRGjI4Gk29LX9
gEpDtR39eX71JJL+Y17QI8owE3cx/0zrrUTIeR6Q/ugDfvonRSVSwB8PGZXDIJBAsfrfhVpU8pnF
y3cq1qLXhHBymaGtgxDJFieNFSTeYDunwGd1tkrwBwACtHA6dqdaoXFlnM3u3DVJQ9tN9HGr59xX
gI/tgfySogTCfk6R5zYChhrUCnb4th5yRT0Kcp4n67ZqzyFc5+5hVQ998ltQoyHgsrSbqmT0inPY
/3k9zqwGoELy4Bvx+qlvFdWCDUBvGvo6LW6oI64a3NTfHdxA1IE8jhCyGcjdpNERGjC36zer4AMH
QcB/turNVidTMEDfvDlEl/1RNGyT2MRec8bZXMp3r1oFD63u06PsDOnRQFoPncMEgui9zIDDJ7HN
1abfP4qkPxNi8/B9jwiGsvqmWf+YFOcttQqmOlNVfVGclREZTDzkdMYHs68X756gG7ZT8z3dB5z2
f2TK41rop0T7dPfPBQvViqlPruP0QIqZ6QTnmo1wbVp3pzJ6ahpl9E+mAI0uCaN4pz1jwkrxvFxw
UrUjaJrU5caSNH4QFnhqfOo9R1yjKxxB8F6rO6K6Iw09hCtRvvtlcZA/JsvWhvkSnKjpM5kbwPVP
Bfql1A/YPor+yFNrSydfwfZnaN+eiNcGOTmcy3s3W8vPQUG08YL5yoQdKH5+tELPm/r/77pA87uR
7HjmKNh9lCL6wm2F9b9jb+dlitDLArcVBwse7/DoVKFfXy7PPNJ2CvgyrW46rSGGOvTS4YBPW/tP
wBjaMQyvXZJs8k1pWiTkRCFYix5GhsHgofIPlRHDdWj+7QcF4udVUvLWoRLg9LVkO+FaAJOdGsxV
T4at8dacNnwnLeCw4mMU0AgghwRE6Rx5NgfXDAXX/czUnp3oLCIfoN5+TBurQXZCF/pk1xH6uYDT
JK4Xt0X65PnDlAIZ5/YD4q8PE+EfFE4p2PTS6EaqOf2ayQQtyB6VjsD7fBvN/O+amo32P5Fx6KbM
E673rRTUbsse3Dssx3Jn0g/3LYnQ0UYyIwBwKMjM6aS9k1DbefhlErJxTALjH5KO7H/1BHDUPbao
A0XlU0eC2MfbLRueJLBvsTaGS11mvTvxTA/8e0e9gd1+Mn3YphMR8CycUlq9v4tVK9mkr7XckGr/
UHZU+kj8TFkoIgaa+CJxaoDdRFc/pkMsdcYcplt5LWWWt+7Q/xlruafYYpP52qX9lM7+tCybIXDw
NC08iAdnJWr7aqJ2/hMxlwSsGTj10TyEqTyKocVgFNa62U1/M268pJlrzIiODV+oioh/3HeRK7km
YxCGjhZ9J09S2vapZIPu5+iWgGTyIadWWiIt59tyYrrw2F7nYRa8oI/2QP7kGXLiKediniUrqdXT
IsU9gnVzl7WT9xk8LMJU6w28cO0DZ1dIIHTnDEj/SHKwxf5bNdpq1rVaSVhw0USeqHbJ3ZREdW2t
uPWWPyHYRIl35W46KjL8A3MJfRuoIauxnvA1TE6Dc4HDRKZy4giFlFm+uGQNmQ+NPsum5e9bmB+e
ePr9r8342NF02pi3y4aenME2mbCADT+277RYhwF9JjMFoD2eQaIycr7kWxkXg2o3QrU8dUZMCrE6
pEJmZ0r/dcG7uuRqghJjvytGwqz193WzwNuYKXkujcbv+amnHJkFsiNn8Mnt3LYAJrU/bwey81rd
ax1szFW1DUm7ezdrInIXW3spnBeWvkzr7FXe/1uyeLz5+qmY+SNZIUQc4n94h8Pl1UWjwh6NEirs
Q7ReY23uX/NgcT0XcuvOAA5EyoCdrDiBnz9Nwi7xpFeSU45NZfwpZZF0LaHdpPeB74af1NBl2wyk
9Bx5F+eC60vJCecsuEjHQk+mZ5E6OHN4nzUXHSIwRHBxYzu8H7/nWqObwXOV3mcvQDSweBYGDUHF
e+iYc3K97iaASvZxVj78rjhinXmIWWrdUO0T06hzVARudbIE6tqQZmO89IYTdPSLw2/S18gyyCD6
QfnD5JW9ZjfX0wCCGr3jQWgPPDmb/bOXXwV+snStO8bRPZY2/FIk6uisyHzg5KMTEvWKuHFTl5tQ
AZAkFuNCH523ymL4cGlTkySEsx7FxgwYBb5YYVDf+D4ysjqe3aDXWexdWp0p6gHqmnKFrQ/guYI4
p0SCqmyHcUYjDcuMvskU/6ZHN4XTBDgZXsmpu8V9aMDOQbKpTtqELcCDI3Mf59Qwm+2t0/2T/6VC
Mup//BpAar1E/4U5YHyATaQhCnpubHGv1GF4bL8uaxihFuO4s4dNPvtC9REiVbBCe0e1Lcpt1N13
8otlM3DzaxzE8daPWaLRqUAga8yL3VIk/wGLyVGVm+PrESH74RBoiOaGlXq7HjH0GUFkvS0MdLuW
y8uLEWb6AnDsaW0SeJcyoz0UUCBgE19QyvJOVrE4Wix16zXy8TZLbzvjeYnl/8qSBjjusgCmDlXo
qRBTNzTa2RVPdOTdGdPYWVe8LTK6ByaVuOUjWKo+/Fbc5nwmLvsk13NjECUQZdiaSb6bYnVsa/tn
RBKsos+t823pfKj88w9QiHCaOtRo1ufekGh2N9vGsFyrITd0cnxQ4+BR/KpfX7r3DmCfeawS1MfG
NRradd3hL8oN8QG/DsAOHiRMbzgLtIheTTfmoZqSXob7oAXxCa5H/En5AnJkSqdsjJ2Kw+8BDOEm
siY3yC9cox1UFdg9GJMP05hb6uZcUNTNksXxWtlAsAt0Hq/99pKP6o1ydwXkwU638+kOey3uVewn
u5e9LeKCmlE3e9VCziB5Uom+KE6n5REV4QORg5GdsuFU0B58K3VSc8h98IEto3+cZpcJ8NXvgwmf
PYEcG1s7r7wOPvhHZr1rpFFaPxvdlBZCm+80MkwsSTMxcPfRv4BQtvL9YTnMnFTm8KMr2Hwx8IIJ
n/aRz0qN/Rt8UWlbSb8pZ08TWOYZar0v+/HgqSCtGWED0jrFmig2ffPCSbugj61mQ863H5Eft+1Q
17QEzBWmVSyLscced13Ul+bNiPAox1GNTlFMN9FGJ8MYX60NECC2aN2lPTBpRCymjn4trVsDigzK
zeu2XvL7+9liYXXUWzf/HnQ9cOb4tCiC3s24UW8fRYi/OJ6h3GuHQga16xSuHpuGSXyWVXvX/LSP
4FKGrVl+kukXJUME/HCGErDxRlmSuORvyKbcDENc4hDySX7c2GwF6qswnTdlieC2CO5xjiVmMMw8
3UsMtmO153ZJC68xXOm8yoxa9vjuEBcLZmYOWoUj6vFljx3SnqG05NkG9gz7YDVFcHVhOEhkaUiH
NgTb0IsFTmwzl4NX7iNrbgV1ZiSqPU3YDEiIXB9fQ8nXRaJRKDRYeCZbROam0Vk1ob3cxrj89EAA
S6/FdnNy8ZV/OCsHKBbuW/cmZGJheGOM9gbJvbz+U1MsA7wX532Vh55CXrgS0eEbTsHS61/gS4ds
iJSgrsCMhqC5dveBkr8EJOBoeVZtg8mmT31P7wv2m243zexz/8b56BL2h9ugNSPfFLET2KNU7DYX
NGKSZho521ArU17NykPTUnhJb8LxsaN0TbyApqHW/1M556rkNtaz66cBfH0PTLXRGjVNjzeSsKmm
SIBUaWKO1Oo0FemIs1sz9zrAKkjfMQA+QjIF9XDQPfBGz8CnjAf9RlJZ/2ddsXAqMPG/SMqtx08w
6Aa71nTOK8L2/sf03Oi/WrRh+8ZfgcXkPT7Ajbeg3vFikVS4dc24MlDG6nUPVW2zx0/rQ9ep+pzw
kbF2YMXKkymKss/VZuRlvNY4mH6tLig/PbQpzAWAnd1SDZLaMKxr7tL0LuLRofuyNKCoiRAN4Q32
O6v/iGXLi1GDobDzcS8NypgayvNrqpjTtKeU8iYg9CU/LmoObVmQf+v/hiDu5kc5tNlqG5TP07aN
rOaxcg+zgUI1mQEagDs4TFOdbF7py+FvCXSqX/5tzk9S/NLUk3MJlP5GjnlK50IW0vcpWjJ4B7hs
6/CBKi259Q0dsrjv9YMLJ33u3DG0jmj1lhPcgKJXphTwn/AErQ37zstkaSROKA3VUmxkS5qxRPME
oTQlZD9LFHYdnlYLrlGPD2beMHpDAExLt71v9DDD43l8GbU1SpYthpf7+XA5RDBOBZzUXcJvU9K1
pZafQUu9UJ2g67qL4XPVXW3TxQEgMKr4Lv1QsZbGWWVg5D4FHEa+2slTeKxbndLaFa0OBLfVM68+
NuTLcmeFNFdNTwk6fViqkYBnPyE74vidE03lZpIYgiZTRMXX2E2QRYSncZZA8/qhsvxjP+4A4cwv
c2qcOhUJHakXEOfu0fPe9IHPWwhkrKPDNOl/6lMpYu7/amjH1iSiSOD46wGE5F39WoxBopGkboL3
h9J/oNUgbCBntyplc4OegJMh2DlIlUcqhfWfgXXafxpD4CFlKO9mj7k9M7aZkHKmeeEJDcUQ4GWd
pZdvuFzpg3u8AK3lEM2YQG2dmNfoOx/vopteSOwoAEMqeaLMtfq/kjVB/wAl5JIb6F3FbeeSc1vc
48VOYQuAl3U0eWNgMWhAPo/FTkBS5lqyD9Fg3hP+ex2GwbrtSa6tPZcXfr7gAFFGy6jX6z8Vu9aU
9HJ7jMkBTpC99WqYbHkD7OwbSNhvmCSJ0VBCL95Vrx2Re/+ImkAC42zbflmfBksw6Mz8GVp1XlzX
yImvLk7BoQYwnfrE4eR6eXaVItRmD7z3jpq+VjW4zjnEK0km4Lk6yWjPQroLVnodWFR0H+ocxT07
bBFO19l6GJuiEndd3TmQvLO6SZOrSUtlrUpYXC4e0G7bFDYiSqd5d+8RsAZ+vdL1jcluZM7ogcjR
73vYpvbPat84GQJxsgdLLT3NVwF7EovDSY0iXP7bRM3IMA5KbWQaOoVOzLbw4MOgE6YcF6sNxWCC
9a7K4CPnBkyb4dtVyoFyU+4jW2/MNUXGqczgDU/sMj0DlqvTyyahk3EBPInZEAObAE2K7oqbTfv/
+yY0xwXl6y5/Gh7Q4Nk1LEGW4InT4Sqf55JLESRDV/du5qDP+G+riR+IyOyvhuD9/GEre+BkBY3f
Ij/egC8uBG0afsFJhpe3brsxD7zURY+7QyTC7UDUaG2R4J1q0EtsR8DFOJBFK7nxI2RGxhOygZ/Q
SLhqX0npmVBYNMQ87yT3yh1pQ8yy+BmpCZlfP9XbMFDVr4pc+Fz/JNcxgsvZ34IBs0mlVhWI6qdx
Ag95kQMBvPimPYYBEsh5EQHoeL2E32h2+cbCAYS2RBC3bGc+ut2iBC1xvp/I4QmAav7PzPlD3OmW
kjuFKyqmztgaa4tlVihUQZRFC9nxmkobNK2O9ezn10eYve/dJcFR99AhYIxykrXFOt7JAt96Xw9S
SwZfA+2Y5z/ZR9nUYqDR0lr92z7qm9seNtCIUfjlS8Gn4Cow7xa3D0EbXlhIN9hE+l3gS4g6stFi
t90/PIeUoEuva2pRlqFN+p6PScTtJewplYL9UgK0SbRblCAY8Ighj0vUroDqFmMjxgkpz12RP3YS
fbq0eFjgLyJgu9zK0RZ8kxDDCtHxnN9oo6ICPow63kNrAUUnzYLnlYGG4R2cNTNNICr9AjFaaArr
vqoXeFa0rtiHDIsr5X6Rm8eAoIE4MzchSWnVf7gWfknAL7MWU4aF8uSROmuSEeh+NI0XsuQcEfgi
KFiDoobaqF1NzY+JUCIjaFI9rmz+PP1kVZzL94Sjv+cztRTIGWQTjnmGYsAZSEcdMi4aW9Ztkgr4
3RjgovHpyvLjk6NFQ9bYr5EwN5hN5MTksOuxPYHETYQmiB5bxQ1zc1kyVmVm9A/UpahCq4jDSIs3
8gaM8EiTmKcgdK2REZ4B4RqYozut9yQ0AUKKnw/U4XaFP85tHBm7JFZzaiRAKhdnumCdLHlo6cnJ
hwBfTtCToFjFvZmootWarze4qn9ygeJvP3iygbr+FzbjrZ4r2OkZfR521EU2fcdnND+Sbyh4jvAK
05vGWDp3CheAjbUasU++6ug3JYttw0hP+kHydKdLM5CtLBh/dOt0Ba/ikhZRE+VPbP8ycG38auCK
UwCD+6m1Nd6VWFKROdOP5LAv6uOD2w++5ltUKoe5YsA1Mtb/m3FmVzpkvfHUECiha13EJXEAd2w2
BmcNFDrfs0ZwNKUcq2x0eeD3N9AQRgwUwyhTEJK6t4xM9rmLOvY0Ocgws+ngvAGK3R8F2NPd445s
zM0No3kNLOT/G0+nmzSPQCq5T/YPOdW7LjImKkoGvFgZUHJwxzLD2b5Pj5mUqhnVJrM7yO2aIQHk
ArdmGx76XzvC7QpDxurtkdvZ5o6t8jiTOfcf728tQ1Pf2iQzdN+ApqyVS3cVBfO4DcOe4waoFKml
pwe0NM+r5yoBnoVmWt8sO0sSbqN+zZpCfQ89ndRamFEThxfMLT6Ph1k/JLhCMeFDERwyhbs12ORI
jY84emaTkpliUyxZWky9ED8P7bKOQ9v8WlSwMzWx+y26vyYv5Hp1HcvQuCeK+95ZjuyaFVzgmP7h
7ztrl7/AHbsUOvGJkpHCYNUk01fR8OWSB0Jjlnhen4zuyFdNRZ+sbwqJ13b1XKbFlfmZOmWt8GIZ
Nk9K4GGLQbTlde6Guso5NE223+LqldKBHsnYN/xL0SIcl8B+k6Wfq3ACNtTERCj21u+aQakSzLOd
bjisgi7PG/Qc5+lsRhvLP8A9Stv+mvnhWU4yKIcBc96ATLc8i2G+Zc1cKokFDZHknhYX3PMyebiT
xqM69EfKEcypzIUv+uY87x6Cvoep29RrPrJQL6GdjwTUdCStUihaHS0QrkfUqcn5XxUIPWMesglr
6gfB0Bi8UKJaMIscJDr+3v2EyZP2zuKsTD2i7+DiTz5+JHGtcLvRW4iTg+KqHn68hHHXXpyEbjQS
6E7C7NHh2UKf9q6kiWe1Kf4iBbqp7vPy1v7sYDWYr0lO9OJV28Y+XWQcUIVikISwlZhK/8axG0sI
V4LVsTb95np1rDLqCLds3PY5EmnSu1ZWQroyjuI0sF6hvSn0YNRelEM5dYRUZwVMB/b6thX9nJNu
oxdf/w8FJ4eZ//78uC2UIDrOyk4yXsQVmbnlRXRQlZuC2RXosrUk4ITMK+A56jSzn2t1N7SH9eos
GE+edptd10T7Fp5a7r886xDJSM8/y+qMbrnripbHIeqqtoBM5z3sgLpdhY6uXi8Q97wbpNHzM2VV
pYbOdmAMNrHMxL98E8hkxSCWz7KjPSYgdnXxGgiR84XKKHIOC4Nl+mLRsIiYqwO5WdZY/cMx7qst
KYeH19DjagpPhBY+awS+mXrF44fI76ALhpE9RFIGbvYTT+nudw6Jp53P36yOWi7YN40ApJjVHhXQ
UeqBcN5rYLPRL0Ma4rQt+397O+9RYiNH3D2k8XXw/D8JFDgOu3t3HYaPie94xCvgXyP0tqN1tmK5
qJpzS7ICaPXrdZaRL5bga25EvoIsLY07D3D/c1yUOLHYjSwbBVjP+9VVNWpDGBE/Sd22LS3OR0gB
VWWj+K4qlh2uwYGQXXGQHoBcVE+EBBaydUTTNp9pdgrUTNySTO3t/3kthHGgi/pWMs3IkwmALaiJ
z4pS6/AA3lMXb6Xd280SGa/VeWUqXGjsoQiCnaq8tj9Ih+uY5sfuQ2XUn7OQ7Y+esRw/ZvGvRMbz
0FxVJNlahcoo0fdO8JQcXZH6NwYkeqXI3p84FPCnvHEELa7pu2InKgZ1gY+9fIydw35XXMAYjizu
qPzIPTTS3Y4MzEu5P9aC3Sc6hVhdV01mvarBoheREjZfV83aIx6sNGCn/7JDPrul/G+m+PWUd5b9
uTR+FK3PLdSfrbCBtWOwYETyHy+vtWoh70b1r1n/oKXLHbV5O1cZWNGGxOhnUDLPDuuJtzMjwzCy
Qj8Fj6DhK2zfZ6DZv6nxSlIOLD+O3ElIhTcRWOrsnsPPCHYHq65cLYR3jM8Thpj1ub9nJ6XbdB1x
16jqJnPMBn5H0r8kRR5wUYWNaU+49n7+flsWy1nrupGcp2tJ/eltPdMAIgjjSaXK0nRkvkb1IyqV
ITtyyk0HXpVDJREZh6ON7q+FBq25HETCx5BA2e2C3EBxiJptE+/kGnc4r/oLJRz0UGchYGaJZqYI
xJiwUGfoNgPSAW/xMw8cSZ3VpPDHFZUhEGeupHeBkxBL6OSIjeOvCfegTgC6aziLUjNZPHtkP9Js
29ODrcPAHElFs8VpxDo5I6NpeJ491pAANuqUAC9Y+WfhJxLXNzxEkBFCLw9o6F+pUvLKB4y7JNtS
jDbU4dGCBPnsNWefHhG9ENDaEEBUO9CTX2yA7NuC9g1dwv78soCxtFrbO8C7x6/3dyTsLUkalRIc
5+6LLtMotY1lnw4lR6UvW5LSGnZ0vYwAMqyO8aRL7BvKdV49Xz7hk0p+XW5nuRtVk0LTk5dMYxmp
58X7kN9LzW1bRK0n+xJrnBhzpmWxd4fJYzywzmc8rL8l9gXbraXnQ1saBzHUENmh3yRYF+5V2V2B
delWMiTXggCfNG87zWuLcZ1WoQ/A9iBzteEN41vQv6607xhTqQsNQqGp1NZeMcdBxq701zoSsAVO
+t5irwGzDGuKTzrAWDbNHoS+ThNUqfuqpdgJnRvdpcIBKSjMUU0Xu/pN3lVCwxUseoyTlPqMCSZx
1JrEzltBgm2LnVEpMd7Ad4JbhRSLggc9OtOGeA3F/M1iWP4jGotf9CXKaFxFBcGXpNbLrk5n6Th2
ZIPaKZI/zHt0With5dJVO2wyLTBpLFWm4FZojJ7zZX/pA2mCcbgQa2s5QSCwDkETfA2A/1N1dvH/
eqaHM0I8EPoJ+PlFWSZwThGAT/mt93hmNsGy7Rj6E1CuRWKYA0Ma5SJ9xm88nunUJikQJyCR5Uk4
zZCeYw4db3yjYPPEOgOc6kcgunBiepLnodKYG7bEUadALli2aeyrDiekiWPF9FIWKK83fOtlcA/U
QcoaY6dNB69BIA+8atj+3DER6Whfdd7akqYVmKwehHOGyt7lNZnyv6iIcw2v6IRTRZ/cwfcC6gl0
4uUElkreIScsKt9ENxsmaASWTArEd1ry/2ruDpG4TEQsCLbOVN2+xcM2V5SeuwNjK4nu78qRc4+F
3vXAfdw2nBRor9lLpYlJUzt1mlCCdNw6kx0lzLZTSz4Jmky7JItLUKcuVFjI7g7+aJEVIkcwDfGw
PF/Ck+qOArBoK0F3MmzIeYsou8KoSvnirl+23qhvnr56RZytK2DrZE+hvVHYwT1NRpclEc3/QduG
OEXrOY3dZlSD7minpqH6w3fnY0fAXrUoWBuj4370W4tVzZUskeC+hQXVCJPHy2FnRUI77IAr6e+X
4S16e3MuSgrzwlay+vF0nH3pDQUIZ0vWPeqOdqfOV07tq5Mtl0G+rDmPr7v82pirt4/ajWe2jc5Y
oAnaaPKHZkAD9wGJosmqHpGBfqUXVEgrk4TSDpl8C6/lEM6+cXX2BGy1bNfg29rxswgoZq05C6Ez
+7BP9pEL9mQIVc3EUKy6Y4yLwYKXMCNAjbMGCnSgloRfdpxNAec2y6DZJMO+1MJgKqIGoCxGzbNZ
HM8FT8/zkWK3eSjc52/YXk9HAcEVz3/ZGs3h7l/og0o+g1rvKT71iqpqg/7eWXyRGzL0XR8ADmH7
ar94oe2mq1pg13VEyjsrOl8dJKNskIjk6TdLv5ixp4cUaCLht0mq3ArqaXdpw2mFCpvjK8xOI3Rw
eAcAHDq9y+i3B6gRkRx67T55sH9W6aDvCCmmBYwUdK3Y09kv98NJS5tcv/bdKDors7w7DdJbQeFD
ok7vo1mti7i00puAp/RdvO0DV/zd+Jr2YPK2L5jgS0uaO5wYDvBH5qCIS3ALb5uI+3bs/PGFcIxh
ABWs/V5cduPDVLqDrwwrmciod5ef0NxeQgywd1ACGMXGwIPBK2sBzpz0otqERnOBcGyXR8IpoNMv
e8n3hZgTa1dyVePcakklh6zw1eyKWymnlAeeeLa+uQcd/70EcIcNY55arjd9uLPvP9TqgN9m6YHg
zMPgTs+Tcyaoo5AunLBp6wZh6/+QZ3AdMOqO0S/mq6b3rl5PcS7UH0P7PR3amSJ0TOrQ86bBEfQI
xeGW6PesmoKOs5I033HmOw+3Th7vnxEx87EvguzSNOaXz4PfutOm0Agefx6ZfHcV/OgDRh2IyYvK
dlOC7pEWVjQUMQQgK73WyQiSEwzMfngup7ZkYUq5DukiYPFJ41HHXqMv4eW/62vQPV9X15OFrwiQ
dJTCaV+oh7nUoIjaAuKYfwtfHpByCqqyj47pMo8UWFsJcvtRvcCO0jr3zzAFr0X64cYjJV7lLpKL
mkZG9O/ci7iSaWgHuabbM+VTPStZEEIbkNPJCAAyWxpNMNjXLA/dka6YVmzkCdHKUVXQfloqumoA
wBZxeAYYMloUJkPEpnNnQqo+hlBOzsfzVOwqmAGLfvmwmLn1Hhdzoxpki2sGHXBOgHtFoJZ8NGvE
E2d4GI7ylh0VpVgMxSXIwBtvMRbC34GW7bjx5mSgZ9HyqSTnxQYjjXko1c0nNM61/MjDnKFDBp+k
57goov5rVg7ACfl35zs4hMS6qUREmLTuaS4EpKu1Nmqpkegg1I4dKSwe3qeZNQ62Z7vwnRYAJk1Y
fsLKTkp3s1W/aPEUNg1KFl27PAFLjicCNo1ZjNRtLt6yZulm8mfZTawtJphax+dymTn6O6vClgaI
Jug8huoCyuQlZ7zs/QOl2Nzo8zqI1bzOs+ywfSBBqq9iqoft3nGIgca0/+9LmiNZKRwENTBR8NFl
nw2Y+mJGM0MFNJcx2RqHu9+OyGUVFin44KTA1WXdMHIL102PDbA14U+lZUMIzG7BlU+rR9T40wpE
xnOJDMJUnJ/c/+u5SIPXgQKYTY2P9uNceTtP8O9dV/VDo32v+3t9jqFvI2U2cHDol0yYXDhqRvPc
/cqcBqQBGd8mzkUG7abr4vv3p4lz9fRDbIrrAKPZmvb6sX0fJp2BBVA1sDMMevY/v/xIFtHWZ4zX
fdLZrM5h2pt8SY2sKcdYuy77aAKfTLWUnvbbnal9WGw/4dzTlTw1pa1YzULWsBKhLCHdUtzjDVXH
FLZ2s6IzD11m1Sbf6xRNlrIfEEVjULfO3iP+lH1YwFjBiGfsXXyEf+xUg36tI4qdMJLsKvXjSr5h
LVk5Z2OsWNT8xOKmLwpAfHCGJGXBKqeAMNE981oSMLCHm+eYsbszHPNG0S8FH31L8u1xoLquC1iK
Ze1ZlQ4CXfJf6cnOJDbA2eNIx6X43FzK32d2VvUkduRpXv3c7u4bsP33C88AtEMLgNznV/vYgvhq
XHHBQk7e0yM5ubdkhdC6TBaBbMPSMd/doYeC04n3uv8eW+IldnBFla+jAByM+izgKBdd+vhRsbNz
p+lzuILiCiTLXHsPMdYTVF9Ghj+5vVOBSrulAzRhKcYedN6GATBiZXONMlppd0s3nKg3KWrzFFPo
ByJfzFj+B/WWmc1LzRNN/sH9+WU4z7bt0m2SUkjQqEeUSe0SpIEY6j2lNNyad9rll3Y3WGjU2k3O
TOS/yeI6WzNuDiYzXdC2GiYKVNd7DrJsgxK3Z7TJzJqt5keNC38xb7NaBXGMxlIViVub1q1VG5FI
xrRd867QT6fmcVz0DslElxugWfSuUQjupkqalH+TFbu5dlsATlYN1tn/bJo8SzmPTdop5ty4WMAR
2OWmS2vouEw+6gNU3JGp+5K+vufX4dA+TS3AVam6+NEAwTusoyABRuz/IVWGxQN8ocbv+jHhI3Zs
xtKyGVnPJQL46eYeroNJGZNqQ7G6XXJuB9nJcJa8x085BiU18VtI1J/A27bMeG/yCne0JXdgGE1U
T6z7aUEiJWl7fbLcBbeLLLABL/a1GmyUp+N+jDIaeJD/JtWnlYpb2wtmJwMXk5bf+UOfJZh9ADi9
9cLBVhut6tW5lWF1WYUchOr3pWQW10DxXzryJkLPO9tz/YH3178pz5L+nRS44QoweOlnp4rBSiLW
K0CYx257T56NlWOmHnRWQG1DmO1oLWdd9j/LDTPg2pzMb+6hS0U9lmXBEt7FD4l2L3ArO5FYFo2T
1JqphwB/Rptm14yM37sJ7mRgY0Jlpy3SPwLMBpj4lw9K6RUq9kZPY/aemnnrtKh0h2T886zHGRQV
QXB9qEkLaq/9OZPM2VqiF3mzfZKAOrkUF+BoSbrMxX8hR0FSWlQjpPiumUHbkoeis7iZZQdXIgYm
/EPO1vh9dohm8nm3gi06xbWsbA6quGLD7ivf9h07ZE9p/N7cHRTs6cCU5nUP7Xi6x8RjfwLQIsUR
/gIsUK5eg2TmRwqgvmxgnKyXgrap4hFt+9cRqzlz60nL7mwb3a8Dtm/TF4Ms7zPd611N4ARDL8ZY
zAUIpMdpkCXtW5no6smYvCVcsaAzndYt1ShUPEWGqiLBTaC2Dkw0GVLiQ9llTHh2PfJj0aEPlIub
KYatUtz7Qe3ybsqtaJgo7/0j98UdCWfzvzSnqbR2Cux1d4Jb8LgaawbKVflSwWupRsxEayvK4Cwa
1mxgoxoVJUx2ura9AL0GDEkU+ryr6Yftsc8tTct+V0r3VGA2kzsV6BCSOk+MtDgUuUadriZkZqAs
D9MCbN+I5+wyCThGTHmTYaw6d07bkX8bBahpxSTGwvINxnAmOW4ybBUql4yydlMjaqgy+XheTo2F
RKnbxwmRXrvpIZgHo43V3zcd/EQSmtMCd7RvcfCOmlHOZ3502bAot/9N7QbG8lNgo4Mt9LJTDXYR
v9hN5tR9TlouDAGQtquVVSiraZwKbpzBxu1ln7s7NiJoEHkHTtPJLUWhJruxoSRB3BynmNa1qjDg
Tfc2XxTm3Gic97nv4+bST9f0VH2BvV7DTac+kUwFEf2Vs5f/rgR2x0N54clCHN9ybdhJWKWMIZ/q
zrphn7jGToyWvq/St0/jNvejKl7AEXfm8oCnvoGGJ8jN6G9YGKAgLUEgtxrcssWFLIJFzbvSoBPt
blMMd8A0llUmYsk46QiW4XGK0RG00aCMOD+0i+VtX7e4WF9WdpNZnxAVKRp0d/pTyefArmPJLhB0
xiimSfqkPgAR82hNvISURpxS8vvAIQ+D3YQ+ghGLjdTVCbGefO+fjf0G5ilTxAsjTb37+nRkZ0ki
rod1Vf31IpzadlexIK086lC5UlF4sp2hBvMSxcUPXSlkF8blLaZIlcagfff9IQlIOrTUDe97ci7t
SlVlEnlWbrOX08D2jF0CY7jDcK5MySQ4FFZWyO75WSrrbaHSKPkwBjg9lzN5VJ1ynRrjM6dMZv2M
f15kuvi4AiqwbeP7SlnUnjkH5+fjLFD9+c7tr9G0mBXZir0L/JKtAef8/61jfLOXRA68gnJpbmTb
lYN48wnayACupSngMWfq+MuJAYLnb+dXR824/ZswhdhoVf0ShBl51kOi+llbfg7IUVlC6AQE/H4t
bvvAwsEwye129hCWBlUK1wjimQtbpvFXmUtoXg+8GKKD+SL9H9+OcmPJr5qFpl5u8IPOabosSYYU
yp22+H5UxRcUPSW8WrkZTR7iCvnEum7zs2mFFvTW55l+SGlXYW3TW46anbLx27yViKz+nuC2f4/b
BrTV/49hmyykoNWyZKjdyqs6b3HEo1CFONLYl6RgoOL3fqKxEZaDOvyMODf0Z9eN+HtJQTc1tz0i
rtrcb//ozl6otF/0z2e5U0v3E5E6SUUj4vrauB2H9SwbmKp8/i5kmthC2tYcwxMeDUL0fNqx4WZ9
jYiXor6VFjqTuTjsSyXu6qjlkEfuZ6BC8kGi9+X0QV78vDkrLrnkZJSbVfgA7kEHdT1vNwS8G/Lg
/6qr4gkeEhclk8A0z6FinkZ0JxB+r9iC8xKk1O2vkp5+uz+f++zhR6G0vQNUsDjARbmesRrhG24H
1dmXjk+T79BQCpxYet0jnB0Yj7Mjw1Lo5Jv2WDEAilN1SeyVTCLcW7me6WgjZiHcM2IdFYZqNxv3
dCow4l5/x6/1HL7SJTLhVpWDooMWLjx9s910e2TwmB51cQyrthtW7aYlNI7GmL8hWl2yzGQpSfYZ
jpU5fzP0JJEb9PQXSWzExvJM/h08q22vpgndANVSHIKWiaJzQL2OYMYlf72irmA0JUzD3F3oGNgH
ypsgsg4etH9zj3B0abVqS392npInWvKXTXNWMyMu6suMqJaQIKSdCaxcMRiAflSowgvvWNMBaXgg
rCWB9XJYkG41DQyiuVUM5XNNnMmZn4wb04FzdPWXaNriuckAnDNuH8IFghAc77bj3XJBmz8zn9uH
m28sGqaxfc2Czq8d3dxOEhcxgF5oUZGty7Rvq19njsBzByBDuHxbBKv+z2dL9VwM7Z71Fg1FJHkE
06jULx+olrEJckZ3/twdxlAZHpgZjO6qyKxCbXPb9oGCod33eJyhpMHN/wYdVFljuVjrEIVKhYfV
7k4DfK8RT2UFw3gUtXlRVrLaRa82hQ7luyk3timJDzA13jN+t2TWlm7KotMp0cjlDCceBI/pyn3Z
vfSvvWtfh1+yS+Zjf3QlzTrw01sAbidT63l5M2GaWlzLVH1+FpqU5y4RT5RYba3QpX6kxnwx5B1q
G4yjzrhkw5lsGM82gpAOXD/clubyqj6D4CEH9ic4R6o28uf9W6L+zpfywHAeCnDianZkLlrgPmku
Jt0ZAoSVo0QEWPO+10LYk6NCl8R8z27D2w3xG5I9xXXYFQj8+ZoLtNkoRda13j4S6JXCcnejdgc2
oVpt8pc5339Nk/XbeXr639HzNY9r3h1TuMCtR271zfQLAQfwil+YkS8Eqn70qZo3KgBU1tDk77/K
Zfl7JPwf+4Phengr9YjylROs4uoX9qzYzJWYp95iNj/93Raa85oepuVROyjFEREVHYCFmZ94DOfx
MVLR69LEgMVAMI255bCiyQhcye5y2wZJunDlJtHBEh9OuLcNNpKB9fCYG8Pj6Jd9xxfzt7n94bEF
oIR4/dDXoouJcSiKw4qyh8VUoBjDw5GiXa/DtDtT9FWE4pgZ6X8+9MoyD1iLk6/6oxsGGfLUNFlj
qJIxvmcUf739IbSbep3C+Ak3yZvhZWa3MRsAaoJ5oZCOirtJVERf3Ywtp4vtsHBnxXchlS7VbjLx
CPVwIYa3SjhP13sGagpRXaxx9Kt9lPomPE1CQZQ7aJaVzDTDuy4f9/31B8sGZDAMNmBhbTGWp34c
XcupAqrIxmjne79fMF7dfIYY5VUvomZ+BUs5z2M+vxbGtNQiRpxTVBRDOsbkf2gH1pamOZFEJDyE
HLTdux3PCNr4ejoK464PX0zKL1TGfw5xcEoKkwViYhBm/CCHCwS0stZTqDWx/6sHHW8pOpAzlI7w
IHMWFeaVW55iz5mRYlyD8oZJ4QcLlYkbvRsluVUYgMQlFI8Mxo12HrFnCb9qy2+vGdQsWAV32pJR
mXa+JQsX0BWGltDrSOZJHHhfKlFiv90ntYKaWRXb+UdlZdw6bjgo0GSU37r4pbuTdRfXx5cRvAF5
98i36AaOstWSyolUGM8zx6mmb1k/xVwy9iq3TMZ0eUuGvf6XdzorRic+HSroo2u/LG0XxLmOKSVZ
yT6/eFeT8riNVkmlB+MnfRUQ/pXU4AfLhlPgVPAY8zb1sgzJKwUvrZAXaaPQqzOYOwS0TElCIqpu
Ywyl/DL9uPr5e0b2TVtaCNpuknR0VtBNI/VaiogUpPy6d6BAY/+UfQ/QfpiyMOVMiX5myNxoYDkW
prLCgNcJkTLeGW3noRcgmw5SYXBnM6XUgf57ycrPq6NIOy8HcoV1uVi5xQPMnM4vuxppNbR/p36g
Ijodpmg0VGXgvQmtRG+ZzNZsTJRrqBPsgtYaLNiKE71Ory2AQLcgNWFFt+xWaPUveScmXh8OztmV
JXECpLR4iwdrBBWrluJrAL/sE7eTD4EC8VXmt0yvRBXUz+y+abBMPgDGZk4sG8z6r6iAalB5JPjl
O3iyT/jiKeR/Ek/pcxsKsAGOPuT6CWsaA3o7QlE2psAX0hqayyPhBtdiRq2W7MGDAejk5tQPcI1U
4d0Xt62E6JP4Tb1vBw/u3XjzKSyZTRunDQNMwOfWFFZfN9d+PzE00YzUg+1tnpUiMmVRybxGuVjT
+/WOdlECfvoMlg5V1N5npbIz0OwRgDOk8DlQHzwpmrrd9hZBTrgmNrcA18X+OYbLOBSyjjmEFR4Q
JHv8kkZSMxCsoZ7uCWF+okktiwmsBQRpfXbk9icO2h48z7f0j62oxh0T8OB0o0ZP/0iFjqZCjdgw
LyVB2e1TPRBRsxGb0hhgtefDAPyqzYiMRvg1OtKothBi6YSWAN6X+sxOR8Ur//NnuE5j3eE8Doaq
QMgLLou1t82Obtavr8llbhfsDTtCzRxpuBqFhaun/z30DtoP9Bhpb2VdqzgAcQ8IVXr93zLmvZFT
jyZdlQCI73Xw1yftcHrGD9AfM4bLxzxZsslMMcu8fIUCmQ96GAgZVO5aYQgEIx+Hf9NZQJvG3VGI
vWqTNviJ7RwSVGywDYxSPGvh37UHliQHzwXRi3ylCLJnuz2AAOsrj3Ax67fzEAuDrNyK0uXGeqN/
D35sRhtRNRN1ePfhDKH643cRbA4uqByj3/D8ZBSjTEqSV9D6v7MWdjDrGd4QQG92uSBEPLu4/8zv
67iUw3cdTwBac/OjyHLQPLGFwof72CpfdynrLif1a1OxeOS70KoglPjxjMr4yiv+MPW3QSR1/vZ3
5lYE1NJDNV830Nura67yNCEsCcFan23Z18eyCxsPlOcZ6j/QcywXEiJiPzLaYyNaxgNUGvEqi6RK
4t/W27lwbKrGR0QIA7zEhmAVfzXkf6gp8lz5JDggoenrbq+S6tdnADYBtxfNoWU1o58IZaHkvzs2
yu6JbeWbwgBrxcnp04IzJ6oe9pn2KgXYkF5FQ4kFITutC2MO5WkEM4PJHI0+sdMK6PqGbQYB/mFf
2LlfL7bWSeTcHBMs8+0KdjMuihcSj74urTCbmbH6OKbVzRCrFdBZSiEc8JSeO/82i7PL9sIUn9dO
LePBvKK79I8SNVgSvNMEUf+8NrlnlE80i/2LNG0P6MA0nMXEbc7OKyNl9QO322pBIosVq+3/d2dC
4W664QwxS258hEMV5XJ0PgzxwDaKJPrS6lPhqv8cnl3wa2pQ60ixk1RNdCBa3q1oHmej1C+stCUh
/1kLph+DP7UjN09f5099iZluP1i6RVp8gOu/1/X1o/9U2f2l6aalIckxjykm1HtGMKTIWCu7t7W3
971lurYSXXwIa7Ngl5Vwu15k6J4YiwccipDuwKWsEI3W6BR6L0PisJ6aCWV4IxPV3LMa7u0mYwin
mDksZUBXQRpiprbRbIs1MBaOGVq7M8R9M6T+P+tQqNv1YJLk1bqyKlobuAcOoVY4lJbIPytsWOL3
0cksq9NalQVzypGut8i0gpICzdMLv4tg1a4ZCzy0/y4bQz65fzIOfhRb2uabQ/vWCbBK94ObLm+P
vaxINHl7TRNTmZEKc4W2agoRGTJnAoxZxzdc6VUX2bj+0sZN6FHVyCV0nNtyQRdbjnhHn/wkgqrS
igX8NfIjbBqjFhi2KLZP0qwC/mynALta6bc+A0t9BhsZFmgMtyJlBLjD0U9I9hEt9ERxz29ZRSim
+lIBbbmMXCTL24UVTeaTzA/abxd+aX0HpfMY+NW920B7qDSqpXbAw4H/ExxYqBcllzTn60PV2hvb
iPRxRHhBtPD4oMe2OjVx+NWUjXshwGDgMJ0dS+uFR9We+ZmxjpMZvolQYhqnhTr/hcqBd8LF/jCk
RorG7PrGv44OmLrpob8eWl/lDQLReXHLzJ/z8w9b5ciNUsqDorv8d0Vp3ChR1CMYfKu/cJCuwhq4
ES9RoBi78hea8e7xvNGzaIVI+JNCmuu3+G5tGzZyuBl6dE23ChbifnltAPVNlaaH+2R0cYnJ7f/z
aIL+OYG+ybG7dB/tEkpmbA4HVDCYl5s5WDdpyiz8HOhKe1LYGBIm3JghL4sQyvTFe2bG0atMOlhd
Etik0mSwQWmxFrMSYA1FMU4x9anA012C9H0rlsfW+8R2hOo3Ejg/tvWudA7bEhYWFBz6kCaEk/Gg
fi1aTLIEjXBanXIgLoU+ThtdRFdwDME0PmJogMS87nV0lemcYu1NcuHYV2rPCQOuRZjfM3PJunau
N6WMD7bythVIjjK7NKCp/XW+JeLofnqiAAxf+H5Pq0Jt0vq6LDfW5JBRZZuFIq6ek9AKSOKgNNua
hpJlUr3HVDalYHavs2+ZFqf6qGB6kbm64PgtWsV/kCsUMf03PKF/eDfAcZkCLeDDtJMNU5DQHps9
reOm9dz0f50NQuRVtXMb1lw9tS4azEFj3Tk/0OUqJ8y5I5Mo0nrGi7ofQrOKprFvNAUfWgU7TvA1
jE7MoKyDWx5VR7BzYx3mWGVp0/epO5oUOMBqZ314oIl9xAcwPBzC4AyabEWimj+AMo7puSDVjU2P
bGVFtzWwepsAPQRvB1cszSvJTBQkj8MR8zkl5msrf00KP1aWMwufIpMlkvuiR+i4MiJTCaQBUn61
w3zC1G+JDRzvOdplhB5Ha5G357OVF1CKJ4Mow0d2SfKFBGPY8k+3AiHawAnb++GoEb2PtxzA0hEG
h7kMf05InZKCszeyWTs9Ti9lC3as6E84TGPE5doiCxyNYciwjEqORcgu0Ee5okkSTN310RSpK3+5
uBU8A1ks8/bPW1KrnYCJAMG+bQN/iEA/KBBkMVK6t+D71Ufcf7e2+Zlue9yKO2hYc7Amrt/gxDRl
nLYs8DESmr8YQHzy0266EEvAeIVBX8FBW7p+eLZi6Pnm6l6wAEfzmNuBn9k8ecgdC/bAog0rbhOY
jVE0ePhTFt0Mwudum4gTnGIcvBjAe2qYYwygK1W1+ohojhIWVdEfm93ekUW/RIUBJdVjI5Nrr2ue
AYSfsMnpgRdEVsEQeJa4uQgG3NkqAkBngPmsBjeENDLP3lm4Pk4WrJHCgiwsZ2VFNuf5UySgdLPt
8RpZvgPcpX/ngFBEzvrJGXOEKucm+7SkYDAYh8Qu2866ZEyhPWjWasmPODpBQ8voinNuvn++2HNH
GkjPN8DU/7Jm55JLS08XJdn/tFqoUK9PYI+TBKyVzO97WJtE0e0qmYx9JKMXLOr3nrTIXpjV02P5
c9A5bjWW1L9xnlTHEqmGWTZZDAf18LsXUB2MbXqCViYt2O3IknGkq56ktpR4stImeC7I579H3UXR
g2NXOHAaZZP0v3SQTsNIgjTfGCgjiGsogAuaMVXNSp1Awm4P4WCpS1QEbQby1jdaJ7r0uKaEqGLI
bxFo6PdYhad3xwSCB4sUk5YQluw8f/hFMtZ3wQyCujGw6Uo0VOW1Hnuje400szjLzeEw2xY+IbuB
VNq5k/MPRGgiHSts7SNoyVh7uaP3AwWefGRtzZIzBfvmFat1/yKaG3GhMRjAxyMAE94ocg0R3x3g
OAc78X4XQWY6dWhu0n5tFZH1qbEERsrZVuBuetBsL7N0zXzaxq86k2I+56h3+XAkMpurjbJ1sfSO
ugf5BcF4Ozns+n9yPC1LvBt/WBHyIzOWXlOUMGo9Sw2DvWKS0ChYbnJZkHBuKpENM398gDOm7ucn
Ho+S8+f5PH2hyVO9bENfu2aecnp5e3D5JvZlrlmmuvRfYyc++BxM9JRVECruonlKoQsC41keyP2p
+wlWcZiNW3BbH/8R5Zai7vTNUYGqkRu8el96a+g1jsGBBqTG9VyEXGlh0IfbiRAOTklW4owfKfNx
6VL+L5MN8HeZ61Hju6HjuQ2k/jAfAyOCvs2TypSMEzAAM9NE7YewWRP+mqFlV5MSSZ9yppiyx4We
ChPOnyI18fD1uhm5gRwhzogG8oJRb4zouG3H90NGBFVr6FC5eavTsGF8Rz2ZHmOf11bd3gnjtuzp
EPxWwas/+5lVdCtKR1ON/6okTqH0ywkKdFozKCiAwLsOW4jA0Z7W7MohCnMDozGX0eQjGiJsnZgE
smp6QURABLDWp7iHNK2bkSP19EJHPGqveC+6whfwCH4dLAfqfeJrT6nrAJdPqlV3iKzc3tyNFaOy
RuYVK54SKH7+L2ExTPLkdJ8F3DLc4mvx2s3j0ByNIzybJgtA3EaPzd0wdpl19QEGpUPmaiqd9ont
/cpqGDWs+CBm1tPXSUvVAP12GOnX1ns7gD4iTTbtiKSUaTt4/oNH29SARKPIQXL4NT9wbODERtYU
SWXfWsJNHSrXvDL/StW3PC5hhwAYDs/c4A/c9WdqmRcL5dTp+mohrTBuAnlZnrpA226e8CUZLki6
T5p7Me+AyNsYx7uosAFiL9c3Ur1lCI2s/5BbylMb7Bixseqd6TyO3M6E0zDCxY4AW47+ke9hdTIC
9iTh2uh+h2EzL/CgHIm6KRqzgV2wmAzfC3D04DwNJKfCz3cocGcoHhoVEdPb9qy83U7Fye9jEytd
brUVltCdKLH5zhunkpSqGm1dS9ppGxzChqc47Ab2+f3NKq+C6q7LN6AiThDxHRrWze0wqhEg7ZJ/
UDYnZ9OUH0ehNCkcOLIwN3wAsyAmhWftCFCYXHcfEShkZfrpo7Z8wh4Sf0FxqzrT//Nn6G8K4wK4
cjkpvZFrk1eE/Rh5KCmAlHHMVQPbrEmZ8zHFZK8Qeqh7sTCC9wu2zKNKt11qUYYWoR+f9KJ/1me8
8qvmCgwwiOaVO4RNsBfpdnNy+QX3qyh9rlVxHjHg1zb+F0TSLkFfLgN/ORFEuWgyzFx1ZWBTutVw
BaDul3vVhM94ire4f3TNcTvbTluWWOdWGAPcfy9tt0M1Ux2ykrMazVeBSkFdkYeL2eaVubS39vRS
07abvbzWulMgnD6IW4ik+EqmHP4lD2F862UOnW7wMm7tJlQkjsVT9FSmKu+bFbbwfojUwRgtLN2c
rqpxSWjJqnMAn7hG8EvopgTzvnl51qgyXzC+3PimkY4WteJ/ekLIw2vqmEnXonxYZBRZUIx+4Bnu
Ucy/9MvYFV02xPI0nXebHEP+/VzaJ7nWNv/yQUUwkr/HDpBlkpSJyZYaHmTCZnw/KWoQunTAWAmw
tQ/ZXXcAadF4CvWFKqJ5ILwKa3++XY1BHw/MTToJIGQgKGYsBlwm58r8FvehMiJ7tvLid8mp386+
IhH34eA5jx5jf6Wu6CyseYlm1JVlbp9IY+WFgTvRqpvYvuMd+mimbcXdWTpQhu14ie4BXOBScWnH
miGyTptHvJsamGeFK7Lc9c+wovTJ/FSacLzTFvxf3THhYn6zzZqGUgNpswrYHyuql5xiBNB8ZLVA
LtKZTQ594+iNtbohhlVP7Ku6+pRboDSIhM7XMT/sigeHH/1uExB1Xhdu2wSESX6KhgfG6bdVF3NQ
fLjImdhyD5GPYPiUtn2NDUO21At6A9XEU1cdkkfipGN0d59lxINNo2YpUk9iYztMBWMK/SMqxQvl
3bzj3vjsYtYZZ9rnOXJW0/2Te9FladDt+NgbFK5T8r+INF5O5OZFoEud7+uOmrLcq6eF9j9I7HdG
fQbgj2kb2T0ubiuLBbx7WGsw9xQs4OP2FnjgwochZtRzJdT76T/jLDsz/c5tZzZO5cZpbElunF5R
BY/xxDblP+FInGeUQfp26YBSx5Qx2WugnuvU4uEr1JbGislRAeJ5hs655lUd7hbdkP7rBBrDCpR7
dAcmBQx1yQgC8grSfktbvJnAlwVmN1u8biviwPRmaKJNWUIJHjOcwPbEqzCQQio6q6sfLdbNRobT
hplOxILen0VJo2Gm6L4ZvmSMLQ0FU8xaH9moYj2RFJvtnUTKBKrd4nB3x2FHrVwUMz6jQJPtQMEF
WKXG+FMnTSuYpcDDB63/gP/ufaF8qp3d2/ir8L7m0x2lrs1aWtcbs1nvzhQBNc69xA5rf8mIaMNa
F3qIg9HxxLSF7mpiS3yhlnbvkL01YR3fvBTfJXsSl7814Z1AHiN3NvHUMjmQipUNHL4UmZoGlT/7
9XCSVFA8dEPyodoRMomfE5A7bUYoDaoS/kG9+0tTiFYjzuGStVikMeSdZMn/kmQraGbno+3AfOb+
YeA+PqN+XdddT8f0Rpg5ivZqRkGPVS/LK+WtWUzucBCYTjnBmcKbqaRMm7G/YLrtVOznLkR+v1Fa
H+KIDWTj/2+r0O4zrbZ4+cQVI81YMWeEZRyJH1EBRAAIN3fH1Ig0VUeRZJZreWciacNUBUNMiqVV
VsRJUOS7RxrMV0atX3RDf3hBPLB1TzotnS8jkJ185I8FC+RsskCF0qOA2hqY9p3jWSQkoJFZIM+o
bcRpcQvP3oZftWgeaYpq7htVbjckNdoQJ+0ONMTU9qIrj20gbZM20h0EplCBPfGh20cEBth7D9LC
iSJCotiU0Wcys5rAqCJLtsu3e0Cf+yqGLvv3WOoYTq5m4ihM7CFndvFg7D7PfH5n44Kbd1avxNuq
W2hlJLdaCtPmhEZitgi6h3sJOAYzB4667At0WgY2L9r3j+MQZ7aRyXACd1fLR5KtSUg0Qi5u9ZLZ
oGfmPO/DL6Iv+ItwLsRqr/E92ykPkxSl1gdZR3bNUi6j31B0iPN3+HK/nG1PHHr7YbluyoJMIGgQ
n3mPExA2TvkOGaVsGyHj7jqnngJBCKjSW7RfbFLKeFyXWxLTZ3du0Yr+NzErlwSyqE1dcJ3QqwII
MWC2CuDm4vT4XbkBrNNB5mrFGoO/OMNsjNYTMvTUxuoYYq2Qo7bE5R2ZzFKTNMPJrOrratkqx3MY
gHC3Y+/OPnPRHkMz6AQ30YIvfnfIRlaMdqKcTuMHZcT8F83vfBfNuMOe3qdRRNaKaXdDi7rkrTuw
hdwWztzIZPgVC/LHtjwQpM1AxYrbblj6h9PMAgmXdA8UL0fS+v5lROUKcGCCJbAjb8fZ0IHCvmVT
BhgBC/20E7svyze/Kfa8AsgExOqxW7S0wFUf4Pg7OccHZn7FslpZj7VhlbLNjofo+uS/zV9cynFx
rEp/q5fDs3zm/Bj+zyPHekM4edLSnSVvTTKYB0pqXEsedpePCoYGgNNGWBHCMni+ROIKTwUCnRrH
EP3lwP5YwaWl9pNikhTr8T56dEjrYPk7qV5rHkTEtpOn2RAcbZT+pT7f6G6b9Dqli9Kf76+s69Os
Whm7XKgK0rzFJyuas1VK8OBdY01iZlm/jvrQLdGk+C/ukYNl/UZr4a5Xh0EkrxO9yqbBXZGFlhXx
hQF/a2VD73aFF0ATbY0onoujQM25Y/ZPtOpcmh6Mr9pNLLDAzAGx+RThx0VocVYxsxVnVGPO9J58
Q5h1lwai/L16jLO4prG3M25VDkd9Cf05JG13WlIcvoGP8FFQRGih1ZxcpG0B1KI3+k+4vAH0qQlY
cSamfiKIfXGn6EIIGkXOWUpU2UIjGppORIaDfQ4MtDfjIdA0QYqqhPt39O4qrNvNg4bvtRWNYy9o
qmxJbYmtCAXLqYutEpTZSpkZc3tt8pYrhMNu5qb57aATP1x6kKn3L7mtFSY91lhD+a9KfN32RnyY
s+MpEWpLN6d6klKUUdSb7ecGDWBPaPrio9E5dNznwKVz99qbLxYsYrMJyXWHf8Mx6BPsGx7HoAI/
KiPxC6ZN9OwL9bhOqa6Y3F1kL6CryaWrbGL4uwzV7D3+OangkCZqS+CgHGGpcTrq/ouGEgDEEKXZ
e6F7dHMoa/v+oygWs6eSLm2pDTUDZSfz/0nGHz22Bo3z2H1maaJIbwhSUT/5Hxht4dYmP/ZYf3Bh
Xk3zSAagvYeGoBQ1p4+1sKdTBsiNSPb+1oXhdxsbDJFkM5hwfYwVpC0oCwvRKKX/iBUyL+FWbDoR
NdvnBIXjYij2eTpIWHy1Yv8NWgMUmsIAll21xE4apGf4pVDZ7kezIBL3C+DA7BbXbVjMQbRBQSio
MiFMVOYP+6ulqIRc1ksONNRpVVS4RrdW1Ee2/nj96hvpL3TqEd1kwjrLuAR/rFDzi5pGrm0pWda1
YOxsm4U5LHaT9fZu82jF/iERHgCFs7jBcUKVuxKqEtHPusYgThMsDpmOLF4O7qNLyEHDQ3cuHLHr
LEoHRHltCP2VWm1ZMFhDExoGIYF1pg0HZ4PMBsmU+scQnBO1lyvBmwaHKqmIYZ6uzHEmpK7xW5qH
9+yey71Nlzy7CoawiuwMNHuPMYEVjqBg85+njncW4RdhGUA4ERvTEWRgpHYcAY0NdxzhkLL1toDO
ZPkIBmdc9sDa+Xok9bC7DZVGR7yGzHatLxigZgc9ZWzW/zS4gFUs5j6ZxTrJBsypxk+e72uZuAal
vLXplI6F+gccrAsm5NC8dMFyhILQP/1n1Bj/pQD1WRO/1wG4NZCu73TwHIRL5rP6GifGhWhhCPIl
xqX2TPWQHE0UpvKa281dHegTn9/QwxjDBI5O+Hw76EfT6V3V7tgZLBvtNvVJ1omrmd80xdHo9oyI
QpB/ESt1aDYy7F137+3ueXvkXyfwnnR7SvG87Jepk68A4WRQya+nR9+ravpPlxap93YV8HRIYEGa
CjLYFKB5ACk69KiBMKHTfFYMaBF+60Y5qJNzGcjhn2zPMkj4GjU27tZ5p5SfQuPepQl/SNH3TugQ
pN72LSAhWIIWmfLyGmjQxi7qZho1aHAAbrRzS+ull8sd8S8hdKTecjIIeFIf6ok0qCXuo7VWaL4Q
bGwgNy8tHwoJK8UFUGqMkIzUepYUyiRIVGDE937/PNvr7+PFi88z1YaT7zLBRwiz22q/v8o85sra
xVXsKwgFiUGLPytQgmx3/jeixQlyoj/ikFD4ayQaKZQSHFTfjjNI7fUyTQqaWoMYXyDnDrBttjnB
8R/2hVs7fTXvgdaib53rgacxCKrvlYnx7MAU7RQ3hiN9Oo2lGq/RyUCEWcyVJgiOKMYIBpJ46iu7
MJc3cPi+cjga5fZdQ37mNCUAvwgY2qohkr/9GEc85acxwlFkCxmdCDJFQ7l3e1SQ/7xKHlbH/a+9
FBY9yz97p96vx8xxLSalPwDIaC9Z9P+cq4+hMtRx7spZhzuMA3SdAImW/ne005iMwytTMqbNLTS+
6ZktzKAqXN2KUWnK/XxaGTTnSSlPEbwmAp23S4QwQEtNLZ0V+CiUJ/mniqP3zRY7aOfxmcBGuDdO
i6OnpOiV9If1sV8Ne3ko1JkKJ/rM2/7TTldbwQUACI2xucriH6g/ZEc0R3UyakD/VoVjuTqX/aC2
u+HHHWosr2ou+WC4rj9kPnohvMDFO43Rv7+8GAhjIn3ObTeJhnYl90LwKLw8wtdfz096BuxL9cDW
WCWgW/4o2asou0sA5BUlcNS/DsSeEcOgWnaG/3VYu2Brsx3xuarsMuJePYzHtohFg4tkG0ZcPUfn
YGlSw1AX6qeAS6Y17DzsZL5oawg0ikBDluMHGuscutIGZEPQko2K4GPpKc8Jn6Sy4Ij4drABFBsy
fwxtFbgwjet97s8pyhs63mcdS76zlgBzOWTvSQo409ThT5jcmn23PvOGnQDo4CuzKqgkwkgMBqwz
OHh1/r1nezIgSyVJ0zJ6vkIoVKmZwUGLgujUnoxeyDi1NSCnBR3Iqa2J6dL06KVI39/DFszE8iUY
kQOAyhooKvmax+MH01+Czi2KIGrG1Z5AwHis+Zy0z55DyzZpx9AH6sfH5/tC7NSQhj60xJbiS1iE
Xmt/hTeDRv2PMG6nT/tcC262up0mHCrKRQ1MGQKazjttNFk0t2vgpRNCGil8cqpPKpmu117tLp+w
v3hoG1HpsRVhADvqBGMv4FPTlnagtpviBQrbnd7LJdi19rgmbMqBXk+rD7KnQ6RWSpdXXNNnN80m
TkBE83r9jp8wctQFldMtfAcTBhYiof0NU0+IgHpHL3xUSUVpbXmILcIuBMRoKW0SuAi3bID56CjC
YXIWMPg90hXnIc+z+MrqhFlD3+7uJvYyAXexHAprJo/6Rk4a0DVspbnjPEpi903ERXBTetVLvzfS
Hcj/CQyryCAZG4eu/q1DqyzRTZXbsoZ28d4DjnDVFG/VruX9y2NUu3msZ/axJmxZ+p/U+5AV5XpA
ZqGfJ/uAigvgqTMkbXzNuexCKkgNjnoAE9pIl4cvhS8x6cyCEUxM61qNxAQRVSw/ITti0xPSkX7Y
I0HmubYoRAvHTsfyP++/zqrNbnT6VLSCj2jkzrtNCw29YPmRPl0u3P09JhPobcXTJ5QHhzFHGPKH
o4cdsT3In5sBY1wTteLUqPuC9nBaGGPgJoLHAZLeXegOHJA9ZIv6hct9bWW7E7OE3C3xlA/ewfCn
BxYKguH7F9y361JgekCiHhLu47Tlks5rk1RIaZ3lZlgGV78s0Ptnsk+K3KkrPdTpK2Y9i1G1tRoe
enSADdV5Oc1N80cS2dqSKeBFsHVP1lSEkprr0ofkqMEsTQeOO3jHoxh6pKY3A89UBLQ3BWkTRa+a
AsGmsgN1kZCgkj3b2F/Oe2ZCh/3QTJYdqaCBwKBhDpO1mXkwUtisFIgD4GlUfPV2jzRN+uDqKqh0
n+meLeO7ZKbHtRWGv7+xNDsW3DjFq5+HWdTrS9hd2kY07nuPBg5QgWqOzXqnfMCSThNJ1SLC2omE
WeaJOiSD1TOdYzepukfkaX+qW4QZgbH+IwjXemKYyDPCIGj07OBZERIxxNT2kzJyY+I9hnBJtQ5Y
MBlB0L25tJ7lbrbX6/DXJs17zpiAIdci3o2qwl9l/nlf/MB1RaHBhC7Sw8l3xlSkqyrp0KAagzBW
enrxd/OfLz/j4tCKQ9jEgsLQPb4eSp+PECy9ykHe4nYTAXvaxq82lBhQTstleKGjbxd2TULkpjGa
+DGT6GmnDFvIBUnfvdIX93/LakqHs0D+lkCJtqtcIlymfP0SZGfHlwYQSexbttpEiadrHYcUeI+G
MTSUWkMU0PO+/Xk2afOsocepaeiAKLQuAOAwRiken56Buuivnq9ZIutLwZn/qhiJ5uGb3eQusiAB
HMMZVQVKVrr0HCWuYHHt6FyC5V5ziEHp4Lp4weN2rH+4hm9dmOr0XKnE6oxQELpxzP7kaA0iJI+2
MyQE3Yc1zGpW29Xu/GKFvYcrbyGFV4Pr2f+A/2bL8Y8RlQAwWewPxu1oNvyOK0RtQ6OMH9FJ56U0
twtUL4vZqVg4aSyhpdYJklPoPHBG3g3ddOjF2XqErS243OEnzBJI5gR9WC2/Ciy++It22noQBQh3
r8u2AANgJRxSP8TSypQwDZkRZz65P1uGw5d1zxx77GssM4A0PNpuTUEmW9yY6AwI21U6iN90MNIJ
MACD2q8vu2+Q4JDWS6/1f2GxgY4nFK6wif/GJp+OTnAtJpwXn/ZkSc+3uunoZaO8QMs+rEugAeLU
S3AsKsPM/qjvMReLmi6hY+TwFLuogRoDXfHzhtuIr3+qm1fyhJ+v1DtjIaL3/yE5f/ZgaM24Xml+
Sx7QjTylJG3X2eh2l7jlK8hozUR8yhnhCreo5Od876VsbkXFKHzndbQ6FpQikNEIHmf/Jn6N2I4Z
XANjGKPKoyI6AvGG2J+Lt8q59fIvZJUZa61GbXWzpuj0HJvir7oQ17XhQs6gwcr5xlIZx7QYhG4L
/u/DSKEjGC6vrfSG6ydOgnOSkEpv4/ZCIcOTbYOdaF9UobS0q4p2hUoZ0dIOpv/8caQe1Fp/3HDJ
pT0e0ab7tM/WOzoulND/O84RfL/YrkxZlw/mHIVxl+saT93BBhISuhKdDjaAcUX7zHZgKaV7oDF2
cFosyoiVh5ylzD96vG/Iz+43+tePpvVkiUwPfGf2zOzg9UKcmUe0pOksGF+gKVR+jh4EfCoKxTDl
wK4R9MTRdtvCCvUu5H0vLbmuS9a3s0jzGe4iuLth8Rg7Jo01c4HOscewhG4wOh2B19H1dzg5if2M
ZhXqiNT1NSjhpHCRJSOmBOYJhRtk+H31RIJjhep4n3ybOMMJhY9iQBMLLCH529dDh6ErNh59N6wj
nnNDoNByHJp29WMnQb1KnZzaeWPsM19+P5rK+64YREZmFcLmBs/lTQEFNKoZ+ee+N8Bt2I/bOOy9
hRrLtcOzTVnQpm9AuBGHOT3ZW9SdKlo5hFvaIUuzUbSyFj3drINeQT1cymfpFUdW8rBUKXWPh13x
ZoHa4chBoBPDEc9Eaet0nziPR6yk0CHzpsi4aZDfTTXfMIEm8NvkC33fY0e+7YEROyIAnytfYlAC
X0LIsS2uGeRiUQn7JBbx2yKqaWxtoMPJLGI/xrkEp4zLdr4GAsHFj7Y7JSfz1O5X1Oulfh0eQ8Gd
+C5G7bCdgqkIQ1LuH2Y8lCbgKuJSxju8O3MvCeqhV6JuE9lzFOvQ2ZNZGbofhaRs5ycAQrCYlo3S
C6gtoNY3QzyerqmzN6dcn7kfFctbMsO/XMsUDc9A/ca/8s2IJNGSbTjXzVp4LdaIeBqdffOQwdvn
T++dCeP5hkBnt0LbN497fpRxGOE63ElCe64FI6lYNDe8HcB7v22h9ukuWRimPfi6W68EkYMo7BYU
FDbIb+hw7y9gYluRAWgDjy+936KFDL5qNMictLUXNqlv6tFjfiN1UnQixRenh4H2MY+jei2Zqf9e
Mipev7pP+XjrIX2lyZV06G5a/KE9K7yHVMLEHP+5y7nRvWVbIZ8IzlxRLUACwgOSVlsUKw5sEtwJ
Urg3dil6B2VLpHnFbaLU1jcxeXWGr1gC4wco6osPoVY7ucmbjcLmbsfmkCYlCZL2DZ89l8Jbvm33
CP2QKWPFluHGipKe+PcHf7eG3jy7oHFcozkkbmFM0gRvUQALl+mA7vG+g6DRF57oZDmZrI8tBt/A
xuxHlSZ+Vx7KMX1QyMFXWmeJFxG++8UidNw4hlMEPpJnKOafIXODJ/PN8kcymt2uMuTppoF/mjiL
lBnZL5rDyGGaXK2MzWiGnX8KIuGm/v9WSuJTgq50qcfmMXDKzJRZbw7WDzDY5x27y3curfIH2jSE
0aRqf23m8v1mRc21/k7JcSIZ3Sg9vdklHH5+Mygxzu0h4gDQGel087k+jymdBJdSy0AnVCxCi2jA
6ChTCsMAAxd7uvdkXD/8CPqSbY+PtNBlNrL0ml7TcDK/WU3ik6+UfxDig/6sQiBH+82kDbP8VjOO
orSN4t0M+SwKO0eFO2rpX9Wp48BkN2jh3/GRxlxY76TMtm343EZIxeB7yeWtXMkS3vZVRaQUcdoH
7VF4eBwfJZgkPaQlRRCErf7IBc+PK6CzTkxNfwfD2rgwZvPeQ95fafw7oWZseiolunSzmHqgrYiK
T0enPWhTdbVBq2GSZqxRiRUux7RW/PQdUy0a98c8pNSeLVPP676rU0Regn6d/RjGexJ+pY8CwnBL
zin/IW8xZJh7aCz7+txl8lmNawZsMO3rkBa0w7VKmqJ0Xq7gBmG6U3IxPTmPv8UnXQ8KPpjLG0Gp
xi3vjchecIJ/3ty0lcaLZaICDbnLEOJEFy+mNY8mWj2LjJSzWmV49QPauoTbmKerGctgyhzccrVH
u94dxv0FZOppxKbFj/I8gCKfH8FvIRALey2VjlvrkPtyorxFXw1E7HRSUeRFv+FRrk/N9jdOTd8Q
9twEZFlJe7FHu1MsfTbWf2m+ue7ERS0As6TrQlupca8AyOV8uXwERXKblyZ5n83y1pIVRmhrRLO1
0F28/RgvYGL6VcPEjr9ltrBZuc5gf/WF2KHQRVzZDaQuQ/MXlrj7mIu9UTE2MQ4jLGdiNgFmhaMK
x6uVOb5PUImNZV20oTouWGNB6OrpL5n99xD9/yZ33MTZEBnAw4wfW/Nzm7kOd5XP9oaLWR5TiD2e
dcoHnalFtOH+GgkcaHLi3PRcti9y0/ybNihgjCrgFOoEVicjthBE+2g7ftu3yNBkKEfyyP1+X3me
6qqneshG/7CujPfcBBahLaY8jNb0ZEcZrkOgYx6N19KpS++CDmWLLbRPOevmgXpYNsaZDr4YTNCk
7Z+/G9BA0AORCo1X/Hh4rBidCQSXqYY9SkQhPjUdCNyyDd+aubp3um7JCtI52alMBkhO/Zg87sGM
AA9bDywZxqFajjKcNuhHTY13cQ3cTA/7Zkw1cFPTyDm9dPJ/qT568VSGGFGlbIk/8yZEdy6prf7e
oq6B3HB6y/on0oEAevPBcr1FIzAg2Bi3ziGVXjGFjLDwGQJeJQe7DDR7PTbzU0Hk5HaykPEeo7kn
SkRf4IJti6vQok6+qswkzTfH9D4YqlcvfzNRbbvlsV2E3VF+9F/jscEgQoPZCdx5jh1MzG0Sn/ZM
7vDADRaNl0UTc1hab/TgamAAnmCiGjZQ5K91++5Ht7vHJbyqp/cmJ24QHOrpZfSwgp7j2yPEPHQt
1106AuZyWWBOtHY+DGjIrxkrXaGn81bzoCAnyZtu93xaTCuX3EbxxquOhpX4JLd8aSBqsMWnviU9
G4p+RAUkOI008aeuEQbu8EOiyB3UaHy8PQjGoqRk9akGQT19QQ9OouphXeUbPfLKZBP6kWt01Ugf
3RxrBcGG7e2u1RU+WmlLOgTlAQA5pJ2oSgb4s+ZtTIs7OomG2H3ArO1WHE9rh9P2DRiIqrRDAEcL
FXgSQAHfQOoZkJuiOdH3P0YqqvohfpY3lqer7wA/EoHfcVX0fCJxuEjZD8Hp3rQyX14t0RuLtFTd
Cb+FH3rXsG1l1Is5B55PDsryt7B5/fRlZTE0i2E2wXExS6ld9revojW2papCM9+oaaUxTlzBjrL/
ZKQHZoWSakm5ozyvJgSqlDAtYkOI2ijyunheecIE5WoUTfeHl4nXJh/Y2KEp5qkYEZa1u3ddCQcz
bw5nAIMpZncibyPJOtN30uVoh+zA/v46sxiUA2ju6DIguGOY5y4MHvsPCu7X7YF6b8UQYRW7HKCc
S8hfa7JZh4jpUM/Cia2qfPVP8B7OEtP8TFmNdigelHpTASQFDitRBRT7ekpbCaLtCg428lT66kMs
MK66iQBo6To1L+pTXKCuR7NRK14WkFunFt97czVq2uTK5G4JnXwUn+cNICgsRdHikkHyuAtgGKC2
gQxiURIAH/2MVOT1zakhSr+BwovQ28qfqguh4yPFLVG9DbfVTjiUmwbadOg15xLWHk6+0tAFbrT2
kEJrAr0skvHPRIsnm4oiesXTCzHq5xm0j8Yj1xcg13MZsXEfbbfnK/1BpuPIHLs9FYEp225whR8E
dVSZfGBh1cqzZ/dBWw2NPCEfly42tvLfg+KL/j3rPBLj6wQWRDVBYlsnL6F5N7zPKQ2899HY7ww9
AVZx/oFvyGyJnonC4ZNrRI7ND9qChEXOzS0KApfz3TAbHy82aErmcakUfJkDoBmupenEqaqqzP+y
GauZ7CCJ/4swZYpoBe+PAl5KaT02vXL6+pdDFifpCRCAZ8hEd+UkZL9j17z63QxzaXo0l/awn9i7
jhD+kcygg1SqtBVqO1xkVrWvq0ZLgt/K+HbJyz/ECtmnA+jyVNKzDriYqf62liie3Eadmjxan1UD
ExXiGbnt3KVqJv40YnW4QHxDzfR2EhS3e4bo/acfD1hMKs0zcNRBFxREDbXWDG5Q/IKqd/ptBE+H
6Hk0EnJoyhccXPIC3xCWp9SVQZOtC7ITRsOSZBz3ulIPOBYa8PJCAek7oNa5mbXtPNg7cKcyZ0UP
voghrY2JT+sYtvgybZHNJSlXZqF9rlPQhy2Va8alHJqRv3LA08vVaUeuP8AuCRRf4lEAP7dM0j/y
gJv0sLzd0XpU3Uwn87aRGn9Zn81uTrb0rpmanafaFiJqF9RM5rz1rVdOqEJs3EAkKVMIvxIReQLH
cxPLob2d3jzIwwJLtrBoo0JkFOfCMVDvidrw4xzTESXasFZvgRogoRtpjL/r74B0WgY12H7Z2R1q
vXVbnMYuPCZhoMUbIECrwDbn08L+7yyak6M6n7scaIs89AjxAJoeJZcqomDdYSBMCGmmVm6rIToz
KBb083uKA1VzIYTj3JnZqb5PILzH+sWLIkUjjptVAVa8+3lYlzrokvk4C8x9dR0xLYKvz9M/13Ea
Ra0zla0pS9XtIVHnIwS9xqcvOQNsXjkMiLhZ/idLH95bovucbI1g/XHokUWunBvjw+txo9UBX2N/
h7vJEYbXZhyIZeI6jEV+phGx1tgzVO/RMeD/FHBNJN4ZE4ja8YmlWU8YKpJW8c/oK9AcLPzbK64s
JurbrgXyoZNMLhdpXBTo+939/eWC7REjOku4JJQBJ7ThVQ5n9/q4J8pvXYlMTTqyoKFN3/mfgn6G
9ZxUa6qQldaufpmvx3XVfruM3iBBxkM3JKdVrIC6wgw63VmSQ1BLZOucs4nSY5EOSF4L6SZDUr5A
9auNeAv2X1PEMSSMOJV7x3BRFrpOoFOuH6HCCitk3lP1Qwn+WANZzQZxOhDUw5hSxoAlTrF8j3aw
XBsiF3uGsYukFklfYh1DWmIKe2rzkj77I+/0dUbpIfOrxVLDF+eyzSKNcoLeLrsKQAiTaeMhbqwx
8l5GMraFHRmd9eyA5X/63uzeRlHVK6CKRZAlzrDHfxh9EaZ64Sl1p4kMl9TOJOiCqYQooKLndNOX
4Tsj1sECWCmsuUNLs5gpukknLOw9b9umchtvOEk4BVNBY9uB69q0AdYOQeH0g0Ts54YVJ5xmCjuU
nQqYuLEo+tTEqJ953xLg7ukr/kEbmk4y4aSc8+zcSEtBOXjKtZGGBQw/a7a2PVeLm9tqY5xZPS1R
uda1UPRDgpMSVE1uu9GjTBMxnFvaoMBtD5+UHNJ+8tEU9GNTOPERuoc2OLIJDwFI7gebXWjw8BcV
Wte+weC38bfx2RUSOi4d74gNrowHU7YP5KDqpRwwdtwUOVJvB01nf+6eyVgjZBLyfSmx4mShu/fF
ZpHNapKNvUGmed0Zer7wd2XI/ANTsJLHuYgKPbFj/e6X68q/4tajRlwlrbnaIuXvyJ/cchfWk018
LSZ7/TWao2FNdReWjTs0PIcGE7CQhSoUDjdgPxL4n17h92kLrTFPNL7kAb0AqYDrBmyC184qLJKc
WcM0JwPGJ9IBSSH767I6X9YX+rCBFryyK2mcP96UblXei0+styl4tJwI64m1mdwB9S6Xsal/KvSl
tOxLp5ELUdSmJtDhElJWDnjPNBXG8fBEtTSA0Mlqv3j4tDUP5jw8pVSkJ9XAzb4COHeTuM4UIAaM
VRXT0ZyVRD+ntux+Nc7c33a1GyzObdxaJLGmYLjGRY7zehSIYS/fei5y8KUIBbvCCQQZzv0vUksA
OdOHbTeahqUUAxsvk+yBs3yqtmcnG0XGUzn4PSO6ROJGM+SHpV82m/FA12TrqTKqrjBcExOrh2cM
N5y6E3Q5CFNjjVel4Yop4JS77i5HzstHANWAq1Xj61BdnqD8Jr7mgQWlOtWc2K80LLRgKk4+jMIB
AjcLUNKgtAeXl/m1XSqXox4RF/tWPO2vqX2QauIINYGVNIcTGRDbO7zWF1jI34PCBpVjmwuzaJ1Q
0AJ+/d3eBC2R+rTy5IivRAbRyfkOLf3KV4UesZithW+gWuWoWrT9uY/oGeDQzvFDKIuoxYJ+2/10
ry60OWHrKHpqBkjiP+hkDByUJEuN1kJd9UMA5onj8D5fIW+HBBCN4n2m36F+XFxT66cqb93rHxgH
RPBvIbvLyKWJzue3ahmUhrUb6HTJKNbDk3FkzspDcqqsZPZq/uyqua81AxardYHx7nq6JRGyetH/
o66/J+8mEvStUrxdet35oSav9N6ET20n1qVKWNzKcWY18Pi9pbRqMAzvRLug/KvdVNxIrOqBp7gV
CANlE+lNA0sDbzqFJcRvW0CR236BnMa1+JW6MjI8+cTnNKJjIcq/ca50oplzeQFVdw40DWTmxNGp
JSvIwKX6jmDJWogtyyrBnnrk2vRj1L4BVT0reduUgwZPqaM1ewq4X7itBEaysvSsB0bX66apRTF4
VW8g4P+A1GaBljZTKtJZHxlPjsW2mDMjxpTrmKdUdSdryjJ8Svt78kb2oa9qnaDiHTltazetxrzj
eecS1vHJgoRkHOsSF4k6YJ0ek6g5QQRBWnbxjdjXljTCV42suOOAM/e5CSC4Qd72yuc2Qs4Ijppl
ZbFpKCe0Q5KUC0SwoZQzQylu6Hk9fjUpsLaA/p0DT/8BVODla5Vcj0b13gukUJBWbbIqt6jZoFCN
wu43+7f6iYcHmmzcTEYwoCnsxjG87XodkerF6Kfmhw7EHg3Jqs+g9L0ApJ9HJxUsAiOHqEGFI2ma
O7ClFH3Jr40vDKheF/2DJJxCEbgHe4lm7H6OEhS9166IlMj7KDr8EPtbLLYWmRob+VRDAweSaqyk
CP1LEZG3ZM0RMwgOW3PBgRSXP9DzEpjIXnBnelDw6NSEbeA3ansR+42ttsvtj0AvTsMPPGUWFrsi
3O+bz+aC6AHXUa5EhAJXL0QoMg4Xv03cVzwz5L8MTpnzh4QcCmHFbOmMrXJTmEG0wDw72R/fpbWt
vmBpe58Sud1pZORfdXqAuIfXF7lTCIUHzDU2aizltNn4ZShR7PdxA5FQ3KxX/4863Gz9EkKwdyoX
J5SW+smyEbaAu3+/slcz3aC0oxhTGbOkm9qPZJFXdfoTtdvXTn6W6rrh/ZH2vLr1he6gh0bDN3o8
RYehJgGKDB0SNRbVxiLSa3mzlF3HPtlNE1M/caDe9h9a+XtieS1jdiYq2gQjNL+2PcbfWhXQeCPD
s5s1xq2nQjS6xE9rurZdjlHbmYDacWm3on1l+Z6XcQ2Iv+ZYWJmekdXLZBC04ju0EE8zTVwCC9nY
X91RVOhgJ+dRNqXRRaxxpj8bYC8Gw2cOflpWgsW8fqTUy/hlIxKbO3qLREyNVzNIUU5hgE0jVBuB
QV3eqqEAFpQxoUSLQkWYJuEFgusQZ/v644JmA5KNtp0hGvP/aw3vK+TULZGmNAkkURbP7T8H+9du
A4BVLFBv9lQ2S1bWAoPrZzQpcqARdAK8El/tqRdB+yohsW8pO9KDRfKJoKHkMI29s8aesJBgNoJL
Ib8qGGXfRoJDb5uNddVF5NhqrmVmsCHwVARgIY2xQ9kxETMh5Bj9Z8h6KWOE8bZiW0rPggeLsLMK
Ev+JPR4lvmr2CkurlxbWmJUw4xE7RJ5qnSt4PxPUUdSMJQgoCRRXxHS+sf6F/sSWP2wuuz4WrQ2L
gRo7aIs3ckn+/AwT1zLSjH4feGUuoALuwimR/3UPIL0D0VF7XnogR2cb36BKsQfAD+DHnbinAmPx
fB9IC4LaJt36r8sGgjaliNZqU4CJ3ZXY+TSuoBxjGNZWSVbTDPLZFOPKrMbWPOuITGnre8468plS
YdVolwGA+ZeZf6JGos4+qrBnV7NBKMWnvTzgZWGoUe7Qxy2SmMwEiib+ArZtldTKzJ8nCDwLQ+nK
1lDgQefsFpWn+oE1IMJ9zj3oimxMBIWuMaBtlD97jTRg7TVCX4RLR+hENNm+8cKf+TGFrXEvX9eM
eQiQfbwb9/2JPj89FvUtYbbigavWu/gE1qakTcKFj6KFiAAmvh3uaaS+wLOy6oPn3s1IlPdCI5b5
3qYhXrzk4wZ06JX2RyKtJu0ex5S4Kd5ZgfriFduO97cnKDSA/shlCl0gCTyks6PBjOG5zycxitVb
olBUP1cuBFKwwoLcsXLC4rJU0+IqeX9GpD18mx/2uhT3Y88ie6GLhcnofXZ3S2lV7TJG1nsrsqtQ
VwqHE0gtU+shj6I13rb2GDyYXmWCHtjeadnrqVRB43zFJ1bkqpJM7yvs2L5rZ3l/PzG39hAEXMpx
dbYfJkDLcoyj1Sxnb1Ra3GQJDaxMYBKgdonWVeURrSS5hgEOnFyNyErrEaGUv78a5M39cTeeanbh
whF4dYvfKLddHzQn6R15eXP5GA4HHkfF4uW9nuEbtV/PxdtTPAOYynwr3/gS4Ws++RwSQQ/LAY9O
xgizpHOpz1fOTOF5zSD/foc/itdkJhfpqNCG6r+3ROfDkcXN1WgUyRwlScx8ZER29WwDmtYPiDJk
wTWZxF4dxgBVjgjBwvTedhqjVh24+aRe30zXzPZPsSbZl/uaMCALCtW1oOPxFfU/ONq2PBnc+iqa
rwER1tvet+gl5G1kkj+hspE9ItNuiHsx8kuGeAHvRe1UFs/YGWKFTWB61w4+Lqq38w8GNegp2RkY
GDFDN3dfJHJg5AXbpB8AUKywXHH5GtaMScAX6NuwC+ZOgBi4V5+L9e7ZkEo/Tp3yJVAzvTCZlNfs
QRftdAvC4uwN+bS3fp+i6j3yrIPlcQmvVqa9lmAAW5+Hm+rEuXjpQ9H5q0R4IuugpgZQvWakPbca
2kAUGj2n4NayNFeDGDe4ymof9bq3nU3+Dutl2/KSNPgmhUrOKuwk620Ae8DNwTq/PILvND7GXT3/
dOyiI1E7r3DxYCX5/PyPVDEXTnBzQEXxIAxv91vsFaOQ6e2D9AZnNeoxHIe9xsLt2ZxabICpeRTw
0iQGUsAwFJzVkgc+yfW/7UXYR5gvBGwS320rIqARjBRZIOWL1l0CdGUBmG5uXyiqlcSTCVlihi6w
E+i8HLoWGrnL0UopsW2A4flZfT8BMnqfrDe35fWrqhkN9RERixBNAPPZUKhvc8osdHbZJpPZwVco
39IBQT21PlT5Tk4rtw69FVn79gzbU4uIG4mllhvc1fuzXhMNmn9y+hoQYp8pKSU0zkxIXs2XyLdg
ce/tbDYtpi+KlixBwRTPUJzny9Oarph+f6JbTGaAe4I3vy6VtKvjnEDVLcvpR33f97zburZP8n4w
EicwN+vtmSItCSCujne5ORkoVZzwMgOHFR6PVugd1u5t/sJeEB7M/Z2yUWGfpiVTTnm/JJDQNW25
TY3t3YKvoxclKNb0803Iqey7ZSeZD1+TUKzh7dSY4ZzmUWYeakcT7ApjGl7rzSOcwADJv7RxlRcR
t95u/1PyX8Jva1FkuUS+Rxx5vhmUrYNIqszGIMiq7D9oeT9ZcKfopqY7u3lyalFO8goj2Gikn6V2
DsrjVku/4YEfrwtqSH89LIVs+5Cmi0Kw2/FA2NDVlVxdZlF9aPItoKv3Gfx/MIvC2K3xh52JBxxO
wro7l3avWkMbd9LAiArpBWVBqiJcE6F7BlXdTACvoGfNsZ60KQGc3w27TGkatBRD2CXhpkZXG8wn
QIN1/ehW/J8vAwdUGdRn/Q8yf5+cd4Jsncob6zLtK8wpWcYdIXnFswAv/xFZd2kehze2GkrddLbJ
gS6JOsewtTk5wowfxhMnGZIA9dh7tfdgYkq3DZLRlevsFGmcVH5PzR4a9kNrsMX2mmewXv6j0hGk
AkIqRZxHKGiYC7Jx3pYMUgNZS/LUUvuYI26qdMeUZpS+1RfENnjBNv1cqrHpKTbue5ynR8i96HkR
oHkUrSQSiFE3/C0wNc8LMUFPOzeYphjIrEHuDf921ASF99dhCgLn6k3gSW6JWWGIisebS5aBb2l3
Fx0+eSd6CfQBQB7vl4uiwxSQ1K8OZBTEa1SEIfN8aji9TeknkKpGiwkdQTbM9E5Cv7pz9UddUujz
DBUHZPhNm0zc6d8ULgzKVDZF2a1WO3q3LVWOS01jWSGK1M6vUzN88eXSG62Cc/q8s6gKGb3mDzG9
2FePrljBoYqtYQvkkfE+n93bjYD2zcgpkxUomeyLQ3zW2TjIg/abPGBWH/mmSWC/adoPBcBX9yeA
vCP1JY/ZnRnCUG5hfIVv5uiwnjNDU/FyPc58fwVNfZnbslmIzlOaPOSwl5aHyW7zAG082KDgdPH6
mV67k16KGrow2q+BKFwfm6kNLL6V84v6mc/tJ7auSVGVKCOSsZDyAvHIOjGbqZ5rrZiN0Kw7KCCW
5TWw9pbCvEa3QoTQ1qP7KanO1wDJGnJjQcvLe48T3ybG6B+Vit7yr5EHhXMR1C255Ztruk0hul4f
hp/wlIIXxZJWmGfBMaQzNn2vd9WFB96C250K0BIedBdVSDQbZJqb+1ejMnMgfsvFpPcr7e1Zj0cx
OqNQceC2N87hZKDuHR5QLmFqO4XdiclS/bI4Yt5h45c+Bh8TGP4COPL4R5xoy/RH99+TnkFq1E7P
Olc+55uyhccISrP0P+wJzKDjnkRdlwYcK7mLhZzNnaTH+UeOw6vKe7NQx7cmMhjgYXvfH5AP027K
X9jfKPrcCz/vKxZcg509ewgwZH0rQYxsRrSCXvlG2Pv3PqU6xQxx2ymfBNxzMNNNb94tuV26EGGw
9ZD1rMNnJGBVU9fLWxEgLYbPumtgY/YLG9lALsEmTjq5IMoJ3xz0NTxSlqj0JcFDcnyAIlNhMXEd
8AYbzOX1S8DMntYbglWib7JxSVzVteXEKiXQcQaGDYj8tR2ZZUUJ5A4jXbsT72AKVkIPLILz0KpE
pmgyBVqRNtQmKAJFbqH5w+Ru/hliEGiMM7bpaR+d+NPDbVe7J0f6AeShj5B9W2iIgq379AGSHzCr
cCGDPe2NPOlFF+Zj/ABDVTEy0HvvoVTBsUw5LKlezfhDPzJrcU0vSV6wusWj6tuJsnoGxnxbkvuU
JEXfWsrqKYpIfUfbzOwjwBzu+fEfYw9LnqHZS1OyrPeWwrzS9bL4IcblveKiZ1RllIwFSfZFxg14
cQwDYoyMJK7gQAxF3HtaMuVFpbOhzXAHJzqoksyqf84JN/AEeQwmdmuxd+WhtJ8ZPkssswAdxxpk
oAAJm6hhr0OTwYImKV4hXjBPKU3Z3MMAtvC6tD/DiksaKm4GnMLyZX2prXY7wX20gu5ph6sZOrGc
Tfi9pRg8YBOKJ+iK6teD/bnsSR5ap4Ysfy2AWoIJG+vxaawgNPfOUnzUTUjSum8oAAX7g0ravurl
eLho5xlzGRFiKbT8BDeG4Br6G3rN4sIQ7iRzz32voTlSocqqQAFjIauyAdk1KI9cfbzohCg3xYec
ceX2kJlPlRVAP3SaELAmOfpUp2EKMbKndWpXUawe8UXJFpvHEiF14jF7Lk9PVxkw5C3HoPA264FR
JBaUCmu7QXlsSw0hudIynnyue0rwWu4DXS6VuYzVCjYqJnG39PnBiV8YXl6C68V2aDAPbivkcMrq
YFfDcAWMDiNBEE0EPGptUS+KEFiCbRysXjQh4h+nItGsdTXdYj4VDKmt17S0cwLh58h3xKUcFEp4
6nRzNnFiJLRuKizljzrm7jwk6ragS0aejlqIlRBvmiQ2W0TuFt9QXYSnqnGpjkgetWSnUM9/0GtH
rNQUERwlj3Q9+/2ZDavS/j0bkS0nIt+rQAUUTukrHq6/3rIBWcxBEoq3oxjurlcVOAzlwlQRCvFH
1/g5s9Hc5INuyhI6uAwR4HR2tEj+oAqdWvvmj2tWxBxX4dmGkQ8nO2/eWf4tViDawK2om36OWvVb
EHfkVM6yPj9o+p7N5ctAUWz+e26JDSjVdx13p1TUeiNtFk0XO923BymduWso7u51nAzaYpT9QOWq
FWgd3ClTykv3lUEW4LrYvTvuTq00f9xFxNlGp2/W5fxMHwYououNKxvtsynE3dOSPpQ/na0C4qDy
i+abJuXi1/lsvENID99K6HHE3ZL3sUm5X02tUoGRwIY3oOj9FZK74+WCikpV/ShcWbdlBEcJ43RB
WGsJCOwXkjV0nmarKnPSnXHiwwBqRuwPj+T/lD3USfCe/DPz9OvIHgrpweIB6DtPRt17KOclXMm8
VPmWBwmVe8c/i8AsdzPwgpZkq4v7u2FbW7CsoeGZ9wwvfAITOgfYW+oTvcNThvx7eZPMisyRGXI2
LyS77iFx4lyrnzVfzr1Pkbf37d116RgIHt3MFAnoPsJUxglovSlSSZVYq9/t33xlCqYajevupP+a
rIGcy1xgZyIo3RDvVbXiFEt0Op3E33CBlfl2LmmU+i8gtJ1EzUXg8CwAKQ/C1MImhYDtqxu0Jzpy
7ANsKOYKWGm3qPnmjDgKV6Y/vbuP/TZHUP/LYj468bRk7O9k/S772UlFluUzVrGoIYMVFsrK7EVP
orSY0EdF52tOMMqpG61Dr5nN/F44UX0I8sE9ldfUGQfep/qSeeqHfIYs8HfKXxxuNZuaW7fExnhv
86yTf8+7CpNLoM7Xt7/4tSvVzaliBvFylJCEHHkml1BpbxKXnJFPp8JIdU4Li6QDN6+nXHNBtpQn
c2afpRMkN9aU/oPKlpiBfoV/5d6vWcgvymlLpsQ3JLz2brtPfDsQzuMB8OcNMaFgr6HxneVzpdGw
IkcyjDaWIm2Ot5/Gy34NQ/svb9OxctdmPEW6ng1+mVZWfOv/Y5rAcdHHSu4fhK0ZT9iW1yGRXnSg
RXonmriqjtQ5jEt7hSQ/7oleo+XchS24ff32KfacTlAzrF20nCbPOZZ2UR6eaGIrFeh4MU9Bl05t
0ZgOCzSQfH0whWKOc6bZEooY36MZO86CHGJRzVxgw9WYm0PMP473Ij8MwLUqmPVwksiG/4uPYr8O
UFb0EOGsJH76Je+PoXHMhr+NbLS0Paf9+ECFjFrFiczBjFc/80UF0wk7aBdOnm8pxB4g9l2T+3nu
fXnvwHFjvu1xMupf0AK9tqeS7iGmXog5KN0QwXkBHbJV/XT8Q26n8VQirDwXfvBOLHuscS/2c9YS
vHoIvuTLk9PxkrIu9P++esWitGPNOnCp9Q51+QVtwQf7E+dW2qogHdQICTyT9a2etKdh2lkPC7Kk
fTFOxpX5DmPiFIszsca+JJmPCjWdjfclGsV31nEaLaJMwnywnnGtQ+cBiLC/uxXHxD0Uhu8sUgbe
hw9OsO3fFy2HjuyfZcYGRDd0DzpCe+/PItx1SZMuUym7YkcL+hxjqtQN447v+pNM2ep626CFQquv
naJj1J6PClycviMnTu9mmxKCThSYCR5raKnmMb45GCMsX+1mE1hjsJCaB4kqrBmvU8M79OeBgc+x
Y90p/FpXmjDiF9+Ul/ZCxiS+0x/1HhVFioQpyO+WYAn85WbRliTSSUzHULkHOulFe3B3AyGgfXd8
3U4L94ROr7sOBlWZNEHppTXi+CdpT+NXXv2Q5PrwgrsSq/Q5ztJWc+sYRZBnvw5AWfz340prDHsS
wHGONMJfbtT4Nmn/O/rbssEQepIiMjvRko9H1G89ye78hW/fpbZuhmda85TOMmEZb1PnUhDBKoY1
1BuvF9vCpExCoa3RhvjYAP1tRAaZo15Hk1kG+fTOXhWjFuNztnzDzA0wUA/Ef1sya4dL/0zldo5U
tRRco0PXmq97extwfreQWH1/7k9RPrRplDLQ3u79hQubl6+uRr+wrUuuJ4uyIeqqX5Mh/FgHtXUK
Sc+wt8K+mUKgLSu/C+UjRYLFuhBG/yyjaz2tSYIrRGVUGrch7ljxBM2atflsXZhXSNS7F2C23VP2
zuX9rJKthPRO1cWLSjjczktW5oooOGEVPFvBCsfbZXIeWkSNqbgCvzd50ym3LbB3sOBu1cxu26dl
llby9oZQmIOchqVfh9+S/8+g69ERdpFKxuki4FsSOfRBB6x3Pnq8LzD6IG0USL2bHcU8FhEgzidG
7pAbndLQWbMgRsT4FkoZBDDexNDfF5SctrntBVfra2uyWVdRdMeC873aIejaH/GgYefO+vxC7iwf
SVxyohZ1HftttUgxAtag0qFkYrkbsj5qusBRQ8xNvi5oAHomNfpHNrnLeQ1bIbYc0oaUmTJnwrbV
lH2yM02rJSkRj6gVbt0IkThRyIzwf7Pyt6I4E9pKQh9bNVNmNOol8C3pQOm3u4j7XcP2ywsiD0LB
ym4JEU/bUZmwwoyvKm9MNI3g1aQq/WxNkDxBLeQKju4KAM6zmuHxKwAxbigyiH3ae0gtt1k9rP44
OY1O5ayoQnB0Uzg8xw/q1+AFxsAj0datbGZLfq8WM6s7T08e0WiHj3Dm5uxWvjjmfjeJ/sszqAJ0
OazwWmqUs+BC2gxJzvCg3mj6t1WxmajVjiDZYSEEW4Dx2EH0nK4XWrjABebhZcXAkNp+HkuX7DIm
OStGcS4zVEiUUkoVDKI+LCvgc6Mik0o0ls3Neh/y4c3jY+BhXCrdb5IO/Mwvn9BynrqNYkpi5wEp
L6/8wEeqn9aJDrsZPOjBrEI+u6uUVahN76OpFmO3ViR9L7LS2TaHzLItF97odLorDGoNa1mMwcLG
JDAxRnr9e/uSLE7aNzae0dZ9R+Kclfa7v1Y8M93l5uluBXL0eMMPphdkZ3Cus9WkRSeLmdCdcfMH
Q9MGQoBhBQrPfsh/q36bIcOvWjpNrqX3XYWZUMtGKNYQuNKp+veHoUhcNHNlDjvtIP7FOaj55cuA
eNr7SyZ2tSdRt0FW+yfDHLBsWGUaoqZBquSng46yeDYkcKz+XwP0c6bLAiPU1I/jJWFr4h6x3SXm
g365GpO8OZFK0jz6qkaot9BZKV7Wc3+aQ4pa2/E2gJkPDX3mKPeqUQzuThz1aYtlW4lzhkuW6yHa
yhDH0XVKw3chhCv7+TUptHbn4hRHCr9XPGmFuPF+CsXsiTyytXZiyiLhDEwIMURag6miJZyJl4+f
X6m7VLVxU2KLFZffmS53djsI7FdeMt5VEAYoHm5bJs8YzomgMayEknzcSizFXtWf8MX6kk3VxhlW
nCAfu7n5lcLdyoDTUlvenA8KXQ1lS2hLSAjpJB16oa4MUahAft3A6YDLNVNuvNFriZmfZD3pt7NG
YT5qPdYBREHGIN5crFuw/rh011atk1b9rGxfPxw770l33N7KoYHtnLRBgsH0oN/bkldzkD1bjLqZ
66cX4lWjFryQuGqICcyWSgMyLSaNPD+kooXwreg4cYxfKVaWFyttb6xdrgwCSCWmBRAk51W1O4zR
20O6TOTq/mjynl49licSOplA9NT6yB52wSFFZ7U6JiO46hTpQfNYUHMLv4ezADsOel0/w2pkNIeZ
qHK/WJZNJhXYaLEaFhR8JNQnFFXvMZkUOfDhtUnImA+lXJzYD5HDCRgt6vGVE+dH05/bOZj3LIqN
W1bhU/G/cf3cJ2jg9AHb0Py/Fe5kzC9V3xMIzFDuerDyL+kRq1iNAlKkaONg9+mfIZKNWUPUex9p
7EUMhXdMvAFW6bv5RpD6F87FBZ1F3CqlfCrDsY+mO+5HF0Dvi3H+7q36e08Zt/kIafm0VOYHlgd7
GIpVUjn0I2lf16RMoMN3wvfUdUg8/6KRaHV9JRcEJO/nEoiqGZPMyTLKxp9GD9ACqh0DP+nSi3Pe
kOle1YwcsHgtt1Pcf6rUlpjDvjofxWP6p3LSkFJDttyiTygkqUKkUbrYOJOHFUKhsuUQ7PhI37A1
pQ5ImJDs2on0f7GnDSZcNK5BEl+fROHLJzmFE9d1XrcPNG9plo9XXNRfnlrv0EKKdgCn/vMz0CcY
jC0gF0HrkHtCllT+DZEyes1hsHVxrPwagcKJoAKoOKZS/aYSqr69tn+yPI4R9BmnUiat0CStdgs1
BaI5T/hZ3R2au6n68p0GdAfKEzhAFpD86S3GCH/xEfCPYT00O7LYmpjkHkTqRWyiLj5YUtHMz5G5
0Wmhq5Yj4U+9CFe5/pD61+Ne1rddj/WpAGZwnMEib5KBHxcXd81vs/hxQy9bkjOQpeFUmBxO+XC0
JetTVwkIehWJwmwTSnEfnz+f731D/xXllCQqxrJGqmSxnMxNQGm+MB1DE/ekaW8yL/G+DUFdvImR
okoFxMfgdhC5SzB4/3PCFYC9hBrnDoyb2R5UPYXW1KMkF83Sfi7VVZDocbK2f8tD2WuvLhAcUnaf
qYZJmCiwT3Dnm7a5m7h6Xw2FFwLXwqR6flHfr0ChWzgg2ikdff+LK5RPgcAfF2dgK0mpW6D+nmue
fnKYmwvyIL7h5iUks+Z4EfZdEAlgmyaBBVCE1KPN5mSo70yNuGqvo333M25Frm9SV5fqu3kSOOms
4eWH53BB3FmzprmUkzwBr+izrnEIoGA2+Fo6XSGOTtlGgTiE27sLTojpBeceGDSntoMCBRYNA+NY
kb8pVbwL+73ZXIiMI8Z0uBhcyBc8bem3vwZvwZ46Imff+jIIBkp3+8jTvD95I/lzsxxIjf7VYMbY
uajSXr38hoKZ54RnwYNHOlO8ly3wlK8maWI249Yup2luumZ1qvxFOJFuaSOz48L4dypejyhbOTM7
LCKEHyuYGweaHfNfJnMi9RE8MXlfQpJGirKAuL7EqCLDlibGdpgj+qnxa++7jGB6JYWYNzWkCgw5
M+uHA5waXFtn8vXCSiYF8kym2HqsNBpQQVKKZMf97dhwwFr1uCA6InhNOjGuFI0mpb/kr2yBCUTU
1OW5zuI1ZegiIghhQ+NVtnIvZhDreit7U7rxKpBGyLlE+pTLvbrZxUPqnW8vZXuXEWLMOexoWsgM
gSLOP/Y6+fPfarYtFzFcmqvEi6Gof2ZUxUNz6dKtRqYKKVlLohRJPdvuBkUBZDcMZSebEi2w1Cn2
k2ule5XPOi9wgqbtH06DjtSssA7quSjbrSlpPZh8yXxie+lvaWcWF2nUPDlAa11upDjMlFQXQhBY
OfMwo31q4ljasXtxZ77di3u7txoX5yItCkW/vkJeOb/FgNHtfLBSVl4yJKiIC/HuO87b/Uvw4Fcx
cs9QnHOIt9a9AQQ/xBfMpUNo61s4h3d7eXw1vg+Rk1Qn2MopdcFYHCcsBXpAXL++if3icaYbKS0u
qPz8kAjzk6L6P3/SKdlirAc9XYPgwRuf4ZIrLwiB0SgxsJJ2JC2IL/YMcprctoA0PEFPMPRu6Z8A
LnyW64N5J5RbHe5RN9hcKD1sic28Y1Cy59eV1kTjb3qbi/6BeR9YtAZGSoIiNOIQAdWbzEYBM3e6
XptTBoQ0ZCyn7wbBpBIgsnUVMr+VPWMQJwk5xdZvsuH6v3OMKZ9s/LKiOUaCwSuwcAW1az7SKyTO
3p2DoavLYWQCgbCjke6yWB7YwuRQF7cWZGA6sg93gh+giTe2tIL0Ka5h9kyfnX4QQVJs0FfRdLLE
7S85LYG2bK4koFXm1TEgFvgU29Z7ZicyiO4zovC05pWI5XAZjcZjS9PicqYPbjTYDelO+kWtNnNJ
ia9LL0jSeBiDe18z8j5EmTozn7cFQA3kZTwsgDMHs2RYzKjD8iOEKvxsth3afizW7bYHo6HwHbqm
0Pac8TVF6SzDUsIUAe/C8y9peg5YNoG0bFw6c6VGnZ1+pcbhMtv+eoR1EusW5CRo2WB8C4N3jpZm
b+x4VLinMm/4Qq4enEgvnc/YjgsbT6Pn3thP7vx7yO1itKrhwpsz7YCHNCCXgw45G9RihGmaNYOp
9SRYzgGYerFuhzNkaDHQ39yvwVV3w2kcvc6ZaoKPAiDFjzkbQy2d91bnqOHmRv0ftS40M6V3uzxg
vpBaghYyhpuCAYg0dvs3Auyn5L+zjdC7RDieZI8tdQ+1b/U9HDb2QG8NeBCHtuVZMCKme9OJZ6rg
xPxqp33wzZJTF6IEBSAamx8NVXUxbS8uZ8GTtDC85bWKgmCndvhmL0h6UOQgcO6OylDOubvcAS14
1GgkZoh2eSIbq1G3634PfZWp+zv0Ze4MB+kT6jVwaunVE1thTvIWdDHS7lDgRYhjSzkQAzNthYMw
6cqsr76CRTN9Gct+sFLZlEn6B+3Ht4fIM5eOLTuL/jfsB5gfHDV4gxK5+plemx6phUJVMnxNKcS2
e6hNemjS92jclcYC/1qepwY7pQq7ygXzRwiLW4/3nNOlFJhowffiepb4vyKbt7P2Ziw6cuMTDARB
S+06YFBzlaN4OamEY8DPLpIcI6cJ8PEY9mSNScS1FfTL7lLjNPzeAV3LWaaU4hg+olPu0chDRZpC
XgP2u1MP7Uy0g6ID6/EtDtzG67G6NluO1ovA1DQUnIA56TaElDJfHJQlZ4psF+fx0gIodnxgn6JA
ELPlDdgYY+by+HjzrtLH0a0T/T46kgHFqj7zpXaZCOmYy7Hn1n1IFU3iYdVaQTvpK3aEdEHrLxCC
jJsH/nx6XaNMEde/x8lynBgi6lgAPPgAU6wtAIMUvN3ejKyowmEWeLf8Zd1HeTRp9gKLepxeOf6L
yc62ocPg74DrE5TiBpYi8r3p65WhwfAdyh7Sk1heUmnVdpCqbS9zkEN2A2wpxLPCaJDWX50Zpmef
mE0phwbMP4FYipSt+rtvAvv036j8GXFF06K1dZTJdXjwAivLKgVIW1V/ZyBFg2QBRpIP/iMUEUec
XB/eS3x8d/bzO6+oFlq93RgnE0OG0/ZPg0Rp39Foyxwkahi9aNjxaK+0lUL1zVvIiSrmj8AaMEGp
wpYpZOyuQslPYVv5VoXU6UcqczkPnzVOxyk4H/xNI8bNk89T8SauBNMxFLewMX2fwMuoooSTDaIX
mWaaFA6DRgdzUk/rXcz15G16u1Doo9n5wE9EezAnbwhDTiQFCvHMsYRclNaXf8REwrK/aRY6y4yI
tvDQBmFg/4MmMDwJoj9XLeJlZi5ycc5tpFbeHlwLWtzY2+LQKrwoHMpmkJFtRtVVpEJO8WSVzcMX
TSge6hMtSUjFozG/D601SoRgliiaAeYJbjdfQD55VqpGOE50sJ1QdOJiLGErAwbBlWlEJEugj6My
axFfd1czBp6UU/UKRE3Gny4I1ExAJ1ylSeoYYM+28N5G/CwpW9mfoD+hVsQ0iYpHldngHAxc0shV
VkLQE3IDkcndNEmIQsMJuQuj3K/W4hSBtNgxGI7ol2w8/5imLXEOfxGG5vBlCJ9xZmvwSN/QtdUq
mtODF4HNAxRD/Q9Hw/ZmDCpZYn+YFrrzhLHANXOt62cbii8QvKuPxhdWAE7ABaHNZbIbFjI+j3L1
v2AN/T4ypO7KR57nPh4Ypr+ogtpw+QlTnqFxFO8IAe4C6peYsO8AqluRo/5nhjVakuB40hsPfXgd
Bl2olTEvYN8HCTqjK1UMVwQIwqYBxS5lm/vzZUiXWtufHq0uUzlIyAYZc4tEbeYnOgWHTTJ/mPEk
7wvmYVxPnXQNtTAVA0gSm7hG+s1CpqDmhrwRFnlA0TG1yTU3Kc0SMIMVyHC5wu38zazeiJjZEh2M
KDJj64F9hKCq5VTo29JuejfyogaaQVnBh2V2CNWpqjAU65tbmlyPg5AF1W/c4Rd/0rYDh/9X5J6K
K30hJxDRpAMVzvtcV+CV8klc0x3/z8fqYOciJxWA2OfR3fRWbn+DqjKq6T44+niguCKbEN0MCmJP
7JpFXmNztDWCiOWWq+3AO75aYM0uMI2tIIdEumRKszvQaC5RrrGYRdOYdkbMPFUCl0wzAcvpM+42
yEDMstdWwjNjEew6OyaTthLxNFHLbLl0sSsb26e2yWBa5DtGSsudcEK7uMVvLYZYUbwgrIeC6lfS
bC92Z8p27B7RQR0NH+hZ9mq30mAFdodfRHTm7VxsV+E2i7MQ4xmDP2DeGyYqvzdjfoBPdPLvmX75
xYXTFk0aDWLwl1aHMygwAkxYlbfAQx9gHrV8aVPl2zcuAszEJ0Tg7z+/zRIK7wnKCJQ3FYAS9t8p
64dt9xG5hfuB9G7MIarHmf720ZkYj01WejHblRXohjf8unokplZznbjbVwQhzCKCBLROVkJhpat9
rXprhZqpnyTd9Zpd5WTjQTZCLk0OR9eqGa0MdlYWAJ8/+JceZIiOW/z5TJw5ykZc9cIJeACaZMvE
gpEtkX1gWSkxxJ0NudgXcDpEseNDRhuIo2cq7y6kDUtWekaW/LUu/CME91pJMj4DoIxXUvW9SY+O
ZieSezg30kpc4wWMWIrm/bKdmQX1C+022ZjhafqTVxFZEj5EbKcXONr8ePtRy7tPVVEQZqUNGjnS
P0366b772O+QMBPQ02X3fm1Z+J3Dht8rK3TuNat/Az4VuGw9hHsxljaLng9pzGKKRR+GTNpZCRUE
HQeUqB8qfkFkD4bxGn2REEKG8Vs+Gq+uchRg+AEix8PRIPUzOVFW2t/yP0RYgOt0Q23rCcXRb+0b
lJ03yMZqgBb6sg1Y+7qrNld/Yn4Y9KnLGo1ap0PFFZr4NETpoiZp2gkFQoKQbmrej3Q4m9t5+DNw
Bffic7wzJeXdx2NiAKPipXRxQAPtVzVaxsOTqsHpc0W7d1KWa43Mgxt7Fle/PUXY85629MPHlrth
ER5uqseTKlvm2WV472mkAEE2+HLF/nOtUUaTpZbuhW9TAZ6S76VM9evSQ16V0w6vYqBsfRcMS/fu
cBXOqYO5yA7RvfoFUfD8P+I5hAYZXVF/ROCXHBFv1+vPonyo24+LiC+35mrCtryDg8ucl379dKsV
OL2gCug06Rkp7G0Nmi9vnbp7Iq7kVqxBSQuh5LMpwj9seAxw1LAO/IXtfWy8Bo/O6vMioGFv+xFU
8EDg9HV6jVl++genuVEa/S1NEuqIp7SNi+6KeYyYJV/lrGWC64lEASr1lg8qw3adUpNcoGTDa2DH
LtskwuOmNwJRhVYrHkJ6P7X8XTlMQaLjbQnDpAruxWwBj8t54aiYG6Ou6gx4YJ/nl6Iq1TBuz7Sy
pZdOMAIhLraKa0wqVARU8zW0FUOKNzte7wJL0jsOfb6Wy+3ausL7TxzCuo7b1i1viOq9ZE8BABU/
qUVMcCvp5xXKG55T7mS8EjGmh/MFBVHN/ceXZwLtKhdzl4QF3eRu3ajjuPq7KBzJK0rFFoOrWc+o
qloGKX/HjPRClIOYI0AEUyrl2bMgprqElozcBmSZmPmq8CE/WOt2wmhI4TuYsgM+U0xsSFioRc5y
aMBb64oxm81cAdLISd6mZGmgTbogMS1Zheu1MMzjgYpGLsECBw/u0O/GTTvm+pjkZFEs1IPLr6WS
wf0ciZtQ0zcGeeiLT4/SJLnPxdjeZF3URt5YQtRvMrn/Acy86jmeOTr3OIwMerVq0a0swhbZLpI3
QP3yLjHB6X9sv1LKkyp/CS6j8VS0PIbx9VHf06cEQcwvWEtNeICOAc3h1WiA2WBlj1Jf6tRMUhzV
MY1HzWmwHqIbwta67GIeLwM5mxYGDaQdH61MQR07oiMKAlDu2ZGi5RzRpabGzFu6Sb6a8oB7G5JW
U5xqBRFn3BxemZNCF6+nHy+T4CTM5az90yc7kDZmpN6LMKIFghRJ1YowhuFqZn32FaAFWfj2fk5G
ZQ1pe60hSa/ZHl9dyjqJDmJDt13XAq8nKl+oO+5is8qSTsrYc+Dd2ofYDegoyEca0mWFKCwKJyfq
ZvLpmzKNsUkl9IwAAMetZCSskjj1dkpglzCyISl64xioKtalPfGJl3tfdg+9V6N8pINvaZhKZaHb
rKfqjcQsZtLxoXd7XKZZ4qwVsBT7abMuhdA05pG7yL2WFSiGYjJNrMRY6FHCzpj+IovgLDxLbIs5
v/ZbW8+Em8e7a3N+eVdtY9JHGUEbWS8nLYewYEX3Bi9vwss61QeR+HwUAlALTdKCJgmXYvU/JFqw
HbFrITAp1rB8W3O74wwee7Zgxe0VntPd8U94sQxX2610wFqPW85KRdTBR/64WmBiEFUDJc0hfYse
sIUh5X3zui8L4RLy0r7Sl6q+dxX5y6eQaObRxqFGHAYrk9sQkJXj7sD6KqDsZBJSnDLVeh8zDk8A
fnhKVN+3TOLG7/GCWbOScKnU6VOU84zRL11WFvCwW141Su0HBRi6fJAZC0fExBvC/XwaR7CYP+Au
yD1+YxVvtghzdwwqL+jVb2HVNwJkTAIgiGoaBkMOIJQuxNCCGrN1zk36rSivzzGQT4RMv5YJK4Yq
O5r6WwWn5ypixMkooSADLvlh1HPUs/9ig7rHOZKqgF8vrs1Oo4rLPM/fdGcXYrSGxJoonvpbpztU
MOrR4iwo+sTNtrMBymWka8K7rgcT3pLDRD709m0FukM5HIseXbijd3Hh/0wBuVsUR+j9c/NBSW60
jDEyiQQq4YqqBucSw2BuIST3vYcFpL+X1TJgwiJQR6hKZE3cu7/9ZWYuDMCVgqER4DWhbVMygHDj
BvrahApFKmFOEeE+REFt2D9LUjeLLviBOJW2gkkVVVin/LwTAw5RApmUAe6vQRn7gE499P/1DvDa
QYZa4Rfj6NXwkBhjio4HBty1/afBcaxIiIRTtHyErEZIGXRQA4wE95RFyiEPEFvujzbE2dEk1CGg
Y6UKJBCvbN8aiOR0uw/tlc6bGee/VXNl06UGg4NqUm278ZSYImeQj7exrLD+VuZur+ZTfneFObgF
7qoNwwu76iVMia5iethxRJrF7Igh1A8LIYknFxm4ozEpssL9uN2UlL9sEmyRhz9nEii1EzheXN2e
iKc1/QUGDU4Gwl/gI1EMyi6Z/Q1MYI+AG/wTNAOlbqcLsex28I5oWM7bKSDzsJQmNa7ZOSbeaQ32
F3IqKNczT6JpWhovNSc/eabL0DGePRBMT3SUKh1CcazX757rV+BTCcU0i5lNTIRnFhIMqYdU3eRX
6kK6VIcILfU6ebdHTTZxWg+ibz9WilycyveUkIyQ8zDN4E/aJMqXCYOmPI7DU4ufI6dDWVbi+0jb
+otVfEIyqFtcNlCwUl8y8FwfteVNybs5NYNk0GzCUFPvV9MmN8qc0BqJEZnITcJinKk1Pblzen7P
2DHvwsUXBZcS6pOd2o9ow/1zlKhe5sgQbuSa054iStKdITAp9jggtbdKyYmnKajSOQLxBgVLn4vV
v1L79gWKPDKH4nfnGS8vdhJecuDFMgnZB0KYoncdxO6HDILGMmH+fHUi0bldARpZBeuTgR3L2CPL
OTtPTyRpJytYPBxXWpBf86VW80ZSf44mfQoPo0+C57itbRX0V57cR8lnP7xUwjs2HW+llaMhQmJA
aztnOVvUhf9usup41UFCOB3WzS6NB4WuqYASeKrD9tioXZ77QChM3Wj7vKZG0r982uSu0W/LL2RR
zX7EqG5vlxRRIyST1hKbAZO5m28rz02My+jTo05hhC2OeYfcutaO+lLlf8X7kMY0vdS+HZRV5hCz
XFfcQO8lq7RFCAumXFN/Uqx/ZASJea/bqK1iqnyBMZJ12+IY9qw6QHZyd+bFQrqN84ZqYmm8pL/c
mPpwViV+liWl3nLVx6Yj7FS6/AjqleLlbZWCU9aj0p+YAqsPnIfHbG+qahKWfIQzxmd/eUDjvMBy
1UFWXqncklfJwxKQU2gEjDfPugvRYuT0JJ742cpUloAnbZpjEt0ZDxAZogIGASh3q2vbCyHjLXYP
/wunFboaagHfrlsGpj3Yv2TSQ6dSuapR0ctUNbNfM4jMtFmY8cWgGomT0R2dbQaEG+1cCgkD1lAl
yh0SrJmz3ZnNORsW/13qPGU5FSXJqsJs6giKXE43wL+/H9YThNMCuuxOvxkbyK1D4A5RrfQyTbAa
cXLMwdO4foUpqHoIMdDs4IWwovdQYa84J9fDnauYEOpuURvsACtLNEKGnPfeglEJ+Xp8Cn2WJY9j
byYTW/l1XeQ0gvKehB1cowCbwsuic0dDugvaSMnT1k+hHIj2BO97Z4+wlfSRTaQMQdFIbjqb3i+q
iY5IFuTrAy80owoEXznLMsgljrI4vqLz0RArYKHumi3XweY8gqksq2Nd5mZGqzbzGiISe2DoSvEJ
hI/lrwdSDg8HgTDMPqGXwxL7i01SS+Mgy0/dgSnFcjEquCbFG8GnF8O0e6FDtSTEfzYmH+QhW//K
Zan5dwZS23YwQlrYShPPQyFecbHFiuIV64Dvi9/xuKGjaSuXkAG/cX9K/S2OokgPDDGHt7qoPr3z
33mj8apSJEP+fDq/rOJfxGi/43IZaNMEFPpeDektJ0Bve04bAGaNEMJsVvSCzU6935XUTjdpHUPH
l3kf8x2zBvoZF6vx1poJb9stosb4OpuMszPRG+xbP3z77vgO00K9roB+UAsY81O4OKRNdy0Mn9YJ
pFa0Y8YOJrjwCVEV7lq4xDqNCK5nLaB6r2rkJwmfSGR1V5DSmfSqo7YgdFExneHx3zUO/ZJ2pM16
DgZ+u+r9TmyYhNX+F/uJZhwyJ8WokL62Jv6tjMii7e+TepxtXSX2otshJ1c7m3M39SBC1fYTzaAZ
2jchXd40Cs7m0+Bt47CjlgtkkrbEL0QlR4vmeF1ykzNKueqG5EHKuRdCi+6WyBHecdxbG4ZOgYiy
+rT4inRfeN0VANtB3Y4YY4APT0/vt/OrPyi2BfUG6t+68USfe/ph/xBeZ4P+hFlsUbGf/EU0RlWs
cCzR16ZSTNBoy1Uvm4CoJXWBYX614xPYcllbeDRSkLUVl0jHC0Act1jdO1ffxxlt7R6PjeDbwK0J
8nhuxP3q8dwvKCJVjbaN1yeYo8ZgS6A7S/xCp9b668WWKZF8jM7/7UebS8Ftx4F4sc4xkfNr+ESY
aNvYDvDr/nbUVCGslDHDAWNQgWNxSuyeWPxbQcvfzcElThIwdZrtwKrU2Hn910Zm252quMPhbJBs
RfP0hICgjW8/ol6dTO5LsUocdc9woxWu1LPrLY4xR6KeGeR3JCImjz9cu5oPbE49vGkTJ4ERiDt+
tkuGYa6S50VpItMIcbZ1tICZesSRaykWuFheVEvhto+ZwzEkFgWzLi5I1+Vut9oraa5S/FZyOEZs
YFZzdK3bztiXF073qn5igEeEbFW8nXNJoZvEHEL1Vl9sDa8wCl5V9+IPV+bec+QtFRrwv+m+RDk4
XTbEbxKCR7L5GqfoKcCnlIvPvq2b1aR6cEd/9gmVQMuroDovNDANC+UfpzvXqdQXpqYzPr4WQN+i
pzTwDvptl+YhdhS/T+Np8aBhtCGb2TvhdqxNT2qNT4tSmjDG8kkxz5xKouoKLe0vj2di6XemVVbx
snZePC3TiGE7obvE66nNoi6+WAdvqsoQ8R98/hTuyfvtJ46S3PNPq0mZP3xXNeBAtVRRp3oAV8wD
OemfnzOvmMsoZSGMhIZUzumJ14zIF1RJoX7dxQB/TLkOs2SMSPwx28v2M1wHbjXQawICCPsXF88F
XYwGttKiZrsy8+ZFy69PZvBaqUiZtDZHDfUDA5NOdaOiU1X1agTtNpFO7FioSWchOuMcX9RwyabT
3A93aodYPubt3crd7MCVQnlY8HO85gbiq8uU9+QWyb3xEoEnQ3qiBX3AbX7x0CkeWLKQgvXB8nMq
GLk03MdrTshVccpcm+4cVhqd/N183sZ6NquT5RPWsH51NnJFVS7IA8P8Z5MHemPGLEinooFD1aoo
ArFG4fxJRY404ufbdj0BfzEzwxTbnqZ/H/+r7j96qap8cQxcP+i/8PTkZ0T/GWAb/R/zGaOqsxma
YDSCe3KrDS5xjRjoiZL1D3OWBpG3nJipDKCGeYWJMIJfOoyGwfbUAptny27zJlk+SUNcZiqaVpZz
hHHpD8PeUY0v3S6MSpusClpBOzOJ7Nr68FPB19yR3plhUye/fyftSQBsbMJKu89SQhNua36f7Nwj
v6Pk8LQdWJo51YGvpHUIohtygM6srU3qdajsqE0deefJTGeTCOlotuiw9NwWSlfJztmslZhK+V/A
oykjd7az27iUKoMGRa9gLoR+UddLLixwoXhEcbQBXkg48/7N2kuIKg8y5FQ/6VgWbSMwRChyU0Oz
YpyQWfgt8tCC7TtiADdPKEyHZhb1004/+3uzG8yHTuUFXW19FLdHhsRsWgMY71woH84iJqZrzJMm
if9fNN7dcZEvQ4maqMqH+loZGXCFF6RaH2AQEsnJdrPlP6v5WoJWE2PUiqZ5VVm+aEw1hZk+6Pkl
MwYeLg/7aOss4rqImpoOWAQJlwBTpf3tr7QhQhVCSA32s+zjZzaadlJtMWcpzQFYIABCRD6lbgOW
pZbP3zi4bwS4u3bb6+/mTzjdVDMftUXq4wdrMO4WMq2h8wI8O4Yjb5NVnvOBbLpe3JKNB5/ElFVV
VPJ3AJPBfnCP+yemzd+7Wdx444u261pMgOW1a3lNv7Ava7lcI5ILZxCSGFTh04LwOFhcYwsfM0C7
mYGT9vtmK1bFLHxetfjoxKM007TnBCtI1Mc5VjU5TrJhvPQXF/qYN7YKab961Fj8CWP0ll2bMN35
ndx67MX4iKLT0wKA1biAC4Z8vo4gDTEZesALujc49CwRSoHnsp7CjQvunHFNhKDUyjcYt6LwP0ZI
7wGXyRzcQQY8Sv59DJ2I05KqcPTLNRZ1azxe4MsSkJtznkVKIf+BAJV8MxXQPymIxCKDifKrgDGY
5Cs7OwWxbPyg++6T8eD55ZK46aANAwVXUe1y2BZccu6NnWJNEeniDiSb+bqvNSGHnGSK8yEWK+va
S84KxRPr2g6jPPbj31F/UpV6S8ly56GVo8GYvk+d8WqlLrVf/0baeUBtZLKKrKUP8blupr/F1OpX
/56xtb3Q3Rwdrtz5FKdimgWrih7Qo7kqz9hGaWhlx4nM0lNpx+nuMxjn6sMzgZnEIb+BJR4WnSth
Q1KDZvnb6EpFbpZARvLJ+XPDwYrw8iNhLIWuQ4SwD1pL/ZwaUNhXplMgcAws3Tb5V2A+JnRqZkBv
mzjLY4LCSiK3/+WfTrm32qs6syzmztr/MRB4ob6nIqN6Ixpdmyw+C34hXdbvi8TAGMSYsLJA6+0Y
1qjWRDlw64w4oX27otrNp235wua5+fuOPOdjuZQtYdYlrB0/c+Od9TN0RxoSmuDoSC562FYStliX
vdC3G/gfnCZntg9zucZMCcrR5KxcKLX0UCLS9ZSez2BtVqYOeKMXL8NXFEWjNSH7LRbAJ25oCC7G
cmjfu2Dl2b0NM01uOv4cW/dzS2lSFfKQTbPTzJ5SJsuS1QTmP595r8hmDO9igg0v6gjyz7uXeCLM
VbILfaLION3iQGXpXQ1QwW4SzV1j/zFWcFd+z8r1ogaPOsNwgdEMH2vqCfJTXAHgt0cRPcRL+EWS
AC1Zscj4vguOVs2QdzLP5jgufGLK8ukHzGgsUkNxClq75a27IIKmLERY3V0nZc+6MTbBlfZ3ejrL
yv4t4Kc9jrII815RRL49v3GlwTV6H2z0VK20q+jaJfsCyf9NF4FL2SlsJyzjuJsXADt8MV5djWHE
5fOoW6OFZ7Cl72012I3Njw+/ijREk2JPH2MiJU1N0ldIx34GPkt1mYNVb6oOsoAYW54hDLj9A9CP
epeCD6Z5gJXTA3qrYYFQr2ugbcsFbqcxeDrJf8SSnPCtSJ0TBYMa0acXrebse6xRKW79KNR9+CN0
rvXX/lz9C81VkMfLh/Y1WA9qND7erk27u7ZItZLdYpAjHCwZxz5g5eNQevssQDyZYqzgOBZ+UoZI
dCeg47i3Z+2r23YKcEqP6Gc+ltXEreHmN7cNrVanFhUsvBqNq7UTH0ZpCslfqEytmKItKMc/IIlE
+pTQpdFaJVi1DSCJ3sHX4C3yPRtVh3t9f86Z1nRRDOKT2OpGrHh6TjLWKJ/ymWOWMOUMl9gwSqd/
X4sMJvEATeuF/zakOqq53UFW4IyD8Mdldmyr51Qg7OpZscrkZb3JU8y9eRKMEVOKcMoNo67M/Fk1
7x6waXLoGf83c8ew6qFvXXCAxDLaN+9l3G7y6E2Us2+OqTAHtgsuLGBXumfofljKBgK3Xqy5/Yew
rYHYwWiHwIt0kajK0ykIESZp/YvUJGy/X4VdOBH6n1u+W+hh75kbDne65QgkgJSBujfp+VvHeGqo
Nry2ox0eTJ618OXkP5tEniyKDAC+hP9cA649gFMJ+aciexqiej1stnVY21u+NModgYghv/HJz6Db
/OAf6lsRzFkgE4ecbOMcNHbMaWGpMypg0isTxboh5yN9ZXbyMl0WKm2yb1juXxq/egCRufArT9Zx
bZuM1jtabiAjkfhRs/Ze9u7yREkyRTwXRhRf85lrfnuWNMcNK9LytrLiMXqmIzFVaEvpMPpaVspK
XFybbQVk8MSGj1LdvjNjiDWmH336/SkOC+q1y+IsK/bJWrIew8nLuoCkMGxPbYlqTVs44zlo0q1s
XR10SPSQnZ/6AIYHHeghyDrJ5efxpAxCWGoUw4JVObsvR5hE+mr5A4eYtkGe6Gvl+dEPDtXlTSAE
iCMfwlCnwoOw9EFasj8iuTV9OCZmnAKwz5tjRTrUBmCYyoLb0KKWv1fTnVot50vkrTIK0u0CaVTR
I3rJKN33OLuNLvHxpcBYVoUrEV51vdWNvUB0NkGoBCNTZ3gs8Cu7L74KWfufiQ/Tjm5QFOBCNb7/
AJcgjsgvUGoIwBOszusTcode3j2xj0VzCJnKAVTf4UiX8TyasRZHJgAPFcwrixz4r1mkH5DyGMCA
23wIwS+VevUPnVoCtPZ6Wp5rTEg8l1iNw7+rgEq25UVPNEJdLT3+MKpJZwp482Dt2m4mJ9kW2EOk
3+VINyXnWpd9SacqzmY4ooFSpKBlLOK73JsP5aJdp+cvGwSF0tM383vLBh2300KqAFM+OQNls7Jt
2T9ez3rzDXkwFB+qntuz5nS4R4OUarzQvF4qyfwq1nxQbf7/GKNO8UnLL1UqyuXIZbhtxI2jPJAb
CXgzj/fIL1RYdCNWugGukhNCyTldZFMkIv+iIdiKQKfl19DU293bEc3iZNfXSFGkR/qw/tsId79Z
buvOkoZH0kjnOSgx+t+PkR06+Y6Wq53B9F03MwhJ7OeRhFv6iZn54KXG+uUKqZRCVi8WOb2eyH04
uX0EQY9eFBkoU3CR+EYZM+pDZ3pJPzYvZvGxGIyAxb5MMUVzkrnbmScfvmI0U77fAntACW+NZThm
l+CBp5OskZjpVuNj2lBwsviVeYhI2ViHZBOnJYeBWAOPScV+oRbOJXFSLhLzU7ZxwaYZPLQy6tB4
nldE9axp0yQv99m2aJLgnoCCXJRIEDsviLTYwaDRsG+5k1uupPHqEP+SXWBx9DmihAOW2LZxmYoF
YY2mrMhCeEo/m6/NASOG7/PM3SlxRpI5ZLYWsfkR4uJtjJcL49kF1aBrM8U6jSysAFXeXEX8k4uE
G05+Pf0QnThNOjQXk8TNY16qawp8eN4WPI1ipg85J/nw04O4F8jCgTb6vj7vm6FEFwMn7+2IOA75
MVR/AVs24aLXHJrkEN3i4xZ6mrpC/cSa2wCfV5NsvuJehEtB8onqrFibdFeBeoBtkjfWFyo19o/m
h5198Rn2esHgnBfZs9fm0w6iISooU6Agx5ua1eLl28zG/OM0/+Hisu+0+6no36FyVDgbkjTT4KAL
tKomfCgZ4e2eqP50VOXpnavmWPXp/V05cjZf/0YYbs3NSXrf9pGwlo/dNwwaiQbx8gnM5wHBFIdi
/w7O1l77NkTIiRmVYj+mzg8WnaHcIyoYk1w+VzmEHlMYKbRCYk/1E08A0eEXAh6Vou/XI+WWElEk
EOFPZg6iJtMIFxsWrdfHc6dyNRf4PAJIflZqDI208R2jaaLZCe3lnQhs0EcuAQzX/YTM3wT6nxc8
TbaCqWE3kEx0BY/M4kD6Jyc8cnLanL6Dec30zN1z2B/XmtvwQ9GyifeKc/Bk6OWVLMpn0jAyLHRv
GgnyPfA+7iyUneRSpgadlXq4Bvy//t+UyBte5h7/kce9tOeyZx1FLDHzismRmbIhimIAgc9DcJSA
BKOYYrLUk9YH1+y1FlmpM75GWrOCjSlxQO1MafSGQMBQ8S4txQWGSqmN01Uka5sNAjtlG/8jGv2W
s96TXkeM/mCXDOPQFbCTIreTiY8tlNFExdFuLbqabmYsjvMUYfla333sKsY1Dm2p25KIJlstFZmI
JCAJ+fbJXcvfplTJHGnn2tVnBWv0f4LBDljhb1pmCjfFIF35G5Wc2Qtox9fd/rq5alzTjvlwrTtC
9KLVyUC5RQI1CkEu02B1HdDhUnuS+P1sCh0joa/s1GwFCppsyJd5BuFI+UcRBozl2Ao4XJx6Bzli
n0TAjq8R8rWfmNJ5QbUQFSz3KEly5RSmZtHKgPkDj0X4V+1MR6g50jhiSaxBYJhY3+zZbHJ239Sz
hZ6dx6kqeBX1ybpTN2d3PVo0wvzVezTQ75rrtj5fNV3yoHUo0MuN5FcmLQgbH4GwsWmyLvLX0qMo
CXt1Vc/Ug1FbCnmkw/aCfYw77WpUbBBGe9jZJdKbQO3Yo35JptmJQzpTrDM2AyfzhJyfnslB1IfK
iVZ66pvHl5ZTMtpG0xMvIR10nl64Vkfl+O/TUQ44vpi3/Wl9Qr02s+VRTfcg+HjlCMklzSIsAOvE
NVeman760zRmcSSmZ3+hcXIj3CJM+QY4QCyASKKL2MZMTEX7gRtPFELOwTwveHyKcIu9xJdJKSia
QECqNf2KePKAPR6AR2WA7Yyu+AA7SZnyHr2zMtqz6e/ygPngIebbmM8bmi6htFZ9w/iUNaOBK9T5
gFRuzVctnK4ZHcmrkyZp1iEmwW5qlvIroeOiZLyK7u9MHlQ5HylODlJFRGL7V6zHIThCHHRwcMdn
K/DtHcNoYRa7JhsBLZMswoa6e3iBpfX1W+XByAAROwSVKVlGg2ikxMZGrK8gHCcwpwS1hJ5Fg0lF
gK7ppZzcO/AY//6xIWi4QLRabyfuo4VZb//M57hOku//eEKuy5tAsmvC/I5DkZ0gNgcsk8VWs8iu
lme2mF6LiEzEhOSrtjlaYs/2tj/BqkV/IZnyVUQewYp2tUgSBuEsCM6hkKCE9DDPZN7mYVf7mZve
XX7XjM7l5om3Spezwdd6zq8hA5ExpophKf7Ea/jIXfy/xbLt907CjRPTSyiEaVd/lt/xdh8FkuV7
usw39DOP0jsKrAmlkPU3YK5UauFiCqCUWQ0AyRHw7axYrYv6YNJ0fu6BMr/7aCTdoisluAfCc3xL
J/TjQF+uC1KF1mCJDhvTtE5kYfsAFhQGpMb8962LYelj+qj9ZCgzOi/NqaVDP29Zr9eDC0CORqkF
Gtgvgbw4PC3aX9+RJFxptVk7+uj1TldnspKcVKcfRd6iqQ5G8YJhAWFoznX+bqSAG1c9jopg0dsy
u6Fm5lFX95JQohIx+QcJgjBbvJK3pcaE9iKiABoQX8xiPbPiQBGDwWFnBgePhzg52i5xPav7eeIe
S7FjBOcHQQGEEL4BLjepAYua9CBiGeP+kyVkUsqF1+2CS4P2XjE/dU7rY9Igo+NA25XEP7kqTIdM
hpuUsuOKdb9Ekecfc1pXjkAqmixuH/2LUijxftMSDBidi819mUQCdZ3SWWlR3x9/RY4PMKtMbarU
fn2uhaATLC1aEM1CK5nKf+6ZHAFxQKYYFbTJbRNxaDMlfcQP207yGNSDCazG2zRQ5FDoFSlLc0n5
D1K8qazXFnrledguofAbbve3ZxrJzpKLFw14s4freHqYLzN4bVSS2He/RzTQI9IVyUScNGse5G1b
r3YRhndIYbbftDf1RTB3JqTYrlYMBxrFxrS2JoqqGJcYJBqhfOCpg97dF4WTkKWBCj8rWXBcoFef
W1FKwsQsORfFOfrwlQeLWlU+gaKxdtx6rjOmltGtuoJ1W9LsBk2WeWI3cd630gL7RlYMW1CevN/f
IMThwJQpzBYc55fTijDJjALQZNMIIGAz+4Y5WvPJp5bJZ/io1k0pGkpPODXC+bZQ0gcmA2T4clKI
NKDrIdHTeQWgDY0Dq7rzb0oK/RWDPompOSIos7kzpGHo03ipSNoRfSzN/auujMGnASwDXYmB/cth
4qPd+YC8/ukbLWMgZ35lkf9Bbj1CsD2zg72SkhQei2Y/MnAdc5QEnPHX6vY49DucJsjbCwUwKxSS
tsRRGVelV0sQX5+Oj0HhK/lHGUDfHRO4/2pZjV3M4NuKLQT9AKzEVol3GDRlFx4O5RGacqvfgD8T
5rr/T+V2sliEJmk5p6xO4fjP0s4ZvAp3CoGAs+eefSz+vJIiL0r7ZnUPTtbnEtA45VjQ8awSFlHz
7MSdysGIs2zNCTLpOpTb62nYdBYxD7vQOuGjUaUoC3VjN8FwxPT3kz2uoTeLSbSwyiCCKluFmzMN
e1snhG+Y4NY6H7nIFIlP8r2pwS041IHZnE1wdBdyDKyRndAJ3BvE5mvnnv/mPWzduuy8gUtrj3Gr
/evEYibylJ/Ki3vh9OEgmiyyWaprkWZuG4eBfmWLtjSldZnJQhTSlvyIO0DhZvuOsdTP4nyoxlAR
zjS5l85gEPk+dKoalui79PVxqbvl6Ds0gk+zO2qxK6neqqd+BcLrLfbxPBn84lrpctg6R/JzvFUt
ChNNAx4rDYQ0uf+hopXgvI/U9pfSQQie/GVKAzjl3XZCv4p1653cpwFZaqhYYuSvu2aQg6MUGckj
V5QrTMR4eY4EgHjvjKt14j8grcAQn8AsKwpn4pZAsGPf/oHoIik+/nv2c9jh/906R+tyRe5Njo2o
7Lhzhb86BqINY4czPM0wSdCQ+/4bMG/EWxQvTFZYKpbKDKigTRcYRupztYNMJyZpNpTmwkqRm7/J
f8pIvCrsu4rQHu6Bn+i/4lCCzBABnGmnphMW49CeKRVsAlaxIZqOgt6XMskDI61c+Hfw5k3JvIg6
1elk8scCPX3jqU4ykscwKKkc6wS/AHDtXrJ/tkK9ERwio/of38OUf1fnTrJ+D4npKQum379GYEzk
PemqPzWsBrViTI+Umur7HswdN9fvaMowDiI3KFPkisWsOWViWK6C/bZzxIbbCFgDi20h5PSIRJYe
ahs1bq0bd5q7hdxRTWSBxK454m5moFvPTo3sM3TwbTG4TaO7FDZuSAIZkkFFBmdAs6N/miUIwnKt
lyNaA3gpPv/jGV6bVtO/pdiLSbw/+kVgGYFPloL4mZyf2McpZUYICsol+AfhLdiggVxyDCBQ4aUa
UmoiOWe6fM68Q4/k7icKnt2zr921uWhs3cC3lGeZUxBsAFGYnVTcbzoaoGW3PVr9tmaSFSWUE3f+
NVyL/HUawJ6gYKuFLaZrD0x9vp4AyWGVOReOPXIPll1jwDC5KO2KIa6DMv7EVSkj8/z6XpBAUMUe
Aw5KNOlXge6ejP4En4B5Vho4JJbX6OPzPjh8V0UuJQ1Og+/oWlriRkNFGU2KUiwDyXKtKc7m6ihb
vWLe3dib20ET0qg2BylMn1Z656K57rWYOskgWieTeifDmdjflGPsfTPpT5YHF76Kk1sW/Ad3+3qq
AS4XSGgECjRouR7Aw1XYCA1jgwc9R1LzeCLXan7KMpjaxM5xI1WJUInvC05EwGyiwzP4WczuuZkc
OJXnbbEt8BexO083i7vqnB/9Ga2LeecW5Q4XEUTnRjO01syVqw2zfX9zTpJ3LwSjx2SMgkWYTNRt
IcApqUzGmMUlnYNUckDSnqjy+khh6dKgGlkdb3JtC1gAPbJ/BfFCdQl5lhO/Anue44BGoYArgA07
3ecVoZuXJ36HekduYL04q7PDjLSXtm8aHuHHoYFkqLIUou2taPcwZ/SqJUlU+JVbSZORqTVBFLMg
27Q9jALK7uZ7NnE23q1JGx3Cv8QKYLsSr9w2pKTVUB//WuyTCt8Jp9i0UkmH127etASGP6iTJOV5
FUW4KoouBG5vJAOsDp3MRACVGe9ijX31fmtjzn+j6CIThZfLZCJDSzSKM6FBmao2HWy2dnI7uSfJ
z1+zNN27DoAfPdB/9qHTJcjPBS9kmBv5Q/ShLD0IRoV0XDKNJq/s5t4cJXYaJ6/AidhQq48GpUqk
rr0iIyxY0Q2L3K/ukhxOuqOBfW5Nz0bR9lU0uZQmPbUmWDgO1JxnaHufyYpkKgLV3SOMEwUo/0x8
Ash1VfASX79ecyE1I34yKcowYCP/6WVfqDd9M+ewQig1jKuf+ZrJqqCcc8lSnl1vXkQXiuYa12bs
GR+3cVZR8OnBGFDkXyvDcAYojqf7B/pgDTm5ImWdpZdQCnYEyzUzn5aqprRTx2EgDf7L1QKIr8y4
wDsdorevtU+FMYbfSgfTWw7YY3JAFMfK1HH+m4aJbsmze8j7GzenTxsBliWZWljwsBCPfjF6iyhA
ANpR5NPXsr8Omxmv3VYBdbho8WYMMjI5INX1XA/vY6sK+pojBsPVW/veozothCc+x8CtShL/8cdL
PuCiMTGYwI5Yu4Oze0aiJSr385pkkB57YDxOyRDZFod3Qtcejblc/R5Xb6a1ARyoFor2jXHjp/BZ
Bw+nxPtuHAZmz8K4BDsHuLI6z1ryU7GI/k5g6TmGTo+meKLUtL+Cf0TxWG/QUzfc6JAihMc9lPIU
KRTBHOFMKnw7K/dqb3wNGF2ttwB9luYnY2wt/zLlOtR5C6J7tHZejkL2wkiWXwOrxNi0XZMTxKJB
XtKEHCW3G84VsvX0qkO27LzcK66/CyYDYUDPU4RXDiFzLlzoTFoK6QCvOLbD6HNL5tKaa8TO/GUb
eBjpmZEMHxPhHFB02GPvlu7KlRu8NqF9xCCilHpE2iH4+44gKlIHYG5J3Klp6J0vU0AKsm8+mSCs
xbbB52r2dlc9JDcw+YQnRDNM11idYZFr9Kp9FMN9ELJTfwDOjpoIo9UJmVIoa5sW03+cgHdTFgvU
fwddI/YZJon4z5zp040pKiNVF60fTXZVg6gI3B3cQKps38mVRyDVbVDcYckSARhv5EfR79GtkfE2
HXPc5CIefjyrybyALJc06RZx5kQGj23McA1q34169ZrwxuiIfNCQKztir7dQEWHHRiLOvXCNjh//
ZqzT689QNw638Uw1Hq+1gXvcLDgcEhVm5yPbjLQPQNDMMkdugdBgHOn8tAuOm+91c4Auy+yRIQWY
YvA+WD2TRxE1/Tp0c5GZDYSqyQFp9PqnCH4TD5ToddYRFA7AVjwJSOIkaaeHNZeB234YtkcqtWfL
t7xhZTNJrJa6pxyWXO+a+jSgaGuyG3lDghH4VLofxT8kNYLd0WIaxKGCjsMUjCQtTxT1WDDlnhKu
zCBER8ogkGtCa+r4ycanmA61ZuuR2EPCaCoUSlHspWXnyKS+AqqcynInHyPoElIAPgFMDdT5AE9Z
hV1E7T5T769XLmGURbdVNIWg9+zHU0nphNulzvFYu8HMYt20AOU2ocYMCS2uErcT42/aGzFZEYrK
HOnlys3DTbTJYtC3/kmRtKlz6EWDGct8CO3rn2GERryOYGs0Zo8znbHskt9bX3wBtUEfV0Kqa1SN
cCVrbDwYOUIt0P37XgwHbSY7tGGKavEPS/pNUX3hC73CM59G8fsI9bVdDh2PSTWQfM2i+ZrhHo1N
9ntekdDDl5GmVZS0C5/1tiDOcwlwQXy6rbRKj7XYjr83NXgMVTJKtmeG9z5f1MVZZ1F7zVRgAR2Q
CS3E3nQ0Zbh6G/Iu//ycHt5ZKR8Zy3pTGuI3u8UF2baotDDGKoQlpJt8GCwT2ojvj8rAnE6ytYew
TB4j5jLiXta0TuPX0Q5NeLh0YM/fawRvHT64KlHwuUkmyAYw8ITcetIw1GYrHY0PG9VLtt1YYdLc
VhS8f5i85o+OdhbI6mykZCxMdZfEvSPfEhwevnAS+xToU9wS0TwJvP4X0t8iThECU4q7Sy+gNT4W
NNCZ2rIHR/jUCOpbzlkYCeMi1Et/ntsw8u5HmeOeFIGSiERQjhYVrnVW0Xvt+h08tMe7MvWO8p2T
QOYFUrqqNGOOdkrOJF/+HoJQTVx4nbANCsXco05+hAgdH4snHCMFfWv83cJpvMjuAeSYCNSqZtNi
/5iKVmihihi1LVUbVJKqsZkiRnsLLzmLVzuKEVvKKK5VxvuAbhJEMqsuhSjTiquZxS5JZfwJmOnt
IBRe+1+jo/cSwtuLK8XjsegyfcPdtrvyowKoeU9otOtKQp1eu9DUgrLzzbKQsxMYqHTtY5CUAMNv
1HINNwrUQcVBtUk2CQTqa9BOMovuaHit2zQzSs8PD25dI8pf5ZmjnFmqGl8QfIErP7PWJ901RSr1
HcCJF08JTzonRVt0Us0G06rIs130akxuqno5St2lvLOxbXc7K/jkWLFRVUsPQuEHiIiHAb7NuR+F
PusINKRB4OgtN0Wjg3GXpCDELXeA44JLLpZBNm+4zFl1BNs/z2hTZ41Qrg27ebA9f7332Uil18VF
KibFfJIBCof3Snq+zLP2W874JFloA9FrwN8zYIFC/RA8OU/L99LcolJ4wyCu2E7I2qU7CJNTb2Dx
uSFqO5MQQHv7j3BswX/S8hgMU+nWTRmUxZRR+q5kpOJxf5DUJooX8XGEkRQKaXFWmMoUAQhu2nhU
x2W1/CfrbYXuI+cvtvvHrqaCuI4IevtafgXhYRyxUJcLAwXqwnu46pNKeVRMqHtlEpmwY17kIlkT
Dq9UMiPic5xHhh7jk8IvnAMuzH3ZRL9cXsP8mb8wLgKe93/00pWDg9axSmvBFmvBfJO48/zQGPRc
cWhEipOqaLjbA3iQLh1NfK41+XuVXd2XeAw3I4Q3L3zIDF7IHQyzd22dkjLTGwBzlpNGaVV6k5yx
KrfHAuNJlH+UXAJpeJY0roC3VyVvOQIeypsvtLsxz/8W9fhHo9Zq6cjxNtIj4pqFjrEnthQ+FMWH
WQaR7bBAL5AbE7gJ2TXbCKFZdgsBJiIRAratdKRCHzCmecIPXifr9WpAJCk9UWf5SqA46Q0yghhZ
8m1gj3SGrifJWXwtart389LptQhpXDQTIaD4b2eBZDYEiOiyX3wv1/0F2tZSRO8KLZ0dFT4nFlGJ
hzTJHyEYJVborsnudVDQnTKns+7ETL8R3d3J5+iOYq6uI01pyuT3mnw9D5Rq4vzI+6t/ZreW/IjK
MAn+544MtEddCPZeTA+TBUuRvSARSjcADf9HlAr2rHlcr12qzlOiyVOwiZ4zGXV1x0Ww2U9UlYcA
r5Qhnfwznk2ThKakAwc53K4dXfEnpWxwGb+Ws7mCd+LDLEJ9ldTieniZjRt+tggL/pO/fU4UBDLd
JVZUNOEgAcV2Dk5HXriD+YetsPZMCqbhvoEq5HfWjoq5MwVBj8DSF6UO/ODfMX5KtZsdsc3ZJaLi
B0U12MSLgN5OBydMPDHW6Mw0UX5hvVcjFzHxh6c2upVIkZVKqvs6VEmBjkDHYAd4Jqq+JfrZXyhZ
yRNZt2itjjxElwEq3ql5anAH/to8aQxiBndxzY+GNhNniykky1NOQBpIaZKp5QXq6gOn2mbH8Kdr
hMQ03WGl26sFi86QLFXu4TGkCMJklJXsCf0F6qtSHskyj+4k1Ru9Xw92m2mAJoHFKMAxONWcV47h
jiKBsVmlL09KA6bTtJ4oaXKkpVHjRk+/4vlFPd87FFGSAYchYW/5bD9NBJ13KRmO6/2k9RWr/GGf
iPIMPQ3q1IUV0wIvgs4oIjoTb/8ggcINkIk2zY21D8V9NeyANEaPCbvT1ObtBhjW2PYPwez9YZhh
Uu1l847SW8fMOg5dlcTgy8FoDwAHVKjDEoWoB2Dmzs5dfh200AgvNROuDLi+oQt5EQaIc3MvMOCu
OTMIBX7FPLgMZjXKjZKL9/JHAfc9XIZ0oxK45AsRZTJlhnWSb5XAwbiy2I/qCWdpLZQVRVpihrsj
v104Y43xrBgocBY7boGQYD8Ie8xraDvvGAJ2tcowspGT1z8FgIEfr5ZZLj+rf8vBaqJcObZu5IpV
Z6Ngspy4JRUTcZR2WXmV7Wz9Fdr/4lh60//Yy1KRX1/yvuIdaIanUO9qHp3ybNJfzQ5p/QeJkpdg
bw6yg5I240Aoq4uld7/J+tfVP/GLiQRtcKzkH/j9bNlMUmNURaIAJFCJfQTgV50jCw5q3lr/PRc2
xeFvqIMFrKH7xudvCw5JEXsGGsocF6Sz7ci3tF+IIxZqUrAR/AFYIyakXXchNOm2xyKYHul7GHim
3yiQOZlknY9FEvLRvccx/VM0nRhdpyhwWqF19nBKRc3MYekjDR+T3RmKIvWzaMMCJOc0T+VCfJNr
4zTm4YVPljjyctsMFpAhb9Dkvu4k67ZCdKoS37KGVjrQB8NTLGQ/uwCHRUlIQn4WtxPwt33Rm8KU
xy9OaIen1iBwmt2dLxwM/bjQlkgshZpACh2HoRIGZVKYr98p0pP45NPxwSNir1EdwfTiZPCJb+sX
OLzebcloxs+ROsSu3lPiDUotNaLNCGWvCceYwKy5T7vhmSS2qzWBnI3aWYH+I1XFsrtpgZqqTtvv
ZiTSKlitzOLFFJzkta5eMN4nNK6zXATVVkJlTX4wFLrnkToZeOQ93j6o+R+o/JFFdx1/E2AOLW6b
LBYd+MEpj/rjgpeBQvnHy/tDFgs5evzi0CkjcxXM2Zv+se0g5tzRgsFnAxscluUoQaf/HszfKdtz
cGUI4wUL6kPRp7FbSZebJwQs2Tsl18sdaT2wATNeiGqcQ891Ic3bHWO6dCzxr9VhkW/1ppXgclpg
6NstI5j6iQ+7NxVL89LbGY3QfR5pLvydfLRbwnzopy2ZtHpP4tR4f74/oq8X40nG3pSaf2HmYmkk
JRh1Pz06OX950tnH7z7Eav9WQIeCJIHbXEE5rMolGeTnBSMxqr2Er+lV1om+2Cb0VwSv7lSMkMh+
yLB2xtQxgbbnqg2YfugezSmEI1Hg4cxtxAKeEEzRdysZwXs3+yqA3r6ZHExn19QEGieA5HRb3Gi+
BqP1N/kebBF94NcqJCXnGrkeGjUbzGMqrUxtn9B14lnIqmJGWaTKWsIdRdF6EL/cBPm8eP/ajF+a
7aQbIUC0Ycq5iFVnrUW55tIbWyRlIYmCsAYW/S8HvpWQQ3XtJPT3gjnuGK86LGmk+pbXUcIR62aO
T6lFd+LYIE06m/IYNjrptqqN40Aw1IHYpU5mGq/UTAS0B1WSM2u6TnsfjZkcyddj9qR/uyiNP+uQ
dQmUs2fvM9+6yL5TwJKUad0CIQRapGn2iaKFjnP/xuB/BcTD7Hfw989mgi/fpNviV+nuJb/7BEWn
Yxz0KMO5AJw51i5E99PRH6wZHXvkQwkyJobYjaWejQL/c3T335gnFQb1T32HZ6y3swD4le0wDFtn
9mX2y4QgMyUZL0Dwsn0epe3C93e0cGGCIp3gM8nxmS4O1kC+NpbWKZKSHt7wYEsBKG5Mgdf4mfl2
ar/kyeysNx+JM2showY7MWo31njRoZkH/6zPzyFll2wZNc5QYZVZngF8zq/7/lxvg7updi84jkkK
iOXJO16f7SPJDuc9SAKdo8ZxGUaM9Maf/ylqq/rwe4rzyda8a2fg4sqvGInZs+eYsQ3uwTcSThFB
9vqbkDJBTg0Fqgw6FJMqCXrB7/4mnqqd+zkCBeKzbPJT0pfETufxWBBmrQlZI6P/6ctHj83ati6A
iNWeZ+aRDRWzRcSQA9hAGExzZh7+CwbRx2POx9VhomdYyGhL4GD6e6IOi10DRQ7pLcgBzQ3qN8ta
mRYlnhF3PkvQLbA8LXx/EP8+Fb0aFqjTd2A224rfYaFqxzCY4LthgH8kZC/nPxvt9GPU4uOETv7W
Tw//MT/Mf+w2JR4SdglcYE9XFpMj6q0J69s81kORNz853PBq7/gHYgaBk1b/SMdRWoxaFWq1O0xC
oYYCgpZUp2wDqqPYIkU9RghXK5csNt8TwNT3mGw7Gdh9xfu3sBRpZnRrb9wxDAHoPgQg21K6906M
b3RllUaAwz2lqfrEloohDU87YmeC4ixKOfq5Y8CXDv+QOXCJcG4wA9WNcsNcg0C1A9JEZzPpFTxE
Sr7Ox+k6ayStLAE4+WjzAQNFEsc56PxBmjw9fw4KJ80ZCJK6fmkSuKxzIB1R99J0MWN0RKAjWw/P
VknEB9YvZSUnfihnGH3GqTRYSvCEMLbSKyMwDTUGZO2j4Y7VwH48aUWALIAfI4JwlRR8hs9Dq44H
TD+3Co8F7LhDTx+BQyXBurpQ+lkJqXxUGlPVMBOwv3wz/pw9mimE/t2S7iaArZjYd5/dmKUANat3
7qdP3g9hx2AsnVeC0Jdk8PqEBfd5JOr3rgxhDgwa3xl5dPdpFChi3aVVzi2lx9l/OYQ7M8Gdu/Xx
i+lYfuObucSLaQL2L6XX6L52cVWK6j3Axv/0Ph7ZBXzxOtmaQiEq8THTttxDODgxec8jciHm+KqW
XzTgMG/O4PB0GQVLHXKMEfbqiLYNJjk/2IwdxWZ9nq9e0rEnEyF9496OpiuMFZUL4vhvTd/Vlx7g
SJK/7zL8ek0shqhkrlzqycEG3cHAZy4rbg4M7Pli7U4WfUHlqkn/61IscBtetwyDiyfgtr8Qu6YZ
K+mi551opRcwtlzqCX4NvzduY4fLb9u1exea/kcCfx5d7diCrEPizb5eiy6kXDWSfaE9JNl3YdEP
SvStYLtsWKrVOG2T83Ifod3t27BM7B3Ui4zLz1klLQZmNuRYdsowu3vRJIv84dtlCwZNAlVYOY9m
s7ricxbMvR6+ct2UovAjgW+28RGVT0NMwWqNBKr0YCNjwKCpMtY4HupcNz9pqn6KmV0MSWi+/Gcm
ThckfXCSrENuIeTsAwrTPOoVzGrpPcjplBQ/q8uS3jqQ6pHo6TjKEkiWmyzbyWljgpwr6KIGSwLK
l+eUAEadbTxDTPtzFYV0eNLCTj92DbTCv3MMAA3BqPdIyCJYBm+yihTOtetuYA7QVp3qbfRJ6sAG
I0h3hdJp9sPy032ELmgNnRCieppYrk4mvOYAJM2ftAYFjjbGRG/8KGrksThUIXf95WpJZe7cbl5K
9wNdR0QOwSUyN+TQGbOK71NxDRyYtPlmtgCfy2YYxS1zhltHNB69f2Jo+4GZCseC5/3DaPMQ8lpi
qAo9OEA6ufYgNE7vud2FIKX7GM9W6g1G+N74eWLBA5nyae62gtqfL0dWFy/3Ck9R4Relvv3qY5Bf
X8XKUd60L8RsJzvxdF4R4gmBCnV6S/VH5RP1VmBPSUJt6y9ORwG5tEbM/jvBXo7A2yLXiwkFxfdp
Fk3Vs05BBzDj9RgTiLTx+AJkYNoPI6EU8DBrFv2a0RelQYzEnBoAB5i8ND/JDdXsO0qjl3/e/fUc
7iY4+EyMAy1OT0bMgoQak5RBYiCCDAuqy6dSvwZbTYePr6bf5odsnqQBu5tvPy81VC/k4+94aT3b
3SU+gPnYzq18BUl7zToVRmu0aYFAwb/lW0Y2cPwgyTv+leWbtjbKnGsKKcZqV8gP+YNgnaV9Nl7V
prwP1QLxhjsQP5sno1R/mqSWIsp91T2LnXTp3OnbOWAEJlDLQa+//eaZlCHtqAvySGc3tl0AJk96
nBSpq/6y3y0dbgL9cwsXDVm72Sy3SCNDS+x5TJpGZnroK2Cj1cp5QfWTvzzKKxMxM/fMfDqpBVZH
69x4FDbOU81Z/VaQzF7tQrfkGDLy0s3Vq5AvLXM4cDOmRZBKiTrWT4NR/Z1H93qUnGL9rD/o9fLG
QgJFLX1ZA5UFPj/rhhUioYehjI1VAftcyBxty91fh7/MkyJ2JB4qYuVLDJDXeDiitGQqW8crrvA7
ZhLP9hHeqUXK1iEAIMWtHzH7E3ImH+OlM6LsSi9aRy8tH+FHyxVerzEn38xZgRdZBxuahAbPv+dQ
668uVE/kQ1uv9tgXwXqrZPqT+YRNr4X1ikXQKmtITHgcxJxJGVODs/rGdFxdd4D6KId71YXVKqvQ
NzRSpOgt3R4YXtOEN3MciZXFoXO2/7sjKhrmJ6X23wEDgnh/Tob6J4IoIpNTPUvVHCme/md9LPNK
C+6ToPhN1WCHjRp2q12RmQXXvnjrgnYA2k39AgwbgpvDOdjEtvJIeT8kvtkJA0xp7ymHNKw40//z
iMkOV+hHQ2euKUbpIhK7PxgVMzh4mkNJZCZe9vuDPzvJQeK8v3AT3JPoh7BI5C7AxwJonUo/w6GJ
SwVf+pPrH/0XZRadi3cMcnILSbitkIG+rVTMtg5TzOpf5izXehnX3/y/4gBwe0fZ2Zc4AE4pt106
nQU8JG1jnW5ArG4aS6INY1FoeuBYoWvDDUT+HevdCuxAG87vWlLzCfpYuLRpY0T7VbfrjcmJWg7P
bscanUa2ZtfvaJXl4o5sMlCnbcoHHRzZE2kDl2EFhmR9MvBPHB2exP+j/y8JDIpc/Mq0SJyAUtUe
30Yp0qrdoxiaoy/7JwAL4R7FLOTEVzY2RnK+hxe8lu4iOYb6r0Gtf2ABRA1tTM0om3wvH4iMq28v
U8NXyR9xrptJ9yyM93HqCQFd2wEUz/4cU2xSQeMPDwvEeFNVi0jE/3nqJQO0nJ6EFB27KkLMZ8Jm
sgFaAfWVd7Md2tF4VHNTUaSk2IS5OpT7G/qIkPSSC3tN3vBRVoGzWB4U71QatYDROZz+wyj8JYEK
fJDwaWixcRqcRT/YD8fmXBg7T3AEtOZ3DXpD5ny6LvQKLCowXzI2m/KTyNpptyrlSg+ymFccYqFc
4aMJikrTsiTX2e5dx1vNSjug1SYUIGvnfw4pPH6GUxuONROd2AB+TUIkLKCChcxCG0klAZxm0VGQ
MVXlgtnHDZvNckDI05lq2Oiy0WZp94AGRiLA2W2rgLJkc/5aaPx5vskPkKAAgtQR+ETe5XXVocWx
D9xBoqBP/XvJnajutzxbxTPZ9i/GH7AAG8PupbB+aYMgpOj/Hrop8+KNdvbygKmCPBKvsVoJvVP6
H4Amue1FDvoSD1JxTXtej91U/11nAPBpVVmYjNfJWem0dJIkZwNqQ42w3/FsZGTey6zeL/zYUhXX
DibZE92scJ6CC17HsWwRpf1lQ9JFS69w090ugaUvB39vK+miz4flH90ovfsTGNt+R5t7mw46zUa/
XVO6QSKPk5GegobbxFzGhbp1X/a20zfrMJXicNsGUFt6jQNXmeYTmddncJVAxXEJiiEvaUsxzFMT
Y4C4TC/1zpH2+YSSkqhwzJzp7mnbnpuycBOQCS8ZHizRE7ydjD2jPSEIBwJsWJnxkp1kc1rIdSjh
gPMztJeUO8WCPUhOkvIFzcGwL0gtBPEW/h7qH8dgT4ot54W9Ma1qxrDA1l0c0RvaFktMMYbR6Qju
Mt/Ea4ZdOlAnFTnQIMwg999iHZWmDlov1mXvjW4JgVNgNTwMM+KysfrJ9YAS+FXvT3lmANW7SuMU
8m0Y2OAglbI99kiLFJPU8Baahp0Kf9A2aLglrDxKtPNQ2GhxqTm+okjv8g1vSCXbP05cpCtWzNcq
LhYeIcTK2pw0Qwd5V9YcDi+9X6Fsfh5E00GrYdk+GZL2lldF3PxXmybry9kUFf/u287WGi9jlRfV
TwglwAAArRl7gYcwOI3qJSEfr/BjGaoQ9wfAssyZHXwgNmEaoX3RyDuP+TvSDfiBdmOGoAa69pR0
tmZfDjzJVQOnLHIz/8wPwucGgrSrx/k3twOkA48H/P/axeIlt1IqTSQ1uazm6NojjPZAC11y+U5X
y6NTfFUsUnWow2VhwMRzyUbOpM5nyn12rokmFeUJtUq5Y4bPjoqlmFDZZpC26cRBeB0L/YgpeqZV
qPtu4okVPm1gX9cjXlAX4ZGdxZl4rjMWSByMD5UJkVXi/SD8VhE5gQIPMOAhJuLkRQ5j5xfH1F9K
pkn4yPEZBxsvPKA/rVtU0Y68VmGnde0PJvkPOPiY6s+7kjaC7zRu+9RJSHxgisoyFntsjSp9QQtJ
J4ihxKnUvFZ7ypNRi+SAYQi7j53zgsAlMCKdGoVUWgthUx7FDIG+gETZejt0xVDpOa12naZHTFNU
UEZNOCXOy5LNla9IJZ24lb5C06Fed2I4Y5PG5YVzAAQDKPY5Z7Rj7aIc1tbFCzYlX+e3fSofUI5Z
VVoHBd6iTjnnFlA2PgDeooCTBWQycpzQHJKv9rGP6+OztsitckO0YA2gl6Q3viAfYC9cXLoPUrM9
2P/zq2CUa09pF2v5bG3uHxoXdiBIDIhPp7lJRm1S0z1Y8VLsbZ1e/jKMPrp7moC0MkUOs9BQ1tO6
B36e6kU6u8OBIGENaGiUF0tSPzHb7WlaCYDA4LfxwV/yrM09P8KNWmXxthIkpcm9snc/otREr2uG
btauCJfZYikNznZtWi8mTjysbFhqvVktrZMUpvVJpltNskscBvjRoewWAFOdEWEXnqKag2XPG+XY
k/Uglg1v322CozGiygjLHQZfWQDCuiyGHljtmZNTVkzF2NEBlKV5b2FsHEv7XthvehAUwjzduSYq
JHGcUcIqfRXxdKdKpthTFG/DoXFwE3bh1/V4kULCKgY7MnHpHykkYIHPQIaL0O/IROeUtUxcUH7j
CCnqQ8tyIE3+uv2HZDeCgtZM1yhH4LvNTpxfH8BP/s2QXevRmc5KP9/ClE0Poi+4sTrhMbaZfWsO
d799UP+a8ugxZHY2Kkj0rwwfwENzCDtNK0so8JjIFmLx0pr7yNL8vudJq+k5t7Mpj2YMe/55K0v/
JlB0KEmJ0zwc3D4OPtLW6kTqmKg27yMYOF9ipjHLm1MgEMlLbk3qNzQ+RhkzwbA2k6wgaaKVzwXe
034ChilrJruXvZeLKcUjT+FVllh5dzFreAOURqv6pzd2N7v2VxsNNiUGJU+M0GxWPA4AQxjM3g3z
Qow9wNyD7Juw7pD1sd48bNX0tg+WjOc8H9eFekW2MRcdM3bosd6lIrrrrbaTXD9xiLuDHYiUa9/m
YiCKubAllCSRnYqGDpfCTtN/rae7aKj518KxA0ph03l2RSk+h9Q18WhVTwsxgar4RSkJZFV9/pVx
2W3RI/E9xy/5/SaDni7Laze8YnjBANiklV51snmG3lCVf/KxhMXR2mMLfB2qkHoFLUFhPxPD8/qR
zijU5QxmQcHiVqO7YIGh8QU9hvH5RZgCuhofsGpwybeeKsgC0ms86GdjR/FftjOFkTOtBwnGE1m3
Wu67XsAocINbZq+5FqJIVONCxRY+DAG3ac6Lwlp6tPT3RQUEdtdOl3ZjMFRuyLfGnssdHiqELTRf
rZG6ouU67V8Lcu7nf6FQRyYhnsppsm0trmkg7xveYc9dnwBYWYYPIOnu95wsAg4+UBdi6uUn012L
bIS24zPrD0vy/XBJvUM5jlKU9aQexKiEYCAj8tQ8W6UA9XiYyibtg/6Paw1x4ZmAUxPe4nBAOfna
ppAv9VWv9NHmezS46xpha2QP2vJcR0WbDQcL1VNL24jCj0Lj4m+NyK+m/XKVtc8AL8dP+cRNw629
6/eZVd1wjmV9peITD+GNi0SRj7W8n9dqWcNoR5eeDjqziXEMP9nves+9nEx/JFYvQQPkg2Dpcsio
NaOkm9Tv42iax8B4ELtkcFy5+4XLmk8ulam6vMEaFeXKgDsOMgOfhhS4G8GnRvJqcpO/q7B5W6Kg
9/1Uokxvga2bk0aVnNdc6wcoYKJyzcABEV8hfrR1YTqTEdDg8ancdevNHBVdwdWSGGlIMcsFQ9Yz
gRNUjJdWa8kpWhga6Hx7i5UeQq/1UvqddTGMdor3SlQj1vqj9VAFShLWMg+tmaNZrT8ZeimI/+ho
TdF1rBrIS+o4FVBrXBMXNSABf+K7bxiw8e4cne7fYsgRAt/V4378lCrPbgqHiFbEkY7yTooi9X3U
ZSsSeRFrO0p08Ik8tm89Gfi31CaM3a8/DcPRxpIq7PVRelO9rdUXrvveXIJoXfI9faru6q6/3lMe
+4Jfrz89m5mZSYiEqMkw/EzmYLThDttGBgKDIfgVZye30lR+kTIbqtqK8EwWapr/oDCqilP7TBaU
C0M09SXsde0tkH1irWwcGq+ifPrVedqcL/LnNKxAtbaH1f0VYYEfQouHHI1IbUuobPsY8argUqg7
8Uw4Yp5/fSN7B3kf+ZKUy3KwD2ThvWzv5v8ip4KsZzHLe2yImU3TjA3NduSVqyQ0cD72L43pQHQC
SuTWvFVNY2Whp1slZkDy5q23mSY2zv0ZyRkU+5R2YIjXbao3EiqkGCn+Y/BGtUAXAI69dd6jld9G
1ikJK4WYuq85LN+YFrU2qHgWgv1BRKecwUvcnI636vNVgTI0ssALW7jm543M2/Ocjd1mNdoBRKQ8
padNKoZPcnCEGZpwsHYZB7+7XyzOhnERTtTD7N527s6glJ5ahyZxWTp7W3TSbg0lZF14if94f2ht
eYF445YH7KvVNkApX2AqAixtkR9mz8ysFkDMYb/tq5Jx3jed3BOCAqL4EdHVM8fEyF5b8/VS4eEM
vPD474l1ZDKhVyTEsn30Ke5TigvqM0X1d2QjlLC9HHg4eHsNSolrgn7xAd9YRPCbUK+e2bSQEYzJ
NdvPIKGUkipgGdWC0E0LnPCOx7mic/22w7cIWkjNtgI8NDGpxPAMHJJ9QBdOG3MnqRc8bGun5Crc
xMRbQDmv7DAFm5XR+Jc4VPJ2wT2YnIukkMrGuiXpsYWAW6IbWUET17cAercZ0gpOL9Hxq0p1qph0
5tQsS1xq67dVN6F+XGYHwvOs+qxT5P1ROpmtlt18TcveNV6L1IWAV1l8ORHk+jm6/VYTcXnE/aJm
/pCXIAt3TWvJWHQ/w91B6KuCfkjPsZrbB/5NqB5bJXR6qrEMindQg0MUqondIjgv7BYwcui34h9D
1URDMkWhLH5bLxlHCeyQf8SIIl71zp2V0sh5l88hFscQhgJkcfUcD24v0Ogk0d+0apPRnMR9GPEA
QAEEbYadCWQ+bPSQTB+2FNKUuxbqGYUuELYrLfiu87qJJJSqQzFCuDTKiTZoJf58Z/Z9LwhegmuE
8ulEt4Pj4AahzmJ70WNySCFQO93ZeMOiNb+NYbum4KrAumlP1jzQNAxq/i+E6lRga5pgV09MLIFr
r3sf9/NEsQ+/q64qlnoeVMDt+eJhclX5aL1N9WfmKcCFt+2HbhNHfEJwRepoYQ6aOXEABbDa//eL
HOUtzDsgVo+t4Mjo0cMnViI4M7gol82T5B457sxxynCXPseE3zDRD7MK638XfAY4zNf9pLZRUYCo
Cx4XiBjYKoCrozSihCz+BbNAK0Enl6ZrCRvHRX1/uTZO1xOJOC57JnjfOlqziBKWRQ9+YxH0AGLw
7GiAl3Kfpv/O9zl0t+bJRv0eW2x3bHCYaYS4jjt3JQQsRuYw7YMXhRk+bR7FxJy6+4+G7MWXvUuJ
nOiY0QR8uxTUN7a6oZt3gajagy/rGYfKyV9xPGnqTcg7stQLaB9MKUYiUmt5DEq0IOVTQQaTajms
mEBd9N+UhSOfMCxlffgUfLsAkNoDt019OvnzrKukMuzaTNfj/CT3Njr4KZWuj4dD1WMD7dyIsuWE
43cTxtFJiVfEY3TQYtOd6RP82gBydzBicadbXZBlDzZeLhwg6qpiGckinihl5iywOzUN5eJG07Hs
JjAHuyTlXKa4nLiY4i8A8r2wyCma40abY2LeuHlGwm1vTi0Dl9iKv0MpDoz6kr/S21txZJv23/ln
tbGZNElDTtZnOfv3wM+R6A6/OAQb7FV72ssjAlL2kYL4gKKteDVxvBjCJ4I50lY57+OwnzGXxcy8
dcFLBgOP1N3AfjlwvarvKL/vVNG2hAVg7t5d4Nf1Y0wx9E0pbsM2d34XhRCW2b58OBg2WserGVrs
OFKkYD5QLyEkb142Wg9lfTZtGgF1CbAl2ruqlROvPe5WF9/BbF7LbG9Zb8P1EXr8mif0tFVm9QHR
ZsLIVLWZb/e/zUPrC/zu8Bj9bFtuXHt7L/yaLfLnaTYsJ5xVxB4dJqgk3/6yhYhTftscrFleIsxs
Q7oPI/71QRUmi8dxE2k4QaDShKl51eiHJMR6PuuF3hGHD7kUw0Icd5mx0o4qRb+l23nHlM2vrkn9
5Zn3c8kg1YPr65Wn4LHWM/+OqPl6CVwRaVXhpncHbV2Eah96MsHrj5I+QZDrjHsHCHR+JjuX54ix
QHSKmqImIpvj0tURyZbljAaQs2O/FKtk1163m+XlxyTxsVJ6pHbgbEnXChb+TIOdvAm6u4Pk4blj
asFflF8n0YLm43BeHJ6Sy/yf2d2udT4am0xzICrpkbV0qaYVyLJv+i9AMqrPQM3OU4vIxRPn3nMb
1OHVLDBJGvdQuQuidUYTtu+k9LQS/EzZ72XD07C0KfqjWziA9dLfAsg3MG2GCNRZGOO+QL/sztDj
MH2TxrEfiJqXF79vpBIGPXRnioxnpNMgdHjs7fY0m3UFd/YI9+nmjVzcvRjT5Ga2iOB0Sz+/JAnt
EHKl3IZiszj89hCR/X+1S9dS0SxQ8+Xfv1k527rKMbHNSCb4YxFnym5htO0zxv9d10vwyG/31r7V
DEM/MeheZyw2BNwkphWS7fsRHnxge2YM73fKjb9d0M0D0RU7VPA4LxT7Ksngl+Nal4KA+qNWtFdU
iDapV9NLtnFC/H5ifSMgZe04Tta7WvxWu4NSyP2TF9OoFRBtgYMVePPpMkM9SaakQS2Isjg0EC0z
vKhzesB7x2mniGLXEgNefI2YzyP/KjwuuAH3YISjcAIUnAPiD9G2HzPIfnBKjZoWEBFfxcdQjb5U
y4x2nBwvsSFT70VD9nzpj36+bV7UGPqjFt7IAYGQHn5iEViOMud/PPvKosvh5ICWdoP71RedS5MK
g56hoUHOqYLItJPnilHNFeKnWZHTvWfu85rOXMq2fuHDduT5GSTNRzrdsl7kmrzaXrxT7+bVg50M
WXJ8qqiip+iIZ96PghTiwFNiZsojPs+cc6lX+/uM5799ZXNAuCOZM47AKjosnCCNUq1J4JKvIyLc
BKiinDLedHPNB9IXCnVRUJlGmw7yxQbQ8X5j9+zKfPzMmX7ttl9NoqjYJGBvfa0AYDBs3k+737Yn
eAwVoGiUlhpjGd+Yx1Lf8vvrZecuUrz9dSOPywkbfzVdxe6Sy2n23Tty2GeV3wCPkXeo+a9TO5w4
6nteQQuzz5FftuBqlmLBfKpUpqq+0UsRqtolgkcHI+akLol8W9d4ouvw/qvCZzB2ab9O+fOY5y0u
HBHgbtU8e+QU6QC2eTAcy4B5b24Jk943FypwNEGCUjuOcvcHnyOiUXjrNHVAonYq1Ud4sBF41QFM
Dbl7vL16cvbQcF5oiaqqHPkgg3gVSsjkJaH5RlXzqInH+ChG+5SVNzbHkveYT9s0D4StnLnSzPoS
Q3buMcxBthazTOL4sb0YZqvw5XAR5TavvG0Cdqg/yTjgSC9lM0LmGACE11X6ySeKWJWV0qRpplFh
ALwNcV79wY83lTYL3Nx6TeohXnqT+F1aD4wj401nWqUNRktdjtpGo3zNp+KXnfnj3n2UDxZpbkpW
MVAro1dl53jvDkz23Cp8Xmqb99DfWc5riCkTehNWfhIh+mHcisn/sdpSu6xSBg1a1F5lu28Y3gJS
/tMPTPRed/kOOGus1sef7M1RHBiaIkT5tBwACuR5m6Clb/sM4IxjLYpkbiQ+pq3B8cYvF077OCkZ
MAOXBv0stSwlOgrgrP38rY+ScjbHujMl8TOPgcLhRfGdncXsANsrewbh1KAfw7f32D7Sk34wWnvi
Rope0Rlovk4RQW8bHjUYkdTcsMpiIfgrxQ+u1cPXdGzgQARZiKe+/1K1h0I48jNkUMCyM44JUdUv
s5X+FXbNmokF+4NmlSqqJ6H0m1cBhL/LGCFmOBMyeV8FSj/F1cyU+I5nZdrqbVl+pnAnJyRTrAZU
c+7W0RQX9y/xS+c0/zOdXA3AjXldY7JbA6vIJAfEqsFBaicS+gLdofC40pm7yWNkOj0Ym4b9aLrg
+VFd6op9KzhEhqDhaGai7ipPZ3u5fY9hJwTEqvOHApniEiylPzfSLP6zuiIPstzlM/Kk95jy5hyw
dweqSjkqHRtGWqG4WWytu7+1ZiF+gxHKAhANo/3YgAG/DC3WzOO+d+YmoYcSa2fBnxes/pvCN4Xp
h2cRUEZvVo6jRt+qcfz9Ry0phAI6KuKuxt1+pfQCXERyfMPcqL+Mhnf1lrnR1kuYUVf86R9iCS3v
LqSFy435FYUuc1gpX4r2gpaET8RshnFrolT+ELrQDUjgTLFvVTCgUHguLG9l4ZcTui7aHumbk+EC
AIdiNeb7VCFRatBJhQWq0mUtefvJIpbY8Hyc/yVanpZtvX8qnb9fy6Wnmim1E2WJTZRP+90HMFcs
qrVXXxpMpgf/L3Eh7fTtAb8KdOHWr/+kWmPniL6JGr3+liSybF9w9BvQofeqko9TWXb1Zmf6awcD
Bt0vS/1YETXEVeqvRWIBG1qK83/mvolT6Bmfg8UJTF/AoxP9Fsh2zvQJRv3iWJsUU/Rewf0gSIO5
AGxnSuQ2/S1GlrFwW4uqoHHnp8xW9v7uM+g/5O755sJ4WYarojE6Js2FwRkxcbaaQiMTDUdAXVCw
uP4/9epSdSYO9HNYlQfnyjvkz3w5VJiIMnwndJvN4O6PMeTctGqMy4jwmz9irEZIyy2vc8gT89C2
VuQnkGhtGaV9XCaFd/KJ5uCFC6m3X/YdC1J4CLzJ15ZMDukzkxq5obpuOD1cpuctJY9shalTeKxx
rMwY6LweEFIke8jWXhyxlPK8r4xcO/pCfsI61BV0fVzgy3bdBiIlU1ebCX/3DmtonMLsE8u7+NXI
mAXgSa3Gy9aH3sqo5j/SnQ96C/oBVezayzDLoluCyJRkCL149clORGBLtsxCEjB+hOeWIl1fV5TQ
kRAj3y04UOXad46vFQAbDfM/SJTMwwqTc5g9HEXsSKsUbXtu1zEfg1iVP9D9IsoUxX7aiiRDe0f6
EAY+l6Z8krYnLXAmEM+xeLvxA2cdePcrVSkwOimddLZmPuRQR1EP56lhUdNMqhr61Z/v+0qHZXNi
aSFTDNC4SGO0EtPbQei6P9fYUPSq/Pk77AKYNKm6DyqsYgd74KkMkUuXgj7K/jyMWJcFJDH+RP3z
xM1Oy2m4XNag+Ge0E8G5nf3x6KSqb7OI3PfcxzD3UlNp2za4ncD+znf2BMQXLcdLfSdCU9jVUc+4
rsmrrXLuLamiv0lmWX80wFe+j1UVWC5Nm5USxq445M4wzCetlyBDGVMSqmTIpeGRXp+3/hV5zPvr
/7pzyhSFGqrvRAFtTFo3LBdtKqnH/UnGWhARsyfiDWYz7+zHLproBjdqDFoPwJDpu9a6CriO0RJ9
kiUUR/xfm6qebEiqLrqre0ED5/8L62bzBZz6qfy4/yGmbEf7xa05qCwG8DZqWbnKFn1GvKgdvnuX
xCuSFRic0Il5zk+26AI1kYh1PsqBghfLQhm6g+gyTuxI8hkuiZK081E9PZSsZC4pvwox7Jcd4fi3
lZcw/ipvDlfVN76Atz/zBpsILXeQTFNHLDUqaEa8iYdhVaslDsgDQWci6BWwyGf3YuFIA4NiMsfK
W5jQ0yIdsc/ExJszh0vWoX1UfSx2oW6bb9V3pFYpFTd/QK+2tV4Dpme7ZnDhWBlrEJj8gsITIZT4
vRptaVGMpRxkcKeCksI7RRNsQ9YEa4GdTVtkT6idDmRq4T/PWvOnblkKjlxYOkZS+DGqgaSLu5GO
deSpKtHCr1sZ+jyHQ2ZJ6HuXN+ikgj4AfIS8tVVGOks0AB7h0h2vwFVz8DYueRedOVZ/QEwIrGiP
18o0T+XTctEhKc8TwQZGoL14+cZXFHmz12YCRyN7E3fQeA31bk63QS6VcktzqHdb31/gPJERCwr5
1IuzrVDGpflsJVNqHyOYR04GSqU4mTM5WIPhNYg1wAGVKGkD/HcqqWxZzqeBVJR0vedDvKZ6TWgZ
sqyBU1hdhyMTWm6pWviz76/TNTR+qzcd7dud8Vaf4s9dqk5dGTUod+73Z+HqwOVoERv0+ZfVV8CD
9gEHQ25g6kc2urJGpZ93FEXP7uqWeUZ8o+n92KE0bzN6JIbTbp50wGlpHX47k9tEn1j+1bl+A56h
YRrvjsc4V96EZAElE+wn4gHYalk7WlgRaGwZXud1fQJ45vW867cEkTHh9jOoyfcXDocb005k0Hkm
Rtkh1GHr984M6tIfAFIlW57xDjr4JIOxEUGNkWvIX72Mi4z01ZprwAaBzKsWXQMLsuh0wmIK7a+0
lc6TXSKQYJDBCKZkKZhLz7i7wJtMjH3/mSIODKULjx0GUkpWhsbco4i+osnDO/rlWq6vKO2Af05l
Hozd9EHmFAYDSE/H4gcMWrg3KCaA/60ql09eId7bb9sCWmrJyakzmtazJ9jbbpE4lsHk39lls1dC
P81wp2j9dPEtbWfy7OQtkz32w3f0sXgVYfM8YFzmHraqPicRR6gKffghAzq8nMKCdN+n3EihCNdg
wij2+8Utxom7bjH5bz9wrSmthDAsLkkwEwsLo/PvQG4L9fBrBuPUgBvS2B3UgS3bFB/o03jwO7wd
yXbGDIgVP765pLotIFvYJB3j4xNC2STIguLOhhO1spY7h3wnIqGyjnYW++sF9OoG8a2EgDtpkoID
jy0M/k/ItCdGnf8i3574Z+HAvnz51VSz2IfcJ+pl9EzhiaxeNdMNw7STH5wO5jdJXCeTNwWmdaPX
01Exb97GCFCpGYcMM5niV3sFmR/7BrSyKBsbz+/2povrdpBtIARJ4EGJowEEcfLbORNxZCsFjnPV
uswo2TTjYiWrGNb18vwC9hq0mc2SaIboQd8O59CfRD/kBtBJ9UBdEWtaDtliodlqfktpqtcdZtgV
vR2mI7md+QOTkhRSyGaJS/8SxIPHcjGFgwUTd6D8IuhzJ3iuGvXP/cpQSMUd+MiJJ3i/oZpFc+Wx
eXB05c0QEbLcV4sPmV8V7OK5ejbMf0QrhKSRCPrgWh3e+5T+EK3DGtWxAzU0KwG5TV9+HPJoKbB7
yQdywuiKCgBBwN/C7W5tw0ye1WKy+Cqk6iwjibkDE16ckNUI9Bo2Oie1t+qPzTKgwM6nWIk0ZgHs
0jEiYZT4gFrXTFDN4sIIQK6LZyYUPHDoUCyanwjEvNOmkh/y/DO7dXL1e4pDVZ4eU4lrQGpTw6V6
rto1EhLWtJnDHmTx9mRa2dULytiuqqP2ptZlDqnYkRRkK1uNpKMSje4sRThOZW8v3KBcHRlfGs7X
DJfJGsKs6zbJ987/UTSxFDx6P1zLs64PaRVCioW6RsuTT6Q2UPywS6lAmvVLQSu6WNkHb+mXctoc
WmEx5K5SYMxYFbkQzqmIYMFzEx14/LDoNYifSZjFEaiq3jXE/OAK4vBXN1FzuLzP/4eGWh7oVf9j
wZt3qNPNUzhGBPcUE5/bXOi5pi/T72XhFZgs/CD2oLSSrFINxAox7IO6oWP4NvkzW9URQuGTI5Kk
bwvxL9soM8Pe4hX0m+qx1FbVRaV6AtZayUqFLhlqs7B2OVTpwvgK469sKSnnE+8qA/J4C5Q87VDB
solsY0bCAdWX8G1t4I3XEotoqAbwkvOX+AjKKuFXy90W7ob7YcWW6NY+BTrNhBaunvWDCXW55whu
Ndt1aOMt1aUU9DFumJ3D/JyHSzQ/zRbOhWIbfLehVFk/dz+wSU+7IeUgMrjWI+ikYgufo+JxDWBC
7s4MlCP4M/OhyunCt5Bxcfef3JVX0jgjzQn3Yko9pxOHFKD9g4bTo7NXczs91Ks1JcrGSuU1jGEJ
LX0QcYOds+Qb3hJCwhXqva6KqKCe9XP4R2IYaodbWrA7Algo0klWl4aiSxNc/9sKD8GF5M5ickyO
lYqh3/uC97ZjZ1dsdYjtRPwsBkNz1bmx7y00IqbZLLS3+qK687e1Y8ta8mrwU5jG7TO7I5bkgnfm
aJk/fXDHGP4EvSk7vD0mJ4GyNKOZv+TJJIs/FuxFANwX0NIaxERCbXAoRJjMBctchXYnlylGsofV
Lz+Ekcp53UpPkGFu/TwuAAioq6KKkOAvEfe8VgjAptnj97Nd2qLsft0RG57d3auye47WyCudzKRU
Dk47WIjtG4G1PCE/XZTxwOBwU62WNnXR+Ln2DGj50cCVMrH7tDNVTQDrLIDQI7+ZdL46l66Nffue
KPiio7fLyecPXu6UdumWOhrfqc9W11UcnBxAb3obJKLwlxLYSqN0abQgTOljWxu1m+tCUNdy+sS4
MeC9+b+NPmk83JWOriBqO8KcRi00xmb7YFIyx5uR8CUyNFvk8nv7QHvKr1Au651ieeI2ynkrpOG1
9+ySXOfva60lK/ur4eJ02WONlUIX/YHTUBd8k9ZfLaRBiBubw2JrXMWBCEKobmLN9zF7ZDojgjdp
mDEK7jrJs3XaoioNeE2UjfJ+gF17LOyRTB2S6fw3kB4uvdqOr7QG/CMNc3QOsz1egfnnWs4g+pnb
s5NuXf1CI0Atc3CMB2Qo7bZBmIcBFAhuzN7/f/yq0ntbrbo3fipzBXBYDmwQC94xJpVTpGLTNhBL
Yz/mz8iw/luWloXWsKy5M8o1b06rk4yqsI6huuoJ9X9INYCy1g5yUeBgoe4ClIW11S4O0j4QK1NJ
inO6jRdSOERj9oZRk2RafgFk8lEDTPLZOewNiKKSa4xFNn546rxccZiP2UGOuX89ud+ioKf/Phna
6cVGwKlEMF3DSzF0Pif3CPJgNABFRZtptXZ5tEQavHv8KMXHQKooIuUS+zPxdEKdG3QvcY4GNv3r
WVA2pka9qjX9GB8IWw3lWo/eMHuRDsAsxnxN+hDNNA4UgAORLkvMbcFyH/ovsR4b9dqu09AJkOPZ
t9tPShi9shvWWaPMC/wli8EiOlGpdmTyhB2KZf3DAkMMzm09O80IGRI6F7f8QUTLY9Rx3R1b1hL+
6KLPp2pf1UNrSwwd2NOYSZOrowU9GzHCrz7L5FmPvjOjhtUSGslvsgNj8XFm3WOJR1vXbtSFmA5y
SmDBJhNxDhccpUrj/XHu5zGxule6/n7zkXmTJzpORV0qTRqszp2Cq1Q+UYXj9tEC/VYcQog42gRj
nogZxYzfc+V4KjlB0UErglL8q+nlbEVWhVPJQO2Lil3d1iF1GqLYXYfRdgux24xZQvaMWdiNr6OJ
WS0slupXDP6Wz2dhE5lv4MhfMV2lHL5hRvfmPf5Yb4bcV5HrNpkSaGbFIAmvpTDsfyaYnjrMAWZ3
GvzIjELQWnQKTIFM4YQZ9dLQAE1FAyAVglfcU1ypUXL4wSWdqkGVpwQeODdQkasZ/2/e96a6gpQ0
pHIo3MH2vyWq2Yj2yAWzWkBZuj4lD6TfzwOZBwFqgeNI6IEkT2Q7EQfSaCEwaMM048ZrTJvHzPYJ
OVpHGH4lThKseykwFoymz/rdXDJjxmRYIb891rcniGG2npsrMuNAZo70Zk5xa9NIXSUr10469l19
aUpDoRWVk/LzLcrtv8Ni9Zxf3F6iZHo/tL2/GEbe46t6g1ZeLLoeXo5G8EjDVoPnJMKRyVxOFLqE
G24CwcyLgk0kkCoV+hFyrXUJqcDDoZbmEHiyfL+DRQzpX3523dTPf2BoiMtMfkzfsO8WssBSajZb
LRQscDpRw0A3t9dmm6plvESpvtcYYGsQEVFLbNm/8joCd58yDaVmkacXfXogzSy23ic684R0AZ1j
Mkkkuybyp4on6803Gz4PrdBwP2+U50bfeN2CyUSzYYV2Tm3bxHIhv1FAMSs29cL3kpwSgsoQHKQ5
6OppgxzrcT357wUURHgXWRBK/dyvd1vnQJ7trrPCR6ylU2XLQ1MuBOjhFMWMlLp0/n3+nckw6Znl
ZzZp7XOSDCalopE5UiXJHNj9rdPue1mlbbheeDOSzAsO9HH0C5DDjxb1OoGu/wW2GcM/iZpHB8xZ
7vyCui+TjyO3X5Lxiy6WzR7eVbNqSGLX9Pi2RZMUX8H6tPLf4iTYfn87cesRbVWL9NTjJlrpyCok
aC1evfraatUvaTSbcEiGo8rp10VEh+mOqPpoANAC0S8t1pe3CoV/v/QH3ikdyMYrsNoT7O193oRJ
tt4YacBb5osM7hPGd8GXVfSVUOXCO+Uk7YhHyXm6ZTNwrUxQa0uZb6ccudQqGuWyquhXZQG8XjSw
OYMJKlbFKFiOr4mN+iSEr6TD+KvxypDwds3QjXRJIwJ3dEzjNFQdApCHIgKH//9mcqZHUeV0h6Ji
yKvmSiCRkr6uOhFoXQkBgI13f6KBI2zFZNa+3lTUCkHMFrSnWVXS2nCDPA9xXSiciVctyzvOP06/
ghqCd7A4weeulOjUpYVHrj/dUkn7irz5rHrJrdUYd+zt2MmX0G2++LVGSc2n//nl8A+WF0+H821y
cvyJSK+CYRKcHh8386QiiYJ6xRFVIaFoH9Bom46395mh8ndcMW4VxRT/xW1Mge4eUkIxIZKnIC0+
9dooOFufQ356+OOAbn/vebRFL+5XRpm1MbM8wO9yz0mJFEIcm4j/urdub+s3FO8FiUQs1hfXN31k
Uf5/iqXRVz8HhE1s21WIQ1ZGkEn6ION/b/xArq49MjD+Pg5KNEANGIgmSkUJFWXJnRcwkk3Bk9GP
kcmW87uSqN5N8IAyjelv8jvloeWc7dWYIcmzQr5dUr0I9UktUsKzIsOeUI3QXF9ZwYc4cmr9Vbij
Jf2jILPQZVVt1fvElWcYLtOMqXtAP1CpdyeYQN2t1+WAHgyu8JdGmb2BH5Vx2TotbW13yKxJP50a
VMt8yHyDOd6B2Yva+g95xNdqs1+DXLHXTfLySQv+ThLssFvFgd9KLMCnPdyDY+7w8RRQBcGGL1De
tE5/mWLDRmNy8xdPTNRhwqrAxb4eKAfy1USfTPKKF1I8TaRXxzIUO6hi7P+Mk6U6k5PnCaojeaR6
x32WG2jXQjPxV6l11BmokPyid+0MOVaZlMtx0jIw7SUF01dF7mjjh+O56aBV6kWjDD1qmjkREBB0
sem6Mav21NIH+EmSGT7zTUHkdK28SFKW1NCpO1YJWnLQsG2OtrHB9H3kFob3VAi87nWebc1bkKdZ
0gwh4/e1ROeiynDCVgzjCMvaO1Lxwt6EvLqxe48mzq6TYdtsl33PN8OgKn6+BMg3aT+x4qpo+Jut
w9UMaEYFJ7g57RtaEUZmnrzpIolCJTp3QUwdtx08iQRuXiSbb3IlFTSXhDH1gysLZDDkeyVy3xtK
rRml9Sux2vxb+BwYEpMR0bIfT3BEWCg/Mbf9e18EqjNxF8i109aKZJ0K5Q9EnRBmJRKV9PIaGyyW
oOTkTdiMslB4+c9+HXYFdRySi4Z3DGGTwZOn4pZwGgbCjdVGKVQ3slNR3P99fcCvIsCHS+EPy31E
QifZD+jMqELu2Tey/Tpb/OjNPBUtFjDB0XFlfV0e0tGP7vhX840IeJwB+8i/7JBVehK/2UilJtdg
uVYbwuRgJsxgd/cTbWeNksKcWlhibP+5gS6rGD7xC4TZFAJUFygmZ8HZQZh71CmylTY+ISukMzBd
FA1yTg6E39J23zWq03IDz4izOWxYHOPg9Nij46NwZOSDKni6R5Dfq4I+dM/+oDE3WINdjeu7SCV6
ez6C1BqRtjfzfaKBS6kxhSydLNJLp1nGxuxhqHGNrf8GWwjdGeXb4VZlqR1AnUk98OnXKxfSz+4t
ebQh0rM5t/cRnMKHV6ixZgXHMo4PT6ngcDA4ntoJNIu7DjY2SogOI6TfAp/jRqSlXHFEjuhXadDX
tbqKMBcHXK2Y+pbnUZkU6TJWuzppQP+OqyJqdp50VE7WTV60KdO4/uz0ZVnCTF8W/fMCLy+go+mF
Bcagn5s9r5ryB3ovdPfHS6r+DQydTK0ZfhbipzDGp2fD98sS3TOaUDZTTSuLUrVyZE1ZnLy+81nB
Lny8JUDw649FJEgKWw4ZY4hk4237uBtCGtPWsWRcEOYGPJ1sJhxR7IAxK1bKW21jKJA7OHm1Uoci
WLpiaN4cRW3MiGpVYekAvYDwFqQJM31LGniOTtjoPa7L+MAnhDezPVXSd5hlorSm7pPg0/z5aAGe
xToMU7/Kr1QJbakLoRxl0f0iJvC96uklkErU+FFzkDxaZJL0AeSgq+b1YfIKbhaGSoXqhztPm4hP
Q6DFPzJeHg/8j7INia94nuCKUGGxwRLcEiLDYEBqBk+LAInpsl8+mmVIfwbkEO1yvPOBpOSjAffv
/nhgUtcVKi1jqxtdvIm2iaUnd+hSxfzQPYCyFlE+gzMnwwcMFrkE/EpVWm/1id9IJo26+gJFjIqN
F3hSDnJH30fbPFLx1k9PvU5Cg0jNgavqA2QMqvPvdEeB9PVWS8tRyWy9AgGNjjKydDbTuaRSs1u+
nbOGrfkknNN2JjgnrNcOOgQY58H4lZq8K1Rw7TjwAFzBBE7FKDRUq1CSYVHObpmxW82XtwhTlBrt
fDCOSTeUdwCDRnOBG9UEv6EzFHyRTxZsGnmXsdJIAw9fxCK6s1A/cK9J40xCbHn4xKoczresl8gs
d/rtU9bnnWEvJbfmwNLoN0fHPBptjpUjyXdc8xvr8k4gCM1Uj4LRvpvH1+qIso60kn99ERPfEbYb
8RBqJCgA/m7oVevZBpC0+Lrj63bSiFHFvesvSZc2UCvVRYd5fk+GCDljTgYxeIhisBBVgW+kTf7X
rZddQ44C9i7WIcvn7kewVqonG0L5fZSr8s37zNfjSrv26qzwq0metbhUVVdUU0KTkz1ZNl9RKfcx
3yRGVOhC/3LGVLDGwiRPUKbzzw17D9UCD97H1XR0IhfLrY6O0Pmro3wGixqx/EWVxf8qdaTz1/Gu
5Co1GdD7h4LmpdBHVHv7FFNQkKUWiOHhwJcjp5ey4WoorUyL/n/RwFBZKMChSA5bm1tzLBnrOZpB
zeeibJmbo9kz3clqU21LlhIP6BwTDhEmOXppajzGyAw2lJAObp/286oqDuizqObboJAeN8gFo7Cr
e2QSuscjECj/FsqRAkki74kOtN9u/KI+2wGczjncmTzvfK+L53i38z8AKCX4axZl+NlUX5ER4S2W
2o3RdbIjC6nEGRqN4oWwwvNi6yqXvva91HDAmIWWmoOEbFz6HkEysJ5imKhmDyi4s4MHr9HjcCSd
wRkJXyKB7TpgXAZNyIsL45koUA7vuzNZXyAMDjhj08HMlQDAs8/MLcea/fxvIaawzXDmBIUvyQN0
oD3+fAzSLDFtVk7laTj2H887u7x/qa36jnFzUoaq6JiuG59JjtpJprcIGuM6BMjY9068fzEZ8lKN
0y80BwZ9oy9Iddq4eTFtR3zghoDRe/0laGxYjIzpzpj21cS9IDwaulXBaIrhvn9JQSL2L4zMkoiI
uU/x0FP/AHM9FHS7diFdT9y4M9N1M5zn6Q+H61N8MzstMk/vATHTV/GmlsgSH7zstUgRNdgICu52
ZnhkVoNyloQPlyDZw/EeIc08X8pkwi3gf82H3Fmp3CUakkHP38Mh4jjJHH6JuHLkjDk1iBYp2Y7u
4lPjWwW4h1TyDzXfE9Qa3inhazE2eTZC9mn+5u1NwgL/D1ngKLwXS/UHoFsktOUKY3PYuQPHWcAM
RxmsQLG02XKyO7kABb+cEsdG/Qn1YxYrp1tSRHtO/NLwBCT0nRftyvoTZ/f3035boiR9DtUQNP5J
BSoNWYU5S14lY33u2dMmSroUvE9ScHr/oPN//UgAinQgZB5NNS5sUyPpDPxtT5/riE4nfO4S18Hh
GY+xKQaBam/vjl0wyUCOdBII0miTLI0DnE31reW3YTGsI5amKkaiPetyyf/1N0VXTWfq8gvM+d0o
6vEF4iwqEgRjs6yRNpDnpu0xeqV2YQpj9SbGcEK31CAqRvyQeIGUXjBuBIZke6XLNNvEX9+2YAor
rV5EnUs4pQa11UZ5rXezehvDWmK4ZXKWiVUkKqzR0/bfI4QyS3xWAzvTCtakkBi5xVuzKKJ/DzNt
Cx5cjQni8cOeFFAoxJVaHLZnzLhBx2K8jzLhMXc8lc6r0Sq9g2/gqlbmKBNzfK9S2wCZAfnFLm/o
H05iLgUX7gowWkpL74msWIOVCvKLH/eteugPV2lq/gRlCbloJHrBfqbaWSmrQIwtNQzqK7yWBvt4
zgvBM50xKhWTRtBoLHmasHzB1Zdzg6AGKeLz7VlqlRthTw9ecPkHtA68CdTayN/CrNJzaknW+WPv
fGdYB5M2rFbOgUa4QZ6G2zSfIJmxz0A8joXXpBS50LMTqmCofCUMhAuVvzQxF66AlDUK+RGtiS6u
F5JjsY7IRW7CRuu67deRvbsAy2wYpSaw8J15+VZl2kxRPN5jEsYzf6iCQ+FZX8qcuwTyAjvQvnmk
QR0Otf8fKMIC5byx63eDLDMOPCdsJllKKnIinegr7ED9E8hGVC1w1cC0XllHHlT1IImW4FbioftM
AS0fBfUyReo//Dsux0kaK7/mFZIeiuP8tfdd32EowAMNKTAcIGOh4hL8dBFkhvCXoke15nYDq1yU
HdDd+jgXGczJwRyK4W+I93nTzxSUSH5kVV3Kxzs6s3Cd4hgZH7IOrRi65Lv8+27qfQPynAZxUFL5
L+M4BH5kljTYM9B2td9Y5XcQ5lyl+gQmZ9xMOT7JFJKozoQ2mtclVxw8DYzBrTXGrSzbAAagllkF
+pMj3bz0vvs+x5v6IGhPVpF6JbBlxNRQcLZ1Z3BnS6w7Lx9MQoux7jNAe6MP/H1v2YM2ROWuYJqw
Lzi3a1hgRip0a3gIjWOSiaoKxavuYT56PPumGm9uP4Giu5sjtcMfP3lgpMbufMJcglyZJ3dToNE1
YDkPkw0dFLBRqfra60f57tyclmDRX0SqmY6Vd8YgSM5SLyivYIuFjFq8Hj9a74kAGfBGyt7QVBTS
cp5o8UOBeDV/Wq15QapFnugAky72/SEi1+46JvBCGmX8zte620PxRZKtnsisVGU4953fqfozfxxr
RNYiJCCV8icjm8yXWzpUeeD0w0l3Qj7Si1orJMlPZgYlxpluQ3fd0G3Mo9SQPRpscrEnbQ8WLHey
tv+B7Uc15dHsPpADpLwNFcbrYqY+GQ2/j5vHKOTpNmEXdqBCcXZF7jE0JVYDlV9KEqQTh27ae6lp
D19Vm2bf42SQoJFRtyeVAMtGAcHVBdFhik1tJUN2rMVM/6B/FrQFx/s3b1n8s6NJKvDmbCNpMwdb
V/lmzTatyruVStTdP69LRFgaWf1fCarzHTlIYdWHDekIgrNZfadcTjIdxiZPPLK2BizuX2vK0chj
NOJCInE5GhQRl7rxfjbDQUjOCTV8BCxM4pQsvTCQnmArFFa4DegkfwenjeETVXSKSbabxSkCydzG
m3hLRXqS/Sh/wJONZXg4xyg+qfwXcp4RV7M04yJchnJikrRQEZXsXqzH0RzlwyVc+pvgZ+aPjbgQ
oHI5INsQgs4L7jVq8jLhZYqd7pIINo/8INw2z5mg54Jc6o37Aoxx1AsJq9hp/R7UbL/kM9ENSdbY
LMJjMnI8zeoDoig238RHHJ4sHQbUR2jsXreSfZsNCVokIrZrmrAcagEAhoSJnSmbZNNpOL00syvL
vqaGz5tALCweX/ea8qt/LR/B1jReqlpPrRl12FMNNzeGWSmh+8b7N+VJYtdaiouGPyZQEhrRS5b7
X2sJSPeCmzeLK03pYH0c+iyXBQ403X1qIsdxAHnjn3Cz/nTZC7S8lIRfLRutK7xaW40u9pagonW1
VXIBw6amt0Q0lBokykRzUTN+9LQ/qD4ga9kutSBUBR+AriOIF6jtoKLnDyvClLIgk5PhVBTyf6Ue
VYk2KMS510YN9ZMrKSBQR5KQQPxhR9gBfNI7Ga9jv4jz5TLwg3efyjzL1G153YyOagUTBeS8CRCu
/KDIpNtZpJikjLFFrWlskTsv2IKAgHNSiZqGpWNLHLp1cbnqorj3Ik7gMlBxZI3ZnokQIJJ82Mut
40DBuPl6roPjq2JZs+XzZ2+wezlIqPOsmCJ5VrnWZe6XC5G6t/YbbJjTW/jjjfjO4amajb+Vt/yj
9HCBQXdg/79guXFXc6dNsltgaXr/wSiyoHbJ58dIaT8/vmEPyKEeYOG+45W8VxuFHfk7+T0cK6By
rATCeLTFJVbhseL2DbL8CCrHIhL/64R24bRQziBN1+693R1CH0NkfLncJgscnvBZ3IUnZkfJ+RcM
mmcshkQPDLYAedVUBdsCfUSYvUAyhotoOT50SY3qcMxls+9u0PyW5OWH5VluN3FJPA+vlb8IUSv1
UISBktF6iPqM0zRyIHkd7hin7U/Py1hrU2gwE0gUQf/ug8HSrg3CB9FsCkNpyomDwXnsi+MVmY5G
8AtH922S9QacImkZhnh/gVmzYGbx5XinwMi6TigMh7K8KoD4VSouDDE4QxSoKg7UOP3M++VdLTN+
IoAQAaGx7NYVcIYTCDBkdkuV103cmzhO7l1xKzfbibLS9mIyuLVBgJZ0/G2aOyBmb6eTLw/knkN9
Oow1MiQ7t/q7ksNmynN8BuHrMhX2u5MTelhMg+fEjYh1RXFhFpXOx9ip1qgw7CJ8zBLRSGgyFqeN
R4/cVOT8mTN+OMtvDVI9S4dLxyFIvGE5rbnQ7ZP28/G+9v1iwu7c038qwcu7u3mIKSTMqkx/ItAq
anlxY+twyTxKOvqbmBF2HLbwhhu+pgLuG6XlvMadzXU5ShgqgpURazcAv8nFLDrEEM6iS37kwrS9
LpmfyJ48X8aXTQdumrovSQPAuq7lkpjdmyLhgCIMpYMi5fOMkQBQRlQUornhCWIohkQsADX/o4qF
+RNsmzmGBT/UN+FjGTGVvL7BuH8dWriaQPKzZU43wdvQ5ooNikyCHXL+4rxRy01WkAdw2Nli6hOA
UIrogQUFeDwqMy4X89OtFEjr/xVQW/0Xwwc3ZPFM2gWq3muTaD49IFQwjMalmAmiV9RA4Ug4YVC9
ovqg7GpLeulDqb0S3SUnI1IjND+7BkQ8gupN1OiRZNiRD5Whrbg6uawGWU+vhPuZaDo+p0+qnmle
RA9vBnZexfIdyrafqmzqgdYGyKGed1dnTTx15YLh2ZEug5+gxRZOurE44TxYDP+iJWMlgit76EO/
aBIycBFBFrk0bSnWS3Qqmu2crXvCENHuilS3+sYNtWQVL/xt8OA4tzpTjguB5RSegXSe72dthYxt
UHy1NZpxgYUgY6PoXornBsLi+Ue/ehmoxAB1+wK7XIEu1gmgAUw9Xx21H+ziZxnMpcn7C4MJa/j/
28gVk1tOqEIhRx8v/bOD7BYBQx0U1dvIvcv8xh5MBwGXERtS2uBQkned9lzbUEVUE3swNIe2lI2W
MT8eFymkTP/mKeRvGSAz+qqlOVUStmCNSZhKzduko8WyK9gVXWQfhuGYetIxk30O+I60JQA1Mf7Y
4WZhFceKIWrguTG9zhVcVRl/SGZzNzirhYhuGNEYalhB7UXCTBFaS+qH/lKB4vTx474d68ujj/CL
80kSSMNX1wUj9Hm+jcQmpsEnk4vxx6Zg1ZB3DREwC+xPpdW5vTCKaTjrx7GcuRsA+tFiesAZAq34
jUMbJ6/XvfLQgKf+D5g8GASUPsa8B+tTLkQdyinTABwUx8Q6Q5OKRIRkIJkiQUDSM+PHp0VbTjdm
JdWVVyu9lnDWOAYsuuly12xODRD6DHXFEi+kkPsi2O6A2C8lBXvc/drrUgt8L69IGq5QKVlnhbW8
juoMFu5rtoAFhZI9L88X53zhgZxQ+6UFU0veRzwIcPbikV8a6lrwwu+U5ekHC0dvMDcG/+6p85Fi
H+SOWqXuwKJx1f2vtRz0fZA4oVk8/L6SRUf3EZmEIovyCqZaTDkUU2qmmIof2TpNl8fqscMEjITJ
kbOPJzjGE7dOdw2M7Tu6Tge4qr2GJSsWVbwTOpYIAtneZFhSfaLVSe60iBtCUDOvSQaCdHXNnQiN
sw1laMCCrrcyyOoecODjrdtIbXzJjxGnRG/AF/Bk1Rbxz1e1O02L2VKXu55YsQjN3syd494bI9xO
WuJduWx4B6SdVST9/SovoCCi209biawo6MUkz63OU5g3S9BFNgJIZMZWWBNRccO740wg54X1bptT
GJnXqsSD72EO7TsADYXuRcb3IHFMv7AVoAPb+uUMYVZAFJXKAd4tBNkPt58fTaSEo/bgiDiKIitF
donVoHIGKIQf4eghlb6XuFHjgftMc5aLcUblz7Oe0kCMtY50O2EHGteyiITObzoluAYNsJOswHxB
+q+jOuu5zGG8yj6wTI1VY7pA+9bxFDOnl+oL1JbCTqZnsKLfZgnTtWA1VTVreuWvDFH9OKlwYeFS
6iu1VepFe+QIdkeU4vzkMmRCLMqxywgfLAmiMA8gdy/0KRzX9bH+tiu4jppQLscc5/vKrArjGREj
Mg3p/tq7Naqa4YBF060sf/SbqOA4rgUFudkETNV0qJUS1dZYuv4ntS82KcqPrMEfLYt00GbaPJsz
5E+gsStwHlz1eI43Rqrk4gPi/BIohpwaAYDRtgtFJZyFkvwzj6FFb6rdWwy0kqU662wh8M730fgL
f6Qd9ljT5AArk95CEsZ9As8MUYXphAAXbPo5afVtMdKhbFeag7gcUlInOmc/IaeJHYj0ZQbQk+3X
m5ENVwYQAcS5haTMV9IXkDXgaTZqxZ9mo0SPkBoxe/9LpbK9Ul7Aq8dsFcKNVJ1ks5pxwsNKudZZ
bWK6VvTtyM9J4NzrrapQu2qn3ZDeUVaVfrd20ChrfeWiUUoNLdcG5N+X4Y1VJlfyvz21I7wYDIhx
3qQFgyE2eQ3v3y5QBwj1qT16SRKILpkOuadSGgFqgFnWxbVe+/dm8B1b4Ma2d0Zu6Li7bodLsOnW
bQpv6mkptGYAeM5YGSJPVXpyhuQqFYE6Ve26mLcSwFc7phqRwYLhBhhsXBD8SYqgtKiJXp7VLemr
M7G/30qKx19tQAX4vDLMVw4u8b7IbSSC5aNbd9O7nUU3pzYZT/jCy27ecNfdycJTHX43BMxunKnw
aTG9J1wcClmvRjrWO9WVIS1gyzo5Xh7El/H2+ooZsyTyOXsi1SczTLAB/NUFJeVzD/qSWpS5T03L
axrfRpv01C1oIB6optVLRbvTPdCe9C79wJG0d9tJOV45Y2aPRxuuQGng6sFPQa6XejBBRXXYDE5h
9PD0twedkbXbVvbNbaHj9/oP8UT0NvTfjT60kq/piDbKGK5g3PMwL4H2xoACeXiCKsJAOQbWYRvN
+1579zrZTkPKrzTy3gW0jnj83PWBulogvRFRHv4Ejof+2YERqFY+UMaSuGoZZ8C2QDA3OfGTZprt
+rq72QPXrrnllwzszbbzAGDiZozfMIkYtMCK2AWmHT8llItsRKdOvnfdtZGlmiFapd24TKw7iThJ
MH+KfFJwcOleOrjllmT7bbYMHy56wE4n4B4LgBhoXngPfbY43d3FZQifX/KrHG6LPOqsQKJo3dYo
hHOu0SmLxOraHj6M8hiKNcl4krk2PegoH9BHrPGiNOiSnzAkQ8iC/jyQNKy4sxPHHDeho8U3N7Hy
E6xUON6qLuFtckSSEbxFcpetQGP7tu1Y1fMJ2vUnVezQQvcSgiB0zS99b31aPh2Op9NzPtm6tx88
RKiKWwTW7JDjH2fP+xRQqqvm2d7Mt/ILllTTwmezoKP6Q2E/RDGahsvW8PS6PDBkRpu2XO2PLCwv
7CvFcuU0uX934eWE5gxIRpPza7erX2+pHc8UUfGIkUTMZWAk5+V0eje6I/MeRiUtu2Jd2KtJ/Xok
dTeGM1MUovHfBfYXz6Gti9beziizAuO8jvfbUUVl+EuqWo36UGzwjv1uzvViG9l+Ao6tVlBv9rPk
ob7DqQHOxUDaTc1vLp3YMGdVg7/0y6/Stx8Dv9iKKdbCA4P9dbLr201cU1z4/A5YM5y9DbP0r2R8
p+MT4P25BYLrV10e9TnHYa+rtNCFFmccT6CkpDmdUa1AYKwdcOb9XdN0Gb1QT5mw3tRwYQ1LdgQN
7W5LbS7pX0jtGPX3djXPKeoVP7myyV+2G0j6OzY9pE4DMac3/8vDHf5iqwMJ7RI3YS7BwGa4rh3D
GuiSQ1ikZL9VRU+duDvcvUvLgGcDDEucv5exbvJW6/q+KnP/k/P4Jf2iGv0VfAaqIEw/5w70eB3x
+LjO9TC+fCYBgACTSurl1hd36PAKUZq/2XaszjvTa3EvbvfgG4i7imsuhe8I2xCexDUYglFTqrzI
W72TVnmnomhpoT+gkfcJx1Ck16LYVN2NgiZabXPqBSWcxU6SC71FKG90KmXfooYtSpyo2c4eofBL
CPvMyZb4xhiqJPahLQ/bSSEQHEj98BNZWYPxow8kniSzhNFht9PLSoofbNix8SuBCBzKUn1Ha78O
Qlq5FXYkhhmthDZ/aFxC85Xa6SM4Ti5VCUSn57WD+halJw/7lI3BIFX/LD5bGAymFMqid0RDEYrf
H1EqpgfqCu41INgF/Wb581M8W7W4eUg25iSWYyT9L06lNgRetZi/j0eYDRLdbbDypNsSrOAZQrie
fOVQ+ns90TnPOz6BYwU6ttc522+ioCnbhkguzwgWaDMRpTp7jBL6jqSPdV9a+MSdW3AkC9oiFu7m
Z01Sanunao5rPMOB+QiI+o22VUnKY5YVsjPEVsvyoavQysPHD7ubsQCYr7qg6RHjvkU3XEyILxCx
MKKqNm+EDxBLUFAEGYu72xlTI51Zb/ZvUXrU062U4/KPN18ubYNQCw4+FRLWV9F1UnTETasHA0u7
XeqzLzB6iNRSaT9N9rRUFSnsPUZb7rmqHutYRHQ/4m9xmV8YCsxqKRiE3tXqg94slXcv8lKDB3fJ
2+CrhRloBpX+gO0k8FjCAZLsTb/P00ZrUttDoaPyJoodepdi67PD+eNUtPSxIAoDWeSXvSEmf4zL
WvPSKwfZBz6W1Xh7kRhxe3SQHaXLTWxwKIbraAfUfqjusuvx3hZ81gqnqYCE0rNhUHmJTAWl3lEo
PxaDtzAfFziLiQFuXTUXDJ6v8vge+t+00BMkkhqwBPJCaujWDfNI7B4vOUxU+TmE8ceYYUpYGoZc
XX7agfJmZjT14FsMVsPIHr5JsOKwy3JMer+be7dthVrsA7/bxKRGRpl31bKYy9OWCGpVlcweA6Qa
ukNTCzYoBdujbQJWSteQIjpWv/+uthLuzJGLu/LvjSNQI1bttizjevIah/1XtanorcFHNP79K8U8
6B0mMHxKzyFGIE96h0RjNikklZBoMTEungPKamtF7EGmtOBp+zDl0hARbkMQHvBDIs7ijjRZ/2w9
Ui9sZeAzXtRX4dIGAsBQB5vVRBE2VJf7m4zpr9I4ZovTehYXhBawhvkfJYYAokhTpguA7jSKqhqk
NIbn0CUAiLDc+Z6UDNyBdmkOub9SDPTBR3M9X+o0gc3VsD9bpFu89rPtm4Y5fiRhn74d/HeN1xF/
LY7rFBldS11FiVa4MWuSkSDSRzuzAHui1FXniUFqyCcILAjWBrUK3xFksG33uz/YkiTP9eCHTLWT
HwJle0qcKwtvwHUr7iVec+hPMYPWzWAljOtg8PaSepmo6eS4V46s02nMD97CFwPoDgaKQ6UdLc7A
drR3PJi2XaOc2FLBqgVNG1haawSrhg7Kg85b4iDpBiuNu6jNZnVeQaA8aDSNGNkFzp9hiJJwMy8F
BkFEgtpfSEirfkTqMOqsNTUGngygOHFuRN0I24dQD1rXRKxP3KHSHBEZ3Zhx6r0YMFGGl1vg5oRU
IrXA70NIrIVQbMtLDQHOnDPkVJamLqyBKX5SlFKsPZe4ns50U+zJGPO2UsvzPCkK1DKEnfW6Rq02
d4zr2thcpZUW+VxVxMSKxqQ+mvj33x2xSjcvK1q5QJehWJ1GxLuPoY3CNkwqUJ45nkseWPl9ReMS
H0OcSZ2uoLF/E8VJQD1JW2rBvVxvKbjiejMjtyRDgE8CdTyB24qmBzqs4e1Lw8nBBTKRdJ5EgI+2
KhOfEpAsL2FwgL1EVkrmeLk3tsyUWxxnj1S0vczZv9oBtqp1tQygaQBPzYtVEh1t+/HcC5sFdQ2m
vhWuIlQa6S0dzyy8roz8kpiLCt1S2HOuYF2PM011s9tJWWXBzl/FP8x7JF0kKbmmRnw4V2F05OvE
a0FGxN7i80k1/vWyDm3jFWhhKMOG2+8FMv6kJaDFeQkGj0ClWXmQPuCE5mWEZ+2Oae48Zj8uJHyZ
QNOx3x2VJMi5AMe+/cO7MrMZpJiOJmk+TarnjEBPFyYsBuxWLJg5ZV72CHj4ZBwSgSRPW+4oJfM2
QOKSb6o2YJ1OL8FaOeKxUzkJjZVsXUdXGS8RBvdqFT6rdM4gi/OfAbnv1B436224dHBLA9fokdPg
TNkLkK+qYNJ3lbzcVTM03+Fa6q1e85oF8NL5hWPyN2EwLGoCgLH6UcuYxE2dfF1A1wlIosL4QQMX
Ekup3CWibd2MPvekC+RS9LdCMAuGJUHyAfa477rZgkVyKbikWZWfgjX3TVyniLnJc3tiJOE8KT7N
OUA8bXmv1DTGuzv3OF3FeRd0Fvz96JMMtzFIsdnVgXh2t+wpYR+n12D4sQ/VDD0sK+/vClAwh/vX
8Ew5z9AMAY9Fg54ByuGkvsa0oMHQ57J8Os67SIANVa29uc9DdQIzARU5X1IbE7mW9Tessl11/2k2
5wRdi8GRT9zpUYtjXkxdJrGuGJotO1hQIaL2E0kFliiqjhcve1EglNM+7LRBMcHB2ZBaVHOh5m2n
DDEN68JnmABbr6sOtnQjKB91VMg5NcviXgYfEdO4rUvndTOGgnkhUGhOx+vxf6Mrlz2rPBF7OzCp
ZQCLTvuZ6JhOQh979Ii+QHs9ZM3K7tDmH/UYoxJMBkmMQcOrZyKRZ2+gMpCGGjbAOjv3TCxCJaVZ
qpVbkbyBRYKD9QwHliEW8RjuXhCZdW/3i5FpZU6dmA8c5bPEVAbySBSu0/PkE127IPkn1wn64uOs
VAaMD/6ccrjxQDVplB105F+LFz2i/AT3HFZQyOo3DNfrNuBejQsHwdFrj504tdZoCdJ9O65BqMhS
FeD05OskdbN3zeoGb9flE9DBP4sqt8DVa4SKCuNUxTCiVDuQQmojaWOwbyLpZQCBQ0R/RTzAuO3M
fTN90Trg5Ki6jLCx05E4o3nZt+pParOUw1ZeRqi7d46yhIk7e51SzARhrm61jgUvSugQTWVNEBkW
dtRqwgqAaldpR5PdoTOUpnq/M3/f9wFi7UjJDBUxZ8KvNb16seRu89m8wSCSVwxjCy8glvdV+kRz
yUjfQ7fZKSrJbNvVMz1M0XmAuGob0OsKfdYSCxFWNjVq5TLG3he+hdI0bHgoldVSW/oBR3p4uIyt
CIDDCpTuh0yuRsjcjCALC2TWI2ym6EclXvbh7jqdr2SI1qrn6ZjOAcP1miteYvmE6WnObZyaptnT
pOI18HDDz+awgc+52YyepOVQtJez36AAN4xtMxF6RI2goaLSBY16tIIRRnNio8q9XF7j+o2TPcJY
k5AlNzH/KOnleoh4Sz7qlm1MnAycRa/ZY/Es1wweZrdWdaiPI2Nr2bkPxnvrFpvKSdNVDUnNmRXx
4lVP27zhZb1udw1fsg1hPNQYKdo2NCzcy/ugm/v9teRmAsnhkh0iR5q+G6BeyINpw9ziPNjrDOGZ
yp39s98agn+y868Z0mKIpBCvyddx8nHjmaCZ8zeHMXXvIozJEl8Vc46bHvCBoG3sch/+Gcl5MU+X
XJ5wqB9+wck3tkPnrIGxtEeYPv+lur2rCYJ7owKXFrUJpcHTUvIvfLWfct6ux7C23T09LsCa+zUZ
VdflcDd8OxXmSbFZX7ici263s5gqCjGobc2WOEOmdbWmjwzDbIm69AC5qnwyn2EIYkeXTtG+QhjW
1h3MlL9CdoXVkzqK/+0KuCFUkYx38H3/muK1NJIOUmD5UuyMckhJyyGTVMXnvJoXFeDFyIsrpcMH
6C4PWMX8T+56wpf+bkKgsTlmb99bd7JAQtKcnvE3WpoSddcNU5kQMDmusl6rm8LPb+xqsuZ8fvME
uqnRLpAFU4V9qqWrvaAsNzeXfNfjl8yBdYfRuBDQ6GmKpqj5eytj5P3EcXoF0TJti8Cbazh9x/hx
znPiyx2GQ5lEFTSZDlpTuL4xKyw+baipTkurqXkBEEQI971bBxzzFMXZJdB02lEpUejqghvjSCWk
5YCE6N6E6FIPRQ9rYOeoFWY8XDGT9UJBmzmOnE1BtoFFf4PnhjhoWVKhkCY8SXwxHUDI08tRyhx8
Zs7JY0r6ZhCnI+M93HpthjJXGcnL+v5yeK0CIhGWNSW9INfzuymvUl3y0RcvfJ23RlE/WJKUWwGM
4fNXilFKK2DHwpmK9XwvV+a2kSZjKUq6xilR5jz16Bf3kHwc97FK+cqbeFDD2ta01haVB3+k/oTF
hJwscIrMjhN0I8oULmAGg0HzfFW6zTzvs0hT+UPw+i7NzoT6RlGvM7rTlpvG5nKaSNJrMG2FhEg+
yuOeNIECVxChu13w+3qO+aGpSkuTFeeq+1qV0o3ar44nW6NOS4MLgcUSXXTk7FwQpyfK+T/d5jA9
EGG8NNlJ8Pd8Oy5y+jvrDVvE3ueP/IEgUDSSPD2/GTqj2xTc3ltozO8+4Qy2MHvtj5z7p32YeDjZ
CtZu53V2U0l+c5zRa09BULXH5kK2Nocm1GyZcHCwAm2HINQ/Lq1gIZfpKxNDd3+8NrXj3jcc+h5W
vKx3aYwYwnCDDSZ9J4tsqOElhSyviTkuMNdACsYwJk/rCdrqNCw3Dq6VcXCsxi4KGupkbb6swN0R
+E+9oIa8ulHfbhHHY9s6mOuQsax5Rd2ITGg94Y9Fz8vQeSnhDsBVbn2AEO8X5aEpc9yMR0k6mj6v
aKcS68as3RB6MKCeHioUwlcl4vygI9rpm6bacFY8+bQTufB4hnMTgsXwl6PjKR76trRXWo3Kur6M
b4YWPWe6pJpfhRU2oNPP37MBs8m/DsVAQMT7h3w1njwxla0aj+hmWcX5u3FjHTJCxBhM96vPRBSI
4sHRs/21arjg0rQ0oYl3faZLJo4GVVWiUX2XdKy0JT1VoRc6kbq5sZPQF9j5Pr2rXB+LR3Q6+GBR
05ZJ2rPMFa2IsphELIuLwKPFzpfp9xKcnRGuLvZ2Ui7FbuVRd9wWrcHcSRjPVVo+GQfx4upIjxPs
YDLLBPYA3FR9MxN0glYBfJdegwf5ALKwx255r8TlTTCEWCLzcIsTSuSs2Y5fCi7qokX/sL9kZAfC
a9pItry6ckr1rwwJcabbcOn7uPWRl+yP7RXAJXs2hzIILgrvMp06bBtfIefK4u6kKbRUoU/+VmAZ
ZPDwFe1+k1Jq4+eP397c0U8gFQmz9qJ7y3JoUo73S8tX8NX2ToZGxdEo9y/cImVflfiQsnEEVi2q
Axh/mGjWLsPQBmEG9WCzuPO2uYJ24SaCF9k1Y4VGUB2gTOqAza/69dGm+v+0j1nBxGgQQ2SXYwAv
u1YmvzC1RJOTkZ6gD+GJj8U0zPnSLaPj78mEib1uD+8l7u7hZBUVBspXrb+HNvkEYzzId4zc8Mix
l0qzKWM/mhNnIweU8n5s837ySIYkpMEcOhRoTCz7LRg+r/xbaucRpJDdxpuFEoxnZpTzGKQEgA8S
wUXMbfvghw4N8/ibcfOWbOdLKGT6FSiB8zzmIz77ZPzutN8//9x5C94YrlL3gF2KjXYn7nhMBy0v
L5CgKo82uJ/oi3yRZs9RI01mi90oxkCHHDIzBoY0N7HylpgEWL38BPMWYFaw3rZp561N+g0a/y+p
mC9yg11clQs0Ga+RE7umi+s1YtkZDQvzP17+kdXmIsVNClORDX2AQ4XYqUpC2P9T8mqFHKq9a3kR
GQjy3+nQNX7yhBg+rtuWoqhRafI5Ha2uUG0PxUqpJ9QHzjqoUaZfxV7q9BGigYjhl4YFocKcrfnk
5+hQezk1EbN+PhSj7Qu7DDnJn9fU0xGFuISeH4gZY9BcqaPlRHH0KowfTS4kQEcQbN8cQu//kWpl
SSC6SEpBaPDWnSuEwMMrsaidcSjicuOAPGPxVjbX6zKbxkkdd7Cyt7BBMR97i+1tPmuLeDJeynww
p6Qq4L1a20e8WBC+TiWTR/fAuvlHIh5hAYoNiVHuLS8nH4ya4aphfkn7RGC9vODXRd+P1xHglRR5
egfuh5Qfg9Hh2u+/8xlqqaCWhOTJGQW2B10JsHmSpY3dZNis7GdA4TOCb2kRd2JOkO/AIKVQ6HBO
ZdlCASqDnYoAVVUx4pvzrs4Vwa7QlV8Ebmo2ibVPNuvOra3Z5QqsTdrO+b7wpUW7dveNdIbzamDX
qJTObRPe1Ue0sirhwHT7zPFm+uk004tjfrfmJYP/be65qr3Wd/RXacoCO50iCHk6Pz5l3ILtO7of
3GYiHu5i64Q4YIVBjCpVnGUnnzeOvWJpcILDEM64er85uK0+rXB4IWgGQez91Y29feuvgcac7JI7
BHwtWSTB3jta9YQKUbcfsONbnLbWVWLAZoIQYdZF+WGFuQG5HXleRWV0k0MRS/hEXwBFmHZbVjsZ
VjtE5awYshNBd0Xue8sksAjIRAWdkG/VgqJ5cu0B6W754fRjDK0BTYN2JoMvRirsphJBboHThe86
1cCI3d4MYbaFtHDFJmD/Na6gLBun4MCIjom/sQjUbJK8oOAfd49D7/VYD/0DnYDDztP9o3zno59p
L2DdBoVxeju+ZNeyw+/Bts3cBJb7lr8q4ZV5YFcs6LJiWoknox40nBbXgEdyndILIL4I9WbROmWz
y7JTLIAiPLIFDb2VTJicsFQlbyQxkTSTIIcOB0Acda855adOHd2f7JMUmcHJnc8wQBcTVfN0lvzX
0BwwJFFYmxLQysGh/9G9Bv9WBMR8yQhSRFvH477cRnfPeqrjkexK6gMpxVL3Zk/ASR/oUfhTHH3k
WjAHD/Z2YA7rw+o069kxm0Eko4ZWADI3by7C4qWEuyTpLe2sjNEFro0YNXzkx9CXwpvPYvLXZA0e
H9BT5Ni4EtkBvKCVPAwru5rFOSfql7dpZwtq4OrW2YAWg/hVL/eGJAxndYUZrrJZrPfA30x765Jo
tZpv6SkQtsaSEh7uyDT8QxbdDRQMYRhkmwBCdJjq6JdO3b1NYdSQ4ZUx9XSwo3onzjMh+ALomQ0z
yJtk7bNJuMfm0QLb3ZLwQjDBk8iV5GRKYMs/BXS+8zRVM6PtgbZr4QCvKmoGCaNj9stoOdY7Nu8l
zxM7hehS+fHChL0/ZTmBY5+TPII3xqvsKp4iRZd5Z1PJWlfV6AuR+K05PBftBS/o7/3s9chxKmdY
0Iikaj42zq5oc//L1eVr8/S54Roxp1f4Ye7uKqRW7vlgcBYGCuyP6oB1HHvcPu+m0ka1qq+HHa4/
lnXE9kLeChYWr7kwGHKIL/gndgtYe3cbWduAFpbxTYvpr+04B9pz8Ptx/m8y1MCA11VMWgiiSglJ
0DFmQlIIM8nNElauJModjd7Pr3+OkM4Mzpz5RtlEUc8tclNgyDOOgpo5JZBI604pdnwUkRcAFcZu
a+yfgAgW2waduCc3g+cN09+SYEctZvocKCe1EaxgAhW2UAXSxGV0eJax9QMbfx9posBMUo40oZcS
930a1C3kP7gDBwmJvvqJgVXCJFiVYiHWQDyioW12Ame1LUqfq5ezfppOGh2CB679UtiqUUhvDVxD
QCVwgyOBPCggHu3CnhLnf3wdPBzix1cqXzM5fV2rG7moNPf7oD1z+SLysd4ZYGx+K6Kd/C9C9y1W
V4VrXKQbdyu2P2Ord63iss77aIDPy288SQ9xOMnThKTv9h+e7A0u3pOMpU5T6xm+e1htADnPOh4f
W/3WKLZPwags54cF6BDoG0zKKClbB0iElAowe/mHZnuFidUdtZQPM+44z/WSTFitc0AhXUAwysIv
g/5mzdCrS7XuPDIp221y550Eh6LW6JUkj/b/Nv+gFAE6j4jjxI75O4yWXCgvbThBGfOnj+IjMziF
dstl86n6q3JJfeZ2USnXXdN+EIEaQR61lSU/VS5uxhHZ9T0VoZmMdq9h1Nu3AkN2Abj9/HUPbZlq
dpVCGyLABkXcvPmOqeai4M8M4OZvNP/G7iL9EKyxlv61x4rrxi/qVgNb8FYegYM8rTyTAhNiUT1j
Ucdc0pZDWBC21laQLyTRQ1DEyhQNgHBXs2TygOH+gfYglJcgBIx+HwMniI/aeWIuaC0TjK3dxKGh
So/YNe5CmmZBORNFD2Vb6ahjomLb2z/ZBJLb0dMbVRHUPQEyytt+8W7LOUcRQKar5rDJMMFTRB0/
GZGZuK/cfDfzRS4H7MwRt1mMNKFgmLKHFvy3Xpov1LOX/ULBn+621TSThEoIbaHKLR2xyBkYF5lG
36d0bM5vQ2ICs5uS7YVqmF6j69wCtVkV4tJoVllj1eZg/xILZo2IDU+rbnZcp6fauYSGipZlVfBe
5/sU5dFLgD5tZ46vTmYuaVIpWOipZ1elC3T4EAf5XPX5s0lEhAfkCoKJIqf9KSKgEn/rLGtZBR22
fgjw4G9zoH1nk9BTDdljr/ChUQqFXtMSdmQk51D2K1PgIw+bXJP4xCXkgdIRMOar77/VCpXMnALZ
av9itAe0e/g3+m2RvmrC0D3ivOflCPELdfCsZRsZ8Kk2TYs7Lvkv+bWqIBUkwqJyGvLtV5uB8lVJ
T1h160Ys+cPUEQCr6jL/ATTRpuz0CQRDVCFECV/x21HE5vkfvWZ6YlNjNsFvUjQbcHiFuRO43+aa
7610H5GA1iFmM+GD878CQ7XeZTxyQmkGIQjpi0nxP/daAv391Cv9EclJrr1PYMGyW9RkwRfieG1J
3L+ooCCyQrwNRtwUSQ+oCV2AbHYly+IAiWTuxPUWdJ6YqB/w1n2R8fGyy8CSBW8LuVBUYFlEWj3m
MiiLr/STXtHMTTT9DUzxtvZyWc3yPHhvPEpwQm4+FzEHWvgZTgAbW7pyLbDKMwKnApPTOpG0Dk0f
gUxisHMcd1odOQd0RCYkRQcpNaavXGvBPKzqmoXR9eCgtFHINid0q/m5prjMFeDiHgIB8M/bUNos
YGJ/r4VdrmGMN+5sklPNNuFsRAT3j1AEA2Hi8xLe5JAJR/gQzxB2N6XLfNMxr5UdM9gqLEuXdWrw
eOOCKAlS+rIEiD+rG08lEQK3bWm39UshZ7Jq0+mlLq/n931Bn3sWfnAB3UGNzfvCpTgKLZ4J64T1
+cittutK6PX6PjRWSIrJiwuAcwwfR/eG9l/8Y1jLWNONpqadFbkPEazuoA98lSE3MN2JMx42MaU5
ng0Cl1JpdetW/YJxgOcRsIQObNzWiGR46TjswSb+lB8bvAp0MoWyDycUw3Wg48KXmm0EqEnwYkEC
kWT9qTtA6B6fDeiC27ychZGBjzOPtlTOe+l5eMQ+f1+iJmVhT1s0zZ6T0e0d3A4/1+paZcxL281q
14Z3uI7UB/OgcoiOPcl8zhG3k8KOVSERe/EzniaJKzbaguDy7hd7SRf51x+k8Uk9DCZPIUlolWfF
LTCDzvFfMJJW7boAXiS2tU8Tmd5izBesnjEsit6/cULbZeB1Le+xi/0wNt+zEC3nxUIHUoPOXgg0
sOGwKYDM8M5hIyXgeZpI/ZxO/nPA5BN6YJne/pQCLrSqwqAw6Y9VbKy2xAf69AbS/W7ODZ9ZtT7c
QSBXu2pyOv7QNKc3QVtoe0JTM3ctmyPtoMvKijQLs2++Kz0w18NtUyNgtDEyVKVwTb85UpIZM7bN
RsaaZP57T152dga55fXEBE1xOIJ0lWEIVKtcgeZ463m59t542oubXR7pxa9gZfgA6QCF8UYD+9lW
kDXwGCQ7HeP3RKylZya1pLGU/dV6y5FDDe6eaqGjjepzXkvjIf8SQePClPAhNtvzIBh3+R68nAdH
7kFfTYYepiciFcwb9lP11MX7JU/ximW4TFyMxSd8JXT5BZ4kHNsyyIomfXqsoMAMlD/DrFSwPIpD
GzItMdjVDG1d9fwAOOdkPTpo2YcrVtwOa4ScF6SNek2cedGBpbk4DUp3u86cylzy37ZDNZnCqr2s
4XVhTDfD7el/yxLroZ3miN9P5cmXezb934rWT0E/vPl9U8EcTAiVNU62bK53mIIe0RrhLncuY2la
60atSHY7akQFgAzJ8c3SOLfySclxXll2a+dTFdV8eCtaC2QEoHWt0knCAB3iZMuVN/iA0Mmlrj7i
XAHUEEooNEzLA3jmr3j9F76ztRKPnym0lHNlv6b6JLeTmWqO5p2b9k95S2k4ghkjan35nNTzncZd
sz18m0IY1x/hMaIHV7nVk3i9CqP+2nZZ+L8WiBeCkIOTyyF/3qixMgepgYFrdZoQJy4u6B+TKSDj
+VmG2GkCrAMD4Ag/zvOPK8x+TIcf6kvw/XiULr8NL9Y5bGKy9YCE3JTiZHoTHuI6F33X5BDl4EbF
7Z8aCyp6zx53t6qIzO8UUdbT1CIaZrHE8/VoVIvvWs2K3Q5DgtnQePHOGexupq3fULoNGhvL4NAj
SwgoZR7m6UgMzDzwJkIkPshvrekfbanr1KsHewW64EFBr09Kty+4SThqt+aMl0083r6DtEB6PRLK
RK6vGcZ7fajrf4V3uNpxOfC9VzubZHFkDr0ZkQkJXDoi+g6a902fDHc9YBUC+CN+8fW9zPLQF38u
MRvkJ+4smdTge/7xecsMSkm67aohSdKJFIVFPrgS55GgmB9JjZH+FG7xNoMACUXhWP75NQAp5UTW
x4HdNo330nVVcFR093s0QxZJnfkh+9dXXM+W68olofZBROt3E4I5gnt6oRbs8//c9S7Pf7xHtc0L
8g6Iz/xS5ttN9EhWMU7pmye3ZxqEd76Zo6JGmLNkAkkdWApqrgfmVKFRbgAHkMlL65WX8B/yeG7C
6xche7ZEYP6a+HfegG3Rtk72atXh9RKjTjmSJ9QVFwe9sDye7tyP49JJOXt/L96drVD5rrXN1GE5
RetPPlkv7wxYJA8ECe5bOM6l2nRQI+MXKSdkCJlUEVluzUwKgMgOsTxJBUKASG1C6lVLJIP9nhHJ
fuda6cDh0VCA2PZ61bdzWQOfOzD9RidSkp/kno0DP528iQ135VRIZJ342KJ870yk7cR2Uqm1NAsx
Lo/pNK0ltCCsPklGR0DlSQuFRVruVp9oyl9jd8ZOokixsXmKRtLn1lNNj1D9NTe9xgCQLhag0vMI
Pk/L9ZtTYPkVD7T0j4ReF85Jb5m/QQhl5ffjW/mJBv8Ciz8ZhLztI2xl6WQ2Oa9XqH41U5B+VuSS
4WeKxdu54ToQORpTyxXSVKVMyqX04glwfIQELSl50DgFcdBMzBokLAfpAMve5LOlHoqGwKBIdmkW
h/y4giSaxcvn0xsSqW7QKqYQzxtukTTuOtZaEOQ8QbV5L3WvDf5cJDJRI81Arb4kS2CuaREANIE/
+dbvIlP7Ol2WZfJj3biowH8OpdqeJbAgW7SPKPV7gypQVIdGCGxEb2kibvH8rlw4avox+L5rDwPY
R6jhpm4DPvUvnwtktW2YntiAIAP5LAEYC8V8gP+Lyn0InktIN8OuyYL/IHkrfQgk6Q2+u8qLewoM
pIVTC9EN5b8k1pLSvG+nT6TbGUagQB1DFLPXOheFLBGQcDsDCCW1aqYVcXw4d6/kWyDp/BHHB/ee
pArDWY0kfcjgp68ww8iNZFEJ2xiUDHQ24SQqu7S6KkiLrqWohMX6f5ALYcHYFwGxBEZ/6cac8Mlp
xPYoJLITR6+MkUQaLkM4PrH3LswQNa7M7WgXsyJWsyfcY7FP65VUhZ27HSx598EzDC+vkNnTp4MK
I6Ohfm3HrdLGHmSXQZKM/Rhi9C4AiyigcI1rRfEHE3r2uMKk0Jc4M4cSakhfZ96sxN8qUrkwqrUb
HMMdtm0QWO5VFY9oYUFsNMB7YoNVV4HpRBNtWiy5M+EJVNpn9ejlt/9jp9GGmmJjqbsa+BCILW4Z
bqunfQ+9Kl9Qog5E4y1JM1aZh6t1MhEOvNX0q38nKBw7uXg4uX8pYqXDlRDsdYLxi2hfAAqSzNnH
9wTlXTWiQQOVIJIao4Ld1d97BI2OmnkpK5vn3zKjwUU/5Ddfm+PLMW4fS29ZM24N8eeMvHAfZxM9
3MM8N8dNxBW+Pz/6z1VsQryVSevBReM56L0PFtBWFpuj2LTqNjmaSuYN6y8/Ctm2r1z5vcjFG3q2
ySISUbSYVyBoWbjlviw9rylSU7LMTlZmKlhfoeN1C7qVYd8XFYb3mjiEdzKJuLAhnXUONczHz6Ik
MsxiLSoIRLvBhb7E47xRNVae13cpPf2q1bYE2XhO2t/nLggGxINBvI4pcN5ueN5wY4SuPAWTQEUF
Oo7H5U/skopqFe9jaiwgarTo5ISVk3hLOL9/t1PWFIyBcn9K0SxRfllIn8EedgF+hwt2rtjFuxO+
GopsmOZH3MpkTbse9qVi4As/mYjbE8G62j/SA19mOrhlVXRAMBUSDOnkyk6JiBkh+wGI8l9ak53v
ohnOFeIY9TrDbzrE1SJWE9j0XleEXubRlFoUPzzqs2yFVq+RgFcpMXJval9EgTNuQoWC7szwlGES
VnnfyW/OQP/w/qHKNZEaNVXhgtGfrIGk7ahxhaKOqJzwgQ0X6+pkNSZu0NSybvdRXO+jxDbhgysT
dtkG8Iz+Ws1ZwuxHaGLfKyN5VjGjVr+LnKsyEIlZ/WXF97ZoWY4Pbq6l3GTXWiXkrpbqdea9ZIO6
NuHYP4cbhlW8bxwzN7rUhBcbC+FB0sQjiZHh/ANXPkxbXoYcAbB1gT0uz5bMyO/wkO+BfKwX528Q
iEIh+fd4prwi5gWfiBQ2DrLRygUbijFbkLQr3WrrJUxVQvbpdIEro25zmOZOmWbDwwtycx0DFPaT
15smLbKY0HPGe7mYmmiphi+rVLSC/Etjy9t8M7AYDz5GK8MgWqELZa2b7v+eqY14Y+CiczDRpBx0
gRKlDS4i7gYPSjhg8VwHRfzPzT0GYrDl1OJ5sBoq+EdqbggMlGBoVLPTgjHHCCxYAZrYlNcSYT4q
Jar/IAOkzay6gcEmW1pUzNy9LfEHVt+6P3+SW80s6lXed6adpF8uhBew07+McSxTV8ushyJjUrqI
KLunlrssYZxLGkbLPg9nQEH6xHeHs+ZVftgYz152vDXhSukGgEJMwwcIIlMr5lo+e+elPeLBFTkv
Q3jiLe/+Eh0Kom7b6OFXeh3OwlrrNTWe8WN1Trn/EvTfKRBCleYl2jo8KDn3PCB+8ABhItujU1Dk
0nuxzronx6adMtflFI4xK6Zh1gWBQyJRbBA7s3Je+kXDL+SeVtC+aUBvwPhH1agjipzV0HXK1I/P
t0mh8a/xQ7K6qgIbJaijfu5cFAC1x8sqN3VZMAzp36HAWvboMzWfhgZ3P++Rp874ceLVHTPKcZ3L
bOfWt+c0nHH/K/9ufuptkB6bCYVOhKQW+f4waI8jHeZBfYmJoQtvWzyNrrZDzurFyKDgIgriI6DR
uNlJezR+dpAVOgcdeKoWca0ro5X+wqi8Q7/qXc5TjpD0AJ+EUkIlIj/9JtQ6sYH5y1qyuUbaXB7k
1sIMA/fVRqjwq0ZGQmNJFYPN6l5HGCZREhNi6KGq7PsLV+AZbczid5x1kUMayqWMYgSe7QTen7KR
EZb4i4CrOnx92XIYUsdCG9Fvfh1vSvHFCvewU22k1/sii0iZ46/LtDR0GJYLWjaRMvTSZxQFIThd
9ZzWlGb8lHP6hE+RovnpYBLi4oRSQYSx356tE+p7gC0rugb9FmGmKjtEowjuPFp804tW7CZW4b1b
H9xt0x7TOkGiHYiD4CuGJp3D6XicajImkm3R17AkskMzHUQqORxuVUXIZ/qHDzNGJgVxNyQV5UAe
u+QaYTWVVG40478mTGELxFKt4l9opDZFCxBrjm5xQtjmQJxnNWRlSIDy/CJXVtou2bb82dmrWU8K
MGrlM0ezsRmRXqEeUy+ZGXA8M/vRN4RFUPdJ+gWaAr6TyINjPaOsNfoRDf8M4A82xPh5EASCh/80
/jjNawhzvDZtIbu0OUVxyJnfKmLJE/6XXFcqFTEadqmUzx0FkERUo/oDx3DqWpOhbFEgDRSvGHyX
L7bJVsjSTPhGk0BryRPyZ9UgPtmoUjYYFYvWZEt8ffitc+zxS+rswaRUI/H2KhAIz+Fgi2XcRB2q
JQxEj9ROh3xuAuTDjuPUVxtw+hiVqlgFo/TqaIheHC1AQo5TtDJ7NwpV8F8J0lIq9ReC7ibJWW00
UrEMmMR9KGcb+mVHigqae1O+OWuyTc5XI/YXYfZJjxGJAMoQ+csZlcchsjg8/nSJknw3xN6vqakV
m2msTgx6yTEHp9GIO0I73OsEaejIjdECpnrEqY23kJ5xvKczIt9sFLBWX2/pw3JwOoWTrQBuJBGJ
uutrXTMHuIRLDHZwVqlLJg7hRfsbIcmxYkV6rdfhMXxZ4iWHP046G71pXsqCL0wbCoMvphttFSzG
VM2+V+oD6knDtqjLSa+txzacCGhCZsjDL8Jtet8xL4+3HjVdfOP7GI/cR1Jh87fgL+vI3iKRQuHQ
RPN5s4pkqH80TcI9/tswe/hXhJW5gsHp+khslB1SXfhiKgWC4BASi6vg3Szz6wKNlhrAGCDX4WKZ
uyq7rp/cvJJgW4qSkmHbpZailO6OPVSV+3vCDle3gntFNcohA+sb1Neaa+8QWcJBhnfbaJ0cPttL
UGhDUnpengQ9oYs4JtqhRodkcGYqkjLtuMGzz+sWs2sX6F6yT4jiz7X7ARy0HqiCYAZASIbAW+Pd
1QGaeVQ86VhKZjMHE6geTiHs3Qok2To8sAOAohxB80mKXsC7l7zjbPn6U/DjSbQMubufhEsgm64p
GpOMdHUAPnLj4Bh5kaDQ3TK8++kmkqFFpNXJ/x3of2FKpKh8m104ueBdq3nZY5JnZkMb8eAQqnhh
td5JWM+HBPyEq2MxsbYdDwH79ZZkU/6Vnqzzpt/vCx8EApwN+viNr+FtcYxar6ONTroPe8/+M79n
FKviOjVdHmEgDmdPwBRMl4YoR0szpEoB7OWr1nXYvSdgighOvEyeLU10BG611oUpzGMcu7VOPEzX
gVVulUMpHhhOLPfzlkh+ycVp/QnB5OBI6oIQMemm7hllvN+S6owfyG9fKfYCPw7znUuI1MuE16kX
gLXZAEBWEqAn6h5SQR+nbEbQcyDIkXuH5oZXUzdBEreZ3f48VcEVOx2mjsEXi1JXBrPJHBYCb7EW
JjKdqjk/BeHt7kmWEZ0Z5h64yqgXuzj4OcoDJCqdz/jeftBMXZaH1HDNNlX5VOFuNJjv+8ROgacB
bblFbRqwG3M9hgFxiCZ37CdF4Pjpl6EJGpzqtX11qHv7mdJFth8Zr8JhSIuQU79Z7fUykqQqtyiU
5INy7bDfgL2bGZBFFXMudiRlhaxEV4HNh1v3Kn1VxajjPNFHmPFQeitYdUOK9XnpSL+lhhDh6cZP
Tqo7+Vm934bMJ0QUlQmHkKV9X82TkC4FeFvCL8P2X7xbIgk7UD32yTe3vSPjoC1X8UtFeP3hnfw3
Kj5NBH+6aFBgNuLlsSbYN1euxfC4qWTrWGvMAAMQleeZlNBrJzGfOgmn5iI0t9VlFvA9vPcIEnZp
0vNH/PENxSnlOXll2MjyRWCaahXreROp7EgrcgQZKe2xt8WX2ixfzVJAYBwrN7pg843q5H4+0OgA
1+DkTDWtiSH4F9MbYon9HgrCHLWFMN4ACbvQp8aasyp0qnxmv/1E6I17j6PJBVekLzsxV3ZTSXz8
XsBr7F0l2ljflaCijnQZv3BnTOlWrz3UquFZxZ7hfYwfTBlIZGtL60jiDST/e6YnmjjhODV1MLtd
gcWzB9kIGFJ95qrH0DfazuciTaXFg4jAYQzczD8YTyKfahdBk0GpE4JFxaR3dNtkAcDQ8uCY0jKY
dNUJxWb1DqZDHxjMF8dN+lY8145aHBZpx/KiYBe03vPtTzXZruqxFHr79KQyRhvXyHtlt6kFzTZh
3SNz2FUACwRn0eVpUkPdlB2t/97jLpUmBvsILVn+mCzo6uSHZt/HFfunJanZqpahO1EHjW6L3hJ5
NTCkCfLCxGo5h2AmnXzoqEmpfSCcW03Isxn1USxPGobMt/vT3RaCm2ZvzKH+ao4c7P6Cwc7rQrfQ
INSEkjZeyjOh2W18LTUwyiXihYtjBysQjuXlIHZPAXlUdQEvwzwYsk6XiH0iDFCQdFb5NOGS1a/N
iimeUcKujRnOggYGT+T4CDlJlBWauel4Yof2QJ2p45+0sL4C1Ifxw5FQ+hFW2Qhu+qW2b9GQ5q5o
leFmzw3EvXkTONtwEllqufr9/KeQ8bVdhqtb172iy9ZAW0AjeBTRzTlmrBV8ng6ZfZmV9AGn2bhM
CPy/8ArB0ajaFRGuuBDTdPiF3H7FtNsE+fAZ+hhQIL8K3kRi6e7TH20Zu7xih+owDgUI8vcLHy4i
JYmBampsKb+XgbZJNFWO30c28xNKPuwnRs5tKMmk/Wl+inB1bYdVhd/mAaB/u/mU/JZuqF060sFw
sUUzFkxLHLvDRNw/4YEWNt7urWQei6Feexs2gJwI3jZ38DTl9GwU5kSzaRT8wHht/6oYf4dwgQlD
+enA8/0W3oEBxB5fmB8dR43rcbZq+JWy8hLkr+Xp0+9viIPx95bwTsuGMZ71n39j7LZsfS9DX25q
T6dw4pC6nwFbI/okPTi16QZ2YYzwGD9WcSptVsB2e5xibUo0AEKNxfsHhL8jXqDw5ReoF0NClAQ8
gJZthXO1vn9L872p53HkYScfJI83lWtYeLczktnQ0PbmmXVhbvoXvCyGW2fbFwCOt9MviYYOFbCS
5rYeI/cZjs6NikiKSwceksHQOWt+IBfbjGtS7QmPqRNFs6ppJwbghOrKPepOMmP719X/5YCoVIeI
e5yvSiXVRNBC7CJxm7V8+lEX5rYEZXc8y1bnwdcwMk+wnaV1RLdYb1gN4NfH7Lo5QE0xILc6U5Ba
h5wAPG1v15adyU0iWnjVX+z7MEH5QGj4pTpDunPbnv5uTY6gwiSNcsjmspCz9mQJShauJ1lKAN5f
hbIaKUqp49kYsK34zEfbsiEsAG+9iQQs4/d9Fb5o9lvONJPOXGGn01zJPChgst+LyOzjHGr21Lm3
Fh4JATeqTF6DWTQhSlEAsW1xsj8z4e2rX6HwDVH4Cvq1L5X7p5fCuCHoQB8s0Q4BDIHfYqVv7fKY
3c27FwmP3Nw36k9TZGLAqxLnGDuxdm+0VZhI6FCXWnocZfdn/sYe7Ff+4mxA4rXqlcxDxnuulszs
zBJuaV5lgUneJQdqBBaH1nRWIg1Xr6/iVS/N+MbtYbnKqnPCghPezMeY5Ha625gZtHmMLCC9Mea2
xabO8Zse68W7+73Nbx6fY01Z2oCM5fWl2YBWyVrpyPNQMDenik0fFGjYNodwU3Fk3VdkuIMTH4eU
tiNCAlAYmP13k/gnaZtbshLndmygrcHu8bDevqNuytDQxV/JqBB9xkgHXqBGodXn5hNJhbqLrcfh
TMlkVPvJjzLkxlEy1EaxljFUECjiEj5yJ8Jv/a6nZ0VucTp/0jxQMWWMuC4BrfrTWebGRymUnrcd
2vm6rOQyO8bgMCqu82hzEo/B66/P9Bc9Ism6Vh8w0WLmxNExp6i1GaQVhAsfpABhsO088+GTVmFr
1+60vVBbzssRDKJOktUhQ3QEmczzzUAFn4gjKbDcDEdHBV09l/7/aBLMEQDpNCATV5X+HahO8/bw
R0wrP6mjMXG+BiMT8PyAggrNF6gMFnxMLiUvD8yP82OVixq229mByJuTe6+6MYhEk305P55VM+5K
+UoGOj8lz3qAgLCr0IO4WKmwpQB8yUmOAGD4VCivdZ55YqgNa+8nrHCPQBA0JqgKFmLuawN0Hnek
+kn9sImKJ3l5FtpZZ/nhGMhpyv6dAuIorrSMR64xNAi3Hv8Y6vFGU6gfwWkoepdcDoR0ZrBK0kdr
iXrDztSF4mrDYx54l6UwUZp4sK3PGA3k8o6aw2cT1SaDXZMaz5cox3aOgSGYLHvZHezImxkVYGt6
7f229r+WhwpKcputnCr9erzbucs2+GO2Q5ePL0rxTV9n+ZuHJX+CXIOVsPjSonp2+ll9Mv8tJwGE
kKArrwzz4pNncHqLDCQjk6Mg1o8BJzyAh8OVuApXd0iCKsFpxceT/iZD8VX0/uEMTwvql9mYXa/K
s5HsS8pVsTApaVKW3EH5R0L6FkQsjbWtJAouzt8JdLna+F8t9zRTGSeojvdxMm2xLeFGxXC1Rel2
l2N6WUKUXpCh7TM5Rpa6BlDjwQTQPwwlYTr8UlTEF5FXj+gbQn9kQtMtjvxUmU+OMUoKGsh+hinX
wGSMTsSSIVqeJN5J87jqb5tS4gDaGjaRyXCa5Io08wFJWi+Trm8No5XVEBYhBOcTXAOjDSwLDjSP
t7NLBoBI8O9XgaEkDtjNSqMRymikws9qrgdcl1q5UAFJ6qM729GglmmG290Y2eBdwBC4atCTb80l
/OWZIDX92SurvaA60RCaLD+tROW1oFIimG7l1GgU4cpbjHrr3PkGSxOI9TjAP6xy/hINZnTjOt/Q
fA6QiZyC/NDdW/I5wRsaK2Ygi48KOp+RW820nA7XMjRHbeoAbBCKrt97vo30WIZ1e+9e7GMI5joP
ZHbiWvFTPJLP8YJbwLpFEZKbQJRKieey/0VqhbNDMeKcjKgmBORHC6B4EZQEvhqZdB15jDEqrmwT
jjZbxhLjQ8EaPcbx52HAk09ZIsPVn8dSNWprV7ON24OBRVeoVioOFcXoasQOmMvrh7xcsoYgZVmw
3P8eley1uGtmSoPeyi/VZ6cFsXOchx25O4IywLXxkNqSs8w/zFAudMopwco5Yd9WaRxmrZ+eQ8ll
nzJHL4VM8M4CNCwhC8Jp3IAU4eRmBz7ZQC6Q5OXzOAfo4d6MEPEOYWp9ocnABjndH9mdRAOPoG+p
FG4wmoe5nLrQHksJakboXBspKLMbxH54ViVPHFVOZ/2FSLlnWIIF6D6nRinEYqx55O9WIq3L7hPr
DXEJWzL/8yhuAbsGAdJn0Oeln3/LDSB+jmMCRKHq+yccz81uvtfM/+oE86WtAF9ea4Mh4Xq/mPth
0h2gfEPRHFErZai5TU0gn+xcRKWOUZ5PTd+y4sW5qi8+4FuZj8Zr1+qqWht07Z7dLhMTaLGqBEus
3vJmMqTlIRGoBq52Rc3cXFc7bG2rW+o3VSCnBXzs2d8q5WEDWyowS/EReBT8EQnW1UVtwSRhux39
rzMdeYECM+A/oRENGtOQ32qf8skM1Jk8PBRnV+n1kbxKPfr+uE+i++lscm0aVvyhU4a7sdrjdIvH
DGKfCjKs7UctsSa9nT/htbmEVfTKoqZ8QIg1YaG+Fx27nGyYE2slummfcPbr9rtNPVp/LLISKl9x
WpVPLJBDnPmwYFcYUuPGsa5h3wUVdnIKySJHs4EAZZQ/QT5vVUueQmQdg9MWvUAIARM95XOqpaf9
SHkE7wq6tjRjzx4xy7AMQ5YUUX/9OUL9LqJwdEQCQnDcNurZamgD+YtlaC6oUAFuPEUpPGgoqre9
Z+Xgx49AWS7PWY9awvZtQ/R1I6ndKBGlqP8NKE3al0O+iGTv6zwhM8rt5aYNvzz1KOJ2PWNgcZx2
8ExovwfGotf8K0YkK1lBMoY4Vv06jceOUgUpsinzHjK2Cw/veQt5lE+0Cv+sq9392y7RejW/yNYr
ry/hyWgeZFMBUOd/CRoBlIFeWdNh9EPO2b9ciKVuMNvsqNl1ocQ2ecs8TD0FBDcbcsDDXlprH4K1
iK+ytBGNOZdsYINuVrgfkTSIuBlsYvQj6hQW4yUv/SEppDJ5L9KleFmPGLcT0+M9YfI6KYadGCsD
sKnE+2eAob82GP8yhREOY/iDDwN5voVOwPaey9SFnKCK+IkHImi2MSU/pisry6KuMKGjo6+gMi/M
XrrMdQN3Spr8SaOtlKK2xG6bz8pWIdEw3+c0Yrtv4P/aAlPWmFtyCVJjFWQUDNAV9py2fMSLfMQI
fvT7Z+FS5B/ZX9OyJ1ZiwRJrWDKngs7B0+MGPLGxhEdZEXTmwTrFff5ezoMVUw07CAskzzvKpdcb
BR0jaZOcy2JeIixcp3vSupGJ8usnEXPt7Zmzkv32nb7pVX5UlrU29142KqitHn3ECHo2BCwNLMHD
pOqCxcw26ZMDD/vYkZwPH6GgAIOW9KMaySys6p0Zvb2nwm80mySxgyXDh/bpnFhh0dMh8NaA2+u3
B15K9smrqqbXPg8A7eQ9C7+KCmKOCOGfJpJec39o532jd7+DGaT0URKHxyppeTWMILTaOBgmyl50
Cy0KxPrsAax834Upduiq4JgxeDEcukqOb/686gXSBPWW8UrmbtD9XHmjkqEP2MU7gJnD2n5GCOa6
XIuPwu6JvkdY3JSDASboILMuwhMLNNgnTCrXtdasaW7lhYT9iYlxcK4SuUIR1pN12FlLGthJDixV
6YTGDeOxuetZO46UTqClEaQKUiXFNwDPsdUZ5Yoop8g/m3udr4ZZV9pCGmVzyyUrfP2UGR2X4fcq
Ek7fEV8JkB25enIllx/DmdXd0lETM2C+J4fWBqS4FGdf0Hu6qZdCeteKwPPa/XkSKv+jAbGRXoeP
fCxTH3h114Bemcp3O+fPirhdb1y6NIHEQZzTxI40dMVd5X6ZHvLYEemVygitiBWNEY817zbFHIwc
EDyyrsSsm6DVPTqksDQwbBtCHdzpiNwtvMgIfcWyrpqygaI0hHhELPdsCAnryfBIYzuqyrzzBTbd
j6dP01vjbZ1n9BhsHJuVil1+laCxjYEL0ACasww3AAnF0W+1v4xWUp6MSxzxINZZ1M/8DAZzX9n7
yVkAI5g3h5MDvzPGkrEywNaqpe/BabBlgSqlQoiFUjDZOzZLazcb7LH5IElBWvor2UJkEE++V85L
TGQR4QwVp6cEW/tm/rCTSXiRrcKzx3svKslB1eEzH+1zZtASUuymfFYhy8tjbd+rTWMAhuL2U10K
WCdXU4jLB/YLu3SetFdSx41dtDgpLkRv4fEtTwN4fSPpnosAOc0JuLbT6hlcwMxw+V8/kIh6KXny
Bjc8VZUi85q1097k8onpMpw8bJTMb5Ek+BvPkbs/dUbqkpUZyZoKXsyIb/1D58GecpYmamIcwxKz
JlCkdcE74TAEyf/XSylz7HcWVJJcAreX7pWNtbgNFkJKXOuhUKhcuVlytWtTZUzQW6ohjiPPFmWr
zVGOz8AYEjtzEPpsI6oPlsNgVpF4e0raaoBuSFAlBWG3mfO2mfw9b14BTxzfNP00EwFwqGP+HvqE
JAy90f0BP/5psX46AxKXr6r+jcqPLB1aLstE6EbZuAk0OJy0EDLkUo/1DvxkJfPMGWq4jJOY3Ymy
xmxCQ3MopU6OybKkfeoxKAch0ESRJVPLnTP71T+3faGsbvzz1AKBvfbyiAS1AWJQJYXbmvrRP2ta
6UHBO94Ivsc6W8awoxP2bg/LEbC7ae4MDgkbskNCNWNLzQKExYgQ/SkJbgkOQgAbPu341NAjgJEV
zP0KWnwuPzxmEbKtTh/UuumZP/KpoCFx20kGgdJoe/E9+ueTfzS3Pc90LqEs9JVT/QFOE4z5ZpJ6
SKr3gUlh9AC0cYYd3zJcFZnvmO/QhElTcd3ln2xqK/dKBd8evGyY5gTFb4zUhC2eiPiZmb5zvWi0
2P49c2jCGy14IXNeJoNpE0Eo+VsE10lHOs0brz3U48MZX8DQdVxBpLPGG1Ov52pRKqI9juo+5Xze
82GjfU9TnAyyWNr9N3ny1SmDBZvXX+xSSt3YzRnIWfPlx1AW7TYLq7LZdnOGY7AuWzot1Rtv+0qu
d/89h6MW1NbXE5Z0Kx+cdE6GLrwq0n7lu/+ZfHgY1fYrtN4w6qAp6bs81HVi22Kbarrz+GgCQMRP
L+q2paeBEMbxgtUHoo6Nh6E+2yByKIgqA1EyePZRJxh5r8Ce3Wak7B0KqmJGC+/o9UdlW0hT/h+t
HfEVpr/KgZmG2GyTc1RIZbi0n0FZI64oiFwufNsIlsiV121yvatWo9JNMpRstzeuYcBqC46GCDmw
CQxnS1XyosfQeJDr/SL4UqY+6nX4qQ5PLRvm/pzUpRSwYqnol3GExVtR2I28wSsxL4Zm+6rUU0ei
leh0KrK8kAgZRbqwGVGmtilctNxgfeXcY5eU1QxiFYfUxDUoU+lc4lrJwQG3CKm/jT4I4gMMHIMS
DE4c+NERu+D6899z6i7bBc0UV935ueH3Ft1Jk8tkt0zeWXYFuoQG3zu4LBEh+CTZxnxKAzwAUgRZ
2bjVjn9BA9jWz1b0y98z52Ubgj90mGJAx2ISa91NrIOG0UPKQI6Ev5c7KQieMI+oQwCMl7P450p5
+VJe7OI4lcxiQWqTSSjO2eiE4i7scCNtkX2iorkSdOGa0k9UE43WjdpUiMT50QcoF3enb2DhPX52
eWQtVOwAi5IBEkLEmu7+94oMaO6Q0CnyiCOgb0ZaWTAx0NsyjIOIuDe5uuLwUQJ8454uWSL7X1bS
U122DViL3K/4L2Je+JggJCWEaUKEZRJvsEAFYY1KX6IxDgGOOLTYaqe82FFrUwc7HN5h/ExQ/4f5
hD0XBtVZbqoLjh17EU3Vs5KcJ8JqPFYWlWPKcOBJaac0pidoYEGnryimCRiE69KQjTZ2ztjIXv/+
14+7X+cpvlU6De+UUxfg+x5VeIMH0wgu5ek8XgJXPnOG/tqAu2CdoVgg5YYSKx7IRRc6PSfXQ62e
CIepAb+aS+AZLkXO2iVuzdoa9hyURU00vTRClO5jHZySegMAshTWjjg9iGhv6i23vnpbsuxDx0Ty
7l6GscJeAeKkpxzQAZJI7uPyNuLa1QGI3lfJs9TdHNr2B9eZsh/bFH+dG7BjewyL/jp8epMq5e1e
Y4i58HFdbJ9BQ3pIAU7J7gGCwbR/vTp1tff4LCrn5mgDxQ+Kfwq9RWLY5I9SaNhJHCcq0aHni7VB
n3KcaFHXaO9fKf0xUs3BKcFx/41tAO1oCuQ94FY2HTEOI+ygxBXpn1Eidmq2U0vYuHnvptPblxsz
rs0GvJO1kQ2EhdUwj9wJA3JbBiXZwiTL4BmOWw2ajE8b7dzo549XqQeJzVL2Z2MKH2es509lW9uz
stdU3Em9UNd+jSZz19HeM/46T0/Kt2EhxL1S/YihpAWxgXQ0pIqmhRf7vrESTH3uevKXPPTgS+PO
uc8qi5Mx8HVHskG1BW2ukAMXiLl2bzLAuWXGoxFw1e4KWfWzgBzUMxgRP+cIOvznPTvkUjtYBsdI
pQsPLC83PCW7EEgyrzt9aqLnkzzAha0402tfvwhg3/bugJLdhoYhZ7f3pbZkfh3Be9ssoT+hDXCA
ZGBGEaqcRnCAXwAPFaoYIK2Qqc6+CcyYY8W3vNowLcE5mqABgSCnL2Nko4TQ/+SUm0722CGOIyHa
GaM3Lafx+3JaXREkY1zR9VDqaHdoPBJgub/CTxKMrxyBhM1reSQQfO5cc+P9jp5TETF8maWCiKvq
ixDfR0AcKbUX64qukDTcdhoNdM1X+R8o1NpxxfQpXH67YJZiMCD5vgsODM6E3IkAgvO/DruGM5Aj
1rC9BE26LlCowowlCrhDA5x1slmCljjfR2jWZydY+dGm7yJem3IlswzqtJgWdePkRg5J+yI6LqBG
ue/V09C+5tlWJF3Mf22CtcdlRmnWYdKkS0CLxXWKho2aRLIKgGCl5Ylon+U3PrBtktBi/Wq7DeiJ
MxNnIGfJktXpggzDPleu3jLgmRkPHkQyzE0xB/7b8KuR7eXLshRfIyYk2hhNlw8TqrjU3kpphiPb
c2zPGYHBuMkRS4Qa2hUOi+eWIGb9PBPtC0ZcPof3ek+krG6R8W+WvVfy/2spS3GshHNHat6/B99U
jn2+i4Ez0fyrDzeivTMC8ZFgRclT8XLW5+j9w+KJGOF2if4H5hovhnvPB0jVm9T7LgXRJcMkoqLt
TYeGsD4uB1GpX8wdb3kOjls7k89guFhQh+RyNV4K4rJnn49HAqtYAoXGveFMPrF4dlyGkV6iUsuV
uGv8EzOnj9DRe8yKa5HYgRrsLnGUme8Z9HSBREQafvJJgCKqmE4STDDkgS1879Lvhvg8Ji82z+CY
EYU4ZkRQqfJug/e3VmZ1RLLmxfbZfg5ueiotObfpcFmDBIjtVtZeDuEnoMxGXpW6H51GBaM7cZkr
EtbuJXZRppzMIPyJf/Cf2eRwGgDOK1RnMY+sWpZb24U8XbcxTqflkWoYODSO4uwCZz6YjMsrYLNe
AR1rKdqJEXKNf9L2467uRJEKC3MYxX3ApKJ7RkKmKgx5+SiXO1wxP5jFoBRuc4rOjQ4pnm5h2ETR
7tCwKm2hpeU5tOfehYlslXnAwGst/Tyww9EZBfkBIY79WlLEVf6rUmh8CWfTBz5HV+E1TF2KAOH9
oxHe5N0/trbW5VD1R9mDu3VnKyXC8GMMRZFs8xU7+GhYeyhRErckc1LSu269N+GpyIqrHMGxBvaH
7zBUCV0voBDX00L9+ZHd8PtbvXFpqIyOiC6OlRuYX5DgU8QlR8pnd1kPe8MjEMgMtZS68vybXDn2
k32UtMUoz4LNiF17DdAq3K5jsSEskmCswjTzW6Kw6hm+Z5oAH54QZfLfmzGFYZrVqcy3/I+4YnKD
OnW97GfMq4TzpLxzRf5KAX8ivh6a72JtnaWlkhz8A53IS5BfpHISIsNwBr7spDVGXGgnqFea3zBQ
pW1oliuzjGSGaoDE7VDQhutgvBCIMtdnYWOWrrkymlmgLG/xP9An1mGMR/qhuK+GJZ2BKPeYQ5Wu
jcu3xrIlVyzzl1vaQc8Nu81NAHJty5Ffj9w77uZTqvzpYoSHsSV8mepo1ol5fmhT4iCY3mYy+NQu
PEfi/HHQnsAjHAit23c/C5HdY/y+wY/jm3KGbBdP5WcNHck7oDCvn0POLeVhSoN9NY2b4KDF/v9g
ryq/R+6sWb6eLcg5W9KlcidT2Zp6/RMyWz2tdsL3aPpPn79P74413BeGe0YYg5we1rpu7oOrAJWf
i0fCMH4KG3nlZpdQuOU91ybuRzJa5Wr1As+DDCVmvM5EE+lfgUiwUuwU9nBnosYR8EhGnUzD60zp
htC2ebvL2CiofbSG6E3b4Ab9ZPfKbU0GmQpOWb1eVxPKSAD/uToLtHXyQZ5R5DHmdoAWVJ1M/gaq
HQm2S9RqjNZ0foTwrskH6GjYGBLnP6jmhDXF4tllOjcbsk2VWJZW3lp4QuzniEcSuQEM/uLyD7cj
ZVYxqgqpQgxNdBayqpdHAGj2/jscmt2G8SX4Gtoq8e+FG1eHTjusvZhGdRIB3PxIVDGC1ehI48lT
QNDIsu2/0JBoiEUA+dItW2iCDR2vtrv0EL7eyra6UvKN17evBDw0yOzaoMHHnPeM3JbUGPYDaSWG
gJ4W9321JeHqmsW7Q/kDuTBlqBsas4bLsR90YupJ2aqZgvVKfpL3n3ILR104CNJLRLFhqL+VhLKr
qtYHyHi3QTa5ZNtwbc0pAzq4yxas3kunYIx8BHaPUTBvZIgetiZticuwwI1PNesdPsrWgRIRnT5R
Doox73TbmIKiIZFTeY7q8H7LPL4uaL5UeNYp2PhVl+SSJrc45ypdHypOzXczgC+HGLUt1VHvce/Q
DKidI89iUmI/cvTuU8t6A+O5zToQtJa5avZrUWXvlFO+oFuFQHMXesBqhYhcHI/O2QpLjADgzA5s
G7XcneMz2romIcM2Q6VudAsvHtUQyf7KPRdr1fp+zUwe2rlRHG5zd2zikep7g/kgZeJuTOq2SSlT
Rr5ZO34Abw2Hurk/ZaGoWlhBKvneaVsf79DTLUoiIXPk2UMH8UJhvOEgjIP487NzaQ5n3MI601BK
cCPeMDnJD25u+AfZpHhMOX6TlcGbo/9rLN6tZPuPn1Op2Wknk+AUUBkcswzwENV+vZxNZe/z+p64
u3IRxCa6AQPr3SP+A8W3aMSz2O/NUP3NwmQZ3/kG1d9Je393O4KGQ8yBJgwynICQWMKBjWVNbE7n
BCmi1gwdiQNGTRMfIuSTzJPND7D2DQ1gXf+T1dex0q2OSa1EXe/gHh0CpM0F+47bAEjs2mp2dEL8
nNUQqObgo8a24ZocR2gKiM8/Gid/M9ewaJ0CnzxBuLh15gQqOQnGRW7Rsl1SYFJ1lTLNkWGxjnCc
Q0JxzBLOQlXS+UWIv1FdsJzmYmXj/DL98/R631RVaUBRnYu5lrtExrhMKd1FnRZKa7kILPqzJjPc
DlGfQSyNUuGq8Xtuk+/Ud5FJHitRbN+TA/++sReIOAsLBIlXeH0fD2dXYwddZyaMpmhhjtnLswja
slOU1aqIAztk0Cjlm/V8mtZ9UCKRe+GJLjobiHub2mkNL8S6U/k1ZXWGcAHSvRnHdXtB4J3vv6pa
GYZFiygCLrPfgCKDubTtKhEjoVeArEbZSHa6ZTCuDcZvJdYZ2WnWmY1qugTKZsLPXZoXO0T6xgxK
SC3gaC81CDKdDBOJmgBk7FhOBRRPYfZmm1U98GzFh8tJijTmXiGcb8N2wqWUGcaSJJrk5CxfzLez
YjSd5qCOIMoEYNK/Yep5RRR0CNsnpjsnWWAJnl7wju1M4k2YZ9foGcbGyZWnn5AqqyH87moBvU92
BLfWmxN11yM+pxTf58r8sGbMIeTDj8o47h+kYiqDp/j+dqVx2p+vB8ycElhB7mka3FQug5hNreZd
AY3PM9Rykp18RiSGBUhTUfjeU+1WYd+NElVsJlGrcqwPzjcBHBaCu3OZL23chkOKOQOar97xcfKp
GZGt1b902HGjPb7g6XwEednu6X3FBmVy2B4gSgvaqIItJjmrmqoPcNemXP/GVYASwj/lziBbSAaM
mKz7p1vmVLIeqlEApJYLAfV/mbZQALzFjALeesr9JcPRdb6tkPNDxRRq0l5SVnkzrK5BOJgB85hF
a2PPUfGDRVbMeOgKuTiuGRwpOeh/IKGbF3nlePnBWAs55PKLCDZd/3D0hqkcm+scvbe8s1cnAN4k
nPhxJh1nNxG6RT6EphuWVcrhnb4esV06DPZEV7ni4CK/P71cPUG4bywowPFYPibm1Q1jT+iN/5yk
sw4A5H6PW1doeyBOD4LWjjseuU1C8I5Z2aUcxWyqUNLYxzoL48PhHPY0i4eKj5DkyiRz4jvJ4xTw
cqSX9gK1wSUH9yBDZJW+N2jNsL1eJMOM7wLaDsQjFWUDkbn+G2NbGbOA/kI3SCpLGx7LupNYe7Dg
71AQFxzZ2CSBcs/SR82MFBmLS0VUWcdZ2YHZNNcahFlek0M7CSc0TH9KoVmaj8T0IopieEpGyX5B
Gc74yj5+pKRE4A2Sz9EMTGaFh0BYHUghQGJUFhXAV0PM+P6IGktwYUwqcJRtnaLR1BvRTENbQqe7
kTRvs/6xkPJYQ258xMUSpAa5KzFnTdv5MPpOCiI/SENzuyCCbvdXj4zicgJilObT7VeCn0KMC+9l
1k05W0olrTNZqMCmjbGciA6HIbg/WelZrJcJVhpKQv6Mgc6Itjfzk8Hu0xSlIQ8yVDyPYU/icPAl
Wu37dgQ3kxh1tJO4mfaR8bfv161IiDiDJxHb/EmqTV6p1+451spfuDrEKSEa/Xgq+yw1gL4aq95t
X/b8yYN+o6VREn1++Irlho5qcOD9X1fBrBWkS0gBo5rjbOWeqdVOrxJtw3QbeX5iRMDfuvl4ZbZV
blpfCjIcshRCYYAcdwJkhfBuNWYN1aICdFO7Fyn2BCl9H6mOFrP/XPjCQJaQgysp+p1GmLNLJICT
4Ud91ukWaUVVRRaTmX8wS4vApI5WeNaezXOEg8oMWVwRGv4rgV7yP2g7C0yIFv38IF0HmZvSOSna
AggQfysHy003gVUMYiZJyIccuxhpaeeXYUkwoOdMb9Y7cjbxnlWoAPXZHDPZ3sXElwsEhicKIRhd
eVqpZ3gaKgKJAzVfZMJ3NNvV+FU5MbtuA1etdh7Zw4Bn+VL4PUUNhkOojkbs2ycw/mOfQqCUEIEi
wQnUhYS4Ef2EhuFaulfrg80k0kptTBhCi1l2T/iSFEawYxmkBk7FsQ0UZlEdBxuffHBKykqHqOF6
n+xrkWupIc12JzyUQSb0uS5S82VD4j2W0ATfcFumO8/uKTppRoxy9pBsgrQIeDiLeNresi2RWAas
FzFAnKZVpEBQbdfQM+fXvBaKPM7P2vKGOaMmdahvP+wV/pQqQVErse8vY109AA2JPH53rEwkAVlC
7y9mrRxFOCuv4zIFa0+xn+jfEae/E2XAto6keolW1iRf37ZxWDk9v5LLXhiTIwX1y+pHVyrhBkd4
XSCx+dZ6b7fJEusQ1l0C8vk6+tVnUUPrwYuU1wYpOWJKiYodvaHXQX8ZP6QxpMk8so4Q/BcaSCg+
wU8L6A1TDeNDVMT9dUl4eYyUkwlleYMkkyowNSzLKB/OA4wRqiZptEzlc9S8kc+70Ham/oqmXFdg
gzfRkNWQKvRdEsgUQMjMWKxJ0iYPfND2RrSnCQOTR5LczLxrRTtUf0cOhfanItX6NyCpYw/2IS3Y
Q21hmS8QKSsakUerAyMhSq4HrTdDXgcebw1Vv02pYlVXqakJe4a1icoAQFIo2EHPZ/N/x+QMB3Ws
LzAtCnzKt3fVW2hJN3F31rlTntRQlYTaJS60J5BrZMok5AWG3/H69hmyebfB/GEhcABf9rnxsrWM
U/2nnxLuXMHHtXVou4ZYfN7iSrNk4nAMEWkaP2+/2xepdK3JT9kfdGRja1Tvef36dqPNOdmIiMCq
WFrhhHHviJ92+MCyhqZq/gOkgiScevDcdS1f76vxz/KmCpDeyeeSoFul6zUVYmNHpud68lbX4AOg
zhg9m6bFGJkMkhlFd0tCcWyApnCEd3LM/I5qaBydFu/quUcEUu7fabEpY8pMCYKZlesELj1NKOiE
oTlBZL7JMeMORlB4qefNtsda2d8dNnhgMbmdFAMm8d8yJYq0Gm9ePu1FahZIpRd7by5jSr+W+DO4
kSRJMsqNl5MK9tREtsOsLSoEf0BUloL2l5j8EBbw/DBvEQogwkCuu04zRIXe9tJrfDcQLcLkt5DP
cnW8gh+Kq/A8LDEayKHyMcibO5jm7huaJELO+RjjNo2xgdx+pkkjyXBcdajs+BulWD9tNpuY1yTL
gTw6jHDwlZeqyy0f4vyc+oNfhFLwx0S1O/H1DWSsB/oor6AKNHWkZRKA2JGbkSF+s4b/HmZdBp/s
PgnV+igf0RIoQWA1B1IcRiKeMEJhJMr84fpSPgT0wm6UWdscHvhvKCPGdxUI/qpC99zV1XXjPkck
UofJcQAGZDIQDwAXc/pYo453Jn/dguElAOB4vd9G1DM8FEFcg1dTAdZX8vCnNTVxB/4rXN99mjVq
9HXr8PORPyq3f3Qa2SNIuMCbB5O1N1pjyqE8LC/DYBoMIEwY62wgVoA4pfPaGj0dNC8z/fhabw2q
1G8Gxmya0e2fmL/qO/L6/aRnE2F13OKf8rQoc550tuvLaeFczaqtQ7laWx1YvG7qAI2gWGuopj3S
7eAA0aH556xUDq1S7fTjgMwv4eqU3xtPvAPqqUGIkL4KMzYePJCQND1Wz4OfUqk1cIvDCmSShiKR
BZkVWzQR5gtgsi8OOnO63bA9nJIUwMcZeeNWBwXkwacps1yotE17VHLVcEb91h9GRufGs6t2v4Ln
xU4mx9+tCCPHn4rYRavA548gH07gBXBlYJonPj8lxTfFWLZCfY4lskpWwbg9HoSLqjgOI840lIko
4f9CHQuMk/1e0XSVRNJDgPCRHGSWhf58/nltm3obLOP50dPZBOdhJPGuawQo3g9Jt1xDZbx/4a9L
yXrc39laskENAVPjwe+GU5yywkiYv6XXzx4jVsvAhf5L+jLfVXHBvyRNMUhghQCUl5J/5942xsk0
9WhakFfuJVa1BoDbonnneWIvCDiMspZPlNivAV/evQQl+tznYiVySGXZgC1GiPQUUeSq6+NOKLS2
FldIYn9m2glFMxTGdJc9LbDlOKHrqgiEa1q7JOk/ZIhR22A+kqwAqAYH9iti2AXcp8MTSskiH06J
RQGYV5gATNnys9KsxDJsaONCQCXEMgb/jfZed3gQCydgehmmvTL9JOHSrAxN0Ov+zH5+Lumb/6dI
6EKiWBgONHTF5sF5DUeW19FpcDfoMBBlXlzB+Ahw8zEyE9q8Dr8NKrNu1W8QnwNb4uepWIafDekN
IBUo/IK9zDJJy0yjO6cPPJb4ewShpwtdRyqYd1+Xt3nbLgR1cM7Y9elwiwgJX99Qoee0Tu2rNiRI
Sibs0MXw3VtWqqTjJj1/bIlMMdW3a2RIYnJP5vdHxKZ7jDNdKUeKPG5uhdLf0v6Yd2pG1BGGUXUd
s9F2/SXp//W9Nz9u84Td6DtlKTynMm1SasfPG+ECszROXqaYmqm0vlFb5XeN+WDYEyeTHSr6DWyZ
p+N3uP10n1j7SkAopxxz90V99vERovRJCFiq1pOMNprmvOGVNXiwc27rlFiIC/aLt1TVXMmc0LJS
hstbjhVgauOw7tU5vX02rAnwDeLvnB0MHd6TwOLTQUZ2eBsuDd8abPenb5Aclhd2GDuAjZ4Xa1d0
1KNyFZiLwJLH/WY5OIsmA/krc2dUzdobgE2SfGMsWcJVPSrc5LTxeKhpc6cquPbp6VkqHIQfY/Ti
ap/iifgLV2DtxEAJvJqpbqRw6sPEYu+GsmNu3y5YD16oZPf2l13Hm1z3kMoUxwpzx0HhFsBTTVfq
gReoeLY5C1XMXG15GxcZitUgOONVSDBS6L5JYoXzwp+uBk9Jzr+plbnFlfUsTICLQ4JpOZnqXtMb
/oNEWM9XmaInGmC6f7zWIm/MHY4vFlGnL+OsRwxpOqPqyPypjkRzHabKHmEsypyndpJnxtqID7V7
ob03DYRbwnC5nE/g6VwTVCEwb4OwqdqCcVn6TrN0ia+QNonsEY1Zgk+1H0D1ItnzGkINLPC1h10V
tnCFD7o/QxOBuFfUEhjbYrAbYDUgGdFWBxWJCpFSu+j6z8pi9/nJdK3ZZF+GwpJQ+Nesrx1/UEsN
4SljKSikx6dl0n+F+c/VZg3V3B66AJbQQnytSbMVt9FaRc/NJ1InhTdzFnN0rMOLPmoSbbKCldll
XpXipwu1pbrWm4pScFmI1J7eqzhAxHrtOp9u5aBUNZAKknhntjlzR8pLlQ++A7hF3NOG1VlbSvSy
mn+aiWBBZFlLadCa8eSVE1PkqutqDVF6f2simNgFHWf2YyxjEXMG7Nfd1O5mv2BeT2DJ+J4ettf+
TaeuA+cfOvZA3TyxKkH/yFB/Inx87Rh2AsUTZsDAGqvPlS5Rhmk1nSm5wN/GHIcs/+QScaqQpJ8o
vFReFG+x3n+xJ8+9veyN7x/slsVzUfQ0AbhJPVD8x4+qFhbus5HJkUPj1cAaxpGYFJ7yvQF5Afbp
owJh3RIa51AOwQ30+dUjipL3SXJp9o4bahgQ2XviDbkEF423/afXB7NGu7YCtDCL2NB1yIAAX7nm
LEu/u8TLMWgDxHqfG53t5ftVl1uY6veYDdAXJOMzKfpXhujIZT65bzSSU0cDjwxpFZprl65XjKOj
A7+PjQnDzUDoFP+WLmGw2Otb7AIpN2L1H2xGBvU9b4rqZRgprW2MpqOHYcMlCknQX7zlaD1UFtDn
GOuiN0cUusKW33uVmsksEnp5ipwf65XyqdrXo/x9WInqvhijVBELM6rnJ4zokLpq2AYIdHzkJ19+
GdZWtaD58GnAFGOhA90G9nwb8VcQCGk2ZIAiSbgg6f4LaXPm98BwuAJNLB/c+qDszU7+9QkXUvow
BwQmRTbkSokk11o6fkHW2apIiWBwUYM0ocNZet06bmHmQ5JpB4f8eDaJDXJi6JQvNYYesh8Z6NJA
UacizESfhLPCVWY9IsFFpuDK/S5H7NkFGBBjyQD+BY5rUSl0igSuODq3l4A79wqLLhHvA1iw8Rp1
Xg+LmWndaxDxlv7bgDMEIAACc+ai+yvT+kN55iWlFx0o2Y4IT1+t/siTTglMeNC8Sdw/H6zy36VJ
la9BcWpVvPntCN5g9mAAHIVHUYr4QVd34wFewePCshehvV2lFJ4fuoIL5NmSQ95nO1Z7Jxv7LdF+
ZUDKlQNureEARGTTG/w9qfEDtF0fHLemjvUU43Ec5Ho8sa+QnufkumFkfHZfJqR9W3hOawFZVKrn
U8/NY87lIjipKX0P1WPsXqZSzUdOjFVYT5Ssyqutjxi+hcJCk/JWw8uYZmP+TQVIzTNN/DHN1svk
fw6m6txZTiW/4ILLDWFAqClgGW0Ij18yhEmdKz2Mq0EbAdq8H16yN695ro3oGLuurdKQAoI+tCdI
FF+dvj1RXy2YAab2glFOd5amcrUJX8CeloRXqyMiqZGN6YmlcehrsdVUeTL+d1RI8GQ4k80o7uNx
ueMnWhdbCL8Uhq5tqL/B3M/XTi67/R3OObjSLmuSFuflxtg8XwbjV7BMA4EP49vKKi75uggTsK0m
nwMS+m1ozMyj7eFvXrkNYMTMObHGy2EYgdlQlTx6bXohz90TkR/3P5mLkRpAUHdrKrVDax1Q5Lhs
4Psj1KTc/q5rNdZJL1wKWtv1PjsoXP6aikHHRW+tu/1rdNQSoS/VkGmjd2FnHJBUct0PWtMbNDeT
dMAkU6UAnHZCM/uL5Rkwu2iQFS+ufp02MG+A+JjhkkBB0Z8egovbje1a9gTdhX831gLzFOAzIKYW
XwohT962VVWsnPfVSEUPaBk853fImxylnjmhTzzm4McYHndRGWMEWp5ZUFduZkwPYXTxKiXq1UBT
l8lIFEEB+YW9Ds14mwKAGXkws06OA1maBlVQAFOVXNREOAQrHtDpr63AzBPb/yuLnf5dJbcilhz/
XOTwOjDHKB4h5X4bk4tnUP8UgQrLumSmIvT61Q8diiGuOsLHphhWQPzPN1PHUgC46zJtoXqIdlc8
/ekTwV4b5YfAghwdvKW9LU5RbLm55FdIMAg0V4Se9pLVLjZ6UqWWWIMqypseegIhOtjKSFnIdPwf
x/2TG3/NKWgp+i9kE9bTwDGznxNWjqtxphR/lWu9+pmDG7EpERwg/GmN5gysrgtkwvjwq8vFO4S6
kfdzlVrzCkHOGmCkTt+szX2W5+okZ73iXS/42F1aU0gmnHzk4g3ZjscFzzoaHYR1n5GM3mWyP+15
qfgw04ER1UudAGCxvOifdxRVfLWeBS5C6XkyvwxeeOhVmOoLbmrfUUvKjmltSA5HFIBd+X1+jNZG
JMvdLrTwgzIi4jmkSqSS/nYQ1So7DYmbXmxfX/r8D1S9X5+GAQEiSDkzBvivS7hlqd5o2bLZEQWE
eXapVo1Vf+agdStA97d9F8Xy6SvgY5XvowQSitImYGmcl5PrRAZDbhargUWZwNCHEIn5mijT4Qfc
kWisARwI0MqniNsR/XNjDPwKsnZvS6792E28d2m52RlNjLQeYAOVGHY001dS4ovDUUHs+vqqBUQT
c+m/AmJuJLzMMbOklPNN0D1uOPJqxneCI1wmOpWG3U+I5erqVUj1MDrv/S3eXJmc7gcVmBQqbMoy
Vu2Fp5YjuENAaV+376HrETWl67h+Ta8GRKeuvs/rAQGc23VLDe/e0y0Rh78iT5xC2Q8tN0yT9i3I
JsTV/iwv36r/D/BY6jeEK1B4vWpaQsanB+WYBayBqkhcwIWViFygSSbUE2Sh+Sbk5jmNBVzZGOUj
iOYY1Uum/wupRrgcEhPf8Jgj1sWyJBcLu8UG6KRw8U5MrbJ1Dxr7NFcZGiePwLPdL7vszEkvLnlC
zXkCb/a2ENvbdxUTp/uqzz9u7YxlSmweKY27WMfEhQIW2bzzWyeTdVfX/uXn3We4Jo/w5W5drKfv
QrZjRQOyn+F+Ixx9+Tp1T1ZJ2BvhKSuFg8JvhhS/kxnX43pbLnmoysyRwoyt4ytHhJblxIfGkCoa
VzRlhUofdMPxl1iMP3whdm49Fp28mBxvV1Yp8rXfEjlQxAZ+i/hpxrzDd5ZIMbu/Zoy6hZdu3ty8
iQM4MtlqOFmT2y15/nG/YE+f+7SPBYiK1Jx93Vl9Pf+R/X2e16cCqu+dGNwvXAHgva0ymnMYGPcT
J9Vewk9CSMqDlrRJpB6HApQfL8MzBCtsxUX9AOVSbtgp2nmpNvUJNa0MuPO/XPWS5jNXHUoFYNSV
HtUeln61/lFLiQIHJhsQKx9FS4G9A6RxxUi8kBR9etBGX4v+FUYPr1ddGWWiOHngfgIwHYvlqZQQ
1jHjOGgFW7utjnQ5BFwFfgqfnNbY6Xqp1ixZFQf7BaVu/jwv22zW8X+Jkg4uG8+YsRIjKkhflU9T
TTAtFdfnoW++ZSOEq6GEy2WMApaLroKcUUCDAcxqq0P+t+61EeiQ/+1TSW/hcRVFWC0JJVnnKRIk
8LisYBg+p6N1G0PtfBuFalwq5Ur/tacmmWzNENBHFyzj8oRo1ANWSrBPiY2PmQS3+xC4Rvys7DvU
TMrtiwbVcWT7ux8pv4oQuJsjjRJmrn6JDr8W8IoJtsGxEMSRPJgaMiVIIbY3kOY9xYF2Y/msSJsn
v1Y1TUxOSAFIrjUKkz+hwZ+W/mDkyKDogViWi6DsXnqU7M7nuQynLoLGLP1f4aOnUrgMkYtbhtv/
CvIYRhnEEMWtVHSpZ4Ytf6bUjmFE1Gjrm/lZoZXe7kAERkRsAs3WaTlffu4Zkm18rQYmvUnxfhzs
ZjyKuDZuFvueCCepjCygcwVTVlv4Yhw++EroL8d0PJfmHLcraBFxhS17kv0zLXHFpp1UWvahnQkm
t9udKtQOi9FK6zYchBRN9Jv588YeuskN6q060TmgCmDdY++AiFoi0ZDxSAA/+57CidvGrlc2sDK+
Xs3hhyY6do7vXsolo4AMQMI7jLO40wdirbpDZwNDp+M48wjUbKjw2cxy6UOYdxcQ1kjbV50ya732
0Q4JzwY1G8EU/wKAlvRpfQOQ94TfEXNjUO3hTXjcoX5RHTy5uBsmcyHeyg7sT5eY+IP/p8WJHYvs
mmtAWtwRC8Kna7FxVvS3xoSjunMA/53RHvuK9YbB41wl0Vbd1qFXDeH//KZTuB4PRwZkWK2U8OOg
cdxemFZlxBWYMnQX/Ol2T12omIewWQgwDJaU1bQhi+apl5bPDDGlHwg4IRdk78oaTMmSTAnbGeGd
cjhx4Qsi/6T1d+Ii+vcYr0Ec7rxRB+bZk3t9b1CWu8+Xg743O3FikYPzNcOQ7s2dj0OK54O/sx/3
DMW10omQQioQ5Ps/Qs1RUUX/yFUyZpPj8P63m0tgcOTHOojhYVbqd+a9N17X5HeYOFvlPod9nHeC
eMna8WmhjeEno8q5yJitXysqyWtP7f3QpXljmfEd9XOA1AYRp945yhcERqpQ8PElh+65mdLf4zav
0zGPvoVa2yMG3nPJ9jvq+TRKUvOP9ruRtOGnG12zfJM1BbsGFD3EVq95g/yWXBvSaoEYEieXtUd+
TQwvD4vO7Hyx6PHerI0HmL/w5vuwxYiAYxRu6PlTvhnEFcpfWyYgyRY2ATkKivI6gw8l/HkjlSBz
QUbL2dLm0GDNHA+hqYIM936A4oEyaWfpE92phy5UlsLLzT/lj7Kis2DeEp2Z9wDQr3dYewYkOYmR
hwyTQogeX/8ZBt8IuIElI6rADz9Ze2Su7iwPcjdEi4ZAjtllzyozMzmefbGIOIIgBZCNTpjB4vK/
QK+XVIjMq+xhaJMm8ihp9hCbaWjtosbX9ByrUAtWWxmu1TEQNTepA0mD974QfAFPGh0SOM90aqW+
MFKwG42v5/rZdbU52Z7WtiDhFLkrVmAhHAvFEKvkyDr8Ho66WYOY7Y3ZMPuYuwmreneDyZERdKpy
kC0KR/96IxrMAMApe6TU/uRYGswPPQbk5nYPw5soXW4t8/XNu8N9BQFiOjnC7O+mllDHatGOBCXm
YyTNqiUd9OqpRktB5dlJiMnyeNcOeToNKh76wqUSLrXVAx8PDc7Wo8NxlGBfeEg8pFacDRK6Kjx2
vpMFLKUbX3U/R92FOGm7BuXzB8awxXMOFrcmhMqy0zY2ShLB6hGZ0ju/hmZOmsixGBWh/ElMjRbm
KxcuDwAu0/ReUAhsmFCzENnKImk1qs6RMDef0vkdshHUDzP3UClebY5ufg4tvztkI+W7ZrwuDgYj
o+VgvXptILexr71Y+YjR7/e3OTGKxdKmHiAt/LwD1AZwhcpQpKvY6qjEdxJrUQxq5z0LjWWadsbD
yUsBF3fXmOthvYnQlXF3e1Z/09wGhMMK1TByR/tt/N4M9ulsaJYHyA3F8VWy0A7XsgegaoxzTi/N
FLGi64iwz8bn1qTfk/SXH7FHhWq7Uq1ObJopTOgl7y2F8HPo+f+G/2lfPGIwqV/dDGm7RN8Rp59g
CFLRPakDVZBiU+b9pZ+MjuAPyZTXeR4oDY5bGVA8lAce4tmfOTH30q/KhvL/Vfj5Vc6SXJuKvXDK
DSwXVOzqjkWBjVod4kbDsUAJ51lWLLBZT2aF8EExmG0elFzTD+CU7i+D1c68xmO/ZzQgr3ByI/Dy
PtI4nIQn44jDp1rFpcKJjoKH6fLJc0PfhUpL8fUZo89rLemxcgWhco03lrTuY1oJkxDXDD11h1oX
q+jI8iEYZFmbuElZX1k96/lE+d43KcgK2sz2VDElGaBkrspUXg0iiwLxsZmAtlX5TjDYLvGUK1n3
ROuBySROwAQ6uPgAvDCuKnTK8ykHZqrz2gUsLm2VGl+G9QhaoeYPzfbjWfGOjpu/27pofi5Vm0Dw
uscpKVNQkQ9VQrvt7yOzbDTvHjkC/kut/6OKz+Wt5kz0e/tHq7Os9xhzd7u7Kycr7Cs9s+Rnbiy+
ANUMsxlOyumHshcCMWs+9saPGRSpadPVQgCt9zyT9E0Z2O+AIgiZOR4jisAgxu2o4hvmz14spCHw
hEEppbYYGcIDn7UqcI7llLqQYbPER3s6NmY2X5FraJZYwqWV5JDOPjpNsmk9x/Kr+c27kNj5lG6R
r8fYU2EJRQsJhWoyyZfYKt0GR0A4Tl/atlEvU1Cp6B3u5rF4NdHL6ManAfMMLd5tUgl1HqSoUGFk
Fco6ZyCgTt2jOGeA6sJttZh/V3stNx+S0iYtR1ObOA0DomOtaCMoakQWk+m4qYrFo+e7WsRJ1nQ+
d77kl2qzy4l/j57ipIdFP3og0N3Lc+sOXYcQR2oM6ibwje4aNHYi7hRcf/rDS/ZvCaT771JKsJuE
NGh7n4OYmPz4lmhhi3VfrJwymYxJCxFD3jFG8cCoIIPqpgnYT6NeYi8IRcObBOQj8Dd6UFBG0tFB
2WE1oP7nn8DVjhWHvfm1AA+9kdwX2Tb4SBeWWX/c7NuUZzcGjUI2LiNj8NEyOgQn06F2E0MsThZZ
RTB9S3Y59phHMLt+SYxOvS7CF8K0LVu8MNMYJTBx3YzFqDK8C4Y/wwhJG2eVZiWm5emQ/iFCtWw1
6/ZkEqlfEeAmGgrBv1efG0yWJUl1x9gDoU+hScRDJvyiInDeNO6yYphz7EB139N6uAzxBAnmJsBW
0wT9xrQahqcpzrARRY8K22trCOVjo5yeDpiPxxUSSs7LONRJIgqiT46W9VwNEX6pLui+N67r3eSv
34+qAkGatPDU8xRxQiRrt8TYbbtzuFiUVOPt5fz5PVCbf6F8mM8I+osPHxoozuZ0+Oz/ZJoDufmw
hXHqui5KlOAoFnzkwPH4QR49VQvwqti2ajbgp6gYuWV27k2jEw3l+2Ev6FkBnOMKAzE6lPdtpgOp
RXhSyRIpc/LSuG1C4r48Tq9oIcnVdk9YzalZO3+y55MSpxhwE/DCVlmaoLYAh+1pdwZJ5GWaqaGB
sRG8EVo2ZuJm1qnh8zL6JNUhPPSxfNuzL5JJUZmd/QdLil+sG+gJFcCxvoHmayW/QoE9A5JbfRbd
AuS9P6x1vybfx83lDWE7sD7CWHvxO2oHQYCnjVNyVl/s2y2+qb2hl+urcbKc32yqw402e5dSRVZ7
M8kVB8XboTY4YhYiCyyCZp0nQ7kjFW3uUmJhNeMrKlsbXANY2Nhp1Q5caYt/z+EtzCSNeuqgnzY1
PO7zieRxcHueqIGcgk22vuqg65aWVNZR4ekTHsFgYCLx2/Yf1FGEIsVKlulu2l29+rmtpmsX0YmC
lA/UFZuqST/3xSiATNf+DnXpOLrQFSKin9ghkk6Ue6jB1UMCeI0W9D2co1W49B2XScs51yGGSDnT
t++8Xr5CpL+/EHtL/l8rRL7BhMF3lmRPzLzAHrOSBpIgTtEZID2i7bIPNPl5uc6+PwtTuOJEt3wz
WQ3Stwv0UUznnKu4jWG0y3Yldc7xacn28+r0y1pTekAMLeEMwYV43/vH2iF98/8EdEi4x+b7AOek
TlPfcX6vk03opHsPS9G/A4fCqnEYjDaRiELuXaCR2qE4Km7t0IBTLcB5fNpF7bB/vUb+69Eb4jUD
m/U+4KRANhpVrL9IJ+MGHcGHgWRwBuD91JYe2HHC9pmN3RjYnHlHk4QTlvOWSMvKDeJKuIN3L2dT
DqKsIGlTj7LyYIFNGWVTzg4tGPhVgfi/beng7Y0AEGuSIOYDA9SNGEu41n3mE6yKtPcq0YqE/qMz
GUzHBEs448AiT9NbNkBjps28U6drSAgSiV7/y8CYNDQAT4ZqKKzEF3Za1AKsUERbR868kB/czfj1
xJPmjTZgabqn2xVz/Wv9LoNZ9ixhSw8dYGULn2aQvpEtT7FQAj+mANrN8P2OqhRlfRc0xlt0XZYC
gkcTcOtWEBkrcHtb6kPVJiAkcNOv9zy4extSjZnkoiuu0uv6L4xT66fmzlCUfIK3CAxsrEv7Fz5k
nQMmY2AC+VgD8QlyedZScU+rr2aX9CKoE6SaIsMXX0qIH3tPEVyVX6tQjv/gTjGH1WAwdDvQDQPA
r2Enyb3CHLGwyI+gARw9vSe4cBf/GTDd8eoNFcVrgFuDvPg5SyI6/P3LZ79qcpqqKZlLTcRPiPJm
4Dn6r2tDzSqMvzxafojKHEI1YqxiO+SSy5D8+khIfhgO58hL4tOx9xxoimze8rYtT0IBeosEkrMK
PSebWU7gvYoOyiWbf+GYM11VhXLRTVtkpmXJz/Kicy6EzFPy6H3xsAU/W0m/mUTGM8vhvnAYhBg4
3OgVZ/NWvJHI55MgPfaF+0QccTcobIjMtkaKtgMBlQaozU2Y+sutvpXmLaRUf1xnKk34WrECOIFm
eKkXbnXPpj2Mmd8IR+ZNdRPXvKKIYePL0a5rIuyusmBB0ZTPUj+E9H4n+zTmZwCiPksnU7APFB1E
yxxAixhBHMUysN6cGZpbc+TmyH4ND9Wtz3xq8dvj/GK0x8s6twlanXwLC6fxfGufmk9cMemFRUM+
dx7NyZBNfnsWzctnyWv92Hn498iLxFD+kPOJTActbqeDy77btsE8x0B54KasIBYgL67lApPndnSS
xLWbSQpaoodbWh+0qrlEtvEdUzA7qZUST/ltVkC3HNjfyc8Xurj8RQ4kdQAbDGWcj04pC9oMNrnE
LiwAqTL2c+LCpu19OqsnQDX9KmRW9xOYWH3wqwjpl0rB12OZeupz+TxWacpgpKCBZEMkSf7vr0S9
KUit8cgluRMyMd2OnTXclJHbbmAt06kv0mJ3qWBLzIUub35kPbV9iwtpnrJ3Qvnyb0+bo4l6ZkTk
uRNfK0DdYR+r4GWT5OZA+ZHgK1KyIVMqElDAmaT1rAngauhiJcSZfHtWYdZ2x/bvTxOXqsF/wNAQ
bdKuPX8dGc4V0qdYTY46fyKazMRM+ExSv0yTrtjzQC2Cl3Xye4LY8BkbmJgCY9INYOESNmu7wdpp
jLE0DylcqPQUuvYOXdU9CWIl8Jkz2y9/xd/s6Ni8cWAOVjCWsoyGuhl4HvIbjK1M4UO5C0DWJx/3
2r0u3SIJYiLw7xvaP/YxzBfL+oWSUpfCIHoEuLnpWmy7vGm9tnedJZzBDnSOhQQZWZ0uFrmJhhs9
0vf7+C5ESc4T460qfWpVD0p9yC7kgD1cqsJR6xHqVG09v6yLdEW3q0oAIsrRw8X/o52EvFehprZP
jzmHZ40lE8aVrolSEiYdbgOuWiReVYVDlGaWv0te+qZN2HNA2UKmyuJdFmOK1lBMiFxqXsDs+DHV
IleVfdycHcibgOwAanolcSP+Ei1DA7ZosaTDdKyivPa60Y6GcFEjEYH0OTGabQXaOQqCxuelL5Oo
nfwo+nhhyRA3s0UYZCGDPrxVQK9DG2ygxZhZHf9gn9X8FUzd9XciWaYoVcmmRWUbW3UZ3xvRkQZI
BHH/YdzRazn3OIn34po6hI4Lnhbm+Dayd8r+T+Fveg57u7N3NhBkWOi4lzIfHLzRDKycQ/hH+PVn
LMVg/yoQ0zc9+WMuuPYIsvu8oha7MOYWEe6ro+Rtl1OHKYUkPXY19/kxiDF+MmIKw+w3MPNeX7u2
8YensvQztraQ+5NjijAan4i0ZTuLLA3tK0zsQA5c3I4UesSzmi8XnsO9IoLntVTXGehyj+kgJIlD
qQzdKd1/DBB3hcZAugpHKP5sNzeSSwW2q/RZvbocNRtc5pdGhsBeklE89JdrjgGADeAvi1cByuXp
54EnM5Teae1XMPgkAMbQMZUmUxq/+QnbF8uz//zBmpJBWjwpr1GNJFkb7Arj4pBrGThBlb/ef5Nq
t7qbijEfhu/a2C+1F82NULi1ja1BIo8yVggLbgrXkC2k/NajOWeo8xZmmq6FzhbZ9fbaAbRqib9Z
tJQ5s9Jz570P0tOCC9SBVs7oJaYPZ1CBkw6j49i7n9Nex4D0LuM10AqHmzE35TTuRh0uSWyb4nzK
IotClytjvqsD8Q4Qn+QIHBagQ4FdQxB5tNJOA62yUvgdSr7JDonJUZr4y6YeRxe2CnsjKnqz9/8A
8BCFqcDjKTv0JNz07BmUaNVOLTWlre0SWQ0dI3nJ5fzvglbdJHQSy7LEGB36YBPW4qrmPRAKoYct
WAmgdi9rRn8lNJAAPmxzotjp5wd+DU+HW+Q9rsFzDf4iYCRhvcAxOktnRC/lsipZ8i9K1B9YaEz9
ZCmmKeAjj07NqcX45oJpLtovrQRQOJNqYed1JX+wS4UlWtSM2jKhpLDn2HYdnW48opAnoWyFgCmL
Hsoy+eJSu1LWICBv4RC9EAtjf97f2aQ/Hp51YZMleEh9HFAY6nlo2wHGY53CWpRkLlp7nHb+Kq2l
nhtr3AH4j9fWM6+k1i4D/U1ncVNYN99zwx6D9DAumsLb6+q1653R00lEYNiTA9pUmnPv/HlrLGZc
5973MxYvBfJlMiZfn1+5qihUU45mcfVjpPxJ1U+4V/L8DQAPxItt9f2peMESuTxfb3GYRfT49Fwm
tUB3HAqQMjlYyW51ccRvdtdAYiBRJphIXXmEm2r+Cbhyz74HwWNLvsSDy19JQPl/M15IYTH8HFJt
MbvR34AtkCX8872WotZeB8KZngFh6Y+lQvCf428P5x3VWyfIUxbes126iB3wsCZDZUcz1GRLilQo
YKMbFltFD2zhYWWPmf+0dkiDcQgqyW9bkjGkVOxN7APwTd3EF5CoRGW3MENveOJzsFZZNTV92vt4
3M4oOcQvZbb0Ar7FkOyj3cMrrn2pz/cJylKEYXKZLv02lymYwPOQzEEwuosRWA9pPv49J/33rJOO
ZSg5qNSGnmqtGLnh79IQCyfaqGN6EvnpNQowkSeHAbpv7m3XXIwbUeTkltt3+9erV9qd1MBFYsJj
78IC2KNAbDMJ8NjuoMZxHb16y9IgM8FZXj2jaK+7fTbW+m/uH/zh59uKrpcBz8InAkwn8/n1rd5Z
J40BVZ7zbcpSVafmfbEGLkhYxahQ4ME9xA0aT2GDm/K6KESx5R6vDF4Y7stCBiW5U4KJbFJNShI8
5XD9FblAGfbHQyiEamu3ToTo3/6p+Px4vtzhYs9xiTTWHJ9EnM1w2hSEM0PtnltUE0UxNSXAJrBN
aCCDA9aHvT3lrQMxguYSSXFVZlCcKujJDS/kg7Q6irFcvP+Cli/LMM/9+shNtaUJplVH168Mor5Y
l1qZIxWtm/BIED3IUYMfIOfI6NWu0B9vQL9nW3VET56e5fn4j772bsNQcLtIsrpdhmmN53CSfvcP
1ONIPJBadaQRVKPaf2jVWYJasMc2i79OrRZBBMOEUImbJFwEF10qc1Q5itN2hYQHijcDZ4foA7Dw
Alu1t5xNMkpvqAy7+eMjtJy1gJKW7BqjwZpJtadPYuq5ty3BbeAiIH/NXofjLHigzecREwZF8LJW
ZNNr6bYUeklOOiJafD9FY6dYluBspcWVWnFd2CynWTqvwS6soHPuNRWL4HALdJUZRaq/4ms/4T9q
17jcUOTz9d1jAQz0pfOZ8gVzwAhi3XJbE48MwYJemiWXAYiQdhIZJMNhpvuOabk0gvpkTWtb5Wbv
G0T2q3sY+eltpmWC8cSNou7lg2wiaDeCdywcYxs3+BOzpSaAUdzI0olkc4QVcOUgJNXN7A56OcgE
UcpaigpXz5n4q2qElN3nzrtE4dSy9Qu+4VnaRb87Yt3OArBN+rWLdV1osTRj5xFDQKIEHZ41nsmj
OydrjrCHL6t3bHGN7vRCbMX2+BfS3Hj1UOcVegGakZT3Id4HwU+IuysW21MUuaozH3gBt4WdcAPp
Z5EEGUKdLRVwl9CauzOAQXHuwIJ3YBiQo+U9SJA5TWcAKboxoJ9/lK8vq3VDC3V/0BpqPiUPG5Ci
1/cAYXzbglIeMN64sm72xnwrlGee7L/siAzQaarWl5FE2lojQXNujm3GGfI+4wjvuSfwJX+QhTwO
0hivMXFgv0YztDr8Kqms1MGqnbmLFcOppuTDTSndvt6p1h8j/rFe3c52F0uFiWuNTwD9Rj33vsR0
9eOwcr8QjMl+ny3N1vc0DQeHROMVgMrU3bjiWRdid4msCINwgYU6tNgYCE27OB4A1CrIJR+srcVj
0iq01eaDvMdMa63SJ/IbAKqfD2cHcDXD0JEeNQO7Qgp0Vgif1BdP1POvAXq22v+7UfZWaRz3XDJg
xIEuVfCvDcoChB+2ZsoO3BAkN0pevkxcmSIqKHF7a/2d7KKth2UY5djScFcj5ZZ3f09hiFize82b
quxwsXbEx6wll3MdXu4k/2qiSy7MI/4KiwbZTkq0BSzm+/UjYbvLWkEsvB1XzthKdkcwnOrAFsYW
BFm2fM/ET6eiEWfalaxWD2mXuK+rGW7PBv+H+r8Zno0b1mv6Ga4cs/M2AgPx3IP3k0Esm0ZJizVd
HzvVdtSrBjZgBb10brE7GXmEl0at34QzIjNW5W6lZ/DP9rEngDf8f8fR8/iQ5ZUxWgoxvcWz+Isb
oo71tZrZVWYEcyezQUbLnbQnxeAC9VV2+5jYjDeHcGDhthb4hujnUgCdW1TAU2IS8Z1dXIxClmiO
ZlfhOFUX/PAV0Dh3kCaVcfN8V5RkGJh0KHEFK+uapGWRfv0LODW6VRF9RqOLr0pmIAx6xlud+kke
imSmnj8GonU9+XYLCxU3b1pMnYe4B0PlDQzOPm1Ci7V6q6jVYjHS0kvdhuKANPYWV64Z7ulCOJnX
6pJEa6OPyVDz1EHUMf4l60SUcYS6n08MoODzC3qDfNcZLmtOr1GkxMGvdNf38hsUspqreYp0kNR5
Qi+3Uk6yKVPGNeHxebdjq9UGwtmBg7/ag2ToejrpZGCissQ+LicFw/zibP9xecL/to5qpizTr7hn
vx0BVEHKXzcxf5oLURpRZDZOlI99IHtiNhA0uM5S+jPvDOjywLZECltzvetVkD4IRUQtPaA9X9Cn
ct34Rp7nkdqEIKhssVROkrVMrJ871lbbDLvIoGVXT5cfJd6r7FqBAHVdUPi2FMQUY6EDjKb9tq0c
D84DUTDOzswrLTn5dUK//XFB57DbsZLHOSuDw70m8yNHle53IkAZv3UsCIdXBwYYK0rAKin/3f4m
8AsOay9HuPO+YuHJV8IGy5aNHe0AA6AF3NdQhhloFrctmTodPMmww+EE7Qri+PymVe4KSBDvh1mn
psNr9FxA0PdbiAsmSEEn5Nd9Od3+1GQKHIB4tybHkzjkpVMlElX53YGk/4z6/BZ0HHH0gaoxtYrq
OeCj3vbQn2aMCscAyrY9NM9rgAMYN7PMLOeY97cKQ7EdQyBm0iz19ezyrIcEsKEKy+6I852NLUOE
mrisxkwnm/B2WrdAT0wOWs0m17joNjKDmadJmhyHDmKkM35idoicAAFBqXbUOnVIf7ptw/yVq258
NuBmD3YZnNXd6EjJ5CtjIZi/ckZnxlqJ59cvcmzJ7HfAZWEHfag7rD9E0yckPEedsco8W/E/H2QC
5MKH18td4l7b9HNRNxjM1yTcZ87yOGYs8YyMcm3i4EGec5kA+NIazwicx/J6oIDNxL+oq2i4db6u
AQiMsWAiu+0HcFQnigaCrRIosL7bhS6Qd3TQ3xK6z7zz+68AMkS/kChos8hgGj/C9kMVUaQpZEnx
0ZwM+D21Rzs/ftYo/3M1sz/K8KEy04mvslNEvRz0qEIYmmp55MG+nePa0H1rW1m26D7Xv1yE+7pl
ObFjgmhY/iC6avF5TImG0a+CIDcPe9aaXnviVdTXR5pZ452biC55aE2fDYAUtWCIP7IPypm9zqeo
/UsOln3HRuSp8agWelb1rYOl9dDwqWrkHm2ADIqk8jSOrLFC/vj8ytbIMSWgq6fqU5z7H/bc/uyK
QQ8MvywnPhK476BnX0wVzhBo1CuFevtHyJkE+vr4vT/dOJiVbON49V46CcxjYvgpJjRsATI37Oxd
WJkIgD/MAhfdLyq7xHJMQPdzh49+ux6pVeZAyOOXPueMbrlyxkfXFxHXH/RLD131zFqhU41kJVRV
dwgdCN1WfzV2g2OAqboAIZ8B6f0BPLFql/C6BYD9MwRUlkqtF3jo03Qjt7gt78RTPDq/EB/12jUg
gh5DsSzfvPvRQZV+0BnUs5qjHZRu/1jgywDhF6foQsqJH82AKH2dQ/gSYFbbvxotbqQeTZc52laz
fq3nd2Vr/V9oYo6Em7nFkrVS47WaooJYX8oAmVjhAC5cb8ZVTt4N4LsScJD+Kb5i+9h2LR8KG+ZG
NvU5utbQlf16I/E90KjHhcn6H0SZVNh5QnRC8aNChXyXl0g/MN0a6FiWqcNCW7t3+/62ocGpmhLE
3gz6e4U5xEP6s6vcsCZkMKnWSAibnFRO3vsTvmrMWslucM4HlO9ujSz4zF9WethqyTOSo0lIphZL
OED6nrBja4DJbIzkvnPef+eekPTGjrSRTUJYK6Y2QwmKSLDVW0sLgdpuvQmFq+VbhO0zPIhvXLd3
5xYa4lTZxhOsJwDKhyzNYCo1pRVRsBJwRk71RciOUO4HQt/OnXaUNdstI4uUtmoRSepu1GRkabHO
IJVeJTboaNu+xjOe636cZP8uINnxr9/5YwfE/Cq4UsqKQCPj+zepz4xBQtVCMSKndTg77tu7ymSJ
lVaMEc5Miz4b3gcx6jeybRNSqeS/tAQ6TVBz8EXsQ2fX1dv2HB3HGNU6HPH4ZNBlqH3i91iXzAXb
2WEm4WS88qKY+N0c85LAPA3aoY+nwNAshp+AMiPTK++pLFOgYu2mpWaqdRcYt2gquCXz8VQ8W/Vm
8uXR2J3edUP/tCOiMpj39sRu8lgHMzI6AQEomiKXSaUOIJdOSm8m/7fGA6JZQb6Gv7bLcHbcZI0i
tJI7/ZCzTWOCLANY+toW0R0lNJYT0wQNVf+aqKBaUbrZ9muLJyv/LdlPniFq6q2PTV7zxhlsFZta
jw4NomMJaXRHbMZ9klt0Fb906pTdLsCp5+tNPYoNcDCjOM4AgaYnswRgWImGK5we0lTY1R2SFaXk
tIQ0qnbtVUli+wNeWx/WZCxHIKkOS7jWGLeul75ux6hWJU2M3rXJhthFspu9b6Tf1o9XPRMVpuus
Sij+jgwDk0lKymaMWtbh5iFpQSTqNyl7WTJnUGZnhxY2hBevm1SQlbAoiNECtVVBM+1AgNXvesAz
CoESgNvGqroBsHZ11Lie7FflU+07dS8e5opzF5QkQW7KVZnGMvZbHewVJya5qBNRTKFKWg9/Mqd2
65yUl7BgoTLocYQGgGNl8H960o4ukJHTJ7uSWZVORrNoFkmMhZyylJ4Be1j0y1ncNBZLQ43rtmMm
XSCDnKPjwEzSuT6KBKcmbFTwrhGuyZsQagTwDxgscQQUiTDZvaefU/Zepoj/vWMmBxb0tFT9k/qr
rYl9nIW6/8Ee3V7Y3UCha206dFOmtv4GRqv+uwQlNPe3xfxi+I2stuxHYgCWfixDFoWp/o1IVplU
z1Isjv9VrUYGTSUxYzuvaIuWruQv9bdE3fKYniT23Ky8hjE/q1HHPv7st1LbEav8HDlkZ4L8enFi
Dt2Vi7az0fJg/i6qh25enKK5aFiYXoh1gu7mJKzdR1Quu1BL3phwS4tyWbwsmdhOimsrS+Jx3gy6
7PszzuNsOsAuEdQmBJ52CgVyizZjpYkcaHx/yimXsaqjdyzVPdsY/fyTLiPr8D2hMB6J17djJh8Z
T51mLU6CUh+1RuyyDGbZemWH0KzHzGyNAocSUbI+swDp66bYju0fcD6KOd12EHmUqxdLOp6TZfNI
g+MUFfy2budLz03RaBEXV0pqEkGqRnJcJhw1jFQ0DafvV7WscVX6Efp7Tbi7PdHKHg8QojaK/9sy
qsVj+xsiQCr3HUF3g4eLSzZ1MRuqRL1SfAX1/BhAxGgzlmI72neeL4x1VGpnUToL9bYG8WoiN2YS
PBeMJqexUgLm+LD4O+q4vTWs3pHbt6wJKV6UsbekbAAo/yZLaghOekpYlaTA9k1ODU0+9q9u0I/m
BoGvXqE3TTK52xUJjUmD0mpzHhQ4maZGzESwQI7B0UQfAOtvnz2LuMxCdsu5rqmzNajYds0DH/Pe
c5Xw7kIFQM9wb+wE3OkrFJz9Da6HD5lNB55tdOBgn2XrgClVK9X78NZw0TaFOBYCZcXTVTAcivbb
P8n4BPcZUk7SetBXvI8wAEw83JgUUN4klRQts1VcsMZvrOHDph28zJfMFdzGCue656CwroYvXNzf
jABUNN+SVjqgHVPVWiRIH+pdWGGg8Xgw5aFDjZf9CyAU1zCn3KXavqdII8T9h8oXtEM3r/42A8Jv
Mv/8JO4RMnBQxumNnu36Aqa7sAwg7aD+PUGJL6wvTUkrm9Kkz/1u68xkmUfgD+Qz11hObdo8ubu1
QeXADkIfqWardDmDMA2CQHdO8kaCphWIM7OLnJJWfQwoUrHND0W3Wf1sj8+6URbDgAFSWy26E5ve
U0zEH5N+7dQLz5G6IBaZk1kUv++rARcat7AH+WNQQWwfSzx6bZBzky8z6zh7NzWvqP7fleWqC3SR
xSDvQxqoytMnpm9wOPb/dcwOrtyWLqH/H9waoQ7d+6wTljUtQ+ok6dDUObfCxh9rEovWTkMswEE/
lGRSvlMLnd3Oo1vDd9bLw3l0gl95YDAaNVGMTP0w+kgvOkv8gB9dhZtI2wZbgFzvJ0buyY+ZmiZF
UI7mdDMN5+JkvGtmD9eu1ZENOYaTE8wLj9D+e+w4cLLfhBR1dNGDz+YqDjk/B05uuY7ww8TUKO+g
LgxBhHJBLwuzPaMW29//3cE0wPWGXaL182LTreFB0a3QRusLCeZ32KnfYwwqNBPfEwMvamTsMYh7
Ug4GTxh1c4Uut2eiIy+cD+tTm3YUNyzQjOj/XNq7/xyTY5RueM+p4nR3nt2GZDc8jp5lBJBITvUQ
UMCCLH1L7F/3a5v8Xw78QeeOwbskDwRCfXfo/WbA6AkV80heaeBDnn6+DDOxWQAmbMR3y6MKFYNc
Qbw5TwH+6QquX+mNlSBDijVTkPNXZClOT9reVjJPf+OsqjsXDJTkLzWbcuD8ZaAyGp2Bc/BVqpXV
fhKpEScmBSd2swrT9WBdkwjX+3Rrotj7MxSEN4V4Nj3xVSUAvSu/gMwybs2CP2aHPYlHnKM9ygNH
xABMcgsiTyou+Vi8aBa2ehl+jOzMGd2P88qW2Byh2x3HSdACD0bW1RgPlHGNAity6DyI3yUXOwDd
PleabubsK2lx6rT/39VSIBpNFXlB4RKKDCVg+rmW80oV1sF8x268tstZKS9u6YKd2gT1poy4uy3R
jmPgjg5QCHoOiXOzn6ObRoaRVL4Cv74o3HOgE+CIriFOXDtO6wAYVoibxPLtHhE+I1t6cngVTnhE
8gvf3Gbumh0y4dEOr2rD7yVaf3CqkMJUZzUU6WOFOyDUKfoe8flKobQjhttVY0rpvsn2TsS6xULy
oRAiqMaXdMnjHSqD6LGeibiCwjAqhq3Gz/PtM7uGI7HIbajXSNUDmSoIrizDdF/Bqak4hSSvV+gP
ZI6s2EwOgXzXb7wPIvq3XOHAOav2o8JVpk5M8lomjpjmqydE2NX6KGfgVReeVDXuV/8G8wv4TTx4
z3SIRWZkc64mUa77TxgTltXln5Tg9szDPjZxtdUk42HYv/G9s5JSQUnyssEoRVmYzNuoK8jjTviT
1HkA+HExqTneNQsiwDTEUc0W3hs980v+d1KobHOgevbHLenTTqD2htlB06iZVEzekbNdmUX8X62u
w1weLOxRcSTl3JIEG2v4Ta9QHfln2bAupdDllU/A5U9/zwsCfBTwCuneLOzlJMyofWhK3Y3TAyWY
job1lnDsEeCVR39nouaGCBj0w5q8x71qZs/6x7ZCZ7rYpEDfQCGx48VqlAhfgKROYhzQVR8dZsL1
XgPca6J06XhzLLAg2Tb+6ggzYFyFDetkP/LDqPO3b7/t1vPUAueYbL65kkF9BqOyeSlbtdUs9hAQ
1Q21AAjJw8RwFkPuNwBGvj5ul7coQLFTOHRZu6V6CMorQfwlnmxA0J8AXd9aqTyNs0FTm6QdTUlb
25DOMi9wHFqkxKs4Bpyf5YuS3clgIIMSfwDItOEZilrlVqiuhE4FM2QAG6bX1lshwk9ZMP6uRruW
3K1a5m8eivu+qeIFA+fmngEJ4qB/zcPCk8axMtyrPhEUXwCIJ4oxEi4fz9QQzkYGLqRIEKENQeUr
pTg1ZpVZwccWAdj+WGJ9kPmZEnNA7F2EFamx/1IK1x1bn3k1tKQNHns5EIMetyYbC+k1ZRxK/QX1
4iD6khUIHKku0h8VHRhBkcJ5QKrPXSuhGijeWBp8w6jRE5xV35p8BpZPcxAYHZQNmo6CozcC7nGl
8ahdKCdYPZC5VzgrpYeH+b1T8DGRI7nK01sioZhkL2H0dRnfW9yTzvYFD+/LL5b8YVyCO0fQh4iI
/NpMQACMS2wFFe1EgIte1ko3y9PfTbfoqo+MXU8rV6Vph9PGzvI7K5WsFwWsh6d1Y9mo8ePjcCOo
RAlnjQEHL86EyvMz8XQxY89e6IoB2U84i+GvB46H7ser/+alTWpUYe4Ij7SzCVzAPlzT1k6x4eVF
MLeiuwlXqzSQ7v/nt0xe/BEf/y9gcbsb5e7NNTqGxArQaAJ1FakTNKcQRsE91VpKB3RcNNG+dUhJ
+1/sqpZQSbiJhikuMtFObfQOqZB2KoP5aj3QrED+jy+q81QE7DShF7xFrRzoJAc3+Znl+IUArjn2
BNniiMRLRk+1hw2Ce9AUnmucQEDiw0EvilolcrtQuoxOUwL/F/bQU25PQDfqwmCAxaE9jV1ygjG1
tLf2ShZRwZu62MjSK/7YY0pLz078S/dx6l2yxa/zsOFNaj8sbl9xrrw2K22KLmyKPiyh3ifwho5V
wZCxvwVbB3DRrvzlyu8qaoXPv9y5kemfn8arP/m7TYCuhLlXsL2FKm25KV8kr7I3eBr7JdKkXx5x
062DJlah0TKuhaCjO1t6kpzwYhfM0eFTDodalOEHhV3i3n63zZb43vIS5xFjhDCelVY9V5AqtMWC
n/exTGwKOqSGDCjc21yEWkR0XZEpesKotvisBZtS4lfWanx32PY7dzrt/FUkqtFpZWIlKe5cneLS
/aip7WucbL2fcSXngOBB2BYMQNGYXzkyLlJAOO1gU5CfdfF9805oN55zqPkkDeBfHNLHVNtl+LpZ
ZZQCFScJ7OaQhHve6VQaweXZm7/+7gP0DJFCCwj+x5b0C3stzIW9QxID+DAXRPqYWw0Vc7REUbxD
0xlSAYUv0JVYWiHJL3YQroBZUxqlb/seyJ+86mjNzMTOnQ227/ZbO2c/ZhnNjkZUqqBmcYgWYF7I
9mrsYZD6LksFN6bRmzpFDapVRNPi9wd9wnYl3DAoM8bhjIfaJJ0c1d/qxqbWaaP+fABwB3nLk1bI
TecC5NHG8yCSlqw15WySAndKtbXUs1lfQhaw8lng3w3deoSM7Bn0hb/atuNDg7a+lEMcmUluXSfQ
yoXA9zkMRqze6VEWf3zBhSt4mQiD3z5oLSjZzjOWAO2BIiY4QtcP9mAU+sRh53e2ReAjDemYijgi
jp6ymYDmG6bC7aoTBfphB1umHBLaKkGb8ek+l+8i/x8+HOKQ9R1GvNTH6IZ+wcS3HyHxyEfmuL2E
5f4ZugHVpwlz+hRoy9imdNN34NsJcP0cb2kGX2J6nKO1pSz/qBVzQYV/A+cEakosBPr4WE54wQEK
mH/JxjBhL0OI14s/yhqyTXGZoPjQ2qAiO8JdHNJe3ZbU/43MxxX3LCxgj22pk+Hin5OsqJXzXckW
8qvfHLeh423xrwfdj8ItVsxLxPPXRiAZGH6m84/J+wT7p3TI8ym7zkCzroteCj6jA+xbAkE9Wclh
b405HXpte8Yus+WpRIJeALO4Epo2RPMPx2SWn4tfSGZndhykcAcnFaqameet45FVoTmhvPW1+9uH
sziRNq+RkIWBaYiP/GkdhUxyoJBYtDqYOz8b+8Rqy8ksknDUE87Ry8oi6OtlvOFFQWc3XBsRPsB5
l2y9OG0A8Z6r5SSZQ8xpZr/HZ1hGtkAqM4R6PZ63tLMQQAQ0cyMo2jWuQr3Y6n8gkqgOdQHCLNRW
++eRPSJNL7fZe/9QgdrCCJZ9v7BTWnNKaopKLJQua03to0fNrBdw93RBFDQzqVnSUm4yhV+RJp0E
gNv4ucNBvamrbsK/GFUfpe8VWp+URY5I46VgSd3flupVE7knaiH0h1iNQtiDJWcrxoH/MfVGeWcB
BnC+v346/FA0xExCA+01ctWsnFI/kYH4W3KwO4xkoVh6Flm/IUjmV8oJ7JHNf2d1pp1galNazuXo
loOiqTJC9f5gJNSNy51ZbSfxSuFK+/y8c+RJeWt0/rwqsRm4e7mrV6m0eGpcexAzAGRfttHwbisq
N2753KkShfYYnzImWF2Apirmq5GyKLwK8lims3aMpF0wuFNZTy4raOf7pqdi6hn3XeOrGqsFAyGZ
I0Ag71RXTL30O0O2y07EBgaYmb3mgTjgxR9G/u1wsOgb2+vKNUeFMHlfPuDMDehUGut+T7H0JfGj
4/1ibpFI3rKBaaoqcfOHcM69HvtanotrxlAk4XWIJHRFrj8bOasmyBPfgDPIe8+OpeqfciocMUFo
4F0oWCK1SZaJpaqexWponuGsuaRkxTOjkYnlfx31kS7cH+nI88M+CMH/RCMiAwy17vxU2BWBlkob
8TRN+49g0srWmRkSV6ajTMdq5pUxYL4a7z8fYFThiJmkMEnjDkmBx44c0XLL4Mg3jJhJhIlcosxo
Pps580rC1siF8XQ449V77EpxnOE2rhvZNY+KjmwPGD02ZVTbYk4qgUk9ICLMl4pPPD7+KL8Er1G2
hL2o19J9Uc5QUAorzGDClUZlgO/vr5C2qhs5SspqBCOruRzow3zIHVddwKdlJPCIX27WVZpDuj/y
hgkpnYfY1kHbmlyEgtzG8e114sLhrDSHO6fbaKeAYVXiq78e1PZFtk5VRgj9XYMjyQWooG+3lezx
Ct9vT/OhYt4QWdWnZMrA4eul+xEc2KOb1YQY7MbGMSQUeHyqk5auHL1cbMu9+Im/wyW710cG9wxN
2/H3lHlLrT401rY2MrLk6p8ngx58Ydzm7pFqVZp6EDm7p7hoHPZ9iK6XFZ09tp0aRg/+Crlwit3q
j+u1yHJ7CjX9HmY6IFeGNNuuzrdo/0ZIn6q/IgeB4ylMSY+bX27FDpqno/s5sEjYnm+TGlLyqvGn
cNEHm82SrOMw0WNpSjHklQH8y2SQc9kYv9wSNkwJX49IQQ2AI7MDqwt6KxebA4YzqIWecFBmWRQN
j9TIJCv/BylnVb1raLQ0+mjMUuWGAWDB8CFVvZ8Z8ZS3JEF6O3+3dwaHa3p0jT4w29E880L+o50I
Bu2nkIzZUhkwNqYCrq3x0VcGd3rTs3xkeHLq/IRq0/C79Qrap/OuVGvJZHjW2DOXbUI78OR2rX3H
XfkJBEcwJAUp6TO99ADcBpgDXYTG1nUjFaS+/eegS/W0alxgduK32k5jmDeRbZuOLzfXRiqdKviW
bi4nahZx9SpOytL66gkVuLSTuEiohK7NOLa72iVbDE+GbUnr+fRTF/ag2O5NDuSeBavX0DARIuG9
WixultPzSZRczCxxWQLezwy/HMV1S/kYWi/AeXR/rc7fz5yTvNN3EbwdoZVC0JlIzP8Xq1107tG5
REdD7OTWy+n37elLvgorPuJylEG9dMCGEkTHp+lsjJc+X+5wZtMhgePK31B38RETqjqel0YDJkZV
SISTh5ouijmF7Pk0YLRjpTIypsegfqC6wMh4+GfoAd3e8B3B1N1XqZXxCrUCSTC4C0/5cJz9VzfY
sixBoaD7E4K8dgSY0jFyxua1OgkJ+0WVyuBzMJkKsZn2guof0ex6hRSPwj2RpW3TW8Wl+rgBVgKo
D3uWKd2mGVOOCdPYwtwILqfTbKv7+RoxCEWNM5FPJUxaxxPG77C4FmMn3obvws/dyayfoWjF+cNz
jFWu8G3owTzTT0c2TOnCa4G3VDl52ab+TYTmdriF61Glnf4qWZ5L0uY1qpB5Cur7sOkheHdo15MH
59KbXL9HDP1PSKKgNc7aqfGzbiK54aeDZ1INIaRGo9tSYx58iTRKqtu3niZu9zKrcGnC/wGYobxx
PiCMXI6sCPfdMWoVE5xYkYj+Wia1BQAjfe3fcWEhU3tibEl0TM7JBqA4oQP2/xBlY7HgN+Oymd3a
PG865nrIEMlcEHMY7qTzrx6HHGEIL4duUfnYpRsoLPoGYiZc88s4NYiE/Bs9ByfWtPlQAc3lN43t
sLbuwh7CpGIRdZfYAEpGG0bBoRWvDz/EUibbQhs7SFEu0jHYt8xjMZochjSVfrpjnGL69q2aIerp
DKIJmzaN/Ge6sl8508JE8RF6Mo9p9vDqRsxMvHr71Rmhqmygt3uGwDgievtvbFXGsZyfi/fVXueF
g6I9snzIheYnEZcnuHkjSn8rXemnV6ghmqMPlhTYjQygDMFFz19MeMNtcMHdT3OccGTzC+DwWtDJ
W5/eobNWjNfWsRtg7uYPnfRMaubkINEv6C6fQnePLUBH7tY4sQKuo/xcu+SXEOXrE6a6zjCcrHC+
FmvnXHFuxcmKzR2GGEW6pYG1NWszDSISVi9YLZZAF0Nu/dJ/iSrjA6sigo7P8GNg8/FMKfIwzv7w
GxE4Gi31lEwkadEFhh0trTjGmGVKLL8BcSc5PZOy7arcGjTBm2jSCs5pSYUPkkFT8vMiQYFUzk7L
FSZsg5Uac3P5xeAlCkbKeBJNFmkNvsjMxB7ofUfs41CDea56D1Od9ukGu/0aTzGDrfh+7WeCCHZu
8lYjV5UcC8CtdLWFckrwMozLZhfb8NRXYXRXmJNif61iAcQrXKeqNZONEofSyjef7MQKkPX1uZU4
UlGNH/Z7mmLrky+KwJXKUpeWK6vblhBJreMt9i9RjkfbnNlJNlWA+wb1M3YLb86iYgcqX8r0AIeb
MG41zGKSpM6Vj3uI4KvTo2pCtuCycvhBc6iwAjWQaZ+iEOkMl4pw5ZSpvy/vL7npiLZhZeDF9esn
JXRPiLB1ZRAd1LVWBw/5V7hc2U05LqhdLnN4H7ViZjbQTAjYNA1EWBAiQFhDkec3hEb0fr1fhwMd
JVCw9lVRvWHkknhfAgcZo9PtLcr4IjGiYNZPV1Tc369s0biE87+WaYTztFkBrnS823ACycwLwl0z
H3S/Gfjv4RW7QMj2uOkX8tyY0JZr92VLtO4q9rL9T3KZUea0zS7PD7sUBiKbJbKSgL8PcdWn3/33
agmd9cCiLIvirbcvFFdiv9s5P8a69Tw15vk/AV3bzgTmEICti6uR9zrcAWoyi1uCCltUPBBPV9Ki
wmwaUd0nKK88fh9HnaYRkWLMhRG11Us0DB4V7u49kxf9izEMZfpcD5Ph0wmGjJjbgnbC+bNe7URX
0Ze3Vwal30S7iRMgRzGTfLJuncZFStDFjdJxL04MC5k5C6YJ3jUnlnHFmf7lC6aRxzcnTB2mAbqk
tV5HY33h5rIT6oaQMizdFx8TuqlxSabmFOfm52ml7a5ouc5I9P7HllcVUxCw1aglQ/xwZXFAv1xf
xJO4EmNOe7yH0nL/v8wA40CJKPDspSwqabC31gpi4xlS+TcwnasPOBXURgH6uqAI6Chpvx/gI7Mz
I7mhNl/v3vw22hKissb6qriZUHWxDwGzQdiRUTfcWZ9d2DwSZ0Qiixt4wS4QqcRgzTz90M9zh2sE
oyQY2xcXYJsw5DXqjrvpPDHIc0S4g9a49yDrZkMET1irAGEL6bFK9KlmbrryCnnCkYGFxvKBTL+4
aOTBNKO3RmVmuFhcMC6CuCAaB37cPouJ3XfTLtiyxJREmwXkUjR5pMPLz+6eaH4bX7dP3DLxo2an
vEebfyGObQ8ZXbJ++rhXg+P9wvGI4YvFIMOeW1ANsN6ulfcN6QQIybx7SqAOab39GP65iSN+9lWT
iILcs1j4LeDoDZTiKN2qamBydXjEL9eS+YWniNDYHSOzR0H8GYJg7z9tRZI9hgMCDL0Jn4kpDtak
TU+b5/GeGf8qrgs8NA/qhQ3kbM4UoFJslWimmqXJ5fUHT+ielOMgpht+S4PJRfQE6qTOlRuT/2lM
ntnLDaox0Y05/Cl0e0cs69kKuFTd9c/4MGLKrYt03Yj8UvrxxiS30H4Iee0jv1cSsyhPFDQIaK9a
qvVQCKzwuc9ackV/5G0bZYIkovWaa4wzbKs89TjAPFeoy/sJwAy8XN/WFPGkCtgYw7Z+vMgBqoyI
VjQISQG+wkXb4eDq+Lj4eGsHO5/Rv+RVzI96p23Vn1BTRzz+AW3Ccf4zeuCubdcnKZ8XOKxO9N/k
r33DV6nhyWmaXCsG9BIaq4GmR3JThCeVdl0rRcakIHs/j3MJFdOxECX37IBlejNdb5F6czKOhu39
rRUqkvgySTMmDYzwEjW0+oraY0q2su8vADvK9gaJ2q1AATO8PZ5a5lIyaBHYwca0w9pbAGtEtCt5
bLtokMjk1kUT6G0q/XOJjIDYb6PWmLeQrtQ3sRK4wpD0laH0NfeP6AElaw6N0EF1mwZZbAZKMeFb
TCKkYO7WhEPZj+O0aBYj1I1GRZS8nviD6bDVrIDDP/+63hUyTFxNPD9tfzZQQnICGxvJ7avloxLx
ugAwbg0Trp9t1k28kFm1jxLgewFpmHYKNgdt8E0h17bbOKbhdXCT+t9GOvCwIF7lA96U717Hrpk7
d3lGi+Tl+YndZj4wYl6+FxMSdWskyV9dZRO+q5ofCAv293l9nC7xywUNrAsTgSTfL5zhJ9F69eFY
1PYrwZ505y624W6YB0rhOgR9qrjRCyDsNmq8s47FVkgKj+TSUzOONdKJVFbNfh8vqOhomuBrofiv
Jj74Ov4v+pwMeWbLX3sfVSeA4JK1jbdXEQwXTrhIitsEQkgQagRU6322Scul3mfpoD9gzNeyHD3O
+xvx/PWXV4amM5O4KeCVp0yqBisuSWdIIgF1YqRAuowWxgOnVof8hOzK4kgfeLswQ1wr0fYyQFgd
MXP2ckWeUwLRGhryqNxr1C2ewT/ZEptivkS2bxwMaIwgxHjMybw4dMdkSvO5y2Hwu26uVyoIfx3p
4Vc1NzKDQsbH1zMhC+IIlaPVDfsN1q5fg60Ti2ZxxKNT1aHhU4gPsqtsjGqNvxEBkuOmo4PAQ8aN
yAvLtl5y4M8XgdrmBU8pN4xb07h5qIOHVLY9N7i1sXmwYtp3Sdp7QZECVZOnIXihZ94R789thGVk
oSQ+jswY98kjUaPt7Htgskirx/g+L6EDI0hAIlRRS9U8aczsMfu66A/nYStHLgNUtnCDEQ46M7Wg
ItmOFfjQZQp/QvI9dbqS7CQcFXJDhSRKt5+0JaDLw/wlTRfyLhQi1kbssUDYmbzvcs6b9VnbM15k
CSo4WAIMAHQ/sFEbVNInzP0SqshKThDqFjk+tJ8OnCIklev7xaPsujqIguc34RcthMDo+JgJTMw1
DRJC9ET2DFd1vbNyrfM7J2WBGNbWoxc8T4VuLkDk6c3XtvOUYVRlnAmgMjclmNs/Zo9rRrTm1FgM
WcdmOwy17QdoG1wcQNuYu+eIE0m8n0J8ti0BXpsvQghc8GUlV8HaqAvZUwp6ZYL7W1qcrdSSu2VF
Z7eIJ82CPtLNDAg5pnvrtPAmBj0+gPbMwo3vG+p4AUveylWpJE7cgVGc6ov/qsYR663ticbl3qWC
RsWsArZadYYBCPoSGl6a5IKyAfoCRe16jfpqJPIz99Bhbyw5Giqrp0adTW6G0EmyaXN84Y13/Y35
7q+xFl8s8ui7JV+lKogwa3OH2p3puCRXs3nvdubSfcv+dSkQFFpHL+2hwEztx+leJjKzms99z77R
I0lS5Y/EupycGqUKIqhgjKTOyF0wQBARmOVe8lPUyk1nGqORV7/yrnRKzBva+R7XmOL6/NycUYXk
PDZwwU7vp8lUImhIR+EQQYM+yhyAab+L0NPoDu3Lfub1rcv3xwzRR5VZtYSLiHNFZvR81p6T5+QY
m1SbeqehY4fbz/cNzhqc24U5EovkPypdi0XRDQvvKqcKcy4Maz+OsGdIDCC3YaAmogt3Nxh3ccsR
WaQ912iHHDQf6PKzoWd+qiwWYRN/QqfrzD1VWpZ6lriJqdqIuejn8BWLwrrPstUBfsKEjJauESvc
rb3TT07BgQKK20p6qL3ms1S+xfuWntB+X7AeAgJQ6v001pg7x8I/UVGlgepucnHpT1/w+jbUEvuA
Xy0gTQuvps4iPL+58F5erm0eeUoC9zMMWni/CM3Fmxh+KA7r3xXYYZ8/uADX4jrxEkTWWosi5MFm
sZoh1eiTUzg61bR3h4shTeQxIDQOY9HK6iZZodAKz0xCvmD2yp1YEaSEkLrwGAsHHR6ehRbW/CTO
DhhlpLfwwIgzIsUp9CRYtkeTdcLAY8YdgUTHWm70mTMcS3iJ0Sl8ui7suadgFiZ994sspvIl+tM8
T4qiESJXWEhMJoFY3yLxh9+BlbGGuDaCdjMDMhqF1swCUY0L3O79AjpB5snm3gQssdx3IbWo+dWY
Im5TAelm1YBAqcuTqokTn6dOagkQXC7dc28rRE90AogjzeHDAKcDYWlnnL6j7g2NZZvIbvPT6rMm
BJW+ev+szLoDjHjKKMbDUL/sFXK0IQJaRFt2MkYShubn3SvKUqxWeX0leKTMp6xfuwoPoWCJMZ6H
j7DRqk+c0Yh2Z4bZj4v2vSmJI8kx7KztqXs/uyuW2AiCBYbwf54CoraRO6jAVBjI2V3TTFsO/2he
cZWbRvG24mWPX8wwMTlCkeVrEuoGnD7Kas+z6p+8yWv8bdjIfzoRWFY2t99zgO/hlDSzj4y5RsvB
6wL4k+EF7IRjD1DzSFN8ANyccn14zqV/LuFoJBEgOIinILKfmO82j50HkSjM3nSCnIOzZmgSak3v
8q6e54pNk3pPqQ385pBbhaQJ+WCoVDG75aqqsc3BMtfO6Jdo2M51AVTimP9n6oOGAwAo1NyPL6ja
vLbYtbdy5EG4DqZLh8ts2nARhMo6yRsxS2HbXp4Y9zBpXHeqgzHW6LWqtw670gXGEkZiyLV0rzPT
msIf43dKzdrwIv+34GtxY1kA7J8ZsjXb4v6K/6hKWUozeoAQ/KGnT0Php4vB70z9vEWiZ3wGnWBt
hoYnvn3SfRicz+gkPj3JtmGs6V9LGCHrL5hxBAPUISXuct6s+YUtKGMi5QgvbddR70k+l02KpG4d
xGSDXCRYl4FuzTGaJI3uznDERehRwWiDL9hDJ0V5WHYyX6eJd35hBC23bbD9gqsPFMwE1N4KZaOK
XzRsdj1lZJkO9jIggroB5LCTf2NsAET0Cit9TFZqNa0uO5BwXH/YZzbLKpNkq//M8Fn2TVkpK41s
FdqZWq4KPG4ulayZcLRktETj0JZQraaEGS0rTRbXB/frmn7j7/4iWhHV0RiS8wzjYGAwbKkU+T+N
/WqZbLldRH4kv/wKNuVLuo7rjyOKy5JRVDhXaPH1/jPUZ2AUEt1ZsJ/zlH3XAA2Xg9Wmf0lPORpg
YgCvwU7/aS4x4xLKei5cU3SpKGSaqLd5u5rygRIPzB4RJUMMVBGxfESzJ4Ueb4InHb1L7kp8lNMR
ZgsHTm0nQJWhVALrJksCGYGjKr6UusvBSLyYR23gwi5sXgZrqdXGIgXqEOh5gDqLYk0k45urY/S3
r8w7MjYkzsMxaT8Dz175C+NyUxYnp1duCLxvglcjG3XFOEOAuveMFqGVTz7T5iddupP67CQeCI3f
SzykM36o5RO6WNuEpS/A7tY5B5WcbQbSyVfj2U8MsTyZNHoMcIe4B+vCpHRrNiO/zwD6/PXcXnDO
nElnBXJRVPExyyPk6cgJHRV3fE9cyEmtjFPBJNqeizqghPJB945o/HHFm7HziRZ88gLJxIsJ9aET
XwNGzZWZEcb1I1o/lzINfb7t4Sh34AUpgB5l3/bitWCCbzjiuUB96aVtHTXTaFudZZdYqan7dav7
fkzV0iy8s4+Gi7sJ2BPavcNu1Swk31UMQqrnHDAeEYQJk65DImWdbAWMRSKvy7Xrlyz1uFbLGppq
b6cTxsDETBNBfOQR3y4nN9NhLusS3nfp2rUIa3VQUDKA8/ijzbx9BIUZHteZ5Lqsr/wiMDhIGzXe
pG3S+wpSwH3DcBQL/deUax7KRW5rl+CXusRqt1ERIuBLFPpEXGYIIjQsQUhah8Qltt7IiHOsEgtp
g64R+SHsl+bS+KjIU92SVk0t+PGe3Skf/7LdgJSlgzBL/uAg8wATawmnjJXJRpvjI7xSc4jTnP37
AFOjJ/4KMUU1ahrsjRsPESa0MRzPsTLvGs6MOYuvaikwViB6HC9/NrZ8w1WOi3YpyD5wL2WFXUpb
xC5ciSc4k0u8wCT75lqDRRI5DBjxEkuTBLfe6Zv72KmT3PF7IVnSQ/Sh999kWvMHjVOZA8T5uNJ+
cR2nKYWUF23xxJ/xTNtf5LERuKg2NKJIFxSvBePmmC/PAAOqxfeLhzmfVDiJCL20pMJuwmhHe5bW
VtOLgDWBNUUNa1zpU4HarCyunvFOhh9o60Ps7b8SwndporqI9Z8okS2SeIrEnBqjdpOU+WukGSR/
jaOx/RcmijVKs0RShCdHxhmiJ5CHYEW07GJd31mF3rae99XPA1eb3zRbcv1W68W4fglDiasY2vuh
6Z6Jq3gcMSLkjF1eu//KeD4zI7dsZdvO4UV7RCVBEofRm8vVIzb9q63Eiz538LjRwPMS6GQDunn/
XN7yfV+FQ21z3Hico6tw4BqOlQf2CQDeTCqFZbMk9oJgNQ0rtlz3XmuYI3yjlqWYYengpuAFnWQC
6t8jLagiZEINUYbxe/jUMG9/eTf3Dqzdp5TADEmFMHG6Vh2izOrDFZY7Gbrp1nCjIJFh24+f56GY
hAP84EF0UKZWXFMxlEV0myoSGb7HXAqsIWKVvez0Fx7xQNQn6T5dMysCwM5jyQ5JLA5GfapdVo4Y
qah8zyZY1J8gouBWtkgncFu3DNuDXi6k0Kja7oQ4wwAoaxyoCr5puVUf5tp0DSMs8mJSeFGD583X
VAiwR6bmJxp5FOVUR8Oakp92ouveq6abI/6HFbG3E9rBnnjba+BHdy6bhAuC4HMJMvNEx4OTwBH5
s6UDs8XBGu/Y4XETbpcEN+Zw7lYxhO38JKmjcdm/u20n6+1SiN6aav/MCNtzpeHQCFidhhTXoXEg
bzJqPR6VqN3g4AXJ0EGMypDSElbyJMiP/BBJT9O2YJnnua75DYgMKjC84wOy+yzoYGGtXbcTOhud
zlrWYW/Kb9k6eHxgIlLL3CWySr8n6f1m7DfnZeR/8jjK5CBH5kBvw11E8aVz6t8+UHgvngKL3q2Z
D72Qish2lBoiwahsrZ8y5Hjo70SD3AkHqqtp+Jsld+TTuN+2TIbgI9fwQnV60OHdWdyHm72PW/v3
eYFLAauGzvUY3/rFeiGuXs76UC5N1l5bIIew6rrPzX4qE1JwMuw3hBMbWRL5qw93SWz1xxXuOCGp
k3PX4Go6AEPvFMePo/hut6IkqLNr0i+WA08qDWHZDnSxtmmVZHyezDdTMRj5x8gDS1YoiNi5saTu
sRapTjJOU6uJoBajZ5cmXDxLMTKjDcNxwP1etUYYYEcwb9hlEE/bqRNu93LKGHzNKw/0tkaDu2FP
k2bTunpNmEXS0NJO+rLhLhqTD5mltGleA11eHylh8Jkg0JTTms9OtTloje16T3L2/NEYvtlIkfnI
OmJDhD2EF6SMMoErF4498+d2sMBMqY0N1B9vExV/GFdXZ0bN3FWdjYtI5fAR/E9GvWRl1A6qbjDc
csI6BCCr0c9pdVIr2xg6xOGiEHG/+IgWN+DsibviB+e1V6GA2nanGYtxFEH6IDY1mK300TgChQcu
hCv5aDOAOAHu8/zaDQh6jKpluyhzvsi0cxuOc0aLi2f4s6bleHfovfycEpLk7uBpcEdf2OMHzBbP
/btfo3x1Nf2f3IP5H9Pc8+3aRmADhdMgFkZRj77JUSojDsLkC/qmQ06iIsiTepdKOBKsl5H3j+lk
QBh7M15HcX4LYd7jr6JT8aPQKfFWkCtZhu91sZJbCfJa0LUJEmbk/q2zxhDOr8ZFGVqNeE71g32X
/W9f2xtCLy+wxs+3L56QrM+9vy7OIE23G4LN705QgHYtJPaHfOK/+vc9WvZThjN8OtTnejSQNINm
oEAmM930hOJMczPeAyMdkfB4GYb4RbKxZL/U7pKKppyztrGOCyFylQu8MwaNvtezPa1I9fVM/wy1
R5ca79+oXOhw2xlmfKviH6eCZ6icWoueuugYIYb9XhCe1LqHYWIB9v/CDa8Gqmz723WdROYFMYWY
LBZJX2skXr//jWG/z9zrVSXyTYEId6Id/etrnuXGDikotmU7O/2vAaH/S7mFAbVad2j2zPBUINkO
DP1KelE4HUJZqb7MyQYB4oiu91XRpip9LRs4c+w6B3DckMJM8L3PoZf/76HSpQpger/dnYJu8mtm
GUs0xIZZ2g7kYtTE2njeRnaK5lDDBsc5mJdQrkol2/QePqH3P2bXsScu0kmbsJn1F2wAt66jHo2k
4ATH3jq5gBe0BSjuSupeEwYxiPfAbMVo5GElQwbWZ7/7Vj7ed3niRvZ1xcf/UqR1mhhmJyHbqGzN
3hdOOx7yM1J9GMvROvnibvmLqU7h6uZZyfM29q4X3qUXlubBd8IDRByoqMRpJxaHA7vbPU2qdVxU
tCZtNRDhpJPFNlipaIGLHI+oQXxPNNpQjRFYoZtcLkYsN31Rl1HA1czS6f3L34S2ZSmVqryW2IUo
0n7a8Q8PUaK/YLlO1Y8oQ6F1JY3p/PN6fpNLPRoX2fFVFKReDPdsNxYdr8nUkMQgE5VrtiqUIsmH
Q2SgxPgXXhRocG9iOTWwZOgKywzCJ5oNL99Z+79t1WFwAkIMHGEuS5G46Ojd7UeKF0T0NlqxaRQp
fgQ0Ywflj5eXCBrlybyVJoRmR57F9ydvZqjSRA2luSs6R8uQqfvlZnOLAp6bu9O1hFAN8Gbcok9/
DJ0lKmPYQPcqdupgOpiTBRaGjQdAS3cSJO3ExOpHw8HkdfhUIeqYoPpftBYi7NtaQfEu2jLMDPYY
h6M69UbChWB1PLSWHRcUFZP6B3YQ6NQRjuQqbJY8sgxhwGeinqWVog1f+lcjkpMu2m+zOgiRNzgv
yv+1KQnlXXCtQXs0NmHGSRmFoAcExTn++4vOeQLZMZysavYZH7xeZqhduTzxIIIglElIUrOqzB7e
8otfo+KpppSSLaONcdS1j6Ggx5gaE1+FrHSEHvN0VEvoBSgJCloI+K5ubgRhUlnL9seTOmOjYk6K
fzUNNpD4X/HZADG78LPRngq8QRkTGSFCv1JA9AsH7D6f0suITNmdDNmG8Cf7UfwM+nNmStOcHtLT
KcJ50F/iCiMrfZoKVyHEIlt0608IjHOUdD30Y4mIZ0P0qy4Lo0YuBvmk8M+/cqeEc43LJbnKJxI1
yn98xcC5ey0YdL97wFGSIy0YIPWyVSa0erweqv9i6ZUqBIe6AkhqI8jveJsVlVD1ozFVaIk0Az6+
KawB/JcovDl2NhrvTGbnU0CXkeLWYZGZcacqtfUcDnRcwglXa6+bi92PFiXP+mTgPw8Miq4wQbrj
vc0gj69ojxN8Vtny6bLhSwaL8TxI2MA/1lOFr4XntSicCbhQ2uKDUJoAEsFnrNMEKlJyVxQ88R8m
CVItnqsUDKXyVaPzvq0ezash3BvqODUc4GlLIvicu79Tmm9wMhRyGCjHhBAG6JhwFrTTicS6uLY/
NYWzcC9vvlNs2q3I7N/QEG2c1zQ4gLWfrh09Ufrj9HgPlY2MXGIL3H0xzgcng0TZjMUsfWfXaWmO
D9tHNldcb259PZlI7jc/AiapHiz2gA93vQNAt9bxvjNA/ZVONJ5QdRyM0E+1zYwrZ8ZuyX6WjGzn
0PZRXoOYeyFA8+NiNGVUC3tWKd/8BAUCmY7l7FImR0l2hFHscMYcYPI/myMNeCIL9mqVLPXXrwGo
OiLMzOh0xhb5o6vmo1hAFX9S+aZUIKKRoqF6KZWNFjXS2gCm1rvSnZ4nvQshl8S+ENNGPV95atF0
P2mJiUuZjFYrE5wBy1jiwwBffrxt0ZvTunRScMCURsMI/vjPwdj95oAnPajOS79jIFivB0ZjWdiG
flnT6anf8CAqX0gYb6Oxv19ldH6Nz7nnNid1Wq+UhsL08a1re2AdHVHy7FrO5G2v4qyDxijTX3LM
q8DxkF2atspNT/xIWrJcRQj7k1jiW/iAiB3zRPVN1GbhBaPTKSNrlEhXoTpdSZfCv/NGyd+LlLnq
1vWgd52i3bSk+/t4TGvmb1+xfhkr/RgEK/r9o/pauv06khEu5Is2PWfGllgNBGgvUugajUXYl0QT
kXAtXZrlWQN384TwVPWryN4cf28OJYhpXdwc39mGP4lmP4tIInfE6XfPPwp6yCNjc8olWZ5jZBeu
s8u7Q/6P6m9SvXfIEgbO7B+66N7Ew1yJT/O4hUu+t8ivxB8553ApY56fpLUD2HdIbIyEN1WLQAwq
Djd0AHTWsvK2cdpt+GzznlAjKv5KqbdYPPLAa59Y+w2Ffh6KF9ZA8nUq9xniyacB7yjxnM+pJKGF
E8LzQMWMI0ysmejE0k39Sh0j7p/FYP/b8FsUdeSW6R90hHPY0GXFUBhQfQNqjlXNd+A+kqJWOUrk
ttPA9qWS9Jp8BmNR0DxhcXEgSUJ1a/yc4bGUytSjLGeO7HXLSE+TAGHtgwGq2aKMqKjTuzlb8Hmm
ovX3idVg5Fq1hqeXYDA3EUsIE27QOXdtdi4rjjzoU6sWAIUo3D25sWnEzZBhaDJVBDCV2Jv9gGtY
cmdvlJ0YURmZRDOHXLJB8aIUQw1ljWDYzNuJctQNxpUEw2INLYH7frdqoJL/wU+ynagtBN3QlKYN
Pfsby8jOTJxhlTqeBVik/159upXxts2w3Zmz68j3z5qsORphhnNVyXRVipmKCsh9tD/1FaR4aLiX
wvmaGdvPjmIfYwTp3JWs21dP0EhzFQE82HudG5Z5eqeGsBgXXfMfCPx7OB3i5SN8bFANeZdqbfTM
xKkqZLhxwEk/xp75/k5NqcbUqNImRblMZ8oE0I6v3lDCd7kaoZCS6LMWY8ZD1ZqL4TAxC72nxfYB
tjK4oDjuQRz4oyB6YnqRvlObeu+/4NFD1PhCKr88jnt939DGF+HEXnrv0EAw0TEjkbPOexVMrZT0
YaBRqZgmrFAs5g/tQ3DMydI8bw+RSzw8HuuYNF/hLEBIYQ+5vbcLx4gaRlY8i5eAbZ+K+VOZbz21
GQOcNrJy2SCY2kxJ5O/Tvpd8yORDvbmIFt4Yqm9Ace6f10Tq4zfWtBCwjmBz/XH4Rug7hBmspbaU
10LkYirIK27+8Ma/iIEf5W+GLFNMFGOrqYV6AHC6oYJKfB3zuJ3/R7J8NQJ4jg0bqVz+aKzyY47p
oI4pQdGAqh7pxBo0FFzMtp3Ra9WJ9QqJzMpyTewkVoj2S1/zZQxONNCpL6wVKIR5u5/pMfHEwwTQ
Hs1Y6Uq6snVJIt3AGOK0klUsCv3c4rOY+tfQF9ANiyYbQeuRoPoxD2XWtd6juxc9XVfhHG40IAbm
m4d6SvlQDfa76cHgvWfDSL3Tq+wlJQ42/8GXFGEoUIHzRJd+B+PdE2riAALQapxL7iJTnT2RGePM
7yvujuX6zrJG8CoNJGFCs6YQeaPV4veTtAZAl3Pj3iZINZVYUOi8HXnMazpafm+mkMsmztirnUJY
ZT9uL08yCXfQts4cHnij2S3pGjQ5wAkuDXiynPNqYC3UGG6glbk+pEjdBcdAbZicnCAZux97g/+X
Bn7pA4pESoEzaEd1eyNR8Ve9b0n6bymACZyv8j4qJQvFHdhtx8D9bW1slX6wGl2CO6GeSz54K6XL
xFk7O+bnqIMRoh5AUzcaOwa9xeY0UFv5wP3MAZdUPsSGkn/GFU6qEJIJeZnIDBSJefD82mmhE5C7
EzJWdON8uQUcqfzzoPtddjQacj8O43FIq27tjXdKWlcxaMJZPl5TMSPr8IulqureglSJiYuyMjJH
BPmQhnQK5Uw3JASJ04JaBI2lNlak/5nPrJQFwgLEuoewYfBN19p6O8XHURF3KPUA9AQcK0zrwJiu
wYaT0sIZfvP4kJfnlT8xXoBgOmFseezzJ/RSGEyNGLygpac82Li6BFRUGIXHh8IqgPDJBkw0cm/o
YfywVt/ohHeaUL91cl1niKcKQ/3dGfeGeINDftVNyH8qNHt7hOtPHNRGIZbz9wF39C8cc4NiqWS5
1kUxzNXdfmUFecV21AOPp72ljaUs8yghITp/dwcSmvpXJ3t1lDQt8vPSDfBcVtV+ZmmKEJLBJLUC
b2vWAVqwMIWcUUQtnua54NoYr0ortGZDauXs4a2FE33l92YYtRvm2xrSTFxZm3vfcK4/t+3ICdcD
PSN2PIRutKdBvOk1Ln8EAm7lDKb3iC1ONUj2cjI2bczXeZeHiPUPjygVbgnWaT0XuN6e6Ko/luBF
5c6+dGLqvxu2ES3Qn46t4IFZaZWHytYgrs00x6a7HJIhdXpfOjOE2+rEmSjtmlY3KI+UX1Ya2S4a
749PkobN+mkoKIMdLC8EK93DgzpH2IFPQ+B8VeoQwycbL341k+RWao4PQ7IiqQPuTJoGRwZyuLgb
zmsOP23Gdbo0uaSejD8XjHjpWCiM1O+ARRbGWA3jDFyuRwLSBfsSoBNsLXCXkyv+c3bfWN9wiPvN
KUQCeDSyPhJEkBRN79kptFtzot4m2uV1L0bmVfHM0WT8NQtcYxC+AmmCHi5TeQfTtzKmeR58TSmv
bL7V8FOR/+By0AIIqWgXWg8+Jy0a14dLe+dT5dK0tFZvQrPoSlTwg82SWMJFnRxAokgUnUTE9YZj
tNVzcyYxrfv9Lye+MUi0RnJ78uvtDnGnGkbO7pbLE4O6s3iBwe7SY6SLssqhPIzDlP8bGZ6MWAyO
kjjnzP1BfyS1OfjVHS6GnLT1nnjr23QyvGi63JOv/Xt4wrcxJS2GdI9iGt8ntWBJ0BeBMglTFXlm
lhX/G+NAGZ/v+e61j0lNo9q0NRGWdVDR4WAeltFSjTwtaRiYMeDHelMzGOOq2eOgJq6FkyphKYVZ
YPIzZZ4sbUxNfkl5J/JJa6XtSJqfvX3Hyi1NSoiDJ3Mvq9HDi+2wsBWZ0puhFLLFojvIejmJ6cKy
bEAJN7RPKBPJWoq3m2fCHm8/qR8gxO/FOk+m2bdLgXezXA431ABiYGvwY9Yf023L0u+4EJK0F7b6
WTvjP/L8raUq0kHdp8m6Gvw3I0YVyNzXHpXnuhKgTCxgWswFy6pNR03s5EVNVE9w9VivYY4fZz8V
ijuruFkvTZgFp0ZGfIHkFxzn3kS9ehDLaeecMyiB044ZW49GMPJKaf1MdDP6l1AG2W4GqTuQEMUn
/rNMd9E7T2wKCh5ZjqfgkF8d5VJzekeiZBC8b1eAX3wYHaD9yzhJ7kmsqfk3WpOTBoHTQF8Gmtpf
Nnd16UyQ3c0H4I8H+MJdKYVomJ4I2Zk9TrBKywkL3w2Zp1bV89376sIO1LZkJJS3hgaNJaZgHt0b
c7rm5oD0JP5MFkgP5uUi2nMDSdYwz4VXPHmC1tlC8mvazdCY7aaadDsEqsc6Gb1lxFeDEKz9pWYd
mGEf1gdhaE1ac1n1BYw6Mb/CTzYAT9D9oIY7FCdowrObpHHo/yBUGWjPiJ11POlTrnFIeQc5QraK
QJJg6S32zzSXgDqQOKdLmICe/ZKCv7ClxJ3BFPmOJmB0JST0hVgp7YottYzR8gvx52nhuHV62+CW
fFs6yCoI27+7Hr7Ce/whjya7DPm71JENHBJs3NpQWG+r8GXGkfpgMirISkfBlawi0M0gxXx+xz61
YcO3tzOMxmFyT3WHIRePhDyrlYRW8TcBd1upTqY58vgUoJpjZkf1YbXQWbYHm36ifutyAXsji/Q9
/O9Sc8cdMNgEOA+4qC7aoDUYzLv25H4irJUlfc96L+n2zuIbUdIvrYyEv/Q092wkWf8DmXlAiC/r
MGOT1wdiF2ksvi4AOdTUaLpEmqTT8XK93PZGQYURWtAAkg8unjJGdbU0Re8IJXfq0qx9s/HYth2w
QEUAErsgk6bFXj/mGuIYsBfRsdn71ZfExvZwkU56j+viSI0xjXBQEOXiOPJcCfSBYwrE6LMP6/WK
IrwdW72h8dkbN/6cG3yyFaOw9hN3LYBo9aJ9bWpuZy/apmWlinJTX2RI+OH2byPEcP389+ImPqxX
rwSaG8fFgdfPYxM+6fj5dGEFvQevrsymLUCgGzsBSCTJCTM/AEXcvGIm4dkhVQZB78lQuES93klK
+fIp2LKNmRNJuFgNTYb5PiLM7P2VKlUS8V0Sqb84Zdf+FoTCBLfD/z/hMYQe7lnwysBNNiZ09g8b
KTEpCa1wv9MEDq6uy4q6ye1NgS0rqC/+zt71k4bw9aCHi1okZITRO55Pd6+V54vP3P+12puarY+v
AMCsr2PtCCbd7XX8B/Pbj6C+QApynqLiQQqA5clqbHVmyIXp9FoMe6jeXn4tlr7OgdMDXVsv+fpw
nOn+gZ8GPBkekBvdMwX6w0Ziqj73o+aaS47iG60I3D0uAHcd/HN4fKUYqHw8CFqLNF0gAHXPAjXp
DfErXq+JJ9D1OEzzP4BOGRWKwY28D8keYSwoVHDk/QvjwUczY5/G/kt/aSndfLlXTjLAQTKtEF6b
NhivZpeYreeCSigisE281rAHLDqdhlMAd+ffjPD41u1XAaHZVjEJlh6xZu6JbRm5/k0znuAGNxR1
EFEoEvi61GmAeyh45/qRNFi4oguO2a73eO6ZBAwBlx7R3UhSfyFNbnTjEETsoS4xTvvZVAgKIRNQ
h20ejt9XAwPBaHW1RU9A/43+xhevffrypVsTqlX36DBIrRpVxMkjY7O8KDBv41Jf4aPLTreck9i4
5WoG7HWgnhKKrg+a5ps7UxBGWzOMTYIRcsCP/YB8Ujlli0XwKWpi0ZMI8DYatULGpIvG/poTdFIq
7MlhjrQdAz8UokiQ2w5jxGuzyj3djkIeEu68Dxqf01V3xtfychVYaZU2qLaHCq/y0m+6QqtWUMME
65wxjRd4XcHUUoqfy/jBwuzLvvP7nz0p3R5uyhUxTuIpK/Hrzli7+VElJm65IV4RuOHiB/mcGvF0
SQlKgP93x+IqvSf9JinB/aPOq1V9shWQ5qqYS4+lspPVEXJzpSNJE/AS2hz+zoGT1jGJsThu8jbe
uaDBpeFfGgzMwQpZ5/7/anFdXR0UacsFb1In2C7m8niW32NQeCDhsizcc0jkh1Vvm2hgOx28ToLW
h1/sllbZRWbNase5hiOis/u3SpEhWmVXx49IID4JncHNVwaON6HH2isTWSLWGnPO6LU9oVlzNwnN
c8wRLRe5rqIbd6XeqWqt0KWgOkzc5FHWm+Y6Attucp2aEyzwzFTSKlcpzUaFo1PlqCs8qEH7AxMa
Mc2co2jno6dX6zwupOPqOAFBA1sM4POBmu8S2ZrxbvMBu0U04p3u4cW9f3klvdK+HJ5Rt2Wd7R6s
Y6hYAwa36fpxGT9rh80oGVOIe38CrgtSS3DiJ7HdiDcGKZ6aFU0lP+wHAiY8lzjpj0nV99wY8y0V
0Gz+tJvWTRGB9UWNlDVsSiBov9Ngz5F5w9TPKEtJW4qcz78FW4aS8XXuSoTFmWdvU6fE2jbH/i8c
V8JuroIfLJd+qrlQy5muxLgOqiJxo0J8THBFAi0ZlDIoxXaStYrRwaNiBCXrLJBYsoWyS3dBP5g9
3KLiGBCN0UkTuhA55Gs5zEa7q+68xFO58sLg1Z5DZ2XQAtfXcredgW94kDYbIp6oPso8vKCPclCr
D/Hi2xi+sRqhfkUzK8FTkgPE8rYV+8CLM1emZdZpwH0d3/U2Wd/jWxiy/x0n9i/cBCB+et3iVurw
yMD0AOLtGkk+twe9bnazp5ZZYd1y3bCXlFcCTT+3p9zcaF7KM9sxSfZwFr77I7jz3dKTvuZ/TOVr
v6tSYSdv9LJHHXtsQmy3lbFB7CpUFHI2yiwNP2EPVGzxEf/BnXEYDy47X6MF0bq78nta0/Cw9ItX
DgzOj+WpiX8VnuSWvMGJZbxU2fw8/GFdQIm1TnGoun8+PFp1KJXoxBtdBxa6yAO5JUT5oFejQHiq
9TvVSYgDt6ii2DotXscJ49MNRh5mGeh/j99Qs46vrDhinwLcdJ9U/IrSzPpZyaGp0XxTSs2d8P0u
GP1E8sVadPSMqeCS96F2ZmWKxd8ZpEmv4CV23N1cLSVjwknqRPI6JyEzdh5GKlZWxGPjKD1dXw6Y
L8ca2CNDHZDp//6IAOPDLWCw4nDhi02RSDqzbfywNL69hlCMp+moUR/lfNHRP7ENvbjtio7kw8bG
k0qelha9CQHkXICIo7s3f/T8haMuRKSgtVVZhCjYdV8sjjVerUadXohebpiDKyVh8PQNx75z1M//
V4ZjO+rpWEmN3w3qz/ZFPcKA5o+eAfMr3bLJADB5B4dDV79/GoBOIlOUGEcvSz8RqHuAECeVllK7
UWtdMujthTBzgRTYGev0Hkn6KIBduPD+hxPEG2i2G1HLw7vNohypti3cEAe+1UqeV0g9ETQ0gcNo
FqdZ1MX022QVx51msoUZyGjB8gSg4Y7fcxhmRFCJNSyl9s/9oDo59t6b0d1HnujDNBx8da5Bury6
RJ3CqZg48PXWwgQwdFLbasVFydeZRQIrB5lXIkGCkiAT5nsLB0RWK4/zfWHxXSXNhSW4eN1NJPdl
idQZ8DUZt6yDa5eLyRBv75QKewTxz866HNLloy+ucB7SIXZ1jb4nfExOsTWm+EfaRjGnoL6T1J9y
HxNuJI0InSS6obeX4DvVFwGLQ355e09Rr17I7gZwmKk7Fa39H18THljfr20yZ+YXTUZF4UL97osH
GnCuywqZ0U875NUXv/CIvdA2LA9RcPjNqplQTHoRLaWUqr8+SYUAiS6lxCb4ODekd7Lsdltqclk9
o5LPDLmRl/4xU5tSJLhfzZK84aNiIDsUiIkT6u8wOdgcjf6a9dRpuldr1kcLF+/M19aH7zWfoRb9
gRzSROBC5ebGAGjRAqz2AI16ySlTQb8wCoUrvw/Z4yKdiZXTBzQ2T1PrmgBknk+UvqW7jTGtV3jQ
KU/k2BWc1tQZSDo2B3BFUEMSwoG3jda97TlsuY4L34VCXBVMDO5F/oK5GORvV+Fz9ZrwIqXU5IH8
Azb+/fWsfrTGZeAU+FuJU0bUAa+bxqIkGVVS1ZtVm4HXqXvchkXOIJIvf7vITqxc2GLq7+US/WJs
5HVwuTjxvl4pCH49EGvcIZC7mAjq7pXXOf6GnddRE6aT2zYR/r6prjQ1UhhZpAok5W9ZU9gtgN+7
5djWQfETbof3dTe+OXIH1qvSI0umd5zALshsLMia4VbKJ4P6JHR2fJjDeFBgA/Srq1asJmFSz3hN
yQWGSkH7JLBTjwsfr1gv6MN3kbvmSc4qc24XB7nvc9VjeiHSWr0JJrvYbbvk1daHTvUkdiPoT4r0
rEkWv9MqbN+dfK8knGGSSF+Icyn+rxFF+HPT59xO3khsgl+z3iX3kSr6nOPHByXYDwBpm6sxH5Gu
5z0P5MAVo33FsyPup3C8uRlN3jbLvvRsFo7Lax9t1laSf9IcmtF4ErhwJCt2IJxaSPlVIN09OG5W
Py0I15zB6TrJylWyaLVT1sFyIgZHtMRpnu8sMu2LLnBOsVZPH4JFKhVTL8NfdvexVHRA76+gPa3N
jEZ4pwfVNDA9FbA4FIM88PiwxAVoYtFhEqSD7sBVyULZv8C2YTqqDeyiLw5+pDrpJT1+CaRS6r6x
618PY2+UkXNrY04itP3hQtYthdxVRsgTUBpla5LxZAznijAJP+UyHOHel51DEIYbBabAGcY/to4y
yrpWLVzVEry3IzVB399RhndXH3eOBDxsOIpnMML0idFRbaeoMw8TBjqmuAhyNyniYMBEmmG9mYbC
dHh3lYrgf15KFn1B99cqryoLklGBnjh/9LcrJO4G6XVcqXMmj1wkzuSwBq3P2btEodmL2tiKp8sL
1y8gI1xht8F41XN8HkG0qNvKeoJR2AUYDjTlLbErIfG9e7YPld0BV8UgSiXoWBLdyC2hTMSoMD1M
NcaV8dMcaEGDyQIX79RBVZt31h7vVbqHCbNt51ocnzojMRty3bHjIT8RZ1JL+47zdnIey5H3EjsR
kWoGWfwvSxNCQ5xweZvfWSsYWV1MZapQBvfoM2EFut1HsiYZX7Wzl/JREV1WnqBeszEGWNXh+Ctg
4LfOTBu+x1Xjrk8rPzrNv3kgvSl7XykyxpGTAuSqVJZPngbbtuQCek75U6o6twuf7VJsQLPBIaFH
POa/LJLM4fdSHqGQ6hsW/Ss0vEQSELRqF4wNjEYhocfDt9gxqj7IU09w1d/QqcODmkNL75+Uu3FL
5wEK07y2UDjGNaFfsICq1ZpisVcSNFA+Q5nTVO2i4HR7RUWc9di7lEW7TXoHlPTf2w/K41gWIRAu
M8EBeIBi+9vMchbFWH7s3AkCCdDi7vuCxU4376ymfpnnzWAGbT2pK3xC/tRiib7xhRELp4GVuNJj
bOjmi3fBHkQHq9LxKTD9RY/X5q00k0oQjiQzsrC0czr0r2PMd/RRijt5qPk+o9FUTiaFfGOEEY4R
KTLTZETXDuUicMtwNt15+MUHAKFmpUcFpKAew8Md/LRVLegrbSaeACFPwcKO1AQ9YRzD5HKpC0Yp
BoND0sBGUDgdd1Vhi3Wv8U7D9YC8Zivw+/U8v/7gkZjOSYdgVKh9bkX4Az5kqQzFi17SEMk1c3PL
dufwcsRuyB2BtzjuMrKVkcvwxkbPWVgW7oQqo7fwjp/WbYyOikRAv2jhhxUwmHXsfwqm/p9Rt4SK
xmLW9q6gt2imJQPq4EVdOq2ii9k3HVu/BdTYSmh2ksHgmvbBh0GZvNOnJCRyeMYi2BfRUqK+sAq9
dcAIYBDeJAjSvrCnMpt+L3mO0zGsjiHuWMMcZhkieVaYWRbaE7pIxI9jSXpRK1NW5uHIbtdZtCjd
TLIqP4rrA7hsqzLKRtXghaM4i5G9Lg2DczkJX+BE56I6aHWM/iF4Hy6WzbjueClkJG90qrFRwzHu
2CYw/sqDUT6fZDppZxDyd3rJtOjDkUatgrZxWueWYvIuahbVzsqsTBnEAm5VnDMCUjzjDc93QEht
69eght3xLO+mmozdbPfkphNP17NddJQguIud2V38BTwjqJbicC5HGv5i0BOZCkIYiEC0E184pcz7
JDbs+r/jeLXUKrAB0jPWhyqmz9xYXenRKZxQBppG7EujpjcHAn7T4Q2ZTjJ2a7vWVxR/iqHlo4jS
CTvvXgnPCJo4BCe0lKnizsdMIvyxsU5WyBqHwknkCUqYpChspKi3HByXzfj/i/KSmBJKqs5/URWn
UdE8p5E7uEm2WoJQu8b9OJ99iZRxpixy8tAVBQYfwKK0kx1H8YVn/U46ObCMeKpTnUmQcQpAiAjV
bvzJBnKDN2FhAECbIwdP6Mst79eOz7y0f4F72L0g0iYgaEG3k2zyqWUWH1eCjTueiruZVfxzLW+Z
6bjrB6maYrUG9ArvxzukSbG965PCZYHG7bN4G3tyjaTkGGLuNFazvhJWSSX7QhyxlP25JzwSHgls
XhfgTWJkl38hrtCkvZZu9Ej20qR4WXNUQCO66xG8PVOghBSYHUIncCaFX8M+Zw+8SQYp92Ey308g
HFGYyS9RefxZ8IaB5HEuzChfCWy11Fl/glMfeCKGHHNW1GZiNC6267+MFQnjHJ5A1GC4rzs36XWf
W+cScfOZfa0eMDYuiN7Edx8PPr2EyQyKarwfqpyY5TVoF5qj281zaII5Uqp/2a4MnQ8+JqH60gjL
ITmqRLpMoUMGm5MOd5n7hg48DmJORoR14A7QniA8FK6dqiiDdhIx23I/4LLGNGNBFLDhoV0zQFc+
S9dZ9DvL/aHkWUlKzjvTDziwI6Z2qdoyq2zir6Dajgk02cErS9nLTfSdZqreHzGoiqzR6g8IOc2j
3evYbGOE2Ta7jw3qTNNCcjdNs6jrIY6pd2u0q9maO0w13OzxWUX9d18d3KKEB9PzVuBbsKe+l/DY
mGl2fDICKqx1Suyqdgm8WIpkkyI9Z6gBE9DsFg/JUYrZMc0vYSWjjsTDxdS9P4+aioedC34SffAn
0vAOfvLv2BfmAibqmdpJ4cOaVrFsa2cOeu5Q3H9bTckJrphCeqAZl6qC/Dar2K5CGkRWLyYZmUmF
kwCAcX+vVQyZRq7C3/o55B0QZF0PO7E+DefjGyFCalld50rmKcb2sB8aFsLBjcqVlML5Z8WJXa0D
W3k41j7H47eJY56jUZjJOgzozUyNP7oak5YIFFE45EdcIuFsRYjfevabFXw0ktBs3GQUuS3FECN5
GIbqU7oJyhElKoGB9XFsJWLWj2FyfDAKGakJ+nruaBpK+BdTvuJMBnKzcFZxfRLo5canJmNZDN72
ZRIdPvHpS/RegaupoBsBR/N8BDmI7ReX4XgNw4OFj9jt4QSjA0oJfumgeR8MR4BEgXi4neCU3qZe
kEdEHV8/hKcYSEwNS3FvcFG84fUeTJmou6SKnLF/Ilp6jmQJzJEE7H72LBx1eZqPOjBNfL+UM/gG
RwH414yLTgiLw8nxSrRw6cjDRlE6612vH/fr/KIi0s89HdP/qB3B1DysxI1JAkaja7ARXnmucQvJ
yK0zHLa22bW4N/FwBe5fnpZ+JDI82s6/0j1EzeXwukN2T/2EbMrpVy92eqXeOE+fqb8p9crBYCIo
7pxuDKp8+mtmYrZqC/D0jcLgaYqNyq0d02huUYJV6VhIB1sIGkUd3LwDVqkqXylrWb5tXmjCAEbq
tJq0JYCq1k/6z0ICgvIIKQAWzO5+mWTPxxqrI5tdrZpPJqM2onjP2py9EjzKzCS8zIz/VbJu0To0
iGlw6WktBQAkmwjeEoMjzsKXkWxPNdpX7Qtl5r57pHZZ7MOiJXNLT5A1YxhLiwB2S0/LyTmlQlGN
yfSi8vBjdwBIKEmoQzbvMl0oqttwXqX+DOfIjyO/x40DsO9R+JWsAcCY1nVXUVyPZLyTXtGI+DPh
ktLt2rIRpN01JAU6K/w7iqc4uwljww3YAVFT8OioQyRZ8DOt6K3MBNtpFDoWY0SbfPk4yYJF5AE6
YSZIwgEc7VxlN6hmIl2v7unUCvI0RKMugv0aM1RDdG08DPuEF3FTBE2NbqeXUiYaiH90mGywnmFO
8F8FJef+iqgrVrlf5MX4Fu846u8ei3wY/4vKtCRQ4X5RIStnjETeSgrwC6RAVpR+x6ZUpRxvi3RR
Tu5aJDGkqQhDE5F16C68qOanF4ADoQOijinjK4j1KtcTcDYnn91KZwBzYwYcrpuY7pgkm09ZJFOx
JRxx4pFtP7TwMGN6zQSR2p60NNR0VIhRuTVTzvThMGEG8fM6Q6zD1RDJ/abC3bjziQvZAjY7FiCu
Tbwqk2tSslE6bGmyIpX/8++ts3rP25jlTmX2R+7I3cMUp2kg+Ii4qPxDerNoFyTm81TWOpqbeEcm
aw0nXsaPi9rjwJr8RVNqgcXlvNZsb2sESuaabHkd88q/m6hP1upL5D4RezI/g4n0lD89W+Us0tPm
lNgt6NkKdGFf2IRI9IiAFWDjzhV2+6N1kyrbwwWjqoDDwsUeEgO1DcFMDmGNsT7nz9fyYl1xvIX4
S0KSfOoPrW41XE5Add5751JzL5erX028Otes7d6FIYyqE4TM3yAGBc/Js2itZElLozwuMr1zQdEe
yrfic34s86l0cTle0I/fyoVJgVxdxDh+xWLGr/OeTi/GsJDk7cyaMdLPVFuhK+WN0QpAIErOQQjO
u8poBLHYf+j0NR9aFTfbOp5w6JVgmua1B4k9ch7IGZfy3XxwZeWLlio9cjoERhBDXAktMdpq+Bdx
n4pUF4R+8Jy2/57YLAEi/PbN2nmPUj0BXMsS6ldTVj6P3YMvVoDcqDwF6mOMrXnXhDn77kNI8IDK
q3uy+zpQsKXlBljWTLBxH1YfiDqe4PVlryg0tbjExefiMSdfnw9PqM0zLc3bYzw5PTjKCgJti1SH
+ulwsI1d6fENwDl66kKWCIjmYpbLuoGGZEJSAj/tjmLruq+MzB/aHmtlKB15/R+pblTkdm3vnGVs
Zo9yu+wX2c6L6w0BslNNYNlHaJS8H1XbmAlZ7yHENMPRBgn/0rjlvhKQ2HGAG7upZgw9jY9watoP
Zv3Hm63vhxP2no9StGDs+kVS9LRkT4/K0UhUbQNfLzW/w94qmFI9V3hmg3S6U8p4++jdSiy+chAH
JiTk+I8p8bZUPxX9ioGJj5ec9pZaaQ1xtJYRFdtzv+Q8e2cSFg8QC1V+6JWZFSjT9tcDuls1WVyb
quP/inYUN1vRLkJE2wdVBvkG119m0UwSP31Nkvs0seXqJslZ0hBEPKnhJYqDIyvLIB8n+swelOSw
pMBUN1tIshPxgQ6gmhPUw0WYNxO4pW7fpdYoFEiGmTUBvsbx7s6fpsmBUa5RdRrwgynJxhGS3Ibd
ucVtLtFfdxy1yMzf0q572CTUE9OFLmMKQwuQPCP0ixDDzNPK+xkT+q35IHiQanFmhTo4PmBIr9kv
CZwNxqknuN6JOncW6NGwnELzxNyqEr4jfQF8IgnxIogL4VHnQZgPLgvXsDGEGo2a5uEzA7woWOdU
NzWWc0tcBvr9CCC5Z16rfyhpDjoe/LlvkrcHtNipOkEBc42VKf80UZ7YnusuyuVrCEplW3MWXhG/
szH6xzJ7IcGlyihDZD1+JvIT881oCYJTiwOkx3YaFs13Q6uCbQWpk/UVZP4jTpkweqonWTkCgDXt
GAgTG/hqJ5E4NMWJuEeHjnFW8gX1lKwpQ9JDAvzkbQ2c8bxchgI3cGTEU9iPNwiFZBUXjwaH0IiJ
/cKKesVrCyJUBF7WdNmx+eSd9DvD6xuEXycglQipJ0Yyloj2/fG24He14RrJG7YTykBZ0XF5Qy9e
txJ1SBYaqeOQbmdyeTU4FRPazxwG1ODwPRe3S5/eI6cDyMK/ZyaIRlefIJYZV85WlLEato/y5cVV
9g0dIMK4bbiStYUHtcpUKj+Fz9ZuZE83RE71U1TZBIS55UUoSRo1P0tTjWMbTNX+7Bfic+iVlNpj
LO/zcjWwGjMIJ1C+/BVCOehUVKzXw6j1Qs/UtWsCVsmfhFv2ixVGA75nABZ2E3SZladkNh9RS1YN
tgT4Vwa9DdGNmJuEJCSqt+yUbK2pz83C099hBjwhjWlKhw7H/ogMf5xkwlOLf09PWOHmiLkNPNw8
rLmqbv6iZzsm8kKzfqeAcmjjIjubxsakZcDajb/afa/gb0gxz+82VODUdrNM3Cof/F38j83tdqMV
83reTwIv1InJPfyCO5yJA0Quc9NWO6Cen2xpPpdkeAShk3BA5cyzo2ePZ222/lwUY+cqF2+92VhY
3v/RrL3SCdEn9XwmXAnExHx2w9f55Sfii/69ANWaQancthiYSM5WjcmAj8LnuGabIkF+u6iwRpmD
/JQ2pngJJpjvdBPjCD5arUAYNl6qcqx3P7e0EhCvPDBrv47qUJcYDKTwsyb3mJ2XxTBfGwXjEvsU
pocwVqJHQJ5h5BaAJI58nD2DU8v5QPEi3BNX3N18KVn0lzLKNAh9h18WPp9iAelnW/pZQ01aWw2s
VRSqOBaNywgJtcqBajwUEDlrlYD/QMLZlKw8UE8UqrFRqJCNyJeVkUCJnNfcoSS8OdCmHiPdhspd
yph2eWBy69+LPFB0AeZK+vV13I5WIdW2rlb8O14vwJNmcdYh+9r3XIh5Y0Zz09ZE3aw8ZjnDYRxt
/Gg2TXzjcmS3fPw6wYWVGK1lQ8In6mzC6vJqz+wTTbctQzarI0v11ZU03NvRKEg0xD2pn/nVAMH9
I4wr1BHFai8qEmNyyQTaP4rMstTKCwEF+jmCTbezzkvtAikqOSXBN0he31mf7+U5f8nVE1efuM/Y
pFXBy/dSyE/BLD6fgkcon93tswIPj/VPS+IDWQG9w7ljsI1Tg3UVVXTp5nEa9NLKjPAeKU+3b121
+OxRHy5/ualHtgqNixvKiyXmi7LoepkBsfUBr0WFpttncMqXyEgkcRoyF69rU8flXYno5AKttPAN
0oDgbaAFIZ0GNho6i59qTyiycDVwb8RSzvC+XLCewVhynmd4iow1OmLxCizCR8LoCnqfXR0wZAGO
C5BwIrl09W2PZJXBcIQ5S5LPpw09Z5i1rorp8+VYVVtgs5U7u01sz/RSva8/pjjNX1BqUHy2ZrIE
j0VvXmg1zbgn3GGwhKIAKKBezZYymAefUFRhjM/x1JKlymBITJQ0f94AJWkW4luVNoPbAwxkrE8g
qGn7x40aiE7GmvU17hNRag8Y+oXVmgFWpp7z/hh1B7tTn83PnDcaApjaYygG823L6/BCKVZxqpnP
Vzi18lf6aNuA6UoEJ7SEaktr68NBQF1JpMMdyVAPaHSKfGUZCB5d1cgTDscFdHvYHx4cBoxAQcEU
I13p5rMqfL9vYJZUWbEmkuI3Xc4m9Kysz7tVo22+p6/9pll4+CLoDb6xrqmGzaRPTE7vySHa6XM8
0ZXmE6DakUrF+eFibXIWxapq+SPNfttDo8g1mG1VDnmEA0Msv2zAHqDdyds0ExWT4pCHAWFe185U
QJEEcnTszf52AXeqCe7oOilvJKA3/TRUJO0nfBDdWL5yn17nxG7Vh9MP0dP0mXE+6jsLYJ8NU3Lu
nBL2mS/nw6xSfq3zzHryq2TVFAr7qAtYsCK5Rb0CXkxBjMcoZk/jEy4RdFTc1x1sQCYeFYkOnVKQ
dCwBDEgo3kuIYZ/21Zf0BzQrrFPpuFC79arq+XYFt9Ksn/Nb7vKatdaXhiRq4Xh+P4fbN50TY77l
KL+sVHvBmuSGQu9odax1EvTl/YQVs8pvYSZN7CHghQCm4E7fv+byq0ml5YcnUB7SfDLEvft3WDNg
jcMF52Quf8G80iAAyelAIrzm/HGZiDJRJBskik72p19wa1f73Vbv0JuUa2pHCZXN1muKH5d6NXJS
FyF4cIr734VJAGcopx0p0gE5bVUnTjM3zoYZyvMuulMpneh3v7dcdALpOfYpLYFU2lfiPFdZvXmk
WIhEPFoHidV3QC6HQNZhOm/DJDNVa7Fl0dnmm7RnNReOVnWHW106dwHDtAtt7EWbE1qCZm72dD3B
RIn0RYUSAjCfouzZP8lxATFrMbgJJ5SmX/HyT0ET9L6qj5yip0OfezXCirKkU2pTv92221JstGuD
jkl8x2krwOVPWHQyOun7HACh1lq8DlttIAcLgXxm2Dj8drIVPF4HUW1wb8kCHdoft2bLHCuoM3P3
A35URqqhCMi57Zevle5WyiB6kf77Xr4HWMCLL+7C2ubic+B0Zf/v4+MDRAJfxB7s+qC3HpmTRvPf
vxgmErauU3Cfb9OzDHotlEUkIxXmTfmRo3TGa2MK17hvKDyzRaCMGpyyk3QS0SO3N+Hs8N4C2cxM
VYHuME4cbURD9QaUqUsQJkg5JTF1RLOz8NdCYPo8IOSE9bNkljFX/HSiryBq9gu/PaP1ZSWHZPAn
u6sSw2jYy+pQD7Z3mjxA+pW12cqN7Qwv6oSL9nCfbfxKiCMGT8pPdJiAGnU/9vGvYox5KvWaAYap
BFmP0u9koCxKUDH7+MveyJ23SY3yzliI/bfT4y0cv+8P3dU+oMDLiR0/fMjY1C3jGZvuJXZrw/LG
PWoT5THsgz8R6hKoPiosee006OMcTo9pCaW4z+TseDxQk2Zfij4byV/75btcIKq7NtDbKus0mwPs
zHTuVXgacbiSTodehARh5IqecgYR4EgNDXophvzLa7ce9gPLEUVDJnu48+FrGbPUa+FBIypKrK++
lUoRbdTqzKYT2ey2SgxwOvEQmBnVpYymx/v+vcXMeRGtXgBEK0XqGNKgEqdm+iktFWsrvr8BCJ+t
r81+xEL9mlHPi2JDPxYs4qQss8UxGHCkgoiMyW0C4d3SboM4OMYxijkLT/odDxVRFVIN/nridod2
PESk+rXCPyBJ7kghX69z5qv+vLD7SKtNfAdE0hLUDLb3cgLNaF16IO47DNp1ykSIvPnKAF9xOuz+
91K/tkBILJYLidigDGjunbNpvI35Em4uK/59zgQqa0w06QHmZHvprWj9pmQvrJ9job6g06kMj3st
4tko1g4qrfrhtJkuzXvQWgMmtX6483rXGuMI1buHW7lWp8veudIpUvsaNyJfLBa9H6w/o8lBk2ss
2CuYV5mnSqhY1V7FlPvwS1Yf7uI3gIF2gL0PFrKXZJEOTqAzihdXStd3JFHQ1LBvRUxu0Cck4Nsy
qnf4tRJzeQsnzLlBRcPcJOn7a+AisAa7dbFsnjQnIDgV52Yfujy8rvX6FTsH46Hr565zOVY0Yo9C
6HS8/k7afpcTuKMNYaRPJElQexgZNb9uowflG9kwD6fGb534J/2/ZO1l+/4XgXziNwZa435cISY3
pajfBAfJ5XoTCH5jQGEvhfUtUFTBOW+3b99cbpwwBgyGKX3OtX4r9Kc/coKBHR3wd5gTHGl6Is8n
Ui3vlPBx7WUCTXtHFLZ9Qu9vWjvd1awuI9PmR4fom3kfrTB5/EiEWDjVKnXbH3L9eF8UuQDxCQSn
3qgFhEmvMwmrZ/jpMj6x/ZMNwOTsnzqKKK5LSiugFXTGe1fHlUQO9k/+Zh161ZxEtkEbQ24aYCaN
vsK7Ad7Zue/r6OK8MkzQEDw+i1TlVpinjcJL/pKguMBF9OyZCk4GB5CRoyZ8vr4HJnG4XjuUHyru
3F3jAd5Q0bvfPVAuwjf90v+lrsOpcKWt4O1IzTB8OP05/1qRCvd3sPaLHWXJp41fgT7wamOsgx8v
4mcoeByJmAuzlZ0hI8kwYvJHjGd21IVEEZADyOh/25ZNQcysIifD3LhxiTWmcSc9Qv2yfByXPKEc
tsdBvMvd34RXiZpL9YjDMLblsOx994gR8S69b+mACif11gOz3Hir4iC0DPVSJIRoLUduGEIlxGhg
HHlnlnqd0thlDB/MKhutTLiilHhnvdM50BYjar6ljqY2/CTJb8HNt3jHwWFnYlvuLTkLAQ7eCWpj
Z77hPTdiE3F8rzU/gdo+KqXaZShq18XDjoFR1T2XBwPRjwGKR6UId8+fgEgo+6CUxkceoXTbxM20
Icq/somzTzJcSfXjYVS8/EYXeiYITtDIpTAgwheTTl+sP+E4kOly0o7G0ox47xA5DU32JOvlPqfq
9B7ozJ7du8Hn0jlD64ip/jfR40miyD8V9CiX4U3PjMhgLq02D4dE+GDcobs8+D6Eb7XzFGmsDirV
ppc5HK4gBdY8cvWQNSOv/B6Tx+TyNcndQm+ylp2ZVZLnuWKMIEiuz0/S/AGtVXxBmRxEJhaaEkgX
RlTvmkk9HOv3BVHmVJ4iWh3kNUEc/8qJuJfIGSwIrLRc6ykmu7KP+fwdENXCxwD5I/Lz2YepPRhF
wyqKLqAawqyuf2DwuYE7xV/ET5qSlk2AlJGMywoKkH8qK30UZPiAbGImzyYTUuoiKyEHO/Ww+rjd
r6gNFWaWivPPDws10JK1z/8Chkl/FYXNjWpeJaGoOUkxxsmetnXEkiE43OpG0FWqpZaDbc79Cnl+
UCLmbviII9EJsePulSYqEXPqKoA58c3YUv9BUKCwh4PMaYBjGGpzDnVjJFw6kKITJdQcCxG+2huC
H3Q1ye5NGpm1Wx4X0SU/b68OA65bQ5BBCcr02y604ao6U7JAmbzoEW9JPv81eDTFfhQ5CPkdKxsB
nbtlKggwaw5zvKKNSH+pbkhRjVpRf3mDS0jxELEmdG6sQECJMTBS/KsvEuY5yIcjg3Usgl/DifLj
e8gfsPDqyhW128hXDlb9OLD7M8to9tKBmwOK7MYl1FoQGFuoYFn7Z4DSmitUGdL1wy2BLVmZeQPP
g54RRQgu/Z2EvcL61Rzeat7UsMwEZ3y8v/P9xYOeV1ELhLnak0OLt0e3JdgH7T/al1iEpOiC4KYN
Lr4b+ku2zipxzpNcp3F9wedKo3GYpJGEOBVuIQP+vl2qwRDi2OBePRUEEvzeDcS+LOEm0rImrE6B
QRNzwmHgfe/i5vJMaQWrfF1L3uLmJIKND/fq9LYFh1BwBKtEkYtIuArDFkQrxcoU7vYMf30QCmZj
41Sh4g8BlyZV0j+eIIln+ptYt+VwsLqpRY5AafJUEeyYpvRmVF4lJFUmYOtwc7JUwHKtPyJK8K2u
g4d9hQsrNeV9Amr9JFZ7jdxU9LsYX4/ndVoos66IKfJ8dZGdn/S0QhvXsm0i77FIgkF4IWeKejiS
mOESU8KzIYuWGksB6F0B+YjpZLhowy06aYPQ8b5YMSabDafZiRz97myj2gFNLAMKPeyIaR0AxiF/
kOO0XJWzdlAr/PZtr4wops+ZAa3HV/tFcdfww4UzdwsURoPQdQ05WnWUUtxOTNpSqhdjF8rf0XUf
UfiLrAIHB27KjfJtI7TumpLtYQEj1sXtluymZ2bmqpKISOCLA/PFUoSKc9n6XCexPc0a+jtNXi0r
w/NxBbC+CCVnl9Rtqm/86BS0d4rzr3eJP4SahK4CovEoNDY5oFtmSC8gumHErE2o67M/G7QgV2K+
i2cmEFdpEo4o6TzCa80qu7v3B2YybEbsigKs/ndb4avwQY5822KsU1q/Vi/8Ju8q0u+bR8XJ8+EI
Ib+XFJCrkJiGN70I5tqRnRHcV68nFMC9vi0Bq+meEwHVrFfdKEoS/a1apwrjOEN2IHPSFAEC/n/M
T2rMN+xhQhkpbR5tI3gJfhYXWP9V/T7N3CKhmuOa02tjMadsEStA8uMfhODGL+QIRHZggDQU9rGL
2Qu9vllrSMdke7wB+/SdVdlDZ3rioANPbzHTjYxMCFV4Q3e+JX8LFa+ZlsSPfBvSE7V0K2rMWqn6
FCv306ezx8ENCu00HyotMOJemWzsdqwWe73ID3AybUl43g9y+YyKZwH/e4G904RV/PILY9kg5wBr
h4b+UqgQxRxzOlKlZHCHM2Z1Vtc+sAaJIOJjyIMEmx7Bv8Sv2Ibd8rYsqEGV/NIEdTL2iNDHSCOe
YHe16m68xZbHUYRyOcy1R4YdFg62P86FXazSUk1Sc/25Sr2pZrEcuSayUH9nxBrV5Cik08/c1ggn
0VQJreEZwrPLR3KVmkwBHTByX9+zK30DfBNvrOyLR7NP4S3CkoW9nfph9dbtlBQg9sOjajM9BBqR
3KEMOHUbDpc0RsZkdMhY6km2TKtA1q+qBKr9rZR9mYx6z3Pf8L1VrCdrfAuKCSZwpCc+gFvz0aoU
bFstcfSvXqo3774vBOT/TObdsKMVWRrMI3gYwB2tRbHrwBGkT+B3O+wHJ8AWp1P6TZKQEwS0NJHf
NvL/tcMJ/Pt7MZ2/uoLOZ4/+ZkEt++L7KsNfTtcFDXCQq2biVDCqw5d1DOwhf2w3J5cuWZL8byJX
bdGhjbuCS2YeINfays4XualjNzoR+srUUQbp94i7xvNsEex3qwVNfRfXXZ5xfbM4jMn544ST1CRJ
pHSegbV4z4+QgetWz1k18uzWiOfutsvXaoVklulbKLgbug+JFNTBDA2nJAUJ7o8wKy8zD2vlkd5v
Wms2bG00BMOJJgUiR6pExtEIknsNw6ErGARh32MOdXC0nqG/qhEw0qdrQKoDiKA5OFDZstS0ty2S
3Q15eQTp2A5PhZ8M0A33NCrLfQ31kXrJXghzJgqyiO5V1UMe25Vdsv7wObhFA41TsYSI09UTYuVO
Dh6vK2Z0dVk+8l2CjlncJiDsUQQ6nSTFpoQ26dBbgHCDVyks9SboQMwqOfbIPpCGdUy+lTKCN15g
6GB1/48nW61D4TJX2FoHV+Df9QTBmJCNg2ohRms+xzLA1gZGxYjIu0sIzGeq4YgvzYtsT5TpNsEM
fUHc3uv4UNhs+C1Th+/Bkg2yAo2uP3swzP5Uo6/8nsuFjQO1SfTg99yntrEkZOxtlOTfqYbnl8xI
zkzezFakVYFIrnUzyh7x5fdSdb9DLepWpR4ahOFsSWqpYjavYSwLAn6iXE9rSyVchgQnac16W0kI
mtcTNvvK6AnqgBCsq2a9wAh74YYCNhj31crsoazK7nvjM1MZXXr9BjkYoykZOlRJIdfy0+hlNEs9
CIdeLy9CEx1a+cuB4W/KK3qoPFz98aKEXvyOqsymXV0MMuYFlO+NrgHYoQ/Iq2TyT6/TNoedzgTR
/Wk0ylHQnNCsFaFUYQWpp4pxvnAwM+CPD6zx6UVdbMhe0keFx2h4RlBMygwT4lxHcTzrJxpX9OQZ
Dn34Sw47TePIMGLnTkIe8PGdFKYAlLf74JrfTaafQPapXVNkEnqFdfZm35Fxi8Mc5Ns84S8QewyJ
ZF5CaXXRB+DEBCDRoFNWeb9s3JS+UFUiIRiqUhPdy2K+xF/xs06jvwxl131+8KE8mejz7O5JOE68
ou53u6+LlRBq+dEAucPnEIXlzCi3PD4Wa2FB5G/Ebv1ZXj6WC1Cs4yeZTgnlFTNKxdZh+Yyq+rH0
/e6VT9rtJUwv28Asy37LuyrKQPC7tmoILZte1AVmpiguuIE2UNNxzjofw5EtiI5KWYtz+1mFNa+F
QnQKXkXcaXi52nugNaK+ctWFFM/Dw0yQCqsep8yWoSMMf+uYuilhYcS2sFfPz48N7yCz4bUbpger
WTsLxG8TDuhcLgSki2wHQwaeF2mTxjSgIexEg8ZMd5/wYpn3muQDZa4OBn6g6KXpJ6S2exy/90MV
2t6fNTIlGoG6Q0iHUJEkshUk7UGrfBOwZNSq2XTf81zc2d0NTFbBuSGy07C4e1T7b3ZrZZBh72LE
LahR4PJKtqTbxwS9vkxFxXyd7wPt/6FaNrGa0RAHfWBv8Aifxvl9/8S79tH/YzEiYw2Zdmjm9GT5
g1oCDkW7KJL9nRJHQXc/nBwB4w/D9o4HwaiUIBAUrqGsi8s7PQvaMdQlRzUsm3/Xzj9iTO2W7n5P
tI2Dwk6xWx2ipqSH9LHs4aAvsvLZ0GHjUhlYw18Yf+zOXkmuDiLW3M8l4lEfYYEwPW+D/2Y4DrWf
7keMZ/bMwyypUhX8XgtdD+lfJMrtMmJof97zrWup921MN4evKC/hVZX5HjCjYsXmrjJjPHv6BD5L
+i23/Sc7ymnwx4ZUAPcsAsYf7NxZsZVVBPDyv1kLfooh3ZKpdyt0dt7VV29uqrA3PUHsVzBmVpIN
4HuB+h4fJGe5l/kPPDc3W/C/VDBbgqCV773bPRN3qocvl2kBzhlFIZLm2DnclwNhHuMOFSz/wMv/
PaHb2lH4kaMqzpoqbbK74AADKopXGgRH1tuUPpVBJxYBwbuCC0LF1JBrWWY1C8WgKqrIS+ESiLYD
5p9HcmaFiGjNT4rlz04A1WsnEREtxEczZHuwLysFe3Tog79iDSyV3AfCxvB2bc/GYxlNQhq/8/9V
Tbj+zXL/7+iuo9V7vYxoYFt+Dxe+UY3q+XCU7FBNisW7TfAzfPYjWpOY2dLT0aduHl3HccXo5Lb2
cENRodGbZ47YAysDGD7Be+hfExWaBn58AvgMqsDjKd2vRjzdWpAIk5rm/xyRcypka3LMWrnQgViE
Ir+u7qS4u7DkrzWsFIW5cP0wI0taKM+RrnnmP7BZWmkWjB/ibyck9G39ZhtSwOTzrRtv/hZZ0vmH
kcEkSfGEevqxeYRNCgswWJZECrMjAyujA4Bq7kxAifPtsertIiHpGimTBnqc8hAZ1NvbLxOhNrb9
SxzE7Pdde9kcpTHligK86cEHEwDElrm6225DXszIQSXBJd64VjonYmZTvWzIwU03wWAvhEC9R8Ef
QIOV7fxQWZf8Oa9yGIeuXFERyIWYkXxx3lmaKPV7767NXXpgmY1Ax0Ffs2r9CzTPGyAbmuGAj9fM
xPJdAcodLEikEXnBHZGxbxjH6xmnT8RoiPJcxzxrQtytCLxbuGo35HMYbPtPr1IIz+PfHxfF/qwd
swxmElFi7oDy09F2MPxBvx4XLXXdt4kW08bVOnGRkzhvg3i7f5IGErXN6RzK+/fJdhu0y3WyYMeT
6V8dJNs1UL2DG4H8k24ecq8zUkgay0eURsBMIGGM4uCc5EQQnKcQsSE7Z0gcP5FVhK+YROIQP8bY
WPwDFSe188hTmpsiCvSJbPxA05ld3fNP5e/wULkphiUBfMsGdK4bkguImphpplvciWJOzOwHp7kf
Ci+vNAttAsUeR/BwYkUAUjpu+gn04joz5ewPD+4Um0ePE0eburOMmidlI87OM2TehMfU8l4HfCgO
Zv2AuRghUJ1RgFQxlgzbeqnSdU9C5siSKgGE0QEIWpabV+hLsDPcpsksU7kShZw32DQvwmdkTb8p
GPx4rbXdrA3gIkPB2fDpKGUwXjoMsUVKL58LtEe4yawHPGF1WLpyrCKDZ3ZnD63v6gLyUEGh9DUd
TaB7M+wx8wDnRjy66OaT6JtgUn209D+IPBJM6JzhFwNXoBBlLyqOwrZBgaxZ1j5VU8uTbKEBj+fe
aa/gvMrMVobUam7OBrjA9LqGEblfBOGF2zFg05yZ7N8QEI+XTFNuGuy2u+ERjF7yTfFB3Otf9H/O
0ZeUgMZ6eYqi5CdjzJMRIrRWYiBqsxvPH59mZY3ujl4OuQsHSDdo2y2s4uAR9qyuZez+riuO7UGk
uLTT61xlXmE67tRoBnSnxrmgqfzm5WH1g04f+RPOecQBmf8N+bj4eRmGyv0mJdB3bqIQPLAhgin3
L8JnJnFlhHcdznNdIXfpzvvZ84oqcrbcZMssrbz6mJOn6TLleQZsK6GMdygO3//sC+jzPMbRU5zI
6qKK2dltwX6zwN9YlHTuUrBC8OyoYeJPEu16G2Vq2u/opwBIvcJEtuwtQ+ErUiFMlKA2+hfE1RgP
Fda3Mv9vrepzbrboCh50HoOJUt7aEsmS50FrUWqkhCc6+p0oqUBqDZB+G2h6v7n3/+BORkGgiJ9/
O+V7Lg/AoLBsAeLoUiE5o07/A1D0gnLvs9ymHtGy4Ga91YzZTZuywRcUQApNjONth+eK8PHuSMVL
0J4h9Eg4rijthQOP2GA1g6TFJF3wLUnycbk8dLgtYZox1irKCUAKV6j+wUxZu67aHT2gbz5zh0iG
wzaclCWSeibzZ9mOGTGYt8A8jPu7Jnazi6N22gIRP+ZxVnrIsaiiFnp1rOhjHx5RLnETD3ghs2+e
MlWXw7pVL2XeWJOBj1MJEGMfubtGGSWrZQKgNBT2tDAIgdpmq+xQkl00JOGsOl0EGk6hydV6bVgZ
jxXEgXrLXj3O014vl0GA/h7eZnGBFLvhWrSMDJr2iyI7mz7Le9BuLJExZn+Lb5uU9sOTFZA+B4FH
ZDUnZ6gcEa7TecEHWUDwVTj4NdZYCClsPuNYrgnAMwprlj7DQ44r2WqiwUrGLPZ89FdRbuamLU52
LkdEr/Cvz9b0K456axCJphBB69Jdv7sUrSQ9jhPRsT6v3S6LqtQFZmyQ/R2EKQxi2AeixWOC9i/N
lfIjKNk+VRddSfPGE8hhu7T6xgEo+2HwQkv/fUQkyOKFU/xFOjdTskUZHdz7S06296IVkfAsYPe3
HFejjiqogPJz+szew3aWS/4YI/fP6rmcQ7iJ1uvtXWzqfRJZI2DdXsSw/vRuPEatTs0Cx4V+rn3w
ZM2+B5rRxS0UeSFfeBkSfttVwFm+gtY4zsGLur9FDK2RmPhwwyfUVDgm7+w+MawbOzRE6paP1juh
9gsw5t0JYRcNBOBm3XpbnUWf92U4T9105599QTNukAq3vuj2XoBRznayMa465cFOcs+Wo3OGM271
GQFHPtFT+xi94ayqPvQLXJrcDstqHydSOxx6Wo/Oybd+dPcBEe8Ghw8BocGYW+tGI7v/d0r3MyFb
oHBzQ53lPWRVAQ6vb2l01ChBhGoqzvwDjDWxwaokAR9gticnpl7sheb2LJRf58rJp7reYYt8wgn+
8Z1xddgsjZ4CTOcFz8sexJ3I7M/6clvWhR5wN9QHT2tJyZku54mbLfuXq2siBVqKaIj6mbs7RTUE
qr9TpZA50osRd2iyeEolrRdS4iynOwUWHY7EGeeHaAToHN1Jc6IOXXfs+UWZ6MubDZz53E5Sq0fN
efxb39Bj/9oFqghkOeDlg6xg5XR8PKksieEjpEynAgS1LNNpp0lwe3/+0O090xa2XQtbPLYUte5B
PSLOX2IG7cNCPgHwgXTxB9ON3mKJFWofiyGFLnLymAdT12hLCvZM4rGzDBwsm83B1hxOWa8DLRs0
rXkcOrbr/O7SqH0wqPWBxTcMxjWqb8tUVQAHw+nQ7ubl4x3+uI3AkBWfspj3c5dQYi5K3VFfdxgW
eep4Pf5IyEgn3+k/zL2v7DoK6dT7La9hxSdizYOtmlGKUmFy6XTjNOe1RWtVWZB4jLVA11eSb/D4
w61yv9qBjgW7MnNkzbZ5JHM5MXsE/SyiN1AgytYrbSSa3fnzLLOMI7eml/vdymdpkL3VJpkKIiX7
9hq9i0303B+fZ7Yc7bz4DRt7gfHg3crh2ToMwqL1Lbawq6cSHgB61GL+AqvOYY2EAlsDZPx/Fzg5
4n5mik8k3eYr+3DyXM74MtzX1X8y2Fvxtt9kdpDuGZriA+LRnyBymzxojiwHJYfomK7UY9uX1Ub3
XGOZtuZvleDmRtQ7blV2RqtF69exjHlKeAIAAqBJb9q0xGlXM+qF4jrj7kZcgY2mupgbby5+QfWf
T4C5+xdGddpzfmZ6K34XKNBnuHzcag1KxH3DlTr7FmLThCeUzZ+7a6D3gnIQg5YuU1A1snUSJdag
98v8UX93VIuiPV23KAg0H5QcNHL61TdUZ8HC0Ox2DaZEdDNaIu0rsMSqkkNCJvXUhCJ01F3m/5GY
oBYY5o4MY50gCaeoOCA8zjICqls5ekl8vRUkP0rOmm33u1Cg3IiCFQ/izzx75Oj8bd5iU3M4PNRj
NJWKdwCUhMs071P0y+zKjL5crQlnQCPIzcbB+vpA17DU+t1vVFJf2zvAsBukWQwdLf+5e00EOELK
uj2gtnNbQJY7piyZAVNJ0+qcVzWMHWyNx3yc5OXu6KwnSSbuFsBYG4gaSmjt3089JVvo1ycw4hFB
Rk5X8ZCBqMjVGgG/PYJWR/zbBtyJWCFPQSjSAIcpZ+io/sRIPhrLnL8pMLDjhmdOmVEfEp4wBoT2
J2MqR5S/NsrH0/YoeRPBSKPvzUExE60Pf51g7KCViOFquJ15sEUzVkQ92hZutUDK9Kimi4TD+83T
DbCyYPBMBmMKxfbV3o0gw7H7adcPLz+RTZiFc8DiURKw9jF883DXOw/ruQRNyTqEf2wD5mDUL1xK
J+UdyrbtlMVfXnyP5Po9fsXWEdtBR7EB6QL5s7wcMU4CD9ysxDuYxxhaVaFu6nQ8Wq3mrDTLbR6S
vNqOldnnL+s0db324/e2lFW7lDVLQWR/goc6kosCzV+51b2uxJPouDnxBKfDEhyhSzwvHFAg9BbK
Fx4jdu+XtfmUh5vIHcIDmr4wwPgMn8deBHH4pcWXFJ4yFx7To1gvj1w+RiH4vEb5dwhFiP836jiz
YPEVf1DwJ7qD8vaKqkMwoFAl+NUAyQ1r4cbF1MXXnkqdzI8drBHBsNvdeoabE1+8tC441ogEjZJP
IFQKx0keONM6+TXATa7HKoWmER1o/LRUiFLDansVBh6hYBJ9UOtWkJolt9pRnV6YSyEaTHMfgl1e
zWQBGNihl7nYQf1D4HCyi4iF4sOJWkZqeA7NYV0f2sCMqn+qTywaF7KyBxVIN9CQYxdL1U2aSLW1
dkFlqB3iZWASlu/zwoamm9JmZdqzJXkfSfN/0i560G3fi/lC1XCEItbEHsbV/Fy2xXoPv03trUkV
rsTE5c3w4spUfwB/VTQL/Teiz4BdTcZqg60Rbnppz0ai1iLktIkNKEwcspJFRabQ+IA4OX1/Z3e+
jjfHYiWP46Fu/uCH+p9eMJqhsyPtj267b/L6Jvy6EfKVg+P8CkFx7I7RZgfuckTm9vxrIb+eWlrD
r5zH3nc4KJhHwSfDtXVGMhfz0I23HTw9wHvlRKRp0t/7fDuAwIMYUu5QEW9Ct5N4lcmzHr23HuNK
vM44tllZ1M79UiRny+5h+yrH0SH9NwHAWmlXkJ4YEMBSgRiUuBrNOl/bJhST6ZGELNLsGM0Yec6+
+UiScJjK4pkz3nSi8Y+Foi5e4WuL/zH09ExVQsPcsgYC9p8N7pmZxtHBuHfKjM3jHWyiedN3g5UE
/gZ2fJzxdZkmXHX+SV81GZ7LIPjtVZ2mlk3vHkU0TAo39Twqyl4f/mA0s+uz5wOLb9PWVajdfCcs
Wvw/Qgv+ENQWvLMjwHEOjA2HsA7+Cl55t4kVI9xkPZaP5z0aXhD+b9+1DIfkotA18A0ime+AHJ/1
JCPzSP5u241y2voaFsAVFqR0juR3ieRuonUhqXJ1ViILNr+BgxTt4OYkOjbyMhoyu/iEG3lsilem
qh07RLYFCOcub6PCvgvET4BGRXCHTR/OEfyE8N17Z6GHNl0YtvSq6DuM6gKp82a3Ocw5Xa2/w3bS
gznBHbLplF43An3H4Uh7CzS9P0Ktk8NmI0Imo9vDznbf0ZcZczFJWeMQ1sT9y+5RJaiijLXZIQmu
I6NtJ6gdaE9dWMaGJW6zVIKeZdWwff331nSF++VkO+ezW5iQM2W+gTMDu/zaylFnp+JttZnMnGdt
2829zPrCObdpSa+N0LV0aCDdFVAfAT2JX1CZH2mNKgJEH7jYaErcp6jFWO84gzrAtw103hJzUSeN
E21tNztvVvV5tZZr7k1OneNMrlUwYpCgX/bACY7LZYhfcfOsR/+Auy5L0ptnG/sltgDSEgZADn7l
uZDgoktlt89x8QYCRv8WtKllReOIWkWP7kv7aw5sGtqMOo/hQ3T7E56yzSjROmTOIFNhX2Y6aHUh
Z/p9mPXviiQsVqsu9+lC5n2X4jRcGiPvKJzJP6BUOLuedc66w8V31YSvCPAuwq3kmo8Ny2dLiZyE
OLD17cKTIQPwCeLuu/x2rX7tliFJRVryxHhGoEvlqzr9ubQASoqqzr4+tOFaPVdTnE7VsQAEJc/I
dwL+yneWz+VJwMIlPUNG6+n4uYhLD1h4DGs6E9xLbEcmwTevP8qQ1fxINyLrDJhG5GDuUK3IBuZw
hnzigkWfnDbtlgsZpSxgYQYq2gkBg0sQfIUEELayxy7eyBN7NPGFSMv18DMqpuL6Z6l425mzI7Al
DuNg5yl1MKWanAnWc2qLZihb3tXNd8NHxvHU5GKHNktFOlv5LDwwdA+6pS5Omsly4grRQEJCwJrW
jQfj8rbveAKPbCmSLlqkyQal/Rcqr3glfE4JPOIZ5Mtqzg8UtMe1hWcCBPhE02C7vOuXm1AOnZYs
0QQkKOWwmJl/tk4OcgRawpJ6j7IevgFTZiFrbXeazU+BP7RkFU5/VJN3w6/x7GidVl0Zuv6sNYoj
Z/79QlJXTv3LFlvQjKmD9PDNbGxt41vdEe4RavfPz/wh22oDBvccAU4z7k00Ib+6s22z1dQUcw85
NlC0ollRLAT4l/qAODGB1g4cYBEhSbfsOjqai5qdJYcjmnTIV2AKcXyZxydg864E4OvwB+SgYt1C
RMSr/4mzmi3oTY9XLjk0+8+Fcj9WQ/Gg86ksw1GrvIYycK/NbH28hje5eIeKI0Jq1eyvnMbuyLzh
tiEErqP+xk87Vzmv2y8iaho+iv2Bov3oGWExAW7BeJ5HKGFwmjyMGOk9+v25ZTgKjv9Jv9Uk/SCe
Idqbd7C88JbtFNecZu2QdB1qaNZQhcd44gHfT6lKN7SVPqtqH2gvPMVhDeZqI/qdL1cL1wqSOvdF
HoSfsEerIQ9uRjZuMnt4hGF+aYZ4LL5Ei55bq/QKfeCsgghj8UC6q6F6Y1FSIgR5fdCtshEAvnFE
2YbAFkq7ultokhA/o+ORP0A4WjF///5vQTeetKfHojW5ChtBf7CxpxwQp5D8y9k96UvQFYlxsmSu
vjvL/BNMcRaV9DI2cx11T7fGEcDNnVmJGmauo3H2D1L/8h0rrtBGmudYFqZ1Zlm3YTnlxCgeihG7
ixzhVtOM9KmbQDs9VglRhYepBv6420HrDtoVeuUefzPmPQVZz18H+Tl6xoEZ+FNihETY0Outx3Pf
WJDPKE8ef1zGFYQiKD8C6kX/eQ47WHsYWqHoAQMAyJ2ZKz45wdQ0CkBfpzCtj1WajattrD2+J2S0
LSAw3e+Vvgcfh1PfaCK/0NqSsJywqIIXdptTHYtgSYDdjUZw4ngOcX3htMzQsBBatvFSNZoisifl
JepNOH+XY/68mTiAT5kgbxzisfHFG6smRInwkWHy8Fy+44ew0h3fM2PTrRkwuNX/gcPgbldV0afx
OkAaeRUiguoG63ysgxinpvO2BYeWNURSC2DnRWqj0PWTDTmfpHdGAsieDvOv+tQy1ElqID7VtOlO
34cH5UXYC7D4Sh1qf1M3PBmMD4ORwIX+BNYy1eYu1efDbCWkLKojP01VlYAsAMmyWSk9tRWRnpF6
QZyhlEoYFQOhEVZ8wN9X7PHgG4IS/X+MQjmbi4TN1+boIZZkc9EgH+/oUeXryaN6FAcU4KaKztG1
KeX5ykeSw2/GV1GKdeJarg8uIwkTQ/tbgBmGBJ6dzxIs1XPF1lxQsWUtduc57VHVGCkPVsW0aBdK
VLEBYJ8lNk3qNRQbjNLBWQF2TFhVxNPSOeLx6zXUEJPCXeiXurNIWhe07ruzBtGVGLa9nt5qAwIQ
EV4pOMFZ4qrHuMixEyJyFZsNQ7CBUmlGH9ONM3vhiYU1IKtZ1UlMzRjK54EzQlHnVvLFSxuX6tDj
M7QnT9qV15+wdt6UwqOGhrBAn/aMUVKE5oCm1F2KqwOwqFG+fpd9HsP3k/TYsZKrKy+n4JBLuxTR
BF3MMA0GJl063vi87payC0Its4ScHNxVYTF9wXhUFBHZj5ZrrPBUhzwpl+zP5V5yYhMzUT7JQQu9
HD9qE24SaQJ5U+5lZl0vB1pd0NZZoAWiNv4DDZYx0NQYKIu1bjEybRR22zEWM2PWADgXFbCT4g51
JWVjVlJg6Hy6Arhf1DPaQwnxPVWtfaCEe+oe0pjPF0XPfzxH6Zeoz/95g/9SbH2RKKXbvITvqbRH
IsiuaNoAvdg0LTa8EnzmWtuGAWMR4GJvYd0WlauJaNSxxxa8WU3FFnsc7moKoX4Mf/uJlNjqSjdZ
fl5LMEvamg3dgNlI1dDu4v2g3Fhd+57sTONhjb5fgsGEvcM+fBJ0Ax6+dhdGQ2U04Ug9KynG6d8Y
2pyNW13KRx+ZUg1KKjT4o0TwKfaMqOIAeuoXdzcGPKSSAn1s4ASYlh/pUABDvDv322v0s9ncb2Cl
1gmnOoTcv3D3sdSxdHJ6ZmatXzxDHeEvsGuFim/e4K4PH9p03EnNM6DP9W88Mox1U7JH57Rl2Dar
PoKgmvls6ADBCVUStMhrEgRTn07Vzl2GODZ5DX3ObaTjDnIAFO8Fx9/1QgdmfR+gY0EVlvMGOIkz
EeRTLbnU0fteYczQfNiz1afDYqbIq6Bx4Eo2jaHsInheXoYakAQBkaERpAIenpPwo9e1tmxcQIwn
gAFedy7+XpMREsR8c0bKI8+Sc3javdXV2PcWyHVsiXRuHQ0qWdFNAoeHXagqdxUFAAay5mkyTg+t
bZfkxOo+RQQO38ZajT/RmSUmebTEGAcyyoLEE+p26WDy4aDG7XBdkDfj+slfhG0GSnZU5ojYzbMN
sHZux1suMfcxZ2iut1gJYk5R6BOoix/0cAU/QQ900PT2jy8HPgNEqMTm+MMQnHmFRbYYmRNdxUYU
jrZMSzfwAFtRgmX+dQxomwD3fqInEMWnsSmIF+e3XpVHxu9noNDKjT+rvctusULFRMVE6vpm+gAD
vHesLs6zSbce0aGU9qWmvP1EB8rRtYHi5K4Gv2NX90JcFzGrYMZmhaQfrj/B+ALwlvOuFBNVRmfr
YfnpGO7+EDdHqIlkhKZaQWCgMlLHfw5+ul1WdIkwdbpv+gc0QEKw10q/MAxuQV0BndENc+x/olyp
MEcEVLzVFwQyKCs+ywG+0hKEa4UODiSNagIWOTzmwQVJfMrhE3INwR6WLAsVTNCwhnUWzUfThwn0
cAG3+ohtBaHOLs1HEYlGkKtZp5XON8BxUgSr5bSFzwNm+QA73oDlDyFbpB5KVYXPYoahgWwLUYR0
X0qTPVRVEvqdFbyP+ltBx3nWcYfQxycmnV1q07dOC2EyN3qJCUwlgF007GsDrl8QgHEsqbMmOCmw
g3xv39P4FfOPnTE1rjXcj0cA+B54LIh03m2FDKWNtAGTyKb04B6DlpnCBktvtu7KQpkeOmJBI4NJ
4AYS/7uJ60bE6celjvnryI6PjcMiCsDWa/19XfcC3Efi72jSeG579yvh2e/fekiwgnE6lOMCagwk
n4bq/tlZRrepFlenUQ2fi33ZRV3+xYDJXC18nZ2+QhY1ARstZfgHiGW4ytLGJpLA1DHsMiy4JkFT
LXc5lQkIc2wNcbRdTtD8ik8nbIB8XA/Sr24HCczCChOopCu6K/dNr2qtoc+FrlUWZ+dl4JRB4vlp
btk+yyiLgYiv4YJ6bFdxcS3V6Bojf8yqCRU/S7gi9VBHvzOvCmAunQyi3XO62ank9fuEXya7Zgs6
8Q1f4Z7zdZLR+14X1Xh0WOEdohAiCX3T2iTjDDJ2B7Vi9rE6Zaa7ZNpGd6F2vRqU47nzhk4vOOhd
waqDTa9cn/50aRmd90MGl70NODzar4VfL23jrlv/YVevNIzqW29EgChlcNNk7UYt21k77shJ6+KJ
/iMWnuEdjwi3OkVPc5UWJLn5gBMiDLeRqkAQstoh7TqwOY/oxpVEd/v3fz+5tqY+JahMcuNkLBBC
CjH9XU+1c0bNEGjDRtomUf7nLB1Zl5aEejidYEOBQFq4CJR3vh2LsKe+k+6AkRerctDNce8qoEUB
2n/dVZ9Ch6b4wEHT1378EDGQ0vlQ+c1SZ/+DHaoaVF5ZlY6M/y77tf1jZg7T3qOc/m3UnRda8gNe
l3g1BkFA040+qIfPNvNXyPiabKWO7HtTjSORyxIeyoXsPBDmiR1kj0pB6IGwn7CjtnVN681WBQvI
tJ4+/XrsFV4XybgowW3OsDR2U8zLJAzPiBlSV2DLK4JVLvAQUqmsZZnVfspY34kuJbGjrEFrLGwh
ke5sZMabBDamQ4YV3LfpksvM611Da2/lV1cEBlCFeO31Ih3WZxaHDWTWaJCr40DG0TbVEf2enScY
B131YPzqvXl86P874QGcaNovljDZhumzmj7gs1tWOtDu+dvEOopE7HsQx0gcb1oIIxmuxWzI4V+F
Ap9e690Q0QHpGegy6WOhc3tZ4mIp089I5uKudQmExKGDa80Hjh6VwXlb0szrqKybOvWmyJVIg7Bf
Z8XSI30jNM3Pok/vdhzpBeN/pkUf1BVr4rMSYe7n+JxPtgBKtpMzYxYYbfE1oR3/sqp+vozmm5TJ
RTNEjnmzmZaS4GPs7IBLiLGuKQE7jUlDbGuZ4zkDAg61lSp+bPhV76xEngaKnb0sAbijV6uYuk5g
b8K0cHxx2XHNMkrltH3fKxSpP59X2XgXzFLDq8cUnnGTWd++vvSLOve3Yjm+oGZQSLf8D3S7rmYo
hGg0ujB0yt2JLWrxzmTxeLcSya42CYNgz50+BSXXiMz7CYuepHoqyyV9/dyxc0e6VSC6bKHn38E0
0ep8vLO944m2L+eNL2ocBuwuCJEMyKeSDiWz8eEEPccFAu9c+8EM1tYhhS8+a+ubx2peLLBZcndr
q9Pr3hgUz2QK2MtxSu3bACP8svPJVkqOHENnYMyD3IxPgy0A8NpgokDpCQnm4otOOMyiOTAwMVZe
Q81Nk5qATl6x9tKmVYCgrxr8gBwtHyY0XHjwYDNdMEQgFC0yAc8l8X5AOTY8z1/ddPh1M+lTer/p
asa6SkcXAHrHcUIjqyaNd93UT75d6Em6MFsTnb8xYjrByt+ETLcVWbltiQlJdHbtkJ43tlGALc4a
LzobGJgAwc/iHafliagNoeSTn6Wx0T3KCDEWq+x9eSayE9keBbk7Y0sNwaeSTv4VHZWx3FDL2ygW
qChIRW2GKUrJJUTtasyqe65/eZXT7SuZNR01SEYnrATn9WI7MesAkvGSdlNJh+dXyGC243J8LSK3
CQyT3yIQa9f/eGJi/FzWjTaKFYfX4bmQbopPJZXK5h361yHSp2L297JWN6gnhgG258rfCydj/xSN
Bw5hlYACZmkP3rrZT1uO1yTwyAMUOs3TkFEhJbW7NfONYGCRZskLXYRfqqWIT/c2LLLUHOlLNRKE
gQUuoQsRLvylXn/BP5t/yshfU7utu9RTUMQg5fqtmkT2+yPhkf8BxsV6ayDvFRSLnm+zFYA28Nzy
WD7FgkDdeL7JCXVRCxeayz52n7nmFwIzXHhzD5h041Qt3UIza+oqC8ksWeQycpju71og+MHlzVft
2pARnH1NR3vaBeGbNrxz8WpCBFHw/mYQVDEkd7BdHqi9ZSIcxKkIcTB6LKcIIlZmtvLxHnKrCqj4
vH6hoSkLzTGf0eir6xei0fv9Vmp/vaWMRYn8qQ99TUqaoFy5qbRZpKLyrsvpdo3EMKGu94MT9ash
wUHk0LOfvIFCViiReIVjxXQhSF5uaZiTdXbtSAx+Z5NTf57/DlBPnhl8wbXm4cusOI6EuDI24zpI
cLSC1FN6sUJxQU08ydX07rpfMnl2l/kkyMqDvJlkUkTt0fNY4EH/4rvXQDloC1TNM+5yMUnAemVS
IPpT9T7K4oeYRK7sRBzPpVzlJWA3pzF1DavvIR7K78WzJgYwzxwpvmMZiZRtBjupcci6c7HDcRJ9
iK88AKzfsU/ma6hEj+BHuOFkqlrQwEjYPTP/rJFQZexEaVM/VFjs3BximbOhbNeGumJXNAvMOuIh
P5f/tXYjJ1bsZIuRTyN4Czc87/9eqS+HD+UoMs+/Et7mrw5bkhevVsy04OG8XjySoWK34iTVSD/w
irHJ76MiOGUXq0rq6osQCMqPKmBZOaheV1HRJE8gkt2erm7iXmfHCS3MVasdvAXCIuvtCH81IJbh
2bJ+FR5lLJIAR/CoJY3BjjTpGuSA9duFDtEx80jWGXfGc9gKKnJW4inmNu38yfahW/9cSFBEcA99
rUOvhnlc8EIGA9JmY66plPoQU1j4qQVxQfdPGqXpwzrYm/8q+t/WN6Lo59FGTl9C4mRgKvF9So67
nVT4Unyn4gnAL+LqEJ5G57pukphd0K6X7nunhvoguBZAbwkl3JchOFXXjrNASUZEEdh6gjAgihWJ
b+fcbnOM/tClCB7cvJWUh1rSJ0U2B82uxPDyCR2FpoLuou+6FUk3WhZFR0RRyQyWafKrNjzSLoTn
M+MLO7pGVz+zIdlTcRLBLniry0mp3FM/oJ+8RKrfZv6tj3KqhGTl7Ar62zT03FthxphvVLvEhAW+
1nZhV7CR9EFWl37e6ORCSR7+qA2HqbjatIcD8mbwnmcyVtIDmuA78F8Dl4ctWQi8gqVtkK5lRLqV
rQfNCLnhxU5DOxww0l81UkmeNkBUEEV7pIeX3jHwrgyUOzEJUZslGjsMhf7Fs+aztBGpii2Kp6Hy
3NBxxCd9oVkMM6b40H0E9eyZHdH6UClvk0QMjAxYSZmFVioZ63VglrctuflXhd7/lq6wgfW2Fb3T
cv0t+1HT+L3YStqRMrs8AfoNjZGFCTSsJ+UK84UOuXqErX5MjvVFGvy7YVpEClA99aSBzQkG7OLk
I3kHoUUXb+1trIyN2MbePzX+FlGtTDd74esFGqX2feVBtCnlCube6bIx3Mbf4rWSIfNAv8pV1lMh
hkrqAKf7gRSbzUQlTSRwoWxjlmVKdN46qFiAJTe3MbQoaLhSM7YKhK6PaAd+xG8ykmcF6yrVW4ud
N933KvZw9tuMgo2lUmsP+0qloY5FC6rsq0QhwVIBWPiFSB6302xIkGk7xBoidwxEz48hDewIY/bD
2eRrY+PrG9Pwm8tRVSESa2fKKtYBg6GEC2ucwjrUix4ddqnmQKLobGDF3ACWr88h/r4gzoI/LlDk
rmQusv2kZpt9EPEVCDt/dmoXuZlVa4xyHEFjan0VxiUlxitTbc611jnT4p9HKp1O0LLaEfjWhxiW
25daKDWar5cZmE/CPqXx0ItM21SUnvdBbt5ekMOXeyguO7O5eNLY0bF7BL0e2di+4MKrq8O/Y4ds
kiRQHKYjqaS6rL0slzPCtDAZLvO8MaMmQyu4U1GSQ6NxX+BGoANBmY5pBCkrURYpotbIskL4tifY
+iR9xZeU8fXhi+1hh4LM1Mx4o0hY/FtzXNej7q0LFRDm7G8vzCeyWFUsSk+lbqxZOv/uUHDVs4LN
CoV25mXrIapN5GKUbQUCMPkAhfiXw3DWRVA2+xqoH/I0yL+7FKiBpPwTdMNadsk/5eWII3T8NzRt
0RmoQCtrIp1szGK0HEx78dTpCJwT4qCrAIdAk4w3iQHhUM1zI0MBADCf1fm2EtdOcPbjkmfodHRW
kBc4X5vIPikdrPFZnv46KtS2nPs19nwvAXAmzNPkVa9hvGC+icfdWXwKeRUUcemwhQd02a7jPLQv
wH7OC8+gIm5tuuF3B8Omgx5Zt33/em9+F1yTDx8KEfC9GdDgsmUfxMvUP7VHc4/+xXAjvqLO66RV
S/SxwRP/2rOx/CagAGWrIyAksz3upKz1g+leVQyhi2Q2uvm6hQlLFwve3Bx/xRudFgtPxf+eNZ0i
eDvE7RQhEh7/LNe/8BsIIy7eHhOIDtqOBaztplRy7TyFv/+zCiCtmHnvg482CR7b8EXZ691x1vTl
tYUBZpnoY6ssDdF7VT2GRExU+aKFUDtDoEDdJjJUdXAGccoDHVGsrLbXnE6cADrKEMoJZmjFBD3J
7b+mag8R0sTZh7ladWdVVpn6gY/+ukXPJS8heldC+tSf9ypd7NCXkYLThleM2dN18JfINpQV/0Cy
V/EF9xVTr2QirpzeYg2ut9tErLXlqPohgXE7vkWrSEn1AJrlANWt3ot2czl3bRnn4Iaacu6QlVDS
YlfLVkRBwHqUaFk7gbzlJ7ME3QA00a+fUGkKhz0KH2MK3j5YGiaMJmRqT24hM+fY2hSBBY/W0DzK
hmq6QnwdNeB86EQAigMJVYLqSyliNEs7WNUOj25CXcwdGq9/rCsWsQU3hyHhnKdP1lYbC1RKWCEX
ZNkElFqB3uLpYMZ7D83ZY3mA4PURyf7NoO+pz7d7lIR8VOj45Ak3dOy8lTBWWrjJEtUKVN8XyEdq
MnPy/Fyv//IEmUbHXnI4lagEX8Pwj0JLAX/va8TS8IAw0YdxjrferVwsBDyAGr9hSJBRRP/l38oL
fJXDi4fHQoNLYqFhu6Z5qpVnCT0fosRtImpeG9nY76lWZMEQ9Nxqiol4VLSxjpJIjMEMT+gXlO+E
RyGUPFQ38CI6VuOM+YB24toXSJsEvAGNIJYKzr3ODwHMhfXzq69Wvrz5OxgBBjqULD6HDiM9x4jh
FRRdJf4nomieBGwNX5N3ITJEhoMqokMF9x+rosHFMZC4hqF0PHxlyrJf0RkZkONGqb3SvRGQp/G0
G+Trh8RJmQmE/ctwUKlFvW+MSysUkX/+MXR+1CIwAlO1wleNPX2mXBNtr+FGNZAYnCMzhT65cXY8
EqRgwoZhAv/YCQgoQOvsQr0cLb+EWHKFktBYUuudPBal8HWQVUApC3fQzPWFDFl3rFEhCIdqxbr0
TeS8qCpGXG3boHgmFMNX2Povcvvkw4dF+A2obQ/wMjtHV/qpMP6fKmNP6aLSF7B/KqQxwfeiVad1
KlCRbbFDxZnA9a23M+aNWi5GPTcYEOyd1ON/RxNPlVtfEOP1N10/xRpJAP6Cs7k/n0wGsJ1jWNy6
zsh6SpvjrnnSAjJBd8lKYgXwsg362wc6TCYIahJBLK9v6JoRu+rKpy2KFdi71/8c2AJ38SV4a6ro
TQqafwmbNN5C1SdTGrJfRCc9TLU8MZPOz5nnVDyGxipcqDsTSx4qhuqDR/IwnrhNyDAmYbQHlaG7
wsAHujZqQWE4JoADC3QmlQyHe1VIMXLjz+Jw8RuR4kINHjUq7X+bpy1Lr7cjIVjmQXJ7R4Ou9r0x
rfyU+5yTcvCN95vTA/f/GnTA1NzvmjbxFFFJ9oXOKP/ULv8ENGvRu4f8XYCwbJcvlZXa1xkSGkKg
mwLcGRh97Z9kV2LWwOhsGuB0wH110UEI3mRzI/KKBy22rGV6XzMA3wPoJXLWS0DjtT4zcPa7g/Sw
UQm+K5DZq54xIAYoQsSi7fdIlvsupYo0AwzNv2ic2GV1mE1CQ2WtlRCxxzldpIG1DbgOS8msPGaV
liXpEXG8j64Rdib/UDdDhr9M53+uR+7DXMlilclDDqx2FQg8EqBEWuUda3I6UgKZDav31HnUb06y
8Hx9ylSq+6L7s7vXFraUaUojY28tZoAy3fvalw6g2TOVWNJq+fMfu8feMgkNKgKmssEGctqD6FBg
P8fICQCzmG5NK5lUm+38vGh778aaXnIkmAFHsRQqiTYxYGe/hBrrZ3hG53V3aYC/q/e/aZzgBy5f
Fo7R1jk6te//PS1PFJAPdixruOFDPpuveIj4ARnBoGDxZRh2/s4CKi4JKlagUjuz7Ko/0wfxydEe
HYp18Q4pg44YzA4ZM2cNtqIQH1IEa6s1nOWHDWVQj7HtMhH+b6Xdw7LgzRPDgO2xhPgltW7w4N3i
XNW7OrEOw0wH8w2Ylx6Va590icAmz2NiwBSc2nqPPviL3zAEpgy4s6esxEUnxECmzJAzWmboRr23
EOsB8koNwY3rNk/XPvUXDfIgNfnzSOuLgcV+J/fHZPpyQsrtSUr19c7xqkHSzN1Zbs/IACGwLOxW
0H2/ePnYKgCyeFqOSreoCRfMsBzZf52zOZ35A3OiI/K+R0+qAr8Hfs/GeWpUcIT3sivv+GQC1sQj
W9nE8feC7XU/rtNU+gsERiLfloKPpjqlf2RUitUia95va6d+Phw8tkuMxoCMidf36Gg1wdQlxisB
GGfHhCX79iCr1y/KDvXiSU5F8WJ4GQfQ36F/G8o0fh+GK8u8snzFJHQGzYH+j/OylrNFdbDpeAzW
tsLqpMfD8J2491x+gWNi0jkfZp/WyobnJvPJDC0QgQg2GzOsztAnM1VDvCD6ngNJPqnHF8+qB2E+
a8+XVw9pFDzCDnjRyebvB1t1PW07cAvxAlNR380aFwexeItri9Wus8e7/z4QI/lH98ZVpeOfQ6So
5QEHxBtBwXJF3lnfG8PgtAO1G70c/L9zLIWD16pD8CYIpdw839fWXAx6oP/IEvNQnKBqm/M3xZLg
TTVa/R47SIgx2HTq1wBakxal2ZP7yjljiR+3VDRn/eVabWnZ4PgelVN2rMTRF7YKOyMbaBzXDJre
LSlwg8cxcwKN1vszhSqH55DT2cV69pIJ2bfRYoKrz59ZeSTxRRi5R94K1wim/IlYfKc0+Ai175VD
lISgJhSIvkXr9W03nJ9yeMyp7Mf4XFoORbguwpAOWgArjhNk+alu+1gz/92CRX1UjCFVZM4AVBTN
YV15QKdJYs++ukdk0oE6bwHgk7eps1WDuTHje1OT3YDsIbxTeW7vrHuv0TmK9MgBPUGvcjhpayax
MJV0wLeOyhegH9reFbMyW8j7J5D54L6vdGU1tDQde2t1s5ZGuwVKQUe4xF7mLSlRQXpRWnIeXiRN
KlerWV6dGtZbj+TN+abRUyDLgW+2fqV4P1JIM9lIYsk96DZ5az4bRRBxTtIdZfLcvBKOLPAg2iei
Aa8UtrRP20e1r8rxmy2zwz92X11pkhvxLuwVGtjEu+Zc8Wl9+az1n1cSdP3F7syGv7RzCI9nmMul
8BkY6hTE8e1DBlW6vZCTqriUGQDvvt3w3dFDqiYBo5jYQsdpejEVULIX+DtzLixaAdSiQtlCcDr6
Jso/WMdCyWymPJqFIk55dL89efrsSGtmeJjf50/Sbp7C0IsTo8uMFXpaf11acef1b07uln3uTXXI
CbSBVvKp0OL0NyFzKssgveTqkqgGuH6hGVzG6Ek9Mo9cxPbESQIDbz9eaA6NLHi+Z2fSz48+Xdo5
sq8QTJbczKMwcAF/eX+n6CspFDG+VjvO5g3ZuVlRgdyc5bfkZhJ4ZdtpIM5nlgkUxS5tlzGKdO5S
eBr45WYvAyZHVk1oCLlMEmqHy1aS++8m0HCgd+v0rSzKclDc2K4T3eDUmmV7uRafXFGroZHsqW3p
PFcZaRLxtQPIw7NguXmrilPOoDIAsTarHN8GAnLIydq91YTMk2Ud+BhovKTpJ7cN4lupd/QXcEK1
aOvc7Nurna3fRVWQnm7SoVilmFDSjQkmiIXYyXSOG8tKoobk44mV6wNe3P5cnJCGL7u4e7er3Q3V
rOxrLh/mrKhxL3vmBvYY+Mp+OAgh1TQyKPBzh8HE7/6WOwnGk6NElDeHTBPCy08JDJmcvxkkj0pA
CjSn9q9REPQk9zszMUY5TEmN5Py4EdO93WAOda1KZASb+K3EMXwXKxKyH+OMNxEuhARsq8JZAAFV
Cdsylra1VX8i3OJiuu/3VRHUj/+Bhwt1o5HXmYN0/OQsaQVdgqyALBHWk20g0je6ARklqsDpxlpK
GBQ6Rb0DXJj4PrN9GdG26UwAhJgnKsD+lLhUuxO+mM1lAq8O3X4teH8ZytufOLNVEkFIaOta+C6L
cQCjhZUy2paiET90tzbh/wjenGqcHJo3XltNdWtCakKVtnPA7tImDw5FVm4y3KIEdN00U+8p35ej
OUSkFkKLEsvQkjVeLmo14CP/OnWo7h5RG9pyBmoo0RNkml8z68EfrbN4Yv6x5N9VaQEIt5/Uhe3T
axCLnAGewtaCnpNy0rLY3+/SL9QylDHSeFRj0/VuTs0Ig6mrA0Ck8HgtFcynXKK+4I2dneKxdS8j
4gku4q3zPzFAiYLNGeoWCIjgs7nKzAyy2RsxZgH8cwMfr+dLMalgU30yUUledqad8HTW/KhCLHGW
ji0C3HrBU3h/SsLUC3Y0oc9K5B3UJYOK1Uema/e+4W+64jHN6lTXen9SWW6bwXsQuaOBw3O8Zr8S
1NomCNcOyfcPNEw/PJS2AWBBB0hqLzebXN5jYMNNM0wHdJRHKY/9mE2iGWpBG1baNcR9PGaT+bES
jp7/USBGddPu/9Rkx8csD8CxqSzl2sk1wKiyAHyX2ZGGyE+ASebYG37/ln7RIhj3C+SK9kxSohHs
vOpI2gLrKwrjV7/vS+jK0icQA5jBVc4ynfjw+CwNJ6foTWjjgdyYDGHIcLrC7LVbWjSxXchD54nu
5SRnA2XQSwXaeU2g4CS8r3l1MEGN1axCBlstLsmVNX6bctQF4qNv7uISyr8d8RiFNO/94e2CEzbJ
NHEPPbcM75WcsbrXNGkDyX3WUosojSRRNaznnSexhDdIrnpyZ5ZJ+HnjDNsdgsKwGiFt04X7F4sT
A4G+RTnYSLIFNEpJSACNF63Pfr8ZGW5vGEw6kS9XCMcHIYWst60VZ2uS2JVsb1/ShI1UdUAort4F
ohuEl+k6tUPDV88uuz+NLglSEQo1qz3R9wRUMP209tTl3qBvNCobSKmQjwZKA0R9UqHj472rUARq
uKS+yLedJDgZMv1VOk9vbqb/AXofjju/RQYCXREFTdy85ol+cKv6ryjLzOEshaHurqr9IuT7ZCR7
hDiuf6h2MNsx8D6MHYe9dJCGK3ELH6bbwtBPDCmSUG9DjGpLuvNEMpinzlYh4dJgMwseyBGp2jMF
wMm/2BIN2uQv0jaOfT7E8oQbH0aINGOSUNqdLlbcvafhAR1/VvwLRsYp+eRWMldP8VCdNbSkFn1d
U4UKn2aZuHyUvQWYcQWP0kJ8i47pwIXANnZTUA1ydVdgv2Kk3r3zV0ZyPZyVvxVUKj6QrVQbTrzX
zyMsa0qjnGB60MdEA981PBRQpsj5QevuSXaq7c1jF47Q3ZmlbWVN8Z7UwGP/2fidwuAfxp1ahOjW
XULrww4AGFh4rPaMkuEV3n6eCGDmKrA1jGAHWkSYaspGvmjxJkRcQYVB9FqNQfZJ2gar3sew58ef
Ug79sLKN+/TlhSMftSAhC3sBrTU5R164jqvolK8PYO7kUmhCILU6uD3Cg0z0h/dM9Cgkle9x7s55
bFDu7vdvOX1AZorDRs/iyW2A7oACXcLCS9DIu7YPm0/FDxH/3/B8DVdfhGYAbhNf1rzF6Dy2xvnA
rOJ7bMjL/QqecB8BCbtvgCJQ8VnmS80DgjwVqkz4M+PyPIHYrjEqB7d2Ez+SVbuUWA0oiUDEzFpz
s7zfE+nJ+Eu1hHG+IctdU5zVmJNTZDuRMIzsiaCws/MtSo7zH7yNQ7UuguTROIpy+RLILBiHuazr
9vJB9pvu9/G+dv02IonfPM5BvqonpQfNaM47I1FVUU9QmjULBrZNxhuvkumjPCWmxa/QiURAxuC5
nptfQk2lsnrcuTAcy+Q3pi3HHwQzzH3QEDDhlfZVxpi5fUsoyCnzumSC8nXU2mvYRufzJPh6y+6X
Cpg+VQEH74Q+uy4PhWBSX7Z4WLoe/3uLDnhLJfKI4e0IjKGBbH6L6JxqIpxzmb+9qQSAtKV3Xood
1EiDramV80LFXc3xkb3IRT+PuaPzbLU85i3T7eFq4UDnMsMCNpK8YjhUEn4TEcEYGTwf4jjPd5Ea
me5PPHw9a57X53jFdH6osZn7D5J01FAJph0GMx10pT4SaREVRGph1HYrXmMtJSeQUZ44StNu+Hb6
frm28KWidlMKc3lPLP2jZ+ZvB7nfP4BiLLL+vsB/qmnr2SyM1mrm2hxjV8yM4xbdacXAh0jKsAiP
gZBIe2g9HkVO09DpLoSHP068Ob3PNujxoA9ImSd0UzC6T9G+GPlaQ+iv4wMhaCan02rKOhyuUkyT
eub4cyqlGYJ0TtGDifsbrfNpdQ/Riwq/UcRZ5Ijr3t30frBsenUkF5WfyRg00IIN7bEEoeQRfAAt
NNKJ95OXrZUCMM9JoZtKfa/X/OZV1a6wDFFd2zanJqOCAuXkM2fEGO5/K1jKT35jz73m1AtAOAvp
4zPavkQdgO6RiCg+aFrrGIaRj4m1Cj913HWCNBuCaPm0cmYKtIK9aPjPUFhV1782TGHHtKsAb7nq
uqTYlARe3E+hfR/u/+o5S5XfnT/tvZAwFK3SFvrj+AGBis7s17hSYiz0L/EbyIpZDOemTDdxyNfq
CU03PM4vvrNjlFDpEYj953hRh0eiJhk8DHy8BZDYqvYb5mnWfcGSdZHBcznFj58KYT5RkfAX/NoP
zOB87qtQcba2Fu+1Z6pUJExfMfyNIr8Vklw0/uHSlfVQTk3jPdjAd8bkCygMYTHWXTEggYbjfJ3K
KXG5X0LBvJZgtOGsV0AAc6gCMQScqaYEiuxvFGrSCUJ+gM7EyHNbDyWA0O+ljA+e63lL+KQqqurN
/WJjkRU4/BKs0HdVoHt/DMaeuxFM4BrjSA37UGMfSQf0Kqse58EYqTix3o+VxKWGghFEPySW0NSe
UTEl+POYJMosD/S6C6FaRUFHdlTGQKBKooj2rKtIf0C+BoEHYVtHBZ0VA+zJ708FhJaPA3A9SlLY
UCrDBSibcxPrqe8/yopg0Bias6tKhi5c8wNmfPOCMN2AfyUl5oBVuDvCHMBEHCXVmpa1hR8pXLbL
jnOxxXOBRPCaZFObPZLGSDHgMbDS/D+AGzHJaAcED0fwdhdAlIIRAGCyB/fuesZ1DJ7nffl7BlM6
HGVTwH85AVfjLmW4BItmk43ntzUUTSzH+dWCz/BLOBUK094KJDXHaM81XFvKndaHA/9E2BuLAOFm
1FJpaHzWVVU81OtCqy3Y4K0Ccqb/Ey/yqbmwNK3bYxLsRqnQVyu4yM6ilNVS0ihjhq+LnQL8CPol
t8YqegO/S6V1TEkkZgdN9pGXmSGKyNAwcGvBJGkSs/nmZ6k9M+HvAomKyVVMidKJyhPNBsjXD+u1
ijU5Pdf2w8eK3sW701HATBglD0QNx+JjYbOJ3xu3b/RNujKngSI/6TZ18z40212FF3VzKLRstHCm
TkjWUZB6vrZvL44yVqU+/4KfGoGqO/X2E0jn28IBFzbwH1PQ218lIPhWVUEJzyxmMsvDyTRSiwse
VuSeQWEDJgXk7Yd+I2wOV4gA6a/oX2+ASeSI7NjNmkf7zS/xN4JnGwtm/xIX65V2nh5VIE92hdpr
SjgnUBpHvvX9iGbE+8PBF38d8xwlLyMgy83SXUq8Ms9VqkWlrCGjV3Q1uOk5x93dyjW4jFGaLej6
fwj9c4KgSciibnzt9tponKQ83g3HZvM//iYOy5QGzQyTO0BthEWIjfIa6WbH9D0OdY5GxAZMfq1g
ayT4DBmlDESO+i5gUpmNCL4HneUsImbGGYi1QgQNXTVrNk7VyUkluGrTes2jj5zykmrC60xoefav
ekDexC+U3X9iPcaAjBgr2uu5s1+dEh809OKDmYFscRgsZS3zly2XnBfT3F2G7w8ksvNHnQWJqRJl
NekgJOgwRcX3yrRUPmCbqROTatr+6xzN19fmxEbakRLSpPztJ2KF/NVGc5emmi8bOTJmW0eyvqoL
C+OCgqlqn4844ErWI0aDSXfoswWcPKGJLj5QQd318T3TON2qxVpVALgsGkefRo39XgbAOzYj822p
kCUxHx5b6qjPIckbLcli2eqtneu6VTp4fe1m1JSbFt3ZvBYF6oE5qQr7lcofyxIjcXWZANPMydBt
alpYiSkWJrhMy9Ov4oR2u/4Crg/0K/2xvrcPF5T3udJTjy4xMvDzqi5qo59v0fiASPbcONDsRSSD
ozok3mVHASaoT9ZUcSeQmSSD9QkAPLLAXZcI7AYbWoxKMUZnJIqO+GhD0EzgjbgA7WS3uZeuK5AG
b6GSERc3S1vQBTB57rAQVcbhUzj/kFRaQ/ElYNR5Ih1IKKHkEO1T4vnPCQWiyc/Vo20zLRJ9pidQ
KZvlv4xSgFN1+yi4fx1ZgXxbej/BUvPzCdz9cc/SnJTtiVfrFYrdPz+E+CqNYoQolmnH90IpeS3M
LTxC0dI7sDUx/AWbMkPyLbynUi19QXJDmzcigVD0qf94NaSrseXvijL8UjClEGrNTBqRyjT0GviJ
HaPJZsTL4BY1+bwHt0Ug8CzLTzeJ6FQ3QJp7PP6CHJVMQVCI0PkNSUg9lenOan7oQfo6DcwypS9/
u6nwTMK31AHoaR0hvbfRcjVlUfbEgg2amEeAqOHOmYbxcGpo3MEQFtkqZIID225JJcF0O+6kZmTl
uj1dKzCVpqd/T4Bd0o6cSjnFBHrX8sUbY1bQ1ByESTnAw2BvXFZ/+GwO/mvEA2WzBTfjJz5Z+ytn
GOVfYjjT9Sx/W8UAyM19ctorMwUgHoT6DmTj7+Z087TSZ1ilPOwTU75ghShL/gd2nNbxZ1xEX7OH
zEdBSj1ghDF/fGBd8drQCA16qlOxLOVg9jYJuDLk2YJL363ZW85Z26htHbC1RxX4j+m07dl4md1C
FB8NV4knv0tic+VRe1ODQ1xBsIpkOVoy7LGniKmS7HakN2BBum32fGe04bd+RpnJdUWIrST3k8oM
lro0xzruAPzHqE7tSzHbrgqKmQB8+Q8xdaNyIynIsmAmPjrhfpe6z7i6srf+8ihrzcGaFWaE9hC4
1kLpb92MPZflf7MY/6CAN6IaV2gUv4Mq549ubay1ld93KPNhR2SpuFBMN7NGcX+GteIwvCT6hzll
vT1fM117q3R6Wqqmfwwtj27VCKHu7ZvABRCIVY3nvQcD4Qx089yDkjAuBAiDAE8utDGj6GFrf/k1
v3qFI97wrRSHL92Kd+03IZN3ZoEjHPSXlggbiBhNpnfcjpq2/VD57xhC4Me2QQhzEQLI199lqWoH
fOOWyBqsZOH8kJ1Ttk3YWaHwm3MGM7ValbG7ZIUD5tRaFuT9pBvVaW0Tv0kvc3LnmsOPBkYz8STH
jqdTog46hrLsAgJHf/hByOSc6M85IjB5wns04sclPDTQkI1VgC4pMy9OKnMRfggrDm/fPH77FfuH
NZ/QmHt9nE4cdJr54i9Pyowen8cDl6pHkrI5T8yUVJpjXfGFBvHRQytdJHAc6TBjLNa29f3+jEln
s2djAKEdWLAbolopz+LUJggYvKMZHdieRDb+D58zUAxN98XGy/7nIam6PF0nYdDKcBB8J8p6xN95
TixXZho42ozv7xnS6qmwp9Mr1sKT1VY7UbmfmNQ8t+qjqQCUGhJ8CCjDRyv4aKMSBKtWQSKlBjLs
Va+EBSl55NuihUU1DHCBPHZKWwiAuBFCN7EQz8idHkTXQbDQBEruOZ1GdlNIG0i3dwyNY682MPBA
ThRCRItIBXRPmR8Kxz2CCUEqRoP8FR1E8QWxtJboK95mvKlABXgQvDtUz0DAwM+0tubp4czwUnjD
+FwKf0h7Zv+J9vIwUHjlQW6lfAWtmPQfHhUqolqGMgx+Y1KFGhfzpiDQSnEm3DhPSCmeTJpQmaQ4
V32wQVAiBcdSuC94gsDtVwTaW+Mzo5aOvOyqWibUyK8WDGWR3maTKWNTifDsmB90Fy/ecuOo61PW
MlLW0gpq946G+EIQ2ZfU/fBN54qX1TQBaXnCAUm3+v+T83Z/cI7NQE5KGOrQ5doAU6y+J0VJ7M77
d6Y3gxxacseKX2XdX0FGgVLM5P0KwznsK6UN7dESbvtDVKGSDJQIZqmNJ8LwO0orGmNGjFhK/Udu
zIA8GTT/EXitHvw8owd/S8hb5w9h5AmKHdz11Kf5uIFBRvw2RJK52vMsRvyyjhpHfPmxd1nX2H4m
V3sV9U/V42qTQLm3S8jBA78RcuQKQn1H737prlYn7SCYMHVPHP6HtrMVwlEAC9tUrOhoPyGpfCPq
P9vF+ZvxuByfk4xCLrpeSZrpGzYtGEydGfK7SYu8A35IyiNBgbqJbW0zGn7KpIogagNk3I004XfB
loaze5RxMEd2/uvQnvPNmUAQU7gKaD2cNLKfheOmV0trF9GIedAf1UH66waYkMY1LIcmb16CROln
YHRBXKjINlLV7xc5wIUtrPFrRPpibWpuMz13rIwLc8wnQss+h7IqvJT0we1X2YcckcNDpzbWJsut
qjAta/vvOeLrar6BdlKhb6j4bTKJzJRFq/M+akObR0lyk4ZigNfE1QPVXjuhRe7fZn+iuFYFKUao
TBHp0VS4VGHMrBNzEOA1w6xG+XhOcA7fqB4Utfzf/KSkdD9CRgleMf8gusufE29nmay1MexsA/Op
+LpKuqh42cCHOPgcYyBIIs6RMdnM3tNwXKE6pbwMTyRPm3OlNSlCCn7dbA3mS0ch8zMh2o7FPD5N
CsAcuo1+0yHHAqhsi0o/zfpVuqCMdhPwEonmFPM+m5i5TQC8yIf27j7qoVI/MNkfXOI4goCLeRdD
jZV9xtkuclaR3Ua+H3nZeImlJRUZZ1JZ3//y9ZU8Vf6Y3efrlOiv/IIJU2pJEJc6F1rYuO1WQFHK
nYwO7mbOhQ5oHXdw0rcj4moyk2FjP8bxMbzWwhPWpQmV1k5xqRx9MHEvJiDN0MV3kffN5rHw1b78
IeGZ9oDMJGq1MEBDOpY2rs+Qjh6L5HQ7qS/PpHDOaL9GjScCVY/v+gZntiot/fInxxeziGkKnfJS
TYezy6hOCJnTRdcMUJdNw9mAE44JM6AbI1qICmTQH0cJfHbJuM9JOZ9jIqliLP7eVj0ZHfu049rz
38oJQcEp3PBmAJ8ZQ+d1i7S2UmgW3XaDIrYKN5sgqESDPAlaICEi3mVGtGHyIaeRPqG5Wde166lH
8XIcKB6LLfZgNlGzN7TDAAdhdaItKvgcBWjjIyZpbjtaQlhQ8EQ6EdWr/uQuWYtdlPZ0sid2TZwu
AE+VxGcFKhm4m5pRANHQRf9u0p8e8/xX9LloTLtNO/RxpgawPjVn1yXf6MQncy+HGwnnam5IXMNN
f4k1BZUrPM5hU9pavoZb3lRDf7V+8CKEi7TxU4mCGgRowY+MvJatErvjWMVkmJ+ME+z1ckXMytII
TDJaIHAMNb1AZFdmtXFrYpBdlccqLwSKJ30/Dfe+7IA+QunvLQQHn4ctOEVEvN4LVSumuz5pAzzF
SvVrF/7jLPOKzOxGW1Di7G45VEAY9Z4fsIWCWCz9Mt4yKhvTxwXkk8SIaObnjqqdWh+MAvV4euWj
9co2gVhARpDzZ6CmXfHxm6wi+ghkFk6XO5YvVAIJzL3ZdWOjNdw834LQ4UBnSdh4EY+EQrLu5pnc
6BRSDVFmfS1QYteLwgqjXh9orSNWgsnDIIlG3neeB/RX5C5xwKGe7G9fhBfKimO2F4g5YzQOrHtd
JParCx8rPvzgIXa2+JSeSP4fte6OgVBBtbwgaOq1RJ1u9ObK5Cp6Z71QdsUBN0SHLp0thzGuvv4j
YOLxx17zn7Ytnw7xKwSmds6+K97YL9OQQnqJXpNGyUkgnxoPykp69wsYqaIeRfjXLMcY+vQ8PIv5
8yXFfCKwpKG4JOhs/VrAfdPsE29CUAk+RVufF724LsRLBH+3Es3wsEuEBARgLOfW7MeBGvRiiNJI
rBhA2xHUnehILrjZin2uRgHxtCtspCz5OHNtz183dxt83p05SE6cPFInYfbnzsFLOQylwLJMEkl1
KaO8NgMFKSGANnvg+Inz8GuXq4kBTLLRZ0Ba9afqKkrFeqo0rlsG8l0Qxyx/mh0DZjfkzT2hO0R0
UgVK0++do2EsShdZXu/AR85tkH+krowwdcOOMNzvjciyyEqOIqpHFE/Yy2BL4yvza+9Wh/hoUv98
A96EsHr4sF2rQbHV4EtYNycKuYHVSG6UziH8Osz1eGJNxMVipoIw0Y64AuqQRZDjMD/1Kc8xEAGr
O8KsLPKPF9llb2toLqkNBvUOJeX2FZyyevi1pU+y7t1f4sBeB8UcWJfWjmM/7fRenLkMXQencear
N0H2r7KK9T0nqGRkYk2o9/audz+XAuYwyrFHf3L8OhOcL2HigdMFTndYLOMZh7hqrR67lAX+cmo8
c+V8G9j5SV0urfjRQ7fR5wMsAPQMxXzT1r3SX6YzhZ4GI2xIb37wTJPd2WUv/R7bjt10icaVHqvO
XiKuGTdIiI9AK7e1c1UYWpD5GzK69Z2pCr2gcHvJeTKPxALUzZ1IDgGCIgyEbPfK//d8eZA12WwL
U9MrWALG1BxeYbZpqY7gcOxnVwoTLlw7alm5jBKwOkm+nGi83tahM2ngd0iED1PamkPzIiDdEoh8
LRbi0N20xAGUjt5tQkCqrX6Il47g15LugvEWIfeFeA4kgse2n8l0/wjgba7eKFZB2HzCfspO+XTA
tYzg3b5elnyd1bsgjmnOr5jEXRzho7CfoGn/en3M5RgM1cMD1S/Vkaf3+RrZSNRvfCz4DRUQ1afF
vs4rd8JIket/tdhWGNvgkS02pgQ1Dqug97N5heQfgSByuSqA0vbMlB2oqWfs+55DlDVKwqdpi/D6
NoZlEIrok84K+NLJ+xT7GtVO7mqoWfabMwiHjEcHIDMxVVNSbJe/u4XTFrLxYHmv6/sNOw+P84o9
mKLqf5gEZdA2RupYtDRR928rDSzZV13vyC4XNTZeyylMU0/Ntc2Lb7mvOMNAOeqT2GB7dmtmdH4A
DnVj8Msrns/3qDoCz7HRljvEmuAxcKae4MuS4tKWBf7UJLC2fbIxUJtFoHWf98wOwJ37KweDw6p+
A/WVin/+W4sEtHl0cCd/h25sTmz26kC/oWXiClqs+vf+Yi+jIkclOpnjPNsEb5laOEGJ+jcRwljD
ecBeUBkMEMYxJMhmD2hxzSsqVDoq6mBOFfW5ECOA2jkfUlM5CvM6k7Ok3OTS25l3RXGfX16fNYWc
QiEEFK2t1cFw2nhKHWjVEuXS11YEyfSrc0FFo/ncbl6hxrKwBJnWGPmHavr+554HrcYrbWRGfi0T
ASdZbUYuk11DTkbAS2aizkH8YhMIMFSMaaAvD4fNN5KspAOrRjyrrrdTr7h+XO+g3+Kr7aI7kkHm
D5nfFIMR3wcv+W2dpt/6kOmRVRZ51jvshNLhdOQRoKC61RkDYRwSf6gquJbuvi/BPC1rzQCgQqx2
1Y9geB3DK4eRcQilvUGvid5F/WM68Fnidh+GBPIBh/70qqeXxT4b12wG2q7SWG83uL2nqsVqmPDX
wI079ey1LKinLIcZcv9iqfFBaQ2Dz4+gHAy6EofsyrzrOX3qeKsTQ4nowq3S1zAODcK/Olu0GRyN
vBzDeL4aZKXYUpMOSRpgX4YMB5ZxRzL9OxCdYAJQbQ4oZwe5C1jwoCNYClTYKWQHpS9Az0i1AhaH
s2wLh29X7jCdhv3t6zxiHxMfph4zcpwR6YUI0TYYXrEAThSldhLk1mTVUBDkquCM1aNTRVink29a
WnW3JKmJGcM/cLQXBJXvDfF5Kf/xQHeit5OQwXO4yomGYEQNUxIg0U9ji20tMw8uP7ABvQ4/9tV4
zIHpiiJxqntrsUJvrZrsr9Vqfr+kOatbg8T5WEBeld1qas7+uzEmcBPA1xWK8ORg2Qy1veXptGw5
gvtOo5FpIElg4iX+x6UAzYXN7dyPyCPvwSzerf7Iy58VL0y8NBtQzFXPZ84I2tYk6QqcvSmbtT8L
szS5aZTy172DS8epsv+WckEs/Db5v51LEIwQgh/TB5uQDZqOOf/z+gLaC3xDl/mcuUewcc+yMgFY
qN+StL7aSuGUA1H1hXVwemZTqmHf4i7wJAsGOcLMchTsGvFHEIXslC+en3skW9QiaPJcg8YpxL4z
WyIx5fq+Ebr1zsPhMmcY5dI3mXOgrDIlgS33cVI2xGUCoHPyMtJbEeBsSJasuL2rQyUkbFs8TTF1
hRNIrlbanjm7SZTjpat9UUIRIAKzNj7tr64qSakI4rxCczZK5qddBBtjg+D8C1N4lJuK8Fl/URZz
43YWlVbNMIB0OOC+wxoZYvxI2lqFeghf7QiUbO34eueB2ShkaQ22cSvRyygbwC4pJEBAkZlxtYp8
GrBAwxzcz/4NVKew5cxrvvHQKaEeHTByqYPcArLv193aSRZEznchctq0yd5x9vuBgYSis/xCt0Sb
fmihHILc0VY7RMlpQDzeM4Ea5Cpxm8XpomKX39EyklpFyxl72NIjVVwExtWTYao2iT0sUwTJcoBb
ztEHLx0QCIKW5hm2jGfYw0wDbEuANG6SUuEsT9D1p7zN2tKRZihoIpxBGOMJ9vQShtZHpiAnKDTC
WB1aJGa4SQm6PC78OOASaQjpZS8rc06PNKew7flqkYQKH+qJdDr/QtGALVHe0bS+x05u4l9Ans3f
vdGkwpHUieEaNcrVHiDPxqaLkN6jZ94fZF4qKOqQu2g3Zmnry8kg65luGtWtvPV+dZvp0RRKKM2L
1OTqM33xTA5q8O6aNpOd1+Dygsr4fwWq1vHm7Pr6OSyIfoK6sD/KFbKzqew/MOpXXFCEWMuXXIDe
VwwIsOfn40L2ZK7jkO7gVD22osJFHSsmFvBrylXoQN/NXpSLVrT7XYHujQ21YKboX8WHmKs75Z7V
OO5Gc2O82/+9NHXUMpMhWeMEjRZudO3dfUArkJcHKC6ue/H7U2m46ltehxbUrs9AKE/XPkhhPiDM
SmXQasAPGoG6hafHihipY0FbF7X5gVv62PPPDiu8c7U1E11ahZr3e17D2K6QSHL4xZwezr5Scr9r
GaOSGS6l4JoYcJXULlPjpwDPex7Ffr9auOKMYUKI4A4+/FLt5/nAtIfWD2zh16SmXUzHSnGpmWin
GSllGM1VCDTXL+KHGDvL3S1yBnlDTdilB+VCfnXffdkXhGVNCC0OfKDYVmB2MfWb8t3KcNpbYAFc
XAqcU9TJx2nXlF3qKrYyolVpfpi7HnXDiPs0IxlOg1B/XfjKp+lgzEMO6QmHLGrHAW79fwHtvZ5U
srEJCJ7cB7jQUZn65QsTl/3rGTsP/lzU9qCtZjCyjx0sSVJ5/PdG55VjYL3LkrVXeIsYLrUHPhWI
mVp6amcUugqilRPcQcFvaSYl6GOTZX1dg215kMLyyBGRydz982QXoIrvOcsOhmJeGVCuzmhlpGnM
hc6rH5TPRdwhn1uER69WQAVlgoRzGSH6a1l7RK/I+dQLLQYJkCn2Bdfe1pjBwG1/LLJjhMw2UKIX
5JdEuiSlgdGlW4yD8a4+DA0uy3RQ+Rm7IlzM0aZcAOuKz3VnXfbufdDKo1FkfLStUKgOigGJnxMC
jCIza54zYQeD1rCKuRCdb0GfClz5KqYG1i6dNFCk9TGMP5p0rWod8lQL070d4uBBHa2ODDT0aDDu
ukcwPc0oVxQCU6etdtY53ICW7KwdBW1hOaUDgVi0+ZzjAPLj8ZG7deGV0UcynbQUSKlIUhfuwkCs
E66ICoap5j4NZVxJ+zP7VSYIYaZg9Jw20/kios3eCRBNThHQSpbZKXF9MiwTwLXmZGNihzEJCWrp
KwoiFcw+FQWRCV0LyWroYNSsI+MSLdkf1iC6Y4Q8UwIqBInAcHbcLks2ScOGsq7SsywJ0WFNFfgc
rktzMujREw0UN6PMvvnBWH937QIjxbHyALZmI5L35YPXxIcCSay2An5ON+ULRk+lW9MddxbJd/Kw
EP85S3NVcOlHEEC2w8ZTIb4s0frEP4eNFXIh/94WF+g0BUhS00c4hiVQdsV1ybMUupw4xVpfiThG
zMPze1dQSYF4+Wafrxsd33WOtPS/gEnwR3GWn0hP6jxSKqm7P16oWAdqo+Ryf0IAkJg7/TdFfEh5
5bFmTbaZUKaoMioNI736qHHFTxm+JblZ6WpBvA0DswcJzHxYDDIE510yfcAfD94TmywqP8LpGIS0
oMHVLepLVndrp65ae1cC6MrwB96k1errBv+UlPCHP+Xae/b/DYKa/5IjVxB4uoS5tVLEmKpLY6em
eRI0ptpKhwI6Dy4zN1+OoeBO1+7a22SyIDf1XUVJ50MDFx63eMN22KVEkuqomt9kdv1mgpfCwG5g
klGn1JHl4Wv4g6yjNxQdfYllMM7CUSoDUavaX3wzFp8CgVjyvYDVYEZ9kZDWsnDpOu+i9GPR2mu/
MsB293Xb9iFcYifjIbdd3EkzeAYRi9ftr9WWc6RcKAcP2m4z2Vf0/hDDoY/RefD2E0u72YbgAdB2
aIVitZ85TfSTXNjVfkLyH/1lLh1cdn6ZPqSa2uTWodE2iE4/64TCixEESecE7qWhdw6Lu8/oYKas
4tPT7OdAcrlZGdQZw92KK5kRhSZRLffPIMksskrEXs5rYo/iVgRUhdHu+JCUmb6VVffDI1nWIqAB
q9avCB+bGGZVeJx9drUWIACpXRSgLOhmFxiw3NcoEspBgSGQoxwb4KhQTUrth/N4b95u0g9x9mfg
dXLWtErvMZHoZpWhToWM4040cgvwqCIhCj6dJfVXhEvIiamR7cr0UpGrdredah5uYJzLx5gDJmeB
3iXFK44YJ959N4XCbY8DIRcyPLAQZDM2kwlPmgw6E+q8xEcHrkDanDwq/4Fwbc3Hl98RBMJW0Bli
PNyUL1j5Q/BX2I3G3WCwFd1q4zY+ngEL54p76L5v1pwXEMTmUOjByjcAISiwwjhRMG0cPSYlrmLU
c8+zOtQtiE2nFaTCTOokFGv3R/CBzJJFJyMrSdtCJA5LkxivfV8RaS5zhPtkxL2A6e9me+v46D/H
GZ5YF9jQHHTWjWs1X2unqF72olbFdvgMkDHWM6zLE8L8OMyd6bR7cpKV9gqTFP8lWI1hRCJ5D7r1
r4POLJhK7jowWYyBSkmnI2+TuWIc8Prc9Qh10jpMA1Jus8Ku3jZKy5XtVLB8RRkKNz4svgE/m+2n
ciWmlDQczR9RwNZzIMwMVRxEzFdz3MK+aAMAsto/zhVlY0Pwk3q3KSI2axD/Cn2N1671rCZGVpq7
ns6Atl/pmZFG7/1fe+RnicX08i4iCd7KdeIGrN6F0f0A0MZ6VxShSrdUTpgSrQlXvkZ2EuJolTRO
D8rxlYlvh7cgC50+FvF0FOqGjIDMv8mV2/mKxrpW+WdWIQxqrkBVWg3lUEFlLGvr/KQI9gJlJujK
9GI1qVmqmQjWoiMoOrlrs7tDP2UuP6HWgVwX1b9Y2A/1sEpl9mvw+PMI7V9dIcMIw81bZvQjM8XE
t94afKPX2ztko7/okz48pMwGxjHnMEEBX/Jb0F+oUiZebnZ3OEq/P85Cgy6R3PNaohTgaTIpy/11
+uCIAFjGYc3jw98coJ1teeRgBYy5ae60vd6TEOEfBXuhp+auIdlx78i8Ntp0RmNWgy7hAvZX4BJY
1N/aXo7UJkFUyNu0UxIkv3INbHhODHAFEl2fpCLzmqZFyX348DPeaXsAXizzyf3J0A/hXE/opgpr
VUjoBwUrIbapmHuEuGwMxktYR1Am7/1sO+z6CHinYO8WrRFQ2hf2LFEUgvryutlw92n65crWKpQ1
HqyUUZ3T9Tx42SGGnR5TX62+OYkmlqe8pt15q5MD2bl/KdHSv72jce6dwQ00RXG6ALAuw0B+F2LA
vzrtiNnR+PIcrGMExPBRXPuDKtX/XRPolVQn5jA8aW7pbHF/DmF32WcwW6DzxXNgzOCB5RZI4CmR
mNvpQwC7zIwZZ6pjAj4T/l93Nq8fyXxr/2R8+cTJX43KjjfEEo2CdX7RyrlmgVx9qSv2OmZi9d3J
qdWNoUdcRErjIMnKEon+VHm1hVYl34YPnjffdr5zSMCbsGZQiyR8sbZf/6Z8Jrpqc1KFKD1b/xlS
h51wR3M1D8pp6Jiknjp5S67QqV6qSIMfU/fVlTS3RsHkePpUHAMd/+bOXr1leJfe2FkYyMnuinI4
cfy/7fk0B7gMVDMW9nFJ9/RivJqA0GUi8FVm34LlGxzgJDNsssNdkdV58DczvgVwzWMTc3SsVCmL
JRn6Pv945Ng0wulYDVvNo8rvtFHypzD/DVXARGOsyBenE30pipwzyAdbm3u12CgyGRwCp+msM2x8
MHfL5axKK5qhYf34aofMT07MV8fQZkdXjV4s2/2JJBtB8qFsevI/AWJDrx258QCzTMCp0+1f3B/6
KpZ2BrKWq8tE6FXkAMbhXFnCGmc78URVCPImjQ+UFOoZLcuQkdDzSjJMVLHaYRm48MtdjamZ/57M
7DlRE02Db7y2yoHr+5u83l9AhVVNPUwc4/jm5A3uj1a221bYxPgHeRuZK3fE4ReROW8H7pX5bnPF
KSy3Kx/Pr7zz+VhfTs2QwMgLJflqA2bU9JOWCBZ/MAE8O5mtXuO/lwGWNFiu/7j0vzpA9GMDsUt0
+3AxUi0fNbwzRE2c2JwQvi2vdqyOaxTmMJuHsl0qEdqOuwXdQYF+vWKxoK1qNp05DwKo6YmyYWRp
rd7iOKwkcx+tf63ncK+14VR/3hmKk3q2MUUfX+beF6ULu8SotDCf4s6TH2/b4E1i0Wcg8XOu9aFi
vqeCKvUO6KiFquBs6q3pCkz33ikzV7n4sqHKmdqBr/jO1/IxR3uvgZQhQxudJabzpbyfljlt+/i/
wVO+wmYL2ID43krFHDswogg/0j26IMOX+r+g/HKCBveRxdOn9x7ts7yI16HZW6vkXeKd3CSxPzjd
FulPIF6ofrna1xkeLmaXzOEW94TWVUJE0KCetXBpdo2FEEZzSu+TaFcDmGMv3ia1WxPiYyqSQgm5
P9sSQLvg/jjLEfTa72otSayvnriaJDPQau9DZydBI77ktAFmtTBo8OXruxQSgZz7x6U7ulbBtzy2
LRUn5b8vm4GBLGfYsmLwqJ7EV8C90RexYjDtu81eJqb66zI2hXbeHHifQho6fgxf2AKbc1cwjawk
ltz2UfFsgn4IxLfaFYQbPm0kZHnPef9c15VElYWdIZ0PBAf4B2hnahmvj9rB7jRO+MjRAi4Cugng
vInnhYGItZKgCZLnA9Lc7nhnhs64EahIf/ERbmSYByJRHOhgG0JV2seR5K9ARV5mYBBD6ljLjEAt
A/7P1fcdSrVe/8KM8Kk71aZegCLuweug1WevdXOCgRS60Gd4BmvyIL9uwOWPL1d+aylJB1B9Fzrh
I0Fz7NxHhstLdjKkmim3kfEecpqF4ycyXONk0EFtq4eocJQbzs1/keS06RD/dj8o6N2ITmvKC4UA
m2Mg0Cj5yxPPS4WuE9fWHY9fCLgpxkjAPfvAg6uTt4U+XXG7VemjfHpCsG3E/L858KLlwtQzRwQ3
nIKLPXE6Sbj/mKp4muqfNni9NUmipLSGQGVk4TbSpHOM+SxHX/vmX1TxiZ2/NgyzayIhvMonyXrC
0V8Um+v4tRAhhqmawmI+PJNMqUA6hqXaEDZXSsoK2mxZFE1J1WTZQ4K32S/ycIowrKoWlyot8Uik
1suA97mSHLzT5vkNLyFYFtE5iKpWqr/dh3fQUpO6vBNBNFVmu052VFg2zlpC7as+433U/G+ezwZX
S60wF+1HooK9r7Hqm/aiJW1rmMLp2w5Rm+byJStrCMegZoUpByPyFCZQNcCQiclsql5KZDGzttR9
TvDgAnYK6qpijV2yE6Ptx33kNyiuUzTtE4bQTSiIvPJ8NGCgASsPrw6iigZopuFI73312yYwjhee
9Kdz4OYTbGZWplhzbYp+36V7bn7SxXxMk4p6nFcs21joQ2bNeQVwRzSAUwrA213+79WR8LHIsrTt
HMLxCtBHDKmH+itG8pA9kZ88fWxhExcvZlpCAcQb3Lf1mU1KZL/skZ7kGriPkin2fuLjLJdbL/g8
IDMiWXpV/P6Bx0IYEr3zxbKgkoCpBoP7vFOQ7LNuL5Oy6hGp6dr6Plo8AmbZ9IA1F8624zmI5OBa
M4vqykpPIhb7qLgh9HnXmgMwNTtSHPhWH9TdS26mwu6TcQ4PpLarK0r8jvxQM0HjBQGs4vXMP+Xo
bZMeGVkHskQZACDMsMQRXPZLaJz5C0/JdS36ywF4UbiiyuTJW6mMrBo6IOv0gNItqWroNyTWIewL
fnmI9YRwl9k4SNWhD9Gst1+m0q8/7c30AZAipoVDu992Ttc+2cYiqnsMJqcH+oEzKjPkmrALEcXa
D6Yyy65sPnyXiXEGtXNWrOvfB38VeQ2BRUhwdMRnCxf9IU2wqO5tXi/o3cyrxulLjiG4exYmLR7d
ICy9sI6MHH6MHqhHxdiHn8k9p7v2yjWk/E2i+EgumE32a4301SPmQLjtezSzWUJrWwjLGExP2F/H
KI+roDVHxt2wf/nbf57WUy+7KJQFedVaGm/Tgpcxwkn5ZLW07/l6b95lRVpw6dtKMQDOMqEk3MWS
Jjku1X8Cz0L7MQ+SOpStsVa9nOzdZ9B3fAuVA8CPVcgi0SHureEPfI2kcqKkJB1TqUq0ZdE/5w+u
Mg16nCH35GUGUSZIVafwvPwpqsUfedYoZSncg62UYmGlEJVPwqBb2ThPBrlcm7HdBk4NEYKjU2+O
hKH2TmwwerQfgzjOYStUwJboQMn8s5GWVglyiGFXX9JCVAL43JxTgMXxr/Qps9l5nVkj0u1pSZjP
Cbpf2D4DCxxz66zHCUFMCUSRUqzWIXb7MNGfDaGWfzk7HARb/khHcpuBKCzbzQrzF8qiM2kt0vpI
4Typ9Ul7FzaETufx4YzY0rIhrSd45FGI9VxdM/Nd02SFRuDwN8pkjACHIuDHIXVmz2wNC5wWPCKM
klNSgsXyfl3NOUFE+NQhbSARN35R3wPvIJ2sxd4hTPvX9xRZJSi3fsp7mlIGzSFLfnPmqbPO8dv6
kk4drjJiAqZMFlCETcdbDCUDTt01RE3WLAkyFEqo2bdpJfa7v1dpzS5HqAc7dW1WxVFwwjH9dAxv
VbP6JYtwQhejsru9L5fSIcxN4RKMtwA7iaPjjLMai+SHhBroa/l/m6335V2RQSwCrnDNMBA2DaUd
U2jeo37rPX8g/oqxl4b9cJ1aI0Wm9bQ/wp1vN1jDcHqQd4jLXWvkBw79XCr+EwMFlHToe5E3zUkf
lqgKozalaG1yVrf4tlr/JIT6bPgi98QpbinFIordGlT+R4PVOE2Jhz8glve2ouswaKbACh03mWRi
WWevik7T0eFngQuLgRsP2op+tYExQL/BXIqOjFQDERsCEl7tPuyYOguar733/q7tJAUZnbHkXxPa
zn1tE+9Mi8gMmvQDXg0GV7NpiFJvZLX3L0n51nhm9ivV/dVGCXitt9NaBKZB/uYxnysozxae/4kI
yw/fknPdztvAolLZ5xQQGQQ0V2+OHhk8yslUf5+TD01udrBS+1atxztLh8HKIEbAC4+ZkPJXhsks
8atj9dAKtUovwWU2UyvHIptTzTHkmv9k5yVBT9z0hkWfOkfMwRr94BUkHly1kHZnqV5S8CSQjnr8
KUHoK8/XlmqkKZ6SWDk7txvgAQ9qWJFC1s4RI8v+ygbKLx6bFVp11wLM9rbRvaJle2+x9n6KUS6D
FvTjNwesjjgGFFLnIMf4nfScOVs7eGY1oFjH76zNIcLLvrkFJM6OAsW9WBcQN/bT3aReQ2OzBeQX
tcnk5Cozq4ZCApvHt0Hi2/bsecWrzkWOblOHf+67mBHB+OvADLDZbz+I3zv8+RhU1XUSO+3xnkV6
uYmHs3LyJ8EmrFSZVbk3Dfq1bfEbNTSEGOZlP79ZlASguZVcEaL39Gvshi7hmIOgKZSaNxUfrC55
ce4Olx0A/yKZFccOKgkTaImHiHfnRoyyqFMrDFRUntyvo4aSKUeMN9aH2t52EFkgxOOfhyWOl1X7
wxY776TBBblE8FkJk6ML+6xy5nO0DXvhEBzR+4/hlZu2uTVjcKnZcxMpTVGkmd2Z5evUyvCFFQew
3gNcsiElCT/BQ6dDu/S74hiuuAGQ1xcC60i0QJqaVWzYwa34vE8d8EH/Fwe2/mh64BnL4gZ12AfG
/Yvw3NWx1ti+AkKapmSHp2L5Qn6xbg+CK9+Ds2O3urI7DJ86BlTSsedMxAosXElL7tEHhc9EA8Ez
j7+FKvRIO/PJyr5ZdH3qfokYn/0qKkzWgSP3uzunPNDHlVVMeBplyw6oTgTHfEOoBtOasPJbOZe8
anF+NaQS69iHPqXkpVDs+gG6eOFIg+I5XhoziS9wBsmK6NGe9TkOSXXZJYN8neJDWOXZwqJ/n83+
5BRWv0vfqq54bBXPNAu1edATXLPxXV/5cq/YG3H04Tsus0OtWO0wHD6p0bLglgp6+rjyNaF+sG17
9QPH4UPS1+zqHdyqShGsuOmHPcymrkpkF+TTiPFK1jhzAfTE92INvikfDmkZz3Utc7X75MpRVGgj
sCcTodjgtuPUK/ATIqLxLN8tLk+Z1JfDZtHzP69ZUnARn+dGxp6cIRegkSI1geIC8Gn2tifUE4Mg
Jfmrd4kEa/U6LwBAWejQzJxm+7h90gJLNBQmJmMUNkqj1RBnCc/glk1HAFfLYC3mQfsbicOBoABN
tzmlidcRvsnvIhQ1mYQBhDQOq6mAwyQ9469Y5FTqB0xleKgnfvEP+BLXhcDzXA9OUBeeHfv6op/U
x6tljXumhlD7DxaoNaNmhwiUSjNHsXQskqLemdlQCe9J5aJE/T9Bcha366YRpWFm1hg8NRxbjfOl
NtO1/yodo/EpXt4MTRV1EWVU82wPDiSisD3mvXHizT33znUknnFEpAVN6VFq7qhiVvlIoSws9ASh
nSw9t0acCycmhRG4ukmk4RD23xZ0sstXIvOpnTT/Hjlc4wsY91sWalC+Grz0qlbOF7kjyOOdyuOH
rNp4u/yY1KXsDXGVH8Pfv6+/QxvWe0bzcusyyju3gwVa/4qXLEbLNsqm0JroeLg6naibPullsQms
MWH6++rEjWdPFNdRspZ7ZTAAiMYjeIzn31SUyRq3PwRsZ09mgnyo37iZbSV6tKUel6YuFwQfxgbQ
v5hvtS+j0iQqylUUbQoQWhgb+8uSaY974jAQbt6BBB9+rbWCCpezZSWdqdGDU4jexWVtG/oAOXjF
GbWoi/QM/JGgaiydVAweweMmo+2N/OBkpY3zuw+W8MQB4urd7hk7Dqf1RJtRg0LXTy2nOkNGMTTq
Rteda26XZuTxzsjkuzGsT8pHMEJlpe2MrMWRl4OqphpAGnAfHCie3SUGUFGgfC6vVzWywYgvZPUf
/zQjJtI6Ism4+G/EsZeiPSt4/zy6I4Z3lDAAp1sFUGa3nXCoFBIse6pzYkuue+GW1oUS5iTfd5KM
UoN2ej3ZffYklgsHrUMKdjzNNqI0HeujzIQEM3ad7k/Trk5banMgw3BLlArMaWjaNcVg1yiEhmyK
D2TpHEuIbtAJJBJLYpZfPF2lgB56ZPd/WMdtslfp937imAlApyljKIFCoh5EqYKjGYopqU1HtD0v
DvPwpB8tEPpgykDKZAZfUgxsklhAi+mQjBHk8XJ0AoFUSsXm64/8hW+Fz2hnfWLKJipdAt4lGAIP
36Q0QisdJmdhLjOEJYKGt5HYXUGszT2ZWNDW5rXYs9PlaUNp5b+k4m610eROT48UA1yXQvyJ8Ty2
Thyn8Bt2fzlOul+0QVpupxibx5tSU7+iOa7kUK3ptPQG7O18AxCXhJdys3l20cgnTY7GZlp9amQ2
23HX1VSVb0ySXSb9vDTcow+140LL6EYTMvTSZFKfN+0LNUMgVr6hQ7vFcPJyRAqKgMzV/AIeV36i
a/Sq6FuksgX2gyWg3TTbmqDNoqbYwXV9IDKHLSuFjr/kcwSKmdjDFRD9M9+FJrKGb5oh912Hab6a
AaZWGIlqJGisPeb405q/8TBlPf+mPOr4AHPonOIHUsuoQvO3SlNtrdO8q7T9kKyi+2MvsNSDO1yR
I5cyTAI1qs9FMFDqVuN98goo1uosi/oAtNHhnxLg1+irEcsHSt26GMSk08GTHu/f720QVcHvSVfS
KsTavRDiYgsusOGVNK7SNs5iLKAAsLr0FR+LYuIo62w2zqIKXipqa4dcdTauENQ86ZgUySoJjz+t
JpXfZGhyOT09HkKxZL5gK9FiItrNjqb+tLsOLaCFB2MplpBupCOz/U8MFO6jfUmr8S8u12zrpdDE
KtPnltYyDIm9/2L+yB4gJf6Vnl4sxzDEiJe0iIr5AupYQi0qkKf5egeuRZ8J5N8/J1qWHPYiNLXt
+KHrazHvfyDctNLbb2SV7BV1QbilBxT0eIevKjgLIaGkEcDRCgMZQbT+Mv3FxZTb9+WyqCnawLx+
+LG+rKifbKBDWGgYwyGQFmAXVpn0GqieZMSCV1xA3qDyMvWR5ych2R2AYjFb7nF6a/3hk+jvWscK
g50P0uch5eG/XXuBHSydPiNQchMt2emrdl9BlsizHhJN4QWmcB4rSPko4N97ESryz6R/a6XTuyEh
oETP/Xj/4kfwxW9GksEORdcELufSUatyft+AyzcQwG1h6EeJBV5WmIfUxKrXA0ur2x1w0HF7bV7P
9TwX9gKEPfKw+Dp2MJy4XKuHJotP/3yA0NqYR83N/GtVjmW8gamPt2j0PgZYaluFWWGlzcW/m5Ms
m4pUFjhEr2WMMVtbs4xXLzmTiD1iY+8jA3a+EuusE+3YRl31AbyIOhOxcpH3e31eotoaQB94pyqk
x7Hxdv1XPLZj9zyj9NfQErI/ZuKWXr9jYtXp1XGYy4IFCSIBG4XizkIZNGgUrNA/bspi5QELsdJ0
NuqWBi3UYBfGeHlEhchwLB++sd9NYAQiYxfX7a3CU9L6TjCNQgwj8HCkM+Vt90VcQjILETryLCmy
71HS0fIQ0hoTEKslriu6IX6frLL0gwuV2IFwVYTmUfd6BCAWFqYgVFXoHuMp/BzfZi5w9exlQSr1
yEcIdaZaj1hbErluMM1PNmqnhh/COZHqYDwB5PU9W4T71SEA6HE7FavUTVK2Nhu98HCntb/nEcF1
Ml4KwdvN/Cf55R+7QXnyXstxiDreXYdZGJWCNx/Snkwtci/wZj6QMgK/5WVj5pIZ62eOYlgz7dwu
tv4BI2FZkbtpOSfDrxRE9gn4Jn+HCgmZemaa1fnuY4nKzJu660Jps2Mku+mrhzutDLjCEiFXbjTe
c0Dlgfbf5sAe80O/ATr63COvcBwTTRmVylkSvNDAqhZ7InxstmWA2RQbC458JALjZxUzdrYQh3tR
o/rLtLP8XVyGkTxtzxYrhsdNNN2HEywS3yxP28qr7ht9N6OPMI88F4JXR9u25lkaA1Sj/Hh7znVN
7+QtgRIoU0VKWTU/amFdjLxX7pbZ2y4RxZnWamzpIITQUIFYdaRs++cOd1+rK00Ko5kPGrReOcyM
CeSzlu+COaxcmv17GN3O9qOKH+pWOB3HhjqwENcM0BEJgb6ZlBlwtXbKTfiRreRAL+5awYcc1R8Y
hyHgX1KcZgMqWzhagjG5RtOnZzYg6TnwbyUGhhM+BBn/WmXLFvOMMaDaPRTkCbBt9mXea2Q4PzE7
fJ4hI1iFCf0OVj7ELCRcyNHsqTdNtqn9Sioy+JfmOklR2kUVbG87fVqib9yFTn3xN5G3ePScuLNH
ga9HiRIKQiqMi7eScgwYGCs2lZAlZqmZOXhnBmsYH0upbUecTkxkGptuR43t/60llsCpkUlTKLdX
TsCN5WJV3zKChpPMA4+f43v02nIvJt6ovGlA72TOfTALmEdSKRycHv98S0NHqNkY1jkPqMM77LsS
yhPww7k8Qx7YJR0sEW39qS8xoxGoxcJI9Cy8negsYxLTgaxyX51/rnEJ9OEwjLbxMnFvvVTRfb1s
ktaz5nUK/hPJ7lqXk1HO9+6oAX59dyEOvXgOzuNNj+Ab5RNTDorHGuC7L+Jh04WdU8XOUAbvW0Qk
vU+RrJ811OTAKReqYENX+YOGY586g5UiKtNh1Yjc4UeY6/b5lxZ3pMG72aCMaUephJG7lNrdRHIM
30KMyUPLPdpXKiwGNpSdjo/FRN6hzEIidx+t0a4/OWC4gINbNraRVqSc8qtxRJTw/kiCRgw/c8rf
Ahrj4fGfXH/ygogOQA17nHHKZxTUzZm9H3P1b2xB/czbFmGhA2ZNDNWupgH8XABECIL+vl72RsIY
2kB+yKo4ehSGIXjPLlJztrHhkQY8vSfzmC8aeUJq/EFkk24HfR3+DMxfT43EJI5xYCzfUnQ7jvxx
/HR41fqinoG7v1ddsK6DtKiTVsnRLkcqeGWBbrTACgcWF+T7IowLiSkEw3ALa1wMgTvhUsdZG23s
RpYfS/wH76G/b9doJH8SJUtN0wRxOeDwWk3pPuMd/7BGGfDxrDmNzjpuevkPN4aK+HWiFUqyCxck
t/k2HT/Zj/X784Ro1aqBTfD2u+Phkc4r1Mqagajztvq9TzZO/qHLCW2JVTNi373GgSXKEG0atAPf
CfARftcV2dhlGsXrZNzt4RyUzyPfxdiZEZz5+IcMpJcF2rigg+3DhZk9G1NnvvhBwhJ9q5EhFlGi
YcqlUnNTk3tSCBmoM9bH5Z33WHj10zEnZJY62kLCHd34euN3yRpCcSpy0R1T1w/asZYrjuqp68+a
rFO74tKhCdVGinhtvU3TQ4GmMfGUrXpdMlKi8bjdEDFUuLHVtMD3I1ZNEwnUkeKp4UM1QYY9gogO
D62So1ymgzF7tAoTaNf9R7UP0sE3hVi0aep4qRCdw6ovrI+KF2D/WJAyI8rmSbR1OW023oe8hrLh
swhihioqrYIqbBhSHSaoVnqD0N8KFz6BXyurTfz7Lki4cUh4JC9O7mNKu8CzI+g8+VPZ9kTDJXf/
GBARqjyAdMKjYVg95EDKnhinF+DTXqAVbL7Mbhsbkt6bzCTuXxfIkryaLG+jzVQoMAqETYkBk9Ib
BaAwOybfDsUUXNUGRGLrsmMABjyuLD2JZyD2fIYW36Vj+zGKPEwDPAOs32XDprp1WLaoztOvR+aJ
dOKPsZtgvIIdrRxEfT5eZaPOCleEWlbBVsbVGORiCMJDPtg4Rnp6jfvYdgQgr2mHfsFKB2AnXRZT
0Jz7+odVsbJG1Q7Db5lMgg2oua2yuHdvTQ/ojKZqueqIMPWFshPWj6NUhUWe0P0/8uRN7LnC9EkQ
ksbMNbw+6jSSSV2QDl3APKOoAB+wVL3pCoJj/edLl9/1a9XqCSqb+cReiWhX1Rh9I8/Y7BKa/j1I
l5b8H5Hl7T/RRabLg8nfzxmfbGrWn7qDwi8kHAC2SwHf+BqwkhpXIeVH3n0ebAUXU5LtQeuk/bE8
e7fnbkR9VolZGEIfMf/JqmLKJJHpQzDVTkGs+nUB8D/V4v186Lt8bWBtHnf7aB2tn1MDfmNdmW8f
gMziehdkTGxxVwlNWajNNhe71WQLhXEUedmKoSSwAZks5mN2xc91aw5JAXtnf7pL2nzflhzdZpc2
mAQ6JaEfxk0Q96482ab5thUjsNy9+S428UfILVGDrltv5MPMsKFf0CHvohm2sliuFMd4xIBI0g1N
E90uJaeRmU9kGYhr8wwAm/oGDuVhgw9Nj8nduIRq6+77m2QY4GMHErbiihepcAsXo5ADtT1ZVIpm
ZXiKsj3bbQPc2rwzEbBnSXOTJAo0/T/4LpU4wNaWANY9+nj8j/k68E4acSqK2f8c/IS1YySUzU1d
clAOMsCr8Fk7QVrA6/Ux+FM9EnCnbzkBH6cUMQgebavSZmb8YoD7kZJBDqMrAnrwusugACIgAgdK
T72bJjQkQYt3R0Ke8nEKC1yCeAq7DodzFI9Fanh5m1ju41DKcq/sN7lVnb3+ucLcViuk6uEREgFV
f8LoksX76iC4xl8KxBooFRoscETP49FBJUwFSAtmDTGgbreLJQf6EySLcADV0rUS9e+hP7/9Lckd
w8JRn5nzErona+0wqNB/PKeMH/2msSvga9jde9vG76hKg0S0UJTDOeMdZmp8DEvIyQ1wzQAzi72F
jcRZUvt9z0B7I/hL/axF6ex3NOtx3PI5YLE503L1Ptkopp7uftNbhxWzGw5ZDAUzGL2P2Q8K0+Dl
i0KUfMXlwBhwnuPQ5FoH+7w/cqEpTWdxc/zDZ181HXvUqs/JiLHdtQzcIbv7Fn7AS/SKqJw8R3Iu
pf15DhLiqgg2joHoR0afUwXcrtwI9N55ZoqDFFFypKJqFsmvmx5YIhE+RnpIbHz2WuzQDx+7Uirv
rpDAOaJyCVSjbtFkML5T2CYQWb8xQn0WjJTKvEXsblq67+wDF8Q6fJYQD8OBdiGQfq4egff3xehX
HSiEo00/w+QC9Gks/ujJiZqTHX4+2W8bkS7FbYqrKRLV9SUZa1c5dIwPdFMKE1uRxhdkd0hfk8Qq
FifScnSgosHO3p6ifD16v6XtMaJWzlom2AL+jJYX74ToFZ4rQYUW15UQ3D6wVRbTYJhkkkgFEJNP
EQ0HNOEpCh1bEdIKgzBYsSJOU8GQ81ZXejX193gDneyrf4rX6FnohwiDUm6/0PlbnzM9D50VkII0
8ztihtb7AaglT7/LSQKxblPs7HIuTfpeQuj//KXL04GJswInWFitwK32I3y6y8glGCAvzQFVWFy2
YkIzi0F5gZM0Ll5qYB4KCeVo1zUhqe6dz1I7zmzWGTQ3Fsi12VwG/NI0cS+Xx8aOPIZ5LvCJRvqO
9MoMMIoc+C8rN6luBTdMjxsSwGFfK13glpuj3UhdflvTe867+hJfwDyG/onK4YhivbsMzg9A8MJp
qPXDhiVlWnlHXP4lwW+XLF16dOyW0SlqEX0XsbK4NJ/K8Ef+NYtHEyUspqkLgN8SplEHwRPIPc36
GI4zwIepsLDF/gAVkyoHvcKdOWSM8uTxpNH6ZetktdjixyYEo+3ehcGhmkexFR+So9QIpvP8+BBx
aBn7x7D2Jo+aGTHcyN5ntn2SZweIThxLQGt5xLkGFXt5IjfRtX+nFt8KuSUyU1hL9MXkmwBDkqUG
DLSe8TTaGq6MaovubuJZ3xmCLDkFP1SKMq6qFHMeu8tfOcjAh9QkzlKfDaAnfVZCOxfsGrb+8SiY
diSVdX2/05Xj7GBjIhz5Nz+4S0RpqpW3pdS8BUbjiS0YvqI5dD1+e67TzB3dQCU293RijUY42/Wh
f/i4EOwJZ7rSMitW9aFoJjWdKOHciqTxFAGPB1CtRa9CNY+a9Ghil6M+7bqcesZ9pqGqKQyaSqh5
V9PMpSpf4ihO6BK1bmmBTbi1IO5plOxU6ATjpeV3qOChZ2a8M9K4tagbuKDrKuFCwcufs4O0+Kgb
zYxO8BGEYLP1pfHmgxClpEO3wSY07tlmKR89Jx3OhYZbGASKHLQpGr+dm4H6DDqEDbIEQq5Govsn
yw8frNn5VfHaCoQ01Zu3pYzraJ/uT0MTncJZIVD4MtAYKwEzNyDEc9X/7mgo7ZsHjvtsEmTmXawi
tNHPol+6XLQX1KArRR5UzESCCuSGrT/kRIAuJmHrCH73ZByX6GjcaVrxWr37wlhRwyrxYJGzeKLk
k3/rNNFRVQN0Dssa2rnjVnvPO7iTsKnd1H5+Pju1+Me7gla6j4v9q9wpY1qTPpK+fFLii3w2T/We
RseTUaExbcY8Ru8iQKHDevXZbtOt7E2M7BeIUV2SOlIcbl09ke18nkUeUFJai9EmjSbXVk6RqEbN
PrVNGuyPkfu2KS9Cps8keik7LZ1LhT7tBbJ0UYJgSph8cbJCbxAM4DRNJbHuSXvwp8WQQhmSahsy
WCFFD87fR5cbXVlmKy6It9OzOf5kQSDFzhxH7OPZnH3roRpp8THbpiMvsMXxvVPQJeqrVzNovEBB
MgaX5NXUV3WSKO4XoLqMwMMcaF9RLNbdpQT15CEWyWn3GjdRfvk0zi2kwSmaAeGWQyxTqH+H3Hol
KCcrFIm10R2WfbcG3fnQ6yTwstSg4LAMZi9s49or2nheJewp4/5IhPgFx3Bu9+HtlzImWn5PoSeX
sxFhHsV6YkpwQcH+UG2JIyWEaD9N+19tZEX+F2t7ac+NXZLJF9GmVqEr0DdOM8PSLftbMonkEh+Q
0DIQg69C8V5fT8AOboT8NXiow0w/x8LUrIY3gMUS3ZRVC+UcZlcPplDvkly0GkWdZ7lSYHroCdbq
I4hrNQrqKzD3taoyaK/8aGXbEGLUhMesLXPHlwU8/BgBSQekFTAiP32tRMeZxKg905nPfp0641ge
jwQHNMSl2bobvAi1mvLGVFK8HcwizR5wECOweP8202hG779LSU6ZVEOX7wsFIcdESRTKi7m9WN1H
ngnqsn2NMiJ0zLpvBw9UmGFshld99McfRvnognbi7W5OKnZySwwQ/fKP7nGpHrnFvRlvE+DYS4Wp
E2SVd0VI/TjmBPT2xkXQc2JjUCqw78Cbne5LU2zh10bJZSFNCxFHMdKkVj2D1rxCI3BjtNdyWsuK
EioPpUSFqoDH9CC5YuDwi/inAJLtOpQ883Fh+iV8UWJyIqkoWbFD3mpQmBlDacGBrcIaIXvjWv+Y
/XDYPpklYKMzo/u/TA2eORPMJe0CGbYGFSLBIP4V5W/ydDIQmmNfDJN7HVCe6U6FBneU4mjIBAiP
pCl7RqACXUQlin104hqukDwz/xOey81FBtagKJuVPBqHe7BLqyPM5HKa26mhsQPNhnzQJa0tnlLR
NvvpL4hpxz71+6wWhIcJR1BH4hh0rAbET553I/AEN7gPHzjE0HtkQO5Ep6OshEyqSVXOY8wxwDh5
E4jnVdhqu+0eDGqRS/cr+/tMwZnT3gb8GhblKoxSdjIa0++yDjPjOe+q9SCgX3NN2oYuk6mnaVBv
evWIelDVrNs3Lhqv8U9npXU88qPy6IxiA53vY8hZKq0IDjEngYeVIlP0rRr48WUhCUCD3G1uOWGQ
OqwpSnRi7cXgdLMDIrGhC7F/4KbtjpXqvYBCnqSdhA2FbVJf0ACbudB1QI7vF2yT7dsw/kzM7T98
XEHIwqGmx/vOSiE0cbG9uYGpMaDJZBp2csheMN0qeS4CwoAzQhxll9JT7x5IL9axdaz+MYe2g+hp
zelKTcskeCqs+7IwJaaZOe48nKGNjnr1LBqxXf3K25zvFZGXUDnjqfYOOkA1khhvCMY+83xJTn+e
uJkzX4rc+yyupziks66CB82Q8gB28pY+on1fGQGtjf4Adti4pFTo4aLWFbTfFdVS+i/1sfYZXXcm
xU9+BEX6TI0oj6fvS8GFhwvNCjni7TXWeuUmsKBzpxG5WE1lIr+gu8S7rx8NB7tNT/p9CDPD7DlC
ucUhhPFqiGmN9yXmGViYYEJRoXzysCPogbQtja9i4sF8FxSGFwx1QB+COSSJXYHarqF/TnRtPc6I
hcW4rtFF8FfpVgWsGStXhNGkO/dNq5jyit8BGpHNFqT3l6ap15cTUvB+LLVcoYh9gSV+W0NigHCG
dP35E1LtCZUgYPwPLx37Bep63Lgk2k1Euc0Mn3pqj4vVGedZYRUudTUewH34fMVZe8hppHxHth3R
noWPvZOkEeinoq4Q+GCiYApssQ3OjdrdpQx4PLzh5qOz7SpWmvzKGVIaEgeYk1yKHRtxMxlQUjGL
li0J8gN0yc8aO9HRC+QAhSwuQHHLSs5OeWJa0W2KBeP8sMnKXi34QOlZCuxjlUG0uCKfViZpcRGL
WLFyLc68ZfT6N+4Vhd4uAFuien3xcO5hlDzvz+Jwu8zAweww1x17LUdiLSr9LyXcZXhSTaSNWmbI
gHxIOD9LC8yPMCbjRsGVgaMagisSoredXCa29lmXFcPHRDajvh1ir+MhM3lFjvXHgybVE4wxOXLn
eQ5dgM3zZ9ziSincPFJQoufLsrqm5cqX/TiQTD/ftHRUOq4IadYYmd6KocmjTMwfkLXlukGRMNKE
LLYOO2fd04ZaDXRDb3tZwAbS9k1jTJp1IM0yrZMdA6+W0rOhr88K1eGM7yXGjTCmHFpwhB66/4HG
Q6XFp4W9sc4XxAMZAZ2xl8PXcEDxfRuhG6HfhFNkgbowxcXJijc53PIlrQWfzJctqZctkgOfKIlP
vohYXyhYirw76C5nSMu/vZvoejetzR28mqeRuFhyzTPcSup8N5FUkbN9+uXIgAulJO/Ry7GTf2Vd
uVWctKdS40b4AgeLnlQtJtBXrH0Fr2ioE4pPav3L6kYYJ0C1PA8fm6iurBQ7nEOO8PhmH99ylfCu
FjykEU24GioWF7m8Q1lp/Y2zw/J+TxD9pXLRGKy6izRerJwxJ4HHwu2t1OETxk1WckK2en18VaZe
GL4rx3Q80K2p9ydY1coGMbVGVuYASFZsJbElwQ/FeTmLsSleJqEAkWK4vsuV3yS1ZijJ8uV2G27Q
G/8HKA7PeFZtpQKHej5nmxeRzIwksf1rxOcHAPn5rNx5jr17OR+PJMKrPiMrbW0ambZNFx5wPGIB
+kNGPAQ0OxR/I8AUfq+a9YFRaR5XhB7u0VrZz66w0UfUmfXjEVrD84S19OLkm34GbUCUOIBZtjfq
xJdCcFTUIpkEbOGcDPG5PoaavOMgirvRHGnIR/1h5gnp+A5MRtlTRAD6nQa4rJZVFpXWPSe09L7N
UHU0Azf/gKite0zlRSUZFHRRrmhfbzXKvkykrzjs4dhpqSvAP8aVe9e9lu8Yuao9wf4IgXoddiIQ
v55cXaY5kSjiAo1uTNlyAVO48GgaASDkUhmC+9A2WjH8Bd3kdBTTyDxjV7Psi7yYSkSjr+GAS1IA
KLINbRnXGioW0Eiv/LMO1lQdBC8YawQBi9yLx1OPh+qk5sqG3jk1klJHSg0Rv3ujRpBLIfd/LtTp
SqiUTniMCwLMzIz8sHFEUcaiQFteoWpkz37CEL65vwkVd12yI5QDm1lSKh2wF2TY8fJMUFj37eVJ
QZzR5Ab/34v5Fvm2CqS8sVQy4pFMHGPJX7w7Y2OCltsAnoZ811LyEOUs0T1pa9gqMxkEgwXBGSpc
7x67FbyvMwsMrUfObVwERpL9w6g/KIoLWHuMREU/PkuweLeScyy2c6ZyLkVbMUx9c8mlhGM2dSGT
prD8tZTzDPXhwmPhqGS9IzDc0cFyMdY0Hn1m/mlr3bY+nd74+gpvy+qLXn3KRnXHWFE+yuyHnuFc
JLNoaswBgXV6oTAwlAo2pC9y6iVI1wN/8+v1nWWfZ0Pv+CgSzDGL0eFGImvhZlWYoIVO0A7gb3uf
NI2P1h4pd6vxWFROxB1LJwMGN6jWbK0YW9Z19h2EleGDUuBpcu7XQc1GbEEGP9MiN39TIz3MY9a3
66EM6sYrgf86v8IQSz2FXy500LOwNjROajOk88Mhrzd8phLJyWcJFcOVAEPclsRP/QiWC7jD7f7i
GAmQVdgsxik2DtCJPjkhMiRxnyTA2VMNmXYj9oqx7QE6YJVpqNkImy52oAJQ4gnqdKDJm5bMSyCr
ABKsIEb/u4UlFxLaE6WU+0nXnFZAlBa1Av+0Uw/dN/B//76AeC3qAYg47h94Rj9nxk2OYlBhzfwE
mmP9UQPCsL1WTTe51G3BmIIBlb521rBtr0WklHmP1nUsmeHx70tZlmuCbmcttT8yUNGs0VSETt0+
x6zLPbCfA195RJmKNCTm+XOfwZTUptREhEYE+D+54YS66oKTPG6lGC6qeEaVRUbp8PaWhdXHJhDO
viAax0A3KHdIIJAuzucrTL1+eugvzOhNlyV2bol8PGHATvVAOova0ulSQVI0Wq5WdTf7UNGcIgI3
wG9nrieYcdvPZfgZxYbgblZkBvZQWYyK92Vmz7rPpcCB63sS4DOjcBLIL+LS0bPq07ZQ73CTLAK5
XbkymJK8jJ12irvsc0IR4PsbeJqHZJPXROlvk7agcyPzgNbZRfdrGHrECN8fGVHa5edZs7f7Zg2R
+JXDWFi9/IHGSjqNGlfuRD93BwBaoDqWhn8kCziOsEubbsc9owR3eGSotmRkqAI0SCQXS6mP+Pcc
XehN7k8s3D7UCURBTM6hM6TeTL6gqFWlRkZ7csFTXiyieahjrw74jv047cRxETUJknE0zIS8tilD
0LZRf45j2g/Ca+7O2WDRyOKAazD8nz2xPpe3bI/bDZ8HjoB+NwK3OHGQzpOr37k9nGX/00/Qz9Y/
wia4ylVic4tSIcyw1gpdKOAzCvhwMOuYwSTW5xLhBvxVqafGN24ryrm/gro9AWGb8UzoWpI4yS1V
9I/nLLmUF4oS6ExJ7S891UmJGtEr8j7cAUHcTRhCA1A6SwaTxNdDZPpaNWSl5f+B63kevVcGt74M
xe1WZALaMYDp9rs7UZA3B412Xl7oUJJnoXg6s+3HkiZT2QpJ6B3LXS+rLsG1kpJr3vcFnyPNFP8/
LDVkwANpKPgvjIF2iMd6LbqLTpO1/1T5DDEzIHeoxBnmwSp0Qz4W6Vbi8wHSpdsEQnsrm6NqJxrQ
VgRVIbwJTQguhEzkU9MnfddrLYiHVl4qft+TailHwUTs5yxT+vtuxGrHEJHlxNI6FdjctL7tSTaB
346Xeokr8m8LLmkjkW4hGTw54/0OsTRMtLvY3xPy2BEZQPvDls9I6Xmylm1GUbTzO1CHaTgYgl6O
n/aNCoLSgVygWiugZHaK+Q58mFUQnOz3a2R67vI1zdEebQSc7ubbNER8JsgX1sWRjyCjIWY2npEr
7nF5q28V05RXphVAGMOtSznpcBDH3BuGDGJDi2PgcubDakMWrdcZ394A/otBaFZhPnTdCJ0Gb1ik
9LhJQXh4VSyrHqe5H1ydISX1VeoUno4pLRkHjRtPnyKluWMadPboleZ6FpZHAbv1yNX6VfzH2po9
dDtSqsxW3QR8OV37mYNLgy3BmylgzfdeFEozSTZR4hTT1BegBKtoVykWx0CODTHLYARIKtkHPp0c
/1ZFFa9/YrMuNg5GDBiLjCswxFmiaLn+aa3JFsHCbULITfYfeUUA2Br5wIKRwsHnMJyZiIDS7iV7
6qxJrnZIUa76v3xD8pHicGbc7gZ0am/XLH/Fc470EBwE0skX3u+S9wymljHgNGbG2TmIMJP8iWFc
8GIgCQG9dPWPaW4kmHPzwACQlowFr1zvBd2pi/6xsPdC4TgJuzw12a2YMBNsB99MXpI7l2pGI6ns
xPYE9+7Z5YjCsqBqeQOG7Q+rBc5qcx0gcW/rhNx4jiW237memDmFOoy5LT71aVnlrxGzVXzTtY/3
hL5fGiwZXZvdusUP+d4thDul6mpSOt8vsB7mht/Zo6hny9dYrecGJ1RlQ4jzqzHloCPdtFpdHIuE
sJdZNGc2MNxqkjSpm90G2MOgMZFydOYPZRzKrgYhxawp5S+ecrd7i88be/7/pVgRmZ3dGeCgaV/9
M/+WWR0LXSlkRNwX53Ay0P07zzAwHv1nrDYDwIshg6CL5ko6vpoD3JOt0VJlMUgLYhPAGX7A6atr
0pfDud9bq7uRKvZWHpqb4BT71J2iCjk1r68tp5qxLy4mZ3Y4N7zy8fzHQXQSRSJmFrEICQYPIv/e
+5bQq9IAKrd3c7XJm5Jec1SCV6mAeKW0GRtD8dI/LqQiN1Pj/GsblxGyimxhDOKFaXuzQx+YXbKs
KNCtMo6z+Rr6XBjBD3KTJrRRvTcDh2oC1FAQs1MJ6fNsw8fkjI3rjFlAdYot6Bipd96URxaOzX4O
uOy83/31CKeHNDxWuiVkgoQkVg/bJVwmn8MK1wWidcXCTlBgQhn8LLAcVkl+8dZ/xqo2F7PxAkYu
BnFGrMdFCw5OL6deTdfNFxvtcU6kuUxg8whA6nKW1BfUh5oD/pUFOt3tE1JzLGkx2beIVIBKVqsy
/b8dCbuV6f43TlGuDvWjRbSR353WUq7B9me0vNWemzfneovraMGZt5ufaTo6VNM5SWx7yQTBhsD0
pCiG8pEXgL6lbgKxShF9cUei4M/T/NcbTegzKVWQdQqQ9t/IchcSiZUG4rq27TA0pvV0Qm1L6SXB
3W2yzwbl1I3bj5mAo/KVWa6dHj2hTVABCqCaDFsj1qjnY5BBXm4pu7gpByNBrLwIrGCfdrQNd9c8
ooy4KfqB+2uGsKrmaGzOwP8TUtfaMkgTipqM1OpUPyeMoBiuI6wmQihDDtVmYkVTzfOP9i3AsQVo
yUvMqTF2PuAINNNZzu+k02axYnMY+iWsFX1KFep3yQFJnSDKTLQ7eu75zLUptsuYJjUEe9k7mpyL
waI2Cmbtj1ojvyj8LrGFbeGWXPYSKUISiswisv/EqKbXl7LUIfBKk5OLgp8x4OqqSCpuj9QrgtT/
1pN6Cuofa5dxS4iAFKSDJgnHVhRCAM5R7KDwlyYqSNikFn0xZ3JsmZEy+NU5A38VMag91/WIaEmJ
eY6ZvHTJN65WQ0m7X5sB0PDv+SsZQTjPkx/AQ0C3zCgb9pvME4qU7zV0sXzdodpVN9ew6gfjJuyM
WXpUwww2Z2WZ5Scp/Tjvns6fA8WgWSKYWhNMCu6QVPoVMvAacMot64MgRY3247A0yQQPIAP7YRQW
/g3g7cQOjEmLUvvJrLpdOSV/TYVK5EL9OiDmnbWJlilRA8+gc/RWLckQNcQJykkv/8apYiGSAKHn
vd1kZOpv1WihMGGUFA2E4Gw+ZFwgGtdsix3fwlkGnjuI3WdNz/TaFTh8ssDAFPkODxV3BvzCy/Op
vKikfg9qbArgxhwkUlRXUwp00evqj6I6cDMV/wUCyx9BNtjRb3Vqs1iEnOnjt99xtcGYXOSfZuyc
U8LeLlIopJBvIKhk0HOaFFSCG/oY3GwWX3wpful8oQz4g7vn2iAJewYMOM386UMbjIBjjZpDqULq
rTlDaMnDjB0j+eMEK+AhzSJeodx+InMq3vmfCnOOAkZuLkx88CKdo3rr8E04EAgzdKzhqru1osHB
SRZzvymAHkilJzx/UmrlSxVFZhumaLGmP6x8YqZ229YBKrscR2+n5boZJ2ePJGu+hkBVGc0/rdmN
Kd7j9tv8XLW9lQOcLWO9WYhGPVB1J0Hv0Z1UnrZ28/p2YrcLlJOnd8m++Wfx2V0crrIOPYBXuz1u
oXat/dwocbxrWZle2hksUx5LtbjO3pTnljUF0aZCMF4WH6bmiyAnU9mblhVxZy8HerhBWY05LogF
D0XnUu3acSBAOQ0vPY5TIr0/3FJVxSdFBHu9lGmOgDu9uh+VOF7eN4mR3KIaEnjgXKHdq90LbiEV
uaFBtYK6csLW6CI1vmvp/m2Qy/80rRhsLj+s/BUsmHWm5LYbBp27K/cqjI/EE025v+R46MQ7pvZ5
fFhNuTLYgGfV9afjV14YqB7f6eJS+7WVUx6+UZLNW/P7em76okpdUZy9/RnLdpB4SsVm4f3dL6Bp
U0l4W5o4PUNIgeSACNb3mKnz0aaHpA96xKnLsMDkLHti85fz0a5R4nXaNWnhuCdAC4DOyJ5Sx3Vc
4pZWchAcgv94EQFYKHgj0YqoU8imex8ELC1Im3XHky/00tcfzrswP4oa2Z0v6u/kZcQMZ61c0ej4
0GHAV83F6qRblmOT8D+yrD+3mZhBcYPQvF7Up3yDM9imos9PawrfWdP6ROXUTOFdsVBcbtdc6pX3
2Cn9OAujStgU8WRON43UvJ7cghBh4IYW0Ze3tRug0I1j7995Gdp/3d/NQP1BaIar6zsPcTit42/n
ZSQN6xer+QSCxLLIct9e3GBGo2W5FQl6cblS9hocpPNn9flM6LPHxIZUOcGDZ8EPW3JsKTLMyAlG
ryxq8JxmfGDrN+vVnLn1ysNhpTPvyaqwic2366VDIDtO+1B0VrnTjzW+CtdbnDd8BimtEepcDlzW
AOyNEE6cf7DYL3P+PTAQ4lxFGBz98DNKuI2tRtzk8iFgYbwDQcBBANk0ZstbBMN1sJfRXUPSqTPS
bEectgkAZZxILC9jX4FaZE3BJczr9KzXSBcAgZ16O13420NPuD510ooVJNfunJrOnJp3PBTLqeHX
ByiFvMa1UONdd2k71QwHPgz2VqFU5gkpb0k6iXkJloYBmxWjnl07ajtukM01Yt9M0FOxBaZiY0gv
tGLXtg6IIKjGklPYffu2CpwojdYv+wq3VWUiD1Dd76hdmt2resuKNEuDT2jxeaHT39nmHjLvwxF7
CVw/CYYNjfc+tFiCpBXUDkB5j1LgVKLxKVk7nk/pgasKihMvToAQcdus6jOuKVmlEd79nQ9XhXJ9
ADiWA1Tv8XQb39+tS2oh5RXXAUuOFaHsPSXkL6jOtrFkgJaSDzFwYSTu0DmYvt81UvVPmT0Z5wMK
ieRmBeY1Q8ARwAW/JUW6DhZXglKzmhZ1WoKP0xkINTte5Cm+YJERqyToqFcIBffgOo8s0CIgCMNM
acCPk0rvhGHAiuVrbPmB2mYBdXqw2I0eBc+DR6ARRMpZz+bzlfpiXBBCF8X5ThDnNX7szAiy94Rm
3EYVpuNbCG/0+MCfHMsd0ODLuDjCiu7CWmQON6cuftUlpK8aWEAXDqda8wEZA41GPplzkRi4Yux7
0TmYN6YOdvF25t73ftMAdidvRGcX/5OCULrODjeN8PAhP3RD+AltnrB7IuP8WyhAPk09Uj3eXJlN
RWoL9p3s2RjIsHj2gb2NQxjU/Iqva1VpzZxGcnikU0D6m2+vfzxAuAh7sFBsLbb1AjbRaE3dA1UL
dmcrifPNyW0t8LOBjZ11IyF6JfIC1MsV4+7m+S1BlEsVS7vO/GGS5ic5zAvyo0ztFWQ8R54B18Pk
CELqkr5qYo01wXM+LQBrIU/3XxtnumDxrx4LPEbUm1xTv1fD+tnOirAgaKMSChFoFws5PkisCvlv
C3xTU31xBikSqmrJ27O+hDZwUofrnc+tuRjXjMJXiE7GD/s5d525eEIRjj7IuRkbpJN/eacRxP65
4urFjsBwwUroaiZRwSsFJL2TPZGBzHCNfv2hcReCxQNI7v87O8xHVpqopWx0+RCiWqI7PE1hYd5m
fEz8W5lXcvlp4aKNPrOMvF9WLhU6p7EZjy8SVTcRHp570r1gieqBMJRH7ZqcuLO70W0DYgvxa4QT
EOcX22X9J1CVrTweb0dRtvKdlIvFYanomU5wxuFdsOxr1OIRT7wJgPWAAFnhobLr//3CpHee15By
mL5lQk4ZqPmuUdtlF6qHM0Gzp7V2zlwxL0rxa8TRrGaZlQGQL01wVDaFogzJYYLpX/TbdGa2MF7F
rEQkMPE6/fRVWh0YqQT98M0dXnyFxY5RiPYjgZMHiuZrGx0/TkG6hFdpXt1+h7h4kFII7tIzmWw2
kLSU3hrwWnS3XiIND3xquAigD4F/cSWvDSPN5A3XcK0qbC9WLG3EY5ZU/bgrHTGPZYugM5R+dBRP
0yTODcLk9eNL0mXeg6QprVXqSJT1HzCd1QDjpKwdVV+BRs5gVED83pHukvU/rgN2KS011SBrE6CM
d4UdqPmMvv+Px+1j6VMssxs5BJQQ6nX2wQvXwmIGZQT4AtduZLO2a4qbu2EwtnfSJ6DZmSEQcgnA
wCiQsAqGwo73jS7Lb6jn94GQy5xaxEfHBGZfkEKYNJ28bxXWF5TFJbP0pogXds21+sMg3QU7Pc3I
LSOATaeFEeQzALfMB8+lnFa++8cBik0Wlg04caHjsg20K/bfRg2sH3sBeCk0YPoStnfBnrIxYrUN
mvAxgGPdMMCYhS1EGE0d50LYhiGAjyx8NMdUF+jJMp9JvZ3YEtJvIV0FW2n+fnUv6m3eJaUPv5xH
uFZZNwx1ZuKsvCGZQK8Rbr3evEPGc001R1/24jJ0ePvFefVIUzqpzfJoCWviYyqC/RaKG62wmxUP
iG9KLFsoAUzy35JYrKhVZSAAnVHb4Ck6BEaOAdl0eXmNeJwV1RGQVo7J1QnufvWTIFmxa0K4uDDQ
rzSSGtL7EzeN7dZ7Qlxi/qrFWaPITEOSYqhvBKHufE6VWeXhUIhiITgEKI6QlYT/DlFpYN6xu2TG
XpkkaQ3U5fbWntspG94OVNsYDtrCZtLt61ODEfcjANMRa1M27tdr1h+B5PY3+W8dpXig7ziBsMq/
0rxeIJ8Zqk4sjc6myPnNPtsjl5xIAmup9V3Le3x3bS0HwW+TSDWSsnwKyv4OGHjvfXMuAsc99WlQ
axNzUI5nzm5luXJWmrCmtD3433AutI4aW7aNhGEn99kF3vPVnzjdjT8D/k5v/UsqiIyu7KvAJLZU
JJxukt6uXNO+UhrTBUqxwcIUo2kxgPNnbCtatKaeMyJ8u5JOs6hkjb6HP279UL8I9n5RvQxozwXa
QC211fzz33UJMWSTcB7JQz0e7GgcAr9l3vk2O/7inmkJpeduJMBLJqulUY2FTeLogjInnrfyA6BA
MynkQjUWw8E2pRtr83hMdMhENXSHXBazH1pw1C4x2E9Wms4naLXxjfk4OlX5LJZCMU9Pk8ran5s8
kZIbu2iB6WlFk6hI3wBeJLrvJ28W3nQ8hC236xS6nGKBjEnSBW3Zw54yj189roT/nhf0PnZYnOaz
FMHAMXypQb4vaVylbRicpV2PrpC9rdhVtzpzQ66WEynn6Yw/jl/YFqw3BtbFvrSuTdmpmT5qKpQn
awKciJdZjI295BZb8rX1VZtVpJM6ezp3fP1M4o1+twvUd461QQQ74+TJx5Rw97LQe2NCnVVGMocR
PP9QYmApV37aEibh48UJWdlwDQI8FWhmZqlb7hMT3p0a8DIYbUsOr6bFy3I2BKMsgsPeIAWhd8Gb
dOKZHl5hqfugTZm0g61SIZPzBxLExAvIZso8k/IvEzOY0kObCcfl2smquCj6VWtrukt+vv12ZggE
4fs2Gaaw8ZHboaVOtlhulzObxrqIy3fMajfLzQNhfh3Xw/Yew0O225w1Cj1mOW7YabrLZqbq5qsu
WWrow0MlHwZBFgkEj335WcFIhtkgJVzQPzZJHAY5TvCDBVIwuQDbPaGSnE5UOiVBfCp/DHnbPdN4
RlzzmK5z00+68K+5KSGSTjPZ6cUho62GnJS28JgWv1b9FrVtMfFxuOtaB0avgVbqTT82Qcali5Ot
xjww+M+HmGSbbwiPgkvbNe3PTenM3XoGzpPXXSBadCk5NAJK7BLlrxdXEotu0QWM+HRjVq3RFTKb
sYh+SwX7oc/X6OrRipbXSdAtxZ1fB0rlr38kgOw6+TZSmhpGz6QDgin3UcjpJ4c7MI39dkaoUM0Q
xHqA+BZwIIkMNHt7yrz6g3hDTaEGym+ir19Od/sJY9L3HzDzmlcK4DzK8n0W3KI5yJ+WoCHmGAYa
98PG+8aW7D2AmXGlBFfNtkoZR8CgREGFlge82Q2Eh/ZPl+9b3jhL9k2NHa0OB+fNlrj7fleGMycW
sMh6Xy6hKJuBa7jmplZ8KyQGdeKuC5gXgHQFdOgzqBI7H7kbnLfv9QQbmXKeWyAmFBkd7AZsj96/
V39YZTZ26OP9NDeGIRfZijElL//z7P5t92ED2Pp5ZGJSxFOx2hsWRXV2LzseGTNbiaxLdi6KgQME
IYafYG/S6qTOoHKqNxQbZnjFKTmTpZ4T5KZvr3h0uMxrH/KHX//ghZT1d0js2tOPojZuYVtM4vFH
nPQ8dNyRzx0Lm06tseDqPGLaMALfEoGlWj73Q+A+f3ZhGsJAacYe8a0nClw6KGMtYQeUKI/rWwh1
6Wx5py11+HmWPAKd7IYux+18ZcArM8C4DrV+PIyZeabeBaXy8dPOwGpT9iN7ChsKZ/Y7r0chMaB5
On0EQ/q2NXj+IFaGbxVlb6kddQCzspX57XTc+bHwIiRcgrxfNvpqcKEAUH46NnHRtI+V0lgMlvBZ
RfIQBP+8XKOrUPTrLY9n0JENSdVyN249vHPciTkJa8H5krJ/ek2GKmlXezsgXnyxjcs+5JucPFql
D1CRD7fMnSY7BSbcf8Zy8JoutGS0rzPHo9KGmtRHk8cItDN3DFtW7MeTeii5m0SIMxJtkX4OTRbO
/KO2QvMCEn3i28Ie3cID9QWtmnd8Ct3RSGXxbQ2n+WfgV+H1/RJSncgZT5ziS00QlEmvGAY0ramB
a9BWdJx77yiuB7C9touLBblrBF6uHTYQFm9LNSGcVkFAjLfLxK9sJWkinqzQGSN0R2kbFjGc+aGn
eUbEYltbaipezsbMpasj5O7qRHIFLzsvu73R4bStwcil/LXlWzp0yv/WBjp8gYeBs/YcIVh0IBIO
5O3c3a5DSycO13xYDFNrCppGLefZyw4irrXjX2y4P7fiixfDHg8aSufMskg4X/OjgDv5VAFeSPVp
8yrgIl2HFK1bczYEvlG+LLzcQLKAzlH0kQc4Teo3Iq7h6qf48L1lV/q6N5bIwyIciPWAFtfNjwN2
i+kyjHSVVGqvmlrUiSyRdPZRAyCT3023Y0LRRzZqKb1w1HZJSEw73xS8IXTz60E0wmhGwXv54BWL
zHD2UIXzmScZq3gjQVFI2D/G2qkggInouEhxOiNXcKEb01+oiDNuzr3EklTss3E3pZsJFWxXoT2N
DBa7ImSBY1ohL9mUOm8LPmBMORbSsxGQpiFQWH2F2B8Xe6/Uffj9ph1FhJpdYPHN0oEJucTpQUCf
rEZTFbA1KKsrrUNkWpR9A8BnwhUlVvRELxuJlZVJj7bZMKy+ujv/PMXykh2Vfbw+c8/0w6el6ZD8
jLFPKAevMMUeFywH6rT+nN1i4AYQg1YWtQq5dZS3TzT+BhJHpj/296+1yqdkRdx8/XnPc4srouYI
FnYLXlEy7W+VK4ZLaWYv1X05IjGUVUWDNBxvdlzzlWarEvg/2eRosxdQTatC9GZ3uu1n+IgFR/7p
NUIk/nT+oWvjVPE7XlFLR7Pa9NZc0Z/+05GpX01i+O6TrBCZVstv40jOPhJRt29hFA/3IH9E7DU2
LhGg0Lvoq06xxJmaYpZeYNIDlVLCclH3rO+qEyWyqT/kBgXGH1SRhA06BQHW1uK/6E3YfPMoTId1
CAiEMB8qc5quf2L8xGrL7t78YwT45ewG+Y8CyMCImdnHR2VMH2giK/obJC03HdS8BmRMre3r8xMY
p1b3A8lUCpVYdxnWwh/hH6wuGifVD4Dtr8u3yGeqJ+5u32NDZ/vXePiYmUFLb9qfE5j+okpOkNLY
slqjOq+qpeMHqZ95Cqhsv/XGHdj3XdKnCUjjTvR8WD68aFr/KSF7DEp8RdHn8UIvuO4AzLo2YwOb
rc1Z8Cy+b5fmbgjITJDiz/xF4ex88HJTbVe13n0BdlHeoQ0vWwIStFTl4jCe4nBErqpxQJ+AAiDd
dzuVcedgCSN2X9+qSEuL3mvoKVxZCCLJWxlEJNe+DeqC7a249OWJRAPVLGcJnn4cNe9na2lDYSP0
fzsp2kwrTJ1V8N7eMq46pCrVz/qg7ClcHDw+8eqP0a9w7AWgaaKBRgO0/tIlJENaLDSoaD0SV1t1
/hH4NwBFju6oiwD+mPzRTmMY5KUNzh45qYhMLUM/gpKCloqZAeteSTulbYgGoLsHBNzyV6k1zRLs
8GvKZsh94HALeVw0e2+mBmhKGRkG2tIztr/CgjCljP0qxkBMqTAD6xAIjB+FFnJExM96AbyXQfSV
WMkS7iJEumv4aSTzj8xRObrICKcoYZ9xtoDfFJgTjBRxKdqOnNcsUj29SJTxbEUGl1QPaMNGMCPF
NOZ/4e9MGTQVGG+FwGIG7TuDiQjGGruBkFBUAFO2+8uIe/9CibJK2+c3vfeL77fINXG9crIKBn7B
Ud3bEsLX4k1qXkfvkwbRR1WSt04O/fomTLOy2woxoZ3Vqrs6BavC4nR9Q+L9WSNyjIRWz7qItxJN
ZJxRHsDGJ4gXit8A7YdNjNiE6ZYjqW1Jy4ioyTAkXFNaJNYzeW0sE3tT4SBqraP66uuFgTW7uqgy
rmRwQrXPqNYLvo01gvs8rs8ISzWVLClmOd31PPP4VjKoaAQZN5oOIuP7BGxE2V0gm7QKuLpR+VHk
4RnnBxgSFz4enRPCbF5TCovxkoLF5iw1I2IYoH/JdQMn4VcJjvoRd7ZGlKETnx5nhxsKfGlv0g+2
VTXVynq3qIlQ01v51sCyse41H8Otu6/HY/RcxCpfiLKHsJlCuY72M0+D89VCm/oDNlUsyFBJRxuT
/3GMKB8WTLYbD9HwGQfeHUzVJzOiQ/cPTBkc2ebOlkB0UESjvMVXziRmfybA3jAmVtqGevpPpbxB
vrPCyPIUeZYsmUlxkk0Q/0RCrax90H5oICy7/b8FzR9rI/QkLi8W1ubsnVKULXuEXqDKMLZHjm+0
pTnhnDFfO4UURaD2z9cLo6He0dErrDn750XmbBDmhqP7c/9LoUo4VeZ4HIE94ebATt5RCFQIj2S3
tZBYXigGStpUoMT7nr1DSp9YW7EjKnJhvGKFPoRSIZLkZj/hfDMrlFB6gLgHZNrv+M2FyS7Gmn/H
IAlHNlwrMzYVxkIA5kEiad7Gekw24TEQS/QWFfR75bktXIHnlmGAB6N4sokwlMCLuFv+1iWOrOZo
UpBfxgkeSsfh8j8ezfWUUeQt3W/5UBARQobTiU314OJL9Id0X8Kv92aJvJcu1bKdkK4VCCZzj745
mPj2DGvlBT7kLIUSlfATD1px5wTfQ/n855As5xWNjaWIf6ivptZbeXg+8dc7Jo16NYmJH0IfZRud
XsAH41RWm5YtW7EXaTY0TR++/VgBkzX2e0mzXB5lvDLnMAFTlNOBKa7DCRKHWCu/H12Zwpfa8RZr
+mBCES2NeRR9ghG/wxmGAydjh8fW0niw2n1W28lMpaM63IQqRMby/k7oTckhbi3k1MJ6c4cxwFrO
PO8UnHxFKt0i4nqa3mDJo8cG1sqIZWyGnjCsycBw8MNwYJ/HRbdLToY/ZHyVSwykUS+sH2jpfL7P
J9Qs4MTnceakLFP0dOYzifGij9pp8TyBEnW5IjIxBeYJtAth0T/pHQU0/i3Quzfri+fcxWFXGJGT
YkE22Ne2432MC9R69cLmENp6bjYPbCVPqBJwOCPy49x69qvB0ERHMHQdbMJ7m5W4sqIHndeb/qzD
LeQGEND93WkH1ZYRlA9BXd17RywzmO/7JhybLxdPfbajj7xTojnZDChOszZDLQXdaPNwJGfy++xA
ofCtw+7pPW1tHBGYpQSIGEedjjmeI/JG5MAlYZs7WhRv5k4bYBYy01OppVVsel+/UGRhbjcF0ZAU
7ui6BXS7VYrvIZg05VIQYbiP2+K/XCTbTl807xwAGXISdZUXJCWxxSQMjn3+4aBUeYM3nGiK/vQS
t131eElr+MGghUfWQh/V30zJagIWf8eHnOB4nxzTieWg0Lq30otkHJ5AdaVaGOz0LjpuN4LnJjxH
thfpf2lAR/T3uvnESVEipTu2MHvTtuTLGnWIL1j2x9vuKQYbhkg7KHy6Vo5u2EaBEQpJFxIOoKnK
sfAEy0d5+9tFGgLWXtX9WNvCfFDx5Qzp2uxot3iOOX7+WEd0IETxpC4QI9rro2sadYJphbDuL8Ij
GwE22qNergbTyWAWkLoCcU0Aemt0XSZnACSIqbiWI0NzCyQrXHU+wEL9iAO7cEVYkZ+xoMqXmfzJ
O4umha3L0RoZeHS+GHJUkospgyuWIBdqXWU9x5u+Atl+ejZJ6DfDWQMU1m5HcBdKj65oYu6R0XYy
x8McaSCKgzeFikYlnzqU6jDd/PTSW+1spYjARnHDZpJdjb+vNJSFekvU7GM/gq72VbO6YYAbEPks
dHCEUIWb3+VTGMxe4mcEEYBgM4kEFYDYhTa6cp77kMsjmqyh9iRrseJNZo98pmpivRFb6q1tEWIj
i/fyUZtw4jp0LInXmN16DmnKWeznYgq0TKAuS1kM7IT4aDM9ru5+I42vVShDtnfUkiLitb80rW7L
obueidJpYy7QDjm3Xd2kGxpR7KK8WWJXHvJWqnesoeof+M803MeQI/KnUJRW3+bG4d7QlkMjvRcE
il80I4z8S2jCoizupUDmtWcHzPEcHNW/kOte6D0Rz7Gicjh1qN7LL5kbMLx4qUy2l1t0JEncbSl5
W3olmpZMP3CwLR8rfl1XlHqSyIBfCsV3z0kwxvzHsahRisJiki64E4cybd4Y/nkv6C2KcSESqpZc
Z+ApCvvxT8FCa559Y/WBTUQV67bPuLtFOEH+tMY5ck4y+j8L9ErkZkgXzQPUN3mSi4aIDwTXb4QJ
godvzAcBCkUubOicnGWgtj/OniyHLPoV14Hh1zRRXgsRG6Qp5D7vHwJDey4bE7+ZhTWg87eL4/e5
fOdDj34F2OVRlKA/K+AtuVLH0PK7p1ombXUavBJ5Ydz+9soJ+JBGLsbeudZdr4EKgNMDqBO9Ke1X
wQEQkR246wIYfeXecuh+rYxTGl/9VykHi6XOE719XuPaCTzjWD2kboJbU9mNhXnD1m0s5TwJaM9x
sShG1fFgeC+3iDQgmH7rLAFLZ8DUf1GUhningzZU5KYtZk92WbID32GtIeaQWtKgQ0Y5mU9r5ffc
jHoXXdHy+Ll7ubgLZmKRZcSJAfbq7sOOx6HoMO6FR2BvxCY8YQ6irV+1Vu47SbUaG0R+0CgHnqrB
sFTsnPzsd0YSmy3zB/PCUCNr1M1VEdlyVvvjxW2x0jRIHje0a6xcS/MgvPQCJMKsLkeZHRQY2wVi
dHVIeTy7NwSI7hG/+/zWnMOy828yf3VOFo4cuoms2r3g/sd0GjZLayIfRQPFq624E4V+T6aG6VoJ
Ev6TKcr+w31PW9uWRtL5bXeKhQPkgl9xyn0zO346wI7JKlYemavwXzt7TNpcjWha8rVzVkyITEEo
AblhSlH4qujpFxpn+7Yv+iHsRiyUFBqxEKX2YbLobLeUPt9QA59a5QFg5OwtDbUIDOIfgaOwLpHP
yXORO3K2VgvHeR5Xk/09NBytddAXylRM2sPcwoG0WDMy0lRZ1w0Xqfi6Oa5kfz5SYK95OzfSzB9s
IcWNsxoTzyR+1hrcfdunbVRfTmveB4a6SCBE1ei3Hh/boExqcZQDz+J9NW40ZDhb0KZio+EVoPkW
7kNYvrFUw/WVpNrN1P7f6qFwE6gtYt6rojttC2iPp3eZN/sR75p7dvT1sD/CSCjUZt8KXN/rmZiT
QL6fXIv4Z+an28PsjIRDMbwOHhHujefq2hNte82CLXh3A4DdHjtJNFH17xkWhIEB8MWKLDhh18T9
Q2cYkojmby7NLOwBfOeH3DmBDggvs3wBuRLKfvevKecqeFxY60m2BEN56zIPGqQNoBovadY8/4DV
hUjFC+SCuugPB8g/FTQXHytvXilfdriIBMSbQjuSDR5YlJV9SYQrL0dX3eDECj4alcL57zabMabo
GxybgbMPKqXgWZ6CKSSIBP6MJjTgojgfIQ0sJo1AOxBOb+djKObrNzrH/9zTUdRsts/n7aFKjbln
+mAIZW+VqqylKzsIrFQt4A0B+c/gbLYf8W9arxBDLUTFPw+1QszYmF3BJOXgUvh+pHU/0qirVVqT
dEvvoLJ6YJQ9q57vJEX26DeNL0T4hPIVE1hfdZ7HH5Mw7/Qc083j5Dxhgww1n9XxpkakrlD4hmCa
PjqTX3ID0Ol8CINRxe/oN/3PGyFi8aB7Nm46KAcoAgzk2ZYoGYilKQveADooGGXIHvhLn/IE26Nd
sSz1cwt0GVcUbyROCpBLEF1K9HAiD22mTonf8EWw16eAGAA7ugdeWR4ZXdfZABzOWYExwXO6gy2G
UpH/rGNWJs+p0e/lMiV83zcqFdeeesv4pqtGQT79wspC/SfHKyeT/Q9mAaBJ+q0rM66pnqlmHuZa
BINNW1LEpSpAM6uiACsmsqGpJ9EGQ8XG+2G7khcS7mbNXiNlL5a7IkZqY2ibjbsAuDna00eyMnp3
SVR/k7fGHRYp3lxNYEEuTrrrwhmUybhHLK2Up1SeE+Aphu3Y6b9hzoQekMxuHBq1vcLNPmiZ/yIl
354dtYM5OaDmmBXJV42KL5S1BWANxJ11AGmFd+dQJizeVkVT/jE4OfWbSSPQ4UVi42qDKsLAIKs+
dudTMr2EOBcBl2EVr96gNhT5yOscReM/VBg+XngwFhzHZHGtAgDR08l2KO/RuchCazYxKuwP6+PL
dfOt58NNMcclRBleoCn2wEAGgAw56SpAX+eOWrXp9oJPwUBNbf7cP3n54RiwaaZO3+NWvogSxASh
LNB3twzHDjmE8UtBqR0FjOCWqGNUK8WcTkLOHJY1SeR3jOCN9BKOJwQXRPf27ycZR8fBeDRaLZL5
TbOI/ovxvnQzXNG0r2q6U9iTHVd7Py/LeeoJImHg+SefhiELDfW7jTxm3+tEZoN409rE3iNUI7WG
x1UiO3V4Aq/0VZCQofmi7NQGZ62XTQRywxHUTIj+bdX3pSYSoqtuLnTuHP2tV7CueiZAQ3ju5JJw
fdOclVfPmJGxXus1Qr/sFiljC9pCTEj7LBblJQAiBM82tSxrpA4LnwLio76LwVEH66hrj8oADExB
pLOO1PnZJkTLxPUQCsTDHKtpJqI7npO+SrtqqV+5OCS3Ta845hOETOQF037ie3ZnmuGK7zURTJZp
N2XFA/jHETTzjYoV8euUTnboonP29bWpOzSA/fbjsZlWB/MUKSGNkA0p01fvoGeb3mTALcHp/0Gu
H+MQKjBIAE8QcO26kj1K8MCHfbXbmcH6FMt0NiTgVzmH14waG54asqr6nB9QkkXbK8yXlAxdF3ZB
6ZvkZY9gwihrMwTF4RuduVb+kJr14Kaq8CqmKWoj9l6VXTDmooyFU26bBmghzaRmM9zs1kDZ6Crf
DyKuCvWVELnVtBoINn4NtN/D9Dqw4+39szTVCuRnqmYbSpX4+Z93r0PSqJXzj1fBudB2R9NAqgro
mpFiQ9pI3ikkwmreh2pUrAII/QfK40s2TywZDy9DDKFVcvB98E47b5IGT9IFf4XWkBeeMzVWiVKi
NpEppGfIS2JxnLX1NofPga5U4BThLs2O6OWCFDnF8/MsWzyCTPrikHaUorCGgvMuJXk4kTKvtH1+
e/x9N5bN11gTpNvMPX+jg9MFkYdm/AfYTevsjR4ZAk2rpEuYAZXyOyU4eUXfzZpUwxtQYDodH2Sa
Xn/REgL7jqJuDpEIInRhoaztCSBVrRy3Gu1ov9lB80i5T8bMMkuqvNmeYbx5IbvZx0AP+ybJwksW
pgKBNyBoGgWrH8cO85bgBTatK4KNDaETQPS7wejSqcWhUuELw72/A97qO338ITkVlo5vwnS1Bqfd
tZT/1lsxF6qRgEbIFBGBgQ9sKsPilimoP83mZsQA45tNyjnXsxYpN24/FkPn8rFjC1LyBslFhgwp
VYf8ds3BH1OZOPnGWpP37wzlTAEQTKkslPgd+IeJauM8iaZ1ya18tadmFUbMwyddGyl0A3Ucd0rX
b2hO3BHrMbTiNBNk78xaCxiyDrbEHbmQm6ZGIsT9nO6Vjewf/DBnB5ms4Gvl9sm8u6XkW8c+JqPN
Hx4fND2V/0AcsYfn9Wqq5hGr5l4JM09Mjb7UmaXa9rJ5juWvFHXXeD2UTDVpSpyzL3tCWeSFgY6Q
HdszDDZ45rPS7WEB8l2CyYWgEFc69eVh5buI+1sXjKiqh+XxpMT4aQ2GVuW8vHQAoLbJ9Viyel09
nDDmojBQkgTHF1MtIAErdwks3yl9dAezzfbPFDJjGc7jRAdp3F3hRikuzi+LcQsULLY+EoX9jece
KxOrCysBrtGnoyo5NM3gxTQDhn+lw2yRp01k7+WKuX0y4G5Q/hOQd8g9D8uC+Ivi0b5o0ZWa5/rp
HZ3GP526uUP6YhojBv0BL92Qul6qa2ke66lSrxoLNID/J/8pDzHmDQc0OVCHFOasEtAFT0PRJifn
+VHNrWL2f46AQXsfnRpaJM5Y9rnaCzpCugv9KjiDFbNCT47EUwqslhRkD2K9Hcs1AW6R5jYqC6Xo
TAMITSdJ9Ucrh91dM/7u6KI5bcc7kJfuMvdix+Efp79UUJrf43UtPMcpxe+GnOyRMdwNFBzZMPsn
smXFTSVPfEhEFKn6t8AqCdeBeykTqxmzg9ImMpaieY72yoOwVQymv5G1N52LPp1GK4FLLFLkKYH4
fQqlFKYvwmFTGQNgaVgC/LjDtsY39o1vaasaLg6aB/95PvlKooaXmn6fK80jh7RkcG4///8M3zma
tZQYkjuORku2NBsapOFl90ruP2W01VqfOfMwgZBPcOgjeFUZ4G6nKNSXll8xVd69qr/J5CNq2PBE
fSuWfvboAyPFA4Q1fNjIYCIbtJiMTf/Q0hgmYDA4qxReoI954ZlBQcWOwqwRR1oXEU0ydDGLEOo6
Y2AMydbShxa6DS5+DblXY8dPech156pkfHUAY5lhH/Goc3Q2V2cOrDWeJ3XYgNKqm4nYzr37mjVP
XFjtcfUiNatoP3Q/xU0H7+pwUIacWG42ZH3+dqqcqhqQyTGjxMMZF+P7rWFMJtBg4Tcf6rpuOczH
1FEab8g2dh4wWanJ4xsHUM87VvvFVphBZs+GrHVJFLrmdFV7BfXOv/T+G58RJEbWP/dlF03C5hQ9
551GIUZeUS7NbFOrUhYZ3j1Vat6BK5BUNgkfkW6KxM5xoXFDEcdX+OBZNf9k9nDCZUE7TjWGpLhR
DiVGZx3NzjOz4s+MVx6PB3ePFz3QVS495+pIJ+1dfsV/iOWOoen/QyMV84lbvNXpvfMgsn3Z3dQD
dX3tmnYsPweBsWqpZwvCY2V+I6chUVU8XuAH6avL+Ne7Ybh9kcohZzKhP/uitLz97RkLs4iD4zcW
jB4CRW/gzClkzAA2d1YfGDT3nc3F+tH6GeJPFvcFSEaFY8RVNRaE0mmybhO9IfxqJeH1N8y6Kes6
vU46YhTEqc3OBrCKmAw68xvkMtH1jLuNVbhp71hL1Su98eQXS3TPmxL2LmfhFDio8L4pJc0yvgeN
G7Xcjf95L/H17gDYQfWgr5SBgzkPtq1+4tN8+zcg0a9xfqTn5c6OAwl788zwgq2a3YdGU1+UqlbH
0pAf/aLkMzrSjt/6zTPnUZvFSCSafhx7TNj7auXhHz45DkkMhWXdwlvyAzUlvUInWhAECLJHUXhw
TWmJlMSJxPdkX9UujaT3i1+Z3Esdflu/pHrlM9VyNnMP1feevXVSagrl+w11nxiSi8K8ay21Hilj
EJiG/JrBImZfQeElUZwjjmIFyfUrNz3UE2bsKcW09MQI8ZdzPCJD0g/oyIiLliDvfmtboFamglHe
sXUsBf+NelDVznjiYgCVffVg2+IcTYqwmzjUnWOTFBtMkxkagk+FA4Ovn0nFiUL8pKY6phPghMxE
pPshochAbPScc67mu0acbs1PyZzFO7sWV46MrEhKGDlw+69mK9BbzODhTmcySwwzcfegTsAZ5PC9
nJM0wDoVF0K6jiVJ7u3E+qP6adPcM0fk8ZsG8XIFtjGWn/8UQ8GJsY4QxXo+oPcCktAVYowgzRtT
sewsjJmGoWuFLhgjfp64uVwlGqj6t/t+3e89BxMdnsZNlqIKvY86w4DpiwICQEDHmiybsMj/Kw5u
vmlHNvun7tPQCjvTz9MIwF6a3V/2pH/1Ll/TuTtRzhiAvCyk03/1apSE6S6sfEsGWzoiE4IAhSKK
rgOsQcMVHM56vxlPHL+ZqbRGfoUenl9oXtllgmmH2rluFnwLBZeqZ4WcNMhU2XN848BQBb3+qko6
QEH8wFLxNL71/qRJ4cV+QJYfoeDPaQCH3DrKlum3eVH8Q+r6MS6Gy5iKe3tAkCDsHASyIJ96E9X1
K0scXhWZLXhAlyCo47mKPuwsTLXsq51ryHTG3i67+YZZbbRD7ZLMJ5crK8wAyCsZEQ6nA5YFG//2
rnQoEzs9eQIPBDpZh2GTztNU7pcp2uRoMTZEhXw2uC6V0lWWENwPeXOyAW0DsH6KdXDDzCY0ko9C
TVUw8MSw8jg7hhL2g/sdXUfB1ELsnTGpAyw4QRKjuC4okbwtm6vfdZ5B1OlM7H/7QKXz5wQJ9V/g
I0LtRoBzdXGiMmVr0g44a6mcIYP4+U/EpTOi0qZWshn2boF/g6y5XoaU+MvCmAlCaIn7Ej/NeIGL
RTS7d73dbNsMemqgaCKVUkxr1cKoqZu6VT2F+Mdn0KKBrz5ckt5L5GIg+G6YW1MfxwHdmjM6L/37
j7Z1ktvVc+dKDKDxRx1Et8UM9wMWVHGHv3jJ3cbGuQ6T4FEffJD/VnZhm2opQp7FOMESpJfHYy0B
xF8IhHyxPvZHNEVLJHfKh7er90IdtMf/D6qlml/GE0qsl5uEWF/Zi1v4tSm2/ibCeGzD+YO4VGlQ
QSHJAHqnxr5+/xW/FmJqO4gf1gjjbxHoE8GD+nb5eKgxWZehQuPN1aYaqr+BiXqBbcjqvgWxFzfi
TW+KMAr0PH0xmx6Z+hAiClb27BwVvImXYQ1FdhfHAE9S3irI4Ee/KlY0nwHWtNbkN6qAOawPJk5r
Z361YP5g4kH/xLjpT06MTnvNq8jtjSG+fZ44jV/On8/WNNooFaAQKr481Ye5wlgLa0lpYj0hWvr5
t1ipHoWZj/21zDyJ6urGdeYZZCALDzMqRAkL9Fa/wAj1r8+ImUzRg/QLtle3Vlpr8kV750BtfOP8
2Af8hky+i8I4A6CDPmaW/BaqgBwjsWXyBdC3rmNItP1jxowSsoifAyv1fL1LonmCnq3SA1U/JlZv
kA4JJOcHna1ABDy50WHmuiMbxE8Gjsqp3/8puGdyBUnNvk9sua0/EUXAunggxzr9Nhcl4wtzs9D8
p5kkxdNW1wxKWJjEl2hWBsIfrcAcg5Zwp78Iyr+Plp5e52SCSpKPih2zfPstf+VYjS+jk+ZMBWUC
z0GZZct1DQBVvLx8YjPjWTjoH5/6eWMohu62cBUoQzOWeQHosetAvEreqIAeEfSa7wLV2lg8koSV
xK67HizT9SzOlZMZePC3Wlg4cSAGh4lE7iPKI1x9gQpMirbIB0HANazGED9ROynYlD7yekwgintA
uZ5JyONvPmysXzybj/xIyj2PJofj/ALTQTqMqvfpc+lLqkY/eM+3BlqKsGn78Mn8lNY8bC0cER8x
JsVQv3c4IMVa4e2/Yqu5KjCvVxt2e7Oimch8fzJ5JaKN3o/qolnK9EIbu3/K/g8l4R1QHtGmBoHS
oXTqM7a6Ma+qHl9j+BhNwX/0NKhJsWA/GC/9alsFZZFx123wSX6TjkuWbwtL3dd6UfVqeRW7ZQTj
zIcVfuN81gvlRT7LV8eKzpDN4OO3jx5TLAvMhQOC4MqJnMR8geMMana62T93SzpOfuQ0i42Besey
0lvzxqjlKbN0CwpFa9LKlmZywlG/+O7QbzGLdd8uesTNhtbxgL0vPx84PtVqtIHSkS7gfUuaD1yG
tjyPu2j+HYJgTjASw4F7qyNEhh1SGUlyxO3OR1mSeDcM39duzsEumzzQE9bXWafMzkaYQHQLiibu
lEJjWmOl4LLdsPO1s/AI4eo3LPcpCb1wIcHR7Ydv23RVrPTU/0Zl+ALcqjnvfTM1DkEFx3mRkcz4
QVDUAERCxKqYhYP4VpuvoL4Cdbdcr7D8xPkNHl8fH5HNF5vFe6Y5dtVSiRnMQalSQhoGLSZVXlF4
WTstVETk2PhUbthfnO70vzNSS/o/Jpo6EqtKxTne3/KLCgnZF8w9qfl9cLRX0jeoE4s2+1noIGYA
tEEV0DYpbBxrA8rJXFucalG83H111gbO9tBdAoMixX+kaCWZhncLZNxFuVoqNRuPzzSJRMCjnqAA
2TT/sJFmtgLltnfJ/PJeddEGreexDW4muV9LB57CVggv7m5U9dW9WANn/4unyWEo1pVC114NMPjc
z3t9+AXE+D4rK4OAvvFd28eHe8p4tYZq0t5UwegeCzvVqmy2++34U7eQ2m4Ma3+B7CZhdJfTfTq6
iBHgnNEFEKP8HqOVYfQG5t58EIJFNdEmcqYqzl6Jl/9qcXVr55/tmbS6mrnmusDcYXkJmg5hFMJd
bLPFdrjJhCRKFb4PhNipFCMXqSMmllccLQ1lyQbpI0IVwr1Tg7yjTYDbnNoWaWqAQD0pgqDmGQ9A
+oTzRKz5CgAgBwoj+88+/RChFdNiUfUMqTsw9Q16VDViyWaAUB9Wz5AUF0Eq2ZjZee9Hh3Bar6dc
6VQZWbTS1jDzV5x64tI6PJvcEdSdJAaGSSYyYCDDMyLlmtmsYmu1ix/RL7Gu0CG3JBX3BRqzu/pi
b52NG4OfFA8AsNiQwaYd5BNgFaorRIoMXIBbpo0Rz4IvR++L8oYNLkmpGMgqUN1v55WhCpOsLqHQ
v/TME4x76ml4HCdoHu+iMg0rr3tjCHB7Q6dDZNtIEgAoCXI6vULDDTxdYLOJZ9D7XomVx7BpNR3F
fdEuYTUa6K9Ju+aGihLBTZtiY4gvZRIeXgT0bQySYOxDvYAo9lS9vBSe6OU6US8LET0CvaxbWGQJ
3mW4Yhbg2+wbhbsm30SNu8WYS2uUZJV9utREIqWRRQPiLnujhzH3EGI6I0PMLL0vYmdKc4DlnfeN
0b1/H+u29ACXZvUhucDZpxSsd6iJTFsfDGVGIOZUjwmW6XAuWGpWQtTu7zVJpz0SjRIU62RyUOkn
DPzjCDRqkDI3ATatEF1ezgZfGCk8U0397HlslDClnztEYXHAWxC2Y389ryqkli7fRXL8MrL04R+7
25oR2rQUOmT28u6TfYDWYmlZFKhsR2+DUTwG0dnCH/4KN0fdtA89dTLOkdohZrhXjxK17EZSZ8ID
TyMvH2gGgfUIYtBIi2mRU2ciyzNAn0PaKCI5sbPiArK/fPDlN9vD7rQNCRpbecvwHWECH5O9bVi8
UaMWKCwodYXv4cyIeecHDyFBQyEgapEfuG4vLc1ZE1Ef/rI1f5+my+wX/sjSlSpQ9w6LzrR7uAzU
rXuzyTE74Z12kpHUePj7oK5TkiIHHdFuO/ADI7uv3mqCMmmmTocvFb1iqUUJbIB4Ba0tj7KFqELs
2zhVMPx846PT2wY4OempqghcauCOFuW1uuUge/US0nJ4Za83qfdDRmRdt6wH6ZFCgL4fJQgrBSt8
6opIqgZPP/J/Glu/CgYov1GHsmTtScteNRiIH5cVYtlOUara1oiGaL4as9lYRVYn9rT/o0soQcMc
ej6jLE0ZdbsCbBYgtZBJwvHk3lZeUtv5UjW7tNpuDtjos+DNYGHunOYuB6OIYTcnwZUtXpaodgg8
msQGIOp9AqNy8U7H9QjRMEfm5iYDYlm2wnOxFTIUe140j6XblpR+Kqo8k+r7CxUeKPYib30wpQzn
S9+Uu8WY1eXprdEC2O1HtG6UUoHPAoQdTx7Tu8UEV1nhNQNgql9JTtBkPWkU5dbxhgTpl2atQZQp
A+yjksDH0+DtQ0V/aYlLNbqtOM4HHfYYJb5AgCUbjr6Qkg/plPq+Z/hUOibWvG8Sn/vKzhPTnxY3
0fEfQTbcrfGaRN5PuPqPhz6pTymzxz4yZ8807jhJqJqjRm/wTfjwxNhc5xZgQcrqSH3gPKexS3WZ
CHQ2ieIDqiqK+di27f/aDnAkQrSbWP3xdz/ilqeq1sT2qgexG5rlEWZ6LPlhDLdXX1KVETem+k8l
lP7ofvdYrnfVjqYtRM4IrUVrKuGzVSdbb8fYMEJpFuguBjRYRwhGQn0Nw/bQb6HgH5HB+I9wjf+5
BIKDP5Xi9btnlo2J0gOsfl/eum/PTtNCggws0ugErA4vY78ISwaz+wP+9xiniFMLufOXMqx+DPK+
miw2yT+bmDwppPu0nNiwEv/XOBggkQvUWX5u/Q75Cgk12DV2mShGiG+5IqxfH/X3xhKU15Am59ot
sU4GmPArLlNaT3On7isTJOEvJ0o++90Cud0eXQWZGpBxLbEAfQJDz7JmI4tsI4uogVd63k3vTpbK
5Jz8Al72TOraG4pe8PAz1es51cFmu/ZldGkRiP7Gu9OThpz0ZbC+68lYiQ1/YqbrAyC/b+C9XnMN
22TsG6IWenO3s5hA7hXorbpJYirYcnybcjmpp5fAgN1hghOSx6oPYFsW027SlXnYyEuGw6iMLVXM
BdE21s5iCus8hI6trx034zfyyHLlmyeBzdka1SBMDZ4eThJWLOGFlQPbvugpHb8gieqTQIBo0B4z
hKUwDphZiiQ+YD3FN0+S8nNLA23o8F97zPFT2JtZeKeCigM08Vcn+kuL0Xio/1mECVPs8KdyBQzS
VGl3zV40pw/yxszicpwNLkwHqhmQowD7vAzjZwfaK4CTpzBi+x4oyDBYvejV1Q744nZCOtcOvl1O
CHVd/HPePtofbtwBfl4TLsm2TbgL9d90zFqZ4D1v/p+jMnQfwEGoRjedMkrZLL0XsD0CvZA7ocMO
iWT3PAtbzlbeT7CIHrqniGq8O9UWnUB/KmpJ1YLriEehIbO4+pUj4hwW5CgdPmACBy2HQJraeMWS
4OfWRhg23Jn2FnF/2GxZkOjgqbJLbGeqsai5TY48iS1M0qxeGnYc6+sSPM8sCXxL+BTxP0hEFlk/
0htERCB06Ls4SSa6J38gwU8uff4hIMcaOA2gQdVEAtk2vqZziSW85YlClBNpjY8ztY5TGFESCABy
u1PPDpoJZWQC4UMOsUV3nS2sdDmI7PQOqLnQbGKZYHG631wBQRYv/z8tvMuXpl9cqRqvd7d9eQDC
T9hv2FjaSXN3ezsXf+c7SXRnSf1Sga6hDKqeHu05YH7WS6T8xcPG91XWjqd7+uBxGmTFMdVE0Iwt
KTQvhNdZpu1jlihFSC0KlZRfwXnVXqL2y6QQnP+iJ/tCjUOj9bpCIukKMhmZA7l3LB9ZzfMrorVb
8bq/mm6BX+NfZ6OCw84DZMh/s3n5UUPeF+Df83wrH+ZM/QFKbq23NuL9gmgyz41qyN4e6JcG5C1V
PC8NHwiHKxlYqTzUy/eZUULZvRHd7isnUPF0bDGjh0DJwMbeF+5W+rnb7t0HtYfXVeWPDtOtxgzL
x4HI1uqNt0wABR02gArHNTo/jvHCIMhXVhmP7Rqf/uhXTMPV/Pc86TwI/9K8R/m6zo7R44GCvd61
TdMi5hrFmbOhwrU1SFXPS20GzsUOnvVHGBQ7UCuB2e2XFM3+QmiHrhvyfSRLBkcNEqiaX95cfjbx
yoPTeoAy+qxwi2goqqZmR0HTUKBUY2bU06jfxbKOjxqe0YN+8PzRevLiO/eOfFzUT+RJb54FOYXI
dNk7Ok7XTDy7Dl8Up7q0KCfgnF0MzEheWsso9jztBrADSGLQ0lYTyOczM1vFqGA9X2gFdBce5BP4
vpBHvZKSpiHOvQ7vIPGydnzgO9Tuerbi++IoVdHmCDtSSD+hBvMzGiw3vzmpArQfSLaJF07AaQN1
b9o/u7T8tt801eYwDTUV5ETC2w5N0LiZKYYeegt2dfQWj5MKnWdVb/KKwkdBBE66+Ga3ha6EMsqq
eM3btvEBfDtg9jaDO5COShy6kCz2cXQh5LcFL3HspNgmRo1aUn6CIrkknqXuSjY8b0SLKJfbkNYT
7AMz3ilawbWGZSXQlAP+8Zy9hum1HQH12O9BuTZt75c57li3JfEXPlUgZWHtHt1x7Cfk1GAXAQbb
WNJigr4J1/Yjm2rGdeagaFNXbAgZIh+H0LX+wtVJ4BgdzS+Rce82TiWHpKTEY/jakNNi0cmc5aBG
quISNfR3q1hpTdVYQ86WVgsnnA1UYGaI+zk7Qz81CewNrO0w4/MSutpjIzJzCBLqvB6TvfcG1j42
o8Aew8iI/4YXElZxO1Is/BhhvZT8z0/G7jDh3atsSTn9amFZCKMSRqjjZfdxhJcVwOwVVjapkHB4
pnCOQjXhs4ME4h16S3OhxjP6c8kimGY5zBgp2N+HnyB1XfnaxTo/PU8cs0SOR8U4W5K8J/j4F1s5
cjiMfUyGG/+XgOFtW5Yz/MJTt306cbAREXQvKOKDlrAejslF5h8YXZfb0MtnRma9OA43uCR4D7T1
0VQUKQBEP+IARI2mqdPHsim2EaCKhSDXFdGUVcKfN0i03e1oMJ7VJsBbApHiaMwrt9yj0xOY3CnV
ds90oRs/lpnVyYhvh3FGlY3UbkPCBgEj6c+T6LbUfJZZAGkRMmLcGuhPrxsyuA7RDaaV97IQ8SWf
gOC+jw8oa97ipP+Pu9VQGZHFeEkSDUpzuOwrsDJN6adYq0aaI0I6jgZ0EftK4o8spQELGoWG4Cag
8u6b4vL4tSEC4xGoeCVlrhxgWqThRoa+aW7V55aZInz2dVgRUxlQimiPtd5uHOHLvIUf+FK6C8Kf
DvjBgdzvkspaYAvh007Ll5G95Fc8kJ9qOXMd5wCRIn4LMgww/h8eNDRayKUtoDhj1qtgUkM7NJNa
oKxQUbR+AEZhdvO6wUeDgh9j1h0c0vLZa4yWLOJtLA5+zvLFFv4H9cw7EtUasHNlX/2/2d+IkXYA
SakicHUlknppkDBYfRGYBot/U1A7ITi2qa34ATtAoxjI0ssHN5Zb3HxxzbY/fkB1bcdDoOjI1N7c
bv57zQg5hDMAjUBZcxR7FRkYWYJnCOBOk4ibcTeBNNr3CXF+ikNSYF5aZwzsEaDll+hgADO2f1o5
BJESO0F/+smkgaZglPuuuQJLpA+djwB2zDOgHz2X78kOUiaU2+ZuTodlAV77J4n2iWH6WSUlRC7B
hNyv+rlF2xHcYuqV7cMFh36vfmKMmJPXCPOMA27ipyWfLNLMz2R6MuXdjiO1KwxF0gxLas3Od+Co
I6jMSL8BaJDQgwp5CZdXsb2XfSWX7WumNm0a+FFMErH6TKgsm+VzTQLhQYcNPZ9ErhHAx17gUrYc
LKXghOuCsywjxr8ffTcVGIRcTtHRtUMcIUoyAxIWYDjeHQNFAh7oRcEAz7DYoV8lr3QSTzkbIyw6
iqyMoBk4SfzZr90st33XmLF4eXYeBIypSZlUrPX8/DH9T3D4T1M+gsB/M1SxkEAAmkmE/S92Nod6
EcCM6qoMBuFGHfOvkJv5Xl2JfiRgXskrPQgszHJVPvtK8Fj9LPyF27XuZeklI/wXlnGbjnFU6B0H
YnpYfh6+4Du2MLqbaw1QbeVLu8PWiTZSgeRp2NDwcedwJFZouG2QC2a3iKJZTpuemEzv5TWL7rQv
qyZREXe8Q5HXpa+UT4sw4d4yyqkDwYtQml/CpqV9pVrv9OZj5KnUq2j8zZumtt6IEwaEq0jYZA1a
xKQ07vzWWH46DSdR6vJd9JQSGAWaqyYB+rvj5RyOCOCzbyOEZNnYwmUxiKJyTXPOAWUAgeGu0vCs
eFsy3CiCNjeh90x0kBGHcaGjx8OVys+y9VLijvH1d749KpBXQJz3UuwDIGRiIVNR9NBZ/Av3MX6k
ScTNn4J0TMfZ+8ROJ21GyBNx7P+lpaXnqg3HIYMSIJ07qVqpfSld3R5Xifuv0ojTgL4P6EGUTNTq
6Lq3pLdtzn8xZGf7RL6Lk52st2KzgBBtr8GMeVwXju+ZxUIC/NnMltSRQOTJaudFdTGvAIwK9uzl
PGfxJSS5tzL6+1q2vWyVHqglgq4ExVhR5LmxDoGmcN4V9hnRkot/4pWl9an7USu/P9xzojPywD4z
lhIp/ck8RsVCr5hjz4cdUOHyGf72n+gUavWpIjkdvAT7Mib9AvXoi/oAS4VqzKHJjl0Y6iwiyFDM
+L79HlMpslsrSBPFtRN3diiYZkeN1UDwxWMpJ8cHo5C8YEnzbKwEVaLTqHr6g4t07VOalQDDJSe/
9ucfm+rOEia+8BrVpHhJXdPVUllXvdakGtcz+VmKWx1dIN2Qwsw8hOwp3ejLRgel9pB26khdEbKH
TxODqG/Ho8dYtRwezeMNrK2IBPgFHcNMS4DuhdjMv1funqodDOrJhcBwrHtLywPb7/pLAO1fPGYU
J/0m6YXG6czlSeIfl+s7sZVGoiDgq8DKPRCAMAnqlDtRgGs6PSeumkwiIFnKlEB+eiHTheIESHKv
4sk8LEneyM20VtJsHZvkOjJ/3SGPSBn30uXh7ZuG9aJI7il6o4mJ1alprWnIIOosvf/4SDc4JrFW
Hn3QW/MsF4CQNWI0BQbfDclfEMT5oGmGm7OaEXwvK0MssheYB3wdJOWkhui79LgUIdWvpOT3tH+e
/0D9/OszJrnzgSdcC2hGv7afZBjPe8K3wXTcKb2A9XV3qGgpFkuFwC4DsYgNV6fhEdheFqhui3Ak
jazUSnk4azD1OGEwtLdzSUy5BeEmmIq7ha4UXN67xS+QyO0iqZhAEluvp0OAxnuF2djVCkqD/uok
Pl+/Pl7ytNOt4z0BWVONLMMZli6O3wtzKQ8/IcQUydm8WHv8Y2BMYuyTOS9ByHRN4PtJPS0q88/7
qtx4hNTx3lGkS5aArZlbto3FETYj7hiDfgtO3zwkqqwV6OCikwLwwFDTcxVdpJWJRqRv1hWk+EJU
EGk0ri6tl/MUdxNfMfFGZGiPe/RhpCK+xtg7vK6mLm61EWmZOdqT9DA/vZAFirvRlwuVvXPCwiig
TUXWzgEQgLt5RaJgL5hveTv3XxIz29aPlYRolsuYUecvxNgYsHA61NkSqPRyUi2yJ8xx1JoodPrc
y/+7LNmFq3lZULPDY2M7ZgRTHqEF4wCxSX/ypKvfK2BJaTrYZA5SUTsTZax/sY58Kg5isj9NNrhU
QBB0mjAlG0PnOhKseJ9VaPViwloU1AZ/rYT5QPB9/T3oOZniQRlr/LVmFeRlB2MUPfEbklZoRdNG
lIraXa1h+UjyDUrQQC241Lpy9CfTHcfk6xapqv7lVojopGmUtQmUtmCLbPrPIl/675iA2xuy7SM8
1iEtumYHWiC6SLAtPXJFmOsg5FfpHuPtNlM0lBZllnrwPDeibg6jsV7M71Fy2z68vSVsTwIzN6wi
r/+TPe2d2lrno3oVS4zg4hiNxfR9INknQzf/7O1VCXCKGDJyRJXRnvazvwiC79IfgiUKnpdbllnf
N/i8S5abSsekCuitH1MouG+7K9SxglrTPcpJzP+bHweKYiszco5BjioTlTDjfcNDnF7+z5iHByPL
sn/o6xk4mL9EgmA2pphPTAW0J65P3eZ+kC+v2ZZwxikQhc7XTc8UUR2s0SMHYB2xj59/QgatQ8VG
//z9ED6kKtyaq/DTxFrHhbLbbAQkCOGNCuyPOVqsw/ObR5sfh4R3vbdDv7tCjMMxWTNcn0FgclaP
jEGn/4pN8ZYi5cW/INUgtvRnWTQRZmviLsicswQ2ow8AKRZJvpMZhkCoN+mt+6L9bZRCQWN6TEyp
XOBYse8rRXZybDlW/iWj0X3aL1wqiEz+wUlMh9bqD99dQTOKfADSMBgaJnNAxmsUz+YEN1KXRNVE
R3gGv+1zP/k2NJosDZinHWpHUBoqm9Uk3My2CnUMdvF3LGfyg7CVqC498jOVB92mLSw7AxyXGgPi
9WwrLf8DHX7czb3kkF+epOU0q+7j5qCWRjko7CouqCRrgZ8hs9Kd07RzPkiIi9ggQi1d9eWgbW/e
6e9Y4JRF6NXSkDUjfS8Anls7Sz6qhR7/DdaC4NvCt7g3C8F239CSrcsJvgIaWlEBYSLQpaENvTSQ
pH3atxc4eR19Y47OZ3jwO4RiMY0l9z8SId8zNUv+VngkaLiUICoUTdd6F61DrCb7T6u1mgoJuDSI
J8j15/hKAO6/O9UIRMLcJMrI6/p0LkloA33F9jSBVv/BXfnn9E+rjNRJMYqFZ0QIoqPDYKSil4E0
t0an2m/gZ7bzQL47x9EHA4JgHpdd98pUdfFaAsz9ekPdL1JCwa9T2oCSLta4zKb60MLim4xLPBJe
F1peCe385z3zHMpafuKdIZepChKB43R6Btr2LeBf+StLyyL8yHj8lJA7l8pxkeJwtqMO43d8q8mY
QQJUfRtAB9GlS6Byfi8HXbnbrbkqEpQSZ0idZZTJhDCOkKn07hnp4B8JhWblA7HY/5YbO1DJmiXF
Ro3xt4MzJ9Q60cDo7QACKojiZiCXnzTO/iPD6UffetZ9+Vqq9i1tJoZX8JYAheUse2KL+iQ0hOkj
SSbbQkcS5FLrthI5QoxlTFy5LYG5627B8VsF94O/3STU/Ztx6n7jfLOS2eXBw7MJiEcSsTqWDXj5
9YUTxh4LRpcP5LuatapVF4Os4cX449WA4KCRS0YZx7fCyLw56uTafBiGIq+axUHITlSZ8i3HTZv/
fLKSNAESVpG7FMBD0JQqAn4mWtK8aqP/FiXpxHGjwrPE8lgkduUe1RB7Ev5B4eY862jw5IsxdlJd
zElFvfuKRk/FNWF30VxJbgLWCyg+XGET/ihkTl9VKuA+D3BpH7t551r32Ykw2RpN6ym9gagI0voC
MbU5Yw0Avo2+WC0koLYjrJvc+TSMU0b9q1FhusR466dUNJrvJ/qZ6MpNNM5iINcIRq4zNvSBZ8kt
/LoleeC5CMwo8tYUleAihiQUd8VoSsJNEABPsoBh9ZfKyi7iJXxdG8AXJk3WC8S+LKes5jWFBSsa
8ZWcHRg09kimgOsIn+gL8ftrfL39Dt/slNDL8RvtCgGk8jMZ8O3Ve0CJ73vEzDTvBqyhsQ2VwB8O
wnbCKbBLZjR1sUAOUm8ByDzAg3fX91mBkJAaFlcb6g04oD4DroP2xQjtCiTlM/TG3vI9nUndPRZC
sBNgAP2iRhgiyGo1HUdMr93gHxjNDbx3QVG+QQPtZYpyQC0ePj/IbVKODZbfHY0806UeGXB+S5ke
ZBi1M/r5ndLq0S5HXCMV0N16jwm8VR25hmHz1ou+d0TkaB4RIkSNnZ/jdycy/BQxfMGEiZdC+wvN
kp/1N2fCYe+hyVBf8jWRanWEN28oQpLcckiUnnEjcOhPsLgEUj2ScTFSqj/Kp5jMlFxXONpqf7VG
4mbCgkiYDciQCEzMNyXwQ/yYAWKytNp8r0cpNftHNbRclvCALiz5NZJEVJmEwheXvmuFTdVXXtCZ
+nSKVgrYJGPoA7Fd0uzlG7nYIqwr7KT8Z34UJk/Qvd1cqyc317sJLGCKTwh3WS2d8NeHxTm6RaTn
amDtZVO8NVRBtY3HPTEoMXYNxp26pL2n8vxsDSiiBEKBJidAqz/ub4lZpEIcjXOtCNKVPpC21YPZ
ayZxIsnbVX4txC0CIvk0QQqFirxiXQ60L93kTnCfuVjExtMCFihqlgh5mxZZwQaem0VVhF84Vl7e
cK7xYzPix7PkjskwqSa9JIl4CLboDEIwN3/uB79Zdf2QgF/VOYqEh/TSclDJqOvg6MYICyZ8GBx7
bxCt8KD+TZ4KVY962jvK6Xi3uFOZf2gGqMQUNYp76dsHx9wypzvx+N1YkdOn7sHw/CBI536Confj
RPbB+JnJ6LwyNTfVU45DexhidcBfyleLx1X+igQXDYi407U6wCK9YDl9ImbbI3Iag2fbWJtf7sJ1
wbJD/QdmA27n2viWXadq9o86C2146w4EUQk+CYRVFPUzpN/nUCd5+++yxLl/cPiOnK27CR5gElXx
sl4QdgXLG5HFxU+j5YzdV20cc0ErTamRzRRA4LWbCogIazi9ebx4UKbKm2SEjMNXWc4LWXuH+wMv
oAaSwkfrPF726RelppaHbY6BmmpfgFimB7CfBPShrgbltqmL0phaNNAjAn/soM+OBQrYctOGB/n0
OwMKcUUwZthV5ioWO3HlOIEMi0iYfl+lkfizwmCACPUAy1+wJeB6cRR6UtSEcUU9TqIHk+hVChQY
gfpf45s+qlTucARU2FLjLUYZuG0M7ArDFRZ02g15fQIku8HeNGO8v7eu+xm/sg3uqJ2KvRHPPHRg
qHgfYvXYaSYwE8id4CQ09KhgTZqRkAhq8fRN3YWjayKsNKCIKzc8B1NveSQ1hyEOBZ81xQkp+xqM
UxUi/+cWcf3igc4Y2Yh+QWV1gITLjf/lAurJxq46BvRzg4GrdVbl91ISOkdz3vx2UFb06/0qC3HU
NlVpKNWObXvg1fo0eEshFIlqkeBlSmJi+WI4xYOjmFn3WuYkaMGRszrd54aor/fh/0g50WWtCmAV
Z+cNze57xiOTkfk3Gj67TRh1NJF5oZVNqJObO3FAG2ZSpmgeObwg/NtQLqI/lnA4TL5Kg+thFKPt
xQ2yRTAjcauXOdtEATzOeXs1hiRuzma8EcFWK6Of+UK1p64nrLKSeeOB+aNX/Ijvfzqk602XcA63
p+8nkbb3E6GVUOdsVYR0eatQ2m/YUjK1ru0YZCUCquUjy1FMOdH4jY9Fvf2mnxhBl3S5LM+Brtlh
nI97YTYquHgWFZbznQCQUIOjOr0NBjuWVzPwNh+x++wCaPpI7oDImusDPikimW9Bnc5myUDOTE1Y
DwywwqQvYKkQRbvMx/DSBeP/aEqm5IYlGJaqXFJcnJWyWIwoLjDpFaWgZlqFqTh2xqSn04ZtwNJZ
745ImsD2lZc5KEQL30DD/PNELfvK/hfhvy+lt5vA6azwfUDs6bMJmzM8egqETeYuKBkryFab12iM
ESka1AZPVlkpIc8Q/hxjVOrs7/5tLCu01Pegq6HMM2IQcTMIamKbqenhpTBDM3qoZ5k1TeTiP3nJ
295in0ke9LqSJ1Gy/Lf48I4E8tHP5uw7bkhHn8ZRfZdH9i/rf3L1GHk4euQzJK0k8J6n1h1/kfS9
moEl0rGZx0cPBQnA2bKCaxjK/7aQqHuGLIQJjkQbPeNiZNZFbGmEJCaJnCHYD2uRTYfzUyUJXyKo
aCsiC21aDoajaS6JPM50Z5zfEd4Ut/jHMOFwm+wES8reUv/jsltGvkbwtqakjrtfR8WzOssbfz8x
v1FheWqweMAZoLdzVQJQgmPnAqsH9Os3Qk+8kBJuwD9fyCfx80F5Poufv6Hh/LzIcnZ0GFHV/7ny
6fCaAE+pLX/ASD41NzmEKPCaumzkIUzFumEDrnSvIsVlVtrO6NRn4JzuOlQIRAvRp21JQznPTw3A
+Hb88YXO26r0Hye0kpFsxx0HuG6hVE07TlPhoXuyH0EG3q0Or83Z7yenod0AUhYihqm/1+OZI2kJ
p6n0n24nTXCOAUXTEs/v9qZOIOROlP4TwHkDUKL28ZRma+ROyUE+s1n57u2WZR3vMwzqjgh0otLZ
3hQk6B4/xqna/ycn1LuKmGcnFXto8iHT+sClI0jTjdeXU8EHAlbjRi/k23PvVXKVsq7G+lYOI7uc
leqLOYqTajTDARhaoDL4I0ZS1Y1NrU0JgPUZbH/BgXLrsQ7PDrV06bs6JA5VDfCboV/HANUCq8c8
fBaejrpomDqA24RDdGm4pMnHXaMSppRnKuC1yh+E6yRcm3NM5vQ9z80xU2F3NpN7RazdJjg+nPX5
u/7jb+C6Cbstsf1EP9LrZjzgiC7gcz3fdrNnhlMz+oDW0BYy3gYbCD6WuiKI58hKDcKpP4nJTXDV
PD8rndgNkdbVo/7MYaiqRDYvKx3F0iioo9cwmR4cgMWWMXwo3ydIY+ANM1+HasQ+2RCs6me23lOd
Qpn9LpYd6AR82to04nddUcGnr3tGsHi/qKmv4EpzHWp/9kxQfuwBNmfIPLQix8efdsIb2f4NtIFs
0gFWVSxRGMA9KGmR9nEFAUyCOb13RL/chgHXYEetyGQ+ix/zo6hbPiFE7ZdwS7AAFOiZwRXqb+2T
qhI1+wgwWSBNS3BS9nGstiD7MEs44M8mFuqukV/oVR8iee4mozvB9KB/JeqlRK1LqMGqQ+vIy4Mh
XNJqCovsUv2KLG/hed9hdNFX+xlC89m+EAR+wTGqm80u0NXS9NI/O4hHVVs0j8dO+1fJAKOTsUF6
11Z/uyf7IKftnGICr/W5682Ouo5YmBI9vrEu/973YYAdvUjLUWMNLAtfrRiMl3q3wAkKn35/C5zJ
gZ2n4M+EmOc6Vm3PXofaLLO0rkkkgDGQIPNxbYJIjSXGwK4ked7prUPkU70xegUs2ISV26XKLFLc
hX6kaL5axcf8xFTqGdmd5KUK1aeWqXIqw9nPw7uLS5jk6plzau6xqbI7VfWILmmLj0wpM96SznKj
MUSb4gogP5YrwUHRNYdUpysHhgIvC7BLyfMaIbws8+xYjDmYHl+71WWxVLnHCavMre+412mYRftI
axPC67RUlMtGRVnYnyNCLqeq4d59DmpmsvZi4JXcAmknFIQp+V3KXoZkDTHXirr0968WMpW1ErsI
8MOMt4owm1tcVD7Q/qXvgFuj2bpYcrXnVi3fhrBLCnwRtl0AsrM6MqjQB1qrsvd1vygg3+c+3JgN
XZSbzvHYxPjHzZDUXTFh1fAd7BGfFl4gY+jqMcYBPXiEHCI7MD2ywvpX1dYJAXhoYiaYe4YXni3l
HbZVpjEIJQFhn5QwZ0MHr9xfgiaB/4UKxQpnRkNw1ZY8CH9Kw+wxQREI+pqtayxaUHO396dttLUm
xTqRarhnNamNn5jXWtueHWxJE7kGKBo5BcWDJ1Pp92a9TlVogaurjtybp88eXqbM0yMWMk0Kpg2z
AsgLwkcbWwVjo849/Z/mw5zJaGpS0U2H8zgHaqwc/znaZPm140RAHhgSpMzL4ngs56NuQQnlkMGj
+poc6ZVQ0ZB3gMhk0fVLlTiw6fus1/GIvdxvk2nUB9XdwkRgIycC5MRPSf+SiBCtzkEe5bUr1hwL
pcb5GzRQzljcdiR1Ofj/fFpnAgLy0PZfDcoDYskQ2B8TrufCjxtYRr3jtowtLGBoiJyhCoRvX/iQ
wYHlIu6cqA8J5fY6QH2pw2ex+rm7ryKguj9LH95iCVED23wW3jbbXPOwNN0b+53ezN2drCKDKO6N
YG7vgXvLZU1es4M5k+YHqZst6NpJWUmRQghkO4pOuI/7lxF/IXuUCrS/ZgUDU2rPn/Y94iQ073x0
nmqrC0HddiGcj7C4uQR+VQMpzeuiTBx1/s1VXoKkmJx8KFs77FneGdRWwJpgmM/uFFuhPzWkPkMG
WCkYMwq53QzyzX5Q60BXHgrzVLpEMbgpO1bPPNdR8ZX2aQ6VKL4JOe1klFFlruOT2NGtMr+Ufjsh
MHz6wVt/agVTlgjPPgCpF9HP8ftrzUeCgXmg+gfsimEjWP/2D9hHNM30GRUV6fkxeP2iiZFWmxX2
tQAW2JgTc5Irm7adwXcaaGBRhA0ivHL4+J1IBmdscWqbv0noUTdiA8te+/qEVqf05MovyXtFAjfO
WE5ei91P3vOeJ5/o2FwkeJUnG2Puv1tIpsGGYlXAJ+p2ilo8VjA0VLRc/hzsOtzA/KE4+teY1ZD4
uqbF/btoxIqPK7PONKIZOkAJnYTh42ML+uDj/Juthw8Isv4X2z4GTcc5D7dMWm5dLUlCpnTKiqBu
ydXi1bGHp/t8b4Fv8x7VQeZ4pXwuKg2FOis6xFKW3BgMQ5s3kMcSDulfMTn9SUYisaMLmVAi/adC
bWvOcsa/bJA1wkqbz4hH90aHZNtoszUslcmCcijdsHkfgje/yk+V4qZy53JDAxr3nIww+6qeZ/0f
n6km/wv8NtFMGVp4948IsZAuhWfnj7nuQQ9Yy1mF2vUhecrTVDlrHk3+rr2GDblVk7QWWaICcLme
WEZsm7UXGzqa1wRDrB+RhI2gjVppf2d6cwWXmLOPRpZEBqjX671iGwV8IBklEHYZBwjD9gekQL4h
NuMfGDR72PSt0MEMRcCE6pTdCNznRGP+WcPiM/us86nuu9bX/J9i4ImKI4vvrc/xd78yJGTWh1EM
APSeJkPUHOiZ+cooTxOG3K7kKb/W98jvu3LIkB6icInLXv1QJb0RmBxMzvOKpA9lGjrb0wo4tJt3
IkSXzfLF/CTg4ibAZ7hV5yG+NjvXCkr+SY1PKR4YCjinAVh8odnrjzeKc3W7Ei3hj5EYeByFpPr0
cR2G00707wiS5OzotT0xWnwRthsRtOEufoP/4ounO/NkbXzUxiAWqm6+U7Eh1nx4Bpg9sUWsRVEX
gv77cKPk88iUV0eZIZ1SRV7v3+whGyHGlI7GRqDniA4QzO9cbjXDxEW2RQG3O6k4cAhmhXqnLk+e
C+KKyh1GVCQXlJUGsclSxO3WVX5KpbDvPaHueNsJ1op1WYQP5FYooV9pzQI+TJGJJSwDKR7yPlQL
0aXe46ldAZ5R+53fWMIglk9XP5ldhuladyHKGj1OQm8wB1zt6LjcNDgzBeOaweUoQx2bXr2SiFYp
MBNw/euFjXyWf22lGRKJu5tws7pu1wx9/mebQ4ykhPKjeCiiO71F7r7wYDGdS9KT35ajcYM2+mVh
cViSK4G6bNXAS4i4X9FxsG//yTO/7FyuyJpX4UBQVFrAZ6PUSoHs8evp+Gc0AlP0DuCnzZ9PYWcO
L22jMlasAAU3PEmUy45IlBzUSA8164VyOgYkaWWCwqjFrsiLFFV7B5l289OTRwU9OuWKCzh5DnGI
dbooi4BnMRQEaysaDigmZMj16X04bJhihKrRpvTuCcRvs3WLvCoZRs0UfLF1O+v87UHHNgy6y6J+
1b0g3SwU1il3rpf3dD6z1kg50JxbeWT2gczchrEniC+d2zQgmPzo9Yy1h950p6T8aGwY0GGbGLXA
VnVCGFg+nqdnAUx8C5kifyv66XvCCC8vzBpxv+ZJ28NGsgiTEiDVXFNknnx/mBxm0mLc7didLxQq
JsViEr1MGK4Hxdtl5j1r6ewpT3XTCWvOu06G9oQgshEWK/eXEsULvBrAXboYRWb/oHIDyaZiC63Q
7TgiuYV0Y1P9th6fvqGOefEud3zXkRTFUVm6IgDqEbx6n1esqhc9HSMqHJcEN0QRu/RYrOs6VJcF
vaMa7bJSUdZu5tJR7/OcfOApvA2Xv5PB/F4g0l+togxqytZz8NkEJ3ousK0UzzNvL+f4QU8DFuJf
y7ox/ghWx3erCehvk7quLFR5JWTmnwjf52mD1Pv0fhB93EWN6Kbd7yFuEatdgnDaB0cKTFwXLOS3
9jRHutH969B7QIwG7PhfeplxNx6tv9t0F6ySd7MM2vtIpGI/9IqD7ftxH5dYov5OsPXXjTyPcfwR
SsGFiFO2N5JGvrzsnoZ85ELOIWZmIwuB6vsdI7Jlh9bAqYijKNly+5LeIMMJsR8SLmPBbKJXHWgz
mvGVXlemvSrxEzTrkh394aNaP+csRbW+RSTOKSU+RWCCH0ofK+B8YgUlPt65cbNgLc5/knkcSV73
wC3qofhbkFLJ9jE24RTb3/isMY+j80o20KP8NFt0IhDZGJab3BMTTjT2Dh0SwabbC0KBF9b3RylT
vNf6skqzPDBVS3i+G6M8Cr7qgNen3BIR3iiFZEynbXGUeW9uq8Pep/AWcuGZiUcLNibVaM4d32JO
zPl4T4WQbFjt93i9puBAXEKosr0bCVj5jDgS5R7guTfJ2w1QSDLboKDTQv1zzSPa7Xzp2dkbjrZ2
H86ugNvFvLbAoa46geSMAWmS+BGg8U0lLe0Z14y6ejh7Z+UkIs9S//NqLGIJSvBMKwJ0Obd4pbBd
j2vaFt3W5VlCEq2q1C3OwhrJi63CO6lmKfh4rmNPqhxROT4XNA9roeVyZA64sltzJPkYvSo3RDSq
RROvQY534M043mm+PmEGmg+Zmqb4kUZ628mTZEjNKQPeE6sKxJdzpMz8cMI8nVSJW3zDSOPOPsPE
53pzeoioQAaflXSSCWbvE+NCTuDlKM8ot6weJhYGQ8ztV5N1r8ST+m5gWkNA3yShhuw7lW4Um/vG
TuIqQXIki0LN6gRZfjZFbY+kbfR552r2mfGiWJPbnLCB1XLlknya71DadyrjKzLmZtCqfwREzcLd
tTTlo99BWEPy6ZES4V5YTXuNuNrfaVeHTskqluMYYrycTbSpU269bw+m752ltwBpGDy9GkzgJKqs
L5nksRAdVWwGIntGmv/IPeoAUzFfOtAnwFKyUfEUj3J9hA4mrLnQFGTI8fGyAJ/Ba5NHzHdOAodb
i3KNZq7pl0XMLHwy532oK5AbpiyXTNh3w0JCOw22JahMr96U5CTu9bk0te3CWQhASMnwKE4oPlF/
zd6g7hI4tDLQkD5Ne7r1hznO1BdCLanNTzybLm8xW1ei02Bk2P5OTLxjn1mnOCR2wtUqpbPZ/jRn
3w+qJyFY0N57beMJmZFNA03gwl73dR1mnfhBPjMxeILCSmAvXwwyouULukjiMLlaiiyrlKF2mFJ5
5Tx0xNTDf3M/AcTK/bM7CK8XwP02Rv5NjZQSOjwfQKcUW9avDIcj8enqcfJ0XVLjwGR0w5Ktj9Km
oJ9EFsZf5q2OHrIgi9X39T8jjy1DJ309imd6rH6CLNmCPXwcU+59MPbiWJUl/ScojgLiVeL4ehH7
j6mL+s9CS8+ioJPbEF5EYj0b+1DQdINQMaP6NaDeHkoOeiuPCioUmsuh7kC6VzcQCzaGmm7RO8rI
J8Gfy9jCybRwuytfCFBOf+lUiLrmLBgUvDpqHIh++uoss4QzBrfaKT+VtDhH0VlEhojjYcbwBJ7C
svmSY2Vl9bAUnFcxvT3YReAS+XJ0gMhe6MzNhUTup9xT449+co60ivCNcdkpwrKiYhUYylLDtREw
Rq0E3F9hGjroAuTMKBf8rdWpEUD9V8x7rP89AfI4kdiuZ3VkLjvjh/ZCfir82+0wTDHJOqw7lHQC
C10D/6caUHrRq0iN0Cn03prGuwHm4bZYodu/H/YMCoRAMHigcdjU2NjcEuAO/uVEzisg9KcHcpxH
RV7Yh7Xvd/MUz52j3oZga6J8LwVdXAjnAILTfZ+6ZE+4rDLM0BMsKM59MBKU34oC/8dVQJGKVkjI
vIXQWPRMQYZXi9CUnIXBu2YUlDlFU+MCprg4A3mBMoAB2f3ke7y5nszl5DvjX7FquoiAp7xy/Lts
FYJjHWxzETp6lsW/cgzeeO89g9n3r6MzhBBSTpHUGKp8M42OnG2j0ynIzwGDjVFxHxRRS/mJWjft
RBvhuzzuH1t/4Tol8D50VnfmhodTh2420zGiBaf3uvbM2XEd6fCM7wMwtN0vdDVzLJPxez/lBhcH
840dblAuTubutNfrUzYGZwbXgCGGaLufo0QXEfHRfwaRVbkN6V5t1VTKpe3U0X5/ul9MpJgoRW6K
quLb0pdeeRayuxrGytRxYIp1sJME10TOTHVVpuvnXaUS/g9/BLP6Xy9hwl3upl9C/obblHRXNaR0
gXMrmaOS0X88tZY6twsvr+2cZuSvJ/IIwjFoUHxWo9GDsI8OeLrZF1CJ75J+O0lsfGdMkwpojyjv
NUm6Cbl5x/numwWCWOrWbfK9Yudf0ufBXVAY7dTm4uAl/Pf+tWJTxA9xJRnFi3BAFAL0WkGXNSPK
Bz9S0aSO9Wiq8HgjcfJ8aHugaSrrjGEliR3LjmX+XRi9SWMQwFjYZqNP6RhdI9weo/Anx3oqCMdQ
649LFMwL4HaL40sXFYWc/Lfnb4v4FqXNSYLbwVgNayXBfxUJeyZXoaNLuUjzw2vtyO8HcTHKBTgn
gkcfhm/mKBvbmtOSaatGw2k8hu5+G0rCQmjfqAcRMdUvqreHDkYppQE+/YXYvoDkHFfou6zp8h/i
4yFfEE6tarNJgtQzDIc3WktC8LWNV/2vZzSXAiwdu5yxCBWJMu0VI3VrAE+63TU3z0rrR9YhFYrM
tS+tzJ5/kuJ+qMbryZudXQF5ca7cWrSua0go8MTJLhWEiC9j9DPAFlxv1HOJEmevIafy5GxaxP0C
EAvf8dmbk0V7gPsKAA5FlALenW48bpjX+sUtidDDdvVBpMPGomIugRTB/MI8U5gWRh6UoLk+CmYe
64frsW4J63yjDl6/1o19tNDu7RK+K3UhXkpvkH8/BZTnZgp5drN7DExOJzKiDZbvBVVXfsE4RB7p
rOhbJu0Nr0RbF8Lv7ghflDtJJ4y5BdX0c1J3iM1JdJ3XV1x+hkaF1cMcAxj5l1WCRNXMoSAGTlJ1
1aK2zSVZ+QZUZ6nwOCz73hHxHm9gBEuFOv3/VaJezeoacdvPaJXFgGjpee1yg+hiE+i5Tj5GXqKV
SQyZYh3QFhRPg8tDJa/GAPd0XgsLhI42JRCqqi2W35t2K48eglUlC7Zk32ePqXEW7+rFLcdDxWR0
ugHqQDshNFIaKN3/qNAX4sMj3Hz/jVXpvwkaSulh3H5SS4JCEtONFblufEsj+O3ewYMGLiGE16dB
oj4BB5bt8mAglxlAT0kgmnvnyE5gr3cNBk9XgP5Jactdcqe0NH51Lf+AaqfSq6/10g5mW1HKo/zM
EUU12lkLTeZdbUFeQCBgtO+j0J6t3sKc+aOvYd2A5DjEPNKRp3PpnZ6qlGQgud6HonJX8HNRbZLK
MNrN40XH1cC0n5ZL5PljKlTGbTvBtkWPsRugfmN0PcjcsNL5I4YomUWb6XnbBPldgvJH5wGE5pYo
ynEVk+7Q2Sh6ZTEb8pKVrueuruyHcMnDdC3Bbkvw7bvEN2fiU27NUa1jJm2mi78ioqzFXRafvIlj
tURHG5hGO4KKz2dgk9tYir/CgPCpH2bFLtsZS+etS8Rzq785vsMCJIb4K/ZdKERZRUhBEe8dfvti
DD7KeAYWnS64WKuzhEjDL5k+hVOtFMRu8o7US7+pzaTHG3D9o5EmLx+lHrxzuWX9ef09pkYXutwf
y8/LiCgwf66bj5tQ9Iw0/ONYMfiy3Ffp/xX424EGZ2N4yHCaCTV9AFaZulNpnj+nJvz9fFWvw6PV
H7ak2riTMI4rlQGjDnE4YZoLuy+hZQauWChpaQk3TTCH6mD+5A9mqhWMHXbR8wAmdUL8QH2M8iPy
ogzdjJDXxu+4tG3Hk6omn0mhROEvT6SO/zKxZ55Zq+ctkKg9TLfxHuyOwViUdm4RXkd4X+elOcCs
IpOIu/4K1Jrjci47LtwTFbIDLf+IvpIioSYBgZO2oSKuRFnz3lzvedzoLEUPqZWMGOq9W38n/dlm
z3UNiBRcFT8iRI+MrwtSl1X6YdmnlqX0vYniADhXkSLuoawX1wxR9I7HV28qbpAEOKnkGktUgqpw
7Jv4V2tjnDEq3aFCYDYSQQUeELYFWkmG1a/mxHPM6HVw8nCACIqoWAPSTmdD5Rq58rIyWjKlcKXU
hq1tEMXbeN+C6HTmu+YOZTefTl3q6UJYeceD8+2bHqER+9ERpuBANf9xY2sSFfJxvypVazhBVm2N
lUq9NCrfdjmKqJy1kNCaErRjV9OhCu5j8tTobRxod2Q4XFKKYMjUR5KC3LEWthKwU1kvmma2C6Gb
5WdDd+ndn7u54ugqllx26KEbDPhVO7BtXB2vUTkWE6YsW1IXAyrPrTSkgjXghqGJwgeY+Yc40R2R
96XiPU0qpFqFvArPmFHtekOjc46uzroHZzANtO/NUQ74h4Hkswe19OOeyo1PvY021aWNO7Yo8UTz
oqsmjgv/VfrgZFUaqHDsRe4eag6UwcaguuZWrPQMXjdncIOoA/dRp7s7RyD27/rf8KNH9qw1c5WZ
llgjOR3KWBTc5KduocZQeXTuj07v/DkfaWqdXYGMXK40OrJlHfAxMR4aQmgyfHBgIsWERGJd4OTy
AovaRXyA4vslKB9i0bQuUSSfY5AZCY1EC7eaoL+K6+JYTq/9ZAmHfyOAyRmIgS0GVvPNepp2afuI
MqImCHnoCeq46sxGFg6Qd4ebLGl+v/DsH51VVHEs1CNuSX3admynXvz7RStHDJEDvxspF/ntmcFW
dOPJZKGf5dtKp3yaSul3FLP5Y7cjas40GytCGYv+1IyCZpztrehsTM9V28mSTQwqoMIlANG2zgc2
CxdL96FZkYUkDNupPs9DQm2Q3ozccYOs3p0rXctcBzDaq93mYvSV+BennJei+siZr+Q8nNt/uSxS
SbGtcoUonCM4u6DhxCeDdrypMXiXWLM799vMi1Kt2kbvyrbT9a7iwSiK8AOCQYg/t8xKUVNIgv7+
w7AD7jZJDfxlws6QGgYWooTJErYQL7tG/bUfbGZH5KDXKgeugho7MV4gPjYXFqQOC1iTkJDR2il0
Xg6GrAhfM6n1TjJemHmgMMueXiUBLu8v50ih301dHgEQVKpimnWCJ04ZKv64C6Q8UrrSdTKRnDj5
2UC8sLSL8sX5MMaMkkFxxatiA/OARfYw0MKWpKmXWlrRWziTAPrl19r+qpD5QorepYqprnVWegJR
ogI5V/lAaQ0yNaj+Nf8TaULNvUGr/1WzUs1Qi3/XpRJ0Xq7YZ5HjQEliUdUojRkBmj7VAmfN8CHN
5CNIwqJPN+ORm2Jdh6rlzB24Uzls7jBbfrvuBp10SVTNBjf0rdsiEyjc54VEhp4MHNUcOZJ+tVwJ
i+wzrOozXUNTfkKdFN18yBoRrlgFhnfH7JBBL6L03naSwnb7mDaytF4N8v4xUFtyjUuPJ2p/ruUk
BTWi4nE+z/MWJb/cJiBVVErVx0Cz/b041OIBSNPauDcIKSWoQ7H36p3yzzIvWfyJ87t7geNTQk4P
PXHUPCwrdClbYdWhrr+Vqx0PCbLIUG3OAo5FZzvdhmvYJ0EgJ7Bt1gdkZuuHKet1N5tECr2NZoTB
pMkgQlM48vt59+35Pr8cIkhpG12BhYnf/6tGNFdjhvFbc7KXYndGTzz327TuxY1qWRAjyautYvGN
uaRrxhMG+1MVLW5dz13FawPglTH/gbOB6npJlP6PjfENpK9L1fNNpgl4aCH0Ir4Koin9q4XtZwn1
xU1eSaqXOcZ1tdC0w4SC9ktviCJ7YIqg1abB6SBP9Mn3iMvn4GJAw09WATYVrToMrkLDftOEQWig
i/jTuMj5fyOzUE9w2Fgd1WdjlTzsjLGKu+ZqY9nazDOHyyosMfjjRdnStorMIzmuCNmRzdf9HDV6
1GCD9Rkcp3HPVX3UBjXfpdNAIR4v2K6qSruNuIstafH5cgMPHL4CQ18T6q3zWga0DjdZotB4v8wp
qoYcbKLx02FVWdfhrQrc78+dL14EREfGfHz/1mPbYZbubmEUEp8no+GtEBoJxHNvzQl/t1aMsmCm
xi67x3kWaYqV8gs5EYEoPxX4gT3LI16xcgZVJSpQbJZRNSd774Cvj3hLlPQM0FZ1SMdo6AE6FWsF
Ict+hZzjEg3RwpS+5EwizNz+8Oei1WIB0zBVfio4sM2spZ77eskufwWwLfs/j9URHsAFcESd+ykw
hawRrev6MTtu0IydEuvLd7HJbOhFWQSK2EkO3hBZqDr8MT7EBVNwgTZzyzVFIjuVF5c5W3ZwSEJp
DrWmE8ShHUNfJVHrMsgPpelplDvnDhr1L5fG3XbDk8Qc8DWtfo/WTqHfiR9FGjFgKJS83xZ8CdxA
h31/DdaW823yPpT7I+8qXcFANeDBo/5ZAo4e6qecDoxitqQmVDSYICt1+j7TBXKzxlOUF+BFzfxS
KCI6tKjniLW46GxpnKvJO1TRROOz5WttzEtjtBAW1jYMffRlMuUWJ3wo1dwchrKE93t4z7RkJZoQ
Ym61cRjwFAq+s/UQ9n7j8cWeVTNFMfdbsRNvH+9hkuEM+NuWFEWw+Fx5T75WehPUG8/u4MbPzrfo
uOs3G37U0GteiBqXxtwGbbF50LCwuuxjRhfjJM2N51eGPrpfcenG3P0b9XNBdO4ibZBJvkeX9bQ8
brdM6fK23mVFLJts2+j61lAeCGocaDRnRzr2L9n8oknGSrsDO32fUTPKFQhsb30jlKYcnSD5xkWh
5bg/KaRbg8r25SXf1sZiNuW/dm/8AskPzGmq1hPce6aQA9zfNJyGjU2LEBoiEIsJHKKDZjlSyyWV
lgv/dlU+dFgA9axm8Zl2wbnMoXUUO70mvJAVWbV1vSRVtRwjskO7kxlGnKlymGC0S+ummV4IgEpp
VBdb8mNikmy/D6X0CGcIguLz2Kn+MIZ0zOC7HthM5sVMDHize7EBNqxwy/5DTgERblzjjLvlFTKD
zt3M+E5dWozS0sGE1ewg9fFA60SxjiOlVDFo2J5ZdukahbPYf+7uymO6ROqp2xI6msel53wsiX6V
EJuDY5aYfBYEnynhD4ff8WfHQsugCtH2k32zVXuHk49Ic6K5/0zlaknvITb45pJOy1TE6rXZq5EG
cPh86ffYXMbmskobV3B6fWdiptS9sHCB5nKDr/eQZh03QajKKmzvrbQ2qBEDgaXLVovMMbFPNcuO
ic57/0DF+g1juuaVhbGiedoTw6UMKBiCiQqI3e8ZZ9uCk6lfR61FNmHV0w9B3y/d77yaGTo4tWot
aCmQDZ9Tm7iIomo+97Ngx8X6Tpz4ABK6WGggOrlqSA4qEKCOd2cs0BE3bB6TI5VIZ+WA1VKLhjXR
vitOZghS3VsguprHEZ8l1pPZyNfjTrEGHHF3xhIRqukykmYw7229UDom5EnHyaSQQDaWOKkqSGWn
pr2L4Ji7Po9QcnYScDZUm5uPZv5pqZvpZl0xUEG2BCZp0Z/wuHTdZ5kcs381TGjLLGF4zsDZGiBp
vVIWXd2LiAeoxgDPPfGXKgTsnboihUDaifO4GuZWfLMdd+NkJcxuu/aeVAfR+7KlqKUqLa4S85cG
WwkuJvvEO/2ylj/o589JvIniMtfINd8btpeRqrAwPcjGIZfToIKDOJK+Ne1eTde5/oHrWDAX1Pqm
I6qiljp9bjROq7WYIX/RKLiTLLIDCx/d2sWp9bsO/W7jQsIGgZTFwhNllitUIGvejzlI+pPCMw4J
DTereHYnYy2irLSde0NTUnUHgJFeXllioVjTZVg7SZb/BG/Y54pPja7wPrlZSABP/Bfqt7KysStd
7pL9ubwlXMhaBkhiqV2ezxfwyqWX5a+27gIBKVj2oTqH8wRPLiASlIY5JRNcwfV0HybUq5116YiF
SP6IwT57Wz4EFli42eenJaaCSECgZfj+iRs400pdADVWvWNvgHHjJVzYrpv0B/dRz7f/q9L2/OKB
W0jp3TeFsDafRAMYFsMfsjSqDDSeD+pKxFUpWUfu8q823FauUvvOa2KnICVdhzXiliPZBrLLb8Sz
/WBGyWVFjXC6TwRZYWbn8twwWCUcC8S+Fd3PRcMxBrwJwT5eNHdOCt3ve71hjbDqzat6P1PytUkd
8fGuiLkrySMRqnIhS9fmF5SZMpucgD5oHcAQMQb1vmIowZ5bhoXUOVGbhZ2gwiNSf/bgjM/0LCh6
i5nJdJAUnDSVjglXBW4vWnYPYcySnBmcflkXwpSbFHzEEFfckyYyXDT4FlTVHDuBO7vkV3c3BiQ2
CqbviJ2YLXHpo78ysr9LpA8q1LpjtWU4DGvHsEQf0IuSg3f+oY6VuKbIFhoNjpYPNBxHkVJ3EI2I
wjXqTZKwv9hOp1UBqu1ehzk4W5Ior7Z5jruHnqA1PRlFO+vpUe3Wbr2Dt9zy5CPZy/6J+j+y1w4g
7062qjR0y3Q+cWVVja+KHmGJdBbvSoze2xGASOBGXFw9xA26v2Gbila33dgJ9FhV8notCFgYkP7C
kT7Tw1fPWyLaGueFrq/VGPHki/4hcQYX4DfsQJAF0a0KAHV89q9jS44vi5k7J4MwZFk2QsIfxdtU
IOFTdcFiaBjv7jcxvZfz6rkvZefx0dMEcEtDgBwgbMKIcS3jtCXIcjpm3bjIZzxBSSsWJnBvfqVR
KQafAM/BX37GXbx0E2v74qfje2IRhBTx/XwyOy9bmNZgoTclkyI+mj5M3FtFYpP7L4nE2VjO+mK0
DKgv6CCSFsxTjrN4evJlCYVUcB2kL7qrWuL8qejYB/sOgqLapNOdsHqDIt0Y9C9KG95A6W76+uNq
ppcYTxzl1NW/WfWw1prptyWlnk2j/xnDwaHZeW987jGHMG4zXnkVLIysd6i/q3OuxystbTNWXssM
rcn33SSsRddIliC8XxsxiKclcPeyTnL0R6id61lhNYzwchiR/91AznFk7DxwW7eXdqz1gkQGkpf+
0uQV4c0JVcQRNmp1ECe3x1llq11IcjcOBp5amXdiRXrJDUBl0wRdUVeXfsMbI3rgAjSfCrEbNxfQ
yGcbLWxszpv6rDMlvH1At/p9bzpNYRKdkmcMEh3/aWTRgKqcPSWU4k/82+gVaewbXEtqitE6de//
KmLwro1IIYvASYzs+OKkBuVuE+QBgZnV7s9s99bNPmozKckr9v5Lm54e1U3I3YcTwAaKeu8sXB/H
tbV4AAFLUPA7tXTzUMpyZWq7eGNOWIaIt+w0Gm5DuQlu2noEulIeYkBAce0aZin0cwIu4NoXr4yj
iAgGANcveLOL0T6G5bC8Jt61hYNErBsfW8jKQNX3qm/yPRkqCALzlP4ObU1GjVOFIT+fd4dU4urB
bTGUc3T1jWs5+1yVqyNr93GYIm6wV19zsUnz3DXJVoR5r3A+ABqd8l7iZyvaE+2Mioha65/LG157
HXDbu2a6sktcFntzwZv71ia+9OHQMhB96Yx9sFeB2nSioC859FDw91Zjj4rOCo+DZ7v1XOO/N9dT
YKvEBkqmpJVLJj+1p13MZCLF90Nk0i1Pds+VGhFTg7suQUqLyV7Q16s2FnSdxru41d4prVGKvPQq
fcC5DfzTncq2f0yQcVLiAIMXkXVOPu4P6V+dOELAsZO0KQg7N3MFQsipcWSShZRIeECnwSdcTRxB
QjMZGBmsFY5darAPiGuTk6XfWvdGXoHBwNwlxrxnJYJn1dmIo+q3WK+OMQEpYSP1MrE0eLrgaIl1
jbMF9OFgL/U6PDHPewq5O/uTe2xbY83f4H5NGZ4/UetdIeGe1RKH0ZGHr8JxRFrOj2WoQe0sQAds
3/Nx7j6vc51WkHStRgzO9sOIAh+vi8QzoqJaEn9VyujHwDYEJmgK2qfKVBERI51ocLeGjOLNvvMr
w2WNwgCf0kn/BwueD+KE/Wc/QeNhd47co8NR4iu4ZqNYSFZKFixZRoTivIjdxi74Tb6620/6vobb
9d7YE5eWvWfo+FYGYcRaEbQKCfjwL93mDJI6WmS1zTw+7l041c77BAxQ05wcNKObpE+c6V0VKhrK
bU8yPTLfh7A2ZDrSBbstWLClp2YGojaWA07Rfynjc0xtpV0/fuMPBlU23/r5uiCBfIdYVu36pJBi
46QzoU5oXVDI6Q4h6scabZhr0QwTjiqJE1lnkwUvDCiolpAAmwxS9p88LW0vf56GSNmQQsaQmC8O
ljBgKUpsrh4VCobl5s3f4vKfLAv/FdB7vPyLzBRsHBUs2UgVCzt04yvusaBuEwI7mf2203DLh2Sf
wQ33Sg3NKPdlGLdn0uX4LFNeIuXStaBazAGRYDfPdbFZA8EgcZLDtSBVGZdBrffa+dAQIN+sC9Ba
Q+ZBP2aTN+Dmp/X2CNE57YH5w8M0TSKyXjctpx3/+xyuTTIUO4kjHtzyyyCWzUdWWIpskHrRIKEX
VU+s+7q761QXtWh8K6UcTHh/AGOnQRIIrQkPps44eMfXrmXTIDvpDKIht9bW/3g4fokVg9oGUR//
HB6t7npHDzqi774aEkVU0A27FT5CggSiwQ+SinIe5zXlw0aKTxomS8dAYlx5EOh1kUbMW3ajpHI1
K5xlFQJNimBRIcPuFVQjSXHIti/qrZ7bxddjxVJIZFMBlRXmaE5ob2CYeeNx/YaQI/HEXkk1ehX1
wiiGd+FqsoDQHsRRlyZbO4N6EZ9REfYSrSdo1R8ZRqPQ7jkGYX+u9TPtLSToLvr3vXz64NQKdX69
LoYakjiiDrnWEKIAV1tBPSrtwBqrTaVGyyLfnrzKnCpcysOnumb1FIL2RtHVQ8iJAwYPxVTFhw+W
BUOFTGPL36qZuIFqh9/Bg97PUQ+jJJYzHNXueBxJhZjQA5JxonpJClouc7cAwdQ8Ot06tJdeaqPF
/PhLyA69dsXVgzRtWSqAq+CARBc3aTYIZZ2RuhznbHaIsfLgMXZ219pQd7i/MoHdMUVxfANXtLvE
l3sPLj0mICudq8q68ZBorMR1epp1lkMQIiHZCGdGDxDMYpiOAkisowsEX2qM4/P3AowrP+3WwODG
PgnZ0z4hdhN1cI7BTMUlrwu62bY6YRaSCStetL3b3lP5OvgKECSPp70ZxcYvi4dSo9nboLT5L3zh
dF0k6BZy0Laewx9EWSBWd/hMN7b8HxY6eAzLzoR2nOfOqRgSVsWcKfLIRYF7aTLIbFhhE+Zm9OC3
kXgmIfclshIyivo4GidHkt2aDYtJgBp/Li9Lkc8R80pTPD1g0ECT29ekGyaIxiIkk858TdYdaUdL
l9XpjniAfyWtwezSCEhVPkEtzJQF1q7jXhXoyI0sMBy2aHKxX41l0ULaOPk1juMNtPm2yyd9WYFE
NrpFtThUOaN1usTq+G0CQsOpCzGnIVkcmXT/FUIrCQpKcxe7i0+DOi5fWHGiaTuUaqzRvD5FLWl0
6tGkDQ8IJMqZOo88KXujjgW0VZOSKIwAGHiMpKvFtvKIcE/JuPXELJ51PRtjUYqFTs2+x9lLsrs4
EUqb2ZO/2xexaO/lsHpBhHdxF/LGlbuXdNlYAUX2YgwUmqVTIbK6WO406oP1kQIuyZ3Iy3cGh/Uj
i2jmxn1BwbJRA1iL8aTeX/sXWCgoCO0QV+EN8e/KHDG28tJkd/oVqvmIuGSUMROamdTV4N4IYfF2
FxTO4iK33S4FDoNuwz4Hjy/seELtIYNU0p3xeWAi6kzxsVmi/TN5DnvkSi871sYiiP64/yFtFHWj
zzh9BDp+88V6hRvD/wh2LeDhTrh77eXtKg9x5YGORPC37AyjbQqSEeTXfwGPtKxFLbx6RzElE7mS
zuhrwSqFGxuaQtj5lashxRg22eomjMl07K1tvuIC3YRTR9b/XFAEWEL4r4UqBIqKMVZcF6OhKoIZ
knkTXt+Fl5W5kdbMgAZeC0CdPLi97/TBNmimXQbcDPk3bmz6jhzNJrVeMF5HO3JMz6JUHgfv+6Gj
Mgd+ExRsdZAFy/Wi4wj7e222lonL25YcG1dNWfW5EvnuVbf2g08xAM5Em4Zm7y+xF/lWGNjMicJi
w3PJrQ6N5pOur1b+Hw4lLQFnbcL+RFA84zvCxWHn6GynaYV8mYT/exUFtFO3n89ntTK2xLl6KXkJ
1GelI5FOosN77S+oax/fVIjlNqr0urf0NAlCo5/ZdjIThGt2GrVMmgCqCnh+jOXX0mEeUUDuwXuZ
PSl4phrsB/JG4isNrviQKxyPyHnFy6Nmks81NbtfbUV4NGSihu1Pzt5y4tG1JijTlS2Hhr0HVQBt
Ms6EBWkFzpt88nX8IIOVTU/lnge68+43ydQ+hu5D60AxkRrlS4Lxf0bEaMrtiPvXi/sXbKvO4A+c
3Kmb162EHpOI/j9O8DW2+PSQwh4moKPrNx7GoZhqjcwHivDQpxF+PjobLdAzv0zEWpgw/He/5l/j
a/eCqEYjXrC9kgOvYcaYuw7HpEKo4X8vUIgGElADkFAcCpFlaiL0QQ4oOBLUC3LlumzueSxUqbTl
WkaNIEPBxM8od7Tbym5KtYYn0oE2d/5+KPpPCAsSQjNOJwN4s/jrAoVN6LHZ2kXsql7BIa7fEtm7
yYhjrdTjlIqcJK1ygezY/rCmQoZtG57vY6K5dN/Ova9LIaVYujLy+ZPAOpl9DATN88JJDbV8ptVM
0FeIYJFxE8nubZ3QYyKqJ4i7C3z0jzyQH0aUgYyEJgTahFmDcOspfWM80/Vobt/YHsNIBdYIVA5j
DV0bBk+GNYp5+3wFemM5bJJEgsM1mtfNZMc2HDx0VsWrokmBaazeBX5rTnjB72rks106V6itqpzp
3KJFEIBZwVzLGbFH1Q2KeAMKYTqrnAewNTpKp18eFNEmZDxh4uR+tlUA73rpf7BmWdoGEnnLyZk5
HaWxD6OhE9vj0CUPSLCewYxPBfRNDPeze90MiGvRUFqV4WWvZCkKJAZs/CLhipkTVKrrcRrnogqU
uvnGh4/uLCel1rHDM6LeA6s8O0e09XKzwgj8ISI2YALsmktEoTS1tl0soObp0xup6NbdAyANOXJ8
8XPuWpGTXVd0ulIdv07LO9EqlSx4MmNcm2ZYH7PLmyltKFcC5vpLizyD+GEJMdWjPd+7Y6LbrpEM
D6w6sopUKn9ppLpSqaoGkY88OutpI67nEZ5x6wy4u/VgyjJ+nHsPZ966MnrYd7AJJiK4ckhlxgvM
sSgeBlt151Wmy0BwbeIW8SJAN8l1g9eipqNBUvhwo2uTJki4Yro/s12qa75FRKBHJSK7XgK6SUd2
00B4+imz1VCc5FyQt23yVkqMwzqLSeWBL3iqmswPQBjnrjq8stFAVoh/yqPHpPwYNFTC3w0VlOLU
uhWHxEcXQC7J3AEwwEiTBcj01IXfMtK1ztaEnaR0mTZsjD2xF2dMuKCtB5jmtmKv04CkYuyR1aNu
SRxvbxPID97x0Bzt791a6nTOO8nTDE30/juoH6PPdbuY/Pnjmqum4g40YjPOeVODVKAzhyqvoz0P
OgZM7KYPw782tbT/IXx8aJr+/9aiVN1sv5juCl2Ny4gD/FMbvx6sze59lX6JXyUmgoTGOFlEaWnh
m8DQQlmrZMQofKdmpreLYdJ1SQjAb2QktpFRTIjpzd/R/TIsVzFqSi2QnAwIl+RK1ZAVHxuQj0Fq
hKxsMu87WTHsP2eBpwlRDjWVfpCYZAgwHxKh/h/Nc47qGqhNisQVymKI+/t+nXOzWDbz0+N5I03m
B58ybyEAPUrTGIv3HnCN9sXtua65Si6undyJCcIzseeHYJccxonqNUArrUwX5h9RQA01Jyf0uNoD
hdKTgIJAxhZqsPH7PNJ9GV82idJyKKPKJd39WPIS5bAz8lels8C1rj43/DFQ2K0k5WbMsdHuAWUA
cC5Rc0yD2MfOQuFtHNutmnooyaC2r2UmyHBTbkj8OgR0TMEWEDzN7q/tiWHPk+1u8sAAm3YuB5Gm
KkZ+ZKZJKO5bdrSvsE0g89nN2nPLVYN1ZIw/chE4Oxy2SknjvD4xWrb3zQZB4JYYZxAuq5YqO5RE
4h77bHR5+3RDhIXZriZEPMCoTmf4gX9y0A+sH/SiY7ac/0Vba+Le5OnvXTI5RC/mugvt3H7dHlvY
m2p5t66ETUzo/gyNIiNqjFVPwWZrQV4B9ugC65p6FYwQOtZa4qx3fOhlReuWYxB2dlic3pbqyEa+
OI4cLJrsxQ9jc/K0ZZFR5LD2fMsX4RPORtNuirdSWDIfGWETwkFDf3aNuqwKxOLP9bEemGrqMGe9
dN7E6Xk06GvJzEgzQjzjQNSZP1oP/AoIMtaFE6h/ODL9eXvfAzhHF1tQHac53FHLLDIev6TQiRgc
HEupZUN1VhO17LO2yJb7qkaD66zlgV6Bw4kn5SCAQYZE+ZajqFS8UUzd7Cfut8lKMoYM+PctVgsH
ikyfPMW/fDmVKu7kBRYHeoYuYjRi6/YwWEi7f/ackfE0Z8Z2PUXyLX5pEyKMPbZBZH0FU4fk90AM
ZfcKwI9zV/wGulfzeQkSmkL2gyKj+C7SdliQqWdFTFBXeBRJMckvoSf6iy1El7AcZviiV+t8OoIi
GoPULEOlQ+fsQojZtlg8cGKz+M4eOkPkbAL55eZlTjt7dsCf7O9T0GxWQg6XPK9UFJFawUmtajur
B1rZqTuG7bux4xrvX9n23vmHI4yjk361WJqFuCz3Yv9hQqbJob/vxxw9JkP8+ET29nReHZNTCem2
2+WPEHYzQ4dCTqiiZRDj+Q7SDO5VQmk3zcLqpDs+c1WyWC+ErtFZP+LW+I5jYCFyIXkJQyx64UG1
8OqsvoFq6b/WG0QPqF5vDIBxIk4a3zOetu6qK/eqOhCrO21k7/bCYrN06jLAnr9GlBHeRPA+HQ75
RND1Cns7S8M7Thh8H/KDI7noCgw860wpCo2eRePYp820T30SkneWceF/qJmEnCkPAeP8QsasTCqV
o2UTVB1Di8BQbpSEKuP99SNiz3UUPPEEdhNwSL2wbfrJwKXhQyKD5Q1oBsCUCBquCiKHM9zY+Zku
uADwxtxShQPITBSH98kL1oAMfv6RYzPQbYZ4SG35s5SJbFkiR8XqVPXgbb5APAzOHxFR6mexmESt
IVZQg18PwbltaVpwdVP8qbHzF/1dZVISbHcEZ/OUTlIQycK5PMD95L3m2/altLDh8lpayJtbl0pw
EQZ87o7pCEFT0ZOC2WJSwo8G5zKGnBBI5jOFC8NEidk+9bJX8PwM0N+TngxGaOrHM1ZZlZLNfL4q
F8lpFEVq3QqgdRcj5+32HgUFCLpXt2Xj5bcu0oATRyAZNDxUJRlTmcF9F7ZCPB+SzWxkAt+GBw6e
KVpVCWdBSPyWVrsWeL+RXelEl04g0F9Tz/drYVVF2rspJK80r/qK2rvyxfxb/RzMx5zq//DqV/Ur
V2gzZx0G/u+o5/axDrp0Srp4+bJdrqgKxWIFQ6DCQC4cDOP8QZOuVDaUf0UTJIzXw0sYjfNJ61NJ
yxyhextrPb/We84dc91qD6q0trSpFYhBscV+E4Nk3gau9b7Pej+7IYI5GltnlEGEwaj/f+RFIWUI
SgAwJV2w0rh2UhalI/XAr+Of15KO6IvIHtVyW6DmvHnw5ier+jkWFVcElyW36HqTB2M4nLVVR6p0
u+ksEZAUqqoJIK9GJQ0+3UrTcGlG20WrFKy5LRHvN5klAhREOtwzee3zcw2KCqH3r0i32hyu2vvE
OVzx6eUFoEE4QfF7zqJz8lXxslSnYYj4y8BrkG58zrcpR8I6kjxJf46TgW88ZIZrxdsIJ+uzYrkt
0PXOf/So6IPVXd0K8CeXrBRnKpxn/2Tx/wvZ2QOtM/WzuhQxN6mxo+DG/U+qrupvX4ngViqq19hE
TWFqnQ5uiBnk8d6ztoZIotQWWd1M8oxXjPdcMCv1ZDOHK4jqUnzF6RqYm+uXp/FjqUu5dUqZANpf
OasZ7nrhk1hdG+9JKRCxjkyWYtKvFOFRsXYJMDp8F8KwIbhUwvu+2YET3AdNyNDCyb8DEKzQrS/s
6cKDuezD3dYH1qEGqxq9RZnRMGfEbZcJJa3iuTzsNdXtd6h7HXg147IKx0WjAH+ExrzmsGhplJ3Z
34GXgLMY8jShe/CjGfG4RSeOOmgI6FjhLrhV87lhXhVLyXEeOS5vHirsaHk/Ssm2yWIFifa7jH1W
VNBCYAnDk44gautjU79umsAjDhIulVRwNbLqkUQVnkzY9jzdo+dQkoIiGfDKBgmX9OJs8rdzlfk/
a0EM1XOuvg4ZLk/13MoP5Nxe6HReH3b7AV2ePL7Cjmo9jVL0gT1K8ZQ7Ra4UjCyBO0Vcfr39bMOy
d2QxhClWDU7L6BkkW3k/2L/d2aMJGef/76h5H+tzQ50idnglQUZ8cKtrt1bKexbXaD8uUwctxrKJ
RCBS/R1AN42PxPkJ1RQ0aJZb9aUg7C73I7ZPC7kICfW8JaX+H/Dk03WrO6gWkmcdXIA7QpUvqXV2
m/tzjGWugqUjYomlO1ZJGqGxg2E2TZsB4cKC0xtQ7ZTEpKS/WiAty3+3zX08ZJOotfrAWH149nYh
XIARWAGc1iQa6Ul7qn3ChombQwmEHUpQX4jmanhouPtAHuUCjnHFFAfkMjkc7k4Zm83wlzAbPmUN
hs4Hs1OOhbEI/oUBnnu/vp8bgeCsKcaFNspFUZ+h6BOzikOA9eRx5dodyTLNIORrEyryj8k63lp2
CXalHFsG21PlObdTsUlZeSFT/uA8ggkhwv57uJjnaggw3om9emwSVncpYxMDi88lRZo5kObYL8I0
8uauDUmD71zZpbaPttkq8r7dxI1Z+VyKYZT5dS9mjJP/WUenXu1JpOZVRhvWTnh5P7vtVUi06MRf
4pU8C7xPzt6SybBs8nEpxV2gf7F8LaxAloiQLuEH3SOKvJ3xIF7u4Tm22+QWrpFyL3ZMaXyn4c3o
a45DoKzunxZ0bkpwnA6MwYRYlf3P5Jd6G4pPSJPJrbTU4E8r8NRfdyzu2ROrk42ZixLvs3ksKa4y
5zTuFhgzsw8SgF9ZUZbEMdVIrjuqnP34GQVymSQjYWy7LGeOaOzyEMhpHbk4g82O17irbqunuZbR
GcH2s4JCCvZBweMU+98PSiJEXkLsCY2fa95VN4HBRL0vLMoV8r7HrgHB7wn0qQ/lLjEIepki/do0
nbhZqFB9CSpYZo9gnxfSGwFUlFWL7n1lF896Vplhd7nFNI98vcmgoDVxCTd897LFUEkTKda5IPre
FE1BWJB4W+uDANAkWFRPkWxnydalyVl7x6xn7qfURLlWEUMZnwyglDRiFIGJkYPteE2WkXK8NhDA
h1Ik0nhayJcPcj+xm4ica/TD3LMj9aUUS020DIdRw+NcLPBv00TaaXwkoNFcv3ZZdK+UQH9ZNxn3
aCIYRylET0h+pocIkZc/cobsymMiAu0feQXPhHnF5ZS6gAb6Oh3/8JZnrLXw9TtQL4m04osAyVzI
ewRnUSbJkFeKwT81gf+i/7/2a8Oj7P6zli45JWGichz5gvPcf2+r1qCXyK7U2fxYTTZ7xuGgQI+Q
NC3Vraacg5HAghLWnlK76B4Hmr14n2leqODWU9M45XGYhX74zWRjMzdzY7a07OWL3rYLt6ix8cx0
miZCnbyFTNDMvUavZiWXKftXQA7Q2ITRoZ8smuyA9vua8WQKFVIEGNBSsMD7AVxalxkNTjmJ0m9k
9ON+6s8z163c9VnGFsr8nR/cD8h1k5tDTsPnJiK9i0hFb9+BevMTwugNCtqF1wPjwwZZTDiEs6zE
pW5qCluUsa+keRd8r1MaJ0JO/EC+U5lgT6ARdWU9qMh1qL+o5pOE87NJwoV4pa0Z9YxkghXBK2Aj
sGNm9J68e+w7C6cG7GnJFEsniEiPtOoI89BI4AxeKKGSKzrMUY8q7CMuSObggSEjHBr7zlE84Ety
HtWVlTclajkANLNZO2KWN93pKVkG/PnmYFgBtaWSMgpyVIecvBlbc6fV1ITocXf+nZK4v0pnTqSG
2uojxIoR13vU/8HFl4xvNaicOIzJMPsjLjMEGLfkSFV+ez3VmxwAFeO4d3jF8uk17Syf2+1vAINb
h7akGYSm4zJ74vjHgeOhpK/xtCCdFE44qtd4n1g8+D4uxPkZkq9x9UCzZg2wdgvF5myMKdU4At5u
CafKFa5fvQgwrM5Axp5i/Da2kVmcNHEjvTh8qDwizME2ioadmOEtwPIKdrHFkRZxFHQZT7Xrv7cU
T0JpcoTNjYESZtaJ/9eoU7emCIVnNY10iEvl7DAuWGYOVVTm1JtVQRX3cWQ+7sPSdvgPKESmtoIH
mjd/4zZ/C1sv96v19t4GH+khCtv4GCB3WoZSmRBzW89acue4B/nUlBO4gY/3cSboJ0+gAy9vWjUw
icjwUB20cq9ow1TdgbZYS0GiLB+vSFK+HDGD/GOe22K6pIspH8ZZ595k+gwqg3nuCCFwHkA2JP77
6uMKNOYjDc8pXwPP8ltviSy4EYCp5Pi+k/FuaiCW53F/GItdzMOYffluAH0gXGW6jq2LdzxraMiE
p2WsylPjNzPcwawf0yjThGRGBFW5QJUn90m6mvOnnvNNBxHdxDQnQFW+0uzQJyU8ElIiFmbVthTp
UXJqPQ7t2TeTbS4SRueCuxgB6+AgOKFiB/c7IylBo/zsxWncREv3g5n+wlu2SmSpRtLF2q0lb5oC
T7elBFWFhp6b5p41BO4N5iJZDt+qZ9/qZ1BV5J7JoDXkP5VHeGpgxMFma+0O8R657Rh+W9dMa7aF
alv2CrU7qJ8Dq4/yORgScGyfXRI9akfTlkiFQqjARacxoRL95rb1eWQ5q6C1QFByYHkuIl5ojVzB
4zwM0AZKHU8EOXs7gcbX1MHsd8vmfPHvAEwkDGkdCVsHIFIl1QsEsFGyEkHzCXgWElpRDyl81VAO
7CUawGoDJBzXWWQ2fUwvq+4WJUnkqQjQYF2f2Qk3lPCk5o3w8dbPjbB6ZFCVJQqIHc7KpsMLuxwa
maOnbkCp7JhjmZrDnnnyOExpXYEG3U6UNicB8aEvDSXjZUBLbTaBFVVZyNJMCTcWNvJmMzC3Gl5X
9uuNAZWhpN2JcOvugapD2GD6J/nraaWW5A/xQzYkJh+gfLbcVVKAgrj+oG4VBAPN3JIiOzmsY+ao
Crcvn5u6hWsAvPG/rknFiGbWI1ChljBeLy14TxAA/52hsr9kKgk2PvLL8jVuecEKIcnMhgha0uld
PIhKneCYR3+JqoDU5Bk2KLzpAQscGiIs7pQ0Z7WL5br7K4Su/5cxi1NVhAQDi40DlgqvlSWRA2vR
d+wO9vpt9rM2Ob/hq6bf2IXT/uKPxLHycCpnWFaBcoVX5zXU5s57NPaLo/bLmhoxyePki8oJ1N/S
M81BS6kUPe4/UoMmWisKiEYywn9cMs9hBOWUF58ecsZC/pNOVTUstYUA+WupigYJjJUFphKjY3NJ
hjamBIVNuPP/hYChfLhF/Nt+mzQR6HPqZQmIU9Jpd0nw+6efZAs8KYUgflcvn4A8v1xBoctrgIdB
x79nhfxrGjbIctZdRPyLWfeg/Re22xQ9/E0PJVaOIQ79lVmZNFJO2jNFvF19NjHAOZC5Ag7bhmgD
fllQbbzqyMwca+b/0XgFPFqUP90+EAtMtAcVJRSFr1Hji6pTCVB73uEy1J3AuLZIbo5M5kgeadAX
ii2Xw1f/vhU583Uf/7LzFdv9liiZM6KqQ9mIo9YSOKAVFwWxDqcy/BbvEIIDHmXjfJT87LLJK9QD
M83N4XUOuPHy0CwGXY1Tr7B4aXLrG+SnXfXVtRffgKMmL7FvLxnDWZj7kzsprP1jraOBkHvXBlGE
gnTj2UxVpYRDitKU51NHO1OLWERV52coIqqqDNbFecExerFl6FlYYifBHf/HC1saN4ENbnun1Z6V
blTp0mUdnNC0MnYVrTb1iqiYwevi4uoHDSEbayx6EKsFRDM6c16ixTb96YJysMDW0aN50lkTEBXp
VUJtFMlVuc1TqwJL6kIrtF+Okr9kW6ci/2rNhh8Gx6+7xVw2MThyK7P9A2FIEG/GpZgUNG6/Pizy
QSeElPGX/MX3EET3QBAmgY6fP54UiLvdbdbP2x35Wjs2eA3bEdJ9NECRLEP8EJuNtBJfDmXcGA4t
Qz1xqkcfpQOEq2jYkZs89Ay/eW4vOPlYI6MlR63ujXTVaZ33An3T3CmBVukdH4ufR3p99ow/jbRK
hsF5as1b4hKWGVvAPTR26naSO18iQAa2JnaIBsw5mvOlhY/lkAVvx1y6z9jnV4tsIpIVzWjdGpKP
GOEs7icIUbsFkACLwJPJ/42FYCCuy8mCfazpK3ZAqfBDucugsyST+gTu1MvWgdIASea8/NoUgY1n
NAGJXTG4pzqnCdRrmmcxuE5M1fGdKgiqhviedF9I/MrJANoZaeFwi9gxHfqczeYYKw1uozHiQILW
CGZZt9Qocgqb5hr+ko1AKHmGF9eh54fw0JiuKisON/gnDCXcUgd5ASkeAW+egxgHgQd/1d6YAQ7l
EFdooEKrDaAwRBZEK8J6gdqGDR9yCVdQFVLAJK2LMTEmBrLyNORwmRgxOfzHYYOiIbQG/LBa5A/i
9OtWGSyFQG9v2c1LS+xcMRNrjkmmllgg8nEeZi1wNmt+C2zYyK6jBDkHxuTVE8tQc/9VgNbjuICi
30mq+RDHUu4XLe/YIF0IFiG5+GomdRHpy3SAgb/q3riJzwWcBkxjSL2v+s9wnudtdqPDLSwWynav
q9JftmliVrlG+yfoc9QAcnunmkr5f1Nd9UBcO7hIFo7dOeUnRYX8al4jl/ODRDzzuc4M7gJOeXGD
7HDPn9Hj6gDBumMhB+kw7xZMm3+wqduR/G4+WVJ/6N5zmsNLPZqUSj09Y1D1tL3r3IpUFBT4op5l
Q78rPWxdtfUszFS8eJDW8vtZJcu0YFzWi9L7VfS0mLjJhDJdeBlfNc9VkKONMEoq3LV6mVx+wDE5
xRVRcEgb8eL3Yjvy4vYl8idwnRQhFZNu0o3lNOXB5uNR0NZEaVgPqfl6qi/iBAVzf1LdCRtjC/ru
glv8FKKTpxhTFsxt8/V6rb0Dz22CTBCbegO1265PdJ1tCaHNlBW+vZLZ/1X2Bbx7fEh7aYTsUccQ
V/01tPmACEjaB2ujPwe6GEdrYiPaOkcLDNxpIBUKnocvngHDNVaOT/4syoUmR1Efon7R3TZcgDI9
+1ulZsDCIaI0oaQ4l6Dvj+Bac/UUGb9ITtS8ckJDBRESnfNjZEuKyUSj+cj4KOpS/EivCNdt8Jty
TdyQWBRo6cWd8woBq+q8wJSnfQzsvJa6v4Zx7FHbDWtOxZZtqV1hT6fRc4xv1Jr9eGRmyr4l9XNn
yHaJKtoaGyJz4j+D57OJjPPaEUQECAw2dUB9aCZRjnKsC1n1nAVeQHxqnz/W27SBnpGbPeENOpn+
n3swWM9962ENDmMimrmvSSCd/3ik7+F5kgUpHQEjfHv54LlWNhxwWWdZwpvIS2+gJRETNPf5ZLh/
O9oLKfzqPInInB03mcWsWpasCEpEAL2OJoh04FdOYNIAEDcU4/kg0gMw
`protect end_protected

