

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g7azmhtm6FcP7uNFjuXJjN8Z6yccOPk3SSjzvKB27peFKmnPmQmov5+YTGwYqqN9LpdyiUExk8K6
vPnJqontvQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MFrqn2K0Cr7TmQ5al162oDGiY83d+AkTWOgFyXPYrTNznygR/tx44RAp24ytphNK9p6shs2EFMg/
Qqz0l8DCWiVEoJ/T8vMpnAn7Y+poGVGS1qAR3qE2njrl81VcGBZJeFaWIudhfr/DLTuuf2T/dWDU
YpelM3KbfYNPPiPy8PU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FZca5XZouG+/BYoQ8qrJTmnJanku4IprIWRkO6VciHehE5WehR0wsZJhfKlqLEeY1oTPA4bXaxmY
NjYkrop4EOwW8t47/hj2kFLI1OKUAE/TAhCGg/aNSOViUbB3dUomG/y+TBuDt9L6g0Arj1vb/5Pt
IChc5ZdEfRr1lJMTpFfP+5qmEH6lePPdzgPZATPB4Zrj0P6EyiEsU1FKBuAKd9iYNGiLCxVomaz0
3/RwK2Nl+/l4mc7PJt5Hso+4s1qHb4s2wD+OgbIwdH26ZkEnKVFpaLiuWQKu9uhDLGnsBMPf7XDE
p29f+mrvP9Zi/3nonA2aBKrTwR7XuH+ZYoakxA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jP68OjlYJglq3zpmKrXOhq7Sex8XNW8fQKp4hUNmuw06OOoKhQASNTnjtyVjAIk/VXb64ViBu1ds
cNMJybDSWBhnChfJq4h9PNybShGJXxSm3NDOo5wUHKf10Eti3fSotB9rVks+tNdTEZo4O97kgfdD
G1FNOqlsYcQiShEGLLiEQ2yYtgJBxJ+jc8mFjIEfPhAYy1ElrvtFEpnhkNS2LfE7xdWOQdO/XoKK
ibeY08pgncTI3pvO6TMbXushf0AX2S7hgfk8ysZrT+0gktqFrJnyR6oljS6VVPLtRNW2vo/cC8XQ
Bzvwwt4cpSo5KLS4XxB6qClZipItck2AUEdIbQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o7jAZIoXlFbFtDYmtXhfRBlb07dhBb6Wp03mlT4T0FXtvccSHWhWZgc+VUNwt6TohLihOwvSipPP
XVXpGL4pUVYNdQBCVpFzhMkt6jhyUgsF5t10yI5Of6YEfQrDHigceoBukM3+/zJHPprrPQE6FUvC
wXSGhBCXnHJs1R+n4l0714w8/WftPQhlD9QGQp1qT2VARQXUKBRxcRjxe9TcLfs0P4xnN7uHu0R6
JTmV+MHmhGpetSZGx+B2Wa1MQofUPURqwE70IwBoUhdXH8+39DT5I6x2+wMY6RcVATnhNd2BCgPd
RzAhwfrcqRiU9aB+eNNdFR8ve9M2nGMmV2JxZg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cl1Dz+fZIDYEIQuUd0pSg+5jknmtX/JERd+yOZ2SRaVra/4pU/eCTjEXMzhz4VFGYB6dgUxMsGBk
nL2WNdn/uaSPpi6mNF0UHQvZik4pUkYPrnRbFveVqW8i1t95SG0RW96uD19206lWrp5U1lqc4fH7
sfKHi8ZpU3MAg0DOO0E=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Qqp76m2aV9ue8Qai7QUavb+lhRYdu/txrnwYLzwTe0vS0S2OD1vxr8VeIT3bF/ZuXlTGm4S/UCSF
bgOPp7VqEOeGNfsSPK+VpQ+foQMENCQYccwKquBDSg/sLjpPK9uuoGLBLxjw2OwsRzplVFXiPcRN
LYK1/FmCP7RJBNgmhh/ti99a+WSl6i2YIIRGocNplQlG8FXq8ZTTHd/x2Gtdf/zGvJOy/fNsos6S
Oq9yJ0rMmbGeWbri5c04gZM08pUmXBsivgOHm2IVEZZFM4SBqrsi0xa52hs2kelc3iKJcWiTvU3X
0fJP9qNFuIjXBPPZvEYwhVtIh6DwiIC2viSscQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
x4pekOA/YtnPkzJ/Rym18Ag1vHoYU0osfAvloYnIeBx0tOIYOv3MsmYyToIhgAZRqE0U+iz4s5dy
spxsTlRO0ebZyGCIu1hUoE2ZiBWwMqqC8lVd8A22IixafNsy1YzINYT+aCp4YLFfm48W5Cuvo1cl
ANMFA6Iso0V74/qM24l667SXeDq26iVLrS7oEvuFCSPYqWzVW28vbeZGhAaurBFt/FzWTZRfHMS8
cWpjHmXqoTe4XDMovEw6hwwB5yrPcYxQwcnhnU1lWT+MPlGf/c9wCYUdjKZdXYsb8QxSkvBnr2yw
eWVYlxMwmjS4vJOPyJik6Cr9fyHSLYOhCZVK9A0/7zLJjkRw8/gdh/xIubq3tr1q1uZjns5XyjE8
ou0Q1uPWleXAXypqQmRDA/z0RWd5e7JR57bthp46CluGOJ2wFnfcdsWEd5IcoNV7fEhFd6Ly9WG3
oTjZMVmq9bihjgN/pOhmW3+26CET3agVlqNlzse2sLtOdwh+SmLfXKLIV4WBJikOLvKUrXZJTMU9
8JFB7hMEGHi+OekkxZRIRA7SYmD+ZkCFlsSO1u4GzL74PPehNRkDoxH9nwI2wSo+Gdu/EOaIapA3
L8k7+iDp7NAWAWfsxttdkswiyzFgXWeJOui0n7uW+UIjCRgQ7eJWy3TABwN2ukMb1i3m59c3fNeh
2WAbBjmlXTGhkAsC+ca31bmdbKVoR442C5MlF2HuXcHnXfPCG49z29hpOK7KmIFcyP7SliDa/K7c
8S3QNjDBLvFHOyqN5LceWkdi1DmpZbU9Ukq35JHEeispY0QKnqP44cjxjulPgdb8CdlN2Rbxro6R
Vsj2T/JnQrjASeEHooTM8A4A/Pf5xei9qmxVZDQG+73E7DisnjADNRgFQoK1fIi1JXOyBkdHGb2O
j+M1BXovigAUpCJQ/bjQYGu3hc9kkc29d2A0HDkSyg+a4IAvVO5IZUWiLFVCiJHlJEaCTam8vikI
kJZlwVRq2Dv/spnk12uXjSoDVunZ5jl7D/G7TkWgqzIe2N15hN4y8SabyD+UWJoXiIRLsXuiQy9M
Ns7FkKSzm4hznchT/RWJQmotYv7TbYqRhV57U3gefxDmXZO+4ySZhGHwTFlQsJbnqAf3LDKO6pYg
ceXJ+SBzpoz0ZvhPcCJ4Gdv+WyAGCLK1sGfiY+PWAKeGBgwoG+xGiwGXfW/2KA8QdF5fS385Earm
pBvP4MTPCBTSPyPCTemakXR+JxdxKYvrCWs8W2a78fvrAZEanbuVCYedKsaaqMN5pRA/naSg6rov
OzN3yDRyJ35qXfQpGvDYtnP07Ans79o0xfomDBo8Qc/HiHDBh1WKzGMjW9SSLNpGBE0xQDGhkDfT
FwvZ+a0USpxrF61u00Sw3ZlE4NsPmnF5xPa05YpORtSV+RBrTAoS6pznO7mdl04LY+rMldiEnyNr
HNQRhrYyU+/QrrkYfBp684ad71cR+b65z55vmLbTFoJx5sqkArYdcaA73oKE3ZXiWwcyXo3JQMRV
kotkkTR5ZPttGUJ7C5TlOtOw/EegzXJN6U2hfqMecTE/zOUtSl0bfBur79rS09USRdIGKPMSPotw
mscQxO6w+sBjeBrJktRZyCjJiH9vKsBJmWzXZyay11iDHmdmJwAM1oEBnhTAZfK0JC/dnayEAGK5
lQVFXhSu4hRMcNNJtEaP/5atD5c1Kh0b8Usw/CWroTiCSmVjxc5vHudH/KMeOm+CTCg2leVqy6FP
blPfPtmvdHenORz86FJTOUoNvYnynUE4ZypuHYGsbKZNSJWOVbVlubtYEBZz83pt4tuP/SRQigTE
ucYAMz9chkSFjoBb+M9I6B+wV0X3S4h+VesMsActJv3xr94YesKI2IbKLEjN7BeS/wvfWlmfARMt
8tR3yn5CRdXlyvjWBHDNeYOV4fPh7lRLUe95REzWi+t86OcBhwpVZ/Z2sI6pzFKkMcjmuPbnJPKG
13xzwE9H3yos+kCOU4h4PeOjrOSFgf5Wj+NBKluuigITR642vD167EIC33XJiuZqHi1GNavdm69V
jYt2xBceOsng9bEm1x1wXehXHvh7U7pKB5AcVRVq5EJrYahwbgVuxnDRfbl96i6bBKgAoAlmmzeM
24+f0G5aZvqahP02qza7NoABMdGf4SyG2xbrKlNk/91Y/FR1qzxC9h9woyq8rVWARTPqNdISaFPg
HsrIIthd5E47Lznhiq22RnuOnT7H42mGarA6Yx2Y+ZFOfYHwsVu8l2xNTCNLkGg61AltxHnTODD8
I/o8wbXBruxtnFx9CNmUwwPZ+j9fC/OTpkvutenSjuAEVz6cuedhwRAN9V11s86yNjmXLd8WTLO7
1Mgvzosy3WxEyE/idbPfHwcrpif2FeZhMclXWtnCoQcGrll7SoqgRxGz93i9FgUAMTAZWhN1myCk
Yt5cAfyffTev0KQAZ7pCb3+YAdD0kA3QSweyYaS34+luY/J/Ejbr0wFDcWN8ZHYhvMOgG6AcjGW8
jkImfVCHTa3edfPsmmlQMtl40n8Bm4xHy98S0yU7xYWPlLU/NJ+2E/P4erB/Oxz+dJDzYwfIT8RE
LwbXWh8BIjG6Vz3ittZWXKgKwt3Nbtb1cYkaShSP5zke0oI4O+m3XsFETLE0DtYRzI5I/g0Gxs8S
v4QAi8R7NzEC48ZQNKkZnjMbTyAVa/cNzDdzfXrCBnbtDG9VDtY0GIHKCoYtnc2vrPxancmADdK4
oxw2QpOUWYtMhkomd1omtKwYDJk7RRtIC5mMbn9BBwYNBLMjogvwhZ2PzlQHSWrG+fT4jlmCA+He
jMIRgT6/nWWZVmY4Adi4VHxL4jdQad96HEk/TEIO07ZdrY3lcOqU30DZ+S4zMcRZw4URwELJQ97b
iLqe8D6tGpGpdQTvuJXomAHhEUWDT/yio3qmMWTGHRlJLrDqQuvzVEwzqB5EFV0j7AvD/xH+4+lP
4VIokJkARBo2s1dyVN9q/jdYwaHMJE2BkbjpH1TldpgtDXLPsyYoVv8gvEoM3wBKd5vzPM5z5aUo
RLXLECbPcwRzeTBOEYrpizvPEYNWtGhpDzWym4gSS+BGHctPiBDKUVc3EbmL0nZUjQNDRpVfvoHp
RmZsubEZ5hQ9OazcbNeYt4VjfiOjcqoED9oMD0pRtdAzbq2XdeWJuQ1+ARgJ7VmQ5tUnI6iiaZBs
BlzulKKZmu217sKzbyT+xv4rYNR9vick3ZUiS0lQg/LvilwS0vN8PiJNQZUPUqYkV4nec1+NZZ5R
Tw6ZvVGoZCX9YNxVZ1KtdQXt2ACwK1IMuFxSHyKjwSA6IO8YSy+jPrWe5Mc1Wohmo7vD1OVw5jFV
OLjBds37PNPc1xF2J6RvtW5wIF2etOIaKN0QdxuDo2hEPPe/zCLFwtPyKelb7G5a1LCC2yGPX1wZ
BffJ06sDaoGifuZcQIJv1i70CJEbkvNVHFZAIzJKJ8cyqsEpVzU0OJ8o0hJKtI0khZIlXpITaOKj
XoXYyUBiZeKXn3Z6fitbyVod+FEnvhqv4uq6bQct/F0Pt/83lAGCeau8gnWOVDs6CGUzlU2FGrvx
zO6UpgmGFmcHZzYN+Oy+9ZOZgS6ZfensKykKc7XjPsRlwDhkTQkEq07TY0X4ULXsd4A8efsRbvD0
q0JZUf1R2Dubufmg+/110WfYtNNdQfwNLSlV2ssbg0sxtwdsKgLh6HHWFuK/FDp5zQui4AXmDJAT
EYSEWjVMwJevnfShwyxj0/R37TAw+wk5D+Vn7oMLCUOaV9uaeSDKZnDZ6iuIkHxjC/iAwLiz5it6
o8aWUkR47Ju6JxtBjfuN2jmRIm5dtVhlqlx7GTZQoYA67KO2XqfOp8/UMGeo1uGnp9jY+/5LTkzE
nOgxhmvG0pFCwRssTNQG3LumDwP0gKiwbvaPxysFjSSuIAY0Pao/BPsax9rWSiM7QuAIrlimsXOl
3HGGH0mftEl+aWadelV/mMsDSWuwH/0COUU7JjwgKKmCeK7wOYVCfpov38nWGPFpDJKiIG2Iat3G
MaDI+bTfZm9DynRs7cWMmSGVvkW5dCjoz8SpTts/00DDfeEq9OZ4zTPYa8P0esMjqdAcC/ap+5iP
q4Vd2LqDekO0+/JNvv05d8vPD+bmjfjYtRHTGpFEIh22aYM4/2bJAyoNDTc13zo2FHgOYAtCYbTM
KshSMy+m5P1P8g6t/ls6pndXy7jtsA05EDVEz+w6X8KJ5QAzg5eIU22ihBpxkXQ4lk/PDHytiSk+
yx/KPiHiu6PXPR5bUy88G0OOXrfyPAOHuaej/TxFxFpzqr1/InXom9dJhXxz2DJrxpa5WE3j0J0W
/qs45iONeM87EJa/CljV321cfW4JnFRUTAcI7l+NH3oH2bBgWIK5v9RhDld6/LuXs4W7ERuffOhG
gJt2gggQOtTLgoD5BH9+CWG6Xq0/7ZoA8yiHROJSm/jz0WuXmjk94kquOWsjJRryj0Lfx6c/qtqI
7badH0c4lweFMmZM/DU8tiCZMWLiPH8WZC2bXPyLmi4V/cVXE0DU9IuhfTTKqvgOw/QjRvEEUuDm
NoCOimvOZZ9z5c4bsMtK2nCdLFBZYOCQJO1/8HJ+RPzV0zUA+B9CfSlU4hKLLkiLRYXVbAqFPU/Q
F8KJtwTlNOSsET4qPhfN9H6wZ/Hz6DTtXMM5T9X9LHWwMOQfFZ5jynuEN6mSmdr7r6IBYKoNd+DK
fCp7mkQUTJORgkfa4TIPk3FkcQ1oIXkjUSYkS8rImtG/a7hFvFRmjRrq4sl8Ah6W09bjB5bx8WrK
UnVbJmoxhDu3WmWX5g2ZnTXPu0P1MVHRDPhIsysDW/a2mtYa+Ityy+Sophrq2f5CIAxCKngK8KXT
eaOeSvvskSBPi17VtBe2vKaIK47QFhtk3rm8NWXHA9EZcT92zcVYmldFcZZkUUadM/gfhzwLPDD1
OggOjNiYnCw9E1HDpba2TnPUiZn2Mn307yq6pGhrap6kxWcgBZ4nIe96Sxt6ax6CfQ5cOR4VLUed
fRVSs6JDUZVwG08Ce69MMKjw0Viy3MHVHkyvcMUhXgurqLGenHiUhFi9FgImS/WygBZsJAOLRKAT
XJnv+CMK6zldXP8q0oFWx/n32SjlXrJXWhbIWt/D8EhFsSozMBbMxt2CYMZ5B5ZpqEw1KVSvDIZY
drbpdyuh/sD+ZP7nglMRMB6DVClcqCb3DuX4exK/ujpPb23ILCmah1HyNFQXUVTKM7MlP4okxrqa
h7ScVBPHFUlt/uxiHui3TPOlOW6TgBZ3dcE5R820UxZsIZIehlwcfA1R5CfYikur9NS0GVz+4P20
RDYsBxEDDJCe+r63IqnD9XTZ4OWuIh/kjlYE/DsaJSsMHxy9U9YpnLRdVyP8hCfxIH8xZYYDqPE4
DwgGnrdpfO8d7dT8Gqedp0LQCoeGdCJmC5pXt9wQHPRB/i0B6FUtvabRwvkFLCvHOcnVNXBHAfOt
xzWHEcU/kDPyp4AmY2Rlf2IxBHJNFLqxPPBF9ZwWJU1WTY1koaTMma3b21992z49d6JWiXpawtFr
4ODTXVGFCrYi56atn/i+X8c45oAfEqQxpyZVhiTIiB4fAMnA4J7q1je2F2eGk5sn/VrvwY0BPTb1
N/s2MFN1Z1vQd4z3bM/kL5TutgLgH3ZtC67zQ9XOplEmg+HBtD3bGBnhacRXj0CifCtk971ZSKLu
rGYXOGEgKKjvxoP8GDdko18n8yXWQ8neIsjUbXbzIRxx1nwJcOm7IjOKtk14A4Kv6sGVTLz/u9lW
d4Ex0jTOPvfptKdF7sowyVy4do4s7rMz4WwjK1eC8xgnvKJtiLw+XjGXoxaWQasSUbm8GscPrW/K
svU2N4w49uapN12/EONoCk1R96rS13dCGZqvx5SLjZUxWrN364E7Ki5Lni91o0YVwZ925fxdI0aa
XLeJC+ycRxpzqzGvh1tMqVozIDIvGE5h9jFBEDqHOWIKr9s8j/buQfDJf4I7rCgTdK/DgJgoLiJO
ga0NUdhUjZNdYVtTxJnhaiEs3SFHaY1szcRzMLA5faren2H/dzUxCV/dY4jZlHA3rMuePPqtX1TT
bJSOlqaZQzDWOFKxYa6dbaYJtlgPmT0rkTcIiGnX7ZuGZo7IHFq4+XACZxVQq9wMBVO3cPjuCetj
EHd9NZTuFcAa/zKZ482igH6qzQa/stMNFB3O22AMQ4TFN6GUHhV7hsno4qNa3B+XRHvGfToVEDny
N0jRoBIzCwlXuqdH2BA3mQ0VCyrKyzIoY9+XVUBdF8OQDIzWDys1vyfLRUuGhoipljdnuHweV1Wr
vEZO/7teoemgU0sGwuz7hf+XsAM7a6G+5mwoZ+RWBdoUYC8q6CrlDEWmO4sXVJF5B1EEbYAn4z8u
Wlf2KjAFm+f/rOJQt0Rvurh9FrzEy9q33t58C1aZMQmWeuAw2GDKVs/apiAgkhT0t06dl3RXzrsO
/CHepjnD9v7n2Mbu5NK3vya3OvjsMqBT+lWH9BTM9c7XnckEEdxmoMUZjbw6Nwmiqr8I4yFB6fMQ
/UScrMdEfRP56uT3QGj1buPVh1G3U4B+UosxtNhLm2j8UwenHjhnndSRMnNCuNcxjoM0xzrD/S6C
nNvXsas7uLru0dvWevEhmEc8QRzXjLPHEjyF31UNg7jAo4S24fJ+T6TuQkGAZ7lbqJc7GIvDOzeC
ZJ8mrNGiyLGUfOQFwkdf62P8MCkqebnZdpLcvNP81FlleStvk9kwooZrBYYki9vXbVNnV/jTJs9E
A4Kq6sSfOLNC/4aKrhgTXryxFQzcIsCnMqrdDNUNty/6rHNmhhVQEkThypfPFeNfmlAHDavZg7sB
XA2we95H/WcVunbOSqA30EDH0zQOakAIoTF1gG9cA1VUdA5KuWQlFZsdsO7+YXZ1iDyMrmPEB5Ff
W1SOoitC0GGcyORNO0Sl+GkST4AZzFgCoten9+Mw2GbBHt760LKTiK5mNgiK9Fv70KhDLVECYpUR
fdqnRr5+tb9QjOsWYfUcOMgf5zZoUumFKvodHBgCNWUGru0+rt9A4ztdojkg/o6Izfvc/e9unSXI
W85GuBcEgk2II+eaP+4QB2eYZNj736F5jzprGCSYhkmCxHyWErVHVwRSpAYdWqgVwt/IgxygDG4N
80hU6JiXgeCD79sKXpEiCqlxOsrj7YtWhZ0iOKY9dkgv5gzrpGFwfhBfDn5sa0yQhsX5i9uE4YKO
nbYJvLjltKPyZ+9ozgPwgEglhfUgaCrq5pQ6W3HZJHtmOjNaULF/S2FVyQGHMh6AHM5cpbXYxplK
Z1/nDjHbEUZtSjnG/JDajVIk2tCicUW/Cp36tcZlj+OdvMml+x/hpKIEXADZjF4OtifCHzW03hJp
+xW6ol0XlHJu7IancCbSR/I18kj3s7uoJPteyYGY6kPdZVV1V6j3rYu2HdJZ5SHQ81sImLpRIRNC
P4WMDR78vWUt3dQ86glQCXjC1L4FmEsVdl26UTbMkhsE7ezo0jvZtrTi9mOMWmNtiTXnrfxHhyDr
EgXuE6yG3CMljAX518PkHsRFquo6pYjiRP7DF5MKxps1hBHX+ToFpIufjT6LcXXiDJwbJAqoIkeP
QnwvGPnnbIyH4qy21hCkdm/vRLhsFOSnBXHSLvdVY1dwMZXDV+bxXxdPOn6qyVZZCZux6PUuY0zh
BVtiMoYT/k97D9k2FtAta2aZt5yiFSPcPqTn5jTve6Q9CKUN7iySdu84UVAbEaXdvzNGh7aCeEMv
TRNDXYDHThsJ7CuCOHFqGCVv45dGAJiuU9gyaAHovU+CizBVLxsbl7anJBeyRDDq1P/6RiaH0Y/n
h95+GzRnzitPvauwBJ4f8hZh23Sv2D9mHrTBkjFweEyzESX/AHAxzmMq2hUkHTAAky4xblwKPVj4
7V38JJUmaA0q/XTIdGAniyCtqaKEaB3T4YMsJYPO4mVl6g8TbqhL5RiSnEmSi9m21EYIE50e6RDC
TNj5DOZ83zNpFtXF12nsS23b+pyxmxvZXq3gGrs8ZZvIn23K2wXVNErQbcg1IJU8adB99pfrQ5E8
YFCVWQv0f6R6uBagNGRU9zzOlzB3o7yHphKnoI6AjqBdp1p4J3OhTxcYaF7NzacehaF7IeloR8K4
qlgaUyQ4okUpWZuCkkczNCf1QFUW0aqJaHOlAZWOfaNsGhmjEHHMmBMmWKQQRQ3Zskz0LmK9HmaB
jaAM0d0wdUEG4hzm2DO1T3TlPCfFeHBAnUvOaA0u2KAvKkdV01WTMAJVo7XFr2AyN5PH+QhDhNgJ
SMey9n2KNp3llCBJbkYBrRZwv9OdeQTvLpWfhM7Oc5sbRcVmyNuDvxi1rVweTSL1st8lcBGcB6uX
kZ4S2ilxK6hoOduG8GFT9dp94zUPb/ExHKF3Yw2GYlPcBBKdfF0yZ4olfZEcVoObUiJ7Fmek/LoK
gTepulr/VaLHY66tKSWKhBbrjgxtoQvKP53Bsu4lbfzSfFpnMBlGmAi006LDvxlpgbQMioi8nML1
WwOXMOpeYAtI4u2Vjsg1nxlYS1xSrSLbplrCj9XpKXTRezlGh5Ba8beoIb0k6nqCt0zYCE/Vw4Bn
A3qulIYSkRQk7CpR88p5c8Ypu7EQfjxa38DwhNVqLXriMqAhWKxa8YMu3fYnVG6wLTUlEDAdsDXY
SLmDHOKM0LETGmtLVLXMslQyvgPYHG9wtWiNBQnyT2Lfs8SlVhhXq3wEh8ur2e4HFKzpRoMzkePu
LCsfGlC9/l7fm9XP6Mt1cNJeCI54FzspTDkqdS9+Afhet4kPkml+wO28rDe3A15lcus7ZqEmDLN0
M8mgVXeOumkXbFdT4KUhiky2MGOz7qaPe0n7Fh7oEWlaIfLylCWI0cCyQt1do6rbMQVIBrva3p0u
/wkLc9XT/73UWniUpdZ55k5igm7t/CFevFMLhQO2Yxjye1yNOs6CTJV+Rp8AbA3yORzLn2WrBeO+
cQ3Q0Hjt4GB2vSF0hTcP2BdX0RZLAbRZbc2DZ7XB8Pmfj5T+WWifB+mu01WLodvObareiAy499dj
rUSu+wiGPcZ5H4jQDelqXCga8lJsNBPigbxOBHSU7Ye9WsN3yolhHEn7190vlDYNZOvJHa3RYgsh
aK3R6iLaJoUqgM1kZoguIqGYElbKgctlFHO04+7XnRZIAEgnYtQ55OiJp6lRsp3E9HlLmVl6wfMN
4ywbAjcJiby9jQEHfjKdA+9Sx328y7lYHmQnddax3CjxTGICYqFX8CNJgvSXaIRrQE0lWRjA0pJX
XGPr1ZkORUJKRMVzBop92QnDExS0ziIs71PVHwYGsFQ1ky+/w9Iv64mTOz1VeSexUi88hvJCYtra
+gknqKCXD0vs7nO9KZfz95yv4J3nb57qraFVA+lCVAEc8MlnkXsnMSnmt5+1WBxj7epirqKYSn5U
34zqmk6RRN+8vVwxyYjN7yYkyq+zHSxHJSfTyJI/gak7QQaXYJScAT2w2zzxnBgrnDAmEvXSB5EL
3Q8ac7M2rtK7pgrbJBEc4wQB+swePkY5kgNCE+gS4mjy80VKgDounSpo2lcIQGm3eEN0I0ycLNUC
rINzlNWsshg/aZj1IrVy0QigG8iIg1AnW6eQBVSdpVI9m5KNlfBErbEKi+Ubwmu1JSp/61LIkgqN
BINhMDyruG66x4E5DbXlmwy5l5yfM7DEux/2STijRqN46wGUSM+fzRPgbO+uykc3lNxGvRnhFBmA
jOhvagDQCj9916MSD1nXdV/YDd7bP+q2jdT+8sprmaNIopFsHtdGFdMWHhDvHqbOMaeGLjUklFfC
2x8jO2vl2cPyk2fHwm0sl198oR09EbNWdydrIk65bTNHP7hCg2DE04SgY54Mf+fSgGgHZob8PpgQ
DeEKRN/Gwm2aaMd3x+rKNDv08c7I006/Tgs1yA+dsiYwplRG0ReBZq2WSa7UcXJDnavKCPXLz8yu
2ogMD1LOln9Jj1uQIyUR2ycFJgpw01I7z8pF6QzlPm572v5rXWqA6U8PatNAVCXMx1PPm8RM+T1k
e8gZ9nhy1z90MK0I8rvMfbBpulzp2i2ax+avy5bbLhD1N73aa3KUrViSyc2ZFwvXOaUaWf3JnJ7c
7lJWXWjmuMwWPRFD09xnghdnRbbrstd1pf+JxenDGSOWBGsirHeoghl5jU1PeMoQKDSE8kymQUgZ
rd4EAipNaPd4Gh8ZyaZj89EnN3m+9AfCXpG9avnGWIHL02o3wOiWPHxoarCNu006PSts3Vdyzkfa
F+PODxTOVxO+I0vXsf/ob/V0j3dgaLsmwWXqZo0NpN+MptMtNDPlFnsPEr9J0WYAtfM93lVAaNf9
ckQ2QkNBI6ewMcYXN4e9bDbv0eoH9qHX+/MLnXy72JabDPh2w4SWvzXNwmjOHLHDzzTUW9b38fLO
nejW3Wm9J4w+O+R7V9AoBCGs5gZFQQ854otND/dFUg+rB2PDI4nf6fVJo+ZllRLYmf6uYUI6cYeP
lMTgSGYAxzm6HZot+zD3jMlvU5vxvnZiCDjAP95tmvgDGARd3sPjhhiF7yXL1AdPqO4WTzaltQqX
AufXfbQ7FA42FdoMsmUHCH9Rod5+4mmuzPwAaKzCCUlDAXiHwOIoAxmrlqUlabge8RWbi6wPeKzw
apCqDIoEDNtwJ+h8eHcf9PT5sGWQ7aGGksC6pl6blSs0QDtCJ0Nftu5bOuFj/3AzN5VmGHKbIfNJ
ORYql1YnYT5k/X19EtXyZE6lHCz6moL9LU+yfLSgjsPf2AXjf6kh6+qMkxpsYP076r2i74/JzQqD
ow/iuLIb5VP6lc1eBC9mZ3N9VEP3EENZ9b1nYssNT9AIOQMnpVDPBOnauEfU+Wtehx/ZUiP+hAfI
2qYLpXE52ZKX17OTpxZcuYYAEu8U4yrNkXp4YhtsoIssny648zIcWBb34dbGIB0XVx4wDfJ9Rrnd
+4kGt1hjQKB569lM9UoOmBHVqd6KYkyYu+4M/VZmdjcLSipViIMLz6045PbH1JcmjGtIEr2dOg+A
a85k/OO7e8fl0Sc46yh2SKf7uvF8n7/P9ygiWlAUZi1JfahDL6k4BJqYxvYDWDgPLmyzstkp7Z7U
Fup68iyaXTrWVf2+Ykbn43RPmYZCnYMy/wV/eqC/OFVpcV+6YuFGV1DDxO9iLt0GDRLYKe93jHJc
cPJKqFHP6f7h/WaMsD6PH7VkhI3zbeMq13c6jrkGsEcPMN9pTiUzG33Xhbf0YdqIErhrQbYbYviW
WttKSmYqpea+uxZPdc+NqbEmSZ5iqnSwp74NW1HYSssGQAU8VfsCBcOv2PJsxzfsUHa8Uf9SR2ZS
dRAITuJXJ2hQ/wtk+JLXp9TIivgruG2yTtIXelhtZUreNnKKWv8HDNUvlU6U4iOBt9hx5MTkKTln
NiM5Bxx11/7/xK90mP5k1Tubz79QqQWHE5LHvvWc71QVMiRNDD8LsQDNylItS3ILnmlxy6yGM25f
q5eTMAc2xrvvD2Q9V0RAdlS/8QzkrtwUFlOMOzFYaLcPFxy91obCrSsG13x8FiG8aEtsm0j67S2I
4AtVUuQd2dot3uAWv0FM3vxUDRpdU3kit8w5+Mg1LPyMtrm7Ww/lqYNML4c9GQwpAilzN5ss3GBB
PFk6g/kfCkGgTWdzXyLdX6wsDLUrlOmqDNufmI3EhUdG4HaKpOkdJQjk5vBicQ3PfAWPRvVPlzJ5
Ko4Y5DkCCTDaZp0mZiLaTWaJoYsAgqwJEBnIhntlcz5PPjr6QyKMHUGTI63ie59xzif9/ZfaP8dL
aXZdhKt8kBF8KEJaW1Azys6eA/Lk9h6drFolIflQi79FRJvGUUSjU2xwKVYf5+hn63BjmmL8b/Nc
PkhV1C55ZkSJZDSh2WSs2fSRXzCYOGhJ8riH6j03hzRFKVMjQPpPbMjQcvehf8F4/2S0Gd7NCOft
BWYq/k/7ViY+BmXrnaG7CdW/w7PEJvLbUObtt9ZZwvOdKX8gX0EqTCeg6D5zlJAehrq04ANIg8tS
gdgLmPkbbH9l9sHy/G3yKZh+oaN3e7ahsVm3QdxsKa+Ia0twGG7cMskwXbjcwqW2wmDdTRnOv5l5
tdpM2WCltTbyFoKaRpbabbfiTI0HHPwDTlVjdAtxjLVoMBJbPgQQU+0Kv3b//oaRp9UEY/zAjHm4
y5XA93IV3QT6Rc2nRAbGJAJ9ri6cyuLT6HAc3vA+YP8lAmiTLSgJjOtXOekd5PTJOWqhBOemPGSS
NZYmer8E1l0kqvLTxvjn14g/Ig+9a8MO0IxPsXmpqgrHcM8B1CiO0PlcdTQ5cHphdaXGASPT3/P/
VCwI/tf6/g2xhHRHeU3R3NXUSRv/jhN87x06kh6DdiP15cuMv82gnatXBVJ2IlSCJLAU/T4mBeI9
PQkXJ44EL9FyvcNNxsmN8FrGhevAvC43M/coqmTS2pTkpj2cIjZMIvuo4+qeB2qoCBZjfIJxHz93
9h8i0+b3peq6XFJ+l6Apw3lexVILxr3h1UeSEeAKKHbKvg8l5PrupRfYp6RumMznUekikD1G5E8i
+pnHzd79CvvF/pYPHPpD8MXt8tBrAfiULD4hvj/s5t3SJvQ7EluDesx5MbWHunL6IZlNsw47IcEH
PcnA9oUMERuKcswSM6Fqdf0/WdO7A1526IJtC9EAx2lZplbdwUmnGmY3k5SeLvArq5L2YvT6LYWP
CgWGYW/AvF3Lb6JozYk5zPJtYSrESebj6yQbsUEfl9s07SxsiNJDnTwQ/wf6xFUjZXKGdVZqKtuZ
GXU8pGhTEMqx56r7RKK6WLY2rnGQR7FYz3rFRpJk86xTjd6eJ6PN9XDVkhKgXNnFZ6KOP93uIIdJ
9VFVk0i9JdTATghpvO/MiiXmYdVfSF2PPBlbitRJw6ZzXbltvxs4H/HSFo2zX6Cl4nmTTCR8ZaLz
cS0cpJDPB11xZaSca3d06p4/ba9YTpURF5nF9FXtdev7m2SldHu/MaaCifK8qJiJ57dvGdPdxNgc
ETLfrlY0VmJgogCuxX2kXEqPaZhRL1rQhbjXYuV9ki/x3f4cDBi6zUNbttE7P6zSU3gDis0P3kwr
TpxiobS/i7QM51M/yZFLCpbeFprS4I/hLMFzch+bHq2ZeaXA2R1hZpp9C9ac5nAoQcfnkd5iOEKW
yFQH+yMCpKac/W+W7alpIYcKC6hMHEUMp9PmATXb/jZzhE/dD8oJKklFC+W8uwjy3cz4AXoW4JDR
//nETve3c+o+hEn/t4RGKpDBrI7qCfLpiAJkhqqHsW1eIwnbnyroBx/cUIAfp5nbDs8dGP3goCcH
nEexyTSSunRB+TLt+O8bHs/j78fXzgyXysbVPWd8UAme1EVhSCfBKZ5QaZ9+pUvsp+qy5APwIHPH
bdcEwgjEmHGoQ0+sxEoLXwP5XuJHNqFRJjz7XM3iujQofJJSd3iXnWXg0OT7d+p/82koKmb9oI/i
8bvPf8sqCR01SXE4/+nxgi4cM+2not38/W4f2kUS5Vn2WGluZPMOa6qGYllyi4p1VhewBILApZK1
pdjHdoX7uFl43lPCn+6KtLOpsA4iipswNDqe/hBajzDqfrLsb4G7gTZUidwwWLR/zzUaxt3xIl7t
wA7rlnuRfUpBTV/g8sED2Zuu1xDzUaA9Q0r1g1Om/i2feBUHJ0C0hcaf8BcMD4SIJJmCAmRqVZ7l
r5OGEnpgqI9pqHJybhauDerR8FRatKE+uqBLYG132IakGIKXNLcidjWK7WgckR43Gv9PjXa/wVOr
to2Pd7KKpwGy5r6hJrOeY+6zGfyCPjglkSjN6XHY5pTdmenM9pZaz8dpAPW1y0DagsiY3LVE+/Gl
34/tA8hAQHlrg8zdLv17GobhJvp0UnLW0Ejn3z2RM3E3tEhOh9YfOQzxa9g+5YdulI9ocBAC1H2T
z7aHBn0HFObaZKD81ZnZrFfsBGMD6zLNBZlAO1V8S9hoJ427y4AlJPIxTwhVk6Qk39v2NohPxY4s
C2uVeXMUtNKwhiK9tgxGoa2bSIg2EAf3Tet0S9lwzlKWfEGUBuwgdijvXjNBowW8RzWL3eWwjvO3
rLQ8/lrGYrN+UR+Nm+hD+jbK5s++8JjN73Y5uNCQ9MAtTWz/cRycZH1UVSOHqWR79V2PeweXjYp3
9sejHbYA3eaTy3eHdFyzWEA0EpauD1nYcaCxVo1HGj4ZPI3ZPJ5xucTTTdx2yno/465Ye9NaR+LS
I4oAiIXr7/4xwVUj43qGzdziamnso+3q1iiN+R43h44emKm0FFio5Zw2pi+Z8GkZ56ITyKhDuvT1
599RNCN8MzDWMnGyYsS66LtMASA5LwE6BEWekwHxcMRK7DGZ9ZKlkdNzCLaE2t6qAjB3l9vELCT8
qpUXZeRXQbyUoosKWudMuAFVXOE6+rK8JcxeEmtCR3FL4oK/Bxcti1lEhtfyi5UW/gcci8Pz7yEQ
bLrC5GIWAqzslh27vxS3GwvtFiBa3zAcDXa2wt6vo+8sll2FiFe75ffY/hqm3pOf3mvQH50gKBeQ
TXrP1LCgpD6Yal2LzMBZ+CUz1b+I8fOnz9Kld5vsc/oHkKemMFTocypwvrf+uzQ7FNFlwwH9845s
1cMhLnrCiDsg3InWGIKq7V4FrfIXOp+l7xAMZCf5jDHoJLQy1rWz/w4jb4QcaC3FfVgfYtwy4PDi
sWvN7k6shj8yqNo85yaCGzuSU7NnErUE3WMndOHksAnjCzOqyk5ktD3Bc4lI9qpS/xDcWO3Vmtzy
iwCNJYyAfT2JQ6/Pnwpqa+oHvTFxZwM0wOChp754mBWzOyB3NGQUB+xAkcIVH+FDYp/Uo60FLrBe
D1+cNM9U5RefrxYvGdE5YeVSP8KJrnLmhINQ1OoUlcAteJ2O32MQqDpqYookHO5unjU3PmWcsBla
509S+PpRhRmLqib57X3P8y15A2+xqtJNertFvZOg2GcAVA49w9jdrxUM5X9bKepyYKX7oyaf9V9C
MS2tCSD0EeXGKl5De8ixENBH53qsfhD/JR5Ar23n/7FipCQV4LlaQiG18AavRLQXfHIejLxdE0/S
eEzEK67/+B788u+xdxBJsQXtQrPCnrV1aK5jdH/JM8O71XfOiSwa+aqv2kqXJiPCpiPTfd4UdR3c
7AA0U0q8V+QAXu6ijdxKHDNWXgOOwpNLUaMtzJRshUomWNyPci+YK/DvlW9w6S8uy06OlXj5ZCWv
A4Fs7j+cYV6hX3ZGxDu7mATlUjyWBp8tPy17EOnGKsSzWJN45RWiNVt6yb/GcmMCcY2V42SYReNz
yDJpL7KEUm2VAMi5V2IE+eQxHzIFNuusYfzIAV6CeiYwoEXVj0Bncl/T6lXLvOKGx/JVYtC5yRnr
EQKh/y3M60InQi6hYWOTQpYOyiGQs9Y36siSoeaUXJgO3Qh8rQR5J8y1Xyiq1AyUFqfkGTPLHtGl
oFpOyXix+GgbuoDUaPupyGtk/YwR6j2qmFFS7dxfEWDEHBJbD4BEraynAYRpn8kdbGn4CeXFdVL8
u1/aqByjzEZQUMEWSX+8I65vO2kGluTao/Rqk/7fK6BnZlevvE5uKoiO4TRLV2X6D28X64ZrrBU+
56EqpwrnMfzmLaH2Z6USLVsjKy1MYeFgy7fRQNUbSyZJMYYqz8PgNrBs82uWoRXFFJ3fC+jBpp8H
f9WFbSxuM76NhWFqF60axJYtr9ziEZg7XJMyXPSj2uqEXQfeskVMEYs0StcVhAtDPHKx3Ovufala
z2QMBHUXACqj0Mm+dGz+f6K4Q8WOoHQzCDzQxT01oUbnYd9JTED9OcyuErb06ZNtJzM2F67p1LUJ
YS2EFqkN7uc67Vi31M3ONmX8SqSm4E61LBHD8s8Et/Gt3xVr3KTp64qd77JxMMXGXOO5UA97tHwk
AS3eucv3MmhZZCfWapSMUtApg9/K1uKujmqlEMEtZmQzn3559Wxy4sYI+OfH61iprcq6ogXTZqmM
0GYY4xnkKTQy8Hnpn0W6uqY/MFx4/FzJnW82HVp1El/vdWcqT/TbBKbl/NMB21WIf2d0ZEYGOxsk
p5z93pCIPS6EO2mrmanPbkaQKOWbXfrf5vjckrtjVEjRJ+lFMVZveL9MhrCkRzCAUSBHfb9gh5pI
o/lGdKUulzWQ+uHy51zGOznQElMVuC42QnKY/aVRLz6QtwV73wwpLSnyeqG8HYqHHryJOsbL1/lt
G0LH6tgkdvWjBTWDSKsZQgrP0t2ZUcXQlhHGWUz2zXDQsfoB2VtWvDMcapvGXn7uIWO39aJT+1uB
o5HZZlIl0kEV6wIMqaYy2UOGsCwn2UDUyR+C26DoWxNluP3J/uU7JPvngjUyHM4Jg2U4k9JSZKwi
y9Kle0YFj0s4EwSdfZVmwkXkYDhMgeNpjSmL1i1nb8RNfiSuN6y1raXsQGFKhP9fYg4aLXCfCmdP
AdoKBjzzKTDrYuILhvLfMssk3WLUYFEz5I9o2qawkNMQEJdZtYNdyukiPvwR7nfNtGS6fKotcgIP
rcEQ1sLQKYHGC4MxSyAzESi4P3UbBnQY+tSEruxgimwioETHIPRF1U0SYSsUFuHUULdWFguIJYYk
Nql1+gyCtBu/HWiWMJPQcoprJ5LTf3dLy84/lYZiEmlVuGzOIPkfphHjhUbfucCiii+TXBxq0LM3
x7u/Gy+H8dCGJtdBZjAyYn398kHOgaxojRQKnKhJdPDDlD5Yi8GowEO+P10wRCawgk/XIKUFoVtB
EhZaHSBBvh8VVqPcbUgF9b5UX2P8rc+YvHJBYG79tFtOz2owmEScB35of+fjB1KnjbFfuNmT6X3Z
cRY20sPsAp2DCzBAvxMADer3kv6GqpNozVjbxF79EFuLG0spb0SvoBp0HITbA+NDe/GUV+dtRcSq
8KM4dwKQFlI/Aq9RnEkXC0wFEc3RskGTo2HmPUJ/3GG7HYNCbd2bpXvPoSnY2QRf6JluWwAIuyQn
Y3YimmG1cc+zHJ0D9hkdP/aIp8XG6+BESp9ZBZCF79zrIkdlLnZqJeozagOnFaqYn+RRSg2JhfHA
1ty+XgZwZjEXI2JNkQtgq0JjEjXqhKl/doMb9UdQ4WZkSrJQ0gNo4haIiucZk6rr4Kf2ZS72cCqD
K3+0KMVgEY6SADK+vvkzzzrv04KiaLAH+tyWJXmRCMK+Q9m/5tO8MPQDLFz39iYLvVzp6+wdVRlV
QqNY3pwFRYeXANsmzuT7nsmps9PkDclpyFy1yfl61+ExgZRVTJT37mg+7D4xwU2xIkxg7dGISseT
vdDNDdNl5cY22de4JqRW23gojBSS7Ls0X3A1B6uJCe2bCOhPeW2IXxvq2vLI40rwiOdCgSOCi26i
Xgyt6TF04CAQXiibIGcxZ2fHDjD/xQvR0KaVHFFeQjX2MJ+KAS6rTdZSvvdXipmYJJyyiEM5puKs
ZCFU7ub+NXQ+SlRDETNnuy3L51zNfgtgg5M4ah/svcIPZqBYIkIWS76NKedXUTc8DTanQsqtpTqq
OhHviYAIe+j/S63jjHpQXCpUPEu32wMTC+qHajBLNHQne/WZCcNNDrgK7epAN3R/rpDgXg2/9M6L
7AsRRYzeYN0VTeRqrwt2OvMNVrrvNf3y2JZWeEVkzPfJQc9qcZgpyTKZ4Yqb7QjMbBrzJjEAR0pL
LL2l5+T9GmZyRkWbGbDPwPR4LhoanoJ4eEHZa4eOXVWRs8mfCl6LcpmNvq3stm7sZbPpUZexum8Q
4ox0KXwRrU92SJ5MRsEKtUkx8z8F2t1M6UrqGs32MZpMfAfDlSg16HvfhadZw6IqVw+LIaXsOuny
9ipact0hKSxTipgFPmwGHqPiTQx+LBSneyDDUjyjbAwDwfHUMGa6NSZH1sMNLBtqpN8mFssImG9Y
cF0P+Tipa013TIJPyHX3OQ3oxIyZeLw1yNVjq86cjBylSZHnFJ9EjiFpGANRumj9Hr0rkPUYyEXT
N1RN0hzs53HtVaf820zkkRfLKo6kYXj86G+U5Wb8w/9SXT/CNmHGm7p423SZYqnIPghhK5qhm/kl
BHO853oRLsNtpgCoIZrBny6Td5AHN9aDTUvFv1mcub6YrwpiPC4B12QGgiYHUNFC+D4roVs4m52I
W9d0g59QEsaZxlsbRC9ZjAGIJN3Hs9ybO0VVvxi2a5MEiWRQUYLD2xH0YoaCv4QUXhd4gz4sSR9m
mQKDhRf8iUZF24JYxaeRetYteN+Nt6U9M+vA7McdpV1pT2NJ0Mc2WVOOLf1FnQZE99Zz8UMdp8ch
+uf/tf1SxKBvdO71QAXhlRdwJnLzslHLook55muoQrPuu1VqRTeG85X1OgBEtew70MUd2fWT60gz
z8YAH6WsMEID1KQ00rUIwoSBKvOrb9wAXAsxwQLj6KKx7Gk/qyL0oAYvhUCyWETridakVjq/0Zaf
wt/2izJ2QECRxTsH8mcbbRFqc/WS0W+Mpd3mCjov9W8ytbrNV9jgH93cK4BPLkexQdQsKrzCt5xP
i0V55T6NL5ZgeN+RSf5cn4cV1/9+m1t54XXZsPc4a9zQzuntbbGraFjvnLLiUM3m9BpaPRRqPxtB
5S79kHf+ED8uQ3tQcK6e2IRNQAR0gFn5N2Ipg+b2ExQ1XXNVovjh1NSAIM3MF8cEUxslAVm+uop9
SFBVAo2/T0JuZ9ghGdnw8KR95XTEGk0oTMbpGcHHhun/+4x66PmBQyfrOPBUyRnnBnHzdx2LxVxY
g2hqpk9zGrYj0nBgJdpSHB0HaH7oUE4kWYhA79n+CiBQT3JzdSY156InL1rYh6TkTDi+SZ8E7A74
aRngwLEyv5pt8bkKcUTGibeon67kwlYdgTpNDccvlj/66P6oxzznLkKzsGxEhU3sOmb1ATD0oyoT
6JuuUgLe97IM6MBmPs5Z3dc2C5x3jUK3kBhY9q4iT3mqfqIVSrFDZ+kEaXyWA3TyQlodDCLOLlRF
KOUtEqsfVVTgX6LpDrxOxRRssswvn1qJlM8CEfdgBKG3mtVAguwy0OcM5phjWwkm9aqogs+rtUM+
IjSLGHFox3UbXF+MfX6m5BBkBI/b65Fckch8xObkRiY8hB+Sdfd/xAkRWOvcbMvcWWNDdY5j+kFH
ZlULPRo1CqwnINAz29HavaKi/OzdIo5K4MuFha6ZxBQNR2+JuV3Gn/8yPDuWtW3DxMSUj08MVjPc
Wr3w/MS/+J+9LPkgBtgO2t5GWCMhZk7QdF/wM/hH+78zK2Cy5KwCS3aZp+jWKjrocIqkE4GVdZ0M
n6NPsBfWpzR6MKYx2r0HcEDCfDZ/Gx7SfUlDzj6+2RT4gJ+zxzkZcjO+IVOoTd70//8XLlXMUSqd
WA8ebTcTYyS+JOJ4O4zscuMizBi88Xm5Tt7H+CI1J6MRo+H3nNOAD/fUOkyWqEql0dhoK6qJx+CZ
ssi5UUPAZls94jUrNvvTBi5YwUeVlVbxC8bcAz3gIYwKj9QXU9fNPM/xWCEnUGyFdRaW5RJcIGTi
YJA/ULJcOrn8KxrpThNO0tDgd3te3LYhZghb3bQCE4i9gVVAIZVboUdq/YejNplgyI41vFepN8Iu
12Q436ryfiWCRc3wnagY7GmtYvGcnzkC4aK3DE7X6SOMwCt0NpTshVSPiqQ1yRJX+wzPldoOhFWY
daa/gFv6zrDJRefv17FxRmhgumlXqjfX/2CZ9FGABdDfFymhAOIJUR5dsfjvSQ/VwCAWcYk16yDu
/gP64LkilHTQcRKPg/SpVzRq/S8prO3yy8VvaxrSZq31jg/fMqiGGT6JDY5R/i0D9DEGGAk6CrLQ
KZOyYiBww35IdFMrIzMH/XWBfWdSiyyZoqPbncGDjYaK+5zfD7Aey0n08G3f1RliK/NNYzV5gV4t
lcwMWpdxBobr2k0h7aJXNX7TMopAVIJDtaBhkTJj5J6z48nVR0KHJz1UAvc9dhSa2mHpw1fhRFV8
wHmYDZlYTrua3KtKJ1qX0PMtAI3c1pLsY7PNDxQaevinwg7FQPkRWASzxnEaQZKDmgLAehj5GtEN
+j1AZAWy6KU+orDBjx7VazecIDdTO63Is0N9zWLAXmhPVvwKr+deWTUDpPTVpgw3D1LxI0LJaHz1
dQYVviv9QPGEAqnyAuzEhVqxmI4YulBqv7Ly5aY+cYBFi2BqYCqynprk4t1+yVOmSxO4dXX68AXL
71FBcFCZ053E65Mr2JYbNBYJh4tcGKtwfkConKUgZ7oUR3IZ6JfOie8jOW07Hd39mj1uR7he62FF
VowE1pGUAdL0B0sf6uGhznsdraD5zfdcW7mPhnZaysDwjp+pHpTTAk0rZoc76CUESMWS98K7oE79
d5wuLb7RW8o4gyC0gMTYiIlR+kgUGasXffBd6siQKdebiwF3EZA6kG0zoj0OVT0uYBXVIPjnXx97
gWoPJ0/PN9dFCZOD86STWvcxf6ebQHTNLcQLC0ZJGxJl7c0mDPhcr5Pd5W567763Ca808DrEv/Mx
ZB7KTXFsTJkZ44m15LM/MNO4/6/3Aw9FCTL3PBAYPnKgaMiyK+HZRsCrMdnUDjSdSLe7Ir9vjfX3
XqAGUpyWTcNXLQRt7bTu4WPrNE3QLh9eo5lsVxpaavVOdIHgnq745oWA5Mr6ly8bFhNaBqkkdFeU
+xO1oOf1L5zx5wkNm3V5xWoBvrhvi33j3unClVrotV3rT96JSwLrGyODdPWcL9z8ZJcOC/cKgNuC
InsVbCHBTUqXjLydiuAM+L4kp9hcETEqqDaYT2ZvMZu1+JHM4BYd5ffc/X7vokjXA52IVTvHxqVj
3lEjUR0EIQWpk1IBXuOAK+s7/0f81boA7hzGRk4YcslEoLTasSjNpjfCHaUW8eBUhot461B96icm
7a49AIWq1oTUrhXn/AMldzqx+LZdvPE11KKrVX4AIWhoL2a0XWdHTFAWMMmz4jJeAoefJzAU5e1B
dEI6HnYzB7NlwP0wDGivfsRa1Bwpl9opuLrA1zVDzKEGDe9+4gedY9ntazPKWYa9i7lZfOLD3lBf
/3S+OxI4qLmQIIqLHX596jachZ2Ph3nI0wKf2nruisTloBzszMSnYPgmlgH4sus2Z2DqvObkUeC5
Wdgv1YAN7f1BrwKwM/diHxIjyGAUAHJSZV0DmCIDtonIDI6D2ufwRg4XCrpnFsKyURYr5hTkvfcP
DaLVDLidGix91WGeUfoLDgWOP3pwnyfEqf5YADu48ccaTYkC5MCLCvOmfObWI2/AuIE84jvS1Nuc
KNat6POm/ZmmMwwBWo28Y/eO/WxZpbGTgyFVfJr4FxXR0dgTIS6hq65gw8reqcC+tZQwOEJ1ODnL
fWQu34Wyj/SFC0/DI4DsbUNGl0hvJM97Z1Ux/2KlzbJL3+gW3q3DVLA0Q0SqmZWQ4hq/TqWDZ1GL
EAyiLiTqyKLJOnv93cD9aknNTOlA69onekyKDs4H6s0Wr4IIQKuiRBuz9deRGwopMSOHBRpDmVsv
sH5zUCIMHBkbjp5ASeMSWcSAWA4YMOnJYRWdRytvNC9btTOSRZNf2YOLzORmP5N/GbATW4KrA+Gm
ZFXR311DTEEWvSd1IhU7Dz+ggD0IueTTU/ZEmPknjEJihEkW7mAE/12YlFB1IfNnYdoW8gIfK9h+
hSovQ65Wk6le35Y12wY15C4RJ2NToDcgYQgn+QPA0KxlzliwKOCCQNlFRTQlBn2MM6c2hCYO4qKK
qVWw4Ce1ssB3Rl4YGUwdI6VOoK7OykjLjf/UnATZdbXB7UPZOGVADkOQMfeS1RVPCyHNadNqeuNj
lPxKA69y65p+SAjpMm9FzKYGCbToPTR2hgOTqqeack5ygx4Q9TPZGrF51VxM//dZAU4ru9AxO267
rj/e+xP44FNPWIUKBnle53mJkOpUvIhL3OmAsAaJgU6nRbu/bE2KS84hUx4pJPKa13WmW5gtCPbN
DCEwuudDPG7p4IOvADOhIVwgLedsSg1CoOnHfFY53DNI57zw/Fc3oSft1eAuz32jM4xLFvCKHusy
y832lEs7h3XFhBSajY7+UHZg5zlHRLx0pi6eo6WIKnDkHUBonPCo/WuHAa8r2eO1mV5CnxQG/rMf
uwsTX0Q9FFOC7DCA05AvKv70L1PKwcEEbR3pkxtOWp++YkYXAujIEwEJ23xcEA18BxFD7J4JTO+r
XjfL5SyAPX7dvhdS873A/4fNrkKtCSneCI0edT3fuawuZCAY8ESDi7WmutfVYLtINX5iX4UvMjzl
WAH6JljsRiVMTl9oUGfvtP8TIxLsIlaeLb2oAgmvkqFwByVw4agZHe1Yw8nbmR3OucUn4GbosDkQ
8adD7cQxHzNLGOcSbRu8IUvgDeh0cMNsRjzdKB3LIg+i51Ffl6xH/kpm45r6muO/wKcZymBbahiZ
bO58uWI8t4gzfCQL9IyZbWXhDnx8MiebZNdKiSj4vKxIzpjQZhZMYXVZvgXB+47SEusSiJZSK1NT
N9lOttysSqM4sLxKjrIZ67xbRcYM0EQz7WjP/mQbNoB4EKCGSW9zEyFivtPhr7aBk/W/c3b9jh/5
k3hsFgPCQ3SWjWyxSeBGk3H7DGsranmOOKlJA8Z3WQgZ489Q21D6ax1644OP+/BWd48jXPkJeB8W
zmIBkOuJFEiCTKIbEMKWjK8y1QrVDuhKCqKz6InuEYiE20GOgRO/16epAfsFmE4Pd2NYrr004ome
HpipKj6BYIDJzhK78a5pb4snZaTUKzUnhdcC2+pQXb6bTIgAXtDfY8ytiPuDRLLPkUWSew5tmK8T
IbMjojCkCQpaJJR9Bgxc2zs1zHGx+PXeWXrp44ldAhNnTDOaj4cRD9m5I3AWvYAPQNv5FW+Rf7m6
0xZsOXpe/ihlArHAhO/VO3Oi8WK12mbomjdkC/atJxCjtbLSjdN2dhbta3irs+1KFCmQP24aFhAf
piFbI0BqIKmc9iP+HCIWReDKsrtkjqH2mZf0ljmUC5RW/ozSMo2iWnz8SNDz30cDifWD8HL9C04o
crzF8NClJKYoZmRmQhucb3EmShM/4MaiptXBCiCHh8lJ0maCPzm+ywnLCcfeAlSmr8Luuq6VAEJX
JRVNAsX32OmOUAbsb7g+rFnLIKQ9SvChnJ4cQGB/ls+AaRg9bIIjGVz66HYOEUmV9qOablRCLjoL
sweYWdvA5QAvo7J41MEyScWi/lRSuWOag7UPJLuRYlZxKfdxJhM+zk+PC1vnrqGy2cN3CyS0E7PZ
iiFzizuSnSrb1VvZGa+wjv465lDismg0ZJMpQSHpFhdXmZ+j+SQpVdhczqpf+63OJBev83uwpsbH
hnajraqcGgpB3SQnQ4pclimMrqjiB1Z0qZWfJ8MaTFd2EG2ouqpxaXAq/jVVKb8ghg5KkcN+zu3U
Wu1v4mzyQYU6YaRnAWkOvyZ4h1QwqFIGoCvFOKPZkEEcG/mMrqhcR8IwwPgWi/SmMTWpFnXBqgiO
UW/H1PB2/D8cTnNjvWIkvnM8g51dsTO3iK86CEGn29cELRxK4Uj1rY3nwH//1QI7R/ZwuQ2xyv8l
qJPLdxebVNYCbgSsP4GzsPmN7CjOtgOAFUOQCdRtjvzvcUPUbXTAeJiBJ3CchKGFXt7YfIZPas4X
dRKxxuA8vi40orETpB3snBsQvdoBgcwqz5LxOj5lUe7tqoXITGNAKapFacfu++z8GcwYQHFUunmI
qODk7JN0G6x27j9vtkaEfAVLBhVYO45v1BHdoHPVLsVzISuZQif0vXEOZKQRKGo/blLD2Gpr+IXO
ibzaQOz8FJ5mWiDn4M8FvvwtJnP5uBcQ/N+DidxaMqpFY5x7kb+zc9SES8K0VuGFk75zK1YiH5y6
VQha2Vx2SAp6Q846HhrpPiO/kKYLrigVVCmX7c+utP6I8UjriOWu1Lns/ZPKCKb9dnpPLcSH1lxY
ITMV7Y2y7zPuG3sq1ICIh3CfVDeHJcUt0DdwYejCE6p7ZGjoa1/PDBWgpCzuebzIjP/dzUoHcV9Z
4gz9gDlAPKOq15lqAvCEVTgnuCFgdc/aZqz1Hos0ocf21aCGEHT9eCUmf3/6vCG9/2f8TSNlDPOS
kREnanAM8hTT9NWniBrCqxIVfsyL8qDFfLQXlY3ZVbiJn3/9OvxXsrodaPvfQJvLqMiBvrtxEMBh
+vs6M1vXihvzNkI7fO9oPYuPnJmx+063/QKoFGWMsWvSgOl5o6HsYMltB7hE65mcx0hZlRklsQeh
ReqMZHzG2myiDkSaUpF4JaZjd+l9gS5OxNpggC9UyNMX1LLpLPtsycZyJjnpkBpsziTN7sHZOAYk
Xh1ObBVjTgF24lAvZjRqR11/frrBZxZhAckIt3DWQM72YmIsNATc7TpoFaDG04CsQGwBtRJ0HgSn
dZU5Zpj7Yol/313lm2d3EVSUz10KBlAPDOXMoZL0qn9vrEGeefQ+Nv4GRSu8Y09N1Qzvxns3mTcW
zBciLAbYrJziMLwikI5IPnbXXO9q2iRrsi9LLv/DybtV/xpPuH7SqZom7FtJJ+FyMCVzjjtaGyON
K6Kj6n+uX5L77ZVjY4opH80Q86Iem/73M8cwl/rU73NURbwXKzkJU8CuWT//SPsBIlkKsS8P8j/Y
ItF+XCX44iG2+T3w8zU21NjmyJIn4K0pVJTVU4PdqZof1fIyrDhpvvXyug4FxPg5kYfkh34Zv5ir
zdSksNRtEkeT1QsgI5SZ/KKrRuudgQ+ZBGgXzP+ghJTRhBjeiblcfwYPwKGJPAM2ad8QlDu/k0FM
RHFtyfluXAoqFHz+uT7YAxe8Hx/zrfWg6y9NAy0oY1PfAS/B79RyAY4AAWPKOe1TzDghIPSMQH6Z
KJIrdXUUp462BdQ0+fbqZ4ecuvF5Pty5NYafq+yjxk+jCKpbG10uupGlbZq+3lyfcXeGdNhyX2Sr
DLHMXICS+Nx0AwjluqJ4n8A9/z9leClNSS/q11nOHtwV1dtSNrYx+gF2EjzWipk6ezNNmd4bHQLE
sU7mXwRuqM2d7tCml9a7i1J9pPqOzMiAAyuvlUBrkm77XMyAAqrl7zeUu8QdErMO7wsXZgFzdova
a6ZA8lCymvnJtNnoYiHz8RAlQ5IEJNhXoLpa5O4l34la9QllKNRVC/j1he6Etk3g4ubB5OQXaO3K
2OF2TqgTkzHjEStIXs469qi/Jbakip/ECIYS9+trTCSfZ9gSmXAVirNqDQCszmELk9/xTA0q61Q0
6KwXkCyFil3KF6iY2x7hw80lkSJWATyK4XuQgQdqpUyelXIbUwcs1kvpWEcTUwJyYqpqnWEoH6o4
7WbYz4I5I9JLNw9JmampGrRcMit7aW7aQ2wiq2M1QIgBddE2NYCUWUYo9irN37KQcSOrmBl4mD+R
D60s5+HhwnL7YV8ZskE7fHrvZ8tLBF+XCy0Mxk4ZH29v1vhzab8jvxUeYuuw6hNH5NscUR4WnGbe
QKZcc18bnv2Cp2wCfqwFWlxb70TWbGykS9X+496xRSwY/4t3224ud1SjxNMoyB5d9iA/ySP+UXuO
ZfemwDgz0Wy7nO4mQnTOAOjlwVerbQ4pHemUjSkcfjBEAbEA0r5NkqiVIwAOX8lYIs+rqUWn/KMq
ZVhg3KXNDSiE8UI5jYW0a4BASh+YBnX81IHZrDusVDUTiPrx1yDsScwnMEnN+UPlf55ZkSv+U5Bw
W54DSZh1BW+uB4J3Py9/UtNbQfWsU6Bi8+ctqRDfsh804nJBeJ1p8borudCoL6IFtDJstBDEcj9Y
p0kio5rRLrPqsIsqgV8HWcL9+UQWxXR4u9O74++BAh4iW21JufCEJHxn3cS/4CzBE48y6cS6EqSW
ng0tWRY1N7Nxwxw5Ylda88cpCbUUHo00TqbDsG9RZ2taMC0eCW0a6kx5h+EcrF9KQTDgA+Zj7SfO
/niCzjdRYg8SrKkc0awZhzNk5qaSXHdmMWjivr6Lh+NSqBVeJuaZWdvg8Yud+TzFI3uOzWR066DD
ekDO2H6adcGTErpdxiTY6zr450iRvOc7Y5ArO2lPq/uVlVI3SAUuxC1sv/tdqNYZBz3/Jgd5DmQg
AkSjIzzkTfzr84vUuC6Lp/DxAQ+HxzHIbz4Q7/Dv0rZsG6hbuYbXszPkWygXLfLpiKPJw91MUHyc
mQkZHQjJheKqEZcsZHd03B/6YuZm1BR+tMIBNWWmzvExvbw+JJNBe6Vvm3x+Vu78X2kIEdqa6ai0
b0UWxDGjULTjkR2wjrTDKtI6KKX+AI2uyVNWCSylJoMC4wCu4zXKkLcm6YZ4fdZZZNKjAloHwGiw
9vjc4tGazCeLW3Yc4STNcUEEXmq9rI/qd+ACsGxM1Y0uPsryELC750F29mkVKJQKlQyimxalSdAL
U1eeHUDDU5qy4w8itnWUZfLgTxKWwWgDRZjt7ZHvoC+0sdvw+vfHxrNixCter4wjhCrXguKeUGRT
ggR1qHAe0Rpfcfxbu+m1MjvRwQ946EDW9oPSfKezc29f6dkNwXl9h2Yr9kDNkTx8TjPGwoPhjsHJ
qjFl9mTmsDj5bmvl/AEpxZqwMsHw1AR2GQAbuCUaHtRTVr0Qmur53Wx5EA0JWZDluxpwCNjNjuId
y5Q1jIKn5RZcxGYi09XpEoN13foYtv2ctdnExLGVID0V11ixT0dKUO+WxCvJBusIoOymaciLnKBt
Kjy7ZrdnYEa5uFwlzTaYh2GbMaucI8Fu7j1LJR3rzdE6q6GE/hk+I2K8/d+n1Avd1fBLK9+G1zV6
4vw0vD5F8lo6xbTksPfLjNYiB2pO29t73EBNUrT0usJsqfw67o6fHGcA5Mgg8P+nDdeeG1Uo3BoW
Xvw52lwh4P4a04xxdikDbIGugBnB5hIqFrNU6JwreC7wYU2KKjwVY5yNT555F17Uxpg+ZL28MEEy
/0QESVdspL6g9ood4JlvQQEN05PjtIKizojtoS/hk7kigxnLDULMjXDVOrKWOUOiL6OYy5vzYW86
iVMNogEVvaHMZyC6u1MZf2mzgjXLbQfYbHcFvQtOKKk22z4cna5leu7w0ux7/2RZyEMeMpKQenLw
KrPvtCBahHBiUG6BWRynLMGRDRNby4LHdMn5yfGqvdozYyXZHXDnoCKGcmjEvapqWp6htMjVSH4M
FurILI0HfNAi3L26Yxxhc1eE+luHDznZnJAmuu17kytYbvcGncgvv/ytTi/X0BsA2+FrMwj1HuZ/
GPxioZw/crGpQT0MGKNn9gO8zFNAItaOn6w7bcdbfciL62TpqWkBP1dBuzEBtGFcA/fURxVKWsq8
E+sT7Xi8sD+Dzwcul1QdjauiVftQaKa2GJW9RZpAxfuN5YqDOp/z/wMdwXXAzYEwd+xkApT9D+cE
oYxSunYviSNTwKI4aBsn2uk7scTwOVjXcMt7k30lUgZ6e/IX8gl59OsDC2FW3BSdhebVAgM5eNVF
E2AEHJeLf2ZD5Ppo7dRSDB0WGkycY032I4wBKWOe3UmBBwrcuMkGJR4gRau/OsJPTbyeFNe1xByI
a+y9OSFUFxr4LV1kVtSNoXpKKVegEBQ/uC9Rg/VRCYsbM1JiNit/UsjXe9y3wDREeajVaBxnU00H
GZeUPeGXN1+IYm587Nsv1NCaJNitlRN3oRTHfdoYvECyiPgnWhDASFU3JtjBA1rSvMtJZnkfMkD6
FDSwPHqmsGYxhrDy/3PJTUrVcc0WR5p21VmDps6lonlkeJv4rttc23FObFXnnPE4GEvSdk/u9YTI
FD+JWFuJE5JYEGw0YObfxKMbQhmPzb9Q4asZW+ViRj+cLb8q2mqyp8VUg8QutzFSuqGWkMqVCLN3
k1QQQrA4/hAoMs1XuRODLZvfGnoJMAsZmgNdbI3dWCbl5714cfavSdlvvpGroO0Bs6hYYuJeaxxQ
FNZHPFKx801frVABy7HVZzikPctCgTTODoz9U6ydReADU1TOqZZiLnaGbqWBhCXeuWHzeJlCWaMa
Bov0VxmEgXSwPz8j6TgIF1ncaGfLpB0jD9GEWQG9Q2ZI9rysNbf325njV+R+5QfmLvnW08Zp58Jg
lsvGImTUeZ92+oupNKkHoHTxAPrz2Ma1zwkz+aBg+I006LCntipAF7WQ/hHtBHW0eCb/+o1RH5JX
MJIR5VHBjI0yteSFOwVLueW1Z1Ns4hDjZ+khGut6SAkps/w5DZjT17u0JtMJmiXYEl1ccz3aIxZ5
12f7/8dC0ZdSFsxYWI06vm/BohwTKERcePf/yDV+B+u69ohvvybQh48Rm9pqHnocZv8L6wuupgrF
KZbR1BtfrVaHH1lhSuxs7z2wFy93bDvPojLsvICDct0N2KXgCTTXe14lAeTzcKk0a/srTAahP0/k
3hwhL/IvoNRoGOBP59/hA8IUkX2mEukAYfG+HRSpOZfHoNGfi+otvQHUCzsUXhMHvLOwywVkouLW
SY+829IZzTA84T3m2plBSTFbpTI3WwX5CKCugz5h9L0Gti4ykAVlX8gu/X14vfDzCz90r5PMt9FN
aMS7IUWp+I6+y3JWFhgSt8CQpYad4rVZ0N9oAygrFRoVS5cL7nP5IHc7SWAb7P3OMpBUTJQEIU9I
baryGOzNfsCjTECVMXc003nyYrqkSnpx87m5/39j5DhpVdE2no1wuM3OVcZQQUJlH7cCnqezwmoc
xlOr3hrr+ZEsC0tUjahdZrVsS09bf6nuVy6JwHt6i4w9rDl/uvtusyLERXbxN9o76NeKPAAMtIS9
zFCUQNz2AnvI7lQaNlWua2vX74PwY55QLq6/vYDcdK7/mY23NpZMv8B96UhHfhstsDZGT7wlGDwK
bziDS+sJdIW+tLyq0bYg8huOy46I1eul4TbJ6Fs182urWS7IAJu75qBAq4zd+zgnOU5VynvviiVo
6tfK10hEQqhcbSbAMBLNuKpyOvp9Wr0M158H8pkMBQBlUBgd/YlPTFnu8FcdrGUDZQBzrsK3sJwq
TJbtWulGLBvykBy4qxQwbjuboY86Aj3uPq5YtO3ivn9cP0cc+DyQDDsPUlNY5WNk3E+CAO9QTnGr
A3Th3PHzDzMoPjB493PAmOOBnL7Gxawv2eAjelxgboj1XFqMD8x6HTPspvLtRcMLFUP2zsSmutmE
5Z9mt7mUDYaQNiNyPPb01PPZwbdL7QDHWX0IkCZKl6XHueKCo1mC1D9anvpat++Ut7DbjzP34wm6
AVIQ26qqHOySfZg/3ncOUBcPPcajMV/9gsLBm/bCQQi2SpmyE5afLoC0plYTnljrQfi+UCoSj0jF
kiQZ/6yhiaPXf7VG+BR8bPEi8gm7RlfgsWXpkF8Ne7z9AMAPGXTWgy+EPQq8o4MpIy0zrMxg64i4
FUV6XRsyKsgI3aDcYTdmyVix6/JuS8BFBG4otPM22hM0ea/AwttHACjmKEsJQJHDFjRGD43v2nIW
0OENpuyj6AFanfT16Hi9JpN/4uTwQvbKvquHBTE91wRf7n17rJMQ7BbZADH/an4MHwE6oe8+nHPM
fxt8Z4wOCWPjZMpDZk111jcp7Br0ozs5hgHdaJ0NsGqGza1zMmXonpcxC8Tew1BpJJf6jz9IkMUw
1kIIb9vZ/HIwXwarRhbhO00cwO1pCRoM+E8pk48Mzl9xiVTwPeKMPtiGQwIzjPGqItohKxCF/JfB
l/7hVoMqLoaRgmnVblfyaxyWe7NJ3zspfSr5h+JCyW0vAhGrYpP8wSHOdIZ89K06N0zKNI7onGbZ
H4DDwbPpscKU4t6qKzvggM8oZEkWn5yL7wf3RopAsrHUbi1nCnj8ZK+mPalNMi7rws1wzFmFAJqh
jKNKUBmW84XRnDcJtl/zh6N77IWxTr7RinMWdK0TCpbDEKx50OxQR9zrfxYrihdawK6OR3kPbGLZ
hlplCVndf/+ki8oklIuEK2ulyFNYuJcct1ZSjf51tONYB3cbctZXq/T5bVwkb+f/Nlnr+PzA/383
Auh0deq44unXhR91MJc079+5rojWIj0/A/fycQ4bTj5h0fuzFafyrzxZuHTrt8imfH86wfoa9dxJ
ks8/hj1REX08Jz2Me7qdo82WII1WsQHv9XQ06bZZ1BN7u6X9gNbVveto0mNaC+NmW0Dye7Cp3Aj1
KqprWeWu2ZkRHrg0NQJiHnxDCkhQzQsY8AwxABQVhn2Tf2M17fhlK0kQEe7ecT+HSPzEdkRiGXow
w/DZRNPzjGEbsfMtk/fzdG9AbX3uZDKeJuz+RhnM0DyncJGAHBf570f+rOZ/iHV+Ne/TQPQc3hnS
3yzDL01b9f29OohqYpu0uTuKnftrAQFVeGxqg/jN/O6Kt73i17J7ghdDXzobn3c/tdDGlxhZDZgg
PC2yHKQ4lt1uJ+xPQVNpNQT7sZQCzlWG+EsdY9Ddnr28+jLqhh/lxO2kOV3SJAxE3KYkz+hbH1kf
NrHu1JPHumHmoJYJZAikJY+e+T0bw7hqQTVmzvb2kORnfPtv35MBdSHiKfHMQcYUR5o9jvRmpmwJ
+e74ksyMMs1n/hTIc2oYscNfsxiRNqPLVhCtLDwuPGTbqe2IgpxwIVikIZ5FwGSplER53lMbraQa
/WX6Ev7CpYcbQ0fo3upyeOHs4B/0SaJ7S60ddGDtm4fYyDE7JSt4P6r0QLzOKEJxuklvGhf6RVoD
LdlEm3VfEbO/GijQC02egS9By4x++ftSs//Dx9B6B2FS4fDPjPsbnM7D83/QIj1krJbHIERyCQkH
JyBHU77A4FpgsQMtmhrUrstZxgk6aq2JOwMm7JWSj5NMNtVaDmGjhQBp0KcN4D0d837xU6LgsSof
r7CE1PhFLq8XWPj1dC4kijmHLlBbFz7zkWbJ7gFh2z799xShT8xppaC6aU8Wyab1Cff5266aHjUc
xbEBHvEau2fspvmjoiNgHV32gnEUci5qgOo2y/iNVZgOp42l3A9mguXiPdUcSE85kyODowQDzU3X
y7BjpoDJ3d9QTxf9JXe9pbxrM2LsGcIu2FlOGbSJQ9dTFmFMA0RRzN7eRxORorRVD9HJNaGFGfut
5wjqqLCCD16aBkTjVz5Zeued5YFtPKayNpxbbZ4A+7Qq/VYuI0kc+Otz8Md4ZYWBtUrDyWNI/Wu6
s5eB0fiKLy3mxsalmAPh551BjTeajGOufYO+spYwXt08psnMB6TTyo07I3qKrP3Mv96Y34oGB5rx
GsJqB5+Is7a2xgeF71zBvyrxBYUVgHnTVh/nvacEqCNCFP2gbLnOAg/WCiSaxO/XdkEZyT/iTvL3
xMfqFaVScNH+zoPqEKT1KOVR13hPHQ3m84YCfPx5PB/4A4V/LfbUr7d5iSlSlHQFuzr8ebvgvAE8
Ip4czTeZN+rsxeaA8CivETWpONWQXHMDdAcje5kG4bZ2N1omrj4Akxoo6Cqp0rYPgjbNLmwvOXw8
vZGvyYQpQkzO0CgyBP1zvikmy9aGyIM4MLBqzBzFXUk/nUVgi3eMisUQnS4Z4tY4bw4U2nFCmDu8
rVAT1WsV7iHHT0GCjDrA6VkGYE2is1Xrfa8tEs2CANQGJt71OIY9v/Kncl+wwi44AUK9SPHPFlXc
1M3P2a3Yr9WUel/pjlt/a0y9pCciEOGbmelIzCnBzI9mtMX/IIjRNqysSUMcPVaaMDYMaELLcjVt
eHZqj4BM4vjT80134amJxHb8lDPYHmcGFxBm97MOBWyUlt83DLM836nLKL14ToiZfLp1P2HuyVjW
Lef34vHl+1cFGcZumvX0RDUoPfGC+x7/whszAhIo47aJw1LlV/hUuSSXvtUiQvvilW3jCqYH+dnm
LeUUQJtPsh0nWOQTriG8Ca6rRHdpvi2mn7MVKwrJ2Nh8+9lUboVI+DNfUvuBUoUqsyyvVTW77ivY
7lF1iwbM6DuAuuV8kSP7CJ1M6/dRQ5Vzp8UHNDN3rHntjJGOJdym4aA/GMxBtqE/ovW6YPuTgAWX
m9eLUGYPWa1rvnSoaQAa/xXFPJwZHHybYV57w546SwbH5XDSEJb7+TgyYd267Th4RCz5ZUrakHlN
uJOoVFUrwgmEclcpWpP7todC1QfaOYhui5DOl2h0WEih9d1bl1PLNHiczPGjU8nRz8P4o7HmRxWD
roTsOP9TUewmUEmLPJvi6YGMh+H9DATQ7/YG4jowv1M3EAcHDZ+XWuMB+uxB32l2pBZ3xhUgegA3
xQlzb9gQqIeZAi+XcqphxlqIUL3E9QswgpQ+atDydBTzWU4r9OkbL1/YHTwepmNqiAzujcxHMIQw
KvUTytReIO+y5aXjUqgNuctsdsUd9SyZw9m2vVp5zFSM1VbnLxHnTTPcyAT4JGy/LT2H4Yb1xUU4
YX2L8cZpKj0DGiw0XlbAglRQNN1bH6QZKMH3/4Ty5HTHQ43Iew34+H+yBqggvFahhU15NbnC3JSW
lIEUDxfOdRkuhs5gWAKoY+Q1ONPoZlY6flG7oEvJHslAOh6j6RBEHSWfWMfc/kr1jmbUeBFtDztU
uMUBZxCbWn/SuI/wXLVLAi9wxBo5poxtlRiYyvOz9PJN+NimEkfmc8QnxEaz78+JnBvIZ9S8xxI4
C2IrrqRUM5QR8whe9Nm6JsYAPOxrbZE2ON2ioLYhtpWnzmlycm6K24kiF89xhu6jPmzyOlW14Dlo
x3+7ALbQR+Qo041hStxvWpS01Bjqot+N8Yx6Kj4TeqWp++4wGhMt0/nzWSIu4JS/2XnvrrLs5jeR
Pk7sNeZh7OktXqYwVbN5U0FBlHXozYIPeLXtVi0MvRmZdADCg88c1o47i83jSVI2fL/WEOZe+1a+
aOlWvEPXui2vCiribEHX28KXNa7PYYjYKDZkssERMUMG22K6Tk+x4dLDzrLt44CANRRD2YbUdIJa
zHNdeIHJWjPJ8sVrhDFFk/LslLePEhVmEce/PVg0U4ERUPBrlLNM0Ip8C6Vu1dD0rfZTKJ06obew
6syfwAjUC2WhO+M7tRR8LhcCSSHC8Qr2G6D+w2J7sCezH4gd1iWHV/6JCzMGxaGeuHDWlkuA1mCg
cvBkDaxLkGbjes5PSr/I1pbYxp48BVk5kzXQPpnyjfukkBpvtEmjCVU/rx+MgD9suZAOIjgSAHP5
LaJeZvanWDQ6CY1za78PWpCCnLP7WSgzs+O6TCVjeOyWsBCWno8PTId5rRU2VnPzz+nWZLK7yklj
in75fQreppk3HhxPMpwFOs5lk2TVKZh1oSj5DzH00F4MlJw3a53PXkRATkYIiLXYQcbg7UTi3z97
veilLNJJsG5xZAQNHbM6KbU7fkus7rPza4qqLLBu5iGLlzHiyUvXApzAlQ9CNYMNka6a2KSiaLxG
uAwqNfeELyOowJaWCI0MZJ/CZGyyvtDRnYGM8N0+7W70su6tJhx6YgdFNP9DVpW2+5srBgaGlodl
Od4I6zM7fTsLXAD7cGoGXfDcEhAYIMVDbS6y3ZsXCiXy5hRiU5i6/HNXkZxPGPe5EcTTIur1Wxx7
Df3vVelhYKo9CRV+WrpeDA4i7AMqIz6SHbSWzRZ7Onw1k+WjPgVzrc0N9GN12o2uC7fu/Dd8XRfL
Vc3vnKZ0j1In+UCaFJJ8r9MbDF4D3v5XUxav76WPEE4w82zC59D4S4Ajdb7AHzDUtz/zTkiD+drg
cKrP7/VgdjMvJsynWc/Hk13SsHc+/ppuljDI3M4vdy+DssPE6SdCtI0JdfQPHekxPdqYCu/JXWOs
bk5oOxCCD8cMEsA7sGnHF9IvVVHN9TXf4QxAHTYwHz/b9lxuFEkyTj5zVIwIuElFimE8rEy5AzaD
NOQpO3Ptzcy4dEH5NJWgkQHiwv1LaDjJTkdKuOIv/PxmpJM9HxHa4yKUFbtuK5meln+7deo9Ggac
1QxTJYcWcZG6TxsSLEXWt3slDE7FgytIhQar2uCFldToHH70nPEXZWGIa1dh/p3Ers/oRxxDWlD/
siitqLTY/ghThRlnsuLZzKpkPZ6jJ3rcuw3t+N1d2HNFdtGhr7mqT8HRvx9Q5/BSeiqrLSawtO2l
GwahwAYO/zraagjTpGW/BZuh2rxYhlZMZDxIYzeTO7u5alhEOmpp67rkfxdfNUdcHNOwH//Y2XRn
OpAzfvEKkVmhU4PiFfecnupoT801MIlThv4cHeoy6+/TBs6z3A7nGyaQwmuIGo/l937u0vjzpBSn
Rszcrme53aIOC1rzcOQuNKltqrbYUlppMApClBESYONw99ukZ30elI0wzEiet8YXUbXiLVrYHK3Y
4iVuHlRDVQP8aCPUZ0BdVQ+vyct69uOuhDhNavQgGNoZbWM1C+uYIZoiDUN9zCJYhRhUDstN8FF7
9fYyL1K8tez5R/uSRHP4uiFAClDu67MbeLj68BvXQ4HAclf1fmilCZaHex0siBcbCgdJ+EtKtyHi
CPPa1IJqOnMAduIYoo1qFFtLMPoGQjBM9gTaEuhGvQHsUfwZ0FJ34CFilEDWrP27IItgSB87dyFA
xX+JV+nKdguCAisIUwL7rfCplEC9IRtgLry+eZvnDfowI1RRAdo/0hLZgwBM+wJrLlhuEZ2TyNyQ
A4kwyzbcXL8TFMSdsyHKrSb6cd4KfqZDLKBZgpyPx2IMrwiei0vWywPI1LyX0azgVfGQk+C4fOB3
KvbuvXac+tZuRNXH72CNq4zEdwF7qRyXrfioENLsGW7SzAgxsdoe1ohQhd2XsabYQuYVeVRsLKN1
ieYRmQCfLd4bnO5saxBwg9ljhdLgWcwIj67gnVrmbJkQ2QDmYoHIOp84HIOjSbGKa1z5SJpP/FX3
MhKVHOLZONGAJi7vgIds95ukv1NBsGY3c/WJWH5y+1Pz86QGA0Kz9ouxmau/Q/FgrL/4qBe9z15a
bkFfX+IxhQNNr8DGrWdHSwJKtoo0sHUC4ZUEah0qW/oHMELQdacK1wBpElUcnyVIIrVXbomXbTSq
Iz53Fglb0Z90YsdyNuBlauSOvSLEQBQP637GcWAhunJcHHHn8WSGQ8e7pFGvX2NsDe/nezrb1nAy
76MiHFr7qajWDnjThltqjVoWzQypF+98SRijfbXXuD3X77jNE00YiSOVyV7C3byoSoptMjtjJgul
nVUBo0GLIunNm44BdeByoY85vey1oLwA6GJb7tFjTOpjsikeM03h0QZrQ20N5OeK/dnyoOg0Kq7B
9MMH29e5H3yyhG8aTsLGzx5+bWqdNbNaBlziTbBoCat9EQAPBOza909cUNTqDh49/BvH3HVS+jko
8fiDkMl47k9CKbp6Znx7UgTJek83Ibmzq2rNB3guXw12JQ+clDmiG/qjaIYPbSFlnstO+oVmy0r/
ozzFHBOkZhpfWAourcBCfF0eF+w9oHVvLiglTbK7gE7y/3xMzXaF5dB+8CCiozyRFVCpQ/Pl/UW5
Oq0B0byfiOdFbTCj9X+4TVBCMOCC2oKnUfBjHqypuSeKcL0xG9hfAZdKwWfFsq8qNwC6ywLPK3mE
yb52q5ZWolMWeeGdCTsTg7SKRHbpzX5t0Z9tPx1mnFz2dRnBu2G0jA169Tz/sHcZOa4hiF6ktaP3
Yp62mxA1vRsCdTAgw+T3QYQyp0o1IAbggY/nCzuxHainB4iEbT7jeCNJiNkuvPcMUdcFRf8MABnB
8rMNxYkwClVdBZ6sJVH27D3CpCg0Gz5+SPFZG3UlEBNujo/KuVs9euzHeGKbiaM1wggY9BBmIViK
0AcAhjAHhp1TjUFv0fDeF+DN/raZ2VPd41eJIvWavJ5pvucfuHQfmOInQ9zwOzv/4Nonbr6fN+Mz
Vz0Uz1rcmiOLWWwtw1rQMnjSt79gRdW2pwuGd/7H1T+0nl53Uk7UP5BNbHY4B13voroX3JQ36Kh9
bu7k63vLzWnHQYMGyJfHv0dZbrnq1DK5trup+XwvUEGY8TQn+4npOAKOGrMQ2nZmEHSz7L5J6o5Q
jl12SLQ8cGpnkIOZmOwXjBGAZzqFCXVNLD2LeKRQhot9FSSIh67EZcNOeRRccqvSAY2s/KFqkL4I
4aU7x9d8VG7kW7oCpsUNrMEQiWtJwSBFNrRHQWY/ovPVlYPIKPAb73i/aaDBOuPJnY0lqvVE7YqG
H1xdbk9J+7rywI5tkKUgs9yWjQNVxUrGOt23YsuzSkAyQLnQnEKKmrqysWinXtR7GbzuqEmAokE/
OoAVqFH6DSb+kROR9xN97RO9o8Ugg5fVYeGLIf0mnAnkmvDin2imKZMj7Iy7hNgcbbL6MWn2F2//
NSO2q2L5WGOBH5QUZrvTuYqbZO2DjjF3HVMU76009VgbGvUdpKG+xsYolbaTK4xe/q4zIW1u8OT/
cA45x2QQ5cYRE3D7vESJvQojKvFiarQgkVTBln7y24dUvGKo3OLPwZN0iJmGgLC32Wqqt1w+Iehw
m16qbJ3TbvqORlEMhAHlraic8Q78QMmU0Pfv/6ynxVEheoygIJ0n91Joh1QJus+7vECo/3cOyx0h
Zn/yXgxORCSXzsyxW64PeqOJDiRYtVMh4wGDFYKEWnUwB8/HqBX1kE5cBrLYtZGMfYy7sPd1RdFf
+aqNwEWjYe6iQKc7MlW7hHZveJ1g33/hrQxzAYfYR7cHG+YvBPQie/cUn1BdSjreCV4QL+OmggjT
gOcB6YCSUoibdbLpXwlUq+KdQ+CwP6J0A7+rUtlyEgfigxzZwMvyiu7YA1Gwkesjv45FXnlwyIZl
CIfK9e2zt8jyBUWZzIBhY/jtBflftxGy9mzMSFIG5ZKxAGu318x08l+Bn89zL8PUbYAzr3xVQCWL
cRFarbE2SGys+4Ic4bdWP9Mtbpi3/pGMZh7rnealfkx8RR3uOa7Lmd3rhfFOIUE78qiGbjNOsG78
7RLPORtM7uaTi5GnAEmz0Bw7exnvUOTojPEslEAjl4wUYHTTWwXOYCRZ0b3bj3wYbKD0asUZG/jH
kg51Qpk9OodoH9B66ZPyz7/i7/oL0k0HPINOII1QnwwkMbm8Id2e4ip8Ie5MbIK0rwVeISeVm8P5
klZSTZwheFL+4vJU469XIu2zOnXtNE4pZpDiPbQh43ixWNokIYTPsUEF4pPCYMXcPb5DrwoUiDr9
gmeddokgIMmTUqBg8nYBZitPOdxslgOG+BC3BBeOx938hbsoTDjql7jT0aP7DQf+WHsbkocTji0c
LrnrucxjUSTUip7gjtwoFc0o3bww3x5mOW7+QXzgF5I5Y0RO1LNGN2lHNy0Bzr/LZ97D5bONwMez
m/tY4Km5i9oX3iuD3st2tJk6oRrH6EN7UxvMB40YtGV1ujJQA+pIGJze8aO8lwCbfFfYwev5VNWy
G+nX4sPUJdSbija9bziY0rt+SA+b+HSh0OuRq1aWzBOhfPRdf7yBFQUTd0wJPAwTTEMKKyKEGZAs
i79kPUYdxO1quDcTaCjgCYKIq3UYoCaXfobItauNRjjjtLvsdTvhtC1T/xxvSvKMIHIt5h7cT8By
oWm2s434cJZ4mNy70TftZEFhR9qKG7WIrxcbZN+TF0klwAJxx+6LYCGMsuXMLRCoUnkNdD7khpgv
zFCTUmsFK07OSduAVi/KIIof3kb9KqC//M0YRbTRi02fXtfpoUxz4qvFVucNDPIHdbAqcdP6ZxkO
jUgXE0wuzPUsqwxQawg3A+E/FDFgsESsebppHH3oz0bG3yYmKN2AQp/4EmHnD+nS8VJXnS85LBar
ZH99auVM8u8HMealM/CmD5TyMqvW/Gr75Dn4ywTnX558/02rJ3NSYl6gkCODl9aLsyI6/BJKpzqC
w8HcNXyh954/0YfCM1dYQKlEhfsnV+6H9xTNxM2rqNvd1UmS2s2LuXf6R4p1thDINX1yK7ck1pfB
daH1Mpxa/hqweJQqHp3CHC5ZdAaAbsZ8omMMkCAFdOfYsrZJrYtMR5MGQII3/7q6S3oZDlpQ+ERR
u6fD+r/77v8dvgXqrTaOdCuzTxtryfN+4rkxglPFW9rt+iwYr26UoNqYIndsJE+/N5fCUYHczehO
i3mLkWGRimgUT0ecWGtmptxsdsNiJDlBg5gY4Fx9lutUzH9G7GCb//eL2gktxEXL/o9zxU5MD7mh
Sy3Hya6KATZIEj/eaZlhIhictaii/2dJ8B38cHFzyB4tmZcVrYt68d6XNb8Fk56UrSxtXMlk1WlA
uh4Q6qnC/5Wg8nOdbCokXVOYqO1rJPAiLMH19SDt08RI8QveNcodU4uQJutd9vh6T2DbieEA3svu
exoz2l1mwTwFmHz42b/kUb6Y9YnXDfxj3a81vjJlgQobV2akkenAGdjvDNJV92iwz67e4kolQUEW
ks1W3eBA61ttNr8PckkVTD7h+b9MM0iwu9DpVChN3oXrUJTcqa0HD8kfeCEHbarfOjlDiJatvO0w
g6KgszpkSPFzpXOh/GVXoPslgiE3Ntq+Ri4kbRQ31Jsf3TtnD1OrId/mokWhLnIwdHlt2vUxgQqn
rNLsIClBRqQhxk3lMdcfm6hQWLEW5pDhSP12+uXWXzwZrSxdE5PI8IPRcp3XOr9YFYnuE6TET67a
12OFa+ZYAOpmvgLIgt1xZ7bLOlpnmAxBFdiCrOg2CtvVqCsiwkaRVyeEzyyEJeKGD2W4otmpbQW/
GjGpdOybfNXmy2o5nE6UVFOmPEugAIF9USoVOjicN0KS6OaQ8wVxm135DBmueP1fuAZskT+j/0b2
AFcBt0HgIDebFcNoLjU8zWi8GlNWWLKTuLvDvvuKx1B8BXBoOo15g+Y0lb/W/Dmxlfygkamo5Wkw
ZKrxZ8qJvKOlWLohVG9x4dY1V8GO7y15c+OwDI1hIJNHPQFXhBTIu2DCCq75BFVkKacOIqcHatC0
ZLpUOuKrMlRBaX9DHN7fmSyqUkxnuq2OgerafiJwdQWHwHUMx/zm5cwlreYzFv8cBOlR6JZDGUaS
rQA/KW3UPQ3LUi6Xps/l/8aKwIz4Eo3yEPcWYXa+EGJXm7Z6GxULwOrN415H7ExIo43MZzHZUt1A
6SAwQ3v908q0xtzDU/u1j7PvFoZj6XhxMoLR2JywV4zFETnFkOhQV+2XEuhy89niYnu1d77wp/Lz
wDzyhI3djySCS4oFRxbm/9M8zzdyKy4pMIt20uXAyFh5R5A4IPtjQT1ILrSYYu64l5IGHCrL4zyT
57zFOljIEF824NwTrJu/ntme+IEAbpDwdboVIbArEQU34JR6/WGmqOzV2H3nKRZAoNIIjp2U8/Io
JMDu4zWVkQfwqwCcB+yAsGVSF4e6TlggRjRhHfFUETAQZR07wpnxa6C2s5DTAyvkP0Eefbtjlco3
3DMABbqwT3qVmdnlawlukQy0fsuKgCRHgjrXu2JVenEgk8IuDCd82OrpK2PsMxPto/1UtUhWiZXO
woHg38C+Z+QtPDXLVu/B77+6jD1ZopfJk5VT7w+Eh9bZ+d4A+/0hkwHK56Asngx+c9GknYQ5e8at
BFprJfKTIbHGD6wlAoOKRmRapgfxBLrANtnNmIQSP+ACoZv4YKL9mJAaW3wrIvbuWke78ODRjp5T
jDBNFZRa7oFi71k4b6TTl/pqnOWCUVH7Hig9WypQckTxt0hQg/1jekgvLZp0UikwABEO6Aat88FR
cQYp1UJoB4wSPJTmFqZjwM835SWr9l1OZst+X3DYEbzeeNTfcy30sbqbL+acWZh3ad5T0S+P6of/
5yh/0PZLSTwZEKErvytHfoZGa8560trpDEG7ria4OxRMvaxCwNTGCCrIYybwB2h1vEXCKucSmJOL
hvpfpfS7RfO0eolKxh5DV2e31gBHz8q7yGJ+NSKLHlG3Gag6TGHbhB9H2XDKg2JYZ4AHDcIYDxYj
Duix5beo2hIJSQJuVgk4N8hRbctBg+LI5ahTn3r6OP7iTJjHROnBmhJ2ndcE5dCl51gd+UIo527P
B7dIcxiNnzBxTiKXzJWPKkmr0UmnVMuslgVjJp2waVdhtpb6mPk2CvQcKNvv6vea/pdVP1Co10wg
S1PbnaMCeNEBrf6Aj5yudsKzUQrXT7VW79R23QjFQQ7bewrT1RUxGyotYCyPn5j+kQ3ULcgsBsUg
LuGWnTDxWwaRDsSt6ja0eNvvvQeg8CrB0VvFitkN9pGC2jK0YsSnrd1mLtp7T70AEiyXUuW/Pqs6
XJLqMPaXJU7lxldm+r+/l1F39G/29kdPiOv/ssYayLLTMzHDqIkYhPwMOkA9yveXVpy5HuMZqgWE
cAjVZjcbivd06iBgR80xHiiDWk/8AdHcschGVCmwNgU5xEWgY79Ct04BEndwCLCwIu0PWJ527Ueb
52dLroCGlyR2NaV5VCo0pAVzM+PIE2rtP5ENtDqlpOB0VtVQcCLwAfu17/l407CtKBEuiosFHxZX
7fmaHPKZNVnkNGGS3AADwBV8V+aCIzc1zxgYEahg/6OikSbxb0Lq/kjuOlh5aBrEWzMlWlhNOG3F
L/4CkLaObuQcd9VjKLxty2hME1mZiS2NWoRqNyK5k8tszLoGeYKVYgo9eowmaxe9RUKmSeIsGfwC
YfL49JujY6NDmZTES7O9U/TaD0CyvoSYdpEioRBo/p7cH6lhLENKMoZtxg55Tld+3RWh17+Nknx1
Oooth1FJ/UDZ0dRNrd92g05GSIBBPB0Md/K0LkGlUKfvhp6uWWmBMhrf1i/2CkvnQLMyNNojc0Rf
7frmivX34p+Gk9Gu/w1zNpVIcbKPFZ/gfY5gDu3ECPvoccV0xAJZJvZWoubyCTWfQy+9xacNdD6B
a3UzlxfNFAznfj7MS3QN1RCV7IGRlGbTnDS6WikgBFMO4CQyI1rBAKFNn2uKPMEOzodTsEJJ21Tn
0XxycxKBJuixTPZ9gIwrV2A4Id8N4qhDYrlYCAynM/2YnWVBr06S6PjwpQaYOtdvKMiSc1XUXn6f
1vltpJNIBdBDRYZ1vxabSd2XiO9HvSRz6qHlE8+RLFOvFUHlorxCZnNEjx2SQ7vT3xtCBmJZTQim
Vh8oayXFDTE8q0Hzhqc8YpFGv3W7kUHRqY3BXgGAfBU+2xyPdnSJfmKR0h1f8V5B+YNW23s6Pt6l
Kw+7LIYJ/CmBnH7Fk9VA09yLNu1C7Yfmt6djYln15KZqR88hyOLtpwwc+H/6gEQ1gfWWAqlj/9Lz
Bg3ZKiIl8AMNwKABSvJwCLgaq6UGlwkrYGNofTDRxPcGyn1XJhcY5HaRvAaA+bRco/vZihhNXUpn
BKMGmel409bk+qt1BmMC7OM6FWH7qcOeXnKMn1hbHXDNcGcAOnrc8pje+bJ6h+QUcVgVP8WYqI5h
yUw3MDh/+X6IGqn8KOdwCwkL8QcLsMtlkv1PduBq497Szco9LhGnzus7dOU73e7tdhek/nkDK3fx
HlwTBldaiQikBh4/WbeILhe26V3fqyRF9XODpjyRIbpBp2qjtrfyMoV+vblO0F8Am0pdglPtUj9u
K16ZNaU8/P194EWiwpcNLln0/qsoa6i96J/Ldq+tK7h+GwcUdLhCCBHwyiA+nPUaPGcq3X5voqF8
94zTvrIxCSowXmR5Z2MkAfpLqcnIRecKzHZXTcgP+6O2KAy/1s5wQxstl++UB7J0VcTDgIsFTwfB
0WmGncS1yuODQ+VwReeIcIrEme73SZ6Oxt80eC/DDCgJgyr2Q0niihuxWT/ELS5XhZ1xhCuhP7US
XnCm5TPU4BrqoKf/ieGBRzhJDrCsL9Wk0lzTiCqB7Wq4SleICSIyqMYn0HSb6yqiOkxPzMXca9up
qs/A6PNJHglOU2rk4eEDht6K2C8LpM/7XIPFVXs+/EvH4DDdB42uVO3XA4piiBBcoTVCsAgGacIq
UIO2fQ1fSM5xZpfaI1lFn4R8dUmfOisfExyo5wH9a13hHh4hB0T3MDNICSeH9nEjowJ3RN284ZpZ
hs/Gvy5+itbclvzjhy7C1mfeVTnZJXDeP3Jqxw23aWyzDgQV8DxGrtHxLwzMbQUaCDh6ZupRglSo
gsUIlU4jsCMotwdMD55h7mmbopjYjnpWUPf7uJ8YZKuT7mko87cjRTMQ9ujv/pYX/tW+COfo8/4y
Go4ZwvIKHWplifjYF/NzollEgx/IktHU1hjOIehvDWdOITxjfQhBgMtL96QkQjDviypyh9rF+hbC
1a6J8NUApzxO7OvG1/lRztXeB1Jf8BfOYqQ7bOBPnA4SXgKjOeUt6byBmAS0UbhsftxmqlM+Yl5s
p9wWEJ4rY5iM1V7fByNox8M/Y0c4McceVLfsHLTY5gsNU82kPV6VE+qMhjO5Xynh/dc22iLXK+4t
4LkLRKts3M0JUamyQEhepx9fzx0YO1XGTyaDSuKyTc3voUcp5BZwDtt+yuJLCv4bovcVMT9F+jg8
1PSnlshNNcnmg54URyhObSTLalQ0h0F3Mp35fYljsFOMjBKts4cavNSCaytc8AMzgSIphKEsluUx
Z7cVa2eJpuufwgkmvcv4QqOKAqP+M36Xc8h0Tbc/uuOYmQgxVsS4dNxpK97hdqs9/Sik7U0rucxe
ofLshnsT+3/KT4+yWNRlFyrGPosNCPYI+gkHYj8pn7XsGYFOI5d4ErNHbf+w/5gcc1W9oS0S6b6M
1Vn3Yt0jRWZGNEjKqdvcoC0b70jKBrriUgb9Mr+gXcW2lxG8EbDUBIJMB1/6Q/31b/YKKo621jbd
V5eO8KHZmqa4stKKIxW6A+5g5V/9bJmL/LdS2GwWJ2XytYLviJaUWsaDXWI6RpiQKBsgze1sxcFm
m+tlIPaEcOjYcmw+n8G1UNClJbo0El3ka4N/ZH/0PZrOF1skUYZEme0XgaUUQgzXSGDLcW+25ug1
yuZ0/KPjtBLc5RpnZbzxM1A2G88stXqRxQTjr4IxQMq73yz1QcnxAiQkwPQ9a0OPvDWuqv42wqVV
Nli4yxOY3xa1RVBVVgHU5yFZL56UqamNn2r518Bt8QHttq40TXqPA7wYVh+kHEYJ4ybHgHvyMrG9
Mng28HQshbIiAf2+PAwTOwMv4RgtQfVeUZ6936jA2w0VcVkL8EXNNs2984KjYmzoWEBKKGOaeiPd
bHMx+CSSKwdfjIykDtZBH0UMSoJefwXbT/ov0UGCJIwD9RhsUxp73veLolTiHpAhdwVuZEdFSAl/
eLrMOTQE0Wj+gmUQV17C0ME/KU+c2SKhE7fO2ctmNMwLEr7wMbxYR+Tocc9sC+oeZaX5aOikLAOb
ypy5pS3awrMKKWfIVbnwerlrTzU2glmbm1n2afKrEvYv1G70EpyONWh+12Ib5e0/yrTmFloCfpWT
vu9BrIvixcBN9zgNPmAVvlriaYXTb8IJmPTj+rQuEXloZx65mXzqVBiHM+C27te5bNjTZbTz78UR
afIUxZsdWW68YI+nOJ06t2zkFQM9I+vS4wsZaQkGQqZL/Uz7WTGeVz/QxPtNKCjl3aKi4cgDYCpU
HD9hMYlzu3l2B4v8AqM95uOycThj6dFGabXdVlcu7NbD4m60NvnBB7VuG+NiBbqhdxfyL14psxz+
2zD2BdiU08p8qNavxP2kUIFQb6s++eBdMWEpSuvFNERtT6d0lNIgNGR7iNOOs/u1J/bvBRKZWMLf
CdixKevSRpHGJdmmC4GMMAdYlBn4DEC5AfdDQQ5hVOb2BRS1ZCzjWPFETC62G1O6YRKK6xj7AuZx
eXzXNRnMo8CdueiNeLp8PkuPOrPF8ZpHNEQ0N0W/KvMtAZxOyMTRWwleQ1y1a11rQnZIvt//6HqF
ncuSZ6oRhvIWBJ1gP05nFi8idxzQzt1heuQENSFdLkQJcEg6iysM1WZrI1ClpDKHb3OCxPHcKrtE
Af9ESg/Czxu2oqWiMx/VjRwom8S5WCN8R6T6ywrzqPUYErC5Ld/mzAig8lySrJbesKJLZi4B9oil
tjfGqF8eboYoILM6X2SPq6/Z6WlNVP6o6WqyFYhL8tUqKhy5KbOLKoB8DY1QwuMoaFi1+YfgKeOb
NmM8opyOjsCVK8fQtj0zv12b1VvIfsTliuA8bEB0fNjAL2lsQXFHEO2gNGp0nQBgFGqeShMzp8Rd
sKwuktJzMRj2IyWNWfTJU8tDLdtBstcN5xJ5VGN6/QSJHKH88Z27H+d43aaIKEtzkur+dj70J+8J
I1WdsCSJFuh8IV3T5vFQ1V9Lky/g9Ngaw6NhZc6dStrmTBi3S6MRi7cWW6ctKp5Eg5vku+Z6iUmo
Xfr2RV3yemaevCX4J/qr/eeFydSJ7dyy4uDjWBmJfM2Wr4uYShZgaDW4/FfwuMVQjfThLJbmoALP
W07Rj1/kVTTo7+K4/7fOgRsmNV1G6IE6T8GG4aT3LHIXiPhoNoUARrl6vcrV2B0cVCAeyuvCbvDk
fY1EXAQR8JMLFyNVHNyaWl3Mq3Lh/SJgg8rYMiuTQovjTHV67UjLp0Aad2iXbdW9EnG8pWHktBZH
3HqG0Ny4Ak+wsr6YpZhmL/eeZMdoPTMVcTC6OgDWiSE/+xY6eCbgkBI+8eRWWwrRogP3ZLXId/r9
U4T+ME9Io0nD34EKZJ0IWNxwTVkxK+n3SZpDIOUqmo99gIhXbw9ka7mSAdvaQ/gsBKr3oxxtzbEu
N3eHqjNPEHUQXtO8bgAfM+pKXz3q0vCUgv9TXjrR95aAcZfH0c5WQg4+W6d2nx9jq84dQbmhq3Sg
EWXer/wHFnhl+H+USNcx29vhzErjR4G6mqDcoqWKr9lCnm9fi7+/A6CNmn46F2OmJnxT00uJugca
TGTn7l58KrB9QuZ/N2AmAt69ag12onrrxUbPxmSZmQ+0f7S+GtlHqCERKf9/9MJtXcoLVYb5tZxm
AKuyrzsM0kQqIum+LKoXDSNM+J4UbGeWgMhtolAkgH1Jz6TaEPw3n26fI3861JwKSVIPp7kLnSIH
gej+nqapgoa6pG0kkzlhwRaQNm08o2bB4JC2AnFbxdbtKMyunIJDHles/JSA5m0A9Ab6hLjT7fKs
q1R+eCqjmh3dCCx5i/XDCzutemS8OLcvdpFH1DgLoGZWZ/VpeI1mnQN3tUHqjJhWdYraURVrjKLq
zLxqPIO75ezqNz687yyifz2tv4anCVzfniWrSiDo1ZNy/rL4R07HwEUNJtQ1Qu03ZmN1IZY9CK73
6os+yCJHhO1Rxczu4cM8WM8XNS0tZAAv7m9mkBFjvge+cLQnQHTTjIA3RetqoreGhqe6Mq5cIxGY
New+H2PaOdswsvMUdmcMYDCpZtGV8sfm66fkmv0l9mPENIHGf6S7974IjW8z6Aa/5h4e5PMAdDHy
tjpASwZ/jcynbD5t0K14rAL6eMcID5p0tUTY4qc4D90t/MCxf62RxDdKtBpnMpgFNJKbhh3rRAGx
Qd8dFgiDWgWCOiP221L7ukg8l8RZS+BtjwQd7jLcrf16epbQDNdwbdia4F3GwY27syNCx0Sasphp
YSZgfi7fgeohJwdz7H9k40jDokFo3BujirwaZDZJDsjGWsLatn/ovbq+9lHvQfL9fZLlFfNJH0nj
R6hRDBr3bB4Q53/TAJ20jI4wHrcKci9ohOFLQQza2UlbN2enZouI6xFETPwCXmwniRn80fNodL2z
nT9acDV+XmSqTV7rabSELGF4ywxfnivwyNFuERuXvfLgAnDEZzbEPcmuTEVKC/DAFkXdFx7fAnGb
itD4iwkdIYOIArnxK6nNdfRIVeGzEmCPt2+ezX8cHedB5Pnvfg1UBmpz22LN2ryOrD1m5hmtvC0f
05Zm3MgJ4ynxXEHpnHFTkNQLO4BIljWE2GUvseJF3n9e8IyQ0M8RV1bKzKbJYZADZKsKLOl1gLRq
MrBLQfBHrdfyvdptNKsPzI24co3rPNFjuZyrR/BhAXEulPip1nbmxxEW0mPkJ+Deex0+GOty5nLR
UUS4zowbo3TNGbpsPTQS3x0fvR/4cL/mFVR2le3DsWiUzh1Ky2ZxVuh1SgDweK5/ENJlgMIM7td5
rZUnfIONX6mlM1iF319tEEn9tWcWgky8BVjmRmkJIpcH9FxbGLRIZHlw4gJlm/fQpQIV+xepH9eQ
d/ZLDhdYovYkI6EKsQFumk/8knfIiyKUiK3D5LYrHvgz2Ke9Bd4NVWkK9zGYpZzNYhFtttCe4u2Q
9PG3vtDFPuCSWisySIfOtTP3ZoHrGzTU0JGo6j/3y0wrM6Hio/X/hTdiEx4rh3LYKGZWpqeNmU+p
vidOsY4OuOcogzJkm1A9V6cCc6Hb6NyyPWgy5ZiFxdoJzSbPFnCRQSi0G6tfY2L4poOdBHHYVLch
PXNQ7ALmgrjtZLBP8D+hd8XmECVUh8mEaxzLbpMo1hLFdiJ07LzS1VK3vOI9fwhuRNGjrzQ/btFM
f1kp3cjTj2+OhWJny5dPTbOw9ms+KU9+rUESo85U1xARLvLMSWWLnxlxDLrGgkgaYL0l9CFQqrNz
UnbpnePDSIhLzO3ebeML//d6ON6u/OVsimY8BQ86hSilCKTsT2+ReHzB+s3S/3WWw+5y8ppu0qvz
BE2Ev8oIKLpQrmArcuyy9ID2JGzQ5jtyj8Ml2BXRKGKg3jI81OXL30L6Coo5Ho97R0GC+/zMyyzI
eOokcni39tGwon59/fy9QQfbG5eX/NBuMH8UIYhFfZhUND/coK1N6u5fyy7KeSXIdanSd+oGgVql
jrruL7hiayMwAEWxPXxeRS+82iq0cRQMj6xuH44Wia4XFadsKNgL0/ugKf+sKfTRkx1NALjbSeJE
SxjAbsnriHV5wAkVgz/TYJW99MGozNHlG/BaUvvL5RKLVFg818O2fngTqq9p/Y9CNFEQ6oeBgrxU
hEyZaKWVTSd1frnZig+mrxJKPEipfanBvGxoBUjYdhC9xVJoIamuWwb7QwRiOXbgqP6IuaBoTssU
KAVwT4RU1SUpjnjGYSFYKKDfUG7/5BBR2nZZ5DhR+3xgKbznusWv2m8QtrchKxHdWrBwx5ih5t8g
8vrJ4OQ1E2emQxrSYNC7hkMuEy8kRxfX5/RCD+Kd6N5vEZVngURB326YxdnIbe2aRIhP0PehUYrL
2dxE+BeKQtPwAgU9v/dI3d4fDgqbRzzTLd7F61A8IQk7BFuu6R6ZRYAOE6ksVxXXV0VKT1yNac23
+wUDRWk2A/fa+WCJJ66L7fpZHnM7PeGWydfpIgc/fn7gpwkvEZhXal0aJS/sVlR/j57HAsbuRGm8
gbyB0l3w08mjkVRGCIMxNNBM55CZ03WUtRLi7WWCAlUINK6M8HYIicVVun1FjbjTdCPnxpA4Do71
5laowD6y6LFN+6EJICfmvP4pyYBIGNO/eyp8IstCIpO53MAdvlHE/JY29k30wpqj1sG7mDHT48rN
doCA2ilK27OUQJ71ExaYxsvlAqkNrcFAyxNer2XbVoKtm32RrHBIEdHS3ME+4p522TvvGwxiE4IL
CxOPGCtAcLvKUA23dQ2am2TH8f4kRBbCC6RfbIULg5DF74EGDMMb1dODP8CCtBhWWt1/NwcMZ4ZP
E9HQ3e49JG0spOiR2FUFwEm4rVJISbha4zNdrnS+OQl4/I9v0TSKCYodKzvhMFfPgHELEmbV6T0t
WGosM9iuuLnuAU8i1XjWuQ4XeHd8bMJVClUGcOFZSwvWnFY1EO3LeQACpYfQh1P3Ou0j7KgLgRJY
ViPxhR5hizN5giXRgSXjjSmsDGCH9XG8rt0f+XdPCh/trFQ3wdET7GBv9ygcgdMboa2HfOK9NoiU
HYaybuRzxZng99LQV3yqPXViH1+MUUdhvySYDXn3TxKi5RfwHQ0d2sPeLwRWH9okr/cBeF3oaKnb
wnkVD4OeOAU94Qcozg7wJPgdlu4PvXUAvnf0R+qB1VOMwN46VKCIU7zwJH9YhnXBtd49kDkUDOig
c6k9rTJUagyAZ+kQlxJOn9FrhgP5eKFcQgGiw73uqdAwTgBWSSZxsFr1WBuDyd4zV0p2b/5iPIyJ
Yfd3yK1XxlvraDKvJ9SjmqLDE3GAuS1C5RWS715QBo/JZq67izxgyHLp7z+M49IcOlyTgfoPpNGu
YjPN+AiVYDOj+ddXHyyLeOLEzUN18vkNqWL2nZoCZ2fypwLH75oDYJmbE5oqCU2j35C+3mURT+yG
aqg6o8W33d/CrGKCqEOr/5S2y3uCFt78yaHfRTOVV6/crASqL8l7/xgBN84S14eX3SXiKgRbGlZD
nQv/dq57MfYvmS/P7A6bSkpx5LqpISLV/52jr6PNN8HSJQkMWqQYgVQ4LqDG9PLa4N7EEgYQ+dEi
alzsIse7s7Rj4HBcl92okyY+Uwx2U/e3dFwaSLOxiZyfQcQVPxzZ/IcY/zs1YQAqhPFhC4a5QxHi
OcswyahSsNOPsycnf6NFFfjXRZUa4Qcau0hQ9SqsswYTIWIQokw2MVWzZTIlaxKs7t5XsZYZqbGS
bIhjl2cCBK1/umapXFyBygSEQ0XDRXiXIiQQ/CYmiyMjwkW4x30jSrFbsWqzGBfKXWRaC+BjaZFf
obkIGQ7ZsCDMG8uFBfs1FgLYuKnqM8wyJ15JKhkj2h9eO82UJCBZZ24B13DrVPrM/4brqDbwfY4L
3RZi5/02uLFL9Pwn8nYKPUugnp98PfZ86lK60BV1S/KLyUKJ6JVGfwaBcVmAoTzmv56SwrGqBvRI
cDVRfguT01aacMO6wRaPOJ9yl7Lbur0Dx+xIX35zbX6UEpy+mGVA6u4xcagPNmAWdey1j4Qhtobo
o0yu5Sb+CzSysP5cnVqS0eDy6kBN716rOD64CKVXp7QIMoxkEYSJv7BP7yI0i5gWkZzlsOW0PGzx
AmtLza0jH/M4jEz65Z89Go04GZKQyBKc8EKZJ8ajrWwyNdHoHgOEKnveMpzalsj70Hyx2QeYV2i8
RV9ED0JEiJRBXEb1tyKVlMHuXHxSFsatLfG9iAU+rBVPD2wPsOG2P0YJlZQkJb55sq6YDV8rL9UO
j7Xug44P5Pr3d0mZYVR4czmU+aMMHWeprhxd9rKsIdTVfyB20X71pPrguZKtDZYd5oiTuEpQtPwR
gM9BOyL8advTXlpHim8KFIIAvz+JSb99xaLtkTWgsTs3VwDY/laDakJtBmVuvhVJEkglxph21bGL
4CtakJxlSWp4A0ppT/cqbiTab5ivoAh2mAryeGBPWwF0Z6iEQMIREwAvn3m9+sYrJnQkFo4CnsNL
ExSIMhiHfzaR+0z6QG4IRJ8VOV6mTTbDDGcHhrIwN9sUW8qHYEcVcicZkz508drkNY52aZ1ML3xI
IUtjXtTnzq/4g66chzccagwIDYsN+1d/zMm5R5GuV6GOZGm/P9Pt6IZ4/yNmVWjpTjuAeBR7Y2Ih
RfX/As+l3rUFNPdPTajUYX9Ig9okTkXhcPEyokOX5KWix53IYjI1xmmsGEwiB3Mr1zAWnp/j4oko
rYMiTvL6w5PJU7s6NhOhGbeeH1dNRsy242I8QqI0SjzGuFM8tLCJqwDTEuIIq6xpmEqO2A40exg8
CWMuBkw6ScqfpMR4w8jH/MfIwzpYATPhs1jo+yWf9ppjvPstYsjFONtXq2mhqaeQ+J/jrPRx6QoB
M2a+vCRUBSMaAX0qjCPpGmznCS7vqjqqioSsekkf9mcqSUfvk1JZs8xJh46kdbY4JVw3u/aQQHe4
qe8YUXb2eXMOgOxdD15zgXfJhCHkegCV1qRZ14aHcRREdnJAeTBJMfoIpSvn1jQtF98igxsGHdro
UUdwFkceQtc/kv8PXYKTkmKHN4JKn2EaqH5bEy+NiuGdv8M0qOp8Mm5FUUcuuAmktUlnDVIsqyLQ
QQLarWeBognYl8ALiTqQKPICIEmXOUV1mSuEVQt2PblYrRdHpPVmj7BlzVqy/qgwhc7A71qaoup9
X4ILlqkLI8/Tyi2bCo/8L2o6QPOz6m3bj2mgv4PN3CZ/zntHC6IA6mU9ZFXenDorJu1Iwk507yrm
68PEb3FTVS5MrzhA/MP9Csxa+wrFynKHRVosWQCy9/+ht6S4r85QADk9rv7wnzj8jcZvafOOE3FB
G77BE1jfsBm/J2NbLXWhmmfGT9NoOkc7JSVNAj5lfT+0XyFKLhQDAye36/DTL5ViD0gmpQTctvLW
SRTr3STj0Esm+V2vn30qY0P63dr++cjr07hWyDj81yu40jzpzNiHLqBCqM5T65KesQvyIl/LI5yc
K7dkUGd2p0wirvLXoJbGsPlkTlvHyw9QGwCPAo8CSzuG98ZL5AEGE/ELIyLNJ1UdfBZ1cD2s2Xwj
SJ4QClZOXmZstVLbA1VyiLJUUPfrqWLe94vOEucqf4mofI+88I8vX6CThwjv1442JYU5yPYC2/Ho
mYp55ea8Cj0UXkDUPE3Ly/3IRH38TWhyxYDorICrjZrB9Qmalo4WXGhxNMERvVuKgG2asFxqR3eL
K0Mqz6r6+iB1PTcjt2/Od9NZlRZjyKshnFHkJ5OWhLvs1Or9tyJLS8HRm9aQAS/SUJ343TYXFsji
WsvVGtmsioLfswUudAE6WN7IZ0H+sKnB3zSVB9Lm/M8VgGCtE1ZWvshnX19shUmQa0w36oz9MZzL
7QDCqNsSGcMsocY6rOXkcJYPRk+OifpnzdhnB3Cv3lDaocKL6jdXgrMhyUGjVBa1QECoILtTNuue
sBoaKq9HxPzJWaun37cLWTaiwL4XF16jZ7GN0eUHOmtcCM7+bvDkCxJAuSJTXsG4q5zNzvIpG2cf
pZQ6nZBiMeNtCuj8Z3VkxAJ2rRvJTxCB/yxO92FtS+bFrQizdR5rubC6msG403FYKPBqUXPLvbVQ
ipyzYBKPSptYhSA3/rkgqMg/2FJidSmpGJ599ELEyHvTvm+hfHXLbms9oaUNn25AxkB/fyjbQEXs
cI+r4Llsd8p30S29fAuo9tgzG+BY5obW4Ooqf1yv/5GnL3rpn4y3EZSfJUdZi6kCUkLNnRkry+iK
2GO0XT4M3PylaoVU3tfAvlrWXlpj/qbvWQ6r4RHG23QD5XnlwZ2uNHiI+O/Fb0hV83Xs4BS1rQJh
S/sdlFV7G3gEQERSGOf/HXug7gY9/VjenRl6tMr+bGuyKeX+K9hOtHfVCk2hRl3ULJInI5JroQ8Q
X8zs0q/jdAK9DBiec5n6fTSfe1jsahOSMugcVhS7gIc8PEjpVRAhpMMyEQZuw2AwUbxzTmt8nfV/
aalduyqYShvEy/NlJ20u1zxLC38YJxFW3wmfBRZY7IO8LRBtcEZLD64njYBBNtFQEuoUYo2Z4+mt
fpeNkeIhaJBnpEKHbc1c7Da/FIVFWW8sYN03wQUokwhSie1Y+tpadVF3Hg/rgWgojlnk7ijS3pPu
FTlxg8tuyZvkV6YeH+oVXaUqRT4rabLoe92ndAQQogXr/Bhu6L7AiBVtFU7TBdtzBLYDvLCP+4HP
4TvzdbiPq+T5USQPcedMvw4n6gaXFxe3cORQDAaWmTX1xhPm554z/XRZu4jhgJ8DewY/kKGy47Td
rflI8vNXXf8fZej6Q/kTVcSHjxGm9Z67cMCdp62mKD/wTOakws1KkppH4V+b1tn1M1T0OvpgmH6y
Zl/1h3FFWgqcepVK86zXRYbRc8Ob/TBPJxQcLWRJcF1PUcxDpwlReTjLVsS7PGf+m4w45/2mn71t
Bjht1k/+QxdUdPo8k6XK+u8V4F8S4PbfJ9kjT9HMg/bKBDj57wqj5wDrJ6Ib42hkeRoXtj6NsMVe
vDxTwtL9Dzy/9qGJWw47Jo0pgQ0S41blgNRO7or6VcJtnD8hmbsEzluXUnKlXLKfzqPB5pAHh0sy
GD4Pdpv+BHrbK2f+hAohI94yW8BJ7tcfPeh2JpsobDEX0FtO+r7XgMyjfiPL7HXbvKBRzehTk0EZ
IHnvEkidNExeU33WFVBGZcKDKiYqYNll9orkBdq2otTF1WG9MfsYpQAlHFdcK5lCKEfHyVMgf8+G
HJmh8UyE7hL1HBOhNPDEoBqqEkPd7knJXAdaWMcrPbKyXzSBkC5TLEK9MG/yDIekly0DxZ86x6Yd
LC3z5RAorRO6D7USMYa6YVc/Flr9dCprFjcwGkQ1bp2WSccwOr7xH2Pa2kZET2Ty8SFoUv/sjWQi
2mJwF7FHSZPnq9wGZxiPHMIrw+Vg0QBw/D5Q+dikVvUIJuCJkrLJJ1BQtOpk56bHjZ280MQ0J5+A
IZ4eRk0FxjO3fX29t7O8l6Q56X4DYRtNDy0Qm2zAF7WsfHksKqAz4aGkTpbOiirueWJyREtk1vgo
nT/LRk3Leo87w9/BRINntBTZW46G5nQ5YzDRDGX2ETb1rFWRo1gfd5DHd371jmgC/vMh7qEGwMOE
ap2I9mlNvSCVPSdp6BXT2skI2xrQn8O2TL2ozZWLGeoFCIIiUJHD+kUnC4pfVNjowlh9psQlNgmd
+bLZxSStLqUetWSG8/20qx5tSIRq5VteA/beAWUvKMR4L4opz9yd/iGezt5wcdjnH4YKS+U7QZjr
XRpzkbPe5IPskaHSsqmD3HGjjAHA1a30kLCbhbDAW/W+eca56vzz/UF6NsLVOz6KEycZCZwASV2P
CyfSVRbCdGC4PP58E3/tIBnCNx0CE2KLaHZSRS9rtauLIzSboysnJMSvYDWVe2aPS8AJ1xoSoAPC
LdbC8w4FyyJzbmvrNJ730AT/DeNOXDMXj0j0ydkQJdiq0eJsdEc9zwWwsJYx/+WOiTCoRJwaFF5i
AaBaQ3Ms2yW5UXOWPEoEhEJjEdHpNOU1rruwsMHooiETUG0ltIbiAoJDoU1o9yAFhsPWJzmJ07HD
5u6jj89mE+hubXLL4CkzxuPN1uJU4LU3fp3UJyNW+9NbzRto9UII41v4mFJumIztWyFsTeLQst3S
WwjePrstJp5oD8UTteIsskhrYNSSjpXKozUSyMjHb5kZwxECrwHvEXx+ofq5GOcg092zwmdB4hLH
S+g9Q79PJ+1SQvlXvCffvfwXAFddwNubooHmg30IwIviozzz5UAni1Uj0TXAbZ9+hm3wsirbS1Ei
deBCcqz3c3fR5NcAwF/lgvcSQAOHATWaa63JPM3naYZhE3yvM5FbHS8t85yoDfGRTAAAJfrPIeZs
xq8ZwENYIKmBckAZAg+S6R5OfC5+mXzxAYM8mKIZxZlc/EufxfR3ker2bcsS+/lSU9DkR9fcdnMq
j9a89PQ0Ld9GhBWW1T3D6vZ+n7P9H7JK04v2Nf9L0HBX9n8SuZj31dQbmWdS3Zz12UgGNd0u19j2
oB/wlctez2smA03qYPavh5vx+L5XUF5/aqhAnzjx1HdPlUA8KYeMLsjnj4vYQw5JxYYJjR/UAkLh
zGN+XsN4y6sUMhrJddaqBaLKMxh4X2azTj/4+WDUTvQi1dfI+HZYBx3JYji1aqroeUimgBuxrShh
1QCb1qLNyLq4vh0aoRo1qhPuc2GetA64DY9wuvKcF1zzUyTNhCXsr9uLyusB7Ubh3Uqkr7Lz1Ejh
hTB1fSy1rTVyHtVYTig7wvKiLJRMQ/vy6nHwaFZxcx4c/1fSEnlRjrhrSLg3Bq76C4HlZuABh7l9
bo3QJJCXK2I55kYQdEelz2zx2Wd5Js0rgRO/ocC5JF9kG6f4CBlaeW6QgPFekcGtDHzDxEh/oxzf
KGR4plHHy57XTx7bM2j9gCo/ZzKb7tX0yA15UseVYVgRScXRdhuOq0mRAX4RdZCnwkpHB5Smy9fb
DVc2AabPqZ8SwP2AgqTH80dXaX/ncom5V3PiX4nKCfsbye46SetUVWG5juv/Xv+AdqPJ2EGifwdW
bvgjG3630QIfzoRjZZk3xMRbVe6DDfEC1DCMEvNCZAXeK7VCcSxJw3mwDjiiWYACRkikNs1O4Zd3
E3BNK1Drt4gRiVrsE7QChAIekeSU6gB+KEmn8n5nE/M15r0wHhLo28LfONKfH8V7nyPc5JfvMjlg
orRfFKXDA+dcGTCwfpB/KgiwE3w2WVMYhs3Tb/VLnwR2ClzAgrC0CgKbx+oxTlOgqMRo3zV+sgAb
iRnz9KNMVo8K5A9egjjqoUQnPCsIXGW+2fPrynfDc0eadV9hvmcji3RtZ9IJxS3I0pNQYNR52URw
Ur9cGgnoZJEJ+i+t5NkxFTY9BO0fcxVZnhHZ5N7RoOsgDif0kLqFfVKebhh6h5BHzaFJeLvrt2Ds
On5BT18cUiDQtiup2/+uIVjYEi+ghzjZdaB1LSYS36jGDxmxho/7NXGFyNNHaK5SerKhMD/3KyiV
KLxJ7fwuNTqTGWEHbvBVr2yFC16LjGx8rPJM9x2t3SG/WegtH3axWTpar+04fVqGivZKuFyKRyw8
uRBv+dtO9HCEEEkrrlYo1XKl69Mqzqkc9PJ6/0DgF7nVh96kp7Nb5IZjo70EmrAcBHMu5ixaxkeO
JeLvvtafPnCcxvqZkDm/lXsiSMdCL3pHRILxjVYNKAMLDA6QbHMYPfL9H7QzWAlRchOHlKvozLcz
85b/BL7Z7H0NrvK2hujX2FG0JkfXz0uVgIW4QAKoEWzxcIEWd3/aZ/LygsZHOc4vlhQHa5YBRzu3
Bff6rsXYBEMSvrCK50nX32NGfSD8PiDI5sOj1dl8dYk/OKHmS/ukFJIpy6su7O2A0SQSQxBGpX0n
p9vh5n6XHPkvYwcDp7r1Rs2DSfkKeW6BIpNpyQrBuAvOX/m2NXpXkwFvEQ06qFTD2iwfkMP7cgPK
wzbGa4vngLP1sRBUO5ZoNafBiv4nNofvSbOv22wDHZhWZcInyfc/IilBkuUADzELY5trOWUabgqG
IpY4XbIbDTQKwmwXZMkjdjkmOtsrSqCS1um+RodB6Gnz+Va1YWYQce3fbP2xE6uOpQv5ferTHR5T
RIJzcC4AjBmlli9eOdtPzbAXCgfsJcy7rMP/ExBqLG8KKcvQWQXuOpUBg+STQjToGzILPsQo7EK1
SXDJvIk8VcsytG63asPDqYROXXdwMo+T+DAW23sEWIiU1Yf6lu9eeOTrJcNJ4Yo+db9OL/5BM/yw
sqTVkIgN9TOSDYuv/DQ+E2V3zF8ZTWwmBNJxJx/f1YaYJNFJ8D4te97sx7RfOZ45E/p/CW/8DAPH
CDAQfS8pa2QwMNI4xJdWOhPvWmIHFpZspEvB07ggopiaNkaoJG3/xEp7UKBxzIrhxHzUXpIFb1zj
KEaBUMFWsnbzgo8u334R8r0q24UlqxkZ0Ljq7LTNkDpxwpwahMMx+YjAmgJm3PpfAlJ00xqfMKB9
hNOktnmuEcv2NuEgPgtoYzjXUHesvQ5D5Vlf5MF5TTV7YBvty84BDvNO+e1y31EIRCQ3sOvd3uW0
sDhlSD5kMYXAcwuNJ1EarH9r6/A8od2a0KDLT0Rp1Dj0g+XPizj46/N4amkzwuHkslD0TjLx9MQm
jEsiHLp3GI6AjrJkHv/2zIfnZmHEPLbaxctofRclHYbrq1xXhJf6LNOIalHZQkMWqW2O3g76FnO4
1qM7PI06lU9i0GiylCAuZvkHF9FJe1CcASh7G5ZfRvKKWoMRFIVF+eZtzpvH+kKYFlYnEJL/xqMl
IXprAvPpuP090ByP73fEmaYd84hxgvb3eWSvNyXHPtVoE6kXjYnnvtuWfj1gyY1hArCyRYCo+fZf
3uKXu2od88GsasYocDgbPhMqI3LRZJigHlAElzqKALwfl80+HM8cnOlFP+UJoQA7/9EMVe4B5fqE
Gq0hsrkW71vk/LDCiiY91FpD6Rqgl063GfsBOKllxDDKpIFogxl5C4KR/BWJy84lwZG/AgrFFuBH
KKPFuMXtcQZq7n95OK5GBBAxBbopykglqb2KwQal5KINmBI6H1YItO11eq4xc7YPg6mBZb0nisYq
wpyF4XOtQmdqmaPyxB0vmKOYZ5IN7zKGEuU6G6ZbMAZypQ0Ad7zqze07xzfw3Y2ZEe/03suyjOy1
5CvEbXEueJYQ5jB8F0ZJ9X7gaB5PbmYn/XsQX2dAc+M/auygqqCozKDems2HY+zKxzc8OjdN+pfd
9VrroD5L+xbSnvrox598mhG81ZW6IEwKXYQBMsGGWjAywtd/W/sreHDz6Ml+sW1f2hqvBBPiKEuU
JyNY6KnxNKoaq/L7yTKtHqqWHEc3UuD055f48A83vO/zQDhWub2PmUVd+zUCo0hYCj6kvsp9vIy4
kFpk366YApSUx0JCDBKoklbaIqSk0R6QN85rfw3mEglaDqCjtpeR4d2cgwa66IednRPxbv7AnZm0
bXkttJMh+emaJxqsQNp1FcfOIjjHrt8qQx6iB/aJW3/dUp4mL/8NXyIOiMYmNbd3cpKelPCvNKyi
/00r5yu5XPNHsLK7uDJnE5wo/5KkIY6ZBKhVsXAoFjjwB5cuxmpwmeXHDblTnY27TRc8VppMmgxN
Mi+zMT7pRCR5Ot2OtWTSpsSfwr2nau7d5/p/45DNuv4u6Oqzh/U5Vxy1CU6K7wmFQn1tm9eVSVee
VP4KFT5idCBlU8I4OYMpatYBBmTP7AWgAANRJBHrfPrOUXxEFqo1aqpnmhhEWRofCl0X5wy5GfO1
/7i5F+AllelY3qp/abWVutNc1luYhXNYY+n62Jhs+rsg/CuNOlgLYo9EdUZxturVfeyORkjqigR9
Z0zZi6GJAL62G8Aj8qUFaL1YnBHccojPdLcjsMPH/CIJHQrvlDHG4a0hp1fvDbrhynjLs0vYB4NL
78KvvfNxa/6rx9wSc9pDCrioWDe58jhti2Q9rKiXe4NUz/3ErFzB8m4WeKjzVru8Kkhbej1j+RCE
i84uB3Ogd3XG/+gzpRlF6LeR5+nJiXFK3EZFOi12oXwPxevo2n6CKbGnAdyJsQ+aaXwAV/p6osfM
annO7jwAx45wA4ahVhvJ60RJy+ytNXMHax1G5qDzyHD0yxQi7++ke3jSUzvqW2Uc7tHJm8/274YD
GIAogO1jt44mIKCrf3jIDX2o1KAaJzJNKnJfEVAo2QO1afuVoIIDPO56ESkeQ5uq7oDdp/cjPwOq
aQ0XZGnxv4cbS4X2+vVhLHlvvDLyOIeG7sMaV/x4UfIqOhDymLgpqJKrAdRKKd8M9rYB/L47tVGt
Ra5IRIo+9ODpBj/e5hH4M/Fl52rb0TSncbaqjEnGiYBb+dWep3p9z0wn63tApr5NDMeinCs+5XVI
OK+Dy17eCHW7rPMMVfmbN5MqWeeAbvVmnfJXi6QeYfg7tora7RrliK4hCE24rdjZ1ay/3+lYe43H
pRrmflRoP3fF1IEx9kCXqcJYbCdaEmazuIfyD7bfQ6d+6NxH/izyD2pE9LDI5DuB7HTG0x6twlHs
HddhCZWcvu+5/FlXyJ275cz5DTlaaY4tFpIrrKvYmqHkk2plgjkiVnBa5PtDULCS5GSyowbqRqVD
RzTNC9yVhlIs3nO+GUrItPEf5LJjz8IsQttYVTKhH2S04gdJGfBTmw27sOOcal4iyuafnVrn5kTo
cODkz2fEAOunIdcqj3V+4/KV469V8Pkq5mN8+QsELG716Ztf+y05cAh7jI2lWp2H7Y6LYRICfJQ+
XsS5lDxxoemnFu1dFqIAzUhTuPRKp3RcCdc3M/EfBou8CSu4n7TTPp8J87Mus3uJ6EJHgWOnthqV
NP93sXwWXuH6fOpBOK3GfdkaDyoG99mcwVB0ZP8BsB59i2OEfgYdOHFXJ2F/CNh6b8hzgelhLIXf
387emtFq/MHfjfMJIxOfMksKF/MGwzJ61LZRdQ43dDOyk5NVSrz9Q7me+Ry9mlmeFr3jHqt9ZNOr
nOH8uPke9wVBMogqaPnn2utg32w18i8yp1AXwsxbJHTC8j3kH4yDJbNg9Sy2bncBi5YiP7CA+iPB
mBI4QDN5gGqfHP2IwqY/L5LfnJPedlOurWnQd+Vt9sHBeyFUC3WAvekArBq0VudDKARIH/DfP1p4
S77/O2HC8oLqCO9k28UYiTUTpnIgL5/FqOES8AUJXQ1Dg7dRwTvK+eqlFrgPgk/tD0C/qX/lmmF2
Mn3BWtBSGA052oP/pUmtle0Rx5xFYQ56MjX3h479dpQCMdVHe7fGdO7SwRt2k3gSMYEedF+BSFsj
W+V6HZRcR42uaLPtPOb8lOv2ZGZXv2wjkMj3DpbrbNYo42WgOeCypI2H+996swN+MEsDOTNDSa3d
M8NGZ9mX9ruhEJYsSNcByyt14CvtxNPCFErWnOKfasmQgxYuyqP4rqwuge1HTenmq9IV0T1U5YG0
hDBs62XBWbJeA8rrDJwLJiixi7G55KF7DK3Pb+6i55PHc78b7DGn23Zw4T929TUPNpyZEDZ3qQUy
cA1vo+8AU+7EQpiop34LtfWzKDCGOSVoU44mCyiZOgHnfUvNflaulsQ/3E5LYUv9X3gIgzQxEvje
vEwjlfv1WflKgzk6wOkKIi2v0m9AJxiO3hqRzM62zxBPfLLI1t9mgTzolNkw76RXD4erPz2rZioo
XLZxcUKc0gjIuyOlICgJoA5HeO5spUaJro24HhFAoq1b9QNHUv+RFpnjxCIlQNVd7HY/mVmR7toF
7wd7bczSI+usZsp/7WrRuKrbVDj7hiQ3fJLp7HdcGjr+6HkKwd3HllevUn5lVHzrJnocLvjiNIlt
LeSHMHE1skSeVIxOQTmXOZHOwicqNiacWZ74QpMT1zRIfui/KPiqBn00+vHKeQ+4eE9thLOu03dr
4dhL0J0wIFdKju+QCJpk5fTzn/C1w9rLFUQBSFGDBAk9Ag+pJ4sB9S6fg3juuR70z7LHpNSL3OC4
Td/mEBcOI9DAcPMTOggNyuZeXnxdcQO6iNTd4VFTYn0u6QAeaOhrQAfDDCUIcGW3YNt1T03zxcss
gupoYJxuMqBamb0hkCDxSpjcBA1qzA+9MKJgn6MCsO2JtEJhoXfsOlwyCqBPvvCm80MUKnaOWH+N
OO89otGdEP3XNAImqD2q+aiCbmSd00joYBG9WLDE1S7kS1pj/RHUKyhEFvClsOePfCFd5v4tjxrA
jdjgWAf7Z4dzflDDYntWipD9tTNwc7HLIZ0TopN5lDB0mk+28qoeInnN34hUEDyRQ/FQewAglEI0
Rr9uSB1F6+XzMiTBBTK3nifTOVK7OBDrOafcMFmdE/3vPZH1nT3IGzPfbFbvEJsM6l0VX9qhF11Z
y1Hci1nEJFbW3xP8Jp342FQGTwdE8YlNCp3mqu8X3Hk2x0n4WmU2eX1prHkTX691kF4xOEFl8Nhm
7JSt4py/2N+O/s95030qBncuJFVLMmolxl+radO1oPnjz1muK5pFRQlbKJgY4rFlSBSSX6OZbZhi
eKOA3mrX9wy/9Z0eEsMkv/O67JI71hxLoeEhtBVfq+sj683suf+gCkl4ZivsjRbn58smxQd1XGCr
5e83cK9GCf7RR3VlNKm1V3Rk9gRMvqeheaSjIOkRelEmtEDfpw5Kxk5iaTqBpgcCGb4ZRXLCuJfi
EWXBKT6GX0rYilJXBV4+uBLqVF9R3oBRAqxG2dCmywNgtHvBNJvjeyioyNYyT8f3XkZbBnoA0sc7
1nrs4U/DQfkkmYLSbjD61cyEnUbCPpo0Dm+suok2V+AP5VYP4fC69HeyGCYQ+wfYmiN/lQnG68gk
JnwMnX85o0HiIE3XsDGWFgvMB6VRtcrGvI6OSbWg/fa1mbdgjVIi2QzaS9tgqHKMvKMYLKv9MsbQ
PFwgknpIygZGNX2qIQN4VcIQAgYbQ9B6oX1fLHH0KGVNDPG3Jb7f8m53gwElYslNn/7huUO4IvFL
s/SuLxq5sdcwpdXWooo7zytbKIY1R0HgzQgFEkcJpwIQxhEn0MqnGBnv8B5eeNQxDHvBKqoiK9CN
weIriWIRF6+/qFnbE6z5Z7Ncma0lmQh+avz7vkcKXrthVYZz87gyn6EP8SYFBd4NDU10vagDF4qc
pDCaGiBVeulVdauFBNJ7WFrCsW9BkKl2gl/KSlX3rVqGA5yhWVqriHH60PgrXNxJRV8r1Dk3mR4Q
qEGF/1ofYcf8FjPvlLpqLSB5H1e6kEsPs0cvZ0QkZ3QPdTANgKJVLCd4K3dm2mMqljTmA7VtdhPc
qYDkJIYBAzgAc1n3KEjYu5xlrROgSOIdKr5QF5vGcLK0ZJslvOmUxq/lFl/HkCU3KyGryikJyv/3
mQWpJFXkD6ftpzSHq8hfPudMb551LkGHNFj8BnR6EU/Corf8iYkrn4clhXCO6cVteVmSRmY7/WfL
vCHKSORDJOFRgKXqXWvFtsRO7dx9RRqfBMbJsinfyfrbVOIRAphwsqVLZNRGnSAggXMi/ZRiO+lp
suetJWCrhPb+PwABTTPusmxzbyYq736lEG8kxPAWWSa+ihSI+8Omfp4li9xItrtb6AyACPJDPrMg
DT5AFWjwW66YfxZm4eVkBTR22OhA1cnrNYbeWWLF7gPSZj7YS18q5I+wpctdijjmLbj/R3PvwXuN
6aBPyA8ORRIhYEYrdkK7vfV1S03XOsv1fdS2n2nyfa71jUE2t7AgSsOarTHGtltQl4ZjPun7lKez
b2HhVJvS4G33umv29VWGqNj3xg76csUd7YAUTIaksNWwhbpawP4OYYGgPHIeT3OU2C9snYOP1cKC
KPRK+NU1Ca3rFdVd2pAmy/GG6D3V02mCPcQlxl4vG3tI+yH9NWmoZnytgU4XZAmKNG9twvnYGRhl
Iq79nJNqMJaT0NunMUz9+5waLY2yS2k2qFD5smf7yhP8ex50BDC+f5tg0xbOnQ2hlbPsd6M06Obt
sLbznOuoeElXTvrNgbkV0sfBtAsB90oLlKUf5Cn8fgkn6dEu8xwnq2fsMI4Bg9UzhKqdrGoLrPOS
vVeNESaf7FZnjKQrxcdAmbJkb18wmGzcwe8vSfWiCy8ZvFnCX+qpw4nzKOjBTaiwxftg2/KeZfqH
izz34FkOmH93j34o9+zXZbkcrgSPn2JoVduetaIDDgE1Euz4r5A7NCAk0P/DG4Zkf5yC+wPVWIlU
sRIBVVPUhjWniPDiV2hwXrcThCkyvIP09+QPEOXNYPJwDbNNeebv3/CrkkAkbnfytPN9/pLaiwWk
pjkLLoH6eM06P8LqRANu8x3v0KbXiPxm6LggchnJ/zRB1A/OnwxNsP8H5rKJz5WLC5gt0wYxpBJK
qlOZmxFqXDJ30vkFVv8g6LYoPCmtDS9A5qKfNUTlF7Lf4nzIVvZh8RvMjJTJy3tTCnqCjK7Aqym8
BtHg1++GSAoIjngOeyJPxlVaaQoEkNWAQjoi/lSpSyU2PMrcWqLAxAo7dRVuU23QbZac2Rmir6o/
TuICoeB42FCP2kpi/lkaC08HTDStWQGXo8iHyAm52P34ZmYcE0IwQ0N7EUdgRRTmuHGbuAa5gElI
UKXexo1Opj4WSLnb78l6FHcfK0dUQVRt53rEiH1qT4veQ/pqHDhfEeBPvrzRSxaE2UtKlaFYCVQe
nSdP3XwVc0As/xzJbrAoy7nNk9roq3Xy7BK9fs8tsmXyxhyuQSbHI/MF88ZX0vdfHDT2ZH78G3eA
hZliy1yBbQMrcz9SrjCXih+TdEWnnftHAHM7SXuIV32ss1yRFJzjmEEvy+5DroY1Vs8tjaELgQ5f
jczzmWEAcwU6H6GOnAUA6fH8FikTbNP9j8N0Nstt2nywtvON9qax3BOLvOCHvPME3vMV8JV0kq4N
gqgv9ibrXbwNQh/lJWInRIsLwrobF9rIwFTlG1euwr0SCz97eL7aZLrg8Ooh5ktNByFZwx3P1Hgh
8S5ljf9xUZqiyDCSYOcBCnMh9sKnMA4gvwquHpMqc2G31BzQz1KfpxoiVtnhB1FRWzwDCVuTMzlE
roES06YlUOrxnUdb/gS/YUXdr8AExCCNLhJigYjfBVJ12BwWP1spsaRSjV3GsHlCCLQZBnGQzfBC
tHCnLifnZAplENH9wFUz4iUxR4IX498ezOK60E07ssgSnw9wyhf0D3oSGbPJMyVcNKSVjd8MhNGt
YJF0UdXcIj4e8xFfKVlenYXCtI2FxTAw6LwnPRzd+BLI6YgQssA+GqwRcXuyvSL0qzb0VEv/FLGF
mlfN6Tf07Ur1OefvICWYuoNMd6AWAy2x7XVQI/JGS93jrQZPlF0TCdonDCEeKXLeUUfkrA+fIxtP
8358lQq788Domx8ZJFxFr+Eq9vMA96q5eWceAnMyAb5d8AUogG7H6Sx3IpAHHyN6K/ADyAsLq2SF
Zs1nvhej4isvH5vvaGhOgP9qIacQ7CRSXMKJG1cS9zT8q6AGTBu+AEf8NZMQE9BsWFkm3pN8hFix
3hRJ/BiXPGHvSq5J/puHI0ACit6MzQA+brGQZbZ6JqMsWbH3JMPZYTnsvZtV2zHpmHS4mI5oElwe
zPXuHbaW1zf3zzZSO0kOuiWOEIkT13dOe+EyvXlaE5ctCN5zHN3UHsKE8FANgiGy1hQJmKCqd9In
MaDX1O2+bVVkAeBB0tWDKLHii6d3IWAcDQvRcfChYf4UdIX0jB9ENMxvtUvOfKzI2vfM5TGAbekI
umj2tTgV1skSy1zOW5RyTkF5LbRVZLXaLkmY6lX6DmNVytUsOxcc9OKdKHFArJ5JyZkt2HoKDP4r
cNUXP72f94TKlXznP1zCcioyzRthRUP1lhv9tvOBC69bza3XFws9gnrcYCBQCtOsCmNBINURR4aW
qH212P9SzWI1YzOHkOJVi8s8hY4CdHCy5vOHY3JGuhm/TrkwD5t0TNFf++cbg4qDCd/1xRFHL8fJ
KGeGK4K7YFZqY49z5psxu8q9JquHYG59XeWc9XAnF+IFlYV4c80nmMW7YFA08YuMQ11dv4K8ayzC
0wxWC3EWjuVHra/7mlOuDe+qPiBt3OekOETDi/gOFISQUlPbRb1NzW7RR2MjKrObYm7sGFtPCCGy
l5JNc37bu5qJBknq1rPnGk2Ucn89WmErYjvLBpTftxSR+T7tRwJ8NATvnV89MYkEAUUj0EvSnAYI
9HOgOJh1MHlgVm73MWl/JS+I91BIU3nz7A2pP6a1r3RD/EVg4EQgoUB636cc7R4lMgtzEerZR+OY
4wcHpg0XrhPdgCVeZfKie6jxeUmXQ6cawckXnQ21CBUrLGqsd6cv0yYlL1yfYi0+Oy2uB6maOdQo
mBxHEbSQJuBjeTo40IfDwDNbCrqx9z7oicJFMywBDKnSZzNGJuY5v7hNka5Qn8nFJobdzzCgjIC1
grVCMHB312dsMKhArLt6rQmkQx1+l0Rhmc9IcbAqC/Bwvfxn3JzAahH7BBKrjsDXyS0UruAeLdrp
jRIKxhoZeDOuEY2Lm7IACZPUmNHBTeTFpPPOwuT+BhZI68vhs3XE37rCHA47lsQ2kaHkU+wPv6Uk
CtDSCC+ClU8K4Kd7fluG8YTjZCn24UGsNCGZOefiNUQO2BHSxHijq/Jw2cGgfBasYbI2TmpDMl2o
DGQAgKpqHAyzR7WVGLGFOOuUsNPbGve2X/SlHA8mSum4ExbwQ0Vw7R4X+xSfFNoDD6Qnrv7kQxZ9
tBoUsF9CdBdwEsN5aPnJe9c2+XAUVLtD39Q2+uXZtuhR0nSZZhlyZWPyy/O3YA4U+CRYnYCsaGxS
Oa0VHZLChUe4LivrvUcWg+ZQdz93wCziB4fDrSwDWMzzavtvQPV9PtLjj+7PtyvIguwxUHguoIdW
QcyfZFWz17D/eG7VWbh93FqWZlzY2fNAcd95fcRZmPx+jFxfMZONr812CpF8YH01C7rKwjQeOizO
LI/stf+mYJPTHwAFTRVyxxDsubZ4CcVLposeCuOilwtqm84NuKtpxCJfUJzDFhQiplRU2qW0dIS8
2dqtfJZOPr2i1CZlb7n/nw1SoZS4BLT8S4Ithcsqc/2+R5cb7svkfK4dgUaWlrNehrR3tSwVxMb8
lYKa7dxtqsaqCHYjo76/y3Rt0NbTvxvkIm7Yzv6XsgWaQBhObcwDOGwh+TTKa9d0kR31jW7ug8z9
756zs3p5A9rfwy9G5thdNyFjPB4lvPJoa9pihW4L6xk13UfM7+Y1RUx6CtApRiTdtYJ6qUtE850O
UwE3yxTgXx5A6trPYUdWAf/OuHfDrVPy+cDV6WCiA1OkHX/0GKiqe7YxeJQd+qfk72hkWHaEyVP8
tFV1KcE4h4nuRrUxtKVVgpqcC4JXiKzS/rzpMd2mueP5NE5fEHo4I7Wrr5Rz9E0V+rJgrm7HcJEP
+5xRcN9Zf8I0GNNnWYxpvzUZ8qQKfhmmiiVevIfmtIfGJYrMNt7A1XHTy8E1SdF/bC08N6HGJzAe
UQXHLhqC/XUedAfS434MBxuX0SOTHh/JZilT6edmUQet+m59b3iJMQiLEIEMvu6RrlPBDCGSZAU8
jB1AfHPEcpVwfJ2py9UtsNEnabIeqiZHm11eGpUOSoGvIDpcnHfl4kVKmBBpVYWHJWFkTYZSgMQi
VxpAx2okxvKi3VEQjlMA1RNxyRb20Cxl08K/1q+CTDYhVYEHAiwzPXtZE27Tq83DWkDpwYncl1rU
QeP/BLP+4IIztOORHOoqfe+caX+iDd0o7tIZwHiDYUdZkdKOl4+W2Xbt2bBtRyRV11WDmefN8FXk
7IOSwI3nUZ6ffwyGsFJACkSBzzk34sNWSzF6skqX9yqgZ1KpBoqIUDZWfcHzBEStdX+4+QSUYMnO
ptKcxp19WM5Jtpi/Mh6u5L3bJggCPA84ylYSUYd9QCxOpR+GS3JY3CJxOuE8Pe/R9B2gdqYTqGmG
eJ+xUbepGPWUNoGCAC8U7hvhbb9rMPrAm8TSDtKgzlGncu1OkJOWZdVymPxDfB5l6HQm4yfG19Zz
u6HuYgLkjtCUuSo7875W6M+v7Mkji+smJv5VmPUPbE1tRThfl9kwZkA2h8v8KrjdOSUZYt82o2hJ
hTtl7UnRcx4gXHp0DnUcG3Rreqz5mq1+PdX4hOe4V7bNBfBYZZkMOsX53hm+cY5nbVAdr8qvXMDW
VOcASSyP7Ii8LMCL3tKdt9AGH6sJSkIdczgpFBihNrdd5nUKGBZt+s8Mju0hTkKDjy+jfQFsLt67
5Tea7fRnvf+7l04ZNfFzkmwrkZRQ7xSzeQgKJYsZAAQV6mzS7UsrMEspD8iKdpGkqu7uJW3krCho
WF300msoISUkvzqSVE/8o7CgZNpDJp82KPpnTRHezPij9IpVlptLJLb3gKo1qJ7/HwsOG1c/lvcb
U1Amf6O46vrbunIxoR3z+gpLNZjm7dMawv4+G4T1WTHq7ASzuudWGIJNsWye43JCuQ5xXmpafAtg
DWVB9Bsas3RoBoOWwDWU1nsKCc+IoIEfVuhygzFM0pqFPNpwBMQa4MvnN+V4G/AqBC0t4FrBAJno
3CcxmnbjrGXgdoXYHER1H5+aVZb/9hDbWxy35QOjznxDawGUE0tq1OyBRixT57/3kErqj9aNBEUK
ed2gOaLruqSj8+8aR+YKFFoicxrGQF5AH2oOOuOu7ePAVWasy/vMU1fec9u5hVzoOoCKEAJ4LECp
euTB9v7OzQpkgFahOE8eSZ1w6KhD4c0AZNDjbUO9ZynWgN7nvipyB2hYoxlxPKhennMF2vSv2ZlK
LseutS0qr+0+CDctbiq823BhbulkN9Bi17um4YP1DoOUZWv5z2T0t1QUxUtcW472lEYpr26pe+zC
sjCaoSLTFOgXv04sPcKbks+mi288PU1NZZj8P+49aI3PzJ/e5o++U8NPM1vaJisoYF3bZOdnYi/8
88fOzRaT67tPVBP5enlJ3YDVOD4GEEkShFFKq2yztA2yIVxtTrPt1JdCU+zkMZnFYT7ZGtvdnvqP
z+TH6qcptxEtoQGLxVKMxLMR+2t3t8fIJF08TE8j10bOGtHWd4LlNbtWcKSHNiktAZjCfm3Ko9lg
GZ9oZyzsS5CtS81caSSIP5AI4EkxzOvSICyGi27nsevhlSuevcpZz/X12/EiJJdLsnMpnK0/IWWr
9l3XKFFt5K/yPd13VfkSeNxlj7XL23PXhx75/rHDGwN4tHNQvPomBtNUxlGNbi6SrUl1tw2e85rD
mHizOdgZL1AEckSjR1KuzuUgLLVKiGkRA1XJeWzHDcqwo6QJ1JGFiOO7ZJQqz7Nd5u6UcqrLF1YJ
Ji9088h2NZx1ksXTsOj6JoaiC6s2fYNSojvsAEHP1O8hoVsD4m+83csefD8UnFxxcCXkMHSDL7Jz
lc8AyfZAwGFXb+golrn85Dd0CBotj4+r4KvOsJx8yeGPZlmUOyVFk8T6YK3NPu7FQMJaZIzwuRX2
WDIofO++gVgsB4w0YXCTL72QY34MChcpNX3gth2GEs2Pp7n5KG2MSputNW61NIr1u9c/LUKJYihB
nu9oy8mjUyo42pgekht6WzW0p1razy5KppFBqtz+aSRFlnACKbIjRngr7o61G7e1KAhAtadrPi9v
VB0O1EhOS5tvm6Wq/74wPvdFYSWc0DFDsYUQeQYZPy6XRC77Feb42JJW26bQhKqhuS+UCIHGj/PX
CRwBriojokBO8zQcy7yo+t4NBiRWtV9JlWykstXtRIyozzsV8o81DbGKvmAM6PJKIL7LKSrJ29Wn
6QHCxDDc2jmZ5xrv7nKuuqreIf5gVr8CuDI/1PuisrAhg2P1WgLP79kTXactduZ723DFPZSu0X79
WUkZTCbdhZPlyjrsgfpDh1JK3lFo+ow1vNn/ZEToOAJOvXMOWY2JFsjrLv1ouonVTu0XcoUVtZWY
AZR5kP5VvfOKLHfLG9lRrFm8/ssaCdX3H9Ux2cAgDu3wAhCJBrJAHWPY62E4yfqk3D3OiqF1+iXS
JMJ5GOGpYoKbhscBfcoPMSvbrG447wU7RlG6GPp1K4YhUHHCwWMdRyYTXu+vCaeGBoBQQRmqqz4Y
PUkpBzhYYJS0kR9xOf6QT8J3HIWxF/Lmcmxk1WDuZEWV6JtO3g4CXTWCfJtLziYpUJEwzw768kvJ
pHCH0A0VYeT1WB8EhDTj0lUnnu4Xe1yiZvXBW04VFVu4TR5rry/OsKQp6PcWE0RDo51LCVF9TQpg
+tX7nqTLTbj6sMq5PjEBJdxqam16bUiwSYbMidNnhOhiIXVlhtclaP1FFAliFIdt+aJl0O98DInj
Q3KPWRTWqQyF15HzX9qPlmCj+d7HaUWIAZOR9nSfBJ6Rvxz1qeL/wnCX6Y37ZI5YfgiOL6XuyViJ
W8eZq83p3n56/HWQrDDGKE+DtTNu20ubiwtPFNit22gxJegGCpp7kE1AsnxQtVYHxK405Hlzj3PH
mUCgOciNxkUg2Rtknjue7plrlaoS53xdJxbIWxsMT2WRi3spR7odISdAg1oq0g57tbVb6w9TXNGO
jX3wp+F/eKpyV/rBy99ECZvjfrW5auZMX2Lu8kAimUyvv8mH5+HSwA7HE/IulotqTubIkhh3ukFu
bhi+dpcSgxzUmo/qI4kmP9r1PjvuccmchOYmA97YRR6+1qH5JXSmNQzH7N/kfSUMyyzghfSbjelc
+O/gW+0ZYLUi5ndCDv/tuGHMHKaRc7kQDVDuqgtWNRr7+88t8uU2vDrFVgUbrUNiaTrgmg4bYqpR
ZWuKWpbMIowMzScUnIfDmIcTKsVHxyDgR72lFrZJMHdoob2tAV9NJ0GcSGM2JzXf+oez3KyAhv19
Bgs0e4b0++W7cuLHQAlC3gmWNaF9KavkD2RJbffqqzXDrGwUHqrQn2dVifa6h1Y7GzPQcT3UjWm9
s8zTCWoveXSecigLTDiD8osiQJ5XTAGBD7mStiQPkmcojxd1mkntmRZNTDu91EXaz6ol5GBC6Ofh
hld0cHPKPdSaT7E3PHfKZbPJfeR3aoxy6L0GQ99gDcijk0lnGoMF8G5NMoyPDnt9sagjMFPiFHUw
eNqRVZeQ/s0znZV649mVTERfx29uB72NVA/35b3oJkwGhcODd9p0gbwy9atneYEP3nP2KQWumGeT
DBhVo4lHxYCqEttQziIcXmI6D6WvCdK/TokClfDPu1RKOEyw1QVovc3a9UM9GuH4dutzGQAzuIqW
1417mbcAyxAdab2VCi/ByL0J0cJ2/5NrcKDMs4nBD4uf0bDDUwfVL7Bt55fkHrKtP3tzj9kwOf96
djMhz+SOB7Y+D6jHa4Iv4hg1B6gFVsr+JQ3VJTdmM1LEKGeS3EOYdCIgTB2D1XTv1PjOwxajNasG
dhHyyhisIrvoT9bLFQ5w8/v6IeMe+vrKnkdT+M2H+FfzSEZkqaMJfHSiLNby6kbNj31qUcSUlLGO
rqPQN++q7Fc+VzW6JV6vBKWMBUXg/V3q0ULY+4Y4tDcvr8BjTJxN8nayWUke6kXh6Hp36EHJ7CRE
zs7vtvaqHP9fG9e0VXQI2Lg5xtx8KPpSQaPzw9Kj69f+5KXVdykiyGtkVao7inkSxkqxpwMO//rC
YBa2hF0TcH//8OM0BTZfTf109gMIdjbkryXxztBYvJL+ohtfTV6SvBeioXRE8ObckawGO+oH2Pj8
f5Rju3uknpjtlawvOIdbswxi0ppcR2YNCDBWrrj99WR+Kr7spf3D4SKu1dXxR5qPMhVBmnfBF0MT
cDhcv9+6XKKLazxTI4sUXUD9LQGiOdjYtvdvxqmr/NPGo0vVFrAe3K+SR0TmvhC+KTDoyCYAYhGI
DH+v+aXPyUSxh5cWRcPcq+xpQcYzZjyKBFEOY51o5C4DA9PvQaQJbN8opo/sJj0TmQWssYA3oNzZ
zN3B19KT0LJJ0USlaCqdcWN1eULRtL6JNtoY48md/yiaIZILuTqSd6/D6R+D6Hk3w6O6n9SuT7cr
ZrFYKKJqjpIJasZo3ZTlRt3o/gXLCp/B+GyPG3rvuS+TNhXXsDgWGBqXLXbVAcnEZxibWNg4Hgkx
7hY6qYAhOr9/p8g+BANWq0qmFQJqj/5jBExHgt3tW/4dGcJDjvpgTzrfgjtDraJr1iGRIWg7510v
xBwymjGlr9slvJYPgBum6GyxCTZvAh3PcUPTonujnfcAt7RZvyIB8Z4uRMlnkPjadycu8qtGch7l
aMKDLi8uNJw0H5teaFKC+oK78tXeaEVmUtG+GqVg3l2vH030E9jcSM8f2xOKKkX4yCoiliJpIjio
z2HtfCKzKR0+LeJ2aPO7wq+ZbyxJGSeWSe4TXSq8xTiimZYA4SYpgftOQShFMWTV6VuVCxo4Pvn4
BTioX13nLZNA1Amh2+NVJ7VJIf7HwxLyWZ6mmo6UsebFXUfvPUOxQBB8VsdsxZAf0TZNQPuxG0sq
DHeeHd4TOJhJtUbPsJ2gzLa/bwFDKOit2zC6x2sdwq65qXvzlYCjP/4A1YBQlF0HtI7XJGL6h89C
Rh1kAB9Kd07o64wXIPbnYVAaoHyBTjFEGWGKXPCjtDkl8OoclsvxmEWmvcMzXS8Rejfz/q0KJxt8
SkIthUTYOeykq/ND1Nk08CP1sx7GMJzMc4l+v59CikYE2zI2H3YCHpM/WzanPfLrOHMVn+IyW6OV
9PITwaTPG+8nikOnHzrsnznGU1m8jkbRG4Q2a9I1C1EVpH3bLR+H9JaMgiJO3CcnFR8ZMPNdfKJT
xVTPD4NgdJhSlunx4CpmqedbQUfsksU/9DWrUT5DUn6ax22pqPJj/1TX10VF7kM/rLXhRhByRHxV
32Cf9VMS/V2RuNKP3Z4o4ZHciD+z77lMemXwI4dvUFscvWwU233VePdl3zwa3+t0YHuibDyKFdmY
K9cgHkXfE5cfIwdhHBmRtvmHT19Hj+xlrMrhXNieO2usKxJ5tzSlBGIaTNlSC0qqBUAHbLaHccGf
TwGKn1bfdeG/KEI5rfimdOOJ/Cst/Euk0H1q1y8zcKmQKEoBxDbZaIxlOGWnUMwOpt+gI3BORWyf
Q+TIP3/LfuxnlL59lbnxoG4S0q+kSexh+ZiGCVFUSrNLcxvYOgJxEt66crbzZXqSsg82k7Uqnn0X
zHyUPRjabKe6D5IJBDUfdgIoRknyBMT/wXq7s5ULhtiQ4L+FOceW/uoEdqFroKSGcFUsNOdqb8cb
FUlOi0E97o0/SIk6VurVoZTmWv8dbuu4Ft9S968pg1X0vvuFsyhu2edtUNRLcOL1fRFzATGc5waF
del9DygGKWCcIx79IbeLgJbyM0huQLV/hQGFeOaA5aQMNtx3SIRq0kagjZf0f/2lGdcON3oWZPNh
nEwhmJR6Wg9dB6ZVfL4JuYzjkpkRZMDeT4pyAe5N1e+NXs61pcPDUynQozYxJPvfOHGQ5G/ZBBj3
DNYg7kfW1pEWIcYa+UyYh0+G9ZkdYBz74FeKcW7+S8au12H/ckybKygo5V2IdZ9PuKIMDQXDsB9G
GMC+5tVxOrOZl3LDWCUaUj3dXUrgIXhY3gTeI4Jfo2fsUc9SrCTU0F0t1I6WP8FpQD1GwfIlO5B5
k3ydEWKZEToU7KLDopW37phNOrl0DRWzRS9jKXSOHD8ACGixpauqCZh3Mi3eUuUYV3XhctQsKpRE
rLnQKob6JTkzDQGWR/wJY5SwefQrPFVizIk1Ohg3VOCTzQ6kw+d9VA3ktOvqgV+3Y/G1ZrHN3dLi
Zya0l25EeRdITK52g2XJgWMcQHs1T4VLRWzzVQvwNrk6x0ZYaOTgaLTv2Nfo90Op3n7oaf3+tVgm
t4yPvFeLEdB47a4ttNT2HCj+AYSrYRImn2iXqxQZXiVVu4qldXpU47oIvJyxTOAqmO0h0vi7QhtG
Tfp32+hUmbFh6wT19+EyOVVxsEGSS72KQK2tFbLyxEVkmv8FBL+sGEhjqqVoYFhR+FipVK7v6X9P
VNGINKnrQxRPf/fWYFDZFy84mlulAO5bld3XlFrW3aqTzWEYB5OKC/WN3MgSTk8hKi4n852CXlJs
KbvQ86UJuxdepiV5vU/zLDZ+rwdMjfYWl0/mgnJMYvgbTZn3USQibrnizrYlAA/HJy6yF0TafNas
ncttETV0O6BvWtpmDGmSGh48RBg3mRc0WVk1HLw+5oxO88XF21HHo4JsutHxFA5gua8/eR5liUO3
vuGpNCY1u6JP211ktMjKfSsyzZiwXAMLX0357d/CjwOtuSPde+xsuWK7i2VUhmZf9Q6s1xa7gj0T
pqXmUBwtAgKKLhHM8ltnAqJw/NMMkTJaK24ER8SypzbigH+a42l0dcHom0lwCcyz1NYKmOteEvOW
iuczjIBxwTcygXOSOmsYa1GhynHgrONFGAy2uwLIgv2tVZaid8GE2tsL0+Jw+TpdOWI17Xuaux65
BZxbPHFWpodPIOu0G9LYhY+8XEHHlxN16qXmKPaC8ZRfXCNJ0J97i/Pz/cCDhKmPOnzFZ7iObUY+
nn4bQjUR+lq/c6y2r/7FzIzO41wuZ9i1rEzgV5dHY9cdrAUf69JaecndOy7xuuT76gNtXtS6N/OZ
fd7bq4ixQsv9VHchlVphcj5t4D37G3MfHa7AdbF+O9tgQ9qxhAzRwfXTIER9KDytNlAqdshonsJQ
hf2clxI4ubl335AI3DEru6pr89oTQrz8K6X9wPsNTjY8n89tH3pxkeibbHYDaZAtPQGp6q1vF44y
Nhn9IhkWaZ6/NRNEioPF7qbJrilCXplIt6pIyXgu6ezc5jJ4Pl+dfgBK0ArHCN04AAgdIo/FO4wA
DOTa2MdJQcibks/aBhXlfz/n8Ihxo02wQ+tZ3nSyAlMR4xcMDj7qGASP3XPO4e34U5hMuEaqJVR7
cgL1VLqgnSIAYE//hsB4pDo2Y7h9q3zB+N2sk5GIAzsslSbWhboSOrRF2FFJ2HhBe/Hw09xVrrfD
ErfVdrvKXs1WPmvlWUTDdhqAAKywDNbhkEzPzK7FfLL7XkjeH+z6Bp+vOi7S5lt8w1a0rAdbuW7u
rPEocUZLR6MDPSV9fAI55f7iJ+cyoTB04AZwYj3z1POFEVa3mHPSO1IdU7U/886SMYyiRadQBbz2
qeqjn5VQj7tkVuPDsRVWGs8Gr7drtHkdwJC/tiTZqQUchoGJGN9sRMRzlnvRYqHlGjorXRqAz+LY
CJnkJeUt7GLsBCUALjW3ZWfcFMbXRZLAM2bD2TnHaDPtPfBKbiNtKBIoy6cOVBMRaboS/SE7XOb0
+7P2ZJtalTJpApx3HRtXFpYZXxB5EJh4GoyiEMHONmMPpmhE0tRtbetPUbptpHK1sxpN6F0qSON7
ppFczjqZP69zXFY4w57Y2ZUH4Y4fzJrjfTYdgR8gFV6ozpNTVEelvM6D4DNjshIBXMgeHvhtJw9u
Euu8eHUQw7lrYAQAglGLVxUYuYlv2Mz2EKwMJhwEw+aaPFFiXbXjIgmWPIjw0XBl4jchLEIbwjq8
xvgByNJZwxpDg3n+GKFzOJfC0ZLZ1MIvcebnTau+6YvnpAPzI1MBsfJtcZ9j4kUchVW5e8r5PXta
vaXYJVulygbaFUM3JP2RnD8ssyfaoNs813tOEhBRxU1TcTJIXCr2ZnTjwRtjC3dL336jNH44aTGf
zfS6b1fEEZxMLpW5I8yTfe3bNiiHlvchAURSnB5VrI2rSYyLDdMxH71NyPVCPliUxUK+g48xfUO5
kZWF5dFHnNKNR1h+/Q09KF09tUKoXZb4g5kiiLNQcjEmjrdkwSbCYuJk5uCsyZKd5DOhtuZ3DQRo
C/EE6rX23F9ILFkZi/YzkezKlxpQ8qJhtldQcIiqL7MBgkg7/i1rTSGTlG1YwQac8DHm0rznqSeg
AuLx0JO8nv3h8wgSsVPqLkd7Mj0htk4hLKh8ksRJshU0ogOp0amvtscFg3sZOUUc8UsULTZkFafc
oXqzKXnzgM7qvyWVKqSoXALOz6H7gN1Cb8e1PI3+eVpAWTlVh7114mJTVClUplu7k4oynb0dbLeP
0px6JFkX4X0ktZHWJjedDzFXUReh9v7PXjI7VMc5lelwlpxf69yZa8T6iaGxoZL7GZJpAci+lYD9
o8tjvz4QNsTfY6nyHrPboZFyKBnzCWr/Ohpr17w+h5rm6uQIJAEO7cLq05oZuq1UNi5IVLFGmpx5
BcvZWvsR62QvI4OVniLQW+51BhIvIH7wM8DI5T5dCqZQdoE+ulMtCdghE6JmaFO426SP/wzjk9Qt
ELo4/OQ6UQU/k2/jVE2vST6P8eRRaUX0PyteuEP7NYvzbx/1h0jnQpsdVDV7plOUYc2gwbVeA7Rj
xUj4eWnJDfStNHtlehvSptkfzC7+ArVP1OsfbpBWRdALDeZR3nvO0PsnCKLKww/7KhQ1vWQY7bWY
8E1ksLAwg96FM9//AGrZKUp/xGLCVcyxL35Vnetg50M/bfQpmv5DviW7H6Vt/ZLztPB19zod+R1Z
ObL9h2Q5+MW2XbYXNX4eKJU0Yb30CgcorEwDhk5KYbHpQTcJf6Gx2JQMqeA882HNvdRJCq4aUjsF
Np7zEM5Q5849hTV34cUYbUQ931baIbtQojmEolaHnqywgaAXJcV95Yr1Guv+PlwggzYxZwcZVFxq
uyPm2hnARX7iPZi9H1Ezu4kA4r4opjrv7Wet67lNlRhB1DAQqZ+A2RlNAWhinBomNoEfVOyETyVZ
/ynXf/UI2Pg7LD9mN4czBEMyZ4hgkQgT2hNbrn5iM4EzaP8FvYFFhpTvAPlbe8mu5+PpiI5bQHxb
mQPiPBGmZ/eik85QZE8Z5dgkIpQGoiZCMth7rmNpNISfNV5GZVNlVrkA/8OlO5D8ThI80ho67gin
hPoc4IElHfb1QDvS4aPTQZ3bGuqFx+wp/Hh592hJIOgsgHgF0SIM1qgH/l6Y+QGYPwLby/L05jbW
IoAXcCc5wztDQrFxam2y6zCHmMGjo+igOdR+QyUXnq9x7OtV/A/8ql+OS7Cb66JXAHiXKUfMS1nX
MeuTKp55U9ne8x/7lDX9spAToASecCGeabTOneMDd8zDDvnQXoArgFjoTeZeVz6yJNqlJKH1psHI
rUqz42afHT+6XoBlZV3maGS48oNVH+u1uZHrCJQt00Q0Sluq5dChdXr53TXZpnuDi1JpXZsr6vLA
lA5NDxg8IYgjmrI37ZVhp14kiQDQ8BCq1MzARAag4Jod8w4fdykkgilcn1wveAnSBJV5uVOJ/CT0
jfqq3s03qjBwj4+L8tYLVoe0FdaJFc9m41ZlCO2w9CVG82wQvB/jRTxeKLIpvWGnf+jOEX1drAOq
dZXPG82iB5tr6famZBRO4dNfyQCxK/Qn4cOL4hUJhS7l+0Zpt7PyMqcWPUdt3MpzC1jOziupck7I
wh9uA6zSlnOr+4AOmeeg3FTO1+3PTgPiCgLhem9LuCLckXUTiTSYUlI9GwNt8jxolRjchOOTAPRx
AERlu9mp3nY4T7NooBFcwZKA0I9EexrsyvdpzVqNu+nTZvjQUggxxyYfOynoowkUHD6AebcGQqpl
/nbXcjigluRqdHXUG5Jge6gYcj615ThdIyJUic3OENnMZgJv8GWtnQdQRNaFhfSq4hyGfBoV63zw
Cfb1Wysc+gnZIBJVMdPpKK234ovwD1wTM6yBiaMyAbqN8/gx3HMMiMwTG6qxTKrpSJNNpiTjPPKR
GzLwd+VEMNjxr7H8jymqmu4M/c1jSnNS/i3Fhh70gLO83LLT+YC1vKKWeQQ+YO3zK3EZfRu0XgCL
BvNSpBXyYYZMM08vZ9SYc8GwUo6SMRJdIPw07PHyHDOCs5urE/V+ferNKXj1x5SWEiENsS654Zsy
tHUpZ1QowwQhBJQLWuSKTTXoM0Fr+zZ4kBiAuy5N9G0XpLl33WgUkFPak8/jGy+/VeIphvYGRtTt
EQY822664OP6ysCjUMKcartp9ozgZbLDs+GXBtmd9PUSvW9c2NK/+9h3rqXILfKWL7phiV+vEhhK
rXhOyUul354qyFOBvnIsWWqMORyYuhY9OuW6mkG8dEc0iyHyVT8a/7f/EL9c88413BIUZk/WmQnB
02UohF22xA5wFnrN8pYy9V8yQ5xOpgsWE0+/Two2tVX4YfY8AHBbZvnnS7xEF3KvheQuSBmeAJRK
5q26685289ewkp+W4mzXcs6yWhFkEKEcz137js6Dgp3PyOSUjy1QRYaXLwsaWnnHZ4XA/LWfbw73
CT3oFkVmiLrKUBY7EzbwekVTIUNz2LPipCIXRWwQLtGTPtXzY7PpUcTkvT2hUywj0kdacDzaQetd
RQML341b1iwnUq32PblOrYrcX8zop3yJNXqIMFtUGg+/jRpKXAkx0m7bG7G5aw1O6iNpWqdOlYf2
eveIqYs3x00U8y8mE7gRb8KdF2tQWn6AstY5+aaBkHkKwNxqp5DZXx84bZiwLLO0uXnG5Sqq7saf
R1fgRWmyINFV2PE5B8W4/ZGy4AnhD7mXzWjFN6+Ca/m18RWSkoZUCYaxbxShEG6ARFBoh+YBozSY
sZTBqLUaDEk9eZALS5S612LOtPU1/Kq/j4yhfs+IcwDuW2Gg9jerSMsJ3n85F/ioFRE19WWnmfvb
x4KHsLfqia9Ob1VR0UuDnkP8IqT2XHqYioqzDe2LlgdXYDsgcrAIfR3JPfVpRXNlAczOz/gCIW/V
AsPCvIlC1CkvJ46mqvpXv6jSTRMzhsSs/0TOJwRxc3yxb8yaSN8mYfYF82bJrJL9yLuDu7WPXLSW
HzHrI9lVWTR3XyQerEW0beybU022NZeLY9FyQc+SmoGdxFz4Be0dgstDB5eAwyTae0YubKkWyH5L
1tN+XkPMG0bEPghmGCvMZiW8zr44ZdGnaUFEIRTVew9mOVF85hIReutEg8aOIKTeriNrLn/bnX0b
4iUosBaJqCBdqbtMlqbDmd8nwRxMWHkPU9O005owQJbGg6PzPBBvts1QBues+l8fG75+yPGgq0M7
q9QZdQG9htuyXVJTqvo6IW179xq3ooN4ROebJNIRGUP87wk/X4Pbz8bpXU3993URRYGuU9Ip3WRd
g8YKVB6YgDy8O+2CozeVmkiZQrUNBfu33J2QhPHpLO8QPbxYMPG+8oBr3WsLU69Q9hhwoU1TVMfL
jCWMP9a69xt4bxWitcUAAnw1y1hW2eQJVxpacHcDSaY55eS4A3wZXJg1hSDgUWk2W3BzevR6luoP
5MtQBcnNQvO6EYkSu4XfgA8xiGIlap1WfMd0Xfp8MYNme+KAZdMKR8z8vw+12pdmWHU3WQiR8OJI
OBHFU7d34Ew6Xcu3wgtNgPYoxteusgww+oNpjao/aC899vuO2xXOhu49CYuLi87z0itqk0qZUY/W
zHpe0Zpfm0y6EHCmuNxvlI2BmJeDKJe5+p5hFDmUi7qUqa4o6dvvEaxZ6/DCwva7Nw+0A8ktGn5q
yKZtP+4IgiDDdcg2SoAvD0yv9QhvWwzsWbJf4xSeI9jqVtbtk8erDf1rH9V20a2ZH4Diiu1lJiT3
vt86VmrbtqORgX3fpU9jsqnCGl0iLV/RXdwmQ81MV4EY6nNsuPEq1WTsAUNk3tDGRdHA8kboNhHx
9O32zLTePbXB/YNDBWju/mfyWwi+k4naU8T+MdN+p25SQuYxHY11Z6KCQIRWT/i5hexek1lciPPX
z1mXmvTFbfROy5ohvgzTvwUz5+lseZTUdMt/9BUHIr2i3qgGTg+GhJ1hsi1mbxBO6q4g6nwdjuDb
8Hn/VfTplITbNIDOWdMcYQtc1DazNMPmdjg13HPINPnHbD5SNGWtLZzB1vSr2ZAaqZNoyU4GS75P
W6WZpFEvxJ08Hc62rBeV9DFoNEFQ+PwbSrmiHA/gpYzELFvOW29/BV/h3vpaSOVcnjWjr48FB2PK
+pRuDNXn3Hp1GtK1iVZVEKlsx5kI+JsD17C4xDvWOKhY0I8X95RsHh8hzA+stYhHdnf7oUV3XjI8
DONJ8Iv5NMmNWAeh9BiLDpFew8RbmEuDymw/N7zK04coR6hloqvja+ayTOk24kWmFEubgVaLB9Lq
aoTE58kGb56El6E17mwX6X4RryXjKDnBYO6rFNL3Z1wNdLlltrUdwt8yWxOw0NIED/Zo8+n1JhRv
YEp22klwZqIN+AAy6hwfKb+pfVn3TC/uq/p49i9CTkncvxbTnHeZZgryBa862ybuowEVa717m971
eNPrTPn4X5zex0VcXT/PpRxTGRGEGyBgE4z9Ci8LfWCO947+8ejoUfX4ACS2a+r+XGC6QbGmlHq0
DzUrG7Cd89C41H0zDUCQNM7j+/0kYPEmYaNKM1vTBBdOe2gI1f9Pod0OqKJ+DOYgB0do7iim4rOG
E8jTjxCGvPBZrMXfyfEeQK84qKKdvb2iJfpcAfMZod2gosAlUlkCOwF3Ocvf9yeUjfI/AuHBsb9u
8qTuamPYzvPOgIt2DeaMhBQDt38UJTaX3ynG0DzuOBnIaV5TfRuTTtxWsFWeekx0GTVbaite7kMA
NlqG8NYUBRoC+c0nPgHze3D4dQq9jFJGq5Qzbmf8etz5dBbQdtT6tCT7tqOzqaReuybIE5suORXw
OttoEW0aRO+lDEcwFqtexw5aVJHrIuahYufL0mlYBY+MV3/QeVkSo8lz+7U268Xvux47Pqr68qsS
egn1egocqwtXi2zdYLyrjNyN+o+bvN9vsfg6d6AorXx236RxnKC0ZL0CSzQtkJ0+L/OaGFiljnGB
f+6lynFvSXwJi4RHH8HwCMwnBUE/PobqCysDP7CPC7z4wpNwGKa7togEBvfrewbNp6T82zlDPWYq
CId8PrkOOfygIc7h7w/AntxGrl+KAHrMjd/UrUnhMIIeZrF1siUB3CsegvUyPm2TPXbsMfyfHGku
L9ifqNjjwseKIeO3rFKDYxqz1AHY8CgndgtOgXA9F6WfW9yAc3x7ukCaUXrxiAc/w2bLfIIb3/0Q
49Y0w0g8E+9sQ6SBYkk8xgLzcrexCUmuO7DuGTb56Rv2WgE8T7wj5KVPk4RbQKxJhhlsxenTuDtq
CG3IyXQxg/YApan0n/MowuPo2pizLi6DgMmWiXjLQAnxH83ik0iNX6EjDSBKei8OWWKcXtvZXNey
jtbrguCXgJrJJFRo2awYWBY7qQRsQp7RjysOsssE/r3R/dACPf5fX6GZMupqG44T0fbeqCZFcF6z
ZJ/k8IXZXr9pR3t4+c/KfLOIV85thzqkjvxr1+ezHiokE0oVQaRNa2+D5jEJiDKzOprSSbFQ9dwi
ivT1TLa/sIJFxZ5taCO/EZQO45XUIucNguTLC4/imkOf188WBMD2jp2jC8B9gtZgCJgnnlFOOWV1
G3L4v8jpdJlq9Zle60SH9V98ehc8bSP7L+01sqHFX/BGlGAzMDSRw0owGuwSwZ5A8cWNzb1s8svL
KayrpptQiUmcTdQLauhV97T5N7AXWTHS83QDacuoLZqOV2TwpJi/ayub1rS1TsHEUPjgG4KM9VZb
VbAQkej7DTTLhnR+IfWh25FlJZUWncH0Wpzfc+hFYfT738AWGK+Pyhr72amO6ZXoOrckDuLsU7ys
RAIVHvafwxcWKsBEMnuWdWpRMMHKj2PYGw0LqAmG4dtxuRs4XJGpZkcYIgzMs9q1WQMT4Tg88+AD
Ezuk7FV/Dgtyxw0uT9co+u8qoxCXTmMfUe5pu4p2stgjZWd5y8vTnrndrLDx9TUYKRzPF+htqZgL
E5Bp8RQJe1m+gxQum8uoyukra+ltPuLPIg8489F/J3nlzW0WXODF81pWQRX/YHacYpSDycX6w+tG
ABbsi/4CEHfaAxK96jyz3ICnLJPbjnzlxqcITsLb+mtcQo/cCBKj2T79Q0v0nfqliYUyU5jmiO87
/MLZ3kvfEQ8mTjWxsnhaYcB4s68cC7jd1iznmYuCUukloM5sM9SdBZ524kvDsUGiABRM5Qzi8s/S
i6KaLu1VHVTqWb7yu/JKWT/W8xLBpQUAdi56R/Mhv0hfQpBdabkGJDuYBx0Y3ad6a4rfwINLkE8E
zJvCRekGOc0RMMVpGa9pFYOz5wl4HhzR9tNlRlawBc3I0z05QMvuI7E/3Ln73II1BX4Lnyq8a64V
R/NiDmwCI0hofpvlAfozdO5P7vw2i5o7DcONqnBqNXwr8vxkCeCpnG8gvtBwKhFeNf82cijCL3Zr
jDWO8n4BFbep3nBANMMbLM4+KrI/S19boqcv2SiQpiMSwUw13oWIH9GdG8/8DhqFJs1iMYEsdZ0z
W7Xz4PQRGir74c13wAmic7dDi/ysdQvdynVFjBmu4XhoX3ltFDrpvWftxYCOPE8xqFk5ZWQWQXqr
L8Jcv9I3l6tbVV67L0pdQLEk5YMt7lbkCErlZQk1aGmjhH51CzWYEADE7mjWI7ciqbCrxTjKCen2
Y47icR2sKQMN/Wk/MIdTQVQM+j848BKvcvBBpzqW1bTk97Uaz3EXH09RrNhMdhaIRp4DyV1/GyCD
HD6No+7BjyR/vYaeQ6Lz2l0BrnhaLmWiS9qdfG4EaPNxrYiLnTlLldN0ZqsDW5cIpcMD3Z1+aau4
bnNBcvlt0aG7U4kUarc01UpNG6gNAg6LClFkhDlCcNuQkVIvbMYgMID7nmCTN8ojUhR5Wb4iOYwV
pvhSB8bGT48pD2r4BnSCfCZMupMk0UMsW7me6iNCOOACMPA67R25soUvoTm9o35gILlsdNraBhcu
D/6fPX4dpKdiWz4ybVzZKJ3u9k+nnSBbFWilFJiMOfqP2Lffag+yTkpCV2/byfz0EupHW5tRycTw
Dqq9i9i01JzagUk6YPDJEorEuEorK1i8G0LV6OudPoxrs8BoKvFv9+pneVFEZpxITBpIjNe2wq5c
c+EcWcGm8J1qyX8J16LVzDbfWcZzgs85KgJquRzX96VgcF+Exb+WHxWf9yCXpQFUFzcD2IANf8pU
PRIZ7M3ADH7lshhJPKGRYaEpLj6J7koGFx+c22J58jl/wpQw/K6ixRVRgCN0kcy3UdUNuDYoHQ4L
/EmybVzlnQJcjE7xFsBCzrYdLEnv88szebKlATNOyAAAhxngbekBS0M+aItrRrukNcaJMK+609WA
bSBmi/5jERtq/Pmxa+ecFli1RhJimH4I9+QVsogJlHyr+lmlPq7frzd5c9e+r6hkqimjh5F2+nnN
1I30RBmjuRoaqosP7E0WTRHxhcqvzKLOHZmaUwDgMBDMQTyvTNovDTvX9KcZ3uxJ6OT4O12N7gty
zJUWEv2Zzp19WGKOMlnYPspFDL1UQy4pcnLFEr0G5vlB1vuLFpq3YVK74OjGbuuyz6PsSfU6BsFP
qviWMSY68WmqzA80EHfycY8ToI9e5Py/2R5EyoEHhXOmbYYJsKW46LdkBIIefAnS+ZvJ+R6F2svg
O1hWGaYE0yj95t/6KkN+razyCeExCGweU4SOYPe61yzp6RfmVK7xP0YbZvY2Cn7+9fsYHRbjW6j8
uctjhpOVxxlyDhiJe2+APfFRtrM17YQWHoNjzFRddX+1T3NHs/WjvjTt62zrGiNsE5Fg51PXa6JW
1AekuOzEq17f1eIG2dMRhVQ0lKfggKsXDukGszGfodV8loA3j+JlH/18cO13HXNAOz78n+1JOFeV
NniUAFKxh71PckiKOkBXCZojVHORYuIz7q89fRKntE5Gt/CZQ15c9bvM+oh1vSuM98hR9yk6uXuU
y4hudpdCCAq6pZIa8BITTHbR5jTMvyGBNpkPSDbPavvuJWVECnMiIqEizuhSKcD58SPZaWzJz7xS
ierLUkM5gdIO8TruGne1/+lbvBIL/C7RvKax/Qu/FrFM3xRL8jywjCJmU0mh7BuGtzgTBZKp2hNB
heiUtBrI0Mrkh994JqWQc5xDoAbA8F9MywhIvvSs2PSSgGO5PbPIadkAm5wQDcPbrt27zR+3sb7E
O6pE75IZ5B84A+CcvFqE/5+koKRbf6nZPfm5v8/Rgri8eMbeE84S85FSQl7iS7EdUdMNtCky/2nL
0cYx5mbZc3CKb5qzZMkBiuL241qGqDDd3mzGQsnDkzGaZX9sLHOshOeauLvbHKQwEHN4aRwztfkZ
pfReKpy3WtMHsV6tJQKVW+fAqa4WEX5gIty3iQaUJpC6EfYc7fkbfanBA2wejvGYQKPMAYPc29fX
XeXRZMHw71/xFsvfs+O65rZXuFbq8/usiEE18mR4iZZZuzzfrmL/LLydlwS4ZS4IE9m2GsefpQ29
JefrHXOZhUsSIxUrjaWXi8m9uQ2XqvbbgI3YfzvSk2/mG2ir2XFOjJzwqe/05BoH+LbuLE52C6jS
GKUuJuMqMXAnEmiz268dhCIvtiPLh59IzSLKuTQdfe0cSlJTiF1N7axgdQa81Z/VayYxIerohx6b
mIHeajMvTED+TQU+jTx3nLAvcC58wMMNafxx8Bm7OGyYCGTrnEvGEx6CWVGHnCtXowY3cZwXYToI
ai7xXBMfSZANUpdrAnEWqnUr41/l2zsXfpmMfiElvsAGRDPSn05tc//VPCKzoCguthM81e/YGAeU
0xWQdgxqP6PvAgz2L3QemyyDqgYsC+vY3E9qo7qdQn0juftLcO7GZhCww/ITdMnhi4EO1/usIYum
1yty/QSKuo/xRajcnchnzOGxfqStF/VegidtOhkc112VRpMRGrxSVbH6tHHZGfSjF8kAjCpgkMMG
iFvGzzNYOYqP3pwUHtBS5Hez4GuRwRUU7VmzqgsMg5sgkkg8JQnbTY+f15/MwJSUzUUm2Ge2k3TV
WX9L1gkYf5095/B6qkgGoz6RKQXKNzHBRmEtol2eL2pfqySuQm8ajWySMlmfVvvtJ+bu6DLC4RgR
Poeyc4FPz58PSRqSECX4ced0wMlyNCFlOXG0dzOv4MAi9QBF5q7HHLqnIKv8El40K+bnmo/QEfD5
6BIc6ZD2ztOoz3hJlamh1xNPttjNdPG7Netlfr/sGPBPbKxA6kPPv9sPW8xUbl9oMjBbfRzri8bV
J5TOucDkTApYorkCDUva4gQNScr0Pmg9vpk/6AAGaNHqhsY3DBCbThS6HRPp5cwSxkyJBMHENkha
mzaTA+Aq6DcJd2a+LF5LEXnC9iIfqxIJZnerFnA62WANJ+gOLoEtnMudXN2UYSmC1MQAe4vUwK6C
Pwjq+ksP2TU5IXNAUAx9d4bZxjPQ2lP6RpOyStbIZKel8KCYRLVtLnPXYHVeadfvoo0DPTFcbWOb
MywAPpjx1RFpwnsjKroWbu6kpAJQy43tQ+OQ1bnQ67uNZ/7cfKBPBWA+J28EyGaqIRRQhUlLSttX
ZH3aByIPIbzCNe+XjbciompP/FC6gOsOZGMfORloucl0VMOqkWkMUssY2Q9qiDSpSkCZ+dd2DSHz
QVq0ZL0bFqsDXSYv+DwEpRUJPor1pLDiCkl2XBP2Lj9rIA/k/+8YWS7+fpZtsdvdYmTxtXUXJ6QY
fsgJffxUkfr1a2U9KiEbDthxWLqrQIhmIJVCs3LeJG+f0fnoY4kdPNVcNfnpeEJNHqi8X41rZ2Kk
VJpc7oMdggXGW8qO33issmLaB1DtcmYQNzhY6M5rAZhlZRf7e5IdeGrmyZQ3vM7hfRIvMBOd/3aI
7OFA7mPwb6K5RlylqiU/OMOhncEyYjKTNdcw4Qqk1jBzOE+Aq82lfAOz4o3ITwIKeAsg5BG2X10j
0C89y+qGZCxowILBi746A1oYvFTAeUsMUoXrqVAEPgsM5smiqFE+cJa1HCV9YDt4gkz76uIUe1js
xlz+oaWjHeWGIB4Xl3RfxDEQ0+kb1UMfBl7CHTzPSv9k7b2BTxqG7iP5Pka1/3cdCv9KWXPI6xXM
PNl3xvvmOb9KxzjookDRwLuZvCHaWyJDEjt94YKsRW6uZW03znzSbu1yPrKYvD0s91m1Hs/68LNZ
t9VHOYYzt1CAWqkaKFw8JOtAibmOg5J0xluOKzNCbgTu1cMcBQag08vy1SRPnOOauXmfdkvB6Cr5
VDRIeQ47JZdFUYYhB9zjTNrFZwel3w+giuFvC9OCaYmR8lekjxMkT1bBqCz9xvtKJ41Kg0ls4aIu
nRyXqRsk0ALiKl5GZfHkenMZeNesQUHsQeR6OErq3zO9OcIbtf/OEn9MXVatgI9XMLsW8A9ZIryV
IvNAbqYauW99z5PKv/+c0xwno0J+RL4No5DVhiWdP0MpBZvteavQVYfi7Vj7YN6eyShOeLG2Qa6W
hL0bmhYPDN6XZSoMk+ebV18HgF8DW5bnwC56ZmR9KpQtarmKiG/I++VHQa9M5oArkLk/uZDYikb6
GmgcrDVWd3LtKd+YIntTvkjp/fb+omM2h5f9Yc8OM+D1uBTbY8Lyj083iCC3LbYtYgeecoA/CNdQ
MNHCH6idxrWoJ2qfcRrT6h7U//tPgw7mNtd+vPjcdYk6NY+D2nUPJB56Fpl+iY5oLz8uo/b0UrUv
oogQTTU3aWCHZ+SceheE8oPHW/HpCcGTTtdbwzRVwzl/45Q4e3vxOAc6utumTVFKNQAQFw2OKj1e
78u/aUkkeeSpnQLm6AQd7eHqE/d8JTcsAEhKdOXEPGmANAHXB6yc0Ao4lC4l4RkFvj87vj+232Qp
lA6aYugxxQwIwEGcXblTrr9J1GCTHi42ha6cEa1pmTejT9eYSTTuF+qSDSD+MlpTLDfVlDu84n2y
4QbZIni426HHDXEnkKfnz3/R/UxaebQdDrUl0f1Qga1I1eJ/yYcxtPATEJxaBrRKM6iDaiHFHLR9
QdVdGElk/uybQhiUBB6hHPbzrhxaxU+H1KqZzaY0WkFyMqhtzYwrtY67AtrN6sSlpT59BkUEBhsa
x2m7akjqxOfKoFc1r6WnDEvdSKUwdiOk4WemR2lBWcI4YImJuIkrHcRbhN/isHTfTSLPBY0eBjTm
lrAzG2AX7OFzSi6lM0GSV4cIFGSlRzlUyi35SRW6Dl7y+T2Fx39STvodQXDnTjmr6GcJansIlIFp
1jsYiJdArsVEXqxq/kjq399sC6HHBVsRi+MNP10S67MBZDo2UEF1wz/3K1ZfeQ1jIsh9mjmM48TR
+R4wSdhdzdAiaXgVvvSzktnc00FtFjOIo2sdaZrXhu+YDBKXgdlJYBGiz2oX2ibRixIorJmEYePl
JB7nBBUuieqgPjxtWd/brE5QEHaTqm7HgwJFixSEdvxNdgZxXwEFGHiwofls4sfIUzcIpFDVCghM
nfHGeudXFSJTMDKhTsh1XFncIDCvPIEuixUkdxU4MmFRs+us6L6nSIB2T2BLLRPGDZHlcQiBLgT5
G9TlFLEs1Z/VWTkqjgRCUFxkTvYTGqO/sE1ui3ngirXjOs/fAaK4eRBSzqLRUtJ9q01uvgSI+OnH
X3eCAE+CVnFQCZ1MqMJYP01k+xIYoVRBnAtm9gntEWw63+jvH1uiAquVisaanabvQRegAlTbY3Bb
e5CAedyK0gbXHxRs17Z6yO0DiqUr+BfdtkIzQZsYCWvkMdAHu9qepUsBHQv3cFM8ywpyatK83LJF
BS0v8f2vBsxYfe2ZW3dkt9FWdGfj2KUum6dGEmyox6cXID1I4L+RupFF39Kz9nasugmEUZ+LIjYq
WcXtRxFchDcCL7JcwanXiuXWaPst/cEgrMGJosvW91xGS5WjCxfXGT2kXYKDB92WT0n2X8gO7746
mxzdHBalxN+9+8yNZVf4I/re9YEveXEhyDSoHJrR+TVf8akfq8krYcXPc4gjRba28A3g0id2FKCD
pDmhnEyJotRvGthMWpNDrdE71uvYNQs2AwqcIda4EkvYAVVn00ZC/m9rZOpIIUA9VncOICHqka0B
KDuuqZKcQZBZsBRf74Kg1qI/BR0v3W0PJHABmMsy1J3CPQfYF9So77vpRxZS5YKx6bjfxqKCANt1
kLke3A2u6zm0Hy5lZ/hxu7ST7Dd47DvtDqnBcWDjUvYIc4ApYAFOXKuRo+Yrwzx9zHc95TfTGjzG
SPG5tqYjPikW+rIRZJQhS7hIJkocjEPhB8nIlyMu1eVaQdg/2SWyauWIBYxKEVY8EVPjbM5ms8nq
73aiwgnAd5C6psxId++JlGH5STlWvCXALG8xP74wuTrAHjBI2rGlqan92ix89ODV0Z5egJRqzvAQ
i1QSLCznz8NyiiJMqS35gu2bavdZ/19Rk9sKjNTaHNem+nl0fJJ0rV3a47gPALUcQws4B7Vrf630
vjtMFqDw1Ea7aB5cQfKQQZN+v/OqefbHfQC1xWVortZamMbEP2vudW2um9wpcrqCtUQbrIdnZj71
o5hGFeH2ZPagL4JlOpFULVV9i1qxaFLerY/2MA3B84YO/DZPn31GME5iy63wpXqWFylJ2ocmcSFc
HSZz9CsIyUSwGCR0pB0kOkv0BTcvBYIg0v/vsUMlkfT1t+UP72ODdHTtfUr6t3FsD+S+VXRb4q6D
x4IpVcu9VPW5os1LlSVMvRDaDB3HS/spC/4c1vYJjJTeuITcjNn0Ie679OiummYtlGAGUDSPrr9o
MMmt3B50Z40wzANu5h1NTyOlixXcmh8PQ6UVC81xOgZtmUm5zU3JyT+dxPl40Bk2BukI+Kmdt0Wd
MOMtsXL3VJoEz5LKTqU/eyiU+PF51nwq1mAgyV7YgyhlT4KItjucX5waqLDZ0VNWNdlmJkLd+PZV
HsNFXUfXeQQilvZJGAdv4bFlrW5kRSt/oaajVFK6TZo+dwbZe5BlWf+N9sPshUrLAIcNs7rfz/v1
K8N9CLwEap4w4LDbE08JDqSTwG21MMFqpCxKY/urORTJmrrE6qpL6W2VS+6YabBY1ldYHhmBTMIC
llBt/9jirt3orehxm/f2K2RioZpx+sCr9TUJBijCqpNu9N72rv9XzxB5YVzOyPfRcP1gzvIbJtQC
Vz1DQEtRErx+D+phhkLeSI2rerQO06eJ4ivkOuUZmg2M7ZdNCHJFHvSo6RuJH4CyeExiZj55pzc6
FpfJ6+/+UiEl65D7ddH5Lrfuga0xcsA3ICVawaH7q/sFXk2PFOi/hxICkDycm/qxx2dKPDqfDIeG
W5Rs7zQUgyLHz17t7+NONXClkdEUvYcZnthINXcinScV17A//fhlDhzISTn+sVMZtCCoyx0lZYA3
GGTlsf8FsZTpHr4SmK4reWkwjJVhLuF/xsp60Dh9i2oP81tSF81psN795HpecuciC63nQCsbxRA2
Nd+VBL2neAwolPggpjc1iOdqKt0sSQxoBewlVPwlAyEr0C6mrXFGA1aSdX0qz7jCOeHr4XCFcnQh
e3S9BsN9qgf+l7of5gB35EtHd3UWsfrwuf1bOivI6UbW/6J/oGJ9XN8QZuAxatP8WLE7ecvgXtJ+
PEgMLUIxKRetczP9vwF7RzigtVyou5v1p5aYj7yAXKNoxXUlsJ0AbMpy2a6CEc3aQCKx4QCgU5On
NtG/NnR6VHqvHhJHutnHGBpBkaFKKULTafRDJzZl0E4j1skKkslcDZV+CR6TXFJg1ltatLmRF7TF
RkHTcmJw/alb/+4M3w0MnWeP1ZIzdKYzfyxl5DZQg6nH8FeQKvKOsTLO57PloZ1QvdQaURXDOnFD
Nog80w6RQ4xPiQU5RkefSoI2V6tN9gOhBVeEjayocYQnOAkGh96axtjIjJC+jc5ggreSUfHCUkGy
rJ71U8bIv9OHO5lxKQBuFLz20CPjyFQ+sXBOhYtQ8ylT1i7m0ZCA8qxMJeTp4WGOlsl2QUcnkRF7
Kd8pXPUwXHUpy4GfxcsruXCbeZTpObwTY6fKyVMWspZ8W5BCsJAqGFb1qZJSazPyfBoxMZwfuaYu
TUz4a+JUFZ54BqtKgi3E9bepkfSUvlO2yQn1JqiE0nLImuNWmOsf0aDn0lmaOfS3ijV6tpsBYsni
ty4giU/QTtMF569zJA0+QFwzoQyf+bkIZigaMFO/0ek6mBjdCbHHgbUFf0MqMO/VEtJTDstQG17R
gR5/imGH+kHDWFMvgH5Ka8t07d1mpSCA+YC3CNShxp/ErE1yiFgyZDW1PctZ6TOy/eiSJovJGZEU
GeqWCOw1UxubXz/0x16oYr223ISZGsfzgcSrmr+VJbl9GxEVgIgcR8Lli4UiJ1aenoMPFSECQhUk
ka8QN233WhZdbF3ynujipO87zRWmtoSMngCE0zHpk0JTyduVGQ6ewhtnDUmXCUFFBS/qVySoL5fG
BtDNwYmEzZ+O2enc8CJFKMxf7pMYaSAeY3Fdk9uooS1JsYCgTAwP5OKua2VESw0/ctSaMtBfoB1r
d9MemPsLc1Nnxx5i0/yLF3Y4vRpZ0Iy6HFHkxEW74gu8G4NvhjgeCE+Gyau3cYVl8ZlJuxRIo8kL
jzFaI6yBf8xGaqaYh86+8yQwdz5WgA/iH3V8lWPp8Wk2d8rscPcTtlO6Ow6AnNpdGtDx5/xL5CGa
U55/cZtIxTYsEn1y4gy3FX6XUzVtnBXnJwJMxBHUPiqxrhytzWvoEWdIgzXRP/ln3bMKFeqiuUch
qM+azpkqdd35gjQXKntgPRmgayA/7PASV/b1b8lFyixoWRmmRMKkNWB4PkGUIgcCenJAcq0H4mCM
q19iAEnYsWYDVPVLNSgVP/UYldhkYp85akUXxtkj8kFuGyKzPjQ/UPemtiOh8/+lPgF9yZ+TwR4G
f/LbzfzlMTEXk1EYtwUtkJgBE3sa4ttjw4cfcYAOVjgMbp1v34f+hXKQ6T4bmhFJNsn7VoyKUysy
6n9FzT7tb45Hyd7Fv1009anLeKSCfWETPmJzNew2h5uulyI4VjQjCpECdyrQh6szw5B9YRoIwKcU
vespYnKDYH1Vnon53YD5kJuu5CnYpbSG3lsZGnuTCYW+yVhrgcjvYKdlFPSASvfVR99No3q0szye
n5xqWEGlcIfY3kl3Ya7DrkT59JLBY1UmGhj1kAghb85pS6tW4Dl1TH8DRZ8wW8pKa5jFDDgspihA
L1D6j3wi4fS1srXw+QC5lr4cr8liUY0gZD9+c20e3zLTij/JlBIeByWxMikQ9/LFveuLFdztEEP5
TqKuDd60NlVWd5spVqeRx7XlM0f3AoGykUBpl6xMVzlLjeHLUdNCbY/v75fSeF/vzvuq3cwsk18G
Z9iQPk9kzY9fyF/zb4r1EBY824yREv7fZTtl6z64W+D6wk8aPdlIUK3ioHT6dn57Vw9EqyA9OziT
rxrMAZt2/N3CEPVhbo0DFr54mxTEFa4jewj2+/Okf6Bk69N9A9/2NRFxDFB5Q75L29KxmhJeynMv
Nbt7sAsnWBwRTqfNfdrqQsv5TGHBNSVIrwq6Z+85VrfzVelTFzhbsXk2aMbHrGfE+O3JiWEpuEm2
zej7BouGFbbzqx5r0GT55gquY83itimINzJZlPubluulcZ7gcneUH0LWm6x5Wh4R0KTSo8ENaDx/
jkiE37RAwxN9hXJmfppyyS1I7CyCXgJhXL96+7Ma/ZbKw9SNDdGqEzriAPRzyS2BedGDqgnIQUgK
qjmFlX1+Ip5ZlOrGmACUZF6pQJk3rrnRMnr3BcFgxCm5EG0zSMcU+wPZeUqcoW360MYqJoX1dw+/
490RhkelbctX3qfuQNJwM8oG2Ln1f9d+DzTiCSVy3Be8OzM1bsmZWuUc/NcSeyeT/UHxhJriOiFW
39n5fjj28dVQjn6Yh2RUAiK2P50Y7RJhkCCKnfRd8X+YbcrjLzEw+psxslI4gg00etygUzVVPq0C
sh2lt9n9z4egLyhElmIhk2Op42QJZA02rXbVGTUOo2x34Mlt/mbyz0QCdy82fk1uUooweRQMLpGP
AxiTn2rXqZf4i8sf9fDZtufkVcTzJD87OpvdqHRZrUwvTfGLtZFNJILrkX7GPOVdHzFdDNNJZlVa
LI0bQV9mrnybxYiOd/q7TJVkrFFECOQ4oTZY4Q5SqyLGwiOYbbDZTjTHX3r22UPQHcaSgTuzF3hk
gH1BAQSw1nyRAVG09uB4cABB5OB2lA79FitlY7xRyaI6T+NlKvsKoYoma220+VV7kdS9f9tXcnF2
ad0Yj/XXGKMTLd/ZpeJ1mqqAPz49EXXcesF4FelVTjFUVdxP9IYjjxEEZ312GhTsWvFUf75tlFHN
74paY4IJ6MiIy9LYcsfPp55opPxh/JBrFtGiTFgnPv/e0ETLvv79MH3tsyt4mZ4TxeH9hcUkmBHm
KFnLg4yCl6lbgA9M9B7GL71XJSL9wvyyFwJxsHYYp5j7iPxveoSPP18iqmBooNb3E6c2hlmty+yX
jJtylWvmVlocTOLvjcYlbsl470iuTeeNX4KkPQ7g34cWT50ce679ooHFjNBhKIfIu++iR3DIdU1U
V+8WsrVA776iSIuHCr59J6SgANeDDfTCtDkk5kieU4ikt/q16jOKdi/CxLUC30lTXjhLaALRDzt4
fTspcNXz60hRUL5Lhy1QhRIuQcAXjgBlFSFJdb7REJHtzItguQogBsM1VY3ANCn4+4At/gKQ7G2b
HN0hWOACBHAOX9a5QL74lRWHMmd1uL4a+4Tvg7HLSieM+OuL2Pw54diKfy3zHarfhhVbTO4DkMQH
aFsUI5iYdHeFTRFR9jQA2Vld8LEW6vHBS9OjgmEB41Uy4So0RJywaxBUV7T8ErR9w5rbvafySChg
kyHQ0J9Src+aAFNJ/MVTxy9sfoIVCu+9r9OH2QeZIGo3bZnz8pYfJwCVia5VGWeHAcn9+jC61MeJ
eTPqI5O5Ysz6RnmtskdSKYXU7RzXaUKXmHi6TSZ7tQRt5cpbcV0ObgQXM8gHR9ZGWc3aigsYIndK
5+oFm7zWZ+U3rP8NU/BC/4WAbN0vIPbO+ntAa3qhyjo6wHqueyJHK3M4JcIDlD+nW3wIHp/uJ4HG
9Xn8FdiRjgtsVz7Z8OmQorDDWoanL2oShpKnjQron22uI3t7LL2Fp4V4/gZM7ex5+O9nL9fG1mRH
Q/ffA2EpPVDWw6kOcJgKlsNn6wt/mY4d963J1Uhzrhl84QFseGyOp4nkIpzB01VcDsh/EQlr9QhW
7z1bYQTz1gaFx7DrGLf0czJSo7NHME4jk59mWyomvHU53hvFTYvEPzIc/mMlqU/98ZtFtVCq1rBi
WkitZ1rokEyecy0jdrhMnZ4GE8odskQs7DKHNvO/ERg90tez1/aSuEo1tivelGt0aQEhmS1THepb
d2MUIYlaxsS3BLm0cSXQ4oW/fKm6GWy1zGJBQwjFITMX3d/zkfaxMpzS1smvkosCulLUKEakUszP
LFKOlaQSwrCT/z8EBJEQKB9easd0VEfvF4wrZoKkgCXZlTZTun7HDiuMsl/tWQ8BFfa79+DSevad
t99yNpxQuzpCtZCsmfrPWLjc6hD9ORWxMjtC5JRTfsjDbwrMhS/+qWcnvz1U5WGPIGyS1W5Rss2y
1SIkTDx0uMaCkhlX4B7L/WHMq+dpIYJ3UYGAt1ZkBd3K+HThLXuWd8LcX8H5i+U2RRJapx6Re9Pb
LUCPSD0Tg/OQAQPzlJmwZ+QmCuIfJutzdreh/Ykew+idxP7eUOrGq4Co8p1yWxc9jsfBkajviCOk
1fmhAlVsSISUi4MlCbyoRNd9AKqFMEwmaVXoFe2wqBfSTStuMxqJ7f71vhXgzILZi909uY72+0X/
/0NxEMoCkxlCniS57FZKnzFDJMz1/CjO5N5oB7xDxlAAf33NdiNKcRsed52GMXOK9tFe+pEQ43R5
L8tb+OLN/59UGMq7oAbZj0sRRxlUMtq3suax3RnvXc4xAvJ0QFP+Hp7UUSjkaYfcdIQXtt6oE2Gc
/DWDGFzFIrsq9gx0pTRub4vjuf+eMwaOWf4qnC71lk3bNLAmsutfcgmJkGTfo27AQHrtaw/wtz24
vqh7p+l6DzYtRRRMdqCVYKMUZ9o3jfn5lRW582RV1zVQKb6oCbbqbdhepxxJVWAlutVg8JXWb3W9
/4dx6WKrH7NWmmkM0pwdgOQH+GwkmJPNEc4Fag5yPOWngTBf0rr0/JUyiJoG7kB7luhCKgTXYXSP
BCBEAEmEfN9CVc80jQLniCZaU1FSWgF1ZK9z0lpHEoKbcMMVOUB1qH0LvkVVVda9wOf/ACc2I2sE
01E/RGauo9ivPqjL17h7rD5qJ3cQb+IuMGy37JK83IZoIz6lO23aDR9E3f9JWlsjnAR3AyQs/8et
w7ajA7s6KbPMSf0iHw+WIAbVZcCMXIVg8y/qEVAyf2UA2rm5wOxsg/ObWj0uaLmqAgLQp5u2RV6F
wsGIqHTLXxgmo5miweyqORQfNw8nXbKxfzkwzNFTIt8XZW4K/znrKRIBpM8b5AKVF8S3BHbBsAdb
d4ibZ8d2QnrZXoOFbC3m5SXB2rZID7r64V3w0o04LLtWTiyV/4FaXid1TTTJwsXGoxCpwDeGJGtI
Ggn8J8dctiqCogJs77R92AjvM7O5/uNsZ3uyrIkwxV62+7x0H1cwuqE21oWnyRmy96BJFG+Bh/OF
94ziFTZmyb28aymDAr14CaWt0+QBPtF+dZgr5g0AmTbinnZ4/NmqyLbCpq8ynMbOpdcuckkgl/J6
CiGiTtAwj1JjktoEerXZ2mBKXeqWBGnGDi/OUuezspRqixkMWAnUsghYtJek6TwOXJ7ZsGvhfClB
Qtvh0a+XLWeT4GporALcb8+P01lPb6AQ7tyhe7NmPLJl3PUqJB2EFUyhfuq1RFoBSZZOaToNx0uz
d5pFBzjp73vH8jKNHwOlnY8+wQ1rncIUgNK66B4bhQgTFSljIHIs3VpWt+KeNqlx5wjAwv+FeWBf
lnq3MgMR5d3kZo4Hzww5dZVndXxspGy1KERXvNQNr7Zi+DhBoIlxlfa+NSTPbgT3osyZTgLcmuGt
F66FJyZ2LgkgNCgue8/GnatjoBAw/3z62lBipYx6snGLxv9nZNbRaOppgIs8iuUlU0TftMhCBAvz
YhO8lkwQzm26hyZKDO3HCb3+vtdh4u1tLmWoaYslCUdyahGwvTMGZ++NGJig96c+9NzeC98JzGpS
Lut0PbLfiv+MbYo0FHrbT+QJPoG5uIxiRwXIxuREwwexfeF6V8IMWbnQEhsT6HcGs5YgRYnIOm+C
8qauhMP9dz3kSP7ZDVKOjLeWyftPGbMuy/JyT/xhvReEcBAx8t/xiIl6kqDX4cLe0k2B5QLUDgIq
Gv1rQ25DyDBiAcSNmCeRw4rL/86x2ViAnEueM6wd+0rtcQq4WjNYBuLPuxWPE/FUPu/qYeNeyyq3
zN0/uOfKEgNVC2lOYjXyNm+uSVGA6edoNpuAmtvaERqcJaA4YV/nXgVpppU7zEK23aas9tD1a3eU
AupeeAB1KoXdeStc2wWcXbOo7H4xj6d72v9wYq01Z2EOKCt8oSHqwLhl0CEQ102fvQcUQ9p7mcxU
egP6QqjHQRz66+yc4iZpdnFZW2BIhssSYsjY1lZwdw+0E/c3E6TvZy7QO0Q35cb/3Pn0AmZkX+dz
DS50R3lxfEEM4EGNoeLq3a/eX0PGBgAWB6XoncUqVhyjX3rMCoGwg/yEQaIf0RLfKcFrUeuqXC/p
srEH2xh8ZNrUAWl5beM1JXCU4RXvFLE52WXbFQwzhSYWcVNPV4Lvpye+Rqf7iRnGqD9EXL45oogI
UGFD9A7mRbrPg1y3T2iAkCwHI6BC8lazOZk2rG+TUDM3bPyv1aVqxB3EufensJ8Az9OFQImf4EO2
92ONsxI4uB6+yE4/oeSlJ2DjMaqU/hEOOH97oDymkCX4hgI26aAAK4R/6WHRbKmuhwo9eRGPC8yh
13SPmqbxHxw88o72XgFOR1IxrU+6X3b9kgMJIqnA4hLKhyspzWVHnfAKxC0X9RG/fSthVtJm+HEB
AyAO2jqYyl63DFOsSIpRNeM0t5EhZV6SwHWfBK3BAVcNDCQv0r2uwzzAeM/BjBG1iQSL3nWFCd6Y
71zQSbuU9bW2y/SyyRYR4SjB/bnqpQt/nt/UahS4ifhcMhTWDV+unLsWx6YbWICvzg1+7OZe32kB
3OptZdIn/emUOZoyHo3T+t+A1DQEM/SvRVGuCfJ7KyS1LzhZN5qRILOSpr0+JyZSy3ciXy3f8Nfm
wP54UHUFd1ExHS9t6zm6Gdlomor1moX7RqoWmcgrQ5F9VJvC0HRV8WiTSnxzhElQWIXxQku0h6g9
aROV4Er3OnutO43HBWya5wqnGxc8SHjdEOa5XVkXLobXEZmhnrZa5rZ89i/o1ufa1LtI3RRZToLi
gS3dphkq8vvP1+JJKlNPdUHo5sbobeoQL1SmoigN+LuEX7msHWzT3qrxDr87gkxecYq77v5CATut
h1N+HKu1eiGx/FMBsDLQx0REogQmunPEmZlJw3ZfRIF1n+FosTelZ4Z288Qz5S7sj9cLtzhZ+/z/
k/qm1xnxJiFe2/MwjUnMaI36oI59KAqZNTQK9PaWLRZ01vEZ+s1+5g0AiUU4cqh2Po9b7FBg6Dxx
ZKFvNNr44ntToJ2scSMm7UcCDd249x092/tj4ol3BdCCmietNDBNW0ffzc2f+lPYAz7c7aC2AUWS
fxbLw2pqHJuDhzxdbxcGuNoWvDTyDr0NzvBCY2iPcsLBIdJ6l5xpdroK2bv6bgRTHpkmhY5frD9u
WTkZ+vunij64GcbrTU0wBCEfhUaygnq/Poi1+F+/6a3jRIIfEF2cYAEl70orcZfVnhU+qCmVZWXR
TP5BYBlLQbvpBx8LtvDQZOfQnVJ03ChFpC3hucLZN/nBCh8O6cKJ9Zebbi8E0tNeNoMEIkMy7mjp
4VF3a/TEn2lp2p5wQCQVL94tSbJCsufiIXqIdlqADtEv4rCwyXgARNeBkFMIW//awCbcErBg/yqV
BlSiE+t6eBQieNdsQ/ynpioP19ocR10k6hfo8SGsyqdt/lPXEFPucDKNu7Z37wDe+HOQGVhMfsag
eCQX+4Y4Q+KIT5fcqNdVW45SxqySbFJqIUVY9FBj/tbzxT8X3aw7CwCk56V+YwBeNFJGeD1guPZo
qDH/8yocLK0KQB5nFcCArTOS/0AHiQmK1RuM68AZOVL0KMd5LUP2msdxcP0u4KzLaxsKPFmBNWJd
0Qp5rYtVMY/rDa2m3KTzWgGN9VwJGAPTDvsmoUBMlaaJ9gu2Xz0BjpmjW2hiLgN8lYRyRqFGc0AV
d3G/9B1Ya5BzvkwVHbn8aAoxT58JrwMktVUlqLoyOi3VFy0eRt9EV4AHaNWOPkZoMd59it2ZLbk2
1do8m9Y4tug5eaqpszqFIih148TDs66qj5RbSNsFpxfsc+HGJciRCtqyFrivmsvfhJSraz+ZSMdI
oCcLyn05O/m1ykNSsGlOtwgneChN9RyQ2R2f5OTWxSVJob/v239i+4G2LqBqzwNAAVnTNu1m11WS
wZOnWtXtnpuvUNa6OgIGheZ+Upxi3l9jqc1l62FaCawc8l0x8ip90nCNfdZHkecPNtJKfKor9Ref
Fcr/pv7aMVucR2gI6enjdjnswuP1Y2wg351i+x4QZBZkTmzaqIFenNP7tXSilyCT1ag08G1Ed3mH
4GeeI4qnJKTvhJ53yPHAqK2eLdRO8dtdNxtsBMkI+OUAzA9x9XkBQKZS2Faz6AYDo0E+YFeahIL3
/4girYJL/NweAksU4tT/NkDwyEfrWyxDuRz+Ju7B3kw9j6dEfWoC40Zi4hX4a79zSlnDCES52Tt1
VYqnf2a+sMgClMAhTap16js6Am8ARCbTg4pYK7QCVhc25a8HYbHmeldgbW1BsRdvXxTjUZQWnYe5
uyjOn8idLmLr1GTSMNhXYCtIYQ8xOLW5zpkpO4L5iIaNQWCWJAk1XWnQyn86o+GzM4BgX1Awf7nP
QLOjdQFFjtRgSXYrOqddxWlQSr3IWUGrYLuBfHqak4r+mZa14FC4n7MYHTXAcMSpi8LRKVRQ7adh
wR4KIuyGAsz9zIzqkiNEcK99cWMI6cvgGbgUqD99mAe97EgfSw2HytysPIAa6ItutjLqf60Bd+5t
HA4hsuRaAjyH3O7+IOhzhI2MF/EzTmcQtDgIMeRkrYZauqhCHXs1eT1a42BupZFpf+dQK3TSP/Hl
cDwGWmGqH1e9fT9xT6EW4tlnxlUpS0lpvx3QZqKS370hkkGqIVCXdjhoszrUydlDEeDFcwJaJBeD
mbqCpdwSbmk4B3GP09zyKE4mT9DLT7TBzV5Gr29b+asDeXdKxJ3cP66dJx7SWRBE2saYp3B6YWCm
5dVrGReM44kKOMPaJSODLqBK/7RXpjzOwjOZofIkL6y1Km95llxbeyaaFrrK0AoONRxfZmmxt1n5
cmLPlbglJmyxfYbtkTtyA8qHRfMrWnq/4mukrX0B3LE9syb7H1JThjReuHVqtw6WHRowiiyw54w8
g/J9GBY1SV9A5aieSlEFZq6cY8oJubFYeagtTwu9fuyGNMxwZiZmXbCTvVafsmtjT9mmys7BPkwT
4S03/3xYq2Ad+O45Vl2v8a3eRpMdcJW5ByJ7YVvuBgKjR6rYBI5opKqzQkd5NR1lfnN3HMeiqvnw
dRxV6Gva3V9eC/5zpaOKyc8K41/aXqUiyHUOPkLKrBUv17lci1AiI72YTPa8vOkDfIdlhb9fMCCL
Lx+JfGJKm+y7Wy+dY2dTAa1emwe3+VrA2FcxfWq8CJou/r9XhkhgThcpicljn24O2Scl8+jGocUA
gr8bkZ0A4W2xG0iP0vMbusGZxUQ7c6QTxuALQehexvoiBNUa9ZgCvlRHlatoYYxga0r4CAzjc0YH
D3EMV+5+K7y+MHftWucBpZliarR51dtGhxRhxxFP6qU5CtsFhz5uqTHGd98dNuKP8GYcOQjAt38z
Rzdu2ismKwGGGuiiraXMl0MJBoEC7GET+STlpGMsFz8HDN9OBfGh0VLAV5WFblvPlUlo4YJwI4oy
jDNxyG+2us8AFsMDIHHMgpOhXMAe/bCiupbpDLUJT6FtVz2Wc0whz2PlMrWFlfGzawa9tM+DBVcp
hbEPfrb7PcdxrxAlEBrwoW5O74O9Oc0wZ4jM3gtY9g2nEeBqyiqdxnR/yfJHmqrjal2ee+n93jls
QLn5yGpIBBalrpmOqC10PAyGlpRJRXvfuf3ngpR7HI6WIk0xKtOH1IAzkHKaBU2ctK6GJFsSwKmn
nLYdUg3oYuuaHqLl9Sud6afJjRtVntQAM/EFLU0HLn2Re+6e/bdGTw5KgdPMYkA1trFYPr/0jw2b
pJRsrxsvoI6Hy12051jOl1eGO/X4RWvYVJwlRBLTt4oR6jZDo6oVcPthj3Zqx+2Wp+HyEyhLzWVi
1seGulA6k/4V6u3IbrmTZzVa0XEXznLHCZ/kDRqMBlnfGuw7M2iOJON84OsY2JvINImADlpUiYRk
KnSSMnv5LrKUCWlPJurQBz8FPl5CODpJP2iLeYQx394mRUtcU0odt2zOnOnKlW7O8Tqb9kuPZ16+
yaDqqVtUct309k9e8V8pyMkmhKPlQBZei0YGI3fjjbnkkDwY8TnwOOxjhQEeyT8n5JowUtGaajOX
w5vOT9W2IkG24s0XSCRI9+6lOdhA55dZvoTomK9WeTCOcc2/YNiQxaZae555aqw0QSMNTrx2N4iO
I5dbSMOs13aVSKi6jDbeNMJMWWE3SxJg47D76DhGEtXPp9+d7w9GDvgiLYrsZ3XOUDoRuhz+JhIB
FdCqtVf/V7acQYmEXrc93RkzpKdZavYf2ekw+njV9jZNsa/hw18P29kwMOIKIxO27T2oh82z7qyM
/DDS8NY94HhuFj5CQSVmwA2xA6p8VejVaBz7i4nG6QWGyjSU1ZENZQMbhH+dI6sckMbr/8WpZ8zn
bUlDIund/u2DPQIFVety1qkm5qcf2ilgyawtxU227hcjgHktgTaUYWUn6vgeNbqBkWROFWIntXGM
uQl9rrY2mspA2zUD7/6J+6TfR6CvTv3ZsovuzemgMgARYmvX9B6HxU/Wy8oTgTsLjUfMMSCSdE+e
mJuwk1YeutiIxvWfbjGleuThLwmRsdpItc/llc3zOrr78+AfMCmHjrtySMmhyGvajzttkHL7Dc+H
po8zEagjRDJZB7AvOKMLM3zYH6w6r98zH4YhYBkZpXCUfmFXRaphEshHpwKHHwTN7LSG7roE1F3u
cmq4ZgN00ixCGvuTqMPOi0QGyYSY1ik4EJ5AVmMCaG5pLvI1+ES2g+H/XGUY1VXu9I7A/B5zl0eT
ullSE2LHESD42SJa5zGjsTTeM1pb/98V8kDF7delf5JkuDbSdgRepPBINhizPoStuZ1ZlDAmTLto
4dDdMnt+6dBm3aNRytUkSK/d8zV1/CKQOZ6PJ/Yin82/NA44TT8ltVH8F0EqAsvDZ9laq24RiwX3
2RSPHi/khwXvYt1DM9YxozIZVfDugLQW8h9stm0193pUvNFyzDkwCd/Yfqyde8EuHabgMfIhOa/T
cpkYay8S33hJSx+mLabCCZfr/J5Zukd05QQMfeIBVCV01smHdb5pV+IkpXeC2wMroM8+9AWJOviS
7chq/B20LhwDraZBdAin16WDd3Jl25wvmU4KY0LOo/f/q7jZinNOim5wkeCl2Qce2H0HVAnDyZM0
pnn65BRZg5Nh9qOR8vp4N9p1pdlONcsJ2sRKwoSkoR22gF0iGspUzgIpnM51tT2NT7trwaM/gZX7
RhVzCTSJtDjGGl3z6qgNLgRAMucKnJotvL0EJ8ajPX9Pntq3/CzGzxUfy9SR2O2NvY3Q7+IkFkE4
uhOmsnLIihodrORn6OWTUIK2y4wsslCjS/XB5tPGVjdpGeOr0Q6WtDgcDslTM9YjUP+L7cz59fCE
co++GW8Xzmk+80l6iK4GdPhq4lHAhDL13gt3c4rZK7Cj4vwoqoNIo+Z9mhCKR+NZ6truzWRXjGZk
DATQQmBK+nqWBAavo5Y9VZqSXHWobRIE2npFI7uE9MkA0+YhGVp/8fepJSnLeq8Pj8rNVrZt0SJc
wlmY192fRSQJcwCHsf3d1O9GsjCWTCmUSUhdgz870WTIxmAd+goDsPCcf8iLg8QRTSsQ+/yJIQY0
yitLfE2nJwYK+BePun/QnGMrUjXnhDTX6+xgErmL6t6I6US1eUWmYqtJmwoecxMRqGsmQVwEu47A
a3Uf1AgNAxWA7c3CpV2DKTiwyCAi0iJJ9/mnbuSc4PJe5XDveXD8vJkcKsK43bEXch6Sy4uM8H01
fOsGIcEPcw3IUxGrmDrWtnZ88zKuIzmTc6K58OlfzeN6RIC5EVIhjAGBHsLpENSh4latdugiF9Qu
AGcporR2Cf0nfT94Rqfg1aDW5HpBXZpJ2XdVATQbFLG+Y4clfJRIT2kxLttVQvoYzmVfg2JWvfQX
cSngmC3xqGK/Ar9ZXRSFnFQIR1YrcmTZxIcXu9/WFu1XG6PUSjHIfj1Q4YnnNhIdyeh3MLDf6sJV
GEhxo56wpNN2ap0+lHu1S6x5ENXf1hl1HNWF+I5eRRTYN9HoHkIIdHTQDZi8WObZjzlizdXbF7Tg
Zm93zbwQCu59yHaq9zWfMOJCjd8KvENyCcBGzj/c5h5l0q1gbjv9THAwbLE9Q+mByCogt+yOLvHO
o+UoeLApjX9Bpj7sokYugqDVqnGKh9fJi049QBcwRDfLI6G/noai+F4ieU8+2fBo45RIndc7r4Ib
qTfU/RAJcRYQ0FEBUveWSG5g68MAH4Rc+qyYJaSkt6ALmCCf+61RyBF5ldwI1Z7OQNhOZq4qyuMm
ZPImYrfrtbUOgkuz+GeE8tDf6h1RjDeexfPTA4r2sEwPp3HbFs1iNGBPZRz39AsBCoQmZG4RNyvg
D2ydZzsZADUT83ydiHmSBpl9zpy0VCT/Nu6Ch8AiN7J2XyuZXMoU0jai3caoker3PPMKhZWJSBzt
PZuyKldl6GSKbW+zyt5aVEjYuZwokukyYg/IskQiBooAyvVmnCQDGGrjT/OJmN/BmwaHti9lt/iO
frwGAplQ3CNnRLT/bmV9Uor/kztzfnQLhV6xDvLVXlCANp1H1znsf54pKPDAbbNA9++xUfnBf5+1
IvlcUXPlAJe+AlIBGkrj2sRD8n6ze4+DAGMWA2stAUzRP9YkEwfYimrS2hFE5xc97wkfv6FTkB+Y
326XhwCqH/A5OzUFUaRd+7kpnV8mEXGG6j+umFqcM+tBI5k5PnpYbENzD28HB9IMIffq+vWl4EqL
I6ldCWVDva05yHBjI+ilBzVkQ98xvB2IunrWsCACPspIBO4r9ZolsVIDaC60FSFBrtjiH7EKLda8
PT0h1K8YJhwGLHNgYUAKkpcbbjW346M/Zk6UxJ/NoshWPxLV24gCb4gnE4wJGA80ULuH23aeeGcS
OV8PKapJ3UKnFtON7ktT3X/w3ipvPHAj7C+1ooUIjuk/IMlTa3iZstTsvZOgzXO+OP/8/z3RqalE
2bo+vu9yWWPdRppRZ5qLqbl/7T69BSfQHUPycyrfvx/8ObIGD12ABThxtXtOwwWEoo8z1V3CF1vQ
0AEmTEgjx8Lux/FugjGcZdz/r5yLUG8WPVLlIWcCGKFjeXufRnTm1G7QxXT3FMOHlH90SvI/hLf5
PqOXE5bimp8SNijuX2tn2DOGMm7IoRXBQIdyQT9XaF6riUkJgPaQ2037OwrA8bHazJwbj27GmdvU
UPnJSv8g62E5d5aP7d2jsT9uIQjeWbgDy9l0Yp66sCE44bbKPt2kuuKdrwHSzfXNER5w7DyXlqKp
XRgVQl4AhR2Yzs9/ixlJSfma3PEGCxoOGw6BGeL5O/U3jviVU/clphKuYMcYp3fXh1Y5Ap8NsBT/
oP7t4401p1V4iQu7pvd3ettT9/Hd0dYOetghm2Cu6mudOu84YTR0fArjA77IqiDo6i7SaBxG+92d
ve0jGeAy+WjU+gIZ6ykxL4XUstIJ5e9vZauFo2db+K4JImNwoBbqdh6VLd/mPUxwKhPByzIUAj94
YzwCra7QsQ2GFu/dZLb6rkcBjSMPxzYGZh45SVC6ywe9VOCVyXDXIDEHJlNMvz9kwfrMzWycPzTo
RhLcwZ9G70mm2rHJ/9RdnW/roKKL90abJDlZYPx+CufSdPiy5z7mTejj9byKjE7u5dDSPGjir8e8
9qxJYPFbBP+HwEKJnPrpLnrxTlR/td2qcsxioPZ506H/FAdtSbOWbAtY8CVyyMI8xJ+Kjw5QFrDL
bUfws9LhNRLVjcg/0UE/zUdV2g1Xxp9lKn1d28leS/N8AgOpVbNwSOq3+kIDAW9usKyb51zv56ra
mWS8/q5yLZR/JPD6pY04/0DktQeoS0y6KlPLPVnqt4Y0TGNQYUf3/BGXp+UBbB3SpifCUghASQdA
4+m60HS4P/n6s2gcAy5coHKXjsc0rgvuLjXbXwrvKu86/p2kIDGwFL/wBD3YYLcwZ+NmiPvEJx8/
UPx/qneeR38IKVypTxMEBIK14/IWaV4QJLUwwTwXDLpwBJiHpT13OUxyoPk/tugL9LXrlR66hKi6
n/z6gsuhqkAPMC994XsuBbtShCE/vp/0XffziJ68uiLwKKLSZYlp3PwrMw7aLgNxqcd+opq4+XdO
+yL79fFLwwKu/xcbSjrPSCz7Mg/4+02KBC0XD/kktAi3cfEJ8iprALtp4CQW2wZ+S8EMW4bG6Uj7
iRp/+8uL1frqZiB2JQ6nffBuFnRhxygaHUx7dVychNA+iuJy20lZLY7kifFZB2bRkjxdQnxrJzst
wcuzXDdv/J0AGp7RhmNN7vyj7uCLPFsgCX+Eyttf6vuMZ5lyjaRlqSCLftglsEzDMch8tf+HBJk6
/OHl94w0/n+4kURjq0lNtNl10xrcXsx3VK917fDfbphdoVmTXpY3Ud5w4IDp6b2u/fqbuHQWo6R5
gdKrF/r8qSGD3XdERWCQKofRwv8jCUazM6Wyk/74fCsFRjo8rAYRcHImZRt3ulh2QYBTMDIgj0vB
ETiaMVRwrT9IuTpDReVeLy65N0SBqwdJIC5I4T1oUdCdcTxyBlvDWi5omufuP/ELW4vO1L2XVIzi
Zkw9CYdAv1wQDx2aGTcOSfhqHHmDG6kniDb7COIVl1AKUkDtuJybAHSbZ/u/7nJpiNPT7cFrilYA
xQw9NiH1ChzwWnDhnIw+m2iTS/UF6Xb0yfdBlWpWw7KIliM+9OzcH/ZGO5LmD0n3jIuQKfQg6LVQ
DKYTwqeuYy6jv+S+kXxefTR5quiHsVtYtayJWqYwOIKkbaAfJ+iAQv8sVr7CtoGmuMEPanf1kZfn
0+rUNfyFX686+ClFdOFi5JjpiLdKEXLnJ5U93D4m0gld8eXBuVel8XjKWr8NYRYGnf2MGKkdNRCM
ylOv0EiMGHmAqB9rVglQx2uKbrUT5mnvKvrEqiMu0Pot4eNZpKam7BvdLzrXjmkwh+mhrGd7C85X
KXCymfbVKTis+0y/x9USr8YIIhXowAGD6DQLm/jLmmmTPlpv0PmG4HHEE6UADlqfHqHM9NUa5Sru
Ih5XkgmSOsShMtys6YnN//hfs+Fbxf7ExH5RB1kGJu7+k2/BsBDOkPy2eQqIA4qUIoiYjy9zCPw8
ujbKxYyRaURGE37ZgonxQMs+0UbA8UxP6YQ29hxWTVQFnWUowk1sZq0S/IQra2O8U7FihjBsLmtu
a5ARQ7tKTcGmB2kmiNGcxC2vbF+ZgZD7vkU1BNPoJG+OgKS5Iz5/8Li/EsRr+LM3SWFdGYxf8MSG
5D463GpuXIimfOph1xMkkiAAUW/Jb4mbc3D2a+99JxJQCAvbR1SCt8NdLg9VKmL/CIlPZJl6TF7v
dF82ZxJIeDeraLJGPdbRqt34rVWBNOCLRnVwLD7JGMBv2XpHyqdAWt9O/tsXXbVTVqeFxw7oa1Kc
CMU1xdnHqVOnzYDtm/UbEZNbg1/CscBgQNGhL+bx64wL9XDCJjLxrglPVpW0yrysOVwrNf2W+kFF
kx1WNjOfspph49Z2DnWpOFGijDil7BPhFDre3fGst0KsSvFANSxaa0sktRci/4qwgbHjCZW9WrbQ
kcd6kYXKnWU456tXatjPwir6U/lhQfCgXs0O52MnFna8AbSasIBCtAaSmaaZvJ22Y4dNEu9feh3m
h3ZjGgjS7yXDTM7ycmazkblwG9ErycLYtd97iI0WABVH6yOYofODIQMaafbsGo3qw0XgrAaN9ZNL
Up1HT2GF8ySLbNu2QSQSFQEYby9BYrgrSrDVLGZ0DVTypXGE6KaYriUQYLE/LHk7Hl+582AaYXVc
CTTo7hSSb11aHHu7PmX/Pfss5fISxT9jICe+0ILSThBN9FdrOP/6E6Hpr2dPRrUBXq9DOvrANNE3
WrQBXmmEg3KTpUzMojLFcxlJfS49VgGqAZ5kosB+Eh0WhQ0aE6WoURNdzfLu2fdpOL77CsrUIaYt
NpHLgHhEveAjuHlJDzaGxJUBeOv5Bl8jBAh7Em+TRFr2iDD9NgiZg4xznboLJefwgeDA3zBOQVnU
lsgqPwivR4swUmR3mN3+xcgr4cfYSTfy9GUI9fyt9f+nWzc5twsXMTFh7+3BkUakCBt5bVfWXxPy
o8tPkdhaZBqw+F3NSL3bNbOO2y6SMSI+uL0YWLBIh5Zc30/ixc5TP3y1ViYQSnluZG09v7TuUoC5
CYova3TDWpjijx9owQqzQhVf2jGu5ogOBaGLsxerOlF6WPuogmNih4W4FWOLE5ERTFmrwV+RsbR9
BjZFmvBS3sVDQanB81nrXdQkpcEvQ228W4haShFX2JVpqXyyKWaR2AEMcq0G8AFxCDzNX6A9z1Dk
eGZdZbf1z/HKpe5XGbWbQVPeQgw9Ra8h9eJ2Ewl0q6g2/dUwGvoMhScuYJ+NwnJDzIsRckpaYlWZ
5XJ5jV02doHv8KyUyh2r3l2VIEFfN1/L+C6owyBlBLkOIbuC09Xvz57lx1kWUULjX9o48rnAkWos
+dKrWJyfFQS/OMl8rqP4u42q+zBbDvF3+e4//Rt8Rc5F2ZnMuR2JG9zOa/PlFOCWjwuqDiMEkozT
CG5Nnb5+01XD/sbWe/DQedNd6YlKfvV4DzWhIUzshUIsgKgjlGBtdf20DWRLQD7B0BW348rrXjz1
P92+ODaGef8vTooEjSQY/I3M05SXOGYjxF1aFpPQDucsghLUVJPb9nBo1nOfi/j6ONQugNc95+G9
1JRQwjDSrkwmRLZxnHO9VHZrw7wIGv2POKr4VtI1t+FVn3K5qtN4uQGMXXfmGSjG4MFvV0znL3ct
77R+XI0YpvNXRHV/aVaplP8tfVkNDcrJDxrleCUgDl0l0MquyqzKzybc63cgS/TIWDTIIPbW2OsB
Dv0XzoGsnecDYG/ztJUJJzS99Zbt7YpROVTobGDIybTWM8UZtOzgTT9+Bs3EERAuFML2oCgudpsf
zE/8yw79VuL4xJzT8mPbt2+7RRqcyNCZxEB595LHua6iXHdrbvKua4lIXHtxUJP6nhXCLqYb1CGQ
nCMCrV+dfNun/lMQpaw0KslOOmohX9X8j8JyIYMGgiGN8bonOJ3+I9Ki9viUTbYb095zZkIM9zOi
UOCd0NZJqJgjcFt4A5Yo0hyoe7kZlLJtg6imhzWHY97/MGO4+Abx84MhDWotFpBBUqraStTNB3wb
y3z7vt8oN6jGx6StmCsXOPcpyToBLmoGP/ottN58iq547selHGRHbNBHmRud9Bm93Mbu8+0RM6RF
zIy8cQGtScU9Vv5eQFQqTncimHA81tuB6jZ85jh1svKu3sDZACVkE1S1cjpgbiUXBZ9FaHeUB483
57Hr+1T+4RYf2Xtayd/1v3POTnJgRrJ2qjsqrfVFsJtUHkCBm5yg4uOntejOiUuyLKLHpznSGvfk
C6v+ygdDLY6zEXceHxs2OeFOufCZtD/1bd0gt6TuzLt9Rq+9O9QC7pjn52gvLgA7TLTkkc64NQOz
abDUoiuvNgIoUE9Ctej1t03bEJgVAj+Jy4l8zmhQgnBBvgHY8pPSCVQeWlD4cdI748mH4nY86866
oR8HjU8cYPmuTjmnP9Tc7PDBxkuCT+ah9YdFH/Grjx+MsYWVcymCPki2Pbtb4jG4ePbmC3525GbS
MO4vZWYdUqoeuU2estvlT0ZMza+eP4c1m1Nr1NM8W8SpVFc2MYd9vb/ry+t2GNN5qEXSi9ntjwVm
V/wIFCBzDUMxwS0tgDvG4h/aXqS+rH/NaAXQCycL+asqqVQF+B2GksXnkXop8IsymT1YymybpyXH
sbgfXAOM5Zg7pQ1sBQBWVIL8oTFQ3NWCj66tA0hZ3D46MHYxx25yi7t7k24M91Ex9G9ysrUBuCnd
z06LMVgjBJ8sNrq7IlH3+zLiSeJXywnLn3yGB9m37Y2kQyldAkuUdU1AVf3a8BSbxp35YL/F/4Wl
RuEAFNyie4O0OB/tbsDk1tua5kM6zOVRE5ahc2quYTLduRSAejUVR3hu+JfenGn7SnwbHJZU+13Y
ilVPm+DOUeyUm2DS/35VtB9gPA5iEtsoB5EtDX5hHiqb4AX8+yvyWhJCF37meeWLr4pxvphJitXK
PLyRov63HddXAVRjknkT+10d02TubcZNTClXan2GlpZvtK0HGIobX7Nrk1szML7aI14J0gcAWUyw
85nXttOqSj8u9LZOWm3Ue4j9liLdtqzMQcboJmg1J0VFqKyBkPuVZw0EUyTvK1zda1Ufj+ma8vr4
gb8vuaUNMDp6HfUFTmnzk8xBx8/Rc0inoCLnPX8ZWLLeVt6LNNUb/t6VYs7ob6NnccGc7InhJRK3
NIdUUrkbJpyp5pvxF7zhsLwgrWCBsDB43umYuP0j/xKMBqEYBeVtLzTL1N0jOz60a2Er3Q6SCiY2
CFPDszTVY7Rc0KzRioZl24r3lD06ts/yQ1R2YgGyQPCrPfvdR+Rnq7DySPFhIANdgaitkdHIFcoe
nnFMLPj0pOXPc/TzGQlVggQzs+hyJbF3LDoEzYK0HW4aO2/qcs0dS/KUmQxUDZ6R1bn4wk/zXlLB
Qv96IR1snBbW9NYA9fRcOHekctOn5X/VavBYSRlaQXrgYWVEpiWwGwuri+LWYVbHwRgf/I+F8HpQ
JN5zqh2gozpWIiSJDxYH6gjel5vSjsk1YdZoIJtf7veBXWdnfXMkUDfo1OH8d1txBBgNZ21g6De2
PzrK4yrNIbX/dzv2J51RdoRHvrcwfW+T2sfm9ID8F7IgxH3QKbKPUxarw8VJUK4OaOEv1m6P+THv
Yv67CX9SsYgoKlshHpYJ0oC5QLznDdf/TAqQOh0iQXVOyjUdMgrhDyzcveqOnhyca/6oe88OT9Qg
A9DKYP2qu3OXCwo/cpLjJY6yY6ZVgfxEttcbtnsppk3urRaOnaJo++dC9AM6mfkzQHKYnNDeDema
ZBkFJE/SDIm+onbYgP/WivV3GHDaU8X8Ykj7tPuJnDX3Ppieasf9MsE3GCGPPr4U73tUkA1Bktbo
wJ3McIPd8sD07l3w1Iqv0kPZjskKIIJXWjxIYevQFoykcRp5IM2iqyYzgZvDsggO9FL8WWMXbMLk
2VeGQwS6hcfDYuz0z0qy6VDmlfcKJx9wKkl+xk9glAx0Uhv5ScoVMAYPI7HVUW/q2+InipZitinR
0R7nU6p1QUMJlTX5Ubtz/GSmTDWcUTns0OIiC8nIu55cvYvBcAWIoTj1+VfK4em8rFhYlMjnI5am
jdNBLt7zVSQStMV+huT0rarYB32LdJtqYdwckekh+bYzpfUWlrrhEt6nrR5NdPBYwrtHKCH+3HXL
hROPF6gXGH5kPuL3IOSVBOqf0d6Gi1XSTnwbKnnPEXbP12skTWuNo3vaJuvAesdctT2XhCmz+FPM
Cv8DHH3MOV9/op8uCsncigkDtvHTKmnnRoNw+QPr0B6drKjPz496ZdUv1HuxIt+i4fu8YFEEfDIg
9W/PFFL62Ih1pLEzAUslGRWYoW2rxyszFbvHC2MNESw1JVFHRCtkRmoWyA+ey61WgL7rAuBp3uQ2
FtZ7iTRj1/Ki/oo40BKdXIWCjgChzZOfwg83R/NZCUcX1sAfq89Mv1ylXNrMhBLSTp/TMtK/Y/3n
ZzA3ZSI2LJU1X/AtWqCfosX4KYzagDKa3S+XekLoUoSoyPfLORkLkHFQNapRNr6MZETeILu2JmeH
bqwzXHfU7H3NHU7eAtRDqZuixqHS+IjlNongLQeoBqrMzEmvS051Q4aHtnwhFRg5ltLm0ABVxQ9B
io9+ixRqz4SZQ8hLRFgD3QvNurf3ZGxoo0upvBXp9DLG0U5s40Vx8bS5mRAulbCP1cvT73Fwi4Ud
CIKYSUQCVdfteuFezSoO69YeaAInEHdNPWZXG3gPizeagyOt2lkIIeJgaO6u762FUno3qf0SNiJx
lKG1RtFygrljQotE7YB7I17olfe6/NQ3A2txc0Hkri2kBTKIQAH9UE57N6HZQH075SYDIEe8DCko
4mxm3i6O66ihhjAbYaMOAXgXLWN+/nCvZSt8DV/ELTlckr2MmFW9q6NAAk1d0OWWHJ5R7GGNrnWs
y6VZvWE377vUBhBMJK2yw4qZCYA7dbLUrYaVBuTOwVF/fEx1rftB0f2I8QrTh7H/d75MtCSuI4n5
OG97psfO8bc5z0IDdwMjEzYV1PEOTAnWj6DI6HSNH/Gx5ef1p+d/IY4p2BNWXrgppCh+nOrtvqba
Wg+jh1vcM7XhoH6WQDnn5tvLHVU/WVOGpJPks7LSOL7o7MTfcFsAtkW9w7rSFeGQYAM61le2V122
7Qj2lRXNoxIhz37YagxdomXzxDE+RchFgojaf+W7WIIZeg1nGWYcAAbgb8mrFcXA4kt4yDfJLpoH
Dk81sdMRUTc65WcwNxxiBUFYk89gv16S9XfSn3DaG0jCjWbwj6hXDQ8X2LEEJq+g9PQE0L1z/UCH
qj8sXdn+4vXe9HEayKFvrivVrq4xn61vzs2JQCeheTbq50fwwr3E3Y5xnTdnOSEMWDR6gg8871pe
ap/g/S0TspN2gelExmij1owJ+iwbDcOkAIy2zl6pPrHt9hSp8oCjr3AWgawLg5m1+1LyFBWLuuI/
V/49dG5sCuhoU99AV3c82VpVw9XUcYFGGNbHbKS7t6ftsSprPS97vi/rrvnHs+lBTqGKKrkvEnFl
Zw/16hDZr3HY0H9kjh99of5ejKy3l9Q3N+8eb/Fo2wSN5CoPKA41ckYP7J0ld2xdIOKujZezWEGr
yqnb5BDHEw2/r4FMueCAnyA3EyOY4RHfCQmeYFVY/MaVKK78YfdhbqDKhUsqmYCLR7qWzepZmPI7
7JdjxOFm17ddOunsQnNsm6OEI0uFVMo989qW2b5ko0KWFofehd0LToPWEBYeMepdQUalW2sSm8FD
YAoiyYMQkYJTMPI4+t46mIPU++4OYHmV8/wHaLgYJQ7HSfy97BZlW8qiJ5K71Z3j4e2A1+7wsYym
vY+eQOyR4O1sNCMRTSCyusK1lTPpmquKDIje96bJ5g3Tw03ZpiFhSTs+w9DLUTuINLVD8w/dIAz2
eLzggbRLqtOfH8oOChSmwRdhRE04saQCVJDJPKs4iaoOcXS+uSOYNCPpcNLJBXwYthvnX5saoJFm
dF7gqsRcp8r7BdMVItxWKfOmLvYUEMUhSYXXLCyfe5Gme/m1ms6u11NIe3KDCBErrEePc68nsi07
Dvr4jYTjXl0YtSOE+YFZsfDGmb8a87giUUffLCy8q3+evyrI4wKuFTcvYrbRSrhScKJVe2B4o154
Xvw+sSsDBn7ITgMVbUgkvl4PMI72W79oSX5LuYn55Ib9A8JyN3FDtNKCAn8iv0DcA378mYxO2pBP
jbzhwZ8EvGy4ZlX5o/vZkwFXkNeSLgsD3NaHqIdhGMTfNjEQ0RqtwjH9cXGhh/D2c54hwFvW2xRp
Z/moPNJABnt0u4fYp43YXHl9oKdV0QbyYaT5SMH9sApbfte6GbK39kxgaz6YpETeAnh3JVnobWaw
rZeo8/ldDSo/klpNnNol2E//CbQHYrv52dow4VJ3AIk+m6KAr7nfG7JLHdqD57YDIpnM0018k30x
WqJRxwmQJmhSwSsfRa7Ljtx/esN2/yV08nHG1daeeyoTM9Q1JWS2tjFHwYu2SqdHff1I8VaKeLsZ
luF1SWyeJRHMK0xXaOJM/apfoTGJD7TU4WpLSmYl1qZdZLx5MGLhLNKB7aDLYZT1lY8DTnnkizRg
rUcHvIu2HcIH/H5z8cOayvtoPWbPLC8DhbrUZEENrXopjH9P5lnxjOa8AzFTK+dO0dzZn51VYR5A
PGXGp7dnKQe7il1l3OE6jfyNfyTw+LZE1FlGzDqaKA4FI/GTmdfxNlGpIo/zgo9CYfVT+rH///da
5R8D77Pz1er58QCl8lwti5lIwu1m7KMfLA/KQ41+DX3as/yXuxbzplpLRFtC4ziNwpISZTwU0/A5
512I3HVJATQ6Vd9LYsUY3niuFlY2mjPWXuo6H9lZsUtKNTk4RkZYDz3Id5lGj5KdLurQkrScO4/I
yILy+pQ2jHeuns0NO+FAKvamNHjghuIhYchqDr0yjDBxkQYsrsTKFYfxN9QQe1kOWfJs6QtrBYkN
ZSqRlAA7b8RhG/6G9S3A8ZPL+w2Up2tA6YmHCzEex9oaCKIPXta4VBKBnLu7EMoUVQUVpkxlvb8c
ihbXEeMBao+1BO58kfrn7Gh1Oe7wcgViYZvgv562BI7UcsO010583DRU7Ww8Wp9CBqXm8DFqEmrZ
85U6Sd8CFtj8JFE2wrJ7ygc/tQ0P4OV+QcsLlp4L7KvEjHxHUTAcab4v7XN+ApQS/fEUfgvwHVl9
THhfFWYEDDTRMzMYNEUyS/Fpx4WvqMj4YrznrIqXi0v1N71LgHbVE3oMdSrmOusG5u5WIGjxgz1C
WL2H2ygZsKZwCVTdydUqYh4SO/BfS5WfLcmL3Z+0phY0A8DyZ5AW8vgIswWGhVlMLLl0SWzSflPl
3S+dTtPyMDDII+I2p9jNZ4FUVjt9jgK7coULMhtepZw9Kkobc1MkFW2HDiRXoS5LmAxljDTpKmTB
xiDOm7IRUi7Xh65XNArnJvcpmcI45yd4f38s5JpayX4NfJwtfy56fz3ekEWFaaN1+Rhd8u/Sg+Tv
/PCBBLrc5ijQVJXbDd6nGCshVLWK1nTjtZX/RtMP3uLCXAymP+ju6yfU0xBMTNOIxOashWc+w/dh
cauL8PTXEcW+ND6Uq9CxA59JkM4DV+iY865cliu6IKI1gXsOSBdqYhb1tpJcytIU3pu5GQJf4xI2
r6Ii83N31oUkVhUo2+EnoanB2MKUjKNkedV3wsFp56beZnZdg9XyNhadMFEkssRrjRgUgLQ40SVO
GysfAp1WooUYa2pbvR+xHuT5x33U419kzm+BQnRuvniiqj4EeU8jjNED5D0KLv92VyCyr1MSmn9N
u2Nv7jErqqd5z6bW/KAu5UtiJypqK8mVAGMac4oNXH6QACePmg3eOT8bb2s5kmbT+SPYpXxpbWnl
2/2CC02iBWNM3meTClt27qZrskMFBPfCpWh8ypexw5PBHbK0N3pVoNyX8XTVpoHm2u7ZgP6c3in2
C4PMswDJ+/BDOWfkeVaf1uLDXXWYRZSiI2MwT2Spy8KVUXPntlJBk4QJN242eUevUYcPYW/WMGFg
ngto6RElip0obdId4diQMJIS2UHkwXVwRCMmKmWZpLvB+BkUt8u4+J9ZBuT9y/guLY8LlYIk+lEY
Xde3YNhW6EB0Z+m7l2p9pbmU3QlInojUBytsLh3cbsKQmWpw7w21P+j2MOM5/k4F+6yvUBdy5k3i
qluMBFegDn9f8tw4D72O1yIbydWRupXU2Lt/fAMFhkbO+toG8/C36v/iwq77E2prLdE4UPy06ylm
du+OqN7zuXnvivpU28TZ80LD2nxpgmVnSzUQLDGn+QmYm4bNiT3TSVcQ2NF7ybFe7pIsxFvHyn+K
HWW3JuYxJqsbZGJk9YWMk21EtybIH+1yV3whRtByOgf+bHoieGGKAfHVWUxl5miQ7NJQHPbOIiwR
xvO6P+lHa2ai7kHa/2M/nGq+/wK2Z65V3CDrGMcZTHArF4yOGTqFL9bCEmtUBun0hX3Jl6rcWF/s
6G6p/CYn4+fmxrkHnFwZyi3lHPbIMe97A5HfnVEvj4xN0MxsIhMNr0bvd5M3hDt9jb5BXcPvDqZu
337jgizgSR5O2yXHxbL4vQPnp5UD5A9S3QnlclDDq0khyt1pAY8jhKg4CCq30lUZYFk/LjUbFKRh
/+ikdubItEN/A1DmF16SAeV8MBooUlXvMPbf2TDeXi336zxMFk2apbPZnlgW5KQyuDf5kBjr+8AC
Md+L6L7mMwc8HMt4u3eV/NS+y8sxN48hdixgeNuu/6Th40SQCDZsd1HKaneEu1GZDqVxAkhZCEDm
Doz/uZDsFSqHbAAL0/fzDkPgejCrew6BFrJcUhzzdOGmvOCHLp/+xNWPZBezDtMtYfYuGUcpTKqi
rdr7YcEj4lxBd4hi/OgHQONs2IzjTM9M5Bu4BHQZt5TXG0/+B5VGxGKBxkkffa6oalrxcyVsmSzx
bUY0r/H39pXFxOmQ3AvgDm63IUX4askaMBRX1xjZnte1+kZQfTCpG+7phQ1G3y8tevalAfQmMdSX
fQFFKzOw9ZD0vhAa5W0jy+qc0c/1Gc4su3r2tHrJBFmDBC8dLxeu5oCpyIuaFI1+A6NMNVANzz5i
uJRVkLYAzLxSqFubOhjySLDS5g18fbNgJveQzuWevn0pA9TVKm1vQ+p6bM5zZlRlQvB0XDnGCqdE
LcM9G2C0N3pQoLllExT0J1NPMxRcR6dSJnOr3v8WIJO/xKWQJKeXH9dV4wDww0fSAiLgv44bASVU
ohA/X6NPMl+NpXQobClpZ5i7ihVWzo2Sjp3ee03ovN1Jv3/mZtkoiWYdowSuKCLarwVF1Qz84pVS
9XFLwkrv67b/xvdLxZmTT+BBGZiqkCKTKK3t8BZaCnK0LvN5muVYFADpQez1OROZRhX5srYdK+bo
pSKVMfDGhVtaPoOGe2Ci82wDsd0yPMfWMlokhXLDKh27BJdJi5Ln06OMkuzDAfZsRIR4e1x9YNBm
42HAbopGK3CCFmooseEcZ69mSOXSvaAws7gUQ8H9+KBOr/vDOOaPYfda9SPwZihE5tMaOW7P6oeP
gIyUCEmOm9MPuR9uGDEXfyZen7jP88/3YVmHKwc/SapXWmtN9K3D6qdnp+SwnKlIFEbKscFKBDka
ybaLCSqaqlmAJ8jvZH91oPa/LWMOBOKtWlyaPuCM+WGYN4/BVW7Z/TudR5gMQFC4Nu4rarYLslyz
Ukejkco4c7mpUiG0XPPYuhAYoFCo6C+cPnnYsXbkbTKhQxnb9QpxJnQxpyHSAVjvZUFRLAKHaX0/
O4XtvkJoJos5WlXNe6TG7sNlr+EMf9z26c/L73aGg7y6Tm/IXTnkcCO59+MNGAGHleFZL11HSwK0
82uE9cUjbzX+60wkMiX8gDxny3H9yhoiH4thGGZiPUV/3vs2llfVCM6pqSiIkUjbRI27t7zXWpnq
gL0rDhML8alM3kYGqkLv2LUaT8Ra70+Hx0q0XGRVNP0JZlPdlYf6a/bviZm/Ta5AW8bBM+7ee35D
ZsbXrLDgYVo/7sojxD+ubUIum8g0A1Vo+ynGyVz9yDheR7ux01HsHP01pdggHTTi4vNMWnOkowaw
ToXTRQZaAMCV4hyKySD8FG1NiP9YCZbhtU0FjdF5hF8sqTlO0ch8z/L76TzOk6+iLqnjm3XItDrC
PJQAlFLP5lNfXvkhh9KUM9VbMySyDvBpFn5dxKbxLqRgWa13IBRPXQ0Ze2hYD4vuvkg+SOpxn09u
nQ5GhdfuoooNSWLpU0j+kQ6FsHaTJrdkqY9B8lds+3rw1snRowkSGgjthWWrzij1CWv2YCQ5Hm1+
wkiEm76bOlE+KEiX/V7Bc+qV31r+oPVGKFMBLI0WM6efVjB5PSVwwMbph8FV99SOPw0jI5hwCsE3
80+4GQwC6PVhBsn3n1VlCdRQXNFbGtSdiMK6ub8jDV7BnPWkbKM+2y7b/B5iCmbY8pMS6rCRNMiV
y6hw0LY5uCdOByK3zJITEp/TeHNma/VEsi+JHLg5ioqpEMjRR75KGrbz9x2gGLwIPvwhimbcRfW+
/O9DgJ1bj1VID54PLXj2Sh+s7KDz9dBrQioA5hMi6PrwEr/3Wx3kZ3u6AmZS4DjPuJtJtjoc725o
T1A2k8eARND7/JESQ4zLze8TmnvY7mSHJ95HMRTJEJ4cOqVEXeiMvaSjahBHSgjvHmXvxNm92dpS
j9QOwszYp1Y/mIYHTCrv+6FpJ9+hEvVe0xJ+4mliv7nNXg1NVNWb82S9hr4FmCiuffTw02MfmBLB
K+90dhMZQPbS9GErvjLCbAq3rUC98p0tRTk5zjOIowbc5Ewz0ckPXll1TpnGB8MbdHtIECo4NPrl
GOLD7l6JRrI5mx86M56lzhX8wMyARsofdczxeM8D7uIZCSLepyG4zfb/+jDQunUOmydnihqvWHet
8eC9e+OqOxozCJ/rh8fIfGzYF2gb40UasjR4w6TpKWSirYxsLjXZ9b6bwiciXFXS7EVr+j7cQDWu
2cf003xss3HTaVhO92zPDchFswowxCt/+JPx64DzUedvYXTTdIU+HymKf+Kw2Equ8McjDXame15r
fSHMUnBB1yLSq9aI5ZOiApD1JMkBIkrrfdZIN5mpILvqxFlbrtRZI1YB4yOPacvYgqe3LcPrHJQC
AoaBs4ZnBjVO68on2IDDBiWyMJdujUYrnLbjXBWTc2lWnunqTU5gE59HEvq9BOarBLpjyK8bY4EL
jEJEtMlxHUPLlH/7NckGn6drwwxt8X80wFX48qFELe3yQaOHvoisgmcge6YhvG6xq5d4DAzuBKrh
Spv06jxSD36ffvhZnKfDenTkyy4x02dAJNnTHhhf6dA3nsvQdQ2Y2BMF8IHkw4wwrPhgigAavUiG
ZBsNZeszDQ6eCjEi1LjHk6hSkZk6ljT9MRPVA1PSgl1LuevFtrGxGV+YsEn9liFr6/BncLo3dDUe
5V0oOOIKD1yfz43Q43nrbfuPnIZy6xjGRLJDduL5sYMEh6Ughd7GK8PPmk3zw0FlLxZVTnIIuS0a
l4LlRbYBZ+ktXQ/zzADKT1fRJETFU79d0hgvX2TLd3RB3Cu3QzDcCoVT0xDsBFRrhxYW+VWN3hhy
gxWl+S++yp5Vef1GjYkV3/K8jw2kd4wRYkgwI0ovi10MNYZzMv8FmbWjFaWbSYytc0jxAdAxshYV
SXzKl0xybUGQtOj0QD/V+gYLCVyp+8S09jFqAjN9p5urSbBN14oR/stMRMHngxLnPiW1SnOf/MRO
72ETFcTlNJoarMxCo4mKu1LWfrxq9rVRPq/0EXmlwGXeLcJDs4mdWG+Rss2AiQY/29c+BD3XuxJk
p7MzDSRnhrlx0NS7wKXXKTFZM/MD13sbJP+Jq9IIdS/zWiS0Qz0Rwg2bq1UUk8nGZFOJVjegFWSo
kFfcI8/Yrl03bT05a9JhIT5Zu5oSnc+wuI8Fa5cX1gNgVmmaQw/KO5SOigw+OLOQRd0oyHTMxCWN
PxxKwdJyruY6HC64HQ2OLp9TUDgYYUdKSkLOqfdw34Jp/B8joXmPdD4ICqUlXMmZLp3inOJDm8oX
DdiYFmOxJfTta+wAIHTOqnEXRl3dBAGxp/Zi3s793JdMM161EV3dNd4gNd9dsw2kBfLqeCDYU03A
aD3EZ0wzn5umVDpXYE6F52fJ7dHx7I3lrS7xRqp1drp423HAjLeAL/YlsF9g6qERKVI/9LmNnYoy
lBb3quBYwJFihkfLsbJQkWTsv9/OZKw2EvAy+LmTNzt/2dcKy4f6CgAMIIWS/q+Le0ilrYAKGsTx
mFgzmESfGgRFHfygdKZS1bLwAiBpEvQvvlTkZpuVN1yYVj4SlbtQqQa2/oyrSc+Jhhjv/F9bc47J
tZXfnQJTTB3CroYHGM3zLAolAI1nygsQPpbKNSdWzcG4DkHAK48Q6GiUbtg2VKcWwJl0O1dGgWG/
uDoblmcSqLmNJ42hYce3WGRWK2ukuO/wy2R2zgl5Z9tuqNjBMyiNvqSUnmYWka54jnq3NIOFRYb9
/phZhYr4vSRgkMdcq6qKa6uFrpsUmD4shamUicqkyCydMVpgFftgbBstoCFyNP18osR047c/fqgt
ZV75r40BMIuPIerWE9jMA41h8LQoIUcWmlMKlb5d5peUlmDcNmp1wZ1+8DBqojgH3qUPalhYnkkC
LDtCNwqRGpYQ1CquR8vtFc8oSgzKhZU5VVru+YCYqNV+PTrw3lXwzNxf8WBdUIoIMUbwn+vox/JX
GyXO7ERH00cjsnuCTnWI8+CiWQPij9YRW1/ahEjQk7awA36YMAzvAI57OXKu4DQZPsrYDwcdGr/D
yjGI4+2cMRnHcY/sozd+mdL+d1DFXrrAE8lQyYMqHWZtp03GD+DOWJBuoHOQutXlPikrzaAmlf8+
/peIB3t62+gyXcT/yXD4zf5sHWjjioCx7+nsiPbT3lU6ZWxBqrVbc2LDuHrq1zjQnTRKesyxr0wW
7uVxcvDn1k313ZO12bquqfYMTdSHdOwL0U/M8L0hQrQekiKesCpvp+f/BPXsWVHhpq7ZyN5DatOw
lFNWL1YZfqdjRjmIlO4+EpRJjj9LxncEDewUYPYRW+lsZv0FPg6pGzIUFBhqcPjtXxGvdFjogqF/
oppFi1BW6x6SQXf11beFPSRSWJ3HiGQr40gFdBx48eWlJN+S1bhxKzhWqFwJlqMr9iY5oCPG02VE
zPlu/dBqYP/x5SE7nrK3qIiNheaLmyJkq7AvpjRPJcFe9Tk7jIUjUQQnkuCLhyPQ7pfBHDwfzAFm
P7z2uBd8I2hHx1ZDryczLqpAYW9/BTuTtVDkKWkqTvT2aNSC+R6k8b1Z4W45JBK3+Rbyack0Y7cD
1YBgAWZKkZY27CV+tbu90+bvbWppE6XoHtePFbJQE5g8cmdf+1JM9Z8lVy81GymioKzipoNELJEL
7LG+8K4PE5NgHDXM+61lmmNywalehOOhS+Xi2LolSOEVNAsszwbO3pFgSPSDmgVFLA+hJiBdQ/mq
yPrYGPTo/GZzed7A67aDg23pR0XhC8jB7u/to5p4DPo7OkRIxfxz/BErAbqnssMglmbzZjN5iSsP
JeL8FyWXEcQzQGO1o0voX+0qsZD2iJQkLzAGV4qRdXJABi3OfDkm4xizXXn7NBxSMk6uq8yUHIKL
hzyAp4CQj80CZce8SRQ3N0IasotTRPBKvnRsbXVyFxWf27pFUYe3PZdqYWluH4NRhlgH/NlsGkEO
e4ou3oMmfWUMQPoJGb0iEJ27Ua99d8WBSFWmd3aSH5sX2urAZzFFgeXXbavFr2aUILuZAhBCjOQ9
V6/6IEOml03fQMedJrrzVFswAG6WpED37lGSnxlHEUqENpRwdXs76IX+kwQ/M7oeCdwnPjw+UEb0
mw2o6Gy9r+T3OW/LSOUhdpROW7cgulvXBO2IuF9vss+E38IhX64qub6ffaL+DWXIOWnyc8yM2pt5
bzTDjvMfwQAILHbTifUJXhXsrovlH6IeWtMbPXrPsvH/5ZUDNOjlDYe5djMuOjD0aF7m80M++622
Tjtah8mWN4xsZftHyw6PmweontL8C/LzpbTTlWn73wYOlKDjkPOlsE6uD2B3JN2R2XQ+5VcAS97k
a98MJBUoV2OaeoxbHDzHfZx8wpFDyy4q2DCAyQ2DblTCD6PUiGS34ishiXcowSJaDkPoDSqurTx4
kqX0zRmIKEXxQ5ZBOGBjwFCWRPoO1ylfY0wh83omplqATH0NW/JoReMa8rj2l/ZE1YIdYTf0C4WH
tC3JbPZfRFKr0dHXlB8CkqQUvennXcJRDvK+ZrKAq8zsH+rNL0Qgb3ywAaVhSXlZQI2LPOvnSblv
RxNmm+o3Z9sQNVjXmqKP81APIZdaiU5GUxOv9ekZYMVuaeZ+DKNkCuPAhiSft2IQNlE8m8wWN7gk
If28b/brdK0AdHngLrH2JWwITHukfuFi6+YL1V57e0J+iJoVvv398AjWbXmlbJWhMpbQ7hYqdSyq
W0uhLp4aqWXHogTev4W/1jproq1LkFewGNr+ehT/RM42fSLo+Dbgi/VtyJfs0rdFXH4/0Lji2/lX
LJizivzU0VeB6g8BCws8VKl67BNUuaAnyOfcAhW4bFR6EIhLMX7oAqP0NAhl2QQk7vPwQMp+F00e
exGVuyEdlEDAK9MhP9asZ+V92FUxmUQ0lPlDrWZ04qnCvW0wNDKImI55lQHEHbCCMTELA9hMD0j6
3LFuPIfChqPrZCzz4pu40ycewFGDno0ImfiJqcpyBqVqh9ZMOp3CFaj+mbCNALaaoSU2HOtOph3L
dgggSDkHvHyNbpIX2EK8Hdf+EFLIggknduhU7dLlW6OW/ADdhk+QmXnZysJvYYPd9RMZud9y3bxs
9yy1i6cbRk9+4YIyh+NrJWXXoSfTnftXp7dt6w7sGgE1x3xQeZBOsmjbs+IoPFkCx6nhbpbh08DF
DDng9tmWHgvZqrsF0jqrbC0SOTmlzs4R+UCkHaDAY75CJtFuubhWOILRD0wKHQ+TJqaxYE3Tt9WP
ofuRL/0rPv6mEx473/bFx+LXhgTRi/o0ybny/N8/tKBWS6rZdZv5MUY8sYuRTm6hwfx4FtrUGXO/
kUNArL4gR+9fj0eapIWUgL7tSauH27fyFre07XeKBBn+G954MB6xsIgLCT1ivMphVpNS57jj3HvE
8J6gJg4Z+hO77Ls2Ek0gjr3BF4AIWc62PrjMnQra2k35XRqMXmg6SqJXRhkUqBhXtMjW/tneSl7I
TBnPD2oO1oURhVe1fwtFbaVIifcb5bbsH6rZNwXBRP9Fx90E/V1OB0gXlXt05x11nZ8rpy0L3td2
JHNNcb02Iume1JKo7fn8kTpsauuEsMbaC1JcuBiyw8xcKczyYGwjszF+h/xFR16+Fe3dtUlPjqvh
7/gnxewvETK4ktzw/1pROEbaW0FWcu3NwOTJs/Zhq8WalI3ORDhxvTllXH0G62dXtcc23uyHBili
u9Obp6boUnZTLRqFxQxYhVZIXAFSJcgV/wzrvvMU9vn/i1iR76KH3iV9Aho4ZiVMYg0ALN5+taXf
rg0E1ThaPmgm2EKRPcZM5DQd0wCgK9eu9p2pTjaVabvnsYo2zycsfVEZO0xp65SZYzhgtKpub9gZ
iwF8RhgDU7SW2+/6b3snsi2fFskPWq8moqi9dV7ok9yHbtq70UBjXMDmAcflkKErt0unsYbM3bjG
VqE8VFZQi3W2lfhNETlmId4c9a9xt+/ttruyE3IE6AGDMIaBbdEm8fMX/swP0iLyXkDHSaIEwBTf
MWaNUJ5GV9RwvyaZ8lHtfmaafYkjH+d5tyabc4zT3LOlfkp6L9FJUhTewjbVodTaOsItrcM5x1gY
sfYNjxW9OViO3DsK/W+/iR/XZDg+LPaoGbvkXL4aiqKswMF8IyEPwb5rZtv5DR9tb0aEGnnIrlSv
HlfDrtQ2twQEQjqJSozMWWWPAamvpk/5CHW2l2GDjTR7zpwUy8PgBvIwkDoFyg2UgWWQpOGsLHT0
JVO4k7GQHUy723XYh4dJd9lqseGsozKMsIswjJRJDBkxo8dbodwIxLBga3xtbNMV0NXDzpGxmf/t
thxLgH7Aams3cTaniNvuyt4UocPpXhipS/QdKNOF7IXDECVAhWRW1n+NctMN+CFIStXomaW4jD6G
dEWEY0NLAAYmOTO2vmhEdTtdMjAGtvnJcYD25Li3UFyY3H0qwcAwilK732ZO+6f7DnFFh65RG3Qx
k6d6Em9ZmHdjs/22HBNJcXWaFtsYZ2gkji/bwIyUd4dm0aSc89aCSOgwoHtfeOCbVTTO2lvxQgbd
poQXlUGI8sJud2DDvMyvTKzn3omYfIfKSvQKiywXghmF1vBF0Q6G1Xg8JCvBd1ydbnCKkABYrA+Z
tTyPjGlbGTjOpV0raQiheNx+v0dEmocFFON79gSi9efjrNh9luHi8JXWITLi0f+ZvDsCAbTmImn+
ND/S+kmFnJZHusMUIb52kOq5WqIheiGnNxHAhspZ9qffwyCvXkAODQHivOm/Ax02vjqQ2wCva1zA
GvgccmAZ1/43xlFXi3Qn5Sy+96uyJpCJPDYn1Jj0i2H8Ue93HMoMrWy/0y+K+JRqx1D55ZtKTEsG
ZBD88wuUB+HAFh2k/EVeSkn+cvs4Sa0eoxsglw+jeLOK0Mny0X1APThJlNlQXts1HNEL2g1W+9UR
Y7+BG6JkmoytQeqHHmp5z/wZys/4FNp2DlPowkFawUnQjDL0Go+S7LKdOgQNJ2cDRptpKiRCAe9p
Utb8cpgcHgqDfhw/1yJOkphNc9Jhd1xz+s0HhzGOeAxEWFBGFcEl/PEnC4nQfCAksX2erHLsu5VF
StfDwg/y99nhqYceUKBU4i/EwEmxIygddSw7tPWn3LR1l2h9HJF+H+wR5pFtnJ1NaqgEfZW6kZQR
cilV621bhifEuPCzljoJQh0OKwtg2zs1RyoT5cPFtai0K2s9KgELnVp/9H/jHcSFcYLzXbMZbP6y
a4qdVZf0xgSpKJdgwcWn8kRXwQddA7I3S92ybXP/L2KscecwvwgrnrRDFUua2zki+EaSTQL78pj5
K4WBvJhhRUsA6f4JIKGLt+Ew3UjulpPPQbuGu1aFB1xF8qQ55gQ3vAyLNi4/uZvKzA2Ojsl67vaN
dYB70ZKieZBAlyu2f10yTFX3ueEZQVdd/RmYlaGzy9xnC1koHYFWnyiLLzDcatGceeWstLKhrAy2
HsJZm2Jy9Nbr7cVFtspYnCc8cL7Yd9g+3B9xnzFSzMmMpWC9klm1BqLmnEBYg8te85s5dUHZYQ4E
ASnt3gBg5YEi3JWN/Ja3mwAvCpc8T63/xo6m0UnKHhguV3wT8g/AJ2X7E5Sn2PIPWmH88SDmtDAT
guqAgHs61dXPihAY0LPGu7f4A3mQezKgOhkmXJasPQGty2J7+1fQdtbVCOhJp0srJjBvoPWHnCyc
JbkZ01mJQppetlD9mTw7a5YWH3k7dlAPt8S/ghavSCaG5J2uwF1zvcpbaRXJMHCjbhlIDMYFCgZ+
bJS8qLLG+XbOumLihODi/mPjDMwV2U0Ea5vlMBYulVad2d2Wz38wSfR1DAkFNuYzstczhX15Lcic
y++szNFrgczwwMeuIyVsYtNppEZXUTT/LSCBqWuYRza5dMS7uNY3Wi20E7r4rtwQu1uyHLvmue93
k7IQlNreTppWJcnkLvQUNrv0fqIlV7P3VExDMXE0uuwRL+AwqP3E5tgyNShx1lds3o1g65m1kWzC
UEOubsILavJIeYfX6tdkF64nVSx3xaWUqHxjFw0yNdydZxG/w7DyrTgWIef4oEZKyslzTVxHO16I
WfOm4teS+aOWPg6Vg/fbYcHxp3iFFsOj8Hqf6Fl81t/HBsk55S2Kytdv7BYkWsePqKPPVzcDFrB4
Zhm/9WjbspimZZc+ag2eP2qCb6OYzl9SZ76QnIESksXyAGEn5fvpG5h1CDCAHGBj5aNNKe47cHvj
O1lEjnIk2zpYQGlu+S7YHQunuTHbGCT90mfIHJdGve0R/451GCmckG0eLzjymOnphUpckH+Ags5u
aXtIMI5jUWFUYs8Ihu6Jw2Q4u1Bp5b6Nzpgn93wp94UEp/yueEij0CBnnKgB0xdF9UDNKFAo2dVT
Tx5XE4ihPq7sYO7tVqDFRc3T4c4XQZ437JgG2vzDn8LqxGsm2Wr6GtqHFY1ao+3qH6ZJCbTjw7ji
LZuL7KLn7J29RgikCSYHXAkEq+lAez962mpQmHac3LndnI/gGcHTCfrm7UZep26+JrcR7RKjU4vs
mTbXIXzG8jbWPd5ug3j055CMeh6tzExxt/ln5svEM9Y1mnAiBvM/fnRTWNzqTJSAa9RS45IJM8k+
X1mD4jwJ7sF+WvfiH4aNFKygVZIjPEzDF6gnfTLfyH7aUIza9m7fnKlmhglZ+XAxJbPBz9CLuoIU
Ci1yw2gQAQHIzu0tw5+uZqUF72QFSLycs4AFThy0iYVO7HN039FZI0LyMS42StUZ8vLef4cy4qU9
23f7LvMu6TEEgquwgsUoU/jB71hrYRKQZh7Jqeah/R2ppAKIDknJ8IfhxZIhif7fe+LZ8z2JbRkH
IV/D3p5yvBf9OCeS127SNKf4PUltUSv9i++25eoLKWHaxlJUXYjKA/Cl7JlMeHUW1/qepwiCQg/7
0PK2n79TAGPtNVzZmfzj+F1CzsbgZmuPSNN9YmRklV5oy6ASKnfRImzr818nzchoxqdHeeclpR2O
TnREZxNhF9b2y9I66EvQmQzsgGkkb/fHxVAZaRt1dNs8dwWj5WQaJEX80IsuO6/H18X0rAUFnbxa
KuiybsYKnScpN3J/aXk82yQ76nYwSuqraMnkfJcSIcHfLja1YN6l3UBreF2ItITumc5yfvqME/wP
kNIpaVxIbm6fArfh6ITsg4XmulmTQl/5Hrz8byIUuxu9ooBCoQBv5T90cU9NcUv9eH9zCRxYf0ts
lRyqo6voA03PCk1tZPaXyC7xtYv1PD+eX71NFff3lum/xKRcCCtWpUx3WWB2e6Xs0onMxN8JlHSA
ZR43Q91KQtsq5PQEpdMkY7FCvSPjvJ1ZegtcYYimY3dh4WyQVJUrJ6gFWcrA7OXyByF4ManpmrTW
CvCgAnfhuM2f1rqPkh5o2z7S/NarAa5u7dzyqnQRhLtrrSUO1MUF6T0D1Ia5j+XiyoncHdG2dJvE
xkqmT7uG/XlyMCxLepHG0igs7Afu8yU9KG8B2ovoP+7BVc/zIqxgBThDYOAaARv8PKhYDJu2Dzt6
0azn46s3fS8Jgwveo/GftsIsl6UJHCvGUaL5QSttGEl5wxCLxrZPFegJOnRTCz/FqxaqkYlu77Bc
VmmD3T+sprB13Wjo17N2VpF0UfCWzGgWdsQQn6F6c+bMC7YTZWCYj7LhaJT9QTOha9SKPSGDGFBA
D5t85Vm6ujmfwLU+yp64xTsHMZIRkQq4BfA03WkjJ5YHl00U9xnNSbv3CciIB2jtroEe53gQNpBv
/6pmbLyXreDtJJ2Yo8iScnazxwJklXS1OI4NnysaEfIYLcjbvd4IoeBTuB2UwfcScopsH96pc5zD
wL52vsur6IBoguT7Zf+XSnB2eJT/w17nPuB8OL1SaeebbJj5FNCVGKQ5Usu6izc0wzPfQ8uPg+Bu
CqlWe0JgonNw2uFDUAsxnIy81bgfhJ8Mgk6GiIKSIcedrVDR6Yh+5Hqs91+PHsaCHH/nE5UAAmzF
V9OyL/LuWRRknnLbVi6vpSIcuFhNpfEWwRDnuSG4wfFji1DszVxIhZHNodnYek0PiyfMJd2eY+ko
mSdzhj5xdJBtKI7GIvJuf1qNH4hH3ntP7xeKGHtZwu2UcHUHnGrsEB05wkjNvlKTezulvTCiAIOm
bDkb62W5bE7QkdPF1eCDOTgiSji6TmIufMnGGKLahE6KLtmGMd5e4mUARmoa+bhmPAXJPSU6wPp2
oHShLhdTRJc/hUV/jjRvTm4cL4HhzvtnKZc9g+NPsSWXCtv7ZpYGSq/uBML9O8lnwZhcY9n5HcNr
ZbIsApiMxlZpoL9fTmuLQhKnT0cdM38b8fMSxoUgoCQP0IcarcCIksKt0Vl5c2T33BWdQ8uGLMTS
mZqVSp17EyST3OeUXfgqFQfKu+C+cjgDv/+9qPJcMUdpsYKG9dU2pY67Q2N8oY/WVql7nQkwQB6V
jyI7c591y9Oyo5kbl0g6yiN0K7OUb1fp3oCNZIjuZPSuNbP5G6eeBjURvat6BPuXnhxppy307s5f
tUzYloAj2YoGr/6NAv5QEXZBYV7FTOxIBkfpK0JSWaUbZ1O2ppquLo7qmtQZk86V93ZHrCtewyub
UHOam4GAk5uByG8OVgQ7TuxFysHJN1/4BneGRyd40ClpqHjuTgLEgu8d8NMWwaMcOz2Mt+noeF0O
HyGhEDqoBLtLzdOhlHUrK6WEz+NOxmuLrwsknoV06RXKdby+9DiVwRWTDZMAV9Y3nWsA5VvkJ6ht
Nqe90RM5cKshVnzDyBFYLKROixnkwUNRxuIU3m0y5LzGKGaJOq2OMIDQczLk2Ct58Q0UHMpIOjya
22K9hCmleRFJaLPoxGQ6jFU/UY2PKzeOJjH7B7AEx5z8YzSsnP9tThAsRzSlGtMmSYXV1gM71Z5U
n5S4TTy6gmB2ZL3SNdle+9H15nE7f+836vY3BHUidOfSoY7wcUMBH+dUy5/HsVfOYlzqGPw4TdZo
mUNqFRo547CZSy1CZxYd759ioBQBzPisJHOT/ru5F5hcqqnXEt1x97UFj/vCXlAUDs4Ir3adigz0
tARzx/vb23xntTdR+v8GxX7TJirl5mylbPkwdrQZQhX5KpBJFNFZdzjJfo+um1Wu6ZGMLTTYxmao
WCGkAtZgNgDaL55b/1vC1Fw1WPxSEJOlI6Dpy/5a/I+FPSluhGFDK/blHez6RrwgK7IuytkKvKM9
VGynv4BjoX3vJ0ppRHVtdU6r1+gSJ+Orjw0UO6riAW5MsXOOSbzNBj7v2ueyb6L1X8ihec4bxs0C
Bkx0aBtOP5hetFalUfKMS0rB1AfFEjsiQMNncrzlmTNj3f9kidOaFP2x0Gn5yXN7GZchzSy/dmHJ
C85xWLdMQVb4JS5LKTotG47RTFOAPnCvQD1uYkURJgJThIG0xXpI56DDyePQ9QKeEwtprQ2HcWmf
kpJs1J5NaNPN66C/axiTLu3SF/U0IASmRwdKrjg4OPzF/nQOmOvCqy25YqL1yi6khJblrJTHCi9J
jdRRntnq/HMoR8Eg8+NbzRghbpG3OnClZ4+H4qunYdoEdARg5QrLcIu50DPcbyI8RM/dUAgvZdg8
b2l/3/24MjzliSmLRjiT2137Uu3E7Wja78VyeNW4PywWIenqTiHWwqwXwkLff2qMw/Sg/zTk4IJ/
iEbNGb4JBiFWUQw2U9Bfm0jAh5KtvNAvWL8iSdfrAb4qJrnxEBzwpn0h9DzVWcCGrAtqfujwClR0
/9ObBVcn57P6Loeh4lANRtg+A5YRy4OorG0bK1qwItGJZXhhJVP1ZS/Tlw0ctZgxNoEeofqQqfw1
WKiPS8ZMaWK2c8n9AizodhknEER6Qn72A8CfmCJxuSoJ63viZxqOxBA1h/15/POYUh78RXeiTxvd
dpqg90RnWPs6I3qvCX1t3BMLy5EClIV/sH6nckmduEGxCP5CYI2id3yg3cP03Nr8lYW+a/USUGmg
fH65w1J/IMDClYg/D6zPx/uwH7KYC3xNe8FGjj7vc733MLD2Ga0atGmNqAtHaeiXd4MQcpFxwLOq
etgaMsDAjyuoMLzoB93SDGAr5UuSJLH86ixsYcI7CBhA6jj9X3LeS/QMnGqmFu3k+zI9ONo4sGbj
EATWgiM5g9deJORvvfMgiWhtRwS+FTU5/R8mhA6/pC2i5iC/rIP7DNTKkXY3hPFsB7C/OwCyknXO
CE/QrIfNfa0L8ZxKOtApoaCiBrfh9Fdq3R4MQWOurI1xwrs7w/90qI4rB3kO9g5CskBJW9lBsnw7
v9W4T3nEiMyvdbGF9G4Pp4LMzDtsLvR1hIzHKwf5V0nqb16FC8zJDEQ5zGXBUm0hAKMkLRCt+AR5
JWEfMea2oWeixM4J9ZMoI02TNpGXZif9vTiTGZx8LMNcyJgjkT+GcTQWJ6TuG7LCZo/mXLTLqJJW
Yv9ksmANS0GEO48F1DHZZpECGDwJKvafV4iSrqlB/uEplvkYiN4rGN3vV7D29Rrpq9STS2RAjvJN
a253Zzitw7AA0JX8KsXSdH0DHDylvfdZep5C1BkLc1jNsIJeDk0+Uwjx9Hh6pvi6LzwpgWTKTFsm
+ro4dKkW599iZdVRNbDrUxx+M3yDmZS3356hYidbJGRy7s3cb8PMpYrVCAeGSB+RFY9iEHa9gGo5
KpVHjPIDoK7i1Brqc3b3r4eLqeSTynvI79JThJuPc5T+XJvum0/X67MDfaBIiRRi+dG+O2eGDI9g
4BozjrCuu2XU2I5lBTUqaVva7OOQvh9255TBeHCCSwY01ZVDd9EqOft0gw3ptaQl0Sv+/089uWRs
OJ2auGNyBrh97wAaYN3EK3c16eSyukNy+qmXkoV2Pa2L7zNYYqLGGo9Q2hMC0imhvaLCEzECCQ3o
bJ+hT9DfGcNlo8TeNEvhlVoWDqVJZhHtA2dH1GwmADyMUKym+LzoKSUN3zWjkrrOHTP0qsXp2G8k
k8rSng9PZ3jGJ5QlH0idf387xsmt5acZElOj3Te5Z5QXM87ATa5+qk8jRWDLWXciUboZBpMxuhaT
tcQWgql6CKHctUpeHPOcGK+X74p++XqNToh0TF+zSzL1/tkLkUzbuw+DB+owJMj08ouxrF45rPbj
mUo3DVyyNe4Zi/FD3HJaJBvb+Jrs21i/jFTwWbveEfI9hh8gPe7JSfcMnTZrE4pwFcPQM2gjN+Sb
HGRInYGbaKblBwUA01SvveuXC6tAqBB/dtaZ4sIyC6YEbRedNdcMoV6mLMFS+peXEQdw0ja4D2H2
gSiKY+NIt+MiJ7d0Zc8U062Eea4Q4v/mHq9jWjbJzCWlNAP6YKLAzTgz8y76WmLLkGtIJR8Un0/w
CCpzrVyRS8yJQB8jRfbxPfndA+KnsFtkL5u4ffP07jcW+QdX52uZwkO1v2iY4Qu8szIwAJylDStI
A2cEo41KudSl9pyAGFjLciGNWPVqssjeLh/qwGJCpr58M0MV4/4/e8HLvIlRHkWsnMexoP+DgaWf
athiQRZCGFsR3S0S3FzXnR9z06nahKB2evrzEKYph8NwIEoN/v0Fu4Gs/IIqyo9z23xIbrh+sVLz
isdnO/ZF7VEKQv06G8wfdpmvcDYYjNJ1V/al954niV/lacvYds8a1DuAmSO6SltzGJiXdZSO8+DO
oEp0dpEsctMjd5n5BRUABVDysYwttuBeJuvkyv02SFbWqevswLMtj7ANFv2F2Q4+1QiTXlRAx/m4
8D86yoNFu4Rrq8yROFgOBwp8nZRcey/OL2gQAHbKdTCnt/aXl4dISK9f73WLN2wpgU4ujnMZafpD
BBt4GtDmdA1BeCB0jEUN0YgnKF6dHbyd2gfOyu7UZa2HfWpUyiTCoGGIzcA/0GBH/enER6/xj8F9
U6tcewScLSWE98R2bRoltdrhcAX0ayohcHIjo/IoQAKrhho+oDt8AjrmfjH4J7DglIZvlGYopwKo
0sEEuqa+PofwK9KBjBalCsPURp4ISs/86o9a0OY7H5MMcYGSyEH+6uF5Xr7mCbWEAizskvlFavTn
vO0xUf4oDBCbPe3imqVvzXWvBaL0T/GRhru+AG0ZOXedqwAXR/+Id3B6uUAQBaNpeL2ITCCKo45A
4YhsxFci8WdNFEwYhNuUuHJzj3I7a6nztbFxviy4VGANVknBLR7ieFeob8Lz11kgwicaQX9D5R3V
zSaFIoqYxBxin/0qn5u6K6bxcnpZzK7ic0QWnfyxdgIxac7kdkOjnHjSB5ef8mM7nUAJbjxQd7vO
Gwk3uYirkTHee7HQ4fCrkob0UTooDQZXE47yn13zKpcc3tCvJq0F9rohULRosWmlp22SUK2rGw+W
IZZwhR5zCRUETbZLDeggRoQgL4A4XyaTMPFyh4hU09HkmzPCN5JND0vGNG7uhXpE8Ux5E2D2mGA2
5KDtUcy5S0xxBvFn05mQtE26dzHidWjHDJB71aHQiI+SfDnKObALMKkeHZvweSllguLw4wM+PRoq
C0LHGHY77v74C5W4IF56I7W9ie3gAasBiKrcLnjojCdAgPqke95PLOfbpD1rGGYQuuHpmJGG3FB1
dGndEmR9ghz61KEqJxKAfXiO+TsA70hEV2YQJVTHHiVQ+ASFpQ+WZHrzPH9mq51f0a9/UGghjBwq
3xyWh2g08N8ttCVxCxWFu75myDrxTh2CVpw3/zEP9WmNE9VxouKvPLVGMfmK87xKBRV5VAAuPRlN
IAAJVc5/eE5BE5HY/oAVp3OLBTa/+06vADHgjHrMsuFHb7SpKl2jW733dfM17ikZhNpbkKd9mHiO
T8ApkHIaTi94mMJn7Z3n3lIterye2dvSTr2cbrsd42EfhTbZ3IJgXxlFJY5nyCuEXiMIaSNtK03q
IyjQRX0gqPD2O9VvF7hcSxnz1GWzrEGoH+jPNXg//fp1+iuxeewAbdD/iihqKG/UOZKmBWA9Qy3J
gh+MLTsRRrU5PiNGrsOI5I0XXvDldhSWpFcphPUlcI84t1kb8qkvXCSkkdeRPDVQMhhmj/r2dgri
C1nfoOY3JLyqg6hheeB7bUdMr91EKAA71Vb+FmWa/V80FyD3AuBrZHcLc/uMnMC5zpatnFYpc0E7
azTEYCFFKBDVIkc84BgHbE6hSLeXsZPgRc3u9YnjTCuUUY2JCBYyfpng9L1U/m3RH4WUvGN27SnL
j0CD4wLxx3r5wHTxtUaCva55p50XddX4HJX8JOFLvJsbKIqT6axut6WpM0h/a3RHu84EAbVIFtCo
WymQemnrFiPRRyxfP6ip7/renUioqQXwkKpI5l3SS8P+WCNhnUgoDhCXr6SYVL1FwqwHvVYRaloZ
YEd9GKOa6qAP824HDuCA6T6whSiwXzTaz+DqkMMIYEHjCpQSAMjkdfhzPmJqd1RNdvR2vyzUSqnx
kiiv/AqdtBBUlAI21gfRUPV/uNAlHvMdsQYVlYinMsydpIysU7UmKUNznw8EHkdFJaa1oThnQdts
JLeRaIXz+NPjauQmMjvrVBE8nyMzdcn0OXcZZ9C0Sd39Qk3SKjaIp6E+RQAadkRvU7tXrWPYBdDm
Agp/y1IC6/xE7BTOxeHKIAAVcs182BG5HP/dNTBogpUEqvTqJgZWAia35AB/T/so7/Jj5Md6VuiX
HpsJqje1zoIAqRWZMnTyr65zikHeIFyEYYj0pM7pXX5cxeLkUqu5s2aFmHMFxWcAVXcj5MG+xV5z
YXaQMTVfdqo4jo0HR/TBaZeTgGvWzJnd+mm4Qz2KfKmUDraNsWYCDy99c32wTdAxMvwiac73kWVl
uoEjjFXX8nz0WikVRWOhFx58oGfN9f9t2B9s9gGzmYBEluPO4raHyN/m6zBSZKYibaiMIAcWN6f0
9vmAvYU5z2kBFf1DEcb35dfpQK1CcBcNPZk/jIjkX4Hf/KdhOSyM3AclcP76VpC+P0dGdOOSMkfY
Do8TxGKq6HAQ5hDdHvpXpl0Q9UPKhoeWRd+H2B/oR1/4oRCNAsy8DNdEyCqA6FQ3isMCzGBe7CHy
LtRck+0BThSsJI3PEh/Pizg23Ee8q9mUuWyHvpiByo1qqbHbt7CAN8/Vn3f4nLuZ+QFtK0TPWQC4
WN8RjLuVIcZyoWnkqqG7p+c5FRKsCYSwwyJFlggWoitY/5JtEibv2JfSC2CCabnt3QqAN6U+j1aj
YtmbntdmT4ABaZsPDBlQz5hAzjkm0gfBCWfSWlvdEicKRAjU1S08UrnK3nj85bmi3ETGQR9oSBbD
VfHm308cccHjpNbP2SV9Li5E2Uv+3/blGwg8MqPNYDNjxFYHVv/d8Ec1shrZO96fOMJDMgslwaPe
rratfFUWLXsQHYEpubdTNjtFmKjKc6BNgBh16Clw1VvcJced+ujdqjpjcnXdUU1vG+3KJYw+5zg6
KbOPAy7ZLNCJrZWkB0QphH0ZeriOd1n32CcFOAxd4xtzFdVn4SwLRcwQrSPwoulMXeXd+Btq6PtP
jpPhPpWd+j01sViLfl2pbJVrafK+nhZOStSTpkklfD/SyAtVBpyF9msTJYqPAVlHxdXdETLAIBlP
CHb3SPBdD094eoOdgl7lL1+BeIq8rv2AhH38kJX3bV6fAMkDYrKCzeeLBr0ZEg7lWKxwgGzg3fB7
VFlhLyVpEGcCiKjjqOUCOSjZXOd5O79uN0iBaoPWiuHx/8xUCctRytd7PfnLMc9NzhjQBJyFIF8r
O1+K2JZqNxb67qM5O+E0mvopcndMGaEj0LYWXEaFdqLS3xobSfN0MZ2/tpBI0YIBCtF5GTo7nL2n
noCZzxqG/zKn71fVEJaTunVwGQju9iSn241B9hEFKt5PEFN4Y4JSaLxVdXV07OcRc+RNeniMc6Zy
WkpKkeRgRTytWxyKNq4S2OY/5I4SW7SsLAnuaNbX0rhbGDWU/OunZ7vPPehWpzaLO4MI+SPE/CPy
u/0rDVPCtbpYdmKyTceB9XF0dUY+vJbzSz5Oxbyc20VTUbLtli7kjLR7Vvso/SBpisJdz9bxMcvw
uy6DxYyXBkpBkcebKEA1JlCU5S8nc/YQbaUQWnRMV3sKDiE8cAGLG4lLr6IKzWzZEKiJhI7AJJy9
3zle4cI0OL0Op3cvf+qYmJQIPFMJ7x67z6sQx1omPuySV+8XQKJfchaeieV6q9UGj1uGsuqVmMi4
oPRhNQGV2ryhIvN1Nis14A4DU1xDp5EkWUvEJ0D/z/ky8BsnD5qLTLhmd1f5U2HyzfnKhh7IHiWf
yEMotZ5NL5t4lzIiS99kUOsaoZT3DHf0gO2nFwd37Y58g3My2jZ/LCFrhx0C1oqQdvkD4jRT3tl7
uOW57L3DAGZ/wqWTIVAoF7W988pCTCrTPKYmMUaBxxs8xILPGxKsPuu4nE9CfLuaNteRY8sGLBpi
vmHSQ5Q84UunnbDeLToPtzra+YDaezzvmErPo2/MvRFGtRKaf3AK+BEK3l9VUComef0KFdCpxCjj
6edgm+3pqy7CyaA3ZwStSr7wUstyThUh+CK79eYMi5ZhKySAdg7iQbUCnbw5C8amT46Mnken+Bgv
GbskjqN/0t3dpXIPbvFAUssSsAT24gmX7bS77ZEbFHfUKia2CN/BlBXWCMMxYtyNJElIbIZbbV4a
ZvcaUhRccoL4yY5P9nHZpqg2lsdGOGmvSuM2wZw/YOLd5PAAjX0uF0ykJpIQxU9gB7Ki/BKv1FVt
3oKhyoXz/z5g8cgyeXl92/D7KNu+4qUWhIAt61yNvn+lnmj7AWYIo3rt1wTbjZ/siJyOX3Aoyn8w
jE/PHhkUCpmCpNoaFIhIdwV/OZUICprgFBNYgjffPDe3BSEdjIr4hg/MbCShRg+x/cf+rTzI4Bqk
sZsQ9380mkbEBGfayewK0hRzhdgdADB2SCYHxzlzxmbW53asZ4TAY/IZAoMmiI3+YRyIfyxusFt7
q5siJKN5JBpk0LdqUvPsgomhTREVm6jhdnCy6RyzA7YZc/dF1kawpM6hhUAuot3VFP/uEnHOSSux
fA9n+4fcKDexmgZbgVp5vgazutzwAqT7GE7H0hT3307DZjPI7zmcT2nvxQLmURuRSbZpaMu3OtkW
LoMGLh0ugv34dnYA00+G+HKdHHzLt9CW5LLotWM7YXwzB3l42zjdZCu+qdp4qbHsqCaOsttSKifE
AnqCXF1S5nKyN6iS2uf6ykUBOKMFeTty+hoUNcYQ4b5YTk6SmE7vu0Yci3CizgkjJz6Pqa/8CDxF
lu5Hyc8c+Y+ecjoz+V+fL3H2+3qZs+hWSHtnZ8RDMpfBskRHk5E0owQdpUFRSXJgZFsG8+YZW0tj
A314t3dWPe7z8ap4BqY5eI4ldCch8+Dpu4QMNRVZDC7c7gNIc0wOm3GrNBLGWcDzpIsm2FTiRqvV
k3vsDMYj49MVcrSOBO34cM07sAj7ghEwM8RWqv/xKs45lvFHoXSNFYa0FAQg54nt5cvGjiojZ3eQ
iE5ZixAVZ+3k3enM4qGsIdFC5u2YKupkt0jGNozXXWxwLkxrCnAPMuLfq6HJDxBglcABR/CAqmDv
Y1tUe87loDJNhnLqGwkc345awpZlG3QfdS6LUP6o2YdPaqxHElO/l/gjH6qyFcux87P3KhD7DqEk
1gPGK8ma71Xdlvk2tInenOPqZE/wWsstYVB3J45WIzKfdtUqRA4Y/ykIZ6CtjfrN4Gll2R/paemS
FdE3Cz4sLGUQTzMuoBUGZYXl/uaMCs8wpuQMbatQx5YiC5yxCOGUdgL1Zdzu7MqNY9n1imuog/UG
57vFAi6q00CC92b4abQndvxgQ9RTKDA3kkq2ixgvFbcPBVqpcmFYtMCOS8tCzFocJqQ1l7igMp+v
hoYTEcuIba4KrhbxPmALo1xZxnvKojdxVPjmb/Z3x6ORPSCAR0u43yfnymepIBHXzM6gMEJu0djc
fF5SI7o1W5WYvgkZauMsYniZVVzQdIsxla15JTRJras4QzB6EGdUDr1iwBDOrC7tVOPBluliawR6
SJQZhBTv+nbOgES4ujNVNL0csaKJ9/KxiPOlZc66SidUSPFdzunSMsas6cjLqmdEztth/QZxUWTk
72aXBvmtgiXZkaP6z6YJWh2cMlD0RWzx92tYxJw7xS1irjM7VkowO0e1xBCFwXQHJoretGbQv7Z+
3uPouAtOzwfryftGdkTz7UKikOvNVOwnTL3wSVywm2J7WBdInMa1jXjToFdSTxFBjfkorY88u00G
RL89zjcpzzQT9FOyS2iHihx2o/0Y7XrFNDsBBCbFQP4RezYXguVDmQLbaUsY1J+mDE24J7F8q+m1
hHtrvwETAE08dIGtQNDD3JzCQ+0KQhPWLcrLcbR4PSpKQn34hix+INk+PLnGikxZag+kdyHNoRZA
Mr7pCQzCC3ZipOc+sQkc75x4wkhuo557uoerbIFV91p50tZGtcidTSgfEys+giXQk7/gz3VWARrN
Q00T4jM3QFH0BJoHJMjtnZHqqE3dd10ZF/9Y47NGb12u0p0ZZ8CTX7qVY8NP6pvcTbG/C3uq70fn
S5H5fVuwOXK2vOCAnjB3MQ9Es72L9eb3WIvAdyPfEnpPBw+k87kYTQxyhTzv5Q1V5pFVchIHAG6X
e2WEnOWkaqgdCPwZBfhOk7S/VW82CPmy42QWBxG/bFqEgsXLrTPSP2gBr7xc8iOStJKVC55/Ormm
E+7HW9bMaWTyy0w4aBhUXo5Q6SiDHQNmJtcpcRHC6lo1E0p6KE3oeAf/w7h3rKKQdY8yw7lrGZOG
LmmyPkQSLXbR1Y6huH0hw6F60ap1VJYafrk9hWDvrQwVVhprlhUut5yozCn9MIhVUgtr8dAlDyy9
nDrYFXRGlAay28P+hRvouxzFLIAGfhKDVs90aROZJtT5pyfuCmJzKLQ9tmj45zgrWI8E9MLVNHnn
hoqoqtd/EEv2Jg8PIDB0fIoImbfFluYLJJw74OphmXgeYi22C8zkNF030vvx5UCMuLthqTAeAV06
Z/Pa7IQyDQD2GAC/VERU5gYjG0iPR/7TxIYfFk53yjYe9Qie9LEziKqTKt7R+Z3E5ZtZ3z2iKo5L
eq6qNfgJDkZhh+L6sXYXep/wiYLI2uZFAAjsD8yLKGdp3sVNJHyqZcCtX76lR2Pms5t6Ei77qNyL
Pwj/p30c+qqrhqQj6A5pmVp9eY/1tu6BIt0w7cwa0plOmFIqhlMTS4+HUFAjVlATh1hOQ27VKZXp
UY1UpvEBEacqr6sGgkXT75JTrpcAwoAfXFbVNZyt/TSrvhew+yxVa5JNBgo+w4Ln0xjAYR9utOq7
PYKy9JI/rC7CRjrtEPmsoYpVwKPybHVET6tKyZgcLasPwNCCdgUqKFLBiYXHPXK1VhWbnLp8En4X
vHtfA3oa1ETJOonDjQo0wWriEtNNAK26z8oY2MFIwf9yhqRqQSEceLuTcE/N0ZGSEQwOdkTeVBqC
YL0PswxSMPe/ASQdi9T0yQ8WkI5Z0hmYG1ejlLUjaCJJKwmEaGzf2HpI1PE25uf6DibcTEpT/6Aj
XKcvSJVV7f0tl8lSKxaREYImU/xBby8TLzO3bdwX4K6GXbR/RsMP6mUyPTWT+gc9w7gfNSkgYCbO
PJHplIKRPQ0/4SYAxR/ICf5jXmuPG8AsJnnaL8O82C5GpIk3WGJwjZ0iS5JZaQO2TmYewKfnIGcV
OKKkUB4SfwId7h47LiRDQmdS+4+c5ZZf/9tZ5QW5OhhPKeShT98ilsv3hK0wY30GMt8wgfM2JNkO
ZOpc9uSiZjksihWwQ27Ltzbsf2FHwx1Q3Fw9x75wDx3xpdEJGUnOMxhJ4V2/qlhekdIl8C2flQvM
O0mHHvOXj86sST4F1hBq5Hf8LCr6GrTUYu5RWDcAaSyzhVSTdPn8pEm99Aj2yHS3MHs0Xs8mz16f
RpCMMe4+Xog8sW9TZ6YB97tlKfjJmXQK1ItJoMOFzG49SLoT9qNr42Sj2TDJxp6eNMX5IaHd6+Xb
OhLAIUGTX8APXWKsTvy0V2o9jQAzN6C+Hv866osEgpthC9fsqOgCXihZyS5uYKQQhzYEz88gf6I7
E1+BJQ8MAFFe3LCN9GE/XfQ1dcSc77SI3ZnrP0DXJ6/EoSREp2Gso6B3Geqknue3X8hsQEdI4Th4
pCaix7rIwvgC5QObz/JZIEh/muQ6/S3Pn/HomgfarI6kLdvAnx6gjsacVBZXbmqwHCAbIa4h1emT
l9Zz08cY7s034K5FL4huxoavPxdquthdBiLSOubhnawXtaqpTdBmdAsMB1qY5vJIFJMbVJaUN+8b
GTKgSXaQyChCx2gn1LZ5KjQbM5qK0DYy6Vh40k+XBgcNa56arPyUwK8FDzx1fPz68yJ3X1pULYlc
krkviqY1ANmBFAhD4dCPbjXMTgo2oQ4osdE//iPshswU48AaJIVgV/9BbeRxkDShtdVDBbto1rrI
mpPSlDy1KYoY+c6hrL0odh64oN8dbVFfzPqShL1pc4pK6ccDC7fBU22sdB8xqWp7COeJED9NLxk4
EcheMUnyGwVvXKHUGFv2PyrFDEzU8d5T8pgD1l+zi8B6WfzWjz0GWDv5hdDnE8PWkTVMmhxt3Hs1
CS2p8/jmnw9KdrKkY1kM0tc64AcoRX32gUFHSLff9ex67cfj+VLLHi+XCAq1uq8hWqlmI+QSSwxB
IFf2NL4fY904JxH9Ql+JPDXhY29dPIY9VRBbiwwSDrdPh/kclZyHdK0V5UYfrXuN80CayTnmyCBS
hwHYGZAJyhF9RrbFI+Ss6pzh6tGCOurRnLPiDNIO5z4f9z6OkEFycn7ZGbgFsLVzEwrMQM0mH6J9
4mfgirtEY0foq2BAsd18xIFvA7XKPoi4ytFEVABvTgWcss5vvBU78pVq621RJARnVckZOTzshKRz
M2FNGwn6vvu5v+JicNbNt8Mjx1wqXZuxCM6VDwNeN5oE5oT5ruRgc+qx2+kq5DOJUSXD6OV/Xv7b
n5VHCwneEXJSNq0jXEKM+ov9X9cwqH5nc2A68LKKwiguSXGIWmbN3McGhJ/EPtxQT1GMmu7RaaVo
7lhhTDQJSyGVJKm1B0/4Jl+bjdi+8E0PGX+VSzY588skOz5Ym79HnOUcfiEQK3L+TG9FY2U7PD+h
ffUSxJ9Kk7W2Qls3IBI01Bqbq96WFiMBmYkN0/c8D3lUl2ik9zkcB2N88NZmN+q4KueBEmB51W0/
sE40j3QFjYGaLHTQRP1fnErgvPctg07Alwavv7kWXlr7iqj7XzbBrtjVjnENaelVZXmbiDOhP2N1
o2lZVIbpZP3EcqoEYYzUt7QGzEkaFHdNmlR20060hIFjupQndI8hPfZ7kuB9Hw33yNBgoe2lVoY/
bJ27enyI2IbWD/ZGks5V7mbTm/g8XJKoL7ZFWk4xGMhW6nqDPtZ1d3B9yE5ARNqugmtP3dfB3wtW
52yidOmmm8XmhzFBK4EVVeUnUkuEjyBqEyPKJQycOAr5NIXCB1aD50aybpgGNIPNMEGhdQxeW5VE
gdKQsfMOqMlQQms5Ke4MI6vy2KemBDKGSZRddyR57i5/aYelZaJfWZh+U4lAdy83VEf3aNbcfitr
+GZG4MwY2xT1IDqR19kBea5xhizYQCluWsw0LRqBEPjKD01x6jRFBaYU4vf5Y3+H69lNra335kxC
JKRiBlaYHAHT2VN4wCPFpHyD602sCsQZ1woHRdwBagWKU6zgHKxYoaLPVvz7Skqjo/hoc2GIKDQp
Je6M3Wns/oQUilhvkNT8V4HLYI/fQ3yeWp0G3dShSjHIG4l5QpQa/TKL40joH1WTpBig1hMEzo1g
5eVQr/pEOr8txPGChVZmINv/s3REEpF/eQZVe4jRsWE9Tfte/jIHzpHBrwfByk3bB7luYM/ix3gX
AjFUhOqjYhPIgV5eH5hiZFtt/HOmDCrqF5udTMfDyytIX1Y2zM3ezE0DhsbbYVHEmd2dOXAp8Z4k
lICvbiz6UPo/OsYtjOVLvdcaabR8U5Lj2LgUm6PKZIsPFKf4jgunUq6GNEjNJ4Ax0fbrg3/ugOED
89fxpKgLgvj+eFIeMBnWucm9uaKcCVCUlxtmeV4pd3g/SU1mVPLb5gRKrc9nodG2LjP2xdta65Q5
dyUHvxrHDiHAJRKbe3YzWe36uDvriKifSXsUvh7KUagJ5+QAJaI3YkmhhxSz3loWSp/Gj7MWblMW
FSRGWnG/1LoQCnTtLnmgdvAKebLcq1g3jUcC29pCQS5I+vtRPmND3VZiWCfYyn0O+i+81HIlPLb8
iTSd58uup2SNdzmfGVtQallrzKvEzgb/pzyzl5hW8iBcP+wOuuzuOisHM/bIMCP5VcRhIL1if4DG
c9SY4r1WyMNlYBqZ/CnPOEqWiPEE+J5j8zUyT/ET0LW2gzndeMvasOI83NawOl9Ov3M66T/5Szmh
T1cTOfiZSv0lgGpVTu5k2wYzTQUFMbBCalC5EfmtYsIlXU1nxQMLr/4yM3lRfsHD8LWBM99T16BY
Dj3fb5CkLp5JvexD5M2fngZFngukntYhu29bJmmq2LXIGVdMNC+0JkVsLzvN8TaVmeGzXYItzmuq
Z0bhhtFwaPBtpkuKHBF9NtgcrxO4zbiFOBLcnsJ9mvOnmU5AOCM6o8QR72hHLcH62BOCPmXgrg08
JtClg5rwlKBVuhqIuWdst+Jlait3Zu+JNY5lQg2XaMq241O/AU5Q7zoHBwIStncXKTlis2SfxmeI
fCEFsDeWvDRcow7nIGve4OB+hpr2Nmxh6TxICVGS8qC6vwYp/uUFBftmNUzfnouDKzUgGtly99gB
CShjsJMB+KLMBvURQLiWtMM+scb0NdJ80h0r+6IbGT8TvJO1Oy45/+FNk8u2HS89SKEyFu3mZfsN
SGSlUt+sO4rOYKQD+Af+NtPFQYROvA40z5Wuy9/cn/aea5nptxt4fF+6PJze1FdeRLaLH6yR3WA8
NYup8exQr0IHb92IjVfI7my+3xKmoPh8Smytj2x7V/0bp95YyE3XW5ONF0E+JZ05/sSULP7kB9AT
euE08+9XNVWW1YIXSJPZ9+kwFwdiGlpv2uUgd1Zw1RKI3BQkjecw+/9c9brY69zfsAc2nrRW4CnH
awPCv4loq/ZKRwLSrxDtA5SU68mVh654QR/otQhFc4VE/pY7HvDGjex6Esa5qKNqFvehHVo3wi0O
ggSjT2VaZcd63Xm3r6fFncr7nTR9BupJLCxf96aAhsBP/h0MTCRE4EnhT6kZTX+TP+PrJej7RBoR
u0/su3RqaAq4xH2muB8AkVFSkDQJH9qevwJdT7TMWW2xz3Mnv9Y2NpPVenZdoPS0PvY1tQe1zVO1
DBzBjxkJgN8xgIA6hTjKGP4jwseSI6JmhBYlb52vZL6v1DCghuGJuyNn4Zk8uqRLFEHy4+k14WfX
zLFoZJ9qxn/5XB97a54nIHZ8gkxeGjtV41EA0NZMYXAZ6IlvEpX/7v/FD9yfsEQqTWU+e5+Fl+Da
CR5OG1Cc3eXv8FJVcMPs/K5KkLBV8yblkUzSAgmp/F7W1SQfPq97dbCM3BaTOwNCJltins+yIvVt
1gMzTd9gpOdEWdd2T6y0Yq0aRBkcpxLnGFcfwUfyEMXPyOmJRrAKZhTsfFiIqR3q6fNpBie5+kK7
eE76sKDZ/eM7uiTE51uSgCz2K7uTLqfpEjctwq4ouTI0dGWa/A3cY7kz4gox9XlvYnFCihFrdziC
Ukvk7S6lasV2qPTljYLyEcuqF478X1uBnqGfxl5dxrm2q5mEg05civHIsI4X1grreOQq1ZDu9+K1
2eOdACUwtObvGN4q/u0CyLWBy2mW9T55/dRxXaUUPVIVAkaOPW30kWs/mAyrao/v/GulWZzqyVz8
slm0X70IVZhrUMBIwSbhh06sLohKShDYJABC9/rPgJ3MhnFlcYU1jsfVKyEgg19huBuyynFIcEL9
ZhqaF0UjU478o60G/jh6Efu85yTfFHW8IK4kHDiLTtxL6qVJnKqBxWDfDKAl4Gg70BNSCI6GV7ZR
sXzILTDttOlHYhWzRcb2buaInKRG6B8ymRJehDVGFb89ELsIGri1VSgcfVBrx0spn/VP7aEUYkhA
I4N+diW1TlJDidVhKYF96xlJm3i2J5qSOcOMvkfv6fF7stm2R2RrLqzY+zc0eMGtsVogJ0Ngx5ip
YC6jNw+UkRwKNIu2zZyd10CfMqIoHatGyc35tWI15edSoxvrfGtn4XFfEVz0Abza9NYpRtvWbPvJ
iVQQcllce63q57Kz6qLaYE+vsc5RZN4U1lij8cXC8c8eKDwQSAMtbAWN1Qg/9DAaI1qGz6uRa7+y
Rgak7oDs+2WRI+GKE4i8162wSoEvXj0Ry8MguDOPdY48HdtxHI3pyeRn996OApn9osiwTJV1hPaz
TgT7ey7V9XsAGpGcnar8PAEAiQKiBQFCIcJccVnm0Up8i7MO9lLfgM3ygC+YaEipkyHJ2nx/FN3R
wB5qlyBTGweeN5hu9fHRwB+9DFnxG4J8M5NrA0T5c5aXtHW/zn9kGjXByOWBIrNJS6azqiJgJalq
YIK/9YQkPv0iQYXI3bS8gki30z9X/eEYrDvmX596/9sAQoXbpiAjxfqrT0TS3oIKrp2AbwnKBc55
6TALLoCVideoTyL8tU3XwvVIrM5DKEHg0giR+SsZW0nZ7PVpnSmG/KDmDNLSKyUUZ70eCtFf+Vk1
DyzddFEBXQmWGF5uIKPbx0AZn0H0t6ZRPBVsOsaPO8+xhG9RmCMQKjrpD+vSG+PDHBzDrfYTB6ri
pyFin1oN/QuKHBtoxnawlf7XWE2oI59Um57jo4emLvysx+HF++LCCkCjsfCj2YaEoUCBux6+u1Rg
o8lC9q2iH+5wsJFOgJMZbWx2TWxYNXw20eacS65Gugrg6dTwprmu93SxzEFII/bnf+If75Hx6FNY
kGOKi1Hf7s+LYwdFC/2OujWpAyRlqKjVYlbiDKNyolAIG1GAu520Dywxsg1cvcbAICYJYK5aZ4m0
r+a+4jWoL61Jqfy8IGQp386lBzjRb/crWd/7QU317MD1phVGhCleNc7rj/YImcsnTOxAote/HkyP
0rKOj/yhEIbjz07oshnukr4gAABuVz4Nu+1UUHh1oLNbi3lRyVjXcW0mss4Z++F74dxy23dZkn1H
q9IPPVp3YlmdF0JllqNnpEuicwuug9EhaJEhNtL9wySOSBdahwm0943zTORu4e+bH7M/lpePXMHI
c4/woGmrCsoZKSG0o7326jHrwvysBu7AVA6oba7m4EjBUE/Ck49w0cvIZbbwAS5uK9egUqOUNUtj
1buqd+FZPheffPBqBjqfaz8j4qfU9bfFJnUaFpum0zp7KngQIB8t+YLwaeltBQnhDlEm+iiWMQ5t
ZWCauj+eIep2UM6aMPLmjQmbd3AUbCFH4VuUh9GNSkJw140uALJZL7tiuubRuCHOzcD9EbVP/puO
Pj74WCMGnGZdvm4qxwWM4rfo61RxfsK5RC50t19vsWPREre82sBJaKpa9v6mS+Txh8sQ7ZvnCYH4
Ya7AxY5DVMAug84zSurhhptfEvKvMJhWCGMIxA1efwu0ZQ8yhBtH7EipvUNM4eup2+9OWH5/RVIa
XhugmqtkwGw7+YgKd77aDUbgvlmHLO4eJ/8ZqPrM9zWpQfYkrW4DJuJfXZ7Fl3Agns//Q7N3eRWX
7I2uBs72XyHY1YeylX3e8iWvLM8BfPTEgVfvMvjI72iHyQRIwDxBC81xpBBpcV5Z1MMkgGgFOslF
Kp8IGc9MYDPDnYVPrWOCI1q+ouKWR1XvmE8UzEwznejD1A65zmdKQkKoKiU6Zc1AO2mXHc5T5t2c
ou1r5y+LID/sNNmqz893Y8xjFcMKqu95fNGDwYzdT6fOsF9mdG2OdG7YnijWlbWqdiqHK+2/twrv
AUhYh34nFtGXP3tUNdyHlYI04DcGNQOH37hgUmSsbNg40k62L2N8DLi2nxChgXN3V2OwPcQ4ec7O
MKJ+hxZyyeIEaMybD+Y0GR4cTkm54ePQbxR/2ZHTpRaZ7eaRKzTfEvzk0ENafma1vBGckMjfbsNI
JAtCpuhcUdE0q7lmoh3coc4w9AJhTs4FsZe/UQcCQCpOdsJB7L5paFuCxqMcOUUzYZnMHGWk50uE
Dji85PACEGmLRhgz0qQn7+FRJB5O+/t9Fmo18sAT0L8wWalJa973bm+PvUekl7bW8/AhUlqc3zzr
5bVyXItDetWBn0EO0QeqtMgABNLZYJa/weY9hst6BO8XyhuqKoleg1BmTpggdRh5Y99t48gmc2CZ
S51q8pYI0R669I6TiPpGoW2U1l1eUxpSRsEEtl6tqWthEjVIBw3r1A0yvrbdQs8IkeBv8wLW41qD
FPcRGAHX6rzzl4Bqmx7phQ0IhhducQPjDckLwlXxY5UHpYzJhQcOPzpnY+KmIPqny7ObOvKUBmAm
441Y6Bp5If4gWhJCNz19vkVqot3+/VjzmeQ5PqWcjDrGIGrZVL3Dws0ubWTXeDjU1I7a1CxTzlrR
cxQba8pKa+tU25ji+xn05kC7QC8W09IR4NwrtL7TmbJL/0ki+5Lqvqkqn6+7dbsDoTd2C+DduoQq
I6EvZ+aFtLCycG+B117L+JgrkEMwtzmVZJmOdm00AdIbp5l5pg0tJNrzDWJa24GHqK4X7/4LebpS
W4r+AhJiNRQZm6DH1Cd4WH/jnhqPlluKmBTrHkuC7kf/WIIfjWV5l2lVWKZ9YPODv9G63CVQBRVy
Gjh5jm3ZZwo2BiujyUR1rIbzX0q7Tl3czn6cEh9+Gla2njhRfVw4QRZREQEYTuYWyMHiZE5GVEyN
af0J5r5vMF/nNJw22HBOd9ASzdRIDV5lQuokDIdfbO16jtGOffKgMIKyI2T846GLoIfOREZqONW+
VAiQaFwp6mYlh+NQPboNjZFr4fW6cV1UmTQ1v6ej5Lr+sTZ7Hs6stvLpbfyI3weMC3GH+inLbwNu
46DS9I3yPNrrJZPceU830aWoQdbhnp7ncCyfDnRGdZhOxtC06vDjRE3KnhRrP0hPXhfFdTrDK7BS
2RxBvw41e5tMDZn0zcJgWudxmv74hhW9xIp8bUHEnIy9mj0KwU53I3bvVraruaPFigTbBXtswDAW
j+6YMRuHNzOJThs0FW8tJ8e50G4NewHQBZXLRMYPeIiMsWPwp9JccwteYfDIq12rWzH7t7B30KVM
dgTkEi2IHg71/NApLCja5b7tj1SW4pdSrC+vsIs/fmtzQpo28lOZuzT2MHocxsJZFu4xXUu+Jju4
W3vFSP0fgomfJfiWdwp4eKKZiRNzfpLRsPzkVrqUwC6z0PcfFX6cbLELVSWoz+7Nc5CY4SmeBTgB
C85pzXAzgetO7zIeVa8AX31XMXhaW1+VXlSNz2c5l9vFjwLPaz5BQ5IJKqGkXxfzels0FgDDdQwQ
w1ySm89h6AeM4hq3RqMoNtXZ/nKStQIxxj61Kn6ZbADAWjNDX3jo4/vu/SCBaHYGWmbpsSXI0NAW
1J/w4yIZ5Yn4mHkwajO1QFxnYASkaSxvuGViXTnsGlCeeTx7hbbECJnsceH7NfdYDcRZ76KdFysB
LIgw8MB1IjsjWxyR7VxLcWw9DGsy7rntZdylFbFV0G32Fv/RJuRADCqMWRDTM/8iCUNyGwbOev7c
9zPY3cjaCf8vaP7RMNSO5yL47xLLnIxkAYSCLEaZdjGS5cRwr/wU1SMJeJsLv5c7ACoO0jspNENZ
O008dY+9FoGpLqhjbZ6CPBYMrNhSpjsb6/ZtQY1fYz/VUGo2N7MFqkDe3LRK2rPGtk7RBszt2Kza
vAfhwJ+jxxHQN2Z1I+4FrUfmLnhYQge4NgBRMBYc8tdrKc7kePy6H8LbAqc9wthEsfAtekClOTOw
upCiuI+Hv+IXs1y/2XEPx8mZa24sT/HmNdkm4tDOmnU10nqfNvReJlGOST4LQELd0+p1Aff/04Hv
lK0m/IMp6/kBxaH7zp/2WKAOIF+x98thFw177rfl3RQSN28DLClI9ID5OQhLfEc/THLXj0MBuc4v
FJavajDmLWH8r2hcGev4ymtinOjK91X2S1t8PfDfv03ClG2k4mW1Eb1uTcZwRCGCwY/t/r5uE64G
pbC7rCBCL2Wgk6w93u/0/LYPs3EtozBfVP4poG9LYsVLxQxZcnHjhOWpMDsKRRBUYgcO0q33dfxA
Z7I/KtPaVa5ASej9LsNzM8JdqGyCo76tZbrc4TT/WU6jNLMA0Ke3mIu7u9lOWp6Kbm+tXTJNsHtV
BTgaI773N09zxA5Nx3r5g2zXDnENWpfOdUOIeV78k3mUV6LtC/sbHo541WUVeYNl0FWeG/4WegsD
NcHjklLU33WIIeTRDmb1bnDLoJmfWUrlto0MSfDSMrV1TjHEQ/hbEWowsvQsxL5CCUVIMX4c4Y5t
rph3IcGCJ9Y89c3bEJjgFbSA3GSpqEPzWZgWjNoGcRavps4U6D271248ND+TeJbSHrl47Uyr2dK7
EbUjWLWVrve26zNY6W6ugrnR7lygUDH7mx3QEVU3jvW/QJOUHtbMqhenxNDgBaIFPf3FI8EIS4E7
gHMIhqTRtsY2p9yYM/FtDnyNuuYwZq3ydr0Qf/TYqUArnDsANEc2Bm1ecjGGlXIQ9q0FLa4icab1
iSE/tRZ7FmqnkvN3gF6xIzSjr0fPnS7At484OBGrV3rbM15w6YCsbkBThkp2x2XuYe1CjbqdBIzF
GtaIizJOPY69UI+aLDNieDXfcdfgfLM3qXvhZGUmzMCnQTt24SdDULjLulkdYihF0J9GzobVGdmz
RYSmKXb4CWp6LCrryaF06ks+Nh4CxwE70SDbMRRb8YbEjMOJbjCbFOXK+vXywEjc3o3BqxK+M+C5
ymEG4Yy9+phQaKccMDBktsqdKHpf9lB92M/rChfwLSBseDPCWN8+0Yi3d9vD/YRhGR6jNF/xv2nJ
gzSGii1P1VfqkoKDZKhvrYHa05bOeDK+MOcZT4cy8mEj6JN7qhSoL2YRtxLJ6wxAyy6T+6WoWEAN
CXvo11UUBeV8fh5h0Ww5oir1u5pi20p84QNaImRGR4kHH+kNxWQe3cCGNgXzJn9Rd9dkzr3ZpoQF
kgqFwwrQ4ATJjVurZ0x5S7lz8uoCRbwhkxrKL/3OOOt1sWnHJY+DX8NwIlZRpmlxf6jx6LWrci06
RUy4Skfcwa4uYYzKC7Vdam/NtfZEbWguMEZnszg9nY7UTvv4HF1urJ2xiFohuofyBddYeo/I03O9
QSAvqY9RDtmLyiL6ujVICIT9JnSvxtatxCj/RPHzoT8hSLAaAB8Qaufz+3vQcESRt9VXf0V+eeDs
vGcMf0rmbsxwXb12Qxf/7u8qyyPE6q+dt+OxuBj295CfAdSqcG4tGuTZsW48SvcB4W9D+AAfRZyT
8/uJZbrANEjrgBMy9KI74BaFkdAosfv3zFt2QWqBbKW/CKx4W7k/JAjhd9HBI0gfgL57Xo04VpIm
VBqPYMmpg7SsnV5cKU8fluX9nLpdK5oJdvXajmlk5P5eNrOHSHfzJXjaYCWNJzmKr3o2LRxwB1aG
LTvcfVJCO4IBrMF1GFaYgb/E7nbmE+WDlQLsB7piInMOfOEB2QUBE8O44n9PuHNgYqbWOJEI8ZYZ
x7OFoynGd9CTZj6pgyuiqFGfxMSTlgVEbbPqfqSNCWqfxyxAQ8kYYv1VLdEJFkh5Ub6CtwEJgQpp
2pUvzVidfiAm6sr2SgvZoe5BhwtzAdrTcpUyP6jNn4BcuYVFYN4mnv4gTl5eD+6Cb37sCfHYkxVF
ySajmg+cOpk8TVzjHoJJW6QgPgurI01ustS8JH8ojYgy5cLLqvx9lBjM4rn4GOYeq5mkV36YMmQV
lNQxn0SqvofYGpYp9TMTsDNbQZpf/mf0YHLdV+FyaLzcvChT2FYVgmgF5b5tXWE2ALyBi1CShAMB
htH35OpVvuggdluL1+K2zoh0bvt/4RzhFwKZSEIDOYAIRdxTFimuNFDifkhm4jpTi/Efz8rF5/FN
qsvRw4ZoNVkkWpNzmcAyrW372FXrgEgwAxgRJn57ig0Cq3vbdrzINX4WjzxEEufznd3ikrJIb4Dv
wZEgiFWz/tUNn3lFEyDZhptXvtY0CkCNOpuMMvhj4vOmz1bktZbuVL3TbL1PoWxbn7cd0eMTrQcd
0grf/Xfbki1AXvfHxyI9PKvlXBilhs+vLL4dRzqFrxFSgsnZtlk8mv2CwkE0rSr+bQgspihe/dCV
fENiBXCXb0bwmSSBuR92IunwWodlMyUhV7yA1iEUijS/LQMkYB3r8VXZAyRz+sJ2XCjX42brBTAY
8pS9I2UNOBOafcDK6P47Lw1Ua64Jac1aUkUHG+rWtVIhyq+juFurtcfpE8UkyhB5VkaUXaW/ofkg
Je/VGqCWOB7d6ecLmKD9NN4/o0exF4OC05n1Mn4ZhIrv3YMqN0Cpfc2q9iwNdY2F4anOKVo2EevL
+mDkMfS1oU8Nbu8QkB0Pbsp4Qu7gm8cGRcT67ojXKVUQRQmjdipqkW6CxK4rDu7+r5dtCa+RUIqx
h04YfoxTRImdFs3v6mu+FF5IprrUYk6qUrVUJQMZtWoqUYY1bepnOoaf8b8L1XstfcF/VJ/L5/Oc
v6HR6sLQj1smCire/M7uCXBsikispIYTxPJLl9hzGbsm1F9rz6QUStPAiMsnVGyEldPdTr2GoFab
RHkkbE6x8S+tdMzCzyN51t/PAGtdd9Y3n7aXoCHI2avGf57ovBKAxfADRnJ/zBCP3uLusu+oBbBi
dgnHKDMpP5g8ykzNJ3Ia9TfrKWKV6ks4B0zUadCmQG34IK2p9ueNmfRrMLnPllbyC91fjft0ImYI
xq/n8QjlwhMF/xRbwCtEh/m7taUbNpPenSsJqDsA9iLgS6EBCXqEgEFgUqQJYyf94B1caUB08rFT
f709+Na8+0gnA1sgl9rAOiY/EfY2IpAcj2yQvIpQ8Kno37rffOtIxGRUEDKMjn2s54uZNz+pwshc
d5agFDPz3VIHS5ItI+NIlkZmXRVKPUbz7ud4nKFeGHe+OVlTVSt8QYOqKKSca17RxXSSzq/I7lnq
d0v0YFnraRWylZj0r6vBAHUtve0XoQQdVFmXnWUTdQw9ISoKIRgbNSNurhHchWWRuMXnZoi3FhEr
KEbzujOTl+XQ3swRfe0InPX1tZV9/BTDCLaMYN59LI8ZZ5wFku0Q2gjWR/Hz6x3LlWuu+aUTa5JV
wN6Oe+TdXZB1G/4I4Q5UFr4x9sWHgTqJGRIU9PGQV694w7LE/L+T5AY4xwv93sSb5D2ELU/Ngljj
GBIFl2ZDCj+t57QPs5gNQF/0Tf4bQu81wZaQy/6BmsIuTfu/aETilaWNJ7EKQ0iHWFfG7GQpGX9w
jhhfaTWJ/T/gped07m+rnuZtlpZQNigiSt4RUqb464VY8HkdtdYw94zfrvPdy5+SiJ1ehNAwizO+
9e6LhCHox2WMr4nQ5MLJpNQADJi/nLNVNb3Q7oE3N1aWl+EpBwRFM/yvAEcNPez0Zm/R31S8tYgC
3iS0Pl2lIYul6YyIVaGxvrFXihXgqp9j4hQ50wPWtboma3i1oZjSE14VvHMDb7PPrwUrP3XtWxzv
9p8b52gFCU3ZLECZZ4YCnheosvgG517oerSuC8moVitI58Kz4yC+M6w2Aoj5KmhCEuiloOb2f3jL
L37NEksXwEk8tPQd0tlSLjNTCa8WkcmbUW2+d+Q8IsZP2Ayxv0AvijO8bSlrsCcqIzHVqL5U/hVD
vt7LlodFq5/ZZJqHL+YvGwmC1Tw8kcpzfFhr7XIGxPdKPdRnYbaB9CpbPhEs2+qTYE1GkDxXX79L
PBeTA5rVWIk17tUBaJO037GbydtEtn8ldAlk1qMjIqPX/IA2wbUN2ElwxGcCjkdy0GZQHOQ3Wgl2
gMY/mRfu1aaNxGFS6do2WJ6VcKSHPfVdukqxfaw9ur2EI2hg6/TJkfXMutLizObIEJVe1RgIkqDB
e2Nd7LQJq6xEOcf7q5NPZcIXZJ7pesaAiuj28T4hSd+yJM4GsHCDD1EqU9CS4yq5dndCAv03c6PB
DPXOHzmQRjSlyqfwl2qA2w8W2NFb/KjEMWWT95fb1VOTScYRI0m34MaDynrn7BXyZhR9uUwVWWlJ
U+3z7crxaVmJtxTc/4chdxL/7RhxTJBCV3a0TC8PLvbSs9hNFMYR3cu/GV+Jlgq+A5a4wVOuYp9O
UTl1m+ikwJvcningSAX8LgnCoR6kcvxQXY7JKf1kiVCeda+FdV+PUDgpZCLoEZxULO1wmFR30tlw
iGdPwbygsiaUhBX2TRArM+OByBj1fYm9nEho1BYHj+TgfYhRb9dAvsWkyb3ezhLGr86c2FbBUFpO
2KKHbw1pWOdepBW30fLPImyYP8qZaWyZuMfyOHO1Awo5YVG2I0KHlqrRXiWLNnZBhdSFg/LmdEf2
EGFm7/9cNooXRZfoWAwL5OvWiKYkPjfYUV5Xc9pTFo7fcHnPjOwl0UMxcZf/t/EoZZ+trAgrWVYS
h+SWAmjdrUGfe9nttFwRr410eSEMm4CUL1o7PHQIXRsV4HyzYt6lX6zCCb09B3MQOaU5TXl4EYrf
rymBCuHj7ySBCA8uXUQJnDKx/+wvMzS2b5M2Fir4fo+PkFKt3vT62DPfg1oQ1RXNPWvfmEQs8eak
WMkoXtTVYUhuG19fKLzoO+M2XNAHMfQMAPgwT81L2PdRF80I0ZSCy5gFjti+W5svN9P5C6i5ynjd
nXCFrOLKkcJEreI8bvOrlUEsPsgWYZLpzzlGBcS4LprIzwGWddu+6bANqZ4ttoN/hwa8LvDigmtX
GCopXV8liOkH/UH9q9R5HO1hBGLTDA61rKQ4zSWhkxXfjD2+AOjnU/XDaZS7WrLRQuoyOQoDG9ef
oC+rugyw/T7pdqAAZ4r0xYa09ksIxNiBvhIIg+yq94WJ9bZNA7dLht1BA7nM3/luXGP3uOkr3Z75
XUEJdgeRC1yMCZeuGeUQjBZUUdKvHyyKCos24/kZtSCCoFqmNlCGwnPdADqZZrbrZAdVdC1rMMHJ
saiiho+jsgDT+N0vp3OAMKPf96rqTS51O98ycY647bcXE7g96N+lzH1QuDWpKMukMRNFQUgojfHQ
c2WXqV6jc8KWP38xaCOAuA7CmLUZS2e+zabzHZuifQWlORc/+In4Jsj/tbYdCD0/0Y2auSJLkHkA
5BPukpMAziF8uNsrkb1DoirCQba4SUQCUa265RUrSx8FcMGhnoK7oU4MafFeB4KPN9uYaOaCe7l/
dv9wZ+ndpTQcljsUs75vuZcOhbERfqDugl7ohIFiVVxZQYNojZNod7bFazXbLLBcTykwA+OyUxuQ
zW7PKqaL+jcqKRkw89IqGRaVec4akdrBJNvbyry7BZRU89q63lIIR1Cp3XSswz6+/Sw68f7ehaBM
9vo3ag5INmLY+/IFE1QnkSf8OYdA6FjrqMee230eKnyS7TBm9DsRhWf7tr/dfue0p+qD9iGe5fMt
lD1ePDyzjGJnGllql3aOWOIW7ql0FdmeTIdz3KURpbJ3nT9vNvR0QIKKXwu2G0OfGJBp64lTZwlk
sDe868BQJeYKuZDsZW6lZUJ8gRARKy8TPEAEIsUYNTRFKM4V/ujbF+JZucnn/U4OXuSr48IXDemZ
OoZ6Y1E8lsTtaNDWnwWtb+oS8h/4v/vDblCLEWNsUiJIIz3w0qJR4raXXy3k5urd0nvwocDhMbAb
hf+uDGTDmpjIyX/lYc4DRNiw+6bdDWc1V5M9MIwXgEfgcwr/5ZirrpUwbijRwKArYuleltd8+Gaz
Fs49TKhs4ILuZ2rzraOQsqwiU1BsPgJjFQVlp4f2FuXjgig3iNORekr62GqD3akEnWfDeFyiWBsB
Ijw9aQN2fz+NuKhRxMDddOT+NMKuy13wUKUVb2KfRCF7bOSYoOZvKqA7iUrzrec50N2rdsFwynZH
dre+6FJ4fULqzqDm6nF+bVrfQmyxiVPyWZRTfZkmcgdO8U+yZ7RJPn7sxR5b4YxjR4nkAW9mh6CN
F6LFoZ3uaEZ8t9QAD4JtXNiyE0BvgCWBpc+HXVbIP3h9a7d1wHGtzgf1suLiLIdsfhWI+4ANaiJU
Q1ygnDkhYY5UhNvfxloVpkQ6jw9bj8l93OsFEGj+1y0rwA0WITExNaT/OHN0e0eNoFNpO0UzhSeq
E0PMj9EyYJfuzgy9RhutZYYwt6tRqv6AjaMiLml5cVUgR+P7RruPbPedX21qqFcAN0dja0+msWZ/
9u//UC3BTK9KHAgOYPsD1abYdsI97llOZoT5rPEmfZ0Um1LFeVlhAfNmmHMfGC9n1+eNGv4bxo6k
cJy8eojOs2Yji/CVzL+sK7c2fACFH7MtB9ySJA1UrTQhlSxcVyM8x0HOf2REUs0Cug2nAhTuJvWh
zFuy0HdgfmJVNQxEeXRd7sJE1c271GYFJJ8CIP2uXvSEtNTuyiUc5YXPVUJskxbco9aCkDX3ovEh
3D/v8bZs6H9GOa36Vl8dnICIpSFr/YWAO0k5ivrJyD88Ie24fdofWgzNB/exZoekKa/HR7SZ+6+w
fXbUoUE7BJRrsiTjoM3m3ShXaMJKcQI0RqkEtY8ljHAN7UTlM9OH/0ot1cjidmEMSsSXIIvzeLu+
/PiExK/wrWxwihK6orGQV+MNEz6Bsj9H+Ce4fh5zeJF9PFWPFkypPwhWj3mZj2z8hkRQWgOmv0I7
uDheUgOKjjA0J/e1iKd8l7GHUxoMXz6hV5coX7Av8npEoJgTH59dmm5Y4tWRvYhGpAzzd2iwkaDp
U2rz/OM/Buxy5stcKbDmbUj/GVsrI219znTEbT3vP492MzLbG390VVSNuqJ60W9ObOlFQr5oAM6m
kDeSZTpGzm2Xx5Ss6sM5jETIUguZwFaLOW7g2b+9beSv8gf8p8bAfQmGM3WN48zHcvExh+ZNJvbt
XV1jXPfELz/yXy52dQaXKyzb0zOCP6imG1ad6V0qoQtaIL6SRs89LLHoQTRoVWziR8RPfAluZqej
on631Q2K32UAXtx2DVHbD+kIlWpaDIcw1brl8Ykyj9HiTG33kqIvwymxNEdWg+27c/ugfA0TDyQC
IOyBNttpVdbTG1zSN5o6HE1hFXaFDcP26xLfjM7/DfEQ+MeVHj1UPOIRtHp8RSmBCxcpnQ1PgeVg
MNiYE6BG6k8S64nsiy7yRFvIgXtCHD2bVaWSQohUXwQKel9G+7+PLDFbgjYi19QJkLtdzEeXucsZ
vrKbxFlD3Up2v1kj1hoiGr9EVAYkbNVo6zPNGGTrrpQfe19o9uqg9JG5ocBvqviYhnlgMuDASib9
0h5BSlakwGs1oCWFctinUXaFVVWkZl57CE3RJ1lfefzatkSDYuHw/5dlfqvB23kq0fkm+EOeVq/R
aazSJIANsbsJKeMe2FAFSl0L+++30jNT9SYkdpmsXeeFiT1l/c3P41+738sIyKS6KFJmK+uIu64f
r1VEc6Si/inOYxIf/wDMyy6JpXtWuPVZKEfWGOvdjfqtxCycpBP6bKcoMvudlQwDaPdHmhe0l9gU
11i+zAAfDaRnasqPd14ELmHJUugNI9k0GQ6PW8zSp5WFt00E4ps8uUPCJiJSAef8FENlpGmoWF6Q
eSKY15USIXC9FdnGAm9U+/MUnOUOC83nzt3JRmC67GyNLb3F4gxTjfeZu3rMmb0IWj4AXb1XIGnx
XCHDmtVXEk8ziXX2HAzAw7zCjmb6vFy7MS1+Ne0C/BhZ/mzXZFfmS6AC7iCNmNMwgJkbU/5UucZV
svlljn9oq12E7JB4egrYm6FzMX5AdPccLFX/t6X57/jyCVmSZHWtSpUhJzGKhvmDQvcVaRnNGBz3
YW+LOACCZjdJNsiafj9TwQ+c0CSThO5asgOfrzXFEdy62rhn4pK318izZIdqy3gKWixixmp9slXs
Skd5jBv6BGiCL1T/+ryoJmOywZXPCNoZqRokU7O54U0RruFGlGKLQDmQcWmIwRv5F+zZy9AkKfDR
FxFZpVcAAnaot5tNtg5cfCtSHFeE4XlIJaNJ84+ln3FlBtHTs6rgBKtCUShRhExfRcC+6snrZExX
h6eWXUNsHjKSBNkJJTleTIQaFc4DsrwpLx4NkDIZGBaC7GxgCBagI+engZQbokGSClv/7qYbpIOO
jtknHjg3AdwtPJ7g8NyfCzCTF/PNjU9z16xPb70LBWGIl0GUnUgozAkBYMXWvhlVWqTB2Txtz4lD
vNoZEjYLZcnY595NQsow4h0tQIvIxqevhwYh/zzXBP0BzCNGEMFOp8tP9W6TS+L/uF+LPREaqTUA
Y4N8culAyR9BK7MF5Iz8EXBk8RXGXKi7LunpOy8krxckCtqpP4BRckweL/yVkbsd+fRkxUZXvAvH
Up+ku7kLAmGF5/2CbbNn4Gqx3+q2XCcVXeWRBsn+LNL9rl10sNi/XyzIpBYaWDLiMpdCJeX9sSsO
R1XqR4sHfKL7+mtPTgkJL9E1Mwz5KZDesfWqicRglWbDZyd4PZ+g4cBK89UmvLtV3nwqcNRIQuOQ
KLP0D5l/DWP22pT2WwSLytCA9i4FVgV8dKvUSS//udDDVbgkDrktEugNbkqwTIoKrWY6RVkWskk3
yM4VC1aByXoIvrTc95vEjWaeiQD/oCt1FhwVbejnBe0FbDmF8CXTGm0zVeit6mGsKIt+b8qaY4W7
rIojBtejjnevYHKDMja7hYaVrL6w7OrEugSnLiyptJHRpp5XT3st/ymvTVTGwWk+y/iROLodDlhw
dqSybv3uYJtwTAhioqwxOqh0QucbpmOrcgijGFRHlBuwdNLT55swSAEdB/H/WSz4M0fmCsQ05QOy
QkKfvcJ6ISZdAtVLAfA9zJhB5B3EZM7mLqBneG0+SC9J+EdDoCOargQUcJhTiFLe8I8SGH5SrDBt
URHBbCDVaMxYp3Kbw+eniO0i9+aeToZPl78fP3REruxsFNvbj1sWyFPFKkmew3bkFPrH4AM5+GDC
RvKAotwrzR41qsB51o0ern3N3gDk6j/sEdAWnR+bM82SlONf9ye9qMUdFHdMZ3UKvVONN12wqrRy
hfL9255jQfkxrADObzT5tU4utbtn+NrAAfzugAaGJcPwGUHuIT0o4fdesgUDLjAhy6iI97EsVFe4
OwGEgiBk3/x+LVv5XLHD/ta91nzvSzAQp5hyndzvOwkH5IeEyW9dU7qjWkBBfHTuqL6TtDOBrw77
6odtwLNLPNRY2HTw+qo1LirULXwDhnzpsBgho5cYz37aaA5qnIl8z6+5Q7QvgnzH6pq3UYI3DZ70
wruzapTZLoSeRNvSGYI78F1KuDURE4j+g4/LU7EavIEAXetR2ykoHVlCY5GvMXeuWyjfJhfybe9a
fhTR22nHG3DYhRsnjo8BYAUL5wlJWqydtG3au1Igmkp7k7nl2Am54PrBiOdgIUHUz2Thne9r5lw/
4d93qT2PydO5+d4ceHHHLuN0VFrqYXF7eCEyXGXsrAr6LSZoxiNCoaz3CXWW85wDXYLCpSjwN39S
baaU9q6+c+4rP94ZBCnzjdNcL16rZDZuI+dcRp97oX9no7RbyZl7yla+lDzCslQoDJI+fMbrY9e5
Yc0m6QDQXGN23TKh6GwWKyF/VujPxuGUXpUCBJKjJ4Vm03KNyK99H1ifrniW+1yJO/PLo0U/hm+a
IPRr+mrLo2kYw5iuYgcIFOSIATSM6kMZrLzyigud1u2nciDGnauRkhxXv3RvgCNeN/9mZJ0kvwvH
sF6W4GaS3rc31F8qFExTln1h9L/DUXAxr3BY2GS7xX6/MKGf9F4rS20hRg/ekl0Ls720zJ/O/QTx
U4fV493lWY47GOdnvRmVgEOLo1MD0OsSTAwGeDZhps7M6XQIQgLpuFpduLo2VTxyUgs8apGB6ZDh
PbqeeXVAhSzwcxQs1YtSa+PUnZ8xd2gFChXSQWYS4zF78o/LexSNn9lHihHN+kv5Prqa1JNE6VED
BUu/+IRMhG1MpHoFszBgBXmIOMY3urecrdI9m/dgOPtFFOlX4o9mZmezMnEadOdiKlYJ9VDhwLVz
l4JTYW4xB5x5myyqApRlawj2s5Ii5BlObVvIXY6Q2hNeEte1Liy4LzClYhh0xif6mAL/xjx7fka7
cPTvwr4cfp0R0gP2iBhkkEvO2BzEX3pdBipGU1nWSsH0CWsDH6apdWhNB5UmiePITwaWTUgV/LvY
cF00lJbU7SECRvSk6nx5WLVNgEp6H8Xpx8Fe/6eK43ErWTzxv9vebuKq8oquFuDESgyFF7aVz+OK
gqiZgiYNFb8yLtJVYR1GE9Pd9lG7EG0OK1tltizuv4uCxAPRSTCsBgB80i3luqVfgjQdD/SoC5LF
lLEA10SKxakSlK+ZrKtbaCxIXT6g4590g0gbz0vLDH8V8HMDB9zohO7dFO4rVMRmhX1AiQFmFzJ5
jbUMUIlqd8ye1supuBA6n5HnFEJCEXDBwzE+xDMbfvSLotgjH/zwqPzEPJrNl5SUgP17dTeTnupq
j+BOC409ckOqQ4sbGgfq/G3ioTeTs6T+2hhRGLGNkx4Nv71bQdGvnOsmg2RRJ0eNXLXnhZH/xwQl
CseDblkp8in9FSjeHKpMTvpYzIKMO4f7TWQfu759WKNHLT1wOe6slf33ZORtNkTMusGSVk92Q1v2
ZcWqZJzXp0yTDH1xEGFy1AWJw6OW9GMIxa+YAixRWN9mKrHENls7M//4h8hcp86S75rrfBkvFhqS
DBLx/+Slokgb4rUNM0YomL9BpwXdLx4HliAO02yu4Yh864GUn4ylHm3AunckIFPtVzHLbwQLhxXl
Dnn2aGrgPMGERrWQbc/ZChM+nMBv/9DN3j/TxMixM52LY1AkWSJQnvtVShLiLHxAR5wO8XDHcVyP
YvELbf7e0+1jdZtO1anBbUCLMY6PML9sFQZVRyfS//tbYg+vHzLtPqYm26q1lHm+BOqkFlG/U3RW
Lmqzg3LnMsMpfZFBKJWZR5VHBHuR3JWEjTpsdUN45ENBQ0dAQ5B9lIuF6qSe08hRe7VJgm8Z9WBQ
HSGUjW+wkPn9x2CNUeG+hG69cUkZIOQiwNyf496XUwzYI2q4950FrQgAsxOn7mYf0eryXjGDqUG1
cjQZmkt6zzrXIBeJJNZCjyJs5GQQlX9mIeNpdhP9KgjfdVi5A6U5d6h5xpzVxsp8aagmCRte1eCx
g7PDfWolQtQkhj2QF0Atb+y/rqSExBkrOSZNeCAXrq4WpjDlrZX1tcSuwkes6s+A5EOvThhYQfaQ
RGQ9lYzD5rV5PDfVeNs9nUk4DVVj97aN+Mko0rAaXHBWQQ0cxavHoP/7TU9QuWu49jXffK4W/HJQ
98focMT2SU4oNRCoCWNWAuoJYr8VSOVKrPV0zI2JOiv+q0hMSh3FKMI0NBs58+vPaWDLMgeZOreY
L/AkLqvPtzPlnxSRKb36it4cyucJyrtmPVNKr05DyFUXu39tHG8ipoK8YtJ3lzDnpF/pq8vbINIi
FYIEVCGjM464aSLjIpdcbtgcZLJiZUDiQQ7MeZOD9C4uZNRffI3qOATD1mUL+MGCumIp2cI/8FWO
j2mDsKEqV/z0oduwCSyOhLG27y/uvT12K1PuAKkzCxy8CzSKY5fSz4kAU5vh0ZNW7VMcrpIQ67aD
FOdTOmEuI7sFLzQdiaPgHQC5xoQ7VTz4BTuEbulM7RE6frYpo25Nq1OSBlAjEOpWvwOuVgC9B3W4
sjOsh2X15n22Gm0DKG1Dq3YASi/+zLYYS5hEg4aTSEmY82QxfOmuHQ2DFCDAQ9Ns+L4IUZCuSboq
itzZX/uDfGCqdr9oFG/A+yTpezO3fQoIg9WYSgDsn46sR6U5j3TQOKywKFLV3Vt6YHSQ5ipCNhMp
mj2cO/tM1yExN2sKUwxzYRQVJPd+C4HQl2Q9YcOHefs9VrIi59YYAJCmZiJLSoMglOQWUMj/xrl3
SLIqk6HVEUlvoaNNS/z0wMcBnG3KrUpw1AJAmsZZOccWCVHGh87yphFhFp2luttFBeKT+exF7g8/
VV7D50HavBI6WtdUH9SpKfXRrdYHC3DdTfda2FXWWiuov221O3aFBINC+30XDKcYEYRRrin8bOz9
Lpc676N4IZ8g8Uv6WbwfXuZaLiMVL7uNxbUbF8bwihkVm57wPpdP71OE85OuzIfvd3Ros/wpJnfz
zXkVTeBykD3Ia7hy+nePlPZMm+74jtboM1iQ37vClOj0bZclEi/F54WrGnscApMYNfPL5vTMuw7i
l0pwENdY9GVw0+wRgvXf9iwTReX7jPz8ok4vL+7YyuDSQNtaZLZ9AaX6Yj8Aa08WXu7jPjDG7GsD
adVLqTwv5vJwOr9aXWSfbv/szd9gDjJlw7ZUnO7HxHMJ9RLBac6LxykFQOOxTiKU78YTbSR+GZ2C
IX+3WKsO1NawqsFkpUd1T11rGdyNiUDVPu0xZimGA1s5lT7lmJ7hsJTiugijrB/SIsQQAArv+igs
oueK4RKspVNrT+5+ci/KzrMYqCsD5TCFUm6SVVwxxU04rDANDYfy3uK+6wp++SlcPWgYtBhJeGuc
XCOpHd4NTmVQ5zpyPyzwd2mEA3udrhYY8eqa2ochzeIGC7ZOao8rT1wVOAVkfE0tL85YliUZDWzX
a4fb/vDsBUKRfWZmVYpkzmdq8QQs/1y02DiadamzKuwNzcClBpRWY4Hk0Rn6UXpxF3IjokLg/1UF
R5AzxqKXcC+MEaJslhUuEysmYqCIVZnBy+80fxEi5Qls7Ob97rWCwasHpopjEo6RBiXj+sB4eyGk
OH36KJNw6FQaFGwhvPWc3EoOW00wVqZeX3PvmuovkU9YwWzSpY51JkFbPa2dKzDLkTu+LrkZVoN7
MoBJ7VZA/mYzSA2lCXz4lWyP/9JrUQu6XTkqwuYhrCVZiqAGPk3klKyCe5gnlmsEmHPGcALPOP5p
lGO/mwTgjW2jT2jprugsEkSP0rXRrtUFFLB6EPwufV3yes/10HzDsSkQOWECX1KdKmDL7c1hhLBj
ShTg2C5KdO0M7KE7ox1ML6EhvMlGaxwiVMfRJ20F7xTiUBv24eQpanTOByIZe7FXnKQJnr8plQVt
rAKnWPwW2mlDk04P5bWLiQJxpuTIhqxPlXne+Z86OWZIqRidOblHqfc3JXyEYQ6C4DpXVzoJV4zd
R/ILQqjflWLQlOGknauTYkm/U9y/R70Np8BsVolfO75pJXsIOBpVKZUPN2ddxr8OvyomC+0hUN7l
h7hnMrxLYTLmNTmnkp7oYAVw9/ohN2evODTal7SgQQckvGGvtAz8zwXi6Eauczr4pzqriP93f5oH
g920C2fm4h7lZHN4Z6C8EB6Z3i31N8jqhBYWclFYNTr+jzCFfb81E6wrx7uDjEu6gVecW0hyrYaQ
+wWLfDtGovnV0zxT7syECv3OUv8WIqvLHteKsO25jC05T0GJNIkRFjn0kYy1Alln9TaNiMN7qiRY
Pce6U31h6hXiFnMXPin4ZGhFm0McIMBWDlnR5QfcmqwS9DCo9DYTXFn3gFc34qiJRC8Swg++EOSO
zvV4EOWqVJJ79+xF6cExfgkXjiSbG/GI80EHXq3h0+7y3+TYbjgH/uzIasW6wVlz9yf7D+agI9uy
pAbFKB+kLGr13KHf8t1OZ/KLPwp1M096N5X0tZbMHxFShFfUDXkHhkEqs/L4TVaO+1/+vcQCeBBA
Rq7ggRVvBIYEtgnw77EB7wxpkmiXW2zF/lZkuZmI5um/wbKTvuzLFo68DJZiDxmfKnA9+7YGMVxi
aazO4bATgWKe5N6Fjte7nBrie3m/h5QJ8LKHhRURSOfk8fRjKz2axrHxHJExztGUcT7d0Vi666wo
1ZIx7fV0noB5EWIEeEyZNexmUMBRotLCY3iaVpQ9d2xIjAs0Ko3q2MLslw8Na/NMVj+CcfaeQ9HN
5RHH3gL/346+NXgk8iwzyMzkzne3q+0y9LSeuRoe3MfG04qbxzcjiSCQyGe6h/4PuKYfg5vXXo0c
PkKCO3IH2ECf5TF6ZFCFczaXXG+XK2k0btSgHHi/bfSwHdaBC8J4pwHpYGmdQDcMDYiM9j1x50Kl
146P44sgK//gMSe+Pu0Ft5JHhmoQnVfiTVJyi2aQ9of09+o/5Avql9OPJq8UyIdU0Pgo8zRWXrlR
LSZtxerzsBK7zouCyerQ4I9+WSTkpw4IeFfEfe5kS34tqXqsCAYzXGe6BNa9hBx7siuR277TAN6t
TxWNWw4pXrFaFWclWhbJvmZXXHuY5USSiALVzl5tqyAsjUGtNDR0oyuuIJP9r0qIhYiVDcg5wIZi
rgr38K025GAIW3kRHlZkb1BoaD07Ia7Dd/5UpyX8nYZbPBYXLD/RW7Yp/pcOaSmPfKRYbEkEgpMz
wG3ba2w/gbO+awrXbJMDQb/7KQ7YeJRQvvGpmDZQTMNg1CigTMchp6JK4q05S7LQX0zZ02IVtHXr
1Zt02O7w2N7wC1YwU5Z7b/5wsJME5agK6n5Xnvb8JnTK6CUYdSOIuNh4ozy/sSA6U63uVcYZEPgA
QA1h9y5TDPWIlfISRV9dlKD3padyqKiGWdWCb96CT7kPyaHwuRtFC7eWnd8XZg7+hEscrry7vex7
x2BLcmffm/PYgv9zyI4db8l2XTA7GcWKbKnYP6azGqHoTTb9LD7sQ8+y1Tq/XF0U9mSKc/h0mmN5
4rMaznsIzLzqyd4GuoHtxv0CU4NZWM53cBmphsj997+pbuOr5Lx0EiHRpL0yjMNjb/6xljKslUqq
niNGYQKZHxAw+xA8HzP3c5GeI7KY3BmhcRC6V4miJQzdPgAIhXCRvBgRwrnQ23CEUh0eJ1VWOcGH
tdAeE5srQBMI6L5Hj2hcIthm/1Jihq2X/delKEMSk1ENwQm2sOMXKSgShlPm07/bgSwkfHlIjVux
hmd13BV/878F29CzCA+mYc8fBFKU2QsgMbQ0MpLAEqk/joo7DbwBPlh0T1AQCFazwgKWckWtlTb8
8vNTXFdwfm2LF0KiTryVQZwO/j7z/VT6/KQbWUF6jql6Uf14XEQ73sYsq21suz2c2h9Us6opofGh
jckoNWPr3SNIA2GpqUtVt9G91/Yw/lBIyw86nwXAEO51/r1hU4mEhZQ0WBDd/K3Zz4GoaNx0juWE
9punlxr650BsiG7yV9eBut0uDtiEt1lPZDCWdHqzge+QmXo9OHAuG3BPaHh4xie8C9xwIbpu8QBc
vC5QHnr6kdOMOamYOk8cIM1OQbK/bfDwvvgbygmi6VI8lSDGvdQBMILrBOaCnfQXPj1h/Vn+tt6g
G9Aw5ZgJgqcDMT+RSxAln6xSez3tdHTmP5MbKFEL3sC9Tcs7rxjkw1JyiuQtmkmOClIcD6AEAN/D
VSsUOmq+q+Ho63Xdl1fiyAIMGub+7+XPc9x/68G8gAf9yCqIiLRTDvYHc5TWMkvmnGl1wJhhVxTD
LCNoGsc94+vOirztJhlWzqo/pDfs3kT6NWzbp6PwCMYg+Rj7g9NwkSeKIRpTglc5TMz4rh4HUBF3
1n5RaDqE4NZ7tdchLS9akoAQeJAGbmp4wv5sENNIF/dxLFZEuEnYajFx7Lqfwv7cIl3HpZv3mDiZ
9z4uQRVhAW3dYAAP3aMmwd1vFLPs72p6Sclbwozd3/AYWDZPYlfG9q/c74gwprCJQLExnubXJEMe
5gi6yg9guALJNRnIyrijnM72ypay9n3rRTpXoPfuCRt/c7A3eyBOz6S2D2wIdHqSogjlkw/QiqdS
Go8JZbm2LGc6VSXWGzMfwt2B1VIDNq4+wP3pVikr5drnb8cL/wEvaYUm0yLOzdKGQD5L59pvtHdw
7RVe7HMSlbfpGZRhFHD/lczz/vsPxr/twJ6YgB7uhZCBl5I8cIfFaMgPZKf5+uvLM1n7AAYRI1Sx
bXJvG03WbSGbCK+QIN8VrCNuUIKLwWD+9rJvMSTus1rAovaXCiOvpUgWQJeJ2UJ5yYnPep3Esnq2
WaOcGyge0CfWuUPQqC2kJZJuQAMfNTTpHjoHza+8wigAWSh/on3SZeGLzFfnxR30AIgQJyZJM4bb
dhVv+b/10YN6K6iEtAlXDWmbueBVb5a4EOHJKaN5OgRPBxjcSgts3kK54EaNgzu6/f7HwFjmyaui
QADkFG0cpRgAAOZLhIkuhUeeXjWFS9VC+VzKmUWNqRTt8cHnsQhA+qxULP+0+1ay9TFLoh/H4a17
Jh78tYdaLnmiYIRxNSaHXb+J2uzh8Bt9z0PsfPjWTWMaQ6iRPpntW7VgU92PydGtyM6LanPj8Skl
rDmPXrEGPY5pTtt10CWGzqt3DVO0WgZAnktu4A19kMguyH5/SwA8wJLppIwaAyRBP/fd/mh9haTr
m7lCoApYEFglbRelidAdrIIrTRhM6cD24r6gLp2yvTbkIUrgL9aVtNax7f0GxqOjd6AmwMl41vqw
EAcb/E/aqg8+7a+5AErOCw4h+GxLgzcMLDJQ8xkWiujNWPFJ23e+0A2SNoqHmVDYo7kOK3lNSWCm
ZOujCPMKneQducOOSqv+aybEEYc4x65oJDfFCthoe/8CYzxAp2amw6pWYeb6YfBgVetzOgnJ7ig7
pIiIJoagxkXgmnVKOjuF/0PckYrZkCiAX+NvtMopQzB+Se3hw0om5teZTUCpebVunWfVwST34Mzo
cFsrboVHS5kZsk4KRBz6w7RcvQUNokLIHKzjzKx7o3A6u+eEDMRwSzFLWpbmHx2gFT9JLWx7yecW
2XwfFr7TKlOmXTWEiQcPdyYyNlt48uTODi9UNsQkiXBQtVCIwU6VmFrwYOrocx+thIOVKlQJj2bc
kfmURm4RzAaP+SYsRE/eZHGBbCdi6I6eZAOXddeMA7xZfKyF/mGNgsjdLTtk89DERAYNff2D9yG3
8I5U8Mr+dsrXli7MWKV+AIxWvQCxiWMyHThTA7NKsdgq03C6oGWqqjCmbOTH6SmFo/G7QQpclhuv
oLWlEq9tsecIuiCgq9rO9oN27PIEHWfUHJK50rodFz4j5gGP3tqQz6h73MIVpU8k9AZzAKNw0qEf
tEcVGeFtg1SbwCDXFzUgJ9ZgzZ9ZgKsFyIDMwPnwbZpI1wTEpzgcpHGNmKtJjfrtR9YzLS248ggz
aV3qOoKYRyGzPjIHwMNrhAuDiWC67yeXxUheQNE0zl6sV1gdx05XryM08gJXjYvVBBmucokw1koQ
0rVT6JDSjEuH5+rfMh3fbY9X5MbLg8+0lwGr5/6/l/a7XuYUkVciHqlBEJTQQ/akIybLkmUf0Ghv
Xs+LaBQs+ZiInbzGrfo9tavrjR/Oyd187Vx+MqVx9AhVSokXeO3zi8ozE7A+ZblKNc4h/L2Chbms
18LOZEbLAEqN6M+mqtf0/xmj8eJm4hhbhgPBEckiz98GwD9mkGqq2jh9190f8ka8xu0wuuzEQcS+
F7fEjOgSJmAdi8w7TS0ZOfHsYswgNOmWG9eFegrbSWe01GCBQU/m7oxeJREsXjHMphnV86q+gEli
Ico0K69sGTTa050PiJ1L3R428/wKRfoGREdzARmOYORCN6QKWOuJPyPdilgtLe2k3cwIyH9SH0cn
TGvQqd7TKFsvH0NCEJfx125xfT3YQcB4YGlxMYVi51o0VyrxxAE9DnQq8Zx70afJWWl1BNebn8+4
vTYDIG0Jf2dpDCaGtQSk7ZX2AKBikYJtc1ZM7/8CG4psFcAB3VCRc9TaKAi1O0wp7Bw592gYH72Q
j5nj1oWMx0kcDv+IyaXTE3gvsO3j9aZlb5X0gwnHR8t0hWeLyiRJsActsA/Kwu8EYOkW0xRqnbM6
fH4Or7eM6U3CxhyYYSMbGAYoCcvsbHOpCMXBk1AYKEjsN0SWrwr0i1NMncDeWNwphG6YS4C1tlGv
MeCc5X5oJxOtdMEcNqRQuZPeYsH4lXRd6Kcwq5f93IWVTOReGk77zwj/oIRa/z25bR5MAddIS/+4
w3iXNL/p/Jq/CJO3nMNGxpm8jFNZESj7z/dWGzCv5qMdTTDVVqqKRoihODrRXAQoyeRH+Mr//F5X
dTwNtTsbe4PeEIkj74FFhNb9arGIbLAsmMAB3Q0cacctalm7And3cRP2muvSZwZQmtdArebHIkw1
EvOv/Da67sddQlgk2TcmYQDXUQ909b8CLoA0lCrk1sMnkvkk0gxYQLL4BelN08tuuxb0koUDVU+v
YvmDnHfQ+G4mkaHcG1Ft/m2Q+mEJt3JSvb1ypQHpyv6QWXyML8VoLSnD+9STQrphH84G0OCfOYxi
RgNV73Sw/Rb3VimnEaOIpe7v2+idV84a2AQiRwv1W2pelKz4j1+sAONrQ7SF0Tao6HxgumANRa6V
41oNpc6SNnokYsVm7CN+s3dVMRNZS9kTnm9srNTz3+GR/f+uWg+9ucYJ50kLfQVitAeBrQg1nMZ0
aYK/4iZH3FuwE3yS8R0XCNLjD1sfAm8zkr83r/gnUlegm4pdlAHuVGeB7rBjwvphPwmpXOqOtXlz
PUg9SFJxlYkgMrYf7HIREYZv1BqxsXorZju0URgaZetMy/nWgdlXoLdBP/A+iZZsjLo16tOww79L
9scymY+wd7Mh1T49vUIXfyV1YYI5AWVONfy+O10VJ9Rp0a0s0YvM4hVsZ9OD0ESVxe0pyXSheUyX
l0E9nzIVC0BSU0SNzAbZUmqYdROgfJjiN7gpj4ze+9aBk27Y1l9jl7tDskUiM2keqLFdeDIpVURC
hGANa7hrraVkrUlP8TBfFAPg7fv8SdxgGJaC3HD3CSFxMmaH3GkTobxLb8RfUzfk4kh//DetxXZF
qY0OfaDUMI8pcgW2nodb7alNJQ8lUHxaK3WmkDxPtoVss6pGLJM//uvi77wEn2M05mmLCMNc2Gw/
a6I/5hlP2d1EKe2MfgeNSesrTe7KpZhUl+M5gPJrjKLZ96XiGXoFtzloSVjPSLD4d+tvejRZl5jC
qHaiQiomHs+sb4UrFd0Qr8QLoIQiNXn+uCO4Ocx6eVHtdVwZvSFhkISNirc1sO3aEV9DLGIlPkFK
gARnEEyZIp/iDJfysvkgWieGv8T3J6mTugk6Z8BbMbXh3TYLTs01s9o/ujub1zcg+GnQ2WXeyA2x
ia09B1ibSZK2JaNWr1dKKTE7W+8fm5yYBILeavmjkVZvtzxhIB82TPKVmN5tXlx9kv2DZRp+Ve8+
i/XKwfJOEJ3Ie1YQJ+Ggx2pS/ot92AqxKoV7W9jMM1wydDMXANgFa/x6wIzVkWSp28o8HwJ0IpX/
3g03xV77Yq+KK2dgnv6vfW/qiOpuBwCPSBKIFfkm523wVJAFB3U/29UBJdswswU5N0wjDX3iEQjR
XQi1JDOwT6lWoNJbvwTSiTr+MW2+hrZwxqqSdz6KlxkU8tlxyI6eX5yNuCiPMcol7SiCieiHPa/M
fQS+UJPpWcY1IdZs3C+jsy0YPDW4oU3vzjmhaPzDIhpij0JZhjBzRGKMSV8LPXLR+JLzS0bRkjtd
8wnCln6GGm0CI9dTXXKpIZAxaDZ+iyh7uqJvCDsxy/vMSWcsqrByI7K9suq4t+D+6JGFbwI4zAVv
Esm13mPNEp2t9e2ayiEpfozARLQS6r77FfyHEHFmRZOGklxQEuCUqG3igGmZh1e9sl2ECDjMHvKO
TFAd1dgQh/IInoTVW5yIXxO7TayKoPMuLX7QgiJra54vpW6F7WasZGaRfMGRIMDPrv3FVhZiumSX
rxOiA0EPt8UvlQ9krAipvtYCLaP/tlb2mRcIgUUw6Lqn5Kc+Q8gu3FVpYGIPmdxIF1sBcYy2hszd
7YGFq9Ur/k/ZexpdU22Jb3cNo81tQBHf6K6HOGwcfWmatyeLcslPdsA+l6+tGimIrcUW5NWCSWn9
BcRSusToa261GdZ2pJV5e6bntZ4SbgwWGmIwEU7eOQ7o4889ZyPxdDNXOXGb21WWsfsr53KoutxN
If64/nZZs6LsoDWkmazvEeyT5gmZVKtK+49VFs5ig24mY/KfnCXipzoE3w+eoZkZRrWdPtU25RNQ
VW8GCeJ8tC4S8ItS/Yw6qOgGWEF8IieOIgtCqVDTvVuDVHd8qBAJTfuEZY5SHYSjq+O/memkViqg
Mo2QWyC3mmLuk2deGBCFW1nVYL1idlDxKkC37Z+W3US7iwfDDf0CJByXZfEYG1Bwa2cbYLQmTClv
/fJTfI423waQadAqyr+xNukG9KhJ7dR24oC22cljddfoxgo7F6l1OgTzi6cUBW435t2v+YrlY19v
FDJsGSGoRxMDE3HXAyP+Ny7n8P3rlf23DnDIshC13UJTtIVN+Q9JIFrIyoMruoiQV94GxN6qGlq+
AzLNrpN+WufDgOyplfqcV56GVFlItUwV+ozMlk35djA2pj0pQy/nV1iQyG0+7yhLHXMI2LWf7s9b
MA6cpfctHZ+ca+3mu28E66f8kgDQZwPFrPx+6rk9mavE69eoedyMk9G2QxBWznwsiLNVjflV1vUG
RQs877Wk1IlGGgKWDYR3EPZufcnXt+o0c2824Di4dy/cbfwa64yxhN2rpkzHZ8SEARM0w84Hc/4g
lJLPPQyQh56MFgbK/ZnuYzsH2Hfjbmvb/VQ+NPWttUxIML5at8md/NYHuAebfzUQsYvNXZ1JgUHW
Se1/GPrWikXHi8UAy0PqmtTsNcqMxvmqiS4xAFyG9DOPB1mSdO9TfOrGcszVy4w57+SgWdVLMoQy
AgYkEcPs5AO8Up4h/kh9EPUhxofAPuFE7vi9trNMtOk6ApS1JZiQyDfnpbP1h+IOM2VFDHTwR/pK
/r4GVqq1O7+40gc04fWb59F66ggvDQ2055JVRGRIgwxdsbIL5yAUHoCSZfTEPQom5eUohK1yBu4f
SR6EpXfQLyfXguJp770zvbH1tz0i42ZdWn68K0juCgtObdd+qSAioJ9DUSj7nwPdUq13jg7CCJzf
bqwghoIqlvodIgucuQfJ8jD8d9mh1Y/SepgEcLT1Zf8gOlklYtM1cBPKkenbcvcXnaCX3PRo/NNJ
vGzkb3Dq5z86R/7kySnpJszAF8P6evZE5yfoSwLbpBGZ4XDkHBFlQvrzpyXOrpDhzGAVai18yRKu
hoS29Mq6QR37TmOJiO2ec9oEfozzZd5AhtLEiJd6rcbRB5C7EZXEw7qTdFzFdJH4UkPrfEe2l0+W
1X42bjqkQiQyAuuRyfy5cFqzbGoihKWM3LDAYEwjBINmTOgPuXwZmppQ/1W2SIxPpeSk7Qjn4jHZ
dsBSOpq8WIRXyvVWsU18aQoW20L3CaEIvlvBINKoJMzrLRDQsuL0kBWXZaeU7g32FluRITIfLKWD
Ba/H45qRkGbCF9dd0+WFGjTdzeNvdWxx2jvzfPMX5UWGk9Yi412tnk96r6u1TRuykFKepWuA12UK
R5YsR/KwuK1oc7h07FQcuQwVex2oKKTV0vSyVma9RnEjz9BFvpCKnEKZ6xk8a4cvZsSa8HbMOhkz
v4meryrhKyTpAN3JTqGL+rAsF7WauEcYrREa57aA6cDDcRrjXUGbpTVY/qqMjibqn1sRfhVQo/Ko
kC+B9u3H54EgJ3tnUrRL9fYX6aj51xYOK8wZ0PVGCtxic8h0UQYvfkJm97TwM1PZCRDpTHjLh+4L
0kMwJ+J/RcpGT5JL2uPo1nOvhDM1wY0jwPYQe97pt21XEgHgDMkG00YAl1QcKTC6jE9Ecb9GcdYZ
DNpNgTHjxGlctcLLci44ie1P2ykEed5CSQ7pl20MXl9n3VE8aBg0foW4ojdhgDxWcB0PVsKZzZhu
l1tWW0PdCKM1QUcsghgDo7N8PyjlRPjF9IypN/gtuTzMUzO4fjDaRT8/+4GWebayxaDsvW6fsZiP
fe11bVj+1+Ydok+L0tkQLcWuHbChHmmlOdCCtzXkJ6vAKiQz74TkJ8itV3gbAdIJ5sYQ048D6L9I
e4OGhCeseD396CmdO/5ufvRT3mXcI1Ephu1DXtZGRu3irIvYAcgew6vW2+tLeAEaFmR+h1rmfBd2
jXTray/1KqVbtVPL5D0bZRbAvl/ejfzq+tyVXYlpzcrBguVyPioB/cQbvZ09ENE55CB7CF322DBj
qiwy2lvt2Vg7IzPEKjGdpy3eJ/xFHTqzOyl+HLRJSHtC/o5BqrtWj5UynYAGBB81NxP0oAyRUpIZ
G3HRvfuNVMmSKzMQSfSJ5E03QSfOpPSns7629R/JhUGuqJVIo6+kWZPcuylm45jX4mDFusuDPnZJ
iMUPsyeRnvDiMei9V73kyXDa6+TaLrvyKdS0Pio2hCshCtvmg5iO7Wo2qXYPIwiEgQdCRyBEocGM
fnjhioygEjNMRr3z7ilHYoBU8ti/yMe1wDWSJ+Zk+OXC4/Fq3bNaVIr8/Ka+nlfJIKR9l164AuKQ
JVhdLNxVweZRiGYsThHi9XSa+i6t0nb7V7BM+wBuHoYi9xSqK7xZir3PdB397X3ge6xxN3RRWl2j
cehY3OVk5zopsCgYC390pDXUlP41zvad9hcZ4moad3DWxgQF2Bdo5vuyo+j/6TU7o035+xGImi9B
q6/Cjv1Yu/KjJ6lA35qLUnTa1mukELp4zzhXsEWI9hp5csN6ySSZbba4K6S2Ov2TCq4Ygivcc+DH
dHNBMMqtNmFEtSJYn2n3tDpe3m2dhKpUSOASDHr4GcTkXfof5usglOdCmN+ABUBvsu9evO0GrHUn
KwntMQZ3LZKIihbj00vl5Yqcuy5YaetVU7SY7Y6fdX/sr9XxzlkY/c7UnJ10BQiqo/jWWFhskUDx
weSxGPJvAAUJUnt0YcGw9TeNCWpO+cyDFbPbuVuUVgmWB/df+BP2S5DqHfjVngjJOVMsG+V+R9oR
X1VQSM0U6gYKBYwlNYzqcyAckLNwSluwYXZcgBi1xGn8GbRy6Rs/RzvuZs/F525yoiaYASKDq7oS
ueif5N1QfDLA3cI+VyoTLnBEUDuuaiddxEB6Dse/wWNfenPfZ6rsi9rXEjAeBXzokXNmMkTuE8Ho
smCtTrBvXf54ZZm/4mPBz8UMndjNNz2ltF1DoyxP0XHqw8pJFqnHAR7Nq1UY4yJeeb8U0hkorpOk
adjS+DJf+9GCj1lXtWV74NS9z5ASCMXiPVbg33hUw52sI3FtckNHwwR24Ktu4Y6SrOCuq1bN4YUs
7L9NB2stKylBqRA9MSYtJ3DjrojDZCsMADBcFkdW99GPetM0oZF4guTQyAbsfIN+VxPIp/QYZoHJ
17bX1BlSYjUOxNYrYXsXLn+1OBfD24gbGoGffyGObzhCBKLpvYGDq2stKhogoWURM982qEUriTc7
BhxiYBsSRlcCXuTsxf94WrHwqwYFCEIhZvn7Id4RIfdQ8kPKtptzNg+UY3nZePkf72wRFKWOBVrV
/nYMXZ6Lsc72PAbTo90vcriCH+qx2iD8kN34PSGgP5W21xsuzjapiCVn1nRFSCLU23KfWXL1/Z5O
XTwzdljP/e/25kTJWv+XWK37X/ZUA8kH8YuyDVZMzKWC20GIRwnUMhfw/X+F0Y1Gl7xWi7xLW61c
qqSV1FofIcXbqggYYIxtqCpWLiMPowQ1FOAme7UgYMBCT56+aRjmD4iyriEtADdI/w5m2EL6tU4n
DigFfqXhHMg34xmQ9prXk8f7mL14MZMqXPMqYymoNcxPCHA3699Zr1N6i8Td7V0wqHhB+9fs1s1p
YPcFnEuAvL3U/2Bmlu4Fv6qle0ULGBb4U2fXLGiN2bd6RS6eUIIAG8uGEYNRJijbVcXhfzJWlqf+
k5iXOCFa5vq8BdGO/kOEtQip7Zje2hPK1m5uY1ktdkccoHYSe3zluTzIDQRMeVhlaQIKeZrR0nBw
w94ctWI89dcfUgn79/1s05p8po9lOFs+tAEl11cRNCk+pxcPVaj9v9jVa9pd5KYuqYujyp9SG16W
AbuUiOjE83V4nGZ9q7MKhQxK4GPSctWwqlC6B+Ysl8PiqShNKPwTa7Mjd8qWuz0fzjQSg1kPvRJq
ZpX6QudeO6eh6xjLmZ7v7jMS12Sh/ZwuRzYeYKMlt0uDhxd0H6Qx73sNjW88VjXVLfC67Lh9yFul
y8zRK4PnrX5KykadR2TvUVpsdvv2JVEywWSJw5oyUEYPBdPcALaJnW/iMQujjMi8+ft6J8vvzNeL
iY6YnzPV3jyMlFjSJImX0ztzpouxI80AkgpRhwNIGQeFjjeY2RdGK50Q3LYUlTYZ0DYoUqr5QhYf
rNQPA63DGqEIHsI2cGwPbZC1aevcT//9/qdnYkuE7lzunuhLcLdxJFU21I14Jwif8/SY6Se6N12Q
GdOMcpq03GT/7H4VjGYzeDyIUt4vUj/Bka7TLJKlGZRyJcCM3J/TD2jfYPQEfdg2pN3NmV2zCkr6
3ynWde57BSj5VIy6U4UcdqS82kVF2+kC8FPgS1ZtMbA0SqayTnpvogGkCL/1FsDnQWb8nLAkTWK5
Wv79MlB+MKrL85VTs1YThhsFdnFLiQ+RioUxi3JhLe4v45NYVqGB2miFTcTenH07LVRCNhZZH2BY
T0CAVqRdDvxyKo5bsVTMNdIygq/CLcJsoEQg4/sgLhL0BTelv5/HlXLzid+hwO9Q0TBjcHZ8ZUDO
RRmsaIvcQ8f380AmSzMp7HMWXiTaVnVvK8HBWjsMk50K6HCVy+y1Q0zhoxNapLMpwS89yAXPI64w
tGlS+vqrQSDI+RwvRLAPKmOQBlVVmgxhuygp71h0/g7rZHEvCK17okTPGl4WWjkSRge2YN15yhPN
k6va41cnSCz8jVK9E0m8P2WlFjsGIOl9rUcc4a5oZ2l578XZd6hCymCyp3V5p3FDwv2JtXwInaXY
cHoNE0vXWCtnoNieu/S2jKMkoz6gjzcVzkLQ2OjC7ZW1G4VvnxAZqOvklRDewJVEwLIWVjxL+X1K
fpqbaDsXAQlC5yUc+Fez7UnnkcKup7EpSv72A2Nb3z2q5NHReJq5GOKxL6YUKDb+AjIEQBmc+I+i
/de9WWTQ4WBUTXotunbTkDLUm2AJTg/JMggDYXvGbjg9itEn0cUXnB2QgVmUsK8f/VM0bNUtXqH3
3ymwiXmO8FQfLHprLlECQ7LdXcYqjL2X/Id6q8Rqg03kxOW1rsAfrX/ZQEARAFILKwkeCzKb86zC
Rm+eIl+tE5UEaPoHB7qJng7asjFkT8n06kwdeXMVOICLmmwH1JZceNfY32NCTHp5xQU21MEt/nk6
XaJnuduS9FHiIiz9xK39yo3RYJrSTsZ52mledxtlJ8YQjrFR1Z4Q+ULtAXbjwUCzBeuAbiZJO9rY
xFfqveomXuzWGmNwO/cEJiJvp981z0/MJ2TF/LsoSVR2OJ0yG1vbt2TiIkYiW71Yp7eUDoMYdfon
YGgkabg6vkbyTR6GRJYiME8dyYBR/EuO1MFkHhSuVmm3fk8lRvqnNtuX5vqNBE3jISoT4vuNC8tx
Ju5IfsUK3JJxl8pZhSeLACwZHYM0GN1k7/oJGefi+GDqJdOy26vWGAirYKy3t8Z1OrccMNzWz6U7
qOVakqXNojqk6Di1PqtEt4PBZDe/TVjlzUkOETlJQZHX203OuM6nEeIXhS3suGG8tO0oigegRDko
MU1lwnhwhNKhBSNYCuFJzSgLMjgpQdiH4qOrMOH13t56niaKt2sScF0FgugR21a6ZPxBYLD2Zfyn
zwoESSnGxk+Cq2B2yEHtOr3t8f1aAh7F6yv6hFvIsoFKFCYb8U9JKlNxaYVjHmhQO/xsikEW9T9P
LWj2JV+ZO8Ib0mpPIPxufpyi4SNG6h7sBrKZQzJWOqOTsWFtLMtL/hpEy1/DUBagfbzq8V0Gr7N1
5CmfhHgvvWzKmCJA67IaLwIHGbWF2ogNSNeiutDNWJ9gMrURAbTm4VfSFDqk240/DY9D61LsEi70
Vl96S46ZdX5k90uoY4EJseHTfBHa9wZDMPlHJgKiJ0XlQffyPb6oUgj34NtyEOHjX6yAzCQYaWSf
9rO0KRnZ01Uxtz/6Re0OLU8XN9lGr4+R3JoscA+CqEEc75fGL+FnJhGW1wguL7JCCv4HJLKHX598
N0aXO28Y62/PeKiIUah/FGgnywhZB1bWBBMl88Z0d+4poEt+noPDU9PDLW27CNOqJPWWzqstoQLh
e0OrRbTLavDOVVAhd67803hkHG+MJd6oNUg1hG58JLC4zl8HFJVt9VF1t9J5EReMFY1Z6NxnJKyd
kJ0c5hWVtP1HUVZXC81nyLczKYaeKpYLHGQmol/m/xj4cGKq/FI37SnL5VZ14O9hC9qVq1AJboPq
0K+rGzR1eJfrJvbFhQL+nM3Epsfp58j68QSUeOxPPyZJ3iFr1qaEDXJEUGlcL3MYdr7CtWRfLUgh
yn/gh4zlChqvbEiYyq0iRXFitRHHQfF2n8BGYDhPeWZeVdNme4IKhlJ/Y6zSYgLFdaWnRFFulzVt
i5Pb/0c2Z4UC7TTCWgGdWSRSkRFV1n8PNo862pgnvkxA69Vx1H8fu+K7JIQwf23XLwdMsPbvT4NG
c31+ivSVVQIdWfV+QZSRK12mQFwj15xgiBXtMTlFZcS5VNWCx2S5Jet+szCW46jdhPrMU3MrfFgW
O6cX4JUBOATzAh2u5jiP3ehyI/THl4G7Lq7gsUvsXKxkQHgEJbv9CSZ/J0Nz7SdcM73Z0B/GTj1i
Cu/yd/glE9wSPgSstNd2xtAm5CEKPdhZRowcUk+Nf+ggjCR5ZDZdaRzgsc9dasQaV66gTpwDt6Ti
0149dxv23wKZLFWDFvBEEc3j6XRB2dPeGNycVBuntkL2tliGPmCsaOB+81Xw30Dia9278KxeX1nX
pujHsTsTpLPEz0fZqZLepp7PyTqymf1kL6d1r/1zljVXefsw2JYmKWuIsf8zUxPvBgbF8bvevS1P
IzOsS7Oeoj2FrFDzLCvikr9y9623jhry/AX50iCcu+JKf199/KC/6rPFNtdpP/WPkb3ZCR/BMSfz
5Ma/viu3l6OLCPt8uyPTcG8jbfTUM9R9gkXci9Sf2iwGLtzzqTeLEUnuP1yQF1EbLi49jHPm+HMc
uJFw9IF300e+fcFUWvjjlLMjzmMdjl0bX6zowuHZ4DJmmCv4iGrqq3VtvHGCeA9eVemWw+lDEU6E
99bEoDj95pupaCnZrjEU7VsZgbkCk3FEUeGFus8rKlaHGlxkn+r6OsT3BYqjJ01IBJMjS1Q+n+0b
eTH0qgpkaEm+1Qn2qjB5S4TO2aMm8ZQjQeieKli0u0mpMiEDBlTp5lQBgNjX66/o7zLy3sLwCfQj
5DWdu4BICbD1ia4BIU6dlCDGHVSNQq0ZwJ0FSTv2oRfEO78TC2nkqZhPy84gUXONA+TW87fPVNEa
x0Q1LSbpVPEQKRBkPYUp+4zsMq4WKR2TJl8RSbjPsSQMfb7e1puu+VZ+TlIVXhHowOHtDR+0IE6m
bi+eAP6W2Nml6Aq1Htx5NfCpnrHd4qCiA20Gktidjavuc+35rC8A6S8pbNwIV/UONYikmdC/CX7z
8nR4qyl3ifqUhnkkSlbgbLYXpZEeA2h/SEdj83otZzYE3GjSXIewjA0Lq8yTrdKuxuK8q4gZfUXY
WG50lsKXMnK1FO9nr4VP+NXKUPPCwT9IdjUWawOe4tBaNycllw5W0TQIXiSY/dbxjkRSZCdUM+SA
C3SDTclkQikLTlIvmmRh4zbIgs71/zBrIlwr/15uTBdBOYvDYgB5QcgsVW3It8em4hDKT0kLEyVO
vKjAWqzkaHHGmeIDgbtwB2w3OnZi+vj5OQ37UbLyzPGzBrm6+FAki8MROTv2a5IhCN+7JCDQAFsK
cILbDpjlj5ykmSs8dGTBCPiAh8ZWtKDkXVoD819Awbs4xMeopqoukG4vOCgBnrv0T0C88Ci6owYb
EdBLFf6twH3NuDCTtEe0p9YVayrT5DoQ3oJ1OVzTDJ+LxdE4NQ8Htk6gC08+tt/Gb4e4tVdxW7mu
XotojjXc2XPmsEr0E7c50Fl1kAUa40oVu7SKUSph5oBug7Qd6LnkskwYMZlGGl/k9YIcEbKHHeIX
JenwxvF13ukpqeVXu0tdZCdhVFMG0Snoocy8FUd9zdYOZN3ccFSQK52J5rmktZYj08edYZM2JZha
3bTFWwiRI+A3DRTYzCItZtWserwpblnHuNZFunP4h8KCVy7bTlAJ6ztyv8FqLwCRFeLToVhTJT/N
xH9CF0+8kDizmToP1ejGla6tjrVlE9EwFnwMP4AoztoQxFq4wzLaksBKtl3urAho5PyriaUr7WTM
jDbLfTVZ9RcjZPro/sUKTmeRmPMftk507LvbKQv2tZOSVikQX0xb9mNaJotipWL90TMckMIjCdjb
skREB4OWNA0QF8HeoYPFO0vU5P18wnv6/qb35AtxbqWg4qcbguxJYL7d/6W6VOKYfSxaM7mARTzh
I+CL8yzMCiCcte/GnaP+gQCgywfSNNwnnEoRd6J2XP1Tm8K+GmWFfuCLcJnj0TG70SSE0UlWczR3
ZCnqhh1fPdtc+2iMDpRq6kaMwMGmXV3cJh9tO9zr6tfzY/MYMKb/fV/TkgR4vszXjfZEa3k/L5BN
7UNCKFah1RedCFLgV/Af2YyK2Dd2TAEjtRkmW57dy0kw5m8dhSAf+kBS4B3GX1szHdU6MUzyWk8z
nUluu18WW+6UZRMSut6Iu/rx9v5ygYuFI7BRbtxNncXwzjOoTIK/Q1jDYuzfAJ0XpTxNI8jxmZI9
pQmbYnvPwlK4RA8vH5FIUy4zPyniU29eRImp2bjlCCp2IffHv24/qutkK/R7YPLD+M1tyNpsij6j
ufpw1X5qkZsTYoq0h5bNYNiu8lTjZ8X9iMfkNN9WpleysjFloFvK/p0mvPixtZJbnuEuu3o1DzZf
vcLAl8nO6Mb3YdzH164ypPmMgi1DyQrkRU2F1BNbi87ZOsCJ9xP0QrDyY0ciGXfHswAuFF189LPE
yb3rc2+WBhdHvq6taAnyC+EEnKpXrniBgu5AS7XS5ajRAULkbVb9HRK6blAvPEbRaDKOZ96CWB/f
vaIAwy/V1USEjf+pOxsnjSGSwSzFCeyVc0yM47vU4wLRc4tW8C6uvKvzn0BssGlcUH4Otb+qDWIG
wEleNzTNJPceyNYlQYbUGKD6jFolEQSFt76wjMxKKgVRLfN49Zbe/D9Y9EBXMp3kjHEDMlbuNE2k
LHFBEUFswdtFxgFFOwz+e4we6AHto36+1a+nJulMSP6GvQbN1NQ6IlUIz664mkfKJjXH1dSp4mod
s/428sfthmqmeeCvrNfHOoiIZeu0x1o5LPZyw1zArBPHrju63SVIBlvHD7QO4JQsWdaT5yGcRy6W
wUybC57+1tVWIMZ3QRXf4H4LEJK3G9ngMfQtsK54rP8ocrovE1fwtPhhQVQ6umJHiT4t4KSL+/VY
lzcwb5jhxIVvk9ck047LewKwJSRpG+CZlUfwyKk46zgQKJWuU5PC4yP9H/6bVk8l6bMVftnCtCHu
1YMTwX/lwrJrcFBrdisXFIHqm/DyAQ3kKRcxbAylPXt8/1pLgV64GbOOewxS41agI8hLRoalv0gH
3QRnS7uSmx484RAuCutLkn+blNqrEkRQrXLtmZAFtyeFKMihzpi3S28O863Mgu9pYuEvG1v9vTDW
nUNyimLzcAGJwpXzKsVeKeZEDEyo/k1p6Wpo5DJhGnecnXRm9n1VZA1yZB6oyMZE5j61E9JEzuxt
8KmVbDtH/d9WOMWstBznDo1MnrINTqN44zhkgOxgOCpZfxaejaKgv2214SbbDv081ben90H8PwJh
ogq4/s8N+IOsKv2ck8XuWPl9g9DpdatMsSyvReadmlImIMELRlMtvFVd1GsB7nGlJvI01hk/2yTz
sTouRL8MLqC5byxB2Jd3QkafYtSX1tA/E3CB2YKZeUwRjG0GH9QbdSgcLS4E/nUZIlpipM66a278
stIXaWWEdoicV5u6R+8UQf/mTa+mSW5XI4mA5W4sh5ao8p7pGLyzZ25SIKrQJLZci/I8HKPi2k+s
v/pymlsCaAPK6ta+Ir9k2m+IMRiy6/q2wuKdIru+COLZYF53+ormmxEEE4edu03Dok6fmZ/boul4
TZ2osCgNfEzBAQSI0BZT1xS4hKFiyC8EHtdMMQ7J4DjJrpoA8ecfzaX4m+fMWBg0zSPgIi5vnwBX
epTsvIod1Ygz6OZyLma2YJ/zLdN9KEALoJO5JvMKNxHEzg96X/6EaK/hG7OrMNRPUYyw0EB/cEIp
bAQ5HGT6kcn9QQI5VR7EJ0Fv3o6AZ0QkgYH6hSXCD8f8dTzUw4H1YD9LwjEzBdPJrphvIp+NCPxe
STg03SG7dSRKCQJuRbku/WywuzTk4/BLs9QC6uQlCyRWy0x+JeGWG8d+2Ceg8K64E1B6kUbk2LHt
RZN5FyWuMwMCCP5Un3p3/XVSxCqEAU2psygYMflgBynRCLUOjXoCxSi28Sq4k/d9O52lc2kyTG9e
mQhhVektqFJHfB1AaCkp9lxdwS/8w+Oh9L/FgRoLG0zctfbs6kRxM8l6R6HRvtUtHWWmAJpKX3QP
LspWc8QePu9ey2vpQH7LUisZThWdxo1xzcRN8mp/LlCErTvtk9nYoMl4K8FfvOTppOt0SbtfBG41
U/xiODcodi99xeDxHyjuQqMxYUp4IDwpHtUMQ7QeOQbvnPgYL8gdZuQs8s+5FXIRC3rUh7vWIJY8
QEBr3WVbawhcuQ4KXMo9M1893cAV2CD7BXMP+paopDtc/3rI8punuDi46kDFqaL6gl6UQNJKAYEh
v9hkY/yKBbX99iKGXSMFlLoDOIGDPaYRApAhC+Mgm7gTGw4AUcfgfkV5PXcDdXYg9/YDL4JQQi9C
LL6jJVbQy6ayB4m043FoM1zH6pK3VWbbpC7OZ2PIwbN1f6yPc/o+xjynLM2pvbU97KP7/wECfjN9
sZfHUR1RabD/yQ1HhRiG1avvbzjB+j1sMgpun8cayHoSlXGc9qeimCshZU2/b4+E8wWc372JS5UX
EzZmoleyh5Mj7ssVDLoruhevRj2SP5Ter36PzJ0YnScHBekqjZPf18RwEd+d6fXiTYop+ukANI7w
phVPjD8fKudmj7KZzzhZ6k5dl0IqSgyyDWS9iy8lDYwSptXf4Tpnp5BQ9fVJY8twBawfbxxY/ZFp
spThj0T6i1i0sKXxVlHOBszfi2GxRRrsxjmUkNLDDUd5ZpOO1pkrVVHQ+Hj1Q/5OiuAhGvB8FV/Z
kSYURavouQcmDhUohFmww9mCvHXGfcuIqFSbE7YIZgQ/S7/4Z4qEbmFEb2IvZ5bUL96ZRVzrZxwH
zlgDHD1evejS4IpmyrC7MbRKLXABRVhjnmI31M4ihk5gpN77bBgywmgZ+8Ar1/ZTTRZE+IqsbaEO
CHOuym64FcAGGaF1K4rtMhz1XyysdwACNWu+gF8jMv2gCMZJb980l5kmDejzqDYDlgAOLnN0a93+
E8efM0ivusMqHcdqCWjF2tvGttiaFxDCxLqDYISc2JQ0ICmQq1ePC5Of/dj7zrd6TuPIlwn3KQFP
ygEgbg6/6qtYpOBZ6hN7da2/I81aNMXHmTGBhEnMiPqsnrmiEoxCdlxxFXKKUtSOq+wgpz15sF4m
zBr51srzcqHI6CqGF1nuHSuw0OKwW/mD4qs0GhlVuEFvzJMP4jEwvZ62aWuSBMZm9wT50PV550wq
+1MnUhSznAHkxc0BPhS0vVyfglPA9M4Rc3/H151SO+wY9UsfVCZK7qrFGWFZywDVorAKt3RHuRRP
wI8eCM10SwO09MWsvONz3fNl1wYKuak9AZ98bxv/oHGUOchDtBiViSO7mnzxR3B7xKpUWIsvS7y/
t+m1EFJRdl7zPRenF3eItdrZ93V17o9cPXT8Foh94MlS2l3i76W+nktj/CZMQ+swCwzVjRixE/ay
LeV2uyfY5bt+YP3VlCDgMIBH0NyCD0JHFQtb1NuK4UAchlpd6BqwaZKpAqVXQ+E7CQyD136OOKfV
7DjQDAuadE6Qtrvmm1D27ezsU7GVY1DjTi+esQVpdyTo9XhUSpJXOMdRozpx8z3QTt8y6x0whY0n
hsxDfwGr0lLQ00LgtsZdl3nXjbhnId5NwUvzwdXxNVzd0j3pzYuvCzgbmMOwDyMC2k8EzJynxifT
J9a8KQQomn7yCApherakDHwM3sE6B0Up+sr1t+cDWyQF/FHIWTAx4fQom2rfiLDUOJsn00MRKev/
gHqIVm7vBwXr+0AnOZkQWDpvC+47iXPPkeS6rosn30eKfMBrPhR0GnKZPvqRbYLEvpyVHbv+b7WH
mmJq4mLl8R80ZNn+QJmtJQiHtkKCrrVqmhOvu5wTJJU3D49zvL2hJTMMPUDt9uSjVfaVqsv+mjvR
+NkckDjNERxJhV0T/A69OtvbeI2HxvPuzxxBWynbYaQzB6gU27Mud+Kn/9W51Hrb4gLRe4J1y/Yb
yDRbYbAmwloM746yqS2fSZ9+++TW+DdHJTDRCTbIr5/Ufa7mlNibHciT1xhGmVseGYlmDqO9EnzL
tXzipYwRPF36L99AURdhvwG1EoVNZXi9IDZ4Xf56HGmpVmNf/NlLlqiS6jxNvsmX5XivrKPSKfEE
wwuXHR+JLyKA1iofiwm4V7vfiXhpEuUWlyomoPAOjtJfUs+Aw5s6D36nRepy1zVMTZHZf1XZNq/J
bOa8r8A2eGjKKVWaoNuA2oTmm4GAh6StxSG4sQZHmSxe8hxqSd8UDqwZIjOosA82qyqOt6SFYw27
Ht6LmOQL7y1kkdooNLK8koocFmxF7a5ppmOs9x4klSv1El710bwQbV42GouM29a7yAVmZ5BJPOua
1ulbrsqbv/h63LaYvgFANOF/T9G75Tn9q+h8G0eJJPh+5nMUIAi3Z4cc3+Z15gPf77Lbt2u8UQaq
gwReohnBhLYqG2lFgjJn7QlNusU2XpxwAnZY+iCSdKdf6HVH0l5opOykCCMkJkBTKnV0T63lnnI2
J++GycwKdbw7oaOQRo8vBx16DI3EhLG51XvGt7Ihl0OmZNWbgsSNGCttD0D8Yadj9ggRlZtPqdqS
DuIK9hm5ItO+blyyL38NyjkmjtTr4p00V6eRdXpoAE5+nAtV5Mg9x+HG7YEJvZwXwAA3uEyybHWn
Ux9y6zwDQvBgSulxLmPYwTxQXuyp2a8/JeYfeVnLT2LREnVMvbny0t/EZ6qXF2wFNTfj+L3/Q+lK
CL7FQOMiRQiB92x9Pa1MnJ0QS7K10I4wC71kRoj8fyEUHu7Js7Rvyh20NzEDuOSiMwb0QjiV/0Ry
b5d4IToHCPuoUxMZsYoyZZy5B9siS51maOPi6mL0iwpB1/cRE31KFvsIWCoVtj9ofNgbkzf0cQqe
luj1G3A0okP531A4wtNEIipcF+7jLr252IMlaraZxt+OLBFEMyzkQA5dyACICCRrCg0KvuD+jBYx
kvPcM8/6Ls9Xxqs83p9rPYfJUHGAy4om0gcq+OlyfE/JtLkVVwjiswvpoRj0EaUZT6c1CNZbd9Lz
bWYiEA9bHW0v5PMYl0LAo05pptTSTVDADpUb3+vWwAceQ64j4BWJEYWhgP+HRWlrPHPGewo0/gG6
6+m3yi85198H4PcZSRnyrt33ixnkB1oPjL5dLlFL6IoSUjw8y2UZH9dbzfDi5T+qWOOW2+KUb+rV
2nhdKk1frOcokZpS8dRVF3STVB4f/PFVEPImwA9rMwZMGYsAwz55ToGEsykK7+LDvBHIKD6VqYD/
6yYGTXfJn8kQdPe6cAkrBd8HpVvhQhCisb1Dcn18rn9VPR/M1591q2L2mjdgRP5/ZAhRvnYgOZPJ
pzd9/XPMzP9uqkOxQ3PEEKmVyq42HXLVcbBmAH1Fzu5AKoRsWM+i2bJtTA6WJzuymAnyM8N4smMS
8nb7+lupcrikHdSDDZUj6MtexD+iDHGjtC1Izy6XpO5+zki/Y6lXYuN0KRbHZdOykK+arwQBjgab
aUz1ohUFQ9Xm1xNGwZdYMYNwyaSQQCtMIVFnG96hY/gWb7p+Azgr/mj/ACThLsC7F591U3iQdTtO
eGkLmviUwe1wdVHtwAvXVs5UvHLLS35uN/91YiOPcKtEm5XJ+gNk7GU2VOWRgtikP/dDXsyOKoHf
NoQ0SQn9aeeHKuXZW3thi27kVNJcsVd1OoiP2tfKlS9jnFyGTH0lNDwIbUKxlzqET6i+3L5cEgaw
Wmg4yLobDBARxm9j/h0W+9fJQ5nPYR7G9zllIxL8Qqjfa+YMvi4dtTjH9mhFu32gaAF7h4h9lSOs
rstyAtN3V6ipAVTSzgOLiCb7D7Ul60alI7rdOCUUfqH4zR3bmzDcI/AXOOAHhsrJ/c/BRd7er68J
vdNj7BaIkWzTZLk0Mp4+K6ZKraa9G4M/cXHkFWP0qzgHdvjFaBNkOFloJfVdhHMluI4tJHMsxlBt
/l2978kLRtlBToLFZTQ3iROQRVRa4NXjp0Fbonb/eKOHo7GE4dKhcZjHB562YErMvHHiKLJRKCBu
qBDYYqNYtmpO5a2YgIV/+JT+tN+KKRESyh0QEuUVp0rpZn/44FYjHLvZ9PGOmI27LNZCOKiYTwnT
1ot87k9TxvpsLyXQG07ysi+0TE1aJtdlKl2Sqjr3sUhid+LrP1DPXPXZCIIQ68Nwf/JP8P+uq8RX
6BlrCKxeskXQQqhFJaK9r68KbWBomwlb6w26y/aqHBs/AqttP+Niznk5bfd8UGcNy8v8QBANCVxT
tIyqMBn15lRtkJ1/3vVd1UPTIeaTcd8sNKSnbsL7IjpcXEeJOjfpTpcLZe8VcaXGQcY1fX4NjxAd
rgCZieZBYNbIVsQNC/vTUNuEHrsQAv17E9TciTNAQLxbBdJ3uZr5nUuePtZ4QUgZcBag1CexG3Z1
HG/cfXp76ugwiO1aEJwZ0Ta5Fudi7eR1hSX+XeejmquhAuWVvPKN2kZPi9omXYINFOmwZdM+mi0f
zizd4oS6aKkcutvWwy250oFx1GbMeq9mPDys02A201RGbXLqERhFAimAkB3+Ul6HzCUyun1Mw4t0
AR7e+1Cdp1YwIGAuqeqefhB+eUrxLwEkgqfDoEf/uij82onAyYatgWscrk6cCJ5iWbEQGpChs1+r
BCcEZRoWcNLdLttGHBThsE5MfDMEPtyOVX33hHr5NyC8ZmLzKQWFGLHtwpCKi7vD5cCxL60qoYVZ
sOoI1NzNcRepht4N8STLY3nVvXEjMMxGBDHeoOZtsSjZI0F9dqbLhlO8sIR1Bvj3gyMUWz2frOTh
DmRyq/+gKFLhZl7FFcze0mDoSwNqJCVjw1QXspdJYUiBvTyXwEyIvwxS1UzF89Pir+PzCb5xdDc5
pHWUOmKm+kANOhorXO46fS9UcIUrsKa6stfaQFIxNQmHASlBMgRIQAJwL2k5d2nsbG+E/cjl90fT
zpp1wGlQmA8sbTuyj7LmP/vdqy/TYhaQA6HCTXMFIqGXEBEGgC031WS4805pc92RyngcJRrRhfPc
naRJgxaEmNTG6EAhIgKPwK4TkwSJlWzbdt2JI+jmLK/u65Maw5FQe4DJ2CtI+ie+AQqUj259S5zp
iBBRL8QHIhBkwFP0iKHSojO1wPDMs9LcMEYLTjRw+KTMzzMvtypxlkAuGL2ZBItPEimKvJLr29p/
UHXV7TE9ZSxx4BcQcv+oh6bPKcW+53rrXt7XPNjqkFk0KC5nbMV7Xmh/mnH1MsmIreHfU3NV7dTb
ShM+upvl9+qKlpdnU4bIi/AmTG1J4mlUv3QTeltymDxpJXduCSlLJ1kD7w+j5CnbbOreP5Ipktxh
EekcoHm3hRQc6uuzm4jQ3/ULSp6VK5HLzTZtaifl1pbyWggx0cYsoG3x1VhHce2hyrTcofKtQMOX
O/OP9vdKT9CVNF6K+PCkqvYQHW1mTz+7lBd2PU/8oZ7Ivg8GvdvPxUu1TxaFj+KiH4/cuxp2QH4M
IfX8wrq7lEqHfFgo2jmvCoKgQzx6+w078i7QhBrDw0Q9FaO4grwlijq5DUBgmvCScyeG9HBY5BLw
D6oEh3V/RHEIxzNzMuOa3VXkZ5IdjszjUXJCqqQoMBfN3zkd+3AvUXviuvN5QgL6HkABeNMsr34B
qVaaQus1bUn9yJftXFU53W1Rrbv8WHi+3O9kIq1lTvMueKV3tbPvZqTGAioWMfLPYybtKUiMqk8k
Ls4tO/pJxOY3ccDMpUaLsEgPOqIYYE9rMKYxjPosfQJcNKOqkysrUP+s2r9bnPrc26CquGsmiCvF
zX2Ig4NI/orQyYpmPMj3+84YFxuqFQ5NEaWMmuhXLkNwFR/vb2M95K/p6o/lc636SISziISKg8nA
DwyHbQ42TAMKz2zvZ06fniEfN2RR+NZGvLeC+OCK3PWx7Spy0joW81kMAQOLtuX5YlmhFP0mUCfo
RTgKkCl0CjM1m9MFC9GMUMWqPnGs3IWBje4lz3clOKtCPMKCWQr5z4NXZ/MCBYhQVokXAcstBMAw
esH83tAeRf6UImN/oSzrjcuD2W3rcr4dlHjQdfE9BiUucbfyW02L1MEcun0BRfb/ILmj5717PV37
iIdZ1uRUZrxarAY1ixJtUG/5p3p5Kl9xscXc7LlfR2q2Qqg1rb/0fPyonBTT7GK6ovczw27PdfOF
8YdG9pUYLc8xdAAmww19KdRCe0nc2Z8Z/A4QmyYCE2bIAp60e+ZrbFwtMGTKrj/fuNgmVOA5YSg+
dORtXgmxHl0PVAuADpSUBqrxNIJhk6YikiwSnD3Xs733ZiDaooZDZ5jZqOsQDg+tkajdeAMP11Zr
RXWNOJ6sd10EI6cgbuTPbpR03h2M+GjJXi7QFApJ2xVpCSCRiu03TQuHvct5V8IBUXAPGHFn8Xah
drOIXX1wUbUV6G71gwUcmmEekX+aSz47a6bCYHIRDbvT3vXntmch+WeqhJs8w0h38gTVTS//mXKu
q1i8E222FmHWy8kB+z6JNXzTLKj+zT6D9n7FajWii6a+CN8Ou9LT4lXHqV+lLk7sbt35EToKymsW
mv9d/zm3MFUVppr/oUaiN81ezVM88ZDDzKlg7IvNZU+vN+fWDX9G8IaB53p5XWef6KMSbQFJYQug
1lt/jb2ldOy8dwgI13Ql0ay/vRQntTI3AXhKj7ql+yj0JDAZnJZ/Mv8r6Ud0u4y2MNDSyXeQ+vi8
q23yxtB9EynmhmAZ9VTaPxqv11cl/Z7EuBRtHQExHrUes4EO6nxCfxQzt1kmklWDWHYta29Sr1KN
QCdmm6B9b/JOKqtySCp9VaI9wYLtXjMp02XJPkKM1fbi/SVHjGXQIPnsd8xJi0em4qKHP7I5PVYP
07NH9DlZTA/D3ydK8s+wYNjOOqmgJ1z5zL7cttXY7Myh0M1Tf1t7BKhYPn048PSDET+syO9wIQhy
xZdFvdt5arImtN+Zq3pNIgF/G8k4gWRQV4cbRtUYwrt8v0IxO4DpMKDx1S1DaR6nOwhOqcBI+IcS
HcYdKpp88482iGxlJ8CAUGN4D8BWcdyOctVX14p6DR20YdoyWYiaPoeTi3HOnNSh9wkAgibBQAXQ
O1gGlX+ISSXKqA8JXO1wDKiG25HruEKrDdfX/vVuAYGEUTciItwOJSHNCd4Oi5m4kqiKsdr0usoN
0klmd4EVRzPuKmwMnD5AMz8Sd5CyBA2MbilX1mYoPbLwUpUONyiMmd+BHLMW5wCIXrqfeHQz5wMo
e/kgeDgGRTQkNvDEy0DpwIDPQ7GB+qW3Ew9dUSju/3QE5/4eP/thYLQRbXk+vl7boA0kw4axfOgf
7LH/UT0z7Jq1HCkHjP8T7lNuAaOi8862MkexTLTEjR8cXGzn+GlxaSB/l9PcrteKES1KV6f/B6cn
bXSFfaSGx7e3kABZW7Yuc0pG2mgiy/EIgZWydwlNh2gNUHmbC6RAbYp9USvhgVb3+GdI2uO3HysA
/KQHK4TMaFwqC1Y9dnl9mO5QzmW4tjrebg98DZUc+xGENYLpP18sF8DQyUanRPXTRMdCOyFt/4yr
/zJ3qCPByexZL44K28prRa+RP5M3lk169GOWybUhSq+oPCkz0EgUcSqr92JXw4JL0g1ZmcX068G3
IB38iCmU/lEibAllMWzBHGOTXrXRhqUz2rf/Md9LKZVB4FxqlFJS4H29IzfoMD9BHRDR7F9ugE6w
dBwg0JqPTftC1uq/SH5m5ss116CZo0fPgnOk5Y4VhS+OJVbTyXluid4ICNqjHs+6JFTxluZtEMtO
4bjUJj0gRgX5CmaBRc+4RLvewnBdix5TzcdSc5iXPwUk71KGG6VsBkI1TdBqUwJD8U3Y2LF+B46w
7FiAJtwmeeml9AGP9tdkLN4ZhJik0aCG5zEZn7xiUCsxRDIz8DMpRtGGwak6zD9VVM+g25UlEr7v
XPDU+PLcuqDYW+esxuU22m9WPgPEKnjl3KnzZtKxWn0Py++i+Qo0i3E/ylc0a/hQU/DS8MEllWHQ
JVg4hD808yjZj1bbjmNCh4LGGyeEqAm0Om3RuCp6WUceVH5nKeWdnB3ItMAVS8/40BPfMGywVzSp
RW+gAEOCkmsvWCFhUcxlvhhGyrazaSySoTL9ZFb/HTdueIVLRTNY9WlVTZk444WGsqJEt3cRylFy
mtJzeIYxx/z1p/cqq5kIech2nHQGlIOY2pTHouxzpC/HzUoF11RmJCywJk9knXdZ3h5UVgV+EClu
fETg7kU0WCyz5ETVL4769j4eO3BjO/hYKiD4BlCsirTuz/B3G6+6HcfYbesprjH3RnSvJCFJsrUx
ZsuJX054HNKdlgvfsp+IEXaFKrz5giWUqqImr2p7zHTY6rhcUeZklighEXdqWNyuzQyoh07877UN
Coy8910WbFd+agG+36qrQeo5yv0SNPsGEiXMydMUMzKzttYOS7RsR776++sagyN/ZqOhKTCorlyF
4A40F8MIhow5TBHkTHscXKel3xh0Zc6XAyb6bt2upeeyIb9D0dvj8H3wtB1YhnpDb5A2ppnBYZUu
Hm8DcpZtjx1OEr9mOjWuMmSawDK+vyIS73nyH16LaavExBR1By509KGdNlfqvGfegLAc9lBpxKDy
hFE/I6fH5PdGoVDpX8/VoCXEqqE6tI3oW6e3/JZbIQ3HSv7kl1owy6EVNtCfj+Yx9xvQ3g/KZz8H
eigQIjYOXHRMy6/865MJEFDHkOiGiAmSz8gDRaujT8wieN4eb7kfR0oipJ/kblQKN1a24kZaL6J6
/1D/6xDbvShKeNsnS5vmu1lt1mCYzX7oM2lIlUbWyOtapR1gWO+1nQCqKUHhrvyVdK/+xKVfqZX6
oXcPd6Hl2EPb6VdYxTvt2/IcJjSZqQOWnkEmFwBRhzIl3xaDFYv6FW220Xk9pT2iPazb49b9gFAE
u9wNVCHHilseCS+3wblEbvNOuIrACHDM6Yc5Cb36Yu3mVneVUB1+JXGUiHqp9c/6/8CSq5Y40MuG
eJjJVB9dXdyUJ0kxmeWjDp2g20Z1novgGkJukzhtX/OmwvGzSgWwGnSFS3njhA99aDKNoWTG5U55
Cjj+xaoOFhXkmzvKrLooRIhDcf/4cKkQ2jsrGuS3ho6Pk86rcM9X9mxKVCvDdUj7pg6ScA6tiB1u
B0UsOZ0AqFHdiqwntLc9TL28lFhzw/XKig3FYhaH+jE4J31P0dJUc5NHaxU3UsCNnBuL1bpXtcxN
PcD8Fo889ln1V3/Eha3Mi6d0w8BoTsH0Foea5OGww16yk0wxijGLc2+86lFK+Cao9u1zHewfKZLE
OfSrhxVQcNPRXJk7vAkom9PMoCXHWz7JQuMnfWnbs2Bi0AHbJNFQMgrbsp9soJiSt1eHmOxUiswF
Nd3wnVd6/f1VV1SSRpzBSt2NG+xaEYYNNgYppXbQeC9NjK/1v17J6vE4Nrd+9LndMePHokf41jBT
dIL0KELq5lbUwqDC6VLptR55A9d3ZKI6aKTVVO18zjrNqVNFpsn5gIw9NIiJtTAlFv8L0/aM8cLQ
RAlN0TvcF2aCyJzRUp4NvW2tRxiClOLez+m2BqsX/e+IIkRUudtd0h85sP+W2ZVZaI2ieHgQ61mr
0gOrDALEqza/JQ0TlQV8bTSIeEFyyXGSmMW/qleehYwTC8Gzw7Q2+0Q1CaJwIYk5xgL3Zg0VVSXC
s4j1m7/3WsV0pFiMK0N1jzU0luEyQywaiY3eefGhegYbbRY6TI1D8Ntnnz3XS/jRyBXzsTyI111A
VikNMYNgct/brvW3M4S5VXkwWI2FIGeNCDWGQ1eDR9pBH9iXPoKc8r8iAJUW40IKTOPvdtmDLkl6
4LYJmIHMWDgOQgNSXqfQ+yRcFPwGeG38GwRQpjQiX2r5im2XwRk5LSMC1XwIW5z/dtsgS7MofOti
xf7eh/SyQQEdbP5KztcvZH5Z+ny+XAOn4+TFS8kj2mxj6QVP0ftmLV7zzygfMV0TtuZLoABRiQLX
dL0KvwhDInULCCvyG0B9RNfR+IxDlg/dqAomX/ALYnaXxlQoI8Yqwh6EcaVx26b4vSm5C3ahNo7v
2KBachuxCIC3+MHQc1TeMptiNforoDXt2O7uaTV+nYQhGwQI0gZxsHraDNU+HJydrGrExwsiotQt
fOkIfFyVit+2fIB9AkBPm83rwGnRvUf1x3w/B0YPzfjts/1T5t3PNdoZf9rJJJ32Z/Pzjkqim4oB
4BeDN/LLZI1gB33QV/kowOMLd31o1IYN2XqbUh2dpWlFjH/eyxpztNcJ7rlSARS16DpSRSY43NxQ
hKGxAD54nxumdTPrTxUi+BfHzeUxeaqHFGpJOWv8O/hvWCYQNC0zxc2iG78MQiP44ZASQ5xUUbHN
a1IMDnELhhv2kQVXTdU+fELe0yEG7Yv1xwOJKbtINheg9Lz+jUk4PpvwvzmNeSarjPXkhDvEQewP
kdDR5XupQjU6EkzJ55DRH/S6c85KwaMfGPIQ7z93N1sVbWMdbZBiRWpNmeUMWSDqLf4NxdXRd6SB
0SSdNMNBb1vfIZ/JmDuaQoOnNV9bYouUJZwS7igcHH5u9oqr1iQiFNsn2SSl8o43BX+IUcOEjgkk
9PJtXKAegfOD+2izSO6PUUikIzOCvG/x3lHt/5Q+m+YMb7DSYzH4fosseDn7SMD1oi8N8gXxQBlG
QBqn+Ww/RpwEEFFLIf/pE/trkAADhqv3FDMgEVYDYHcfZZEb2erp6kFufBD+l5Yz/tB5pI5JwHlD
znCRHtwEjuuNxfrHcsk8k5JS63kuFFoDKC4tMrQyPwNXxxTTs+EDHrQbaqV816NHkFudo3uqwWDY
vPjOe/MvnWUliaDDtdWbJWQp2vsViqCxPSOmaPsSaQpumWUpN9rXuVb1GxxrG7h2hPbmt0SwEzBC
0Bber//FEjWQenyUSSUJ72awhMPlScSZf3Ktz6LHgYc4N0hCMlXtApzuKmRT5xTN6cQy8cruqTC2
ZGhKi6i/JzkiM1msLs1vuiWGUKM+eqGFs0cpP8IYloQYpU3DVUoMH5nK7oMqB5r8G+IWJPNVASug
ajoOdARTVPZwx3enNBR+1VSkV/KOkgPiANwadnTSuraq9XHeppHfR+Fi8uGjotghm97XWmYGkixw
mwgrvflCDKpCcmJfOA3/55JvHQP6Y6n5vh7Vp4Ch8kKi6zSoUbaxSEYBSPgk7ekfxUUW9SIMKqWY
gU9a0DVi6iHwhH4jBWu2yQ5i4MCUociYWdrcSVTxWbQbWHNmPREhu3TKXcknSOlQgFd+J3Gc2FuD
GsxrIbO2QxeE9UvnelpdVFsnulO2bYKbK71JYCHwTCoV/defnyfhodgq7+7+VlFcbpBrpeUY/L4R
6jxExdhDhnwEPEZHWOm7uyvmbhnJKReHqGz2nGr1yDfOUO9bYHRtYibGzTd/H2M1SBBEZ/5NTvRW
h+j+mNMfDLIvJlEs2Ls2DKQmTDGOcN7gkf8XSCci8naaOJQI561LNzUq/gAgakuqpn6wOuXcc1Aa
1nsPFkW6KKDkuoQE5qlrOtstXKMXpFbmEQjRMD/0Yk814PMK7syOJX/WSoqXvqbS8E+dS4qvNHbp
OiLjD9koG01jE4A/llmtE5gRDKfyXP4wfXNV6rb/PmUTCEjQJ2WBCWIXGpqQwZsXF0/Lcc/mYQZx
d1W0ONOKlAbuVcSIoUdb/8MBSakmtPylcnSDpA4xAY4A8K856X8Saf4dc1ZNez01dz13GQYVgD9c
YJe+q1r2rTHtTtGoi/rUOwooYHgBg1bRWaceYHtbbOiB6bz4+mUU3+4C9VY4v9ihfnCDs/Yug3QW
7UA7odiZ967hO95B7D0zVENkNKq0HtP1jy0m/oCcQxpf4RZIcmeep51EoktmG4K17bef6KqGeH0V
Y9say7QKPi7s7d1HR82hzleoU8f1EvB+C0uLAJ5xqKKAHfms77pKf+X3z31/JhvShPpYS6U8NqsL
/3KIuMu4bJ3mpEkB4TMLpsIsXDrXSJRlE0AkPdy76vglLqGCzbDnQKz8PloSN1hiGg5nvP6eFZ0S
npowYdSkQd2dKfStEmq+QDMmGj+9Zg3U7VeSM9WsvWtFHJQ/TrWjxX5xXGEIlknUfm7XYe/JG+Cd
AHyS8NpWitm5NZFx4yGCTiHifO9OeiKBr9gzP6cJqBrF3aD/4zmpG9adAfG50ZneQNbMhVNf7vzI
G/haCuVUB/WygY03tHjChaZZPTGNFywPVbYOXM5lhrIMnbP6nHnyVROhYCGEQmpGNghYI6mv/nnV
fwkVp83NUJAcXuoSzuN7oeMI576NjapM26rq3U2E2qhhAe/rgT4AVFOKSNLHvxx6naLoHMKVrYNF
LB8mw1J5CC+RJHwrtj7X/BKeIkOQXEY9cBSA+hStomuoaQq1AAvpV2N9kS04sJoBj3nscnDdG9rf
uQcaU+EI6yGl7PWeOIvFGvb8yBgaGNETCWhbLLdfdnNV6jweodS2Un/1deCmngg9cUzXrAhcZ2ai
uwvbugn+ZEyXpIZoqXg9bPmI/O2XjJgsvxmzltM+CgWxn2f50ojOE2s5DqXf2s7qwreXgRpzwCzO
A9vWBp2Kvzx98MruV0qf8maIlS/z18mAuXen/dlMUmzupWDHwbRMqOM2q1m+UxG3q0wXiKQDjyf+
CNdwsItCTrPCzuoPcpQEvJyTD/GzpsbYQ0ss3xV0+Wlf+pZCE0O+2aU/bEwWIeHu5/7euMxSUyMq
biqeBdze7AlmhppmlYa63YY6vYJWzER3i68oce2oqA+rNDlAiTnN6A6cMSGQICqxw/0TvwEGVPhc
rlFqtY0jB03Q+XuUhnF1ZIRPII5nnwVJ81KsaISt625bHYkUa5CTgpJwEW/UE7NQdGCUh4qzdWNr
YFuWMaKQUeb/aGG3wBWzYC4+eNhmqUAZ81EPqt/Gu++vth2nvZw5NC1M4nhlxYK0WfvPgYhsjvS8
DY2CjR/aR3z3x9umPs6ZZ9tBK/BlgvyEKHJP2rk+/dkxKbe3bd7c6o6CbEy8/rt4oEAoSJRWTa3q
KRgGP8643wL1pCGoHEJlTEusMWGItgFSfLdXwF3bGjBRlIuZ64D4lTvQCxk30BUinypxJRRFOtzK
DhbReL6yXhrIutArUPLFeVGY5nXFBH16OQx60QAvBkrPs8l9GgF9svi+pjKq8qH+A8Cpq+T7BYKZ
pozWCZ3X4rtCJVBTvBTb8cwxhk36OpKitBzco2CSyFW5P1aQ2c3zxu5FznL3b7Pup+v2qgNky50R
Ra4Zj44AUtXx4UWKc4qhh59eWw0Qha6Lx/mtZ3W1mwwG/d+Dko2z8GsyU1MGujbmHKd+Nk1ge4R/
frwhH8T4SVGQxeWqY7VmB+Es4UyuY+nf2XrT5TtblU09rSVKsxcfsJXgjis1oYQoVA2xnsV0stRd
1Pj9a3NUWNqmhr0jPMDvyskHdYBih8Sj++wC+w/F860SDQGgGLnQjkV/tmvQFDt+WDh9xC4LI0sb
ozN065Ksin+Kp9WF7R/mFQNdruCtMiXey5Mch0umlS2+FG+NAMFoiVxOTPsQkWJxoJS0tv3kxAE4
YXxmk+LDGqWtbk5LEZMXztgHUf89ZeJ3DsafUwQpajlO7bQyZyHaD7Bc1W2KnErXVquvdVhsIn16
7EpjT6mJTJwKAJeL1xfi2L2VI3ig0lAJN4W6Ocsfe9QC6lUm882Ga0Y2Ff4itfNHaOsa09bhpi5C
4SISzbfZIjKdaB6NgUBPYPJaysEL6jHwiStVpdF4Yx39wc3JTFf/gC+sdXVAJ8XPYc+1wdar2OJW
hDoidJgbcqUuFt7QOZtliEX0wQHJ4zFcj/MXRgE9PxXpbOq3kVOFy1wtS2KcKy3HNpi71Cmb4PuI
hEcqkbhqsEi6ph/x+bljk2jZpBx5Bp95WkNXTNebbvS0LzlOJ2FrvV2VUaoz1LqqSvkAZ9KFDoQn
OP2oHZpyvMw38VzNHC8fWuz6bDLZyEwCbh/uCfdk/ypqHiZgobFNdP5QFq+VbZglf/c8DM7fl8WV
9anRIeuiNgtHkevrcMsi4IW4r7iZgYlEV3otKiSdP77YLx+9DPvmuAu2jfpWu15cKf07ioRD9AdV
CDAuJnI+ubbNO9g4PJpIOsi3dvvU/J22OVaMISdgCI9V8uEH9mPe9kPnFrKeP4u7AXz9kq6E1SRu
W3eiYehw8QfvOVQo6nzV8Sm9ry+wpeegphRokqBTeu6DqbLALUXd2jFCp1ExJmCxUbT3gfWneDbD
48dxNEr+JmQHlBca2l91cd679P8B5sSJBuP33P3Zwtw2xasWyNYFhAZSED7YZw8OMq5RaIS7E0QW
6hcNIgRdLdYTCPpTo4IBvjbbTMW9//BAmDjboc7/+3DRNY5Afn0ZPDL1eI/gguHjxkl09Mh1qETu
41Pu2n9tZ98NanUKura4upqXZ1AQxGBJpfF6RHaSddXEUnFlJu59t7jfGh5Z/YGV5jTNqhSWxVz9
jJKFxL0iGUpxaVfvjDihO83Qvop7D0Qj8pcfjLDsM+5gemlWG3xQ/8FT+yncA/xC+i6mFLrRmkl6
QakvqU7dTeA0ahA3Nab2evYohT/VaEk36RxeklCKLuZH5WxxtsGXhwN8+dd2A0tiTkW1clep9HgT
o952sCqBoRwPEMLcqrjmajR0RUsVb1Z5E1ggsP/7t0KjYKzaSZIvv7IIPNk7nM1aGrqoAyGo/R82
2ctTjPE7ZJg+4XdjHV7MROYW0Y45jYL9LPQHwspjXu4Mkh7ViXD10q0GZEBw7jYUoTcmnId7M0k8
w569mMHNRNtKCTJk8l8zB7YrVeAReCR0KzL1tWx2xGe/lToVnYvF1cz2q7ruLqbPN2Dm2eJ1Hn7J
sEcdniXgJiETPB1kWCIW4H5jRimn/Lfxk3haGAxSfggwXshlLcZgzm7Y8rSNHYnGj8iBScokz5yc
pzveMK4IrqWaDBE5b+kvARODHzvdjuNqC3y6PeXmJ2isiMJdSgS+/rJ5Tb8hSvAzm6M+wiWlHyrt
GNEtHKKl7YU3btm1vYZae0H6uzF7TVkr9y/MRVlyuKX+E4MP999C2we0yRLPeW7hRBHuLq1uxWmy
BWyo47GZfdAh2UHOCW3UvPbkUxeCwjSBSH2+jfD85StECjR4CY6k8G+z+8ZleXa8iVo3q7oJRlIe
uIqDdLO4NKi2dgbDBh4WJJ2SoFbHcIkF5hNoVszUF7oOPw9LJuz1m7HXvN7UoEH2NJR7wz9CLo5I
/R2JQYOwyP9NTy+Y26BbdNtwy9IVnXhZ3Sjn7Gs7thyRtHecbGZhIJdoJ0H6GCfQVTA4ciwtyeT0
La8I5VYa7maUXy5td6jYcf8m2bG+Hm/hienQ+WagQhuprp2IiZlW2sz4lIl1og58BkaGO6QeoTCk
AvR81eIFxpWKMrdwsL0FHxujL6bY9NE3aTyAnbUtA6kPjD0mh6hNelVai3Nms/TKNUBlhYz3RFX+
lGBEZIT1/VgRpLPJpJ0k+p8JWYC3b7s52SFtRv1oiTHkhc7dJyDyA8jhRfEDTjoW4HdzCiStYucf
hzEgcaC47Wo37byxHPWYwVHMog29GNR0UOIlTgNxZRDPM0O/JZDm0QPbjzV71r9gUVZYNtKio4Lg
TJBd3aPrDWsvptzhd/RSMNMiuJr41oPHNL17skV45PoYbFB3Okeyp4a4VAdiP3MZHxl35fzU6qh8
ZRsoxo7w8TfPWE8qRVLQ0RRblANvEwEWu+Wiq2S7dVJ+NzF+u8z+i2b/49t6mcz23z/0JC0npNC+
DDAAA82tJY7Qi01ylvpmNlPHtf7cGm386LwrVozf3oMyeuelDK6Ba9nvGCzSYXG8JKB9Q3xTs7ce
k0tEh7nSz+jhHo0qTAQbzvrwP1M+91oyAun4YqwwRazTvttb27HpcEAfwo2JYjzj9GWffSmsxkZC
LTgmiCPC8obviAPO+LSEbY39U96pEUwr9oDhe6KUzGhTcv+M7+RbuE1HMO/8l0Hlb/IKLWxRpEuF
x/LV7iWaXswm9njyqmO5FKlf2abBQy+KmRlCLGMhr8XyPHPZpQx7eyvmRS5SG+66dN7LkABLt9Rt
zhef8yBsrJ8Asg3/HOQvhKigNKgP2o0aeSDdJjIxLLWYSBOa3noYjP6j2AHt395+DkGeGmch2CQW
e8umkZqOrE2Ts43nL5jyQAtZGQDxV9ZbHrdPvo8SZ8O9xamKL57OD+ta863v/112BynIT/Jsb/CM
rT5eQ/jiMz2fbMjZVPi1NeY4vYy6aeVrwbgHzdbNYKctimlNtpr3PeX3fRpNGUiCosofXw0LVsuG
5hcdU4d+EZ1bjwHWz1Tf/cCjhaf6jNgztTmOaLTe6VEveNKtWI3zTXuGf1q6qX7NN5IJZwQE9PtF
Zg3ikLa5fyqqrlP9+JXOfnBTizSpE2Beq1j8jQ6ZPPe0N6onklFVGRC3tv8ZkqvQaQR4tqKEWc9P
OM7VqaurMOn3KASPruvl5FtjK4uWzQ/ro9PojtlE0Dcq+sf3VEIyqeNDoRLxVqCdgykF3ymLd/ml
mmeEGm1V/SOchFDiQcugwfdqIE/HVGcWOR4+DIVAl7EmoClkehykuf4ao9mmXPVFWbvFz7meQIM1
75hATjNGes5GtbGTM2B/xBWfTen3K67MkYU2laUOeUZcwNhXiKEa1vlxV6QqyBrfMK3t0YA+QarR
rIbNU3AHaxxof9L+oaX1NN6sVmnbYIlJTBiMxPKJzHaygJ2K/nFrYOMswo6GtPxOeS17gIyjehRM
xZkguFmzrsetwINONBrOVoZ++HsjrW6lerctM65Koydma13knTgqK233EBAb9XHjJ38YPNIVtMV1
0Pa50EpLWGCDhY6WEn4UYxf82zLwg2ETZCx+2DL3RYvY23dICGAA4qrT4TuQOsoFFw+Pz/ASl8Cr
bYZKFDTZ/z9iDIP8v+hSekq+JOWepI06vvMy64K9nNCMlvNoWqJ2moO6tdRS05I84wJaXpGAQQdz
4BsWingVT16Jkz25HCVqpdcIlTADUsxZP8nu2fCAlE2pDXST7eghpDjvzliJJoySxoUbjVO8pig0
MFdUqC806qxNB/e187uddVPapB4tQ6M8zzmFf7cdboKUR37N4oUCUj+fkF9err/QfJHmuMa3YqjS
WBZ5ql4WRFh3WB2PXUadFZNI3H/UGuEAr+HQ9zoVmClCN8N2V29/pKaOOgBV0p9JDfPqzL872LR6
YsJntuDDi/dTj725bPSHZyGaYLmksh9yRcX5utoNRlS8BDMRC1rlNFZHN8CjWUI8/hNUnrHqNaKG
geOBjyzwiUtWSWeA+SCk64/VXGf6oJWj/zPi54ZW0nvO84T1hOZWTVMfZM1yDsfKjTp702xGHJEi
h8E2UfkKNjlD0zQg+MEFijqx748vGfSAhs1UAGUrMKKHyBWSG0tnJVAi9tBnCUCII/wISY/J89xf
WRcUUsO3P7/R3FZnQwkR/498DLBR+dUt4L+yIN0E30m4v5MUV8lYuKXoHHQON3SMtQ8QUm+cmNBQ
uxegxO3XFbUlm7egsCmi9rj4T+F0t3FbrXlVgOnLbg2OM+Mj/DQ+xsue/FqTMfQbbTOsHYFIHEaJ
/HNY+SIq9/JUdPFt5hOINE17j0vypGoO1SNYXktWfA8lO21J+eGr3Ik7OZ7UxPmKTz+Lla5MkKgR
6NNcbEjarbN10vuyjGVjhPqfLd3cg6tQbsYzDjbgr2L8G0gursBHvCfEqnTU6ecRHVUTEuf12Qgw
sCD9zIL8eDgtXOPv8EjzmlCdrF7i8+dwCSLoK7jgM5kYIfJKLVYLU/EAFPxUZRWnrJ7UFv3hKbZ1
l3lPJ6av1iUWc2o01E3wu7P+K5sAmyhbm33dqVebfhXTVt271djdyaZWOJs57o/3mUMAx+31MBQ6
9dQZYTbNTcVhj8Isr35Rxtzfp0UaIZuSHzyKPK9TENutXLBUJlXWf5dvWjkFo80Unsbix15wCNd3
+zsM6MS2ADP9iw+1agwKXnDu5xqzo0hfe+uAw4+eHQzn/rFlyOCUfHVxmdHArJrIQ97HO0uim9J2
6yIAFXrqnvGf7pDL9tn/JWliy1QmlxFJeNg4qcjQOsqEQxjro9F2G0y0Qc+TQjin8EsQ6cFG5oJW
/I4gwAZj9QZdtJ8pQLUf0jDxsez6p2G93zagZDvREVGNXTVnyPTiRkN8g1T6gVVTDG9qK5tvmpck
CDE0F1kxCPReZ48JOTcl+7wk+x7AdvBDvP2F0v/PMaUNuV2do02anqcnaqIzC7NPKqFqglpqjJbP
KNa30jQp8xJLrf8TGsX8BYm0IAhjxA94KrH0iHNYWn6birOqCOmCLQKmWj8I5hjEvd7nMEhBoR2/
f0jKkYxE6ggC6/2dVQD84rc1+EmNQwvHneIBkYeQQfi8kjO2rZfKWSRFjTlaVUPF04gGg9V99y0/
N1t0jDbxqsMUPPsYJbZO8dUXvXKJ7oaFjNnv9DEMfOPmVa0soaz7xc/DQAcuvpSZN5oiQAccE7Fz
zHZ6KB/XM0y3LT8bLkTsByEjYuNIi2QbPER/5wpz/LWtAllm8hvkYlYuFEyKto00xhd30dALmcZ+
cwQuPzUdn/slsftf1M/N70AKIldz3d30yOr0Gla2+UlYb0lhClUwjdJy0xds6ZICNx1PZePL7N1Z
F3dsSln2F4xUs2CMRwFQsq2f/t9qZFUpFuvHRDT8Q8GnLU3Mp1d/tbJpMuQLiS45G7aV2cypsK0g
7dOGQTDuZKkf60ReAIEoVmy8UQmMRGYIsRW6+zmiSKTL60zMOsXrSA2jeWiivMffdgGBU4O7mHaV
zqC7NBnLZiAyu0DqJ4iyUNzQeDYnmRUhmiutN9lvy/OX9ed/mFRLL866++fddvqFg/cG2Hx5Nbr/
iTNIROuESro5vvaQHfunF9URIPNYDvr20cxsS+CYgM79tBInfAHXMOTNL1NS5xYFk+DRNm5VL31h
xJcScYBdmyYtRQB+UlHhGgBPCU3Kemoe4yjzvK5ce0uMc1lqhRmwQTOE8L1Ce6AndkYbu/V8ut9X
RBUdnem5uJqdGR2kYp4QpUhxIL/tKwY3s1QXjz1DgcTdGrRDPXomt4MjmCHrv50NG2yLRMfbNQav
vdKGSvjElCJS+WZPb9PxU99gOt5VndQWPqvkToM8i3bG/1qNxHNh4cES0/IwLXFfvc8/fEFLLbsg
TvAmBj8+esqotOYcZ8LyHnbic8K3yH6xdsb/iHULWdP9UZOSmwt9Wemaljh1i7UShOtY2O6HxpeM
y3Gw+2KEWCV0KUWpRbjwZyLvkZmLyPJi2cS0wtP/78bYImN2A2UEzNpl0bEpK3shZnvF0uUBHfJa
7ry3CRezb1qxBPX+HA2nW0G02+17uu6mBPYnEauhss4WuyeWRmjeLL/Ymk7TJSh1FEqWT3ZI13l4
Fle1cojs2yWbMfkKFZTn3tEFo9r6RaOyrKN8VFbM0VXcGmz7Z5HWW2mkmsFMVaYSGBu+NfktwZhx
Sgvcv69xYH/88UzWylzrSKyKoJ7MTk84vaCth69Qg8EETpP8gz3jzuf4bcGj21hRyrRt16fUTLs9
AWxfkEzz2gvOx6U0SCNOKWIWZqK4nZDvN1fgf6Mzhf7R2ye9TABzm8rCNWruvAbSqQxamZkyvA3u
1OrfkiaZ6PPN+eEYxSYg93203OsuqHU0vuthpqtnYbnTduXheW33WAgwas0ySiO/6Nvz77RnO1Gi
zUvCtasCift7qjNLxLtzVpsIx8oOWEeqHnjUtMznR6nyuvpdGjCNajJEeLP5smGAzBIrmzArq3V/
04X9dCDM5RYILN0M+MiIFQxWuP7CUQlT25gZotb4LfvTlJqRH3LJ4UOKukBt0a50J07NZbNK1nkA
HdrM3V2TieJbFhyjRbVocesszWXUNU/QHMWsXlPUtafAwT1MZsOh2WKcBWxoBm4jQFNvKwjiiaKd
mMTSu7B+5pL3wCL62ZDsHiY4rtxv9xXdeKHmef04WN2sNERqVVCG+u2TcMibA/qV69ECIF5hWZ4u
LkYFYe1cf0iGjjA2w4OztNERYZOepQXEgevEYq4+LS75EPDkhj+fgxdEWPwqzNJESReWJQZJYajP
10J+xJQSmcyYelP6878DddYjCuhWwLZwYx93uRBTyxg5IKer2PmPR+s5kY+h2eZi7+t76cBoHcFu
X3o1q0mRBRBGacLw20mDJq5Q8kjnhYECpuDPqD6dSWQdjg42P4iOfP2fqLQiEKvvO39eAM8PuTa8
rzUIQ+KI2LNH42Gb4cLO6ERraL6N+R265JuPAHirukLH/015yMA679EDM15aY0cTZ3TVY88R684T
mdbi8oZt/WQ+hbB/uzCsFb9Q94LTcBsfc3D23IaSGbD9z0ruAVPS87WylVs/UrkzZBxockqv4jiD
M4HVJi9ph+sgPbCs105Wk80rKdCugA/qoBepSY2loUSjbLCDe0ojmuTW3b8wTJ0utK1uDxySBuE5
KzRGGRqj+BotU8QDSP7IlxZ/ci87eTE3/YJQ3wCxRqQlruZII37D/c6i+7qyZqCeJqKK+GDXFDn3
+7CNHlD18htfEDIW7HLUXFPXxqngKlehv4y9qqOlF9r/4r+A0jnQIIiNGdWJyo948rneyMxB+MsQ
rym+zhwNxIOichk9GbcxVjV473o8TSpeozmlpSVKK4PJj3/pUjJM4s7uKXKVM9U9wYNqG/A0JmNS
MEQ8g9UVrKoqPE6KGQXdeJ9gLde4vK0X9RkL3TKKaj2+JL+0q7nYKhbk8NoKAHPHxutfZpTeqI1P
GlU0GDO/aHJAVvrYw5YJcTiZtHOOLnfUl0f5enyDXW1Nx5/qjmi2VaOqekzjKV1IATo/rb5zmSXE
1fu9NGopAeasy1WAmViQC0lDIqvEvTa85DQDSDl53bT4Pa/xdSSoeAWoS4qWpWBD16Z8ig6v80K2
PgZhL+PsK+UlC2hvGKyu3yJ+6KOAQARG3qz3vXMLX1Cl+TDJZSZtA+28rO0M95sWYBJes1Nd865i
sCiUap5Cdo/S9xElf2lD1SIVibwq7d82ZBl7YYXq3iVGYyDMYsr0TbnQuu6Pj54H8kBpx8so3J3M
gyoAhiaohnIPXeib5crIL1QkBfbFbt1ygIaB48wb0XOLPL36TT/i1EPD2Y+oIZd2VAvK08Tz7Q6r
7B5D82RFe4S7bIWgsM5HSnyZrEAirMlXdHDv7Y+PMVpbUUexmCKW+KHghwcb+OIf8KX4Zyr2Uw+i
JFzhV2eTuYGQ1MEuP8WlrhIio1AC6UytV6ft2PVLN9mABMXrf5GgNZRVSplVF75cmciPIzWyvwp3
/scbmzso9//6VErRj908ttBtOyShL/1JkeVzBOxzF2MxTCWQOSVaH8/zEbihKektmlJUht4fxY+6
MVZaTgRIE86Qh6CpGW5ONqI0ORIUgyTL6d2B6rehHU3kElSt/vBoOZcRPA49qfCeZg+ZEF41oc82
uGiUnVWziGPAq+bXkDLIO8RUP3FF+zZc/5iTg/wEwV1x4A6FZIfEhnphFyoLh6irQC1pZHi66i/l
pvh/k/FrHZUe1RuhS3sYieqC+jFxWWSVVpZyNfwxHxMSyOOjVLGyEkVFuJXeH4fBVgyL4ezeq7jk
3PV/3Kdx4QMVq/sR1Td+4ztPV4acTTwBIC8MUXqpb9x1ymDuxPAp08vhrceZ9pbBGVDKbzPKHDQl
BUZIMn+BEZm75gM/8YXglvTcC9vkEV/Sh4wSN8lE1HOk/U/6YNSPnBYGViVArYoRnSwEoHUb2rVU
qWj4M1rAN03Fq1qbxGiesio5gcnvQ/aZqezG8MHVSSyG2ApMUVoDruDbXT0jg0aH7e6N4baKSleM
6oK6kt5pKxq0IJIeSJzBjN52cP+Ban0wFqBu7PJDgVmsQCy+AqOzclbkxW/D3dAuiD6NKUqWac/N
2NkUz4tpY3jTZ0LkMg2Fia19EhrYDLHz9yKpBG+vS2v0acVpWJhY7tw46gQC8mqcZO06AW7H8KXp
BVGv6wlOIh4YWgRrNvfBxxjbfldhMll+0h3sX6jASPHGoHe55z0sOeU63/GRxtbKkoLjN98IKlZ2
I9vP6xa9BjVyp1gDbqpe7GBr0Pb6Gq+GBNWzpQVds8mLs7uQvESq/jSy56H0kY7yai23bqkb8KtB
fWIBsoV+cgVGsK9U1nku6/UDmh4qd7b7IZedZODDWxWMmIRXqEoqO96RL2iQBInbh5aDo2IgB50v
cG10Gkd7kjXCtBALWOqxBgO54Q8XH9ueKkzFEAkN8jKxY/vOsgkYc3+OrzIXOVP9ADb8HyGGMfvf
FylHGNW1WWuWWKBe96dgc6K50tX5y/s1aJKvTilDNIGvI8Sy4T4q7EJowLD393T2vWLmgaPAtZ1y
6iFNtEkWH65+j6gc4NS1OB+rqdZwThK8ij771hinG+plKO/gZBYRBKbqbcMCeTwAbYimBH2gpo8r
FyG1cvD5EcghlUqLGRCxZQ90cufegYsrygOWmvLCPMZD982KJ5eg+TMzt0fgp4H0SOQbDB7UpU21
kzcSI2t15idnHnJK6JNkRPx45O6qac7GibBPgW73oS9Wdk+Ih9Ch40ZKEIgLOpfceL9gVd0EzafG
gvxmyfV9KQhzZCcvCIR2b6UOMZnmh75Rbba1kmDRZcU/qoOhfYVsu4k+wy2oQuJMRsb/iqrVEyXF
TBQucyxKbcBQaCA2d/3txeTNq6y5NdqSvtjcqte4bua81H857r+5AHwTtanK0/Kds20udPNldmHN
LvIpSiZ0bmRA0wMXjL8DtNE0d3KytyhTSJL+TlUpAnMWukIFW8h/2wGgs9zNWHuaB0qE/5d3tvKc
7QaMZAMF3w87H4mKrf94HELoQZcIz9J6Yh+KHrSIlUtR5rbOAML+fYiCvJb6MXCabnOGkW2eiLHk
13Uc11i1X6qLpLme72vrtLXfOHDn140xgsoPzC4VLJat9eixWTiyr5SHu/xm2w1Y8Qiw0mvE4aJz
LdTxUSZ/+FXJ9w6zmVDoIXzpnIQOAOUJQLR+mHxR6TAETA4PVurH5QEYpkRVm3SS2QMs3/FOnzyB
HAl7wb/dxF2lQvtfqzoOiwEbg7U9XUSiSWz4Jd6jX0uoV3tnYUznZ8tlsGBeFDttlaZ6WOX8zRf6
OfnOW1vOqs8nvrh/1vjh6qN6nYIuQhj5JC49yMiD8q6xFdxNc89zL+SJnkVj9h9QmY+YgXb7O0TM
7EtNLMS5f9K9Ujcwf0PPW+iWqFU7798cvIxFqzKRbuM3foObWa+/VNGIPhkKqWpmbrWCBhXBhgq9
tHruVdoBX64TR9Uu55lgw/lJCC0BHHvgLfnCcv9o9h5OaBaLjAUjT48HVqlzzOoRiM+Hxx4waDaW
m0G+WH1T1oShJE3DBwJGJcotXdDxXCoU7G3tyqAZs158fuPAcSntRDTegpVUMu178/gi0mjO9vLL
c7MVDejnCAOPmvxSz9k9ZTIcI3sO7cqLzzOyjJbOmQ25boCpkLFpgTixhQF+9zCWL18iwcUZ1vJo
spiZtj3IzlxBkglKJZ1/ZnMUqkU8SGbZxoXk87rZMAVr+FAQXk/KQaVxNOViT4aLMLOjLVJPYScB
6jqTjeou+AmNzFFxTqp4cyS02Y1mJV5dFN+3mN+2S7Qb5yas25/GMKSObeKrrGQs9URFTe3X8kYX
8Nt1UPkjFIOQ1UsP2elggjINpKN3ZCR16cho1EGS5t2vMtc/y/FmLIgE9AmZcZ9hvcAt/W5Xsp4s
eAYjLMqb1Ddx4kNTUNNaXLDs/RpZTVqwD3LpVNZooj8xX3mFIeXvwBEd1IqArYRLqFPjb8wyFcZ4
TlsMnE5mozOZOwuh1zPOuKl2pGnseES0SapTQy6nz76We9S9+IUxj54F7yy8wDozeXcfY33WtJGT
+Tzt7ggxdDjqEstL6uWaqMOd/YwxcK5Q+D1PyOsPaTFy8If30EhyiKCEdRVvuKgdO6SVBR7QDM/a
RWU0CVtjn06anw6yPbvmNpzyc706WTSwDAf2NGYlY5LD0R0nuaJ79jB6WvhLKHdpF+TFxG1RMkEp
nVwTQ5ZwqeI1ce2Th3DGgM3DC3XH/k5C6a5CSOS6bFVK0vMaFic0ZAwuoY1Nxu6zv2wxtfHGHW/h
0mZLy43+Ut3f11zF+NvHyq6Xks+JZ7hDDUqwi+Uf0TKNtDEdqy+wYP9gSfoyZDhBR7Ntzjf2RA/7
Gst+Kr9O8RasCTIFySgh0R89tECNPEDoFA2XzTRmzepWtKKnoT6ASDOT1katP7ioSlQ0NYGj8EU2
4H6RNqWHsNo94rwTRQCvd5MgStw64+hLcXlZ+pExxynmWy+59hb4M1UInbMdDeY2cGcBI8Hc42Fa
8GnRKOuhncThLf2dsri+fIHaI+4pThK1etnBXp//A4+6+JFjD6tdNrvbjMeBqF0sInt54RupL0GC
WU4gSSDeMcDPg4qSQ+BgVwNVnl/iR3jwzl2a6iVjg9++S4pCTpL+rhIJuQszzQV1JyQv9kwF0VI0
yf3q7pRn9fxOpp6VNMJ/BAE8rmzfdoah4P1j636NVZicMuH72YvYYSepi6qWJErNQxcY1KZR924Z
miWgbwYUBKlzw95KNJ+A5DFz51xbf+X5cBI1E7DIIs/NqGsbqoNTDNMh3CnTf6F6Hja+0aXWVx/d
cmlCkUdcYtdiJAxkMSmT3YIMyqN56qcpLW0eH2bE3CAhDwwIzoeUD9eUU6DpbJQ+nOeZ5VXx3s00
ykK2xWpWzRqpLy1uZQTQcGHFRQJX0ZiDh62jf17F4OOOeXVRJcGQaBATWBl1yMbaatpfzZhr/1si
Fkj9Q20wMdDIvsY2t/AZmXodkw0dRPSBgAe/yu9OJ7dYEGTvf4V+SlIKrgsm+og6P32KLDwUrT+f
0QVBqNkr/mhV4tTzSGQrTEB+rZdMtUOW7dkN2cHC3LdUwFqHyd+e9aNFFOQg7iHazdqyzvVheCp2
8vJuPjSqviiRtY7a6JfBIk+Fe0zV5lCCGimhDenwXu1u4675Lx3RKbJjljAaapCV4Dx6cSh6amD/
i3KmVycmeOdvhZRMOAFUwdrClL30z22EqR7zQEa/opHmt6XFDeKkAx1tHTGqyYZarVFu73WdgyNN
7LOpawoS1iElCQ6j8ntvhx1AEmwfjrzusekImPy94z/HnRCQYc3I37NMDqTDBCtaZCJJGmgPZZEh
zxkc0yext9bL774TkQFhRGWCzfyNnzrjb9MkxCvcxfROPg7qZsoaa+OtXbhmhKQ9xQGmAHBltee/
ieDexSY/Y0jQNcoAoZdidi+OCWWebKg+BTaMw9pVIsAGDOSR/O7uCFImgIBzmaWjUYkdh6njBjrQ
WxyT2/uv3AhxZ6m2jZfKXev7LRfKG5fOt427Aa9fTAEjKS3d+b6fuHW19uCGRvVtnJBuO4mFKAQd
+TelXGgdcxGIjO7yjUbfxfqmftyhUW87tCgVX+9W6ysXN57bz+gTyeYBBiTNhUPXudc2d2RdzOWL
5NqkfhJ7/3Rc9GWhyNWYJS0SU1EUiHIXgznvMEAyxrl35pzcQ1xAFY1YZeGH2jIexUjbURrLWMXa
9ogjmk1TMe+9LYnd313XmnrEnWU5P1eMlgkrREIbGhXmq9Jzbkg3E1AM0qplBMv560f29X1Hu6Vb
ftlrIfo0k7qZUrL35AaJcByxl/JuIz8Wzo74oDS3A7T54FpDBNXXFE6FvQ/c/W6QpF2KDLmtGV63
cZ7qOPBEK3O7YNaLTa/MQ/1j2VM6wXzYWCmUvPZ16LFqAB+0WMJTTTz60b6uLR8sEpZd2oZs52Q2
MQjCTMe1eod54/FsV1w7awZ6YKEJc4Fqk+OopvE3KBNWfHz3WkcuZAUPxJFHba9HNlQun37097Z8
Kyn3JrWtgeUOqVNy6A14xPFwD/i/5EVqvch+LmO35oTpCUM0bVeVgefZWjme5ZXzvEN7z2t+YY+p
xqcDb1oXqQUKRa5BmCMFqFlxc0AzGOmLnVniO/cDE0ROz8BSOLR4WutN915zdF3ED2t2eEqbusO8
e83Mpmyzn32t0Ku/CRO3MyoGH9KH4pjzdD0DRwzJFsOwcep315peNCF5+l/b+iIgDLlf+ccHdBVq
L7CvCVqoq9+VIFxYcN/N6PEoBRYfAH8PorWBf/NQj0sXwiY50414Pr6SBnIGRj2JSElJ4N8G7Grl
LgMVVxAIskEsVtbnd8DaE8rQisnXrIzfC8/wkBasnWOahFrD3Rp0YIUgvaqutNdzorqCQSbPJ2j5
8X/kQ57ZDUfQgYaIRF66HMZl5HbkGsboS02gX7P4++VknnwGwDEyhQzzAyjXDJRODDb8Kl828KOj
DlbWMhXCI7m0wWrg74RpTGTlGp1Dzz1W6aZc3s5bf2YB5CASuZ4LdmUyOXjKyf8hlFRLn0Dn6CNw
GJHQ5sifR3l+v9mTVaOgSXnxVqNhCPLJIjmTsLP2KeAhQt+/Tlx0R4DomjWUDf758WpUPHbuOSeL
/uiVeNgoK1NyZb0wEPyQTyukxrn6Y8xpyYQYB20s7QRvdIUPZGX5ZnlIW10Oehr9hOHesTG8oBxA
c/GJNOEg6YWc8hofeosTnqVvLt/f4ozsePDL0AqFAn4lZLZpoOOlXX3J1DAUnOnG7yqBRrKTkYbO
BmzgnW5yuHO82RU80aN0wq8uybR95mLf0D7xBnp+YY1nmxPkyL/RVOtFUZLJANXLOExA0b0gn7G2
su8XQrEo0UuDuMfFq+nu5xi4oz+2jUVpc8cd9oxRrTrOItFZflaXW3/HU1lBJaYsMEQhpxdMi+yg
3BSaBOlB8N7bFbAnWR3jQB1RcEeuEWq44VqOaG7waeZmuNHx293yREAqPuDi3VW4YPC2UUBKC/7n
8bFjXetgz1JG59efUeKDorCsf0PhwMNcH2z0/KZEG79uR1HluyRMzFH90xp5qerG/Cj5OP6XgWas
qM3IRfvgOegyUrLODIe49vOaTVmeT3RMXW+hTnXzs+ji+ziw8LLp22IVOlbAicya0+aiw1YGG/9X
gtF3cBB8Ka1KrYPHKmimhujJ/7o0OTK3HQUkirMhSysqcTuODsSa4WQBza01SLxYK4fJJbm+cwml
j1JfYjt+Z794SB+X37/f9+5cYnIMDxGhPRcToXG77NPJQpwB8ANgCM0iddTFJdOeQARd2I5sQ1nT
xokKqGjArHf1SwN0/hdTVz0GXov491T4odqDRQpzAf/I0llSreC3m4q97D37nr37PZB0QmWSGlOc
4j72fccMspgUXHUSZNz+i8I5NV3jFDqAsInzqKyEqrgM2qggDzJAbi6c5x6tGOwVh68vI1nXSfkQ
JO8sXBbZ916ySqu+61X8GYwTVcBIqyv9CObHl1/CudKhxHLxO89NPmqxFTvqER4iKdBebbJOC3Jp
FnLxJ89+pa0KNgxOAkf5bKJvNeOC14xlECuIxr1cV9Q+0/gtfvsCpR+VyULBDT1XHetzOBVZ/ufx
uVtVIbzpa5H3JpXxSkkG9hiiD4UgyUJKXkmLvItYBucyhQqy53G8gVhhOmpbXjUao5eNo/MTKrlJ
f4+AEtZl2K+I7CaeuOhiARRgxx/2ry7bRpJ8PmzvnMkj5XwF8ZPHyMXSDdtKaOp1KQEXTll6y6Ff
i6MnoAFhdEVM9TuQ8TL5yiNABNVFPQ8p3ZJ9dloWu7fcVxNMMfPpUHZh6sqSGvAp0YLLjn4hL/dJ
x0tBx94FOi6Ww8umjQrNb3kMa/FMsG19ADRsdxh/LmLmXsB7sQi7OP6+669/13DpVPWnQJ+BkPsq
l9Y7zvA8CapLuVkKprs685UJipfz/Jgjl7FiZnjDJx/Dhq9kNpbhXJHQvsshCA4mz83GCVAIjxYX
jEKmiMp6rWk9LcHCVayfdRvRfBjyRJiM1wIJYyksHAvGndvCFKiV1NLMSlZT/K3t1Qb0/Q35kqZn
1eIl2p4fac9KmLJPVc6atoHm+nMbjpv/MwdCJzVZGs/xrfYOANMGHMVANvto6YjMk1YJGYupNKUJ
jUS/gFw+gaspop5zwH8XlITD+Xe42JVqyLlhwaloY9YGMkVacAArDnY/lsv086eboa+rSTJnCfiJ
W2i9zX51ih35u7grWBAJDlgU1ZCIC84yy7qhV4hbIiAmRfhF8s2bLKaKPI6PMYNLI0ko+U/I2LoF
S1LcpS5lsM9fo1gwzbZLklGmbjJKoBOLt4TZAeW3kYbaL8gZFaYHfIsOGTmagUfXQPSWauPd7x5P
Tz0mgjH94RDs3wDXKOul2xp277VYT8l8Zjiw1ZGUW/JqfCbAbtjXLKdOspGykXSviDz1vYwJszYA
sHTTmLSWbmoM25brAYThzXi9ifscM6yNknoAzvKvFg27vMChWGJTjSHa3EJEJAeLoK0wPLLOQKoc
YAxrtzKhzUGtwhAi5v8Z2VIqw6L6jLzIIgfp+u4io9Q2ndvVISHlT9bChoHDwzXyCX9APQ7Lk8f7
nm/DCmG1h+eCwUcQ94vTQKdI2/DW2Qg37t/XP+FSAm0JSqqYRFHa1BdRfHfLcel3iohLpnScPz0W
9gPPhc+mZsWQ/A440/FTarU6UmtnWzP1mMOcLRXJLJxe8MggjN9yAtBuxMq5NDLakdctxxGxhFKW
RF5nKm3PuHLt1YkwxMQQ/8G4zor2QHpIHlERo21zVvgXD+khkQ4MliPKMoF7pN958OzjpOM/2OFZ
KlKSesq6Y0oNOqUdP+/exzTzDU0FTnO4t/8wIaALNKJcQ+5VKW7PHjiLc4dfou3BeJJp35OU8ZXA
YCeiGTvF/lkR1n6b5OUwmMEmIjjS/+TiQ+UaeJbAS5uotL4TM8tmePDGrGtHzHbPjf9cIiO385vV
8RBMQREibRlbRbavM/VYUdxv2NJrjMsWfhRKUzYq2YdeU6u5Z8EH2It6pqpKIxvkHqV8oWNGbYNJ
D9ThRsNs0XMzdGapiJopK4bcBkpq0hyw+594bQ4Gt+0WkWIGuHzqerl/rONqsjTakFrtogiGiB3Q
1gUfde5whFNGZWoZYJoXtls284WBpCwPOotF65h32mjSFuPa3DuWx+aoVWlEwaUqzJYakP0CLuQw
/hcKr+g8GUsYsdTFQj/526eqdds+DacK4HtKPc9EI8zJ26yJFpCDsnqPsZut5/yuWDNKafW/qPcZ
2lVjtkFL/1WBA74bf3bBRQk2zWB1qgWrGVU2DILNuZFeuf2+j2XZZ1fAZCDGlo2k5iQ4OZB6H4ux
j2dhK5NsKG87/eb6WD6QkaJR8yHIPyECj+5htijNlApwj+KaoDb/fg+Tp0lIZZlkcCbwERYJTYe4
2eOLbFdY4H1EACHTRp+Zj+V6JvrxAkb5va62XzSzI7D4OSACZ/olVbwGXfA9L78nP/GYLpFX327i
7UhZ0NO7WOxTqqhFg6KQqFDBmZzJwRZFIGP5GAwJqnVtRl1Qn/vqVXcJrkcsPNzHOUBNox/mWeL1
PA7EVChvol6jtoyE4g03E9cdb71CfnzKqx5jVIiJFidDJQnk4wmECqGWJjVustgRbPsf5mR3dfaI
EF7jTiRtIVag46iEpm7f4ptuxj8+ubs/x2jy/uUKig+sxijbcbG4d5/dcA+N3g1XyWgdHRlhqtTp
ELTDXEEwBj/GsYa2JcZb78O2Oo9uTsr6QfRJ1aKbBkVdiKW6v9QUtK9YBX5hJBOCLC+XsjONoNgP
YaW/iOuYzf0mdtdUJWOS7oIjd0s2UilqBuLo+nSbAq+S0KypCMztDcWqY25z9+5aNPGcYO9lracv
8KNGp6SO8UF4VuQ0VMBYOx/ruTm/QwbQLyFKNiaQFLK5Q5w90zmlJ+UkkfYQH9oSITTbhpKwgjq0
ANMQgWQUdoTAW6ouwDSS/SrURTpiH+uTG/Q8wVnl5Wa98BAIe/cQYJOdpV/IXZOPenJBUqJ9SAgw
P3i4VhIjmSp3TwZUSptNraG7C7W9QvWPDA560r6xHQ/JM4wNY4J+5qI2bPlqpe8EiEt2SQ3b+/vx
1/858kzvJj7h/hc3slVhOxX7dhUPTTN2F07M48O65V7ZyWDiozq8tM28rgjPh14eX+pHfvWwPlhd
YX5W+I7ecStdyziRkCajbsdcAR4SyQbiP1DP0gLeauNfWTiga8tdZydQ9yK9WZjEnPuEpArE4sm6
WIGkIZbde6p1SCaUhwh26s+hD4le4urSQrz3tVTUKVDYsyaYh2tffM5EiRl1wOke2KaTD3SEbdZx
UvtXmTj1riTKW+KF6FjRETsWYsCdL/oKXdrCP+et8BVqsEuA0b1LVpwMl9lL3aGmaZ5MSDeHEl0r
sJqwATKgsYsZyUIj38smg7lCSE73pDQ249BKzJreX3lr6RHKOKH4EFaMCojt5NfIkYzIpe8cDe4r
j/6HVVYLKKJMvDxjtLSnrLXHE0Lc8dU5cByHzkwXGJG11WDTiYRh3rw5dD76PU1A4j9Os5idEh+O
RAuCazWsMWUmzuODVTyvuhCt/k5jRY8ZbGLzEYsG8mshOaHtmXgd+2/xPLGj+tFdHKZiWYCIaqZ1
B45lzOSdXEs6Jy+uNWZ5RzWFJcKEuFISa+GjQ/Otw849YuTdDFIJR09FbRzZqXS7N64fmUJslP9w
NzG2J7HjHGzwPf4Muy+NpZmPzT5TF5YZkCcrL1PEHtuTgSY3fsidbO3cDasWe2k7C566aYkTySfe
S69LSJ23UnkiCehcNYpR7rghCsMbZMzVeXKCXItBSMIjWFSDBQAt4CBPN8ZO48KtMmAosPxlxvZ7
t/kC7zGvQeM1/Cf5lT9lzUdz5RMyxG2dkCIyfcTtQJkKBKjI7qjVw4rNxsGhQUaTHNE0vtFTNOLs
UDdYxz+rnC1/sEXtche8j5/3+JJh53gm8qIXJa8omDo+gGTg/9BBmBKI0x/xFzNnNOtESlsj8EWp
H8xUT3o+43yKXz0cmZXBKx3Impn3CIuc3p4SJAQCap/fkGvwPZTkLEX+Y88en6souh6OVHTAHsuR
DsPXEQFOLg9iIakQABtafv/UaOeru609fMiIajyGu5aMrwxKVbTuKyNP/JIf6M3XwsduwmY5c/ZZ
K2PBfs2pX/3vaJtIG8jaUXWsjCJZx1FZJ7ugRvMOPHTsHTkgcY6PxfuYbzUrrm+tFnlHdpML6wzT
xl2hdPT8hGg5FpF/hBKhMAvZVOig1A4OB/m2ynDpknFVkdpchxaPbNoRRfLQpFsOX0UuUQZwZQRs
7RBgY24iD27UjxDpP6b2cSx0m/XkEUUp0thl5rwCJh4mnxqp1BZ7mYBsFtACiuDr7DZZ6SnGM7Ft
T5t5MyH84jjJZFAW4Rfd+UqlBVjBHEFsC7aC9MPc41//npR7zLG4qCUHhbAK0BjbkNGJaT6U/NUi
duLoVFnXozA0vK/4rKiyfA3hroF/3IZomCazKI8bOo/Hx8wuxjfFoP7ch+lF4BWqk9qLnQTT7iwn
+Dj1kVJk9A3TRqXQCH6VQ6eWgou759oOhgRb0XFijmECLQyUbwjVPzmwUbEvUMzoquxZ/3WpL/hd
QMD4O4fxJ4b57mtUXHYyI39xD0U0lH1KyWBAJMO7F5WtpUlwxwfAjARICr7xi8uhkY5Oo+mhVX3n
UVhb7XZN95+XtazFaEI5uuVdlTua0bQnEvIE+PO96v9NaWeDEy9U5CaQRUMiFgr372jr9c/n8ajD
mc4hRSmBzTgsZv5CyW6QvZesfL/hC7/m1YEvbGJ99VNanOa5Khb74aPOY+L66MU79EPLGr4A0gEJ
ygwCGdK0isHtAfdizhiA0msG+b1XzTaoBaHJ0odpoxGqq5pIoapQnoWd+gzNXEzP/GTjZD731WrY
PokqVE+vgUPHANx5Oc7+MmfbzQGksHNr9awNO2GYG1oaadg9L3bv8NU+O6Cc8KQNVVPTNYwFxZsN
Fc+Nf2GJCc6eLaeZu9sys+JMB66dxCP4DVMUoPbdqo36yt/cq6x+6zMuMClp5tk89pjp+6wfyjTs
FtZzBYFAtHAxPFmSAftZAPPb7NPMKn44oztTmIpLJ8XWD3mCtaYlsQtyI0g0B5DUmPDGts0FHGlp
CVRqsXRPDiYB6LuBSv5Z1gBfa+IWq74eOnjJh3vD5Loov4elqFM1iVTKnuzkVlCZkKlxCO//wIRh
xouj3fEEst3e6AfKAMcql6bcFLo0lmIU9Af7lg6nlBD6EbjeM7dvkyc4Clt7m0mWHiH0Scfy+Vw/
0iUzkFx9ilDHtIQZrLRUJw1ZvAtMrsg1wNCG13ntNwO4+c1kvE32o7UrX+AKTHRR1ju3WSU7zwm4
xfFeJNKEnVyekrpZB7MzRsxyg1Rnkx+a0tGxynqSisGSpvJkSc4uOVOBfFKkZqmNkpvIVr5IGFLU
Xm0iFJ6IBiI866UiVXUSlhZ1VIh+FG/UiFpSyGiPcSZLgR34xkXbc9n6QuXYOcOFkidJy2YVZEK9
OlsLwvqEGLaHYttbi0iQVFI1C0T7IaIrRkSrPWG0Tk8owR3TQt/nW05VK9fnUa9SCjU94wWdIUnq
PNWTrAvlgerjdWeexdBQarYgkWdzV443BcfiPHcc0p5888ioFvOKKuyuPQ1CU+FzB6I9G44p/Jwa
Thi7jyaYrJ884NWcqTNmFk7sdeWTLjYWP0jXrpfBGT1OlYPUcocJT/amthylALCbWVuIlSfS0YT/
YPn3BeVr7B3qhaWHJFx5Yu708ZMIb2ceHMbLntvVrCVBg8gZ80UJJPa8tBCEnlo7qrDpou+PiWD9
gxjQ8/6hq+KFdEFHbkcTK+kfMvNLBq5GjEXWxtH31xF3LiQlrm1agWa3BkIx5HQqK5z6+VhPCcNk
x5ntbBrLydI3mIEh2JgEoajiaGE/ZJXtFP3NHXAC2ZmFz8TwcXxFD5XvgpREFF8JW0TF7ByDOsTR
orS0vPnAaLckTmM+aVWpdw8rasDAw/yESaOLLOOtdAHbABFdtmWxzBujah2/fMq/lYsJjfqsSCI7
MMb/ocFeJRPtuPbmu4716MB66hMpnD51wf7arH1r2nEZkE0wRZ90Wk+PDfFvpnwj3NVhuwedVBKT
IVqXF6eKCKVIuQcm7oX98RSyOrMJE6QZ89aXpybP95d69+NJyshGQa6a8Ojr4zWI70Xw1s6kZLkq
JNMUyTJj5tfFm7n+8/4hHdl0608k7opcT0jZqUqEpkHkspWilkLTaIulBFf3n6SjGpa54jtwCP6a
PrcRpiNLIyaa7o73HkQzCblWDYJSpscwIHTlNoGj7hOJcQugE4bKQjeJtABF7InwKf4QW/6n/mF/
KLD9uVQVNIERXvF9G8fvALNsdIbGNdDCma+uEeRjwEtwZ3T/ai3GjgjAvFoKdzlNXn4CvvxcKO2z
LFo7NAm+1CuMO4qDVPIIV+pSB73M4RY7cr0gWKbcE0e287uMghQTmdRBqoSHYvyEIgn6yD/xbEDw
xVLqkfbwftm62wa0trF3MUmVb41asy3d8SpPd+DACSMXeZprRIsT5Kdg/FQV/dhzry18+sGTqHGa
2IKBFqeANTqxaiHZaAtI3y9ZYb1Bikga8vHLnLFbRHlE6lONMGmZC8hlu05B9UINJITk7ms8Jhcd
ulXN8nQkMG6jBnnk28yOGzUiQH1UAOkg6YSSSjvGcIOwJ0KokeIcIinQ0oONHJr53rnltZc/RiXa
+WO+UGYw5j3y3LxQjShD1mTVtQxwHIPmogDMZ164jmyWcX/HxXie4KNP+8EhvZ4z0MxGp1jZYZMB
hfv2RmyN0YrMmEsZjut+Ccy6vWfYaeS4OpO86Rb6RXD+yRCYWstqL/C411+xrLvB2sgSMClS1d9H
byg1Mn/z1sP6KZ19CjSWoILnw+DCewHfb6LjwYZWYAwBLO1efDHFxaN/KkSh1Pj4SjAkfwjIHQl8
FeKiXroUC8/gCDt7ANE95SY0lHA3LPWR0VwZaYeXrSKzvnfI5LuVHVBbgz1BbvnsV0sQEHVbvgjr
cU1kfmyIschzk4IQXZR5uXbo5RYLF6tAcfnqPAR2cqPh4UEdtzzzGv1TN0a5rimN9hBckFqbdzzV
Otyo2iojNUOH1W6WkgetyDpbjAHJxPUJe9sddOx2MuYPAl1UPYuoo4CFikbP0/k4nojfcrsHqjtt
pmLRGqfggC/dg/RojR617QPD0qRing+zfLlxlLG4pWZkycoRtn9oapbtQ79vShWSvxIxFVNSVisr
jpzkijIDcAe7FuOp7cLqfj9QLBo75cCsNuSAFaAEXNF+TwSXfd+g9GQggsAmioEZltc6EGKMDzsh
6Jf7he1+0ZngcPKIKl1TBpvY+AFbkPFQwSQkBWznfN0ZNMTj7VAPutLmGVGZzBHCc2EdozHH4ieT
1mQK1BYIvWQDprpfLJSHnDVZ/GAPSiTh1TsqXJiuj6CN9OX9UzIqFMxql/zH0KV0KPJxX1oIPIsx
R12o81pwzgIzeQ/SOVnGSsorH8tZu5gHC00op9RXExEFPbwFsmwK7KJA/e/ULTxWtEkvBeeY/wDi
FS45i44JCkQnNjBVH540k2Yzh6FoOKiGlTxoIo7nGk5fevQwSV2INHwEICr6/NmcpCR3kGEr2yIf
AKJ3vdxSgZzxBKs6ffPdrjwU6kN9ZJmKUzpo440ux3GLehuGFkycfR+Sh+oo/+SjEBhkB34y51Jd
Ypu9wRrow/ebGuFbCqPgJ2jqKhksCSSZXAxLOnRvutnIzS9TdMLX+qrVfBVGj9BkhkUW7DQVJWLa
FbqFrldTOU0/xyjbI994XL6eKttInhKCqMgJJXZ8hITHEOKU1BP8bJdhZmmDKgqipZoliATfYDLV
ShwBOyJETguWEAZEy/hmtc1Zbemup5gB7QpYjtCS4mU+vXaR48ihqk/tzM5BTpAFE9PxZ6FYdeth
l0ewUJ7cvLpXAKEurrtIExb3lSezvoVZgLdSPd7T1oNEJtA4Dp7kaQ5cvUmzzAbqmLk5HNwPyczH
iFN2DziGTCrG4kXV5IbWbEJkSIF2HwI1aMy4OaiJEQzrvn+oEOn16uG3x7Yxycfnq75NOkoIi6e/
sa7iWMHMTUGWUzd8fDidcfAYskikw7Z50RZWdxkT0Z7jRyZcL/+rIp0TPBz2h3ByYbbyYqkc6hJg
PVOM4viiBhLqDVdr6hM8rwO6Q6/mu7J96rb8AC7ND9Z14MAHR8r9G1CDzwjz1Ent9Q0yYW1Bysk7
LpYsuvinikTRUp7I/e0cfi4dRr0yRnewHtfCFvUHQMzLYJRjIIgKY3gQ9J+Ge+UowPdpNvLDxekV
mdw0xJ3ITWOJh+saZzS8jBt8SLKbSQIhprA+sXmABVxR6ei6iJde7Md5aY2Ar1qncy77GL4REaaF
1Kj0LckPHLdMZQmCaP+9ydPhHY0vje1Ag1A5WgGr7d5vSBvYLynN2ZxBYDCrU1/AY6gd970cvx0Y
Q4UvN4729sSoAiXkcF6a14Tr81hyafESPdW9c8i1nIExsgSFm8nMMXPHErAyZaWsgKNScKZb2KPp
7MHo7rh877RPdf6qhnQqgEiVePn5/Uz0p0f8WDGsQsIsUbmxSFw7i+MpkrrbpYuGu5Juw35rE+t+
VZ8yF4M0G/i4V+Q/qGWEvRlDDQAL1ohZu+79zTxAXHYw/SeAqpG1T1CeAhukN5TlKbYILecd8RWA
yCvU0nhUw833My5VK8Rt0eFw6MQmPun2V1qgGFZ8DrHXpPK7k+9LHdKXDwLcCIchW32ZwtJB2u/0
YyuhPQbgjmtKrttneo1RWa5GBPvjbGC7Ngo8HKuMMw9T2017m4uUnICPSFTG098ZwZ2buzdiU1qF
TBPc+cpJ3AybxjqyFBGCZnYOFIAPdvQD8rFhJbQIxl18qKC6xLN6U3fT0IUpjMSntqCJDtxb9QmF
wsa0+iTYkQLB1Uql3oH9RYIUKt4RXbBW7snj2roDX4ChiFxZJf2kq4CLBYILXGWUCHVwRhllYQUt
1eLGfrH9/Q5NrJPmDWvRKW/p642aDzf9RALaJ46Dg9xq4VpEmoWAPaJRhdtEG3MN89twnguTtwRy
rldiBm6JNpHmnp4OPor4fdUiUg6xLaEGE0Mf1HMnSG7l8lnEO6dDrpXObnyQnbh7w639e46Niopm
HX8CX0lG+zw5A/bbMLuV7GCFuunLS+H6G3jsiJU9eYK9sWknTP1efQR/R4eM/lbn9uHHK1BcGiN9
tAmT76b8wBQeFRNhDfEk1QpXBvVkVxZWuhz21kVqv6bI4fY5RqV3UKOy0NKmblDvbOkD8ihfa7Y0
I8ZdwqvHtatpptt3slrQE53IZgiHpcW4aCj//A3c9uhjucolgXNQK+fEKP0Mkb7zZeho9EodFy8j
3KxSMOcrMGEF3kLiuw43RtIwW0bVWM9bdRq1A9mriYwJHxLjYBffZFcosxeg5/9Ic6Rrv2vSr/GE
V7PjMOhO6t6tG+pwmvqYOYAqAO+jMZ+2nseJLjudM6TC5lA8pJpCmnBpgBPPg37jvg6h+ulHhFyr
sWydZw4Npcsow9Ix0wRoyVmNcjiUkpvNKlz7t6r8VqCdZRI03X1vg/31WxsO22hM5OFXi+b8WGyC
imw6XuN/X5yKPtNIRNQklEkWhICIkSoc3sGFOOT7BNklb7NwmKwJ47gf1+kJ3fSGUjxpCI7/3cOR
o+wJVDAipJPgbdLZX6woxmmXicO29G8JGrs+UzeBQTBMVKMsh5wrzpvtLwtHZhT9KvO/0xUCtyIj
t1DtG7hEBbWfmh0FnpEtpqPt4lOBF7SnJ021GTGK1Okb1A1G1DVWilmhxz2NkmBJqGPJJhZrjnsF
e0aDrKtjdrJAEvU06MM2wKg+dkS5oQICt3ocKmwxuXQs7SX64NmjETYKuGtGyqbr4khOZL8s0o+N
ygT8V9/m8mbYi6Ic9sFoYoTUCLjEBlyFy/3evVWt2hMishpK5wZuNv6Gr3gpEu7WtbxmyqCfm4fr
NXCW6btiQuUEdhy/RRPyNXfd/KAyZLkyvikKCP6vb9SVPNIdgC+w180Qdir2g4zXgWElpNhnIMlV
hPZPyT5yaWsc1DAn9NnYGln30YYf2GWiIgj/U1TuJrUDl7Egp8eiQX3f1Is57OMKE50+QaTle4he
92QxT8I5dFrqKzUoraznDfltl5CCjFCz4EoiwQGmZGez7hDQPdQKoefpVkngdBIWxMTEYf8/UO9m
+ofZ/B+mAtWZTH9VldQ9i4H2UVB4jIH7v3xuz/Kf7sZIWc6wsQ1J60j4D3xm8HMW0dQKA0PXGV24
i6khdAGp5EEHgWn2MKnxogtLwoohxnBiRU35ji4osmJkNmpoOfIc/2H9lsMRLI5+c23umgxWvLVv
WdvSKFcUNpENXOPdwx1lOmkHbYIOM09O0q7+JyWDlcJjvkxROU56z6j6t18wmSXeddSxLRNvH7TZ
6SVwUyF17u89SmU6rj6FTJ72On0ckE+xyQ6K0NFWZGCTkwvwevv5GsWo/7HIFH4+PgDwe+W/epL0
Bo1FvCvbm0UUfU0K9mlNIDcnNIuJKxPV3rlADjyC0e2beV7GrVzF3ZX34lOYXmCVKuDGcwYZpRez
SxIn96u326a1h1eQMhxuyy86YcZFP2AezWS5+z/TdSBEwFJUmfpCNBebzAxIV3CmBysyP+vBGIGy
rjMBSQUGdGa0wbFekRwGp7F3efU+DnWVf1E8KfyXsJcMLPRvLN3LT7Rdl4Vsq6VNpIUdlg4WgLqT
vq1jo1gjEwot8aLJP3lU+RAKHh34hFS0FGxn1yjnLATt8ft+Ir+8qj8ByrYX2tFq5UrvM/8Hgbnt
v4rFhAqocW8vjLxpQwt9cZBDcXl8eNcEPml0evlVYSVbNpTsicJCdV0GfW8ManOqZpwmzeI1E+F/
VhyOa1Fnwc80dZsWON/3WcXETJPMJUC/GGw6hvOyHbTAKQuYLVgdnlqmcJd6rVyBXlg55wOfTJ/l
2yhKzLxh4W34bCWfOgOHfsJjkyShFoVpV1/hTJgdVN/dLf+iJf/G7rElyZTBfPwVE7pRD+UQZnUh
pGD0KnhwWTf4pKLJHF1zitxDVZY3RgeGc6icaDUxZo1Hhpxch2UyVRmNNZgIUWbvg3y5D2546i9o
5iclEzDnRkbN+mLhnwMUPcB20HjeBH+UvgA40dQx/w3qN+vKLT0g1eaWnCzU10Vsm7p5/JyyYUDx
sULfkJZeVhC812VwZ1oDwMr0ozZg3CTXa+MKtlUa9rbisYQ/jGVH6+pfRoYQjWQqU5oK4LNXgK1v
f6NACUJ+GWMSnbVhswt1fzKjVo5wL3Gf+HwMHs8u5yWOjwMhWQfVF5KE/YJKw/PHBGH+WGg8s5z6
2L9kquMmDo7D39EouLTNCJMh8z9vKRMlqFYCdbaAss6rT02IfCT/cTzmqNY3BxZoVMbX7ahn1D5V
b7CwkmNHnUaKVBi3gg/EBMz3tUlnOJQpl0ne+KWbfyKFfQrKhTUQPO2G10ye84xV1rKm61G5xdN2
NDeiC5LU1cLYbElZiUDcahuqOCYrv81yCAS+JB+lpZn66L4TtofMr2MbnE6dTZvlh3/hciCZ8ia7
6t8EQybWMB4OU4G6iZbIkjNPS1GccPeQjx7KKIL0ieQ8XaMt23tQUfy2AliBSnAm5YGZZICdb3Sq
NSUvWXSMpQVQVTlnh0N01qHZvWdSCXt5o4LujhM/MYOXhgdr6uxhxejB28AYPoHbM42Q7QTJuhIW
oiQZl6HuVkdn+W8/Y0KUBUSLnoyc2QhSiYiCurCM3iIxvhWZm8xsDPphy93ZtrQyVrbfiUqOdzuM
sFJS9TJ7FFUcfAIai+xiddk22GRTJlD7QsnOQ6CRkFgZFHiQ7h+/zxDXGqAHSJ1ehKC2+2x6LNf8
tu93N2aBLZY4VG97ll7hgMjCUgTlJkOvcO7161Qq5qL2MbYU/VBaibFJVXf96wgOwj2jSCkOqOXA
PItKLKkkXR2I/kaVlQgdeBrCIKxgd0VDTc/G/DcklGamsRFJ6Z1fHPw9w5XhvzLs9eCXPcC3Lu56
8srAuNdPMuOQVP76dCouKnFgUlCmex0/js02LCKREhoCnBj/ipQzPZvY0/jji4GClzfA9tVfw7Tp
Ew5676RQjGASfDpWyb/hXArufKQ0h/tbXHFF9siK1k+P7JseCZqeMMmviDj0XHvPErD8bT5vM68Y
IREEQc4pHwNclWvpGUk43+cIjuPbBMnaiqsCHi2yFVHeB07AqRYEMKFvvLwIV2UsiU6f7O9BRtQG
jxOKak7N+mYAVHQS0zs5pFULYHnUbM0pRVhtG33+QG/pk8NEYk7bg24B7Qu1/FesbiChFKSTES1B
4+nfXisO0tjTeQNYSK+iQN4FH47twpXT09RQ0tPQfNwH98ZavM0Un6nkPC01DOBVwvZQ+Nlr43I9
hJdcNIJMrvJOUkfpuCA0/KhkoZyB6A4axjl6DwJxQcnF1v+bxImaAIkJ/ecQx5Fk8hHNXNaHb4+3
HnB+9RINeZLKobhOYIxE3nNsbd36vw1C3LI9IPaJl8yKZPw8San8cgHa35pkHLHm5zwdEjSg8FRY
uQ31wZwkx6X5AFNqZ6Y1lQv1cwdFQhHxOu3IvXH6KCQTtxtvDpKJ+TAJTmVcPQzex4i4r3n3Nhke
SggurtD+ta74YYDNdJW8A0+MhUAsCTWJEshk+/OWwHY+PwpPNxjA7ggAWFEAVPjED11ER78VVfvE
0rXDcBo8o9pqbq8AK8470cYlXRUMQHVYtAybHHXyJ0UT7CtNxEIbPSpqmVRsCUmnpp9YOf5UeBAa
CG9yy0ns6j2xOdZfQ7MCk46889GCAhZOvIebRFnkqQc4uGAWZqHLZDxm/H3VfJC0kaAMzx//3TpQ
lVF4nCUUN0sOR9x3IbRP82IvXUiNig1Dr+NFERTSmfHLjRQ3aYhzV/mHRjZEXdKvHZHGby/YSi4P
T4W65jpofYG8Z5Z9kME8Lk/apiLP4CS/VUikRmwwdoh0yusGm4nVQWl4hR4ub243tf5GTXDxVmZB
S7XINQGCMXTvIZHSOQjRRQMZ1ROzKutiWE7at6JUPtl9t6mPgTdY0bgXigaFGkPGShx31gv0ZrGn
e9u1Nlw6WyNPseZcuQoiiep+qKv55tRC7r8XXW9RcyG8OHCFQSpN83sc0XDrPVK8zIdcw9iK8cay
LxLzAmEofO7g03xhaEyiKb3HyzOkFnFSLmhGz/NQutqGvL0JUj03ZozKrabyuZEX5uBfJG4aILDC
g98RU7nGetF0DiMn6PBBIKw9GZ3XoaRZemf83Of274ceRh7FgUZ6bpOTFDQify/pgSG+oW0ltD5E
BQF8k2haIRcS89HTM2sTc+nd0AKbvjUGzqiWEwiBKFTDx7tzHygEc+PMhApA+2ZdVAbGUL68mMu5
5zcnHZ6r6ri6akw3flfQX1IvglPuEZattBCQsz0BlEJsFajuo1sJOgjZRjqd7AVkGWZpHpwLT4JW
zEioiXFQ253HUQxkcCNWtbCzIWDP7e6vNTR6aiv5xtB4Ke6PwV14svu5ZEw9RDXJv6Bd5yGoFQrG
+n/KVsGHYIM5d1NVKarLy36TIzNy6beywysTXY3c9PSxzq50XjWaTy7RQLlBWqYKpypl/hATH3Uf
YURVF61nqH59AKsOWzJHG9YgdQosh3TgbIvzMmJ1YrRMDcCecW24TgpL9uzcfRcRpyAfQZacQBFe
di8Aaz0WMTqCxaTZbsXJVh7nhLVHjmN5+nE92L0px5C5Qq3tp8OX4/kEcqwkNBr/sa2ulzKh3QCK
dZw4sBVNndasDAiMRSr4MHdxqJAshq/iFuHjxxTkNcTh7sdY28vB3pkNZhopbZ/Eb0Ynntbimyr1
GKAOsOghKV8G2V1XJ3wbccmTepeyjsOV4eRVh8bVZFUW6cjEYfNOe/nKwwhk31mRgyKpLnmcenLS
AJtQgd634NBXsW1kZl5dQ0xEBV43KxWxRoZmzK2PCh6o96pEH3saYjUQHmr4U8VVY02oPA8qHFqA
8hphri96lqZpG+zwMKWZ+JtQkln+/tqvM5eF+Wf/N+fVfN5lQbn54hkS06iBVgmN1mw2qcDchX9r
EYFU2VlNxvt+3h8nCiYcA5hc7AM54xUcNBJIPr7ZUlkBVT77De0zY91mxc8dzNaX16CPsSmQ5vbV
L5c8obm99hy+zZCU9sh7psasZzw/7EnKY0cTVnfF7zOO27MTW573o53zlSQ3gEU0xQaZMi6xX8mp
s7OhvykovN4M1V5cadGkGWPcD2VGafRzpN8GF7Up2aissucxTy5A6g8fLQnwuY3cRRPPBukPw0JH
UUFJbWExBSe+fgAUZ4TyBhyjHKVcrgJH18q7Xv4tu2W7hO7H7L1ZaP2DqvrdG7pJ84yHHHml68w7
cKOOr9pjpmNsnFyBqOyvUlQ1TQDwS9O71W+6OLTV8O2PnwIiUNtxzz1Gy6397dYdBaDW6cZ5DraB
8r0pT2OeU9z2fLZIhWnr4n1gjfUOA0vvfZoYBGOoKPSpT4jhjVEjS7tKeL8NFDEeCEyfYgzWOkOl
g9PjReO2tm8/qC3SCm3jmiw/TwK8ef5fovjStOy9lqx2TEz8miviNLoZ3x1sEOe2ATVCX1h+IULi
YMHamw/fGojE/aw3fLb9jcny52Ouzhs5cumybTJpedO2x4lDNjLQjSb12SWznHc/I1kVSdL2w+40
O9G2Pxg3ECGrDG+dClUAfI3SUEg+aOC0SLLI+XcSdvdLdyCcaN621XiAIVFToWPQA7l/9N/NX0op
kLZa/zFqF3L2IvMpA5icIBYx0phmQbvvL+hNQWS1pN+FW+5vuJXlObiXu380cADY6BfgQj0SPJsz
eCPInEPli7Wn8JtK3HS/pMwodoR4nysJ3O52fAdkXNKj/QmgdsJHyYCShaz5Gv9KxXteZYWZfIjf
4hPSEIEcqnRsP3GOtMlV2zp+DDV5YHkfoH878n4RwVRleYJjPK8J9jfAhkj2glBrFTPYlntgSBgi
vKJMbGh/1M21eg47xTK0D4bl6c/V3ixb18x38yFVMapNckUZev/AWk70coWW2xaZXzDWH+ftoird
EDFaPbDafiy8MLTI6vI5qCGstHmdj0+bb8CF7f6ACSysBuLNnMc8xsqTOBxgctwAkSRgGmjLolWf
6eqv5BgBGoqbbbqWYrEvFpjFN2Z0fVUBiFK/zpCZu3JXATr6QbPTqLEvAwoObtBnFand0GqOl9o0
pwJMwQOoPd08dj2UacoaQ7ggxeCYUPOyls00fmUe8zPDUFrUpfL88FQXGWfuEtlptpiaZ3y97yQU
/pIlxz6Xe+Cd4Sc1oxOyP7hejWBOVKLp6aSLhBQb/arj6l4MvHnT1IJRpsWUaNzDe6b/e3ZY2eo7
7pqdrfcQD21WBNvpkXAVDkfGc8QiGGt15KVzyxW60Q3aFG759TPjzmw+2QXVAR/F3d7ZRkKqhqhe
rtCsjs4MxktZ37XHSAAIBI7Y+8wsnmRi1bEUKZ6x7yOF11Yb86KblyI3ULSlbCjWTZXh/FrQkEig
eFDK3vbjun2w5yv0MrydEGL3agjrBRvjd9nkt9z7GGq676vej9Y+trdTs8AbwZwkPyMJg4/CZj8a
LBrnw/mZW6eLsRuFAIXknckIZeF3zUVNPbmMRPvCG9wtDM6mmNL4TsjDIC5lu6ZV4gtn7ZO1JkTz
Avr81TeWyQIXiTMr6zy1OUHC7BAhqt5hmWC7xO6l/vtyzMUZ17M+FFxq8mSrIND18QM7LMcZPoLW
GC+PNpa6MZeLKzIlVMmmetkOYR8HJTxV8pnieosI48U//NtN5kPQw/3eSYLzhANR/Nu9UVVCFUfb
2JkIaRRSiiBGxicbAjV6DINAlqdGEy897VQR9y+XjxgGsM4AM+OXa/q1m6tghlXMKM6d0KfACrwj
qsFoOgZ4J/GHYC++0B1gqheNsU3Dl8fbm0bLDgpT0PKOh0XekU8p8Hb091jx80eo/Tj+2Tn19SHX
zn4OUqJEvjcy6D8YHvWEtgpzHNfy6gct8tuZMY5puejS9nrinChjZo4m9labxq9M4FraU4WntCaJ
CNks1+MLL52VHLgjighTIlBU0oiS+ZMYqKZTPSOhHo9inqNRtUFBLw3EC7h4KjTXYLPoyP1vGfuK
fkT4rtUtvElMYNzYJowOasUNI9ZjvsxSgYonimOjZECqP1Alwh8oBwhjV/SkGFxzjGu0h/kI4EE/
GpMnT7ppB/QLuNgpTjfIzcAefN/YtGwpPTJ+GpqIJtFrm559uUhhp5/R9W8yJzqARxqwrK2PRxck
cwDRPPFea5dH+hPfgqV5NPXzmyMCij0E0SOh0ZWCcu0QijWSD6OEeL8AJmAyznhagjCvHSO/dvf4
xdNBsU+XidTj0BRkNOOO6oGAwm+e1mSgac3zKpa6EMtKat78dFWVGfQ3kdMl02vaflDgZZ1VHQy6
5/FX6bsPHveM1F9ebNVx3vrClBUGGGNHbD+ZUBQbrjV/S7dqyc1dbfuq22tYJozaK4TPySgk4Jju
GImqhjFrnWxo4rsw64cMXzVtqygU1SV8cbvHuADoJjjKiM7fCjBj8C7kPp2FWDqtj5XnvNonnSrc
lryms1L3ZZvIIj9r6x8fWHmp3GbWwoUAsXdBlATdLOpaa+JS4CdKYE4lSc32dMUlczLoLtM+Du9H
8pc9QCntoIVHVRGlT2fnWXxX59egdivOw2ljtE4hwA0+8244oyWUHevlXGcjGVlctGHxxBfBtmwA
jIA8P3Yw8++LVxV7Ild84J5aOrKjJ0sbAY+p3nTZjdXQIW/9zi7fRP6DBycWJGLq0wuhJ2eEgAuQ
H1jvVMxwclhxkrVtiTAXC89su2pADA3LCQmXqony8gqrs/Zo++plzz1uJvYzixl4pPJrI0/zgjtd
XlsK7l22GWuHwZp3MFi7mAHMZvv6h2nDMQtX+jf5beNwtpajStem6ciR3oOFqPGgOm72Rjpg/CiP
X+tMCrWktu7eYwi9n2lEjGomHmLxApbcRQbqVLkQRZfd1+3I1L1wYmAlSfhhN7/qrj/+MJ4IluWp
oWCIqXBGj9zaHfEDHaThcilgz5JJs4rJZeeqlSxG5+5HLfhXIeOUnruHaUBTNh1sZ+ANzxBY+/RT
VwrIuz7QniNL6Ky68Gp5aedR3KH7rUM/x0G9g6jtEfeUAmJnL6Lt+PT6/7yBtF3QLl5o1WWCQElg
Mf6ofCv5SoJMOn80cCEQSP+17F4ARSgXb2a7bcn5niUT3Z1V5dY8enDrFKpH57/vgvTIegafQBPQ
O0Dk0U9a3jFze3rxJR7I+Lc81c/w/m9aqRVK1VX3/dMMB3Qo1xL8Q2zXDvwhNwBw5ADCTkMTvES0
Y87j37YnvCCgySckKt5OCrxrgUrxidvvyTmTdIM4ZJkNL93Bw7q5hRiMeA3b0xTYmBSihl3VSMEj
zN+G8Fv2dEGXazFUmuYkMrwF0GTL+QrNCI0pgvjsRITaim9CSWEMc5PmW2OtRrjzDm1doM1qCvC/
AH88gnOjwHAJ6cRfsE7a+kr8Kq9nyJgE+AZF/Z0fD2vgw7zMPpkOSZDio5rlHJyQU2brXDxj/FuN
ofhR3DTsAhB8JhSmWreaqBaG5J5iFpfeHFafwIqR3G2hR/7q5bpdYsH5ihgeDWtPcZfo+5LPaEe6
NeZoAvD19ulfhevKajgFvrq2o/pPVWSk0XTRTw9EIx8ZQuSbLVAXnVtaj3JB58aNIA9cvvg+biMr
C3mMWMriD1AiiSBk5c57HnAftEomaENlmDqsPNnVSzAo/Drf02gqYtABFvrvo7cVTa5ZgAx7Mhbm
rnF70D/X3aFaiX1qv9MF7mGYO9EEDA/T89RQNyb5GTmYpFtJYM/14GVl72tu0ubZr+g03nsw0y53
8x4deOufkigfwmL+D8wJ1gIAEm6csLfEpNuR0U31Ko8dVpr3sduyQXDXltkpwn1MrWjOHpIR4obk
30O8NdY67ZlMQ7nQ/n9cqDb2xygNneBWyoegDJTMrdqvoihtPukdaCJZyTyWKb4PJc7R6kuqEwkC
tthgDGl4CRt2UP37o6pwwS/bXP5vxz70xsKYSraATcx7a1zVeFkv/ub+ez/kxca0Vx3783tzaMOm
PZA8RutHJWkuyCH5rzPczlogPIypWpBGsCpVsJa0duaZl1CLx+DZucbZgfF2L1Wj1vllItCdqw0r
fL1K1peGtxMEeHNk6I+mHqwit+SeVDhcpwMMlkAF2xEiTSBk6VL4OqElD5baPXr+2Qlj6IrLoqYn
ujSPidIjaO6yRj5NmLadyk4XzClUUzjxBYRVWU00eTcz8AKra1Ujy14co0xb9YMjEo1a5j9/LxCd
auCrP4ZzuNhkh+HIzS7S+jM89qQ8zmuq6u8TVyX8KircA41HdCwxDmHUR1w52o2WsGmgkf7j0uTv
3muSbKMEBcmlvCrppvaEA//Rhrm0b7KK0ZTbq/BndS5/4ECNx78cVfwuPTGb2tBFtKTqRc8+uCdG
TyLoqOmrlusu0NeiEnjxHSXGllqqZzpaMItQ3UWUZeHE5ULlScoYEo4njZROmVzdkVYHM9YD2uql
cXpLKsWL+aMSiRUyyVHKCmOyjX6BnOGNCMMAKJlfIECiWImHgU3lt++kTxNg680PU0hvnfFdDWBB
ANufnbT7tcj6M214F9ZJfWuVZ/my4T9YAXn0nM+woQ/QX9yjQfVWmrX9AF4Mx1oN66iQtukzvVBg
N3279zUIgRbo93PEbvmKeAfcztxbUAVEdcrGFbUSAfAE1k9ReIrUZuIaBBc2OEGgxcXllZ3o8BCV
Uum+JeECfW9qyropPo8PN4dDGDvSQj9BMv+kFnOPYr6OnROVx41DS0+AVTlcsqX179eX6/haALgU
R8UONrJTNhOLFTYbMO7iRwkyjKIhlmm4NQ+Rsk8LVjKoxTCK1Ma0K3h5ygYdop9cjDEfXwRakkzp
rJgIKWaH+DVrWMpM6rI07192hUES5nIKOyCj3ufwWMcREY2E7G3YdgeBxTKZHALk7hPA7fYSFOyC
xObyu4AniQVTo/6QKGKH761FBybki9BGY2xmJxBJJ9Q3gyBY7j2qhXFx7Sx13TBIYG52Cu71zuZ9
4h0DBgmHCMNx4YFkOyeFpYDurLx8MMHpCL0psg52Uln7kHeMRFKjr+ENrGln2WaNLcroThHg0BCW
qizGkzmdLSf8Cthq6gb5RaDy3h+tMU8BALafVpMHM4dlpLTG5lltt3a9JFxCPaNiSZ+WNr+s1VE1
Dy/fmVfDB2sYrP6mML5pkZxhGjLY3yke4TROkgWdvJuSQYBGcvTZZPF9nkdI/oIH/wGjHzgEC3HV
93/MxS6JMDMNmv4i7nM6dnCiKBn/dW/4No8+3K/YHoEoRYd9c5+X2SQZcSXRn2CzJO9TMcfyFFgJ
iLq4FKgTMC4FL+UAoegal5cfEPhVEhRLOuptnjWkl+mTtLCZ7ScpLq3qxzuaeAvXoyLB4UvtbdTF
HrHfqo40an4sOUmKMrW7tDAtY0dZCqmzTwmEvA21SI300/mcO83MbyphRibB5nMlQesJ/WX4SuKt
6xkZWPB/gfhcWKCrncuuUfz5hRKElnsUnxTIJM7NUmn36aQ0xB9oLAQ+JvVRhD+G/Xb8KDO40iHC
aHzFLwKDU4NgtiKqKKgQmqTlMJeYjvDSjAn0PeT471OPcrjXTJ7auW218ilftBf16zAXqSja0Tow
AeSAx/i1E5iVQoC9ALNEtguzKfCKjkBOKVVLv9ecaTLaxX+qUsGvdVvNTB5bIpAWbYo2VYfmqDDH
WFFL/G01uFYARcFlCv2Rd1D9lmlN8JWVMX/PORNT0EgOjQ8nSXmz/q5hK1kDUDMjAruA5PCdgAxB
yAIJhxfd+ZOgvUqPN94XOTa7+WhuJy2dagLjDmnZE8jNZe9c97soA2tEJJ+3O3yD4/Y5QuJSBAtm
m+5sPbBY9fZm1lCVoMem/98tGuLp86ohaqH63/IYtBtdjdh+mP1YASN4VoGsSAX8hzRcW9WvrZoW
7u5VejHvtswVrKuiYgmPyJHaT3RD2ddToXVzfkOpAzQsEpbeUCMp1Q94raJy2BO2AQqReW4dd5LI
Uf9ub/dIFCy296JDWh6wdig4rVxb3sZDg3ZRveMxRSlzk1ecj8aQpfaa/LaaI2OF+X9scuA/Cr9j
XJtlD46t+0nzMuYP5hYS/jsy7p8dovbfBdbv/hUAbOjpjjBY1RsgL4CW+eaorwVb9ISoXaZul1Al
y2kkRqM6iNx7bmw952+bsMH2Zuptt3L7o1UBI0BzckwLDualchjbPmmOGFZ7yq7/yk3tqTYcGjUa
WPRg0ntr3ttA+OSgu5TWl3DK8itz0d7QPh2J6HCk2N6CrE3pXrysrLy7lPNIvJUyAdyL2qJsNDMw
9lhJq1U0e3Q352bsrde2louk/1r1CMVYLqgb/5sVGQeLhlzcOG7OfVQh7Q30NZqRAsMh0vsHhuFw
m3Ab9ZT2eAXuqJrRbIa3DangOoxxrorLMwFtPqQdVQE5q/tpnhtzbIRBqL8tzY2GecMhVMPZFu8r
uVJQI1Je0yupuFSL/0lhOC7v6OrWG+ka7C8oXdTqHUWyBeqWbCgK6bxGIGAGv/xn7ZDqs+1q4sCi
yYzg6tPclfPDvxBmIfMiV86xm0LlwoUmMvle4nv4Hjg+AbNPn8GSNTkmQMDElgmB/m4uhwhksxts
vm7akXfIcERinZqd6LI9zY+DzKlKoNnzyH90fJB+aqB6nouy/O2PF+evuC+VMxSzpY3thE301r8P
m4Xhff0fx2LXiRYYpcjd/G/8okItG86pMQ3Oorv1D4uVaoF59th2ftRK0Zo29KjmHEf00Mii9Clo
JyYGkCkYHPjU6UIFl/vwt6jJrUYVLTuq53mXIo4fICVSB1rW+f7scAzoOMkSGWKIYouRvNs/a55Z
/uYYC93wc3ZgsLdJLaEad2F4+hMVPMX52Gq8ymB3dsdedTDSmlEubcFjGPlo0lXdRx3lwwSaieZb
dqUsvo+ip4VUAWCseEV6Zw2o3lmP8bibHXoXKCzGDsoPh4+oSQ2haHlhaOEDOF41Ufe47fw3XEdD
+EiePRkUq3MRi3K17BD2erbEQNymERpBoSBc/6lrMSksm3XD29oXFrFqZCJQvmezw4Xf+b3mQOJq
29AOqpmGf6HwFe6Zab/u/P/ExOhwflrV6O90Ta4F0XsK9jUiEPCTH6TAHc3rxvChx2ErDoYj1Rrc
h23sxAYGuFR8BgE1vHnmaOvcVdOP1dxRhQsLOxpChYikwroC5UQBlZa6uFcBDNX//9BSXjcSXk+l
t944VRcvRzH3xHkM8EvNH5z8RcBn7rAOK7CH4FkHh/lfqhyppPaI4hlCm+vcJDFXCg4Pd/AtGSvL
ssRf8Olc1XBdSzGHbNkM57fRbR5L+PrAN1p4ho6HgrjZqx10bFPun9LT2FNruMPkgOgmKGP5aGDn
KxBVdjQDe/MaW7KVVJreuVf5VTjK6dBv3Hppf77+r9FOosSjA4shjFK51Fx5etcsh+JeukL59GRn
iMNVscV6k040m9JEopdG7YwLHiaUjo3zRq/3VDPFcGLbxedGbvfTNHDUGg3+IQN3CEuGS0uhtchA
1Az0J6r2lnR9GWNYdlJrRK5vESZ+kTng9TdYnz4PU6wfEt9UmXRksa2T2EPsfBWGy+NMXXXvl3ku
vrqkisryagP+58mySDp/2YOFELvvFkv8Du6DFFzlcwh2XPy3mJxEqQiB9MXRP64FeNTiTv+h11yn
WjxfzurAf5vM56kPX5MFzkpMz8b4Rh7r8mj+ymVzu4Lf5/8FjHHP0ut51cSNWdWPhCTccc3hLRBq
GUt9ZcNwGjywSuo+yjpkthJultK6Cnc00G4cKRkQEW773o+VzBlg0VeOPTMfsR+v2ZkSkne6LWrn
2RCAjdqWAy5SAktcq0fSy7sBeD8USiEcXdzOuFTMtBSXd/AJssai57kEmX5nUTfOMr/1C9JfdU7I
od73x59xFroPtZ48/EbYydpxS1qULUdq15X8YhYCeNzy0AvGjptArdrOhfafKNM5u6EB/oa3M5CP
gXQh/svuS4S20nWaQkBpmyv+Jk384zm/6/59cW2ieKUaOxYgOVk4pT33/B76Jo7YxXwXZUgJqnHq
NXqh1fpt0lKzLOkgtof7IaX7ke53TXdoqUdY7VmGi8JdIzOzugV8p1DfLfV4Tov31Yq/dNUGvSnf
VoQcDz0HbhGpkBq822g6OkhQ0Hro51QTWI3ejaQVDgVzfSW/LSFpJchSBevn185hGjP1Sg3dh6pw
/598Q4sIvOtk4G0aBte4zzE6rY5ChT3j8ZJ0u98Cf3RsHubNBTfPXZdvMxVpS5Cb+YscV5xmqgGb
2vXvqqKuEv7N3vHScrwIAgYHhAt3XTXXteMFjLmTcGhwDej1Si1PU5YI5UV7kvEKuL1ecPxMb8WU
9W3plKGhROU7ymCACYq0k4oRPGfxtwh7/Tj3FB0IgT9CBuaVousIr1nP85VsnNmMnS1fuL2SBV1/
S2hRm6lyJiRrHA3p4t/NWzz6CReit9C1SBjKsJ758Fw+UnPKg5Y7Yx1O7t1eewn1sAHQQwcSXPTr
S75XHPmeAtnwqd63o//sf7xUxh33DjLV/l2jFRzoOaoD4ycxHVIAT2H9Xgdw0wGfDlk24qf2dDED
Iv5nu/S7QK79RzWmhZSKaQIv025SY6oj1aH0dQaKx65dmiJnYcmjQkd3PXtrNvStmpbX0J36sl8J
vGP1cw1jCailqkAUOOwmF+tW9bp8VCnR/C3i8g6Wrjgp9NIlOwB4dzGSFbUJGh0Q/FWtLK0p1P9s
ofgMQTtcNW4B0SY5BHKFnCk1PXGB4ST/EFkzZHPDo9SruoJZ2dg+ijIKxx3c8XUwtXTuFJoqUbGr
GhlNP5sOB0T664tprv5RBtVAQlSbbKHE2xpApjcQx2CW4zU6BUsy5y51i1OfTNvmG7A/ImQOU8W+
+hzPI5nEBjgU98nhXIlwmD8jP+vypkGDz/3bbDp9UfcMfplQjt+ivnH/J2OVpwIpt+mbEHXMYHSt
2Dn5IGKRZCW32lNKS1K5Jr/B+dVt6fB3/aWKRWdne5VyJLBvpZqkHsE5IazsHfgvsz+HIaMBxpsg
vssAORapNOQ21f+UbqC4pOR1/EbGRF/23OL/XC590nSfzpLONO4NwWuau90YOVr/iw+nHi5h5jYg
jFL7NUCKa9mRazkwPlyUUsXVLt/OoJmjYgMlvul+me5vE5WbDiJ3nubrRtCMlFAQCMNIJPsfyhQW
2OWVhOJXrl7EwOwt+bO02HNPorB0IUKetVy2ZyMDDME0Qz66v/14UBc8NYNOTqEWgdKXSiM/qn2o
bRoP04OLsLJEe3LHIY/e0M8wA01cfW79ZI3f7wWV2Qnd1sM6SPa52X90exOm+oqPkFv37FpGzXBL
l1Sdj+0GK0qh45TCsmvAOSDnwzk5EgFf0mklROkwSbMMnL3MDycse+C/gWNwhu/AEaOdV7Pboe7/
0AQoRpn/4nViCRQUmGbcZYLQHvlNklCoLQLQP3W7mqomVyLeOrKU3Seyv3XNeXhRwhVtwUKoOCYf
QZw5A4dHkDblU8tB5kCzxC7FoolDBjm6HeKfwgA5nxkYfSHzUZ7BXnkOchQ+eFwh3Ij+eaWldmJn
cMcxK6nXEFY48w5eWqGAUI9QXrqV/ZZv2uHcQCIqlykD0IY0py6teKR2QPcYbUl9j2WQ/yLIXN8H
2QLnD18TdjzxFmdoYsTyW+iHfJcAeMKigO7T1wg2d/qt+CFm6qSGPQ572aRpP9+8md51U6iPQV+s
G0CP8LX4zKPNVfvwD8jHuWNNz2XOiMK5l/fOV8iXVlIeH4L4JNyYavk+KPnp1S5va41g66xEO0Bi
RW0TA5VO+XDVVCw46dda5D3BOwmeX16wOxDZtFw2G6Ct9wntPit4Z6IdIFEVAsJ0aSJC8IYB8LDf
BKRw+7IVrcfdwYzoFXeO9xutOF4NX5nxm4bM/i9MSsO3umalAgsdoDS2qAfsGbGqh2WZdS2a2lzf
Omlwu0kNRiceU2SUY2ZZmr/lzCLky/tA/2MacrInY032TkyKrW9y+wf8o1aI/cOdSWJtrQzmjxV8
HNOQVkVhn38PxEf5z8uP6dnHW14Q31eqfBREJvF5lfJlw9WwGIHNHzm7y1ytMPX/5eUwUs/UfLFt
S9lUiXu/PYqSPLyf9LsFqNa1+1jTuCHpgJf2K0Hj+ykRmZ7DPMgLtXQlZjQKuOiu89C7e4VADrv2
HcifAYoX1C9Xe89iPKA9K2+FUUlWQcLxaTTJk8AqdrvCNhm9B0VQ/rKT7ZTxMiW/Rgye5qF454C5
g/JFlgtoiDuTnr4hb0wFo5c0aHvVueCV+6sp8AKdHvq7PBaBNXwC2q1v/dlA5JbSnJUmKj55NCIO
fK4O1+Bx+1htu/2HNGRGwKiak5klBJF+qsBD8njcYVsp3wPY6ZzGeit7gjYfbisu1v8juVMGOa6U
gFN36rigjuI9NH4Cnbmso99Oxc4Qq1rkj/G5qf7AoJBzdR+4o+edgLEPfyeQKRLjjBZ2Kd686Ph8
6ktI/579JoOBuBRo1Ms9KHcPeQkMvKQeoBOfYGL17TQksIf7MUHBXHCBCnFPm95jN+6ZGTdms876
HeyoNzOCGMEzVCRAkfUmEXsIbsHVuU7TkxKE5WRSiXVh/0l9LEenQ7ka5Q59b6muHGbdCoXi2cKX
CserRrFn1zcqj+rbDvdWAdbqhUFxYVrM/IpF0gPuwzxW8XSik9bLY2OZZ4TmE0U19Vul3GoS3zSh
9oTc13Yy5M0E5SEIZTrJ4jz+DDBYgxencoSZgKCm7O2Qm7elmGhz7WKyQfFb+ad8veEIkQv8gdFJ
I48VT6ea5ZaN2QoQpvNVnm8wJfKH3mradug4Y0I/1CsdpwNNuGwfGWe8lwNA+0sWvSeG90EUMT0L
UzDcqNS1YSPOkumwn9qibYVpQyCoj80kKeSzmw4baWdabsUo0ovrdGAkbLiemt+pE/Rc0SDezuDn
pRfNEMChyujtP1myRE1HUYSp+MCsq0iKAK9Ycy/vMUaX15ikAL+2uUsHSnvosOIltuWQdfYeU0AK
nyCekiZ7fMcmKEgVuUQnDfWfn/FO+9TGfkShTHQYJxFNUN0zk8vR74pvi75bNT2q7zPv+d7GF00j
c80LNl/V5hfW2mkcx4goBqF3J6bcQOh6vORJK3hhtStnqke3G2b081QBsB+gCZLni2n0StCsaohU
kigJfE/aMV39O50d/zh14QfZOGxtoeO8wzIkXewF9+bjZveYJHXEGQCFc8ZPWrSYI4c6++Ml6uQj
9Yui6X51SsrommyLa5l5AcvoHaIqaYe5qIoR9RVUNLJbInpXogFld1AbPqmqmQdaNZ0gC86k38sg
UHgNHVSQaql4q+TMi4vstJZmSpSOKFIoCbk/kOcVUmSdxv/ivO6w8t/7S334uX0as2tlqA6t0wDA
WOzGLPhkQuvmEd2L4lRZd1SjBsJAyY7e0FQA249K1QmgkXiUA2P6coa5zTo4cV7JfKRmc5VjHiQc
BE3Np8aCxiwmmJlpKk48AnPqqloBKFBFmAS0uy55qJJHrNF3+3xsbgXJGzNJj1NbDQXxnFPJtYMz
e9fqMvjiKYDA07FBSAJZbLQ1b5UF7JcgyBg8QfkeQc/XLIH0KrSQvzLSwddSKUVBMhsfV6U5vgeY
vmVofWgA0ZClDpXn5o2ZQAe1IttZa9VCVTY7S8VMliA/rtfGUCB3OTJRi38fKZsCi8AsberhORzc
+GlI5eT3wMM825tlYhVV70QuekAdufuWm0ITzO8j8Mq6wjR9itPEhAFktZAhjmAyvDNRFdqgxJM2
7XNKA/Za9czch3LwRKGLBr2Zm6nT/RHymiqKq9mWwB/2chetTFC5zO0GYpuTsm4UK29x71OvLxAA
6Lr910Kxjjwk/Rcb4efeSSQdtTZzOrxlxaUps5pewS9GqFRnLtW3ld06xoFurxp+uT3usmoySW9w
oyhRAsCbxsSv6Ra3x6uYplOv5Dj9/0+RiZz3NXox1YZuWnAhd+mx7a+PGLle5TJTWU0bd9gIfIDK
C5VLFIpU3zNt0wXYdDdSO9IGW93bN7dJnTHuj+4wuQxOvZgmy81eoUAoiu6JqHBCHVyq5hcUrGtL
bB8yhm8C9wq1Th8mOvuAivWLZQyaNE+dSgI54AFvpcacvUsTZiv3BXOB8yDec/aVdnt+vWI0AE1O
y6JcrCdOwbZHcZ2d33dJ82IrfPdHXN28kigSfS9t+ifthBQ4VC8NolgxmhTmER7hmXmnEdonbaDw
7lOrDBGAJ1UwTcyFahGnvsXYJHyzAgJl25S6WLZ3NGf4HKmyNBcUdsJWT03mA3VOb0Ig8LSzCdje
0io7ANgVB1w8efYWKz3I3jssj0NgLC/YjsEDfzcgkhVb8eTkzjtPYm02efGNaoBsdHPztE2OlMrV
7ULrsezYWJMwU4fCA2y/g7Ia01b0FmVCn6OWq8SB9/RyxQW2FWqfV9y+Uq4hHLcRQ23KhVl5ygjR
lfy57NXw4TOWAKOgI8xg+UBBZudDG9UaNVualao+LHkhIN4UdC8tJGK/Pcb/q3egBJLvmAUjhDTD
g+KdnMgBsPi2oxKKxVN6nytB1eT147R4vjMqBXS5HRk7S6+aseMo4mAWrslB6/dWVo0Mb3vAh6hU
UYoFjbAHP1X6xDoQoj4Sn1NKkJHnHxeneyF7DiwlRftSyZXBoSiEwmUBrrVJn2+kwrQ/hlPs/iGH
wTYXxBzJwTCf7+5I7ZFd+TkL24lN1QJkFE7l4fiRcttIinABtH6jI/L52Bbru4TGajvd+jf2cu7A
m1PtwyRKpFh4UzP/sMrzs1pcvjqCI+3Tjo148FJSxAspf1uLmWU7zKIDlbj4AoypRmwlgzdapNw5
PVD6ezMzOGDIP38sWTq6VWsRIvQDW33Dtv//qYwQvH/+4Q/TZOkCgRnstS+tPLpw9SXDAeQLckP6
wMlNSAuiHBrfaIn8qeBQm8zb7te2JOjezPsRdlvAZujbMLKAsgqBGG1GOEKJUMhEYjbTJT+wVf1g
7pEqJjAKpxKAY69KKY0HfQ5iTiZjOsuzTzwFAB94bppDmroEkayYMB20oIeZjO1MNJC1nGFLQ8cM
GHurEkWPQHtinyfT6V2i3ZsspSieN1ofjEvnU2aV1rU91YKWey7mCoUrrdnBZaqjO3mYaPWKlQ2C
fwOVT1KwW+/uYuxyVcLkbdW4UXAob1iSVyDndgW08vnMPXF6AfFK7ClBErL3KfRDJ7p6q2WUt04d
+QAL6tTeVyxTb66wsuWitX8+IfE13rXD24bUZS/rPJQgSZwAXFjUoJjlS/hhGgO977UhWvsDWMWq
Nk3hHbi+L1Ak2+vzBareCDCfWq6zu5naefAzc3Adld3V9EynCPj0T0if/87v+isbvnXi+qVWEp2+
JYb6HQLE0VzP8qBhXieQGx1a3fYM4F6IILquGJBr7fHyFO4cOjpZclMo87NPJNgyh4qWtmHE1+cR
J/0gxPUsNYkaUdRZQHyteguaaqXpT7Cn/vJJZP7lHJvPE4slsdkjX7FTUPWwLkvQVnj9ddH8llvj
NtUxVMXCu0UBQ1DMgxnFO6llRBeOxbc0EzE4OfIxKHwQZtr+ZraLer7IBkkC8yN9abCoXLWB7e/M
1/XJlRnEBAyiurdScO0BKiPR19Lfo6AKhavVCyACYHoCjsEuJnZoqvO9FAXBY5OhDBBpqfcIClv5
lCI9krvwi2Bh1TgaQBa9qvX5g5d5GZe0UAG3/XoniDgqOiu+thcEY4hMqQBIlugt5RDnSdJrcRya
UMY+v41a2S+PaNqI72b1dlW6RkD8DP9BpCZP8oAGSfqiMI/8nojyntcOPvCfyx/lI6InTQ0I33b7
THr7a1bbOocw9Wr8mOVtKFogoJOZS1b7fRZVr5b4sp98kY9bCKoKrnVjwAP2ZWS0TGKQS9ezCsPl
1woWulRou3efdeFhDLROIyHViZKDEsUspKM6POuBByREDerSU3MY4uJZvrrrY3i24CGV1Gzd7Wj8
FokQVMSzdHqeXA6zCW2ZtM/9lu+eu3++UmhZPWKKolyUXytM6JZ8vo0GZ7HokFAM0WIUqRrJ5z0a
dazlthUvTmiYbeH5g0um2Z0tkVC4T4m7aOiJjjUUuNZ6B16nuoOceXsuNeyaK/6LlB/sIrOtXAL5
VTP4YWa9K1I+CnR1PC9n6a+PJzvmqPeKOJDaJu52keXPEGXbtL/6sGUWZtGUWpsnHaEh+2eeJUTk
ntuPjJI0tYIG3/0+2ZShmTIC4iLg2uiCwG0e5BHiYFLvHxeuK8SaY+2K0ASSmySosFlOuexYDkgj
oQQokrcxSR2BNP4sZOrzQzbW9ffrCgF30gdybUfDSan8mq4nyIRI5Gu6I9/JoyP04U/ERQuBjwPx
ieq5d9w9nmEHSG+44SarOXSsTuOrHqHOiXCDYUthcJf+PgdtcYBz6cDbJG1OesblCQAZFa//cq92
IAvNlVAOsecMrg/zBnZYOIQ5vHL3hCHJGAhrKTvhLCXmMCK+m0pO5Xy2U0QdyXDDcoUfTjfw7XLO
42FqQ1SkHCFTewZhHE7VItnjiUp+F+f8Q/cnfeICXMPUe1UC02jXFNDlbYASsi3vv5M/dFPQwNZt
VYJco2sgtCR+LvgafEJBxMKl+lgG2UPyz0kQzMH5NuzqwWnb6SdKULVCEoqhxiT6mXsRRbCI+teW
MTIaNykP6F3zJv+TULpkAmiX27YafZCXQyau6FMKZtCn9KXRq+FQfZSnCV+p8s4tSdCXIEiTGzHs
W/j91In6gphUFvHl4P6yXK3ao1pFPiN8VfyqJXWTFwrO75rFdjBB/tVRXwd1hI+Yr7k8Yy0fzG0P
h96vQ/11t77JbbGzr2gLqPfGaSTgrRdfWoYHYw/tAYt027DJgXYJvTyRzOnY9cnDM9EB8J1hynwI
2w6xUgZW6oUCpTI3LUGAiN0FQsF22sabNo7+/qxjNebx4swqqcGWvcpY9NK+3z4lChWNSR9+3jfN
3XYzpGnl1Y4Q/tH4/RsG15rxAvYLy6TIGVTAgqVVCnuCeTmLafW76mMzR+wgU7CZtZxn2h5PIJur
m4eWOYCcmP7WGZKX0dgplbbSXwlJFUHmQYUuY1gNmT7GQy5Hb50BtnkCW4/KNFLjeXqGKmABlw0z
FmopwhtCDWkES+xU2M4pVgeJkCUODoH4R5fG/+pdj8zdQMRpzFgcYc1tvPp1xSbfgHTdfh3s8M9J
+IxkE4CBArnks3Eu6XZ4xLuridorWxU3j4DyAB1sWEvQuc/rV5WU+E0lzqfiSmv4eaAn+rcTqLnU
NNy/7R8b6nZge2q8NIAv7RzPsU86rFtojRKVprKaFogqLQlTM2p4uy/NDZ3dTBcCvmVWQRYFCu1w
YsNLDvMlSGeiiY6KTyTDCF9vs0mRQK0lU6fhtKglPcJtIdTVU3vMkDE3hFuyZi8t6BV4WD0vf3VD
krN7ElG1+5vRHLcI9SpcutsFIPudarmzCmxptUyoARTC7tZgi3tkoc1qKtlT03Wj1sPBQ0KQO1j9
kPle51pn4nwqTj9Bh656N16bF2J0xKK9ORoFnHA3r1/9DEjf91H1/X2C58+UmZf7axcUrlsxn33K
VSJUJNlTM1vfL7Yee2ttzJ4hrQ1yB7E5WBkYi22BZKGrzJaIO42LxiYjT+Bv7oyqxj8bfFv8z4eM
BMPWU/w8NxXZ/5RR5da6xdwwkHw50MJw8/ntGULiJwUhKwtMqfFwuPHQrZIvMUMcJwvXnWtXXiu7
xWMBG+Z9ZuJNhue8vilmUBWE7w+RlsUO1cCChrqkLZAfkzqePBfX2uwQ44qqzQbIZ3eVaWxRGCwa
Ce01Rp2WPbB9f2cRl6OBn3EXG/4WpCUF7PrMYr4Udmj6UvLx8yN5ADJ4MRfc9LvjiNpDOFKRowFT
tkkNGISajac2vBvQivzCFLK3XNnc8O6DmMbTvYpRCiHCy7vyyBwB1IgIMm71MocngoAg0cTZJ/7B
Z5YoTFD0Lr50Paw7kyG5KSZ1mq+5W8TJG1tzaTs8E8z618UtLRR8JVNiMGd6jUk09kfiCcpNUSFQ
hchFQl+nCNYPh7bRBD4v2WBoDBWMQdMOAsXYdaWcIJpa9kH8FVsvIb5Rp61ACowtUwMkfvZ6uMA6
eYQNMRQ4EiF43r54N8yoC+1kcEGxB2WNHweIc12IPpna3U2Fny0g6ORaXYuh2lbQXbbGRRAmQbUo
Eaqpuj7EtBf06iZJbmtaQq69/NeVd5NlGuzOSitZuoRlXimh5K13mjabLxKdfhoKDr1cV5Z36t14
Xmkg5KBWa9FlqbnZLOXdydxi+0reBWs9X73Aww8MuWqaftRz0S5aPYVYhN+9dH87irHmABGFzNDb
AVByx5ttr8+OEivshJtMc/hPQGcrIFjf91uGu5wuJKHOp2/nJRrHwiitm6Z67hKOZky51znGPItJ
otLNN7kjdbDRzWEGHJlddGaawZjNeAibmQ+qTC8IJ06kknKxL9MbhKY+HKa9/K35VKh/rR5xIf5V
xN0zEBEuwlb4ere4U437PRQ1e3sC3/N0YoXP72Wg9CGnHxbOi+6bhC5VTYdGwUMY+LSe54UIoojf
lmoHjM5kAHn4dSOF+dmy3imzbfpoVxUrOL5GPSL37vEdHN2aIwtr2bCFFnvsxoTNhI9wALB6B5Up
r3QrMAcXvzj4S5QGJ7GRmJeUuAAqGaepDy0WsgrhixYT5ANyyqI9FCJNYLVdgBlvwkJd5n7gv2iP
UEz/iYWI0tADL+9p1HMJUKTdtnhIogLzHntS6qqGCXe6tBdHsOX08qNrCTfm3AIzuUMPtYS7vhCC
nDcRp7k9DhqrbS5PPGzVB2JN4BUjA6Ew0sQ92a6GSo7Q1MAFdDPY8xawuSCSHcKOgUCcXTC1eblY
YBMRGozWi04wpdyv8Y4/2OD0I3OcLE4cnRUtG10gBgv/zO+xTH/dyrYg7e6sfeWtO4nL5z5gKI1m
PxfSEbO2dMIukyXrjJ33ZCkW9IfkACXvsLp90WHP+atGmVZVlb74nO1j3Ovzga03Ut6Q95gJtJoa
OY3wMkWnJVe8Q5VTEdCFHdgWE+Jfpv5EeWIl5FaHf8KKNyAjGnhhLAKb6ACkvzGaNVbT/GQ/bkKZ
u/JKuMbIbrc/0D4PiePIZhwXEkfIPg2yaX6jRLSnQRHmpgKRDc69NyD9jr00yJlbBZnhY4TlrhBm
4yzaRKQLDHJBGM3mGvzkbwozp/2DBfXSZGxU3fQpiRr0jf862hjnDh9cla1RcP/4X5vRuvwHHXR3
X5KtNksyFHwr3JAGkxiWha0bcr7TADU62eUn2AWYlEnsHHpiG/oxAwoJd3zhUilnuNrqOhF+OXfA
BoxkagOAzam6qzx7Q00/1ZDCsSYTUWJg2FIzcD6lK1CSjRTt4bhwGLwXgbiOBA2rX2ZhUXKqqyXw
mZ8coXIE/SObS1pcZGOtmGhJXFZkCWpPamhwm4FGKlb7BKwMsdw20CYV0Ggxi5kyWQVn2Y9JlCEk
owFY/E/FhSVel8aAe6ynrdLvyP/okWLCbQAQZMdiKiyjYPqvpt02ESPbanPtF8PWOvcCjn6sEWjg
cf7oHthC1rUDoOTj+BOIeLvfQbgKjiBrAwhm5vKXFbBzALJcncsH92H2qTyWznujuBdSQuS1QzmN
L0rt1o4XnGtfTDCgtFOOtwTlo2aGO+zPJoM1aX4aewFWrhl82kstdrEy/dD3tHND2NVolGcXGCFa
7Sa2juUsIi+cFMlj/0IJIuvpmCjcstYhQjrv/TiaNOjDwzdsQxPQG7pA7uzwosQTHiyRpBmXvZlr
rG0CByUjqGBHjejLlktEgzAqv3cnDKgf8GbBqXIakhAhWDYTW/Th6153CrGNb9JMQyfbloPU/54t
4x7RuoVYiYoHEJIUq42TkAXxvBK8aJCBz66L3XUJGUP52eI8DFwN50xoQUxgvG+aZ6Opa+0uK1tY
1drHQIG+X4BpM9UTuuReoU2sqiahQF8FGZssXBYRudkAYJ3I4tSctY/4E3SuHqEIOgGxBby9EYV9
CHFYi2UpUbbG7at4c3adOBgKh1o8F3uBCcK5iL4j+JUIPK2A3NFcWBTR0s5BRpWLiWMkQp++YlL0
3YSuPyxsBjsB4jHfs7DL/hPaybKPfY4wQebYb1/S4CEP2iu+EQ/1kfIslAfWGckbcXIFKKfOG9lP
g7ON+bsZloPp7vWYR4aPC19oBg5OFvtDLmv4+7+N7LVXyMRHMRVt2tEDfPhF5k3QJz7MANY45/A7
JnRUxtLuGihOtqOZSkn6aU/58eu/diVpObLjnGsQhR/x7gudXGLxQAhs9PIhuM7PsDMSddisqkhO
LJbRNQIR2J+FGD1mPSYKpOMNjBfvuuLI+2sAomxTWvmds4oTxlVKjexYND9nypUcndEFNZ3OdPky
on3oFc0A2WrppQiIM/qCs/h9UsM1JJyEIyf/EvT2eAVr495X1i1dLsXL7Fg1aTV68YIawGYYKFvE
2nQs7uvSE28zpX7FPnsUPFZIQu2XUo6gk+be/gTKzKAFKAUThJdexVP5xGDlze4uzuL6p793I8GJ
OJt6B3IsHbEz8N10G8J1lWri3goa/friiHH/sVVxXuOOv+mMatGaCajpcptySxzc+tlV0GgoXCbh
nwsFeXr6WJlrj4apmat1N7naNKd0XjVwcIXCF8UHJzt2p/p9EeBeSN7qJJtD3GC+8CGfwTn660Sx
YraeGov48gLelPMpiC3kE4OXfKG/Y16/g+Up2Mxt34ADs/wR3Tkh2tEVxVwXapxRb3r/jkk9GGS9
vWp/DST/S27cdoCT0BqW2S3nJ2uNccUoVBdIH0HBrDcxT5HQ+rMjZT97uQvE7Uo79VSBCXghm74y
l/IAMhO3ZUEYWS/bKEBvsJl+kjUDnOGIRiGXkHi4l74An8ew/ruB32tZdmoT4A1Xa9eQQRNDMwpm
St3nnJzAIGqRZDCbOY/Ht4BSBPXE+f7S5zhkLV1OYjBH7aobD3wEj4o7ZplR09Ibb/lYbEV0j8Xm
q0RZ3ad4GMmU2qwdX6VS/q6jBQngUmI48HXGCPVd12jryQ3nw9bUWUxnmNTTZO1APq48MzlEWla+
AbhB5U1SZOuwaK/5wKJDTJ8JDsQHWGiCw1X0yv8TiBtjwOPJLYfO7NWWn/KZD72aez328t/QEfgQ
KWxk1H99odiXhmEgBsuwxHx0/t1gh99uVvjkWuYdB7w9yjxM0SNZw5qpG0BBuHNIskLtBW6vKU0n
eM6HCborNjMJwKICu9foqkRB3x7zRXmyIaDmNA7/S0Av1LtLL0QtM80dqlzBmK52fVVGjnWJD4QX
TG2lX3wntaEVbGr2uTNPamuE81Ne7XM+DAokx54G/aS/vIqrxWROcUf/eqAkDXVPH18jhnVA33PM
/dgcJUwjMVZ1MLgxF47W5pfJO4cVzomplqHP98g2uf74fm1aG1vFU5qxEUtWPSfQahuvgAWJk7WI
bACUVr4mOcvseswozaGe26lNyP9v2icfK4HLNUSN0emmMC8LvvOnSU1qfF2GV87KlK+Bib72xnqs
nNkFxoRKaNvWLSsCb8S8SyU+MY43SbX+6AzYI1GnfomA35GXQ1uVxLEyPI0vYc/snGzGQKNQapYV
9220oG1Ma80GGazzN8ZDTlt39B2G/FL9caCRWmpMyD9KoZd2uDn4uAiUQM9Lx3mVkEfXpOoFNqno
VxqRjTsK8zZH7kBQii9vk6k4fn5oclkMsbqCoTBSVgaWITxJiprysSCUaDlCTneBw4M+mF78fuch
E5dgf5H9yRNEzCrgMo+Pg5MYs/hrc2Rmta2NkLd+s7jlP/7zop24QOjISUIZu8s77Iy+oK54TbeQ
nbBwsb19Vb8lt9vbJulVLci3rWWLPKfAlZByli3eM9F816EPndYGPuNK/tfgNkZonwf0rS5sKVtl
zz3D0TvqFN7FgeW2wLoL6d4QAHnHrRYy73aDJdEgCDchvgbMf87B72/uXIpB7TJUvoQPvYbUArM8
xe+fQ0sG4U+Z4U79ckMFYncpjKf51l8xR5kN6eJXDxAGVyXq+nVTD/7HSKqRUsHANzgMSFKippwW
+NhDRslsOtGGAMkrAlwYBWjeN5IeEtcHeseTBUtKT4Y3Kr3HDqdIB9vCvIqfVFVso4MeqjWicEXs
o+DOagOxqdLi+n+5mNSnt56LE+1QmaOqUCVMajmPm4x/UH6nveI7CKvR0doCPcDhfef9Nqp7Z1x8
S2ZIN497Mv+lqVQwwka+jusdi1VncGdbycBr3/TVcIIgEUrv3a27GArigsfY9n7mehgKLUwD/d01
KP9EWvarvCZqwaDhfMujQR0tIzigSgbPclRwtrlwwX01WPmZoMYyImE7xw6qLXU2HpGDlmOkb6ns
n7ctHO0fC7anGBM2E21KGmbfy2OL+Gsdmjj9R+fHi8Fxb+qIjxTA+M5QJqIuLdi9evwzELUj3AqK
cqhAHxSFQXZmIhckutfPnTQNgeQHjJQ45YxxzDyAqhQsmkiciz3Yl7ob3GxuAHBKXxKMK7oJbF2P
3PiJOR1uY9TNFOKCo5Sh9fWj+URhtNzWyLL030HtGb8wSlmitBQJHYgUOaAcdPBCz3RnDXJ/0R+3
u7gSh5reCjV3TEgMFdAxDj2svTl/+jLPkEP6owrfPUgR0vDelk+xTJWxsm8bI70wvZP0+38PHKpX
vuLsyXeY34Zbv+wIQDp6QDClS9XfgBaO8EQIT1zcvW+ruCMYruD0BL/L0ti1nioyBhPyf3kMSleZ
g1shXThZTZZeTddiWtdoJ9QlAQUxZH95Enk25lvoHS90R48ZNSOsG+ajVJiqbTQSVWrUJA2ia4cC
5SVmVxt9aNVcza3NxLejIB+EB+/3d+W/35NaeDlz6pWxrY35kDUccKeNbY7ye5Iy4CyGZ76LlpKU
lVid7reKC0Kp1IJUinkU7fervlT78LvHratLHtRvIrBcgSSnka7iZcrfo2IlNWLr7DPM0aDgY1MS
ihM0Z40Fjcnjy3bMD9U7Fs+X3wvgkpXwWAtgg2bbE7albrOIjLqkTlHtP6jUFFHm4AJ+z+bOHAww
sEnTi6ikYv+IkEbXYukAhPxKRGFsC2eygbMf2hM/iahB6/KEeHOSP2Wvguyj7LUBqn6zmCjKDh0X
HdRbTWHTZFQjCf2ElleTcfff1z5xcdQzLz9T7Vh6PRwzcsKLxTFqx1vZ4Vi2gFbugZMcK+exDVD8
YjFa4QTQuokyelWXIJ76CbplNMO1rAoDhN2RM/+JAlQYM1cOZGCG0dmVzjsBu8oHPGv+KxCHsmWb
7FjesEySwzJ+WrBcRvMyMaufzrtQujhu+JLytjTTqa/t4a6RU+mbahUgCo3Afjc1Pudjx38H+t/Q
npkpSWizZgyQx5jOM1VSXhrqqdWFRIK9B8bOLIj9IpIsXMkcDVUbsW+UMGlAX03nDcu1qBSmSxUK
gEaokFyh5HBGzVW4QWZjEJqDeztMQSKScxPDVZO6wnDLL3EyWf5zTV9/y+MT5rhv03HF46XUgelI
G3t2j9IpHzoB8EQ0e77TB3YT5beBD1PAXpC1V6USYiUGRZhl7s79oFWPYtpwNz1rvj1SFA0k7XiQ
xbp1xOOBxPOS1X0vdBndNJbRX8yHeemyOCLPSPe9QOjdgUx5ovebxEExbY6rfHtubyVse7DcVODI
acos51U5sf/1dEl3CNYl9P0x1eQTedztd/WRKCNJ88CHSgppP9m+98N5AjTgwdQlJz/5DpgaAdjx
VP5N8H38eOWE0UVBTS+csDVnHH6dejV3kDp7TskQehYAUH0GMP4Oph6YAoTFxoZPfyor0DorNoTO
nsNGqZZV5cDEZtEmCxUcxqElhQGbuE2hcLG2fvB0ri78EIVdWVYVU+1ErU0HWJ++nY+/+05xF84B
sx1jlfeaFfyawlJLFbn2oIAQLw0xxpn5qDcM2QNko3tU8DLd7J+7UzrCeGmFNaWXD94vDSJj/2t3
vp3bqqnMu2MPAht4c5Xogk3TYz8fb/QtpMlKpRU36G/z2+RfuP7GFEwTaxnyTWY2lZHScfotb5zr
lLv4qO9qOnX5y0uX59sq1rtTieNhbRZTa2kqqXhoRGhb/9SbIcatTUAopUJVh7B6kq6xY+znppOH
viTANLyDENJejUkcau5BbECf4vxyWN5czwvxSWysziozReWMz5yuCop+VkCdGNEO5Uex0cGOq04c
oek386OkS7L7Qh7LCSJhYiS3bxmtzCuEeFuDNZKAJbQvNs0nVDkyBxNT3ljSX4CUmu53kU31Od8/
AP7c2ZJQgausx+7a84fsAIOjUFohA5xxD6ttC0/7XkAffmhKqledIrVrTC4o9gZKTTiCayDweevg
EpPqrz9ILKrNJE3bgv29WdVx3iMZR/HiJx9YIZb++ma/wzf0og74ttadJw/FwFLKMx1DIPozIDhh
+XAFhPYc/avrHbauR7Z6dpu+but+hcyEA6tvTmHwLUG9zeBtMVt3hjgWZ0vu0wnYJWA0FWGz3yNc
fSbp9Lj87tY585vQIlArumSu9AMs2r3ghCeKYyDu+vSjmEKGW21bPLoS79fi93d6Uim24hdDQ9LQ
7YNUlQBLHzKPgfRLQimBm483CFL6FElS06LS8fhy2QxAiS/SI2RCYAWEK8sNDvWc7HbAc2aNrXbk
TJNHF7IqcSv+/jBl6PuWQELL/4j8IuBmBwKrkq30vTRk+uPx3GTRWaFq5MC8xYf4d31qPVJKeut/
7F+Fm+Rf9xnnRBcSxtplxYH7Evqy3REq5G2le1RTcuCso6orizoVTeh+/U7casjeYFye6Flts1B2
3ItbuxnZHAUUwsjuE+Bu+HzTO86ql0sDxwXCxwTckaOpArhEPrrbqgZfos6t0aPGU75cZ42+zw0W
V3nV+l0SBhL6bGxJsEA9ZfO/UEkCbSGcbzENuEblbR0OjPEgUZqpnT4Wz3vESK1XhLn0Oaob3gWH
KkD4VMVd/86c0nlqbVxbQGO3Ngwe71g4F4Ko3RUNFuV2U1yod5YDNl2NgC67JFt1dcFl+oHEmq9p
yJvmDhVrcmbZMYSEJ9HNpcGyndxWdIRB8YvnPiwxHzUK2ysTuRbPezohQGYvsAfk2/WidhG6GG99
mkT8HvAYjUXilQBLb7efuP8xbbb3k50Jr9egMZu1RoD8MHNlz6s2fOTZczYDgCLKmaMp56EcT0sX
87Eno+5tYn+PDtZFjJ8WpaOo1zzv1dWzpgtX9aOvbzWnN13OG3QK+bQPyf3NI3xX1wE/2/8W7CnK
1Mc9xVt+bSns+zCR1Ha1hDr+pYizVwZcl1aloGv0tsRkdPsh8Egde7DAR4wXKrtihzJhO9Bq7b/h
s5X1UHTlhxKit08t0fayNcoAEPeVRbZaNg64VJS7DsvLZJBKCo+IBctQb3UKeiM8V1QLuwgcRUO1
EDeAkDH2JdegYAsfij2BGart+qwCaqLnfRlY4im7N4oroCKwAln13TaG6Ut9SEXAAZhoI+NmBq/T
DZqZbbDx0AY8AAhPusroMyJpGI12WPA/SrSvzn2DZWWMdxY0RWyEMyAqhd7Ow1L9paaAY5a8d/IZ
OBEzn8xX4E/TZQleGGkQc0K+UvVC/ZP3rW5jT3ruEnGQdxWIFyRySdycefOxiQszeRv0iFBjMLtD
8kixlFiD7wny77cQ4CxwAu2e9N40qm5ygVgE5K9Jvu1gP6S9nS4nMHZUSBGMMrRLZJK+B2JySGZf
1305b2SSyoVeHr+8lEoCijJ4vjIlUAqQqmzoaasvKBpVzTsZqmBjWzRc+nCWXjyQdU7xsyXUOitZ
niIh7OhIu5O8OTTtMJKph99+8gXJhqsQ6nOkD9F8vBv819iiiTGOLC2hH0pRGMfNibDb3raVA+zj
NIiY0eYR+2fXB4rhSggavQhoC0B/taAx6kzqOL721cdDN7s6yXj1DJeeZ/rSjw0CNPcfDMhB6qvr
TSAa/2ObLKxEMlm7inEsqZ9tZ3Fy7zBVY+xCRoMk/hyHdkBRhLaDTB9j9y2HCOGaNVsiP3Wi8sQj
EfMYS/5VJMdgj9UqI0BOljmv9t2nCZoHloEftJ5B4OkbLoa4UvSSdIpEc2bX39jIApQRspXASn4l
GKQIVNZBabpheUSnikllKrUrunk7OOQGqGjOUgmWJaC12qtSaSobM8B37/MAqj2N1UAHCjci1DFw
5MJ1wsack8schivULvn5LSlmOXw87BhfCm+q3QoSFTaJMfM1L09M2FArVSX4mzQcdJgQEGwqSMfS
opteno0+aLrgx3+rLSAS80mDlcFeDVI0L6eBDbLiNOlGHY82OS8S276EZKIawHMfhPlMgxioK8q3
vXEw6S0aoB6Z5qo48JV5l+oS05jlu7+NfOWVBz1o/giUWMaeJZL+ZfpNuUJqwZRb1539tnwRCepZ
aez30qeIXxAxzU5Od3QvZHCFVZEkPyl/zJaMMMbtZPRANfei0Y4U95H1ts1dsrWQUnTBSkx9d5De
lqyUDmmvPCF8rVuyPxho5NrDVd0YiK6tCZsDnnAA/76rTz36e8aDWwmHPDMuO/3Dw415jd8kKHY+
J5JP3bh38vd7fXYls83TTrstCm8M1x62fyBkNamkTJK/fQnAf3zkxiXxahCMtCDmYbZFqK5mCrrY
XhyW11m8XQPmhvC5ghyKqIKz3Bz+cclFKHuXF8ziyvdhcTt7YLw4HXSykSgqQEw+1GUa8F8wQHWe
l5PUNZKg52HPsDHWAGkkI4a2atZbqo0Dpg6DaIyUR9GD0T13PaomCRlx/3ric4GDfUJpg6o5qOXQ
cS/fshd/nfKfyZkcXpfC6RFCrso3y3wWW6pZjPxL8vqxBHVIkjLdgqpbiA6p8G5dueOe7XsAP5bx
xRdnsF5KWnaRW0zctDYFrGZLll1CbEODk+ufJEESRZdsxFNdmPABVv/tUWzcf5gLIKK9VKYq12gv
wYxo7TRhLS7b7QUbAyeLWdiQulKTQp5nR28tGUpqYdXcvps+a20d09JpsiHROQSPT+xSKJ0ejE2E
zbrOPIfJF5mDj0hZuGsfUoo+rulwnGOqaFd5vO0HtCFNiK/1PDeYl3PHH9GIK+QihE0UeSxXyxSK
00t30cO1TZlAcO02zH1CQMTwE1F1n5Gr3wFytP85XS7p/fJw6VpiPuoOiSl7p/9+rySth/W9GwWo
+gOfRllR6RnsSSYuT9TE3GTsZpacx/ZeaMWT2tN0AZZQTCphSb+jPMH4YiysJg7OyfoeuoC+rD7P
JugJwX+WHW4yt9vdu8JUxKzYaGro4i8MLh6E1BHruW1Q6Iwn7qO0EhXjdJXHN5RJQO/2O/tx0teE
Xx1vDxxhHTBk3FDGo0yr0QCn6kIR/WzjuZ8jiTfFvWgR8r4gh2MUmtq2tSaBGHxd+yI9uS1i6ysg
PZ3IOZofQNOXpH63mW+LBIdRkzKobtzTuBkAnoz2tQQfPNq0o58WWTiFlUqWyjX8OCoqxQzCQQvx
pTgiQQuWMMCHHDcNvAdBXbJ+dP7XVnSRAlgv3jFuZG3xOuXzwmbdHwFyeqUhFC99X5pmg+UNqe2A
T+oYQHNzUYWkQrFEtb+tmwlTtLzSJceAR6o86DbL2Xy90C+pDLEXugvDPLhYgYlKobRKSRhhkJ8I
DaGhzB5pP67HZp0cggNnS0nnU18LiUMZ6ISySVYju5z/By6LLT/FShu9kl5rG12ChJQgAUaAIB2Z
H6mZf29XxlFwlidFmuCdpVjRmJoaukHtek3ynJwSjqzDXdNpv5f/3hl0GVnKvzBG1bli6FDC34tX
+Y2jufAgSjPvLFVMgm0hy5gB4bz/8FhsAI+2iTk5+u/7uMlfk1ZP6/UEBpvnjUo93O4rEQqOLB5c
sx8TWn35KsGP9/8WHN55dN+XaINOHZijdrRtoS3rQ2SDcVmGrWPWthAPwWKXN8IxEfNxuLhdq9RR
aRLVkLJtzKkpk2ylAbAgRBaotKI4Pb2LOw3akOb4HIfW9rSkd/hFkbY8qO81a4DyJ3VlR9iPF6ZT
p7hqTMK16DaRLfHCP3QKH5PK9Ub/0ShB1hr/sYvSaxSJ5ZVuJMXjRZj/OY6pRzFoXvcyyo/ae4Gr
ACN6Hqb+IHQjZjwWpydm6KyGYAec/wmemuPXdtIcPDNIjowgPrL/nXW01eumjEyPOovSNqBKGTX9
Lh3b17cFhFEZDLhmUWt6B9UqtzX7668QDFr+GDQCLQt9eQo5OlxbCrKALqYmL/OMg3q682mlnuuJ
uiOSnVn9sHvgCCsq5mMHpn7VkE/xzAkhk8vWdTVxfqLgTLj6sFzboi/xPXrDqv0DAt+QNKsvYDP1
ZfJzGmBJsT2V8Y9CGO43EWSsc0LJ+FX/KvN21ucUl+fsw9XZ0m5H+hddH/mwJe7f/KVtYhVX00PZ
buZrXG0CZEd3FKoiEzeNsQUSUg1A77i+m27F+VwH/QqUpqkttSNn3wN8Pcu9N4h7c3Wtu8wiDi6v
D6uGyl7TFSr2c5Idxp/UnUFvtcklurmENVq3vvsnm4t24kInJu1zxrV8O+FKut9Ls3Q0gVM7MCn0
VtRuBcAO22vDfSyB9HGNDLchAKO3Xa2ZbghH0A5VHLq5Eenkm6Y5DLcwD6H+RAs+JAd67//kOZd1
adZZcFWkOw++eoCjJJ1Vgr/MJHYQ6RLEc6KjNYmhbEITIAXwtwBaOMsy4X6EHuCnCdo7sGWbZqeo
fT6NPKhaopwA1st16RY6vM7+ZqGOkIIYoKHLTSI7tTJ/g420vuWbXifMy/7DJnTdGmLmNcQiih2t
kmekTZZMJ0qXwc/6leBhWr7NSdEhTo/itWRWUiWthv0abSmFR+3UCcmBPJnzlj0Eeu0+fI3xPWtm
CxNHtoR3zaN+9oSsgozN49gfH8SsUFzMkb30Jt/yhX7j9JuMYBJHpyuh8F2JrE5zQDsYNRylYnnv
5owbaN00/m+FApiDdxRXMHKLA/N5ySLE54mAfzp0v4RvoYCT/GkH+Fv4qJLiERH5RBlnHDyeYW1V
uG1Zepa1TBMuE/ukxtqZIPmyLLFs6Wsu4jR4SWvfbR/R4wQ8rD5ZOcSXL3GJ0BlYJJUB3AAl8LJt
bTtDbdSC3lyF63Yo4Z4IS/38gpUBj+2RAsO9AFGYq/Ksbb9/qjIRvPfer/ZdXLW0Zs/ZTwxmflkH
tM+xk+ILfk5FSX7kF4Hia1ObvSgMdF774zBSsK97BoaYvxMnJub2LxSG+c40Ne9KNOX49HCjnBwZ
KnW+kIKfnFWQVf0PjqrAN75iRaRO/X7YOipcRdKY0ObOyZ+t5ZkU3kRoSv6oX/mV6wok7dqVWt+M
XTbaun1clVBuiWBI2rGCRVB8xH1W/eRLfBT+tmm8wYdmrkxEhHv0K3IVD/oFvbB15vvtzlvUEdEr
63tR0Owd/rM40BNzJJ83BXKlUkFJVXr/x45kYudRfhuQMZ7hRuNxLaKmWOv8rn9dbYx3uMiRTUjk
GnHXK9z4h4CNJ8jLrCbCe3WHAsIpNbCJ6pN+ErmaD4EKa3349krSj+RiTVmybyOxvykgQN/PwexS
5Ou+hly/1dE4B9P9s/ugEK1fzxZ9KYWatdwlyb1I0NCmR6uJO7IJQ++Ldn/iCmpqbAUTNMU6e6JI
v6sesYqu0Up2Q5NMabme990ojoB6nqQlXgX6s/hHvzYNPxYTXE/OJV2ES/PBYpFdCyyaXQs/TcIJ
Y2c10fXl0uXdsow0sHLxoVtBgla82UQp6qqPClms2NaU4/R9jG2gRHGTYPCbcZ7C37hz9VAi15tg
75bbswesZzaSh3lpKqeOFbsYeamBix7zOh+zjY3VV61dUegz83AI9X3T4BjEU7cWUPnniYT5qI1a
itaSCnyoUJcZQ1m1Yl5oCqWIY66Atpl9EWeEkDzpwz+hMxCZ6BkiCGb4I24+KEID4jNoV9Z3NNJh
41SPVAuTZZcpn+/0DGas8jPH7MquWF1N5ngEMas6r297lfHjeh0hwZ4UUG2R4MRHX24QKvHHtfTw
gQYZRTPWDUgdanxb/FAf9VAjDHTRPRp3Yt2wvmwLQwFCFd2yVFbquuUrWmifId3Sfy8RhrPdW6Q9
JpcngjfjanmGgloLdXTfhFwfYiAIQT8R9fYHcLB+Y0U7W/Mi9MdmVjAVn7Yvk2RcQYj+sWWvpDMi
w9Cgjah+usR8OLU7YNnLgneFfodk1Ew1gnSAzSTyH3q0YDIneqLiFyFF5RnhQqb+el2Rq1oKpSj9
I2dktYe8QiiKjQRnqWclHcDucUTUsFew81vqHi6fjY7d0xDY/l2yoag7TMfLZ7LFW/CZMe4OGYda
/yIf5DqaMyTAIEo7eG3gGt7ZLCFclZiHMCQC23SJ7gJz6YUexaelvOST/2C5L2XHtxK3L0fADjo3
jIITkRAbQtobZeP1mIlmGq5yVPkWTMxzJRbasGiY7SAy0QgLlCTGfxxOKjRnOkr9Ugn2HzTlHLEa
LquW64n5kij8NK46Ib/Y+IF71B4HLfrIOIEPn79C7QV3LQ6VWo5DxSssaEGnK0fby3KfIxlHGPAv
Ejt2ho+RWYqhRfseGZduqanPYYuymJwrfuwmSgX2Qz4s8t5A++jQCjCn4SOpVk9KvDkTcvSsIs/o
QZp7mTI0T74JMLLEvt6oqMjigwPqmCdCjlzibBVMdxHxDZ30aj7ZsbWly58qrQK/XMww0+hKMTW9
VUFK1uNOkKEhemrK+6Rz8tIva7+9xxGN1LabwfBWbtAItvJ8AHRsha8pV+cBgocWQDQIHKUtjMzj
ww4010b4k4a1JKBMhce3V0nekePn2VR5VWW1dX+SycSPYg11sUz9PGRB0jWGN72Denc+CBbX9UpV
3dF7x2eOJjXz5iaG2VZJnFL6A8w5BhydKvscosrdIWCvcfCXwsSBe+v/h/vuTldsftHWpMLhDjuD
9dwXPXPQRB8J+EAt8O1cKsoEWiwTNrVWjK18QCDvAp7bhZyO/jaiB4FK/77kasRRsfvQIfUHPbsX
CJ3J0/9gzt4AavycnxkPkOL/2IcTQ27ep4WqeVazMbJO23GbIMj6moaMHsA7CVxsSAspJdmVxGm0
micAgu0b/9fFKjMjVmRTKPOMwF+xO5dazyBCkj+n1aSPPrfFtgqelE2x+RNriL77oy09G2OGF/e0
ZOELmJP+aTrE9axBI3PHLUztE8fuyKGkNANNXnBSQq2XtLWckbBFDDj3dVCV8PVXp/Sl7mmtMhfB
HF7G6ivTr8nD2QIW9OZpUbhHyCcTDOyNp2ZIps65E+68MwVlNdl4pjxxD9dgdGVlQQyrCdwWJfq5
5V65YcVwxmPjBPx6/oz2SBImwvvgylr5YubNcekLxKj6D9VpsiQ7/jiqIxKurJtBXD7XtfVA7Nqx
0Tld80gFsjw0Ac41DuHpCT3HXFL+swGcZWGXDQgw6WNHXCQQGZQJV2jZC5RFqc/VUrPMMZwD3rOa
h9P2kYAp8pR0cYKknYIDTIbfMo/l4gRZw/vFprjcUCOcVO5e4AHThUggKMIla70IP7b87BniDOYd
I8mkEG7ofoa7ig9QkrpEIqTBIkwGqj8mf8SyXE3Awr8+OZLDywdd6rprWTt6lLfLtozCxy0CppJS
s48vBAgtfsWshK6wkzNlrLHu3Lt26Oe+4IJMn7hrba8/pTRdX+VDVd2aebm895ags/LBp/Fp8DWF
OFaKHf64+IAXSjp08zwTLMNEA9bH9QOfrzk7car4kUc/ahKfxQtBqkb6pZ8vBkO/6lwLWtig2wtq
Ed/3psd615mmnWvmBBs18OlIMjt7lrGa6XiPaK7rYlAzNL+iPTQ29L+kjZqtcMZVGF8ENiAFS91L
B/OXbnt3PbXi4iw5744L7lWiZbeQFRUg32vTnLwvavPm1IySNBluNx3bATytwSsxe8ZJZkK5a3AB
fuiQlE+5p41cjRStNtWEkftLiUR9p00IAkIH8CIQm+1wwCPL5w3RMdnRSRLhkPUDhLo8X5wUCj9V
bJdb4mfvckNOu6mE15IdU5bRAQBRsSyPudKibdDGCFA2utS8BtT1Ybw9L5lP7dTUU9iwcY5zx5OK
zSk4nDcYFbfgfSt4ZJasQ3KXm5QnYdR0bMZRbh6QAq7GkH8CUwk3xAlfhDRVoE6qFdLJ1J4HhKmy
47YqrTV/GafZsmrYk76SbvT0r69RGvWlJg7lm5QGRV6wzqh/eOl3RZsO/HuymAi9nY1W0IzgysS6
x1zl18ghfZpzy8UH8D1PepBKQHjPLFUTvvVUuyqLXQQfjgiLE2zYKHXA6IzIZZKXv+f3gA3SS/jo
wxH7g9VVjmJ9k5w0ksJme3vRu/MePQLgExH8aN5ELRTr0rtVqJskLUCmWE9r/hZUY6vVN/CHsTLL
GvlBH+V+OLDmwUczuL777l6IRuGsgFaqsWjet0Lj9eOpjOpWDeavLQAEdDH+Dy97D8XMlKSeCE8I
OHBD4QFQr1HS/KwFSW2JpWhdyNpczblWH3b7vPmE2+WNKSe0/EghySWg/P8RCZ1VcqrlEbFlw+Cp
8y08+H5aKwprtZzqLzQ2c2Cmt380cFU/XV5SgqCoi2LO8thXWikfMPgjEb7Pg3NHkVC7y9PS40Q2
Znh2zA7xUCysTgfOPKofCD64xMJvTB4dDXV7ngAJeVw9UIc4lnSzsVupzdaY8M+i1SO9Cc/vsf0H
wJPkI22nODTLwUTpo2y6Y5kiH7/bGrIBjVr++Kn97C+f9pz1ZdESpeRdutOC4Ak5YH00MunLy2zR
x43OD/WUxN9NbGxVQZKS1HcdCxt5tnt8kDhVcl22tPcqykcBPwhwRN/ZkkRFSWB5K+wEXzeG79bC
dnC8aemx92fFNny93lX8nQbC4eBLQU9mq3J244iBhSqWZWxPCgDFMaJjdMpR7Gm9/G4SRJolbQFL
Wcb3nkSiILRwGgzMt0VQP/fE17muIvpbLsMXBenpeuiBCo8s1HiFt7hRBOqOJZ8+m1LINTYRazMT
Lr8EQOyEMeygDjGDwIeBPpBDLVaedFVSbNH+Q6Cr2JU/9qpNer3f1wPnLvSTpU1qpmHeWCHHLAqS
ErdTCmMIdPTCvWbynu0TXfAZnWeb+bH6c5liEMxzG5avcleHxlgC7WLt6rZKoC1qbx6bzFJ0rXbd
cnkeOuhycJHkTMddVCqFJrK1O7fzwiyxWY03IF/ICsZL3vIw2jXO7M5TAUyyXnRc0Lqnc2Ff3mcg
uKpfX3Lh90kYqk3rY3GtK36KVgYuE0QzQ4LR1BtLq2p3eUUHuiNVKgos+1JuwetfyMLRP6YrP0jU
L2Y7Jr0EN9PMnjbm1fMYdqImjUQlPz2uC++XQ/Rpn4zM69s8c7rQSmkkQc7HQqHDGtoKdEYSJg1b
6nCwE/SmfVz/bkYI2PosjZngbZS625kGuQccFtoBk+EH+Xs/U0Yy/vmEhSgKj3nojYKbl7ADGV/f
tetlYq9GiUmewC9EhNA1UE9NzaT65rjzg7+wCWlLU2Z3YoHLcBGoZDOQ4jBtM3LzsNej3u9UvJbH
amegy7QhJ2EgkKYsNXVofxdLJSts6lDTfCZ0Vvs52hRxKj3u7brTX6mj5/rN3g9wMqdsG5q3CSDW
yAD4+d3VGXqMaNnve37gduROK1zWXWbPJscT2KR0FaQ/GMCMBpbs8qELQfbgRTym7Iogz9lfWGbQ
nhu79WPu89Dx/qOrwiSSQIObyR8YPId6tWnHD+srjy8Fl4XWy/AfBJaM8OtGP7WpiPMzJTgfTDxF
CAdX71eEZ2obSie+c8tNzUJsgjj0E1/jpLb6dtU8sGxK03FQDfWVnNrqUKZso4lgLKMob0d1rzvy
ZNHeccou7B8M0rWZeOT2dbnvUdPCvCPd2vhs61o0gEQRSjUFutgOkMPmJ9A70wtjZlToY9bIUFOo
g7bb5lak5Cg0RC11w8vOiQyzt1PGxbQKqZBq/ceehgHieYfQj4zyGzYPqSObnyvWH76o9ypz367q
nQOe9fuyfsEyMoAx9zymx2lW4FYBSKakYkEzuqH98n9ceRoGJlsXDDdJ3SGqaU+A0wtziDmd6YWy
XrkMglEVSE3H/98ChWj5za2EpHmC9v5AFBeYhjscxEGlJP0iTDB62lt/H4E+YrC6F+mOXxfdnL5r
jb6pTeLTSWAm66zxydG5Hsbd81Rnaj2fyvMWNL2Aqt48RzwNpbyt6F0tMGiAO072FoTvm9J6QDuP
2XR9ellpwyW2yflkkp7uhKxLcKJEfTSAHifw3ALWdUw27zxv3Je9ZismDr5335V29PW9tqrnNSme
P7RcBvM0L8KAMBiJjicgRR1D4z2/otHCElZxqlAKEoPG3VVvUbf3o/NNZcNMPR0Z0JuYHeIQgMyI
rmzz6tasqmlYKgvXp5i2GN6QAeasS+hiZIzLlb/iC7Yr41OczXhEk7hgTjQHz+eowwcSW4X6rcAg
Ui+uEn1JYxnGaGai4FZT+IxvK0c1dyrmLATR4rWI3b/FLo03f5Eej83fhDsSOHhkh1ZsK9/lcc1o
L5rgY6ohJ/8bi1zjNwStpQiUddcUl11imhicAUYm9MHpLBmeEQYAzQpfVh12pd8qG5GbT2YPpfxW
zPATDQ6e5MysJBE8av4wEV2z/majctPig7ImH58QpqGkPr0xQuZlpoiZgMve3ZsMpzjUObycJcUf
MOOPFf9Fflpy9MmE3t6mh7QDpE/82o4Y/sCKdw1tFdpaCJbsoyyFMzwEBW0wFKRhMLxNggdU7AcU
fZfxN4P3NLKG67r+56Akovpd0F7Xv0M9/1pQ2mM9+2xlQfPGwLboBO2UnzDFXNBFvi3lRdYIka10
BOo9losAxNDlBqGt2xZeEK4J5eC3I9Nx/hGjGaukk4DiSgglNFMv1QtRWe2yslcMeoqa+GaI+JvW
AtNk7mZxgRJS/w4DE09SCRoaMm1XRneCMOwDPNDPmgO/XQwws5ufnkKk1dCGi3tzGtDqAFlp3yS2
SaTr79nADOdmTYx/KdbwhA6MjPi/h2FyevzmMkEOD/5n61jf0tgwVxwIIqUFm2WUrO//HhPRRweT
ejtBI2PwTN6gyaeQgHOVrtmhwDoP7LHQefnc/wRPUwq7JYOTxnpKYtaVNr7MPCIg8ynQVlsDAd3v
22ejyr6fXFX7EmhFk+KR6uCI7/2eqfz3lXENV0030eQCOZ9uDjhcel3W3IdpA8++JRUMlfCkSHl3
jmKKBHfrKot07e4BPFGh6wfibrWjk9unXg9ymT+GUy+JS67f98cXRX16XBgZacGmzYwf6cRmhU5P
p/qfdYVZ1tNOhzrJ8+kRhYiSwDA5W/rkEYb9BnqPsAd+eMgnUY5Kr15Lvm0z0lPbxvbPDs5wpQSl
uCmQUFAxbN34C8H72uGcOkFP5uqYaNPA6awqVjVYsST/GSUoLdUhOM5socs9RU3AUq6VE2WOawKe
oSSBSonhvNduL4+quhZJZLwbGv/IauXISI2/lv10POVGXVYY9Yt1VfK9obl5IgeYGWo2ls97cOQB
qN3oCgfazIWpkhXIY4nyWzx4njaZ0Il3Ct3sTi6PXlv9uTdGcxnIaRae/xOAme2qbkCbvJGFQPQ6
cqGoBsMff7mv7QEQPgwaABHVJ33btLXNOfq0fxGtQnYA0r0xFZ7iWFVd6GbxvQg+GBglDNl1dFIm
7tfaHoSITAfWbTN9ZcFyELFW0JTUdpFCwp16k5jsIhLv1n7x4jOb2MklbOJh5XShnUV+CQ6WXZho
pGTS7UYqPh2XiQQwqDmovEZ7YPRGpLhvOmYFBNZCbjZDxaiMlxklKrHLZD8jhgqnAp4eV4sSEMNN
E7H+66p2WlZ2fRRN0gca/FVHPpUBaGWz8ZCAoiQqUnIkNT/InYh1xFhVlQBZcAaxc3YqGsgqxx1V
yH37wTdwltbiQ2qO6uulj+y6q+xqExNrTbl8ltFREEGuEPyC4a4L87DGbaEh+ZSFh8zyHsMmMZeK
JYFZ30Z867RdHCOknswjB5z8/l6HSxXjmZo88wR8DswizBxfMZ9i5oPtxXeB48avLYEYJXxUFZf0
vAmDuxHtfYx9hjN3gVKEYYGg/6/xrfuE83IzK4MCOw80M08EwXw7g4J3NXvWWBg7IuPhehMf2OsU
U9h85OnW0JjxaIoSzFO/dyCTS0Gn0fFtLb8PyESFI8PBrvGJjZtilye73PfyguP39Y9MxcsVbwSL
txLQRHMr2w/5HHBjgpW2XNhOt4sv8Uy4Rsaw/G2i/6z+j7gi/rx+Xqr9kD5tNa9OxwB3yU3kQNBd
aZFOgZiFktzDU/8YkiHOjF+NFN5elmZ+8VG9xneEh4otBH/KKTIa+ru/FdJJyly+vLeFSh0w5b4t
C8dfARvQIYPhk2LIQNqnyi8dXaUFd6moGyVDwVbIVSVsxRNE4ScyuAnh/F9LCNe3Ztn/KAzmtGDB
x7DZUwNxCZUvZkzYc1vJU5fmaCbpelCN5I9gH5wNi1lowuTMc/0vSN90k+/0bMtyaS+jQlU73U9f
5DcByyqClL7SJko21YS3nyKeQYRMj3S3TO7vPyTvxkvuWfRNSJznfSI5js7Olu8xAFDQNXJIaSK3
9B/hnP2aPwNGXwJqB5LAUJYjAKHUEt+vhjlRaiapxg2TfzlYo8QaIX6jU2uK+K6ODolvsnJx8NiI
Lxm4ItPtGZvtjXGHZOkpq4NCskmFhONcDp7kWUXv7/1ab/smye1HGNSQVp2ThOARrBxCZEGrBeVi
MTzpCx+66bMdIcEBaXMFUWrZzswtzpz4RYSBYepNd75FMgO8rwvtthOKIjbE+MLL16NPGIPQEIbh
8iE1t2z6pBiO87qLhtqpQUoVBJAPY7CClPnsKzkwGfNe4KIQU9fPnNKes/mwoELLycVMlVz/8tzq
ih5h20F/K01BAb9fN5Lg4XZFTwUJb5FUdrFwIhyw+QCuN7viYalws+i6/oLWBS6Zd6F7DdK3Y40q
YyiPCMvGr0S2FrBHOoVdSbMS7meoo/1/48Z0FjQPJQtbjKDL7P3OpPou3d6sbxRL5rpeSECEp0eW
bbCj3uEBSbJY9ippS/+8u28qufEHHqbAdgZUR4HNegyNagtA1nYCHlw9a8alF7Ks03NJKqLU1Xfm
Ye4M35GaQtwkYjohjp0sSGqbAhYdcais4+J1T4HneLvMICMc3ecXSQ5tyfKqz51siOUOvmMShEtO
YE5oBmWVnat5D5y/Ns+WmJVDgbFW9mx9Vj1BKMdkBd+n2PN2SGM01N6R9g9DY0p3RLRxlcQx8kBr
DVw/13AGeRC1+exj+P65CeBFDilHVu4PQG3PsqK/s+rTMOKcpXCA0XkSBEFfZFnSMnHWOSwHV6Pu
uQi8KeYf9wgDNYH6Us1P29D3KXDW7WtUsI/Frmk430TaEZr5gVd6xhZeFI3f2gR+DDJ9ulR6RrWw
Q2cRswpDg3Zy8uNyozF5LT2CATrtMkZlEs6yLjSTt/jPu1n1LgppCLi1EsCoA4GLnBFRtGSJfTr7
+Og8baPZ0nikTG7cWTq6vNFwupZbcxlCDqEXH/9Uvr9Vg/xJDPkh7WydRa71VLGV0W1Nes1kkh1n
vtZ/xB1d3WcGdA96tfhtfS5HQXGMkrl0HedUcVdY372HnYkqe9tV+G52A+PNH16v/xs8lF4JFq0i
Y1KHX9mbLSpgYtAnlbzAe4j1wtvOc8yHwkc5Wxr14jJA2cNE0HK6QYCp2RM9ZjnTB9RcHvr76xnw
+E8IG9F6brLCdqAsn3BTQuRrhuLKs4xR6JPGYYCaHcqY1wVnBUAc1EGTpLGqFpuDaVkaIVf2JuIo
VvhhhqAOBUgSFfC0DUMf975ehqG2JbXc1yjDd3Z3xobHX1hQVNv4Fj9jR5b/ztj56meD+v9VOm7g
GPugaEtP8+pDHc7qEjFMJA0ofsQ1uSFj3ItbmY2jBAiQQVvHy9AZFrbZKjEuCKF3In7DGNjnnmKU
l8lSIubxBt0NfcaOYU4/Co6p4YUt7jaqdw9Tq1ca6Hl/hcJv0PV6Kzn+DuPM2lDWObma68Sm0wJZ
S+UjqjaYUVatG5XGoJ914y4FRK2OpG5wcql1Y5EBwIQilU9JNZYhJBln5sFMIcQUW3HkPHQCp0Qi
do6MN4UI/Cshi121ePQLm3gWIrrA4GMfch8b8syVzQQ529KXdEl5nP/cpyEBTnf2ACFbxzWzJftD
KBTCAyjgyVLNK+bbNQadJyv8maQGRuxsN/2a6EKFqB6Ca4dOn41O1F++xZx5D4rZ2atB84sXpRlr
NoWpwkKg/tQFC3MZ+BnsCsZGoPVHAuYyo38mYeT51IfIrzwxdt24kbsTk2SOkgTZ61/YzDEgWhiX
PQkJjPpwoBTfXABmc89VJICWKtppTIYhGGIbRXEETpxQulce6UVQFN7qnINI0XDnIJYhHeS5V8V/
6H87pcgEsStR471S1Hi0FtoEgJIwpk0cSSemaoKXxwTE5WzpAGk0Z0O0k3wzc2DH2lCxkTGa7KMQ
vQnqdTSpGwf+43T8Fconya9RQYpybINSebQa8O/X2GmRkbJYzvl+Nh5TYBnUTEe0iUELrQIogtc7
tURFs6Ke3hBsRjv3NqGkrEuNGehysz3csXqoBixirksc+k1Av/iHKWY0GXh2cr7PQ8Ke9sSZ63Uw
VrIkZYRTA/16VL5axdPHMFdsO7mlAWuBFdxeSwGWVNNhRzON8NHm0jos1Qaj5b74FVk/P3cka+E/
RgPVjAuTcn7ztPQs3R4uy2kdxIk7Gxt9BDB/R9SHDg8ry3C7Bwvm6jo2MVcUHpFSDEXZvy6Pkp96
WzK3DTQX8ZooCGt9ZryX4gx2q94gMhGEjZ4AsDOY00WiCLkir3B7F9YqAUnWsKu849aW+OdkNEdA
af7HQUxMJ6cjEgeJx5FaITaWbZYqpmeE1MVu3aK5zaOF7rcj8w4sgQxkeNzldwRp5k0nSXIxIySb
WP2/sSlZbaITvTgGCHW0mJkLtnf0jBZ7rqotnI2PjEf8m8iV2NdUgdOvUWQM8Mb0eOfbRq75uFPA
y1dLZVywdxJ3e9wpkxM/uMXaSq4CgQjvbghuTqwHvZsskoslfh3/354VRsBTt7Z2BPUupgDxiGtt
tS060eD7geka4aDwT0U0n0UeYH4LuwTLE6jhWwQTh25GOr3ojoKtsBl8FsrFpdGNHc3BKgoHsrVk
oVl8gPHJb1SQ8qQAwJgUHDDWwF166u45ndfYDH28TZt4z/QrebDnYdUslhRjYsbU8mcpDlaLfck6
i3BcuRrMRNq2dARc/EPGO2bmMcFlLkga6ZX3vTbz/mi02iwZxxLOd+5IFKNFNhdzWjBV3bmWQYMX
k0UYIqGkvvrFFqjnY4sy8Nn5s8uH311qSKesSwVPhf2C3L9FG5pdiCEYY+uSMJzAGnVCAKuPCkp/
eRM0inLaMe7Wpz8arZ3POhXwV0uJ5gQ3zHk2L/jkC/moUwPs9nVjegUypkkzGvql2ZAOC41mZMH5
StuwULaP2dmzhvXKOGhiO2o0OE3tEI8HSgejACNE28C82SpImC0XZDInY9ZkcIajuTARCUfsnJAt
NMVstgF4IhrpAkMLgpQ0KVuQ+VX8KJF9Q0gmHhSGwIP0grzlElHXrxNjVHIwTPA5lzfBIwv7a3c2
xiNw+QMmXqlWJ01zziM6RW+a2KjPigzqIfZXo6ZsHic5EFRdsPnxmJrOjLkjWJFc5+2/WDYNbIoy
syyZYFC/0E4ch8FZJ3N/krpqHj+LstXNUD1oKLjGWq2unJngBE/br1A6CIbfN/WGzNd/died3LYo
yUHi2f6PAz8KSk1/EOHD8eshytwdv4r3k37KUAqKUnSLv0byjDC8cNswjNnKe1HmweOnlIpnvHsC
w98uA8yOix+N3NSgB+33/RkVM+ZEwFyba/41JsPLaqbtFKeevsvl1+Z2b/Is0kK5EsdAwC0MjMYd
t1co/NHKOQRvQFJNCgUb2txMFvKAgWAUPhApsUF73ElHwt3/DT7Init3Am5dYcOR2RE+29G5DLdH
EraHBeslh5UXJW3ZB0XuYRvfH5Zg+eE/zAmgLZujPIL9iUqXPeMeu6WGqOlcWf0yVFC+4ABpiQFR
4kC8l6EJ/YX4nC7LtKLN858XFWTVWv3hELsEnrVTnRyVq7l3dw3Od0qMzi2NWagCq2fjQ6mOCYks
PNkvclQmWGsZDxMsFXJHbbi/aNSHNMJvS3m8WMq68T+QGNa5pYinrQ2YD+wrpmthxuCDQyi3tcZx
Q/U5r06sWGAsFUaPwDRO5u9X0eUdP+82pgV8wHZfavBxQ7ExQ3w1jmQkaiZMLd9XpTCbq4XlHS7A
INgN2sbm0YdDyIYnn0GMOYX/nx3czOMBJR3ze5kqDjsfnEPpTUSjKGgETR1ZLxeiHk57+KrMC5G3
nb70RC5g0OgO1oBd/QRS50sASkUE9KBI+RZPtLFC/1eG/4+tZe4+t58eh7wRwNGkTgHisYYKoRDA
XzGfiX24fApg1hWew9VoWH2nguGc2N666DE/au+zsHlWPlPcRR1BbIHG+ddZm+Sl4YIt9IWw3Lz0
ZU91xn2pd3nqVfN3+1PvG4sQs7PbYjnmyk9PZRjs0DUWWKBFirmuC/D4bUI3tEmXMg9+8wS64ffB
/B7lIVTxvvgZgQFpJe1gCRGOWmvl2FS4KpuRgbdtw3LnFNAG3UugPgMXR2BxhQMbt7+maNolaGvU
KWE0IbP7XHb3tbCHHRK5cZ9yPxUDenzi36cZXSLnlt+UpeN9Cjjoj1Wr4BOFGlKgUWdENydHEWab
I8tbgI6Cfqlw6a4XVMyw6ckRtj9CGgxh516UZntLjMb/+GypedR1rqnEnb0dmGLddYohtb+P9PPR
bf5tWUw0E/kiu/2jozhPE9EKO/H73xVgK6G0WdDAcIPNgWq49CAYbMMghg2BVHLUZ9Uc/k2UXKFQ
4iUorfUjbqPzYVrzFQVgbB9yY0Ml47TqYziUkLQEhTW0561p4KvApvPQmz4aVUUjB3LXn87QV6MP
UVD/KhKytKkfHUglL7MJeYGVDdy92Z0H7uenX478iux3JgZ41Z4yWml3MYW0Jh7AtNihjvbSXxIK
Kqi97nFiaEjjnliqqNgXLiM3AfN8HUjVZZrMZcrImFfrnXvUDlbSFzhd56pauULoeWlyl9xGML2q
N6v6fdtbNt6Bwz2Px0MWlqJt+w5BTFE2l3CujQeIJSddKcn2RjqYhLGo87+T1MCCl/Q8JJ7/YJsK
FYMWK/HejqLB+3mlQYHJB9/Oqwf2baYYonF7AY90sWRYXNPuMWD04AqJrJUWjQkXa/DvAHVlCZQA
sV484/e/lSmTvDwCVtRKMLuXT1ffbKqs+xlnzSeaQswnM3t3B8xTzKGZYlQ42yaqtwiaKLqS7wK2
+QTP919T6dPbnSvy1tKAG3miyIA+7jUvzxcnID2lbozHJZtgHrIVLqBjApmUm7SGBuyNiQRsHBiI
Kr7gzZ0xJgbG6SM89Mt25c6tPUhNnWwntfmC0zVZupcPzw4j+3xEftcUNfd03CMdpfUShYHhQIk+
qTcyDMtUKfUMqjpxAqy5febuMXxdcZd/t3pREGecn+hkzF63sT0GKfU0hmk4EqUCMhiaMOQ9PfkZ
Wn/ZKJQI79u4UeO28pqomErUj3EWo01BtNMl/+vWa5fETuM/6r97nhYX40QpVnP47fvzht9FXjYU
+lmVPUsPAFgAy9UgA+UAOrDdSRDw9Nb2ZA8RHeXRyq8yvgd7Lly8D1uLQ8KH6vynUWusMirZH4o+
fuhA8d2ztaj1dgH8py79OxBUdmNt3h1qF3E55qJ41lYEKUvsYKYOi65vROT8Y4h7VzUbmqE/pIJm
r7AZvB2Pf7EQ/1PMhLOq8TD/MhBiqni4tLxcMBuA/4ti1DMU1vUTyU75Gv71x4F7UNL/xLelikum
5ju6pSlmbDf72tpxY7vzrW8zLTVPPwwM/KP911iBZil7Qs9IeEwB/gA5/qDiOvo9T8ZuHqQtWvPN
9QoDfyOuZZtiZZ+2Ad/Mjdnluhk5rWUMYjzFHjXC0lwqWFslh9sXgQU5UISVCghHifaRzq2w0YbW
oRYeqjR+QTcXsm1pZJvP/aM5CKP4xQ75SXgeIeBlb6cKgDYhhFhzEnTixPlIOypsXufTOC/2QljR
EUnvKt0wK26LEdvg8IDveR2DOZL7QlRWFK6BBCs34Wkh/LqXtosUgWRO9F+NubLGd8vqsBjgm5SZ
JVW9GsUSjTsfgBWWO2lMhabC1lLJCJjazf0ZD8X/SSrJq/JCG1+A1scEYmFAm/h7UtjIcDsbb+pq
H3FUJs0yiSZwa4j7JAhrQ8Nppkdb7LaEV8LeTmx2BD/PGvVf4s48iii6uZyHRLqrZ26rF5HluHtj
TNQ4un7PGx8pb5xRV0R428CjiylkdlbZ0OAvp/pgFisU1Wf17seNyNlNH0o2PdaW7UIp1cAruWVa
Lnzw0CEDnRHrS+TcMlALymXlWEXGhZhfSf4PYl5p83Vm18QHFADs/U8lwSUMe7HKJ8QZMlSvoACp
FFMib/GdbWkp1Pu8ILXvBqZWSpdXp8m1btpIWf8TMfzhd3cj5JMZrehB5ZpxpTlHJhg/kUFDASwA
Godd5STW1ETeWi7/As13EoUai1ZjPNaiLjU0Rnj0PC6geU719rr3Hi6oNvU57w+vh950e5phCsX/
s175MQ++Hi7wZ3jLre7oxmuKEhuzDDlF+ecWAf3kAdkx28fSOqXdDsmhCyWvjZqSQMbn1ARaRQ69
lhOInf0dEb0zDWpaR9m1gRtozxC2vxLpha0qblRaiRVE3BX9qvlCxQPdas+KlzXNoVv4jaIgEx9r
ujIp4aJiQoT9Y7Y3AwgS/uXBhciPj6W1+PiJmcgKteStDlXoC0llY4XduS3WRHCXRCc/HvizogMN
I5Pw0Z9+bPj692NbFLTc69QatIO/92GkktzWjAwNDYyLe5J0W0LpRkMTP8l2lGAWYckppJBV4orS
Wm4+1zM4Ic79kX7Zv15iElboExT8PiQP02LPnFH1ZLBqiEegeonZIveC8gxLd4WzjF9I70X3N+Pz
lkf4PzjP+JHk5A/koWmneK1jOyeuMV89tk+BSI+RxtMiDaBWE/3aiJ2LOq+er2b0XPqRF3UZcj7x
z/RaFS0JMLG39aIMgd5ck7AFfB+X8JaTzguDZPw5U07DWOoP/9yWFTRnTrahyOSB7ddNdSd6YVQ8
LF+hbtJPXFLkHICUJQY6UrV5aVwreavIzGXnzesVVOjACwy3U4NVHLv2E6QEkdLBUa9OB01Sam/y
sikQSu5E5Pyv8I4gK7MWmExgSKzerFve9LvFpEd4Eisg/kkglAFPG7o1biYtz6plsPek4pcgt4t2
ejK8eVqhIl2g4kEyUmfNrZ0vTXZBJw1gKHLG5k3IPeVSvoT8kXu6cDJ1whL7yu7Q3uXZuH817GiW
Qvob1Qz1M4G56f5GH5K6s8YUgY/CPlUl8ZrVUPLuvXhaI1WlWGmfOqBZvnJpTr+0fZTBflLhAa/q
bPuGWw18lOilc8z8XZPxv+PaanosGqUpMfRagFLS9al9g40xyVTc2/JLnmJRqulhDzaX6izQ/PXK
LFxh9RQz9a9bgCczu5MyIKpd83eBC7UL23k+j21HVvTUHmiH22QTL3kHg///9fQSfk5pqCMPNyGa
rfUulweVQCDyWZfVf29hJa0bmcdz88uMeszJNPjTWiItERMGSBBr23REvcn6v8hctCvg3JE4pz3v
8DV+IU4BfYGP23lF+f0yqwBJjp+rfRB304kTiGC76NcY/3B/WsYwNhBhArk1Pkte9nyzzODiEcb1
KJwlPzgUYjTp/Bzqb+pJ/DgAt3jx+zdTM8ZOk0JayxkHXsdy7ChIM3fymrJ2yAwqXPLPQrGtwhip
k9p17SvurTyTef6wfUh+6GhEdhfoe1Irb4LkHN60yWPHLrl2/AbPc8RD/l0f1LfPhsrw7s6sADmD
Ee+AXmATr5iscm070drnQ2w+qSXcBIJzQf2258fWk0Xp84sTwQ3hlxaL9yvrSsAWB0AFbb2s3hWp
pHqgO9y+GqfWdwE0FACINCIwCEJfax1+Wxj9HoM3gXSteBD38E89mLEs2crB7GVBBhqAhGr/BAya
U4OimFeK3StnIRsgp97QRLlNv5usyANa8Wf44HFkp9GNOoRE3b0hLx3T9ksFGVHFg72lc/pN/yt9
hadqIxknMZQe5K1XUY0qa0rjuaU2KHU2XeQgehIQNsaoDt3shfxIOAetk+lWbJU953OoOJVRuPPz
5iPJ0gL5UWPiOkU4nkx4SFN4tFbCNsDOflgekV/TYkjnz2UbAnGdbB9znZ0o6H/g8aTb7DBgD28v
H6JNXdaxqmc6/qOlob24djMkD0vDkp5wZTAqlN6+EA8Rox/Hi5LlIJggdHOuYC8axzQD++XkLTUH
4RBH2e7ZwWmET62eH8FZRlzJ6Zvb4W11K0cXeUwqt1Fc9eMNsfMsBOEgrdNCt6e1BFabrlAR6Wp8
iEzENV9sqzp0O9gvW0W0b+nZMt9iMKHx5ylWDC75OW20woNsD0y2QFy9dSTUmhsPQpGiP1XQMOZU
iw9nv3QmYsRCzVG7+TI9t0XvllSB+sjmFrM+LxfYU5D6XNxBOB0hPDqYYUrhwlJJFQqphFLVg+rH
5ZU9DFqDfo8FH4ez0sI/6gLh7S0h86dRjTrtru06nupYhsqQlZghciktwi7crI/a1SkVqSnPXp6C
EqFW2bqbFnymrGsd0itfz4+RUzu3+9ydJw6Km141pDaYVSfIAP4qVzkMZ4QuYripP8IZRwryhiM/
pZJ4/nlbzs6SAtkGpbe+aISTE04TfPVgikxzqS5N0bbQqreWn8qFWDh+QB3DDWLUePI1j9d9I2Xd
151r2wjcpQOSdCQYtOUZVvjHU7btd5FVgC2QwWfD9dIQAmLDnBUUZIZc7MUi3icUuQRkbNOu+QsR
8QbeztsYCUCBmN4ZBhBUOCmRiGDKc1+Caw3ozr8bN2WwYoim4MiHDz4OtbBfnkAuKQ8dHu47cYzV
MA4J1yb+E/Bp4mg7GCuZRNVWex2iofIbYdz7ohHQWyD7QUfeYOX8VbfINiE5rP4DDPZXgE57J/fS
+Fs+LHGocBnQlgDSER+THIJgHu7Wq0m9ikQoCoMixvhp+BGTVfo4bT6RqwyDH0raLRLPZTrHoMqG
ExkdwML5Lda+MTl22J8wCowSa+gR3OayiE+zGahhd8XxB/n0rFo7zuZ+8ZV6SNYxMPdYGGFkfn7e
Izl8EOA4HMsCxsbHNZZaWFm9LyW9bRDJYKlvQVLBj0aloNO3bZgHZKBWHiRTuJOb29K9dTixm365
anWT5ru+AmYTayMqXjJZ3YVlUrpqI3Fw5RALKb3oBKOn4iv1gN8oBHOhuESkMAHG7SycTerJJYvi
ca1bgZiTEkaqztr0TUiJd6w0HB5zafVXAq5uXHn9ufWKOWmXDnyF2lWshAREQ1k2K88HO1zTQfKL
qeqLFtPCszhC18JPuGlZfN51rVRKI048XZET6JzHPtX6OKCJaDcvsCjB4/RczIeTMyJNwmrWGOx+
/MLXFfacjJRAhuHGEoCWuVFbw50hsA2sJhlsm33CamAfHcRWMaEHJZvEwBBgZ8tqifVps0i/KOdy
hcikXiCxm6oLQBMuh1QRUx2LaJCVhdcfDtjj6CNZ6Oc5hNO5TrMEu9bYxKaLr52S/PM7J9IArAQ8
se+P9mdZFsTCJt8kFSPsiOAUe23GTVw0FhEdKuUvxCA2vx8by4Z8HrIp1Bq4aLLuMvuyukISZJYr
VCldA2l5FUEUcsl8ziDKYCddfoASTck2A9IZRVO/jCmvO7TkAN+4UONyaBdXpgQlfuBmsPd1fz81
C/Ur35f9v7guWkjqvXb9x7XbPlDCDSe5Py6nqZgRiAkNysXEIViZzOXQWK0qH+ULMK3XMVpaqTok
HwbUiKVfcIPNGT/VcS9vCCD/EmxwZ3vnR2H7DxHAPQFpyfx/QsZ9zhwKORYsgpz8ZximJwUi/aju
YQaOonNK/BKB9EBYKG0FUbx5q9veI/8YgnnECqQNC0J6IsQKDYd30pF52PPSgqhEhzp4/bzPLGVD
30uMXqpP7Wc2SMCaXzNLz5kWmEnzyNm1a1NDrSWjhGR+eA6uTB6cSQxF7cZ7o9bAoKiXJ4/to6vj
mu04YC/KC7Bh37SQkp4AFpzZawFj07FdDeVTyI3Ux3wd9AE+aJB15qSSGxQRNYA3z/h+/zzat7gY
h6ZIs8kLxOA5jCD3j6BFCHiN5T/hTDmjvakPyvsyA2d3x39R1yd9ELwUTV2tQZ9UbKxdAE455zHM
BmwjiCsiujVh2OaH8ACVv+gLv6e5phaE91MNuDM1AbifPPSPY1BqUrcxZEkdPIhNhzYF7alztywv
gCE8wox/2LviDuiAScu9YgTwfE0tTZX/oF5MngTmeC4+T12SaWFrqz+Oq6a2pIe9+apNFJ7kt26k
UoOBHX2fHKpTyevKJOXE80uhN7e+D4NDDG4r+1qfop4gQakUsxyR6GCYDLXjZLZoQVZ5VDfbnTGa
ICE+swtTWs/dC72FF4kI+dMQ32Cha6n1QrCscOloL7GIUPw/aqu3EO9Dpm3rtR0pUqbpR2dz8V/j
/nTU7yiWZy4w+Soi5uF4ocoBe7Eum2RiSaIJgq9f7Vds+HT5x+eLqkg/cM3xy8u+h2daD8fZ1ZJZ
mG6arXZYsBmg3Z5ImbhFXmUsMVIVIxQcHSD65ELL2POkzO7nEh8v2SOgZc8DnQbI6BwBWkS/At/K
xTDnCyjGVB4G+QhjkiPbrDIsPGEuFk2G+SyAx4yOHSnxJ91EvZhRaBBLayjp/zH4+8P/0vFbMsDH
NHq+Q+dzo8GdgWKXwnMvp9+e8v6ybHvMv4hVnKN+MKGlfh5Yn/Zw+mF+N0pwFHqNQXdOMf3Wjx13
WWD9e5xXGMFMvwlU3x9r0Y0oXMOVBUrCJS4d6CP+phqutLykeYqBfauMipYWJ8N4RPdjG7CBG9/S
vO608swDxtSOyhrPlHVA2fcmb4GyCyAZ/xPhz7DpqFx7qeMb916IG+b5M5yynATLDyVFpqtsxPr+
6tySLJcEvofRljHP78ej+21fANeKUQXb47vhs4Iotw0JLMjS/+moIPW0GRwVfzku8PIdNZ0Nmu2G
6nibiBs36j5GkpWhNVb0cIhks73bzJmOr6+6yiX0X+LftH8tFz2uDx3kYHHtqHEcTqy5FsPpkl2F
zl733JFML01Ld3IsOlobfScFybXLO/Hc4uuc8h+dIoVjfCIdBbSkirH6+pUcFKPdNcz1lwtygXnt
U2iHWu7N+9frTgAVhH/N+AoHZppHDPH8+J/Yukr05UeWWAaSzB/ck48+P+kE9P1ytgHdLcYLYIRP
gU5b9wYQBlH81SGbsvE8/B6R6K9tc5l/Ch+4oWM+9s5OQudMdJRLaf6WZvoqk1Ju5E+9O9ETJux3
0BYKws2+VIAO5OyxgKdu+1Y93vDEu3cAw/hdJLS7E6A9ZFZTgBOuH9ztSoZxv2nIIWsuUHycVsnV
IOaO8ozvkxGJauxD8UHHKZoKfPuNOa+M2ku/9sUllC2bw7SMmYpBuMDoA60ghi2K0d4qh9MIj+V4
m9C2uuLeuEWOZsQfkNWrD4SWysAlSUFlH7ekBLpdh4g4XXbwN4TkngGbdK2tiuAtEL3HT5rYaiiB
jD9XQAfIABiccKux3mrHyczHn5CAY4ySDU6CVHj9XbP3Dw6jHAkyoaiCYBuhBA3iVMHzjtDRjxec
CKXYjsSo6GI42ainyFif6DSLZF/1ALJtpmCbWz5VqR8+ymLMWFUx3gI2t2dsowh9EcRPi7vR217p
yjLi/skD2vi+e85/pzyXoq1Z0zR9Ro0SkX+QXAvnwZpgHAlLCbzT3BsPp0TploQXp8aEQfpCkRp9
0q30K6+5YEEoEKaaPIjx14kw1aLQyxbgyRZMKBlR2KIXCZI/M+W1pNtNGDo/P8JYj43NHoXXa0LC
+uFdrtai0W9QlTzMIZE6k6MlTKKSJqUbM19w0hPO6ezQFsz11BXfTuyzKUOOHA94Dr8/676ggm1n
T5CRmFXy/DVBSc7cybk2fF1dLulZKCZskdx8Bl6+dmPYc8rlQh75jcziBAp54v+pmnV6MCAGZPL/
x1j9QWHT00V6v5/1Gjt6gxkWm8Roe09gEynnJi2QpxIPi31OxKUGaEQFjcJnFTgISu63n82aZiXO
5VvXCthfEeo0AqWlPEiUES+z/63jY1OJAytNpiTeW4KzUDGRE+1TvLt8265mfYMPXWYdHtzGA/+l
NcbsaD4NG/0CILvLijs4vBYA2HXk8FFWZX2PAnDF/3lmNlbnCZsSppZ+D6+EyMEw1LRkRrarDmNK
a0bmRybvl97uoWCTNCq+g5QIuxra+kNmDM1Xl3gmq0EL+JQ3RILomRIvQecJNIAIdfreQvJfTr7f
4gC7x3P+Rv/8ZghF/z16Bm9h2yHEhNsWRRpXWziGZziAdWnz6/cvmGPfvjBpw1OQpw20xXThR6Tz
ADgnKgm2mLcLp8NKssVkeRCONQtk+vTza5DtrupYiIU/3U5wLY2X8m3P/xaXufH5m/IYaiSbOP96
xc6k1O9hTc+Qw21jK/sUGlCwcaXI/dwN1h9AAb1k5+pKYixC9XH2BFt0FgDrrTWO4BOBdO2GjJkd
juQ7RI+BdBGiaQUqm5SpLs7YVkvSljF2Cvw63z+K7+OU+w9E7hJBM9kJXpBBCnVXahhKyqUXTVoh
wPb3hdP9f4KDVAsB0URpjDK3Lp0CmGUaDz77CtdE1721S2p8ygBLwsn5VNUfRcuWIcZ2w0aAHHK3
IlwJJdPLLwVG3uYoUA2Hvn4GUplksbQmY38nB0HdsCeVMMN5Z1s/99uHjI9df2NWpO+Zl2kI/No8
wajv6gPUoQ0AF7BsWxyk1VDscHOkKS1Kahs5SZ8qRWoVOfXDfjPQN7mmcUr4VJOig0gvo0e6A+Z2
hiFaOILqcsXxVqsBY4Xmf3mGnT0ldF/V6IdlpkHyHgteNkixetPhudeSBCnwmXtx4yerqgEu547j
hRD1Uu9mFiSN0nnBmQtixgg+MKx5NsfPzNQqiF2+1Nr1mLDISTG9MORVUzEiLYXc+wRkrhhefsXx
NOhdf7AsOc9ZolmNRnG4xsTP+BCNFyukbnKwn3upg9rgP7hWvsvNuhZOAVLCHfZzANOgOCGkF09I
OiPIHijfCWf1ynByaWFLqXwId7gjYsfLuFvucIT9wfHPTG8g/n7enGFs2EWb8D0rT9oh5B4BaGWx
rlvqO3HL85UtjBG3V2hxp04j/x03G/fzG6qk5EgAeVSZBLd18t3N/fZTk4T7vl9aCPkDAqtCVgaX
hZ6L9J/BC9D1ISPSxEIxDz6hL58PpPZAFSHAR7BetdPxnXbt23dWn7sSy+5zk2wcB5QN5leeQjK3
sH7sCPiIDuZIm1bsxhTmyXcQ7ilmivsTI9pBn/FLqlKqXspHRUDVz/UE93iJHEs9KksrysanUIGf
Idb2figWLCOkojtQBAu/g5NRr01vxII5lhVwLZOdSSU0evRKWF8CkxY+oNscybTtEz4IicLLP+wc
oDJ9BYTdRZQERN+b7I9KdI566REnsDvnBAf0tAkhOpszKP/SGKr3fAArzhsHXM+Y/rCBsoMOfFiy
LWhGpyaXT/02GH+3lg0Vw05prbkeUR5L7P8XoPEfMfAPdIq5Wr7fW+jB50Iu6eoSK2Ls9XWXxxQl
5lL443WBzrr0mPAQY20lmEWks6mN6Mar3D2crrv+Rn1XZNdAZd/oSoT/aUel8ehYdk50xen35kA/
snRjoFZ9PWvg7n9RXm4tPK/k+wEhYO40JNF5zGQWP14HTfVlYQoUetFmoW4fTEBRXhv3/s2VP1rA
xGR1ZS63PVuDvQbUOSJ6VMDbuphDJpXGk7sCuBvBmwYNSOraCaTFOYz1LPtjb9Wrig3Sea5Yf+nZ
Vk62vYMPV+v5WK/eLwFAi62FLyuMe3ZotZrbBSOI9OJ9AuM1eFNS5U5sd80N+8n8xUvMLQaS5Fs8
Dx7QF0P/kXhhP1eRARp2z5D4Jdf84kvu4DO2ttE50OpN+wyqPIi5SlT2hsb4qhkZqKUlAPvdQ6qp
s8qZOut39Spi+Up7HLXS5VeEnzI1uY0hcdFqadVdrN260vd9wiK5meM6p9afxhMjnA1Rp4891RRT
3bYmeZihoX5g+mDxDld/ciWTgN8SENmohmy+mYPplZXyHVEz2S2aTeUsMYctVjnWo9FDzjVyQ3Q+
IX5AegRorejsYH3L7MSOQiUsC4fMhP3X2yXOtDDDUVfO6gClJgtxtdlYVYPXXWKEOFzgPKOzAwCn
SIY87vpdnGbuLB4+1DUdOgZXvY3zCadk257eYI0jM4oTg092MDkF3Drhq1aEK+gdyqtFEofmAU0e
78ZZChgI70xzofzySBNDONOWEqmMA7RwySnR9mEkpAwX7VowuVlUMJYZAduZh/FzS0dgOGan+OB6
N+lNbYv8QXs/R89FOUB/ARh6hmC7Yf5VAerX2zBI8dA6AQUIW0JDFsyIea0XKHyQgSzDKWDGD+63
w/M3GgBcV6V6jz1cAsZXA/LjAw/gmqrHc2Ijw6zTT5YYJx+d7Cc1W1kBFK7zUj4fSP/mXFM4K05x
aP8WeTR5iAGcv5x+oeVIBcUlsS03IvRUaW9H2FE/BXgZASFnmmedv3Kbd4F6WXsvkLEwWL7QiTlj
iRF7NU0Flp+h2wgrilRxto80NtcyXpSoo4/uuMNs/ja4ZSOwx4H7soknZLWBhAYE2v9gNd5MkIx0
iuCptoGgOcdmqmVgdYIoo0SzZqJUn9X/S0LlG9mOnQhx9ypgn3ffH/F2A8+JvOuJMsxv8xXeVY1O
RZIAAHZPYNqsEO+a3+30zDcxUfMNXT8jiQ26iaaykOMgXp+Ye8x1aL4cSdC+m0k7+nCVSb9Xcs1u
+2qzB9BsK3ogkuKU8liBDsVkSFH432tYdHTj+t2hsek6AJo6MDUt4X8gr9T2dUFyEfprhH40redf
RURougEKHFaXL7pnfyeNKhcMrmIIgLR/Lwmdq5V7c2NU9qb82WstnqheWCcvmJD/li9DWec5dByl
v/H9+kfvK6wLFD4wsgf8m5+ab6Ub9eRDIwV35FAN9KlhQJiDvv4bQPbC31ZF/SUf/ni8OtW1Y5zL
/DlWsNPpR8XHoOu+LtsXZCfWiZSe5UiTs35uCv7TBEuwlxh5RZ+lKRPPoRwWYFYq+Z198Y1lMxCt
hgZ3z5fovaoWEquhci7xkoufxGLFXtn7w5xXob/DLZjY0q0PL7bY7+glAOH7JImPYhfkgbTcbAcX
G3daTNz6QbfRVu0N2q9PlqDDM5nHz/4Nv3wUxlgWwkKH6eoGndZg6KZal2AXxje+pvbv1dhmEgHm
YIXGcH/j60uZc9qxnxn20hy1sILlU+h/AB7R0nIJdU3e0aPTQYxZ4XmXJf6qBWCl6BW7KzOazKRl
lw+PDabSGe4ZntVN8XSW7qe/izMdq//u1fRxjzwD7kimXaIDVp9N/VatZmHQJBkrHfsAR7MYkl+q
akAwdmFzKGYA0EKm+NG06tgHtwETbdmM/aFUEXWZNv3sg1+fok0MqdYLoX3vkhBGox4/YZLth3HN
+CgCLE0XmGd+1kN7qQDALaM+QfOn00g5b2lr6F6lSLbLyAQkt0znoOMq/o4Oz+u/0DjJPtUlhkFG
1/cPRZN6R84Ul18d1oxN+cg1A56NzANdWVrgqe8PU9NjY8sFbRTX1SS+K98w8jPhLoV6784161of
R1dIFbEI+9565ibGVcAmhcOr7sTg75WXXsoJPZp1Ot4Hfy4AvkaMjxjmvF4CPUR2D7tQnHlnY7C3
XOz88jLFcMREElvKwbK4kXKOluJTlpbiUYyxAvJ/CTv6Ovscr8p9E2UcOfRhjfMor1dufjSPKoBJ
SgDc5/2uXFWCvSc3Wb6/MDEgHI1bomZBk89CjEb+vZSq1Z3nPNvev0PkP1EDqsOFyQ11rp/BGN9q
VQyr6NXDsYR3NX0yUqBgJeC66cU2nibwklKsSitfpaB/2jv7jHv1djeaFGR25pnLiD1cEcx21gkf
fX+INZzHhfkIUTLNfbhXpalG06PFZ4GL87omzIzGbNMpYcOR1gP7J+SjmDj71gUGyBkzYvDHWE1C
1Vj77W+QCJqk415vtuGCQxpjFSR9d2jIlXa1yPNopr+Pd8Z1iAk330EHhT6ojcYSd9pqdufPrNAs
uMhEXzPDzyjWTh7bzQwb2eRyjF3VUJz0kv+lBds01PdqFgcSxtZlRt3vE4Kg6a0H0Ujb04SHYvCQ
ZN/sEGKWRgwrfvokN8vtUJtlyY9pP6VrRXYU8KSGQhbKeHzJGEMVt+MqOVYLdRfsvJG3jPJpoYqC
GUdRhjXwnjNFoczK8+G8GWdWy2fKFO27w+i2Etfguz3qExlbhYGb/EMOVgmhyq3A9OQpW1x+5SRn
9XuM6Z74rVlvD7j50tiWZEyAy7IIVYuiclaoVss0eVWFWoHdnabmKaqUixK/Pl6BU9y0xB+zIXXz
Tv9+Kpg05iRUbvjlENPWpqAIxRTmWaw8MLJZ+I6J3Edmjh2oXX/VAvQHsD/vd0Xkc51QdNbFNf19
ntAP5QmT3N+1jb+iF0KLojc/JsAzmTvz8Kt+Qwya4J/x1OkaLLOBsBnyygxYUrXrHoO+ayoDYTgc
x8nixZ/jwXlacnU0WhyGsyNOhGndZQRiITVBkk9V0wEEkenaXWzK/laWuc4kj9fD60afH/uLeqE9
EbpiQRPrTPnpCkst5+KnbJX/H2ohBYKd1+BNEV0c8+lDTPuqyzUzuHT9UCDmfF81DCW7Grvu9HEs
aeGf51wi1+X5BXDgPoRtL1NaG/q9H9T4JQJmA2UWkcufLHjBu73xCpY5vk5/iROBhrcOi/LtgBsD
dWc5C3HXTydmE3Q0nk2CIUjuPL48rpzsoHMWpjakBrm1fy66WmCzsMyDx9c5kvwd/KmxjOqQSe6t
ws9W4q0KaAWhlUxmh4esnz31Q5W+HBuKC2/EQBMBgce3sJvl4rvRVPlg7pffg7YP2fTvAhKOF8Ta
cLd5Uc2p77Ui19iAfcurbTc2kWe7fzjD0G2CFZRMiPwWbxS2qJn1btIxx8d+J6RUAHXCH/ROLs4g
lLSswKALKZ1cY9+l0cbQhQWB2YyPLOCX6RW6EtsmFReJQrEt2wj1aMGqCPfPz/Nhm7oIzf9zKozK
+CIj2Q3AbcCO9QAzQbYk7mDhmH4nYVOLkD2ZvUKUAdISqC8CNabXr0qHOsvd8k4xAesOyiBUHVvP
+LSQUJF3DoVnMbR4Q/gGhd8MMTCujPY9O78JAP0uaJsO//Mj9omcDWg8kjB+/hMzuQzXbsy50v9S
bXQ1PbxUaZrjSH93K342xw4zUuDUe24eXGKKjYef8EXsUPVREQpJG4bdTM8px9vHTjS0Ac1ND7TS
911ofAqoyICTAOWNS/hbzGOZfl4NcD1zj7hFYSjs5553wjV7nPU5rr6n/S0nC0cHLyU2h+geCYxx
DZHav1/Ir/seCeF2+FIXJ0/mlDdz4+c1ddMK7X2x2XrLxlf+dCvqnXRBdd+ghP5/sWez6+7gFFTp
zAQp5g+WnTddudAjkgHmqA2Tkm3H673DaQSpbvmhEQT7NAFywyyFlJ3bYaUZsbSfQBfVgFHPwPlv
tpgRylHCxCMrjI/VGbFRXhkAJ0hySOT/PFjUqBSCl1JcnGQVlc9kkPT5Q+DOc26kDs8/cujz7Xcp
bxHHoKlPFGjwsSY21Bk3Ycl3dfD2r8dptG5AQufxCls9Kk5DStLOmzYzdorcj4aootcpD4Tu5SXo
QzxqaARA2rhHvK21WqfYdc2FvbmYPNXibNFc9bMtHlCtIns0F73Ce5EMyCazoflFplgZIn8vxaDm
lHWT1gmqfZhNhQi+4l5IbT31WQhlCeN4DXf6cj/I6QI9FP287x00WPYvFxdTV2npXzw/eYDwwXjR
IqhxvyiEng127D9/0uPLKpKkRxSHcjdVpKCL9cJZXXGltec9+0C4jYwMC7G0ffCxBevxapJ1lSr1
v6Xo/alh2zIZuZovIdRH5QRAubfEiPWwXq/Ke8KXuiszWkTMDnuaNAm9rlT+ow2CPyLsJ82+EHJ9
vPWp2zIGwEalw0i+hzwUaOEfUAZb7KPxZpyqw88R0hcUaeoNU5NIdGdarmkg06X++/ecSDaWG+H+
67i0k7D69yjTlC4Em9kZkYNFk//Q692kv41f1/n6YjPSY4/O+zTm+Rab9CyHoMIuWX5K2TCAsSaZ
1Cqxaj+vXkspqo+3OwF3ZYet49yJcRanRVLutPMtzDA3G9JoLBuvcjzpe1l+/tdmGn3f3b7tJ0dr
M0utiksOxTSIMvBltVfN3YgmtEi7VyZ1a3JiHRo7BNcQtyppZF5M8BlxsSjmCJEVJPDduGvUzeku
x3hRI+yFGv91PjFN9mfHlf/Pgi9zvtNDhYyMVlvZD+RSJYzyOVyT6XfoBAw6R2syLLYa6/l0S42t
jUbq0B7EXc9kAthSTo/Zc0URKsTC/88G2dXfv3aLVajDqQtq1s2QFB9BzSisaf++RqzqJwUDtOCh
oaHyfz1iYi4PIyLa2oCfYvVoeJg0FoPRaacMlgCJkhdtIDcp+l9sB4Qa79HqjGar4JqclaVMxQ4Y
hVHsM6IZYj2h6+36MOJD5kQazqV4ZAfCblIq3b61nAKTV1D/k7Zf9uQPIO7olp+HW6uiIImrQiNz
8tEeH2tb+B0HkGdq4cuQCmn7BmzHIkbmP5ofWbc2hPLJSQtkuLEAmwTAsv4TudzXenDmzdvNnQ16
/dcQ9Xf3LP5E/S7Xj7QG80xz/pb+TXxNvCIiW8tdfFJudzFRlF8G3+9o4UrLdLQNWzCYN2Q8xHoq
cVHHlsxJbC4G3FctzNoaxtIuXDyOVX/aItd2uTZEcBWUyCzE/ycjgVvyYCXk0fOHwkLhOY/y4mfL
UL8Vj0SmO4EXYtmFYzQom/XE+d/hmyVLiOFxpn0761/Kqj08OsKqXR2YkHUxVNLJ6wWJhzrtwULS
T0zp5Oy9by56XXF00Vq0HgzOiOWNfoT+uKUIbfq0hsLaDKlDlxoQ8fuz1QWZ7IHddE4l6+Kbjoey
A2dA8CwabhWF8KYlVxqcoA3HyEbtf49fkPYf2bEkSW99TOpS9TlTCM0yrEdj08NkL+urteoVFgpo
sai4JXfO0KZ0qL4KZxKYKpX985K+fUQT6jATrdMLU8CPeia6r/v/wm5wuNOYgkhgQC913QzmidTa
purXjhW5k67HeoLN0emBY/su1XnCJ/wRfhCIK0sNsKBiCUDwb2nb+LKUlCdZRsvrVv7p6O36DDBr
raG3cE+zLvK0kKSwZ7FdQlqc4HstvXKA1uyzM0NveZ2eSBKxJsBXrI3/xqgyHWcZn4ppc7lBQrP3
RtcZnDMn2ptPWjUYR3z3KyhCzhnLD0eMzpF+yRAusaYE1lBG1whJHpF4alj7A9v4N09bR1vbUpxT
9rr6pVggApC7l9kLy/LcWrESQ9H8wm6rQ/L9VNfyGmwsYkBABqC+UvVd9uvPMBYFgf6Bq6B5gOH5
2cvpXWo213ivDo7NF5jMQFve44olY10B8/EfoanyManqWaAXtCw7wbQ/3JUmLhCcgU+q4us6fBrJ
/9IUEV3hGOhoIP2wGCDxfnq4iYmRdKgEQhu4ypBZocUQuK9VjAZCwhhLmKz9rztzedupx4P2ZFVK
SWy2uxjovZmTOVFqvlRisBDjXT3LgJoSNDyOGGnBS7kAj5JIDBrrxn0fJ7Q+G5WwBHG/z0Y2Z+xk
7v3yraGEwz1j/NE5YucXRBE/XPCqnKyIcfHn3WDHsbH108KjbLOPdLXenDYA4H3f4xou6IcFHWun
2LAWN0EV+A/UIVr08kXH6y9RrFHrkAd15zxAh9mvWuq1RLymfojHyKqt5FTMSabUjmet2Cu4b9W+
JqJHTaISu6dP1O6zOzN8Yx6O2nXAHdkg3LwNhC1N2c+SWQTqpU10EIqkJ2ws70af89fKuX84jrk5
w9kEMZWDKkgvYx3/biQMYQ3h3nWaZ8cGvggAFPXfo535JcUXkp+EoVjBv9Z2S4BCdYFuwnpyt1ur
OtelWgmuOPB0taq7wiGToJpO55cXprbDPSk0K2TrK1slyN93AB+Wc5m43dhCnZYD1HG7dp4EK3GL
rwXjU2ro1vC2evMOvGE1+e98a5Ux8RA17JhN5vB/vElfwpdtlm6vyA9hk3RjH0ncC4yxV+duMhhN
0h5yGWfA0y55kIfDoJ5mgc0dHQo3mH2CXF6e1/SIRjUpa1+yuAiyMlEfT8bHkhR9ruF64A8Yk9NX
eyfofjA23+VhkNN+LLETMUiYIppX6cMU+bjA3eWQSSP2KP0YmhjFZzhXkpGSUktiu4EBjkgqbMpx
/zPLfKc1cniQLlSFr9yhLh0UOEelmHOh9DrhOhYDXAB3GPSiXYDkO7SlxnUhjr4qbELXncYNtr/1
LfcoXImWxJ4x5AbUS1cPdGfoKFTQTGV4Nkw/9x9JPyIR2wWLGg+xcwO7DerEiINhCTBaI6BSC4tP
qSKCid6/vujeySsEyoqmmmORyOz/vIwK8dWY+oylhabMhLUOdq/pbQqJkJBE08MgEa8XU5G+/F0j
33SsbNkbxanHBMwrNT0/uq1scAudo7w83EZLRnr+1MCOijmoupX21HOF0ACtX8eQEqoIvVjleUwk
e24X50bpb1ig8zpiq3IRyvl41kQ/hmHCFgoB2XdsF5cLXVTBySyo21909CfcWWk9SnheGu5WCeYZ
HEsfUncudhZ4VDPS1W/fb5eVxSYAeXOxG3Z3U0WnumnynJcIBYNJ1XhUL7p9dqrp/JDeMLbL5dnR
vm/31RcwK6ZUthGOmpbaOQK+1xBclBDRzAAcyPR9Yh/DnQN4VQlloqtYOOjCW2yPu+wPubGxwDu3
bUsgadKvo0fa1NoeQWD+qSWIBy+CcuNdN+e+Tdx3ukQV+U5e7iYNmIB1GsHPRpfaDZIq/N899hv0
n/3e101BGMirfU6/ya7mzZfudnU6feiEMyIg0VAGwJmq7gGNTrq5V9fVKaOuTt8ZZKyRLntUpm68
6dQ/f4xayjdkFTLUzUQsU+h09Z+fHEWHjGGVx3u403xQU4MDFmioR4qufV9ClbNNoHx8c7bC0h9E
tWrZwZNpKefyCRMHewR8FgyE5JxFg6V5FU/kPqKFO9eX9wuyxDWX+/X/ZRio1Dx+Dr9gxa2DI7HG
3cGDFNnTaYxO9bNJ0aS098AA3JjJZ6mri0BoFROQYzNbAKc5JUWKp64WgD+ZGmJsPIBCYZ2K/v0z
Tb3ihsLRhPVYzzQD2ZuGTEJlolOF5ABMxW/UJJhCXdEaVyQvwG6GRH0MpJy+dSr6WN/Pmk1fy+rY
B4i3v1vYbSoxItHPZ4427a/wtllAVX3I0tpSn2xCNgaQ/OZXquWUDuNvewIyeQf49fkZIc9HLlJH
+zN14HnGP03kn28iBBXtUybF7UcfKPzUuYQL4agzfmkeoNnM/3mtBOaw7h6VGApAE0w+HxB3+9fq
zGO54G/NdUDgOSrtGzZF/8kTJhZe7Ppi5UGbuNxBVI5nsTC3mn6+uqRSPBWW6/2ILEH4BSivbTir
W186Wis9yVCOquKhIANchs+LhAUa8AuSBMuN1UqW7CSLu+udSz7X9UeFHPxyy7fLnHR/tMIAflRH
min6DjtJJXx/gtG7frZsBCwM2irMaO7FIdmy6tZcQumfrPxsVnJg+s8T7DaLDI0X6gUT0vaZ67s7
G15htexYNeqkVtE1dMXthowKyI2CqZFgehcqu6MLq3HPKFVojWf4aN5hhEWESPi/2VrCOWGZVDdz
HOyl2vzenjjzvRAIAnX/S6agGrJXeaL3TKUF+IH0GAnVgq1mzRS/TqKcWZNHXzDL/0+v1qQ4yROP
AGX8dY670yoQgGHmm26QCmx42p0d+SF9SmOxaae1a2atYvqnjVJbEOIIYZRMzv2afQEmHeWuLl8m
P4BMJLt89sg4YcwAnyXPii6VdEdbEIV9A++ejNIgEZIZIhK93n/2kkxSSLjTE13wlcQPsmw5yReM
VcMtNIFyyx2g7gdQQQ/1vFugmuxiOv2vZiVt/Qky8SV7Ojv0ctNTUhFiQinaoPqanAynB/A1rB/7
yllEFY90VsWzbeurb6I2T1LicKQmmKXyAKOCwTtp7uHb2nelWOtqZOffzxNe5zwHDuarSfNzuVbV
lENEMsIapu+HXgwCOLRVRSqW0dutf7CIhYX/DTKvxeGVLDdeXLhPS/4Ni9iATOgtaBBG8poSCRzX
A9JhGT0yUUzDYyJ+1SJn200kDlM2RmMDgrSJR43NuZFf+FK1bEKwwMsn/s4wq4Gobne6V/owVxQm
IZ3TqMEMvpRrxIRzCEg/RX/WljCC9oaH4U2r1DmJdgtZzaSGrqe+dqsmn59dyh2124XGu4bK8DsG
3gIkz/+MQJPm2b3htYpAIgC/H6g2TK9AwXT/EhYyeEJ+wyMHw08nNUfcyPDM0kFtaFSKZtIaeDoP
afp8U50G1DuBYlVQum05GlaDi19wkoZAcXQFYAyT6r/cx2drSsMO2e1ubKNuh6Dj7pJI/a/gX8lJ
8/IYjLThUzh1lQDatF6gVaVmfN4QqRu6x1NhaYDXK5IAXNdnjnU4SWHPNcsEobabe5c2Ngs5oaga
nxs4R3pAL6QSm8VKS/Qo1O+Cpk2P7yQ5vGTF+/W0x/fhg0w3P1VIK/U6wQb6P+VmIwzNEb7PWcmu
Ogqv4gUjj7SfdDl0iSR9JRFxchF1h1GKGAZws43fCawJQVI7ZhiCiDSDDpNp5syqzlSldqqfL7sj
7J8mDdfAtQdBBtOkra0AgbQbRgTkVwiSvJovaZrhUK5s1OQumNqTA+mtZzsHEa36EmxDP3lMyxCh
3F4eF5LOn7AKE6jDA62Ab5BEmx2htdKYUc9Ked9QgrRCRDIuwpgEEQ/SViXhMH3Y/kKy6e7rnUbc
W3cfPAmJ7Rpfpp3gKtDUz1k3LONSe/1RUl2Z2KxRxeWHw3/vgECOa7AhDpE54UIJ6kJ6gIxkd3Wq
Nndehontb0cSAEhzoUd+C8OSYBO4TvLqPUxg2uwrq9olJuYKOixXnDc2UxdTU0xFgbfXUXJST41i
Fcheggg2BFLcNcDRO3VBSoEysFWNDFKeiUVEEt2jjYCzTiQ17jPUaKiT7m/hFnbF8ryPyi1U1G78
jkd7FRX8u/VK+fXzS4egHx6HPkphOBz9s07ncPmXlZVTppF+G0qDofapkxK95M2Ffn0afdNQz297
XwS9w2nM3jAwg8+oLvFY5LDKYj527ij+g+w54AVimSLmo6JNmqMNKSHZ4KRKwmip/6Yaue2EOPVF
OFbJQNIAC/DL6l9oDgodFfNhm5QPbolHMgMLNHznRnirxlb4Z1FZlVxFf01nBWbMaOvcJRk7Iw8Y
h8Gj9cEPzD9IAlSdUk/dA+BB2QAtsIOb/Btg50+Glrh1gsKW5DeOrdstJqGZPDDfXylTDVsULhSa
nAndSSaeHLAwH4DUV8lGowqtel4PElS0U6Yw8XKZKk29p2sw4JBlLPv691oJoGZuJ57RjmLFB/2P
+6IC73D4Nzp40ZsWBcPB9v5qdDvuuEJ9gGKTYRWXo5SS22XwHHLQFuQ+UUcd4V+Nqj+EfcN8TMfW
R/gxiEBJUGij1OXD1ZqEXk1dhL3feMenulfMSSnjYeoX0vwlOm73w8mYQ69NhxbxnsSdpILXKt2G
nupUZmtmhCOhikNJ8JadGQKt5ClsMwNxWGBZ6tcEMhD4AdG5Ww/NCajWzbHGOHZONGn/PgeGVw63
SLRPAAVeD6oAJSLwDTyNRnc8597T9nxYBHttC/MaMZ1/qB0UnSAWtO+15AkF6a9oOHKliW7aBgJe
52/yK8qHOfF7K9MOukWi0nWNOcFITe4LezYGztSSQlnF9PvvbYolpj4pI6MyW77BUuvAZRqkOCH9
kLOXAK7jNWg+UNB+r2Tzu7r5LHI5BxL5JpqOm9gWv92El2a1IxDcwgBVY9YuCYlTWOBv/DXVrOqR
MlwyW5/ZVedy22ay8tDRtF9cscmfY7T+TIlH/ZLsbUKFn6p29RpA5NQt54uU6n4/JdIwGdX/CkyX
1XQ7uFTyInKmuuMPWd6G9ee9fzgyUtZEp5pr6n3jimcDsPmbe+8pj7wOqRuuapSH8EeQ0lxDpMRO
ZBaJqPw941Em1UAZqFp1OiOKb6a2tCYLoAIYwVmIs93tJ98ryIeOJUCR6vnxYdHR+fl2GI121P6K
eltdqsome//gcJLT7j+zLMUGKrQ6+xhnqMzf+1rRxMWuwOc1KnIEIZUvl4WNvjGSJ1t50bHk4buH
V+IChAi19VhDkUB5g4w6gnv/L9bQwVp+FUru9uZKyAJTr3MP3lb22tiBfCdqaCrEHq1h7M+6qql3
1rD+OE1yAlYZFhRno/IFg7p+UtVW9MQT2O54tkqmGyL5amFyHAY+U9SoOp841ByGUfYut1U3Q7yc
FM5u9HdbfVMLuId7qohd2haxbOQwg69eiz78ZIOGm5vwFnprtZWZ6qSgiFoiqhqXDTsPEphj3sz5
pglavOnxnbVykH0IgoGf/IZm5pDOaKquhu9ocVDuW5ZPOsHM4X6FKxiDlG8gefNIa8/YbDRucl9E
7YvcfWiv4z83ntPX8/wM55i7HLtfWwde/N6GEBYos2rlG8pK8dv6crPvBe+n/AastS1Qj4GGBI36
jVugFctCFscJiPV34nx4oiKhzIgvcexPhVA/1DLYy1yE+md17FX81VtB0Ujc5r+KG3vlgcGhHOQL
rhmg86JVHJzxn8AnmopZP1uve128cOOF4huEZkPXjA2sJNWXiPG0CF7cR+VGNjPl9XZnqkuCZWKb
XgVnzqokgcfIlKJBjtnqiPM9K77iXCuqHCOry1vl/AyBHrKMuNnaT6EU0PTadqx5oSvE7wXdUJXi
sT1BrczBht5+CxOEL0Lm3PGm74dx6YA5UDCnchU5plcqetNMb5L+SXCJ2ODAhuz8LsQoZvbFnISe
iGoyUL3gbDJmsxZl+w+GQpZ/JGVvPXZftnl93AljOX4wYthKdEqrMWL5dA27BtNImYToh13UJO4r
Tsu/EvDSMOvYMvRXkk9UiX48vcmTwaaNFpQvENTB82JICiPg5U+M6hKn55kU5PBOzvYC8WLUK9R7
fpEgO2OGd23L9/RW8d260iErlk0P9F7d5aqvkZEx61zwpUCp1x7gUitCmBecz0B83b87z9ldcdtZ
sKAZEQKyWz8v3YayZfGMnmtcVt7uvbjOBFEHG09LFJCnVA9neSvvHojTIf6KDCn8Bv17p9/OI5Yd
D6fEQPJJDdsyh4mMjNCCngxR883YG5FqFaqOBZmdW7WM+cyn06ujvpel+vB7ZbMoQ4Md3cFGZCs9
F2n6JsKE+LBej7Woy6grLeNiN215JtDrMr3t4iSfFlVi1GuttL2H17uLOm7nH/e+MtndNpR1a/Li
XCIQ+pgRyiNTs8f7VVQEuC3spKztFPm57ZeA+w5M2Yqav97f3E5aBpdorNgbkKe0GPlU7iKY0ds9
RclZUu+NGoCs6wyiDNXTx3BGmcK3BG0vE/xEBkneFWrcOg1muggqRHu737yvKTW1VwhNxTsPgGzd
KtPK0CIeQhSUXDticyk33oVKX0JGLiCUgjavn0lb5mn31e6srGYNvHzsaEwdDzkIXDU5LCMCHOYu
tzo6MZHunNHdjcn8esuihtVYWt8Njx7N7ID1EyEuIagNqjpEv7OiucLvavToB5hJresX6dyRqzEZ
Cj7WFq2Dhod5jAE98qb5sTSE4O1cwev/i2AjSAt28p4b98NlMPmf8LoIJ3x24oONEmV6EDamz49g
XIJoPDXc3d/Qqz7bFBRbHWPa6GWazahKxjHKgDQI8hDHCNlHibjWN7nAk0SZvbGZva36wRP6mFB3
wAA8668TedQHYaUXNT5aAmFajuuY+eoWBsns1AWts90PA4MvIYUZAq9m+gfiIeILHQTNzcy5PJ0U
AhDK28wuj7NFBThMrPJ/8kQ1c/hxTZlAGS7MG4C8U57/s7bBbzukdVaEfiwbmCOq4PG3GwxSkLAG
rqQIpbkIWf4YBX595oavELWyjJtNO3fejWfIyEkDp48SeqNOhMv1wNCQQIIdglxKbCs8zH0IM5E0
5h49YK/VfKc/BOBae3h2x/CzlSP6CoIpib4qm8lQAMZZlDwYbO3pamrz/9+LVXOKRjrBHz2lNEh+
pv3cbwWaKNS0AUDyzPRBqxRTiAJQm+xF9/pqfSqPiRQjyxnwethvSKaSaIN7SKbVebI39zj55Eda
1OrhRp9C7mpUncZydpkIjrH+3bGXauXmzZwkAeXflNTaxr45fRnZuxR+MZB7wZfEmfM/qZus32Ks
nub7XG/ySDsT3dfO29hpiKWRJ67GN3t+IN1sP/b12ZIJTYSh3b69b/pW5XD4+cpsql1oHatsGeWi
6RbtD6hrwJKCdO9ITDHIxBnIwT5x58F3q3x/gHSl5ZcwnskRfkysPLBgXXghueaWBVtbOA3Jc4UD
oFmhdBBDG5ZwtqzZ457KJN7I4qkM4a/IX3K2NStzOPCsnqDwrhm7WTMCa8E69f7ucX54wxzQ+I1Y
ZWuzNVQyRXhKnUOZh4jhgqrAmIrHPAEhfDshc8v1HQbinbvhZXwmf7AEKfkJHKaUgX7jMjcePZFj
nn4YN4Hc6hbReB8572XvjBIZ5olHlXXajMTK8xQyNTJZQSkL04dlzNuHzEtRUgwOuiv0yhI/LQpg
vt+XWLfyvyaV/0AgzNKDrTGCn2IOvtY7MWxJuM7g1P/NbZHjl/kyAQ/9iHn2VMVG5sVBopRE1kSF
GXN4bIrfy1OTtPA2ug0m7YH/FVEMSNGXr+FhVSz2WT6RG7UgfnoGXgVZ6H0DK3ulonsfPc0FNpUd
2wgpcPyZp8/DKsFU3NH3eygSlLcoNZziiaD3rgGL1F8ltthxYjDTWijHipLWOTS9KU6xT2CCS5H+
1zfdgI9MlJfek/VyuATzOqLa71Emj8UV5Y8y3CKoFxxR2+J6NkVm3r53vNh27nDlu+XTWpFnVnyz
eB9+rYpWWd8bBnbM4m4oHxV3HQQLzXFGisQoRqBTJGTeZvdI4kScEpiQLny6QCwC6zC5ULBjZCmP
pVVJIovOXqesLraJLGVqvjB/zVwJi0KafbICaduHwnF9jv3kQ7tX/hxWLZDkyizzUR1g8boXp3FY
2FETFM3dq9f9qtuxDJS8HZSrTER0WSblfggftLJ/NwwcoO/Kd2o6XxZqrC86boFmsB8m7L2g7eaW
NKjPCZ0K4o5ahPzWbw22ACJXY6x1PaObnn+/4Q5Vo9fbGVgiyHZ0017MexEV9jVeePXhvYGiuv5D
MIBKIrwTle1WI7hkMyA6ONbLfkAITd4EX/ooQy3deQRLaOjrTRiX7oufR/h9h+NgOO4aXnnLNHpA
+IrghQp1YCOlo88EVwE93nMdt4ml7Osyclv0ohhcHIOnCJDJl4HP7935aH/w6UvMlffYANG+AApP
mTPXpjYdI+Y/Bx5vbceMwFK/LinpzeUbEEpPu6wmOA1c/ssMN1wPPTmO3c10Mt7+B7g8bPbxa8re
qadzY3iL31oZmqEmjGW5NAAM0Dz6Krelkp7EYoqtjjJkIyLZaNyg93eZUAauLfPSc94GO6y3aShV
b1r1Ptstfm88suaKmRz2N4MgSMWAGQsQDuYOaKtdioUzBEHjMK21mxzIJaDRN8pUNbSfMs1zFmZD
lMXRn5Vft545XYIUmFsH4O9D1m3cd3aigTlg0zFeyjO7uUSihjk7TurJiOUSuIwapdu5b14+k/In
cG0U4tAIgQ7lqAV1dIuAGO4rdzQGs6xzpsxf2g/I7FYUbEWIp59X+VmSCyHllIUhq5+ktgBiMKQa
CE20Onxnjrz8uLra0lT+cCaCoCVnBBHon9dT2IrVhdHDy5kRqWGkkys6S2JlCzjrluin/JT4/eJF
XFL04ROO0t79m8pSCXPIpifh9PpsTesELSHl89bLk0pH2UKkprNfYY5wz09XUbO3PzQBSuTvwJ9s
5AA80S05HxIslf0fjO3j10ppmRcyoZD/yDRPGIUJiHN5hP/QY0wZ8hcNNffjUKBWu2x1l5ID5sUx
v6Gr7NLdcszM4wlXCLLPYzcdv8bM47AytFI532frS0AkoJl3jUvkWDCpplpl7BpOjDRXLoUVtRiG
zLwSILjsaYpaPjd71/GqB+XqKvcVUDLv/rugiprO/limlWdnP75z26kCIAqFj1MS5lVNcuz/XU87
enSSaaJJpNEijtXkoX8N437JZBoOewFk+JrdE8q/Od3hjWskjMg0SbziGCNAcKhJteRKzwZv1yp3
Hryx+MoCpCCoXHmCtEFs1tWpXC8NBJ4G2BQtePP1/cZsJEQkgM39miEH9xG+KeK1hR/Efr4KVFW6
GYDdaY/jwiEyBGGagEo6gThI+B+6rSatHtYLGeXNnXooyqo44UKbaViM4N+9psCMmbcFeXdYxNAT
1rKpjtJlYuQ2ezBc6GDlbn7hQm6NnXQOLlpbIIZbYpZ5cF6oelh0d0CJYaKRHhDpql2EOZ+bgdoM
MULUMFBvIrdBZ6KelapUYFPpdCKOdQVcrNYe6o/WJI4m4R4gBpVEo0qHch+IO3+/5wAdRI5uFEOS
hgCrCgk0Dsm6UloMt3opUUqR9PKR6ttCjEly19M7YOY6GN1LDz2w3mG5vwBeo73sXzWAnC5XKOM1
NvCNhQUaBdN0agtuimd6pMndtfEezgl4B5kaekFYtk9N0Dx0j8pIvIwoqXRrHUdztY9xnB7g9dlD
f0AItFlhegrdlPrrRDU1FhRl//lnEqLRs+tMfYS8FskoSZ5qSUWRqEHkFzQRsQEjOPHv3qO4ElX3
VAq7uCT0c+nvqdWAEPFDFpX7UBpLxRws1otzOl9zR5PX9uEJLUwPKf8JL/5iyFHC83we+foa7o4l
yTVv9cWgRRblQfZWhVgv+Awgu/MACql6BaaVpyMjZn4qiMmgsZnic3Q+Oay/XkWdx1fVKsweS4Mm
xqjrG6RNtsijvNlUqG7XcXRQnqrGx2Oi2HaVy6hTQQVkAIjI2s/TK9kEFoSVSLanswyf1YWUFlXB
1RDzsHn+1jn8yaW2vlKJ92Crx/yjgc20vDItWASf+S1/3j+uCprUcb7YsNwx/B2np8sXrIHaEyDx
rFCDqSINRzhKPKb3TJCfJb1BP75AOAkGoaImcxsYsOqyIm+/A+vpkgK/YHunKMxVnWOzmlKWFsWk
obA3xv5uDSUqGo8Xa0HpaFUCGiESfFX2iMABkWt7cJDw+u2SzwETG506cUMudQ08xFndWyYrtiLq
7UMXM4d467QA+d/vm12LkLJ5PozPH56KjZNb5FPZHrQ65HQ5abHhL6g5OQB16IWAxvXfH26DoGvV
k35cMnCwWDobsxw1DZj9f5awF1avEWyxhLnYdyFyB/4tiCEZmLwQJSVW3J28Z9IqD3T4f02Nx74q
vLo4vHh+9BTu4misgKtqJKj2xl3HsfU6yGA0pjnCR6ztl1xTiLq0uPktSV5mhi6I2st2FdhrTGOG
U8xNyY2MKxabYfqWKo1tba/XSBe8Y4MXP73UkVsPxtXuI92UVtX8v6jtv9Ygzz5mLX++Rf0XRROT
ulKT8FdLqwRsT6iGMDpUneq0c4J4utBSsqSSuWX81/aVDzo7eYGZEFKaWv9edOHUWtEF+VRK7ubB
eGd2joC8BqAiWFYoUcwYDyQ3wXD0Obgw2XKNRCHGT0j7oLXlR/MGbwuXXHFjTCXMEcCVQl3vZiKU
D8Qc+X2r5x2/AGiqcFQ1zOr2F6Ze139GFHSbIONcOnQKXvq0h904ejKXbQ/Ec4TzcvOUMJ6zleDL
HTOd7e4bXpR7hHbqMAVtiRmPMCVAff7yoT+wydVfBNh7/BDbLLYIWT/zQ4Sh66ufqxYgM7DuLVc/
nn0//1bo6s2pi1wAi7glW4+hsfi6e1yZXSFDxE/2QccDL1sVCBL3IcNiXKcRcnX6Eh242ciw5ArL
lveOqYQxTn7oHVauXyIh1z/hkUn+EWNZhw8YU+fsVAhr1Ge6ngSAZE5vKlgihT3AUTXZo2dMcvaB
632SMoKhtFkbxvmi5WwV+YHcpFD/kA9XrvtcuR2sQOiIPeoGznLKm9zMt92aUUa+fh02CRPvTFnA
xl+e2E7TqgQ3vfL1vxvizyqSpSlwinZ4ZvAf+Fxvqh2tZyI1f6VPQILjq/LwSb3VU0XB7a/lU7zn
ys0KfGNWLaZvSmNZTWt0Mfp/JOLCKaoYVU3NRItP1aURxvXyZcFZKC7aVcXDpeeDnLwr828tpofm
tcuLNxVpUtWVemXLJWZBL+XJznCknSiC5aJ061SS0+vWXFveHRIfYnY+H1AkmhSNV5zg4MAOv9ci
GR0JDvZnWtmnDVTCOJlwNlAq7bzfc78/E0a7twQn+vATPVpDst6Q6e7KGAEAdUmShrxs/Fqgp+wt
qfdEiX6cX1CSHQGQUUTT5gA5JfAwkYxSnibNsYNle5qMfThfVYMZNEZaqxoeM7345/ucv5kHGAIy
SkK+r0ZaGIVKxJ5j2pyMkLbhez1plhUprbem9BUvvj8jZdEpn4NT5U6kgAFTigNKxNft7pXFciqS
YRI5vPuOcnxgsAk5KcoPN2CE3UMQemmaKuXotYW3VanYnW3xshxUA2YPKHTylTPdATiMbyg6ZBfz
UeOtC+v/Ywb7IPZBVmdi92Q10sqxp6ANw4mbkRWA/riJ4Blz5UCXtsz7qE4mdHiVmN8RvDJ3pEex
9pmy9iChyAmekBYRwgiL+9Hz6hmCXwQ5xuL00GXQ3DMeY1A8ro9jBcJ623vncO279cS64h5y+ZWA
UpxG9HVI/UslwXwgufl+Uf80+Di/JwXTx8Ck9lgZ15OyxaKlQqZuUAWWCB/bAV6B725A1QSG3PZx
fI/pDN1Ny809PHRIY6T2144vyz4c9xbNy11r9H7h6a4Do93cMzkzFyuPtUrCtBpgU1UZLH9JBdHY
8H/7Z/hqNQu663b2QV1XDDwWb6bcIX2KAiXLyqK6Fro1YMnSFX+RrqYZzEN5oOMfIUVfSj2e1VPP
4j9mCU/5KfX7qkEnXqM0M3qTI0OJR+JHb4CqGRGQAzVoSjWKsi+2+Umu/Niyo+SSWjYMGMZjYwtX
SPKqj/VbHBg8u3tVg9LX/mEzG28ZhYV8V3x59s0OF2nQApzQa4RfD0S5r/le4KTtz0TpyMEIjmpx
Zdar23s6RUou7Vbef0XpAxHVHOnTj7TAElja34NjGdqrr6KEGFw38zD1UFEjbu3sFqDnoO/xLQn0
NftlvCaXIg0Af4enQafXrimKwTkZf1oz8w/6ikrAyDUfb/01gj53lXIAGoW/xrphIijD7Hy7Z37b
Lc6SPWohYE70emIKnIhhOUJpJi+xNlfvX7Zwu9Infr5kJ+oubTf+kNsNDQEjFgyC+1/TSU7UoZ3X
aoCLIuwP4xc4ti9SK40MCBAB17KywUy1Z5dz0Z0cpW1LkmZXBWaO/pR0BlJ0imHwS8EiIIr79sHN
JEbfImg+TBePPb+/R4pSjo/0fJB+ARTCTLqtSv+X6x9RE5JKEVrOaoEHHo0cHfiE9+gRLj2qKLdM
BkMXwUiP+K0VfvggluTDxzJGtm3V17l241dtuGVxeu8BoBE4u5Z41nrn/NDid6sh3UzzoSwP14D6
VLQXj6HmAPqo5H+cfhGYV2bYfNzi5cNnCCrotqDxaiaChB9U+IdEbK89bsgmf8z+qPYj+r7spoPI
wfDKpu5UeudXgyEdWYj9L6lft+eZEZNy2LBITuYNyyI+6wFuIbVn7kiUilPzzUqg794WiswGjUsQ
DOAuixO3aa9P9BZZpNMMvFpc6fxc3UfkAWo92OlQYPfekkkihkZsWtqjG92toFJ0VdyTIDNwV23x
8p6wgR+jufGnFQOv3jYMpHQkgidiqyB1rwDwokQRsPTuDv5zQVsTvFxa20NQUJx5XClu087keB2o
g8k06Lx8+CbF4hv6+HP/A7d+gFLR9TsFUBYVyELlAqwwjPQTeVTJOPWdF/B0dZ5mbp0vofKmhV+b
BUh2bTp8eG+GjkrTSg9TufNI71TLBXsqp0A2xovbk64OnNjlkSnHmwYTASpYLHremNXpkq6nbi0w
v5l5QOU7Rh5ho4nB4LAdGFxypvJWNY+CO2BvRYetnHSs+GrCtWmLFsuuNbE3RMyDFRmvW+OoRqIG
njjf31Dp/7lXAUvUdaa9OniRPiVSdjezeLvjwl0HJjvUYi1cWu4Wj/JEBdYS+u/hmzrqnO7j82Tf
TwZXA4L75+U+gi4nWCrYZkkcZJwqMfPpTlJhiQpBvp2EdPWTDqF5P1qxz8qvpf6TCCn6RaPcAck4
3MJvP/doKw0lZuPjEAu/gx1oawgTH1PCqMcfcUGQUILmmXs4Bpu6nfVxHQDC1KMamRFCUM6CZQgM
PewKHSIFDHcrvVahkHlKYpmTy7mmB61Akizew5GyQ6ugCU/6gu7giJhoHVG6h8kPODxFudXNdj4w
AjQRNrRw9N2jIqA6rmeudWmJri6T8tJ/AGeMfRPQxTaJ5XyudNNvt0mD54z+tZVIdEnU91fMyCjb
/SOy3HejN0VsZ8oa7RCCu6WTDOH/t3ydRrzqoVf1MpwTiNWSGf1hAMcJ4xCp/5S3EkxBBiQPaEti
IC1atMvIq087ZSKUQdDfRuU6wYQUBKbl/AkncPToRTKFsbCz8dJ4nkOYEKbauv98OhSHRyr9VJ0k
2SZx4y+v4FrzGtRJ7XGpWs20rwIPxA/fnby58ScntXZ0ioff6lLNk39AwbhxzIANXfGSh0FKUvxk
UIiUz1TgkFdE08BBUEV4ioACEzSUlbbqR8/N5Ku1R2RBWF/fNvnwmFm+dU+iT+svUzKk+Zzqd528
IxTvB7O/mLbAY7j7XqpWrS6zPeMzlCe+qp+V1iN/q2I3ciMqSF8MOg2yyUBGTt9E+LXG68cdggRk
t1jUD6PqxYME3U7OixLP2Kemy5pXJNbDv3GcS24EbJMh64DS4GFNPywZ8A+Opwf84XcNswoORhVb
mlBUWXd9ksW1pp+vdAKMIvb2AeZ5be4VimHynxf0phwgNyJAcsEA/WH9YLuuCFuprf4n3I0F7GdC
qWU9kR7AhLyP31sc2KROPgxHBPXCy6YaUUjr5e8600DJEx43suMD56+2/A3iS545EJnZTa+3DgHx
/DucjPTRTH+HGpr/OdSv4wF/S2i0CTC2WVcGGtAQBoB7F2Fm6EA/qAP18obs8odoiuG9+novOlds
S5fv+xqDyZ8gYtZ8+rxY9cEtre6kPEIRzUi9+5Z3Fq6kBR4rI+9Z5wgKaaoImMPpzABGWwuFHq4F
mN4qe4JqJmmC2gknI/FVjnWcP2PeuejpTPDcItaG/zBRMz26zYowVOx4wH/FnRtGiRFoxCmSL3er
jtrQueIMycPE4Lnoio/l/oW9UU3XCpAc3xH/XOHYKM2I9tZa5acVcQsewkB9JdPgWAbwFTm7xgAO
Q5yOqv1cIWxQ1wqysXbtLQaapQJHE41lqkx/bdO/6L/+e7/03gWSiQ9QLIxBBi0UbhQVIF6mkrmM
9FYMYEXXUu0ptKLJkjYkNS7uCcDhxSnbOGmlsssQ4gJFAxFbsPU7ftHTlJZpLhR7+r08jFtrOILZ
2O4psRHw0/u5ePxRWDi+oi7mesLmFj0G/gGsnxSqB8uU1EgQloQFMtvTN6DCZyU/MiNhchVU9oJV
kgIRNDEtdVTOCaNSjdA+2HLZ2oS6gpY96ZxMsLb5ylwT0WMafOprYOuVU2nY6xv2dfTkRTrzUNPe
gojTmoGPbm8RqFEjdJ2c6Cqow5lxppbXgs3YcXcz8ZRIt5BecWR/UqAvHXkMPhm+bGMRk0A+RmCt
9mrNyzN1DFdNnZoejRdNf6aGCr4x7l1FqhDx5cYg2bXPn1ymaaPR49mOwUtw+Dew5hRZZxZXJmIz
IYu2SROSY23gDe9dJ2OMcb7Blf7dGJ2GC0zRR9MpJB/claqI2VTue9XZpStcc4xSbInNPwqde3b8
pb7/zBnGLbwh6tXD5dquioCLumHBjD29W66ryG7xjVBMekz72C5wTgCSw/Vhz7NxWMWMVKya5CEq
IcLiB2whhS1HlpyDzHEfcki9qI32RP54Gh3YVyvPyxwLmPZaxfFM2pV1rSynbHBCWMDcqRlTsRkF
u0hFYs01zbcUJsE+3XKRcLZ2jOdR5wJ7c97mWwRedkpX3l/WcLDpLx2h4gbJNZE6ijzajVusp9JJ
y/bpilNHSBI7TNTrOTIP2mxcCg67HZ8BZMQdN95x792WaQI90SqYwHIrF4yIuPSbJ3YyKgLqNEX6
C8jyPocHTE9rsLZfzyGdUEqgyrGkxO9ittBVknj81bfXXCXkHI2RjKw0yUdWYtSL7XhRjec7ywuk
VGwBVz3MDnY3PXWr+N9IxRHeLNuGYk1XRaQFTze3DSci/7iywa6KqVm197joZUlrp/b74dkeZF8m
i4iPll0MWWF74ntIoW7rC50dJchCxmYm4V2zW0pQ9M8Ejj10XHUE+u5PzLu8wcgWJme1kDq/62CZ
HkWTk7JBBMmku2OhNiE67gYgi3Je3xAKreUU8axR/0x94JSS66WtjNWMnwhnbOMdaqQIjsFoAUSx
mE8r3sM7Z4OH23Zm18Frbvkk7nQ9PRTm8ktlhKb0ul3Rh0nNTApaMjuJlvqrjxxKrjr6Prr/YDa9
g/sydrdbd6TAaHPNwVAuyNMbQp8lkKaQKzi/QG2rtqbD2aDrDmX+yXVH9HdsD1EGa+6JsPs/XkGZ
iZeIrcHtvAABibvj14Vdbv8Cu7ByC55EeRn9J1b26lyjU0Rf2O9xBDxrVlvTjd4niOiFp/BCxL4i
3sBAmHJJ73qTwjU0JTuSV3s6jW2oZlssPlrL41Zwju9nNQMsqPbrUTk3doFcO4UE1YIwTWM3yL7S
if+QNVaFken7b/AOohY4bzPc1KfqJsbDHTMNQ43Nwqj3zCcrlSU/6oSDvA7Dq8/9/RbwSNKZXtcc
rsRRRzhSQXbZYCv2y3KB3kXPWGzY7HAxZbZHiWfLbLS3pWUJBTX+v4yMXnr9U+xuxWq3Hvs44BYZ
zk5lnXn6UYKjdY11746tnkUemKyXmfGqgbe3atkWcbsrO2z2gPbFPLQ1UU4uFfBD56zQV4x265sP
57eM0HOts2rFPd4WP1TXF+BwYGUPgZsBFVumnraeFu8jJDXIZlYJddzuPMcaUYthUldHcZArOc0z
tu/Jf0bYlIFGBdE0y3BA96ENGtBNbR3YI6jraGJvpJt7otx8P1L1/IBu4In+jruOclAdqBZFaIHT
FJrBXMmJLer+m3bkCQz3vof0u7h83BAmrhQnLkCiBBy3eGLRv/O2czjPbX8SFE7oDh1l75NpUESv
IMWjPfnjP7pTOYbl4oo2++kIR0t/qcbhTLdCML/QWEtu//OzcUmrgbAKMbo4/IZBiQtPtgEv/w6m
WpUSzPByqMwQKYPaxF3H2tz1O2e2Uet3XpDDsP72m7OvCZ24zjGWnNk9JikeFhiJCAK3zxBJ5kxq
9HdRUama2MUW5bulvDgCJjbq4xWDuMNmjci2iVgH+5rAYs3Aq49b6p+FGq/E1NnsbTWd6SnI9juW
DhxS4HAgwde5yqw4QpkZoUBAL7ptjcqlwOpD2xnWFoMxLJLHdH/W8jV6HSz0T29ll3BINzrOPD+I
6PfYbykwLr+yC5o7UVqmjtu9cEdw76+aEqJhJx6Iym3ah746vxssTTGFqUfonwp6sAp9IZWCbz+m
1NV42CBQkT1r5sSZPZ6MlPgUxuLTniA+z6xze9enVfDM9Lf3wNIOs9/WxaEHvWGJpyddyCMi9GHy
FehXBfHAhEGE2qWT3YR+fA+yHrsRc3cOf1sQ/ggPcomvbJbPy/StG8g4rJVIcofRajzjUtNIayuA
6/cGnRTM6LADhLeXS0TRjDJPDxI3Cgb06LHvf6BIEUq20uHa/BTl0FfeWwPoZceAiHkAZr6fJqk/
6aO7zs8IRgQ+pr5NXV4Am51TzY0s01k/FWzog+NAGp7Q6C1TfpztwRfVchqjCtIFPtPuzPUJL+lw
kp/NLHrgyxypEv6UvoeLOcnS4uEGPJmC5MTEj/vCy57DpuePrreI5OxeHfnHn46TT1Y5HTpofSg+
93ze9Iko64oGtrEGCuywJ1VqYOExZQjZizMrcwO0a9M0KMSdeROHr5iRn6AQZj4CWH7xmbMc6vOD
xQqrd19qoMYoIVSjJQ8t7kmoYu3L3YhVox5TJVti/3WM+aZ2hWUxOcOg40tXhAxj5x37V1hu+Qft
z1nssKHusF0hNCXDfJtsTO8C0+zN3efAtXd0o7Asc2ZvskPi6L9J5iVrR7t0tts15oggxbeNWAo0
WHSsHYgK0r6eorhkprUlKltJBbm6eNCveyiMGB/N0m9cg6CLM97cG02GdnbrVpWHtcIs+8eLbS0B
/jy2VtPT5twt4CiN/RhS3yrmGDs9EI+6GzibYWrzuM26Rq11kDdxSGbMDTVNdnC/axScAvVycYK+
xrMDvuH1JqkkzykKT8Um8Y46i+ElBvsEc0Sbjj1EvVKWVAYycQ4ynskVDqz7L35fYXqnWOVT2Ajv
kUDMnVN6xtaFP3DIHBzep6XJJSsZvUzO7ej8ihjnvjE7gDPG0xkrPgrfsAzBAGM955hLVCSmJ9lu
K2qNJmIXpyjuWaZZnrowEuV5RuqnvEu8ngohs4MP5O8CV/fGJXYoP6GpGwIsvmloMfqP2lOlYJEx
QMGo+ytv5BXtA26Ru5bfyVZPm3KTtujIB8r+CE/q9C58tg1Cn3jR1LPGzqK1IRmwtauVKv6BM6ow
w1h2Jv/wEBsoKt8N5eZK1Ec36HuMQ+zmMKt8VSC+y6iDyzys7zqc2seU9DqYlUFd7w+pauZmttT5
K/j+aZTwKzhx3VWwzZjNmmXlG3+A8Fye3oo77igENrXR8lX9jXD+6ngTziy2WHq7RfpWhl8LbHPP
WYgofqxPEIGtbs9F5FRwf9QERMgs+hwL9E55KabUESswiPZijkIgftgzp+l3RyRQ617Uk9PcwMia
VLOvRODQK7ctuwcTzeFBu5I/4qlnV1h4Rlwpyxz4PFUQ0jinXk5LuY7argSMK4yMajQjqjm2l7Q7
fw0FZlhhlDlPjtQLJLStHBwbxrom6jpFjQJNuSzPYyJj1g0+D4F/GpC1OyOZLhINm0eru/oCUZJP
UFqz3MBegfzUUI/xvltklflCZm3gAYo9BRYBqYU0viPB1JVwxQvD3BdX7qCVRnAwJxeLt8gV9UJw
1t8vmPArz3g4bVPRxB0QpA3JW5A69M6ow3BHsnTdUiTYKafsIw2OIa9TjCEgJ73lznfcyjsCJMDo
fk4wG2NHTXxo6H4cj96YuRZ1o0M2usX5v8L1o0uPL3TcXZCd5mj7ZefbV6n9SFnEoA1GCsWEw0Sm
yzYq3SzUPfXK3Hq5bJnA30ctBJVew/mGbx/i3FKI9T1gE6Hor3gyNw6LaJQE/VGYtMsg3/mIBptq
+9FkIoce4Bp6RElN3WKWOH37fyPQ3Ghgko/vKBTxDaiOnyE4K2xbI/b6tF5HSV9O4NpMzrRELdCW
Cb3gipwp3Gwneqqp2BA1obwvxdYXltGcn/umRoHJ5MV5bwNnn2w7WKNzZZg9kcWerOT7p1e/Cz4+
hXqNHGrm0KEedJCAWFKCp8QDy47OekvtAB7s1n+MFbOjWE0zf94rgp4SJOFEGaCx/B9k4/9Ao88V
UHRzKZ800JfkEKmRuKA+11+9f7CNMAF4Q3qKGyQYNLvGliUUliipbVWU98FZcnYq906hqxp6SXT3
lxe58oiW23ajsq8OJwhhdSjUwEBNrgMSX9hlhoYmJx44Sq49WhYAN6l1y28tUVYZzudAmdeh/E7V
D+tTrXoqaKSu+7GdGXhgkLJis+cdD8qbangfD0l1UrQOj/pci/UJ7gw72TFbBHjNz5rFtwgBQaMa
a7Wc7KIjqbNVZ59lheJtyiNYmkp1x8f1cBCzohWSz2zWVXbdfMhzdQGJI0QosVsZ9tFp8S+3Z/Mz
+JDU6V5lM3ob84xlqhbmCL+wsT5CrN9Rv5qMDLwf5jQXqS2bMjTzsQ35bpA3uX+l9/18kIgrAr78
8eDssMrDj0YnGH96wJn2Ojtru24EzAPp+SsJVLDWYmPP9jBmNnZqDZvgL1TrfqC7YOQtUfAODR9b
nNagc1XU0Bc8J/fiQGmzoCab9xVN7OQRxXClSImBUdQUtEKj3KcxzdAOb7E2bWW9SJICVge+Ahbh
tJmJGHXBGmDkmNMAgzDC6h9qPVT+0n90Qvx8yn4/HvOKksslG2vP1Zari2RJX4KUsoDtLMpLTDH6
a0np6GxHGOSswWuVS2UgdaE8BFFJnAV+89PRKLsAOBgIFxiCIgzJkxo3n3hOILVsSpPp0IjSaXcl
YpypybgjTcGHCXYG9yzw+Q3nm+z47D80FgGc/Brg5LIlIATeFu+4AFTv3wYlLuoqyS2u61zb65Mx
UuaLUF7zo8ikgLC+sy6C6Tj9Yg+PeFKGK9IR1IjrzD3pQ+nrhSZ9kFHZjCz79Fgmqg+eVQ6mlcQ/
fepJKLsif1DI83GXMkg8qNzn9+ORQPDRvVKA4G+4SuILF2gSmXnAX8uI7ldPmW0drBQBU8u89V3C
CSWH/kEEUHHsiGzYXLajnSrgevzSxFzpJU0/oa3BLoCWeQQ5mwrEotuTp2k0bs+xe2Q5K49z7M73
yJsEYaenn6oeTbBFhVj8/2WxSS1JZxksLYdhaT0nYpkhttWcLi5C7xWbXIrYRrFwebBoZhm7RTTZ
jZjbSNGaC0uCl9jKMlt7fYhSYocb16Q73B7OvlDoiqk0cBedvNW1vvCpb1yPkd9PoqvZsjulvfZS
sFjb7jMSI2XX4uhTXrWMzMJ+2VtQGhVW15PLtC6+ah7LEun9Cj4dbfYR5odQOyQaHVvlhbIzac7u
N94N3PBhh3fBuJXEy39R6EDbdcaFzz2S4xOKUbO2naxMkzX5p5T4Jg2FJHGQl74IpfgQOp2u8tLh
Wt1r2mw2e2yd5s23z1QkDNBm8NrIdZ7n7++X/lk2Y3VK+Wwx/8Q/rr71IqDTGUL0I3K7lqhZfebD
qUU9RaMUI+3FFZFSs3PYX5yGwKIZS1mMIvTfJbO4eoj4VTjnlo5PPZC/xuD2qMCbZtloX7e0bjrS
bTZIZZX+Echf/3vStE6S1BVKBYQe84t+0g1GToONoBUZ710DZ3eWiIsrk/AJQY5IbHVcyYfmuF8u
Q9KCMZm2yV8pLKQ4tm9x9/6/zmrgaA3/fTTPpNwk/rl5LcGt1bEruxvTMH3wi91MpXH1tn+aq/CV
Sx2fm3tmOLvH7npnNnb8qPh1pdyLrCgMPIQwK8y0ziKnpsvYGc/fUuNLVtyDewTbq94r4pdHX5sO
GkIbcVOBanm4khKV86cY2NJXWOscYIfnCo1M5aptOExBSywSK1bKFl2xPlGuFt5OIfilnq9eyXkG
mZGHh3eYtGKkxCxtWZREiRhB17iNnrQZdxOQB3eSly7bZG8GLInsydciWuwrPoV/sgS31hudgwY1
9xJm/sXW6tRlqXL2V90Aqa7WSB15llFWTsgZ2I5WZ/TArG0J5TNiNDTpg09U1QrIPTsfq0/Z6MLP
K4aTVTor/8BGv61FpX2+OcHh0pLYg6BVMWLdkK/xfX6wFFSxqrTSaN0csu8pemCwxw1qeeVUO3jv
J6TJptjVNzlwd16QVS7S8gVv3Xc7xHrR3TdaL0GGUKyBDIbUcIRK8VA+ajVyLwmJySvGH4Zz927p
RIVi9tyd0RIQxMUdfru6fdTeQvN3x4r2K02R5cGLxR0GMUsRlAE3jE9erFF8o85iGEJibqNDTfFD
yC2EENIk1AF1a9UCo9AvdM+XQ8SQVgfZDarU1tFC/PEs4EfWloXTw70PM6Id1npJ/t6piRqBsS97
NRGjoEgtKYOW1JmhfTSvVSYNwKM6joBrABaQH+EnRod2+OZGjtH5elPKKZHa8t1GKbxOjFROGp44
jlncZ7lv2pk+Y9ZzaSrTPuBxr7DMPZgBHhydzdP5XTMmp2pLtb3dyVUzvrFms+HGDbc7jeuqiCmW
DDeU1Pt3hsGyuXyPhs+pP0tUaXySe/IGDUGFf+2eE/9X+KJzcaNxg49rnpqoO1f8hcrhXVztlMfa
G8XrXAqq9lWEedYUh+BA7W+sQ/REYdkXDhcyojFtAZ0o0z7vkh/NF43GVtJW9qEdU2ubE8rWTnim
xCRhfbjzKak2tkSvNoCCQEllafCsVXi7hXNZfIhdOsR8zmpdtQfR8aENXiIOX0tgvrbzN6MdsQoD
iZbK5d5wipVKuIINCF0zzTSfUa04t5NJq48U+jb1NEmcotKyevNY9YEiuKjqXDie9HHBwYY7tAnG
LlhHIymfQWeO5FGwA5r2KyhcoWxuEuTamX+Vryrg5/V8vtDPNhONXvowB3CVn4MYwKMNIDFVi1Nu
WoGjminkaEo4vDZm1+kfE9hHVGlv7xB7GvrY0ahvfjHC+C1fob5WUF473eRaYH1Ifq2nwZvdLDnP
tiu/gH2EHm2fnXHdyppjNnQYHXYfPaECYbxMVnPPNB4PdTRiLbFdA9eZTqt88b1gWXg2maKI9vVo
xr3om+PzVNf2HsS1lqZkWB8mVly3CCQpVqSBhj0m+WJL7M5aAx3dF66H4wBdZXYjFCKS1LBULWLc
b1bDGupKGGtw+Yc8yKFVdLKuHRoUMqmlEjU7I+m0Hpt4PLfKB1Pmc3OSYuq3qhPBhA7JuG94b4nq
Lm9pWp6+GtcjezyK26wqx+KYa5EmmARbpa6ANDULz0PsBepBcEJuZGXh1nskd7K0cLdMtPDZV3Ha
diN1JrB7EnwR4O98QRwLe7agELs3pT7s8HG3st4IlvNnp8ZQk8vNauiU1LgglS5WnD0kU9Eif2ce
aeZCKbYdsAShdFdl+ClcA8gcsqbw7jFzhv1Ps+CWtXNwCSPTBMuSEs8MLD8GIFbR/IF3BYY1ihfZ
KknIC/SLmWSXfNP/cMOZ0lnWVZLgdamh+3eG4loPIbS3MDQOSdCSgaM3/IyNri9atPm4W5Qp9RPh
1oyRQYOEPHYjL3SehZkIocX4Ew1yTBy1WNd+iakjnYSpsHdWDgl+Wq6v/VL2SDAfZrR1WkRO2Wxb
SeNoaRaRijO9330yk6Rn6W3AsHw68iTzBdo9mdjBOo88ChUR4sch6Jzhxe9ucGGnzY6trhHFPzGt
sf4rXrfO3m1XJp2U8yDXANeEza+8miDLvah6L4C7cvwR1HneXFlKW326dFcBtKk5S7PFyzx22Nso
uxSSvi/V8b2+bR5gp36byu9FXCY4gqyvPvqH+x5h5Y3ByFXpwcKtynt5pVn3X26eOK1TQiOPntae
2JLwl7tULWZj6Zx3KoFjBLrY01PEYpOxcjgwSnuzCbCJtvjnIl+7W75ihcqOmhmRYZ8eIN6Xpm+m
4zgBjSA42GOIBWntNgyGIkfVMJtJPRl9004Po43pZ8GakJmgAS3XFnFZ7uqv9yeUv03LL2YsrOrN
zWP5Zcfivwo5c0qbmrv1jTSifpBE+NV/0nFDshKOZ7kD7ClgpfTXOC0yUwEVhD14Oy+oeECQ6QXr
1d5Z4iENDM9DyU2i02WPd3r6+Mv7/yLYhrQoVfXQJRi7qfzIU99iRZLojqIHlXGM4p9qOKp1duFB
yF3MF+PIPyEz7nXojgeCjA4dLLBRUBibYSHrIVaYIkRSGBoLzVSEMeaafW1iGRADWhBwAllY+mGI
bld9eJH37JcdDs8De+niGWGztm/UPR0dSF0SeX8afP3AP8X1E50XRvnwq33ABbyPgjc9Uuh3X7nn
UQ7o1usJcH092VoDKoPhyNeNY2KzgzwmR6K91KosTp/b414RBEyZNTlsOvv6S63v9T3tohVRQVj9
sMNQ/ONYOGw0JAMzzFQBMpXPch1G0Z1Wex40yDQ8FrKIXL/eZeggGTpLZ8b1h8/6FaanSW7nTXvg
QLsX9cxYCX2CQOChY58nrKl9OlojFnm+JmTcWEOvsH2nh364nqWC6kvw9Iw6Egj05OSHM8Dz+Y/5
msGLcl+YMfJWCrBO/ekXL+rGqHrJBjhAZPQ31IsYTF4JOYABScpthZ7FrpZ/18bjMZKH2c/yO2EM
ft1i+bg+GO04cqIaihYBgZ9tRUTRo9ZJITqdPUtodi1Tp54S9FK08vY73FLOACGmjxkfc/j+sd4l
XuNeyTTc1i11WTAYbjaud8aA/EHV+Up1AeutqAqHp6WmFsenRRxDVyz9nB2Jx+4ImBtvP8OH/QWE
drEbc3LCjtKak0ghCMaviNEStdpZV39qd6iHeK262aH+xmDjA5FRf7rmmv2hgLx1y+FiBTJQhNFU
/uvhEBjyZSgaDOc68X6rQMSmU9hOSVYjBiE5+oaHjbJ/QHVzy9SOUUAvYiqQ+c7Jy8fDunp8izIh
XZ9874tK0V2gqgcK0mwDBoHNimJaGq6UfRwLdCPfzRCvtgjDaISaQPr6fXkrCHOFbnEAowjRW1OU
C9a5o6/zktyyTrWKs5/D12WRf6xiJRr5NKgE2n8d64ZSkXcDkgIBmhXAS/CTAiMcaO2yweIitGVn
BI2vWMjB4UrBy9Vc6dszKKG+59zZ1AEXiiefmPUZp6M1q85vt8zPHbhpzvEaQ2IJU3nVRFoQuAvE
9MTZvc54PTu+F/pIPXwTH5We3f7EF8RKKtmv1+xU5lGxV3bwLmAwcQ2w4VU53YiRPEkxfjY24p3S
BnuPzWP20f2FJEfz+XvMF/eT5WYER/HlTL7Y16Yjpr4hpc26Vmk/puCCBsdAPIDB2mmjgVDAmWg2
Kn0/dIdTBt+Ij/6PWWsroHFLt4sLoxW29gQR6ywkHJ0VrRlWk6+nrpuuoYE5Tm3Yisnpf8V7cEqG
w1wUCFer9RvuF8sd8qGMSo6ObXmdOuDZ3C2Ikfvt23PZLHpJqaD9Q20E2C8WmAloLIgO2nrFvGdf
C1fo99jHeuB9E7FCL9CwfUBsF0cXgk/q/ZcTXREYrYmnLqTqNPjNV7LK+N1fniHX7WGYaXw1Mdsk
1vAbFaG4FMi9t69oAjrsbj+d+KPc0a53OMb5nt/m/iPY3Pzpwm88RS09lY0JrRed0MgmjzILAesg
n379UgiA3xHDk1pKE9O+IXZRTpVbwpz7ij8b9QtGAv2Ww4hk4LgxdIAfmhh+aPMfR02AMb0BoenD
bhOHULQpJN3+hgzQVRcnSIxsut3Ox0qt/bTSK19WpbN+Z4LEcKs8Cdpg2NrnA0yMx56ON6O3gnJv
fyZ8KaXzWf6cmG7KDLiuJPAmulS19/IRhZKmPEkm3bRFYuzDZYkFTtvP3lGbb+Dndjng4idPAhfH
kgWJYnJgG6e//RxlGBtksJsubjOhntp6Vo4AUnGkX1Zg/VxvelHvAaGWcxEGQqm0luqtm0FTC98+
6E/74tIcjhTa86b2xxYmD8qqKNOJm9XEQODS1wgaT01np5UKnshlYa4TLPzmweP2+vsI0dB5Ma2g
Ii3HrH633x0femUE4+v7bFXP3Ji4njb4hq3Sf7uiwf8L+JHBbqKyqN4F61Dsk35SODOftJyZP/k5
Xfek9h1GYP3IZaRJdzKb9phZqxSpXNCm3Wt2ddP5OUVkKsMQffsfz0fVmz5fyUJbg2IkZedqiqAw
VExvkTNY0LZwG2M3+xUatx0SDWocORZvBeXgvRke3DkiMjPuYznaz7OiJK7XV+arOSNHX8s602SI
qjevUW/eNgEAN+Qvc7KsQofHzKBL30kgmeogmAap19dUsjxcFTJIfHdmCV3uohiZBoEzIEhSR7n8
hHt81K4pS/8M2f8VhPl/18WhVKjOzU5kDxt5PKqOOCmNdu6fuRvQD11EF1TMHYduGzw4Dn9blQhL
Wcv6eK5iHamyuJ8MADcd0XUELaagnEKBDa9nt9nuExahYExb01W6sPV3JSLinx2SXcBJYkQEFv9k
AaG3LwFPAZiCsRHT6KHO0ay4CDipTDJJMKv0qk1otz3rTcY7qzkR6Kobsj2+lE0j5mjWsPXrrfGK
Y59GHfHvMTP/f+zjDYLNtzb/7Wx3b2SlKfXm3Vp+bkjHUMTSYl39gGEo7CtJkqBD+nE7+4JXJOm4
kQWINtd/GltMDUZUbHJ7wOwdYcsr6LtOElQJhTqS7wc/aYdwr5RSbimPNb3gWlfFOo5uZKwbPtEl
dKLx4gbcRoo5dy5zjQp7RiFLMd9BtwjG1Cpvcax2pDPaY5c5IqX6SWBvRFk1eYr3pa3twtygtroV
a6ahtetgwufmbpKt0QxvHBGppGxwwcUT13pMno6UfycS1wraGMcqeNnekWRNvDBIoi5UM/xrbJRy
3A+ryKVyq+htg5e3NKpnzTyBlv9UBD9NpAztNqw/xSMThg7jOMe48++hi55nUyWw8dxva7jaaFt3
D9tU/Ln2iNie3XNdBzc8MPSskrkHLPG6PTPOm18E6ICjtPESSk4be3vNx0c2504n3BvSEwW9KoTz
/7AwZSwkaIi5ptoZih6ckWHd+nphbLPb7f7sM5/vtruNKyga+vox+IIRcdqzBSpZgomrFMnZk9Ds
8oXd6IBM62Eeh+9brg5GzkVGSvZS8ToGgTbcQlaXOd4aHRVI8HzWHHOafrG10vAVqYnoExRLIRA7
MHpuaZs78inlkpxQ0M/jVQryl9tzXn8Y4KQpv3/fTeDA655t13S5wBYdLuMOUjUbtlzOvlRSr6TB
ai8Bz4NaVVw5ysQEpoRC4lCmNXq7x+QjXXfjsxAFAmZV9IzCIsHp5lST13XXz/kN1RjWiC6pGZps
YHUEqiFXlqSs/x2TZbEUwU0bVGDew4eyAYrGADzhTG952bC03tayrQrCryJcwa4B1Fvr4qVmGtit
fp5yNVtPQwNDP9iOgezRFuw5uIHd0aATLZPbBvWZib//El7Tcv3PJGOuBmoHDh6YrSNQ6VVs5Xma
SfUPoKiJ0x5vEpzNHKuBjDs+82Qr2lJDWcVq2Pnp8X44qEVXOHlRqC0MTV8fS+BIxvd+1xAks4ts
kdVoJCFRdbJerk7XHDK3lK9LypejtQ2U6VBeQuhWhM3Z6b3GC0A8JYH1wTHDonq3DzWtibMCYEkJ
Uj3q69xlYw9ejur8xnmGuKFjaA9IAuQMo+ILQDSs5aA9L3uhq0xd6tRvTC9iUlCnGF4c06zwmSnM
DcQn3b2EH2Wqgan6tUsrFkknAPaCI3emM038lhjz9SOWNwZ8FrR4W7qfQFQ14eKriI4NmfLrfgqf
E2hTkZZcuNnnyhoqHyDzcHjDkArvADqsqe4QfnBfwc4+Eu+Z25yKzVx5wbdeyP5/vTV7LnouNpNF
zkX++LKxnL/Mbl70DfQxWnioaPwGu5do9lF1mo8WSAtYAdRE2O7pcoeMvEXkXft5dC2k/AAkcRk8
d/vbJtaU3eZP4174cHmOK+gae9T66VV3SNMgf/gjDC5sCVq88nzf/Zeh/lql5vm9F99rPZKBw98K
2TgOepPnh7kReNpZKiGEJxmcaREccKvZYm9cqFcaqyKE8wLOucB4b43dpkC/TD0I0ih8bgihdKB2
mHjJPjwkKpLuzjnZwV6NpTqX64wH4lKUQePVs5GqLUUIJrQq0Tn+81CmxgV6gfAOcZSXROFSgYj7
gkeDM44YuuQj+ETFO5NrK29c61R7oCZsTNLe6RnFovSoobcDL5rLFx9sa88n+P8vfLuNXaeOyRHd
Qw6f9ltqWHZABwApztPK3Z7lhhXJNmWTCP9F+18ektFvAnJaRa1cbn9k1fzjgG9DFjvXgPIw06us
fwQlrX3OfpCMUrkuCZaz5m29flcJk83SgaF+pZ7I+wimWqJY37gC2NXP7bsxiFndzSu/d1JmVGes
8+yu3BUGf5timn68UKtc4MMLw6jjsp4HYOUqR01sQwib7MRkbH76UyhixL10zDnNvNzoDAgJx6MC
zuBOTLOxUOdL35VGzO7J2bagh6OmJ8IplpJYQm54gaV203rfWzBeJWDnMZssAB/jXCPrYRxIXzrg
/XfqhnAjAg4Dxf9XY7rHYxOHHZk1XsW7iiqe4ppG0BNXQQpXhn09oRpN1v5onmjzbozFe4eDx1FS
v21AgG5kH2GGNqXMNioNzeT8uUlw/g5QBp4rlPbS3wJ9RLl9KVDbRc+acYwh8PXhS4N9WTlpiT0p
V9cKnSVDXdbmBMescz6bSqz//6aZ9MF0DXuK8RDItqq1eOewuM1Lhdd1Or0+3W3AP4RFTFvF8F0d
MZC4I6I/h/TrgmZigeMwdlOv+0dsDfORbBMNAV4z22D1kbDr0A+lY+PKIsdTClPdFnK4QX+YPTAw
oog9LGyrmfm17ENwgaKNDDtmKsqKnvxAUFs/QxFDHwNvq18lAFZIQI8CnAsZatUQituU66ADMhut
U0RLHGk+3WAH3ulrKlea74YguOqfc5LJV1CJiRm65U9uRo72Krn+FUwuSGnhNbwP9HAT/7gKvbEs
QYc89UEFiyKjzUW14V7NVTFVFu+NEurTKfB8V0+V9tN0B04lfNuPL3hnKbO6MUbHnGgaHmhs+lDU
/l2t0YP052aongzyv+7fdk2IbNOsfR0k5LNSp0fdYV3m2boipAnZzhGb+QFZxHAzzqGROq1yYm6J
Stbi7NSgLMBZSvvg8+zJ2VeiHJC5Im5IiFZreU1hxLBKgJt10WgfDmwGi2mFYTgPVXU49WVOr/mS
sjVATFqV8bycjoxOjBS65MimcD/830+88CdZtpLQZtFb/4dYO5Cg2SAq0b0GnlaIldviTZhuv6qp
NbKLhi8M6Z96dQ+qTY8sVHDi2tUSS6dJBRTInM7q9hXHziqD8pqtc/ELmvhMrxc8UVO1RZfkvgEX
+G3VF6yxy5v5IrQ4zicAG67/6fwrJQ7TIBCxTbHNeO9Coixu8TlJch2q0De/u9f8Q9Uq0y3KhG+c
n8vTo6sHiCGdCX89TNaXjs9W4qh1Dv1e6uVRplcsZrVNqiMwFWv3zo4ImBGW7LAwJ97A14fuBZq3
PwkwyOAtViK7/r2ARJiheYpHTQcYNTJSpWR4856v8s4MCknFZ2x3Qpdy3KALxvTmJ9eFXBhJyfUs
Aenz7i14Q4ue9/5xl51hteB+shTfMoAngNt3O/8IUSFFzDxxXSQOYnWfyITWsI4uqFCB+KqTbq2i
bXJ/OJ/sNCTGR3XDYieMw5pHM5fbmMWk70cc1oEWIuT+3k8Q2uNTiA7xS2n2XttyJkC0G4GlIlRU
4+Pxszv1P0Dc6LQoLkQ0xW2mKdKmuvdH4g7LUvh0NgDTIoJ9KKB/+Ar40FQirmTC56jaz5wxuvfj
e3slKg+aR6NJxcgQ71iEurbI53IPB4X5bYyaH5O8AX5Vjpxa7mZ4ZrdHrcjamK4mra+WpxGV3sm/
Z0h+thbTHm5LPSRm+YovadTX5VL/v1vy/0FRb5ApBBVWU/yaFy4qnjmjLyPfWlPsLPZfk8j/Ft3U
lot8T7Ee2N9XLYfdCf5FDdG7FJgxBmLDo2N70Av+vfF62xZk1ZaU5R6vcKIj2ynXlFRRs82oIxv0
NgH0fKsBUj6jIoce6uQPLPARnfxa2IvQ0JOT5SO73PTAT78eNJiGZJTk0pCtoSG+BaQQ7FZEMQhY
FYdzHZohxDWLuelARkB+tV/GBYR1FmktfEGGm9LbMIcr+mFKak12FnZbqx91x11XttKXL6O3NpB1
LKsmmAoxr4iUFyh0hJtuzFL+E9p34lGpwZOcC/ed1A4hFsxxKnEo+ytdOai9uBQArIJ6cX6sIbB+
5aV3ynXE3lJ2Zrk30AS4z4Jho3e82hBDdNCUxpcbSgMD+shmiRapAVYWw8K9M6jGqfondeQGInMy
2CdLCtvEshqmgc2re/vsjHOXTKBLTyse6zwJ0AOQUOKyB4mowu+6pMJXFO6r/DV45fjWeOacJhZ7
qXA8MrpBLwVpretQOi+JLwiCYYj3H3RnoBrWJZjoQ2rb0hfk1t7yMMjKrfhv41pGRc3KBeuUYFL4
vwZzBLXi3jvd8jIWCPpwwQ9jmJZJl0vODmfqw5orQy67ZwukblIbfCQjQt8/mq/iOZkyuCW1G2ZT
cjLY6fWKwg6QNZGql5xNVL79nzFLGfRW+emwqdgMS2976awIhx0BTnluc9LnH4Alcoz4BDHUOxBz
4mBXMwZAsbc7rZ4Xi+0flWx4xml/5t6NqhPu/I6obcgd2CmNJc3E0NroxEvUsCQKVTW286u4Kigo
nZbCGmQHp1dFW+hCQLz8ACPi6vVTsmLTdr/WiwD+jD9XtrKDOgjq45K8Jjjf9LdAP4tFOGgRUpYc
ny8q4YywHyg/jGZFLVop/ozlcHTvrkAirq+E428Vnqow8eGj+sck21b4pEzm8tM+JKm5Uhi9mxlA
bHZAEayYPJ8C/evNWKadptf8gO7cN1Q8xX/1Qh7vwGlwKOiEgiXCvCJyL+otMQdeFwpVuS3W5RFy
CPSrmV8tzJuDm4PNvofvDs5rWXQAc127cSFcX5UQxHiwGs7UVvRu6gOE7iePpIo1HUnkqhtB0g62
Gr7HQOzYhFpVTxKRQjD52uCgvnZZE6fj5EeWGhib4uETd01i5lIGyuKiho0nbKqs5neAMe8a33Y8
kt3t7uDigf4DUoWPesqHoFJzdjduDfvcG39lPzFSZDK/JzAXFmjZ8hP4WGy92V7DhDCYnarWYP2A
e6lOR7fFBlggE/qjQKGo5kmd1waqv+B8nY6AA6X1veI1EX32Js4F0egY+JSrFE7venh4Cw6FLCgu
tnEuWN0d9GIiTWi0zKn2+O/0HlJjJrrKrZ0VqgMGhDsFn6JPIMC3wdJKsOpSePM3s62VpheuHHxP
qfRjGjQWkSP1T0m4tf1JPmo4c0GNVcP5tgKrCALSeSArFttJhbqQphVvgrqq5TgXIX3HvQ6mbYrm
/zh7mnliLshaDGR8aqavb8Edl45xOS2x+kPmkGPugccxpMHnQtn3OPhcJ86kCgarDSvD5KqKeHsy
LYy/YblFXBYElyN/Jue+jhcijZfjoDtSLoLpPYHgvNb8IxQ8q1FOPUfwwFThZw7/VpH+REtGECbW
XbVUsgqQ3MOFYtE0b6kToEuH8mwEWQs5IsE0affqXSU2BwCAOyZu/EFuTyMcbRIZBmB4yCBPfAqj
CJG/Y0PQNQVE3pqvfcAgEvtFsXMz2HMIqQTLC3UEzpLGv7/xOwRVRYUhfqo4JywpF/HgewiiWhhH
LXQUrrpwZi0/nIOqh/x5ZC1WJh2hW2g7tF9nYYkuaMgIYeezDAJWe+khCZAmnDqsA6ERSAlR4Vc3
fnBRyMg+EDBsgue7a2Ye032ET/gypFDQ4qxTTM5aJYBVngcf+tDS7VY6EMi8ftssaV0yePPJhguw
hVl1yFMhhIN7uI7bxDzVpdq2OwqZ47lBqCsWQN0kUZBwYhcEkmgqV/0RyTrLboCILcJyoruZS0YN
xIBOHGez+X8liXtDM5Smm+T2nXr7sizDJMVj7h/cFF0NLzdUSiOZ7tO1X/nNL0uUgWUvnGHUTfO8
cNknsKeNhQYfs7bPHvsiVdQvkK4HVqqdiXyJHpjwIXDXHJwc468Y8i7JR13LRt3YS6mLK8yGGYS5
/SO2gddAIyNJXnfaMpCJk7i8tpsJDOvNrHsUE95JV0CApXCd/To2su7Z7S8VO+ljnnByBkLt3EYF
c4t64HIPzxEfnHJeb6qxPeXRytvNvbAw6MaDH1O2yJDx0wPe59UspRD8I7//phxU72RcGBWweXkS
AF8xlpFjgVKb2ZkJiB4vHyJjHAdejx7E9/rDxlc6KZ/lblL8JJMMVx4sgSgBQFhMAyx2mbBNtcQH
FbinGUTBWxjxBD+O0X8EKs7QM3FvKvZqalaSU8lKYetwOk/Zl8dsLwauBlFfSR2KbexeQKGjv95R
kmELGmgAIAtKnHY+xtRnZxfRUwesloigXpbDRUrGP6EsbCHiPOHDYycmdZePobkEGdZ6aRDwK6S5
bQ4FgXKSQusqLyZmtU11Gcgsp8h/ZXOyGUm5JCCQYSR5Wwe5PdoGWHOsq5LkTj3v/gcgPgPN4Yoe
SmHBZvLqUVIUHmW0Yr2qXrO+BRDVstgrw7etzsMT1tsFx4Uid0XG9fc8KEZQnYH+u2jB8B4yiGjs
fYz/Ohbl2yInXtOHXq+UuQPJa/aK72zfjl/0MR7/+vJFsbTInAtVAGHAJcxpGA3tyCFXVwQ7+b+s
gjuNKC772GCNIb3w8DoUr3pzZZKTNyQ/YfB94WFCnRD5tirnw0TeDC3UVhWtMwJvaywrn3cM5fdc
o4F2LDsuttHM0PoR+G0prAe2WEE5mDs9pIM69BFIwqnYixHnw2TIx4CCzUZmtSH7ErWq4xh4T/6+
mfFu3fQq3PeIx+AUq74Sp+roafNv1Zd2GD8+6G0QsXH5HrWai141UmqyBz05vleB039gvAOT1tdn
ebmRKQLNGjUig/pJ6POmP7X7UfG5be6AYvq14GpWQGI425dH0Z6FEzniRV57v/yOglYo1DWKKfmC
cuGCen1CUNGIrxtRClvSHfPSo96kXPx6wGpgboOKNPoQ9vxtqfALHkjvPH2wR+SJXWauhjbocGm0
g1HeagNmrrpNstA/n6IYDSVvevUjPtCrMtVO0k+oj7dEd8xSfrptiKGuSp2ZeEY5HkDk+H1S/lsf
/6RXRncykw4Lq2g1odTGsEn8qx9l941ZDVpwBMcAropkCtSkH3HyW5OGky/kaWL8N2d/f9f/POC7
23Ee1RQwnmayHhPN2o0U+tqV4C6K5WR8dLWqhhsZYtjPeTdxcyvixMFRlbBDdeaVZxQtTcy6jlBH
74inRAKFC64hERZfnbwVbL5mkD0R09Q7/QIA7qqqJ09QwHWRc71vN9H8dV3TWL8idjcf/fMou94I
3PWAkTOHPLh+ZEypNz3pc8mSTtIUC/1itM8Q0zL0U51k9nY4Q61BKvwHi8KDIj4kwlNQZRO4GY/e
mec3umticxLBFZXpQeBxSwr1PYqLbfW/hmau7pDCnkC+7DgypZvlp8qVY/HHKZB/z3dpMTq10cL9
G6Y5Co1jvOzn0AH6slGFedkz+54w/5aKzJXT7YpZzAQO55S7lJ+BYXKdTDR2CT1fR2yO+UUN4nwy
0i/6yUe1C5sDtRINsysPfXES+Gi2t7VYLHAnyeGxShyI09b99UMu/AS8UFJ/ZTWdwcWhDlULwapP
gYalCc2v0uhHYRuergzk51pMrMj9ZmxL0onljWWjmnsVXzvQBkwtZ0IenOhN1QKtwBacXgm0ga6p
HLAgROeZqXcZkD7QV7sBVaXpoCrqmJYIwTmIPgxJ2EudL5eh6r8OF2wTQP4k5RT9F+UfM6Krm5W5
ruREh48Lyo1Ecyv7zlKLSggq1/h3SBYOXBsc5P0fJ1xPIK8ELQdvEHz6/I5bdUU1mj+aB8an5wC3
eJgkwouGDQK83kDNy70dMcIleROD0KqcRKAWPXtAY1VgVbIwPUDLDgeWcXy88ry10Ngtcxb1/E1s
zATeyBPrpx2xKPka2q9yc7VN3Bk9sLecuZrZGevVOYew4YiM/iYrSNezxPW35Vl/DgAP6Ymw+68R
zA01fmVh8NW2Qv9WgfiDKvfv9ao512+eCN6/PwE/Lvm86AKrAL+kC/dfM9a+NhnHU5OBZtQkA6TK
M3lT67VCbtAN9+7wOb7OcqxAQ+LfR7adsfOibowj+gIVjCZC0s2Q/F3kqC3XhF6ePNAsyY4SgOfv
BNNaxcU5nAj4h3ob4Cq3Xs+A1e/T3fM7EBCfiewpsVwlxYlaGTxm0uscxWl6OCi6fUX3Yq7zj5ZG
+UiStr5JHm+n939+vRzCnj1Mk5QoI6EzzMpLYu4+GwdtYQT8Se9wLea6/HYvNFw/wTc+ylujqXpi
lOBgLahjVm0jp519lqN2JFoj1nJIdRXr448+uDcpiza9I4UUasF9AbMXIrLztVUFIRgGOF1uurAH
ONSp7nHAVnOcAmrJ5zRN/wo5ZgnEHWQdjz//0vs0GrS8RXmCgHOFGKcOZ4cX/GyxCSsIZQSuKPXt
LZ9f+ES5X+xVN7NYC2eC0aSaSDyrubmnfnx3L6SYoGDqzbsNK7G5oFGkBCxNcqXlrA1mn1l1o63t
aJweN1CN7cpRgszOLB851Fu539tydt4UsWxFrsF3JqxPAxeTt5Y+EcYCKa9kMKIHLq9FIhsmjbGM
/OhUAJ3Qx4ztP8SwnZWLFgpwRsJPH9zP6ozXC1k1phTbo8IGDit7G98KQ860nX2QP4aDW77MR8l/
FhbStB64pVM0Pm7/koh6rV46wKB8StsSPUTYpM9KSWvnG/KyzZ5tL+FPc9eBGSy1qYNjlz0fOVNp
QTcrkZF+DZWzowiySgeFPFAYh9b3titFL0FOPkwD3e8Fg53r4jzyYXbK5ZnNQKh4tq31vJWB8Vdp
S8mPmVWtS6O5GbF6erIyD+mHTP/aR2PAIrRw8nt2QD3ud+WBH4rS4BqTCfvRwoi41hG5LaUtQCmT
w8Q/6ygkG+6WefqQZjN3di48szdcovbMLz2Y0WwzTEwbPVoXK3ZCzRWY9tpNQmUs158A8n9gYncT
1o65RmtlWzfMTsZ8/BWkAcQCgBil33FQm1Uo2wcmQ6G4Tc3n3JA92PX+JRNTmV68g87o0FnFl7yj
MXEJfsUo0cECJgpc+yDgSsClx91s9J4PE+YjbBuxNlai8Yv2YyDT8vSHmUuXZHhwOSRQ2m1Ukg1Q
AkgiIQDFutG8vnALRjn2OwlhwoiyMLsF4LrzvHmzeP5Rdkty1DY7MH2XWERnpxIDyisoiyZ6/d+/
O8UTqvfeVp1GoXr2wSNIBWrkeeafc6FA13HOohHnxpjs22C/DAnTC5Qz9NJERZTezy8HqWXpxXQR
GSjUVxQFtlstUUgx51aZeovwPRiX5fSbcmfIeaqLZXB1MF9sOOukPUy3CtZo3sD19JH7dxCMz1vI
Irknez21Tp/E5+vs5z5/+sukD/92oZu8ZvHcr47ZewJA4EwHoAbHMkluf5J/memcM3vy7cL0dnhv
u165xqMrT6mfT4ZkqGbjcb50DuTNHF+vzofoNcBuvK+WCnDaFxv1tblWOTuw2Lu4khuG7jDZILFk
7X0BFm05F9KRS6G7GpVjS4y1eq+V4sykyipq8HgvA2hjNor+1RM0gIssJVxCfVhtxlwOKA0Wast7
8KlYCKFhxo81/NDGEY6kwiIUU9Y0kyj71gN8IX22OpsCsUHZfNy0nd0aI6j1lCJe/vBA9VJ1Vd6y
8kOr5YCBygnBpiwb7xmY6EJhff5H5jyF4mo+MmGC7ELjmhELhcZ0BEKtFvKun+ToTfdK36RzWisT
hQXpApCZxhr76/Sc+bdOCp9IvceFDr4gawifGo6pWgQpikH0SbBwXo2ITp0e1MbkePEP8fiCA6lo
9edobfwekerdxAIo4Jh4EbzV6ak/1hYZUPWS0KvRWHWvO3LRSXD5JKqTVr/3EXiyUV3Q3B8SYwT/
dvTP0y2vnVQuCM/fwBJTWRqhzJNsIVNCyM/Bws1Yb0kbHzVbfPJpaxoCGslugMiDTOTfKYsDkq0P
u58QgoGNh+I1JL74jM1d+anBm0mLlU6Pvv7k5xF8eg4AUolHYU/2YkCqnvgwQ4fAtCf0pkDeLTiN
0QWNJG3WBqRaAsO0paDHZgj3ZNcm6Ov0jtGsnALt3GKp79zoJMWX2MKQbWSfRj0fmkoMXzCJv7WM
+m6SCUj5uPiw/89VatufizKA/Emzmqhr01FyG5JNJbsjecyY/gwZffbbT1EcBlT0r5iIKmQHYgPQ
7fSeDAT694nNyR8ZnEOVJif5jayxoHDMekkXGru4EVrviEcE5YiauJyhWNNGZ6emtcGwNIwUMj6E
rrNuN7L4bIfkqdvkQDNQFrObsSdaHs1vol6ASVeRgcUJ9B5323oFG0hqMbffBxeAEfFYlyZi7Lne
o8OGqb5QF1AY6/AR9G3p2Zw1jBTb4PJicO3uX6lOtrgDodQt3m/0Lvus6BSMshPApMzQJWXdZzw+
77lIK9CYcOuqbHkHasJGjElW30e55CiL3oZk0ocZHlwqEYxcEfPeWLnndHgESDkwuuoRzqE5dpAJ
03jtwpG+5gELDi24QtJeYaoT6cGeN3DHD7H/n2I+dDuJdLvWJYzwkER7SsTKOqcLHHFT8IhuyguO
h1QMP5YBx+iEDAJhIkTDW+9Qc7GUe6cZii1eGgV5qrsXm4G+9qNbM+mq0n6ACtOE8U6WjU5EoCgT
lwsNbIXgLGPj5da95Q5FDCrGvEe1PTqRgd4i+PIGood78UxyX1u2ZwSHT65IbRTFRkv/2WArqX0z
Y2tPTU3LWVXnV9dlSDVqqGrT3bATlfqh9LBfcXPaW6LEREDarkeSK1cKhGwirXRNu+CQg5IPVEDS
SwESnpoDxILBX9K9MA43+zXJ8wPvgAP+CT/6ntTqR95skqphsGP82Lk2z6qt5DgbYAEJMV0cZXQP
I4rGiKNzafChKK+/suGPPnZkdRKwUbLFTVXp8C6DnIBidsDbRVExTVldglu2qiH9IK5orKQ/LRnS
MdUO1dwkuUZVjPqDOaH68r7n38ydfBJze8vjuK6l9WcwINQEojrzibdJwdtOmiUGlRvl2ZO+I1w0
MWgRWQGdkKLtq8x/0fVp6OVFtoZoKNLWITlTRQ7Jt1bUKJ8+eMvnqP6Ac4V8f0+xAjkjWrNoTjbD
ELNTDwHQdioGFu/QlbCJFAHUHrumGKAdaC7TmWTgmHEFNfq+PylBjwGehq59YuYeqBkO9Dxtktph
9qCu+H+rom3M3ejuca4tHvKgWg6saR/YI66I5cQTOJSqflmhN106TQWNhhtiHB05cUmnwc8CW6qh
nZeLKGBSCN+StgobLdAab0BjgdzAO78oV/blS0qpodRVCZ4VsbqJZ7kn3tOMU8vYBJxdX5Tk+Zo+
02QFoCm+WO0IEy9aRO77ivo2GyqeQB3Fke0KLCfhbQ9DQCK1qJNdkmdLUf5WgVjLr5mlv83a6MhH
mmH6KAhXIaJly0dNaxovkDlZVbHt23zuyn45k7pE5B//yWYhHBojnyMBrqSQ+wfcAN3PE1s7kSkN
9JLAINgxK5a7lSnZxbCHXOFebTUNxOPenll1AkILzVPgHHls6TAsmR2E56HAhtqevfZyrNmnBAWn
PNdwFaI6WAJp2JmhPLvaIWhnlYWDIaPIXiYorW3zmyC6aaflcGG3fgmOxb2eYi336Y1iMn+pcwIC
bBdv9jX00RHl3PV117uDaNgcTMN2NdKnWnkjYGuaMN9+092YQ6Pjm0rp9krgGXvE9KWzx1SC3G8/
Z7rkP0eP6OHtGW+sW7Nb7A6SA71RK9+WmgCHwYL7byfBp2SQ+4sMK15Z8/IfnUJluom/wT/3W8oC
cMiQXdGOwc959qDzyGd37ex+H1yEcem4xXxqRCh5QsYwph3SJD77XJrxLSwAbqwPVlB4pYPWBr5r
tBdLCXZAxEaoesJiaICviwdV1/bbtLU2vAHl1+nm6k4X05oHdavQ/hWg0j2ICUkyR0sZ3PfjMO/W
aSdlIw5whsu850phXIN4r62SjGZOGbYsZxci/hekwRVu7qyhLVT8blHIPpcT7BylwPtY4G/6yqHs
Anp0eJ+AD+NBwhVE8RTmTgI1tUMqmR+mgR3JGMgeA6/eG5fb69s/PAWfK+YpHxgGzUE5ZY/j1nT2
vn2924Tu+dH6bJQOb9PQmb3TQYdKzsR88fwhw4j2b7+FfhHvPfPP6CTBjOOmtjX1BPC0+TdxyfgN
0QlngxpF+3EgXG1gB56n1Livm776Klyd3/TotFRj0id59i7Frr6aP3o+MjsAqp6fJdeIMOBiU6E1
gm3VBrbOoXm7D1VXV/b76tolbs7/XKL7SUFKbwV9l7RmgVu112rLyC98gLq0Afunv4XUhRBfCnuY
Zr6rg1gFGJdG3yhVJIJAUwTy8nS4g2Lw5u3V7QL14QoIBMtsHcVXkMIG1nDQvtmr38DTO6imfqmG
kATZvsq3w9/88Rn9cyqN5bkYlECmmt2bXWLhHnG+jzhmO998YUKf6Mmq/xHEq6tpI3TP70DT41Cz
tqZuj39F5GvBlyOkyu8WuJEaR7CnxYnsZca1L//80XuQ3J+rRSW89D9gMQsiB1LXnJiBkt1m4l+m
xMejId5+VAYCb1etCiFWH4JSD1yeRyyhw3+/OtiDJIbeDszAZip9F5myZk+Sw3HdXyikrwX/9mBs
v8F8w6OyJ4qL5x0f4OzRUpZQrPKyA6Wp4DU+BvzCSOVXthzmhSryFSPP3Vu1hMXKfWhmTVmdAlrL
ykuoOLolc/hyQe+MRHjjl+TdbQmC6+EYX1CgVDp/7L9qvCZd3uxIk3ip+vS/jRnflSlFIZ5w2+PM
AS08LdHWwJm0/w0ISy1jocrIFI6vXX6dR3WAhR5oP5NASO/3AY2HkjhBE6+CULW9ccZAHu8Ae84c
7cLfdtdcSvEs9yVhIXmleV86PyBUdq6xTULRAXEnZtFLUoJob36RofU8bd0hjsWOZyXpct9So/x8
XrK4+dh3mPDlc42XD2YIs8N89b0YpDD5xEsniMzo9MahSfoMfqnDi4kNiaJFfxaXvtdf4BBZbX2h
uU/DZNdAtkE0nfC3aZ2660hV231ohnnXzPKFZd7lpHjWbkPo78k6OKQIsLw2KQYrOUfKv2peXVgW
OirFasQWqwyIEWm/SGEjszjgJZVXuQkm9dcrIQmnl7Lnmrrv45zufL7H1FssuJCq5xYV85UQ+jTq
fA5pzTZMKJXZ1/LaEgbPsBo8HUP7NdH9pWkGRXChxewEmvMlzQEZWVyoP22S2XtOPt4Z1h+MImS2
s6Z9GNQtTxkvrfKPkso/Wmq3/qly3B2iNbzGS9Dd3klTY029oRzJ2BlSP1TmxKF5/o+OqwhCRE1Q
RPEiQ4BQ+b7pBWk/bIXktQQOCTS73x8DC0kgDcKYvZOn8LnucdR/TvO9CgO1Dq73cMyqOGp5RKLw
pKQGG/XGSESJspAg4WRVd/dm/vq9VNzuLVfPwIYUqt/KOlh8CoP0WRbzZU72muW1/AGErb8rsb5Q
yXYkCNDMKvr86nSnDdmsepCbIFYLu9as1v9FreUekrvRUblGlrABgpg5fObgpLEosRUfC/mkFry9
KWyFRXXvkSEZP/ReM7WFXykj+Qgdb/d0WL4zqMVsv3mAzh5eYWJYlgA9cdJWVXPBhp3baacgU39O
wSx42e0zmYeQtGgxcbB9tf/+zPpQK+fQ9WqCLAVH8Mg0JqYiBopem+Ly9mbTSqLPhR4HsEvymoAU
LBKywnqWWVaieSVInfaeeHGimfBLp99nvDS0g/RvhUB+HS6jJjHqaFMga3oXVAcxmgS/F5ui8JUD
6E3P4AGyNOkOjYB4qeFVLuQ8BpWbBDk7Ri6w7MidqWim8wSV9VldnGU1a2mBEw/IqyZPfOj7uxlN
EmkGKwknEeHlT1HB2IeCN+Hrq6Av+R5AW0Sz97M6f72NozgMjK8TrPRO1tyyfjoeiDzOiQJXiw5S
I6wLHrNVYBW0rg25bE3q1eVvRI0tArlwTb1SRLku2CdulSeRdfkKEnNNlQ+KZPJh4/3mMMfawJFx
yBgLfedMAwhaT3jprxAphNHh6I7GXssibKrSSW7mGJLglJWuQNmasM7DzGYFzrO/kHfzJ60kK1/6
GXAdjevPvbo7MmDcgFe6vube0ArtuQ71MA6HODbFhuAD5CkNZp1wLkCSgDLTA4pcXEDBSB18fYfb
y8/BkT94ix4QTHPFV/RIjQ/iTucGN1dTMPIBuE25ZD/M+3WaxtIOfrggMqryJ2h+GO6m0fdIpGBR
XOXldcsFTeviJ3VMPuYGHCUxEVfONI/MYROTb1QZ5ZmyEhP6Hq1VZtTvoO4cugOqnkjQ4edxPkiA
1ftmgWkcynnrYCOWrfuzhgsQxDQfFGTd/aF5UaquarUAmQnvTAg1AUr3HNumzBhVZTBZiicJtr+y
HyFgWYJTqJYk0ZNKunYzaN+cYzalQgcZWafFxxKjM7oLqZUd1ZYSr/i7jNUkcMNJzoPBijOX4py5
Qw5lDZN9mvGSoK+kdM1Ph+lKzXRI3Fcmk3OhALi+xxMviQWFzPpe292o0djTYKHDdNUx7vYOZ52z
CWvZu522KOkuDuY3g9BFZ3Nt56jcAFluHF0Vb4CyhK+mVLCUl6YyXJJV6B4iXC2CNGT6lTwW9RZY
JCRnH87WhPRbbLmK2kuEw8F4PtcAg7GggKtju1dEdDFlUhPUZv6kSWPVnnRNXDhmZca+BExl8EdZ
6SRT9kslRlCdX7xvzGauL9PXqFiltnLpOTD7e8s0YzOftmFG4MGOtCVfKrZ79wNj0M0EIOKtWpac
TXB0m7TsweF4Lw4A/O8fJZDfDVd995J4C/7gJukn7C4hN58UbrOBWPnKV6afNcDiEAgzpUhZpd0z
oiE+0A1A7OZtRIkc2pAllyjOCVWevLBGeMq5+sv+khKHBQ/CfZgBNMzYtboW8LB5QSjox8rGcq9V
rpeav0qea3pf/qfPir49lXAmxMGLwei+h710/d5M+I0m7VMadhNHHkZTb9DHuP3Onb7RYsrw9S5b
uN+YmfYRHlDwEbW2UgTczHQNYKza1QvR8m0AtjdltQhL76vslqXDD2DKRcvmUlfSFgDyqall6qN/
IvnZb6kNymdx9brrwPZbJdv/Qu3Hl607B4QkJ9wNiobFbF2mhDv7JnEyF4VzMS0/+n1lLXdRiIFn
lmyUMRHNaHNVAOpK5xK/AkJZItEEDUAFYrXmGaHk1oOHft6d6JJW/vjK+N/cAVEf57CgXI6gexRA
4PZO2HQidq2EPMhTZD6FF+s/K8lJGNMJpSziG7mDD9sQqbHFJHSD6aSSwUD58mNs+tD2K+57/ZA4
dcfCLIzh43TJcYTgj3wzuv/O8aB2N6KJzuWFv8ljNcmDUID/Gwf6EC/qFJVCUtOt0Frix5PsIDHx
yLwoTB+dk27bt8j/qvSPpF5Vaapc++OIfgeHoyd5rJjkQBlv77mPT6vsGu89V1XI2bGpA4YEMGKo
2E5931fK+qw8RBwA4uuDwwNf1QdCH2Qetd3OhqCRow1zCLudlY6inxjG1QPIWs/9C8gCGNAnjmzR
kXe+7R5J3x9LmLpNlcOy+sokPq50Mmvoxc0JaaahHb/LD/C0bTxJVL+wS4fCzzgf5ejZrFCaenU3
Dc+aiGly2o6GfvtWkXKNHDP9e4lqwqki77Wgy1r8N7B6JJKi9b63O3QkiK4PDcPiy99wHHE2OKCU
AGz1YKywJluWI3WT0NiBMCDa7kyCuiwqQoLLE3lGeCCfWYnwCm/2NUBqzRoTumg17zplG2nEimTh
eLsZKsdQjnFdxGGkLUZJ0z8tR/NHLolnnU37QmF/Qs704S1Yi1PneMLL1qSrJByCJSPm/jbAx8GS
Di9NtA+d1dhagE7K6uvkHJlod/nM+Kd6vc1/F1JMAv473sjzlkwnmahltboynyr9+vqxu6yPZFzy
CeD3QVzkaH4H44+1lUbfKIWbnqicW+Ab+/sf+VdK9LyzFEWzHR+kVF85EHyN8CGNwPcl3r17M5if
K0N9fvLN2eTcL4xXvBdKFmuzQfD07O0u4LKyWpMl8Ivs2KN029D3nN/4zsRuD2CU7+mc7pOkH12N
09LwOxcaNnR4bpueCcRmMl+wSPgtspBdLqIVkdol+rpqbe45TyklwEV4oSf1I14ZjQRvqq+DTLSs
ysvdLgRKFSF3KYtuuPuTX9Czsv6WgNKUnA+/GWO0A9xrIILZwr3mLtHI3OlGxjQlxmPW7B7MXJzR
IcDuPDYkSTCPwyYixkPzrl2wlON9w8hOV8WQMLqsHKLWphFnCX8M51sabv+Oi6Ng7LR4DAWLuY39
0kLtcsgEvTTW8eqM+ykU/r4QFat2Daltpg/EDhlH8+F5O+zMQPsgLaT+OfaSsdOkSGUekiDXSiXL
Io+fq7zyrrsIEdMOVVD3acWa2P7V+S+9XR+xYYjAPIxgWNneqathWag4Pts3FxuEa1kd5xBBJSKG
sVDy3d+K5WxzL6iZFp81KiLtxxJGhen9kaK82JDAKk4sNcciB9sIPzVzuk1LAbhclh7vArdW/xGL
Wvvr6w5gMOhecttske94dN4/4fyZzJu0Y/3wc/gzErheNfUmIYiyomFzFlu8RB/71BAmms52MtXf
1PEz1wro2N/a272lBDFgpJ/6C7kwVFWn6TKBSCKtryeZkPv8PzCRNEB3wdSWfRx2v/TG47k6Z0+W
3E1EOLQAusOi7GThxbj4SpfH4dDZlUvfZRBU9NjQ/rF4AZtFiW0o6Of+Xh3HUPg/SBZ+38bK/wtc
GUU/bKCeAW5XLDOfl9sLtJTGaxB48nzJROf37SnvMlt+3lakpXrsH8JIhr/S71K9+AxhtQT4nc3t
kGH7dUYjXRKa7OtOYATMmqnBMDXxausf6AS6yfE1Yhjm3AFg9RzdqLjdaPTKrLTMdCRgpMq6T09I
N1BXMwYeBSJudyrCh29QJuYYjfS2UTqmVhOEmZwVUmSMUuz+Mt5CuMgcR4ALpFn54jvXyhzghZ96
1FFhUhM2cCoOfYtYrhpR7LkHbJiyLCbYtPlxL1dbmGTeWQW3RbJ3DgLBH5kngBSWjqCnxCxfFaIf
K+0kkj0Kn3JsVdqxW9s2O0U8/nrC+Iw8wmTs4aOOlJyYWO3H6i0FNVvDs4qIWJeydfMN2H6Lu/YS
GxKrxE5/80hlsogJkSnDHr1vE2nORb8m09HW6oBlmr2VpyrFR+n9Pra5FmBcVLkTwLuO6kmYZX/J
xXpPHwXlfua3JqntkdUuNaeiSg8wT8+pP7P74y6snh9hc79oh+fQQVjcJSvttffAKgyPg8RLj6w6
KxnEc5kwmWmYypJqFZf79z/wflrX/BWK9iMtQMwqqMgrH+irkZZvkvGspUgPnYteVvhfa6FWMzmv
qSoSEajjNZuHwCUnxfxlobBMIkTCgo/MP2fLc5XLRgIYrZjInktnzTlOqMyOUbkmvxQxub3QELZY
jH95WkA3LND8iAWMwrv/d+/4L0EpcqriraB8rqw8zBjKqlkC0aXuSSXwOAQkQaVQZaanVplEteKv
LpQF8ePpb9wTO/tL4/nt1xcemqARRGsU8//0vmBF1isMoK2x/W279dbtMyjamWERRZYKcfNrhe9q
0X2tZpdixN/1Akk51Tsek7hlYE5iS4seNMP9aLU75cEb8Zgb+w2KYPMMipJ4GzngX4Aacdaet5Q2
CSzfvh41mODX+cYcgDn+1icfcKgA9YivaH2bLFiS3bJnZgd76X11yGPWy0hz4Qk12p5jHCNp7jGn
rwwjuTUev/UB3F4cDp1BjS/kKXvv3TzQ8AkVce/rMYpgQaxCRQPDexYSo1sflvzGQbwjWDuVmUKZ
kzP8KFX7tXlzNyu5vSaIe9foKsyHJ6eiiJeQMQb6l+P9iaDDAdz/cGnI7uExd/0IIcrGfBSij5cA
c6B99xNItU8dOTNRKj4qoaiAaydta7i5VjMeJRj7zUQp6DnZYe+ZgyoIOn53j+ErnGELeDzP7pne
Ov9vaFPXeGUGavz+ttcZPx7mTpp9nsStFdvsmiNXy2NH4MlSkO4s8Wt+Xq4q2BMdE3ugQ3qaQhD+
vIGsx7SoDHJaFGBBiEtEDi24dpy4JtfWSPk2tkHJgdU2GbsktsQUmaxV4esV46dGBC1/St+lTVwS
6zy2Rku4t4dtcsTP5d+sNoT0qPribatcXfW/XwLsTfbADAG9pCtclAnsVQhjCzKcSjjciGushPVc
Iy8gi8eVucBXFia6us8a0YYdtd6wErXMgyi1ZpIhtK0RT2TBImNLuRVjVZ911/FeDHW6FAsB1R+c
wdRrXDkMHOjvwf+j5dMlerRR94hNR+ogTN/C9xI8B3oDM+WPTXIwJPwe3W1eze+YorlMzrX3n48n
TVNJbpsPpoompxUb2Hl1tUTF9yXtSiju0iSovOkX/QgWwZd8nUuSxuHetwwuof3hbZ1+jpszuQpp
w1JwJIjzxhgdQZgwgqt02Gbew6SybihFyeE3sAYr8MsIF5cd5GNGJkd0/Y5ZGeV6q+zjQdda6yqE
0QqoK+oXZZ59UY79UmKQ6WO34uEfNKZlhHBEHNPEmimi8c9zlGpbxpMkna+eBNV7/TtcwIV8Lhmy
3/V/ESLtERVS+02CVo7gEF7ydRO21NEcfWfYVapIsdCPfjs8y2AIywAxGpiMvD1JXvEumJoFRzA2
m6gav60pue1R9uygGSExH/dqum7bUplfOUwu0lEvsg6l9mCjLS+Zb5NgaZJjA0bXhY99yqczmdVi
qSj/RM+KuIWDQFfSVrjxT544NKusgvuXcqssC7O9aki2eVYfbzH6Hp4OOpsmi3DDZzzKd1v0U25Z
MvGe0/ROU5zoCtr7LAw+0elkpF+zuH/CgswxyJD7NqYp0kDPnnuC0TCkI2f5g/ATDu1TCIx9NXbd
9AzSEK3IEojAXlBgO9lZiM4R/dthkd/aYquor5WFJ2FiKeu81htkI+ICZCoXcKU8RWHxRytFQMug
tn13FOxyhwA7hyat1OKBvMYn9w9DXlFlYOmG8VwcOcO69fAOeiu1mZLZ8Vy+aiJOLO9ImC69vGyo
bv6sZOD3nACZslnU8WcsfmvuBGeJgckhDFQRP2e6F7oz5LtKreOvjSPXGq/HOyyeBmMLvb1zlse0
FkP2HM+/1NvDHEuA3JmUUSAXfc+v0/9PeFSJZDqm2DHk6q4ME2U1ti6aAClCyPoklgvkKBGgTU9P
FDoh33SPkiKwHV8LonYMsGPlmbR5WS299oDRwKJmc4vPTsLTnlCoHhsoUfRPTn2R5ogB6tBwgLi6
0xqKzVzj8KbCMbMVaMWDFLYK1y29cEO2BDqZy7kn++DtM5qFos2Xp7hSRCqM3e1sKbSzOT17rU8A
R4zlm3oIVJ+Lb4WDc2xkErs9rmjB5+obzH7I3Cp1fAohpPvORQt4pBInmYfJYq8V8WImf1DAW3O0
MN/c+mFJe5NveTX6xtYf7cZGNK5+7HieA9S10eZK1aLE7my0TdQ9a++gOGwAejiurNvp23ccH/QW
izV//4H813LnrSEqNw2c3PtFenY2usYeKyIA7GTRhCquE1QzaYMAM52OmUpIi+08eLEsDQfa75EZ
T+n9LlOZigh2ZOaagTuRpEkWsP0DyHwzKyr5cQ/zYzOySnEGwLVHnN1qYD/YUJ2g9mvT3sACCeoi
YoBDy1PP/aR8dyxUDu/ejVt9ijd/5F49x6rkdTeVrOhEBoXJ6p9fRLmakGl8nVBwMHJD4yJt/6PZ
wFI0ohoF3AvBI8dHmmlPqTq+uhQdd7fhuvRx3lOxFajdeIECBpWa0lWeL+12D2C1Nx2p/WBecQoC
7eVOT1+Km6sJmB/zrLeWAnMBjornmDVTwCOdcJIYViJdchzmER+ODDMXB1GaYKoJoLbaudwvEv6U
FXfDRgpRPxW/f72ltNt+void8pl5NCzuwJj1KulAj7/A5gugJPWsUKpOgWiy2D7bVpNzbaVTNNhT
gExTIDWohBwqPhkcwA1G1PI1HiXI5qHDn07ydU9euFgjdZuxvAGkz887cSJZSYd5sXrs+JYj5coY
5v9ytgY7L9no6t7b38QaSkKNvEYOBtqsspkiottA3I4H0jAQdeHh7M2AO1D7iU/i6O7yckkM5GAI
Qif6kcAM9WZwVq0u1J4BMHBswnKHg2K5XXUn1rErpu9M1MsBiOixp5UtahXs2NSD7CHxpVW3lWzS
p0LGKEfyriKjp81yjgjJBAwGsCPejqvWMf4Q6/aId9fL8vHKXCXB0JkV+eEOj8GSAsoOcHcWcNcC
X6GiQNkxM2ry7WJgBGUoVFyJybyk5l2wFy/m4zTpQ0LMPgO0H8yunVvKa27Icrty+6GPnU2XHJXi
2nuCPhp8bWmWArOJzX2U6OfnUVNkror3IB4c38QlI6l29/HEN/dDxiGyw5UoTd+8Rg0IfNrHfuEj
LoVcMUCVGRHAmRdyRFNI/YoFZlYMe0OtdBIriF03P+YcgQp0nPr9z3pPUfKN4Gpzaofxq0Il1cdE
cvSy/cmpw1/TWjV8862IAC0N4UkaR4aQ3/6IWvNqmy+2HtWQ/OZvE3hA29tCJBU+Q7eaCHas3KDx
M4l9RzwjRZ0s9ZqfEnmUMbSdPNmihZ0gA+f0NYaVmMoj97TuC22TWWgvHwxPdkihFYDsodZnmfeU
C8RnX+4qHXwVs3WQCmIJbrVYxssqgwDUCOUHzzsmyM2DMFHZ9NMafgJmIb0TqxYzwUCj0q5xI6fh
60DEXxO54yHOFxNmc95pXxhQZQh22PRtI5+NxBsmL3kR5Cap8sZN6MhDF27ZFvhYkoUxBbVupEud
CTxIzfi5n8JZ1qNDzVmbGxMGtXfMZqW+f0ZaoK+cYlv0FEgNi2/6InAwFU4GT5MXhSGfTjOxaLM+
1IUYpm9bDB8Q3h1ORbNs2fWLSFklMFW7jej9BnyMo5hK05HWedngspFlEtO10t0TO0eY+iJWDzww
V5XuRKtsHecaS3xozMnhdxTh7G0IIyGga3Z9x+e3NSiIQSS905ehHvA3/QeZpKaxrE4pjHsD8x+e
MeinelWVWj7EALit+HaAkB0ZfxQoIJBVOO4TJo1pCi6G3vl34oJKsqiJYyJGI0jm7kow5NzSC/D4
ASAncnZPGul59EGKmF/vkSz6C6zV/44aPE1dbmpr9C6zM4L11YYxknvt9pIjtw8JIJjbAN7soN6s
SzLhpd6ADW7scynCTi4EOnG1dMFK1vUDjRpxxDwDVmvo/Ro27g4+1d9impa53qlEv2QhaU0zgUxz
L7dd+i0hwv889pyBLJ68M+/Y9wOD/oo7uNczRSGUdED4E8WOEVh3TPO6S8KqiYP5EsA5RcWhDnWh
05SGKyqNQzAQan6WtQHa3zR6TrhlLFVPKzMTYOJzDGZUGCEhnIr6/a6qTf8jgDjnIV4rMwTESB9E
K8zJe5YbUrhPsYqXFP/vnpbUsn7gFuSBdWJb5Q8wcdt2xve+0yYXDao0wAcXF85G2wLrUOJNAAh5
rEowXCBNOU6KFiiBQpxATuWne1QIsl4MAX6d5coKl7Kho31mxCLVZ8K7nPgyQYYwPB+hw4EX8iBA
2nE/YqZmBgRRPxLhkp6FAkIWjULd2gRSWVxrsT9bsHl44nudqdPOn6dxlSGQxXo7hPEjv9bPBE+l
1sFOnjDamwY/7LDx49AKwhCnYrgZvlrLx2AN1nGY0HorbUBb6Z3DLJoWq9ZkdcCifNpQ7WjTIb31
DNvMXwMcNUk50TVskiO6tlnurw10nDWXpKoIPcS4YdBJ6jlH9glJxEmufAJUeXXGbFctOGCUOTC3
oPwfZi3nYZiuemXxKuj4FwYokK1cJGi/GyEy9QiiOV8G77XdGxByH/2V4etCamgktAYvhH96Z7h5
9zAjhMXW1v8QnDV04otbet2dkhKxDDV0ANlIlZ3j+MmV4JHfvpwV4ViewyIxyYASgEmkseO5F4kk
wLiKgmkPMgBWvuXBKCcBWbo6OGmMOomiYsre+FAdqg933FOAw4mDTW7Pjs/QuWPTnrqQ+72E7ebJ
3yaVOcMIlYq7GAgsWVmsv0e8vNgghebyb/l7E3aZ87vgfsMYqAuZdg0YNx+WjW2ImWFnngQSeTjB
xAD5w9GBlDn7WOh1oLgdLbcYVQQKEo1hhnS/9etMbSd/aOEDKv5xPDgwV3fc1sjhJ6eDt64XjzH9
nJv2BvM4srSdYaZbg+YOVkeHa/KmemABilmpdB1lxVTvA3Iuw6FO+0OrugNKcLNm+4blZ67OLaYC
mrxhc8IRV8D4TBLFwLm4AdHIUYkVRxwlZpEQje7ULEADHPH4J/OsP2Pjgv2w+jgxhedz1QvrW7i+
YR/rgEwwPwfxcjtnbPgczQZjCLv3mEv6Cqxx1vI9IjMZSA2kqUcBDfxAs2S/+0BqZq17EHO5jKcj
44nM07DlufxTjP76fjUk4OcWkTNatjBYDhU4MEOrmrFk/YsEF9cku+ewEPKlsrrW9nvz+q8GchVL
Vdofxe4K/xonmfgxQ78mBbh8wmNdfOt6dmDKfJPJ9kuMb97Gi7GwUAtq8ezK2D21X2I4QgKzIxGd
LiADOaRQ+AxUV81YBCuCWmt+ammWq0jNPFqX4aC5+hQDsmy80NKzJjD7vV8eSvGe3zfTZHFj7lMn
ZP/Z68Ajk73D2DVDuhcnGW0PiP1zuAAtFwfhOeuw98d0LE5jtCqyMsQSxdsrommuOL1JnuUxN8IR
qVe1yTxcdbiEOl0qoml8R2o2lx3EvmvQGQIWDks2niMHUfQgxD2hsrZwyl8isyNx25waalUKrOA6
sCVrckJMrAGRSrPVqNiuiUso8na154qVjZTsxYQg5aXJWYosfInyVSNpwHFpkt1KHqmoerOf24vu
LLFW6idmV/cFRk6wm+gI5Cn+dQNm6ka2AirGUS2z0YkBldQY9CJUsgQmFLmKlPejZ89iPAqMKLC9
hyAKC2DV/R/73C1C3CD5VzPDXM85LIo0dJhYO+GHy86zdxdUUbLJb4PvoJKqSPycykU8a2tYyC1x
jUTkPfQzkhVMGG9WSO9gH5Q+nQXSTGchCpYPBqCMyeVVNvVnQK1esF38/20afkJR8y50TOiPx9Yn
jt1o1FwkJkguxBPGxrnlaPJF7daMzZyr5ReoafzCMtOjOozPggjHXksPWHOtHpUpdt+SbJrqg28p
buzKgLLPbQV5sVeZKgbPRW6Hk0Vyt8dPtjRbSa4ATxCAl4ADgFeGUFgkUPSS+JTAHp9wZRUC49AR
BSJIvhQ4+vvhXqgIjX5tRxwF0+DLFTUddQvDtLIAygKTrNTHZUcf1sAAXm6WgN/w0grIc5yPKl+e
XlKimaGHwG1Mj/6BHuYWdIqifu4C9YQY0tl8oTgOgphoDpaMI5vQn0UEeNGYlxQuNG2H9YCnAeIK
UENiIfb/RuhBIr9QrVadHJHE1uWWq/uFMN+fRv2iuRwQq4YZjveEpuWrRfJ0ydz9kdc9I0vut4qU
GushvWc2UvHzL9WgMBoc1/lnKK1Y/zoNvb6hVPEnIEAfsF3wKQFI34QtJ94A3nj/YvfumOE2WTDh
xV490Ihdhugzl43Z5Ti5zzYzT+kZem5GdttwFEeX4mPcxZjtADj9lqj7BX4CX11c75jnXpkjcjoQ
FSXt9zLoYfJVxGm8FKfwnXdYWcal1YGomtKLB3LfbiNw/QRmuVLfK17wTpddqYy+XTrY9SSCfiOc
1Vu2YcziXRPZlKwk+Tu2AvQNLdkMrXYnV3MhI1/H2Tv0D6/kUAB0oLDmC4pdHM92oYmGNruv1rw1
yZbYV6hiEikXXfK97oeRRYrB6zrn/LYjumMpKUJv2R+CLqJ8mStJPOYfsLPogAH1DuXsCW50e0KK
FF3rLXQtUhQMiwh3JMoIMBYFx2RgRXz+eXXasDz1N4PhMoyuFsnFD2zmsA70SsqdhxvnSiUZ/EW1
9kewt9myqeJBge84hj6ZpYv/yNRYwn3ExVxWx/niLyEPuAswIAieMJhB7x9msd38y3mvgMRnFgAR
fC6oht2OWxnAG44WyAa0IicRvtmNmCAN+Yhqe+5jVLuP28KHYN818Z9QMi2YaZqHeMiP1PbadGx1
BePXgLYK7a31CEEtk5k4EUP8g9iplxyLwygJD/sPBsHCvK4cSpJSO0AAeFMCqENPTixHP7/gxw93
yRIBx9mAllI/qBRhisnQZAExRO5GDRC2OYDBMlyME45iTimVKguCKBfMfhVrDV0hCSAYOTgaflAV
/yUX1EP9MY19hhAUqHnd3xY2//guyeunNgkY5BZoOOJzP98hX5fVDHAvGUjgqPLelwshj7Cw6Eo3
lITHnA9R5hIfi2DMFsDgFfgSyMqk9UudBX2FaFwxs4zk4JsBT0b3vDtvlgTLxk3OyQueMywEHzdB
sDMpOsI3kl+oStargc1XoshnIxunuGVTGUcl8RYxZnochg8KS5ROo9zmtfXu49QwLP2RhkULej5t
gKXhDTYRqBZv8GTj7GyKZfRa5DjLPiSz0UW7CEiuaWP5/JYpN7tsLFEdBPi6qT0Rtcrs8NXy6E6p
yzk86Zx7C8WmbYL6TH+0jU/IxIxLMBNaHE7kV4LAs3Nkxnz1flWSvd34s5edqy+Ts8vXv3CwuWmi
CYzDEg1eICsDTu0NoJIP2+qqbgx2mn+SwfaX8ohW9SfFMzzBE4zUkb5BCFGw+RtG31H3FwmG6b21
kW+/8ApoVgHqQXmGbZ2sTFrdTK/DQgEiuEgengLsWovcD9/+ufWJZvmUJxW6p2Ljv8jkdT4Ovgjz
sNyRkNTKBhyjaLsL1UJY5xuzIsWqfGcl7M7eH4PFneQ8HsGQxPhdQ4ypzE9VrrS8jFXATCbvCAZX
84KlNn7RV9E3zMPoG5uD703wFowv1/1VV4RYBm+hL0WPbH0XwvpclPCkJp7XgsU+ToRcHa3GegVE
VcCekHeMfCWGoEGZiIx4//1MNkteH7sKRW1DF+6Hz9F0+4QhAxYHA/sJNDaefBQI2rOuaOR9eSdP
UHdvAeQWOunmiQ1p3auYOBPDfuyfYUn/ERAYLVbs/mzJVvy/QfCLMrnxeDSOVdXCfUe5cU7EOUvc
MWD5XDQRNKjJszBBqOeGTfMThhS8EWlY4kooaqUh/0jlBnWqfWDuTYcOpJy+GXndaL3ooTCwQPI4
plB/UtJnHtnCqXyTtzoMZ/2H4cytgmgQdLRiyUGKhaDDeJkGbbicaxCl9qbdwB27ULzkgJaGuUwo
8vpLVqoOL6/nJQ+x1KOQuFzSJp6tf+7oB9J/dM8skD5nIAZG1sU8LRiz/DnG4+krp6Wc92lNSroH
5D/ItKjCeCjb9nY+S4GWKb6DcDGJyoBEdX1Z7ZEl9pYj6D7PiwzA5MfoJXkk48+hYCNSnOOQOrTt
VLHOQsLJ0wuZHmnJo6Yg1VxkFBm2+Kucu6L34zoSm/Ak3hlqIcz0xPw/ckfw2+LcaTGU744VuPDM
prWv4J4Dq8XJCk4kWaRL1Vvu58YINy8nlnkJRrHV8mDCuAyqQlS7HkrqWjpa2orEEPkK2VH8sULb
h2XC0Y3oPX5RnDc+62sfPLCFnsqeaLBeMUL1414lv29hVYlPS4WyOIWUzqkeTncQ3IsuYc90qcXF
b/MEBUUHXn3vHlteW+JeVc1oilPGNA3QldReGIUPGRFYp1KzCZdWCrqpvRr7li4DhYueE23/gukv
QWDAJ4SIQTapFKVfMN9oxlC8M0BBVD/t1JQGrgdmFcFc4GdeLnk4gJpVIxAa0o5AJ/+woYakmAJ1
/28fhQZTs23Jvr9ZQ+rCEvpeiwJwIfoP4k0b/zYCVcdIm2OEdbuNfH1HNCq5q58pdTLu2mwrhEUg
alRcF3jMpqBaHfq9jNJrwQem+O83TYN+Hr68RDlIufQNV3nYaHOgcXDPAK2eLAAwgXuZm30eNTTX
QMmDo4l3pJet0iJAsJDLFTgtR+OZ7bPiLknivENzxhdSBAYfVPsejkQdxPGuexT26JDuaOjMwOvC
7Ed8fA3M7eDfYcHqrIP7tOelBFVmXgWjJWtF0wK3Bz3vLxnJ/QiWxC3CNnDfANfwuc/1Wvwl4FRF
Upw9fUBJQRs8u7fTmd2rs9Nfj4TvZ6JQRsb4LIgG06sjdMMt+3yVwMl6ZQ4DGM64OtQs8be/nXZ9
b7aP/lTSNGuj7fRbgJg935NyMaxui0DuUJWYqPTqV5T0P/efbhAHybcpCT8Hma4zCZlyAZmnkkYV
jvTAbt6EEayzReGxpkMRnAGrpgW2wsKrC+OfPrnjbJWqFUo0CxxusAbW3iIbmhuaZZ3KlY0FhjZA
+ylx63tUc6Awk9sveg+jpOoIG9E36anGShh0xmO8jSh+4tsFKzFmQruBc/O/FSG0vyluIh8v1MoT
1WPSlXwK1Sqj7BQOXmx2LCoPz1WlzGo5VgaqrVcad0xDtv2AJWddvttBdqTgb+RTWtf2kd1XINyL
A/t+A3mNJn4bMt04medgibzJ5pXiT8+t9T7Ly2olimGM3xCB5Z2XdtzPanaT6erUitGYXJx+Bd/L
YjwhGxyY+jXdojEfHAb7+vcsSat5Qne3jraOeHNGt/GU8Gepy+Y3dAhH5nP76b5lYKkGjWJSyyEE
nYNa3aqboIMfHOXUk+FuyAkZV62vTStA23E7rRnczOZSSGOLjGUWkfz9rSHY2SteIs0uHpYEKTeh
8iWHdZd705i9HLS/mc6pWdmn/FhNonKep0g6s0OHnGJnLgCHFTFyOTZA1j4PwKFmyLsrVmTB1Hb3
09+nKotkPbx+abI0iGS2NEWUaQt+ynffWo77uOpesTkpI8vUcFlNCSEBpC5DSUjvRBD8hWP//RZv
pr91V02n7L1Oj3Qb9tdFHynzzCVptjpHHM+9N2Xin9KMBFBI9Z1t0kdBNTGLsRvrJ+WWhpzqacMy
LaSljxbqnWTUxASZ39lVAKC0NQQ4NXxweZv79mXs+Nb3egPW9ZTSc7defpu4ecKSdTOcKQeeG59g
iSvRjlGkCfD14kdz2p1yvwkeJi8+6QLSTyUXrU92VUioPS8isWvaBDlQn6bodrlYH0l0OvwfuRdC
9JP/AspYUz30pBa7x05ziYqf0rkeT/vk//vinU8I4q1B4Y3ieh5khByByUuBBBO6Xl1wHVKVeipt
5sjFudSK4cYoxTnxikxU36RIa8oQiICOm/GzHvh8MzoiU7mWdNSgNjUFAeO+rxoC2nY3Xm9hDnuj
59oEHMzBfD/foEWqz53epMrZfhkQRS0mVGjnf2l7B4S0iC7I8TjWR3QZwhkMAQB2neAgX6egoXSK
9GRpwT2H2Hn1BvYT0H15WXX7SsEzaV1XQGZzokpV2xZjj6dt5dBdBzhzltmq/s2dBh22Sp0sH9Y7
wV2t5+WERdEkmTza554P7Nbxuy+H/L4+tOMMcL6CY9imGbGcVuEdUbNJ6DuD+AZY/c4EBMPsdPxQ
yKmJrnshGJcecc6wrkFuqimDhbkmrBkfIiWGO+V3Rva/WjBlEl5Ju8o7eGKxu86dZVGOPOmMzFAk
fWr2A7YmDwmJfTauHNaSZNnY1+y2Q2vG2eGTJ8spYQm/JDr44QQ2vwq0fXgpl4nqrFPvcgnHZ26a
H+ogl+04A7njc0xRJRNXExX1eHtnpritT+rl+XV3Rbk6fVfOrsbI0GEieIgl11QmcEXzme362qgl
JKzSdrFpPTn7MyqFC/86Cei31yfHw6NJ4MpSy2YRAjKxAcSoKxD6NWChy55Wpep/LY19zpFq96tE
/z4R4BJphlWICwgqGC9GZ05oeHMO/s/QrNY7Rph+5UI7oKsSvLOUD4pLecmEWtbzLjco7P7HaneO
//b/sZ3nVy4ZBV0ZonO3qhPMSI1tq8rR4swSvWsJg2qx1YUGMU0iqQNrjjVRBoj5Z54GIRh/a8l5
y8XuHCITQqtsw9KY/HRba47ck33zJQnyEUMVYPKbwiqv8vrXGXgB8iHBDWYjBf6wodCKC8A6jeuR
q065WBgW8qSpDp8WDR6+MVHp6lS3HS03bZUTWcVT+DhyewUsg1FeecwxxsZweLFViLW3prEQeEzo
eHDOQ0PLdibbkx0FjPNpYPOARjo9OXmLWfD0+M/ej+a/XxZbg4HRyph9yNTufdyUyMIjOm1i1YlJ
G9Xh5SSFniwfpsR/vFekbtdimvc+vCMuinv6RirEn1QxNRDyh7KkAE14d1OKvBQgq/zHy+LriWhM
XlR+CigBKkiic+xpfPufpO0yGKHFkhs7EDD1bQCa8K95yswxLTPHhLB7LLs9WsUI5zFLnAGj+z4n
BvbImhWBCgHSIMgf2EygUX3b/ZymF1ZLee7oW1LNXqGljB9HAW6tbMcZ8N6vYjPMGRVbb6UkJG+a
Rjcvzvzw0Pj4FhwzuqDeEcVpqxruRcZPiFjD5AGjID22wUTeBSPP3tfbUUGJtxvBax4Ig4zQi1GU
ZTk55BCfFBLMzXXr0E/obnwvif2ZPzCiPJ8pxjNl8fnnkA5bK+VMhzTsu5SvhqBi58XZKuCHnyL+
3sjDnDmsraEjz4PN49jerRwLmJs2pW6yPXEMsbxrNClgkykiGfGmL6yh4UcpWX+OD+Eu4o2t07ri
oY+hLQpLIaVEqSURBPv/y8yZNgQNhCf6gJVHw3AD3MKE3gMWI26spJCupw+I01/zUndFalY7eaUW
kwZtw/RHlI4zKD8LqiF2SuMizSH4D7KC8A4hJL0HODLmCgA3gduhBncdEv8M25u6T6TrMrbw6U2l
7SxwgCp6Wlsq2ATJChZVyGuZAIAzdye0FVYuPuNQCbE4wKrv5rfvFEmgJvOpd3peDIK6Wkr3OUke
OUmlVKwdBSfIVLKdolIUjwmwOXplEHq2c9j4NsStOyXwjPw3ZOopau6BM+FlZw2kB953RB1YCDE4
GWtEbjCOwvDvLG1paXERvugsOJMaGCFAmUs5W2Snhuv6D/r9nOWfqoiH6YKknpCkhax169C666H4
/lEqSNTHPBFRdp31EtiotfVygYiyvdSVxtO0QXxjJnuv9K4OJanR8Dr9E/FyggBj1LycSAuDXap6
GzQxE6sLJ6BK0TLlWcHL9pqVwKY5Xr0GXFYCdKU4vxY9Ir8HYCJb+VzXNp8Kl6BbGzxMFy2G3xjm
JTORBrBScbN8Yy3Vqi3WSfHFnaKNpwFe6jIqAwkffZ4Js2wfaHrymWgaDH/M8GBbOtRSpfZl9UJw
JhlFMGq2CWJcjjqEaMJeaTV/fqV9EOVNMkGKdoS4f8FxM88Iizhyy6D7HXUnziR65c34XxN3Vp1J
s8Ymmk1/OEVsvqj5VlWscszt12UZpRQHyvkRTzqw91I/6MwrW895NGh9uIVYTNv50lbCYp7ZCH/I
7tWQl/NaGeWaetpPY4GeM4CGcokF8rnpJ7MPwIoNK9TNtuZwJdNmHJxTVPRS8jrDs2M2i69QwGGx
0LQFEeif59G6WZnAy7PIN5l9WdV6HQ0uR4NYGin2cmdaLRM8XPweQG0E0Ji6wtgVVNEoKtBc+c7L
PlXIR0zsNfeETEItLcqKQ67JKlueyYwoV0VfE2LrEriCe9v6MM3c5tVPdycSltTGQ6JMWBMZgaG8
fj7wWx8S1ioJIVG6f/lSyQ4SL8ydoPRizOrpMmJe0TszTQUStAp088A+agIdiBugYWFsTJHDk4Vk
37NEdUeHS/xwRhAOgTiFyayoMAYX2mmOZlBWk9p9jBXBqIYXhgs/Sy+Iu0wxfqBTgRnwlpg1UeWG
xjnU9emcijIb8ZH6zJs0mEiT5Vuadvupu6wGqt/COpbd7bcYwOgid8LN/c4MxAJVWtyTgS1yagQ1
t2Do5Ob9b/j2tsi9WkiCtMZUhvZKXqgh3JPLrOV93PltL+swtqO45paBpEDZcC0y4JKjzF0IwvrF
/ZDf/9/97uqAzNQeMDMEwKjFhSgJBvzY8xC9mhLrlhWQKPdZzFGVtb5kndyctgqz3IWnevbBMup/
IVNOAVwrH8dlDmWgQW/JaoFj/pE2m67v1+aPYb+/tvYW4uCJUdLwMJX9ZRk3xhggxDMR3TS0Xe6h
uULPc7OMfgCAsedNen9e0QHB9p4uAy4u/lGasw1ULnHtDy49wRwJpU4EZlQjbH3qJaHKz5W46uqc
UiWomUjlYyJGqRFbVW5TDWr5NvxPKlp29e6FjzwP3eaBggEcVEj+onNAiOZKICZk+W3FU4330JJ+
XR6h6XtTv4D3rdI2l2GZnCLorNGb0EMoqGw6aC5IRV13AKOoaW9NlA0XuF7fmH2rexYN+aH4D2wK
q9Y1E93fADpDLFOFRbVhUlnFXn4HNFV/CxznJYozrXY5Jfacza42P9d1vpDH9jVGKAJyqnX4BHKU
UqCNxz1XX7trclRjsMjTRwLzV5Spts0pYMIVfNpWfpKkbJ3lB0KQCPj9HLOH5AKYDCAPVgvhA7hA
ei9dOo2kn07AYwGrkG6I/IfsWX+uL1B/GM45Rr+4+VNideudlrYtRzzhgwGpW8DIaCz8yHe3zU3+
qGI19MMOic8yHgi1uAsnX4REO+AU/16UMWzqHp2Xx56UAQ31/+5fROf9mVl/eZ0vx7MDe8FeuiHI
NALSnIjJWGSMVGcchQpSh/gShtaaNlUb9Dv5/saWKzz/k7tAvJ9Q9fmlgfV31WZbLIVsaQfZVzzw
KWXJGuoG1ab8tLFkWmDGaVC9WC/O0CNBsoNaT7ZlCWvvaq2ngG8W6VQ6TknH0yYsfUtsfhiYmcZB
osPv8o6gTk9O8ZwC1aOPy0fMNWAr8MGvnmWl5UPCoXxp+ovfeqZAFK8DKQMObKmIIaDWu2LeOn1e
+n6Pw99oJfbQz29ahznVlN6dI9fXtDuFyAJb6jIhjxSJ+VZGAhYdhfP9Avm1N0xGcptC62MvGO72
NrjGrgcEZLhpMFZsf4i5vL4QoY4f06cbpM8ZFTEfnkFL/Yt5iE2ShBp6qduvSvNdBBPtjpRTX/IX
6wZMgThNkD6RnxwXk39Oih5ZaWI/48G5cAp0UcR51kHdNPVM4pzkrxtHF+F5oHlNeySXPJJS2L8i
7gJt/okczu/Q6TZUeOGIc/Icao4JyE6j33HY4WNHTgdA/GhQkCNwJAGauLnBhk2Z+o36cBjqfPk+
pYca087I5x1aeAd9kqgM8a4R/jTX0CVtKnu4gPslapIYXQ3u8Z/lcc/MCwSzDpu48XzV0XXrmvfN
0bH5Db5Ki1JWcgVxDaIaSzreQsFcvmxIK6eEJ7RLQ6dzpfQAPVb2DxKeD2u/DztWPJ3HndwM9Gv6
6znLpVs1ISHL3RslB/iKvFxDE6aQ2ByKt8s4pDVHTrMpGEA0XJUx5/91IKPzO99tjxF+suXsez2a
1pGCwTq7CebhIjcriNNfrDX6TTJBG2o/F218o9yYzQ96711o5BotdAThkBly7chmNE4PrP9+jvg/
OQR7NY0VN+23CmxlXW2yIPyxMteiv8i1olRSvG3pMIDrgbppuRD60FuCCxjBnSbu0l6hsVyB1hUV
4LMxOU3pPXP58sCTUat5/su5B5vFvgoTkzSkq+4mXlz27ZHMo+o/kwwHzPsgGPWtXGshsTC1jR2X
4dtFKrpMhNBkUs/In2Bkbq55F2NfrdciAJiyQ72ZmPE9ghm9gYrs7uSh/lgS0MmDOc8BtEHZc6RV
m69gp4VgQid95ZeyETmniTmo8xM1C5/KEYDr5Xw0JEHZflG/QfVfdx3oSWjRyFM7s1MvsnvD5eQK
tgr82z42kiaG0qLXxXhcm1INNITKjWtqMbqUD1GK723/Mgo1Vi+hkdlNQyDmol3a4Y2wUHhI2eUy
uM14PdqVMzwEYQ5MwZgRk8vySJHafFgexin5lluGcz1ikFnjL1NeHplPN3aba5umtxVFdcp9dnVr
OvbJu3DOWPEDu1eRpMgAou1gs5EZrBvibJfVtZ5yvbGgMbkz7Kxn209LwjY6MoaKAYH6qF8mCE5w
ZrwLvhqKb9EAFqHrg03cXBa7jrtHsfL+qqRAY8o+1Aq2zGsQWo2IKQX3cKHmmFlVrNDpofXpFMsQ
X+3ue3l4cRJgp4lAmk/b39078vh0WX+k1qN3bkhsD+F2YuU98e6Zu5CKlyT5jALVivZ1wahbdR4T
aNslc9CTpuXnk4vQzqQ5LvHlMe0ZfGaHzzvyRjdm6w4fHYW6S2RdxadmgXcEjemzMIIDyjsLkop5
lZhC5mid8NWhkAh6vfMfLwDRaBebXK+Vq6qZfZv6aox2uavnr3YW+zEOhSw4hL4/I6NtV41GwnUg
71lOP9Xl7I50mYrL756Lx1jxe4qzZBIA1q7Ce4ffYUxKY8veij5vuPZtNHumOpwUPcnKDHlC/9Iy
l9tiwajLhB116yF8Z30jzHW1d+VqFGpmM4ZDpR6mK6TPbRSserSbf7yrL9KNJ524YHkErTYvjyvn
4M/sSlEESw/4OfM6kN64jwjgg3g216bEOqtHtaGWbHj8Ezat8HSdfNXYuOCHzs35yIZ4vaFls3uA
iaalDD1/FQbtLhILrHb8V7JV1AK4P8+uOXLDY6/+b6xEivtrMobQwjlIrp/1z8CwTDWRQJNFe/NY
ugBawxVxt/9sB9IndjjuminznQtRAaqy6krOorJ1cNlFDYRG3FemMHEy63pbOEX7u5XeIAJV02K6
VBaTkUnx2dGLYApyOsN8uFcs8auxBOz/NKnVXoGOgVp77rtcHmiJUL0bfwbwgEpctcr/0FHh+j8X
ZRyPa4yDAD+vyPII/V2mwCfFysvzIUJpEA2SOl+o3TI/yvKqOK/+6pd5LUgUBnHiwBQ5oSZSYZRS
A5MJflxjfZ7xezlNRac5UfEQSNVYGc1JUbF6vKZ52rV1pZS+3NEHyAmtcPzFKWoPSpM22WefG/Ta
A20WxQXeTQo86+2pvVvgZSBPuWSVl9rjwP8vWAS4oBamklnDm8K0M1lah2DRiNzsI7q4jvgtuGLE
gwBgbAOPxqJ9kuqojXcJj3CcwARlNhf1RRjmjIRtSmKrpj+JOqb4VxTwQ/Sm6A/BoXcADtKg2P4U
c2AjVXOvKJexSGzg7RPYSdTA8YKso3VXoSGQAWjvIsD231i9mOO6Gp/0M9o/08vr0xey/SXjqZwb
1yC9tq4iV1fh7283TLoM1Rl4vPj3ty1/yFTOO/G1F5Mtldvv73FXqsV0gz2Qg4C7m9qOzAfmSC8x
S/uqmgrGnOe3A8h+cmp3TjxyImk1FJSNJa+ZNpiLfGipTuNdcc4XPL9Rjx2px2DJg7fxgZVylPUH
obRAo3GbFopBgtXMp1/YiOGiBN6/Uex5ujUPBXB+1Y9OUhVu6ehhx5Ghn2iviqQbSwoFIMn4F9R+
JqONb5Wpz7kHkW1q8XsDT7M1/CSN30kiXUv7F5oPyfuMF+YQ7HH0GVJ8ldwWyHwcdOkKXSeebGFj
bdCgCwZpd4ob1FIhcHrlf4Fx+IZY8zME8eeku1YbIQ4DJWuLakT3yZVowpAcus9v1lE3azUvyo0u
yobfEqazntdCSxXzT0a/0x+zt+zyQyH8lxp/Sc28T/JjwH0bvB4x2jfRzP2Fz9d1aieELwco2xpK
LESe11ZeprvkGv/dkPm2dHfVjcLCKhfb+mnQ9h6Zw+cYSHW1gNTxRS7YCI0UMhGW+JpXbrXvvZsG
9Y1OUg08xRLemajIAx2lAbS3nGh5xX3B2spwQZhePxz+UfnYymqjFYjO+rQ5UEl0QZHfv0Jfu++T
u5UrnkzR5Q0j+BLrmwBEr5W+r4VGeioWRvLkUddc8F+oLyiRLs3Wuzvq0p/++h6VFt1z0XcOYPcZ
IdcRf0RZHpp9TN0Zd1AaoLfW6Hvzz8U/WOhhlIUyE/ouxPbBQwgUZMwYbAYyy7ccvjOEKs+Wk2FK
xIdxKHR8st9xA000rI/eljoRMMBkereGzk1P84qHMySYhwkeEZtmjz/pYbpyUTodTpNPvfFnrnnC
FdOFoxPYxY13/K5BM8nUDBTRxf/I/lQUORcZ7zmI91DRzT6dvwi4gk+dX7E79xQT720H44RtY753
S+L3jnfqAaW17K8JumzJJDH//2e6z8I6aBioCkEtWVI1aTLcl4xSwEFLYvBDA+BaEgaXQMPL6/aa
L3NTU4VoiapEwBKv+aVOKQnkhW7X9aiQ0jAadJrJuZyKJCOeL22pecd7cTDRkEnZeOYVR6BdXCr/
JRz7Qf+MtT8KrynAHYbywIgeyoqhzkhqTOKUDR7L0PmU2/SCE/vp3NT32mnWPBxKWQnACDipQR1M
ErxaDeJOF+x2vTTyOIC77SLXkjpN2ijkUBE+N2zFT2V2vztdb8C7EwvcPEKu0oa3+pfchZMwR1kg
qKU//vpEvfCrm4LAtSUY9Jl8Y6UWFJG+BPxMV3olUeSp1YhHsua9CSUC5k3mL1yhvks2rlAk0FLP
IE7fvbzrJUuRn72QAZ9NgrG93kPS+rDprk7yzWRiSH0f22x7+dJdh1dR9WoaDqWdgwHR7KdQx2mL
Qlshpu+gR5mgEqQnZ3hn56kF947duinz3XQoHGSs6k1YTHKAg/g+prCsknDbVbHETqmLGsohM/Yw
Ba6HjITp5D3IcyV/J9aobAEFMEAIGR2z+/TqVL3f4yYscbNYzTC9f7j1h4mCWjBQvo7JbOpbZbi7
0cg8g4s4QPFLZYQWQfz3VTO4OLJDP+Eih0FXKZruRzY1aNxPJN13c85BfY0MyLb4NuV0rBGDJtcS
8UNZ4GscS2mzL6dMMDgYfx+eW+cORG4nDFveIcKjng4zPFZgIoVykveGqy34C1iM64QDYSmKhX10
OJSLkkeKnodAg4S9ooYcsz73G5NcEPwTWJn2wlVCfHa4AFCMcIy7UPOkL0zRR5Kj9FUA4X/rg/Q8
o9Am41DU/4DWfTGuUIM+82a5lrZIoLhARRgfFXvsznGpDLUO10BruQM3YrGsAlWICcupvjY2I7Os
p0OHhCO6TOKbCdcnaaOFS7CgJdlVzZG9LPQfM+yxCvb9PohRMBBkttLZCA+8pNwD0d/4JYVJrmTI
jIgotiZqdvnmRiQjRi8UIx5FyYAgQlWcz4FET1tJhSBzIMPwMHlwpwXtmmq5Y/AknPKSoSK5Adrt
+HR5JFGfpCWu09rvodEFbyEl29Yij5nggxmgc+MI78UGBLZcxZD8bX22vibjgVKFuAJQ+Nuodv1N
nO6BL1Z0/vohGQ7Od3SWbgIEZz+puQvXEbiGBlZsHFh1XVswJ/Jy7OzJKhXGlN/jZy7mCskFnrFu
0MWA+cIWe7VKAyKiNVzHgKGPgguyqJNRVVYblvLUz8ilTUvecTFaSHKj6YNlGYz2GYAOWrzryniV
/J2SQi37s7hGTUvBtlGtbeM2hlL+1Grw1MfQ7q79JRpwQNm4+AdScN5ZJ/XLZsNOn6+AMsDkf/GS
kKxNAFJhXxcgahPtIABtyxGcmmEkekb6t7Kns4EC4iKxsJAQLPBZdsADfqpFGYgKIcUG/+cEQP/t
kWSjjWfMEe+S8ImFmKBT1iSpiOvMs8Nh7f0qMZTvKJKuFAZlj6mfW7tNltIHVlBByhFfvZLWxWxx
MojXdjfWlWV7Dtbd3uKS4nLICAzuFgiqJVs2RopizFyijoNLi/40nolU6qKJcPEO/3nyh5bcHP1T
nWGZY6D4gNP1D4R7+0tWC+tMyCDqbTz1pDZOM2cqTmCvo3r1EVcC+vji9fPoImHcx415XMeIV3DH
lwDoQGD+iXPvbgouaaRHWB0a9HncCJaXxNiD3sPltqnWd4Q53ZAxgmxCj4VV/5yXZCja1FP6/afz
DHJ25EQy7ldtlBROSv1i1LlNWQu7hrX9JMxc3nKO2ZTwMoVXz3GKsRBS/lSYLF6Tx3ewSdSw0qLm
a+by8yNNbdXdUTYnbWJcYSs35C7gb6kDMkM80A+zj0MQCsQsSJLTZgJBVXhWy16i1M9AoYUQvux6
drKlaIYr8Xiw+G+Drr6WorapFnBLaLl6Tge2Tv4BRrwYxUiSMMzyUEx2FnBmw0IybarttLLX3/Xl
V6r+STeXDwwMCA+FITC0wgim00yXhrW4I/hAO/LD3fcShc5OMpnRKmSHJgS/3x/Q8nFw/N8/PeOX
ICd5kPIQaNhrR+nfOiFsTtKvW8Q0R7qr4e5oqObw8ebzAPLj/uxROlrythXtyfmUzh/7P/YF7ksw
/VCMMC5IiBIeWYF6xQcKt83gIz7r9i3LDWN2fx7sMF47rzDxrNAGGn6pcdrlh6+ZVrcxeuJmeZx8
+jKCDYoJhWjGsnHNhXzCKz+CscIvSrQWgX3bG3Z/kG2TAHXqtKNtQnaxad7jXnKOKR9SlnhfV+Qz
DN0ANOS0yQw0aEFZwOclc5ex4O1XyAta4ufhm2Ev3cqqBbInHtRRrFqh/QBvwYehXzHEs2bhE+1l
5RG2F4WAllnd5mf14YGquYVGXSSvJrNHeNhrxwY9AHWw8bOyOt8iQh8K109NiVv4Sm7G7yTU5sr+
3odTn1cVgag6BozrKdL7e8vZpT7bYnd3xgO4ZnxJaUIFg/t9Kr3ZXMhQk3cB5rAeTk110mKi1Qnz
1EnJFjAqAaErTIZ5G/JxVCvEo84A5QWX1tpbe/C0P63uZGvj4ttS1g8kja340UbucWr/L20WrDRw
PezMGK5TG/mY6jPMnhFP7gwEXsIIySKef8X+J9Gi/kQaOiWW13voJzF66Abm14buqBp02ZdWPeAo
uLg7RWRadtuYARPuLNPo1XvKqPvWdvF0KgmCciAA+PWqUF1SqTA5d5dvG9bhb1QSPrQIfOUTomuH
O6rcD+VVSq7ar9cKaN1q92zJMDrKNHA31H6MnXNnlKuN8r6PM78aj3TiGUPf0DLVFfELJyPqBx//
nCg8QZls3FsYBqK4ott/x46XmXG5TxpzYGqQJqtSRQfaYiW13dNPpiy2r0efZ0X2G4VU20rD/h0j
KPPayNRmnn5s4bI6INRkutRGECZpDSMKqVovoCPbu9y7DoizDjdTmUTxdqzCDXJVHzx1ZmM7t+T5
SmOLbP2PYpCsw48BukdEelPXUSbY1QcfjrK/QpXJ5uzbBgt+18Z+KVEJsF/zK1gwp8YdA1MULrpq
zU6TxDBHjczvxg/nuiVSi0yaEWEz+IAMnZuKxyvduM5l0UGZDlNZe3Q4PgPTsPSC8jMJToYE4b8c
zexna2Mkhu9BJJesd4BPNbiUiiYMLVyP+xls2KLL0T7U8LuOspIqN7OQj6h2xia+UpnJ7xEsBxKk
IPsebPcIItRwliJy4CEJlOAfp6gCDJLWU3KfBlQ8lS1smnD/+nQjbZP0K1oUcCILH3WQAztuTCyz
//ElHXqlaNQR/76KjZWm+gY4SQnUzn1UvdCNDoM6I7p/JbbKpVFUV9G6SoWy9Or2BhUTvCnp8pn7
amt6aY7LHvr32NFE04ENEva32I2IdW3h5rH7YM8gobizdWi0R7oi0Amn/5/LJGrGgF/2UhNKabCH
9isZhHMX1u+AqxXHnGAr+KGpMgWCq403LEc9zzoqRm8pAW8mqVQGd/6PMjiaYM5z0zKQiKKVJJEW
soPsKB7k4GJiTSaSj+Ighq9XxRs8QzOMv8RxQRKF4wVwSh62lZuMZv+PLfJzS2z2+AA0t9pbuueJ
mqeFMrdwIyOeoLteg/lyCuQyKEBeRh/kbpgYRar6avxO8Ljtwf+7tcMdC8gHSGX8KZpPP2SMzlmh
vrWPDdWyS3ulakthjx2c/4uE0blBqRWYZ89vnXpDr7sF+U3ktq+1dl1wIejsu4VNISzFPmfm0/2Y
z+tJRDFzLmVQSooRT2swuZGt0hHcs5cV52ukjwg/6vk5w0uSuuSc544OFAgMdH5vzSKV+kIGAXkU
clV88fQWh04HRgNsu/jK3Nx54nwkpK7ShYVtRy20LUXw4d9TO3xmNXBT4zvkAz6gDLobtWbp8ZrV
fGUP1odBT5sGIxmIpi+pI+Ngkpasnww5e17XkCRlrA7ZwLxsF1epVoF5sSzhn54hi5kslAd7pyoM
5+hd6nQPn6PMzWsj8+MXV/TGicGjThyn1StkitnzNjVbZ+hzXXk1QJGErLz6ELmKCYG8DKiiPgQX
xSQ30otm9J1+sKdvbgI0Pxq8MjIfSWMRqfscMscGqHhuee9K+LNp4hkSuUliC3DhO7doVgH8ZY3z
3hTwketAzFglmn6TXG3Sa9LI9NNoOQXgpd6SBE0Nt7BOMQZKoqGIFfdPfWgJ60W+bl8Ry9QjmqN7
RVdARrSOu/rTCWmpH+MCESEFimpI1iGhKJuxvU3egbRjuqNDZC0NaSj8K8kfShsgPcf3neWgSnLK
5cloCIjA5FydVELNyWkDJ5BG8+LQRTcdDBXAl5IzD0sDhvfsHppdVIvD7uRpu0u82jp/JyMeazBJ
8s4jJ9W43wd3YGUqb1rgMuABMloJbr4ELCOpM+T/2Yo0MUsIek3Z8GKVL0wek+cdRH4BlpNXuSkL
qWr4DBTuPtKZlMeTgEPyWerUY07GKQ0eKDysuhzfbDM2tjW0yAP23AuaETU8NmXOdtXu2Pdv+ndt
cjIs///gqdjaydUUAMueUAbpgtBSLB1h8YfLP0nBn3yOQPq1eVqEf4cVWDjGdDn9OL1cs3lT8eTB
k06m/dxdS+x4HG1SrFeMVKsd9dnNs6VlXXWUf0Deke0U1FQyw1giX1bfPFSDcBV6I7ckc1LE1Zlv
I8BLyDsSi4Q/r7QamJ84OO99vrJU0OwQQC3uxnVcHg/SKALJS/zahuFnysloYqbm8wDKWTVUTojW
nFgqOArCsz4atHFtIQm49RdXCS/4AZccxEESsZaouAeY2h8qeB2UAl/4v08czSLlchMTEMcnmv2h
dC2eqaSSooINKipiTDTFV2yBOZmj/cCiZaVl/CTv4lw0QjWncXxRLpsk7RvuRwcQT0ArX1UoRwYT
nZWiFNVtA7rptqnvpqOCzujh3bIJiYrnB4wZtdYtpYJS56oBXwUgIBCwj9ecqjsm8TxCf6XwjG6a
73gH8s0d7KSWAUwPr8H9UqSbN1Ygenxmq6ADZ7dvqs5xKiwtE9oSrAB7pXduRaobdYyj9vlRtG74
Lo9MUzT1E7rmEUMNWXbGUuUBIPaN2ok3yUQr9hjAARVjJ/7Cjxg8cSF3Vbnn8MXyJ0jCgPFMobN4
+SzljKPWZ6ZyRVQT6qWQM77RyhP7ZmbkXAAHurIYuIsQPiTRNJJ3PxQDOdtV1GX/nA0Jw1Ctm4QG
4VrT7rcoFB3EfjYWfkfaeuL69HzcZi6TBCUCBGAVe3XH11ar8Bv+PHPxzB19uoIGsRFLtwcE0ZAv
v8nHf32IrQcaQYP5yzboln9nrtrgyQ3Th0y9qVknXOul77Z+rI6rvKi6J99xTqGzkmoNbJUePe47
XxpN8hhi3+Vxcb0kLxuWSS3XsUBGryU8KxwQlGBlEw7Qil7C+7jbszYgmuuhqGKnu3Z9KLsUTrFz
EMPtnV6xowFFfd31kHaOO1OcUJZIpA/ICL6hXxl1p6YSeY0X2ZY4YtZMbhOeNly5kiZcHF7tC9vV
NzHH4TOufHrr1SD8/DyBCuKYY/uCS5sRqei5aXSSBrowTUSgdoZc5AJAJiOxaooX63GwcGO2gOJW
jAeVAHayiyGrtgGCcCjftNOTSDJn0Wg5hHJCeXa5hylN9s/Rse6B0OGYAl1qsyHTpfEeHDqQbkjP
2AeloI/Ja8tOZjxtXOG8fjJapEgA5tA262iJzYPOX2f5YZd0gjf44MrOfpnT3+yQbZaKzOKjcO8V
ADSDe4mZSa0+bVipQPhuDWVhpCfle416jm4twTbla/CRfyoBSTN20Er5jKzYAPdEec1BlgT6I2Lp
sX3IfttqpMWfBo5zM3PgUfN0Z+pCZm44yJYP/XRLrJTOWRSUYdue5M7lhJTeTcofU9qPUfv2ea3o
XUX366Kcw4TtZYkQXar96g69g27yIwA8clyBsHDzKc4nvTppCUT7adzuGah+sgNrlsj5ddqrQGlF
29Q4hvr3Hj+ckcczFoIk78ItX9QxVFt60IdAfxWQauz5McoW3vKgNakQO7UkfIaBv23IqH5ddSKS
EUydxqKE9r1nM54R6TnCq83LPwwRmcwboZ4ZKPpKsygIBgum4Vg8Dd3y9PnLbKK0uxhGnK0RsURP
ghFjZaLdtM9Q6wz8ojK9mEJIKWglaKhJPZax5q0+7Z0t0UGjfmB4jkYG3uXbGrDoblBHSVPEWul2
kxZQKBbp4TaogM6qr2MDi1U8f7G2KAhRCMQ+Hk8gfbsOPqCeDKV40V6cYe9pBZ1bFdGhVkBxlEY1
59ezVf0i3a/p4RnhJrGGv7oLy8+U256TM+vWnPTnLOe/IXPcVoIDedMMdbemVS1oCEqm1RJlxOCE
voOkDmSrSrMIna/yxDjGsQ8Up7OvoYyvCBOGjZJJbBU9d8LoVmE8v5mCKPtasPBzoB/cQ0x/RJ7E
9SHTynXy+7EnA0O0v6tXGsSDGQ7OZZrY3gbc8waPhewOxTLwt9mUIsVsdjduvY92rBBnd4OASWnd
qLsl3dM3NwR+vDGS56YocZh710989LOxjgVEywQz8N3xLto6bPy2thbY7hoxoHljgDl2KYj0k2nS
Y5iIucIf49UgczaAta4GBDFptbdZRfkqBrq/aenrMAetPCh3OGhgG2BbMYgQymukYhvu4w6o5oX0
Gzc9CiS+Tc7v2bduOjdRxAsKdJl/SfQneGwyKOdKMd+QY+m3sK9ubFg7rc9ZB7/SKbOxF+HZeCdI
ocqezI4vIxgQ5saWdI3+4YrUhs9RD1kcEOETf0jsM630Mr9CeQs7EsNKkdZJ4hr/1/i3IMVcEZin
O7axDZAB79Bz4uFP+mR6WhGxna0DNb+BV5nnktWXQKSxpusi3+sdLAEdyXsk+g/ft3hecX6kbdMd
t8YjCWYXycC94qDcS/LaA0l2gxnxgDcM7UyQvIjzr5NjdlyTidSeng/Jwgg7UnB7azJO3nctdOJt
Ul0/p8Vb1K/Umhjbp8hOfKSUcHwdn31dVbwZp0z60rJoGcPOlDrosiK81SwIetD0kcV0bXU9T0bY
OyibsaUAOsEu/0pB8XUvduSbOqJ8nTBIVTXnSeDPrh8juHjgtZPIJKyk9gcCcj6oY447ezq9Ib8U
U9yK60EvSeePyqbL95ErXEZiGUBJKkykirf2SsMAEh2UeCCn6RLTfFGLg8prYn+Qe6SjPVB8OtL0
btk0HjM7SstyFeFp+YzxTjzfnt1WyT0AkUTC0e00Ut9nftuj6BlnPJ/JVrELyHnbgIpWV1AkSuM/
0GEBWG7zy09Yr/yW9WnuY1snbb2vPfaLQNDbRbK8/kJNZ/rBQs9atQ4v+/hwImGSt+5hdaq4CLwZ
7lEB5XSllrjg2+2dxKFfTgEYbKMvHi9oWqFDTX6ZV89gdiwNkYpbhLBWyE1bazAagwekEbJ7rFQo
8/kxFOGRtahN1qXqmQ9g4aEbG9Bx27Kmzi3hynz8tT+9ezIug0+UkxBak4K80lpkECGnKWSeQvE0
jdY77IOGUejt/IIOvJtwSLHt+PmlX8O2EJlDymzrHHTlevQVT4C7xu9B8yqynwryUbuo9VtWPIIV
HyxbjsEKnIcp17p4ny6YxzCv4oL9CfBn6rH5vbi+wfoVBYR1e9gu61+gxr6xYpxXXOlm7+wOjuJB
/xA5oVLEDohBEvEgHa5yC7bcT3ZC0lFlAO5ZesdOeUa4dkGx7cf0SNcsenIFlKLlJS08AhHuOjAs
pf6oD1HlWBtDQTIUteaajD+09CbZEiVGfPSJZc2Yw8+hPtN6JryAdDNdq5kcK42cTzB4glXI6Upl
Q45IGPDdrq4rWtEWEr+JY4pBP0m97gHbJQeCwnJBqAClYELXrc8wnj+o43NpCMwZTtj9J+2pRHnW
7k9MeNTPpCN2y1tpOZI16C+e9MwG/BPnvdQfcfUIvRq8F1n7BpDINRtflnVlpCN69D8QtUzNSg5F
FThgeN4ZwqZ20mGvuhflwvA7DkNjv0g9/mMIdPbk9LptIelOA0JtSrFdOmPGLSkj4xZgV0551FG3
YtoxGyRddD21gQ6oLi6uUYHF3fwFYrMsHwLTNdGDf5ugd3/sgzzv+CSbF4cJd8Jy7BN51PYaJ9pa
ywuCArTUchW76qtLCgiFMTPtQ+Z26XzIVn0RIOBO+qtRYEBMLV2rlCDcQ8yk9z7wNJ2UukKHeSpO
HQphdTbv8JWIqD9tndXOLA2iAgjXlhdcHG0+iYF6Qg+L+nHu8TpOFBUkXZGU20aanfGM99blt1/R
T9VE/m15WQzUL//9o1UnoI8t/uVoUhb54lxOEzpmWCZ+jIV5JUPU8r2Iy5DXa3LT1kKBEs8+QRjC
bCoMhKBIrVa/webgUOZSwNtoXRb9y0+js9/qXixOcdETKvHbQbVxvr8x6O1CUBaIP35iEBY3Hxfx
i2iAuERho7qO5QJmP4yhb8NSUmbNAGhCP+4jDk8ZOTLQaHzgrewucYDlpNYNAsO9OzvSsE+clFe5
UKwLTrz05CiH0Dt8byIlI9d2+4IG6ZRFl5oGPhjRflFIbaVAInh8r0YnL2l0WGOCJTDiuykPYHd2
nDugd3z+K2VSFsKpwLJXt8xywdPm3k+tAvdfAyfn4pI8JKvYxTq9X0pNtrN7j2AOh6tR7/PKI461
pgyX3wlQNl9oeWcdI9KzYdYkSGcjP7G3gL38eJkUhpjTp1jGhx1Q2I44peA7n29mbwY21AbhScKe
57TIyCjIa3xDa2UXRIgeRVwCHjhSqQLVWoShEdGmlGUMrxpXQ9FpiEXaYGY74jis7h7586mBNR7C
o1L/I+GnVjtQCvtcEz6vSSOheITAxf9Ci7szTz4RIPtgGSc+uMBSWbmd2zxeTgI0E1ma59W+OFSl
SD5lkxMHI4ND6bjrORXkcdbltB3JxydRB67t2Z1ziBTvT2kc7Teuv8ZFW84t4D5xhEZONcxyQt0A
nXgXJ9kG2ufqASb17M4M97WqKwW7ggs06FjGPGub8fcAt+SXXbn0fSB9giomapOKb2M9QKYdRRgi
LgfL3nslGFjEKCGxeprjGrMtwxlALD5frQPvGOECzcSYxZ8ngTvoGgMIaLjgousvTrry7KPcaSuK
CWQjrmx8MnpWoL/VWYzlFUtp3GFlmh3hn7s9QoqUB/5MxafWtEPbwRW5NqA8kBK/R+ujZ9LSMMFX
ukMueP3EbeZ31CzhcNBwwtWXjtN4CE1T0VwEenPGGQoJbc7ODvcaxaAlI/z7A4uPkpiaH3iW1S94
ba/klpcIyY0tRijpGiNAKFoPLLXCc4R4u6MzxOH3LniyRzGllIB/6jiaXJf0+u3KQoksrI84MUdU
j/SWr2ybq570j8hX7zyMwvpEK6egPAPhmOc5WaVNvg9ZjhdA/cf1Hokig2DRgREyO2H57TgWaC81
A+qUwSc9B14v4o8R5Kh0kMrul78UOydkNXclo+Q3ftiHb3OvvS9T3Y600DF/EyKNyTRoLq/4x86h
AWQDi/WGrb2XVmlaIU1cH3gtiT4u+AYN/CUbU8Lv8ywyc5Gwfd53J9HOjWTp47ytv+QkmjrgG8bp
EXGSCGC/BhEMSy/aRlKeM5CRyCmhQi8WrGuaMSmdCOoAgEiesA9ZdFe205xHyblnuF8YHLvfi1d/
69vZeBzj4utxwPZKRZu6U7YM7Gv856Z2cqwco3OjtXwmLaFiJzOjq5zs1fivo2UJtBO1OPe+YxbV
Hsw9pwpT7lsmxCImWd9Tl7TQmwdF1SVmVnt2rRTJmHNaeH9Khzpkln1W5ZvQ1LrtAAnp4sZbZvbt
HQ0nnu5UAosEvz2PJPlY/b1sWj5j/sPTbDUfRYvzX02PCFENzFiH0sjJtRQilVRDEj7jDUBMdCJ1
aPX5IimGrbe8EEAxTqE2rBO3MIaKiOJ5UA9NVjd8Gon8RdwWvJjFvFmYFnVFVAQ54M4F6GySztJ4
VmTPLvYeUgj2NcGTEzU2KxdXdOoEtLJfpln50b+JxWmZQsG8xepqvO0sePMQOhEf8lb4WgXPrpc4
nyqxiiGtPqYmdlvtzN9YpYDPtR1vWHvcfhsk2kswnnRP9hNU00L7TxWqxgrFIGePqjewV7vIo09s
eoADh2gePterAjJHt0aOuDhl64laEFw0iarXlLYdYbkzT9QlZVOLbVNIK7keo/J5Hd9L6jIDYqG0
OyYMI+gi68hYNTOY/llaU8Ue29fui6vCKRp3K9zAb6SRypkAmVA7TyqR0WU0YSZOkXKPdgoYNvxL
zeL9l1UmEgNYPjjPcIQREYIRCm2EoUDL3zyJBs2z5vFRvlTT7zYmIR7rjuMaShQkU9mzFemjWhsu
7FkzMmy94etqTKgquA9541sayCMDPt30rJxVX0ej12D2cuQ94FSY55VNyoEXz+zf49BzDBsrhiKo
/0EHlIluURkgs07j19L212NPddLlUMJl9gHcu2NBPGLAacufYgdRgpAfrKb6PQYi+2u4y+kfrXJz
Psgm109LbYK4NbGKkhJolXuFo4/p0/PLnOk0Zq+gqmTLlR16DKmIep2MIE/FUyM1gMWwaJG7TtuS
0n4PqdXRrfzMZJ+5cwntHjbb4XF+P6s+lqlK+5M3w6GixkWrfaqj4AafPsPzBLJnCZYQBzTgujLk
tBj2sbxJYy8UZ59HeYcizkJ/Kn/leXf/1c6/r5GIMbPdupWhCJkM0HFFg2oBhLxiMRoYzqJEhIoX
RRxFlKyJ/A2iEUULTO7klclo28xI8FHIGAJ0HRqablhqKAC2KhKmwKkltj62TVsW526atqEBhlPo
WWsnd5/EyqI9/fvaV9zFK9TSouqhk3vTiYjtdv5MeyJjjSduuEbCBqILWHnMjE2NgMeVXHmsAcaE
TFaJYOIMdiZntCkObdWE+VRdF7hXRajfYRwupkHsqCjh4kDXPpGvnQm41sVTkFGvpBreHsqAHAmC
1g5tncujsJYHSAQLnPMrnXu7risab8u3y4pQ2ADEtSVPbNIRtcOod7u5aF/pZKY+m0XkC6X86kB6
vwp+IQQDHIOvULw3jJQzflk/o5e1pphLHHjZ0Yu8n67UzwMA+RVS0FifHXQiyYieADjC1DNuNvTw
W8ennJNBkI6SE7dWiqFR4dctOQ7jks2P0UXcRnhG3sbwL3xJbrMMbAfNMVQ9LnTBQ/kSoLNTxbry
pkItOQLvb7+Dg1S025aimfNNouJV7Doe38OLO2IsX8/hV2hsfkOWp8wSjP+foBoV8d52W8bUGbc6
JlgM6rWhBj2vL0XiZAh1H+kr3mdIZYie7nODa7tQlvaclCeM2UgOChTjxxQ1+ot7B5vbla4DHYvO
NloX9ZoxJ5GZ1rjwJKUQv3Hdhu83J3wKwYsQV1niDxxFVvoqFsoGWfOx66/jzvSSdlJ+RpkvyanX
dw7BsGPx+rUKGYc3hNVaYy89rFLHFMaQt7bOOPqlQo8AjtAhue3UKeBcHm1YpFTe4lcrpgJxsYRn
VZm2f8K9Y3NwOBFN+xjA5Pa6yGFonaTLinPrHYtg8j1MxwSgaLFQmM/n3qnzuIk1/qdOF+NQP9wG
nflfrantLqF4MxRZ0+oxpNQ0szuNDGn5sWUd6wIGrbOy7W2M418m4HlRP4r44TP0zp7neypaVow4
m6/DMYYKgPd2yQTNPom9iMJiRDm6WWBRmMKtQBPVemHUiLsp3Goed0quqeDIgnSVWAop1OsqnC+M
bVuPUs2pLzkA9Z7ewwjRPMDV+202tBwCcaH5qC+qKfVl9dX6fsuPrWKW5gg4SlwFvwl1z/KoXe58
3tvoQaRyN56pWcgzs9CIQPdHpAl0Mz377C7MVvn3oZkEB3987+QNxKU46Ign4ssxTrvoCa3zVWfT
UAVWuhjqJ+r1F9wX+txPdjGHZ5TyRpvFFXanDRCZlvql54ZUzzxGgin/Ur4rGMLdBddDK1B2eYuh
v/zR9CLjbr6UJUI9QY/1eZE9tBieYTkFFR9lFvHYNae48kj6W6JNToUwz5QHOa6Ub+L5i4VzmuUz
0LbNgGrguYybdpg2+mUPCjQG1SXlN99qLLaTe6De0VOEu1lSb22qz4b8DCWYARSzq54lZzAIdagp
UFVVw7s5gs6qtfI4UhdArNL122VaJ7aJdp4T2xWSTbnFWhxrLdxLw3KjLoeOZkWAQA80vnPb0rfV
AAPBD58iTaxRI6MAJobVBObLPEXBKrr9xYL6CosRZi3mKY4Rxx6L72rGLN2NPI1nZ0kaYnKIyTro
T0rnPYVDDGkH81/6PgaAYD8PcujrVtli2oybVt2WsyrOWQ5fumnX3DVqDlI670iZAZ/Arsjdt3r4
OpeAMnn4xoFTs7ZdmIW0Yjff41HiJTWsnQkU8yAXigLJcDC+5MeypqBx6aPsk9rP5OwXSjnmD0XP
0B4p6XjIym7HZEFyV1b6aOP8onAeWkdmCp23EWtBT6WYXRbv0Y66tqrQ8alLkQD6c5ujcANv3kqd
kHMBYFjLG7VDMkYnMNnYbQp4fMA6s84LBoriNhPGl1emB1AZAaohWQhta50Fks8QMkxwPIzJt5YW
964OW+m/UyntE+4kI+ppT9eT14xkPlm1e+chv+of/BxRKOcAa/pfu0WlTegQTwWcHopzglPJPM+f
gYUKRld4UHK4DUOusgx67gqa6D1tdgwGdup+0Fzx2MvgaWBtC3NDIYfNKDqNcOiABE5AbMJshwp4
zcN/4Blz4ZQgMa/SmKX9aI5Pc1XUnkomBSu8iLcteZrAUjDCtcFrwyGCwxm0whV68C4jzuNhlJUr
Kf/FhrGWwsC8OUh1uCIR9d0qFCs/YMb1XObgsrNPWHg3GrKEPEEDoe3zIfLatsFTPEOn71KJsUYi
NBc05a9t+tIH3DJhS7WIU2mjHJCTPRQcz2W6CCMMpcbnX0R7BavGHvVemQfhJu8TbN2kD2HVzcNR
yx25ObZNLWsKAZ/ekw5Jwg0GIrB/XXPdT+45ZBQV4tNajiGRppvmIek1WQRhTAEQdhGsMftSNgkk
ct5UEIVfkmKP/13GNAUrahUd6BDNTOUZUbd8GsPUabO9XcCBepc2CKHft0rMWUO10sgBFZOvO+b6
y25w10hwQwA4pLoHEXYr7HEPW+EqgW/nrZMek4PaRkEIzGEvSh85Ynjxn/K51Fgz41KnY1FELUp+
FKbU8xcIq3tQ34tgYlB5Stm5TOJTbMDd1YnaOw4gw87SYnoK+Kiyp0NV9DyrPjgRMMx9x4QrwjMw
jhKhfYtvVEt4h9HOkpAFAyk0uIcUX9hDKIplT40p52lGdhIOJ93EHm8HN3I0coC+TaIIk/foefzM
5CGeJ7V8tB2ATC18vs75k/3pS2BTtbFwKEXMI4/nnkQjFlmhub1OkMlkN2ifjf8oe9QkAUUFhc2I
mVIHB43rMooS+J9CE4+KkLvayYbpu5XvoWAwKaLdVB8D6hZJ3oJunbJQ51vvisG6pEFl6sErJcYX
teJyVLb1EE4SFZgjrTxSw2py00Cd6A23KeXEtEGaedhQIVNEV/CFfo8RxjtKeCCDsC0GB+hucbWw
Id5gSnj4Ty6oo9Nmte7Q9PdusI0N/zlEA1y7zxzWU3f1zXHQ+XxmDknRdcz09ZMEa/SzlDeU5t94
r7Ph+4s1h0MAWlilLZgJc869x96L8nVwJBp9WzJF0SUlLdsRDroJ/TaNt1Fpl0/3XXvodv2DkftG
EO0VqcRNoeIk/tDYtsz2ZGrvVwX4wydSgjxbj9c8fG/Fi5WNJcsIXETyfep7skkfAFRo0mF5xFEs
FqWJ7BbuFJoFnnftJw+UP6EtRjY5CBab8ybr+20Kq9KXdtX+wbfD8Sy/BYPkIGgblOszTy92p1qq
sOVGbRHhYxhLUY78z65sQKQerFDA9Cjpulp2/P6QFnU2UlSB4KIBS7NIvvHZmB2jPYQvp/PGD40n
E7D6egbp4Fg18fVVRuOhYwEu1U5JJEHy3LqKhG8NT/qjmYni8YvrPXgrAFEoneiNBJjvDqrQJa48
TribGEKvn76+8jU5+7Lapn/VzrDw2CDMW4PLfFR0qYkwyh0v10pwycgUb3vZPCM4ziJ/0o/yqygY
j0FeV/25cYkedakm9JTIjKPPQ+tyJHC5TJZX90T/Gih398ybkHpsNigW54QiNlAtXH0wXKT2VtIP
nk2ZapngGG4AQKnxTSDdbQ3YWKxriObTrTNtO3/ZnVB0TFabc+S+AbYk1BO7Hq5kJG5RSR/+BFzw
cgxYUMAxFZyXQr5ZqlARf4sDXvrwzbzco+fa97e1/cnCoRAXo1IZr5BBfdB0k38alWpwJdEfiF01
Hz7naAUki1EVgdAUuYRXe+fxDaqMwkzTqx0/XFApP2ESK8zCNaj5pedYwHqnVrzqPm5vYi1WNvpE
Q4dCQ7z0DEdqcoxi/PFkjttIULvML3x66LalFk4hHcZMnpJj4mLbj04qv9ThUiGMwV3E3xpnRK8b
I8kwY6XnzY/9118lWkGYHrlsohiPO+Dubm1BvOK8NcFbDM/l4ZCWspTaCfRx85+2Kxn7qqincE/c
ARTOACEtDymZuZTS7Evwr5oBbKZMlNIcZyOlLmYnyugqwvPPHcAqe2tnQXP3sl6SEXsmukADu8UY
vLJb/W23X3YHDOSGiyuKzEy4+2h074e/S86V+HOGdPByOIbTK5ioRtw6FjFinRBxJCjGdgDv/G79
6/VP8RPVOAo8tghRBYE7Ng72QNCgRB9yQceUA8c0Weetc6usoh0/ZR4phT/jBIpe5j42fWj4gVK0
rM3B/I7J/Y1e0delKKE7e8oqIXgGowo7T2FInMYnIDv0hw7IwQqdntg9QVtZonDN2fQ6zWeaa9LV
LTdn/5xMnNc4kOWun7eB0Eane9qtqmipeDoe1XyR+q+hz34iFN0A2Quow953mwnft6diHKGgJUlO
Bh0rBsEVH84DRSgTmIuIkhyIvV12eHPk24EonROXUtpFfgeJxVt/9CLPnKfRCCiHQ955MRAg1rsZ
DIQdgvC0UkeslR49RcCZVv0+Nv57HAdm329QD6K8aJePSXJ34574v/uHNVrNQfz5qzYIOeezP2xv
KVMXYtKr79CgM87gmi6ShejVN9H8Jpn7J8tPT8WUdeS4JCqjPUOaCnAzDp4igU4az/C6R5gcqf8G
b6fD5JXt1ssjaInJczDegG4WUmJvke3yLOj674/9GCPxYN5G4A7pEk7Z1MJjoLjWc89MpGEP5WWx
KAB7bRfCtQrV/1xpFUB5dc7rbF+TN2Su1AJJT4Aja6/Z9IK4NBeBFOXprG0WbrLg+nG4wGyw9cKf
gt258myR562FQUeLpl51gjM8zCf32l5NmfYPGUqssfsGdPj94767T6/HpSfY4HXMBZ0udeJKjzFu
4spNCz2s1OdINq/38aTsl83q13kzufnXjMPp8BVxN5fdyfaMKFzGS+awpb3nzCP5eq7I+zyLLBaW
90Ve9bR/jn/e0fN4CAKgK+f2E0Pb0WrBVTEBk6Jqn3kYUIo7iNuiPPnQGycG+T9BWDhsj0CaWXhh
31NfkMSRGk7LtzFFGPRyEGs+LW6rbn6PMGC/J5xvYPcBxAxBeeeIjfHq3Lx4UR6tKyK6Um6ZDvG3
LQg+jHTt1sEevHiZ/x6AA58/yfh+6Rpb3/x7SrXgdDpnv6452LbO3DBQNhysBTpI0VIXZkSfqElz
FEeXPsklQUify76F+44kqEHPvBy7++tebdAPxX8jE8ySSRKbWfuD//O42Ym3ZcHL9LefQFUnNS5r
a/2LGh8K555CXvcPFZemgFibr9evqLpOkscZqT/nO0CK3Heq7vbCWQgRxaage3jq+8BgMs5M2WSf
kusJrsZQLtnlZx304n2J4Ap1ToXAlw4vwHu2h0B3wLsqBKrvmML3YOeCxjbKZx+jMio1lLgvCgKM
hPhA53xDjWW19h/c8nGMhE9dErW4yH3bTzUurWhRouJFBAaMR88AxJ2t2yOgBYE1jEdaRvZgNPe8
PsxTfHcwZMZ1b8Ykc0djdWi+NWGciP8KqN/LF/8UhKYOwZ4tpTKAmJYeFBL6feCvtIRQ4sB2RetA
utqZtcP+sJKYJ9fvfaPrvNUIckzyBqf4bbN4XPBY/EcX65TVTwPcL8XGrSV8KiJ6BCQsPCSvF9Gl
0ITdPhkyQ+7mFkGlnjJ4iK1RX4Z8lm7Nslr+eYfwewsgEDnX6050P0xtjDsB/qWS0+OqVM+BXDnI
gxfG6RsTzf3KDLYlfaETt8QhskzIiva4m3+ZO69L4gwMHx4DrpVgnwidU2VdPr8Qy823fxtaGUQy
vyKUOi2czCQ0AlfCwVaCwODn2OMTxE3Xj24qHeWS3sBzwl6nmS96J/nW/QmneAicPB4LWQ3WAf0V
sG2cBBm0ZpnZR/Ua1LUSnjHFi5kQpWUUHfwQG112OqdvmsdUnT2l2tgWPX6Ihr4BVmgv2olDQtLp
G8sYIp8mNU0wRJSxlW/OZnAyA1y2MCrCKbD6+Qc/oDx3Yy6R08fpnPvyR7TiE0VCAZ5u9FOs8fpp
LwBkXx+gu3XsUwX1PxmvZxb8V4zkUzaiXr8I3C07uti/SuTkzHi7LmHsURRvIMY7iEc8W4l6WQB2
ca94kcdjo9ZVNeHSyM8PiOtGtV3+c4/n1NxF1ZvQ+zS4pao10llDs0FjvRzgdG5Wc5xxCAJ4lkV4
hbGr+IghF1VSRsrAttow4U97e2kcCYf+WsgqBQXBiRB174mq7t22sJeXXTcD7/FTM7gNUYRBEAP2
nBZw+IMtIBe1StxgQN3a0nhTbu+xbkYqDGubOmG6iHluZ3QixOtgjWVtOghoTWI0YjKJm2jeWyoZ
go7pxIzIV9HFRZF7mqCu0UblhITHLp9pvdzd+lwhmVIwIZcTOyWlYTsFu/63KWkaraOIXxLG4aB/
/Pp+azSmfy4Lb6FImcJtFBhe4mrFdGxaPwB08QT6kGjuWoE31GraNgAf6OgvUXhojFRCBnOAVBRr
MxfBqFtn7w3XJb8R5e8tG1sKi3nwGpNfzI7ipvZfVw4Em23wwZoF/WQqCkPIfXKDmusnAV5vhJhe
bbBenejkxjx049/X3FmiirVaR3Fq96DsNqMpyFiu5k02dg2Ymk35pEsvyHtj1BzvCf1U4MnwnMpK
UX9W85E0KYEbuiPTXguxU12AEy74nhnbx/JZXA5oRNOWRU+ffxuxSD47qCBsPMDG35c4zA7HGVmQ
FMyFPasEEOcOVPEoYwbXm/0gTQzoficptm0BCmh34AcPp6mlsRDjj4rxAPOYYrSDISk8VUBeYQyi
eRExC3EUdaAReJlStfUsjCeIDSL7NTZjFwH+DwJDovnU0yWWEc/AjK+Iux4Y9+cZQeGm8V69B+2Q
zmF5nJnDlFtU2HpbQ89ATJamnVhsXeicVJWmRiq1bLaWRADZ1xviKtp1SnkkFLqtM9+MA8+lBVKZ
nAW88+h1BFjMvrJLMpLQDMr7Gt+iCmhnp5aKQ7bquu95kt/K/b4xyPjS+PaKShGu7CckzNMiLjL6
q8mbglSf/dYZV0qhTlQGNw/niakSknMQXYfEkmccSjYpjN7D1GtJ7jzvzlY4Zy0OxL+52maQcXTI
GYixMtCO1gAbxm3gcIL7xN7oq0fbFZr864Bxvu1DP81lBHo1BMpsmx3BVuwn3lMFA6Wf01bfEOjQ
eUU9msAg2wi3ocveESerzEKerw3pH6aXmeZuTkU8SGKoPzN/nNseUtt2MF4Gzo1xewQEP75EDzKJ
NQ0BaHr4Jhe37Fl5UfKmpauWMFdkWjWbo5bmrD10xguOUEiE1ioZ7XBfKqwdT1YNSp6c1c/4/FGS
pwHE99gHftj14SYGJT5RcUv/5TDsNjsurTAOiz7CdCzLmnnr7FSXQCk6mlgSUvImTy90CYnfomgd
8M6IiJOev2jlk94YrE9LeY4XfxQS61/a23eHtrlfuAwxu6O4L1zoUFbgWE+kV+bxnTYElBDnq5We
Gzm2r23ST3IwZejGv8AGiBKb4yMZ2Do6q3T+QfNJcxaY7cTMdR0dV03h4nlu3cbol9B8VHLhD+fv
0oHxlga96p4Ou56jkixqsvGhxs86rKU0ikaQmzbBiyuu5Cn7Q8STI2hsDwPsTJxJgVJm1T17nGLZ
bs7M6p5IdXu6ga/zriuUYmrRgb2DCj1vUVwlhoNMFpzKJx8d8Tsb87Mj5QoFE0K0WcMk3J89AigI
Q1FD6N1yyR+ALqCKYhG79pJ31cEYezTSlg9KWfOa7G2geX6g8JNT7VP7naeTr4dpjxX0PbeM/w0A
DbtVucRKrBGy3SVfYLDkHj8ByG21RXLZuausqDyJ+RBhwcgLkOSR2epZOrlfIAb33sCtgv2LS23c
1DuJFIPPDvduk0McyyZ4zeOKKsE1L5G/asrDF5ME2l0AimHBV+32SmWsP++QZ7sm4TKGPqw0qnu4
g5RQrq/GOc52WywI6PEBEJClCSNlq3M3UEyS+lLAuY4ZdUOTjwiFEoFjulQDFS+2SMb7DdmDsJLg
IOGf2IttSe9E+ve6+rJ7VCA5XWIOYL4ZCDM9wOkCVcxWXkLa6nchFP8NnmjC3enayk+q/99fb25F
zzU6vHuW2ur6+Ui9LWTf9SJfIaBusovBzxA2fbBCeuNjvyOs2BfcW+xv01NIS9Kke4tiB0KeJReY
0PFs+E4RQutJKLl6pmOkFVLcOS8dGEmJMn1N+zK38JwqGmWXEbAQu6etBU5CsAXUqDGNapzfoAlr
iJqUIwTMHuY97mcsqAWShyWH+pt+YiJj6zavGTKqrgjj8dZ6XoBYOIRtyo6ICq86q/UVmGtsG1VC
jQk9ekjni/CoJlosWfciga7dpqTlGEcQpMNuHIhcdU4uf1XCE7ZSVLOqLOnOAJxfE5lkd6QOk9OP
XcaNZdiwfdWT334Xwn16/FMuKICqJCHnt/0BU355DXys0C4mZFyhH70ExiFeBzhf1ro+7NvylUh9
BoVTqoX4F2jo5gTMCyqpr1C/vz1Z0nsXDcysrCMbs0LSs7sKRT9ntC92ixlp47lhndjBTIrQDF9c
zEOUtnwc97HtQyg1Ez7v0O3YBgdusl8OuUw5I5p2I4CeyoKRjqEPBwFP3vEq0gFuLQZUMeJMCToK
hhfcLlvqxfqv1GklnPoNCXboK5pDfDYjzQZeuuZp4QNIdPT69rAsAMJeqxAqTW4UjaOTEo/OoSsV
asQUDKEDp3w21tfJOvU0oDVE0GFjQFBCh+Bh4EbNvudnhocZO+Z3ec/vbGAQjw7fjjmDoEGiv+kF
zuHV57M+Vc4U/G1ykzA0R3tWMwiU8pWjYLZRPtYH34tNcDAZGjzlmk0BHYzSPhCBb5c2zM/iO52m
DFQcfyVza/o7v17mCmDnF5kMBx6CNaaQjS/Bl2yPyaxZiegCd0AIQ4f5nxYdITHR4OVwgluoPOXh
TzIAnBZfQAz6XXUosh6TcVB0v2h0ngAGlOgOO4yuYmEpi0wY5i7ncNqwf5k4gb+xsTkqKuMeCQSB
VzGtN+V2lZz32jnsqBkR/hMFuvck2KkXIohzqjUQK5yojJjlvRZG8tvR7db8zyJRFIaxob2dvGOw
ep0ZtGeKwy8jSR1BBhU47UNtBlq5OipsgaQ+dhZ7HCqwSLkrTQLMZwi56+cmUNMY7Uudv8Txo3QZ
iAyWinN1tQu3Hw+pNRtW1iDk356ZIKqY0IBf7bghM/AEtzfGHfkjATU45VwTniYjQAAmtrRcPls4
rdsJ2dB1EhimBFS6Iig1M9T8GmwId/HRNl0POEEyHr7NRlNXZ1rO8KT9/t9/rt+6fYR9C5HnFH6D
V1b4rgwyNkzX78k713/dN9DfVr9e10zPAEdtgLyg0jHka46BxNFcKh7q+Zs0nm2SPF7UJoway2RY
NSgQMTd1lVBaKlVZz8mI5dqfOLjuZG2l5OSlZT/MW/77H7joV6bWa/xob8Mn6hoT2uhE2wMS/Zox
w525Izmxh+A6n9u6MQcAcm+SmYSbRSEua6r1Gz28M12tZREjBvV7ZIsZE4SW/KdpgU/8KGomtAmF
r1Mw3X9nuLuh9deSry5PRTGxyBBTMxL95lbpr27RnJzwMNkl8B7Tb9s8zHceslOn/pqAXX164x6d
NWbsFWa5bP40Eo0cEwmVDjXBm8HA6nWlm6gmX0WZBBoCwdDMH3vV5q1jtt7MMqQaF1ti6YFVwSvT
2hbx+jM5Q+xcU5beuq9d33WR22kS0XsKEbBA7slr+arnZGRJcHIcScJ+vAwuiTog0T2V9JoVVY7F
+s5RTAzYpujgrGJSwEFxnCkYzCog8h+IUZ8XbXYPV3oPMDd6Yj+9XgxdrasalOB4imYN4guURgWV
KO6y3P+kHdOWf5c0yIlcdBuWedP8f9q2iBs9TNIKvYQRX5NXVaS2nsWftw01iFJQNaXqX8SUYDWf
LBuS2VXQMRxppWP7KQukglxHypG0ewGuw0ny4+7NrLbkLYk9NCFiRjeEIhYjhZk+gv7iGWMyj0tn
FeTmPb6MwcVxaWrFHsB+ZIBEoV+Xz6/td8poxzzAqUuGy9SlOgV15zxDge3ZnuwP282WVB/hRru2
3Q5hJWxDeF6r4QJ9RZTbpfXF2rd5XvJkAj4PXfRKNaLfFmjgf8xZgs1CHxnSjKjq0P4fbbYbnCt9
P6wgQTooiNzUZcJlfcqmbr1gp2t6f+lsKT9htufFoTA07KOw/gXpSsI6fa8RQppqw5FnahzVCdfQ
yMxVPLl3jXzbNybQhydEzMd8y4Ue7d9HYlO8BKPwZc/AgL7ZEtljTLOAPJScLS3vLWl80k/gt0JA
3kGyHU+mCCwadGxDWSmOy4uM1fb+dbGQ9JVbxlQkqZ/4sMau39kXE8cjbx5CTXnx1ch5z81sBCbQ
zrHrKYvmHNqJAOZT6oCfCEDKO5QA4I5Ki3J72H3prpqxbc0Wobv3rSoledYlc7En8EeRU/uircfv
/EirKshoBi8MW/cDImmE0N1/h+o0HvADvNLoiyyK0l4SHDkJEPlb/RBWgjFb7dbIPU/7YeqpTD9N
UTp5Tzc5d0GntQCeV81ErmsTOSJXJjJuOulUZi6mjz8T5c13p8/EDsyX2Jcg2hTgu01qme4ebJeT
QMY2GVAXCgvdmTAn4XjuUNoQlNWCMOiW+z8xfRqDH0CtqS/WyEJDUrIG3nOKON3rKMsyBSCqQT1N
vM3+2COyZfBd2j5FPq1zi2i1zB1m74EouLySd739i28eWhOJXCovt37y6VPY+5Hn6hE9uKQHqvnV
/YltD9SXBWP7o+dyikaVVmTWPBKcKdRNva8eCqDB35R1GmMY7zdE2hcQM/LFwJiY5MWlLQiQJYWh
ohTkucj7xZaU3ITT7whbLEpu0iZHVHVMFSYnyVCDBLT7XoTvLdjpuMWJIHjC94Hkmo3uZGdaFovd
M3SqTwt4W5VacFivWheXtsUpEL8Zyc6Skx9m7mTRarvc2LV5wMwpk/2qEG8NVvXBeTxnZYtCf+ft
Q1JNRZ6SfpuBhw+QfKgV93Y9SvhVX8w+S6spUiExZ0VMBSP7oM7uUmd5WMIWDWX7bVkFZWfG4r8T
eCDwK00keNmgSEgmrCo4wBFbh6DKo4D47nOd3jaioXm4dXuk+2IfzrVaI3cz49r5cwLuLMrriM/D
xexMOnJUGrzq1rB6PrQQOHMpDuVyfRNZiBkrRK8kfVo/PfuNcSn0D8Vsxlkui3YYO3Vpy1qB+P44
/vzefdHdogq1coHUC4tmUy0XX+MDiswXAB/gpPfZgDj3QVFujttjpyjqzek9/a8BWFFsryo0qp1W
c3osEpl7U9kBTUjOiwPJv4ALiL1nOd5FG8kivr8k/ixqL8WELcEfzB8LL8DZTv5VqeFXTrMeLPdL
Jl3ldh4NtOBohpSy9G5J9mCkCGAZyVGzEeqr7ruDfUpCSTplK0/GG3kcTecOsTV1vWG164auYfeV
XNnEtWpfrAF6l6c5PkGGoBnmZmNdPGM5KLYEWzaAhf3sMxQVow0vXan2E07yC0la7vDcIClHWb9a
jAWepx0ou5zR9jEnqtuJa0yTq/8GDpAEaK06P+lBM5E/VUIptvcZEepJYFhDH4Pl6ZUte90elJzc
SI4T5rRQsKBfYVR9jtdzkPlc04pOqBYEnT+KqEwWAgPHBQ9uAce+/+mjnAhB85SVr3k5w+Sm3KGv
lBQfJEya6q3nO2AsuXMQoLoG/QXA1GsTjmg2XvC9u8SwreMyFh9doY9Wrt+mibf3ntG00s2zNa7P
0W1cemgUpgPz6DIQ8ekFHtcojIsG0W6EWiIvS7tC0aWgPsJmT22HFmlWfuCfXrVk2t2oVQG2JDWp
bkaueZtKC+pmvRcSfl4618b+iCcR4V2a1Mm7HwlJKbsJNtjImsEm+W46JiTCzikYGb+EvxISltz4
Tq1H99MIdN/j/k36fKoQX1m5jayQz5RQAQmkgGKCIoNw5Cs4Q2gDl+36PnCypowC8dzyLoUPrNA2
sEC95P1oXynZ/4Dsd2tao/vmWPjJu47o/u+T7ZIFOf0iKQ1IWJmYmrvyEEd5eSzSIiioEdEsDrna
18qY5OW75Y5Z6XdqLTKzmHf4o32pvsxKHpE5xHjAwdw1+LM16T9Y8LZVQ1CLXP1XDcCHbD1+1T/n
boyIao+CsdfuuOO7B9ATjdhPwBP5rWmq6P0I/JdSVtMiGHyvGottWk9pXWdSvuFSPLXyR0jkfH1G
ihJ7L3yUplCgqbXGbHluIS41SVaNU0ievv5kpnKA4UBCJ2w4qzGJ9MIAgQfLijYdKUB7Vp/eGn1Z
OMGDgypnakBripTFnKNY6StpXhwLNkumu/FuoG4+XzgINvjXy7Ic7R3g7VCn1Iw2xLaqm2V7E6xL
mcUN32zArNRkcYB/8BSw22oej/oD4gEXEax+0MtYXsj+bYxeRxJAK4F5Tm/XoTRkITYjy+RtwaV7
FDklLIk4LQco+8kikE1fLV9zuuMIB79nrInj55jLZV1jM9fcZwqSsduWNcoVvmz1RDYH8XH79Zea
Ul+HHGCsIdXGIfm0ti3mGGVnNpR9+n/I08SYZkhY5pWNitvE123NVlkRLyFD6ZNO9Q0T0/fdQg/K
WV7UyT4RQ2RGsEUkC4WK0I3psGP+WeGAkZDp8UsrjxnIpSkBLsy2hM6TD1hACQF1bvaAscMf87Po
muzSWrP1GlRZ+oBe5z1ar42Px9/UHcMEjqBaLilRQOjFWc10sHej4RuUM5Nytn0rdjn5bjXE8hp8
uz17fmDdbRLmPxCdOI/xA8DYEMVRojuRhvomLXgrbuFqlLcC4xuH2g7jUfEmCgXg+8Vs0845yY7I
xEqIkOJZFBZ//0WYhcvFoa0FizSU06R5leYrS64hPmkqqsANGC5S6jYurp8ekLzqKyJuZ9iNXKBu
VK6bsa0hZ+LmigCefOztA6wRhk0CS700BTfK45zLOm/7MXWSURA5x0n7lt7m+Pefh8pkzoKne1xa
8hUVe8mNNZmSjJq38ZsNKqGYl4OsvkJul+k6qvasD0/8I8lcyPsP/DwZsbltKM/AmwQYCM+qwIOW
LTyrywTOGMXRqK5Bl/piuNBt/APs3PFU9Kz1pwq+F2o2mJwKw5q+cQbcQSgAwTKp8gzspqHA3PJo
utJo452p4VR9S04fEVMKhJ2BsC5/XmoEr8hFZcRawPW6KUan9eaOfHwOpjzUGAHUvsbw0UpzuEji
x3laMPeXQ7gK8NA/uxEgZ0ayNWMKEoTIXxmAeY6XkJ5yMEJxplrVpru8kg63Jj4TnYnbSn2qWqP9
UeHCdGgfwV3aZW8FkobAmm/pgXVBCMCTqZ0cH4+dowpceDgVw5FOQFDJrKmpFEWOpRB95Pslo+BA
qGDtG+/onPqGXQ4gwa9bnMluXRP0Vg9JlrvxygQP+dDUIkqNRmRadKBF3AzknWe+jyHOCdcy80UC
hltSWJ3uD+ozRolzdevi6B9MfnlYnktJ7S25mEm4cRS2OM0tghKHwUn5nhFVmbExgkPYtNNh4QOs
vxUid6u2tZHG6z7rs4GY5QnqmwEC5v+pk4bBvlPTO71WlJax2n8hOtG+ITOmzHevHJuHWr+8TOYv
bg07zzkWJixfewSPmuKLqdXYWD73i/YX8F4QT46+KKWZI1Xr8ye91yt8DbXMmSv1kDIJqsIv9DkV
a2o9hyGx97c9uDVpkUf1JiWX+UdzsQxA3/rZlvAFPAveFNM8xYI408mOLaOCop4Yugdq2mXVlY21
gDbUF2ACAhOhUO53YNIM5TR7RV+Sdf0BPZ4ZTLX3CC1RVPMbBhvSrAH8IxI0FKrQr3PNvvTo6rGx
bzdt99UEVInD7lc4F97qEudKzMzDD1OUAtV/RA4I0Ge5DOIrrKoLsXiIxIbLSIIoSnOZTuWNDPJ9
IFBHMPQ/Kdl2TlRo50FTlZHGuDtq6FOnRuRAmCZ06m9BCVjtF1W14DFRP87kRfOHCUPRdpRtKf+n
PA/vv8AESvxyArqqJNVvutHQ3tcRdgnJH/84gsPrNTeb503bnEGqS5j6+yRBPrDOACPVufQFUs4B
YCTo4RagLlOUh60raf8V+5FoxRTYdONpD5JcZvIT8Y+leB29mVoCJMd8c9qbynFkfbJKPcMB0xbb
f4kyJ42CvUmKdvBdqyZTW3h1jiA/UdyvuHgx5O4e/OYCNlNL5BR196kp8lMR+CEfpqCFWpPfg6cV
dckvYHZQ2uvAwALRVmkpqBOSMZuqyMyZtclaz2q+bStm/E1lpdtZnmfbLOp2oRkxJYQjDbTESVE6
9k+vWz/emVelNTyu/o6FFnBYtUn5tP7OHE0FUkagSTw5gZLvn+JnDVV4Bx+oOrV7RjaRbRfqRraS
WY09W2MLNlMSpj4oQn5atSkUkasrfHynjsNuG+eoHZx2okTbBA7MKaNX1wkgAfnoBQHFN9ctD1yh
KYEoCM9WAdBO/uVOrrtGq/r8f/IaRqtzA68CPplG09/ykx/ys+PDIgWdjNd03LjqY0GcgVDlq2Ct
ZkXbaUWvJbXwExVKouKTthi3NrKxSauqqeIDNy5deUAa9Q6DDAiB8MpQRBqna4ldOY8hdbLjeXw0
d9ko9V9adoKD3gf0TpwGMpAYtr7DflxMVcyp7AvC4C0P10ZvV630RcZWPl/vaLu1HEsEOivRyud4
6NxhMVTw7vFthjdfcXMYSZZwfAcrDv91AULk0kXWH9CsVyk//PL9vo5awRG9NYOwQ2i6oX6i2aMn
DDMx8JDhEuPdsn3Mlf8voBGhLWpRhhSE6auh4N12jRTNfurkihEgTYuWw1B6TzNRx+dLxKaPDzJB
n6Kx6+eNOlYq/NEx2FayEFfv0H7zpquDQwW03VvTcjZTBhWHPClZDgusV6TD+qze3T6jnETkCfIH
QeoAwJ4Gfrt7goD7jVYYhTqzL1ocrR2gGBodod0OJA9ucKn2CjHd8lWvfbmrwm99e4Tq8+XH3Ahs
ofgDPA/35pfgH7OSYbBaieI530O8IPYptKHndWi8jA+1/Wm6S4vkcghl0c+UdRg1fek+DCGmRId1
7LZCP5aKGfJBBls1GyZNEe6U9jf/xRhIDQ/D/KaYXMJLfI1W5BtuVEK3Q9BjxcrdXHTi0ZKI6GW1
quT3pNDLShZBOXf5pWNC4Xl/i06GLiwvW0ydFkDt2tjmRJmpUzrtKTYXE8+FA5cMGY7PFP8hfTAE
WDMiPX5Vf2Sd9D6EX8KJO9072NITk252rQA0UNVOZLJpOZ+gmC2/eQWWbujVPLb4FjRCeA0Syvm/
w/G/KRYexVonfOpA653sHmWTgm6RHZ5YuZLN6VAUZi9MttF0l6aBZ/+5ZNP/IsydsfGiHDVnIEem
ZtNOl0kj7VSxCIa7bb6wwYCzQ3/8YWnshHfgu78G79Sr8bSSxZ7b0FsMlwDY1hmdKuIdQ20zPDhp
PO3ubAyMdgJ6cqfRR1dhWYUVGaMOhs8L+PrA6RJoxCKujw2BtV3QMpICPyaKAQtCVI9I7vr8/4Vg
6keJ6lF6C4V/NjEOnECbfdUOwFdHaY5gQyaaog7iM+gq5AImMosW3lZcluvKRY9apr0w2ZZqt6sG
rYIQsmsCZ4lAb8CIqTElGwNMLY7NjC0iqvpvUdvpSiNr9XnkIGrUhaLAlick62ziatw/pgk5sluP
/GM9snEW/QCiray7vFMYE+oMIDEszSKQlig8OuW4R6D3T8KqrC8UUhQ1KookGwhc7z0YKY0Su8ms
c61hxLoTc1HlNwIT4CgM978HPYT2kH1acraeqCJUwLjcGV5lb5F5Dt8NB06Nqm38VTzcgOf7pLUZ
emcSZy+SiNgnJkJbra84aWudotjO0Qd3N8mxhsq1ft/9I8kZCXaxTZuNcVoAd5qM/463i/hmk+5h
AOqasRTRL/HVkcm/BtjfQBlIyyio1G+cOt0cVjlcV3lI22X/yKiNfCM+B4RUwVIG9H0ZOtNNHDFs
4HwRP+Z9wPisH3Cfu3npSYb0eTx217esKfcJOXdFnxWepQwKQfclOZKUtJqbJBrx7MMxc6tubftW
ii8ugy4TEWv+NvR91ClZrIXbr9GZgE/lgW/xjzY59wehvyxWxlOmOorSxZPTmpbbQfwIffSoHzlK
wRabxTNU5YqDMLWM2F99MlwqXvQxPyIc9mWPYwWkIC/7fq1tzm4KV4AgyCqvlATV9hjPl2j/y58u
B74qytXVNWx2J3NHAmZ0Nh54VYVPCzvE6QVNZG+ZoWXnki5dylnwUv5m5+YrksxhZmqDLJcI/YaE
E646HzdXGfDNfJ2zNrGlWK3bMLRn1a5vrJheEIHtO0JkDP3LvjOy1SF+ZlovvKZKwKafBYD1ergS
hRSyPqiN1/FNLbfiMMRQJbgnulIQZ4616+WfuJtwYdoNOV0HLDeN/xW2JG5HnH/2OAwIzEvKC4Oh
VfaF+r5JTx/xBhZw1UN32AO0l/39UV0AORrCY4xHq6/Lkep6C+xP5OWdM8kvYwp7Um1saFl7BdYG
j4SBenYAHmgzDC0/0BAUCFmqffALjyfy87I5mptvMbufZ6+hIlYjyiw06OvQgGaupyCBPJWbNpIi
078aZAVRIw9dc/RyTkabKH7FmmzTGhY2XIsO6UlwlrpymvjMVfPC28nvsOeOUa2B6TDxXvU8fQxk
5gOYRLOxL7KIVQ/wSCEmn6Qx9ZibBfnUfmoCNYuax4LJ2BjJzHeAUQqjiyczTj6/7tVKg61RSRKn
3B0xYuup9bPcd2aqf2qPsOpox5LaMkeYhfyWKMJ0C277UrSxspaAFcNA1FC1mMes6cCKmFLi/gST
07A4vVNZ43cg9uOMzeWCD0Bju8a8rEWrmtDichH06vaiRxjhhwTR8AabSjBw5JWrDwOuI9HbMDWy
7/pUtQsCYy1QP8HBJfZQ7ZGYwy7v7nrdxgDttZDHTmDyd/tvqqOOt0XyRK/2VcB1ivl8H6WVYbrP
YnGSwagvs/4iskyR35yTpi+lbGIBjUn2ohFyn1fbhhPei1qYWvsDHoiFT8gvnjvZHBYbUafdJVje
KO5yKI5pWTVb6yeYpV4MsbRDkfqJXeCbsDUTavbeswLxObzSLZsreS37Vz35MFuOWfFoQZu1LwjO
FJ5fUKxp7Wa3IUBfxUmLHXo6U40YE4NI88rNYHgKvGyjIzVd2MM8xkjHvRoc6D08CJEiEUfM55k1
fa0IJXFvHcyoDSBrzxClp76yJKki7DpqyZFoHBDcM2hSiLPQCTpui++wXSd0NGDgh408M9PIqIYq
Sj5x0CFO31aNyjtpRB93wTiq6cHIV7UGWbBpSiNXRdGkff9Ps0YHgDwA9G/g8bPBxG0xo4lNbjy/
ObNjj+j58gRMBQrRYaibiNL0x4osjYKeF7VK5vMu+mqxBKuCz+9zynLc5mG9Lh7R7rTpq7CGQm/O
Wxv29G/i4XSL5BWSw6gwildVFDMoOtWNjdbBK5nxstJjEyvzPXf+9SUajwDJKrJ+4lEDIo5ANmoT
4JXUFxJB+tVrMVOsVmflOxgFc1WG5/xCOf6/EMbwM7h8lz1iUEP6XReEAnmUb1zEbwcsDZO7bgCM
JQKjCrYwJNOxWTcXwx/QkoqlBmJNpz09RVorf8FoU7UtN6J+GxxHo6hNKH8wn3SAERYoyAk0KWyW
G7Ri0YqdJ2Oo0Lc5ZK0o+wxHKGddAgFBmE4ukSMCcGshn2W/wUuQK1B6ODdI9OiHjczJfa2PwIAe
t/h3HKUPk2uRi2cqIHiX+xO1EqfLfa7iQww/fLclR9paoBHoxY8BxdS3A928niYgiflhDK+ySiki
XTSrIydRB26XsTJurHATcV0GBeuu16oqiL8CCPavrOEZgj3XnU/sQmNZiaWC/C2QkDtNkAAHg4dO
yhm4+haYSlCSuH4PNTqiosKvpVLqvcc7d3oRsSA/y1D+XUnKws82roU23hQBqi07J6hFfficXt5z
7n75k+tLj43CIMcjwME9mBdw1dzEIqquoqYUMSDdelwlv7i3s04ZhcBWtqqZRHBndRJJbuscL+zk
XUUyju/SJQMSCzJ0r94kIDCrYLynV2S70KOA1Pp8/fG20CM5XBlk8oLMbTeyncizhwewIsYdctMJ
y1W6s1rGkJdv4hwsw6wdGzajtiibw2PfVGSSKvzgbE/Hr1Afb/4+1mCWP+U29+UwIkUSakiJ+Pkx
vN43OU77NnHwiZWLKwPCyyoSwMJ0fm5t1xQ8/wURAn0lGB2rXJ+5igv13yyTNUM7bg/W5G420Jey
ZWp4VwNdwkwSMWIDbZOHn1waURjdfLCR+//0EFuz/gRUg1GIXjHS/f9HlYWonhzcVT0JnzFvMqCM
N9pm1NgXf2F1eFz8wJilPnYinNg1HU+Kyn7D4PUfda6uG6uiZouJkELHNWzT+dLGLU7jlCQj3sao
rcsTfEmTcORZHQsq2nl1kiSWUVG0dYwsjRIbl+Baxm1jCFV16FcQcdZyvWj90iuOIKDWqqFUfgr1
MuYnMoyuKbQnsQbeUs7oQ3NOEtTf+bmhsdEhsWSLVmenvat6Za1kszhaNbFrv7o3bR1N3XI0I4q8
Yv3iEFU6fKvcHyJy0tp8Qw64uk6hIM3yIRoB2MjANZwWHK5grJzVMSx8bRyMwcNQoqzV4/Wj3lrl
u8Ya5ZKOv8GP30fPFBrODizl1eqvkAu+CaykdQKaStM48AGh4UACYSYOJ9Plw2FfXAwsuFVGH89v
ekDpwhArgCS46JEJ9AC0qdTtmGC8v0Ftqfb0betO/OTgKNFfvaWUa1aNmwyjQCHnd+FHV0Mvo6TC
S3g6vgMsjeh8P+c9PXj4NMEr0Wc06SwdDTaOKzCspqWTFP3iP3MNjW+PTdjBeZygmmi+JNy4YBQM
nJAdaw9HrpJwTovGJB0UO3b764nzrkxrD/21h7m0CS4Z7QSZgacNzXroCapXkh3Gj3BZPUzNkFwe
nHgAyjEnSBwuc7UZfL/BAr14YYhPZNv7JFAp4fXCLD8m4gU/bDiFUbZhozRAGT8noJ45wr2s3pCn
0AlRb8RJLijZh/+/hvH5P0aziYSkEIpevrJfCr+Fkr58OgYtJsNq/Sdx+aD+hsKK+pOxQhIc+1Z2
emvZk/3CIXxHZN/p/xfuxQTugGtZpc18cfyXxE+BshTG0qFcD3CP66rjnWTwu1OUyx7F2bf60N8D
5OhKoGPUxvuFdm925/6i8XIMxdAE+wjldjZxTf8Kv7SAB4C9cFrZsKXHFDut9TN6UA3duY048j+G
QMnitmXY2W9o7BxKNj+dg2RC9roNZwqw+dWckXlcniOTceie1jGBeEpfaOo/edrUyz+sULq10bT3
xmt5jsACDWx853DnlyWlJEMMR9s27efz/glosKxPBtaxl2Ag776rIv0lQ8Z76o7ighu3KhxKIZQl
yyKinL4owIBqehfFxWHpMJgwP6QTGfkH8NWEmlRXfvu8rTfWW33wJXYAD/NOH7P/PTWzDCFcCWWp
+E2fvni7bzqAXMtJki59WOOjR6Vy1lA7gGBeZmInWfkc1dalEU9lKKpZP1h5WFVInnQahujykAA2
1AHg/+1J7GcKt8xJ6B10RdHbCElxAU2OQvvKLvFrrWBhf4af2IYnf7b5HtfY97ME/kiwCrZbIv6r
JAalcGq8LdkRZk1vuZ/314uo7pciCveo71JDNBNcPQemaysyZkWiIhYySGKtRKF/J3oQ3jv6b287
ZKa53t8EB+yYRPkaWMs+qh0bMb6IItT05rHzjA8N5FYoRath3DTVjOG4CKnnTBGv0bQjQL10kOM+
rMYjmq1HEYeGU6wvQgvR152zVXjUxISfEIjK7f6NCwCQBlHu3vZy04dhNRF2s/m5luLmJHASqcre
DNpA4TIvArx52tHRoDFAZctnTZOXyOQ3fMBMdyrl3GUNboAOU5ozjq4cil1LJdY+pPX7eD7E89E7
kuFkeDbsHT23/KCDq0W1A38MTRD7cNrhE4FC74GtWYOaUyRNxIcuyAdOPENioXKjO0vhl6sWElfH
zUtjRIZJeRVJIk/WLTWR4MY4rXu/FpVykaDsGkQjPx8v8vCFb4g/QWZIg1x5SnvK4l6Xd0pfF08A
zmacC3vQfXXBkos37Co6+NRKbRl8aqyre14W2q4mtG58FihF6yijBxHrRcn0I6O+Lw7jkPWhlGO7
mYFRpms8E4qJCV+/BRXizuvYtxx31Ypbq9qwG9D4Yfz9hm+w+RRyesi3zGAS3sXUyyMyWDpyUQ5h
JcmfJ9zAMWj2Am4fScCKOhLmYPQbBe45VoFFTp4tMM+d+Hpj3llkJC/3LwHjf+K69TyM0myQfsTG
nMWsT6BxRM4qynK0X74kcsRK0TxerfiQzcmsMeL7Rp3NQHcpOEO8Y4TiEQJqb1Sdz4G0EBx58w7C
HjITlG0c04qotTpthQp+1PiF7GjjtajRf4dQDYO1Th7KvvhtVPKF1s5vwP+jD4ArqcLlUnZIQZBE
6A8jMaAbpJiqkeSKPXAj3XBdj0ZOImczRvE+NxmQaIGqz2pCenzX0rOGsCBxwIMGuaETUcC8Tw67
T/lE73siDdeXibmJZ07V4ls7xb+Xssb5hyOy/U1/8Wb7h26G+OdabkU4PQXKLRoxtkjm8XWZ+/rm
KFOaJNS+VyEZCoZNsz7SSbJTcIJTXPMTGuKr1tOLT5aKjecDwhQgrdUm4jkDcQXoDtfzRjbwxsUz
1F6kgrJIwue9iNtsckVUcoNa0s1Ug1o4z1n0bmhy23KD7n1WNZOVvfzzEMSxbRnipx7oGNj9IE1P
NqfUrnFXuv3R3mLjfHYleQYgRoQ6Wjp4VIxXaUiryxjZsgRaoelhUXFA1EdA8h/jUfhqxNefyTzX
55tVJjxjVELvidGvNDYOKZApSObbcidGHE1G8ZdpF4k4Zif21KWlTk4+ZPdu3uBA3pVKTdyIG/dl
yYBensoHgQTYaWNO8hB/ldgi/B3pZgpVKQK/MlfUBF06PNCuDpbB5+ZQ0QEVP1ea9h0OnCrrG74C
v5tQQXt6CuYCqk9JW9tWTKIgvoqeRsctnBHAA01qdgsRvYMhHVsJ+rOfUqxaRaY1SJmrwwRUWe00
h6Iqv3wG1bhhNm1FDxgcs/DwA3gn7mJrXNQP1dbGqtIcE+4ixz5WQVAJyca+6KZ+rl5mZwRf49nv
dwmRHiMVFXRFgp+LyN70Yyd1jqJLTeyRMyqDJvhk3XKsJhfYaPOZgiN1kUbiFcX1k98gcOzTWD8W
8H3Qh9/RKp3ms3S9TpPJCntE61yzMdzhSzi67VY5w5tYO9OZP26hX7osQ8BhPKn/ZcrIFQNMM2e9
hoxN4ixF7xOUAXJTKQyYX1CHMyUCgS8QtvQSivCFwRuyUaLveYxeJESq8mxVm768eyMNj4gAJYV+
E31RTlWn7/Zfw3D6DH10P5W/pRc/nMbP5CgwQIPyAIv6KLPFdS/WPCSU3dbYoKfegAhRvi73moSE
GE+1tJx9Cocc1Rrgx5c6G+gBKDBFgiW+1gRXeOMmG3xucTPurNBi2KNEuNyB5YJl0i/UcQyXtHAL
aWzqnT5LLbjiJCG0UmpftAfYkPKunYTVwe/V5/r6a80LQM6co6F+OJ75qh8WB6K81jup0YKznPnn
5wIbQ1y63DtxPdDZ+J/ScM+vyUxSrWVUlsODCCAV1hGzb99ykVVpV2QL5PpBlLuuabwWndFsMl7r
ToPut19bXeBYSGFARpJZeV86syWir28x4djiA/YDceO5mEEm1TUu+rslYDjnvnGnbNSQxKw8uYTz
FktVoGW8JAJqhDD9OXgggMkv8vXHvoBdqDFPPE/9J1nGlSPcHwquJf56cktiI13tQOeIqA/6ioXA
INxea7119AYVYOFyWy5TvIxjljSRPU3pajCmSZE5Qb6c/iS+QRC5JSFeMQ9o25AEFf73WqeqnX6t
ji9cl2z+Mf369N/Y4vY4lrO8nBDg4uq0QdOspGvuoT8EvzQTMKGdRdipIqgWCZT0k7aRtA+ZFGRx
WNcfGjpYKROTzYldE8GAJLGFgDRPcfoyppGu8gDBaB/Nyzx2XrsWZ+dAJaP5PnbiCovX0gfPJamT
hkdVOiBZ1GpVn1WKXx9jMSEWkeTqEGAkGyx/aG6ThIrDHhOAgzUVIT4aY+jjm8k/ZMiP97qRm1Zr
ZicyBFo27X79KQ560Rvz33Yl/WcLBCGFYUKonqraomukhOoIfgfJR0tsz6qSKhZ4FSTGzbDvxOn2
K548Onae6/RWWlfBggBRV/2JKJPuR8LiUfkjCcEfCcePfbp29hkdy+Bi737JOoxPYqqVBofwS/uG
SIJu6PTo2MPCaZsYaHyBoXDAofGU4iaDlwnHiOe0LR9b8K8wmIgTnDzGFIyKI9owzkFBEIQ+gN7i
H0bq5Au1BjewNbOexxjLfsZaSSSoooxEqcAmaExV2ZamEKK+rt/+KFnvLFwiCtxjIyPsX6KWRtu5
mCyLi3impCtm4EKoY3CQEXlq8ZMRx3MctRuB93DsRmmJBxOgYGB4WsuJeX3XuA6VuS8sIWPQTHAk
JxILyQQyHIAvzxTjcdh01aTqJ2cBN/JALjPdSJ+bq+MB8ajvAnBtuTk3ly1BX4trji55TVdUjsMc
/xFUH7qQW8GZ0ZAUdKeDsvnBjgDoAc5TMQ2s25prtUq9Pr086PF2C+OjmiECuLZ/t7pni7xuNaMP
oBai/0cGPwh2uMPI92OmBcjzwF5rykt3srt+yo8VfhCd46exmCB4g1lE7R4jh+Iz8RoRV2tUsVyw
roGtNT/pHAYxWW5zlQvJxT1adbQoTjSO5I5UUV63lRC3cSv+RRkFlP7zwfFXwryut1onPq9r+aeA
JdjYN3VPf5LJ6qdV3AEr4tVULOPm5Hl2zy4JL1vSo8rG/8NoFUjefXTye3X/8OOXTZ48diCLjj1A
5r3Z3vcWXuwx7sF+h1PC9VrY8iUS7zKgpddyJOx3Y89D5BO8JQPbgoZrvsLEACB8zTRgmvUtRule
cuvMiflOoE0Rfc7aNKOxJQ8AZaZ5N+EqHL/wP/9oGomFsKCocpbiO0YpSxU767PImQDC7y82n0O8
Y86o0LkfEkkuePjODW7YniybfWWZejPa8R5FEaPEe2XmP+aQsmeA91XbLrheFhKnoPY4xeyMWmPE
Ut7Zn5YBv8ukfRlyTsw8ULmZq/8y8GoVXTaI1b/RG5wUYdjR+igHm5tgPUOkITAjAxRzFTpjL+DB
SEukEjnSyLThKHpaaLVV8utFbjKmX5kkInXvmm4r/Q0N+83U8biD6jIPnM38nFdRhSiZUmn59Ypl
HEXCG5C7xgeUyetHrn9DgWNW9zKzZdYG6booeIw9sneTZAfhsbDcOsR41Urb4Mu4uRoM8CN/LjDz
ce1LS2HsXDwCKwvP4tQlPBYNuU5j+pLyap7sQ/v8Y1fqojG8+jaak+3J7hVenBP5ejKVyYqUZCMa
WXtr1nMBU4kVCywrnHKJrfB5lstumDKF88q6hY+sWCOyx2MeZ+Kp1+mTqOLLGYbOxZYuNpqiyuDu
Vymhd/kY/K3NnVbr89yd6pkcosgV7zHmVkplZ430CHJUl1VbHior0KHt1q0WK1rATdDPz7Kszd8y
Q1+PcCqnXDRGzkTfay4QGvcnXqd+Jf4BLzf/fmlnsq0eXs26flA5zyG+GIz0pWLbWr3NCWLX9BtE
ArL2p8PWks1kiyKxWo5AqseiAAbB6+ZSoBkfbXc7bgBAt77jSrB45lbITwW3XsAPhpO4kia0EeAQ
UsUHp/E3JNBTJIcJ0QSIDZOa07fkFMtQz88x9vM7cUmacE1DqFTRoJ/nfsVn8E6xTZonhEzcql4b
WA8yAN7fHILeD1/sUbIFXe+QA6pF8TAcArjrCyNnszk2EnnqPh/zo/+rTrdZj3bCkozAEnsHVv8I
9Bjf2GruYFTNnAmrlwPZ1b8iRps/W+Kdvn6V0rH0U4RfGLmIn8GNF4cPnxhShLb0gma6QcyIwQWr
hzdnLpgxGFX9Dcl3LXshw1Lmc77tIcn66HoNTm1gB6xUwOLtnW7m0bSrWsQakw4oJGNt2bA31Cdf
093Hmci2BOCj2W5eRvGLh9o6xczSm0KddEe8DyGerwboT41iz0PhDmoS7LUaRfL+A48t5rAi2B7+
6eztFKg1P0Vj+74Yf6zPfVPuhLzn+kPrxM/9fZi9Z6CbwsNgcsyLIVhpgyaGTKq5Y0Lv/Aaoy785
e9k4oa13OTtNoIhnFmzBHFnyPqgglCNbSXhB4gN/m6LkMMbP5ed19nEE3xu0X3vmHWpI/6FItnor
8flUz1CYtDRjrViWI/Vdz50yEKffj9m5WuRyDB9svwXITTsUDblbNo59QfGQYxlD0JYOF3TAHcth
XvHxSqP8dbd+5m5EWqRUmWri1G4nqFTo5KzgPrG7CVS1yw+BS02FJ8cma5VHsunTg6+gROnP9AcW
XsbCiRwA3CUkdMSXa9d1bynF0B/v+dYc6OguFn9J4o2EnvcJEdzmUXqSkXQdh/wJXID91dmj9FKv
NqPUo8xiL0AcE8Z4PTYUhqI05KgjsKC9+BLh8wkhYfhXDDmVYw4tv6rTGJS2jLUcPhLRmpn7bh8B
CS23n2a6Os09/Vtf6NGIqwQXzwanZoHmyFAveF6Dg0aVkmBaYIbwP88h1OYq4EqaTCOlENjQ25E1
ioUNzmgYG1YIJrkKZysKu4k1kdfIz2pjU4ZTM/t+rJX8CBtV4pIgpvdt+0r57JygSFWjuQW5W6K/
6a+CkVZpRPmKkokKcJpHMJPyd9RWFJShEVWkUfp+mIGYCHBHUbfsSfqau5l+EIIr+/3+TnjQQr7s
bGPnoiolBQ+VDih+ToQNSJB77onMdOGI+alcQvZOBatCuIlFeHZVRBcCrAh/FYZXU1RtJ+ubQb2q
fNX7XiyQeWrnZQMrPDYTzoqpjiYADni+Yin9duiXs6GTJBmg84YVPNVoaVvbCbPs33xqVIGOPSnP
u8fJUrGX520uzrPF5innIbyMxsc7XT8JpOGJS9LFMBrVgsXxCtdH9We6/VbA9ER7yFP7dT2ZiATz
geajtyS2pxHfJdCAiT93GN3Mu0p1MQIdrvSoMDBc8/t9ID1WzCWMv68xrn/ofEtlloNhLggs9nGk
MfU7BB7VQ7OEr3WHl1qVQGFpCQeCIpl/APZcZWUx8etEs/Wo/GXe5bp644GaxwXpC6VqDCyiZ0v6
qNkXuoqBdLwrGSkeVzBhA6EeyM/X/ssV58JbeX0D38WqX6x7Yxc5YZyJBTFu69emYm4s+e7Avgi1
+sxkrDi743FeK9w1MYIH0VIN66lORvCfO4tTDNQdMWeIF/3LYe10UZTT8JjMNGqIeJ0Q5yj9UcLz
B7uxFh7jmlYUJgmAISX6XOyaVgodlpIWBGYmXGxhs0erkgT8pYQYXr8MUdMXAkf5pkvWiEx6h4CP
cLiQri8o/bss3t/J4ld60i9wC+KOu68uw5BLZ2B+XO55m9BXIlnSOUm4gSqlGjrlSUEfmLI9KChH
2ZuaPJyeXbuCrTwR33WbOF9LvabxQTSJXuDtkVJauQbr7U3ZShBTgLSgT03HihwlTi0ouVcjaJwQ
C78W6xWx5T3z+s62nxWUB8Evr8IMqN+DRzGxR6TqH9RcTgCVeaEx4NJehtbCFAMPCKFO80DaBJre
/bCMXNdCqRXVbY5BkyLxwQI+bMtaBMK43LeUh2Ss3UnP4H7bPn28QDFeJC9x8WCCuNP7VyK20yhs
dQdpWtr6L8j9m9f+idINcaIuolywxj+lhJx5aelFwgJp5a7tQ7qA66ENnngOVF451kpRPHncagFb
x38BNbxEulbKrN8SCDC4A3SmV4/fQcltyOmcA3qR41HUwHITGx120rP4fyMTBs92TxI26yMsCKun
C3XGRheHoZc4tS1Z5KZi57mgs/ZwVN0j65AoadRjHQ927PYp0/7rclHEonS81pFWSHJEEtohvMSz
3fPL2wcI9XNeliOEh0Uhpab8MTu0pQc55wX6sq5Ga48VzrN9H/rSlChmBP9l8Px6vSibV19Nu7fs
xTE6b2asQvPpwiqwIVkK+TKGTLUMp4ndDmz33qsE5nHdzAc9WJd819m0TxraJYAEjaCzJ/Kwtz76
JbCRULkqn3OS4RD/bIDo9onKsRT6qxbBRIHFE3J841s5GMNOdh0dBcfkAUhW5pPSzrFP9ZN5wGJ8
z4i8pEyHXmrgwA7q39RxYOSiKO+q6QTNLBZXEzxiFYXHF0CWcBP6KQtk1GuKwZ7rg2QJCpf9wknb
lKLu3OSjCea4dKPtpJfzGFXSPArhy5c7n7MEi6xNlA0b5Gk2T4fDc5MlJSuBDOWA357KGDFy6j7O
ehb6yS9CiZBjQJZWJIi4yDcu1UtTHrRfExxJfNwHXEkSPjkdj7Jd0pZfi0wB+XB9/GpNq9X5OtpK
pW4h7rZ0Qjv0wq4Hm5mKBs//aY3D8h9CU7RZENsmIU4pI2y0eUjfKQXNBaPXePrD/mkr8yUwR8Px
rReMJ9wKdRUNuOMZsmBjJBwFD/kMQujEZvTfR4Sc8wPjfnhKAMk/ffzB33+TNS6Yxhr0m1nYrVgf
jwO4L1AwRW98An4q7QJdJQw6l4IoVPD1ToGGE9QmRjX0tH8XKsNVXGyDScFQhXbvQUYByOp3luoQ
1W3wGSjY0bNutC84bDuMbWQfSdjUUQB2e19GrIalMOMfeF9NWDx1AYcBwQzO1u5mHWvuItZWqhCV
79DLC8px4Z2HXDdc7M4pc0YWx/7ujuaRNGg54Jc3xdZXXCw6iACBWgPmT+X8ScVnQZJRlnIs02TU
yijukQAx++98h9Uqy9B/ZL35PIr3Fvmo8wUnfvHcJawQJzzIt2kQUZJsvZVlz0M49UiCXe2TuL82
ClCNNGj/KDaLB9nYPW/B+Sil1vVv0N0MraokJPeTovUawGc2pZmgNylG5WPgFUxnMVWFmGEniwDT
wos5rMJUk2cIym2wXFK9LnvbLlvtqB893ub0+wE82BzHno0hVRuU4tlDaZpwo+uuH5dur5QHb1pZ
ZPTqHBohd0l9ebDM2ll/EppzWutqGOcc1Og9MCIZfRdzNGq1dVNEDPa+xAx1ep0vznkL2C2Ug7US
9aKeBqoRnyoeuUT/uNT3Um7Md2fl8GlaVL0h/QsFENzxKsMdtgXbK8m0JaO96qChhBOZ4Qa3pu3u
ltl9YxJJQ34OHX7k3cAdOiubdvlW9Lv3lW8gT9YabJY8Sznq5fh5KZgYKr2RaywPZxktsiGQoAVT
QTi+B1HUVzcnrfpHzbnEDBMXigsGCJnhzcEph2MMhh1mO7Sawm7hdQSLp0y67USWU6p0s1v795GQ
3OcIKvVVJd3oChkCuUuGQPoTnioKTPIFBpV5k/LpyeX45yIgu1u9hEgs/4iDUx7DiEwFzFggfINU
bqqw+c6YKba2RfDipi3Hi9QY2MHgKCwrIYOMgdnA4ybPPvS+DRkjzODLxGVavB9L4vBYSqAjaZDv
ppzAMrRsCpN2vACpVVeDwuQ/wM+816qDIweigEgpYkJ3U4+uFFM0dOOyzMiJPcraq09Kk8WYQ/Zr
SDUvX8BLcEsZYmyoCw/w3XG/5jb7pe/aS27PYzBa7FjQMX03prhws+CaIhZgBJlFpTn3mOsrJFLt
8yquKMGzzDxp/KugiFl+RtDKfRVQIFciG+moXKs24edoetltscsiTfCAqQ9qKYYl1lvoe0t2qSd7
FsmVDuU1qz6Ydrmj1Bj/W0RaVtQzpljHTixaxNZlxrvKzRIUvK7zVD0n+Eq8xzQDEKBK7vGVmeu0
FTUbfMjOw9b6aSa2gJiO3d3RuGpxcD9rCQ92PHNdlgc14U9wqZtpljaxa9P0WaZSSsSbDcyzMKTe
h8zKTD40fJz9adaIJFVYccelhLY2G0btV0oUmkW1lNK6cknPjEhWOyZqS5lWhlkvrsC/x3vKsCCo
X+H4LwdgDVhxNj6ZDgTdZdvE7h7dxphHdf6/cpNrKpChtdNHqH3+iAA8gI8Eg/g5Lprf9tMMbh4Q
kNqnsig9u4F+Mwq1n/YMGfLvLvHEUCDT+S1ZX/kM8fmiUBmuFO1jOT3N79ZQN5MRFnxMJX8vsvxy
nlQVS/H+OcmGBmmyTr/5XO117fE7oVcvQzMRx9uc/JMgfaP/Eu0z3rEb1hXAG6PDAgimNxQNlvdh
EzKaUmvp3dGOyb5lCGJl6+j4qWHLG1+zqwUVHrviHl0HI8YgjlRSzPE9wm45Z82ADp1t8WTTg3SS
FVBwPALxg+nQMJjzE7z0NzO+RXu71RXiMULtrM3VnfvHsRa2kkaf9XUq48nZvKwV0ND6oMcAy4W1
2JcBsgwuntAzGDvl9mVK0ztnBNEVPR9yf5MMxgkHlD6JCyd8jZgTN3UWiTnbXGmoX9IFr7X0KipJ
gRmHe9dSJ0LstaaT0LN9hzc2M6Fxzcqonc/ep/bMWELmgycGC1QgDYCBzK40zoN6oybuZN0booZS
wQAgMeutbOaFHmvzc4XOMgRUeqtiNtdZtTkihRRYhsC8xpiywxC0T9V1OBCEMhvH1VFPQ7hx/pIO
Kp7apz5YPWyTPzmrhCiYcMHx1LeTYEJp+RlXGa2fD0HXxLviP+cBYJx19SnIU/RSQKJoxmiPWccL
lNlRik5/Q0yyLD4ehcBmUDn713e7yTJM+N/N6hsNbGC4dsHnjfx7fGhfj/UOOS6itVAJKqJ3e2hP
rJTGmAvcQik/4kR02M1hcBxgRRlFYp/+mWRB3ewYM+tzgRSN+30ymsZvvcXgWzqhAqprukEkujR4
oECLcI39ZQXZQHWUrsqEP5H8dV7ptiO1UNOtSrkLawnDJ1i+XIXHZJ/mFnIBMh3JDPzAgzt90f2p
S5SM2rQ+zliePfd3gV7nDT3pXgmvfVrT8dz5JMWXnPXxu5AJFy7PtwJqqv+jflFd0smbSMSn6QUy
0ualycucHxfUAH1j2gQtXurFxIfDHBOth0uBbe/o86Gk62y3vC1n3pEq6g8R8/d7uwcUKd2u3FgP
Q49kg3NSkO5dMWEp9004Tv4wyuYwPmAzFCpNsFIv7L4TmAiBxJKbfh6U8YjgyOT909RDN36ZXlF+
da7/6szFBnvlKzbhNTB0bjVDQTcuRg5JmBTh0Q79A/PuTjKSIF7fbP6V5EPsyoh1EBfGf6EtH/ap
wTcu374K9CSuwmsE8Ha1nIo95ZOLn/CbOLbJdJ5vc7J6tjYlFlmaLzcvQBNPmJEmdfm6be+sQkvO
cMDhnq/h98YFhAPugfzliHP2lx5+otGrLDSZLl50IEW0zYsIMydngMbyI+4OHqfQjeUtEYnfNmYD
lNevXvEbjWERZLfmARbcx8QJydmVyDZiVI4fdkq2m5eZ+Czf6r2pG0EvRl4wjDt+5enZStrzY5eQ
EtN7pHr50RV8O5kuQGgDXamQ0+g0FWJpOw7o10JjwWjumIsP5A62m4A2iztwQ7efoW29EBsFBilE
JCuKwNFCRi3I2vYpYZgxQRPsC/ub5zvLTN8zNdYKJFB6w32oR5P6ECac0cr359GLGiQ4d101WJSM
kWTiKDL7rnjZsydsxIu20iCzwkYklCQRAfPFCXUPK5+xYdSKqv1PWFpyAih7ZSpPLF1wvcCBtY18
XdZmWnu0CgX2Pt5yqQQNo38GYtFyWvSiorWqilJ7YVXHCQlYnYvZRjBBTj3t6mViqGYCfRojr1CB
mrS9jcBWf2I5jqaG7GQrDQy66q7/yvgKeEcuAK2jNzhbnGZ6HKSX1fiYcsRQodEJmEwHRe2DCu2D
cO2xXzJXGTjyhNWaQYCETCaf3ySn8WkWZm/Ylwy8jfZOlLRrKB4E1/8mTVviQ38Nr1yOzM9GJfyd
R2fDKYZjcsMDPI2z+PszGuz4vzacRqXojLSu5jXQIGKQfUxWNo8ZNpOHoMpTqSrImE1gJiRoVw66
ztKCFQSmsvstVaEw7zVuJonjbfQVkzXcipK+Ue9W7UEiYRKR+6uk5vmZ8KC9ykplp2hzEKQ48jTW
wilYmn26NYE6ZXL/WMT+7Pi2hzSvXcHIJlFJhNKn09uCBSHIEHYaXrQln4OIrzshRxS43o1aXKZy
u3pAuNXyi5bBa/lP2FW/t484WQaIAazjnX3dS3TNt2nqMXFj51lAyOhMlO5nCkzj7Onxu8EhS6L2
Odz8xGme99t71WXTFbP9euL3BqiDuW+7vHZ3Ko49CZ5WTuijcVoNkh5c7y+UZuhyQIh/qvF+TOKo
0t5BVDamlMRZTOvQWRXBHCSEqvAOar6O0vDH9YQh+SiFmHH6oFMdgZ1tLJIBJTVXvR7I0vXhJPDS
7tvpfUtXgoWz669YaSYowSZakksqohX66b1vPXbHM+JHysbla8H3k3qGkmigTqUwOz9WL5phuErS
tK5M3DwDAUUM5i05j6jdj/GUMfsjG/bh5FBMswq1dhv0CMohtLI4XOvY4/Sa5YFg8rSqsKgEppgW
pCnkz2N4ajW5n7xny2IZCd4cr7+bKN4bQT2mqz88yownZMitJQGeq6BUIaAbaRn3CQ7DtzuSX1P/
JruT3tHO8/aSo3jTa4uKJ1tb4RGtqZTWpYvldawB3/35BXuoSbiFCC6SfMaZ6OuxaxR21mRUKqVS
li+4ALsRiQn5VmKFn8UVOkw1+Y/A/BCc4M3TtFeKq7iZF6nCHFb6lg6jrzNrg0At25fTo3SstGAZ
xjUciNEMIRCwvpU/Bop7467Zi3EJwdaAawg2sspct0XW0F9MbG3cmKKbIVBTiYMluQ5XrM7a0str
Vr1Wyt1GZoI5YZ29jviQLhbV5wDXuEyreHcmU+6hlcaLvopKdTAV5VdyTyzMaA9EQeylW9p6hDci
K9BkVTHYVlGizkM6/v5dS9ZbfK2muDTbAPptw43TMZhNNDZlZoZuqzcmhoLrwCpc6Anja1OyMKmv
ENJLi34qCe09mjTi8CvltS6SF+/TsYfX4Tp3n7Bssqwvou8tpzUGFO2dc46hHt3wT/0xCv6/LVEB
/eerFbjaSbfvsQQzo9RREno+QjQ9PDfzKMh7AqNoh2/yC4osCrW9kHAZ6HshjDeTVbZdiaajWsFy
iUDjMTrO/fVk9d60NU46f46HHemu9FGvL5l8uu/JOyMKMgQ4sraXFu9uO8ezsGQwKx4ZKW/AiTfr
DHzEvccntpZw1Vux8dkJZgwQVK3AIfezz9RunQQGONTcEAlqb8J+Th9N0zU4WFiMMKrmZ478q3GY
2jlSq2ZEIqlUC3Wss8pkxFNZ8aQGuBV3EBr8S07qnh0vU8lqHm7Hi3861IhXaDey438SZVTaTq1k
enY9LWhEsneHVcO6hsKb0O7nzMHkI3whFOutlFFVxtrF3KO1M5QcjXDrfxfsrHQs27j/eGeWcQWt
UJ4vnNnDakE8NJ348bI0dGXnZxlAIEXEChGq1B5dQ4XcFJKJEDkchYL0sUqDh6cwmKnA8r7GbEwH
vIhUKy9gmNUEWzYLr5SB0zTNXo3lBzDJrxsLeuRlE03wHTWJLQWSwOoevfP1V+7QRkLirGs0VcfV
TEjMAmLF5zSwoWgTh7v0GPQKKKp26K5E2ZmPR0ta5IEx9mgj13bqS6c+MsLXdUxvR2QNWo0L8tZ7
PmOCGnrDehNKxGmXZjY5ou6Pxc4/R7uvjHf0kwv2yxcOmG1pCzU5sQkHXWSoP1CdDfNwLLupc9DP
QC6Su19QTBvEZM36rZyyS9x6jfCRIxx07SqOyjCNT3cf4tDN03TbYREjo0YsRBnmWB3ldp0IIyYi
keg8Q+bnCDzuWlO5QB6GUeShwAZmVCi2xFAxtZvcF5jF6awiKBeKZiUX8F6dfGfFEtQvHU4XDGDL
HqOjpmtIMKNgIQr2CR38c2rXKb/ahBXM0KkkfN4wvzVql8jGAfRdqZDRcK66aKodyp6LJbkN4TJd
1qz+po56UI8Dw/5GU8R8G/90hfstxNeqn0jvvZelj8hV9uekmeTu1GvPTrxHTFJ10naQ7tiYdJal
HhG1FeJ9q6AD0t0fUW8iKkZuSLPKPQDlbXevERimfQ4mPEtT4Sg9FdZLaBKPyZtBHWyXvwlfmGBw
hWIvCtiy68YFYGHZAJgPbgT/BJfxTRJ1FYNNIBTzL5Pau44zwO4bj15g8eqCMCjqhG3/Qb5bwBOP
7eohI+GpcqCqP5gTkPo7/nsqGiK++2bP85LrUQ0mru42f+w8RjI/x38Lk1ovClbYGBXsxKtxgTq5
ClIw/Sb2ETDmNmqrmeQ5EiEpgfbds9KycJW5vjqvMxwwuT4IbaQdEMhDe4x0c658qLsvqWhn6NHF
ZA46/wzLiFxOvyZJtYT1asww+k7B8rD0xPClVi/MjE0AUmMlLhvUNM72fYgmTUnDu+IF5i2JC9aV
iXpyN7JRiDjLkoRqhPpa9SWCUvjoOeuKRvsAkozdEu5dcTZf6wy6PNwR3fxWyRst847sTPwsU45s
RDHElCo+0hBqUKsApkW693iWKIPm3vnQarVfzzvSsCLv8C1YJhI1R/A7DSTrqDudE6dvhliCjEVK
jOfuIFGXxi40PREAzUy2509Bke+9fsXBBC4PJHidYdHH9Ifggp+4oB02WR9g7sGAnw6SnU+BcR75
l4YnJ1IedZwofKvjExZqSsx3DWLCAVKOPHcompra3AMqpz1H6b1FSjfWT65FFO9suEFdDEu3HTel
uHS6J78Z7beGFx/1IF5MddjGU2vRIvByZabw8OCiEarBU47huZnIADo2o/ItfMhq1zDkoQoRZXEE
MvGTG+KjHCw6ylEZjsn8D2CK3kVsAYAnSdKLsV7DGMZkr2cF1iKNcUJLm/Pm1Qesje+cHbA1biZk
2c/UcYhZ+8kLv4vs4shJSHbrHgaxhPDdEonpM9clSzojVD4cgwUR6FW82fabbqnjSjpK25MmthuX
T0nTDNCMhDwO4L0/fGhJGv0w9g5kyrJ/nw29j0OhHHn8qNzoEyzmkG1WEKldOvS/uYC6nz6zoHxK
5cjH+Xe4or+bZYJCV5bqJSokjsQnktVgkDTCQxXCvio4OLPuy5k30OfbAKaggWl9rzHqoULL8FQW
DFMkH7RWKpnxFWOfUElsxASbFbYjSc9cQR0rZdAwm/XGokm/seDeSMgtNd8m7e1ZQ/Y5e4ri6Slg
l/u+4lXtbZKzWG8LIohcyM4cpB23mDyaxDJc3h0QW3lUJ0wZUUZtUlEWcnm+vtHhpX3BBvfhE09I
nSdwQoYX6q2RpENCk0vNGy7zT276r601de6GWDHcI3lMw51C7wxM5ZrRt/PhJ4p8MYbHBfuP95vJ
YUPmgWMvwNRFNMuP1byr3PSeMsPs57DKNX2Bd97lucgZnWD2wsdiEMeA/k9JVktpVLPuHwsWZjw8
xcGF7R9eVDt3t+IliFFtyz2PUApYXVpP277vlpZ2h2dcjJ1Cfy836xy7vaqnQIju4eX/G7JnpCWP
YxR3AWaND00o2J1taFQeXjbN/2w2TN2OmZYdJ/VoKiIMr7M3DNfll/zEKTRwVC3Zch/TvKYcxnJv
CX5G01vT197R8WH4oiQt5oQNqT1Ry9mCpNPN2SJXQ+QqbaI8EZkOQ5lC0IMN8Vutd0xUKqW+hVKC
sFgnxFvqv/vmVKpSr4nqvdHlEMXDqWFDRFEApt+6jeljuORPme0WKQtBuUUPCr+g8HP8adFRXcKV
qPoDyHQ/51EU1wz2j61DqHgYzmrlNB1TQRKXxhfJRmxHrta6yD6pgJPJSA3VfsXvJvyX3CEwYIEW
/15AN1RqWy4kDXaoQzcoqSpP8fF35sIDl7QIkOBa/0e3PJpnAxzmPLRDqFGvECD/CyelZvYNH501
xgjnRqsRXUwwMD423MMJuTC2T6F1mBro1XHTDuCbNIUKIQOEyE82HPMvX8wDZEf+JRkatIXCSXWJ
QTKt5WrHqBl2CD52zGXslsYYK53zttKFUQVsAJlqjzytAxIh0pIJxprKzLPjt8H9oimpsQSTqArK
0bH+K5j0SS4lMPwLpox56wZks0z+7V2H/1alAdQ1XqGJCXb9QVvRHFoaqQetcmoshC2F2lvfh3jc
LPQMsoSxL1zTaJ8lY3CM3fsMegKSEaKlMUNJnf0iY1q1+P++JqbPybq/YTer/e1im2EWn5Z78sQE
Qj/GO1VG6+nCCLLtUSKHLiefj9lbWccc3PxPF6yIV/RaMQPZbVYyy346UNesqrJSkq+vEsLz7Cb6
f9EumRpTrT0nxAldUGKsTFvpBR9KrmkVAwDSWysWFhu9KkO/aI3YffGZOQYBNKluH6Mp3QjLKZzL
9Oz2hyKshMmaBAD70vBZRO//jmt330uZyacvIGGVTkhD2Rk9Xv5TzldXqFiqKjGMt7Vc1iZzjjOc
fDp2+asus78KGVuAKiN+UHY1BUG6K6pdpHaso6vOxVNGD3WrWF44oFFx+0qhqZmputMkwFL7jmhf
0Mwp+bw3S8b8OR53eyE3HccBV58Xy67Zm55u0B0zbWwHg3fQWnel5B2bOKfiVdcY1kNaxG9mXOmO
F+d8Cus+7C+jZMlqp6vx5A67J6QNeszbOrJqS9s/BE4mloOsFmhlHXYwhSj5F1pg4+WPS5gWdiOV
TzmzugEaxgf0obWY5QA2uLUvWBDiNboz9+j6R48b1bZ06qN/uILa3PlzBnl0ETzEjQOS1RyPyFOA
Xyu/RXQJ3sqpXIvzkG/QJpX1bojIaWwjIZ7OGTCDyAPLtAHHgYXb4wDnKxkYqwVbna3Fk0yfeMvT
cZxZKU1ysh5TgVQIUyAEuEhbtQPqNsIUxHBCTD0ILz1RZ9DMMNCBBeg30PkyYID2GNX0JN5Ypfx/
bz2bDt2fGpDFiEobHQRo9uaaM+sE7vMQH/JGhow9JEhLdOd9Rf8537s1Y+ZMYKh48SDcIp7cCghr
AluBpa6wGjY49aBhPXKdc7Zqb7RavYjZ0HapdnPCbtDgluzrpk8d2KmcDiyZ1pFG73H1p2fKPbLp
l24fh5CqKcesq67fpjKIM9asGAmwfw/RxuAYCMSN9XbFQO+PgJE8j5hNmnfwvL+2g7s2xtkmNuL2
dHALy6o8M3uGXlNEQQJKGT4wiSFR8PgQ7YfkRSmqLGjSmKntv8bJGnZhohet39Ox0OiWowiEOri8
oIE0SY798lUA1x+Kj7IQGaygamE5LZOk6szySVwaE98vNam9PuRUjst1Cwhx3k0FPQdgMn7mCmlT
lNYrWtcySpelrMWzC0xhUK/RClzHPz9jEkhh/uuX8x1g2kKj+V2uobfPr/CEypKskSI+Cem/ursn
vNRDEZ3nbrQEa4EFEfHm8EdbyC0RAWBQMIBrs46ed6CS0B5qwnBE0eyt1oR3C6f/s1J0q0lsoGVV
s9Wak4qZ90A3a4gcsXP+SZ4Bp4KuPyy6fr+T9SkxkXPBGDLAdryKsbASevrBceEWjKlwFxcBxHL/
3PCyw9nZudHMBTPdlFXYiQGSYc4t6S8Fh+tyz+Qcf4Nq0nasYis062u0Nw2Xjd83KFuGPkNtzDwr
xykqydWm6i02T2IlPfgWCyfCiqOA9h7beEUIBkAChXL1CTeiKbx6a5gbxHdjR3yKGXSqsyqCZkNH
f2NU20yCdT5awwV2iFmVvCMs0ck67f9FHCtiOUHMGens/zq+g+2IOoD/qU9LIS73zXdZC5a6equq
X8TdgwGFacvvkjACr8O9cX3RUkyKVu8UowyjzwfvVcLQ89xWBdpJ3MGTqMx683k4J1QrNkM66wDB
kEJLemIXF1kEtr7gI8yvIhFS+EGQidFyg+i/IMifiodQqIzVNBxoh+IG9ICWyBYjcoJTQOCOb2ex
+6z/sqzjsr7i5YtT+GmfCkv5y5qeZErL/J3wecnWTv2gjfUgIl2zOZxa6SJPNioraRP9EGizFBbH
vcqgQcGG2RtT4qFQIeMeYq0K0M1ZMGx3MTjZWEe3ytQXfoqMkHIsOs5WxsxVvkbEdbX6PwT1Yp5m
BfI08Z8qHqrKdsM2OzO7ihfHTmkHGriEaclcdA1s1mbh3eXf2ung2dsDusCeU2hlxAwEk20Oz9HA
IuSjznKMn2xQ0e5CGsLEpV20lovKWqkx9trTloBJUVzx4usP0AEDT2FteeLelEBx5g2l2BwXvH4s
vLWn//CxGi76Tr0aKMv05qNafYcJ8GX5tH4fj06Vzjl6dutkGzfHaiAd763gxru0NyKBmbsHiylX
6zWeTAkPArOY6dHJ0Fl/aXkAm6O26jL1LnT0ZBgeARYBxV5BZFRjvXh1C8YDZEdWXW8jrwekwyIy
sCvWyeUVeaLmQTafVENA6LcuZahSGIG/kjLBll/k5vGzdGPvq0JSLZ7r3/RcnU2ePtqeRexyU5eO
kZC8zHXJ5Q6HjH/QvMKaU/l/dhEckIzNE5cTgQJj5Lggp74TrzlUc1NXASzNwqheTtsA5+BU+xmV
BPTY/jdyQ3i8b6bABBkCYqG3e7snu2fRoa9ijZEGSt0q21KQ6GhU3uBdR6LJYlKWE9xf+lj7Vnsp
8XeZoqnsXTP5dICk5jOn0ObCc29CGdJB9KtfgO+R2kXqYMxbZZDN52JUTBvJz3/x9gr1yxqz7dOr
Ij9asTcsITR6nVtgPanG9Nk3bU1TC3oOELRoL33cK7v4x2wZ5rWZapR/adx8D3hMYwEWk5Q/3Bcv
B3AVQXyjWf67BGkz5egZkFkDwPI4ITr+HgNgKtFgioQgqH6E/UonNxUhReE3Vsyw5AaYpTS2LHZc
lPhPZMqClkfeImc9lCZtsjY02kURcVXjvmf3jk0vPmtrOIHgkL7I/Os2whI4Ffoos/GwmmPPBAGf
c0XRhBy4QxR/k28YcoZ2e37AQlCUbXkRwtRBWVCpovXagLvhUe5aWCeHREPl9HVGk+4XYRR1f/kn
1hrOdzojn7FBbRdAm4rbdCflEqKnMnUzfFzGxMmmrd9Lc6nPmsrmPuMyYR3UzKsORBoeRnmQeWpL
ILatiwfB99mRfdA9/0RxPAURMc9SYigxOckiTKIE4rFl5WHNVh9KuWS42mHMpu+Bzwtl1jM70DcL
UpiHtoqqkI5JX6DSO1w+7KD5c3KZ2JDF+NfayDe+ceFpF0RMfQwt2s4JpaM2LbQk4h4IiERri6tm
pkAjKGa/JN4KYbk0JZHBjusywvJPTnXlC+E1Pyyj+WvyDytbQNKeOADtvbcwvi6l9u+yV0CedmqA
p9wg396nfY6lJ5iGSeIQekteRyUEkFI9QFCcJnO7zCHZPPbFHXYOP7WwltWRE3/wLZ3LWOv1I7bs
Uznd8taEv920kKzSZABf8GqfEujC2Nf89O+PYCqG8C3hrmtVkzxuHr7GeQtDvZwyvhCHQoLb2VBq
/+Vvs2Pw3LFSeqX8xiHH3pKp7h31d8ICmp6OM84iX1pKZEtIhlO4WKqooNRNNZqLmMRCqbSm8MT3
0KHl9VIF8SPYNlayw89+JT95GnB7i1DkuZ46ivRJAEEdUbwQEwAcEI+CSbQ9Sqc/ypyey1jKnT7P
6CYcFxVKmo65egUqK7G5v7yvI+XKzFLcHy6eaCmTNRMCJwRT0FuWk3m3vhRUGLhblGSgNQr42xil
oAxCt2e1u7Q+ZmdjSeezq0Otz2cY2LVaRWCRrm9KEf1R+069XaZ9ziAgOeifs/k20zxJINWZITgR
WezOCDrrOkL7NglQkLCbiVYPifK8WZxxerxLxGJY1zDHmFbjma7JxjDJBISwXQHDZ5VbkXMjkIs9
PPkAkFT6LTqWfCHKwr/SF9O9LKznZbbcoX0Wb5ZwPB8xPrZb8ny0cpYhN/Quc7wskrKm43BqX2P0
L3B08eR4+juhXUM8+b1pvhOJ24fbLiM1PyjOc0nOTDKnrn5RzkMdLUKWwor6+D55q4P/BlFa5w9r
7Rvny+P1R6tbH6O8Qw4iASIdFdcmqLKxf48a/Ci17y2filEBnZdBnJkTi/VyXfHQQsAHAjXnrVxw
bfxG0jedwKleZjk29lrpGTs1t+r5MinTVSqtBn5ozArUHneD04ObB9Yi1bvJ/ltrvvBoeSN3VmWa
97ZM60+QZDMqVJOfQe5nM6vivif2LPnXloNpGqA54fT7R6KnIoQBUqkLZSYiJPhjUOZ4KEsv+5WP
icWsp56de/Hj0ofGVRBZqkqbBWc83W6w93JUAuEvSCS2Bp5HTh9ilkg1t99ZUy4BX+RmNlCpUylw
YQZH5TJlLqBE5sygx9llP/SRtOyv1lXgtL07w39Vh48r68Zr9ia2spH0FAqduJ32eumF687xlXjQ
ftkVQN7FdLesSSykgNKp/qmni2+/f1rvT6mAre2KnWhA/lW6ePnh2eqiJMWnEsnC+UxUCUtFpINZ
zl/6A5tZuC0BDU6I+JHXGgpOPf+CLmuTZ0YzHvaq7fu3GRtpY11bnnak9MN7ZjAZ8UDv5NxzYstQ
9ZkywMbKKB7Na8T+HqvWCB5M9lITWTW51XsfMjp/BALEezOFu8LPpsPT2jSPaA8gWB8aJcG9XQbJ
CNGU+oRt9GSEsMbwnkhXSuTwqIucW6cGhKL1wOhLGt2KltwMS+9UYsYi87Ed8ldPFAjrGfD1s690
zHC1mfcGmfNB2q4QQTNUc8GN561IuiL7UK1s/dzAgMGtuKXrk0SUA2W+QwjvpdyfoKuSJAXeac6M
wzR2WDh/gRZq1BrczqqicQqgDh3boAWowbew3LXWZANEryKAxq9L8I7EnSzUIOuRCUfCYC70LbA3
CL2Vp+JMNiOrvPQP7xpQrK6YsGtMfrnyDMTpQ8boO7Ciy7YEx47b0EXArdsZPsLDoyTrV+GxmU6J
wuUZ9mX0ZEWEXD5zjTUgtuytl51/VsEHQwRoCSJvZ8SnoSXHnZHzoQSbzVdyknHfphYUo9ffgAGT
neeQWDeszFUHEg7GPgoK5sSBMhBvf24Me4L+B50ZZhYpoowM+EDdfzxFPNqp4lYSZ8i43PubEEHa
9uFXOq/NPxy2rmDDxdIuU5GxSVxn/e18Y4maLI4bnPQXNb+JvYIMfOhR7/wiBE4qFLHju5WGC3rs
CXwWVTggX9+GBo284GZvinv0nTYhy8t+djj6f3UrymPJz39IpPP7+Q+0NoFcl0mVa27odBudDrkk
aRu23JzCeM297WzsVD59YJCGo3FF986oSXv0mcnfht/kXL9C7JhePXl4CXCr68qV8V73meU1G/eg
CEVwRk6QASfIhroIRwGBLPi+FbhukCuV26IoNKVghAL7WNATK9FCZ4Lh/m9ERtbg3TwGnGUQVdIo
kiSv8i/LNez6F1mPm9KjbiMD7gJzryGfr2cabRebxFf06GdxVcQ8SVyuhXlg2j8E00/OaxtPARjY
QGNLFiyPeobvg6msfYY/6omo9TpzL4nhgwXSyXjO+NLZDP+YWGibaO9PExz0ioDAXflyfZwpZgNK
5nBSih+EYHqHvLuF9X1YxpecvOPs1K5NskajkXiWPW31J9TP8Nbri6w+gIWC8BdlJd4zV/XDqY7Z
ZrJx8orywarZyjBaIOD2f7b8cUfPqn0VoQBw/Dn145iGsHBn17XhsSpiQwedN/+D9HOe1nK/lD/g
93B5yF2bnZK5rkReQVxWtXV/hLmI2Fh2zQXXyTVqpir8LaQeMXEYx7KvYr6ci13IcXt/a8ICgVbG
ZiqtP1hZJ/3h0tpdTcHX4zYKTDAs3GItmwSErI2KhJz6KjrGpPqRlMhB1VDf9rxEBEMINcuVj45r
QE9E6jx6pFUa76s32Jfoje4sy7hcIqsafbFU5nE0tP7p0EXzP9Q0Di3GZE9pf7Aq2dSQkWxm9wBs
iG5wPTGlfevCsgtFqw+PeU2Z0OCAbS5OeWBFyWWb2IZTpKBpEYTZt2/CfduibRJfv3Qe+VCsOFGv
vg5MjWiuCwO/5Enn4AsPeZ39ZqgQQbkWTa+XtcnEnOHk8CILd7mPvWvPCuz5FPXlULMLbqjoG3LS
i0kCei1mUzzJxRXYEHD6yRwOLQ/uUolpMIRkUByPy8YNqdVRpB+SqQEtmhM2j/kiSHVhgv07x3Eh
hHJs8U9T2adoqP9VPTbrIZqEIdwoch7RLC3alNAgarSz+zjwMv4m/ENMoHMbK9xvS49a0oDNpRiE
PksoNwRvzioJSsFs/O/wuAO6Nlee1kBEUzbjWdzip421ZDMxhB66SUrzK0sXCkJz4l0RBlaXjZkf
XkLNPN9/TZyZXF51iHODrt8cr/KExyPZ4fH71LxF+F7nwdoKzGVm8Ts2Mv6sakasaQuHRiVa73Ph
R68TuYwupnUdHrcwXvePV3YKzqoQYmPc9Izqaqb0tqiwaX+smpyU2vl7IOPGUIi7EmAAPlYULzhh
37TnuUCFSZZ3C4SwQYe+i99E/5+EXdd6oP4XoA9rvEVo4uWsCGUsDRIp46gXux5o/YzV3nf5egRS
q74aKm8LGmNLMKGaRxBeN/Wf2OLzGFqdL3EmJY1UKYzuS0Uf+GkzheXDLCK0KCUQRLvfl+tFGkAe
NURBVwWYJphLGA6BT5n4Sh5eT/uDtTyYFI+LRAi3HIYkkxYk4uWQluFf36ihujX7+vkr6iFaO2Kg
seeO0Fi6o+F7nG+jJikaAO4whZCP7RbK6NjICNwOrLiHpPIXPXA4WMjKQPlJrdf/YMuvAVBjBNpG
tVyS7F0Rqzj3YXGtV73X9ZHTPDDzZAoMt0g+rzYlKAy1Z6DV7e6EE1q6z2dhCSuUho64LRmWK9Ko
XdpMobc9AhPb3JIpUpDLK88lJALcKnnkLrUyaJoA9mMy0CZOFiEmkADEKo7JwtQO39tYJV/EohA2
fUMAitMzJ0zXZs2FDSMNodfzff+PihtOteo5Eee1fwx4KUAgBHPY1H4jVEx4uQR6IfZ3hI8EwrX8
BgeN+bnQRCgWc1erHXxxsZ96Gp90SfiYxxQhbJITyNqTXUY+YwxhUjFAmLbCw3e424nfartk9C+8
AuTVpO1y815COeN6xrSOlkHACRikmqzaqUVNlvO/3ZqZ6DmFNpj1Vzh8LCNbDtItHdkQvoZhH4yt
5k/g3wbBcvPaVy5KVqyVPrIZTQBSUEG12dbLeTWHgyQNNIp4t0nuJ7sCEsr3q10wMgZL2Du79o9P
jIRBnYmqRgaNpRSKfteiUNDuntvj55TPQNRV/IAMVnsGA+ZRG+pToZM6lRM/5fSlQnY3nbJOHuda
WrDdBdurE+XVpG2okKG5HV0VmSgKtyiGYbj70rpGK5NON9M+bvNunbuasVLznXuKUkZIkGc2XSMy
WmmRL6PSZxddBqJT7Fa5GWqtmiT2aY6Ws4cpDbisz2gHIuALR/pmMzJ6pYlFLyGHY35GZ1uzI8N5
WJSDcKydyEKi9ajq3AycOPT+d9aHGCTdQ1KFuZxTnVYiKhRn6RbNzlrpqdWb7f+CgBB78yFUpQum
PxxbE3b4/nUqzusLH4g5jGgpPnm87gp+WQaA4v504pqYVw8wNMwKJNFZRnRh3KEk964hiW0jqukI
n4BBcJUgX9yyk+LYEyHPr3BfsYhlwjgZYFZ3g71wcPH/ajgmKl9z6qcKYj3yWnO2A1TM4bR0RCnM
K0N2RSwcCNCsl8u7WyvPFurrmI6J0lcffQrG8pGbFL0ksbEDeHK1K6GmYik32u4sQQNg352WVGk8
dyc4ykv6wYs8tbRBwQ1hMzZpBnBTCZNO281WzeJBXE8JrGmg2qkf1G4Dk85AmZ8kGKftMKvimQ76
nTKq2ezgDFYGiamwo8a4zLQZNrhwuBRcg6RMJkh4AB14WQga1HcaMeI9dfWAZNsMH1K0n8/qXlPC
3q4SgTxD0s7a609xIM06tFty1mUTU2gBA3NA0DUljJNEEZP0qQKPek8EvJzF7uHwpIY+2qB+rT1F
WQbg0f9Uv0KGZJaaDhygWZMyytjN+8OCBnRf2+IUyYETikxIrwOnurNwPih6XyHxjIqjwO6CGjUK
e0xCE+06Lf61KMAhoExeCgCI+GH03uFx6kKbOvV42QSHkVb1X/GblQciqkEW3CklZlXrBCJqKJB+
Z1Cqb1BbfpO1MWxTLai4ni1xAnDqBEkmXs/e7O2SDdLXmVfO1zwItUXK+MvALSGW2tY/wojc+XXf
mebCfFXvjZAUAaFWfsPqXDQ86SfkYTIenh2iUf2xooxyHNUydzkLWyPqienkgAnvQR54ptG8irlJ
3C8B0Sn5d5gOyTERN5US/+5+XB5JgWdfTdqSAFMzChYb8v6ZvoMvPag66t7eH+uN+Ti7qDcSXRhC
fnVRFaG6UHgcvrHZPTpMZ7V7Peu/2Wa58ZplgBskBKy4zw62iZmj+6bz+QrH9HI7Qs7GvAjA/JRU
aSRFxlxUNYAuXUUf/V2G0uh++nTwl62CV0bWWWEwcUmpxN/plBP4ji0C2W2YVgaVWoLDf5O0zFXb
DD+VJrZaSf7x5z7I/zrw/iQfOv0ofqjx+qGe8g3ayDxBukBrjL8Y1OKBcsCkrbeniZ/MoArIO4ap
x9McL0eLnaPTdmsAndaZyCRtzYSMUM6/xW+KX5BtBcLK85jdZWkdtdmLFSKs4Eqsm1aJ4bHLaZyI
Ofiqar8EoZ9ISG+rlPoYBXvRLeKhDXUZcveDNdfbp6cKNCr/s2yG9/WYutpX3A0fN/VugXgCU58Y
SzQE0q0s7bqnD++QfVp0TCk8SX1J4E0ljKDSx7rkXtOPM/HLxMy/4GDB/GDRXMXmXUUTdmswChPa
rPD2L7z2cfDtmzjpRD379blGJzWYXmtXF0FcYf4/cpXg81iTjWmf9KhjWY7jDHdggYK4DPm5CE+u
AZidTO0g+edJtauZEFaJDeuNPnICrWcZEn59rkjsiE023LehKLkHodoZ82O9/Ds+vgqLdS7FZZMK
YsVtY/V/7oA+CE4O4QRnIE4xVPPN+VvVvuwFpqZY14NqNLs6+g/eotWNtnsr1xUV6xA6Kd1YBPqW
Q88ONUrLCRB7YJcgmEPpCcR1KFfUy5uk2klX+blMAa70qo2for9BA2NZ8xTXl32XLlvhQnWjlt0C
BrDsVcLpJj38WlhjiKMQqPNRelXsiYU4NM+uIh+mwmwIOZS5d8lB4RxT8tj9IjxhANdzmM2o0ReA
NsLpnu0jAVm6iPxy+UdxTykqmZH9wgsgGexVTpzaEWTL+aCtjhgqY9EaFO0Lk5sID4xbWQBK0N8b
vyY3VCxgC+jpV6hNQipLN2YWzcWwdQfgYuH2Kg8pu0/e/vzFLzuSrGz6eCGTcmGz0dVw+EOgDs3H
HQazOuH2KkU30VrhFZeqNfXB1+FNHJe74cmyKlyXLNa9msQ9aXigQBJoMs1TlmvIo2nb35bi7XR4
gL1IlMgzsZp+tUQ3keJiPjL3vZE1MpqUaV/7FSTNtacasj9FRNwvXagJElBaPWR/w7xEBSb3gr6h
bdaH1ug+BEIH5Royc1gyOy0to3OO9yWbtHZAJ+QqoGvk/m7A/ys0kN2czsY44u0HzLsY7SZauXDb
Aqr7Zlua/LE8KReWdGwlxmjt7m0eLtd3HJmdHMDOrjtsvmHHAGa6zpmkjs1pU8lbFhUkiFPEds1b
b2GgOUxm3UAVCmaA4IP4tJ/dIMJ81uJMJ+UhexilLLH7qEAsBIEFeRKdew+b1KiKziAtL/UL6GM0
debd0GQb4HD/QjtTC1T29CxYtTOxNIkvMzw0d0LQMLDuWmIoxt3aWkx3OM8+qcop63vO6cZBUwlw
9V6+ayQVrVJ1JmFLP48ZgtX8tcMwh0m4jvS1YpaOugUob3AxvLu2iHqxjIDMPrdPZDZ5wFs1hPUI
WDVMzCI2WTqWTDZjVFA3wMq3gUC371FTPCtQeaz6u6piwkIsnL7Rp6E3Hrw/bkm3cAApm7/8ia6w
TlQdFaF9ZL6TW2pgjbAwx617yfqYrCaGx+be0kgPqYZkzpRAhK3hjFHYmYRtcf+ZIjRtNghl3brr
50CVymj279lel9T+PRcPg6EjPKNqPmTmA9BqDykNZu9ANsKW0lC+NpwPRTpKjUBdk9fNQqQWapwX
fNvZx6Iw6Oz8RRja+pi0/Sw8PpwnYm3Rbb2Ow7xYeQ0xRhT613e42K8Hi+K5/hFf7pwpisiQJcy4
ooG3libWGLS8uclhmD6UXNsf+R62uixKJc5Z0F7SSFUaPhFqVAsYLuPtdOWJI+EMwJ6KF44MDUgl
ignAWxWQtQMtvNEyLinj9jR7/d5HjTW7z1oJ0Kv/OtVkC3SkDPwLgpkmxUm1Fzv5Q+sveYiTbWqq
F2LGiJH7Awf5CQeegSVXN8PzrVk8X87ZlBsRtjalj6WNjG81kC9QhpfFqwYcDzuHARWe1e98PRbJ
sFwDQnJXQC/dsnxU/oSXloCD6M5xWaenPjovfr7Ku+VSmhdqhfkXoj1vADRQHk4bCp3/rdBVQ1mb
sfQem8SbUM0qE6jZ92+E62WjpB399A5fszPM3h0okrFsZ4f1ODDJtQ29XRbhHHg1wfiUriDHhh2w
HS/noC37FS7pnKZsj8LZMNeqeDQW/tqwbmx+QSgaiqn7AzAbqQEs+zwxVJZAKB0fLllnQKm+26Lp
U6gfFsFBDZ9XCc7yQpUwqzVnOWm+7aXtlQxzFP79O98zz8+0MxbA4CxOEWn2NW4AZLWF5EmEg+ee
5QFtOEJB6ThNG4JlZXoD8Pk+KZUYvb9WQ8biTtzrTKih5dSc1+OMeniutrgty9V0mg0AuUZKjomP
sZ6JqQSbWSdIsnbu/u7qXSwTtM5fuy+I6/2gadwjqmwMoucyWBzm5PCUOHFzpqLLDHO5oDzJrfDK
9BKTBJURldMpNWa44QusRBnrlDSy87EibbDO6m0KRaiZDNIcBSJ4MwXLOfALZdzr+cFAogmID6fQ
9JGygh+bbjHZ96QkjLeqcWMqN1BsOyqfEb4xWM/8rZvJf9bZHobIbcvsx5CrofBZKHPifx6/Niva
9rLxE1rtZeOhHGyA4dsiRf9PkLMZFaaecSWbzx7uf0+0MxZIdMSZPdRYE6v9uJ0F7oqSzfAGG0AB
wqsvLcltJSBv136VesDndUErZAjiix94cSTJeMZght8pGMT3KMIUo4zv0NhJTQ96I65jsbWqjRvW
/mRLrDeRgOWPHcOt8LQIxKWzGPPUU8Xx/dqmHFbkmUCdocw8GR4guih4El+xRzUuKkD7BqHC2EOS
K75MDsmkrI/euI7q56TCwUjtyVp1MDcpt8J6kDvYcB7sD8nCicAFLnxO42UmN+dL0msQIMwkyYjL
WPjcratmG/BKSlEKAH3B22Dd6a1REuyFH7Jf7XThz9KfNHo32PIc7+BmKBzb4YorzW2EgknMcS30
XDBqgnI+ehPBxyRoZtxDa1PRuA8dyjXfyh9UAZ8jReEdDEjaImDFiu4K0m867rtocSIay8LlSTAI
UZXQ8c7k+OW9yNCoPgmfuOiNgWVrTjthk7/UmSd9e32yRZfR7mKFj8g9DLdTaGMOyYpsr/4OcPja
XJUfvvMm78lgNu0C+lKlNhFjdf4p0NoMeq0FpD8dk19beJTu5PwQ+SmKw2i05Rj+F7fFstf4bh+L
ey2Qs4Nf3ttODF/AgGct0xXrSSJqvBIJEZtaEkswSn0oK0mPFRVmo02cqsFp1jkES3NGFpxSmyOa
u35M48QGoAbhpgK92kZsexP3EjSDxBN8ajD+bNSRXRiNUTvVEOTxy1fCGAYaHasX6Kbf9U8AV9og
AaLV7UtfJTAKoZYx0hUwTVv5G2fAROelxO1qgKlSI2KYd3posg22UBlaj7gs3qbRGxFc1aRCAAdU
rsH3DcsUWR1hVIlqirHmOnjrWOFtV60xOkpUIgz2KpG/TOgeY0PCghtiYD10qdmWaEK+km5UTq8r
9Z902alVTGHdgQlXiIc1HCToKawvUe+OTVfLWYCAR2TRr10HS7ZxRseG9f9LOk1NZXvHBzp6KFcR
fkYL2QCfQwFrCVpF9mZbQDz9iYq0m44ilfLPx/FAwpmMYJA5clsROA7jPeBY3ATzm32YTOad2Uz4
7OxBTfjwfRGsuIx+923jkkBoesB3/d7pbk90l/kerFzfXE4z7zF4RnFkPVJx4AvviRoS+W/SRNaL
NDqVwm+fSbaGSqU8+sJ7+IaLqTr86z7QyDPmxPwf/9kqU7KOBUJA3hzfEFOUTQNHvvX5qEXxDavo
yIYUUvJ6uJET13TGqIQq1pu8bdGnBzSI6hflUyZDoCOvqH322qxhnL7gWxushDZEeYDhGN8whAP7
XWxtqf2K+SRSNuldsUqd1rGz8IDtrDya1c2hLQi/2sI9YoYBmhmOdGtQMe+1yJwvMZvFvHEZOPB/
FqgydU1OzPmKLXur8wTwBntjDJz7fwOxzal+OsyImBRV0Oi3q2MfzNZKzb0CiKoBiNUUSMs68yJT
dzX3iH+du2CSzVaEFJRJ/tUYsNiltr7keeUUvAiMyV9Z1KSGxSFxCIH3cSzCO2OtjVSNX+Qz32/3
q3RZy7cyLIdWE4VXGD7Z8qzcC2k2iIXb4JTNf+yMg0IB9RrDApeq7W60MwpI7twdDTrk9bkZLDHG
06os0Wc1gOsZHhOGaRQJle85nrLNB0HcJcp9bm86+4uixhDVXSt/gB+OhtXrpHncgKrqmAuZZV0H
NvKteiacAYnMJSaGRvIkGKCrFrszj4MYU1QXHSa8u9ONaGMZOXMSUqzk3fi4P5hgCapq2YGkX/WR
XaS/fnfYova+ZTDvLZuodz/HuxBKaHS/9vBij72uA3wMKsVMbKMdFMPwY7DEQyEhVMJl2uROIlaO
S4gPDXqU30ANJRXpcfsMrmLP3zBH5r/M5A5YgNvlTcprjCHaJb/NxdT6EHrUDmXvT8TWLKIKbtjW
IRIJHAE9sxVHoYNOf6T9C94cZjl0DrUiJRB631bBeRUclMcKhBcN6zzoFGxPcAOQrwVcd/9DQOHO
OGpouhaRdpEVHOkcsIdm/mjH5Mt7GfBeDSKsXjpVancGH7s5ATnktjeoTvVmWidUbty/DbguqGQt
n0jpM/zNrJSvWVD6Z7CH5YUej+9Uafw7D+WwWMRqvBMeKwyvSN6flrAaz30kZ0iv1FChe7vjirTs
bbXYliu5xv+KpG9kNkATYPX651qeYgDzuD3KE8My5Nx3AjfzD5DgaQ6MnHi111Op5wo49v2YaKFr
nt1ZKwS+MwcnpFEm4O90GFzYN1vmWeOLscZKNJGZK/SC4KcEQ1kk/DPKARysz7oHQAA5XxJLgygS
v+zdCev8qxDjVBqmq9yQVvRzJqqDg6PP4KY+UHUP/9onuFgaMPhaeEVASYBjaQoGF7HIA+4HMfYK
FEnzy4erBxWnu21WS5IWFt4VjZ6Oajx/Q2pJGoVXnWzjkJdpp62Vd7pOYIoVRZoI+wSKvVDKf3/f
y0g0Pdom20tzemmOca8hOBlBE6ZvrASfu8SJSgrtUFpd3lmLv9f8zDqwtSGlfe5tZ6bKyd0m9SPu
YZ4Pcn9Kecg/5OnvHGSBkRbOMJUizQUw0h/et+HrhZMEnr3LJz8R8eOyQpOJopvrd7KBL+vXfXId
Uo0T4JP1H2Qedm9ABa6xK6vVIcX8ttNCKEIikjv0kQSDThhYYCbD0JrLglDVDAS7eS6DKq+iMu4U
rRn1Mn5h7nGs0qGx3hMLln9ujL06dMsv7DumY72nDgYSa5R6TFqo+nhn5jnKaoy/to6wosq5xjrH
WBrG2467HcLxrMplqup+Tr+XitLZGMclyu8GwyiHy1BEbkamHCraXZeH4HzN+3Zm9iwIPI9ewquV
Pm1Ou9HCRmYXDuCx53RPN3wB2a5IEpEQuDCQvLY+qtEUhpJ69ntLI4izw0Bog0BuKx9TTL31u836
pe6PPm0gvaRetitHpv4/N5Bcd1DCQmqMBk8jKxfWX4u2GYrCtUE1x38kBMsnCsw5xY6mzcDWO+9l
tefKMpOn4q/eFZ7NRj2VFg5eCpJrsONXEy0t9qtytmPUPCSmusRx7hEqnrk2eoJwe2lc7fTLROn3
tAh8pHn2gfhE+SHVIoHd5nqBxecoTraSR6eLKb9u2/AYb54ptWJjAnZjEXiubSmyUUEkiQb3xIUF
Q+n2iuG/Ho1l6yZoHEaQp7wHu1Gyzw7gK6/SMN6ibSSsKapdoLrS8yC3rk6EiIMmgMjPjwVhyYWa
IJ7LP5Zb6b9+lD2PcDHBs9zcBCsYsKZ2cr381+Ln58nQT805KnvSHkgHEdPMvRDTpNtbQw0tvZpa
LaYve3nerWLb+DFvWJ7t6IcwsZL1lj1R3JAblF2B1c+o21iQYF1ZspViRm8DDl9LutDwKMOkAV3P
LyzxKNX61Xs12BC2mPI4/1PNHncvHUV6V2ik0WfZ+Jnibya8tGRmhkreOcIEYaeqECDOHvcSTLsM
/6TkpxCnhX8c1ZCSTCSTujMYA4FM5xqImaygKtnP5xieTGZNqihH6gp7n8ViaZydcVINDrKGI0Ui
D6txhlVdX/WrjTuT1Shedhp2xv6pUh3VUFAZ0beWLo0u+Ro6H+iUvkZIeMag9tFZy//cH5hwjQVh
Fe85xdkjM/AJLcyuWKEKxUHyJcPaMhrnGGl9t9KRlB2ryV/0dIWS3xKbdq17JNCCq/b1FaGzs78L
9D3Xmpo2czrR4akHxy147iGnzSSSH26Xfqp7DecS5qCY57BbKiXJJJIkJg0J1izPMqg6NpvN0bBd
dLCOUhosg5qVFdyqmpNDvYayUCiACyWFf+Q3Gqj01ZlAmzmclWuQqi8YwQUIakzGydIpry85xLQ/
n0FT/BKDUhVopr6FNkeFEKR4P4AL/sJM1LMO/qmEmsFZacXDIQfOEAXAOH9+1QZfWIRbsjJW7Vj4
TKWM/5mpZEe/odrJsxBhGhUtTw1q1uHMPn+rHxW3pVEUjXmenp7tj6/ei09QhojDYjUQb9bSCRMz
Imxu+YGdVeU7+Hl/WKWPjOo1DiHdpCDnnJgwpE9ct2pyTYb8vdlFBubFB+Jmj2aRFdr3/oRIaWxA
/0kE13XlW5BRHBgZCbvkyQNdOlUUD+7zYRZ/08iy6B1y0QaW9UcoXR6zTHKfPBImnldUrVB6YXbm
vyOtSsewghkJPQXPu7AXhSeDSgjWXSNiBXw5qtKlsinVb9H/yIWZmexihw7gJ53IDmVhRiNx0nHN
cNUrwj5I6XCBUPUvbRbNKSyDcuX5rWVyS5kmHWLYSc20jL6sLsgs03OdUnJDrZBcOi39dC0e9Jib
u78LP1SauWFWDBWv1Rl2Mi58VYN8ojPvXgymCpFGJlMLEH2mawHnm38JmhGr3OCWLqzykFXOimv1
Mkeq4NeaC4M2ZqN49SG4gVUKgmf9laGPXxZxHnsqnTBWNA6pQJXaeOFMBEVzB+KG1NaBTBhw3bXt
/pdErSJBjLzVN3f4WOQ5Bo4sCU7us4JIXYhSlARPGySefAE767bUtOxmENolMCmPZXvmlb6ZJle9
bXoN231gNI4YxwVC6Nd0D2zxnz9nN2wyYgFbIz0gWjUFX18Mk1TtwrNrm77C1/+xD2Cpa/cUcHaB
j1/rsaIPMuAfASbSCUzK35zYMEu8JCURoWiCy19+nPaijW13sA6yU7Eg/Af6YB3AouR5iZDGcM54
LqNbEjdbKZDgRSpNm/l+WE8U8SKT0hhV5eURGzwUnbh2uTPo1slAgEi6KBGc/FwURvFO+CM+3FGC
JjjvMdOOnLjc0Pbq6jhuOPjAmPRmsdHAiypthBn+6iG8Im15ijRpCEmRzl0MwuPxZBl6FHJpop5w
MJHo0DPtH0g6H+/LGKZajLXxX6JZOmSskUKqlpOb8YW6DB7sgI4dtzmHfgLhB640MfmnZuIpzxor
x4seVuDSdKyHvX4Gg5LWvYXTIYMUqRjo7RjcPv13ib8aIEroK4NeCtDK/JEp8haeQ9Zi9kUpnECd
PCynQRAEd4VMuU5gsUp7sEGy08eYvwTcXgMfH+iafK03xLWqwhHf7OyaaCwjcUhQKJGH+KSbbxNS
kcqVsqsaZnRMdKqK8ckWEXnHJLURFyTXT4L60zw+F6Otx4JVHiHUXSeb9UjS5G5dkFWpqd5qv1Vb
3JhMZ7szXrm4p2+ZwM0Mkey04l7k80X9c3JU6yIPH7KOyi1JUsFLNHtUYPEv7Jt5vNYZCIKZ9/K8
q9QeX/7Mh223wDQTggWjX489mFk7KBNow8oSTwobP6dGKEimhmf+lB6HPL+Zjv1dr40S1845cdcO
I9fFA4QmWWKw18GAC7B+CEN/qzXdd8tOY+GJuOkjCIV3UhxElZzAaZV8PK0E1I4INCCzXJTZsIlI
0vD8HjGwq67/MXgREi5E/182q7ilALzVqC8yZjLxnDfHzqMh3amE2D5o3UGzENKMC/6tfx8vGZM6
c55ZyITWMKJRcCVxcIIbsn1Cn/Jd1z4LYoAZmyP9Sn9pAHVu3unPxSeO0km0YnMm/ShkVIf6q1lO
PoKdTRln9R9ngBxmBHA+AuzfMwcrqe6NmvPPMKwPK5+LgZznrrjzxXe71+DSH7gMey8NNDayhvGS
8UqGiMi0vcuYFZVW4V64g2TIi3OuNz1T05MbQMe1LkDe7nJHsochJu7UH0ysrdicSULtbX32p1uo
peG5YDWHXiAH0u0fefowU4lqI0gaOhdWEpGZxAAxESW6T8mbGJ4ovmSBFdRUiKCNYkzNoRFmHbJS
3RLgv0IJbY5dlSxWw0Jn3vs1xO+anucZFilc4GaC4JG60swwqj3sENFKNxa9pfGWxyDq8wmmoSsA
MNAcj6zPMpkUqjeG1Hr42TgCuTJCU9twRUW/dJ7iqydmywhoYSXNkUxWFB/uuA0OnJBTDxgJHL+N
cqPxVFov/w+dzuIFeslGBgfNQMeSkUv97emNCOT3mYPUeEJLgm2h+lmSH5wmRmIq5HuhykjBdovY
PxeV8JGzNO34dL2S1ux7RYa+Rsl8Tnw4iezEQNdHQqalR/TcmY9d2uUTZZ9H8teOdNrVruQ/QYKD
BkqYLlTJwKHxzmoaPasOgt0x6m1WTB1CRu07xiNAxL3mJM0JAw5z5o4JyS4JlnvWNgxmC1W7JdrU
dDh69J+t03tcTbfM+GyFBs5DhYf2yvTql9uwwfYmpTlL0WLbF/qtBsijbmDcURfkymmGGnYXW/x+
LhvpTcOiqfQQVFYjqcxlX07MB+LaS/cx9xNeGr9Dt5+TBomNZme37zlZ+xHQr1kK4QSO/yh9Dxkq
rU/48fjwDIL7CV8RhFVW9r7noI5B3V9cnEG4SQXpLhTk6aF2rHcF5bTVChCQKITbMlGfz/zu5/u7
XYutWKdoUhEWT2JlUOK1ahLaT4O+/Q9zK67vEgP2TKoLwTpVnjj3DwauYF2ZeMMLFL7yP+ZZyR9K
k8D7QhWfbCG6QLAFRe6pNKv7t0nj7R+MvsBE8cytHqvaFDlpmLA/Rk1DEERW6TG3tRP8RvxjgLsO
hzwGFVJaco+bpuTNjVaUQe8dkoy2eslUYjSR5vmahRU/9WOmJsrIcpaEywhefx3sVr/mxviLheUo
Ga8LnmmC3YAv+Vkrq//zbKaiqgab6gOVmpRIOGVlZPa41MNONcjjbA0e8/cjN2aaMh1bGUimPZmq
OxkFO7bJv9KMTclhPLsJCJXdK+AigAqZJag43ReocBqOrer72HrC2AMhJ3Z+BTpv9kvzALO9mSxw
8iI0f/zg+0qezsMbvbhAq3tm30Jc3SB2KCru4V4afAcHS3qKm7M6SQmQSDX8bChYwvwLgi48yCXY
y1TrOarh2wEpaKtWuybIRU8ZOEgXqwMT2Y9m+jU5jdXM4lrR2q8+J3W3yy+9KZiFaQdotlRkVqGM
uwbpDteMOqBx312VtNVnuUtYO9do5zpjM45kreDvACr9wTDBCZGWv+8oK6WdhMxnU5pQ636KFbAW
q/dlWXD+5ULmN0O4bnplghtzoCcXSw0cQf/Yh4kiQwXrOKgruUWWXYYcY7EbKv2eTBVQ0vV0XU6F
GsyKtXHOuAQv6lDDUoX9d6udN/I0tsOCtyjJKdDyGlCed/X+AFgvMkljCjtzcCLUwykNUY/thp9e
mG7M2oy8xKP6YEAEItl/YLaOsSZ+UuOkHIvFYCoa9q0K/rnDMQYc6x+ZeTc50xn3BueUu1wpMNvH
InGmWRy/eQNk2AIGuCcWVFm/SwlFlK+hdNFjdP7vPQf2bQ4auJpso2KlmYnxggEXdNT6Wm4qw55y
fYNKpTp/6Ed+W3M4Pl2BnaNoOkKoR/EVr5Sq9C+C2XhDnB5C27EAKC1Yj6uqWes7X2ZKlUVhFq6i
PgagNMykm2fX1vRFRMpuXjExShYjuozlsJOO/AB6sZExqJfigB84nvvyvPdvtUTrlALcdIGzj/ww
HgqGeo3nXpkRAL4RPkQ9Yc6ZPh8MtXR46YsMRLThqe/yRgFRzVnk9OIlXuFxT/dpsnUJzcYB2TcM
6XbxvKpmnw879ieEojo+oUf+1Hqp5W4cgVzfAytgOs2du0uIx7ekSQcvr01Ikbl4UtVUGRcwZO4r
3ckyL36qqqTZ7dGfcpSZaCFXRiqGoUq1eEUdNLHkDO9Wt2uTYQER73JCPQdWdSPH0OgXt8+7RlxE
hVJWrhL4jZquZeRtISYPxh93jvId1/LiR3aByznQjUpPdihMyLT1biPkEieSXsRcQUctohu1SJwj
MiZBCRAhZTe8ka6CDbY9jBM7lXyTQxcYeV9OHAZtgG8f7zKcJ4g62AvbFweCZaV+4Ujt99S35fB5
3pf6pVvGWBrqld1ocYC8Ul09eH8/OZMzrRO/9lOglHP1CoY+Oy0z7FqOCqOlMBCfDF8EN4QVqAct
22HnldZXp/4JBUo48CmHMBfljWsTftuinJdB5phd1OFgkCagLHcIY9Kr/AKzj1AdiVuR1aOocwqO
JxOZy2oRgiJdIpTPH44mt6wQGv5c4unUKQWfSPKym3/KwOeKR9wEAv+2yK7elFIzw5B0DjSb5pA9
88JoAAA97Nz4GxffXcfnqtJng7w6hi1iiMbnP6YWKgglYqA1DX5nzYFIN0/59VD4u/jb/GbqXJCT
+VYDpfk14sH85kAqW8CiHiX8NyLV3AuRMl7Xv3x8iYAntw8LxDTW42uHdJyWYVs13SyI8hOXqgWA
dIE1npmxnOiDXc6l/uPbhvFesMKqVbuF9A86Zu3N2D0Kqqc0ro+KVvHQybYt54B7DDz3pmx9acB+
Mjs94McGyhCy8jxbHVugvVig6nlOX4dq59xrkUlhzF7POQtX1MerU5IhSPb7yW9B5ZYI1Cv6bKU1
LmoeeKDhSmI1I5+jhosDwRW/hCD38TXPhJXnP2/js98Tpu5j9lk6+bQEFR6uMSmcDJCyZj16Fl2U
oQ9KdFkjCXMt4au2u1UGnSRSkUo7J70//DhX4BRCZB2G9sSC1BgvnVT2V58l45qxBFyZTBRoPb/8
gOOJIE3MsQXo9TTDGpYzlCVRQz76LER81q+2HoRko26LfYMJ340b2RDXbutnz+Z2dh0TkImBoDPZ
hmBiyOaeP2CzgppULGjTUzO7dLVvAsrmXZajIle3pwkP2KpEJUPc2JnOzwCmG6ocVmgO6JFpGeFc
K9JxM5iE4v9HyDlmpzv0y5/oVjwxYgsO2NwCUMkYnL4leliHzU9fpnXj5Tq6q2xUg9QYWEBzpWsD
iSIGU5HZzfmmYsRmJ1y67GYo+BGYrgY3XwjFX+EHnaEKz06Rd5u4AQR7z6vT0POHlXI0+Ndps50o
k8PbciN7+KaDMjVUWvnVf0ZwSqEBIEKegPTUvnSq2b83Na8xGuPw6ARFLlwGws/CKCTw8lZvvteK
nY+yb1ypj1jl0NOsQrawwiKYW5O5N2Vesx6M+sdamQFtm1fRu0bLhCjP2F+R6sHVNbft4e0GdrVU
hinaCEDm1N9dk4NYEiqiwPyN38aBiQHHxvhNz/kd1p1f7ZiiNCE0UNGh2izkIfQrNebpSNkeG0Ak
EUSy2h/EyG+kqjvBhGsJYnh/QkVrHgdq8FDUQjUqkxLhOeP/o0xlTNsvMC51fWyxpvM8zi/HROsq
udseo7WKPhwOipuL8ShHeTXZm/nn4DWzDcCvEpkDZoqgRIrMUKtSjVhOg2nh3Rf6fNyvv/fAlCs+
Qc0OC9JmhuPrX2k+5cIraEPb2dJJlKXWClMoCf0rx5RcbLMSR7DrvEliKeemfkszkq257wyue9Io
MrBImD4L08y0r9FLq1gFQQCd0tpELGFlrToVOJ0fm4k/t3IuvDdIAcfMuB0wQGXFj5S8GbfWsq9T
EyzCSvSoB0tYiyJdkyvZ7EY+fZUofoDDTv2IcgWJe+4zX2AMth1jSMkBoidTWIxcTMFhkNbqhlm8
dNUHXl+fFCjRh54aUk67hpZKEtZQNRs3aEvAoFL0NR63GL6oJhPrsBhsSd5d+TUtHu5uYWzVzE6n
7/uMWvNQbPBdvhFz9FWdkN5vUOGPDNMy/SntnoSmTUl/WyW9wki5s1sC9niXxAWxPAqpBWGi+yId
mqSRBTfjEETE3O9LTfYRwuvU+QK7UHTPaaexRUdQjEgnZL/JHW3OFuCfK4CwN5GinECV9QX4+Cd3
6OvYUvKjSCEX0hN9RsWRsxZBKoIBLHZneXyyU4hnnkMYA3SNxAezYkzFQ0Pc6C6ny3O2AcX3ifCQ
ubm9K0kOxsXN0q1K0uZP9Ev9ljwhT4jZxjcXodSMPXtGtRW59vSFJDC+w1fkbpC6lv3sdMQEfoJA
Ms9Yy6F58xHsTAx99gR/TMpXXbktnZBXXbuPIp8d7JD4mrNvuDvsA+ATDmc9qtFA6x+sipwPgBTk
Rc6MoAxcACUIInCZKlMAaYL4IVG8mPd1GYe2ea4f01hiVsUMGMsM4iUUK32df4XtEZGZxbaodEBm
YPl3CcG0RksWUH6eXMxZIoz+jhPQMuoClIPGicLcrPkz4VZHOAAD20RiKGPabhdcSA9ftlnqtYWs
0OLAbGqH5XLdzQUGSovr9RifPVVdkiN9ypiPD8XwIcdbG/U1iNb/8bhf2JoDerCzZAqF69Tmc7UD
ahs19Y/1FfoKeOHh4fzUq4HVhKmyCA3vARKesSIb2z/M+lKIaNUt66rGHxc3g5xtLGgtGivXSIjo
l3X+y2uR7nGdcBLpK/T7b9r756NMponoLJ51hYndMXue9YupL8y0H0QCLXc13sgwx1nM+WeAUmt5
HSRrsn0voMV3ZUyDMSShzuUJAhUyPbs0lxy4V2eLv4LYeXTLeKrG75dSo82DuPY4UGzN58hleMJh
ChSsYrR3Cd9FCz6Z1gsls2EIlPaJFY4hmW/G+QBZgwQBNTWpxgxaktdxrBTXgJtlNCKjpQ2dPnUu
l/hr32pnGHNGv47wwztVehYfYt8kWilfl4EMpcesRz5EdzeE+scsMJACwnR+P9H4a4Mkruh+Asxn
PB42gb8t+7/W12tjWYzCwwEgrlYCJUZpUOo8bhCfxMb7aBcIFVj6LYIUbx5jpOMZBKLZA1i669H3
Y0hIUpNKWOCNhFTo1l0Rih3bpW0TtV/I2Dyli08mulSm/OO6Q7hUIBWA899XtDcD+WwuEzmWfsNn
kHfjF3eGfWzFzhi6IMDBx+Jp0CGRzOij8T4+rAUk4gPaH4Soqd70x00DhZzH11JR1Ya1t9RLW8tr
hJeOvOeqwqW9WwNwBEJwcZrHAya33oQ3fyzXtQqIJLpRaaYXXfkX9AsG36Z2YoANA9ThgsTfd/zq
9MUGYBrYGWuAHM3eTUCcbYgccNlm29xPubNetHHqp2BXTq1tXYjswXjRO5uoy94iu35iSNefCuSZ
Pjc9tqBl33hVx6mroK7I8wMTy9N14IldCqFxRi8X6JWt89tzh0zFGuy4tQw1BczaXKp1vFGUwXaH
xPyQXgezXfdGcOPoPyQFb6Nx64tYx1pE1RPdic5p/Nz9XFSiHKIunN/qY/MkVvSgV4qvvpjcdLUV
kb5AV6lfkduAUsUu6Ojyzh5KxoycOoQHLtKEqpwucerubBDeWH7yv6ByIsMFmUB+XT6ns+9aee+4
KJQFqj3rOsA1R4L5vY6z8vND3ZcYYeejrugm1j3EYnW7uriapiFRe3wJutMQQBlsg6pGv8ueKJJM
yn7zubolMhGUBctP7LcK+l8+aCscYGu7Lh048wA828gfMirLS6fJchdU5p9xeSgh78+m4M/isqvo
N3tLmVOdwHGNX7yRsOwfgpEszySlMQzw/Rf14Xck4roL7PgtcXRXrptAqVDFUS0EhNseOUNXt6WN
s4Ke5mPaEgPf/Mt9ewqUZcnH1MTBLUND2c29QzZi+CQP2eycCbtuu6yDpguR3E20zWTUzx4omsuR
FMJqNvowfjq4A+az3myGCdWNCesUnq+ba4zoK/8ShcdmgWXWTY3KSVWMwzU60XXwnWeozMi91Tu/
/1EeR3riJ5sQHBWxHZMEmCt1f6DQOsp5PCWrZRLD0Mne8dlAfKom6xJD491qAgEmpUJE7ZYo/E1R
bNKVZ73zT33HAaOZbEXDR6ts3enF+BYwwLh3i26Cq7H/WLHTHuMrq45apGZKAlEN7wDYH6uiAnGF
WirstU5JRMXcKtFmCFgX4P641nf7+sIUBkUbfu234kuTUk9Evpwyqm3jiUa/OpRs2ZTMAMsjwFar
jsUmt47CD+88LslOkuBo47HFPLEW3fG7ZrVG4WufjgDMVXfRpX18U4C7jZWWh8vQQ45imIF9m6X4
qRj6175a3GyIEYG+ZuqRgs+L+UM3D5fmRiiu3zZgcxcdUjw1woPfx6YTAq3ZjL3Ezx69mp87uApa
JDgRkTs84xrrQItIko9DU5eQw1/xm1s5hZZnGdxeweYb8r8F04Xc4FANlXz3m3Wj4+kz8C8SHk/O
4ZYPlMw+7sfpHUjTbfJHJiYJdEr2a9dKVIl1ZOHu7WkIi9AVPBIveGmGLNdREecxrPSYSXXXQQp2
syKUc3Pdy4ELlJ0aSXTIAzdDcnAff3emHkWYApvIcclY9zbgXe8d5FngqfpCHuN/S0eNAyjeJ/U2
STcIhSKRkCWpjTpsE3BVtPgip9XQVIMksoS9fR1lW/QUhrDU5ESUNYnnHwJsjuEEIB9Ld9AJ1INH
rXDc1ysmh4bigKmYp4+rLa9/LCF1p1yZmkXs1ypOV3mCuNB4rLs3Uikb4VNIAjnP15jiIPov6COn
EZLlZVNzpfs079Vynu5S7YLFRO1Zp7OKu+4ITnfcOsmya6/AjSXrthxQbWoPXhW+2y08gBR5U3xV
02/D+ITvCPXv7FYXJxeOmP3RXABMh5ltKDhBlSn92sj6Jy6hbe1jY0/7xrqHI4J5RL1As8pEVb/Y
nBS0Ok3m5muby9Sq25n0JWU5R392pBxbQA46OMnlsCmW9y3y3n3Pf3oN+kki/GHJQp42pYbW49sE
KWIE1Q6MPm+eSSBdulza1C6+dTeYJn3FdO/92l7SKCIvDBY4BguIgxyk696Xm5a4dtwrqv5puUDY
gontMukpocQOS2P6B5ptLoK2pE4MWwVHYY87t4xURv5Z2ObsSDvSoPRCWejwyMbKVRaiydIx1xBr
CZ8aX/PsLPT4+uSnexliYVRlzd07yI5DKW7UwwtJvHJzxIDIylQTGg9/7uWwvXDXCqedrCBb9Krw
iQOjEsmfoJOhS0FGTWZJ5YPt1RVyQen+lBAS1poLdR9Izu+0P0gVPRfKPF3hsrH2whw/Pproyq1G
abcmGMfcp6Ittues4TbejhIHTl4kxDgF5i0lrgo1YXDrWAOdYJooYLdbr1xzYOzXs31CKNGzDJuf
peKe6Fk/2mxVJ3tp2//Zt2x+1FDmw0VbgiaUJyntsS7v7ZlcqpMnFXqBvxZFD+n0ifqCbPPZ3H5l
v+4rv95FNeNSbiZnAjpXqTQUM/5q/dUFf/TkRq1i6SCL/VedAhK1m0S1tUPH/ZgCP23NYOvMpJ5H
mZlw7R9jcmyrSBTjfHgZkM1tRoPF5XKzW1GLLmVFwQDzkUmMnZ7QbT4SIqoat20IF27Fu/Du1wCT
syEtoEewCDCDKdUzFZn0uR0gcq59HvCI4crSqeNss63frwvfuEdE9aoIARr71UcUBxacPL9V6dvY
YKx98CsEczLFPAlFguzO75KsaePAV1dbDjTp/u0DuWfj7Du6NLSaolRLwPvrb+ydaO6ARRP7SBqi
gcXtVYDIM/Kg2DJhPerWlmdG44hnH1l6skGyfyaWjbj1ixavs5kXg/DjHxNz7G38q5S5NsH4/C5t
D0emmpbeX9tuhFvL9kQNqOvWNP0mFMwLimaF8AHA+Z9XVKCQ9yb4OTaDdKkecJgKANwqDxgw9vA9
VlU5UB/R23nCy+OItY2jMOncsjVS45oO6kAAcirxjn07vMWIYrXB0zi3O806R31MfTXx3tSWrbmS
DKjNFvfAwf60Dnvz3B7u/ck68YXN9mwVPvXnL2Vg3a6IMZiAXqTLbtggGTNPIUPWc8YvHF+lyxJc
N2DwPwXtlVMj+tYbV4lJnO546QDL6jLBK+UJB48fC7ObNwXGouu0yX/yyC85YJs9utEG03iLnCui
KMZXxYtIsFEE/d9zf8X0peuimKsFc1A4X4iRVPe0qjIQZdAhttes1w6Xp7+9G8e4oLc7YyL+Wtmn
peTnwLGnmjpeLfVEvABE1KpAjINRq444RxMU+/cIG74QJCJgbWjMzp03LHiSWXsY+HJ1glKkrkof
SeRX2v+Rf2e+/7NvGzK6BmiYSD+GX05bST5SvEXOE/XjZq54B7PmolDCc2Zsy/7tHFTtw/98Fo6T
anfqIy1n4DMYbu9wS15uaAMWGMd34EwJLMpjsIslIGmqm3eMF1rEzT+yQp53f3j8W7EJIvzjsv5V
j+wNHB17HrAGLyoeTWVwsKDngnemIHtSul4eZix0n5JIplQvPjGNOBxQ/Tx0iSxwYL5yITURTlmu
DmXoB6lxiZGv5TLSMd8UsABjmtpnH4RIAO/O/8FPKBHsj8u6x26+q9AirLJdf5u4+D0+FYvW0S4w
4I4vpkMgcJ65w4EgQiEKbZvPStdRrfXbBYWLd9nCTl5jJj0HYJfHt/N23STnL8uICFgFO+iVLZxR
8poMNVOLEL8MFMdAEwucUC4bYugrs9ChUITviSg7llg5wYEo6dMhWu4rzUBp3V//psG0bXypYK3E
NWEfhlgi/F7dfBrBXVNwoj+MI9DWDv15CfIZzhuDqec464OThcNu68J360vQLkkL5aMkr2oYBVas
oq3iehsgxkKg4cT7vn1uLWFhrrRCd8QXw05UyI7PWJ3ATIonVVbbxI8/t9QNN15Cq2xkB/MP8iLc
VMiww56h5LU49dCrKNhHnFbXzgDBZGXAd9EJS0C7rIZLPNT6mDykIKHgDcGBCRvMQIg8ScDKRLxJ
i6vzJjdX0wpWI2KSvPm9UyvXwez+71cPBM8G/02mNHjCKj4HXQ6gT1NiD2dfwjkW/nMrke6SDML/
j8hf86WMgoiQTcllh8FmzJmTbQNC2ir/s/nidmNFz7ERNhE5RRB2MQqrb3MjkPi03iRVeznFLopo
mhSrDRhSwG5TN8AInmCnY8TYA3POqF7RielvWw9ch/wq3iZitk1EojF6czPbKKO0wgMP1/Km6LnE
ybUOH9XnPJosBsyKjNHQni7JRbQ2TLDfLSHCxAedgHY1QKhfYqoAjHRKEz+/P39C0cdGuLGUzYHa
VFtxbDGMwaaIJHp0SHkcPlyExFox+pHK1LdGA1TjbpoYwUol6WmeKwFR7y/mzwI514k7Q945La1X
FiWbPtbkuheAWDGw75Rn132YMZaS22eiofoRARqE4TEeZfvUa23cabz0N9/esTqzz9G3ISQTvpXw
PXmj3m9lyh7myo0CxlPVhV5PXLlns8Xf8qj/LT4KvN/pNOG5FaSEC2gah2n7Q8z0EK1CCkf49r12
LHt7nUu2NXcJzFsSIU+c1oMqiEWwsusIe74DqWhfwAV8eK+00X+P7jwUpJFVcj0G1dog0Erp76VP
Epb8geUjZNM/cICMc63Krdq3JB/pKIhXbF2fiIQ7Z84V5Ft65xRLr5s1PoRJqLcgFtinEyzb0rge
0OZD3UiX/5A7XKMz/FLHxRZ++dyzOx5aW6153xDXvrQIDODZ1MJSSGru5C011V7QWOyVBPuqBcB/
7TbFjYJfy7lFmV/ZWqLT5rmkO7UAV+v2PeXvqdixC09n7HTTz/9KPUhGKzVSNjLi77Y9aZc3QUKA
ITM2PeNEIcqn7OxQ3EVxksEc8+l/446wTqg0sVE8LB/2NXIVB1ZrQKqKcO24X/su5+2S1AbxvUz0
ox4r5CF/iJbvOaNXfvxZ6ShvUHQ6G5VaVgX/MVn1I55419EljXebt1kaoq9qFpo7MSni1i76n/91
0lXlKIxr4NGQdQWBKkOgz1Bv/JvZvQCoToeM1HtLSmPAeab3ehfUaiN3N7cnC8PDBiuKPes2ArJS
0ycpXD5XWNqkSKQLZWMtpB134b71iqmEaB0ZgEDO7qeY6go+W8d2Xn4H1BWIrxHAsSVpsOXa6tBz
9sNu/9YWZrU4U3uA5kPubFST0f79Hqd/HXkSRp83HQ0LhJGrQfs8calIDmHdh23SVJxbvjvDQg8L
vanLSoGCGM8NPzzJdokhulaFd4tZGK5dEhqEaGgaV6dvLgfxxK5MwkzAHn635FqvSFRi5YhK4YNs
ekpPuRPdrs+IQDuGJfeAMAqN/AbEgBIHT4q1nKyhvEeECizHNgC3kExUNjvLITDr3/vpnMAuFQm0
qcEb+A90nbNN1IJVgox79DFPGxCwmSBTO/UrFx5SNN/9SIq3UMHwcqvF6CqXwJyZQmfCDvrNm4/9
uSgwdGUr1bpwupRk7YWRZaoqqZsS+3a3s/29cRxsuT8G5VxOgWSVBAqw8mTsk8t7G7GNiJLr2f/j
fivCPRBc/5Tph12G4ebBRV+C97owzGCkmkIPzCclJXzCkfIhfDenswtrPVnbwcpTihOy9m+i8oPU
Sn3dgn/Miq+x204PnwL60ev6sf3c+2E14N1cbNf+pBs4lYWKzINmXoSbfWSxb3HuvLogW6GhrDEw
qnAvszFbZxvlZLxXSrrBVKKDXmc3gyDrOfT753iHt0ucoCUIj5vR5fBRmsuHdrvniO0gMEKLmraj
d7YJirDEiBqRAAzxGTM63wFBAYixK114gpQRrQCqGYjXzlDp2agS4BvxT7wyrvRKzHQHKRGWuHfF
I0sUqDucuDXtreENQOoplss8dAJ/JeafamxKKHKqsaT9CLSBmA60koZp04/kK/vLo/rwRenykd27
k7ulh6Rsu9cXh2buvFGuUVZdC/pUvV3UCHr0NAXRlJFjPA3gVsSl29BIAG8U0+T9tXkZvowqxwx8
WQBffGslu7HZ/+ZqG3oAm2g4nfTEpqjofvWlY+zgCfAorTgin8lxxk3tgC1Iby4buet1r1hfB4ee
97ZtVG/2LacUsvmZK6/AOYjBblYQLek/PfWVO4wp9M7VQ+qIRB/2Q0R7NfJXZjiRyXcO+yGOGm+7
IK1p8G5a3vLD0WYCONPDiwTFktu2E4m2cwZg96bLilMDNNo4X/29V2Y8MlFRFHqmimCVxo4S2yro
v6fW7VY6MkW4oy3jXGprRnb9U24/cz/gk2R7aAQbfY4kQ9fUz7yfX+BpN11bl+46ShHTYklT1Rhe
2DhZN3b1+pig4c6fkHcJQ7RZzfrwfxGjNo0bJ0lxbOcKW6kk0vHWz1Z5eHuz4/z7rFwkOZpQoUCX
BUKPXE1+IBcmClAtmxcbUmm+DkLiYHEd01pnOs1nq+9HjX2csmEuJoMRptV8f0Kguxmb7+1gf9TJ
JWGKHww3ZFvo+DNnpH0wHl5QVc3WVOs5QsLizeNrolMNmI6UYBNF14Z1MdPEhMn2KL5qEMxrUtc5
QD7JKxr3sgH8OM2/GwHvRnB678odPMZqFRBgLhNmbstdfj8BxY4/u1a7EYXzPuMgRD6r70pAv5KQ
c49CKKBgM/7iGACd9tu4KpmQ5eIh9kglPOhrbqpBMlqku4bqlOISYL9ZHHOoYRs2SaR1ldDyJtf8
OUFr2aPSF3TUArRYHweP/35Ik1tdjXE2oQzFhQV4bGLff4Os/TIxFk8Z6GJyq9sAyCAZJOAa27/r
6dcoio2D2c3txRrW7nxDoJT51xNvS8Y4KhB1dL9rwAYiUfzKjM6IYsXVKe+NCgP+e83E5VLZeazm
lA3Az9cxpzlQQxsknXPlyFI5CyK2tRbbqCJe3J66LA0OyMXsXobImhM0cGj1CrsxDi5apGVJDNQL
Oyu6ucHnCIeUCjJSEbvl7Z4iUssUqBH+Jt+7tWqXdv9MSgFjhGXgRmlsHS0iajb+RV5dVXNHh5Qq
t9+0oMsq/YuKC++ItXr75XKV1AXnGxSdpEC9Qt3F88zjSXRtHIs2sQF3+2R51iQ3pUgDwtpiKkoJ
UR49Xoon1mUBNRaDEkZDa9H6ELGzwIgS6G5VgZAiBug2F5dZg0nL48DNoZLi9qFC+fiiRnJdFiDl
hpr5GPhWUf+MY2CHlSxdp02OgwU69k//vAVGMejpJEBEefLGEgRW4wzTDUXgV7i5hCV6bhItMOIg
4E44OCMEGKujaK682ae05sdtd7OZhrKvHlouTnXQJF3tzgtk37e8f+Ipdb1VKYONCi4UGf5Z/uKZ
hBvM8FSXwXDhKMhVyWImWHgF+7DBnOZof+mYMECJW4KngsH3+g5MlItu/nU5uvwTCzRyCY/cOFTK
MeO/zShjhmYQkGW2Yp5h/vhpxGBYBqs4og/WbhwycOsj2VWehzGjEjwr1sVncZGwTn4em4sR/CBy
4WK1hq1qm8ubPzDs2pU/OHiTtbQKxDTQ9XbXMSbwNal3oUBwVtE2aIvjhBd8yxDtd/HWOrcegkAv
hfMDZbg21AV07YzqXcwXpTjYGYJrybesP3cJyvc2BxE1A++S6Ofm20dEm+KKNVIGmSECXlWWN+f5
dqAKtBaq4VUyeTEquNQoxNnl/WWkJ0I04co4pc+odey0swJdjFTIatt05NuCxFVQtSGE/5xdNBnj
YQLibl5nUKRMegrQUBfgj6veqkbZu3IkP7qM60gDvD8OGqrqPILSx7iXpLP7wlzQ7PDWg1jKHAxj
GWzss2bEs9hh7nKVphrTdnVu7q2pJEUZPD9nsmCt77/qTnmUDFZL6SJpTV/lF6MAAHp6tPzLw98n
kKa3lxSbsgMVD5DXik435LL60/cjGUOcp67T3sDK92Ar/tVtsX3O86N0nfBdx3e1Jjy9uV7wz43B
Im8w9rdsQHquBBw1YzF97NyVIttSKKtwOnJsWCttEXd0y+fOqpTeCUiR5lfhXWhlqa+t2DwtODvF
c8fv5eg51GWVUKK1+1F6lhq4ErkkPC9FevVqPynyfmO55idKhuqcAw6EXkUuezxVDBxBdCCpwVWi
/4R7xwRM0cbJC9cbDC8rEMfQWJ5ZrxGCePW7xzpsZrbymJawBk2oJzA9TPrc3+r+MK0XjhUcRThi
Ssm1hcdn+bWTOJl5bmKqIo05s5lG28KWGCcjmp4cL3hqY5PyXBpPahHAME1X8es5UJgObOoKRJAa
bRP6cZxLC3Ag5uS5NEfkZ/zg4slRN0K5kOHMUrTRrNiAgfPgOK3hHbccxjs2vrGPavNzawC44X/7
TehUXWxADZ5om07sJbclyH/jRcN68uRffW8JPMDh0hfFy5xtlUcaq4OTIbCUKpK62UZti1W2ta0b
ne0+wbzJqaz9C7pK6Iilp4dF0jeMdIOpzIpHrnXrczwpLo5w+LF3MZjudtoLkm8pxKiG5EupFlIk
KCl+U/R8P+lwY9W1i5muXJaWQ9f7zATPO0krkQ121A+IWN0hvE2AnEguJHEKfTFAxpEzPIWt3QZ3
g34ZgeeMeCLExh3Mn8heaB+uyIjxP6Q7vxG7yWnbmPO9vI9NTGKeHDsuCTqbjTbeiHoEx3M4Wru1
WSXzsvAMCnQTdvS1JpSmzpz+oloJjFGDeoAVzW9IVDyVWtv5CKw8foHuFB+QdbPGEAqk9N6J/Itf
pTb5ZG0DbisccaultdMT3PCWFEEKDPFoXcklweXQMXemuBD1R1JKShrmzr/GQ6tIKa4GUjeSOv0w
+OTtpD8g1Ou3GIaK2F6ztn4mJSalXADdWaIXcpwNRIuDOzyiA4XpMICZY7Y/UXz7M75J5xEKVFQ3
6ZTD4Mm7GXNDV/z5GPOjUOxaPjJ2NJEZ6LC/mf+5+F/TxImHGrw+fxooxOCcQyA+iQ1JdjgGEB6+
qg/cG6wfv+G91CYjdA+m452KIR7SNz4xL90W8dLK+J0ZueUzvB2e5HY4jyuXPBZMwllPNyPT1kOw
wUgVepiX75pBuPT7eqWyFdBV1jWTapNgRAQaMEPMEayewl03XzFPc9ScTLbmqQLzRG1VjHvAN7lx
W/GPTcgPFUtLOB0zYNigEDLMzyabp4LUXzog7X0nCoB1FnF3VrAhtoiydWIXmWdTD4qn5m48/TDi
n9GLf5anQlxW0yUGdLYfD28K4oRfoUahCQvDNbqBGS97LZEuLTIC/4Fd6/Eo3OSxvJvfqidVdjrl
D82LVGV2x9PEYJmPiI0xGpQq9GzlbE/dXFRTG5OA/YhTr1oFjhhwpiXjMgT9zMJ5EfZQpVWo3rOa
XRs9zHHBs3CTJpFGpqBBiBr+oD1eS8JBaFlejykxIBr4RL+AIY4Cm23ipZgaYW6ydlC7bKFKeyq/
0TF3nAT0EqNjd2qGaGVclLSEZ6VRb45SHYOxADY8HPXG5Mm6xbJauUdgA27DUoubtxUm1prW1G2q
M01dZREy3iGJP1+YIh+NrjEFUlob6fqDWoY4mYT9Xiulps1vQnZ7eycOomg+5xOaPZa06ZktdEbM
fAx+ZanQ4R13sJRyV8VH5AbeKcqdb3F7522l7dR43CVpCOBm8i+Nc7A1GuAKPYrznP3KhYUoe6ST
Hhqmagelm6gXQUPCFIas5ZeDGvSKh884a00KljARDcICI5k445u9w5D7EdqZt5gDimiU0XEC57N3
B47wZ9N+EFWlOPDMyu6A9HSr5DuXC7o1XzMPJtfS1jduIiaAECR+TeiYY6GPK3vf8qpKS73/ohRt
rObnGRnuOA4memliTsAwBZFB5cambYV5s0PLWV4qUbUz0H2FspBAA4BTHB+fDv8ySzaPLB0neDxS
PuciT2J7zviYNkz7qCdypnLDa6jyGlBMUc7Gitz4GTxScR3FsGFDeM9L66Lm2koQ4mxeumgx9Vk7
sDrnB9kXEDefM49M2TBBjLjp1gADk7NMEYOTisVXrgadfRdsB1GHIiXyzFJWC73VxhWEB0jbIVVD
KRnC5R3ibCpUlMJyvu8LgvkIzr6lXnJqJqMMkkY+jR9CpNmpq8fJdDq3/cNMUzmDNP5Ya3RASflV
25yHx2PKNhaIHmP7ZnfzyJAV4buo5SiediPl3y4mvyPmcWG1e+GXTlMNdtdh1c8oR4e9zao6ab25
W3KkntgGTDscGmm1U+HKFuah2ImA0VcdleOuT7NmiQ694a/VUxLp00sxNV5gzDAs68vuvMMFQKkT
yWneCgHOBcDOVRsTneLTccL9Kr0SIhIv6xtp24wi06G0XXFPCq7upsQRclxpuQj69/4mq31HRK+b
PE53qIlrc7I0NeQgkhF63ofiiwvPoavFm8tmkFNnlZB8DjEs3YYaBfJBa9zEuZq4Fn0aKb9uFpgW
qqDf7qwwLjDxolP7DoqGW+oCgHMOFoxoxwCh4rLQkKvO96+e+u+LWtlICdsJgyMm3gohKOJPxoIq
xl3yBeYZWiZmZQ4W3QEGpf7PMSYTRy3p7PNw1FpdHko9mdas5XzMUYGycp+DqQpr/memPIlcgV3J
E7Ud3ryRUhtvsZ67nHNw1PJekbCV4r+Z7UpOm+cMgf+3aJMd+LR3wS6w2MduU5FzssHHi7D+2L58
cPjDXJPqAv0okVHcI+tmgIAuXlUIupkL/u/OGQRQ03N0lNqQs027hkOrAAEEq2nKyHgu9bdzS79K
seHDc1xfrxCHpvAVZHkpeDrGTi3n3fUFhI+qi0SE8rwC7vteUDKQ8dR9+NB4evoP9JL4eccAAvVe
C/YPxFYYn7QEuSiVXlgYqweJgx/SW0jL+ekzfelri9I3LfDZnY8pyYHK8g0mPHdmnk4E4BDvOkiV
07Us6obK6kxQeYbDQG2XUMcnqQmAIZEWFUADawoSut/HhDzs3cWKY+GmEWRP2735tv4TE8INI2kU
Uyk9I6oBq/DAU3xXJl68xllMcTk4pRPnFiU5choxYmMy1LBIRxyZTNeGF4GP+aql/OpdhPVkQdf8
dF2E2fhIE8LJL6NS7A9Xdsfgl1wGirtCRzEzr1m9S5XcSMzDW/sNAx0ZKH+aONgBis2ahqly7Gzi
lM211kfa8CWhcEpljpkrPwR7kgkfYY56sH05hLclWlO1zX1VBZhUyKxZUGciL7RG9LEIQVesx2VJ
oW26gta6W0xjtUImlXUDzDs3b6xeyRlvZVIA/NdTH8FKI7jShYHEgktEJZBC21pNTheKNapeHBws
T0M5uCivBT8dx276n1luyzrGbU0mJRgrYFUm3+Fu+QjcPQMA45IhKndCvXkGdyoqa5BtG8m0P0Dz
gOUpieRv/4ZutPvnlwrGv4ihVwuktMLIiM2xuHOzZOKeToBbFY6Fpj6+/qOwifQqhaA+O9xaMABO
FO0X2uFQomX6KVPlUGZYEHtL6cxGl+5AHukZ7yA3f+8fyz3HZm2IHhKdIh1bFI2J1qRf7l4kdH3F
zeX6JCaQr++JXEpcWrp9VvGlKZXa9RTAPZnujMnj6u+w1bk9Vq/3idlgo8T/YRUEVis6E0XV5i8J
HFDwVZIgyHvBgtV8n97OJvIhRpGx2HN4kfJ+A7ReWbskRQ/m9Y3Jl80oiTo323J7JfpqT/bi/2zb
0nrSj1kuV2JMZvmP9sklHrsGAqmW561bBXS7I+RNj1aKK5T23wfdgBzxOBGUVbjUxVZZb3B5aLpR
zH+hO2GW8JoSprJjmLOwt9ZAv2djY3+tN8I9auINVP7xcprL7o42ClqFnjGmZj771kRbxQtFc5tR
OxNXNz7Xai0OI13+nJxqjtAQYrLiu6U8TJ3U473xnDVlKSsuHHDUv/ZqIoBlUeyt4yC3JttDaEHG
lL0IM7twMW6Xoi2h64CD/Ecq5onqm/8vQxfMt9jxRjNKj5hnS5DE4UNR4rComqs9BjU0/7ZcX6nv
LRFeYbYiuw7kgeDzu20s4NJWpikR86NJtuFhTWOJX7+mrHe9dqqTtD73jSO0Jx4CO3lH39wzHTby
0D2fKWZZixumCKiElEndG6Rl8umgwBUddQVYrNQeZDjzkmjNkCQr6+ztxASuIcYIsJMW/87+BWgl
q5cLl07U/LQs6lu7ube8OavMpK7CfdLYfvIhjNjtJXbf522gdEQUTPy8WKKykoQPWhqbjnNLJN6g
nu3125+URpX/ttd26mYyGI6B3WmEC2xXJImZepr5AbohJU5BZsGuUZsWlYBAMej3UjjW8KFLjHUm
F45TDKmxV+iePgSWE827yhcWe24uZVqKaFjh+EiQWh0fJgyrIP9aDTJmDfEiJEo6qjoxYNXrsR4K
WlXbGbE9DEx1YStJ6qKN6L4H39vggt8f/8FFvcrqvMYJl3974++a1RyQErs/x/DxfeX9df2OF9DW
CmlOL5E4H4X/Gatijsj3JWrHVZ6j/WA/r4sVJng7KYryrKzM/DqYo7DX1eVboMSm/tmBDiIeufnH
ZbVt1zfWy1AN736NMzvhbMm2ZF9GsidRyTvHrcSaeV272FRYMOXejQIi4r0SLRLd8xu5MY31fsRo
yOFYfqQRNvg/NHqlCXjTPfZC+lkjHC8804JAiKsan1CZ6TesLwYvpg3modbrPPNaMoVImMy9g3yY
DotZBcvoQNoI3Y6A11LDOWGiuWhDrpdYeKNUeHrH0Q3K190+Xty+9XfgOufwQKd4ogkjGHASbFET
VRAd4asYPscD+ypu110/VXbt9QYeGRFF5Sm0a8YCEs81YhNVZUfifrenDZlXccmOEGtxIuCUfmLU
ArrmqqaMxFimtuH/uyOMfzLW6q2hPmtUi/lkVu6AeIqVkBVu2Ui8tzs+30MlVmpbPpqgRoxMCqK4
93X1xCSzX3Ypiq931hcHYhT7mLsgLgHzUW3v6lBJEEENUe1PRCf0AND57uvThGT+jzNUXZ7+ZDAC
KButVb3YAn+uVx/LxCo/ml2akDNzEQK4STqIcdnRI02Rc1yNb1L7N4uyox6dFmw3eEDPWXWK816O
l9euqdhOLvSlHrEtPJDdTDhwaXEIL66l5+l211GnnGZNy26OOwQhPOAU8CnmQJRXgddqlfcJQGaw
irAesmQLsAOh8hzr+fg3YAh91O00oA50fPaWkU82K96PS1P0W4bASJcsgfcUjoUnKEuZNhMoMzxk
DPYSgfqocc1OuIwdrifZbZ4KHGu4kofd7reQSGoQIAvEEJrZRP2K90DduikTBXrXyJ1/8ODSgH7O
RLEd/kdFVU3jSU02kmGoUZKUjN3tK66eeFZLemgdIqkiDzU9hlxqJQEL8VZ4lsdgi7BdrVMORmEC
yTrsp0qOYJa9nLnX/KYCDyesRVCaWJQVq5J2N6A92Jvz70gmLU1AvP6phWbSqsorirdy7mvxe/Ma
JcQm0dGyZhmd7u3gbnVEhNrYfIW7zXGGgRAsra0UptfqjbSBskD/lRd1cwve7PQllWygLYiGlRik
gSsLmlrX/jFes3DqDZlgTINc+RYf4OX97SsnHkdLDWROJ/pDyWiBH/GV8N/58EU86rHK7Wvoj2j0
BjH/dn2oI0fXtziRlk7GX26nV04TsjuN4Sib3GTQwAHEelhn0boSjzO96+3kTjcz/hvDTvqXsJSI
cCBBRYQaIhpyjuliIVdR9Bv3Ukdzz/gO2Q39Dao2+DNNTi/CN/7MoNtIkBWWFOUN4xCsFUbthbwb
MAaKHd/bQHSBxEUZ+q8WCEz3+FC14y1P5EloDM4chtBxwiTuQ4PgkGb8yApsfSfjafsrJ10fUw3U
vye7hKqlzLkSPAgfvKagYw1cLOOkCjZSnhCLAAI+I7fRy5o0N9cakE071Z7a795gxi++BvW1NJG9
3zPA4fGPHNJ3HGiEsl0ZGiLGxLOao5Tbdl/NHsdn6308kj+UA7dZ9nXlMRR8niDw52aykI3JUt4x
iBjjw8icLf5CIMjifIv7zEPUlbcQN/FDoksAxOnZWxUEn7Audr84h9IgtSHccKjQU0VVlfNWwj2K
TS9zOF19YL1tobiN2Ln8c/T5xE4srHjtqAWhgfyvGVwPQAuF4Bt/uZYzz8E+8AwcucnSYDBephji
j/FA7xh+qfug4L5d5zlwn5PppZ3TBdkTuaDPsyyFe1fiUTAm2ePuMVPp3aN74HWpgZdxaGVHUVur
qQXq7D8CBWo0RhkXRD8wT3+35xYg93AE8RMCCYnRmxnBBUCxRyoJ5+TgJrGzIrsLOrQqUYR52eyu
Ju08XiZ8CK0Exp9/CM9nkXIxWSVzOSqlCVKsNbPPCjhuP1YqA8+pO1pbj33hYQV3KeZNKVskz3X8
teDwjcZUXZaCRsQ71iP0dev9Jmm1osb+T+AEkTa+7ajXWO84NOtCZg0ji0UOabfK2cCw9UPY39YA
DXf3TfGG/xSOfGSQK3jE9/JSSRb8QjH/OjFPtaK2DCvOo3cWitOJzxZe8CdvfE6ZfRx8+3Q/4EYt
35om3HRiZDNDr809NaksSZ9sAgnSGt2sWKwAAANEHB60gWFzPz3v9RcJe3wmBr8oHClBAsxkdWTC
DIGQw06GJdOzsbw+Va/vWP+XHAHDRSpo0AmAv5mxU95PGeuEvT2BhCxW8EV8h5JUV1AGr/n/snnQ
yr5w3//84wADhEDt/U03VNxNJWuTFzZnREe63tZqKTtMgTehCVngtoWqOVywlXt2d3tgoeiLYx2M
tUZMeBYusdzIc2uZ+t6agfyEP2ogAEB12lrgTyGYXQ3/Qe6m+xgTpfYJ3wlcZmq8JjkKHXsr2Nqr
rwcHru7AeeczopRIK1yogAjV8jk7W/4t4CI6OL8VKJxkVGIK57W1OY98BOdgAWTmVDQd2YyicDzy
HgjxnKwNTDyZzNURlAqFyC+NV6HoA1bNGbalVBXaZKayJiPRjqOBtLCJ11mdhPqwyGIebrwl6KBB
4is1NRGtH/xyu1Efpni/n3KAqBVUEcjJN9BwrBSJ0opKfXwVIRm4jJwjAFVjB6b2TAlZwnn07CsC
hzZc9f2ZSDICG8yp0LFQBzrXb76fZ4we0hXtaujF0yQ6S4RIwu6DmV+flEcLbUb+V7qPRtZ64/O6
KH2z7a8xck0CaojTQH0Hq3wSnWtSuDWkMwNP3LVWom2ZMBoYXfudh3csP+HaOStrpUnRuljroFjX
oibU/wKJKai8X3hlhLLbXSAp3vrfIJAXidF8v3x3c39vc4k44V2L6DL2uYOtJe8T000Ulmfq1vz2
AolktkM7laYhQX8cxl9E3tp5qbicR7jzDbduDkOen7SiM5a+sjvX+iTBADpwrhss2oQAOLV7V3EH
/WncUmUzlNhRWW+Z7dmSpTVF0T1pAvyWPKaggU03/7uvIl5mEhMKtSymDkeB/4ekn4CHm4EHYgSx
y/gH2JLEGNCuvcBLx10w4roUWIbi0wymVTSu5XGMjVTW9wmrUxehVpydgHRqvI3fGU63svpTOY33
XwUn8pLnYvh5dszGy0B2maqt9/dahKAgLgiwHiu54avvftyLgf4fBdvodLPKtk+IhDuvm7nwMBGZ
YaUVMJ/TK84CYfe/YOHohtI1kzOrl8dnasahCWKOTv7zyw8GG+qNW4fM2ER58WmWkBsApIOkwvul
0XrgWyvmPa7oCb3sU0B5Nj7qrOKwlP0gsy1Lvmjw6vhFViw1fAB/Z1Kwm+BY+Iw96y/NQXTNsb1r
7qpM9mTZIixMl35nWIUhmhyU4NxD9u5+rS/h1aD8izh4ipIm+L91VufCQyufUt0rWMjlmapp7qnB
LxIkY8KrZU+C7X/NLYvsFQNu1EtMPVwVf4RPOByC4DTpeB1/7vn9rDSx8s1VpGtQOM91bztJ+USz
pggJ7wq+4eqHtrn7EIM8JP4rJquiHd3jvUxSjatT/Bl/a8XIaoH5Ouqo5SZtHWQiU1KmEOZpSJFO
F3YLVMrc5c+Yhc1SjNDH/0cmuGWBprYWUwpFOkE6j6q6WwidNjgEvradAeuWJitciTVGHOPxjcaB
GRjQxjufni76TUVdvnfOrHMjHtFSpIXClPA8E59If/vOaVcs6W3h+EUpUBV11s3xGfue0wNwPA6U
nLMTYA18A/7FocMtI5NPD5PSUDA20dWECt7RxLr2mqkWxsqrednljwDT07kZWzivAXu/qtt8Hj2U
ZlU3dZvnznm15GaMolwpCGmX3s1Zl54yV1re3HWf70gmWtw9O/zx92BVNFvd0qvJYfjdl85PufRD
XOiqe8iA7PuaX7t6/XLPMyTOxIupWBQByxzZ/sfLKliSB1253BFVlGZ4VSQMyoOc6BDTp67ET1bD
IbtjbIYE3NjTrFy7tjhricOCsHE3lbdw8PB1ytVCa8a4uoMEjFiMn+Qkp8buSS6yMJdZz2ymOv/0
4adfncx0nEQjms5AUks3Lf0F8I5VskHmySlNSk5VIJQ1uBPjKPpeKipvqvKYitIXPpNVFcRf9+ZK
7Yb4tWVm+xsQEg+fJQDuyaAEvmEIai4QtD+wQAh0GUR2YjT1sc5+nTllSIa8+uQKQvko9Q0v7S4K
vS6NSR+T1gR/0jyips43ZUNrJASLyMRJDo4AkQYk7L32JIfMaR03hGRzkYvDPY7eg+6cbmkFwddl
M484f/iOlF9blCo1sfedcMbwcrtEGXY/AMRl92vBaTYVgl1wUcNrHnffkE/iNAaczgJKqnBoaomJ
S/4U9IW1mFhQq4KYTwB/WF2bnfgwE8jPDeD2o+/dmi86AKc8rSqFc/hTooRNYok5t3cq2koO0FlZ
LIjcEncSwjIppBFiH3581NfYDp9brg6V+Id7s2380xIzhNK67AlCq2RVQ1DV1thxTv/H9SryaG5W
PVy7ZBUzv+kUECQ63uiyhO/ihyJxSq0ejS2c5n02cvB0Oi0ncCOj/2gK4+4VHqo7MBwoaKCGX53L
XKCQnRmRdP1rXMYtzfVjmOBD3ooo3BxoZdOruE5G324kgW96CJLCF3oDCyuB90CFsf+JF/uq+aig
xo4JzqWLP8tChaA282I78VthTiKHdUem7Kw7tibhy0oBe0tnxNh7SDAgOUzhDTHiAmjm/kvP+Fq5
596j/yZ3rw++73GTPpuv5t8ztrszL0NB2KjqAhIFsIaMapLvd/Yx7VLgmUwZtiVAORRvc8w/EY0c
NGDDcxVwTVZOvFAl8X70V0u9gMZu7rinXEv5p8AO4s+cImgCN+k+EzckOoUDjz5etE0znriEPRkB
L4aoZZukwKQ921JC3XdK8BYEbFoMgp891C4sE0Ndnyri7spGgF2HHH8P3SRBufziSEBUpKjgF9ck
JqF+TIeS5HD9ar3NwRRxmqPP3zBH0Z//wM2U74lV+XINrVZPJYMBA8Ik4E4yYIvfjSAhw9NZObSy
hJ8+omma53tww6uRNnNxjhSeJ6tCKPNcbGpl2vFo+Sl6OU+xSRdW+R5o67GIR50m9y4RyTP/xu3s
1oapPDhVWeRPEDoTK8CkjQjdb45ypUHaDRaWqOilRwmyvu3kGTBuCvMBH8kPqKeahoerclJQife3
GFjOWM9AkzmVlOVmW2ItNry3rvijuEqzjlmgXp+2wgQsqzV5oN2V0x54wrrsFZEQ7X3UpimReSAb
Ml0G0Tzp5dKPWBQJhVL7gMI/o/QB4Jf9t8EF5sjen2OjgQDB7ZMJpM12HCaG4FeK7UHumgmmkfO4
UuRPmisNRzjZpkINKr1BIvb4yQxEsU2hLoFlV4BlWnhTdGBBzTxTxdznAX83rP275qTEueVJEcIf
mauYKbWQERyrfPhsIYOPOm1cofd6Se7DozEc4OI+HYeydxahGkvDU6JF2+q6Qo1dMgmi81DPDxHU
6VMITMgXg7MpMbMJMPf3EbJvODeEDzVpPffuK+MubFrlJvRSgrRoNFoih7xlXvuejT809qXRl1F7
YbKnB+wSdl7I6EyXd/8Y5UvnKBqgMrCLN20GQnPPKIEJaGQdiFHr5NnQuDGeIaKD7TMtmhTggZ3s
36hgKtNmbCek9vmczsWrx+4njMScbImZo2Zh/hcSfoGs/L1GceiF7uW7uoCtbJmzsxl/HIQygQW9
CECrBBZWC7yua9ZgaM2dYu//TCHOZ531seyjY9mSjg+1nrhGXeuXBdFmHmc7RmbgxAPswaWJRjcb
NGfiL2l3tQwdyxNVGHdAkpq4PZ/n/rqt98/lvXip0reI9KntK0JgpWks9uV/QMtOqSTtYmzhgK/A
HrYxgpaUp+3YX9MnS3gbaSxgsqFsFQ0qUwG0r85E1IEZI492AvU+2gvrUS7R82kMoep0cNFzZlvZ
0seOa/jsmYPTeIZtZnEckyYJ5a4okRU402Xa3ZMZYDTwlMGxduHw9mmGh1gKV3c0Zl1E9E1aZ9lG
y3nQeBAyeHpNwKqXj0hEiCxArOz99lRHZMFRqdfcTDtq+NJKgS7GxMADfhPuTjnePbpRYSApCnnl
+3EiNAAQHdDQJqF4zSM2YUC2fejehGiy7Z+cJppFzbKUVJxx4zahNhv1C2SJjBm+lEDRflkZKfOp
SjU5bP7kITbOK/ZlNopwsKuBDDP289mJ2LMWuj2BWyaqKf7vH+ZenhUpxcwlszwWta4Pl5UViWLh
ARwYS9Y2YdmpS/6hvaLmuDrD7I5dSyG2BHdfbn6zxrQXC1vr0ZC5PR9dawC7TJZAvHtZ3l34PSTi
D7zSwwVtOBaYBqleZ5wbAa2CJxo4z5mIlI4yiO6NJWesqbHyIRivWjQNzbeiOl1I7HXbzb3/aYrl
yOK58G3MaNAWf6g0/KA+eYeEL3643wPjjUAm1HcrUT2rbdNPGkBDhWvcXH4TbMz39KLxGfXYrkJI
vFpHlYho3hjJbpynPNi3T+poXSo5kDB8dprVWH8fNMFwiqm5xc9BO42WpU/T1laA9gbqVmpwoyUo
yh2GubHHq7nZ3EzAWZ5FeUPlrkjqqpB0tX/nN4Zvu4A2lTJC+E1tEl97d+4bnVc/VV/nMwJo2fw5
sd1DUcMhwX78X4XMtM8ixWQpJYJrug0GSTjpsDk/Vc1NV4dgY79+KkDnJOkVJf0ZJrNvHQ4aVxds
rPACnL+Qk2OH318w43DOKQHXHC9DkQKcHsFNbBg0dvdP7PitDttznuDjA714rKWyuBTWaNcCsubY
vBH9ZdM8qSDIhKls7jGJG0KJPUwsEsYoJmQWfoDz4z1GR26ESKjPmQl6AquzkjCb35x1Ww9+kWHD
bci6VkbbFneIi/Sjxr+Yx3WLK1Fv2c8VfwNXFKDATI2+TPrsrbbI+3lu5fH4VPIucbj3EHK7qTtm
mdSkr4+JHWVCVUsyaRfHwhxKuH4mqfqpy/C1gLJRpzDpEdarOU5lCvee91dCHFnJlDmpaLjv9pPA
t7rr87w517IlKn8pElUPYHNhenwBgjUDMYdxwGKzFCFDRqU7F13QS++zP2G1ABnWyweyYT25u3re
1M6w6oa9VdD4XFce6SMsZvjz5/jlbYDMsD6RWT8BRxDiQkyyaqL+rWWKraDV+PMfWkuk/0z7pem7
UzIeluRxAG4fzvlbgdEIqrNAXNXOXs0N7ZYHqSRw9h4JeipjiZ11pmzq/whjPS2XYNGnLtHpEmIb
Dx6HGjRMnkRsW3ZpO5FH2JsSr1p4VK8+Y5zsvypVBZYBd0RASte6LRbielULDxJ9wmDg19wyXkgU
UZ2l7n27GOlPsKumtk7RHyNc/W10o6d5cKKHeqa6N8/Rz9K4vhramU0i+OF/ZSayqpgx1R9W8yeq
t80BXD9FHpVQaNPXY9sQ29feCbCPuxlXOUA0U6zo/FynNnVemgkstKEPIBjOcHngY9MG2mHYHVSL
Og+ZOmsF5U34BD0c2CajibNd0YemdfAeprdyKUo25DcjzEEFDBqWQjt34otb7EwMb+j1PBl8wlD5
1PIfsuGbhT0bzg3edyrEz6zMyZ89rpTHmpsea4Tj8cjNXxicpsgjRmntfm38y7xeFiATw5zOpkKg
YUDcwuHfvC53eBBxCB5GCGnQ7P8iPOFzEA7bJ4eFxtUkES6Er3nOIaqEPFC0QyxkuHiNuN8qYZ8+
2o2a4XYBtiJXa3AlMfhTE4qo6/Cx15rj63J0EERbdg3A1YQJt7+9ix52hZRrK+fBAsxPfQY9Zrxy
94/dZ0GoSiY2uy5ZvhyloOHo3AY78VqcfnMMXopP7aMkE4UZomPBWggcE+jdEsgOImm9zUKsAnVG
CuU1W35bvwhWVWQwDE20C3tLOS9V6lPCWmZUNmTc9PFw4xSYYTTJI7lNNHFHtttxJA7bzDgz7QRk
MScG4VtULqR7Yyex+eesYjxTP2r/VpVu1vew5co1DqKRVjgsKXCigW27kEh4h00NMdnL8JuCo7pB
J/2vHegvsRUUeoxX0CCZ3te/TSFBbvN96NP5Ls1ozdWkex+pwjQ2xKhubdRwd8oZLxoFghTWw482
weZCo/a1bQAwnBDz+fO48Zw9KKlgtj/4xNBcd1SqMhowPhpZPjxkxEuBSGYTdHWkGPgjO/ftJ+CG
jO4xKWJtj2rnLs7kb/T5BYy5g6JwGBwcBDa1uFR+o/3zI4r2TydKmGBYs9AO+8t3zzAr1C0+gYZF
PNFSSc0js6GI+NdyHm6lDD1RmXxuAojhwvVrmRdjeZdhZYKYR4xHrMRZnSz0U7ZtUeVNoMSpb9mj
e2CpR4tD+VZa2xnYGL3SP98F9UyhgUskq1g2beNB1j+MHv0FEsXcgG5CBjZ3b2UZPHoWAUcGziUP
MnXVg1PfUYPsh0OE1af8oDsD/eDoi7M38nuY8RnIxaK/0qg1n6JzLSxttIzvu6N8vP3N0af7eav+
7UmBSI2KP0j/YiusieWnx9h63R9ljh5WdmdjQDlZL+fP9gEtq78RakyyaTQICoDNjCUD0KgKdnTp
JZ3n43JFFp5qqLBHumNHChrMEd2LcBCF3TdVN4MhgJRLVjUuBwrbuT3w2H+lKFu84xQy2Fk5Tncd
MojAKMzKi8E/5XF5KevUVW7IxAlz+SFS58ASqWZ4vHtsjEUvtKNvR5xVGb/eCVLQQ36wa0KNedoh
5RlvFSbS8Lw8zwIIaVWUzSNdUscnavBWpgZoskNvSZsvnn98lb4O97Yc3895rZCHAXDBVIyTPdSJ
1AJCfHM669zfWVDtOyGMYNWMt6tn1h946DGQ/buetJs4SO/8nFVJ8GTk9Z5A5B9qbEabUc5hhTMM
iyF+dclEFswXNE3VlEfI0o620inwT8Niy/yjmOGgGQYdItte31Plga49+uJQdDW24R0FBfzSdK+L
OcFvCDzlxitVPRjU7j6c8Aqk1iOJq1Ja422o4YdcuVac5jQbfc6IG+kXsGXsTDWQnncfnBxvsA3C
H7hjZkxLJ1ec0VyuHHfTw7Oslq9YKW3u4VsDPr15S1uxWN6ZPBtEGm153XvfVLkS9fvoVx0kJzpr
ge/aYWfUDUmYrZ41y9//E9ISJGPeTov7kKa7mHo7a/oaTdJbaE2CBt10hiBHwHK2dl6JdJ+zJPfX
dk53d3ktUxUL6l+wSWlyAXNf3UHJzKHqlBxwNeTYpniKKx+FIuDTglrFo6kKO3sKPb61YCyyGPfy
ug4NlgC5l4iHFsR09YA01D+A+xbzRxQjr0nCwSl6UZqk8yrC9+e1q8+jjjv32h9ZXcU+lI40jBrt
u5huya9BBjyVn5HI+VRDmdEG9f6wnIF9dJ5pizs0m6T2GxNwr+JJLgE4bmEusre1B65A5eOsnQGt
rXrtBxCpPGP727yEhakDLjLSWxo3oqlNIhBG+AeiKVqnBog6A6rucJNdWPliD9HbSD1jNDf2fqfv
nyifAGiUiGmIMbigweU5jDUBYzoGEdSQixDVFMRx4rV9/HvTxJarrdd2FlXrS5l4ziuUDq/MfrCs
0xMIvfNfNH6WDFHV5At6B9JNVGFblCAhYngt9PIgCgx15DOWgsxPf/DcNeHBYmOSDl2aCQ6vb4s0
v2rp/+omD0KHq2OMoGg/DCJrx5NEputTTulOCgKeVQ5gX3V2DBM2Ex9BSAFRfp0xFyCtFObi7zZ8
VxD9LJ7O5W7am+NBjbkQcp26XeKq2FcVdzW3+9SONaOljJnfZ+g1tDhJ5KdJEzgVWKy2q5ote1aP
eX0+D31h6ZfGdfkD0p5FiqvSH1jqN1WFjlbHTej6Ycsu++9E78kXQ4h4EJgg6CCuuDNehLpFHOHW
5YlcyeGTAzQ5Eb/mwhnpPgxCa38MrReaOx34nHVIEn2pX+OliOuh/FNRppPJYLN/RbmYIXNq0ouG
+MvPH0TuzdWxtS4m75hII3m3OpiPFdOEk+zjyIAC86osiHbLc2HlYnubu/eMMTJUovQ1vMiAwxkg
Y+7zTahwz59CPOxLDTvEzZ5mRm1q3LVJ2P0Ad60HS5yH6jxG5BGxuGk7rwmJJpPoCTyNSUpfEJt+
z8LbTKhA7CaT1KS6ptSNQiWtxIXhrd2bTWkuPgNCWQV0/bYRXrX1eqZwhhLS8brGI6GPvuu1UaYa
CGt/60GiOqen5AiCqALrexWicrgXbacelZKqDRsuDs6K37ImJgqbnt6Yzh+ton5MITEqcO0JIiVP
SCm/Yv07MZ0k0DV+/02sJj3c50FB+hefucJ1d222tHYOmY7kPZBD5RZb9cKGFJO5D2OTd82FwKQJ
d+QqeX5jKFXeQt0MSu4S+FsUgiq5Tpp361nI8nxR6qrYSaRD3MvCrnMEEqF146eHR6c5sA/o6AK7
y/5Md3Mzkt0cZmx4Vq3raDB7PmZZIRZUiT/IlpOe4S9xHL7HdM0M7OrGTj/mEwe+Q/9pFpHv8UWp
2iW6Odg/poQTojebuTRhJ2teX64Oo9LhtvQOruFCj6RoQIDkePjI0TsWs3jxNfI1vgR8nPvPbqZb
dhGMTYknH7QsL2Bhpu3t0eKB0yc7xf9CRWNw1K522Av0eRmzjABoo2fxyD9Qi8G6lFGoHsInnByC
RjUO6yvkOjk5Z1LZyF5MRQh9jpHHiZXi25v/U4Fh0zBnny5aOFKBlFcSQh4NTlUstTzYJKewAFlK
V0AqwP0+Hs90GvqMlAIGEnYEt/zDLvnI2/WHiwsobfRPhQEfxukCK23ZpaMglXSQ4cAKvy1o85R2
Goja71fTm7V2tw0nu2itAeT3rwGcnl3eGkwqtIWkgRxxHpFUdZqi4JsliRCuh16ux+3vbeOarH4l
dHhx2MB+Is8lGZeP/JQ44sq0ccfVF/A0Ul3g9zr71aUzoWZpRxxfJ9vSvfhHjhyfAnXeM7tP/9BD
9JAt50QBkIUrcOLRpfdtMggdqsz5GPsnKR5dBMWIrbT9JuHpi9pZPYrwxiu9PMVhODBr1pV4b69r
oDR6jBW8OqT8sSycnbvobxzKMdF5jv2z5Z9y9RG1WoDtcTpNlD4R2PHGh+KWJ0uNWCCdawL3vkiu
hUcSjgGQDlPyYmFqtfRycJOQ5g8ZPTLgLJHpToVuRlR3tUUesrS4DilLOg67BH5eHiTqVzn9RD5T
KVEfZH6qy/IXhuqGYAFnQ/Gyvl7TpjhFIxOUJkiBxGeWPrC+zPDRvVJuKtMYwswUm30la5YqdQW0
Wt1Nr9WdTzlprTBZJplcgfpGHNF0OpjoDjCgLfhSpI6r8HKU7ZpyaVh0D3nOLVo5g3uLJCrIXWwN
7N59DRIpd0KP4Y7zIdPJWCqdCQz8wmpYLiCJYuWXpolfdOloalI2+hQzw2HI0incEjPJQnKO1YJc
hIudwAIfySR4oQ6xwC+M3IP8NJZ83U0F4VGOWnFdn+vvjofA2Ijk/SWGUiuFfk3kLxMiUG3sbTR3
qpgZDQRl6lCY5GiLEQi0m4Mr0LpJ5buz0Ux8t43TPwqZRysCjw9P+R8hQVck8KhngEEibDaAI0BQ
qaSbltWWywNqDdHX8xUfIQGNLGQKnTVtgf4g5Jtic51eL0Yaxk05bn7eE9nVOWr6xJ7j9FQzvWlG
O45yL5Y4RReDWMmyZMyLIVQSHKrb16zutlZpTiHcfdbKDQAt/elw7cgA/bo38qe44a7lwiU4r3bJ
P62JzOCSKfPI7/fJC0wXPrsBhBIIPyWfB8QtoSZ2NYqeSRyHL3viilYLdmwIvqKgnBtPX6T30uB/
0xez4jWFnzRIr86Wl5adnLtgu9lK5Q1F83Lz4e7L06YwJIIZLuMQtKzNngFYTl8JMv6bf73kxnKV
IVR8Td3PcEYuAGaM2Id15XDEvq1/OkmtpsQuIJoWXhFE0yAZKK1z5ak3n+KLzcytm5DtsxMPB376
TNMfWZJY8HwCk++gwgPBVHI7pKy7q6UCSo1dOxG3Ch4D8QV71AKKcglR2RPHazkizELGAU/sJn4C
dVoyeTvS0rXUeX07TC3ZDSseZry9XxojSkEzaF6G0OTh0JuFYVEyjbvlX86zRHgEYEgbdFZsX9jD
xfeEjL8U/CGWU+/n5EJYVfILvcZoxGjYOkr7Mn026gl302F0DLln9xtrOKFaqXAq1THduhnMAg1p
XUxssAdVl08TRVVJE5ljIEZjZUDQN2FdE08kQtv4NfclDHDGhcYrWhTZ8oAoGuAAhZbQf8xROd6v
ZEj1TGY1SxdxuUzFxr3tpE1hYsy2TP02WE0RhT5KfDLo5cwnbMRcH9x5OQpONMbzwxLMxZuSWxjA
krYU8b1j4IayOSrSML/yKTXShv42w5vysory8DnsR81igi6fTdCzrquqTDTa0mj1aBMpDW2Sk/lK
ydMdqRpwBvLrlpAoyXL44CpvtFGcOuJSsBM53vvtjpzenFd4vHPK66BD9EunOfr89z6iSxFsA912
X9xl8X0ef0eWb6leb+9nZF+RybLU0fZEykfW2ldyL/wlqV7o7QtWIZupIZL9Ynx9XGM0A7Gl+7hw
2lY+NmUyddPAg71dyggzljfEh+ZrkrDlu54J/TsxV1QPAJ7JuO8Zm3CMcNTXTFQU3+Wu66xvi523
MIoI71VbqGhBCli7qcFP5hgcmuu5peHsVFJLSrzglD/A95y6Orcpa1HFoFrp5gzF2vYSE6ilK94p
CmKB+OAMnr34IUO6n2mgovjp5J4VmJ5RJMlxc5XPoIph3tGdDCow6MOpnqZ15p7Q8dCChnlp3R1f
RM2QgmuatIVv/twcEbmfg/rpgpkx27O4Z7B42pDBtffxPVUXNxG7Abdi6UTwPhcc6wl5inizd4Mq
/ML38279ZXL3veFVhL4z19EMT8g//gI+WNg9wyw8Y7HZnqgVeiCn7hcYW2z6reEcSD+QHrqJIT6W
+hfJlYaKOfnyzcg4OyybD9FZN8+Li5JSYzER6IiefiCfSD4WogcOxP7axmh0A6C6KiRlL+D6HKsu
A4He12ITordYa08j4PZ4NaGn3ueoAtZQpmAa594ZU75BBcmbIv46zIwE8FAa91IA82ztGxMXj+Eo
Bqayhelf+BQEVMp8BT4XPEU/SzXv55ygihVUymvdf9uedzv8HTuGXiEbqyWkavFbXrl70QM37+N2
hEFeLOeQ2Ov/wgA8iyHlhkqMFsmoxTvw3wyn5xCy1DqkMP0GC0mlTUlwvwevqaufSWvAiC8dkjay
O7hMCi+r/vG/3ffygHnEQ1wss+H2Lst10bszaFO9t2e46zGQQvk+oIIHoP8ghkbe7SixoTYFOmRA
Wo1PPNa21qHItlkLXy0UtT1ptmTggJ5mMmGHHe6GeTaz+PVYQvti8G1Wkgxn8+K14HUOLtpjmaSL
BXIGBHfsneZb624STUFv4HmSGBddoKs5sEyvIuR0qS1lHQX67/hIKJc2IF7V5W3Wp0insD2gGJDl
9ASBYYQXV+se4vSXEbJolOPBXGDecgCcsKphy3II3wXRKMStyJIHmTEzFJ+vC4J/8iyP/cIT90DZ
db76pBW6rto3R5JbTisYj/ysTzJs11f4bRg9YPj8Fpg/uTx+AWyPv3i2OP2UBrON6w4BDnfneeP7
esD4olGAsiJO7yYePoYf88Ti5OUO9sE04++7VhB59we2BD231y7EWMH4CWYHp1XWJKbbNHQZnHUH
j23q5kO1QpgpUXo7wd9ykhf3UW2n/H9CUA6nQaLrgiptYtglwz8/SrYs99V9dhUz7b172u51w1L1
GQhX/C39C9Fd9YsX39xp47QNEQlsgnsSHhT1Ii+HnBJQ2Pc6PotvxKQwWjD93nel2UspRvEyfTn6
fkZTBX31AHoxFSOREjyO78+3nsP2LLaqu7a9C1celpvJ45kpb67pJ41H3a2zhGHIH/Lk/w0N20Dy
HcIqDib9vCcdKQUcTPf1IbCw+Hkd94j7wIyDUMNkSOIqja6DfK/yMMIAnv93O0S2pupRhJdCSH/9
yxtVuSLwHi0iEiIAvMq64/jAzrJBW3D4H+xjwTQqfkP8OA0xeIeUWLL7IxyV55KccNs7ic4LXo2I
cL3j1Mr4RawysMKCe7C+Rgl5lAshR6b/bf1MEqKcBc6Sw2j5+wyT8eM8D1ep1ie4bqXahcQ9Vxli
gk09r4+OVn3ZMinopvnWPLtpBw0jlVK6nDIm9E+0Iwl6T3cogoYeLqbpuHYilyIfRnrZCb2Nat/i
XqFGr7p5ZqD0hPs4KoBChOu7dOoUACdqmCUq9qXp+YcXKrI3L34j4fxiQwCu/4qboud5l64amR3v
8IE6Ue6O3snJ8y21KvlRTHRITnTwMjwrtEk9bOrfHAIsWLYVF8b8dHpQ/rNWHBfaEBr3oU9k3//D
idI1g4RPumPfk8EcdEuqxYDv3/hY96C6xCfclsiPIjIivM1pY4gyDyUKTNJb7/tyjZN9uLHfckyA
eWTVhJMVrR3NewyN19kX84IGXMIrkPEGx94pG3UsHag8GeKU8H0NHFcWoL0lOn4RpLMhdQuEG03E
QCyPyxsYrrjf2rChzZeRShiD9reduiEaYXoQEt84z2VVNwGb2cQYC62+efqvdEHbMCEOhcKNVAs/
hZKCUeovYVMnnRkpiiDU10PlCC4wJx9KifsOU6TBw6lKDAcoXbYv3tRubhKherOiK9WFaM/CEC3j
mTilKHYvdggJZrcDYxUyORR918i90ShYprjNwCWQqT4Eo5NLnq7M1UEsZfcCF8OkWEV7ohglcL1L
tCXc3Wqx88fattE+yeZUQkqwJheN6eEMj8riZ5bnxQjEUq0oqzcNyfQuNpMAdkBHXGlzqlBcGqWa
zvDVZnb9c/4QjFb5oWD0DLQK7PvBMWADLKx6AoR5aZSamxkPUqOlYU9yjLq+z5GDtz8kZPhSnx4x
vOHXKXDqQAtMOMND2A9KojWCK9vk/eRokTNKHTUpEtRc/CxDFx5tl9nDewqP1j3NQ/3EAtuDfTBR
KOwMnX/1o/ovEKP+Duxl008vogvcOqff5TVzRFqw1foOmi/OyGRp6wOU3SISF2WwMXXOkx6jyMeI
NQjLVL15hlbHv9jJzEXWVkyuQFBjF8cBcSCTUeJsHB/SOnY90K9nWu1h4MUUQpesAlJvzQ3SAKw+
ICHC+FlbX7BA4MjHqPXKSu2y9JD0dUI/60Uju6dYV8UzSpkfa2GK5tK14jA8TwB66MGalfs69Vhr
wo5x1yhrsGKofiyT9iqycX2ugPaL7jqbH33/PiO1DoJZtIHwkB+XHJCPneOq+x7QylrrQHFsq3lw
avNHAjIZjwuirGsYlsunXN/cAAXzWZcAD8tuEIaQVMFrImzpMS/X//v/CjMzIIRgx4BHbDpM05UB
OAhh4L9qKwQnAE6JVFJu10omF9tyKufdVVP+fa8uC/yWAsUHhp+JJmTZVPl+OuuPyv/7ACiRlISD
1cLpKvXBv81oxaAj9IaMf8kqvRdFxS06o9Cr8BQMCHf6n/f+p0/95fTldbCIKdvyEX9L7q2spvWq
Nn0h0bclWADBw1T1PH7dB2IWy9aaVEfdm1p2CSMZB9bwNWjrz7cjyGDtQYZ1bLjS4JyzVsl0px5d
e9wA/d1tK/IVa2/r45aNXGIcadWzRS9E0XEahtzLByy8r3HBhD04/atAYIP/gWBSoYu/b/Dg4gj3
j/F0U1fToW0QF4i5zJeLi6KRv/Ftf4TeH4y8pT5kmhOtO6aNJBAnkND7T1nE6jhkwCXFpatqflRi
RpPL2Xk1eA1q2zMxE9Spx7eFQMkOrvbymSzgJNQMj4IlDgFIaCOGM8h2NEyfNlkLu5feNimqCX/e
Xo8k5AKgT5zov8ZwQxC0dPIsKWpK3ZcmGIQVIIyeZzCryaVkWg5lLPJ1Wy9alULJ+oM6jEexgDPX
IaHI2WVHk24az8yJ4nAsbxvLSUmXtBmkLpy/W2l7NdZgpRw8ZnJhqemU86qodHNLCGuAM92aRW3E
+wvyaTqhIPG7zRSz+/y4KqcEdqjBOj8SGK1aOzPq/8KPSKy8juz0dv1rIrNsMu4l4W5/DfONUbqN
G6PqKgiyJq/WKFaHjYYHw8iJaMfJa1nFoUDWlCVC+62bEjX27hly+iCLdI1Fm2PdOdMX5pJ56Efi
E9zpKu2sk6eaMkWKycgUO/wcfIBLTfm2aUFVrpSZz83/sGf6IyBvf4mHVl/8t9jHsX8YpqqIoWJ7
hYCFVy1u/F+/5BLYg78cdpeLS+ZV4uAu7FuthHFw4tH6dqjXafwqhNOXK2JQ2YvLApN5zVaocP9h
5LifYVHhhDyUTgCa++b5dr19gW+snJJ+q6T3mtTdw3cB62Tba4/LHPIjHFTxHRs6iTpwQ1Z3Y14p
0mCNhFp86lIB70/p6N2Nq5RUCBpTyQldStxVbuzzEGRNuH30kiealIHiuj6FobFsh6AutUW+yfD/
fb4ChgoSCFfbkVTvXt6R59+UIU/AEhtsGEowmnH0uc9jhl+ed2XMWP+XR5tkizxN+uwvw0QzJPmV
Ds4WsWdDvvSjdpniqULHKVg1wvQH/cqPczoliT6f7S2WEJGcEtcLE56nY3qvb3eGLJWxXRfIXH+g
DgDiaAk9aQ12FfmhZXLHSraJRFDoopGiQzd/i7AC185A507/i/fL55EX8I164yWmafavNv91ZqZG
JBuNqgF+HlZKYzk9QEG0THFqUpbV6ImJR04a3cmT8YjIU9JFi1s9rX3SQFKwqKLoa9oSzPaWPino
ELWeuN7beCPTM9695vXnS3+XeyPV2375DnFDlbZ1fighfG8KcEdkp6/dLjFEVq6jDEGS2S0TCQ5+
U8qyUVGRgtDjjnOjfhc3KE8cz3k6sdErk9bV0Eg2x25UUaQxBPorEvsiSrqRXLRMloPxUl9LLOa3
QeDnvi0iBejIbGY5hZdn9ckjrtljM/ddl8+QTg+94f5dtm2fmrfqoYEDsLKezsvNwlv/5A4rE8Ip
oJ3PvRe/kHvhCqXRSz2jw5omqsrBwr/cYIcMTjM5kD7Kc73oRmEP8qmiGlt4w763DVS+x8IPTkpY
lPfR5lc2JYcBt/dVehNJuWvHo78CBR05tKTw64oWfoD2NYZW4OJEh8LWyxGgX3u/zy/i/ueA15bW
hzJPP+j0aEAPqVWBW0K+tRaWtN+CJwTW8N9wmhn33l3EsPn3FwKTRJNhghavb/7eNbtgU/OxHIBT
4Jlm3gDD9WA0h9mOthpb8fGkatHQC1f1Q3hmeRTzCugYIXX8L2cMBdLAA4BefrMiyEfNs+mnhCsE
rC7OLxL2jDgRwgd4HtPGBXnjsgBZJZKSMRjLALDeizZ+r4II0yhGah6LfTW4bb9fjPDhP5ChmbUW
vP41GeqVVoOF2GYTIiIj8b+ufXcJzTU6wZlOHhyipr3qf72mMt+udSelErDC8faGdttUTX1PnG6C
jjOA8lpt/9AnXAhagr8lYZOu5Q3oLf+vttTzNp75DoZWHD6B1z30MZ/NKzpdp4iVWslDAl0m42Yh
IYTMXScUKBlFuf1dXEWD2jJs9nQ+Pj6ZYslykbg+XZgN00I7EhAW1K2WNpzyrB8lyhSI//0qRiEn
vOFwIFXnhC0HuteLqOzvgEIYIT64ghQ5bBwCwzIBBqlX89UIhB0uyhu0SRo3D6RvT6tReb2M8nFE
a4xVQ0MrA0eYlbo1yTggubQ1lR1tRaIQCXpzFIwqhh5GDbhMTk9EAdRHsx/XbasNdsQWMdUQbsoF
0DyvKYg2ZhmlDPqOKtKqtI2zJ8+2MCgOJxFioKMjc8fuhFNKdkw9qY0p+2XIn8wm2jXucV1uWaxo
Tbz8tipxGtWTOVqJGGPUU4ob5EVr1Nn5Y3cfAhTYCFYOAI7wqiludLWsRuRw9CHfeUo6AsFTvPeC
ZypZ0ljt9O0T237+feBddavx2piG5aS18YiWshuYiEoxim6Kbfko7wCQVYDcINFu5mMI5UJKYVpc
NYhGHEyzRCXwRuWo8VOCNvpMXR5diSlLpVBkkjoZbuO61oDTZhZm4nLHL0oLcL8DHVbkMrwHVq8s
QWLFcSmDVOtPNHBL5rcmzf/yAvynFgmK5hdFohaBfuVlWSfN5D+SduUTuPZrR+aGbzc+s/dZwmo2
vHFGpGWoUzN71yImyXUDXMHPzKfxOIjZzHiv8k2O5KnFQYqQxB74UhY/0kIwLKyHeP0J+7vNchp9
SbHru8geuyQhS4uuxKidQAZGz0/3bN3pSeYeaROEUN1qL73gjny6fgcDWUsHLtoSChWcaDy8t8RH
K1fYoywW19VvWYGG1bBe9EGONPWTZIvrwUhEPIEqf7sx9tVgdxiqTOPVFRjC/snlK17dnMQnfX9B
loMM9hL6MiDyu07+4premV7e7jBqvV86PmfQpu0yOpuHMuaiO97h45XeDrwJN4pfabyFiaPVsK0W
msTTMTq0MBUEsBqaaC9va3yTYtBcI6VJMD7CfJRoBHytzg3M8tQfEfxmFdx36nKdO2PwGkCqfx01
iVlx8HU62U2w5BgEho5mzfW7XBB8P34UXRZ27f/GFtuUqSHtXnB7f184SI+B7TM4Hf79NdktUPvE
OCYXjMhIaA+6ERKl2Q14ga2/jSBRKHPcj5+wdBBVArKlexB2RRb6xHX3imf6Cy2kZGzM13JJdzOO
Pm+I2/qcQniGULkKvMJH2LcpaSpUzY4RFtfwJTZjOlIITzXGkWsw6adlSZJkV8YY9HeZx9W0hWyG
K851sTHTxdstdgQ/ztSJDiY9Nh5L4MFhi+FIvODaJrXHDsxkTCvp3d5PSdFRtcfD1qlhavH6Rx3g
CNbhh/g/5YNG5Av2OrA8nYFgHG6HRj1/x5aTyxvd1/wC2OosbqvlwlaAJ0UbBXIU7ikIwZgX8aeb
SOtwIXhvorLLgIL+a/gJKx9MVAF3zVnYa0b1UAUH9YqXGTnfGQla9aNEBzUm0y0cORdAQO7AoF7Q
pgOrcp8lj2EmdmrQjlr1INDM2DNross3XMy1dj/7YvENkH9/MCW3W72Q7l2iwOrW5YMsj0eodnyE
OER7l935T4yw4o4eh9inO+xDUEISZ2w+hWEAWdejtISEBjxC2qyAT6q4nElejfUeb7rFKXsYqqUF
6U3vYONLGsyV+apYtoGeGSxgCxxSQxrN2nRPBXvXwIGNOzByqLkKpMreZLmL8qD3sS5j7dCvjUyP
Zr0rt2YPy8fpjnhvq8ab+2jAfB5x7I5p4bvlGIvvlZkA4tjb4QK0z2A7JGcHAgU2usiN+Xvf+nea
n3ICjaa3D1TPUT3Pe/OGnIyqAzGPXStV3OhfCHZLeS4EQSRjPYMCjCIL6nXcUXAZ+DW2tyN3rduP
onssbDL+e1oLY67gf+knztRnbmDv+Rduoy+59lb9i/gtepqL6xhVfMjX60Z1d5l1AMGagvCu/z7j
NIeS6x3HAS2c4n+fEfYOl5ZVZCsthRjWDupr9mNNy/9CRFwv4w53cWYpabjRoYyqk7HUeny/dxHL
WZn55dZQ5BXRV2P4Cowtj4MzCzwRbPSKKg2flTIx3l4aCWhetgZNpi9SQNgVEs2oQB61fcGQtL6u
+RotB76GjsZz4H/SqiG/kZqrZc7fyGrr2nVyw9DeadHAIobVNCB8XU/Gy5okhpKBud027IbVIqVW
xcfH8vNs7VXIPSpnuEoTAhzD/SQusq6Yi8zEDIE1mKAI/UkXlIstxrClNYHqTfXNDbrTmUDZxx0D
/IeHWn8y76AhY9aFQT6/CZ3wqjdtKYwSceVJZOPuHlVbehzjnJXMBbSvG7BgSFk7FfLITKGy7uFX
ujRYHMysskK680VHdSXJexsAbMZhCWPkFa+FKnib7MejK4OVq9JExsyVa8Sv/v/WV9p9vgBmcEr8
a3NjGXk/qBIaQfrpb1J2210hDOlStz6lSb3AX3HGkj75TAJzl5wz3cOf5UDi99R7lWGXsL6vQL/t
hAKh2zXRs/RtFZt1OioAs70006LfFP38aJzwMcdQRWCqNqSiFQdlToZUkXa6Nr1qrp84LDuPtKTY
rYASVg15OROGugjE4ynRY3uQBldTR3krpxW5a4D8maN9E7zo4XUHLtUohBGOtv2c81tGViXRks/K
nSv+eAdh5n1tv0fvHIsFWJsPu+6psSPYGFUfDAt9UtQ+x6j365Hbv9czQ0uIuYkh0E59NGduhLeW
t70GE/E/LPgs9VaWT1i0TAxhhQnh0R0XmmoSyQjN5+JBHzwCAJhMVfMI3rFREr7kGFxcwD8ZduZc
3Kz+F+mnGcPt9jLGsh0EpuZH2EbNyiO1tNkeqT/jvFT+r4dHJaCMz16WGLqr1l6Nn0VXl9PRy0ka
FCxt4zaXnNekqMGK0YEZ5G3K6LRAV+ft4N+yzblau4jwXZfuWsWMnffYjcIzAR1B+SR4hDS5L2UK
iaRPCB5EHn36ElYRdVGuy/uPG5KKHsxBgD6z0m/kx7dp+ic6bEiAwtz4e5qLn6YlRHUDSbGtz0EA
3ejEs6+qiNlutd7y6AJ8PBTmC/KGrC/NJ2TaSWVaCcXaZ9WKhxkJc3+a4rbxNfdyEyp7kOnI/Sd6
+7ZNgXXZEO/aLbksa+nZ4b/0PP5O7frHFJMmtgRG2h16SUulQxWvD+4lMKuLW82N4wZWAZCcCdD5
z8/mjKu2t6YiGFIx1ncSCXqyT7Mm4k7PmZWjrUhxtVKY2uxs3u2WK2ErPnNX4cTxc5lKT3Edgbap
GFOdz1b/gA6lqsJRaP3BQX91pqTRsqXTKCNAqxf4+7/8QdP99JI1EdUnEDzPLqeDDGJa3hMOetbn
vB+qV+EaGhMjlKc0g1Y+Om7iu7enTqSDybzSEmHjmjtC/o5R1jPc5Pp8lxOqG2ilQkGKjbmFZ0bw
gsKO0gbyxII3Vkiwt9rUjMlUUia1Th3Y/0Zaplo6a3Sh5Ppf4PqbFEuo9+oRkMx3loTtE73tiup+
RzUIB0V5ogy0dhgxMz/PW/2ym5Vq7HCLgCI4OcMpL6wWlj/eKSIiwpbEavAoB9AKxoozmh255ih8
b8Gm5wou83R2O+I/R11R/uswzxwe9pQ0jpxN5EtBm5L00MTyk0JgHcmnCA92cLy0EANed4GRb13Q
ssaOQg+L0GJVLGXRUBwgvuWuBsaSSF4aOPHkeSzLEY1IcdggaxBu01UCGSi+jmuUoMp4Q6K76O5P
yxyJL3KqWv9Dv3FHJSGTBUoSk7sz67THiKZfCY7sFFmwSpa5fJx+tdyFVgxhxhGp8LHRKcicCcwL
h9ieYAUP3t31llNs9L03wLiljdEXWN8vYYLuFxVkfnYk1ZbfJNPnGYXZQApxFcYe/MxqShEWBsC9
T/RhAr4qhxO8hE2FXI9ar05PLp90Y9crdrluAfqKrRqZTWzNii6w/xb8bfH48z6mwZYU1ESkTYXS
pvJTi/SuWbCVYSpuBow62GzijvuP7bOOLtrqmmoUoztLJ3MjgMbAxxtvq7ni8YdgWlCflQjDcXWM
QeDZLXMSZK25f0PsoEAtT+yb/mptrxgs5Dq5eUKzCNRFP009ayY536GAVW2HzOOvlqNfHLP+/0xU
cACp//tc3J1UWCjUvoYIZHmfEuJ9WgkwvZW0B9YT0qokTrZHafpekLfgmn0YSHiTLsKLLetEyeKW
husCpiQ0ts+abvJI44QmfrDZIOUbrAale9UfTow3XSqbZ1P4IYams3rEczRpy+6ifpoqqb5nXWbT
e2pIXNceMW0kv/RZbhyLoz79VhrtvKh2CCg7YDvKa1Ma+ydGh4ME/8nCpDroNBlLjhznCpdb5s/n
/cn+Gq6wf4Nl9RyFXkhRkcCmun8VoasAyENKHx1j6SLJtlKm9sZiDlfajhMugJ5BnIC+3ladiBpH
BWOhhu8IKRnUSK+N3oWeDArEBDcYOESI2wh02M5gJIuvMSnoW7FvwHMA1dSIUNqX7KhiyPI3bfiJ
8pr0v9UW1nZ0ya5f5wnid/8Fp6RCRvy5tNeNZ7RxSruxm5L0LWX8JY9OStdcYPfitMtvUU3hcUcj
hqfWRNsVa6gt6f35fpzGTf7fvfR1Uoyyg8kSznmVGvGVob3LS9rAbL3MREcEn1INrR8yspvjRiLC
RsAGvZ8KMiunknQzhHX+ArbqzgkqJtC1tZeijedVrkcq/aqEPiQx/RM3gzp5xoYZlc6E+/uRODpo
ECbe2jnmk4t+v7jzQQ5lLc+fy7F849HK6ysyyVwADpnsx/8Y75O8FvNdykPfq8AlgXj6mPWf3LK1
0cAKNaCkkwGUcBFjOG8zOtrLKvHZ8ULGhy/O1s6ruQkklmzV5LO8j56A9t1ymBSc4ge8oxVlNqgC
nQgETgFw05mh96gXJyJmavkzyE7EtwJzWTXmtV8s1ChIwO1I5gbiRLAKFXw8voY0/4f7RPi2ZwHL
C3B7U0ifb2zV2rByCAGjiGlr9yRORj6Xd03tkuHG9uNkF67hbgcmOHbLuu6wNe+3TEsdmgEV7V7U
sDpxuKLAPzNTmSgFU8jn4s8xawabvda7I6toUvRObbaIlRTd9Wyir7vaU9sJGa7/tUeEfi9LMGzt
3SAYKTrt6ZIBelH9mprurhg8FI3eSl8z4NesuB9DS6MEHjyFjnMsp6l6QG3olmwiZLavdxqRoq08
ycGbbKOaWMncCfcRbuaqENiuZUxKo6rETNgMDvFjyWXFAhRAt9G8nSLk82HMZJM6eUsPscfoIoj2
l9FZoirnQzSQADEcA0efQvb6kspk3VEngoVqH9dh35p+P+jo71BJVkpea5Ettk1LLSTc2Z2Q2P/N
mGkJ/5XnHqC2CRKFnr/fKooAQpsnFocsKm0aDcqecjnuJUmtnMiKGuwpyG9Li012dR3M7GvMhSgQ
63+j1nmzteQet+d9MysFxyepHnlorR3QJsHB7NewGd6XYJg4KPz3K7eWAzCa1x91zo1Sf9PxPWCD
p91a/ec+jNYpn+LH6HqxquarSjtA27iYvbPqumdpmy3cDtNMzYNICy/ePxM58KMGkG28sHyVgh76
ujgkoh3WfKbPKK7wwbMJAw8fW6Q2syah21ZwQuS47Cb0pbxMIh6jKjOrcrymFr0v2rhV/sJdPtaF
O90JbU9ULYX3jkOyMWc1Xlol2WNIRBZpjLJh0IooKZQ7nFOmZBS3Qi+k7NdFgwIhNPs7uTOnjx2F
CXBpLPpZfl9kAyPwcvTwbFkHipwXCImYBKcCYoyWW9xVzfYr9UstRbr5hD0ENseUbc6M/+z/DdVc
TYacf0CQwkoGJ4XJ2pOi+W4ZGOqrt7HnX5p6k6wt7FsTXdv1WB9nEePHKBaLrgOe2iG64bD962H0
WLi7l6Bco8xTH/gbT9sD5y9ukfmEXHJW5AUO+7Kh3GoQF2cnHPh4L4LTwEiDEiOs/cTnay24qA3+
7kNjTtvGObocvLR4OtVxIkJdWjTHVwKUBM8CGLLLQE+hPfsd+5soB9Qqkrbc+8XvDZDkutAznax5
qQi+Io81WrzoMAYvtW01FWg6Idu8tPLSz9wYeIowcxn/Mmd33wlUmZXNneTWdeSSLEusYAGoRM4z
3/Fa27uiYre+9zFqnfZnVt9b+ExqNgNOCXIbD1HPH4t5MTSHKxJ+J3hx4JUYU5LZ/bOOKS35y9OO
RYn8CNmZbhD+IloNrTXlg6yShiGxj1VyQ+lDvxumAxk28irVOsl0Nsif5J+TXnBu4KVj0F7nhxlv
6n20OsJ6LYhKN8GSuBspMPfu+F+ZaITiWqTvjktRs8tyTcDMUIt6S70Ol/n1p4oxAZknegS8HMvr
/Z05raIB4F3eQHK8MAgrhfRR4MJ0ffkCUjtuqO0R7CN6O1bdO8Mx9iiKQochis5L/0flCrIuktH4
lmouwiuteIkJTQ6ARE2OkG9sj/voDr18SGuHSHuTFCrnhe+XFCBTgUTomjyybuTTRVIfUGcamugK
6lRgwWayEbgAh2b7jYD8man2/N56IFsy07Y3aRBcsXf7YRyI1c8q+bhBBvcRIBChTJ3/JqP7dQID
hecJI8+E8lA9VtJeacdl5HtiZcsDqhu2os0PNj3x4Rt9lzHLYdcmeZLK6/iCo1y5NE2qik5vMcC4
r8kerStX7Wnv4HAfTvJgQUl5M9Fu4csdQLmjeie6w3azxkgdzoWfYChwHYQdr9vpYqPhyduZIALn
tnGfJ3PCoom2nd3YnYevyPnFBhFvqosCPD88eUgas/J88OD8C1gvkgW28qvOi2d0E1EM5ADrwmPv
zQ7yx9+osBqQXpH6PoggxFotuYHM99upSAIOEA4IXHAJjxuAwIKebEZcuehTB55sTdQ7y/Hy9ev7
HqTTfJ4mRn0x7V+sdtwGCEx8FtorfPreoJ/M3hQvdelT8PrYZJ4lwqlwz/TxhOVahTWXxuBO7H0N
JqEsEiP32WvA/8vmlXEfGDYKdRF8zX1rE81L/OrLGK9IuIi5ltx/ecOn8fVbsCM5uLyfWhvIkNRK
PynZfCCsOontsyNzhIhcCoqUA2Degrsa9m4Qlx8sTuLOGNnX4/Ucl3ckzc9stt3B/G0I21rmzJoS
6CeY2MYpS/29ginq+hDEz1nolcO5HrNdsLMbfES/I8JLGAJZgPYKtu4dINHQHGGXsMyttkId12av
YmhHMIlPJoZ1KbTwAq1H22I5eJV77mktzB1BeZgNhnlJLWkzmiyNwM6+okXK3nRmRJNc7rQzJ9sF
v+IJx4HSlAOR2CYCTJf277TnUPIeVRZWTw3mA52W6+B4DcwEpvRP+EUT3b+qudS2cga/ES3zhcza
r1HydvWvgXGva1NTBCnv7/r8j9I+KKNKW75otQuyB7esZAjPZm+OL6itTz+xY2LA3QC4ACmYM8B3
gZE01dvUOITY4QX4M/fdfYODO3ES5V5whB430WoZJiTE5JtX1NJxkbXc3wRE6OFVsXDvv7usUB5u
817KpFAsI9EfU1rghpeGDJai1ik2Id2/EgjJwkkFVW4pa/iv2ENxFiI1q3ecMFfir1P0zm2749Eu
k2tHGf6qNqqbsozxpF5yZJ+VS8QoT/hE3dFChXTqvv9AjqPtWTuAfKSjk6wqVHJTpJKcAjadrKGV
RV3lfwJru1jCsTsPVxpaDfWgfEFxR+N7NY8nIlRtaWvGPhwuJXHYw9DNm9OctLv9AxEHPoYi29x8
//uRuh9RmRt2tJzDtWPdHrMkRtkLTBQpH1J703Du4hQJcSVX0N5lkz9B+NXW4NcItj0hsM6ZpLm/
tIVAfn6NUlebnLmnnSDVKZqyCRraI0qhkA07jgckqd5bCv8yUK8R/mX8djWWjLg3as3UDpFBAfnp
HKmz16GyPcGkvCWWm5f+sLrsdDr56HJMo2PGuBlfiCn2PO+dL3n6gWHFVER6sjTO21pHBvVWM/vK
grEVgQvh1N5HOMhCQWBkgLi7euq83KVvrcVyF2Gm2AOI0vEc5f15/WG8UkeVK97+kIWAe4gukaMT
TMGgT7Z7rOkNaSrz++Ud93/DpDAnOR98iaDdXEZ1eUkP76+9GnJdruRetN6Gk4BiiGv4Z2hfKU5h
xfGnMfXCzDT9htDCJDdVNEuLtapJ1hVsJD6YUzeIO9ErX0dZp8C2omr/PETZG/yVPMn9Pq64V+06
BCxe65ofXjQW7nfKiLPBRAZ3/Jrf2bJcT9qT9OWIQhHwZ/mKICQXnUQ+oRkHegXzTxGtzixRMmDY
Zp7HfobQwxnLapScRQ2OKxfThJLKW7VcnjuGklRUAQqvpcnz4H0SAV+t/V3GcJr765Ar3EuJAPwt
IYsCmkSfl+YdKglTglGPPx1P8dL5msWKcYX/zrq51glF+9kmPyoK44ulepM4YHc7H8TPP4SbmPc5
WGCMZzudyEkta3/po9/paHRDcYgJgrYJ/80+6GGIh3l5tB8g8u9ZNbuRAmCI9bnXcNQ4vENt6tS5
oMlvmEnMzNnqU9atOykqQuTrP66r7mcA5iEffOfhay8nqHcp7wHwW+J/xl9OgLfDFTqkJQVX5R/Z
cvILVhfl7jD989B6U/hlHFJkz6XT+PIm6YHU9NCz+ObqRfn/QYbJsS4cWGtWz5CUCJepZDeYwtd8
5oHOg9Gy96/Es2BBFzkhWbnRYX8NpFS8RiHr++hKaNtTQ/Fl99tX1Dlo5kMOh3bmG1L0arRRAOMy
nwtLquNYFmOXSIKcZp1ZuJfb3qWBsqx6qCoMD5ew98hEmgwOASyti5mGtelNStVwUVmyP7vZUpsP
TlCq4P1Sw899ZgIWaR15LcWZO4dNigC3gGiXfp8+1ykVDpa1mZ+CXgPRTMHx9CtY+So3rQ4/aQFu
rpny2i12cNJPW4ZmaHGQKuJPHXCnY1Gd3/bnwaX+ocGngxxM6OQjjJbopQeJu1lqwE0jWELOpaTi
vEHSftLERPaPzdfhUZd2qlxeAvJ/VaBFIJRioGYRpRZzM0Pe3mO64BuH3xWMpwxCKiOscNhEv/fy
RpNfr+LzNw6bpzt5oetv+wdpoJKwzMuojh/oTL7+T+Gn6NJZGJNWceVKhm0MBTJwtVfND6VEWJyk
0KKjOioxHpVewGWEl7DnTATOF1t3HCEJpqm7R0ipJ/ckgKzmp4bdtQJhQVZFiyF42yVa5RDH7HUm
YV6aTUCQPSsvgJ8Qx+vaZe+lYPokw5bD4oSrMv5qw/zT8YNJyaD96qdRBUMPMSF9+CvAMT5H38lA
tpHOr82sP4Co8IIIGTdsIkZKwxDQcxgWPZX0S+sQ38voqhA7UdN2ChOpt9T5TdfjQLI0X89MRhF0
P+su4/QHe5MOpndzprVn+3Y8aP6FBPjfzCcviIGWVUoKEEbaaem9qaphf6oBoTB1dlEHmPsmNQFT
patSzVZ+AMaZS0bjXG8waj9MlUePjHPCgoXf8dJbIL1UPO4LEXyTVTgzNS+2DCoUM+fjpnWK4c5B
mkGZUZ95Yc8s0egHXILu5xh7J2QDGXbcthjY7/3ZeRdY3YmCL58DiuOOhbp40lBype7zYDhMgAAl
+RLpltnpMUO29tzHPfmHPnxccMVt5kCuELVVw/5DPpNTf+FxM+cPN5Qq6+rI8MKWB1TbRtMaRo4j
bTS/GknRixbsJ+YIeURuUS+VoyTHtP5hQf0PdHfjfPO609JK8UwO3MVjm9uoM5O8GM4nr6scMGkF
szGIdwxNbd+jdrQryDa9iP0hgB7jRiNlzKG35wwqnZgM068TDSrSz8FqgDW1UyM3DOoHVS4tLWnS
1dEhArrsg4ZgKTx/quNQJ2efpf/KZGsy2ZUsH14YVYhqwc287lFYZmCSTU8eeADiJhcMJDOKKXLa
7Ieoz9daF9JrgPSUOjtP92ootMcECR11S6MN9up9Uilyh4UGz4bQIEfJTuPB35Ag2RAt3NGkWG+K
j257AmpMHMCuIBO/pkFGOxhtYO1cdaxM80BKVhjCIqzB21g/iGSmVGdj3GkaKjA5ykpvT7ZpfJgk
Y1be+IQaGjXW9xkZ05ltP5SYMPm0YcpRcwAUCkG1maTh6pYAd9Qk9Vq6mex47D2P2aJKADT/Dcr5
5/+tos/UQixtc2axuQPRax7xrD1cmtH/BXDZAyzjRAElGtm/Rt3B+8rdFfvpDZ/f2yFBhNGv3kT2
mfPMS8R7i4R6HrT5xq4ZvzOAyeow/o+wtYeEcvCvTZ4+yFFrb7lVScVd1R/aYDxL8gVdIU2QG6l+
SVLDyuUqNZJYI6va+xPa291H5iF3zqDWVzpYdHpijGXuG4iPM6h05Rnx7/QRL/32JWmbC4z7fguj
Xdi7yZwU+7aFjfhC9K6/7y3wlG8T/YcQxCMWK23kQfWbqgU0UkV13sb+uDPVX3+U3P0j+ChoHtiz
Mhzko/GtSBx8RKQv2j4nHxxORMUGTJOtRsDJFFqpUg0BXuSvHywGHGlIOUwPbHe6EM5CVeXi4slf
d4jzmtaeJWoCG4aQAmNeawXmSpbWLAHSufXM/sohTVgktjYQuMgZTVgIX0ezPVpQn2ds8uDc7NIZ
3RVWut6+ApArKbZDy5daKLAYqLLAjbzVHtsDdzctbllvTPeuco8LJ/icN1MdGSUkyjdVR1nS1wRS
EgT+ON5rTyH+DkPpBlo6dP2liA02Z7Uux+KAsquNJ9R/VXxx/hHnH37y7wr9O0FLrExRXPNosgAr
op4S9fX7U/7FghLH2sLfR4/QAnHGwa6/9BDnhLlaAJhyfrlZD0cu6kQo560qWNT89frE9RoBwdij
UHWdTNuneZWzpzWUpkuDaCxKBocFEJ4C5RaZolUjj93GV/Ut9k+JAyc8QaTfjC9H1tyWIRw6qWT6
n0Hutk+lPABo2yscxkSJxBInjcv/yjWHlTDteoPQV/co+c/JEPo4orPJnwmrjxxYAhqbKQrfY+VF
GUs5hXVqFfZReEDPK/qQTDc5N68DNlwAaELLp6Fy1ji5ATSa+n6osoTAW7/eAuzaE79zeocX/mZF
YgJ1H87vCSZCeIYjSEH2sQnW447ZvkVThrTghgfgGVHNz2f+4VN5kFyd7bzLzfxTVyDWbQemAZnF
PzL+UddffjXdveHrQfNhe2ZG01Re0sTZsVjFVP7M849iozhFNWr18L1KGWKpeVwfx/Np1I1eV4Jy
bhkV55LpBevGhOaEUqrLwsNM2YMuBHErwBhowYH597qYCqK0igmXUtE4y7tDkDHyJVf8FRfR1qTG
Hl/Cl8rQio8mJBN3u4YDbjF70sYygiFg3DpP3TBU55puFBP+ukFYY1QwknEWTKXSZwn6+52mfFYX
5SBRWJMCAALYGT3CtyWjeN7UfjkaZ9HhvU8YI3j2J2QJOxGuLSBb5vywqjOgI4a2z2ZHzdRA06NN
PbtjM1z/9ZUWnLxedQlxNtWfqygk8DFQQUvtXr5qNLUGVw41HBGu8XR6XgeuabXKK3ScrIR73y3v
Yp62ODbcanV/OOqt5/7b/z9j6n/wtcjJpm1YsheNoXh0l6pvulVfI+qJ95f+fQJRGR0o9GMHastg
A72STiCFOit0mYLZr7svhsUeIvxbmXmUKFDfv130j7F1y50nQbmpdMUPwa8q39kXLKt5at9tMNmz
KYBfVLZlgUKJbLrmCK9kQInAfwC5sVzi4yNxM/58E2ulPhj1VpWk+Qs/JD/lKk80BvZJCxfkSTVb
8qhQJha1Qlr2wPn2oC1H9LNhU8Jr4jqEyTJpvu620RxU5UILH/2Le25mmuZqgoDRxlv42LSv6g8S
ZaixyPyZpbE3V1WpOt0vD7UbSDVMdmKrZJp1dyntsB9G6DAA2RwX3UvCT7sv8bwOSrKexgYxsofQ
H/kTI7Lne6dIfzoEexTiI7GcfVejGYz+Ku1GpLrrlnt0qaJzW22vxym3pb87cUKB6ovh3GdAWTZG
jPNj5vDuiHtP5/4bEIvYklNPXX0w1Asfn9J6D9PyRhghBECgYFrGnkqjxLGamOrUdZcw5/WrZLs6
6PPgCMH2Ax3RrJGdeDK4YMM4Oj7VuvaeD2A8fOrt3glsioWssHXns+OYUQF+8A7rO4O/bC/BqfuG
dKaVPiXiNDvqhqV6U/8+J9z/EzHcq2Cn9xJ/q7wnOOyi9x40PRcrZxi1ti989fyezNTt3HmJPaHD
IcbScUjhHwDyDgn5YiH59TXC3uVggnq0k0dXiMzralWBQdLMgw+OUegsDjI5+E+EJwTTqzHikLZx
pAHOY/+UHV2TVO9NuBjrZ0eoGJuAl7H6r/dalgXEJV3ZP9YlTKRZmD/o2sCTt4zqKxL0GC74YoCp
S9olxMYdYYO7cPJ6G9H3OJaK6yVDTWvTTpSQ3g7DTeMXjfBufGHeVM25mtXBVguz5yrvswYQwU2L
FGrvHCXAMEZCSw2NA835fAVxlf8qEi55ZuhTC+fq/Btg0TWzValG/+/40uoyUNbvcQJsmsnEe1yO
kkB6IonrP2Djp6nxoVwDI4dvmV1P84DcQXchezf82GM/6ytfqQ0VJZ4RwdBWinOhkGbqEjErGILy
O130Frwy0hAVqh5Duv/Dt5Dp/9Xhg0HeR7/r1pRT39qoB+vi8KSeXWRqSmDyMnCLH57IaLDdcddx
uHorrhT0KREzjdi0SyanA++krWkIsq0p8BceB4+wzNGcrZu6gtA+eK13pkyi5IZlznbif9pl33nQ
0vk168lBJwnQUStekOHqK2PBgSPWOpYOh8T8r1XW8bdr2VSw+gChdhmSgvlN3bGxV29QdMilbnVV
X23/w1Nbtt15L2AVRMMHFO60asv8NV8gHfXBhEyTDRdZNdYZnHKaxOUxeknvPSzw5wn78Tp6rnXl
LqZvUPEgGDfpjdFE4SrrwdKqBYAxk/cI7qcGlpO4qx3bPNltYTC+Sna+uswPbS1efonBJATEfrhk
DjSYQYO/n0weCdtkBPO095KyfEuRoUL2axv4Jd9MnXhcSG9FfdPVMafjzSKTedh3sJZENki2w5xR
Te4zjBIMQK14ukcM4d7OelE5DBU5EKefH01dDkUBX5jbF34dZDBGEDAryTuCGeO0PEz6xdT3TrGQ
bZQYo44Z5da2xgevHSbZh8TDUZebC2oChSCoRJqyXdMY8by1q6vs2CumKa8M3pBGL883z5N+EZYJ
KRk3X17R2YLumN0B2ORBDdqtGmT+wcwwTOZwKrTecTi2h3DzNyb8M8IWMslzbfAB8+S8cb2XAwqw
jg9wb+PCGpPhi4HWdWYUaILyDrLIQjc4/ARnM5YDyBFvmlVuLYr/cwU8VtPCdzAKBvc37vk82NRP
AHwqb7fDDpz+L1VVuGJHgblxBKvq0XpEl/OqSwrK9c2MSnZ3Meqtva9oWfYp/sleqnwuELB6VU/1
DdzqQlwfJbsSurcIAyoUaM1E8d5qQW4FpWKZCEFWpT4gInaurIpXsvm3D0mhzwRliIXnWO+aLGFC
d9JU0qv5SL0MHoW6Q330CyKh6ksVLphtJoofq9WW/MmGB7j0Jdcwajncin6nnziajBlv9b9KxuAB
rPY5iRbpo0HxN+AXul4+nj1fHuYbBSLtfom4Y31YA6KqZFOIZn/6FXbWzfXVb8YfCQ2utHateFHi
CWCZYXzsxqKCXhcnPFqFGRLyt3WHJ/m12S6IAiDZ/D3MkmD5RAS7nKBqBsW0l+6xI2WX2/KI8UNn
LeaXzdOGKyxcc6sySYXPkEaMXJdu/hGQ5fQjppXNaMwrNmgGUNonWCo+3kARey1aJy3viscYkXm8
p/Eh34jnbWOA5G9tH7s5222+5ce3NYTTszWhusrV0jXPEsU0ugsX/bYNRsvGBVzxpLOWkbhTZFB6
pT1D2O/JfZwdFG0kPMUwllKUTrkKVFXlb2zwxKJ075wf0E+O0xZhfF9Rv2CDu4D59RVNcaxKjmPd
DxrIEhu3+zSewziPGjgNTnUMbG/FizBu4THmc7KVmEVO3E4SNTZir5QjXS3r+CnENoXJB/WUF83z
/vEaX5+v8LB6+LV0MM+yzc9SuFtXwO3uS8Ag0Wncyzp88PobaMaHmiyxC3e7VuyGXHKbxWzppGTV
aLUKl3a78uBnutlD28mMmpDHZqGCPx/PQ+HzZN0MpdgrUtHRrLZbpv8wVZtdh8ckPllvTrN5YAE4
hHR8c6kBKmA0j2YvqfOK3OuA2Z0Cny5bB4RZcNL66/tifR1pzxQf2viiHez3kr+VGnVNnXLbrS55
21b4egO1EFwVB+px4VQd9NOy+bbp50l1PGwn2rxj0KscBuLpb+8VPuFRnDWxGAxY+0Fk84W9wZJ5
IZQvWCcQvh6iqeZtr1/DCbQSDZgU+4c81oAXj48N01t5fL6AMuecgn2sNFMiHYAJRrkMw3eEd7X2
6MebCTwE1qTy/7psIvnXUx/tAzfqU715RmFmAevGnbJZXJhMu/mFJXAzRuzrCtUpC5eWGuFiSyq3
hKw8P1gjBo59Z874WfogYO+pdeDJtVwY+GF1xdWgANaSblODo6I19FAYlPFOWiSxKIrtye4InFz+
2KAuNgUO6IV/njVpPOJkFJ8fNVi6YamFnfO5XyddmJfv0Ih4Yor7ks0MdVQTDkTCM1+M8A7UAxA5
AsYtCB3Ul8z/BpFZtxyGE2ifid5rv5Y4QIuMxr3zuDetpAVxI8IsL5wjfi/4t3pNzkPX9v0roy9b
KoPGfPPc6w0gY1gyYvyiTryt5BIhlgbblywxz3gqKxDmHI+0WsxKxQa020amKuSfzazyv0bNiXep
8pe1cjDCAlOkwbi4OU/XGoO0NPK5mz8Qf+Pyi33nbPMlSo3MHi6TUK/QeIU2NlcaZaZgOuVkk2fe
tEg0IVyXvE9JgzhZ3Qsoxz+mQ2Gq4gtJSj8CiyKM54VbsbyB7JUe5KuWCVKCsjV1e8RH069LQRg1
rwn74ewvVDW8xXPmvXXTIe66eBnGFafP6QkED2olZ700YDHOf5WTLfo7MfBIGpnUu7GVC3RcAJH2
Ac3bslRTzGVQxrrRHSGUxVDXAjMWNQIpYKXs0B+J7QYHrWSZTFJgbCUouyTlHySOiKXN80QRSFu2
HKpO2cxxT45tbGXD5KDL5tE3olqNcAXwFfuyHaEdq2ofMAKoPQ525P4VY+icMWY5Q0TYynapeaZn
hc5X1WRJlYltiS6PNhfswjVRhSzAbqbGEFwullrU2R+ASEilhwk0YTGI5n+vFJvUop5/4Z3Xip8M
Dm/naD0fLXz6kZreNNJGEgkt9OwUvRPv/KOzpwQ8MqlEsUnz29j6v1oYfeGm/pPWeoNTXDMTHnn6
fFUMOAAU46GhChSv59Bg0uSO5SA8UcB68MeSVU5bij6zJIb9QlgO7+D5VD3awU1sFI0nRTT1ecbL
N7daU0F1Znr0InX0YHHRIqta11oB27D0tbe7MmHyN+9e5PqzdUECKpXz1FVvfNoWum5wNJjxnMEt
PwXxc5SYhEk6Zfu5EMPJrh2FNNR+zEwYSW00jevfiP2LVtxogzrg1xbMa6GReGe17kVVx/nUCpr2
S6WEgOOtbwF7sXB7k2j2M3JpEKI6XGceFGADU6L2OxyOZKWBhb5onZ29Anfwvv5a0JhD7oYAD284
WvT6VXYoVj2uEwf8b4QkJVOZa2+71hc4LGJ60ngoa2M3cMRacD+jBYH5RswCyC/n4slKARxxcYAQ
yvQEhIACdY8B+FDRsdPfIierKKIIgEqhMS0gzglOgYhcZ0an2DBaO8LlsuCF8uzxh9VDCalS9P+B
L1vjPr1l9DePNKjyAhM6d7UBXE6PDu/vsSCQyTP4tungmFnQjlh2zDeBwxffndUU1vigqH2E0zVd
4cf8qa67Tgq45N81pUULHwVPLv23mJNWtrUFjEerbPAH+Rvv9KNeZe4yRa62tkZ3I/OZ1fHRlZ4a
HkG8mCVcBZkZueggfrK3YjwJ1ToND+EHsG/VdhIh/fkh4Fz09ywtiLGGFltcbW/B4Xnd4sjkv7w7
OrkQE2eiBRZmZr//IjLXhYnLQbIeYY8MkBu6/0SCKjhCr6dpw5NTYL7XRVA4fxfj0IE22Pgr8qhe
wrOhiizAN3Xc2VtC8sqobDbWAOLXy7RmdOQT5bMi5HoXmzY8Cw4vUJrTBA89c5WNhOXa2GVJjyPD
14mdVGeMqG00e5zau56Q0I7bBbtMJt7lHRFW2rkOl5bHK6P64fv9PAjnUDwH1r7/zOylhWNB2ibl
UGjsAjpkEijTyy2j95tGGWiPD++AvciGNABKo0CUraBZQ2x87r7E+aNBBxsxlEitD1x18CUFsceo
uvZgE3O/40aSYNTc3KHzPoUaDG1NU7YUsCLsFqFRwSuxLdwBnPRtCjH2uDVhkL4V5GYEOWaR52dN
96KTFchGszJGbrw3UbGUXZiuT92Vy8tcu6gOKUA386Ga7RqiW0WT+LduNF9UyswKVjkTG/ggQ0Yl
+3BL5dOIRcr7frKYn8COi5ZzpZ68Tuamfvdlx/1iCcYakMIXwbmEZtPnGHtXZwlDuIn5ZlE5Y5Rt
81JHHcxSDRBpMnz/ujaZ8qUJwQMKsgUs4SVLSBmzdNkEVHR1lGlO1vSiQ2drWNPFPDL3moq+2WjJ
aMOPtiLyYKTy/zPuQJF4K2deD+YnEpg6HhPNc2FDdowEsZCpLfy+mh/74tcqhuIUEgdRY3Ensla/
7ZjtyFmdv+iYWWLUBw2uOuzMMxYdINQMo2VScFx5f5KEYZLWViXgWMY2HUmH1xR8GdVLgdLFN+eo
s7sAFqCjPCecwmx+sJviU2ZJGJXIe/Klu9urzysZYNc36KiHijn6Lyz4o3eUhtwcwD2lrxIkBtfE
jwUJWn7mX3VZhO9N+Rf6bnw4qAiyvFhtH3Tkp/DvF0aCRDyeQ69NNDNf+w/hE/UDA66/2xm+fYFc
1sb/4JDAj/atJtArSkicMhb+bkwjwi/KdUmRBkNCFhvAR7xj6O3bK8qzmEmP+Utci46PbV0J0hb0
7UrQ3AkJmAn5uSVHk7VOB47KO+pgXD0gYe41XfCakKa2QFOT0KtZC129T6xdx47sMPIi4ERwi7r9
Hs9ebcvEn4/yHnHOHDjhN7NTRNJScxVh88d8EBgeUyfTtIn5B7DYaah0vWPSTxPbed+5HruDWY6X
RXC6GR2b/OMMlx8G7Wa02qbBaWHkdqwDrZmKzj8K3bjMlNkYwPTjFksMZvxHF3MrDu866s8mRIcU
rBvQcdfaFDSd/IoXDCY4fyPqQFZW+XOifzsV8MZTnSM4su5cwJ2rTs4LLDLAABRQoRaO99NN4x0Q
XxRtKxFLMX4bj2h5m1Y+Q80GZk7kMUUXoA+rCX0KiRhk2+d/a5bv4FWecHuCgi9wHJ6V/heJzrW3
k/I4YYmoxKBCF9dnDEWtmCJ9Qkaw+bfaqySNKRno26eIcxok9tytCGPEFwmWKaUnmomSvbZuqTcY
QcyKc8b5jnfDJSzSGFzh28yT5uUhITU4pWcVM7spbObWJnrkvfz6ZZtgxqLISktseDtzPSGY5cla
5fcI1TsrgqouG+ztG/6G9Ltn43mkeHp2ZiIf2Slno78q92ZaNs8JFcYsFLuMFKNpaealJBLAW8sM
lhp67yGm9/DevJ4NbCnC4PSS5MQLpUB1e7bqvfotS69ai1vs96j7rfgPlvKm9uPsdQh+MQIWBUvp
fDJ+o4ACfbqPEnxIekFGE/A+xx4WYdYzD8ItxT8fyrYucCAFJv9MQ+gCqcFUlzQB05/orJceuoOI
hiVfNkDNB/H01CO/1SN6CNQLPO++0ZccoPQTQcbb8PhOVWSwH+qf9mBcTo4X7fpTYyQsmjZ1ZVaS
o6wTEh6w+rturbZFGbbrLzd+0nkayF/zQUV4QMidX58Rw+bcEH3uQrVR0jxYnANZVHGsusHDJU5+
LlF6GI2+8QXK9NfE1/0IgBn1H0vyViVRzDfgRqTUQ9mjgoIKcJ3RGc1AtOuAC0XZrc5EbhCqp0a0
qCBzbz7aLv74rP8pOQd0tUEoNwt8L+7IRQTfuDasnydWe9x5hZvWciE7tEk8YLYUY1SDk7lHqcYi
Q5+1b2CbwO5nSK0rXebYT3jDrA7C2a5732u9QqwnZu7UZ86iXnIMNOuTDjDq0BzZ5To0q5b0bG/o
horfm/GwYtbT94hUPSYkCBuVPDYO4zIyn4EnLFKSZ6LQh3vTuJiLZaMWXW2rUJuytPz1XEO6AhAT
YdF+hDPrTvmYLoSD8R24eJaDDRpTI6C9vljVGzkFYiiMgvGOabkvuMPLYUs9oZHC47A6FhccR7tO
KTOdgDqs+y5hMRKlT0uZnrxuo9LAHZkUzOfU6t0WP+2F2TJxsnpcuckYBgOgVZ6ZhCTHZmCADStI
FhU3ZEqBFsKDTtrsBtHPWAIEgemy7NDj48vC8SBX9MW+4aao+19Rtb2Jw7iJdFoMDs2ntWPyg+Tn
u22FfbegyX7VZCTIKgQ/6PAX3key3wQHjtrW745HhINR62NkoFbaHiChh7OkQN9D55G3TdxD5L97
Bfg1TeApjyZ7C2IectOog3mP/Ew6/zzonxUPKyYv1ZhTIiXA9oSApST+r07AwvLFK4LOfgEs5XPD
5VD8VtJRr90P3Y2oeEzaoDyYJAWYiRZHF2PtsNVBG9umCQCeppvQaW3j9g5BCJaPaVl8Erm1EanG
iRPvDrzg3cvpyw0bVuX1wxcQo9Zsw9fgPrZUIzbP5XUPM8qLG+OxtaftF30T3+NrHjKxNNsLj3hi
vt3ies/f4fXVX1PqF/DyZOGhx82hsinB8hSVMmECRUTZ4BfW1MrlicJH11o1+DSQ1ZZshNZNgf3X
I2iK6rCM3wUXRZy9XFMUtu3nPdQM3o+jR3rpsmLCIBiKD/UNzcvMvKdlMOYCoVpeB0p40OvqaZ37
Kfnll7GK+BZzR5/z7Bf78yKJU+zpb0So/oUFtmt8IPhkBP/m+49c5Js2PgjrUFMR6mnAJvb95Sgb
GebIfp1mq7Ab1qd8laTs5Gz5YB67USkM2J6igVeoIWlvJCi2ERybuJFxqRhSsvwyCeulTH4vmew3
AsiTuXBa/MEqBmSBX2hFCmtJfKhFyemHAS/niluKPw124VULhZocELCSjBCRDHdeZ+IuGixaiemV
mrBTtC5KHDtV8alCULc2jo9oD/ASEwkkF8pzotqpsSiNO1lgq0dCtV+3kQIh5CyWU4z/LJ7klngs
3w45qMEVVgXCzscwCVy4+aK8yb7lEpSyc/WzW9VEEZMZaFE70C3Z95VDULlDSQueDU1ioOz43Ro3
eR8fqu0CfzFdz2RsjbSKYs0ZR1Va/vvHFO10eMtPj5VdrNbWgpZEgs81+oggUpge8Qy8hvALzBoG
Bri/C432hjDABXT0vsUJITbOYSTRRRVyAMEt5caOEuwDHzTAiE2RE+kRT+j4ZXfObAUkgIQBeGuf
aW0UHx23OjnfTqWb0b8SIj9tYIKlF/7wFZOW+VTQA51HyWh6vdKHOWNftaoYiF0GF5NIRzvLBMBJ
dNmRBgMPqyokvlHJa2WRBkg3sUqcGZuPxqckCscVk46sXZ47HL3uwhzUfEver6tlN5cO1Mw+I1Q0
F0uOrZLTvFkc7CVFfqcnf303UY2d+s9dwPYMEgqp+w0VKZvSLOvL1rkU7FbIofypQJ6HLlwioDMK
lnR1/7KIcJosQozy1MEkC0ARxI5HL85jXLzrdCwziObmwBwrq/LpXDW5sX2Xzy7kxioqhUZkqLsn
A3VFh33WS62m/0RC1JyOgtqNJHAXVjCSS6T5S2fj3+LC0s4rcjKslsSCM3PlDnOGQ4CblT7QRYcs
exNLIznE8tvXGRQPJblQrMQ8OPGvSPWsYTZwouwqg3wZ/9ozqKL5eoVNcKKGtUtsLKDRSIFOaNqC
cWA3NIgOf25xRoOFdjCD/SImKHSlbeRBKAIUbABFLnHdANQ0fCj2P6s3gZcu9MWaNw5HQKWkxRUM
bRpRXZTkF4MBW9D0Nn8XkUdsz4d8p/WiZXKVy/5FjRUrF2ZAGFTVxy80hONyHHArJUDAd8UXWVbF
KCsmjb9rydbsPCfhmOVQmrbqtVu7BzO9xXmjAMri2/zc5l8+IJTHtR1iBOO0BsuSPDK36IJwwFaE
Rinbr5lHc0ynNUYRM9S+YXNQ0OpXIEcGsVh6qL4qyrPv5gWDm8YjInOiKn8TqO5NZE7n1rcFTrKH
JFkFUiv36wSNfQdf2aJ2e57JKWq050SAejXxY02NtfLiebXySMtcZbx2aHRTs0RUnbpQqGtpxJDa
djbfhOTkt185KkzpAc4gAhwQqWzi1INYkUqQYUr8inCpLJINCiagqu/j0B/SfXf+3wdbYM5DrVX5
UZOlFJNFY+CJvvOnFEn0y+5zNXw8D6O4mEusdO1ki9uLdqhOa5niNqoAAY6d6XhRQP8uOdwvayqD
gIKbYo/qU2Ztb/CfgVSMrXrrd5NyLavDjYE7+WB2heXPAN5gZk0792HBguiDbiKuMHRfnryke2lA
VknZyAovu0DTgzCwWPcao8jh8/KQcBIKCAbvU5KuEhcXJeGdaGZeHCpNbXHyMplEArFK/mm54RP9
45A8NLi0BuinUG3zIRLNiqZVUuvZdiP3imlgnpwCDCXwiyVERdyeRZd2iUYtnkvv9T434LZs8Jj/
wJls4siV8BOAn7ifOTY3hg0/1PAxH4TKDWwwkL+oIbWUExa99GFFpPUPBBqMHJrwr7LJKM1UL5VN
yFFMssZcoiAHWmyuhmkkHHOcmO3p/1F0CdB75hZOZD8OOGMPUvt9+fxMYjsZmfkaRzPHgH2CiPq7
+kphLYwO+BTg2BqBaXH6WFrubVjjAC1iVayNNfxkycsR6+Xv0Wj4jvJsxa87rMVr09VvSEP/ZNbB
HuDCbjPwJSsOcKT7E1GeVz9UIRrH00i1uILFTo9LLPGtBV6shi6LG6obUJS+TnJAM4R9GRG3WA61
AtYLKz5UqCUSEDpc4KjBZpa7BM8we0JjlLMSk17oP6yPXsoNeG3UK8WbHZL6qf2KK7iaauXt1T7i
IMMLu+eijPCjGc5VhIlPr5I8stKMbC7CX5sKfppwzAw7itczvAzmZPyqZ5Rmc2L6Lg+MtykHK+Hs
HVBia2EOTC03CvCyCQdZQZsfTiPEA9tsIwSGJGDGnKO2G2kJLlPrxIXBjAPwkn31+TiqEPsveY0x
2KmNAy/UES7pJVFSuc5UvBfYMfDUCtl2WrvYUNTxOOTtLre3PGYe3mTwdXNBrWjm0kBTO93RIIb7
OojZNxA7zx2fUXRPYO4RdAvvwKrPY8BwI7pwzRy1yfwr6Sxi3kzS/ngraWTr7r/6fcmWac4iSSJ+
v0OHjYlPSyosGctaRPgpNgAlXoH+StjENGdXGa0R9snJw18xsoR8P4ea9kMSjxYcxuF4M44HQvgH
5rb68gavju8YEcSv4Xlku59TDoyfr0SDnRioWEIJYzJUqK/kimpZdFpXeU8vbIINg2rqsNvxYksr
xGl0aCDQTN6RlGKdV94r+xLi8UagYt+xxKhvC0WXlE+F3UcV3/02q9f4XL/wVQ/SL7LbMAhEqAau
xL2zAtyBiZKYOew41ci5/Ju59ppnaC2Dmnao00Di5MOFyihNhBNWxLq3XftljKeOlOwCz7OoMlFP
e8TQmPKxpMap/wgvKmbAar2w/zYzEBHkh2EAM2z44RmUgLAn08VV6Lhrh2EK2q0Ka6SIU5TiRSTS
VjCm3viwrM7TzG0icUeMZeZB7jHKelMdGbsJsIeIeR8IgR90lpeCT30u3KWzpxjMejXiGkMFynPr
NvV933XzxQaMRuInzcBTbWSfpvt8BLE5mIqLPV+8G95QWjVSZWx+AEOTxZlAARA2W+VUgvxlLM0f
bsUsOApAQSEvkVHzzHWgJNrLoSFa/eog10OJj7WfAUmh3h/hE/Z+oCMmvE1IqRreinkpm1giZG16
eUaP0bpkCtbze9Fd3uUst7sJx1PPCHprUL0gUia9N6cnC7gdAB/bPtGhO/ZhxPh2oCx94T/Pj03u
FEbI1LxbT62BIaYHusKDAfGG+7r6DcfD/VBPzaL4AE1JKhb58YQ5NNR4LZ+C42xAXBqYP/bkzwrl
hQBcAhY/f/I59DBhxrts+kLUE/gfGriVSZc4Jw/5YyS8xXbm84b2ptaeAC7NhTw+iEw24EQ9qAus
F+JwEf9TRuc4Z+W/Qt57EjyGlBGRUAA5sE8WkIqx/gowl5WtqwTgKcGKtzzIbAb+qa4XymsaN3BD
KJUGIN1d317z8EuFdomAHIbHO3qILpfM3nMZhOKXhgHJq61azbHsYL/SeTBmHFQ8qXc84ytBIqOL
S7THnTUlcKGFi+Fx3HrlWtSh4yGY8oYDVBhAEMMhVm6rdECmBmsWp6yGBn92v2NG+kz2MoSb1Oem
Z/nFal/c9gahE73HZDmPSkdqk7qfbNPUVR3Zr2iFXSn/7ewrv8Kp9OLod6DeZvpk2C46jbxwRvXB
EZPklY5tRWvUhsIYCfAIOOiGdzYIg4bygeVthF70soteNvCV0f8caIMJKZch8aWOHO3chJA4nJrj
ib+64ikyKXp+RCCs7qdNQfYLjXPPCei3VLbEJdN4W4fP2y6SvAdnzqLUTpKhUEz1mG2cmYqreatU
4yQXDAB5aykH27LDB6Qi9ubG3zselVFkPg8kWQW9QzO6sPwnE8YWox4QtbqOaSZbKe6Waz4GlVrL
m1OI34IQpHKC69+F4IhV3oRwzgG4qK2OFLxcNoOAQzawUHeZJJqKkGdHu7o8TCIyu8CkfjCFYUu/
Jkw7wpc4s2Qlh2wGBQCYNUshug0rQnnXIteXmRUHWjG0aUYEIAa70zSyeUU0CvAkjIX7R8/up2p9
1Z19ws6MfeJukEx9Ot1g7wlR/zad7JSvfXpTT3ldyYoaSqHJw/fvZ+SuL8r7bFm3a58A+PSMK/7p
RN2lSZL3C+qt9O/rXQw9avTghMFs7wGYdZ2LGhN905EnGGmBeGl4bz8MQRYcZbvVxSAST3ixYinT
vo4dxctmZ5gLMFcoy19aHouxumRE/B47wJGCmupMxgZLJOPjU5jtWBuwxG39iuA9DehPNtQZXieP
w93YpRamZX7d6uqZIWS4SHqw6aEHZQZ4ZwNpaTXDpkRZ5Nr6VY7wHeGw6U5W+snmQ8dPgVnTrz5H
uFCqrxod+86G9ZKdBraExiu6W/2B65fGGSSUYxNu2ekvztDt6ApO6WsQDKXPDBz4E5CNpiE3ZxKI
IRWuFbW4e/1wjXbDcRfUnaggFBBm7vvXck/RGWtGM4YNhQrb27FpOU57RYxmODjrjjPQ02T8s28V
4VJOOmzWsQai8lj8lpuSiUnWwNb9wn68nKvaq+UkJnlio+VM9uF/Cn1aCWUW7zyZBYB9W8S02oTG
ztpwLSXRvWzc2lg2fzJu70ur+GLDdPEU5Tfuew/Cz6tenKbigg9K+3EV9DdhhycPxnbXkKCpbO7K
FvKhG18ZLQiCEdauxyDUl6NO2feUA+JVLoQHuUIdhnUFcdwQ2XNfs0sqJVRgjJRMLvwklQkWejgx
9yS0CUmlmQMv+8fZn7uF37TV+PFlAOeecqocID9msDGNDDlrqol0DValo8ksVOq2kHDB+aqQWv4s
W4Xd8r1mg/Sy3zC0XV9pmGvRK1mCxs+IBxtseHVzPZft2QSO1ty4jTjncUPel7CRdM94h49TUCht
9YFNrcQ/uA9fUJ/t2Gh5bNBVjPw0Pt76ap98Ov14EYz94HsmlglOYGXGMeIxgJV4WCkHrd7e7Kiw
M6UtsMtKLDTIkkgEZJA/yvB4hjPP1eB+AV94JWQ5yMek+/cTG5QN6lu0TalVO4RT4rq5BLu2WlSj
Ifam45qGCOQsyqRNOWgIdx8vZlrwZgCvB02yI89KjyYolQUy7jXLZKp3sRnHsig+SwNnFv8MvQVX
bgKBjTXLMGxuIkgUUSgHOGGL0ic0lhgb65huzeKNczixx503B++oYA6XIyBEMcO78kqdn7H54Hac
lzVYg2kbBis2du5lsFeO+mqkigHY4Q4wYbdBZfWtu6tV2a8X5SGcVj6mwlEED3AxSrxuII+UehxN
gCMMrEqXokLGwyEuXCwjjVCRSOltPTDoghRRXlv/0oJ421+KtI70jhkx2Fd1gF6Ib6Oee1xJ6igk
CJyFs5LFRgmu3JandSrW3yRP3tMI3Te/LSArxCmmq4jqfFi+wJLnqqLDE8EwO6MvVE6rotYIpc16
m3fi/vIY5b5oks1LGLsCWOtGSeuq35FUz3mNqScWoB9PN6sirOS3vWUjbCKkgOs6kyKoIXB5Jo4z
n4/il74Pru3mGkSw9/gCwhH6Ngwh6Uqo8aWk+npsBDzr+timO35dFYe0geQuwHaNMXCV1aQzqBUU
PXg2Xri1HGThNQv3OsRNxMP9TW3vGiWkijg/ndhPyUaTukaLL++L0oXXlFrETG8G+z7sCZ2YW6cT
S62KPZ48IKR2PYhTwIvObj2oaB2Drt6Xs/pSQunEBLhdM5H4sL89lhkAUm7AYTO99XWvd2U7C/jw
pNAjWrHfG+z0eXhiTQMsowtO2gsars4aShopjVxXRB8DO1B8i85/XndX6LbuKoOPKLLz/NiW85NJ
Uykb+CNe1iJQc1lCKIy5pA6bAFRY7OKl1HbCVWdEE2dF/7cV+cWEYaJxooWhbFwEWjLPnP1sAzIq
LMP2biB+WaNx0vhpGmQV7KgBjEqXLV4YEOel5aTjJ4JixH3Pr3yreYyxu7dN6DMwARaB37N0x3A4
RalqI34xtSiV31ZBmswrEvx1XXgkgv8Ayd6JFGmM/jDUEntEsVG0JsyAaf2OYx4lyn2q8YMdSfiQ
iODdXYgmEjbsfDxrQTab8adCNmovfTqHN/f0+Lw+5IYEqyX6tnNzmSDTX+Y+xA1k0AAxwdcIjzIS
c3uErO8grZBt5xf3GDiKfgAb/OU6HY/Rgx4t47nYLbAeqifs7TH/E1leNXUyDbOIpj7DuZkQEPXs
LAzx0x0ygKTX7wmd2u0opRz8iwH2Z2U49CPnyEdOV5BsxvAlLqPJMkpEPtb5Tsa4VcK6LC5DXzKh
m7Fe4LEifYUqmM1C8ppv7l+2NstLJaBF7QkpaLGGUBukO89abhztpnP0FYx4LcfDFmsrTC/69dJs
0qFw0EP88ecaXOjw0rQcOtQxvBImvROp3lblJzKyJsnKNc4mcj3U88z4XiJwFT056PCIjC2kxRkQ
WPDRPwkllbdBMXIELU33W2GSbbcRRAZdgBvUlRx/j78OdLnC2YrDxIJ0m4wP/fIbff+xApuoH7np
a4lj047CXs6LJD+kYn9ySnj4XHSVxvSYEdVwE0fcAomG6H29Ia/U7CM109+ST5ZCtbI49pXWWja3
8aqYJX1YwJs4BsNqTjN9Lty6rEQ5CK9Qgwbuqm4eQHxobJYdemLcmuE2VMRp7XaIBkjrpxDnh6zy
9zXqp0LCU3VM4tkMAgUegDc5bUgEcDpdhL4N2hC25Sy+FuiUHuVukEYk/fdMzG/jbrNCs1t9Da9d
bcZQT3POwvob+CGjQ+B3JSn6VsxX9o7gniJznbkWTF5ZEY4+eifT053t13zqu67zeakhJ5Uh0Nzt
JnJoLIr98+qXd90hfS8JbjKSIuqL6AcwQBSgI6Y6rmmrdYb/z9KjAHpgEWU4CN14u6NQJNHNchRS
x2YS4WgketfVT0a+Oy9lAztWWWdxY2cLRQj/eQH3JqsV4vf2C12xwh0N3EAOnc5x8k2KCcU2Wbpq
n3BVfz4nPBJXaQqtHLdYsYyxze/K1JJUIwPwaccxC5nxQwYOr4smS6qU21lQeX39WIwOtSrWSIvE
MaxhnSixwHTtOjuj/w/hIV/hNXZbbki9Bh+VgMjojdxiv+mZdQvMTZFmHpKCneH2QrsyeBlQSua6
bbjaAVS1Y5k7Wqu4IAQuoVvuRQqaIfIyU0lf4is/xkwRHNAc4MhZJBxQ/tlZrQZ1UCXzsk3h2h90
BDpMkWW3cpCs3/YfIOfxXf3zv3HnlZ9Af7WpMkTRyU0USv1GKs0A1dF40ttGi0mvir0Vor+onsU9
hYiKLQcturnK06Jyjr5wH2pI7qngk/Zig98wlnxsvwuGjp9aqVJQP2aj1JCt9oheETGg7RWVEov+
FK5mMEdG27H2i0TUfctqu+rUIT0UIVzgxCSaCBl3+W4KDkr03TIiVdGpA7Yyw7Pm0nZeSiGmVOFT
dC3327n9O2hDHxXxbno1usB9diGbCc+xtEkf0fc1EspT/AZXbcxiqGJFEmlO0yrIhHO7EbGjLlJB
oYmUQDXyik/km6YN7MKtZQYb9Yb1CHT3rBhzhE+uEkmFBtD7OBDlHEHXHR2z4B5fNZGjaVPzihl3
AQ4rNPjVteO46W/L9Ut/dFnkS1dGV9Mho/gzLnZe9UX3jvfs5oTGZCNSNjeDKwMhS5S530rIyGut
JAgobspN8KUnyBkPYmLFJ0twSqGClCc5oFJuD39nlnFZguPktNcjQM1L23EX+//+sIlFOSicA8vm
QPfsoERtNgPACCLv0JGRSlpDqglVhEnXwAZsSpwtBMZnQH0LZMeEZ/S+PnkWZYxhcc6MRWjJHAWg
WrIwLfCgToy81IRBmy8Ffl+lhLrKxviMXuUj7RzvhBmWlAALLs8twXdfuZsiXlnWaJKup0J0ELxx
ZOvJXWLYFsgx2vAhPQ0gRwgeSejMNyi9lcU0TEl7YDaiUZz8wSrQ7zi7I8R2ecN71dBrUSTknBCE
SHPGzIDW+1Nn4LBtWKrWLw6euAt/dU2bSCvIO8ods/gkI++8Fo0H2nIE9nD3cHZw0NjHVN/YMThq
WCGPX7ZEEeyN29aRahHHae6ziBlm9CNSMGxyZAs4z6SWmG0ceI6MM8QUEJq4hAI5GhnzYKGUIhV6
l8VbT9nX7oh0z/nPrlYMFaWUSprE40cBWfA/Mwvktybwk0xqFE9p1LykR2tJ6Pe/jAkzV0Q57mTZ
N+BB3+8PLj1EX7qhUaOSjeU1dwVdkR4lleTTAztwUqkBdnz/3ODS8PQAxWVfcARVdXC5bgguJrpK
99nruHiQoBaqDA8q/bSYcemLg10PvV13rlj1FgCO+9tZQYqrSkDx/1kXu+fEXdDb6yS8qQCWOBD/
dq0CoKfbhErkJdLfvNdOZB5XO2VuZg3M/g8NoT9qL0qFClGStaVDYne7iyFirOS5dvMAJWh2fatm
HgjusKxilUF2SwOtMMBDJ1fc9S73hmhoABh2kCD8dPMJFW+B0kV53gcF+a7ikw/KOch6cgKAoiUM
/VFp7WIjYWxdBN3HDChrpI0UC9oseoiqiBXo5ZSISIsfJnfl2N6KZ4KYrFcn7oPZI0CwYWiYyuRW
Q6J9AAzODRqo+xjVWZH89URD/BGabSJCRwL8vk0qyCcftCVzEhDzBeY79DrTej5Me8g+T9725/AY
nnVjT0v8br5YBdIAlGjqca+muyX96rjUpzgrGwRsVKhcIylfjUEqysDcD/Hc/ZDtNM4A/8zhqV+p
MYuRTqKZEoJ3bj9533fWwb4fa70bLTiWrEAZ+Qeq/IkQlOpPa1qiG+2Q+bl2kVpyR7+9dMWqWetW
hXX6JoXK3OANXf4hGZzp3BgFvkq9FHI9lerWOPdctZoUJm1II7N3Z8GTwoa1/1O0f5eokLxYsphQ
51timbFhygIWxbMePTFLt7yONvyfyb1cqBlt18kj7CqOXLNxUQZkpfOXSmVhkJBd2rDcpa6iTyOU
4e7bBQSJjqOVz7pVpkeD/56379WPkCzP9ufOiDNp7R7JeMvfPtXTtiDfrbOvoYs/MfZRb81w3WJH
xX+ospYhCECUZyodVwl0rJfIbpo26T6JBhNMDlBP8SQkIJB33wF916/TnoOExKakJnOC/dXL0Sy0
mPrU+7amU7z7vqOqJn5pl6Li0pvpcNRxgLL5cfsBJcFzapXgUtGqwUiEGX0xnPeSmU5Zi5PJ71a5
S8bH/Dow/sCWQJ/o95BQHVdXErgRXCg3q7d7kf08rRpdgd39+Qcho3hhA1Xj1Y9v56KoXqc2wZVs
8aQoHdrTN3KhWOeA6Xfm4j6ep+IuP2b/wBeoaQY36dpoTg7QbaYSrQ1nQn/NDiQMI7XDoOhIq2ls
/AK2eQ9vzTzXJn0J6k7ZP5szScytTZiWDlC3rKaHmYa5PqNqQafxOSHDpu3xt/5thjD3GS1NPUTI
5UomrIoiGx88dVERxLdtjxUIBz8tO5jTbr9CEfnboBLg+epWSRvl4yjIDzWIovnFbAMYozT5v4n2
5FtSI/BtODI61iVPSC757Y6sGZiGE4gOeUjMGSuL2YmdtsWA2aInEPuOs39zx2UqZl7Gq/ovAwMj
2mnUoPdF9LL7NSlhJY1ZZRZiSeI+tEP1rT7eWnL/q2zB1QepkZLriQooQv790jd+aofX2dqktQRU
NUOx+2OGWxNeKiQoTJuxvzbbUbyxiMpIjXuXQoCz9dwjYqVjm2d6naYMuaokvnw80VMCMpjGIwbf
oKUY5hoXjT81N66ug0ly8RStBKDH5Yflk3VzE2Ik17BZC8+Ges4MpRZGPguNTRfWez0K10wnEezJ
TQAsakkO8HlJMYIXN35+ukkgzrmn2paeBE3W7IlC0cIBuKFXnDQoPUeZn99fZQhdnolFcTdmOBQb
oZX8zO2SLnV02RtEHSRRNQmpKzpqgiqsFj4ju38zFhDB93RmK7NaQ3Z8KWxZWJxqUg6S8iAsWAbt
a1ORpzbmrnH977w1MefCB3ObXolthJaK4J+MDSqyVXqUcYAkiIFqaSTUATgweeb51tTvyZ1KFuzj
OKq5mn2/u7Nm2yn2yVf1tPLg6WKSrKO5cpzigJMFGoq6A03BPH3gytc+xMNjtizcFphthp0Jn1Id
bRExod9+W7hNrvFQUFXBeMj85IiIH8QNGJj+QRVNNnEAh2LuX5eluC564QnFu9ZHFJhKyMsj+MP2
bX9pH/7E9fiu/58yst2hM1qb+GRF5xJh22uJKCAGGk+tD+SPbzO6AyEN8HLS/12gOphV3KKKuAlI
vcyoNgunvM668pBgLyfxu/WWah6/FjDJ1iwBtP9VbHh1FRDlJZ7Js3mYi9RHRnj3fDtQmxNiSbhY
2NEsMIBoYa5ru2dgeA/WQ58DN/tgQbyV7MlROAHKuu+txlxN1eywe0F3R5o8nnIc7ubQY1bcMGo7
bIQwnDYXyEmtuPKuiYnKhx7dXnkwqKXnNQ2TTpuss6GmjwN2L6U5wkrOPiaTs1XdzdVbBN7XMqzq
LsZ44coGavS/QAnEyEdp05w8w2EHPs1bjprx1f5w1C56tOKLWpy0i5yppVEmBRI1amBLZEkkfqFW
xLx03Kh9gIXstbwZy+CAE9uTHmPEOaGQ2kSoVIKt0HYXIQGamvcU94s2BPIZ36XKsIlw9jydlwgv
G+YT3zOUp4u+psOwRHe6ZYl5NEeybR99a8NLSHyb4rCmezsKjlcPBa0gjAAKQ/sFVYrcQSqfJuLt
asPs4sw9f3iPmcO4yDon58jVduMrGhDwBF8KNi7KwFliCbXLfjDGZzt9w2kxT5Xtx4FA7fb6aA4x
P94iHzV0mPyFIrdm733seludpOopPX8igLy6y5R/N5jEDPlbQKOSIhPHuNdCiycwZs/7U7b2UjT6
JK7LYPW5yLDfzeV54Nl1b8h1mY524SkYyPKC3O6WgIBj+dnS/ikDSEJCTwtHz5KEQCffb893URzD
5RLtpkXczD77FgJZqkzvY76sks+cEncllUSWrfzko1Sa3J7eQ/HP3lhINyJ3y5E+r4zVAEPiPiRp
SoX8AfIzkfv2a7Gj7kNYM7nn7XCd4cellrLtbwkgXCsA8CGMTJHXlijYjKMsZ+BkrhF3t+kdHfV8
qEE6SDG2lwZ/JI7JRj148kwghkL909dY303OsUiSa8EaZL8fVhOkDuDItzKknC5mEuq9j3jtuM/C
JqwXZANLWhVH2nIprFfnyLzBVLCCxOIA2g3U0bUe0mTQFidJai+6oKF4u5i4tefEFpDsZNwOTHV7
zkWuRir1u/H8cz+aT9z7/sZ/7bJXyRJUwdlbnjzlNzNFo33XcV/3rzLt8/4Fnv7gt9/iNl9qReQz
Lp+sLeNy9prb9M4/URmExKgrfjrQr6wCaV8Cv+XFYqJHO9SvNqKKj7USNtYcPBg2rrfN60GNEW/Q
6IX1FoMr0NCwfm9GnmfR0EldMfz4ueQjVYsXY7H61cKlc/AK5VpHevR/bASzXm5s1BLuOde9Oqwv
NJUc24h+llOBYv+eQV17O3I4yJ9cCruBn1KqkGvSlcm2rrA8FjEzItEis0FN1gUikKan55M/oIpV
iomQ1OlEa322QcXdoswbJDjeOPs0vGzyBjfBIMDwSx293bs0DSTmmI/9zJTSMSQ1ghlD0qHk8EBh
E0fGddzfOgTX1TulhCVQcGeiDR1rMnjFi1WJKxZa90cBI48d0546GLaT/8HQa8amSyedTHSYn8CS
/jyqpTPOYtD/LFO56Nf/rbjRD7QjAWKaSk07QUIVK6AQ+U1VP4UKJtQdgXDHJfAbtDNgIfMvf9xP
bsrwG2ucrP93RRI4BwtfsMBcf4Z8Xni/UjwOHDZFkMjZop5MKMrXkhBN/LoU3OKbigeCQb8OVIzv
ldu4FWRrPo12F0hCqyMUCtMUTnmDIojZG8qkBL/JgJRgyZC1L0yo3438ArxjP1RdK53nzo+/CS0t
2yT/vc6tI0ogdVQS8CGbQ3BhtiTNWwxdPEE7O4qCJ1jy75wrtDHjuTxczTc0sUXfpa41IH4SovRo
5IoPdPI9n8+GkPxBnpVn9HKORfq994yNTNMTwHm41gH5flG90U4BiY5hPBtBxIfWA+VJXU/4wNQG
rhGwg356+zkfMySjajAZGDlv+7G+CiAmpb+oF7eW+zd34Pnhr5zcFfOCUmlraisWlU8S7GQyQc3l
JGuvlWldATAbBt8HVjSnKYNPNbtntLWVChzfDrJhb4AR5SqWhdZJCMIVBH6P4iA8pjbkXx89nEsW
KiUtH12aFtRRmhQqIPRbw7h/XilPh9u9M2V2VouX2VVjTA3Qj6U4DpuVK0hwSom+qOgynmP5uJcr
5sFP/2s2lFv4ppHGQE8/H826yEkII2ExK9DKnS4fy4sOe9SP7Y/6e16rIOThwqRIZxCLXfygBs5Z
gBPn8b1VAUlGAIc0BAi4G5ZfCLp3dJCV4PVAiqzKcU1jzaJitKVQBufe9DBblCmxRTsCbmQ8spo6
1AIR66796G4M+ranr9rzTbTrmwjRQHizJXLNBMiRfnRIdvgw5DpLMR/wAkiTfJ2JC3VmGlmKReoJ
nCMWnbA4v+tYGDDD4JJ13VPUSMHwmR7GJfYcvuj6W1TKvhx3jdzciNAeGsf11Weosb5pI8e1m6z5
ol1BsMXmwKYRUlF0DfyDW6M0UCmDTAR75EeF6DPchOzj/1nHGEkDGWqoqf7rAgmdOwRSCW42Skzc
MAOQWTk1BzLmlxGxagW2tE0vmrV9VyoV6dbVV7paYuqvsYLHViQQvntwmqCfa2fZS8XyHAZtSY9H
RtuLG58ZvZdT63lUbRM1lNAU6tkZaWSesXb2bk18pFaEKTLs8uXPOe8DGGNAhkJDs2K6Tq1Q719T
pp+L6UbK+OTu5g7/5ny1ZzOpLqu0FANgdGqzeLB1X534lK9lPdI626QLv+urfE1g7tyGuh21z5bB
wrlqcdKMhZknKdokw7GhMooSQcGebjrvTKMlXNnHmfu7fOqvaidM1K+g8dk8qZ5RG49oct/6OH5s
ibh2YRCJ6vJshNp1OWAIhK9TedCDJvFM9NjQnKVgjsau659SRJzxb2mLay7iNCFrgT4/2S8Kzmvh
RrYVVIW2j33aRpOxcr/nkW/ubwNTKwRbZB/xU+bGsKw7s71iFwleTIR8usXQRKx6QGS+H9PzGdN7
LYsalJfIS3m4OA29cEzvIPXtJu7XvpwuAGZpY0OEqfO0rOFRx/+oGUf+eX17Ayv15vlQIsXL9y3G
jcq4odQLHj+4dB84bmelJYNe1AwuOnVRW8tnfLXSwzsHESLuqVMnN4fnwANmkKpAcosj5u6ZFAvo
f2C8DbV3m2itMIcooKUd3xNg52Ips7RIabxV7MimM6TBGMpLGOe8CPbwnFMMc6SK6oVm73XI86NT
UsCfit8/A2veNDQhxNwNzDS+fzeUWrAKSQOZIUOHSHGt9nxKqGUUb+kEZgw6yb1asgnmN/f23hwu
22J+GkbZMN7FImJj59kuENppuDqe8nNvEhOy+2W0T/bvOpebhMLUAOxw8iQEbOWB9njDATrbSv/I
O7AG9oQi/65lIQNQyCSVrMx7OAj/XA5kZAXf8jrFem7lmf+sn9F9MCHFd9M+gds8JSN8il7QFHq5
Wzgypz7Hm7QptrSH7qJ2M/ldcNW24kcqM1sCoa+F3/aBr7g9U5SZoU72UxyZUskrimFAOdCrdmJk
UpfxQd9C9LwA/mkpVomQPLft+8UJKBmV5LX9EWzB/5aDHkUwvE1kfGF+NLxOmNEiRGAUd9M7oUu/
h+AFToI6fQz6i1DTcVPLxp18z1xZsVSMqtmOLdJ2/HNzsEsKXNzMBZU0hkvtM0Jwd1dmMY5x8ulh
WAdcwDHiCL+0OKobHGMysomYUeCT70rjFcvReMFvMd477jWd1vQaCrEsj/xGR0pqwtqdG1kj12TX
5zTnxaXQ9m3h5lqo92WKK0CjN98mMWPelVrec1HRVhljPkjFTl/uRKORTxSUOV4JwvZ2UsBaIPg0
YcR+5ImSepoD2mL3bPgnM1SGvLW9TaPP0N16CUhlzYUuGoYY39Li9z40q+dnT8ecl2oRQ8NKCOhk
ECAKRGBWWg2O7BgAt5MXzo3c3pqQ4lfLKVXVWqWcW53T5KGsbTPse9tJSDEDPz5pIk/Ae0lD7HsX
WHXuaWD5s2s8pk61Tp8v+OqlfjT/9cC4RstDIMpWKmdii+T6W4hMzDtv5t9a2PpywLYDiqJP+u97
C9x/2vbxX638o9I8T50dG2EjuTw2/bz4RiSJLFbMG6MbUo+liu3cYFHnU/pkuOK51k1X5PdHQMcS
4YPoTnqJk/Y7sRA3kW29u5MT3I3jeAnB38VxYJ32XA4RTPofyFjBIyUD8BzQ+MKQJAy0IpHT6SWb
WQbkthj4DCHiWzUyQpN5RGZ2iuuQPs6QDslojaBKEG74UmKsbwhDQ4sAwkMtuOfQmlMJUNklUHdd
+4OKcCB6HvT29ARJRQ3JFgYvnAGR+w3rgPwTnpBbwIhJtucvZKPVA6B0SpMrUypoPBFMAfKtCIi0
kiQ3aPWRczv0p9jlw3qmb/0J9lHayFQluv6jx7fq7VZGAvohcVMWpq/F6aygCAsvgp7KDFYIWa2E
1AKbosoghu0JERaNR7ibmzcOZ2TEox2ZSclhFP21iaGT0G0Pk4BnD669X+OQszrAPL1v98Ifvy1H
tpfYklv4jxlF1q5mVnrQAZLD0jRuCRPKlmcK6LQm6gKdZGFeysWnonaqGU/B97YY4OOzM7wRSf3F
oQKpVR5e+0SpY43boer+JR+z9y4hhfkfwvZ2/AaVE6eVPJL/gcg+l/OUov91P8kTuk3oHYtLUiyb
SsOXuAY5LbCxbhWUFX9oACyCfVhp9KdinVsBmHvuHhC5dgF/LWRCmsRXrInKIYI4ObXNVdNPq1cq
mPYfR5GNi6jBi3ca1DU2o35CPwwpzRzwVlMH0tneHrIKikfM1Bd0JK5/Yu4blBb/WVOGcureYZB4
FjCu439JVquWDvHFWOJ5sG0hY+qxjdrUXCwEJ+BnmvQ4+ENeXaIlNnH5aKA9qMBRxskSgzNBtALZ
QeCR9uNKWuoHO0wvYBNWk8JzfeUPDSTr2f6UENE8CG4BHaWGM9Gyg3F0+0L6cWufFsDIG+sK1A4j
p5vIrmWEN1bZPmlFvyEMKUvx5N7P/36oDjLiyVwIEDZTj2Qp0WxC/muGtFoT+c27kpVhqsAid901
JwsHG5tB89RnRRX6nWEcdYLT2d1ItJ/jgKCFRUKgB/pKWaFTm+voj12Cz9GRNVlwnZ8MzRfnk61v
jR1lPa8n1ZuTFYUvKjlX161Zxd3bGzW9LIvRpF5x0jT3q7ga1wQ3axCdrBenr6RkMcb2WuFs86m8
lmaV0nXjPsRJrrPTh4bf26IuXHrygYadRLSmCBglO7DHZUxQfHteTRZdim7RK86ySfLOnGNHusua
wLxnS4E4OP/AjJkvq9YH0Yb1a3cWYSQicnOR7F/v9TKdeZCXPgPpXW3IPuztcZAUrNXdiK1DMZJj
tIIS39e6CSbsF9l1dimLwCNmeabSvi0syLMMZ49pg7fCwJv4YRrpHlNYO1mTGKvZNPQN6Y4qeAGa
5JHZz78FdZl+8POLeniTdrv9hvLodwXQSn5YJ1U33pU0paZWoTSrcsipNS1Yw7/6dpdaIAoKITk5
phI4hvP+ypXFXQfvYVp3lIl4kGBmLfLtR6r98CX69mjA5KhFXuqswXUSwF6tPeaJwQ3POOQIJHML
0rJiek/+MQNtFzCQ2ipfxntYvqsbS5zt4RCVC6xaxpQ2ES6CuF8ki0x+fkg34AsXigoFGBzfsK7V
DDj2/Sfv8gJ44KvpHkP90PxG3Dkzf8SgYWJ8T7Km/UvRq2tXGS6JHoev79aOfV9V7H67LGNv7XIs
Xtrcha2GoWHaejfg+sZG1VU5yVcfAUR5zypcQyQENjIlQg8FOk4OyBEZiLn0zFjAZUir37D1ooV0
y4eTy1Cemxz+E63GDG+caHIFa66OvitGKDe5kbs2zuYtm/3D3nTcvXTE04QvkOZyHApiU7Utp52E
7ody9esPUc+XAizGHksn+CiwflSmsS1Cq6rSvMxiLhV1iDZtkKUcn6v5S+WXjAGvfXOfHbggLDaO
eTyunoqpWG847w+YwNb890ywZEWFtdxReUtRjfETFSRBqm8IXGi19K6mvvjrTlpYmsS95zkai6dY
myfvB66PEA2gr2wLQt2CoKp42C/JOmB3m7AfzhF8tv3cAYgiVrgBhq14lYe5JzJyz4jwbZyVn9ae
ci9ERiZioqLorMRB+GB44mOBNoZU86sroLglCSMoN6Q+hCQa2BuRuvDxbHJU2y9xP/KCjRx1Qy8l
QmKGJs/ZLu/lcI6IJhd5ACIDGW+VpU7UpKQbhctuFx3rygew5LpbEVBOHppN7QkgE+/63fW2N3Gx
lgP6399RuFLktivvTG7z3xN/vopIgvGUhLXv4LlXnZjRTrmISbMSbI0qvxkrmDSIpGif/N5W/5R9
XwsbDomc6uJK81PFkQwXeGxV1bwHG++NjIKFXSC0X60HwHv7F5p8ur5AfLfNx1jFxqVkzXTBDw7S
C9LBu82taAVsEKqunQndKFOrrK3Oc9hXejZ+hRCX+seXDA5gQifzFJXXnZ1Yu5+vjv7GRh594Luh
3oDGu+njBIyTbjlUTsa/yqkIfh5m/aBQoYIpHrdeMVqJm1NtSV7QeQr5ue4gD/gLvc1P2/BFQnU4
9DBKZgUBufgJ6KQVmoL4Hyu+O77m76uzqC3/n+ygX1/bYhePdBcE1+thgAgIYMFuXJEU0Y9sHjnr
/EcxibFxGNtbRercz/3QQqGp3I8EO4SO1Wk69TiNv+8LVujecj9c27a86x8Inor+YXWXvO61Jjwg
UkcrhqqmB6e9NPTJUcHYCn8Ad+Jz8rp9mb2QnW1/xU0jyEBMY2Q2/jzS+1dbYkT+MgN8GHeIPRN9
yC4ZuGAPBssQF8NFPOH/GGAu3Ixgm19J0vi0de5he+1zKIhHXuVLR4kT1ue7+Zj2WUSX1DMwq51S
PPn9ATx18OG7PqGVn+OP6IJMJzEyHKxjDpil7xvgMFo2cb4vmv1LMv2rh+vIaQRw6TeO2FexsPq8
f4JqqfJxcwi3hY48fc1DDSBmcC9rv9FK5AKZG5tjEu04xUPvYOodnNgibjDXHPNF8jes5X+BvKyC
il3JqaYdU3y75WunJt8WpbMfcUMqET/HIUBLwocNtsUSoYvb4wD4BPnCCswvY/74JZdyzGL9dggu
VxQtjiuvELNRsTtZVGCE8zpzbPe1Lynh7k/SMD/dTwj6+DpjakSMBCbOEzFS+8fWEg6AxmJ4sTjJ
CPpxeQCONf5qYVlDQajyINCP8yFXGWv1bz/WvijN5zoOejMWg0VcBp/C+MoGOv0xiDxo0ZwBe57k
szr1OJpk9ZGsnouH5YuvW8nktp7maFzASPAA6SdeGnQ2lymsppLUqVuNbMjaGC555rcaVc/537nB
bUo0oYka4GKbliXJokoLDANt5SbnArr+gH7eqO2GpPsoU8nsafJBt4iIOpI2ZSO2yitCCinmTH4p
/5hM07mcO+PipwS7JRQzRfc8Qm1vlOygJ9h8qtXW4YwnYKvsee67h6H7xeQSJBQguNTdBxw8yjCt
HaKIK9+Qt3D8QVU8dqpEMWE5+dwh7ODkyqd+1QgItuz7MM+1xe4HNK6l8lW5olfuJ/0mIC646Iys
45DmR3YYGbFpoB5Yh5AScQLptIAWexjtz2hSIJ+Ns1DPfObEbpSdJ4KGk/Az/LvZwYRhJ9+jAl5w
B2EvbfIhin0syEqyVcYGS/Zu6lqlEc0bXzDre98008Ho3N0+U/ACDf7WhBDKHvb6ie1lXV9dAd/O
j9KbNvnTX0cytwUk/QT/9MFUdnwWuMq8Chz8+7Y3Xz3mp+eySNP5w+OGSB82+W7eM5QiUbzkzvWN
5iQrzQEV5mClXMJwuEqje+u1Q36dgvUmyAPdS+hvNw5hdBD0Hb1y5zb7baXZrQlI6iZOAfp7jtfn
ywurHJM5nTe1lV4PWqsnsIRauBL71tdgI3WiNSyR4J5kr1TO6NtMTW/e14mWZPXruH21HtmLUG1q
w5M4fQgZW5aMzwAJhCIXBYZQXSn0QS7r6N0F+43IDR5XJZtTAraGuegnD1tGmwf9/pgsLQpralBt
hkdEA45wCn5e11t4FjlCbPdb2hF+vlCSYHGTa4ui4Ev6Ez3h1CtMs/3TjaNciZLBKONEGXaHy2Z1
ab+bpbCyFbtQBh5ffqPknmrqtaJcQueifSdYucZgyLlfdv07ddQBb0gRXk/dp92xSzSDyaook5s5
pNWX1s2+ckQXq4xPuxc4cljAG+nHCzdaQ3E4zzAOh7vNSEPKq3Y8uS08YAtHyKW8rYjyy9o+p64v
/q9USPpePA9V+PcEHbSy0RbsSxvwAIeXqv0tLGuHfyVKOgJvX6rnPBwz/ArpvoGL2QPz3i4UZoS/
C5ZDOT6oGmB/digZ97RoFaQTUMeVI1B0bz9keFZS+qZnU+5dNfRLOvf3FiUt0nrHTjWrPFmcJsab
UTM8qB5TtxCV2xvmFnmTHPwhPJGvkWOFjAqjut0yqggakzsfxg0a70ozxGBVsEHuPb/7YPQyIByU
S1Oe/S4xzXmfYBNGyJLOL9grdEyDrUriqSa6JEDRmYkTOIH0xAs5LGq7S8r2D1V5q1zn5ce9A1Yr
etX0OGl20ejFd/u2Ec82jvCC7X3PdSVAEwSYOuaJFXs9ZiR6ggU9pHgaDQDNGDtF0N4WCF8T+pIx
7aVportNG1S0LMKzvcTq+36IOHYq0aPufxTcuP2Q+iRazFdFW6Ni6t8AK7bgzqs6iXKn+6T4e7Og
vSNz2+YcHkcNL9svXXygKCBTxZ3UfiGQuWrY7FeSqAvecSS6z0BrzX6f9YA0ka0LKKAk96P6biFS
4vjRnAseFSklnvQAFjV0VW0IBvHH1PZJBKb5ipJmYek4KgMmTRfP2rdjdI0m12GcWqylfiOlO33S
i8s5xb2Um9zV1hlb5ICNA7T1oE46tnFW9siQpdQOpBuySAApq4HQi0y7SS7I3zHWF6Ba3zn1GEjX
qb+6Y80eLCykXohhW5j+PfO1Qm2Uo2kM7OCLxh/iWKZHZzVXhqoR4Uios77fsHVaEYLIbkdUZBHv
fNL318v7ZC8Lga4SdAYHFizSLNkW0ykNjpDkGhXxCDTXOV2xQ0iCAI8yLH8ww/Mfu5TKwFoJGtxx
wIhcFru84K0Fpu2Bn+PiHgez6LNt6qTWR/E3zLdizB0AA4tSuqwY9W47pVVTsPdJxNrwGEwimOwx
7IWHMa479TEDN2QUBr5174sQ2+2HhA63Bjx9uQONMtwmGyXsJm0N6rwfqno82XXQbTFuFq3KScDy
sBirkGFon2dMdUeUZX+YmIGUwYfeJ8yh7BVij6n4xI/AXWBUjZQqlgw6M2hHgEj73y3qWWHZ7TT6
FmFRJVRs8d7PT0GQLtpfyb/fdDZbVwigSMw4+pz90YblfHVoyCx/fDVxS+JwSOHhhjPZPSMlcVw3
KWXWNwzjzRdo2cDS+cTK+4UypedEGNpn70KOMSxzqndk4K8fjAOLpmFH5qxQdGVTkVciu5T3tPbC
gZ0XlLAp8BP0YajANg8fX49uzGtr2id+xaSwEfYA9uDMH7yoJWYSBm3BfEZHkJWvQfx4XwluwKlN
47KNH0r9/uYsNAitx56MlJZxndgd7CnrdppAvHM61uWrcuYWyj00hs5kXWodmZer0qblY2uFwop3
t82WNQueRdJ8EqoSNf8JXM7i7fiYWDO6clRv/6vwRPSj+aP23F7o52S0r6+eXCzyZHKrIwuW2v7O
BiJuSl2+cpJL+6qLo1e2JtC78wDa0J3Z2QJv5zvzAzUcYBKEUIVHBQ7YYjd+H9AxyegtYRH+C+NM
Ys711jFF2m9vWv0jsOpUu2hUJ79qPZucUnRcD1KB78VjNfxDRck3GfLEERT5OerKESiw8Oq/dqPO
fa4IVFOR3Ps0W3ZNwSb5d4OlzHcytBpzqZ2EovbgbDU7EDaRw9qVudYKpMiooP2Zvqq4kkUsn+Q/
e+pbdZwSWBwwpwJUSZK99+XSRrrgp9PvFys3l1T6VP0/ZWITweWz8zjw9QlVG4cXKv+qk77QkjMf
9KbZ6F+O+uMQc3JoSe/cj2TLThudwmbkxWK/SICx0ZXMg7m37SlKEn4UyclkcegfjsdJQ/53Un3T
8+8KOKuvEYu/I06sZTQt624osFDAXOek71+j++jLiMwWAJwyzM8JbNYWi2GuJCy7L3ju+81I5jcQ
zHHpKivC2xgDuDO4f6sptGruMuEPqAq33xkVmFeYMqudDJiSthCpwxSbu+Q+PCV4Z6BZpEFw1Rg3
tBjHSQ9qis6LLT5gKqVSdAn1FRvbw39iN5JmTaqHiAdWA861uxlO3lreoW+hYHqEz9C2CC08YVbT
27mLK8VukBfj8vvAZjbJLWsU1M7+rMrRlxmzP2SE8QgEKhaNeqEq3XCV/V/9yAAxr4CbHwhx0pGG
ZPszEnmINK39tIyQE5ZKv5jN2eE/D/W/oXEfw2Uyl1tMdulFmCgTSIqS9S1eCVv5QymfC4ZLRiz6
sm46T7K9ZZcWvoo7qyD8QkR66Jhq1YPTLJI6oF/ao/VUoaxjGDrRNdCXo9v8DdxnePFHSCfOEWAQ
4JMYfIBxl8DtEM4nDmbtV0b3fMoU+y9oRKyMeJKSnb+sgS7bNI/fLam1lccnBbSY9e3cDZIyq1jC
LSb+Y89sSvqwu4YJTcD1X39fanhOHSaccNHYnhwG8SYQifcIMiUf0TTBCy+HCVZJ+AL6RWtYE698
KKmq6JYN+IKW6LxPmWTBq3XGUvCl0h/HHmuMF2hzj78H0sE9p2GtsR99HEsp20DbPT6Sb3ve9KXe
mcXcD1C9HrfkxjWiJ+vBWQnqYswA7h26WinS+GPgL4bmkrrQVDwCtHnK9SfZqvVEYD+5UG/bwjD9
2qPEdFjhXTG+NAFu2Qcll6Y+nrHVM4ZcWPlYYQfRaksQ/Y824aRcx6kSKKNHbrr1Lmn5pFTVgaz4
5vPCp4YhahC3Oxq2xeUwSnrp0qDTfth6UwClWKlcj0MIxvLDVKsl1Q08pgNQPZqJoZetjE9KmqHm
bhaexIAemFi1vYTPFamjoyr76RuF3F4e7H/8deAGAWUPy419Gp8aD2G71v73I2RJiEBBk8eoTfhy
pin3TfGu1yjTHAl9HPFxCh6fuwhbp9DmB/Hh9EoImlqkEOkaknLRvMmVt4If8bYTemzU+XEZP00G
MRoiNQdjrcirwHSd2wPwVmwktgDSQVV+bb4y+TxtM5eez70d9ZsDCU6+171l/iNbN6eSFOLgxgZ5
JU6GN+fT6r9z0ZESr71sdkRFWyoDm57A7HYYhrkVb/8+8CdjRt2OUKJA2dZ8zazGj3Ovdi7GdWur
DvlfhvnRRLUsr4xs0/Arh2Id5f/uye8+BQ2i8GhKtofAud0ZTgCcBlVKK5h3pC78XK1oWiA9EOJP
glXGGzDLklVSLRa8fh0e55E/9ojd1Y1ELPzkoQtXIAhnqJsRebRQvQR0u4Eij/x6zjkcMKJZaxke
roVRpCV50vE2rRtw2Z+xFwIMF10k7VHXx5fl0cJjquOEanJZmRBwed+RzAtbx19bHfvvo81SU8Cx
vWJsJYnrmO+CPr6Fp2oDxdvp9bHi5zL0WMAY3XOIMc59Q6A/QAGK5VHj8tfKQdWUZBlgCD4nc7Ci
VGIzTmdOjLllWWdDN/pkBcU627VTmG9DDJg6v6ccK/+2ggA0G+T8XAABLNqaf2BFE8aY4MQ5D3Bz
p2lgyvlnUClRtgNiS5Lq2NN6WqOB4//9VmjHJx7gB7q1K0pBG97PfTiRfP6T6/fHWBd+W3aZ6tRE
29uzNTiQVGgRE4fAFrjdqdcMYuKnG5TbAKfX/rGe3mkMeArFkmX/8TpElEiGDgF7Qtu+HqFP70op
TxCNX3onazPElq2RDz4GlM3qE2qv+vmxvzpY43N/VQTQRqA0NzWkWh7UZS2dz0p2B6gIFU2kR4Y0
AYGif+1dahSkrIcqPYrg9vNQhZVVb4DtBJzyvITcYnw9t5k8y9NngcuvMigeX4zlR/x+583vo5Pw
FCwOG39wE+T9hoP5Fax7pM6SCCdonFRKe+wTHi2+oO1HkZJxmhJuXjKWfqm2U2te1JAdm/rQElQV
5IdhFyWAemGCS6khZUniDxEW56Thb0AgUAm4VoDwaPHGkvlPBjf76gwFi+GoJFlXjf9FXfXWk4yq
8jBcWz22ijuyWb4VGB0GZo4u+dPi/2AjxLwiQq5d+7ZzavBNN9N4t+uIjcpSA2YTfZ9v4Vr6oxU5
O3wmU6U8KXbI8STTTJxUPj7Nw781hvOS1g6UmD2w9Ful3j3knMTcoAYlMrF+rtCt/BhGI/cuLNQD
KKGFzr5fKBmok+uGtGQTl4yKLNhRNi17s/BrfRrkkt/kRmLIywJXs+SFXL2J521isCDj8XqbGnOD
/ppiMaVIZqyGVT6N4Atky1quATkQI8BAIvpxG+Q0zWOu9V2TJEHGNIrlyxWvHC+G6ejNfW591by6
5UIDuzk0QADM1fpnfjPVDKG7tAV9xcNsg6enUYe4lyDKxElC9WuK2zgJwGBMKpdBB9wUuLesUY5R
G/IeWmUaWOknzppP512VQJxTc1V4l6VYG1v99VsMtQEA9zqttKCf2X3ZvoSX5aen91Jo7+tfG61E
0ARSwEic6dDbxf/CZxuqY4Yc8VyGVo7lGLWIPMnm46qHMzZT9Hc5gYQZ258V7xV6YHLuIQ/4Yc/J
AJWWvLsMdmA43le7QbSoCek3b9lAKlYibB04329kV3N9RfgoQVFWzj4MVUp0TgrgnWaeWJKa9puE
h3sYqWwviR0FakKpcAyEgMUaycnV1qOZpPrqIQIKy+GgInrNHW8CvCCa+R8k/9UMWwyvZmyhz+yI
cb84m9/2xeRoaZqu6bFcuW42v+V1JRP42kMGBaFyAInSzhDWyi81u3ImCInvaub/+WvqoydiBdNV
t054eTn7TesvRwByDxkf6UjW7+09Zdjn9W5ap49VJ1jGu9n8/Otp1rVtUvifLV1yTTYWhkhYKaq1
RJN5Ir+fXgibaY2MBClmZSwlhKwJUw92iHBRwI+l6QwJgkoJ/rkAuqkyJ9vbdrVGb3FRybfPBCnB
qLHXLbJlk03GHvF4JQheGdQWe+htiKLSwZog9u3LeX2W6UkfGG7CTc7dWLqTG8/cZvU47EaOdDh5
ihfy1ZFA9ld0EdUpin24BeoT3yOCpQo+ZSljH9hv9xS6pBtU6Z8NntXs5JPPmhDCsSgDrB7I5Nit
Aw6msGb/hZe+BifbqdOynVULFaLKYTSuQHbltbcac1mIYhNeRv2M+R7D5KecZ6TTCCOTRSyFJyIC
slnMwjRd5DBxmwamjHV/HG0zEQt+kAwRndJ1E8db+5YYYtUnfWZQ7yCurAR/7xvC+PbN7oHNQfwL
T3FRIYKbEMXRofjAZ4nyqCZI691QvFAhi7j+pNZXACAkJkj5rWbcCSLspAQGvpj8CsTlHzIVVI3e
v0nLTXKnvU3YTrahq1G73MmvuhumhrNHjeWCURRV8izX6U36wMpZE/S4OSiLcgPU7U//YcC9rys4
0bvgGU52zvHqqjUPTaJiDLbCNQiSOaqZRC9UsDfZCpXw1XdaauH+Q7CquughF36XkSwXjYgdkuzv
tHaLfVCSsGH8LlUO1AnZM2+EdG2C64oj52VCH/mZXc5ZRv0i6mEJHXW0QK8rTdj6Gd6Y+S7RqxVb
f7pDBq5WD+1nFXlY2osf/ar1bljhKTT1005r1ceckXw7zm2+E4VS6WROSw+0JpN6BoJUxLrp7wga
YzxxcvJgSgVpsq2vErWTF7Ryp1IqiExmGufg0OcyEhIed1zXciNHGMs5gT4qLzjb7aguBIRdrLvO
X0RiSrUhCODmwjGWNkANpmXQrBAsxhHER3ILQSY83NPi8i1xPfE2KVsylJ825PGkrCEpffqTv9zB
EJevmCpmB9Xwr/bumb3eAOqvZfu5sLNIGDaqI+ATYSfr0Ik1uZaCbAgzx2HcWDW9+lkUQxxZfcbt
USGqOijHVv9UzmOms7mD1+Aa1RsdN8Tf6a2sdIxtbV7YQoK/kGgntAGq9HL14JIrLVfD1K05ca44
Z+cTO3kJJlbprNbPut/wWLa/e+omCXvnavW45iVmI6MgVAP0wLmO6aIMt52tQr5clrwOowCh1UGW
kSxOjmVCiviRyf0FouT0NquYYNQWWMJ0H/MOzt4SuJnAfKoMK5AuuJKZ8Un6+lO3YlXTOCiuQiiX
ZYSihSw/UUzpgRTgDBbglYCUE/2NbzIoy+8uUzjoDnDpK7ibBitrsiAb9BBTip46XjZ6Tr/1qVFi
ij+sMObkDW+fnygHNNaKwJZHYY3l+PBhVIQPaR0GTOyqnYEq6F8FRnDizzbBIK5fCYwf+pL60xHE
KNxA0cQXQoecabxWgG9Rmx8Tyg/zhJWnhWZBnhBfr6Zl14HbvtXpdc+8PpuvQbB7y0IeN29ciVvb
x/QxEGHj5X0y5RfofBkAlr1Iv0s9ypx1E3A/tK5nYc+SVSUeo4ibemuYKzuVygYqlVJOeQ7MThwo
mmHGPllBhXNrvIMFSyMzPacOsHLWmXg2lghm00nLEbEHEHG27LphcowlyoDOoEVOvobKC6qHeFl5
XIM3ULnKQnmhKCMlPYVPYEtNW5TD8AohQyOdq13Dcn7fhvsiFgGBMrn7C+/Iyj8uiv0fAXDL0nLR
qL/cfzNpVktiR5h4dEKCo8PiVUQPnC6F77vIBUKFQmTgcR8cbs0DJ3NW8vVtfuu0JfIN9mGHUQmn
AXmWgUO8uLetBTMzZnezky00w/iFaAX7FXW40pthWmwEoQvnN9IBi4dT7BcB3lBzHUlkK/sp5VtB
3bNTCCDmKwbqRz5wszHqo3h/n4uKY85ckbJ1Hu0A/cYgb/PQOiAdNFf1+cVCQKb1JuAdnNFBkltK
RCHbfSx3iQDSZIQ03qCC1FngZUjbCtgWpwDuglCa7qTsPWT3ItbaEx+j+rl5sRnbfvnLDnp2i6Oo
Y9h9peZu4TmxPrTCKc6c79hYoXl8MU6ClsEoa3Uqdh+ASo4zVkBB1GjFjYeNCHeUo4VxJdGPp3RY
Li3gweqXxAeMziL6mYRE4dhEdBlY1CYr/xTYycJa+mTcnjsAaWoXKOUQvi9d4sT9Utn+6qQCR7Ap
qn378MeXZKm+LTGdRa9xRVkVhcXlF2qUKqxzIy5wxtNqrtzStf974fjVGKFIBXAaMU2Mymw25jHE
yU6ELzL1EozNraR2gndbSQ4cGJ4A+4CzklJIwTR4g6fS8jXOBPVnHp/rzcLorvAuscd7/d+llLq8
sQbMAKfHp/7s9gWuM0oEgV+g2h0U4JP96TV6l32kJxADp0X2yqoyx9jBGReiuf29ck3MTw98OCOW
YhGxJh/IdZzqHTfeagFzDa3kqTW1lQQSqk7kHxaFHXjyEjkKB5ctE1aAXCRuncej3CfTk4dHy2qi
NplZCIw8Qy7d19+zhW8jhgPOBJbOx9ZLZt40t7YxGv2fOu0A7lG0488hEJF/kGa6FvXXv5pPhHOw
OjIPq4gb34qIxvrbL0KUhUDD0t9w+dKlibtKEGEOQoF1+i0mLFwFYAF4Lj0qVpaLSiH5hiN+UA10
sDP1awFSFmTvaxcw6KEkynRI35LICrw8BBSxYGZ6OTfYTh+rySN0vOei2IfdruXAjxDZwnmeV4x/
7RCZelRBMSBvPgDFE264HQPhwWxdYe/6ibu3f5iXPGL55EwvtUo8XlqOuVpLPHESOeY0+VqQNC9n
mB95ojzn24W1xAv4VyuyR4fif5rS+3tgT4l/udP8g1qnd7LD2SzpNI45JPnLDzbzhNcg4XnX7Wqf
I1RdjuyyAgpvm+V2i9FAUNDrgKl/UnM/YJLEc8cVFLHFK+PnE2xY/QwZfk594k8PKDqCdEo80pEa
jEw4N1ZgDLnM5/9ijPywCh++csjR/ROd2okxM9yWKR0dpKXPK4Tzv46EWxDewqeA5UgiuYbaKddk
kTllGolEMO3ib2SMVat57HPSj1DHorc/OzyIBKvxriAKsJurwf8frnL1each2xCDhcntdM4fNLgM
MP0v7xKeZUKJvIzcF41YDYy4EyNRwfBrWi88kuw37l9a5TV0NVbhJrJN8zEQNPHIgFDSQSRw1ZGP
ex4FOJjonDvQw7nHNqDmwRvJZeaBhttKC71IO4/CSqAjPctftTlxX0juVOtQ4tl/X754fZzW8fIn
tJQ3NGLz7f8pCVPhW/tlnQA2cPjreQmZeXRQlcOW8sd5P7h0/WQHcw7oytDAF/dqAddn6tYseNPL
TJn7vbTAf7CsiZGzrvCIpa8oCpKvyXzmwMehKhCnhj8ro5OiCVt7RPNcGH0m0UuCwS+GyDwhzt2L
HYXOBtsT1lcrYElilLXn9GSs3Hx/oL7GyvmvehELrmSktMxJ4DU0O7hRqZvvodN/XqUcqStT40NQ
bul4fRjUMxMUSPO9BkMHOk/52C4B2Gjb5MQ3weqvP20Da26EAjddqpXPTClwXxA2s+2+wbVseaui
pNvFswJHPfqsrei0I76FmEaiGhv0P8LSGCnL9BHsxrPKd/G8cweTdTIE4Rb1+CH1R1WFM/XTD4Cw
tDOraA/vvUx7kmz3j6A8bbKejAZXMrKFNCNYdRAb8DsMNmBIcrWMMXTRo/RxjJEvMb8a3Zz9LLlE
lADw9gmGAotU6T8l3uo4ZmLrhMH2qYC1+NILA3bBWz0ePDiXhpKjSKjT2UQ2sFsAvQSzy9dHKD8h
PsrZZI1MZ9SyeC+7h7qlsdlQeBBRfIsi6ka4NZK2YrQ3tkuy26hdtiT+nYqqQOfONsk/55eC3jbR
NMFcF1Y+dzUBoonRw811Iv8FXTk9hFprd66W5sIkXn8yURj0dY9vnqIePtKggzpiib4diCXpRc5z
s2sW24qKa+VC6f/AH31Fn4gnUsnUPO7Ihly2158NP/9//IZuhEPOkOweIQI7Aeu+dqT3Ni9x5ytg
7MVLLzKTyi4TFVDD6NLsTmvbAddmW/5MVh/4rtzI4PtWEJg+MCJsX71+MvALuEFqWsckzY2nTgp6
tqq6ceKbVZJ/cAiSA+p+oMFxUT4ol6quvzk7nBdZq77pkvaD+qIffpers6k8NnMLst9/CTqIVYgM
Og04XWpUym/BCp0wO3SuoH/eG0z/nuJX/fX2Lv5J+JANGSYp3+rbpOHJziu80pZesmTtpoAQry8p
72gzw0RB0eayA/k8kmnfuRPj78yCDhQBjTvT3Fw03QxhpxCj6PrdFx/j90Y7E3pTRar8fT6KJ7RZ
aPFy7tBD8D8VNREZm37uilB6wEvpySBxYBBVyrXGCQq23Ghm4+RWBbMWDUac8Xt4DXavMRxKszj6
Psiv+5vWDYqacJelwuAOdxEgu39uLpMJrDlWYsC3SI79hf2dfYwHa4lrV0Fs2eanfFSi6W8FYC6j
SnBueABv5DQE10tW0l72tblshnA4bxsi9BeYBxh/eHEw8ivFnSb4NWf5rjcWsytto7lCWkdpBXWk
ELsLStjW5MaakmUzK2TRkl9lIa52W3msJrtK8socVFa7VLka2UGnv9ym6oHRuW/yYfGW5fdV1HDf
9ozoCmr/6gWV4V3JaJYp6PTE6VusX5ZDO+F6pP99baOZIwiRbLLRGRHdavKaChDJMx4kLzTrtJhC
zPUKV4CyIp1pWbyQzB8RVBv6TbPmZ9CIQspbXA0fpfDuUdlDmQBipgacrQiRvSipEX6uX7iXsCOb
G4Ho2suwCOiqTm+qkEPbXsq+gr5pu3kJE3XYhjTWNbSfhn47PRObdV+3+Eesl70wzF3qNtCccLum
3yOKF482VxE+dVJ8JlyLqqcWk67g+hL8YMhZXG0x5DcvRr+O04+x+oyFhs059bX5GVn5ZAPv4QKn
Y6QBM+k9i3ivvDgOuuPgB1OvA1xcZSq4pCT0tucYD6Y1P49B674neyLTxtvUiuIpfyydBCwRIz8Q
t8Yr8AQaFgBKD7eOb5ciIi7n8fJYUCapypK8dF5vlMuQDqabOiLHI/IJytQJBuYZWnkN+XGjuIph
2krp37cfvppXctx/S3TzNP9Utscx35HeAZ8qceSrD9KThbcp/zq93vtivI8QVR3fWSWYCVjOyTFo
0fvMUXbgP6V71Vs9mm6te28eg2hfgBqg6V7lDSBGq7d0WUL98lle75w8EBb6WIwZO47H4PCfybsA
Db+O0vNgyrVPeGNaBzgDkZhO8DetP2KDIgLPncjk8ZMZWOC3fU0/eoEDQVvzTMX8bEWWuK17/Sph
W5b0YwiaDvzWDNTpXDtPG5RCk1CALpdOmXyHMllR1Q+e3+NILoqXdTFizTcshmXViZ4Ktnh2ojUL
/pH1TWx4+cZMMpI+kV7ORGW964Gia+3melGShEZw0G7hlYOGTAK0kB2ywxi25I3XnbGjxlS/M2t1
JsJw/dDvFPrkX/pkuVlQy4ZxXGe0dfOAXSlosoA9lvlMuYGsIySZMaXdJvTAHyTYBBXJynqReaQz
DFVWIeOFQHQEptSpv+jEof22WIZ44T8/ayXBMbqDFW6Hb5RtlpmLECzYS2m5SbbhhwFpntQDENG7
KVFVNgRwqbp77YKRV2wtjvXgMb8pAjXTsuLzxGH0v3IeSgzClZ3bcjwVRJBa3oepbx0xObG2xbIQ
ujtNUcU2jasBikCqL1vdJQpRYR265JUKPZB2PlbnRES3PmUBw0sLPv1vNZ6pKo2Vgidn0H4/BlHf
/LLIjmjaxSNBYFJEICi1289ntk2DapQ0H05KvwEHhBF9nwrF3Q8uvtD+ICdgwzrKtDOpxz8jHdli
cUce7lWV8vMBb/UqAU0WhFGKJAyUWxKrhU4nvKI3LYvGa049gRRzO92mYQr4JdFm8NIyBUa2K1TO
q/IzMLPwKSGLP5i/41WkLMUCGEdwABPKlAXZHT3h055Y2vGREoQxCsOysgwNZo7l58uXMVXWecoj
Mb7RYj6ZbNbk5RSs8pAzgt4+LpcD1nhl4pYFgG0lpoHBggnTMYkcZ6c581/XTeIe9F6tWy9ezIlb
fjrSt/we/Eoej+QpCu9OGjzIuIcq5Se7S50wBb012VzqHDSeJrViJ0HW7W4hRsvgotNyM7fT4BXN
tgqfNXexcVF6Nt1mz6lvTlE7Ft5PQf3z06HqN8AxUy6bEURhgls3IV9SiPACwsw5p9JZ32kgn2Ac
bE2DKWZcBPG9Y5GvJtBFqtyVZ6QOFvtcZWA1ea9cjayS7ozQP7M2qIvrS/X+MNuuQUfiJQkZf1Vh
mjKOTVB5aDDHhZxMXgKZ7o9X8E9rCSyaQMEqSyxGElaxDTFjC0xya3rGz3QTLNY5+3iDwZRyTwD8
dIG4+ay5nzwydYLiRGqwjNUrzd0f+SBxjEKjAbjoedTP/E6BWoA5RCzQdDpaEKESkMeY9+0zDdJa
6JWwHz3OzuQDBkE17LkEnSiJnGvned/H0hGzKwKr0HqpFExm1umck7HY40bTNJC1xJUAeDFGgaL/
A4OJrXUZl4CIN7I7AmWHHaoSRK5bFPJ9/N2NR8HpmhBBcrs0L3J5l+Ch32y16Poft49g50YFLz6v
yTA8OJs/RafsgR7fCPFkEkc5pxW9QdyNuOtecz0DuFW+iB/gYzzNUBanatcE1WdGa5rCBhbfozJd
7Y4+eOOXio2mWPmx23Jt8nS+A4GSYUY721+X8ITbemWHbXewi7EbJCIDCh8V5rztJnZwMl1UzdSg
lkcUg00UfSeFTjKTwtYrtywjcDBERHg/HtbmuELkInsOgR/tA4NmlGzpkcTJq7tXNddpOtE2FpCf
Ve3MEGOV/xWCBbRU75nP4bmIaKDsw8DSgwHQCWzncJlg5SbEBFIBua2p+983sC8jrvdo7q5tSEwr
VRrGmTBwNEGHWi4Wzq0FTdZDYCviQ4MYhrKNd3ybWRD6eiNeZ11ECV11wRe1VvIHRSGHzOSgHhrl
3Lt1kAEj0dPTjBGcwVz6s/VQ4NoYt6b2wp+ENIS3XJB6DKTmzGELnY29aV8Jx2GY6ShSZh6iIi1C
j6j8eI8+iO+oSTS9q3aXu960AdLUlL2x08LRPDQYlJjrv5f6mjYE3jSh+DIxh8nl+wmAmiAUkpBo
RcJCFCESILItyeOtG2nEqaRY3bKMjrwZ6tIE/jrLEF5K7fmzo4KPWGm5T9cqmea+n+UmPZMsSINz
XgvlwYEx8F3OWWDRzDAl+BFN4KhNsSckao0/h+1PBckjKxZ1vkg7FuUmGofYwsmTVw5ddkqtRjoo
OVxsWvEPKkmpzJ/wRTM4jUoCWUgquFu5f3atlyMb8lQnKByfqS4jKQSNqjKxTUKVBB/YOKCcm32+
tZKXpp9X4IsLNxLdYcwz04MsvhbaFg2Vro3PuDCCwrejvwF+dbGlCCeXL3SpEA3nBjL+OcE2J10x
0pGhUPciE2QXjyf32H+/pQonkdLWMaW4zWOxn+0hRBd900Jvdw5U6LqBdF8Vs3seXEwn5hGLlZ6K
+HgIBHhcIrFSrG/KZGJCbPqcUCdBua8hd4aAr8T/YUqbHyzbswavk5fp4AtNLhh4a1QL5BR82INj
swtBJhuOUYrYJMzDDlM8FSGLL+grHl3lHHKLk4gt5KlyKqJ7f+SqPJf3LKLHn376xsicyAk0aw3d
nWxXFEycXsCPEVz6gSLY7Ljbu4sYGtOXOQv3Lt3zKUgiEF9qmTl8Y1C5Oalq2cyzgPHDjnVKUcSv
eHsz2nf9YUXqsThg10FK9CxYc3DLTj+DJVzugAmbr+fwQOwbozwHuM/rNjxi5VxXOphbJUHY6Iid
dTZy9jspwvmJGmiCJoN/lD5Y5KjKWfz4aY1mndC39IFiELgRqe02wIH7QkyU8DtpvaVyW0yfmTNK
7U2JkuRV1I1mEO5Dj4sGjwdtA5G9IZ+MFgSutBQWl0BnDwjlhpWKnrVBYYDws3XR9RSs7HW575Dn
4cPIK7iBg/hqeqppwN6GimIWEW1iP1gro/6FB03xynhZJgFz6OzI/XqQy+PVS3WRNTQ04fHs849G
lNDobnUpvXsMfFHblZ8u8TaMxTLonV9YrrVz8NghaT5ptNirwrMoe/seT+xveJJd6aJ5GGc4jOqX
gdhglPJHCQe1b9HW9s1bL5mZcjwY52z0X1z2ixCXIiINO/tpmqiK+2PAQOP+w2mXcr38Qae3WsR3
y+vxBRR9hyArgDsMlDDGU4qnqXmO0TWUuX8H4YcsWSeoKLkllyAkuZJQzFkO29s9Iz49vR2YWb38
72xlslmcQuybNmzt1O+m3TKaxiwtSRocvlkRUN0DCSNzs0q+QzsgafD1dLoaiFxk2TomLgigVMvi
SHq8lkuANl/frIKAp2vlEqPasYva+g7DG7pCra0JEPztHlwnqM16Os7gbDpHuu0EjdTufm4mlfHv
aildko1Qcsdl1cP6FlH4RMyV9jB5GVqmEqtv6utT23ByCejzDnk1v806q6IqVfu0EZ1VWHMW0r45
LwESWkpW3pzjaIpDxdbYwuusYzjHOL4LHRUBDM9lySJw/gaV3T/zgcPPPlnNUKhKSh+o+NB1k5RI
0a/twvzv8Z7otl2YXP2fQmeyCirSBdr19bmV/4YzBhiMt71nnJundfygGDD7GEOk1QXrR5eBFIk1
Kl2JDAe4zXJYTHfGWHAg+QoayN8ttAi+yL3q3LWk2wy5qxdkeCg6cfBC4qjVEUgNYLzE1japsYmP
z9gvvdVg71IfbgYxvmXiOKNZ2Og3eVt+a6o9UEUaCi5/cqC92T49/AttoVNjZl/NXaCuJgsHLkQR
2BmUK1AlVDfAP2o8Eyw+R0miH4FIMNIuS6MmAcw5fGepYLoyaPw6vKe6XJxVAu1C40T/npESHUZf
ogihA6sPvCS6p/491gyoUeMKe7pOviZ0h/EO/EyKRg+USlWXLoct6F9ou1MDSwBnRyKj0HO/AiBO
iwxW+q77GjtLwpBiF4hgafEfkc73GQGzGmmbs5qI2YfjNXtEIjZDIvjZq08e/ww0P4oqBJwhrawO
q68fJ6H+duBgSHxCDBy82wpVP3X30oC3skvX9LTSYcYQpJ1HqSnxM/W+8I5e02FQ1VSufVoUd+a1
mPIZzbSPlztGdYwMC5GcU1WvzD6LmGJz5btqm4lQf4Gt3PFy7FUMMLf0OAUfLG3Cexlr+WW+49in
ZfRsd9zSZLi0HyHYfycm3pS4HCKcNK6U44ohapwDSv/+Uf8MCCkLS2TaGesT8Sdv5ww1H05pLvz5
lIrae/IEgHqlJDgC2pzdsipZPEF0QO78pFXb8AwoFr2Lv4y3Wdo9uBm2DOmOgB8nrskr7suW0FUS
r5AutP5Czka+wlLJi5xBKJGsQW1UcoDa2DEUrTbTTYZzuAvXL3ofk4rwIipbQCo9lo0OtK+fT6bq
KdTn6RxI1gXinLmJ/Nf/WjY5nmYRSULQvp13YJZo8UnMwZ0SPbBI26olg0moC2s3LYdgju5kVMrd
+V6mpRrRsbhTSgP+swwtEyRpVF1/VKF5POsEB+OZ0ok1NpkL8ttVR0SQMrzwCTVJYzexmb4JPEEe
nVESu8eUqn2tT06YAGw15mCHWsjJCnGIQhSID/x8UCYtEvCVg8YDC1Y7LUMYCc33VxqhY27iad1Z
RDbwcDKkObjN4b4y+tfr2RbSMbTi5ATitgf4Wd512VB67RtzkKzdSQnKwfh/okmEl3knOK2D3w1K
iHfzK3AGKCTEwpvnIEBCG7GJLc26USGgfEj898f9hneeh4lZKbg8EW007JOtiDVYYPbKis9oIoO1
HsyR4LHt+G21JD3S+QbwY2PZMl0EVbmIe97GozoDy8Kw+C5Nk4qt7QqwHFM167muFCYTRzTnuuSl
mglO3TlWQwfp7+G8OkqlDBk4muAeVQNDQJRbjb5xag5UoYKEuXA6IDaBzvy/7SG8Gsg76u0esI1x
x1NV5oJ3JmMrbJs8AY/htJL1BXvRLICXTQhl+3wiGiw0bo9Fd5t4c7Q8UpPKaasYe9b1igq9AuxB
yy4dfdjkKiRML4ZhlJhwixoXjQEaaL0kTd7tsOZKRgxXMsHFWw7MiS+zTDEgMSHXyq8GDXqW1mSJ
iHvZhs1TQnt0yOP9sQmiy6hNfZSiaxkk+PE9SGDatxfeJvRVslw+EIODul0xJbQpeZDOV9beUvsU
Dhar8qpSz7sRN6ieL8/LfdpDqqbuSYFZOkPjRK4I7m4OI/FdCpyHHrKZhrfpOIlycYeQh+T/P7TM
QZ4Kl6YfENM4qcpIOBJiCnv7vrtE9TPZsRrDH8puY05nT2tjbJMLjtDwABdKk2aAbobCbqTrpSrQ
3p/ZItAn9o7gZ3/auBJAJ/9qfWIANKZnsej2VKRZJihXDkP0NEfnaYDi05QuItoeGTDzPWDE3XzA
n9xL9GNVr2NzdBpWdelWRV7uarkrexh01y9y7QTq9P+MSMdp60TLMQRuJ9L1u+0Y1D8ez8s2HSK3
4uMBD3qb0+Ab/aGL9Zzt90eVs3wo6cVZ95ziwNafuvaOOEod/Ed0/aHL4wXhprd8wdNFJqgpIf8G
2JDh5GLYURPCdGHq08hKQyAkTRY+mghnPI2F68RDzXps4Q6TeHXQeiy054QtYBbVossqwaSjaIS+
U6zS4/G5neoOq0Iom5y2KbZnSRKIkKW+Znb3wIpDhYvtJLyK/kI6TQtcdKtTakenc3D9LGp0Y4uG
eaMUUQJXjWxga1K/YTXTKtb0h8Seo8v4lkOsp9vdsioUgRtR+0zkSaKo2UkqllUHMa6xj+zkn8tK
4GBcaZGM1gpfE8EWES6M2ZubaDwCtxuLAp8FulJbN39aUmAdlOiXWU04qP/fCG2RtCsMXKpGCLcJ
CvmkU/0akoCsOy+ZNx0Y+pemFU9KhoBst5S6PkWCrCficf/DlE9lI31YnuZRomUihiaxqmtVpPtx
Z69RIBoB3UU1VkoKv3OwTqPxc0pEHyutCquArCLnFD11DnO4fMEXVPDPDE6B5xwH+OHCPH+LEO6Z
hbly5Z2TtaFvtz9H3c6ca73fuHwp6FMmbbem3SXb65jnfig8GVOEm86NBKr0nRwVyZ6s2AlFcZKY
Tm4axPVOl0UV2ppEdF70lEzcoSZHv5dN9dqafJqVzabs3MuUohmwH2rXmLz0qPzvWABMeXo2+mRv
11fbjK3o9ktWbJ7iFTaPu2hVRK6ieh3w8+Yt+WqievWKNCgcfGpe5s9fuGEJo4ZofSXJpB3Kh2DW
87cHwIDw7bA6v5rRApVAo68nXWGwIC3SBbxVbw62bNfzj8ZnmA3gfW8XKSxaOWijRzJbUpzvaGPA
JrShce/zb6JhycPCQs4T809l6K/B+c4gSmvJRoGzY5o7/6sokwPUVuHWGsjC9y/oL1vQiO6pQYfN
y6q4fIK/a6m237S9sGtng4SxkEdiTyNQfWghMnsGjnUW/0Yk4bgNtw1lwPFpDlmtfhuZ92mQhG6e
1/9ZhUxp/qAIsprPJ2xUboU0Ph2unvmNY9mhRk2VaPRqwkzE/A047Y/3YGnIKfvVzeMRlwSdN6d9
UbW4txxQHCmvbcXQsG/xGSpO2FoQQAhexRDq1K/sg9oxi8M2iDaDmJu0DL4l4JjA5rU1aSly2UJ8
EuiIku4F6KToNg/NShbmlEIXyZc0F47HWM2dH/cL8lXxJo/3LhNpFooTOPGnst9XsmEQbjFgCIF0
2dt500U4h0YAf7e9WOI2Dt4/pE1EI9Izpo4syvu8PLfneWQDKoPCFvdWxto6gHo0JfFIKgqSyXw3
gYsDGRp8PqzdsrJQv0JjLhYRSuuSiyaBzsSPdpKSp63xrUP8/1XOlpETkRQZ8L2B6+0XTNBBWAIH
2OSSR6tV1iszD5KvX/qp4a5eFtA3OyYneJugmvKJjYN+P5xsvYb8jGd6Wf7p15sqJ3ANb6rlr99l
622U0QebGK9749qtRKFih4j6zcleVGdDZFjYL99Jf0d06zwNPzyY/3Kmtv1VlQZf+Q3+TEFUpnKR
lBeFT1Sc6WfcXHgfhRFYC4ksqT8ZQ4+Y9VVbJqUFS8kAtx9WecyZmQQTwHtOl9p3/JBNVVI1gRvR
LAoepQYGDmGIgCMBus3gTxXKq24agNAkRATma1D+pQTh1sp4Hm4otVjBWFLTZS7xaSP9FTJWmP9I
8Snv82xJ/qd56s9TV+v8XOTyjZGcQqoda/6c18PmVG2gW4I0E5zManYgY7YlKCzij0O0HJ6ZJJ8P
GYJFTE4yugC8v3QxkX6tVyIUScAfDsloFs4mNbvd8yzvWoeyp8u/PsarAmjnbSH6uONwHUBCZLsj
PbnaZ0V44m35tcRg/BP7SsJr1FTUwahQ84wStL2nW0/6slzOuZNXNx7Xd8o3OMY2SpYdArib837G
NGvrCMMbvenoIlG4EIBdxTRLYharjB8MW73/Sz14UT5otRg3goNj07y9picDCf6doXJXChm5aC4O
K2zamVdBgv+Q+5ug5/cSSvbDwZBLAaFoml9YYTXvfEQaUCZpalXm/3WPexPN+K6MSXkglV/COeoT
hvbK0p+l+Y0Eyy2FdrDPRMCWGNEa59zBlOqfmu2sxdOPLaYciM2nDSYW1WMjgsouB/hyt6BfDXMJ
1Bq93gwNHK/nyLq4vCQ93FzY6imsucyl1Gt2S7rx99uRKEgNxryeHjNVEsh9ZA1FVk5uPwWNX4nH
R2BlZgranuJHwPIX5W1NhjzXKvFzKbJE4gOlZ+2fFZcy11YD/+6MOrYQ5HMYo7p1m3uLqx4TMQ9o
/q2k7L3PrPtwNKIu8aKwk0vcWkS8gPgD78jFiE4bxuYqoltddWIq8xxBNJVdES64oUKO4J0Nhg/Z
tGQ1SQNv6kWTwAF98NJ93WSZ6TYKVtTfO6cCm1BnQoU32k07nANBmBPzk1L0O4XE1s/bL6KlwUy6
uTcSf9QwRiAazngp4jSf/d68xyTDHn8uJn+ZAJCE2jc1iXQjS1DbGJsKZZth0bkYlUlxZpAh2sgR
iDZVBjkPLLluj45cIZnfxu9XSG9KyMSUIVTiW/DPQ8+k6dNnJG3u1d6UshzbSfdH75Zy3Nu4yW8a
8b8j3MufCM3KAHcVqHD/YeUxtwPDJfApqt3LUOLpoB2KnQcihbv44ZFAOeR5n8Qg5Das8omySbLa
XXvgGNBX0psFfjiUC0DlsUfb+fgAXFpBbB8riL+L9RUBBp67eT85553TQH+Q2t5vi+oDshPl4G6i
LI3sw99x5Vj4jp28yrOqUIetr+mu3Ew/s6xJC758iauL2Im+kivJZ7z0xB+3Cu/xcV24CSYzvG2T
u0G/2OEtkdtgWpNvIrWE3ycPspibT/TTx9J6k9L5FKG94lPCrUM4CI7upJ9GCktajxII3J4aXCkW
WG2KiC1zRUk42N9N5ZW4U34ntR6TnYuRFqb1XEzSUbBt1PwqXjDND8SlK4CwM5uBUw+UamP7Zqr4
26OPztgCt5UaUzdeIJ/3w0y7TmGm0HjOX84SLW3tLvv2yxB2GvhFLSxSGdWCqj8yu+Pj+PDYtA5+
VSFcIaaWDtN/BgmrapeWo3CmhYB+5RJgX3ed/OtxiXiwM3FvSdb84iqohxQxS1wKl4zqc4hNu41N
bTEs/d0bE+RThLA3pM9xib883L4Wy0T7AgMLfL4BnqqcIvvvo78TfJrwP3WQf0dJCCCiA54UAPUz
EEQkEDeoHMrwHIm/B8WaJvXtYS55RjEwxP8kKST5hG4cYhPRgozklzwCqFpdupb9Q5PGbAsrfDZM
taBw+0LTjAuJJGijWLZSswg1sjGiTsa3v8P0fXLxQ5MmNIxH9LWSH9joNrKKqpN2GTIDrRQ6Kpw5
j8njTv2Ta4m0+dN32hecKzvFgBf2bXyieiQdQOKBLIhflA3+T9Hh4YofClHiUzw8sI8IDFsa1Wj7
XBUDYe/2G5wQxKjpMSBxgUfHnZIrNflyMR3bQ9+uosstb/0ZLbjRr5ga9rAbl+rifp5UuOsJBltp
dSFCPQz9Lbda0nlYBLMrehe5kMnNwrAwOzjhRQs2yura9VF18NsPCdt788ea6keM1cQkHiJkuL6R
Jnu//MakDCdYnLpkqBhJToS1rDO2l5Or26DnzaC6wervoFR9hhXTR9rJ3zGRBTA2JphS8KXJPb2a
pvLOtl2lkdF0w/OqcPVYq8R1P95mwsHlAXw3TG4ybOjqYm88MdU6BzCCdtQlpoA0v9m7//mg3fRh
GwB0Bx240LnbZ2zTsz5D3T/SMZSbISje4naYfdO87EzvFjJl/F/FkK8lCfbPZV6R6p0aiVT6SyZQ
IGICa1IMFh0fzxfoWzSZZtzQcEDHZTwcQZWRmslbG58AKSPlG2gGrhepp3/xfLxe2E6shE0/2U/K
WN4LYGc9A/AuPRd9U3sHjSVl/EIMCXJsVNWgXwW+/VyN7yMAxFDTDpatcinPBOBsx6caYkN3TheB
MSe5Ay7yyKzhjOAoMCHddx9eFqavPWfxDVwSdMggNz2jcyfyCJFwY79rzMzAbnN3/VeFTGIZDVLD
8rJSp6Dj7LPCAu/DYRMiWrdcLunMtHet1ceelCf2LtvYBdFzzPeP1NdA3VDuLoTx809iHdvVUMyj
kZaJV/v1/tOLjRXcr9tXVDQQVvbGwUDnGO59sxi+QN8QFONq56ZlA4hhltso6n/ng/MrB8AO3cJn
M0owh8c/tZfk/3feshhB5mJFKmoLVNeZ87hFmOge/RuOLQhtoQa0R2N3yClQzYRhLVlxNKHl5lh1
+UUFNQtuVe/9DiXRM6AlTsL58sl/rHiW9zM4cpUfDd2POZW0VgBRSrhqVQSIPcd9AQ7NZt7kg4AY
mmQPz95xDsNXuT11QRRkZJsNlttBjc8KKbO9hcsgMmx0spkfYbnRQu/P7ryfGjHui512HVBGcqUQ
cAyvjXM9oPb3z0GzTf8PLapcVghUii9SAN1YcBuSt/PKWOh7AZ/UbgbhsWNqZaO1egS+eHNzxt9N
wS6QXeeFIRGNaVHKxU3S0E9kCE4KOB1h54mTCl7ZPZSrmhUOgsBZsI7/Uc3yI7uFDL/bSb/1C7BL
I/K5kQC3giHaIR8khDAT+Rmcx3m9toGyY7Lz2A9KP52XQHSPD9V9R+R6dOM2gE8/pbIJiNzL/n6M
m1CtX0qUpG11dB4T2rV3pPsVtwBIIe2/QFT85TCWgFneckX9IaVOdlOToyMwFM8t4v+7xGIPiSZy
MU0JznDVNhVvDf51593lXIB8ZW8b9ilh7l4TzLpqBXpwqg+abX+aHlO+F713ISq/QJ9PMxWTltFz
FUd2tg1G++z72H8nmBJksFKY4MF3D+kWYK3W1VWKtmMxcBBeT1ojyJECBb/irlFD24cN+wYFjg9f
v7yD5SoFvrNWV23PovdM5mVJRqBiAJce0v/MpL3RZEElQE7Gn2PR0OjdCa9EzqbKmHOT0wc2V+6+
aS04phHb+v1JEUW2RdrrPAuB2g1AuKQPPVxyIQnHXOiPPvzsr7kINf6qrHG9fJ+tzVwfRuryun6t
GsG7nAb19T/G7Yc7K9e00YpYS7zo90+yCv1iSmBCr/+hFTSouWg8cQp6HqS7JgRnuuLPOn8uqexK
ULhj4cbmve6ZP6FZKI82AH9r10k8VhGqndU0WApmFF4JjrEw/FjvPCkTHSNLE5Aep8p4b5xuAtDH
EpYNdqB7Rr0Sed3iCx3Zb/K/XHqvxhooRLQqhlmFNMV/4013olWPOuB2WLrkalsI7Pk2rDWId9LF
w2RUW8IaeXuIbirL1NGoW12vDij0RfJXFd82pbfHZHpvO13tPy1wsskgsih/6Uqg/briIP7sK5Ty
tahP0rm4N4qhe65OvTpjhQR6BReB3xP2m8M2axXWfueDPAZBCo2NHx/Vd4KXIa+gsbbPBLJPNbI6
oQR94kpIoRCgndldSsTgxyV18kyPCllLv1bH61jeyAV+eYePUx/9qP5hhbuX9PZhEtXUhl+PWhx1
q/7HCSYT9gvoaNeH1lPZT8+rRNmuo30BYMP7hQ/eEZG0NbLFxG0TsrsOSTFueBMfAAtQYRd4ZOOa
QNW8G3/y8NLRSdgPa5gfNbFoYZw8eU3d9urGJjWXVL+mrXf6WW7xEoq+Zcu++uM1ddUfgQ9tpuIc
u2UVz4SiP7jk5MhZwArPvPK914ppJcEtSsyy3M8PyGIKPEQeEaoN//S6cXZI+pJNQEHyGw+FgyBj
jVPBhhcFLMF7eG6vBWCR9tlFtVfcDTCQW3rct/zKIIal0iAu+N8NdK+NgjbOmva6mNJ9eyUt+XNg
jXzCbN1dQ/yre1YsWtxktxxYZ+wLkPS7YWYtprFLYJxNbWVB5ftY1OEPboseZa6iwJoy6ylgM74h
0XXQ157+jd3RblDrsZpmNp4oL1YCpCIDgBtDo2jPOO+LM7Ix/jzSgJsjyrjHq1Fx4xZgaUnCVW5g
OJCPN3i1/vOBXum5nSRKfsfr8YEgYXXsBkBd2DQ06//lMEqnfWfe+slW3b60DbUiRE0Cqy6G62sb
cjjwMOjXbWvS1eaGho4bKwzwKkcl0k8jvqbCEhdRBHnYoQD6Y7bRksh1r1uJ2KaBSPoKl1hLrn3A
4sJ8uv37y/oVsESM1kGPRSt/5UdyxqJKk5WDjVJtsM5/g3v/sZuVRmqK/nLdhLdTeO5AEvQ7aLkF
ZlJ0WK9K8xSOeH+q4p7E/BgWjYxS0j2Yd+ONez2cyqHfIv9Ab/+bx6Lbu2nAS1n/m/X2tw1H2oec
IcbEX7+XyQMA/SjDaL0oE5RUX4YCPzjIlTjd3sRR2uLkllv4PAcpikKN8V2uCBdT+gxeXI8ccMgl
qnGfI5U4ccSpC2eb96f6OBCQ2KgEd8O1uetsuSgCiE7TWbvvoByozjsqOX8y+Y0Lb0Vl/am8/csq
ktQDP0sIsThx/zVtQWdf6dGG1cZxtTFgRy3jhCFjWNm0OZAf9K3QJef5e/8a0Ds2xi6dEUOthgvF
W+bdjy/rzov4/gIKcZgrNf1cscV0VK5xnXqS67jIvGCaL8rRUjkQy4RKteCxA3acnlbUXhPKaOcJ
INsjOVYGByGNrwOmfbYDf2DTJGu99iIeVo1pwDtIody26ZeNex54PDEcQ6TvYXz/Al+11f9JewlR
ReN633QKVx/bZLHr1h97dw7kQ0NGAyJsEaxWgFVsJjl0kxKIZ9UUQ3C9aJoLjQvKFhXWp6bK4tGv
evRpughFZ3WHNk9xjo1mk+PoyhWq4fbnnoB3EqmQqy6GsRNfoQ/9/zMH9aKZ2/CGFkSrSZtQLG7C
ymBmVcrmkcRSIbWXfwRPHFhxcw7zrzjg2pnHrGpSxr9pKSz8DYsjtHXmOjuTTQHI6lRIXckIDbni
idpAMOL4U6aYxpfRFn0dNYCW5wJBYv1NxtEvqN5EGD8Say5QCrnYO0m/pDbZsgRMU9OinIkucA1f
MzYgB/fPPfUqv7tsKE+TBvYxp+dm2JEcpFd8GagzBub/zgUJ8Y+DHFnRI7avEMEE+tEzVo+2tjW8
Q+XjOpen8RuEMurw0TmUDDUIsrOABReSFbWkSx7AHpcCDAIxBIGsGKW4M4IEvmZ0arg49hsU1Dwd
QWDyt1C8LGCsiCoDaYIssKyUHsMI5925DQS/06Su5EZuYA/OhyyOVs2X7eLpji+utso3LnEpvTi9
n2OBTRRlaWK0u8vB1xMvXcXPjNLGRqE45NRTSqi7mBv7U38DkaQ6h+kO2Ooy6JStRq5IIcJigtu9
ByDtG4q9WFCIIH36IGiZTdb0jV8wY1csDp/D7Ls4/wMEOQHsIOILXYztY2ps1QQGc8eX+U9Zrqjo
wFMWdk30CGvaZpFvp6lr5P4Mz9mYtYngX25PwcPVNrLppnAIvZyY+2rM6qDGofYiwXhg+XJ0LsTl
gG1Vb4IiQFaR1o4YmE5fZRGKC/I2wjPk5vVZO+9m0c92uwH0sh72wUZ3zqUNI9Jo2ABYFu0gmvIU
XhoXRCrcSFENB3re0tv/NQWn9FhWjkj4RQJxPIMTwC39/gHNH2knixaLk5klLsFNgcoK75OeEm02
HswWEitGd4Y5rcXl+pNlIErn1OGFPR/TXZEKf2IWhM9OBEcs10bvBa7Wwgk0dMl7WfFEYTHSLNtA
QcpO9KmkLsQjk/BQRtTE9ROBFGHQ+1ozuG8G+SuNKMH2/ogU9n/lQNlmampXMrYV2v7pNFfIKM8I
8c/vHzbaFpV5euqWjlXPxEPUo95QV3f2X/JlyNNsMUUGwGq0NDW/lByo+FiaSdCviHTBEhXqPVWf
vbZA7xzqjYqJpewtmJUzVG+TVB3rB8BMvJ3RbKC6/VZCGuV5T43RbReFO+BXibdG8X5f/YMwHEhm
Ik/cZrF2YHF/OrmFFR6scjLZ8riGVBwypAfl8qf5aHB33aer2jk+ccPnZHklDadzHxQk0Rsvh/y2
nRyWtqq70+gIyLfTMzZkWfWGw5/TsOxPjIjeu1eTMaPksQm8AJzpNh9ocMDyO3qaBD6EPrsYxFUF
mmsrk0Dt9hJhFJAZ2TArHmHJRaH3ZlCQ/fQP0KreqVu825fjGrdpiVyP1G8pHwI7ylbc18XfJOHX
10sJ9JIyqh3tmoPqtY54fuCV6rFFgGYLnwlB14xbIMDHJ0Hu1ES2ecLmpGQF2V0XD9RyeiR0bVOM
a8CQLII8ehzLh9nscqoNsx/d9SJsfoq+vDc/XHwfix+mibvYSiY0vq9nbFppJCvObonwhMVDlINU
vwZEXIdcw4na/Y0MoOmxUag57tBpcfUKXW+KYEyChnveekI5iOgvFQbPT/mos8YlTQCDbmK9/OOr
zeqtphjvuBDhCzqTeYt5dqOQcBKfi7tiFWrnlGAQMKXqRZbwQUw+AGvaS/jQP8j+dTC4WStfT0gd
3W0hnQ4DDnKU3bCBmVurqJmhwPXoJYqp2uPv308/ECSKYULTM6VJ1nPSdb6co5le07BCbj+6jB72
2Q1Nz0dJr++MDK/PZW4O+jQ6IyxsM1dL/2U8eH0Hhz0QZGqnCewqY4VjDCW7z5d6wY9xhuMZ2tfC
HdWLPznng+jDlUyVIy2+sq0qsVziXVJyFEAlvATyKv/aCdNLiXN+bNFRWWIhiK+7dbiitQmSbkF5
ezw5NbQeK1MHOEe24MEInoNEZZN5vwdvljMF+HJI27USEYsf0dbvSOuB3dGCFAKHcp7sPKaY8E5U
4rSiwg5iyhkgIgsEFnWVIDe1dI7GR6iu7ZNHNL0hNutAdnQ998ecfe3oeBcx/2nbM5W3Snd5VbJ+
MuQqdzUBECf6vZr7/P6CjnHbPeqlBdDAML6LE2r2+qGwPjazXW1m88gCk3psZZyTncsoGeS9E5o/
WXKAW4J99Zrl/pbZAf6MjVbaLO88HaUjI8kHnTaN4p4U+i0WzoNxnQ5L2PTE1N5eN9p/NPaSzI3G
m5ry7vb6JRQ5660svlWZJ4CinSmnedUizLBxYP7WqbA8QafZn0pFAtxnwcvKa6y8+vxOUmwPda4d
GVNembsmf1eoawTjT2xAed87CpYFe+V2KAQ1hbklVz+YMyjZzY/qvaDQQM07Ap0H76pJa/6nrhjF
vk+hoeKQLIJxwZxPE4QMi7WMLevJLu47N67wy31Qs3gIzIb4/fvqroZ1ZJ5idOXr+Szi1I8HO0DO
YzSi48BfKyoTgiAm6Dmt3HQiw3/hd4MEQFhP/sbRYjeGvK+JIWGiWsgCuabSpEYdQ2nIjgrgC/bR
aXrkkEvnY/2SnwbU3aRHeoYO2z+pHy1Za2uq4TsgOPw5Fa7MSMyy2Cvshsfu/PRp+NfmWKeZd841
VEuRE+sdRCgtMTnmQfQUj15FSn02lur4rcn6HCJcRxTIqiu42wnxloVXt70JLsSXsTS+yj1dIosH
gQfp1zXGDy+XDcd/t2zNWYWQsc7mlBvoOSi9MRTXK9KwjocKbxFYv7tDLFnbij2+OCiSdw4XJmGQ
c4zujDqO2XXDE7Hf+b/aZbN3wQYZiBpAervJUderMCxOxQXW4XQkbCXIzwloWkfPTzXCQJaG12ry
NWry6afn/dcT+GtYaeuCJ6gMiQ747wukGFqFtqCjkKKGqFi6syLMTc7sntTNakD/u82tcoItUBDo
Um3neX/NnA2b4xQ4WrHuchZB4/ovOyofYGrSir9YQ/jnwDT+ONpY/YSk1jlSq+JCWogA2XYaTLe2
qSHpOe3q47+zRxY0+erp0huzV/CO7bMAI+b8eItITpuLtTvNo3SoNPre+ViIf8orjDhIeAzSp/2a
PvZ82FwszAMOroC3oSOwgdx2MvW7s0QrybdwcVcHN8EK16IA86NfbHTPwFlKTUVR8F2R5OU29I2/
7/oEOTNeTDxYwYoidUT7mCzvgIpLLyIDYcBh86bzQon1q9LoArtO3V80ie2HbIp/NycbFqEdHINT
/CsWR1avcZV/L8t0ziAunG9U4Am2SphcjcWM8RD5zDR0oTRdOLEWXXuGzY/y92FQWWQtpPJDCWjo
CmzSbWv7SDLck46fG1yU6+PGwvBaIrYA2SYKZmv9gyMmViaFS//yLTPE8sKSAXQ6aZNpHjxRBkwQ
nsM/sgKw5gDsRfenM7/3YztTQC+i5T/heZMDi4KRuwRRU/YUXhCUKKYAMNMMoOb6u6evIi1LhhMZ
Ux6rYe0N27y1r0tpO35ZZyygdR6SGW+rGIrz+/7TZq7qiM4kjsRQEnSCrADHxQuJv38YfGrxgpnz
0RlwehdrI5zK//0oiwT4rte2AWw2v9cggIG6iyfG8PlJ9+8un4WzdbaP1rvVVL7HG0Lb0jNVcs4y
mCAOwi52AP9x+taKHzd1ubBa7QPaZio8ibGLMvuLdYdng2WsaXDnJ0oNsOe34zx1aHPCENZBUKvw
/pzkX8GeDTdHSHcHK7rPRxlqILXFtEVy1UXjk1eYsDZibIPGHPJQh7fBA3bJLoi0litWk6wPRyJK
XcJsTxh+EP1CeVZDeZtPr6+m7v6+WoedwYM07X2HJmKJ4vp0P89iE6MUgFDeKlrl4vvhzo970ZQs
1Hs9Kgcgx8MYUddG9Cukn3IDBLq48dmeujDKLcgEq3XsOVfssx8w/oEd1CjS1odEcXLx5GPYiaSG
r/HBbcT2ny0ItlWpPE5dxeQRiJQt5obnDHn05J3wFgOhRiMXF6hexqEHoq4JtgK3ko+IDtkZ+oCB
SQ/Gl+rZjQdRtR7IQsxr5IFEwYIOW6AAnhp90qB8yJceL9oIMsDCUJPbw/Dkiti1TfPTN1y15VFd
Kc8ZdPcjv5BqK0Fds7zPyuG/COmppYSMrwdWSWfpdk5F6VqFaymtHlA8A3+IjDYcehRvZF1CNVef
szQNUV013VvlJMl7o++JBsTTuW1ef0n603sI9gh/jnSTq1NLHbuulgI+gMT0oJCpHz2v4wosr/lj
XOKxiK/OBQWvvw78ODIoNviAc9VXXtiBJSPz1t8S64X0ep+dwlml/Vo8F83NH24eJ3eVDosebUBn
Y5RFCpmVhoyk35lZcEt6F+/v7+AtBknH2FjUDOcDFotONZbCQ7ckIbLy77Nzkhy7unWqoFU0vbm6
T3Pg1sc4LuX3G1lkYb818izFmHyPzQZP+BIJJRfgDCWhaDYcoW5LNVZR9DQFWuCSTt2+B9g/kX8r
KkC2UOHOVNiN2Cc+7BxG+ZaF4pBYZXDh3A5CHn9xyGy570IzBSwSM+CJFJhdsVYPeNOZ6RTcowru
7pGYMY9sptu27lEor91Ex2oXUV8pXhuglre0JhTI9fj3pcFjqZfriVZ5AwSE+TrwRoq57eMZ3GpA
4onkvuCmWqda/k8/5jbTwaV1QQn4wzAXd4ZxtIU/mKET4XPoO/1sIruCVSI7ztgGBL5SA4iXeYh7
6m3UzbxnOTRi5HQPCC8MvTp9ddzRPgMhIM9Tv1LK+Q25Or7Czgcan8iwajsDiyVWIoIgIKykcCYN
BZnVm863f2YH20fZCO667D21mZCEY5ihPhiYkQQpRi7dQEqXnE7ix7Vl4UC9ys7rS0MWarYA0Vnw
uEJTesYCr7Ayn0ib1G87eujacta+SJOHZH1sUU7Tchq48QqgOUZPiLjPPSMZnJQoL+ZIIowaSYze
GO+l5EctaZjb4/sJCKpV00RttuqBLMD/AZpUCvoY/PWw/jwzIUnYSdfJ6oiJwVXvxGhdInsUx8vo
T6B+9M3OsncxaY6bW3/FT6x5Dv+ftYLJl/E+GL7uFt/LQqicpdcV3eEj/oJYbmRUcKDsCvjks/gT
/Q39xKPEBlnw4+dmefxe3VusksKDiq+u9R+WhvfEiWhVceanIbstZulOMjvmzNR69D1JUc1rU04C
py+ZpGR/27LLInQZU+IefylnFIgAWAyLajCiFCfmXFSmNkuy3Fxe+MTKjLpSWz23Xvv52J0d4Ng8
pN2GczCEZG3EMlcrfFlC5QkPhSGfrt4vHF8Ea+5t+FgYEBmuVDentARBRWVvnwIMTXSUmiWVqn7d
fj+hYdOWMIa4piXm9eMXp87uNk2QinK4pzO77p4KhTTqZpdM5V/521MLlZ6vBZOAuWZ3WkskNpSN
2yXa55GojiawE1BEgdgaV3ZOnHB/uXe0jSCikBjvqyC2mTMM+H0FC1v0jh4uPQ7kFy+Ewo8FlqIb
GXZjR7meXBnqjyCMCveTl900iZ1q/4Ie6I9lLE65NP4SVvafXHjrcr55ltmEGiOcDF3mC8ZZzyK7
HaCgMPaHMvqb8VxubWnRDVHJp1Qb089KbS7lF1E5O9AOBEVwI7HIDoqpBqs0TwbF3FJMJM2H+Vga
MTWRPV/794X0oeVN2oA8rt9ZcsPWHjwHp9gwmrM4+6ISGOiT3SYImjCcgTO3JWekKwjOHI3funLH
1VCNwtfAVX/W9MuJ1pv/ifEVXyUsxS6jNavt6sLvarRsHbPYy5ySMMvISuNd54uCn/pnoQ2QNz8B
mfonVHqbMw+zXkdtZ+bgiQXkXnJV+lEGC0BBF5jCE/I7OgmRr9wo81LXf6LF04zO5MYX2Vm2iBp/
LQFetQj2QuhF/cAlTLc4txhwJ6mxtpHJYY/U6M37xxkJ3tzwQQnoLKieT4KP9vLmreWuB6H0GTQ9
lzSTmZNxSegJVApDt26hlnLjmM2yOEWqqrKIkcSG8znr4Y153d2ItORDA6pOikelIMCAsu5H5Gy8
hDWs2DIKJK+yDjUY6pdUETH9qPw/+m+NyhZcyZhW6TdwzJr+I6twSePR2aMYO6Nf+QbW6CtV0W0H
43BXWdAUj74iB1v/rGyyacHlxLGO6VLu0uPU+21sGC6v4i+xqtodiyTvYZGt3wHv5andqxEXbklU
9Q7ohGqtndQlYRpEuLOhGPgdb+A+OLibGobjFqXsgHqLS4g9xZRZ5knKD9kUW3AqEhxKaTdanOIE
KqH6aNLTP+Wgu9W+TE/UgQzLsQqHG7y6WIBj/oTsjP31i6HOWcenOoiVBGSjIO40L9GPPEemJKzS
/ln5v/UerI6gw2+teS7iRUwDhnrDHhgU6qYr1Q933aG+iFpjIsXCgdMDSAvTWIEp5ogLW3Jbyuzt
lXGEeUHXbuCoHBdWCmhmsojQTjgkX2lBhYzIj46idUa9ue5scY2gLedfEhkeE45XBMl0Jpu+H2Dy
5bjG7VoeyPvQyoHjCwva8rqINzws8mrhUoxxs4OjYGQRTVRlR/oEFJ4AJtBYYLBs/Yy/TpLwvE6P
EEa9JCGruiN4p9jpeWXnJKg8ttisVCqwIM7tOE0IMP4bFdK4opRxrWra8dcsFNEtdKUzWqslq9DS
j35cT4bbd9+bODaRH55Af34bBKJdQoSP8qJ52pAqDD95EMd3YlTxiKE/4k2UGx4n3zdM5P0/ht2Y
NI/PEmFFGejQZtdRhM2e0MGngzJcRdyk7SHH8oKqgNQtW36nLJ5yF+wO2m2i4FwsWZJnlrhfwjYU
XJmbTJDTTB+qCQ+KxoNGWSfnesJr4Dgrlg5KBAgcVqpsRtoWoAoNCWbq23Oo2nh3OOQiCQAC4IPT
HQptzLVFByuGPeU/HhQE6ANPXkRIobJsNDZhQKa8YTOAnV8r8rKphZWYxNT0xUoOVN3SRIu4pYKt
vTBGqAAsX21EVD9emXlZIG025sbfDHj+Fl8hOJANC9xW/kZB421OtR9mu+GoxQf3J+v3H2rmULoq
roiq6aWp+1LWfhRc6W25Qv+l9TWEZYBjmjlUQV+zqXArfWPmk2YFodoLmDVGIIVO/hD+O4BE9zyH
K+YgPqtr2gXgNiKGLuuK9xIbbsy181AdUA8VkrUj4TcYaVdVumyv1lSs77opMo8+VjekoggsYfGX
1J6OKO6wL21l4nXJzWkes6VSdXWV6x9wntkQn+RNa6YZAX6RZZCAhwlPyl7F/zqosodYLtaGq60q
EKqkXatpykJfOutxlndpOyoll2YjMlvo3Dl+UhX3vtjP16qKzQuO1YEXiRTrXumnYkAWL6lT3gQL
xKvGx9D7HfvZqODEXLAeO84dUUJxJjayDfRRlrzEjEvm93opi/AxXTkFJKrRHUlOHLkEh68SaBhT
PSyu6kED7mRxC6hrtiEC16OzsNA9+6Ou9f/lDJc3aJWdXRaoTEGPWXHXHorsAAAAoNZhAh0NYETw
p4hbQYVuYhenLPPTtnGvPWmeOtw7CGFseLIu8fzYreDQxMTrntAVefTEBOjlee6xAuvFh0ltQHn+
aj1oH8yrDepHdtz9YKMRdk2d3HupirSWf3c2oAmhIhxSMHTj+HUCTG9Ee/WDv+AVyHub8DFuodUi
YvyWupDAltbdFMIFbwJw3RIxFLpQVl+bDRGR2i1iJ4PGH15rnyvEvJ6Hjxbr8BwAm1l57JBT6QvX
+wmEl6VRi0CC0OSUb9S9qBr98Sx2hRrOpFsvYldhV7ExqmLXnk6Z6uWPG1vSa1y42NS6t5quHSIe
F4ZQuGBipWSuQQ42UrxV8fcvGvjosLNK0qzCJSyxmll4ldj6QaZx324NMv4NZh/HU3YxIKpHaz+s
nwFzEhi6U/+Glw4Jvuo2w9LEoy7vo7rboEZ05C4mv8CP4HrQmf7KyxoZ/W9NaR9jP+YjuTfmgVoO
TRI16oSjzC3GRELMryr0dUTDKwrgj648dJL0qvhhouZ11iFfF9Xt2xpO24Xg2AK2nSgIIvQdPQJL
evIAmXHr41SFirLIZ/Izc3Y3vLP3D2ENQ55p49YUn66gu1JvVF8au3xpaa6OnnO1UPMwHykxTRf8
1ctetS4ZHfzEVGD4UL6Ibf0/IjDae5u/dAivp3iMD10TtDqDjCHhMgfFDGDSLCJNVkQTRdvC36eo
sfqnzlZGrO/sH3L3fZOiPq5yDBgpRXnF9+dA3a1W21ZNc9ZdpdDLjccDAHxoyxdrleP6cj4SU84T
NjW+9+tQCjoswFyO3A3w/eNW0/wuY7xSxfUWrsSI68gwlPUGoMnVadXG0mF+N+Ez8hxlje86rzts
jwI6ZIYJi5hSqC3FosoXRTIS6NB+P5bGnvLGO22Sd7WUCwMtPJK7I/OFqQEYH83D4gOOkBTSIM2+
lSOQ/JCWpypz5589kGFLCfWung/ZHQPQ9LKQPUzA1Es4s+rFbtkpTdguCp04XJji3jFChspFgNwB
eZ9s9T/LTTIO5067CyKzEa6tmeGd6zgkdtADtxlLZCNuFd1j3/a3bRgVPAe/ehabYab8jeCSYFLd
/1+ZsiFjYc+Bk9Ef+4kOP/ZvDp8Qeot2RTUz4a0EBxhebdaiayRMYDaW+ErYmGSOKLM8blRCCUKk
uxn15MHMN7zaRW8CGFx9J5GEQDDBVYiJ/ALYnbuOtNXUkDPDpU/+ckubZ+idNB2O+kGdhstlQM2/
RYqKSafNqiJXOo+n+EqWqZWr3j1li0HnppHLjUd/Mvyu/qmWkD/qttoLanJoeab/yYM1a9xa2TfR
H7+7sZeckkBPnxtdbgXhxIckb+eYx5kZA9dMxpA9pGDrvyfBy++m4+NS8zAJG8QGr1abIxpuKpId
PBztzjeZGvUyNkf5x3hjBgJbPunkqtEEMVvewsO1T4VGkaxUcmKVJF0UgJ4w+mbZveNlMPA8RgA/
0L/ycxyOfWg9OgZhiFfWUgJh1qPZqs40FX88naNw5MfCNlvB3apOlsMc2ZmAQHKnhQM+wHZzfx5O
NfqCiScnyo2COsbnRSA5igpszmWiulUs19CW7pVHu1FbrDV17xngZWREIWT8NgC5bzG0gOPBhyAX
c/96klMKb3Dhr3HYIFTNl8ehegduy5nab8ACPjMOTXnUReEnqQn/p4ILMtctOLBdr+fpMo/AtAxR
Aa70rABOAnzcDBzqN78E15vsZb1v6haZ2QbZaSzeSyVJcYFqm6nrcV/5kuLjpcTdp+88kJcbAMRa
+hUBUpV7oqvorNw7z+6+bsTxVUbRWPnn/GHL5Ec+2G6oQMoqMoG8NeGrarQNFPqGDIcHq+x4bRYZ
sn4hywUj1QFFUi9lom1VGaYk+AUhzQuvekIYNtrtf0FCp5Fun8zkP65MIeXeDw3RH/vZWZJ92BT9
llIP5l+C8YA8ZAkbpU7ex4u/oVA6seyTO9qv4mbFz8TUiZoY1P2jfxHmnfrioft8vAv7z/VakrbD
0M71ClCW8p90OyK2oQfiJwVgGNNbHAAL/Bp0/I2XTyoR6jA5LvKibpiv/c0od9LkcCebz8FMi9xF
ietYsmuf0sbh3yc0BgRv3lHhUDpO5CyRGr020miDeoeNFyypleTOTIp01Ouv1TGmOYqKgp/xSVGm
Frou2xN8v1k9rkKv6TNYasoXN39NMwNJxl8lNKyRG77pfxeJ1ur6OPyMGx18pLLqiuGEnV8Gy82P
0yHNkF69zI9UMTnJzp2pd30xSxON5F40mm9XhIX445B6lkVjRw+CFBymOEvgbKt4Af9G/ACycf0N
t9QMWz84Ne8I69u79bue1tzieG/0zYQ2U0XbHAs1JLXIA+Oe75RlYz3OoJgtsm6aHx2J0dKIhP4W
Q0lalduUpeDFiQQjdWgLPIXzDPvW5BcQYpgtPqxWDPeZ/J/YPFF0ITZJBSKQf9/aJOsaxFLLKMi6
J+4efUMxipEKKb7nJZAv188ZmttiuL0czeKl4Xmu5oxfeuCVRF3CwYHdoabli5jD7Ij0v9KkTRT7
jGR4sT3YUe9i2aiZXTIhfJNcM6/xIWCi3G/twTrYnAydAAxM404P3Rf/v9jlxgvjKDJFmiuTBb3c
eV/4E5XFUpPBuPQN8gjixsanUFn8cqyvMJ8ptdx7MdLeA6Evoh8q8wswnQmm1YzSsefXy6Sf8Ppy
cBsA4HhN2uWunhGY99Ek+A+IGEkTgWyAkH2wkkviz0wX0sepo8ADhnbysvOKlKvMTfgnOaulgNLj
KtWVL2ZyH6gniVrKJEW9Omk2AbqQpoulovvpYL51ZdN/c4CWwjRUXA/uc7YYqHh+mSsqFP15OzhF
sM0utl8aoiSkYZq0xq4ZMFyRARj1+Hzq7aAqUlqkX/r8P07l7Ey/Cy19qFxVe33/PrWsYxejC75+
KDmI4rvChCBFCoZPeaNDgleeGR2zqFlCrtIqQ0FXrX7KCLX0lCIA/I+O4Q3P0wZvTmt2nXd0wBtb
+DFijFmj2ESaaOafFaAjvxypeNpLpCQcfxSyftI2OvZtIGrar7adND3/2n/EirBnI6L7d0nKKCzd
4V3GKzL0nXm8udunubAtzGDnaFJrzmvYCpV/gJX7ulbCVdL9eUnV5AmyEiM+a+qfUxukbfnMA+Ke
srHDFVgF9V9K03Wgka14NVEYy/C/ZDSJ6yFM8N3zxBNyPIyS3K37B4cMvSbVmVOq31wVl1JvPxKY
vG3O4DWuptgEC1gwQcTJZ3KghLYpqdP3/BINbVOx/GKRwCx10wRmqgv94Go3UIt2guJO7C+Itfai
/GoRZBLO7XgCjmme4w1fy/JXw+mK6xJt+02etXAAtiJlzsmCYT8PH727bt2JT4Sg3Igy5zsS1vVz
IFVeDdB8zKI4Iez+/Spj8+szMdJxdfyE1sn+2CsrNvkwb/rOktLgnccpc54XK25A5tMg67hbUm0x
CzEVbzEfWFPu8Vr0nLtQhn4MWKaMeNb1TDPuxMSmEXTRS49DnlJFfH6ue5hB08d2YO88Hu2C4Wiq
Z53J01d6zlRPxFZfCp8IogNcBSP4haoTyJvTw2b3vQ5TQOW9htFYkoWMMX3I4eUYwlRStw0mT8yk
8CTOo6qMBJpFnOL4Zg+Z5XuSHR5o8rMS7Bgrnxko71T2mGl/qKJCZVZK7s1qblA1m1mmdUu5Sjix
b0OFj9/jRDLla0P2B2kfVoekYavhyVQQdsfTq+ZplXPS3XImczqedLQt8QbMYIZ524hVTFg8Vg/N
LEWx6Oxj5TvI3qgsQ3qccC6VET9bVLuTrGJBPFKdEuZzlozfjEtvMrm0OCGEeni1Ac5aUSflzsHX
ywRs3PCdWz5JpGV1xeQQGGN5gNVdtMEB4DmPj88Ns08nu2EEADr0zZUMvmUaOfSS3z4hIvUMLSYB
jTrxmdyrP3RL4uGdpwBu8YJJ9haUgd6MRUuO6kMIODrnXdZGlOW2+O2ReydhXfN0G39soaw+w6F5
lBdflCsz+VptsVyBzc/ImyEhQ2IsxoEgJncuCVzgcD5WvTSbFgDDKm7ohbu69P3/CIYM8flrFkh4
3EqFU1Q1VbKlZlbzElPGIp/SPYsChJY/TrIG1R9pHl7p8zIOG5bHHfpL0PPIFyZ4d3SCWtp0NLle
GwDH/AReMNvTnh6ZwCNPltoi3Hn+ysk3CiYYIJoMo8xZhbnMIfS4BgVN+vRf5wkopgRurBtQbeTC
foj49x80D6gcFHBAHGv+8ifnR74vKai3rKPPKlTmsperzZp/J6K1P3vPBzXDz8MvZquXXvQmq2lh
ea2c/K8oi7HaMYZ79tROqDbRwloUS5izikZoBUSF8bjzbtyX+GkhqAdTzdj5zOaH4k5u5+gg+fkn
X8t4+pm6ga89wIFKxKHNoGE/adxAw95VWgWBNfookW1luaX5gvOb3EeyRcS9nGMFi+TLSp9Ye3u6
FxsvYaja/szPUsABr66KcKUhp02yGuMVzJkqpM8g4DNKI2bvgbDrmiN7wbrFoCwKMD9VdDSWBrDp
JGFcvxbDo8+vbWir6Df5M4GfqGRmWs9w2ESCoBnQoKknwS2Mr+K+s4864xNEqg8uzAcw3mKnq731
zZOWv/VqjHH5GioiXLPyOK8odDhdotjSg/8snAgdRUOG1E+h2h0v2a16bog4tBZo80D4fhX53TA3
tmKeRjgjHH0aLwXPTu0KhTYKrVtES2WCLEn5sab72skhvMC5QV5zv0G63ZuKVb57H5TM0+TGSb9W
fRcYCpUBO53xEXqnAX4ZBqMXFA8QSbjOt5J2N0YUmRyQAnAleJ6DWl1wIaM4fAaHD0JhqzpYk5Yw
+ua+irV6EQ/8C7tGt7NRovdlfDPLwM6H5+GjqJ8WsOwHS/CIXQvbGJlyYn4jdRFbAERh4802PxPM
gdVld4rN0xUCCGy5WcWP6d4DGQdBQOl5q3e71YKcJMBBMKKW1Af5Z0rHrL0hFV3KYvo59WsmI869
OUr9D9jvGBdGaXvYo2c50iOZNCgnuYmoQcQAHHXyugYmnzNJbgm5zJE/ceZ4+0Q4dHNmWITXl7ZD
7Ycu6VtdgSuUfurTBSUjBgY5epca3ycMjpE47VjWOpRd8rxZeRufHFQ6VjfR4IHae5x+jOMjN4zh
brAY1bgPFQKP/ln4gh503NjEMQ0I4A4e1l9feygmH/o294wxtgvvi0LGenexja8oKiDH0nkghNhk
uwowqwSGyC7zy1ZLW9xiUcL6/ZDWsyrOiqbrL5tv5CbM8qSKufeq3ihjpu7uhXMLFqy/hyejiUW4
kx8j4K5N4RudRFh0sPefKVXjHgnYwi+6+EEfeZfas05bJe5Yz/3bn9EDwMlAQsJy4GBWzPBzMdkU
iJKZ46k2fNrMSrb1uFYU5xQ+PfkXekFEPQVxF5hv7Hm7Kx9k4BdhtVYGdNoh1iGF53FWSkSdKN9n
KpgH5gkp4OYMgXE3noolKyXjjY7ZCFi2rUkcvO4ODdNmSsRgs2/5D0Q9BV1a9h94zT8sysVnfO0M
/KIXEiJhRGJdZJQQ7X27jCsnebLH0td7OsR0nz2ivAzcFwNWSl+WEsPfHk1dSnYjUriZ6vyJR5KL
/nNZbsYp6y0Wm6RR4XANFuqv8MBX5sNFkTo3rocLXXvK7ueCdnpZENwd0j9LC24DkZncG1MOQTMh
LLYKMzskaIfAt1yMyZIzBTK0zz8fduVi8UlGQOEMh9ojNYNajU0SL55FrBEYh8OSBnuT1QXuSsPH
YT0OqUBp2uz6ModOF81/r003MsFDKJec+OICbYdAkK4UMHbe7u1JWpiSR3/TVw9pxTA6gWuMd1/i
z9IQCx1Ey3mD4NJLA6mHgadVwD1MTVTF1F3l+pL7SCLojXDhBSxyRNzWByv+qVstytc12Luuxt1B
j5nMCz7P4sMA51XNvwQzWty+U4KRk48Aysc14jEJEsD3DDtiXU7BR1HnB+qSfhlgEq5q+C47IuoY
Kra90uXd3dDj+8VLNgx1kxoY4OCtDcgFAQ8V3GklqEvEe9tmkFwd/RobsqyF56hWUYNLoA+lyF/N
N9kOVM+w6GYqhuKsAGFh+fps1NdfRlpb2We0sbZMxTI69fb+JmXWxqNjgCrKIrTN/r0YemsiS/At
XpzyXlIN2yxsLg3Fe7zzlec1UQ279sQ35MES4k5ja93UyiMxUM1J/AcjgOheAaTalOc8pDa3IhUS
8dK+6JGrADprD4agGwK4geme2jsogSAYsnBdYNCcxMDDcWIAIGIf8Xwn1oBZATBG46JtSmHV5byU
1jG4jrpIvG+zGxygN3rC2Xkxtwze2ry737IZpixwq8dbH1fjYPg4h6aeDAFhmEnJtNg/LmH5auSR
jAFSfdKRgFsycF8P7WVj+/4onkbKDbCZcptaLGWi5n6BVs+d1X2aUfJaxNQ/yUnvBANRdgAe5nns
zn0kZoQmdUJX/yXdhw6Hj2JPtj5mM1obBB7xF/ou+tTVS4zGFXX3xN8nryayej3NqIZBDJb/OaBy
JNRnNn6dkKA84xfxB5HZ6nLIiY/vFJyORuFRpqhbhXGxwAOYG6O2KXHCPR2z0drKaaU42neWScbr
R9Kl5ln95mt79wyKi25a2Am6lzOLd92IH+6haXcBQsJvlzGcU4sVpAri+q3KbIrJky/ULmsePL8/
jWeDEyIy2YFe7GUqzgR81aYR0r7HUfk4GjCazfUfRT6UZy3kZm9g4duJ8UvoSXFdOvACw0r8SgUr
UjBe0hjJoNK3qV3v33UIcVv3yfu5h8Z7bwt4268dOIsoS4lTLvfd7Mah0xi3gKVNe/N3jtpMSgDN
fw6laNGWn2wrNgoQofw6+l1LOLJCESYH8K5z9x3Ozn5OfCjT9E6xM7Lr3XCyz3NZvmkyvjIch0TI
8b3jaJ4p7gX3g1OfaptsEId+5QXdGxgoEOcY3wS5SRTUjRArscpvTHNQVhwSsYzcSJ17/OtC6f6u
sd8KhHfBHahatMRbdJh7GqRpt6E6CiyAwQhs6aItV93vRrpX5SDRCeLpssEW5LsKKO0qLJCoYout
iu8lnurnACjWHjukTDqqhsbxWvLoZCb4UFcRjfyJgWalFxkVfsM/Db1TH6yA8iLYyfnzCaGjdM9D
oXFk8IW1VSXraxMakxuCBbr09KUhyAcpUEPGeoSHvYtb+arzijiOtEhI1IVPXJAqBLoU9aCIW4O3
UY7XIyvPQr5W5aK6qw9LjgpO/jLCM2N8/RDGmgBQWw28dIUVrEKwm7e6x1U3bwo3D7/gVk9j+ydx
1qVzBjLYeAo7NdO+QyG74uMdSiGxZA5F2VwUpoZm3vLArZ9nM+ZDK0jfS9FVDCI4n6lC2GNDFmBF
3LV+u/Dnskc+2l1EiqU53QckJ3DLbyEtdvj51qzo9B1+j4gMWv3wg8GWw//otYsxwYVtovAIo9xm
X+ND3ENiT7i9iQPnmCLK6Cn1uIHsT9AdqKP38fUoXNTGPAx9hNS4SpPZexuVECDiIIjsv1BvFyIQ
aMADsnmmrvo9WRkdWJNy45HpxgtpVjEN2nwm2U57uNnfG8q3Wd3rVda/BLSPNHlP8FI9YrN6Q9SX
TwYpbuGSvSwmh89gkVOaVoSJi+gZGis9jqX7jl5M4rZvP4xoOMVtCPGAOZpzqYiWDYyamTQvM5Zo
U3hB7qMgd9R06j0lwAfqUScQ4gEY7Bz4JcNwGgCLmoQf1OfLSkxWhJBM2pQ21MBiJLmsO8ziXMZz
N/KNCcyiGjlhZMVd6+Ck5y8q9LwhYCywEBaalK0Fhdpl1khKs2BeznnivOmvelL01Tx6/IO2Zts0
0OgbYsOOAgI8uDb+jUCm/ICeEdBb/3DbR/9lFDQ4mENXxRLSzDajL7r9kqOxroOCfSfbUf/KFOTv
dQzdKK8esBQy/AaoBqINcx+wDy8g8p3rnr5P6SEnIHmDqEp4vuscuD1YvIOENvYBVOH4AZHqO1yk
MINRbVs8TdEEhlubI7Vt5L5ST3QawdmMpTlp5OmARAVUcNVhiuSr6d83egs2OFrbhVfvnVltE9dv
1DtiG9/fURHXxOMdBChtUCETxhGD8UKeHyWFkADu5bkeOAuVyk+DmBViIIfvO6azEcy8SABKAgoC
o8iAm8q3uvN8S1eEzfuNMUfR/lXeXNxLevtCAXQ7aNTLWZzsjaqZgaeGsYSVSKF6zAlmJh+ZhYM6
BXoD3VZzn3eyk+tGsn5exh4uajSERTeK1Mov+/wMMvgyJ25scDLQ385izZn8MRyylFJoMjokIYJF
5BeIye6JUuhpOpVEd25RgvlGrGeO132stFKLrgplX1fZZxShMbHRIDGdKY5hcn6ZMnggn+ECLEDb
0gKUsXuBQSfiVJSryuVqD+rhXWDxpXB6S4wZPsEizhKEWEaeAsAxcajPyIFzdsLRvpe/FbtGOjzN
m00V9C7xtFu4Ks2EY9XIt9bNTLwUsJ5WkACjgxW3QJdnb8mIBcRXT3FYVdICUIhzWHrAfmkaYh46
DQNbMeGnDiUvK/gtMg1qMmgb9uTydxeQf5xH9a246K9jhXTr6W8s3VeZhaFngsLiRPlK6kPA5Uc/
e1fnggRtjkmB3AyljNZzyp3hFMIELOmhyVNM2D2lh/1kFjXIMMcwQorNI6xyu+h8ks0uCSvNUmew
CBfRSzqP9EzH3K/2RdF1qsA3ZAvFxM2G6QFHSPdobXt7x16G1jPprIWmkqlwXlNURuSs/SvJrrIg
dd9KAb5AcgcO3YO0GBuFjk1dnjDAaR0KkvO935y8eM/jOTe62UGso4nI3pL4cge5um7hEM8dr5j6
/AHI/Abqpctio4AyxeRwyxudIwV8aOJL06he6ujGVI+xWI7nUxh25wcQX7WmoANAt/mO9XApALmP
b4+96T1g+TWLPsDzj/0gUZeBcl+MeJXrKGZ1fKcZh1+pQ/nqH80FpxbeMcL1JQGu4YzsgBYb6b99
pLjGKYtLEDJy2ZBPS9OhNiYU1pDY5IDMizd9i8rd9lsqp1xICvVEUUnyy1ctqEQY6VOyI9c3+F7O
CS6j8atXu4U8es1HTCmx81nZ76eajDp4z4UCthDaLeioJ9WWxFaRwAbUZJHO+ne/1xeTnJfvG/EK
saw8TFKW1JKAl3tJrk0VMpraEYOqB5f8AS4eAJG2QAvEuid6tq/NWwTCITdgKHOl26gfV+wAqN3x
tZ6RGevnyeEeI/+rsRmZMGFOL+fzsrywqSHm9jpjyMyOmoittSxdJ1fgG0JajWasON8Ua0fdgGPN
ZbsvO80YKwPgnXHNJin+Al0sGAwWTeGWlT+BMpWDbig8iHqt/s1YlSD5ccWP0sRaLsZ3UWbdvsPk
AK226jd0c+KDn11R4kcvLoYIsF8FEq9VykXkbggr9ZArOSba//qIPKB+j2wPXOzFlFGUDU45nNzR
Wqly3Fu4rF4bVyusd2gp/562XF4KevnfIL/58btg8QYnSCwQS5XXQn0GYuq9KxDSZWGnGd+4mLRV
GmIimmGYZlsga2OVHMM2pmbIgmrHwOk/Vq8PUwQEf4u1/p9h7lP+WTf4uVDargWXBoGVIDqaT0ak
dNWrmrRdmIXC73255/vxiTorGUZWkNQSZ+N8RHSPdRJooWyw5vrFUkULOUbazhv1HBeA65WtMzyM
Z17vbqmzWk0aU9uEGuP1XJdbEMvQhR5Ytm7whv5z4GIOEqKjxnqIVhXNuMsEpm8mqvYXka6NDFFw
EJDY/TEHAhzH9iURxzuo3oEWQVnLEnUzza6O26UnbgaoD6/tSy7wJnPyxjjOATI2WP/KM9H+01Eb
r2Q2qLFy0999ffyqIb92NJwxtObHgj7zZKTBcsDW8L57+iuaf2pBbkGZeC9q5WOnv9OGtIuhDef1
qnbMb7G1jrht+w/jT+j6ShvuBBiTlfUbQe/WFV5ibn+Qn921vLTKynEEgx42SWz2g0EGipRUbSC2
g8GB7P3adsGFBHvXiaOEOxu31a7JQcVukDLsyJfqjWiEv95Hm2PHYVVdmX0ngESCkrJg0xy68amM
WlkF81qbbZOPFOUjSax8jlxfnKDUhaNYxLvmIrX2Vh1yQR5+6GuKnuwJqGf/01j5nc+Fz12Kf8ir
7bFyJHkggyHmvpsmyiQU/tVhIWnvxSsMvOIBAiUs2P8FqkGb824VC+ZnWByoXlidjd2LlpKGvX5i
0gDW00TNx8AY3QWTAa6xDgTt9XBiL+NV/nZQSKc4seupipkktOCH/YgQkLGeaFN4L5QRHJy6QLuP
+eNoKlp+qoeeqVJ5e4ze5X8B87A9qDEwM4e+C7UoIimKa6elHEWpCxj9oS4A8MiSoFNsPSGWi8qp
QPb0joxxdQ4VWESZa5WsM7JrA++kTHWzenhrD02s7+ZPvUE+CM+jrR2RF7KPuKrvVrWHRcqZOaBF
ReNihnRmx/0Y0zBdqqTak2y3EJxsXIGmk+BjrEiNvOVSMyCpWixOpN4okaj1rjQdIgXTG79wC9IB
Lavm5dIcYL1vjLflWPmzFO+IUa9FARW4n1DvqY4RKpUPtWzWZv1u3di/C4AJyJWpge8evciftwXR
PboDOdaS+xZzmZCGlZfjAN0Ge9Rks+jl7ezpgkOX2SYTNUtGD23SbyeqQdABf95dA6TMhPHq00gM
AWkJ3MAVDvF+tYWONwFUri6Oghgu6bHYRkihQ9s6p1QZ69SOCcxAALw0jkCO9D0LYZIgh9d2Xfjr
8RLihwbIwzyUUPFLfsrHbOWBOKKJwpuL3KBvdSFsJ6KQnYz7UvpBDGxmluc1y8tRjVN5HFzDwJEJ
n9LbWrgPxI+8hKxmYe/VYnn6jho2JhCuZMHfgpixQAOt/tuWxQ42sfDrW9/gnj5jLlN/gkdBTH3C
RznWMmyUhvYIVFvIPiu/CtqNVb46pIqB9XjSx2l/T/wfADfOaOVPEWruJFXmhdoy3DzeDYZZ2OzX
9tVPZBOy/w/wO/9ICc57roqRhb/lG0uuNzhwSizvCt25QNJDDyWzqdYpFbp9IhQVAHqhu6BKAVtk
6Hc+OtnZibr8TIu0DF7FbWjplBbVapNAi2Ln15efu17u9jnVXuBgjm9WNFh/AjvnamEgKFikWAZ5
dw4lC3g6NuU9EIeRSkHhYZvIweKnRilMxR0hTEq5Ik3wST41FjHd8Ftgj0J2G789e5Xd5+DfIBWe
lEtcHEHYcdxdg3EjJejiBSISgi7ACasLXjgXKTaGu70Tjski1ZkXOJ+E/S4k5Y9mVv844VMrgeVX
pXYEo+ol8qV+tqBpNDdNWnGRrmw3+uutzBuzpUNypN6/rqm6WGZELbNRZllF1OgJudow+i4/eDuf
N0ENtuinYHbmcx9KmvBtUk+ggNYpfhzD9sFJG2zvLakwciYjRja/uImyds687a6lO57ZQkVZ6kGA
ERfRuB0EGko+LOIyCTiMQX9m7dFslq7NnWY4jdv9eLnuw96HSiGbXXexcT7LVuWr8K3L9SEjf5Ig
t2ufDU/qU5QwI1v6IGLz/f2Rr+Z3CZqhvkx7GDGNwB2vi6F/GvNXERP5BYwJptJu7TK7Fxh9nxpI
JCp7QnBzxCo/DfpfkGSLbNIFauXDkvvdgVwdqtdU5X4lSwfnOERF0/IzNndPjqGlPMjT5aweG2Hm
1DlSjIKfpFeaemkmcNE5CwYaHS+fNB/k7xENa/AVSCT0KpDDuL+iY6G3D8tbefFWGQEL94BA6fbt
qcZhB9UjIVEy3HSkNYFGd6Lwsw3RjsJuRWpXdP2MUlq4HOeVaeYpDJYN7zXb18FqKtoyKUNH2yUF
xHho9j3OlT/QrO9VGPnVQttffZeQ1FEOJXFhRS3DdyBvBCRYytHKZLDlrs38OCahSUvwt/qsmOPa
X3BLLyXTpJz6E01QfEbuIhdsBz4l75bbY1sCtGEQb7AoMlFQ038TWtdW1TXwsGh+CbZyBNm+jwKZ
7bNCrg4KCCtM17HVMQEa65prqcgGf5zlWNm6njsb2yu4U4f/nvd1SrJ+2etn0w+xnJVS3WEZAGUn
sHkmx96dfu7fkbhWD8ZAKl9h9Ls/3sgwGblr6vTuLwnXq5eePm39y6ZtTRreXFngBKwsdGJCDP+V
bCDYFU78tGRq55Bmf5KEfEzFVpgYhmg/MUN8nF4YtIcCOmxrIzH6nojImN6bi+y7N+jGIrm5N+aC
sOTFVYV2nsz/jijPsCrGW3EAtmRbz3v073PmuLtoM10zvPnAs8q6dPfAKqjuyuLwV9H1BHukmyDN
RuJw8tcSNaAMLDucUy2LReBA/FPI0yi8eMHapR53U9JsvLiuHdQZA4MD4G7WgJ5mni3ZqZy7ByFK
+B9WiCUNKb73dLVHYdLFYBvXh3zO9pgjWXsiGxmqxcJ3M46Z9sRA6N8qd/7Np/Hz1gDBFgOzdSbG
k/PK47+XEYjd7lWH/A29DAHBU61byT0uugLuz+ihAMTQ9xl0psJwjCXjhPrOrbt18y5wbzOQv+7o
vtTO/rre3zqrx5U0yD5zqvHXvOC4qMHTitFZTpBbzJr8ZRRUTXSTQXDuoh8icXebnhcMdomgormG
DSV7Mo+VbA8zQyEHDKsLq2EI8afn5+wIHdPVi/w8HYkFd454FWrHyobGm7edfYduarI+dwDeY/Yh
bNEhchWgAYBZBJqbnGJVbR564Sg4n/uiUUw1Z3eMnd05LsUiMGC6fWhud9pPH3huqMJ8SwKhCxAj
JrbSddGjHOvezgERAiwtOZzLY61t8P+xWUFIkQvGBX/IU80bE/mnJ9V9lbRQwKNQ16VbJ5yaqVZ8
Ti/rIXGbTfKsCKO1GlLwuDJnST9KvoCQx3zLPk215cuGGlJFEzr0Agh4dJhaKnNX5BVWiR8npgDr
OBIVIItCRwMfUbsrYnfyC7YyNyJSQaIv9j+7ofXuVSkNRyU+WdCgF0xHIXyRb1fWdSt2p2hy8kfp
g5Nfi5G1KzwUEHZztbnfVfeN6CXyUoinBan2ENIY4csDKXhZhQ5cteH7L6G/bsqI+nizvHQP0Tzi
KzYBJxQbIqA//5lqSdUWMMdSZUN1ZR3aTFYgBLO4/fa8vroas+8/8VaqQ4D4RXt45FoPS//3+orR
ClJW/0I9g98VqEj9odUK4hWsaTvViv9pKU0lwtb8uFYSezw05JziuhJzFkRQabABItLBCXoRUqfM
eLVAxlI2Bt4kQ/CC/obBmPYjVPjPNpkVgBX/aYEgHbYzZ9HCt+HM8sTBkKZUMIzsn2w+zmSsbeHc
J4ZX//EJMhC6zc7UAnmBEk/3wAJVmV0ZgRL6JrPqSMcbxnCZk9BFz8JYv3LVGcXD1wdKcFaZyISw
zxVxxsqOW9e/PNuCbzaAE9cGgdnDzsb6i3AaIrfHCuAO24a+C00CwFMnULqZcvJGwaIs+8HTE0UA
m4X/AjYcV5t8UGCSAv231q85WhOklmq35xewI5Rep/VMQBFRfKPHkJwASBOe4BAATM8mETRoztwY
YppKgBn6Gi70XItyajimcL7S2yDJHRDNnMTuI7RtIuJ9M1TSGIcehHrB49iRJZu+k2Mzk0KetjAM
vzZJMSbVT2S+WU9rsiaoJiq/t/xvr+g3FVOs7WttsWGx7c+oynYwBv7piQ5MhDLcwgXrxCFUlt5/
PFjyn0DKwm5VM4IU3PcWpaXiymwBe2Zrtg8jBzbegNIL71L2jQyVeNDLU4SyG7Tkf/E1qN26nme/
+dI9cC3AGt4tOX8ONHh5HDAUs/oo4v99xh2N88zYfZOPXZeWrUU6L7ji4+1U5EaSUZL6AvuDnDGI
v8lZ4cj0k2AcfCytr1149e3HlcjDrscV+awD6JmIzAjv2NH9IpsWXVlbb3hxrwTG5ruCXfF1FQT2
yCPe4YGGVjwyFbab+rYcPoV9mox0qv0RFCLIshoUcQlsni5eH+ojuCXxelug1b3xcbnguPrbc0nk
rKMSypqIQzn85AZOoSfv7Nf0mzOg4DKLzit2rs61T99MkMI3iCJgrpa5ZWMOG1WjE0QxDV/JGr9e
CwQUddfELn/LGcn7pXcNL23FP5pmubVWq0w+7TYQY8iBX0qqTfzL493I4Swyp9mU+bf8HFECZ7+Y
9vX5FL+khJYyd7CBheRybeelXkxEQj8dvAZJDxkUzNTpH6YTIs8WxGTiAt7wpQrT8HqLMBUOTJnb
mBV/kiz+csOAWCCS5FPcoKsp3ixdxnrHNGLFEbgN47Ay6el2wfnLZ0qFZZJACZKLshg8SeDsFkcx
8+hnzwggemoUioX/jcNSwCZqm22O2sMm3604wa5GxIAHLSWvpVsHHp9V215wIuwcLlGIi9/4Gtzm
uFT0uLNInmdQpcG/pUGgwrSqzxZJWrkxJQPxHIz9tioZVjrT57edawQYTN8IywddczOH1A5M8W1G
JzEPZgNO73aOy44Ja3zO7HG8GZ9Ce3rVZ+vcQwSLUADNji/DshxAur60iUtLLfw1iC9lfDxIvQa6
+ZKjHwNXuY8WD1U6t/U65fhjLY1WKJFklFVfwk8IpQaW4ywL9BOaVnu5ZTV1HbTRb4zoGK8oSIDc
s4M+pe2kB+cqAX7/0vVMLnwokY5UMyW7KNfQ9qXrlLIcqsUu0A6JfHG8BeNpBI2rbAW69v7hbKnz
0QNEpIwYWu+CuNRV41ka0azJD5VMom25tPKKuf0QC9591o99vclByRsqzIEP8ZhpWj75WLV2Cu5c
EXnFfn3GeqTcpjtTLJsYEazvPZ3OffW8WQkv+VLXP9BVLy/avxZK40IbwH2Sc5h+fZxeXoLqfjjp
Yn7vvO63EAfIm/+E0GOb1kwYcNF99S9Iz5TlUfC8CWiWgIKW96HzxWnNN7jiDf8kg2UZh1gFLw2M
FLqOtVKYm1uWmEKo54SMS55qC1V21lZw78MegEEe0PdpIzrsS7Ka6s6gyvboD969BPkmMUYJVwOM
nqZTl8jKJOY/+tSvY662tu041x4wLBnH+B2NCD20EJfVPG32o2uurUHuK7zVYavDD6JedhnSNk+1
FBpqhrPo6OcY6NhdqDQHRedG6F4cm60rhV6EW8Ybpc/QUcK4zlOmruEubyFi4tMkGiLKQT90DVRc
YJ48130nSbt2TuMUnDLzhWvL1PIr5to8SSYuGGntUgOaNNfbtbZxE3QmEV4KlQq3HxRLrEv4z1jI
r6/QOl1HN9Lz4kDeVQCxq9zxPe7f2dklxbQCfu6Hj/vjKMOZ1V2OGxehyC0sQzmMEd1+C4euxWgu
ZYfhYJPADY0sRqQILe5KZRBMWG8e7Tj1aUcrKT7wGXT6DIR6BSPgL5AbEkilqru4Nbh92HC6Gsum
18LZaYD8qiU2VK9wRDke0JxYgMwW6mmlbNbTOBGmRWkCB3KeYYPQnuoIEjSF1zfM6cKbV+1ggnAH
idEsxr9AydK1ENMeVhxjWg/0rPa/9shKu7qzv2c4qO6jwdMwP3yOQRtQVBJ8zFgXK8kR7tHjuexh
ysHm5f55EZr5EhzBrfE05299x9sRDgTWDzR7jpuR21y7DLkOTX8B+WSnESMxs7APtaifHyNfcuwl
jXjRTOTyNuUbit95w/LrpGCTUjje2Zr38aR5Hb+oQ2qFjLAEnPJSBrAGMIU0rKwpkx3cw+u8hBdB
o6L3vHBSstiqzbxJorb96AL/C66fAvA/j/r/jn9lY5hoPaHFuqCK8ES9FCGJqvHmvXLx5qcesAyw
k6hO9EytrwP9l99GaWrZHt3D8msTSlK9Byg+3uSably6+P5dGBjoexMzKUjzSJnyVEkuj4DDdx9l
6KLgiV6f1Bx91POgcJCQd4WIuWZXgmmiOIisuDZBzHN8SPdUPpybKTWemMVGlGV7G8wErIzpBpT9
UWe6+PlwaHSZghwNXH8oQ4sSWug5Pzudcj/NkWxl4Pn6nMYgRAVkEHi5ouCeSgZbrzSwV2nr5jct
McCGSrrrWQih1/LQrdVdfK8k7l1VoF50fT0FUnnT+1LwOB/Ye4JhdBepCB6XRMYNSZETuVm0eh9i
3gmgDjIQIvsYR3vurLmqvcgUNb/jG42KUMvxRDsWg6Dt0Dh5gp13OkwfpELZu0+xF1eV0hw9eeWg
vao3JnZdXyHufU7nfOTXr7qBD5JwzdFZUnIHA/76MJtgPmM9oQy5BrSAJqXR/uO47Zv33/imniPr
Si6TkqrDI5y8D8PtMbWCohzdDrALAucCusa6KjaD87sBJY0kH6fl4pWbgrJP3Cua2T5T2MXbLzv7
y+tqMWiFlR4eIGIkuqUKqrZVNOJep74n8pr6GveoPz47LOD23g8q121ljTmhMay/Pk9HnyJNfyzc
MXxYwn01A2G27PtEW4cGvUYI/3CPHi2MnPkE+pSz4XxDEdfAZ7rn9dxlrR1bC4b8gDvhumpb/PkK
GaNpHmvQtjMhXwqUcQfWPc8n7UOwMiu1DC5OrsWUZ6cXQlU8yoL8PWJA/u36eQgxnpOB2i/X60x/
qv0lusPQBMldaZ9GZDK95B+kjh7iQXcRqGmyNfNlVAlrEZtxJ0dgn5ceQeD7xw+H/cad4RfAitwU
ievJqj0bbNH2kDm72vNvdAeq+RoQlABGKh2jF6Ceykxtfz1ATdSVm3OEHNYZvRnUfcXPxAoN61HT
TlIZNB5qPDMH5aWDgJ5E//hQaXKklOxt6jSlEFOB4/jn4khjpbSDaZzhhdgU1pPqlsDUfFFa6Q0m
G2AgCdjldmu8MkuYR9cXGuE8dzOTxK14e6m2nBpN67//PBH/l2xul17W7prkfMua0G4oV8s9oInz
VQRHBQg+DmFXsfC7xzq6UA4FloYTBE7UY7jFEakduSBHhFs/JoUUNXOvwm/wHob4ukhGy1EHMjds
1ESjvE3haBr6wCe9wSPZhOPkEyllHCOky4Fd2+fLTBYA0oVWLUo2de1tCJxkLKusBS0UUvsvwL75
UdBqagHvgS+vgmSYin5zyBSgWG8i2glVwjgVhcgxgEkUo5lAvvwPP/S9HN/XEczRHmgGGZnKiPnS
uFOYK1PbU6UClo+X5cx4H7c4RCCMFBHXt9fcsXzRfNs/9qrinjdzS9RaQuEc8CojSJK1KxRbXQNY
fNNG6EG8zn4aiow1dWKdp519NFOZoLCWg7ObZVaCmoo8lqP/uZimCjN08Fyejj7NEr9LCgckxzJg
FmOVsF2mqn8FIUiodbhy/+82MsG3nyGbqSK8ssFbU+l1kpLyLDfNAeQ1kSi4JfgbWHMHN+d2aDA3
QozDrcFtAMw6vBvs0ScdFUslqdR2ylyWHt8JnLF84kA/gQZpd2dufn1Z2Wm5LY1+plB1Ay2uZUOt
+/11tIkzH8TW9ZEca6zVJbhgj/oll1mBI/BCiL2+sa2kbqN+/1feMZraulq7WFN/fpdlhxyPK9ti
DuONyk0ivie7sWiLLE72O7zo7nvZZXav4Q/A66GX6Imo3gK0JusdX/amaUUVyP5vDmdF4BjihLOk
Mcb+QsE1yIV5gDU9EpL/dN3BmauDVbHuOou699idhC5WCvY1FGDMj4mgZgfq2qFP42YFiN3z87z1
5zLKsOi1B8OlN8aNerB2F37a4ib76qJ+H22SAU31IGDPvNV8F1YnvOhYzLHoEr5F9nEX8PTHI2Z7
nfTyVAY3l5zZN8NMOqfB5ibkPW4z2TsjP4sTdhXE6LSte3AI4gz3XjvmoTH3YfwFbqp/dM9NH7gf
TDr59PGf85FOFDLkNZrpjY6oCbiaTBKByktMnJOXcdwwLO1lQTP8AtSb+Dkql8weum+Ib0OyJVpi
mexH0C3db89T/FSC2960U1mgEbzCYSHiXcC8XFq60+mnWJEUqYe/CnWRKnsN7Khz4zhRHPqRC0NP
RCFZnbBaK8tfHU4n7JsvAFLYSASd3SpmI1qov5fJUIwZwjaP2kN4E2kgZSxe0ie1Yo8NQ+S8FDYK
Vn1XoaaMQq+t2my2rtrrLrijrHKKSaIbeTI9JJlOH7y57vhHqc3/HXhqBhv1R97O8AjMMnMTtXWJ
MrOkkvInPjMJgne9+bE1GjO9bDviz+apYtgskXBjRux/uy2bXVuiamN0WUWeq0qu5hf/FihMpEI/
131ohDQKtISaY7QYVqStySpLElDpd/zU6ILfhdYm9khR3cM+VX7fbHz9p8pMu8rSK7GEDwtHGMEY
Ow+fAMcoEuXds7SNGBJfIDnVSmNvG+Ttx9wr0QYE+jmk7e7n7pMp+W9xuVOamd9cL+S3p6qrupLC
W3AN3mfxOHCP0ZoIBolSsxpjtiPazHOtDLNAKcSnC1TSJHgsczI3tg8RZQ4Z0NNg2xeEjWNV/OxQ
yixL+wM8QYJApdx0wjZGypU0LvHsMDLJkBc9dbEytDKIFo7FN35QhhhXCrqkWW1237lLxYkX5O3O
TFwYwDDESpkzwNzFJWkNUp2QxpOppMobrhQ620/KywIGbBRh3CUZoMwBOHYG/F/vNoOhoJwDw38w
QU9ZB7kjfWYnMpVXauEEPluuK3buzxZz3lSQ2cPET1PNB0eAs/CzAjR5rFMoqU7DdOEqBRfMyhN+
4noawG9RCAC9a24Af96bfuyaWwXD6DXxMvSU6WZStgVhbIGe6a5BaVDk4W+M9coPHZG7id/VDV8z
TmBmqYacvtYNNMMCzpyXOIqJXK1PGUv5tzG4WNtDTsZQGC/uEgIUUY1IYx7RohpYZ46DziUKB7BP
HW9qbxQbPrbEI9I2TjPFO3F96422ioY0gHZ52YNKlWLkgcEWS8CT4ASMcddIE/1dOvZ1t39unCBD
Tg/v0zAHvfLjbOD6LoZEmfzP1eNTxznRopaiDOhrEp9pPLDBlPeCHxrf5iPYESg7pZh6IkiVvp8l
XDExRFaM2/BOr//Wy1f38TUXhlJaMJTMihKxEOWPDSZwQcOnpcjwzpCkopHZ1kwa1FSyk5o6wGe2
mEhVNbqI3euZLJOZsoR6bYdyOP3B7Q9JJ0fukkWZ2duxiSC16797Qu7wbA2T/GQxsFoLH6AC+mHE
TIDKXNkkaopua+R2rNdXEHB46W9vEFLQg91Si1w71Qhu+yJd+byFbcgKfgnx5c1LrldKwd4GeHC8
2TGW6oj6mO2Njs3iTtidjagB2D+8K9o2HRZHrb0/tRr5nzxwFGTVA6eGNrY/qCedabEgTd7Ag/lK
Kl29GxI+NE99CoVDK6B5mzeY8bgAbm6vDgdNIxiB1W4u/oRTpIeKWKCaKYnsiqh5eBHbLk8Ygx7U
jz9iZgB2qVMIGHE3UHzgUgd4khVf1hZ1LiggiHqKXH4lsxghFd77TR+NT43rRVvyn7a7ZeGaWGpU
CPT43/FnWkpqS4jPu9mXz3zcezEmpvL5twzvHBDb66OX3+EfLXES56i+R82VOsNG0kUUtszjswpp
dZY1PN/Y3cTZB22ZcA78imITKWZatB1XozpfpPKD+qskE4eFaFUnM3s79D5PvY/JhkdCvKE+lin9
8sgPcBkxMd0zTgxLNBI87ocmC9cOa9sElX4ixD2NEIJaICffNX+o79RFAmHfttqhQs4Y3tjyccWR
SqBmqvu3hytx2oaNqwHnXSTlWmwdylvX1YrmQUohYueHmvhCvK3g9p+gKI5hZUcUhQ7ObBjtUVD9
F/pHTRRFZY7LntwhoT91aj8U/dAPYZ2daglQCjoGEs2a34RogRbFnej63AVWaPbfK2oGABbP6m/3
HMfguo1hU5VfLkcO8UBgXAyVtb2adHbSvNGZ3Gjd/neYwfDhfwFwScpmc1po9UNGXjiVZ8mW7giS
gmnSgFxey/S7snHbLxVLkf52jsZfT4kc93FLoiaJpO2Lb0cW82tuW6qvphS6C6yTUpabLPnCQ9i6
EDW3sgiG7e/t4QOmj87aWICsS7e2TuANfVYfqE3ruL8vzhOOxYuIwcVyLimnhRM6d1q1IVHP94m+
YggaNqlMdZVijUrv5cRM4kJpxYz18SYwIZtFBfL0R6uaL/ybNr+Q1kFW2g/JGKUpMM+iQtyBl4nn
ErAwx5NvzG8wIIH0va0Mpjouy/a0O3Q/pUzc8xAhdk4XPivPc6+IqR0oBBoC/B/3cUPovr3jL8ob
QOoxdBsR1/gazgFz8GHOTV6TmranHHd2BhOYkkAGwbQyIPBSUpzDmnMQynfmXs2fM1FhDVzh4Ea9
hP9SQoHhXcmi9GdPMc0JjngO4F1997ADsm7WVT7mkVo2VJ05hZyIvgNBlobWrZkDWIF2F2VLi1/X
7OqQZhwKX4SGXbK7W2NGSbLoBnOHd2EkfuRtwUoYWEjrmo1Tu/r8qMpUXDBWXmpVXyusZwW1D8/U
QfUcbUFpBCvzkHHKDzInqbFlsRu3fkhtVqa+YAb+JmIAjDMmuLUdZUaPRlpHKqewdtIvG8xbKUWA
uXRMvFQ5y/4uEZoSMsxH8haaRp288aczsS0hOe53Zz08yhX+Eu/h0zkOthjuYxr6OqgrNkBT2nTf
HnaZa5UlUc9YF0rTkpNlCyQkOprQu0lQpr17NWJGcvrfXinpwzcJ85fonB8aTZm3oHzhSgHtUHJj
3AoXaz2p2NrEV6hOyM6AUlYCDv8E/EG0Wa8S2NH5PEKc6cf7QXJvbKEKT8uMhRkLkglkarMn4bl4
O18fh0tlrHO0RUHeDXJ+NBXVeCJAO2HfUzhiHJeIaC4tdENy1sAFcx+tHFFDba/KRlvi8ETy0Mtb
hC3EPrDL8NWNuq8TnWU6f5+pXnXanmPEUcVv6L/e7kVlqPK3hHNzVYar1E2NUcFgssB9oV460TSX
03khfefKF4x1I1G7/AUcxFSs9e0+N8UnQJylHjAhWOfTrlIXrB061eMzyu+wXo1hGwEZ8br/8H28
yP35DmRZqjuKFGoUh0chuqplduDQHUbOCoyNDyPGcNiO1P0tHOqM2S3ndA8LAOElQGuSy1bTrfbF
xOQ/xJ1kMeSOtqkEUaTmLHfZ2zQIfCWZoWMFQcj0/0cFTVHKsfRNMLmDxKhD24KTw0fripRS1qVI
e9L7xG/8O4I00kzynslO+DLbYkjB6dFiUcvMbkRdfWzAmxwOdTwUT9FiHaN7r5o1bs/6sxdjTo8H
B//kybx8YjUWdOfT9B27wzOOIO6Cfq2FI/wUrcxiqOv/XU7VOMEnp/5ip6oXFylNoX5/fG6vIrDR
JSJTwW4Hcr2+eIp2CdBv8xutJbnfebhrMVVe/WplB4djrKeZi0NBJPEWR/qg8+BWtu7/5EAd1eLx
4fK2J5brMfQOne00gzQ/SwrZcXnCU2dYyFBbeeq0HwpA6BnEwoURlIP55p8PKp+fZvqZh8y0fbXS
fP8u89KeLAJjFqSBxzLtekguHh9+7v0pQYXdg7evUp6WJm/p7ldlQfD0x74ofOtrmYnlQEr+lyZV
48Nl9bQiLX5BGhJRkkiNeTnJ40edOXVdHzN13s9wAllkG8hKteKx/bpQSBU4ok9NXiDiAwoXDKx1
4qKwyMCiC7i2lr1teHxnzV7sM4ctbcfvRqDJnMuaodqggkr1PXUxOJO2QQhh2BGaz6rdsi9pVZwH
14b2k4Vkv/uVaZ7E7+RNDQl5d6m3J+oVzt9caJsH+gZFu9JxsAk9aX97FEoOiIWac2uZ+l58Qh0w
L8TI1vQomWZHd5/u7r3W1gGiuayIIupqA7nGbEjPPWPdSv5OA+BGb9suo0dxon+k4tP8CKLT5yrb
V038MqnP3ysbXnQYS54W97UI5WA/gtnD72Tq8c3trpnuXpmF0m0JsjXrxXhdT40VKLfZGmvRDIR7
q7kd+W3K5efG34epJQJPg4sBqdvzpIN21eiV2+qehBAPmxYFDPfYnLDTgyGmw1jYVOnk1h9C7oRt
OyKwASkBv5BUtAi60Daw9AcksQEPtXVSb1OqxMXAxGN3lnTm8fs0lCPh58wU0H8brK+/V3CGQ2sp
kuv4KU3YEdluHfHzXAVSWD/qsd6M4k7Q6b/sr0ZqSu3FRGmsg9QHvgqBT5BVntwihAb5uloa97uo
Dgu/ES4ZiiyRQLTDi432wC7RyyuRjO+vJx/kywj0Q81SIo0wFT/Set8TldZuQ0ebhdlTLVHUoPKW
H75Lif3p6Zo5inST0yFfNfJU5evfvMeYw2Z5g5rYJzgZf/0XR5nqeDVEwK6muxuhTR1FO3LbyLK7
ypPkah3ukmoaYZ6VW0i2ae4wwx239C6kSP/dhzMTujDT2RLow4vKhh+y/UAMZcZbOd+8FR1Zkv+W
WOg3Xnfrb37YbdqvV69kc8ovAOZTD8lajKuxnqxcy2ldy/tT0wPRTzW9FQoN8kVWbKoz7/ODL1e8
3bEYhoKOUfiG/XsYkDb0vRuvAvr+DNcxtYRa4P8fEl4AhxrdvgiNqdpxaoe10X20rFlifkl/3mRU
z6nrOKBdx7uK9ErHY0EorCgY+SKtaR65UEMLG8p9vGpWCuncn7TvRratadn6iozPWWDfGRNROI59
u021yY89WDkdbhBI5yvPMQ5NtlQNBU0YeDH2w5i78CGeRiBEeQHWkBeVxt/FTWO2FS1WffL3nS3M
59ZTNqzGPvmZPsO8GsI6H6P9KBFybT9b/FHTTCPVF6GNSbphDJkOaf3ShpAq12Q4NKoPowfbk/zE
JANSYKQRVq/hC4slu/cGbs+vr8D9t86NGOKKIN2qeXIszTMVz6U/bZ7GTg1V3Vlch0EXaR8+E6fl
pEhHQHQDS4ndN5dkintYkr6aV5QAAxbwT+YV+8lpsagEOorGhoN1QqeL7R339uZ7eDfFkkPc5lKd
9m69iRUVoh9GlJ0tWKhhpxHftWGy0+PWNqg4BXo6uN3dEMsfXnF9VcEGSTTeBXPIfRfjAlL6FHzh
tTcsLEUaah8S/b1iOPt1NN8/VHaTsIQqYiMGzTfxTOzExoi5uXCggCMXGe83uYvPk4iWO15s2nfH
BNJCXl/1P8sLOQuloejXM3GYqaWZ/7duMxstZwgUtr2EiSn5jYRiPDA/bv17hB+zudwMkqWfz7AC
YDy1PLt9VbgGIlRXOPUMgNIVhDKjHsR2cvm8eCDkZfdzaGS4jKACDfFgPvw3/19kLtCDDVeH9AuW
VtIz7Zncg2DxZi/cNBEQdWwmbOYOF/308KbcsUjr6vYF3UW3oB7jpQRb9ZwpfQleE9YGz4xbGa7C
YmCSCXXwv5UsZYmqmkZ45on66uKzeavDo+MZfAf4xdyLpCAra2OE65ejnP5FPpDSCWBvMKXmTUy/
SWZSXJSeo50tHM0ERb9LqbPO3snDh87ocZbGx376skYFgmULH2piq4T6n6Cye2s/FTim7Ka4WJC0
1nveTxBnxMiTkFbiyjmz489T4oN5LoL5Myx3mEmPs4fqWqKiI+TGMnkyS+0dTfks6WfQpANPwr4Q
rG3urvJZ5AQhxJh3oODGJGcu4/Fx8CR9xJNszQcJffmFAL2VDiJxmBfngYNOrhFgTpQFyd9Ichug
7LNGMydKkkwMDaskETiUbLI+fSpw3/TdCafq1bRQrdOR3tW+ymNPLM8rHU9ww3j5vUn2uwbt8MAY
VRiG1BlNajG5mhItOqwH3xtw3vONhNZzoFLaQ3pl9XhTZRb+Q+l+5Tk6LFpXD56brvYuXDximuLK
qY7xNA17BQmw2rlAKmhSMeGPzquHdqukmyDU+hMlekGznifeDb8sFsfnbKpsYRo50q42NuhyD22j
zeWxY9qsjYyRvKmwhUApLBiEgEq4b8bw7b/oQRGhK3D0SntRCITLsX+KTb7rHqwE/K3qgacbsgnh
3OX8Xc1XZ63HzC6cj9VU4xkBq2J4EEh+cZh1jGrJbkNEetUr8LE7BQBcaCWTXp+/VPui3r0pJ4fP
wzv69Axv253z2a4NiIscs9Z2SQF//JSBhRu7ulrt8deX/e3S93gOIORQ4YRN3Mh2h3+6/SqLuh8q
SE5CHAj6aa4VE9i1rLcH/mSKWeLG5VcCf21bAJYHgwRmQYSachHl/GDQaive71FtV0k2VlV6dhix
540tr1CGW36NwWcHgnd1xIeHpSNGXOWxjcqR73BiRMQaMjpTXAlp6ztnMwrM/ErGsvPxNoYz/bVn
TBOHATilVvSAEFbef15/geSsRRvjul0ip1OVshmfFMp/0WhU7hYVQUZ8V5R3/5oWgoWfxMm+mqeN
SFysEf/LO0Bt9HtC/x1WHwWgLwpUC61rWnjLGgqR7QonpK7C/BzZ30MQnBqfMh6sRDfkMJ51JDb4
hMIOHQMCemxycsgBGtfdW9hWUz2GhY+EZC8sZTqdB6yobw9y08jdHdPCX9qKPNUBf2DPKmcnqEZM
HK7lIuL/9VIh7t4TXLuWqs2eAj4DcAyApdxKSNPUxaWAwHhjW0KIZ8FcmCdDiLNeb/rgUO+WJ6jQ
U6Ab3y1gX8uD9yZ+hpAStXKhbatsiAaF/zMI/tRFIhgsVOFCt8n9PKw4Nbj/iaIlBk8g8H7Q7xaW
/hv27o23HGimGn7MquXpQK6GMx0LgD5TFME/qgRYg2mJWxdVDxoFwiK0IJ36dSW5zTJCjW1xfAKI
2miqFVQ4FnADkjq2KyBDXn5JsuiuRCclZqMC+NRYaaGuMiAX8Xhc41pmEVrNEarUyzyZg8csiex5
u6TeVE0keMpZ9tbLULdGpiTitTWkLasV6WVNaR8d9rhZdLhxJ5EDlH57+ksTLQ81i5rnr02On3h/
IMquVN1venxvyX661HrZODsO7d1uZUAdO+J/rJ+s8C+71Otz2G9PwCxMk1OOIgbMMfHbVEBO7BO/
OyhEJGuDmD3LymliUEII2Ob34ZgQahyPQiMzbo/cV7sr2almr94JqzATz9i6Hy2Xh/uFojMk9CHu
tIShxk1wQ3oAjfVWExowbsqcpOc9CGhEmPmTGcZImhujTX7lx2d8iqX8K7nx0+Pr3BjRrtZX00Yq
qn2VB8Fibl3MrcJsMSCvwgkP2wE3Ga3bCRnmrIMUunJ4PAm7I/B68TUy7CxP1adNoQ4Md45aNNT4
yPxNsD3CaTPniCkx7IHaa3mWLqFPcRvnjUWmD7SMphLSbKIksegiTfubvpcgGsvLt5+DTkLRqBxN
/A+HA4Yhi0xBvegyjp4ETjFGXYFV4nd/AG65NyEkOhnUkxwQmBIzix18/gh7AJQCbnK98Et4j46M
5QItqfTOrT9ojQoiMXWq73rVUv9FzUrGnuWtbhGycWwrP/AVzlBTh0mjvqAVOn2RZp7BWaIa2y+W
MDHApKefMqFvY+obXTLjuTOhd7tfEE51c10Mb4kJuu7YAVvAu5blwC1uJ1m/obPHyuxZSk3MjuRQ
mXeeR9KiEHXPjAuuwzoLbOtL+c6gh9GHa53hCoELGxErxYcqkD7RRROOHEe5eDnGrI2GgtMHNNsx
dttXhVzpReJHwji6A9iMS2Y68jYGcBHllySN9sDebUCGD936FeYIAp1iW0khKLYSIHPDfnY0QztF
18GxVOLbIPu03FlPbZhTA1Sail5A0x3qv4d8H2RXVHHSiTAA8OB478s2qCuWth8USCZiVFRYZ23r
f2DfkweU7kdH13FItBv1MfBVh67e44+6c+wefpE1Q8AlB1YkrTu6q++PYGPoA5bAnq1wS98/w8iY
FU+TudpqSO3SOQVnnAWo7W6Gq6/1d9P7B2dNePFYe9DPz2BnXd5jHXlB2BCnTyIxXbER3Lf485tf
SMer3GKRWVJ5FkdtfovcQzEE2d/828pqyFiX0YwqBxV0XRs68Jeo+iAITJNL41BA7C7YUTsMUtx7
ELIaFBY+8HuhMFaKV7p8Fk2zJ3vSJ7h0j9CCvYyXyKm3nDVydXB8WDD8i6OnvIR452Bdsd5oBkql
PA5RyCJZgS00CKcX/oE2z7vgPylszM1PmLJ0MiEvv3yvXKYPSyeVZGVkvttHJ/X4JB2eSNlVIRQz
/VHgWK//FXRbvSaW4N7s9MIO6hBAWbvvkNApQDGQyeAMmuzjL9w3MKgL8QVrBnGuJ4JMj15uyVQB
sMVCo8u6OE8smdIL5aZ9A+/MmqoNVHKIRWJGP34Z8k8LLvS4fDVT4bpDhTfi8DtRYn0Gz3nbT2ak
UBfAENXeksWvQ/pqcgoaZ7dBrWL2rwZn3WyhOlMV2O8sFVBCWCW+Rd6mCKjXDf9fxcffHN7KOGhU
t6KIfNvjOTclSKBPO9YeINhTQqYoKJeA96hb47e64CzQsEGDkOVs3wF+WFAjdI1MWiDfzaLy+z8i
Tzz5ex/ZdHDj9Ul0AwiKdWG9Hu923kWuA3nSYTGWw/Ip+6tA5Y7vioRr4N84waDZU732bnzJBpMn
Z/Nzve86Fi6wHHTKpkvn4439HI92CzFgbK1/DU0cz/bpzmK6HfOxNUPE/yE083M4Kwc1E5V+WfZl
80Ubfr3I7/pd316c3lu/vUbGq+a6in8CyaTC1YEZWUTw5tjtW5vjlQs0VpTsCH8ah0T/zJV+DtFW
0vHvAPXPhCF8uuzy81MkYjCQLF0X1LgZ5eM80hp14HXpR54zMjtBZ1L0mC5XLGN6o37qEGVrL8J/
wdfN4S3OhP/FnPl+AWpId9E2b0ilxZb78r+yFC3vqZWlv0GXSKNae69MnPyK1/k7GEkL1Ikx/1jU
U9jFp079BTb9OlyKJNKNhx4X7nuohamwZgESAb4g4MrMuroLink/SA+YjBfcmO/dca+GbpCQBYDi
tJbyiBZyQfrEUi6srF42Irj0dhiZSszcz4D7ABD/QrpQWeDWfaHpY5N1GIhLqB5lbhkJiSZ0AwhC
LUlDqU5LXVL7cGFDATApxH+tgjeu8eoCr3lMZg0KFSGczypAlZTh+L+gLEE4Cc7qSl/8Bmg0nTa1
l314BdY3Oh6Lr3nBPU8DJL4/Q8WXjmF/YUAknih/jXmxe2/Ii8or1UOHyeFLBwjrY84FxAgIQips
iRfFauFsm7T0OstQIOTp0nrhjXX3gC6Z368EaI4+BzdsKXeEV592IzwMTLGIqPtCRyz7R3O3Z9qi
c1TKaISpFIgnOW3UpRx60rFSLFP9Uv2TAqNWUeRVubkiiKrzgl7NzBy5qGc2uWFYzjnmenXikiPV
0+RSwc3GACvossPAt8I35BuoXFmY6LNyTZt9Ucxopn9ZSvqgb10D7FQRfgXWhYhrk4/6h6QcOSgZ
qWg8HWYlZkDIPYFEZuoGHk+aF2lDnauNlOf5JHydUhux1v81prr39Of9rvBsntHxPKA9bZRTuhW8
lJ+5KLWuR8kuK2y6z6YN1xEYDS/gZkrJl4hh14AayjkUKMUNqok8PIuScs55w7dR8D2S3BfFZKJH
Pqrdlw/zkCjkPGXELe6HXsnPyBUq5J7MxA0H45mkR04vKwsxv4chI4/kj3JGNUVbWoTWTP6UpmS2
nxq1vIZmKlsgFEmRPKx5xpmVnjtbKdsLs+MTG5qoTuMp2+plD8zH46BphDToh1OjsEOCis+gsoOZ
ZXzNP0uQ38tZxmmBeoRp5xYfdCk2Ysy54X3GliadoY+iOByUmTeOlQFf+wjii+fn4QmRojDWls5l
tNNRhAFda8E9tETL++fh+n13LkNyt6OqG2vCM8/5TqI0QjlwF7JvjWoiuschRRD+XIdPSIUCEuM9
sFIDk61vOJYOf8I+SDOiXdBXRNfpcOBd4foUfO7KB36Bskjh2/38TEBdOs2sIDqEJuMoDPqb0mhc
aTjh4HzMbZmL9dVpq8WfjoIsQjLrxMKiaTJ8LKpePT9DBukFzZUSYvkf4AI2A2HyjY8AR206gSh3
N5zPdwVKRUxTgCFHRlVOSSD+MT/bD4dUdC+HDfyEbuQKS61SAZx+SXBzVmQX2pFf+bwz2uc/ynq6
XHh67GTrkZUFfH71vfGSNBqSJ3RIwQfMDdFKqfuMMMYR60jfTC1ALVgYdIzRTOy3gzYzktes4lY3
yVc0RgBb8wXnbHDjV76fE9UIlM2cjP+G9eTF1sE5Zn6i5zac859IKEiMZNl5YgKxHWjVRQRtEmNI
YspFkaqG8oAM2vNRwr/l9z/UxaPYySCQFBAjhyGa5zeK0AJJVrRiX5p1GpezmIzzUKQA6a8BBLmr
cPBGiiOvh95EruV/lpLnjjd/phIDh09zsyo6o6AOCmutgGDmYEg9js3L1yJxHdF9kj334isdbIgH
oTieMxGahKNuo70qlzIQzS4Jr2fPtgrerME3kutMmhtxVB+ZjZuFzr7l+AdYyFZxpRIRs+Hh+YDS
FZ558ng63M0pOuM1+lj5llUFsAwiC4uBw2FgoijYjyZuP86NNHFVNJ7Qz9/l+O9vrf4CtAScuw0h
ZsFse13SPbTqXUxC2s73d7HpgcEQtRXb8aRD2rnNWkfg3XM/BzHLjMjWMd1bQzQIpfGs6Uh6cUOU
8FqZWroaMA2BU8IYq7V/nG1ANJyJIEmDyVezOt5ZLNkEyEt4G/AMVyKSX//sLUR2PbRZZ78Cx5z2
fUBeIxUHxWzTt1yqSYRXlP17NWjJjvb3sifvh7jYP+WEaULlia40p1fWgggWKGsoD9JZgH88iGHD
CQPOXa972gizqD8SPD+Yn3Pcnq7oDttejY7/2C+ki+5os84+EgrfJhufb77+5sjWouu9+5JjXaJh
wdug3CasqoB1bAAbKvpyeoVjX8n82DUPH+u09+u6/5HjIcjXlXvjJweXuSvjB4jo3DD5ST7z6u+u
2OJUqt7wYN3NXx4lB59K+IVOWqbdxFlDrpwW3Ch2Y9oc5bj/krZZR4Qc1YZ30ymGaA9riTKc//bx
lgEYdgLccFya0GWrVKt+oX23KITvVePAxM0t1jgbext5VKoPojEv5nsta1ZBIJehIq6aTD2j4Buo
T+gVSHmaTewmhYjIeGHPdU0AtfGThXziEqW3+owbhS+YtlRJpsBun1eFIkzqzcwfcEGstmENCIjv
9excWe8qPxBpYVYSOPrPsHRDNhwTTgNSWlQ+sukJ6/updWS7g54E2VrMcWa5AJFM5z/1xqVWjAkS
RP6ywWKQMf1XloVzaClrpWlJEtXW9g/nWFYCEksUYX9ho2LEZ4SOOZ2duSBOaxlgm1YHCZzKDdXR
Bu1sGrA8F/xKue19kXorKBDEl6j0RV90dpH0T8FUEEXtTJkAfxA0OLX7UzWozXphJ/X6LwP4UT89
D5c9UYKdybNDKzUseBeNbF9mqwGYFtMbxG4kqCr00f++Ig+tqnbn434B99MXSofhhHzqNzs+fIEJ
sdoXK1eWPVwV5QZbGSqZ382xT7buWlGof/8QGIF6p5rIEnUMJZXDPlpbLmwlTfL0j49sAdZ6wTTF
wsHsp4a5wQ0iPjPz8kc9Ga2kIR9Jl8qCpW9sBP6ZbDPeuaAs6So0lpww7xfSNAW0ethwXP0USnSl
/Z+VHsiCmwoAs/WVU/autdxtmDA92GYuMIOxPsccoO8BwDYPT+2GdBOCZiJx1Cs70sEqHAGvC66n
jfocPpOU/ts73RAUgIMxMvzto6yrngJJ423QFX4lNK06IJZs/h5NxNOqN8Emv7EsLjAfMoI6kxj7
/pf6p/6lvZgst5ZytWpG2+lfKzq5DCFjDuBFsMxPpDVjXq9XXnCe/7Ypl4wUG1q2+Llkg/iOpRtx
R2RpXeAjs2QqgHJ0S/KoZjx5+rX8N6ob94u3QHCyrJ0pDK8n5ytRySqa6uGncl3detcUChWoPFVz
XuhUVKSFnvVL9y/n1IIaKdEY0D+OpZmCkTAt4jjj0XNjpiwECKgBRWHEp8paWIyTi0ZsSDF1/uQk
U+KL+yfDVHPMdpg6WKxnoVBMpBMqJu+ZhgPne/tN/rOiAK1WYh0p9cEqOk5gcKdJuEaGiy1UNNnI
72DYhyvYBVl5//coDjjZu4evSEdclz4qUaZVygVAsmVn5NgUoMxhEJq0uSny5Spou1N4nSVZLNyS
UAbm2Se3l+3jf4MqHblagkPB/BFN6BeykkFUyQ7S7VTJpMXIUekY2ygfQgQa0I00SaYR0TSRNQDM
sCRyWjDf7nXDRNQtTlayEeEoWaJRHnc6+YqzGvR72d6BmAH9fqxcdhnW78sKQNpYbjfpRQQE6GVW
waVAJa8br8uTBOcOc1gG8DNSsOBlN3uqmC92ytHlxv2B/e2PwCojzau4LbiYhx/N7BIpGpdxtw1p
76TJRWhVeuvrfbJQZ4R7fSQKaV7OVEv48AJ/8uuEgzSudB7cRWmut60FaEuhfzBiUXmHKZkpXwtD
gPbzBBBQQgfwsIiqVA5vxjLttbeppSBLvhZigi72Xarluq3hGNLnkg9pvE9JOEo6pC2Ikp7CAp4Y
ZnBWv7DsEi8KIIOeT4RfEsgYkJOlfhbUMRz6g0+j5aR7oV8qpwd7fZuEZC3BQig/iwm/fGcVUoDI
KNxL7qP+5vS8b1hIexiDy4PalRaA2FcT0YSjUi5KNxJUjXSkvlgyjraQbtRvPBhdrFUqYn1h2FPB
OO88wPvGibjsxbJ0IMPmq5Tg4UKqv7Uqzf0E6kA5oJPoC/SiFb/WoKl4xIn6JcmqSEVYkponODo7
AHdxVeo5A1ihZSMMtTOqreC0k0ZnC2GakpFqH+dIgVIAu4AVci6GFXxKmMahM9H9ktN4FJXOZqRQ
xK01ZufV/YKgFGUZG1LRUvxF9wQC5r8Hy8fZwoKDskLX060SnmwOevjj/oZilk2PhRWrzzhfgnXN
NpcaQcVmpXvzHtbxj44n+ZeUJiD/bhKWVXqbzQfPAjLzn4EsZRQj+LlqgJAjHQEDJ2cCuYPxM8Jf
QjBlUfflQfcfkOERSNB1mMSqP7mr+KfqusBfkCT24te4UHJ6jtgC+M7qxj+1zVuU45QdeDIGDagj
lRsCmsO89MuaB8sIJG/eV+8+ZMjT3qszdANeZ0Czgk+USe/jgJ5Ma6L3k4loddOuRgjFVH+Lmyka
7pk8yQCIn+F/HmTy0RTts8veUdyC9zGyv+YA9Y2/QcTLAmgecXjiFbHwCIZ7FWbZNt4ZornZ8M62
MEd1OhjVwOxOEx6Bp5tESfV5svUuHsB4gPXXYxF30M7P4Dh5d63cUDT2m/YgYqGDaXDxIb6Jiqfq
kfYOVm9gs+pdMBI3d0jA2sp9KrfoaLMVqB2YXrBU0nvS9tco/8wsayXnz2APZKNFZ0XukrHYJ/zY
/H8pDejJJ9lserpa+E//MXCRmRos0WZCN2+CmhLmGUo7VTtRyKcBKS7f195VLIcoYMOCTugVHNdC
ph1Zsj4XZ0UhLtIE0ewIQekuCEyz0fCE8J49Yw3yr51+CXXsEVWExC1XSZpiTrxjqOoGuWZhamoh
Z/oio4Vh77e82+zthSsnR+GBruRhDFoxJdl1hbOYSvUZuLI7KT3J67W4l0iNKFabvgAnbJepK6UV
sU+KytFwiovz7yGRsRFxkQba93/2W5glfLU8HHA188s8Z+Y2+jtH6XO/E2N0TCdMRcHeIO+pU34D
q2Usz/vAEVNgYnLg22Bv7k38o5DI297LYdZvhMVeYfQjllL+lhWmuFCerAOC95ZUjrevAyNdgksA
+WSTMIPZnirPoiMU8inxhhW6GHLghF9xkfQboqCnKAXbavC05ZebvfpNJfiu2CnBevx8eVnCARye
N1U+YWSVfMTZ4/9hkCS+a3F+XVkUqNYQESVEpooIsMD2zRU6eHSZ8A0/gsbiJ0bU3CkJVIerJl62
2ubwUrfLpXW66Jjegc8Ely3Jyf+arQRV6oM/P1BFssFZ7ciJj3cmwM6KkjEbuBOumu+YSGO8eEEx
qpIdtqNBI5MPTV42RxsApa04ZJNMDHrQFjxripOZd7QXJJ03ijQaa9/zCIiVmBTZti4KdwkNpv+P
RcE2RQDxMX+4ZBWucyIucgIDszTkiuR00RIwf/VU6Z2vD34KFxiZDeJSt2u38FW7dMylrq2KDVQ0
V1LS2UAdAq6oxyyeW2hNiNmVfCHJgBAuG3UhY1ofvlpAttQbKYcHmwBd9qWs+9avxB/DN8rfyxbV
jiEAr+NRcfSXmmE5tJBaxuLoIQ7Y4z/BlSNcQlCM5C/AdNplCC+v4Ve/wL+06dOf3bJ143z0j+Aw
Rvn7ZnY5XYQUj1oSM6mEVQflRtpbSjx6BEIUg05c1DJ+eTmuMaqKBJy1+YSvTZb2Yrf2lHrD50hz
Y7BPlPLfbmkF7NcssyFPXCtkov5JhNK8cBq21/4CuAo0H+cavljEiODKL3bsQcXcZI2agM1Y4KIL
twC9NOSpovRKp2uM4omXaY52QHbETmWrjMzZfICsrPq10QUeNHcifn+mbVlWVRvrla5wJe6FuRAf
/YacqB4IAv4sHUHCEzyBWODy1r6oLrYgykpoz/U61U77IwUVXtpeoJCi186n1WZNZwGnZUfd99yT
vZs/sQXQL081i6Hyfbk7C7pbBTwVsLryYn73JtupqwPGbd+YHviup8cHbWant5hWQqJuihICNUMD
wuA5q4zmjH7Qmpj4MyN/D/VXXpwMG1DDj63daP6fG2POAn8gtGsC48FHtakGByxlGMC+njmxGCPH
IEePznjY3E/NTAs6Rfkcl4UHPXeZE++E7GVypxm46gPZRy4x+XNMqNjGVWt84SUQjURSopibgl5P
H7syBvotUiYu0KFTvm+IchqqQUX411sOTQTD3SfpFdQgeD7sop6pvMWZtyQxPrIuTZDmsG33d8bF
umNjAMq/uzHaFwaE2o3aHRpWw78q4qeQCoraazMYMmUSSTl45xHKzt1LtXMmlQwiBWuUmd2SMsrB
JBPV4gTauMvtNqai8SkL3YWYdbCDdaH+Gvt0ZEJJmZ1mFkrlYdLaslq5YWP6XWXsT+gnOw/B/cTQ
EJiAKsrjBD7yKJv7lbl5jLBxaSTZkE3ZUYo1WmPfsOwC93vnu0LPqtjJ5ZEutP7WGhf6Cyokqgng
amG7X6oYZPbl++IlqY2ktBLhNmOxjgMi3TzJLHDdeUvLC6KKtSRmxAb/f9AeR3XKMMx4uBWiSL4N
I5ITNndTfxLqUriHFY0GAfnsJPdoj5AjUKnz5J64fw8v9T08wQBqwX3DCpLCxgtlgPwU4wmjTdyg
QXkrwlcm2fzrwRHdQtM6BIHUChLc/+3Rvo+3LVQSNlrk8Jpg8Oup3GuTN7cQ0a9jrka+LtpOZHct
kSylv4HL4/OLBoJg3J7OWl0m1X+z3Y6wd9SGKUIFHW0KgqZfZYS8kMhDoKTDk3/YLfB1V8s9G+LH
nsWYPQ2FZc1a1vQ9WZuGu8SffYCSqT4gSvLJrQVZvGRmV1Q02tmNhE9oBy0qS6Yg7SRf3TP4p3D6
OyjOrfxY7h92tKSUmr7VaRjL5w9ZYsk2lwuCpLWf1YCOQttVhzZS8jk55iyvkpVHqfvkJ3zJwNdh
R1j9upMtKLcwLjJa1MZ/aRCJRwSP3I53ukoGFqlGd0S01Yx5cFSjODnPotR5VNJzwLqWNSH/jEAU
81kmeIdjijV+ta6cFBakUgKHAaHmwm/M67xb0NT/PUhWZZ6jJruM2h9AnUCT8ptuqScwkROZJC6H
PGxeGR3KEm43VEbXpqgzFxuKLJiv5EDdSAVFBTxDa38R1qCKv89w21soUAIe68YhnW8KZj4LDTbq
qo3mPeRdyVSYaNzegnDKUq47VFfZ0WrjlZswCUx9Q178rLWEOw4TnhQg8h4OONCC79AYnWXjATW9
1pKI4HeTXOujxDI4YZNbnM8OWAE6SIRCGBtSeUyVknjDX59OWK9PYkyPnD12HmowB7XSp4PjQU2c
1lfS5gEXR0cEuhxZHjnwXOcaG2y2upSqIm1IVK9hgSiCQKvoK1fcuYhY6wGkuRETDmwKdB32qLZS
3sqmD8J3KAL8SHlMt4c9BpFUtFOdfjAP5YEbG7W61XwG3zZ9p8+gk5ZaJgl8urKcN7+Qn3dwP9Rk
ep52Ln7XNaLFN1jJreyNeY1RcCAhku6JzvPcAPid3WM2Te9XbDR1nrxERoznt6PNh40rqPdp0VUd
fn3E3kEdKtbL5k+0gOrvAJYWlzwVSPvTlJPLJeSVmfxPv0R7HtLDFc8g+nF4qw5MW48xDYpWNjWG
4ujC8aD8R2FZDPEusdt9maIWY8IGWRJQ97pa9rH8PBB0uWUKguAJN60lPwZv9vLekwaB1hVnj15X
NHmaO706H0PfRyFVqq9LJAUMB0YFYLUspzN0VZM5QtQ/c1tNooVHS2Sh6jZJHv1/xYxtwoBkx962
c164BIh8tsjJGVMOaVOwnRfj+B8c1MsK6VaZxXH7c5VtHX0d82njFo7/GtsDS35glwkYiKk7Mxl0
S65kt9a0kvYjqWzIMWTxRkmItEtc4f2Osy6LcCiGx46o6qgbaCyBYoYY6h40LJYbofbpt9lICifV
zFRx3Nj+QX0hroCI5buCvTGKjbdwgbiyxcYqtwxoLPoNE1pKfXcQL5WlMTTfiJ9i+osCLlNJDqv9
vLf6AgSpKDCwltrZU/3caZEmWCkxS/U+5qMudTfUQfaVtvLvt+DTXYJPIjiNb6b3TJykkj+fPymN
m+WKsehvfx8ZXYT9eywyY83PX5dD1V7Yt3Y/0+ZMW66eEm0szRno0udsWYJi2ImwbfUR82CAmZC2
H9Eh20hzWfVTKBrO9lzowjsAQgsutEOre4M5/JCcBhqcvToryrvL4Yh0FHN3CvZB6L2u6ztcNTfu
4G+GgzCIZjAaGfI7Se2XMU2wtWC+BObLim/r413jZhm60Fnp8Qhtdx/KP/IdhYELCTYKlkDm+ToQ
247TQIY7EoymyDsqXgt+3tY91VvOh2GxS2WMcRQ8daktVkqCunwZrM2NiBPko4iGU8niI8XkoR3t
2wq2kt5pINCOMKzhwQiyPavJAl+yzHTaoCuKmAWLz7A3IOYyOoDSSSx33ZMMRAablYzHsgo0Jl1N
tFIQ+M0lmQQ8HNSnBxhWbLYA3h3TXoCh+yVSTUfQAsl35KihyuekQrB9NbNCc5uUnWS4SAR8tF0J
nCbxW7SmrCRHcRdubyP5Z+AcgU7Dp9rljVb+aGYPG522U0LzKfK+x/dR0+xCagINAsj+OgOiM85s
aIp4jXkF5C2ibjnIdbiignHSru+2CvNev1X3QBtWe7YbCaKfAl3FMmK/QOgFu41JdKnbodNy1fs0
bTZK1+CrtHRihkHCo2HbWo+IrFnuHLWun1gJBraJENUol8ItfQdRFmQ8ijY06LEahIqS0ZRMORNu
hKHsiPU5Jthmbx35Kd/YZyArqFOYLZ7SSGl8kZM5PzFmmqCxlzFpzcrIvvBS+O90Ed3sGqx/O8Lv
qRgIZJzPytq/oZ7FfrrW3yxpOUllLQRRvWbMFUSOu5jM9KCJyVlnrKtAW5qYh+Y/gEPlSBQApj68
nBAIN1Z8zP/4E1W4TLmAK4P8aKqLERJr7jimctKxdtMLGWY41wcHEdVv8E2+TvAyd2UT5qTVml9n
eOnGRr+4O/w1/n3C6VFMosRJP8i1PL3qsmy86Mp3fzM8XxqaaqDDDt4h03BXysG++BXk04UebURo
s8S8ZrWDhtT0O8tCtD2Yid0CYqbi6VBycKr27B6e1j4cRHWHXKIN4P8ZWPG4disoIYIk4TTE4+hN
EvLj/tLxKXQ2XJjuEm5S6cBbGvtg3gu0wEJ+O9dGsCzU/P9cehs19PeFnD/Q3vI3a2gKa4J7GKAI
eWK0N95Pl3WxfVYx5mgn6ah0b1PVOr301QOkGvD+XRiogLrNUJRoG0qei0gbj3/RS+R291/TRFHD
VsDcw7ubj7vAPNswf69Hjv7ZBOTiCYgI3VpzYvq5j3JZVfPvMPVy8S5l6MBHvOTL0StQTyJCUUQZ
AdvAvNBwNUxhIW0YG2M/3G50LMP7LX69YmmVUwxwms+gFP+COrdpe2WiAGuRrIjAaLZG9jl89iDR
Cdgh7/BTww6fJueD7R2TC4FI/FMO685TyjPHd8zkWNtI+pj5oyqLxpDqbmPKX9YldZ4ewVyPz22x
N0cbg+cOWHefM/R6rR8CtEmx5SAB7htiUViTIXB1/yVE7ak0tkdZM2aPS6IvlmizSb9NN6799QS9
fd6U9gs5GrZjdmFu6mIaRGRPXBbQrBW7argyRilMZmIyESPtOObPabjnBH2RJZshZhlItBuZ17zw
BgTUL9RIp6L2PtHVJgT5/gFNQ9CJJfPwQlt0xKJN/tL2KbToGPxMnqDY3eoymBORkQhSPP4EJ5U+
1+i+HT5kfVUH65D4XG1ToFMorGfhhzOgLHwDnTWtyRyCR/gBEe2KcBy+cqrv7vy7LYbt68Vyn4rx
HGhcTk9cOELGdKBtZGGsGhaBFgZ0FIx6ERknzQVpiVPujaruD5mq6Az8R6ZyEKzX4c+s+JeEH0AA
6MkOd366uQVtBNECI8YO/NGeZQPVMhTzZdDTDc0zotrts1BDgjxeNC1Hz8JLCq+MHNvzrJkrfpyU
VgqgIXotJ/Kfde8C7lxEv5/M3B4BvnfyZ+OIc8n4fYdISk52oN7yz/jGMHc8jr1JUhYn9SD6TAPw
xRCSsyF3L6okoAAw/tyiw8JY5+1kM1ilEYI2zto7ZyqeOusdx5bJG/QgKbdpjQS/kJ2tQwmxWOFW
OPEyqQC/CJZL1Ke8Sr01Oe2XIH9m6jvm9U5/3auUUA3aN9HrXChm7k1xnHyl7tfUfCwSA3EViBF3
1v3HFlJji7zOedr5iKuXe3PZmOK7t99ixJuhsVs99oaeAkDtg8elxYJbMgZRbJWwsmhgnnS2Xu0o
bAdQAI06eIhWx5XuaI8pT21H1mH1k6iEReOug1lKoPg3sWb3Q2jGDubDSZl+cXPJ1JQUW6gHSWhL
/acNMo8XKsM17HIzcTbQdgFar+tbE6eeYLX3oFFAYo6KXGlJj1ibPBEKnodnOb8ko+79cOY0i5Do
N3Sav7NnBoP3njdP2yysXockWqiotTZIhARRGOAvEksHSvS5TwLj2oY8F+9HiLuAPrcfml7J/fAe
hNh4ajNPTlqZ8m508B/md+3yK4vOroMMhBCwlYYWhfF8hPvI6dXzAOhhjtwOi2Br2tH7unImqV/H
GdSjOE0R+Feixu7vum6wBADKDXP6NBqZmmHJ7Zz525z05FA2pW8eHef9V7ekTKlmO44QKYA69BXj
X/an/KwfZjGq7M3VsA0QFAPA/PUL91noqPY2gnEe+WSA1Mpa46nQywY/LnvXoCad6CXZL2fv5TR2
skBfyAeCgST+C60LAQ27FUcYAGNQVdd2I8kL4FERrIRuvG5hrEd5B1lSJTHb3QQcqRpfyvgDojZ+
jm3BupRCtry5A0XPcmzFBcGTvko0NQrVLBUJAU9HZWnl/vhcqH/l7JwXEr+vQga2HW3IpssaIxeQ
ln26kup8z41NqgH042RoGlavm5FE7kI3QaPqdc2gq/18bpVEUU90TO0onTIxwwoB0NE2srlpjLEZ
/597tCvnhQ0P9PnDzzWBS+T5UJWqEs9C8f49E3huOtzlu5xaeV/HzFpx8Uchv9XtAJr5l02Vxrsn
E/AgTTyIeUk/ylLftZuP6U68Ysx0yHhTPmACxADwtDkofAieX83dalSQDXzL48XY1R/ATA4FYysC
HTCgeMxoDEHyLEMr9RGkkWn84Tph8tOmbsLT/b10kfusObzQnrbY2fCMDI6kU9DtE8I4EY1DZXe0
qFq4+5A6rTHrwGR4+FCfHHZcV9JATfU2UQR/lErI3gdCnCNZowE4zQyeuuY7wHnjTWLSshu8KsqC
DeAXJxIQs7wlSxg3p9GWSnVPIUjwcMOT9k+gVQJ2Cf6PSljU3UZ5uUjDO/mXWtEUZOn2lVv0TUgF
3SMEZUGbLKwNXd+CB+KZ7k5KaYpB85TDHn1YrvonV8aW+X+3sDfKdq72R9JpaFG+USTlv1+U37er
USOdy4z4iofVBg8lzHbL41tNEytaAX0ozkBW+TJKyJ/iwafFCI1UR5sbK4TikUTlyry9A8xdcsH2
DRAKgux8C6XgRiJS7vkdpUmlqMF+QkgmJ3uCKiA1n9w/+Wzw5vNqq4rOYvJaDohUCu+IJvMfOONx
1VK3VLm4h2uZh4mIcdFqpgFSwE8B+k/sEkgBgwK0scDdGw4VGXw/7KLYq9XTm/M/NL2LchnYQVum
gxI1sbZSw8ZIxWcb7PPeZPf8ues4JwVUZUsVaLB8kIVVzUv9U89/DJLMnswCozKYjRz3nmeiQGto
D3JuO/puxlN4FldpYh9l3oW+r7eP4lWt/6yxlCKoat29Xc1GMPEf6AH91wC6hbiAS7Z/Fs3ZLuit
FLcGPaRyl9g+AFVNsWr4RO7qUDEQeVyn/bbHLchAtpRtaRbFw+boLNxuvtbLd41pPhcXF+n9Cz2s
DxCxRCoOjRRecUHAB1hfxpAHk5N6jGm28wbk4gBGTXXuEccm/3AsBnq+IO3r2Z52DPKqqY9zHFmH
sZS1H57kgWXc2W7ZTeachwsJUzYkn7AEN3pieNBIHCaKm7Kx5kAk7kurJNhcNE3hRVa6Vbq51STm
pNbK8UjjwEGauQbXqexcyaBj1E5yiv+WUszs5D3U6Db2uaeAUEZ098qvLY4MboONaWTRh44+r4Sb
YjgvlQOsRqzCHv2q+4228JNEtQfwKgCleVac0jL0cVlr6x2Lb5DyyemKCFb830u1c0K1PrZMzfpT
ep4ODlfM0zeisyujqrvQoHmu8zoncf5wcNWHGbAPKe8p7mxyOA64r36pv4ODZgDK3LQIm1c47rb1
sfB8Atb8iniEHrek1GgJQcdYywJacOTemALYwE6Jy4QrtIqfAQJGKYvein10pgBWsESEO5XyrKN4
C67Fv/sIGxaO2GWp/IVSgOJa2Mg3hTdi4dbMgOJp6Ktn56nKfKAPWpvidv0T/FYsA9B61fOQGGKe
0uoqMFVXCS2ElSrj7Yfdr1dpG44YkAZpQlGZj9d7QkG8GYn8ILx3iiBtlDuNbXmEFCscaUxaVsAK
uKGqj8bqF3hDgqouk1N/+C5nZv9aQ33ZJJKF8yZfgNVab+mSJUM9qr55gSdbW49lXGT2ESjJe5D3
wUzKUI5GGinSb6n6TfMG+XWJEeq4s3f9pnDKRb2s/G6jKMZ9EueM2DKBDtqjFzogB+LU1k2SIFPo
tfXW8Ryr62lKrxwP51LYb6H7ES1zYEHHEtSCp957Pk3EwOlXFl9GYUNkTmpWD4Z8v4/z5GDAmpQc
SRJ/z/RYokIA2vR03BBvb9QFphb78b7a0VtNtGQnfraG1j6Epj+6ZxrcEQ0SU5L5m4rrbpVAdEy0
nF0t3KSsnmNVy6Xep7Rj3jCFwOnwR9j9aWFaH6S8cxGpIMqf/8LWvw+X+GTaT/NctnUJBLyNmZb8
Jq9mxUG2gCDkTBCzmf6Fmutp0Bm0HI2Y8VffYzo6yWVARQWLp5g0oTrVcmkQpoJ9DHjEnNHn4Aem
WnzJXTSfIAlyE8MAKtCGnse0kLzsDEapvGQA6Tcv4xMvzSdXnlR4eRRyA6c2BC04ahbUhvbJPjW9
vuBTxRYs7aqiGLqE/7LSRVSfdlAQpDhZlXnq0te2GtDs6z4duzT1R221cskTXTs5V0QfZmk+Vxza
CqNta/awdw/PN3mhi9kqfqtDv9SNGjS5enx5BrHKE9AJp6oA8xzgfMowQSt+v+yObfTZV7Ocno6J
zF+A+8oxe1e07Q6+y4/a2RjAptOMXf408bPv6YmMdxBWLSOfJlw+3ZvECT9uaOvyWltzTLBkjl/F
v6lhDgUzNPVhLPH+ofwZgRio7iOkW46ushu9xJvPKK195pQaOxn2yOe6or9i7eoT+xUxehWBql4M
qv5z2Zu2tiVinCsGwtQ5ZAUyFzTWzjHd0IOq5KocA67PvHfy7pdK99LiU5oBCWR9yQoawIKCUk3a
uBmpLwRoywQtVrMVbQWp7rdngzUI1ot2fsScrQylKdWPn9nNkD6vZrgnlql84BqbZ/Hb3mVz+iyc
TUT+Y9vKdn+BHtvPAWP6QTCfp9rpFf1HdL2hvTfee3ied6NXHuEfR1f3teYgIW+ngtEBTIlrf9wS
ZIjzkxCDbXGSfHr1ypWelxuB166JrCCr3yBnz4bHE8H88x4URTUc8Xm2Y9qDqMD0dQRrlw9N3tyF
ZKQPTAIMcTVnsI1580/bFtswS4EZGqmy0yf1QJQS4QHhlf27vL0LLEPElRM+x4H2pMEY/O2c6Tqt
EaNprxMx0xQYOJibJqrsl2458Bf7KZcQDt0dUDbohU8usq38Sy0eyT0H2j+Dj4An5NyAxUFQIf9F
b+jZO66HnDZ0iQQjr51oMwYBbyIChy1Dz10l/g93gZlEnsIWe1+pOisiT4NHAri4xWUwSMtzb5US
5tdIuOhiyt4J4ljGwCmjhxsKeNhIqgthSgDqUfT0eLwpV+R/DxkdsPnuTa/5ZpULsOWaPKIVIqDR
xRHY9yicyf8/yAzYkLKaW7j/nFKPiB0dCk/y9IljYIJLHeWdg+z4h6VQC4JX8I0s6uzLa7unDT91
4tUdkXa1yYvfC8iaA3wr3LgEYHPfzI4hu7rwuG/+HBiipd550iCTYD5ZbscRBRIvs77zyMHao135
VGD8788WDHvLMarWSwhxmJEcKDtU0sKK/olqwhWGdiTNOufTB1AIDRlZjhzpx9Va7GtyNywbWf/B
pyasnN+wdogX3Abfuhs8rBRtBMYHjkGv5WomTWxfmMAtFrtulyoqYSePS5zP4Jx0caoFj40SwBMZ
PiuVtOyERPT4O2RZP6mKvpciSO0MDBmNqwpFfQFipr8/8UbyRb/hUwdZ0YRYuqzV4sA371bTlKOV
t+J+ruAgFycfNZHZD7yUCUlffkxjzED64Z9iaynW6+lelrm1uSx8MGxK7IcXiausTMNme/TpGrU9
kv6JvzeU53mJUQnMf6yVBe+L62TW07RLH1rRL/ZxfiZ56tXJ01LX32KseKTJgMKIkmERsaP+5UyT
TzDk2ITSYxAg4O+eARiY5q3vM+uZ663JdasLnZWlC3cBkMiwyqnXu1xVzxqH7IQTwPlsGEfff9jO
yf4k/YbqIr2LLLimQT0XPSFdevc8A5oE9WNSU6dczFqlta6TG/Psp/m6wAM4yMRp+J5Efa/Rg70f
TLH+LQnD5eWxZeEK0kQDZPUa1mECAA7dzNnC2PAfXBqVfE+shsBVV80JZhCibqv/m4ugDHBVvhlf
+8K2ZeT0FIKwQeBcNgHra0TOud/D2H2yimLA6TYnKR0ZW0D1ybbuw3CCHvtO+wNcJXQw5vp7OpPI
QMCTFAnugx+w0/cCUC+HoNPgCAgEqGinT/9yYzW79e/aUOOpjmgyup65qZ+sQk9JQGEjYJKdZdr9
7PBDtzXmLR/ozC/1NC7/he2NkxFy+bZ9s/SFbn03SKtA8pGBfJKSYj5ghHLtxk5o4KWr2+FkhN4k
0DU8MocWtyVyYACzqMW2Njhy7raPzd4DL3TTDp9UVFXbY41FJD30YNDg+uYxQ8hNY8dis3+YkLmR
HgGfFrbK/Z8Q7Hn9yffB1m6ODalTflNolP4F2pXz4cEzweWVYSTBx+lzm2qBO27Ac+pk07sz7oRp
qafVDbATqQgDCsRX2O0A5RjFCwbB9ypWW7iqdLoNU+muf3dybWk3hahvQnO1x2nbkQIXAY9/KbjO
rKMEBoG/p5WFR6ZTjOX53azSvhJ9iZmFAoi9p6zGYGkjq9M8XZIP1mOScS3Pi46Bx1SP+JajB4J1
ob4QwKiXtHij17tesFFIZsDkNyk0vacIaS/y761jLJ1a717Jh6xtLsMlSPWy1B4jS5Hm6w+Il3LP
Q14hPWOycg5QbAaJErknW6TdD40pWhG4EFyJOmvM/qtewgrjiNfNm11zeb6PWJi9xYoNOmea5oh0
4L05pUI8mUWcEG8hWZMeot4nchK8tgNjrfrKh1ONhfhZIoEF8ux9Z1UHV/RuywDKbbcrocYsvVWq
8QhKLbuxM6NV2nFIjekinqOv6JgKKOAdadR2r9kJkdf8G//dl0SXokBC6XrGgFamxMtfwYVLdWb0
UjUTPwJOuJotfOgNTgi5QV662RIl9JFAWac3hFy6dzvrxdoa34AqmhDZTTa/zqVMqmM+47I21nqa
uTI55pd+FwhlzBUiAVuOIaTexwn9YRZe+iSysjfZOQxLuyK5u3KdTV/AoA1ABD90hxNizgacYr7/
idoj7Pv4QR+FPANNFJMNI3w/zAAw5glYfFYLDC0AdluEiOv3t95nyEFHYS/6fMxfoiiXkxPuh7Jt
VURx/xHXgf06R88dk7eZGqPmyJaKYGeluXT41kiyu7pAkAKdGK+Rbhgk4OCtW24p8oLWyck5fPrm
LObNj2vLNJhnpvzh6hycnKmcGiYrHt9iht1ilMNBtTpw6Su6GWTYzlghD695gKnJQiXdb0rhrLAm
kQ/m//tjLY62ctTQ6OBhXwg0l2rYaVWIoYOSClZVJ9DM5Cmyhtj6SSnWjCrpzB8pM5ocHXuIquoN
92lIWs0SHR0Zd6kfPpFPmjfov0C1gC9WRT5UbherNX6uaU+8CENXcneMYWj2BOXt/ok2JwhrDnB6
RPEeZmo7ey+v0PCkK8XJBg1rH7br+AqMQmZdTZCzr1u4W8COzS/w2LlokfEtUoigVhHDa79ruabC
3LWx7Y4DN5tZOvPFI1KAE3bcLyzXmS5kZS4MNwE3mseGqyOhfmPx9gJVRGgi4s5mJQApUqPQ+kJs
SHqyyt6qYPyDbF4wEscTT6ftBq4Ajq+XiRfYA5gJ9yDRbt+Ct81YCwjnBnyXS0a42KqZ5PLTq3qU
xYWdjMiodDQj0u2ynZ4j/Wryosy5+d20yelGfNYZaqoGB/GWYE86AX0KVM+YE4ZTyLTTIZXBOUQi
JNRz/RURo4mRo8GpEc/5yacM/REA2TXKEa4CoSSWVaQY9JnNTmFnR7U1LI6vOX83nBXbGCmmoRmz
dUWwV4X6aBu3EDxNpOBbWPmeGdif8dwWseKKGmPMhEU6pOuPDsfUlY1P47gNyiJbqOY3d9K84ZwG
+dwCG6o6JRmpm27PomxKY0Gy5pHJ4+DgexhhCvBUiSJVbXKJ+Ez5YSYw2K8FiNP1pyLYNCVq33+6
H993ZqosPVzR0qWxh79+isCuMMYEK8RMm0NkK4sNOgGWpXZPlhW4ko1bBG/Bg/2kpZkMs7jbld2K
EQz3qQnmonpd1FW/NsrSF55F791bBXKvowAA81H0bHbnEsELrRank88OrdaeXa10h0S9QsS4lUzh
Nz6D0hORnLtm/m1/pzRZ5BrMxmwofxh1YiHk5kaWzPXdyjYd/qGCx+sME/VCYhpV7qVlrj4uOKlX
n6WUoZ3zXgfWYS49WAy/w6/zSfa2Z0lDealcaooKb04lv4qFF0V1YIes25uWPNAZZxW2kdqbH5EC
bLBIM88jJlK6dxbYadKAzlt4RgEcXLFlZcj7rFtXvW0KbDlezJBVBw9vBoqnin/42l9vf0KY8gth
sXwY0oNvyZzIhdNKI7coBh9IEGHpQfezsiD3cbhRQcl4SlvGPoDK1QBZmiU/xWG+y5GreALnHJHl
yniRLpzJ2plbNfRUkEXqy6j67beI+WGtc0XLvM2+GJRbjo9MW1NQMTGC2uv5CuOskwzIpouN7g4e
XIvXbBH+c2BbJfTAbe4gedxjMuMnkAiLABys5AdOtJlyGV4rRaBrMAB8CovLJF3GM7kMH/7PdqFo
jeoxnb1Gd2yde95qEY4I+nfHg0UYSRGX8aEQ6Ex8woxsbA+vJ9iujlxR09leSsmaF2ItEqLi7ABf
KVHr6tnw3dIMoeC4vgukUIcQ6JOH6zrcuysl6BU1ENBICCCFd2x0IV0Rkl3AjsbS1hYjeqP24CI0
Zk0HdlVNZKPlB7QIxy0cXBjvRXD89Y6RkbQOuhYc2xBgQ97xK9zv7AXU/7Q4FL6RJdUh14FkeOif
ncKld3iqq4TVkdUBRtygigTmnoOzPME/tU4OBlsuJ7pLKG/U8RAr2BZgjzciNgSfbwjMhgNd9gsF
gL+zIIfu/mi072FxIDQD0gwPLfVNvD4Lo0UKvPPWbu1MqbRocWYdzxzOxszGl7PQH4icxIZU95wE
Xk0v2U996MLfEIi9iXcCz3e6mYWdMbqKTkIuEhaDoyrAqXdFd9/n34Se3KaF5vfRYwLCIhaHQI9N
5qxZ1w7UiGbg/OEjYm9fkxo2VHbdelDsCoORbtk9RGr6xtUfkg0QQMtca1MInoyZhI3xIfLrBa7D
nPgOTBwI5YP99Ae3mb5PEfHwxqjZfeloL5w6JbbEA0nvdMK3WRO+YxhQhxMyYK4fNiSS1hdYohy1
5e+YrADSWeoNZ6BJGWc/wHZPKNiJeNwZpj1qYeu/l12Qt96+UkydXSjUbJCgcfAoIXIP6awqkVFq
qyZfcOlKhnikoFRMNcP3oETbVsVkQEvrY/mUYxkTjN4LxKrac0YCEGIBkczKDomyyupngVf7lRTD
YYEuQmvkPciPql6xOvvMvtrbM8h/M/83n7fINgkXcedGs+5AS9KSRtmCFRx1fiOGUV6a5ayL9rfO
ZcvPwhb1tJz7Jgmk2oJZl4vAokSyGwTlH7GJIwGVpaWl5thuj+NCbc/BXovEWsxWFoWIgSd13C1m
przW6FQZm8KqKYgwk/H6BKLFVeZJjEgwPUHzonlLzl8U7gjUQWICz5okkqyNcoJke6Jsq0HDPlwa
YjUWojXte3pCg8d1pL3BliUCc6UmUj+bujkUFhz6x7l3JZFZmpMDbYdCxnig9SYccp6q4IAIS35r
nV7dSfAP4LAsjSHQEKg5NBqAxvgLeVUy50ocHfVvyIynnzS4kx2hTw60vwQP0FQB4SBh0wT5rANm
6luHmNVGsemDaWNkQvxZ6vbIoyiHwTpRyfrH6JlaFKGxlB2eVq/xAxJ69NhKyuUxTorGFw/zt4jm
OWovXyjUXOJNHlGDi9RB6Ql4ehClcSGAXtVW76hjul8GQhTU9b2/1ArnJ3zPbksU/sEXzEQdrbKT
1AtCZoJ5Qw1mLb6l3MUd6PXMtaJwd/WpzLTh0A4tXiCPbGUxS/fV4wmX/+L7q5ZD9Rp3+2l/mCS4
MnbCqmHb/Ie5OPKbThDXQhsrgbZunpssUABaYY7L09P6qoUjpDw2qra86s+nDAV3xOnK1r0frFRC
l3UesQYl06+P7ynijUlyuJV09WlAUlO5bqRC3943muxKtlgD7n2E3POxKDN7P8D9ii3RdEduQYQZ
F3dOMoub14V8exEgQw7WGAc2Nncy1YEPyhtJM50AB2Tr0R8z005h1hh4b11hv8jmg01hEnhD2K+E
4h7vCm/YXC7X8CmxuQGFgwR4798Oe9+3bApXUbOgD7k8eDcxXVagZBDuVl+WOlkUVtl++q0/hC1C
Gtu7zTY+cfGa3QdIljBEySK1MDahvbIyKi4FfO1AsJZK8aqBVlyZaB3IVL5A8h+LZX3AerEwLpPo
aHybO9B5+gaYVcmNjre2vOXDyNaOeks0dRwQxnEGNGlM9dBqwXCu1IJFuFoTuBa/Flny/sD2Nz1V
+PCTFZ1+aLTIba1EKauzd7s1VC9CbBwxAMGsqn2dWgJKwzU5eK7W2uavl7aAZ2aH3Lb6nnH+Jp56
wSuuaJDhgTgNmiPgiisYyKyoY3luEC9DdvThSd2DGR+Y1SuZLfEO4bFY1XGM84oLBmvr+lb3dsXG
r6zXvIddSFD2Bzi595DgTFyS8ylw46tn1mpJo0BwLU+KtBvlzM0h6PICKNnQLO6Blt8wauBiqDv/
shdqusLtOVQdE6+pmd9ZRTJeYJ/wL876JAu4DFRqNngQbSpP7DVBKdAoXZWAfvIWi85JZMyOKKDl
O2ZVC4V5C6dYX683gI1rIJ2O/+lLl2P2JTvwbwpbrkVWR0i9II5PMSRjXKXw9rHu7XU/+Lcuw9g3
5tehqwDjmJKtOYE7p4MIa7jmFN2qHyiGiipDxn/rM7jm73HNgLnB6OM/zzzIq/9lIomGFtUNmfcA
6arfQS8sXm0Ty55U0MddGuk0IE+rYBGM8qD3oOx6JkuFn1BrqSY3zG0RwNYjHo2d47Pk8OtJZ2/5
IafcB+FPbbp5ISKLNLMdGWn2+vrda6q35zoVlDBFA7qCMlRq/WbXnU8BNDzlwyqYseSTOk9Cu5+t
uSkzMwsaWXrlhYNKnebrIRCNzJH+AyYHlgC6rh4Pa2Co9/9vVN8ODLsxD205AnIEKdtaAOyqrxCG
AoVuhelff2Q1B1BuIkPrY9n8I+vhQIaJCOo6VMNeT6DpIiZxB3L0sgqBKpM/Mhr+kASIaB32R/4I
8v1i38aPefNLJ+Dt2KTIKoXiC6wdwgsCjefXcl/sLXSp5LiFV0ZUoOnWcQt6uxyhJqNp+XlSJj0m
U4S/ft8Iqs5WGS34ewajYCSbI5r3KlCkRTiu5i851v8As6nbRoBCsOaIfKCpOYSHx02ZO5YsinX/
/Cum32UzvgeWeX3H0fKcs87fWoM1SbmO8hfzterKnl5hL7dymA9QSY1N714ahsPunxt4Duk1OywW
Du7Hepa+vuzfbCctntVbAmNaFWpimNu3V1Ho0xQQflsrV8gXp9dJ6h1yg6xdUqIB9Bcpio+8K4kz
IrKLz8bLgf3IjJ29W/5HWNP1T1HWLlGxEBD+Dqv4C2psx0CjzrqUEvhWJ7Wcfpc0PgfBKWEDKEz9
nUYTt2wom0Jczbhtwy5ruZGvmrVPKwZH1f/mn2lMxiEPHmMlHQZ7ujTxowF3xyXiRzWdXBmDBR58
mGZiFkp/sYw6x0bLnkgUEnBHwIJ2HnvGo8WltrQsunj9PTwNSIKeIv9hd1vIzmpTDeoiWvMh7Hiw
WgiPWGQkhXJjJi5q1DBtzur/VAL4w3WUoPxEybGOTpls2Axqre7kyuBBz6NiTr1CeaRYXZNP4pvF
2S9j5gXpALPVGaVbVJ4TH6f3P8qZXEp4J0IwpXqngTTHPjDBBF4MQrkxxiPW9dgDVyi5Zfg7b0/6
Q2f8b0mAAgL4ylixU/GLWmh0wGPKvWaK1Kh+RZH4Lkuf82kO1+2dA6eI6Xj2gUr2HZhXZ948MYZ4
pAbZUbC0PfbmGesMzpMGZBog3+9aqk+XUl6Dopa1gq6w2ktySuxCVDg9eqn/TSOFt/fph4eNjA0w
NBl6BZVcnxquQpHL5gZ6OLONHJVQuItTXcWEP81mcXYkZEDTBFFXQdN3uHngXPYDUbcF26s23uWU
ugg8xBLsm0S2WgjvwtaGsQ7iP2yXYhsGkzI6obvnOWZbpMnH1Krk+ZD2jpoqA2rBhpe7kF9ncn9t
vnLHA+W3VVXRuIPJljc8CaKwXsruASd6MKj3OCq9SevuvrKDEHseMmdJboX7Eig5bGueQqlvh5AM
Am6+E+o2ABmWcqaObxSQudmKJAVFu1daKYKOasJWuUJBrw35PsFMfZTakVmXbXKfIVSy6c979GOD
gNYY0ePNmdah7dZWAL0EX5ubvjsG9z96XzNrlBsDdwbDO095KCSeB+k3+I1zyTwVpU19QrZtwqcf
IPIcfWZ+1X7EX02pG0gb2OHxHSBaaH8w/TRdG5e5nAjyBdt7wGh4dbU/CSLwf83iqxTnRl9pFYyv
uQA6ht2FJ56aDPRrU4/6WzxvHs/MqF5eXLBYH8Sh/e88SpS4OkvnDl/2DfKjTzfzQyJ1ZjpGax8F
s2mjxwQJAnc7zKCG4EoOXMpspyHwyHiv2K13/R8CkcFm+rrdypwXNUWAPGN8iNH/ogpKnGzU/aME
q2ojnfUsdj446NHNMiJFQ14l1lh2lNzeyCB6izNJCcGknfe5g7Wa4wkM4GkF7UG8iwdVLrQz5QNm
n0A2mGoD5KBxX7FiomaZliyw/FGjVfWVspjtn476yqkLttujMMGyvA8sVgLBQLleoI0k9s7pHMB7
gXAnTgAldRgzqa+vSamvNZ8kXDmQqSTxpxnRBWhNn3bH5kZKgaG1yNfxOqkGGvbl5oiMbecJHlGX
ASj8V9lrXhHoVReU+BTQWQ5l/BD/xCHo0ei0kUPrgB1Sbf4SL7NYEF/5CkFtGp5aT+lGi8JdOc8Q
Gxdqlef2P8em8SyoN5MupfHyTXBhc0vqu/K2pIPU+DS3OskJTBUizgn6uvNOI/fx2mvrTSuLfPV3
eQ+MKRL5zLaJ58N9VPS6z48JEPIQC3yAu042KAZsrw4+mUdq31bNu7gQqSvmYUbCzrOfRFpo6gNv
vt87E2uckPGnmxtjt3HAPT0Mf+TTFGV+NfQ9cU5XTR2o1wXW8RsyKi0s0FrttEEjGa/HYfTyf8Bp
Y1lQIputVrGfxjDprEqqOMhJQi2CRtFDOxB7Lqm90gErAcYbBF+g7buDXoZnEcFEdeUCXZJfBV5g
z6+vWQrUeUwieMCPhDlqmCxPyjXfnRAp9wTJqeSnao5avPJsSvnsdYZ7B9t2s29CjD7tpW3lCwUX
6srf6eFCcqNiWpC5jgeykZKKNvuRWzIUdEkENQMvbO+ohEoPv86W3wDvfFdJyEfP66dVxo+aDTcV
t4uOCiBegpNbqOCQn5yWK40lGO55daZV6fy1R0Gh5GlvXt1h8nvFt7uvH1piFh+wWj5WxkpA+rmK
+79v3dpCiiwskTogheGIq8B8js/bnD+ZO/WweUCu6wdu3lesM7un8S+yT8473towZseiX8Sj16cE
OGmFcXf+Tfcmj8/WycpK3pA6LyaSCX+V1RGjGan8AZvOFr4/dSwlQYjOx5DTPWs5wk0urrtN1XDh
Sb1GSJaQcZlXQgq/ij+8Mb/jGc8oKA98TMqS3SEwN9bgSgTwpjHGxA3cAGRngrtZxaVEDxHv1Wfg
zVZ4HhjYLhxWuujBmFmRzCHEg4MWtLX+HaOJO3iWD+6X4w545z4Yt9NJMwWlgz5NIFaXf37xn1CP
sTvhY6LRsFvycCTfVW4OfHFHQ+7yHjAN015tgJKkI7uzmxGpmjdyxB9jeIL6bCvu7sSh6FTlepr1
1f6yeZaJhgeUwoJllfUwej1e6nzT3aiAKvlWMt0kyag1o6n20kOTnPZ4ABNh7LF9BjuPULvK+jaV
Mpp5YNSBR3qUDgPG9IShBvAVa1IsQHCqor/2JqiCmBdQr9kwJr8vhwQNq+Ushp9t0ZwIpsdsWjeL
aALIUyjrpZJ+qOOyRyzaBZ6HOqwBKYXy9YnuFiKBdhcvdjf1b4iieB/JkNelPsbfRZ521KwmjMdE
ZL2YlzQHTtpfgZJBM2NNIm/3fCci3a6Qu9Z9Y7/fTgpSQk6jGzYQNMTkDFJUytYrJmlzv6B7uiXb
hlfu5gb93Hn+rpyLC39JJE5GmKjZ79CGJCoUWQeTc+CHB5cJwOUhHzMZ2ExjRk1UUHWEvNftBZD9
SSe2Km6b9roJz5FoYFxbbLp6HDDsyeHhw8fVWJw3+UdL6rYZ3ldAqHufSZ3hBRRj38MYzlkRKhpE
5IGeRJGsYSxAYvyPn7EWfdroRLuZGWu9zgzipuH9hRWq1CVf5nq8+QBt8Ptpc0WnwpruoD7fBzDr
UDvJqhs8IfMK2q6+TBqDKY2k6w0sKQJcNPdZVfNkeZJzV4lTEN3FPK3bin8roH/HdwxUbxnsjLNl
PhD01oZAcErz6muvIWQs4eVCAoKse0LoUIRLEnxn5uwcFYLa38N0PLPb7H7Yy+WPm/GZtp5h5Ken
EUuooKMpMYS1NvnncMQ5m4EHVKW8PTORVx6D5FpisRaEDgasxHWSP9WWp0kfTVNzuNJR8ZsTTYzV
5xJxahjOKJlIR6SZbQmDLHbERmJ3uLuykvSBrKRKR3+sQS6sE2q49dMNRRbisC0MLE9meaMaBt0Z
NBh++/0JxbhisU2k2lZmoR7mqNb44lRuj09U2+x4Oec9QGZw26V3aPf7A+c/mu+XvXNscDU1y7Q1
q7XphudOby9CrckGzq4IGucjmJqXtNB9kkycgj1OzSJc5s8baK15g1Q1IF0yM3UJQODHjA7Og3BA
KXHNlxXQO4A3vpj9BGa+chuyZaO4qt+choyHV+iGiSSZ+v6FhTuHrI+7JK9ofX/J1HQIdzZ73/l8
MXwba0mCHkOAipMcRp/acD4iZwJ9RWFiEWwxfQcYTGHAnJ4Noc/D1nIsHRrPUThwRxgbh6k8ntKW
GZTMa1+fzEcZ4GN+z//pTndXP4F5lTmJRrVx8/FD8ncvZRuVEmXBUrlghTMbzMsUBV3KA48EJjir
KdUvJtLx47TcG8q0KaZpTpXJKHMdueDAiJJBI9hDL76WkIOxXh+bHyRpTMo/e2NPZUdF4TXuBvQG
FssZtnmfr4ZI+UJ1C4Zn4PaSL3Q0hpqDaCtio1RPtAOv2eULXTIEZ1bKqqqCKfh7drRYkilbKzyM
CzM9B7GWfZ90bmajtER4Qx3rsjcoF1F5XVQJnJ0y9OrDAYZv2Tzw46uli/As7bfuaVvC7/sjjlJ/
TsegSqT4CfzzHWKbrhRfWj4I+QfIttPGMnuVjSWvTM8F7qJZbk9zOb3YefYLjZZe+ipHsIR6sa0x
8HjmjIVsHXBvfFGojU01FA2R0aSaboN0D+xsuFsG+9cVzeQF7AY5dJZsMaq4GurrpCDgQqxDFbjM
Xbe5J/JrhcZsvAIR+BkcYzSTsnrkiWqSovT+4PYrdvD1C4qeSbRbvQmJG/IQpAwkezCh+Mykeb4P
AmTTKPoWiWsHeW1AK+bBvr4pwNXEKWM5dSYit0i4Roj7v3q0/jS9QN3HWyq5Vqmtf3N+9vTmlBvg
gCgyf7GJuMyxRO2cc6fwZCN14YlTwjqls510Boa1l6kgGBHbe+UVzoNMxhjTuuboDrT/0YZLrEjg
qo2SIZX09nz3OE0dnB2PdIunOwo8ZaOGieTRMMuK9NTHtsPsS0gyzRPCtM9LNfG0CklNqMR3Ix3m
AzZMNvKBO5oMTIW3+NhSrnOx9xxSa4Vn0GURbjOf6Jm0iFSpWQlDipcoq3HF8BoIqjiIjPCcyIOg
Vc2ZusjQWx2+S2xICz+gPBvOYcnNsnlzBijX5kJRPPYG/HgmWhpIgHjVXcayhysx1UyTJyapdG2O
7EFddaSqfvhx9k7099PhPsXcPnj7yl7FRoSSeDpSGNPwgELWZe3E5DSFFwokcGpP4mtCYHQo5ulB
FKUbFQUdiSXAvGY+rWlntqG6LODqKV9NCZBCL1TqZes1dyOJGJ2k9lvDI4rBPlue+6P46y3xsB2T
Fs8EL5UNgQxA/nG6I7JN6cmyy+0PFWBfzRFpv9ugQUfIcQOZXNDNeyxNga2Iu8jMrH+QH+aSXcTw
gIDSKeRVE42Cbzv7fod8WusYhp9wLjS6qEQdkynkuPWyt9S/YqE3clTlcdO8yWOr52zZHzN33rCG
tG4aONAnze7AT6qnZLQX6jcbFyoT+7zsLRlVp25bZLsZDGaKp/Xmvc9/9m6nbFqrTVpgS4cOMYNd
CNvy8GSI2MSkTbWp85Wb9Kx9/jxIWsyzJeKdbrOl6vUkAFSnDAxsft/orOf0sBwawvTBlsxkAk8m
NVViwDTRNUYqrizBHgDWwwNH3HZij0jjBCX78QjR+v1teuNU7/s0T1qUwxxqeIWSzULcIvAxaUE+
rb7fjDQpTUg7gKtupyz44M6Gx7rwz4Im1cANJK6AlHTtoIw/B9aWMkqwRCSmX1DZypT8yvW17NL5
C5kxjaFuKvJAqzk33i6zmRUodrwQ43NS1nBWdnwduyaYLGDzztlBzgeUoIMpoPmkoj9300i9z/Fe
uov53hYVw/xNRvhmEweYrNLpw4KxkxLDKWowe4Rq6xPgoolMPx34AGsmDH0NLMVjuCrYeros0vqk
HclKkv4Wt7wCARX7tYLuyIyGryC1LuGJsB1djiFIHTq3nNnvdb59ZAu774bEHwpffzgti5eVZQ7C
gpfcyCqQLW08rxdCggWchO+HLs6Rf72jBZSuQlKCawd6KfacqjYLf+VZQFFQ4pdPVZEqhHt6TIse
DN3WJfcfp0RV4lcrlKSpXmlhOujRgAdTxmrlNAwixO3QIWBo1YzsckQbHeILKVsENN2W6JqAcXd7
XaNA+pvsjEGo/32BDExm+WG5U2j995s3oGUFJxiL5MCsPtFaR7owBC0eVgWSTu2sfNLpZbEezbKi
UnMEAa8ko5K191QjGajh+t1N7C2RfpLX5urVjk7/rJZ5KCkaCLMqCG9VJ18d68JjOAcjBnWSawx5
UUWJx4eno/niXJVKPqy9U2oOq4pvTj1CBgtK2AtDThCDIuNrve/pJsrYLn5DiAbViGDn9JU6ODdq
F7etl0eOaAVB30jEt9YOoOHPYT571xTZwNNOFLHZ0xmKAIzdPKCMxNgQrH+Bn+lUz9IB04JYwoAo
gQO3X3xGaX96SY0ZzTnjV1ZNpe905p/1c17CN0Zu23b5gNN0iQUX1OGBsvJELpoin5gMR0xWApMo
j3EsVqrDslzRuKPL9Fcu2HOqW6SH/KFmEMs1Aa1Pyfyh2GChl/+0Vt4ncKzdB8PryBIhKhmEXbkI
U6xM92LE6X2cRm4k5NWjt6bN/wVp63rtD9kvOSup3W5Zbhfj7CmG6V8yBXARb9Hp5CWM1OtClend
TIXm/KO91XgvkzvK75Y0gwcMa/xUOcc4FPRH1m8iDUtn4lKDIWSlGp1bgAR5PPGoxK8/VyQMI6Fm
E+98Ui09Y2CDwoWz5dmiveMtR4bqvjh61j8w6PS4ovDsQ+k8taLfftiesHoogDoa4V/cTUn0edV0
isj0cNY2m8bEl8nrbBmA9kFEqgxZ4F5DjcLfO6i6wkb5OXezDeXt4ijRcd6mZVktonm6HN1RWyL4
SKDdG3Fu/kRC1LJeucKblaC2oXLo4Cf2zE08jAEN69wH9R/5HkrMyINPClgz3gJ6NnqgOXoU+rrA
2PZTaKHasgYLv/NHh/MSzRFN4NMaEQ2ZjoKBS030LHR3o42U0vA46a+7L+3L8oj6W5lpJ+CzZxfs
FqL6DNRr3BIHP1DqBuqUWoZdoc2NLRAFJ91YNJ16SjCPYA5hmiFnWhnq3VNcAM1ovRCVG1B3xDqb
79nKxuXy0yStF9H2e0qpJQ3RC/MWSqE8f2B5Pg5aTGZmaIGIkZkbcG8AU33179ZSpkjE9NYR4DFk
bA3tFlyuZUYNWsfJFuqB7w+A2ZlC7hHWXWb45XdIkOEbhs3Iej9kWuFAct7B/VDQ/o2pBGyPohMo
iVpbTJqw3tBnHy4Elp+K0Zqs5nwoesVsv6E2FSXWUJ4TbBlMRBDg03A22LxbEcDObj1NsJx4rO7O
/RqQtxG3sgIV2ebpNBtNJalqxi+EOHzrsH7r3+7BtPvmnmWRQAPCvuXqGV0wC0rSszTxxVEjGb7G
X64zhkS/6vserS394b+tHomkMb3zAJ1e4ji7YkzOl5g18ZZTpJ8Kc/mJG9b3LrpvafvXMgjdy9Dy
rBFEVyiXyqh1dAEjTqa7BFjdSAxfpj0aC9o+BCO9Gr8vzokaeLf3CHXy/BhBGYNlt7J8t+k/3KLj
8z2OdN4TnII9IJi3IrZPQfkzt8022PVT3TmnfA/wd9Eq4JHF9CjT9dk+dpVh+tAdyNZ9vVVGkpNx
eN6EHqBZw0QOfybxA4ESmfwi9n7C0m+VLMW2Hfe6RY31nG0buFTcIP0b61kEQpWtPlIkumbLfWtS
Q2muM9zWO1GQH4EL760O7232vYLDdMPQLQKzyV+7xt5tY0AK2BTb5ydIIv1Y3/UNht9f5buftjOm
dHKJUpj/cMTO4uyjpU1me92OvSeCxCVQDqtf9AZpVrfGX0d33VuDVUElpu67GFQ6ZUD8DeeXF2DU
4MIJK7ZnVVdqfSrYdvD2jDPKKQnqJvkyXqHF6aa4Vj2+3St61j3EGmfXbEoeNrcexbEzX/iEJq3D
AUzFYbAZ8up/UfKqpInBdHdEQH2C6530f0g3if7L0002i8xf040ScA1qwzenOexl37Yl0udr0F8X
se98Dnfn1IvijmqnygKcPyUclu7cdRZRikWMrTf1GZcx5bWdkpD/wLxUZaxwtgvT2dE2a9FzL86u
gI61tbiYLNjcj5rHkO24m4QeCrfvi9V4EucucOzCq4CSMO3rbH8Z8CJZa2xqUCl1lwJyqHleP3T4
Yb83vODUXV38uJHa6DvaKS+raek6wamJUeHvMjw3GeLyeKaKVx9WtuswvYGBRviOh6p1NvMEIlI2
PRACHY4jnY3iRUmO2Q+NGANiuxdU3CYFQ0A2AySbgB1EfDQeAnTJ6TYoRB5w3+tVAFcpKAAfMX07
YR4Bpzvys+/0R7R91Ttq6D+AsWYMvdXL3nVYUIMNyysy+zPD+ifMk7FhY9Ny84rdODBs7M/pnSu3
mH4AM0VzNXmXgF2UTIdKjhJVQwZl3SNevCUrf5zpua+dJq37VnL/ffuqSIpQP6ghhOMkjxerRzIg
XuyrxYPt5CVHSD4PgH2G69+/EvFA/rAHlYwWg/hZeg9YN4IKpa2vmmgHNAo33uKHYt1A+oUcP52D
J/FzfqiAt49Zco1FIVMRxO8cM6ejyHmN11ne8n8sR4TGfcPf3WJuyZNfpQnmhC/Ny4DIGRH5XR5x
C0DoV6bO9mxWSOGOwxWllLDGkCROKAS1PY35zo/tWRqOo2XQfR3JgJa99utPjPAxB8ANgz9IV2BS
4BucGjctIZyMT7mfg38wYzWlz9HPWKOOQ9sIzRyrVFE5dVlcKaAH0Ki7wkv929DMV1NTi3zLI29/
B/rXl2gOb6YlfTQt1vXU0XMWR68T64E4lBXrze5SkryjV370aLN3JTPMa6K4z54fFQ7cZzlDKKWi
4sI00OwTz/lPw+iRJgKuVtjPswSYnkvvIjNKfR8q9X0DCFhEhyduV8FpMSdIwmsIJoVkMyb+UsIY
jvmULpoDRugOaWvvLM8GwtsWl6ZQfuhvxICFUSE4UOGVgPphX0Ytqjrw6XxTwIBGUR73N0xmOXeB
gMVIYf/YxEghs6go41687wAWGEkWVhSon+4kbRmhnGFBgMq185QKKxmkdjOGCGEP09g//ICcllTM
5iVtA/bcCi/q7DCYeLrWBax43k9RPOyH+V6M+FwyNPHmCmYeA2aaPnqi9A2sIBioST47lrjS2Fen
tBYNOHLgfpKiaGTaTLwgbR+26sxV6JQzLsqNfD1/TWdAITKtHWGekVIjDRRm2RbeoCRFeGstrRkk
Z7miVuZTG88MM5GmhvJ9dtn5AULfcesP5MTNREypgNEe59wQGRiN/NTvNo5qsyp2kd5wZryFzSwj
hFgoRoVpK6e/SFFSNJI8kbRrjTMzIn2B5GTk7OG2saGmeeBX94OEpHetUgKLUT5E6oel6oIeLBNq
hzbHyL8NEpnJfVt0GIYmmGmwrdQFvx1cUDCyvgsC6Rv68ap4mJj4tLVkW9pIIZ/d5cLX0TEQsdVA
dU1n0qxwVRMhvO6iLP4BEC74NoDdpgpDc2I4DGPAkzRdj6dbJJj97jAZIp6DK8QU0Da3JJGnFDSG
X2KM8+eIhcK3vsPkrj+Tr3mdjvRS6OQq6iLNJCjCQo5/MdjXsRTLRpwl9fZGifJqc8DIMSQeexfh
axysTe8TCWb8M4gIZdGV3hGqotZxpYqOM6Iz74UaxiHNm0UwX4wbPnmv4j+w0BkCbzqUU5zQBwkr
i6TpWgSiZpAfX2L5IEvcQwGJN6IL3McoI914qfr1UEzldzSXPlxMIeF9YwmcDgdwjtG4Y+B3YZ9B
lzAdQ969Du0l7V6FNlY4wZ7lmegTnAq6te9B6d7U/A8hsXymXIaiEt6jfjobVov6JJ+/IoN16Rc6
ngeEHAJvT5X3vp8JB6UQPmoTc//MYdzZLwi5whhrepDr/Jx+x+IVU3E8x3eWaS+J7BhuPnXqhFPk
/sfrq3/NIPV9urB27m4e719j+EaP5pvXJe4tLVfr+sbR5zydWT+iktqqpNZiZziQPoR7ogStohSO
eCOlCKJfmfMqqJfZ0zuwjBQ6KkaRtywfZHGNuDz5FX3umQMQVEkqD95KDNREPzRcWmHjNkQAe2Fl
xqYfKLFfIoTPET8R7cM52LBEivSZGIdO79JbdV5tGmTYrhQd/f+h6xOC3NC82EfGFCxFVH+zhFLp
4QVdUNd48s7VwO8rzNo0MfoXmXkc70RS5IdvfkfeizOiDuKJ7BaiTUvEh3XpwVBYjvtGrTKksUXF
KrGIohg2Vk78KvVQ7z/PueJSeD0TudBlvJ2npkg3pYMGtTXsmyD8IyyBXbsf/KR32HGTBzEIIAU9
1axqUfC6hmEVpMh5VoPfayyOBoe37Aa4+QaV79GVckt/0c7Hhe7rEVIFCUKI4wPf4NhBx3GPyhe9
Vb2JgfeouSaph5G64BaPKmgAr6Q4kDMQZf7v8Jk4O3Crjhpjp7kdl1ZGB/GtXfnIBZcM051hPMi7
bl6ob2xB0a4+CV2txLxnPdSfVRzFkgfy33evfYE/qv9lPHl3CUaIkKFA6CFgwmqQp9Yjaf6HbzcM
tsF7VAgz2h/zB/CzLMOl+avl3xgePdA1aqwJghefBix8ekD4ZoQBx/jxwGapOoAA7i2e9Uq0hp+/
P3OGEMpBOv/VQSOL6VzGjsotn3nkkWPOxthws1fKtfvSroI5zSnXSwG2ZHOQVw3Bvgz68RntUd3w
U40XG/YKtK/Nn2SBFd7a3dsw6I3uvEdhWoxAjEMDAusrnHm2s5GKkJ1D7pmgK2q8akiSlb5P2yTQ
G9Qe/NdjRqyGblQhmUc4/9uUrCMhMFCWmuUdUREvdFn0/FpWekc+X/JBvarFDbwGrLUROqezVZN4
mErJ5wNRuPV1PiTy99jbYlVhgaUH0VSJM8KBqPNEapI/jrhNZhx2Pi8v3RTHoNJvl94q8Oz9yilT
umWihsJurg+IqEFtEWCw6bj5Hp5JDRqjhxAWnxVl0VTFhL59Hvx66Ip9AtkrQM4KjUNCws5+0TT1
3UKCRMuDej56p1+UA9OLAQ9umwmEnTj8KZB2JWwquoJ8TbB3GGU2c7B5ln4Ss/OMNFZDUtweLqhC
/jElYKoi6Sk2CYNdbRl9st6SQy4nn5t2HDyEkA29fVxAG2vvr5m3UzAGYfAZdrAt+466ZFBVlin7
de5iY2vFX4foKmngKCHwyJvQYq8p1GkAeskY8ujCoaAYZJDQob0Fd3+S4LBXx10l5Re/JYoPSluA
XTXjyGneCsLiWJnpsgE4VeIPzzSYHBkF5OsnCvSi7jE7moVJQwzpK/XMYb1hP+zEfP8MESg9MQWs
LYB1Tma/tCeUT/Hk0R/qdr57bmYSi9g7mztcmYGx2aNqFu6JlRpba4RZKYGPOA71ZhEUPJeS1yUp
ClYKiUcK3dwVzKrDA8tT4MzwHrEaXpMMVN2t79UOpqRTo09ZuDQR8m6+rxMaDOtRyFkqJ+jGH+x4
Pk5K831l2iq4M72TxwLVkDgeXwRGre0ptpVwZLQ72OAKwmxhe19qMgevF2+3yWPPdGl6dMk4cnS1
5zrQaVCHr5T1Y/PhpiwtdUKFv7bHFlDCsJKI/4IkQVLxXg64wWtMOF7+2SnuqdqlA28u3VWTLfIs
9yRBjGg9b2xU7AmKrv2Dr9JQxdCwA8FNdaGSlMCeXFdIOqdFcU7/d9mva40Gz4u1F9ZBPLw6Ck/A
ENTWIyyIX9/soKmeA4XGoliyeXTd4HMu55OQsgdRvenK/vzcOLW9eZvISD0sSaAxdJorY/f0iFlE
EnW3EG8Y9vdcDFfRbaKnVKCNXlnFq+CntTL8oOYh85tNf39t04vUO9uheQ1hKUS1Fkwws090YOZ8
jFyzfkdiec/fJaW81LbTuoy2KgdDJrzplhWbzJgTqeznxqCEVl/RE7VZi9Vmqz+g0sPX2RF743xO
Qptv9+j3zjOF8dZjeiGg0/AsW64ngJX66nY8kLFgexX3wYWtS7fWPjing/tPIoZ9oAcl4UUJiQ1Q
wKkRsw8z91umUFJJAW4t7ZgOZ39oPKR9MxtdSqPMHU4XEm7900EOjhkVSO5/u77xRwQimfnyqLEZ
NLiEylW6+Cgp1VgfTQVt4ik2YLBZS+KTnxNauQA+rgI8jat8c8Jf2gxmnWXyDrNLY/blPJ+UaVgF
MzoWhOWaD0N3zW7ttsqiyG8AyGdmso3vtouQ4dEHrl4/1rkPlmfFH3ubVRhzchd+s82alTMvN+xq
KXDqBsUWP7guWgeTkjLl1EDlVv8lfn7SVqvQ5w+GHvjC+szUvj2V9FNkojP0TACMdAKBCWzlbLqE
gto4Rh7jvV50HfwESB9Y5vWbDGOKCQ3uAlgXtZeK8keEdcoBHboIBHppvUphxgoWpdQqr5v8hK1L
WD0Sc8zHgiGDZI5xw1hXc1pBPFsV9GsWLGfydxx6c5cOcPGBkdVKu/7VZkZTOZ7nq4fI3WruUtYG
/TZYUQagE2PZ7Gn0CENPeTM59tc8WHn1g1JYK/tTNLM1JWbC8Lr2kv1hncYhWxdeSMhBbUcUWmpj
N2sa6BY4cMXfkyyFO/DGf6JFzkb3byXYhLH6TzgqH76cK9SynOCV0CehOACqnsAEQKmAts/5abZo
6DdjLenwJmhvr+TbcUTj3UjBx6897lGX/iBuUEHOXuOYkM384LXASCVk5QQTX/gm0V1m25XCBenR
uHL8ZwZfAiBAXEgIQ/5cszat+oZADX+3l4nbzyc3qoxmQEKqMUqZR1OJ38zXhVD6XkqkpPLrdE+b
SBajlwvwi5EvkgziWOoob3Y/4KzT/5AFW8yDjs56hAD5XaHKjX8PLppOP+PTJecM1W6niFeTbNfO
HmtOp5Eam/aWnZ+RIvHV13i7R/rTXJdYqz9nDL8j35D3W8+RND9G3q6K3ZXDXbACX8545HK0likZ
mg7jGBMHbTlOc3Dj/jtfYQ1Ag1ErBe2KO53+sbMWXnXpw+pXE4WBDtwftk5WFIW949Jrim9+O274
5XrBbd2NMldtcVYk6aBwi0GOaEONQVpT7xUZRkBlZr3H6pO79wg2mWXfCoynWludfO77SoxF35z2
RaE5Y6ud/4gfHH7MMZlCQJptAyprQnjcr/WWtke6nzriJJGwIqaD2VzXoiLoV1sZHnqhyjD04YDy
8nXJUTWs3mtBaQ9Jw7TWFL4M4ejTiCtBOg0GPXFQO13+iZgMPa5ynoqzRSCcbvTClBVAcZsK9nfM
XqRQJyWprLo5cE6f8/gY+JwJPjXEERkSunqFXldWpmT04voMpCzSUp9g5XljoJuoFo+R0om05LK1
k8Nj4Vw7/W0ovohRAlty90YEmNKTNCWw4TwRbkyn7iQu/wh3VBhCN+pL7GkvK9ykXFqPJuRY28P/
ZmxRWLEqoK7slHwwkdA/S2syzxCAB3nxrWQEjC51TaEfdAJlzYwBO9IBTyJstcZiUCvl9OOILB8J
XMmZ9+U3CmzukAiHvt6Js9T3CAbGMejLdPmRsxu6Yl4+dmZzhdHwE+w5lrOMtBmFf5r54AF9UolI
9OO6nuu88VpV7s/abgidA46+6y+bOegr7j3KPyN78yrRzZ7Qkn5SFLLU+S7en24f0UMoDn1H9WFq
rnIhjqUG9HwdiUb2zwsKmzBR4aCJU3CQVrUTsmgQUquNWlpJkBzfJjBRgr+q0X14FQh5tz+3xSb0
NF7l4lA55+r61ZglNcZEOdw8jtHiBaSmaVEAxsxC7HVYqU6Gte5jbmMfAIpi1zTYfFokCrtg8S1v
oTasBdNWrvSgsYPOlMFmUIL8aD85L6pfC1mK5VbWuTskTxqfEpXSJhjPVPhT9RYNit0R1WXNI0ay
mY+/VutSrWKzv66LB7mQ13/xoH/NAMa3o8k1AhLfIpzv0oF0A6bDeXUx1LbgXW5kOqg5lgkW46+d
/iUySGwYLBIb4EY7C8gbDWtcwCREGDkcfeltksns2Cj+HVLgoAO9s4ynxjC9dmGqDSQ6OVLZUEbz
4AxAB+H8RJTvwzQkU5t/eIinWNdNwLD9LZ6Q3nOCkNahnoYx9wEcakatD/sqwx5YM71DoPGZ2ZBW
h5VLj0QWT0/PTI2j2JqFtjGChnPcT9YFSxRVvhXXVdzDzu0jnROC0UqSZ980BrXkPbkjSpJySWRD
f0f0PziGacc9anEg/YSchCGrHkQVO1My0bAyUxOgGFmzw6mUZSjJzDTsF/qTIPJjQeV02NB6UMeA
hrP6q/W16dIKu2bRvh0p/YKZYzVLvltYiiQU5wcHJWClae219XS1bUlvfR6BhWUUmOiQpzWHdVEW
O+yxjIWTUSupil4pqBwcLo9VLOmEdoVVfi4EnecQ9poyKFVauoPEj8xdjAa8NfnjACWT0t6z9BAq
P5v0hbCVDaQpKTc7qJjCwFZ/+QhRaILPv+8aa1ngHRkjyZh5qwi6jZb6TVi4D08OTKHomElXCAQb
xFZa22RFMHf/0HDMQoi1lEoQLfVRKROTBTL9S+HYyGKMeRxbQ9vu2B/WcQWgxUNOZajJTDaaqLej
eJATq1KBBmOqDA311E0Ji4Z6fUyDy/tG1/4UPcmZzrDOiog+lz7s/pTnofCssZoydcUoYUTRa3Cg
nfnFugjvwui+earBFnFM3sVf8bwTEO1CX3UHu8bgJcSfyFSn4Uugzms2JFeVjL0CFpL8KzcxGVeI
p8EUS9xIOZ1h0WdLISyyno11TTtJ7yxBMBsUK1oumPxfIFdahPUXt/MxGdjCT6PfZdZhGZXNurJN
Ve2KX4ST8UA+CMuiN0hZOjRgvosMczF90bwk1UQVvXEX3L4BfT9jppO6oY7QUrmhzx1GR9H2Q5V6
HP4EvAZb9M7xrxQlr5Lg/+n9dD/If9TmDLFsSyx1G8b8MA/G27+9IXOWd9ws4rFmZ7FkR6X41scU
rk5TSPESiAavqQr1JVW9ZFIveIXM5yZhSyJCnHSeoPgjKlKzKIOWj9W4d15dD8vzvy4i40z7V9uQ
j9mx5sSjP3NG40+BPd0V9bjQ1MjIVCISZ22Gd0ie4vEbJiNCwUfdk4fhyoUtNoYab2Lb/CiP1jEE
Pzr78r9Z952RWhH6IsOM+X53lLgX12q6SnmyGsEmKcNqOAR+cAgaFLbGVksolYMNLfwBV3kZ/qR7
oMSaz2Tge58dv3tlAf8K32UxzKWnOHXK7J5guEEZ3lJBON1Mok3t25qE6arVynoUMn7Vy1zHHOg6
bDuJ+NeBR2dmQxku8KfeQmZp1vnmgesIISabN5oKV/NZIIhdUOOioI1yMYC9u1g7BJhp0SKe4810
hKqW16yEYCkOa/943632mAD9jMXxfcALPiUbdPCG1kGFXvSOUBCRjLZypAX7aLCao+KgP0t0ibo4
pTHESLvQN3u/95dnCG6dzf5Lgrox6FW3r5V8eQuMEuXSFDzDE2EoaPuZ0uplMLQqZ5GAoX0LeXLA
gQ+9VfrajKZ4qoXkGWkUxHwnDanb0HQZnuYBJ4qWkAC/EXTJ1kA0ww/q0HqNBq/EOQY6IsqmueA0
L3fBK96CCKglEMp/0ylGZBBHbU9Egq3Tyo91WDzI4rDMtyYxvTWeZOBmjn9I6RxGcRcl4b9vaZDX
YDuIpg0jwYO72GGcU881bN8AFjcLbiHRMO2L5Ddvavy6Way1n36q2VhzDh0n15/KKj+JsTaGIljT
rqXIV+hYdar8IbmTcCxtkrJitoQNLhqZ3mv+yasup8EUQmjgltgwgJnKBibrJm/05HR7upyAA1rv
uAeonCuaACJN9hVlfr5c7yWHazjfotEw4lHWxQvlmLwARzDbbBMrVIkL6tcC2vAm+TTSE4mb3LUF
VXQ+IPq+EOI4aI1xOzc8wQXsHJqtjcEAjeEklNe5Kqw/II4fDQsguxcQ+wQX83ghOf9sGlA2H2qZ
66RWQ0AUP/paYcYAPBVfxt5eGoCxUrmpRDAvNGvG87RNP5enUrbZ0kERxIzgdZaOABKjewRj4DZQ
CUrqTrdPqhPmVood39pjLYb4DtSS9P8hPZbhnrawF8GnyqLD2xQITi9Og28j9/G+/WyXEMxei9Vw
oJbHlbBzRf7zwnwy2avRLKCWixerUxKsKYsYYgg/0qoCqZ5ZQdQYgEHc2oBgc5t0OSV1k7IVyyZW
HEvKm5aw9cAMWoR3o9mrjcnEjsDZBTqhvVxhKx8kKSIkB9iNjX8H77QxsXZk3XPRNmScqPk0bLET
Eg7bz4RMuF028BAkWy1zIYDLy8HMNyFG3zc8CcEFofXD74IYNEN5md5NHqJ91fLDxvaa5gvolxrK
7Wsh4NJjjeK7Tu9oZ8DGy/5VGWY7MHmF7QqSGVheTq1pLXZANjJcHzKxxOHxL0VTowraE0CnMD7a
OTEp0/fDl63bFStKWNQwaojGD8/jD8JKqN1f2l7scIdwiGkGG+Sbgh49n8p0Fmd/SCW6P0VzD4qc
rqqSItWcnynZlTCkVOap9NrIHAqmxCwcLB+0z2FBdL8SI/RfDkM0xCsJ0TCqZXTNy5T6CYOLvhPf
qnQBUcfGON4SJv2qpFH370YFdZfVS4Nx9tkZ1hmPYmjHQ4dGhXZWHiEj45ZpHyj6U2drSF0TQgo0
B3UrFgicGqQBTjXheTGPvHFcc54kBtUlxMDTx/EYhxXX0MrCdHVpSNaqbedUalOUbRSE/ioC0cXI
U6DO6pyNLYX5aocaej/+vdrPl1V047LfUqnNVA59Moyh+DP7Tsbjb6mp1GZjbznJtteVCWW3/sKu
tcWwSyy4jr30AHh7mv4n1e+wTS+FAU/x5tI6Yx+5gjc8Ybf5/HPAEX41UXA+5JMeN7Aw19temuC8
0mIGAIT4V2d077G4HKdRyXMC521+mLmfWaFuRmC8DTE2izAViwtvdR9c5wXnoLzIR/CrwFq26uaR
R+y1Klw1xIUthRCYW0lqWXO663gAfYUzBjCXFkFBgdM98w+VlGkn/6Wr2PwMB+f+PcGsLvbnFjgO
zvsYb4Pz9hacPZxi4BnwHbDKKgpFOKFL7B2nql4Qpde/Ay50vID0sKDhRrZxNGjfpMYgTO/Qg4rF
FhundLMl78giMTPyV63clOPycj5dNKliIyu+9Lr0J0CteXvbVaLE7NC0wloFv95WORvrtx/y98EC
eVfUZs1PSFNiEnz3B1GT4l+OHzzy0+gnxu7dsohQqcnm7KVN+qxlz8Er8FV08N+NOjWI4WhzoQAX
7CLKtxYtZgDuAc81bAYdFjj/KreAH+j9byCbQYlc/YUuk9QFsbUL1xOwyQeN1s35RaWBv8vZFwYh
6qPMNJZZpS2xiDOXP2jsoLb9vGUyyZGAFCuPgN+n53L1jxxygZbC3kwzZw7H8h+gA+f4TPKpLM3q
xiG0TH0nCo8yKW/+dMkmUOj0v50vpO8WSaWjMeb36+au04ykF3aA2F93lvwx7S5sunzg2xgQt507
rqer9/+9KnAHaaRCEo8CmieN+Qsn23A2jo3HKuTwEHAJ8Fkbe5ylkfbFNX02q8uaEQhSzFrXMKFV
qb706kaHMTmMKGwtMb4WuHMnRGpT/zwIpm9Wv5PmQB7MNpPnRpDTuOCOw2Qsw848rEt1FXYcGGPP
niwZWVn7R7MbyQJIUrtF6UCxsQZO50zBTB8bP6+NjsjAQFDlFWQ9oMLfyacr2/XJtc3A4Qeqf6EH
bInDP3VMdn5fxf2aTiu9Kgr3RB15KACQy/vk9fT3Ff7hD8c92q8xuD/kecWM/WF2dCQ7XWBG6Eie
cYBM9XbLUa8wmi/183RqJKwQM6N6nOEZ/54Lj0we0aSNGP4VZLeMyDI3fNfn6+Ih5ejjnvkbyX+B
POd0YFAMSbZqEDIJBpn8alouBr+VYQIQ3IuF4A/YsK+4LosJFVFJKUwLkDA2syxB4szzIVbr72vj
I+Hirp8TMxp1wDxHL6sBRTRZ9H7+FUIvYRnqd170RJcu/hBTeEr6acfxen4WX6prpElVSAS60XIv
ucjlKDHN/0q6FLXKvfDVCylJuj69mIL/XPfZcxhpJFsfxCjShuEXsUelyV4asQw0frevh+CVxlDe
5u3N7+uAdGhsvlcjmumWolM5sdax23nYLJf1/JXxff/QsRL3n7EM22HghTWnd7yDH2VFQHaU0vXt
uRmCWs8q4MWpzfyx8UUnfJPR4iCKR0OmJPnYEg5kRI3NJblVVU4suR4d+Eu7gVG6899qiWIO9NZb
4DH+0In/bmnPDSoDLJFPvotiqeqGWNbT8dctO7SSq+BwXMCrkkTaw6ILG7MJrvAi1jGH56azji1X
uoE54hg/67oDmZfCElPjnjPt9hlyyDR7Y1UExTLZMZHnTLzhM3aqB8NgPF0NLJdRlG+4msfFgsSz
LPE/hxnfyFqaNH2oLsfo1Pwt37WR9DAicX1g68nwQl6tkcZ8u5PGMYO8GZCAXm8BNKwAQ5F04UpR
z65C7a5pMjDhyB2B1aWpP3B6qgx1upV0l11aEcFiLEyY0u20Dc3g0uM8XDmLpq7F+zLyvip2Bau+
M2lLycDCe6oMGeepRfOQ1MLE9rJbqbIy4IKGODKd14ZnDux0axpW+HDfEgzGbv36F44RjjBMNmpB
p1YkwbOshtzk+l6d2FpvE+r6eUPqhC3W3ALstqvgvhNPiAWtSM19fdGLQ95js4cuiU4ocTgpQnZ/
VGe2e6CH6q0JNpleTGnt5IHnsJ+hJHZJUAUfqUs46yFweHpzR3UktlEjmFvbTqGjcskoBGBMyG3G
U83kHn+DNUuZaFIFFDBDkTtEaLnJX87zJ8gFLL7qUoqQ/0I20Iis1e0tQ1hNAVDGweTjWRYYLMXF
Q38K4XD5ak/0ogrr5HocuBMbkUsYY9DyClMKts8GZPGq7IwVtMPEGjqwM7wGXkmXeQQpF0VL/jJ9
yfjdNNniYJcbbpG9hdatPeo512cuP2xgA8c7RidFkAjxhavhhjxHD6v5ReQHQV2JKsRk4PGviKyE
zpMT6RemxTBBYO05ei6XkdU4apRvjosoliIzv6hbyJ7Cp6UHdmqB4ubyKHl0XsZz1qkXETuds+KM
BrcvZ44Sv05T7+VDyzv8P4p7Dn9ZiNItCUa0teEP9Tox6zynnazI6llzBhlm1y0HH1coYqpBH2AB
RkTe8Q5MqAioPtf5Hh1Ikps5tYwnYdvGD1c/XDDUiEJ4HE2vo+Z6lVLMgAtzSIEKZ0uFkWNzp8Aq
mPrMlq6wAtQdX1ynYTbEWxALF0i/ud1XD4WSsQGI8qvMpluxtCNjvaexHPeQsWEePLzwh3rVZHcc
++zf1+uC+eMCmUQFfsgRhNdbFsgVGxIepDmaYZLedtZuQylFltWnEstrDvuJlhxCzO9V7xZ144vE
4yXzEnfk6oCDHA+NeuLLdxSbK0SP7hlJ5RTqSQKnrhf8AOJXHpPkw1C/HOy4nvcUc2Sr3BCJeMUQ
MHsOW3sVhiUXLtjtNN/ul/bZ+z4QpeNtiT6f2giqk6u4kJ/2NAq4nXv32wL5dztTqiieOSV39Jif
wLjUgyi57f1ll+Y5f3t3rDY6dFE2+QfrGjJ8TZce2bYX5+I4irx4glOT2Lo/2nJT47+ndGu6R+Zo
E/H9CsOciQ+Uf4CEkzVgRgnz9EfBu4wpjDVrBS9Y6sAvdGFvxqe5OgAmR2WvBKorAdFMPT/n/Ugb
sSmrc3YNDGEJRg1pJp0HFpTLQgnCgiil0w3g7GW287qTFUKfxhmd/qtsMA+1ifmqOIq0GfMj7UHy
CprYnNAlHKwsWYdn42KBXWnpjxmC3i4NAZ+Nh+ZoeEgKzC+jo/jIAoBk2rBf0Xje0nN5OkcTZ3+i
StvtyRmI5r/X1P4to8b9nCIlK1CxCY2dpjWR0chW23oqoPCl7vv3b9/rYS2fcIFcENBXuYAxzzBy
O9JXNtQjaEcPElk7syq88OpEdeZ/2aZ2I/EaBAm8hSkEHyEOzC5phx5HXInOElWztNGmvBl79edV
ixx6hcnmZRblL3Hx+eG8TAZQ0J+mQCIWJNntXIUwk+lM0rMewQ2TX1DsF7meFQe28RZsSJLsdU7F
EYTkfXbsaZsjbDGHjvmqKeZFo6UOTiiY4T4WjfQfC12uDkErZC66XoRKBv4RiYY0rE8RQLeeH1Ox
f1XbYizj/DclfRbsLniLM8wjjmXpWa4PTFDX7c4NolGsRw2yXmPak7vDga006ymnN8B1IcUV5WTS
IglnDRt1IX21Ig+Xi0vcIIxktE/vPcsF4mm0Rf0UFRboykX0FAJtqMKaEBXMt2W/JHYUDp4kHXFX
FQJCU+vOtQtShGs8wkT/wZMXMbabXhfU6lS8rViG/Xw4o+69qLXg4MGAkwpTC09frwfv+WaPlOfb
2SshV3c0YQI+Hn0GECWmp46WN3G1/smaKGS7TaTnATUhgG8oJi08R5iOfXtjmIQDt2T5JO/sodj1
mveVxiEsKdVgKSOpAcR0HuWFM+wuRQJsk3KVU0oBLLPZGgUMZjIuh8BoHtVfQNeDLH6TBPr9ffsg
1EtLc6vD8Ik1BW8AYyPFyr3xtEXslbD2LWyR0iODgm8MOpk90nCsaVK15KSd7/iHSMfukJbB/yHj
+1HB1csRrLR8pKshNH2yUunCjmDmQ84xbH9JuxC5YMInoeOUFuGsGjNpf1JFEU4kFw0vX4uqsp76
jSsXdoGWp5LYDjL8zzGis9fnxG8sp5LzL2eHC0hkE/gtrN3keI7/SnnEBAxZrgpJDHzlq00KNIw9
bPs0FmbjBTTCMJOkJ4casg1FATJglfTJdbM8IfIirTnewM0s7lYNAxcndQZ1LaXyFklZsyor48+Q
4REC93DlTPCQ/5mWZ5/xcUrQHirreKzqGUAQhbyFbiZLDdFO4XvRXvIOYS/Lbsq7jTsDwV95/ZsT
wUTvcyb+tUP/r6crYh3u3exU5jd2X23QwopW6NADta/ZN3eOJCTIxt3S4BrC1408hJGOjImbLtr4
g0P3b6ZZ2oAhisE7aLw1KYRcV9dGJPDaE4Wa1G5naKktAOTP+UoSsGcQYX4606+bQhFl0XlN2/hV
zaecs5TNjgyGiNCFv+ZnZFKSViLF7BWpGeJsySV2Mdid6Orxowk9qcVvUOmasJbUlTyxDu//nOUb
jXlX4XVCwM8RiJj8NzCMoHhlhAEaJ/N3GKkq4K+j4ySa2HXI7wr0ClDzQtspSqX8yVrDYspdn+b6
j42UJsH8fCBCyVlxVW9SzlxOGuH1NL9uUaYTW6AOvv+03AUfw70CQvb/qYv7vHlj9AgopdENP4VR
+/EGht1IFmjt6K+NawaF8NL/CDJAuYR6nTJLZ9S9v5Yqx5bAoXW83MuzfTAVURjFv/57zzGx5Mfu
J+QLy4gO85Dkt8LMUa1oCZXvB5rcMKwz3JtUlsNbUSC++UHHEKMcSDpn9NpP5U6CrEqrH+xYbuZD
OOLJ3SjWJOZOeajjd78VkcOfFFJ6O9o5pswGOl07EMykfS9sc69kwljXgI22ONe/FwQlA3verV9j
FgdRyTd2xS4A0iBnhtScpzFQWN8xkMJpA/d9hIeBCubOCX7GohIReWTRf3R1bTTqyPbOdcVoLl2J
XYaouOn7rxsZoZqBK4UT2tELqE9rKnkfH0k2Dl1Cp6P+hz8OJ1Wl021JwvhfK4knetl/hNr92DmO
thQbkHXSpBqf++SjZoO/agVOQoTUZRR1nliqT6GoUBI5HcIyDcom75+KC14nqzcgX0z46fdEQYe7
wBDpnQPp45xB3sresCoDYWGKNAx5puHEGFGZshYEXNeZd+vN4PUKcb8IlfOZhhEk2nigy42yWVkO
gmHAlrlvh1O0tbTZL+eDfUfmofW8JtGeRmlph36YRreCZ6E/xIwsWHhHYzClG8X2JHltFULZ+bZT
oOxEGXAanaIpmN3/Nhb/X1ro+L3V5dQVChfz+nkdXmKZBS6XUDyZtEF43Mux0wKyKwofKx0tkIuT
N9CusaRhk9Lo1otmsBn/gMOHkfP85cTjdMrEMUKdcSnjyYoa/AgtK5rOiceq6Wd72wK5wfStm5dX
7DMr007Ak1RlmKwoz53xzMe9iCBejtk77blk1LJQlGqIrKr82Gh2BU94jiMtKPoWUA/+O26lMufh
EYMzrLW78XYdLIEnEqNzsuJ/8M2j8eMg5r/S0kI125NB6YpvuyquhuskKyzX3lEF9qZgfMEJ8lW0
EF++5DzKs7zoXf+k6nJzKVadlzFr3bz7O78V4YmwKnU9aXYBfPsZEsNEkPLytHOYUW1QrCxZP8rf
jHba7aBFjyA1r0zXsQMjgcpcQGwh4uXovlUZuo/mF6kow2bVg552udmXxm7I9T3lteaYZ8O80C/Z
+JxAtIla9XadVu+AAT8iCtV2d/qnbZyhTvirfq1VURhZ2bcDoZ/sMGJY2UAbyY1ZvIyjB+XahMEZ
smQaxsWPncDrj5dzykjOOhvW7aMuowN6rJi9I4YfpGOxUUazaPISHvTeeEEyEQhaFU1DFPCtU8oQ
roBs/mmcXqFzK4ZU8Hf0KSiB/a3B8KNiJcmxOHQtofIRUXAXFdM2G/p5lvl6RQM+1ubPHhSIgNRd
rH0kOzyubgUvpaKjRTP0hG0PvQwRjjthGmdZXK55+WNkNFm/zSh/HoxKLQTbgKxrFc+EtY1E4UoS
aAcNPxwyhn+c3mwmYn9L64453BrRbPf+uCuLs1P7Jvucw9Cn+ZV+ZTVdgvaLsXhyxXtERxYpePo9
6VfZOn0nope4VCSbRVOaq9U627jjC0/nirRtp7CGgk3lYahvQzxZ2jMuyEtruT84A6Us0L86bQ/n
SGXYFUb0mpIdBTP+9OxAn3Ix3HQijRhyV/lxcAjS7D440quU8iP2PrEQ0LwGr1cegYHXY4KivQw1
FjeLlIy80oLZbt5dt7wuDu944+N5M0GqJ/Wpf5ezSoXE98vt+BhitBQ8HORb6ZlG8OoK20tPH1Xi
+Zfwo/7dDMMbW5vPnGzN2LeBMD7gIiKsf9f4gMsGFKkWSksBMtZWU5Zso9Fb3Icn5FZgXO+mpvIx
uQ0hKKacw9o45A1VCjZ5KyISsOdWYMU3M13HsT594xg+qzv9EyY7PSM4Rs8gMRzAd+Txjn6iepCc
7zQ7vcs9T8FI4gT33kRmNkFPfGFdhUV9m3nPrJCoawWYKGsbjDxWEDu1Sl5FyLEI5kiOBsI6irj0
92F0lL9gDa/Yh+/wi3VHOIKxmpexRAW2UxfUhp4Wkqy1lPoDnwG+m5D0ZPV2MXiVdgvQr4pOhOqh
bFWHxA534SSmLasF13eZMAOzOQ4Tddmz4UxkVVNDypS7i0EpHuesJX2uWt8Vlksv2kv7SFz1ehYc
bVnBiRyVJMag+o5m+BvSp2Ul1Dbc62gGRl+u/i7ApOfVxCa6kmYRq8fMEeNQ6RPjtwaevSMCUtTA
JkfuH8Al7KuY7rHGrgxOuRucMQXfUS9N7F2QeJ/ZPDKAdSPCNBlXsRNh1X2/BNYqsVQzh/yG6Y9J
uHA92FFrkjLj/LzTrFmHCXPNZjw2XdpUtOzd3tdImZVov38eXIIFN8qdjIYYMpZv8ApvNHS6xWLd
ueBeOHbl3pPx3G248SmEKo7+JADYD+hFPDR/nvwA8/UrS68Zkh1seAErVqXqkCiBUl6UzVGP9O0r
dvw3gfSVwBDZbfw7zSoyN/5Vzgb5oVrjsrC/uo2rfsYwU7UlbGGhzu3y6vva42G22LCPdui/bV+r
liLBUMbJm/3N+fEs12ZVRzCHTN9T/49Og4Qc9hqe+nzmFAz5ih+/R2fGF5WQ3TLwi3mKHwAmUXVz
DLYoEYfZNaEjGUtPZtsyTpBBtVQ0g8mseI7fgVOnCyVWy1/agIzyGE3F/H3xurlmvRXAI0BSQxO4
4dxMD/ZQ2+oy7SpchE4o+4yq2aZeWXN7X85XNd4JunEu5Uwp/NIN/Njm7cGWb9dzc9IRn6xyH0L0
tlTecJEjlCjDegwjdo0H+Cpjskch+P9JNQuFb5TitSdMRUej0vuFRVwvve7Kjp0Fik22sppgrvqU
Rou0ElpHyBs0oCct6Ey3aO3GORUVtGFR4ZtCIW/Df71Td+7QOOMbJJZ5CbKWGxklixVy775NbEwM
rUc6PwJWgv7SXLn4V81e4Em/RMtXs4vu9+pnGBAfLg1OK9T6BfVtVO0ZUmKo/SEAtHYnFlOERLYl
+osBLPLQWRbJryTrQ3LthbdmF+anEt8wqN6R4oCD0w7Er/mNX8KwDDpsHcUkluKfMQAMPD/YmEM9
0Stf9dLN1Yaqf0KSHtiEincPf2TJQtAER2KV4ypuTBP99YOWZdVRygZVs2Ub3iZ51xGCq3TQu4aO
Kv13k6ueFwD9cBh6TLMqWOZ1S+KVBPiS0bNNcU8oPq/JTWE5lY3rjBAeN9revqr1SKFmQBfzvIZc
a343yDn5jDAfUgYZf+PR4hR4mCiGRZSsBibmKGXIEJ5cUdTAYdA7dBadYXJzQEJgQje+5Jx+HJ7N
VTTdD0c34xWBcEZUGuUGs1ncHRrnruQCKVgUay53FZLSM/gDPIYo/4ZaGzq4sR2IZQ9VTMQXPjR1
//nau7skerXFjHLR4RwL85MDxybtLc9ZOtv4AO8vIIoQRRfn5gLzkiRoccTtgA6cAIKXwG5mMVxy
r0HEIM39SVAim4f4e+qjUwG07l5jz1d3Id4hbVbkzd3Qq1v6YQgOsrLM2mxJ1qCMEQ04vhfCLZgg
kGHg67L6tr92IPxHbp7p9go9s8cRvnmUfgTN5B9AzujZiQ7KeEzd0OT/UqNj8gMV4ePxJT/hYGz0
rExkttLrCdKo4/9b4sQYJ2Bzij5aWoWAgD48t/qpUabAlTMJcKIhftEemeLKlYnj5X/phBpVittP
58ayC0alYrJQSZwz8HuUDM1ivx/s5h9quOtNkSkKQzrbPFwmCeS/LGaBo4Cx6Kwkea1RHzAbQ/Mg
kr123V7FXZkNlb04U62j6OI+NH9j8eOvPBJcDP8IB4xSg1ZlHI+YN7mPjKDyyxTD4VJJC0i+c5y4
/1QiPYlNaqSf9Hk3C++O4QlyYBjcJrKuEAXLEy9giWn7GMF8SC/YaINhm68amgRIL14MY+CTlhZv
DtR7mwGWgrPfx7XWGra2q1wPQNNVFhz5CMtSDYB/M94V+I3tkZCG2TESgs1/jJ1QRXYgHEtJ91RH
eP6MDQiOwCdACbC6F6pf1mOXs0uuhWC74iZN2d0hdBJVrVAYN+mGYIfQQNQILYzhi+PiwnqSQSgW
HxrpMBzqqs0yJ4jjH0joe8eeFz8a8yvZGxkJOD6/7KECuoDdN8XkQdrzAUooh+81xkv/0IRofBl7
3NAEv/dNj9CHq8k5WoZuyy2aO7D4BE9UeEFJe+GbZ27zavhMhIFgtbOnC4r+AI7FBfGORkdMzKey
K/3RQjvVgXXsLAjMd/eTUFMVS3FJRQfjtiPKnG3ftMX5Y0mmX2Kd8rr4M4JpF3r7q+rscXY+rakT
dYTGcOBfAxfFmZp5gwBY4mGhQFsczCfOf1f52olknPx40Ko/edwfjEVuvDp0IixVIk7Kk/uEwDkq
h8DnP9ppDhKknBr62Z5K6OLvNxcoDJycrWHHfJLNkRjKfL9x4KyygeQL8D2q5ukFYtok03eyhHXA
lMkfobkGc5A415N6mvT9YPPEd+gvvI/UFh7SpU/pQaP8bfzOyBZbENaMwrN7I2HzX7G+p5gGWbGJ
MPME3N5xK2ZWYVlJEmT6krr+nPsNWqdnAioJ1+tmGxZ06n5SEpuoixM4Jd3VRrttgV4NeBrGUdL1
IAWRB0VZcK3WF7AYDDu0LFpu7S0jM5X4bl9Tv0o5wiw+XbbO7AgG1fLDT7kbxY9tQyCv2R026EP2
5G+/nvlVtH7J3cLSydDBPQ+QhEAC1O0lqVU4z6ak/qccE0+F8k5hFypn7FWQMt9Iagj9QKFkgbia
KDO9+j0FVqXNfTCeWY3nKwFAZaWhSAJOND5Ody6Jkkr7mLYn1i5gkmO/92oAQnT4+GA0/WsfMtLq
gJ8JeKiZFiyM/Cmc+vdHXK8604ONtFQ5YVNiI0XcpEiYniTq0xNAph4zLABxAKzSouEssWEbZKvt
gtaeDxgnzVgpvOs4C0TiLEMiRMAzsu4y2xbf1jXOZIGX9R6Bq5TssmUAqSDYGc5MR9rsimVecdYx
Q/AZmHWZ8seGjAgk8wWYaOw0GSwG0j/hRfynB+aSnLba/zLpS+1zwAzhmseAqoz6ChVVpFF4iXo9
pZrJKia73GhFJgeCa/HjV+OJXltnrtxSG723W7py9w6j4oML+r7432QLDPjMhhxmARf17tFe2MN3
nwPNvltqKI9SwHaoRy9geEMKOlUxt7Ql3eWlYuLXxg7m4fdf+mfbZ8pT5jqlu9yURCDumMNw+xY1
p4/fO/d/l49m6sJzTAfZo6C8hs5L7gax4mApzgfT4S1hHGxYH5/w9a4IHj22UhfM/UWpT4Vcl16C
ufhMdxWlD3tYURVd7jq6/WYTlexcGra3dfqKVrj3gFb1LSDwC4XK7AP2zSEcpE26e1hyzIemV4Dr
8r8w2/z83NLNwpYfu0oXFi0hmivnfYDTHCAKO3UkUUb8H0cmiIxF5GON8A6kE1iLT5iXZpFFDX7t
49lCouYplmHfqZskZB344wZVRvwOZVpLxYSsrftufhAAKrJvVAhtFBlbvd6NVbVhjwbQwEPkuInK
4Gd3dTQ79Vy/t1AvL2m3hjjpOR4oUEL+4P4A0GZKKG3Wzzj3xc04l2zOaWouSgBth7ckqCLFZmLd
Il3o+u9BdftCs4hm2NsPp/ssLoLhZ1X8LQ/0QppKn01HChEhMMY9kTJlZ2Cr14nP0h0vfOE50xzr
BGO2xWhazGta5j5p8rOta5KzVBmLe8WLsaWQVv1WByGTH3umQQHvGoHTJNbOEsD/uN09fS4A5XDi
20xLL7T27N7RtxsOViWH/RMWnBhI5e/5nYHaW8lOUD5XFZpeErDifkB0s437lwiuIscgw3WBu9nG
98ol70G48Eg/yuve7Xd3cu2UdWExGZf0olcbyAHYmq436KBWvwOW3TqFITAI+VUjm2wLnfeqBOHX
6duOzRdVOXmwfEZCNBuXJKqKKYZJP+DO5vgsaGd3p+RNfuX2QTKrIRiaScfQ/mUkE8eVLq9KRmNx
TtGbHCUdLwSqrjgLmfqiY68lEpQ259fDiN1+rgFNPJc8IALJeBhP18rVDcoB5OrIshoPRnz32HIw
+Xlmyiou10/IuGQbGW5/UMfqJUi4Gs76fyTYFbO/kioxdKXl/2LIUGIH7+5To2kLG5eeJHvMG3Y7
0WrpCwl3ZyRE77XlPmKnb+gvA/2JUYG/aioP/IUxrdOh+inyyA6LykBEb6c4qedlZBlzbL5gUqy8
26uR5r4CcBZPLbU74vLF5elLnWtV3n/4VHB6kj0QoNclbVm4qqQj1wk9eIAKTICzAlRVxAmu2uZM
cu4zMELW6fMF4B/eLz9i90aupzRKH96eESRAjrEI0P/X2tF+1ePLwpsv1IFji5CtUyuolc9uk2Pn
/XIdVcrhQvGcesDYJse35F2yNiu1D61/wppnDhJUuQusTInflZfJRkNDB+zmFp/ncgv3ibBcMB2i
+CmH2YyiZutxGxpIs4p6Ch66q8bh2GQNbwA2sOGRl+C7wJEVxSO4kCx5t1T/Tl20aR8LgYdKsklH
mlGnDPkEEkNggrAOPhEiq37zZIELGItYYA7UxrUuA7gunbXxRQVXdMhU6bO/BKzyf80fRD2Uu9K8
49gHp8Rv9C2eeeXYGiMwu1JDHPrh/foRPuUXtbm9PnRZmmoxVT6mda8MbSYh0rVo6kqR7f+VxUFa
Vc7A560CCMXOoQJ9gn3M9NmJ3U2o+kVFfqH2XO6Ekk397e1UFjqLPNbtYLH6PKrYBkdkpz92J6iA
ObJWgDM/SWhhgIrRg/VuPdLJtKlObVTAhynuzPeAA8h0hZ+bMB7gsR0GidEagGhPkmGBde6iXEwD
HclXr+cbWEi2Kpb2eYeLISxfRy6UjMu8exqKXabc2iVazGPD+fqT5IIvGMgYxuBH/A2frODSIRoT
8k6Rd0oUTo2DZbDiQ7Me303gs3i76PWQ9z4zoQhdhS+gre2cyJEDsKUnXS2XZCwTOM49D1yLcJzE
MExwNBo4u/r9SWw5CJo8zTKMa3tmMaOyA8BfHH+0BDFe477tfoudUn/z1arVs2xJmCIgmNZ1AMKl
YePpZHwJKVBltnKekfXTkwB6gkosKtZpLXP3SaQ+ZTRulKKOnoseFlW1z8HfeZTZTZzv0Qd+sBL1
PSZLZJk2HuE4Wl62z4+YeiMqZoLg3iGRcZJ1DE/z9TP95DoiTOuG8C/dgnJt2HaXPwfKb66AO856
CS9NKm7rtADyY7MUQ20kSHRSq92081yTAvq8iY7WS3P7cewPVKFmBQWx3qKjOUVhzh+m9OYNtGfK
Ejo8IK20ADcVm5gVcdrDdaDvBZ/ekOkruW3BRF9Yh8D30disfR9hQPoa9+kmlLsOSti/ugI4r4Zn
TSbIhYsbyuCFOHIvQ93Z9WcEtnG4aqulZosOoEMAVi04uRa4UI7nlRv2lEJkPUsRAhFfL50a7oSP
OOF/6ko/kSGDtQK9/ZaS67dzfjb+3Oz93VosOp8UrkGeNKKPTmtqWWYsREKQe6BQYGIRJ7Ke9d8P
Tua7mqK6LGDi9gzZ5hzhflNBgCKIj7HTCxjR347TrTLy9iD/Rv6wpcv5u2TlNywAt9zzCBqh01W1
GemR7ZBndfUwBwCi2GPqmCDLzn3QTcarN3tELo1h4CopvgpT+50veFHYchpMxcJbuzIwH8g0NPf/
Ny4Gd59XXWsIQH4lWTbI3Lu870/8svX9Eog9nkb5/JprGHejuqhG1VYyDyoXlwKI8jD/lvFX9SEs
mYvJs0QWU4UdZ63GiSQqVe+bLyNGCAFij30ZwDFq4mFukyCo5rqZ10hLTSC6dcawjpOl8xeOn61e
6n48lRvUToiGHDWWV3YAmu65lSOkh0lPM/RyP/2EtpDrZV6qav6mjMO7o6V3nsIFjMM+jROGJty1
7aC5Ou21Z9iahAHClpHqKSXHD2WzyP3txG9icILDINSsfL0h0Ry5qTMnD63nTgygLk3qfG5tZcFj
0IuIUnaE65KIznzjKU802lWCbA2g3dZ2V8KYXuE6PNDJBNxKeBL6SQdPipf4gmtlqvfPI68iDOZ/
dN40gWwM+rYw3fEx1/JZ0z1qPrTbTyMEIy/FQDFi/o5srS6cH6J2PMlhUgyZV4ErgsM4608NjTtn
4wdQQP9Tq9A3TUafrY5iLjD2KxD4sIs7225XHrY8V+zctuaqX7ow4uhOrg/t8HCqRCwu1EGbh3DA
HWTPbHPUvb3W+/oTJGnCO/8EgZB9mphK70lWRGOGBn9g4yDojArCO7497LQ9ISZk7/hxC7HeRZij
twxJmu/+Uysy+9OnY4Wlxf+LsJzF/8SOll6lEt5xmHykl7i0Ao4fZSa94AaPsIa5TYBz6quBn93y
ZSxgBfPSyLk4TlEtBcMpaNcyxFe2PLqntMCi3wXm2BMu1gecdzzJfcrO+ZYgSSPGfPyWzd4/XB6x
tAZasCP5yxvbWJ8LiNWRPzLH/nDEh4b39WY7dmHYwKaBnui9H/jplLGSbJUR2Q798mch9PKt4Auz
+gkXA9LGCbuMDELXMAACMLgPVJwfEBEp3tmSJwS5r9bbyJop93gSG1kmYmhcHxXSE6xk6PArGpmZ
5z5ZOiNYRhYTayDq/Mo9zb/zQQjOKc512y6QYYqSn0PVGtlHonDwZYta+COAP227DZMVxOFTsnKG
EE5rLzK6hQJFSM9Yt4lVBck2ojoUm+GGkx++P3eUYKIVxZRbTgO//+s4qQNzAKcoicAC6Vc9jfb0
76sTn0GPnqPyNKN8K9TH+UHELVPWHLtThTdWtniV/oRfYaZp3eBnTH7qzp2dtZWAHkf2L8+z9PUv
9oJASSY6/uxvQIENGtQ/nu393P+7YMFfYXT5yP4Mjs/Z3snQOYGJc/F8KqudDip4zYhwuu8G615H
VhfwFNGRXhd2TxYklpXu+2qG4+8rcKI6UZZs4lDXkB6f+8dS/w80Lcw6AAU8kEH7nl6a+memGoB6
gPQdWGd2Ay7r1Z92waJ30hQeWCAcRrlBXFmBJn8DfDTBu1oipmvJQAbZWDdW9bO3tzNHVVrGLboW
tbH3p0taSun7S6PG1+xMQViB790GCYr9JADbGIOmBMhDE/8ve2/qzZD+kPMmuT85hCSb4ddf+rf2
gIBJZWXozcGOEiitcZt4pxA4yB+yBhrrmogFEA/04q4exSauDmhruii16P7DNFVyHwdrA2jfKD2+
ATbtv4lWo+d3rsVe73MqZxaO5o5SxULb6NkIeRWuL++Lfj/VeVUgsUPt7zBbM5a12G7d1jEyEpLa
6F/NpWz7gTe0ZRdGtz/pLFAZrwc1ZfmpxqKj9mzpN03E6rOY87VHT+iTmrgNmET6ISZJdx6E8R31
IDPIhn2hHaIPqdKxPP4fEkSwp2nIlNe5DcYyHl0iWe6ENTLE43TSzwLwQRNKjvCGC4zkYlehkZOP
L7p8qw0kOZ5eUsBC1/V6quLHgb7l7co1BqNlkLjbnIKFvIlrzQ7/aDuBJCPysiFUaISC//RASsO3
NXfCabL51PuDXQlbmpyz1e75ewKHRY23RbvbpGYbbHBLRatUqELAvw9qV5Hs++hzs82U8WgarUS7
Y+6D0uCOsebfr2LYyrucGgziRrzAF/4PDTRrkROsc9Ibb3YMu1nBXPk6VhT4bjjaYzetHSC7xJyC
PnIiTojs5Sy2zFDPCl9eXzWu5zyfpzptYyUheexZyKeWO7hCrExx8jOyv7BSpwNXiKTySok4Ko6J
DfAPjEy82uJ87zeAfvoEOWfMNpFToMcOoP69tJsGUQHBlvqcU8CthE/CRduNk2SAlaaqUJsZFNfe
T8ikzpwoYiD8/tIVRey9K6hkbOKrtPe7yKxKxdkI3AhxscP1jisOGtlaslys786Hom4mLNGxEM27
AZabCMOA7ZvLa95Ul6wzVuYNHvvsazlGUyY8iUkzW6JJ2Mrs/gK1nAVJQ39gJb/l+gQu3Mjmzzot
vd3zgkdpM1a2fJarQTWmPT4XtGVWvI1NWNLisTO8dQyVgC8PQMMBa+87Q9l6PM+7QVwzpSQmqLbU
UvD66m1F1EClOrNc5MvQXN5rHfCLZoNcmIdyGZZ6giBj1JN4C9S2V7hXU0mlXP5+AtGx3VIvnizi
n806se+efuFT+kOAN/SP33JbFLBEYGtj+tRIE2Or5FHbsSBJ2EmMq0vBuC507ypANLIfmfEgnxbR
ib2Td/dY2bYKF50QxFK7+uVhakCtzIcKLd9Jz56TWVqjdSsO+2kqwMUl7cbOdV1Fv7Zxxd2FORrJ
1A30jwjEvAYoFhpWu7xUsMt4N/JX5T6+Yq2ohrxHw49CIf3ttJNE+F/Avih9Mt9tCKi9qSxoX2Lg
sH2OdtTZJ+RDto4Mb2Dx90Ht2w/JS7Sm0NKn7jd0MJKWis36Lohbj4t+yp4nJ6VtpV4gBIH9NtVU
yTj2KZMl/OVBJ6bWblzfMstlBxZ94IzVxY1RuQ9jwUH4mhI6JL1VTT7H+TuD7XNvC6EZ9Sw3OPdn
xlVUtN7oJSHklqKcz2fLVeBtx5SdqF+yyDt4wRfOOtG5h0WTUn25kRh4K4FbcgDz+oxtNNyvpsJw
kDUwjTsn3OCbXnwb6ex85YX3ktjjA7HlsbJbv3nx9o3tvuS46YDiulQEJ6Ut9aJDYxGSBDmIH2Qi
607VKjBzc98ryVfWTpR1GWjEX+jrQ40ucbr8bQznmE+2bi72f9WG7jVNXopb/uBv8bIDBcYCnPGP
2mN4TL06m7ZvXtAIdRURSwZOaVpM5C44AMZ02CMae2Rc5w229QohOcdRE/5CtcdznFyOxxW15Xs3
ksp2+oeZYtW+MOYdbCGPtoDZLkO9d8/3c7AocM/w8HfhKTbRoxRng/OisMYJC2P+lAOP9npgA4Hq
4qx273V4j/8piQ+n4KkEmP7AIr074FGStRYOl7IbCwMHpZjuyk4c+3DqTXRsaFTKX7VqG00/PGvp
ArUTQDMvjkMJTkZSO7MH3LMjzp5BEwyIP7s4m8/yb9yRsSRDPwJoA9fY6d1A02P9gezZo9iQA7Zb
MleJ1qBty+1sUwP/O6q4M4ljLi5Izry4y2VPhZSx61JEH7X6SE/+X3meRIoHq9upThFv8Yrfeu4s
ZjyIpQS/RxuoreJk/B3cuY2BWriow4dmRmZIO1q6fI8VOljcmCFrYulZV1OClNT8bJPypL3gOTqG
vrKPCPCKZDMcjt/vBG890ftk+UUHK5tTKFyxSZDAwbpZS/UM7i5ZRGXhqx+gIkPhyxVv6DuciEim
bSFYc8JUN3epbDroJo5lY9cAgS6PfGQFZ/YT3ygP6jYRtjg0yNXpnghkZ7GBTuSCnwTEkzU5cH7L
JWCeFP9iVHo7DEumibJNyBzUK5QJ0WQ5zr+hvoqQZuiqRG1QehpXjYaFT/srPpOSdM/7SLNDLoGq
Zi+EZ5rwcKTlzjMI+4eTgTOrhH/KPETOaTZsDNM38hgCG1+ttlzkG8PA3viUpItk61seKaPImVrV
ONYupj+CL4ou/SoJptT8A1edK/2oYkxrVsrnhiKNd+nbVF9JVrlNwrVxPIN0iM2j9FAU3OPKUns8
V9c70eFHOV8vBQd2YDHKm9bePPBxLU6Q2cwW3liE1Ijru+zNxur2kJ9kUjWGQurWeN2Uwn8kEI+q
Sd8BqdNmLANlbimdDzD5LgNcW0S/9CT8xnB8GZriNTIZjtvtat/IkrH+Kmo/PTNpleEi54/QDYga
5ZlxP7sIWdVZQG1e7mF7mgjfrwFiebO5J2Dw6sXuJ4+kyXODealwwngezw1+fSpzDEvWWr9CTxCo
1K5H4RvYh+ECjWkR5u7LR2Hs19HzH/7s8Izh2t6w2OupcVitO2cQqoopNkI1jeqiTHfaZ93iwubJ
/DuBYJwSidx6piZ5RriepuzcwbUTgUy+MLxe+P1N/R3AHkdROu1S87t9jCOgQ954Q+TtytpzXVrM
lqkungifWXayTOjxEBpFMcPCD2uqMshiAoz0Tdk1Dm51NyLYRpdn9dEfcNdUWrahVfNzRlc9KSYl
GpiU5f8LUTvlLikGpLwQHCuN2ihrb6O9/0ygtkBQNCKso/guZbkrFcD6DnYcOM+vxSBZx3v2BBlY
BO4uaySp63f8K6vY/TePUBhBi0IPKsjSt5uJ9lTpKE9qOMQ6xVdzF7hR95mLreOLVbW4ooSRUVPP
ABMemiVvTWC0GZRog1oepiAiwM13GW1QJIr+kn5mYZq4ezW5TotXRaWnkkYJ0mzzmHew/gYE018P
Tem/DrJ34ilXfTXOGj2n9kGcAAzHHjrjPBlCGkFGERWfQWW0M9cEvhoZ86wp40yOgr0Ob6HdAJsq
R4XWnDCz0Q/tMOiGVOg5Tr3ss1ZgDKmvI63opEVkTlKg8QIoDAGVNbSBHkKidXRbSHjFA0liY8aD
dcFaAS/womgVlqsmgMy6ixIXWl3W3qvpw+29Fmz8DTDn3r/qbu2aSGbGJnd6oM6Am+Q6ZgibGRrj
E+c0DIHdj+XpIce9crqGBCjsZ2CBgCoUPjnCShGRvaUMUCXl8pFDAvSMuR88K7j2AaSb1FJ60hnf
M+yolFBr4iDbEFcCUl7n7jFyQ6mp9IZ7793pz9zv0DUWS/W5wcsC5KBBLyCzwur4skFmQHeaT2dT
5/a3ofq31oRMRCVwEso7nh2DYmTkrLe+uX4VU22UaQ5erhf4JJKn0qSPg3Ssf0lybR4jmLLXCxjx
qhiebxDzv/Orjcjz+uoQH+Mb8c4n49ApGKL/X+nPSjPIxyNuc974P9ZezFrC4iRvo0a+F/5P2NsH
EAVNsXNZ4AbjcBp9tEnjXeh/xr/MpBp5i4kdALsY/Fe+7jtQqWSImzVw8JtfAWT0C4zph4q1b77L
6s2QTPG+5D2cd1YkB7tOyD5bsUQegcV0bu60bX3LXc2Fy1I8jnfhFCLAc5YuT8kUABmTmP52FUqu
OkCUVOhbz9hrSHeD8UDA1w5W1o6/9g8ruTHpZvJmJGuWdX6HLkx++OP7+Dl68UJx0TTDa1bAWLSt
/jfSHBtZ+5gPcQUNnBhTWkpbDCW2OVDIs3aH66p+l4nbooxPr6zxCD7KgjetaSRd68OOgXzbyZd9
aLdRcyHcJSjaUVJCkWH++LttqfKdBIdsR2CJZEYeobxT8DZY8EDMZAFc9OeVop6LFpDdVTcuHe1+
8XHEIj0NInIU0LZRF4lMJ5jswLoJ84m7NbCgW1ssZDwIjjimCOCrIMnoKKs/A9pd9g4SdJaaJhxR
pUMblVL2HcYI02FTSaW8iVsx/kS+4m7rYAOZR5I28a5joKAL+XYwTCd7GBs/GdAH5jCj0JGhwDMl
StcQQ6ANvLvQCBwINGE0cKZu5znq6YEU7vNJP6OYC68n6kv6h3zIWqUrVMJAOs/E1TA5+qQjpHca
/+l1ToZZAWCOl6GjdRL2jXO5RONt001NPVEOK9HFemq0M4HSCRJvhe8OtFc03wzkXbAEDO8anmW4
Xewefhtd/uKT5Gwnnc9MyyijFz1YjDbxFbeHgurCfLHoWZ+qEtzG+02I+HnEaPchrunEbzr260jk
p6CKY/KkF4bXxEIe+yllBHy0flzUEOKp5GAhNpLlmu0hlEtnLzftH4AO6O1+T7uuZALrs88cYRhl
q0aXO/ngRVFXs2kpOEFuOzccRWB8fWkGesyGxsK/VX2CfpGQG3h6h3FP3B9p8soO2n943jpgpM+s
tzYr8Aps8C2KTZp5Q7R0gZut1sAY8J4SX/KKp2D2SJ/b/Mm523xao/B/l1AmOjsPnccz876KoKgE
YV7sErExv6q2hVfGiytH0267oQuGCZlUqN54dDPN8c2Xw99ly8WrRJVmjydsFW+EPf5W5EDs8xiF
shQBt5/CKr3kvUTdKz2hm9iSUXyPNalZo/ldKFdKBUQ4hZFh+6HwpyZ97Hv1nvMQjj/R2n7BSU4X
oMrlbagATnrIJntSO4SGMd9RCw1Ii4SiMdwW0s5jbp1RknwSGZiXF7Hy6JbLY/6sKCNd9OSqdzcB
DW+jshZZ+1GK3sLP7jVeGP8AvfOQlBiyOqUWU4pUPpWHrmeSZdoJUsF9GGhwKJxHh6jfWpKgeYa3
cGbJHS6GaN1kjQIl/NplDlJ/dlnS0yDl5CE664EJOViphNWiW0MTpbR+wq6COYIDIYW2IGwJVlBO
vx0jHr7UFII570dv9zXGO4FSSkKNWp7PVOr44jzRVZtdQB+N80KEE5xEINtCA0UaJ8hSaEDdvXrh
2vBNiSXRp8KFpEKnBNmD/zEYFETIBYdpM9i0fJKCc+LEXfCpYTVJrjQmIM0HrpPwWtLjLFR7zwTH
iBmCrrgN+sx3krm/ed0/aTj0SSKY144uWRCj9yaxLu949YhPNzfNxg59KNVCAIj0Z+MylfNXEyEz
z02gNCJHJXn68BI+s8huYfFY4t+zgARSBf6kT3DS/Dc8hls5E8480IbS35dA77fOARusJGrY6C/Z
GMtSXudK9abiyKMr0miQotnb6OGUq87TFR3B88JQR7nSr/gJLZ1U/T0BO/eUCjI6/MfntnIs0vtG
o5/eOvZKtVhn8VIOHifI8s+XqSZQ/LGE6pTOlSKp5PPVYCgT3lgWWogrFnpQSZVgKGkqE0QWBbA5
IsFZACgvsySFGMu8HCTfaeYN/MMVCCW4FN/OnZkvWINmHTS2GxYZHrh8Bpp2M//z72mE7Kgy5RbR
7NxVGHwgCnxbW4UvIp5QOa7i0otwxku5dob31ydhVbFTd6kRVUF10Q8LwzWdmQedBkH677ScH1/L
gxsurpVlSijGO7GDpchGNmPbnBQ4XdwAPkEhgKiLko+NHmSubsQfvJ0sHATi8oMYG1QmaiV2yzKb
uh3w7ZVVkz69rlqmoF4hgi/wOqhtyooC06h7RKrRUtVqGWbwTIECvVSoTJx8GUfW7lQNYpNYvluf
Yo3NSS3JAP4gwLima/8zA5iZJjtl8d6kpgkIQ+aKNmkG4aExIhzhw9nlyk5Olxe6amLHC5q57PPL
nHMZGXyhJEYVKXUsQyeqx6KLL9krCSAZ6kzb0lr7B3jN3fl8X+qSWvnbJxQUMIBcswjv2T1VbXFJ
j1tJj4y6B5KELP5ASBgHF6ISuO3gcJw39ztehoyyZDNsUUNbugoJvmtw6ZhstABWTtTJD0UiGckI
7jTsFmGRRBCdoU2tg3iQxQNR4Wqqfk96XDSFDsHIFutCA2Uozcl7UqQB8PEOAwzMPsvDqLg10PvL
urLKMSws2i9+mLUAK0C7V/ikSfTVuN4tTpOkpJwcE0vC+MriYin47jFmM5a/MTjSltzqRZAJQSD6
wEL+AexAvyuIIRvPFIaX3w58khvNCGaQ7WLOfZOCbqL8hlLnImp1Z7L+AN5Pt7fRk6NzWjaKYVlD
Pieq7h8lFVBLzm6sWuS1V1JwuMwuTcbIGa+/C6m+1i+KSspQJ8on40mO10gnSIJtZ/ymkMMNKCnf
pv9WV8u7OzDWQVgmBqZ/9Hos55YCBD+jZv32MnSIQJZGVHXj4l+1h429uCk1WGgHtzJNHHXspId7
UdLf3pYPASDWSSAYnED51uEQ8Tb2GuB+c6WEf8SVMXNr9p20fYhQilj+6JlJ1MmDCPZ93+qnMuJu
lNSSRF5W7ffVmmkK758+UvvhuBgWsrV+VYru1C+FH/R82Y9y2jM1L6ReuE3jOSq99tvthPbunWAD
04W8I/qhjXhoiAUKjP1J7xOhDk66Ca/u1Bx2ZiOA1uDwymtjFD2/5TW9kMRIcjBorfsmwUsBqHC4
23Y2FNaRUT1lGO/kJjDxskgJ7v+T041eejxrNrTcl8arrc7WdroRdBTDNYif2bz1ydjUrd/nqB7f
Uc8IHdIEifshyNzJRqahroE2Q6J7Mfd+PcitgETBlkTr/yDLLlcIODsXlEoEccalDEiYTclvdQ31
VYU3iBi7NpSyTchA9bEDXxoSFzNKUTJuCsdmE9Lb+AFOFdi6Sp4fso2xF2ULEU1ATL6GXtYUn8ki
ttIuFLSfxwsExahYkxlM3SEgQGN/lkrpE/+w1FrgEn8Vl4xxPEV8PEwroSpccKDjYsM6S66SKtvn
BUXOA+tQEPEqqPdnRvEnLVfSsKJzymAhV8scniNvytwSImZEOasZfbrrL+TtYu97jKN5UEguLbFs
dIn070ZPP25usTo0C36+Y9PDPtOiEPZoZlLyWM2DSGrjzdexFRvH2UoGfCfJsbFmz+Yj9zVmhj0B
WhIu4TWOSmP4Bp1jFaifZ1yk5fqUpmBdLAxyPTKmyg0xIrds0Ost6L3oXgyAc/fOZByEjmHxFPGT
Yt0B1LkWnVSiWCb/Mx4qci+WOxL+1r845keKZmc3ViBEp9QIzuLPNU3eJ5Ly7htesPHu3cJ3x1cJ
5+PMwsFjnxOzJkp0UM8mfmF3uslRMWZmEWdCuSvdmBM35NzobKLahWbgrWKURZdQvEbaReiHiCK4
/yYCqYopUuppJf0uW24t7dnWBqdtnlaE1upTJ4pcPywMNJjBrbUHU7S98pRnXyrqsusvOtTknguh
BC1BAJt3rBuSpcWAPunq6TJFMXe/VCM6sEO0zJf1P4iQIUAqTYho4/PWCQ4dQ7lOxRQXq//faM+i
FoiXMwi9F2Kc3cLAFp6sOWUFv8K5Ri3q0ARJAqepTSK+KAr83kROJ2Lq0kGRV8Nm6nfV1q7GiJzx
hH22qd88cqxI+qErOomTFPInVjQWqW3NZY3U7AvZtNCv6M8Xr69Ec+9TgQi1qoMyDWP4j3nQvLdV
ouaGfF+mFLyo1Z61kHiO+5EU1codwV+Mq7SOt+EOsIGsLCsL9oMB/V2c5F8jdqJhG0/L3/2O8qCJ
2sQhdPkSexvtE54mHY2X+sURJOTxQNTEOdh6njMj9pVelPU+GgIPaq+gLk5dUu9FklEpJT0q3cal
Ocq2ysDDCns5BwK6tW9UbCtwMrRadOyi6fwq0QQuR5/xamNHG20EqcLjBnfGn/IaMZf2iLIAuliX
rys6laQAyspJ8yzDnFWvmA3cJejySzWOEf0rgKSrHE6oBt43/R5h3ttYTL7Sph69B3zQcVnksdU5
YvnMXOof1K7Vy1FWd6XGN8t/5hBmsOIqGKvu7NXQ8hs5oHhd3bBTCPqygvd7FJcM36evO4Gtgixx
HQcaMq7okLiLohaxByg+G9plccxkw0qA5DXyeDpyZxaEz8nnBCPI5PMd/g2AW3sXG51fxXOa6zyj
NwqXh3MhqXPd/MSrs7Fbvu29+vG2IZC6yPXbelDzDO07TnIGFuusbtLxTYGgz1gJpS5IgXB33xnm
Ff/eacu8OcFtM+7xfZMlIFw4h2X8eclbLMbVRksaVSM3bE5n9ppRVxsfep+TYuSkJICcnGOm07yF
HI8/EbVBlpzrWiMM4DrjQ8Ni3jlyio7T13GCAY2yJHlyKJfZXcizjv7ZytkESMwGNMBy8Uy/8WSH
pgeygQKEHHpBQBB8eP1aIGSZllzvswqaFw/w2X7u5/qdMDVCQDAsx4dgGy4Gwd5k0M2cs9h4mYnj
jQXA4kmuVjO4ykRvRywl4wG1dTmzpYehSSIMhuFRkWJUD5q14KscA8eKWRJbuRzJ2BCiSiswePuu
OF+yg3QmFYYwREfBj6Ul5J14reZm+J0KUkM660xThZ5lnRM2+HFOfaovwulTfSij9qoPHj+El6q3
wezFP0TQVkI3ON1I6cN1rsmNKG+piVecY9iZ8yW5dlOdrBfmsb8ejXhooNLiAFNVaEHJAna6uYEV
yN9MzOq8rKfyyDkyFQP7M1o/MS4ajqbQvSkNqapH34eWIVG0ZbAHa+9MVuNxJtaTgHNQiHliN75t
xo6xwuoOk2GqIkSbSW6J5OUIKWfULiF9CbQsigOHeatb9InH6d3GEBwxXuKVyiekGiWewmAXRJI/
O2u61rj1e0EypSLQbk0DT218jfnDPwQDFqLs+nsLA3d3QZTSYZytYFIM33s4IPjGv4zRYS0t7tOf
XxwSrafOWbjhSGa5hlR/yQZuSuQGyQS7CpZY6fe79dlLUjbciK+fxev4eH6mvax4uvCveWKCkMaB
ETdJR03YdKggLdh9ZtSRoq4z9Z1XJYz5yBSeYOaxpOp+RgyC+2TYiPBgxW9GZAR2DnQzHCR7mPgM
tEGALDGx7mjVNoSiRU7t2OA4Cequttgxyv+OMYRz/bu/b7rNkcd9DTyaqoYPClhLNYFHmdlqRT2S
FzWTj0O/FxLIjMzWkxOn+/roK/WNhwgRrRtApHZcLTa4Y4Z+/qgQHQ1IGJosykOYDohEzkR+ux/7
GRlo+7QJgyYbRpfIwNu4/Rn7n/ZPbp6/VgSPvCVOzGyG/s6TZaaA8EgOlmhiJ1xZ5EGZwA8q7lHP
knlrO1DZAFqBALSSKhutoFWBHHuZeo0XpCJQQaLTCT6ZwFxAKHdYrSWNxnlHrqQXL9ChAO6s6HBR
CicI/HixowDAzrchJDaNY/4XMY9R6WYaJ+7SFvO7DR5Tonv164WHEcgLHz56Tuka6cKhjRiPxROu
cqO8bTy8K+/hxhR9Sj/90v31VqEfS4wrLrLUHhfTHOe1VVpUHSxL0J7Bf4l0+DIo8ZCffv3aT3vF
5nKdq18ekGgXACUs35kNa3NYAquTDS4CJr8UcOdH4+glCe2H1A/gKBWu33sJc6DMhYW0fOaVRpK8
sBEEWY7lizGh91tcvK9BBv7jDNRPfaGg6ZBzJsElY8YbmBzUcKgGI9vVO+hfyXVc8+fenWuBIaY2
sM4dldufL1ako9ebU07OEXSe8aKhYLuFQAVYLww4cYwBSCXG6QqFe1XwsHnNlBPGEfcB0opz1zUW
zZejaA1uHsdy/+RQbGOkhS+mc24XGJz2YrHnIeRz8g+6CXlZNZ/1fFbcuwbfjJBW3irJ5AvOXxvY
YlRnTVW1X4MX3pAEMwuxJOyOODvXIUQucTkL/3WoIrEgogvqDe408ZBjljwnSRx0MKnYdbLq4zAF
gof6lZQv4oGxfRDMmUnMq2fXrZA5aCgs3xhXM391zj/6Q/AfnzyQjtUQkYShvm5kwUzOOMBUlWty
k+1sdhTldFlp5u0f7E1EwlGm4ujGCdjUCqGpxTKBQdo0MR9PmjBMz4r5idHoEYNcZ+QGojxmjlqi
IPfwDRTaXZj2n6a5n/02PGYCZFIjERCZ/JFNDG/on/6pQUMSeiOeQunTf6LYkO8vQW1I8+lie/u8
+Kv3qc3H3WtuBQqoTYZNO3BNC+1kp/Oc6yil4wJca2lgHUJkiAdn/cj6B+aFYMt93ZYA2BqdOTBv
8hrDjIrY/lVfiLGtAl3pNvKGQRYfY79DCymD8sgXRnzlGVO87qeN9+DxNHABh/iGT6XL8GezoL38
0BBPr1BOsDYmcsBaVNAylsVZHuqlZiP7KmzjRnoLIpw2zIuuSahOTVyPjo6zxWfqAVxB/7JdrkeX
iB37WXwOQtXrtPl6Dy2OeaOl7TxWYAe6yZ1yF1Ua/kN5MJABn/W4+9c2cykLZrQZii2hgG3s282v
q+TqKceV3U3WVOkiIhbH0PklmTGQpZnTkett34xIHOGVb/kjkQYah16yf4q6OIDgqZQMNLOsruFS
ZRKFw6Iw7kJqPstU8xZRUubtty+pGj9+UFm8LT2kkY/Jt91YnRqWI7iaqzXnRr72OMw2y+UNqOH9
jN+evlTNA+1D3Cb1Uwqk6Lnj5WnT9eAAPVz+ilAkWLBKopFwPsrXsHas6s5UeytXXLeYWG7238Hj
SvloF5Zs/1veZWAXzKAiEEsOB6lBK5AF+/zsNj2bglnrKUrQXWuqC0mMG1b7Y5Bttp/AKwLByWeV
foiZZZFC+3SLMqaPHyzQkdv17v+wt7e9uwuM5WppxuXYaL3FRpP4pUGdTXbbzCrsXOKq9ocTdjzs
/BsQtaBnndZqD3y3A40XQ3EvQz3wByW3zahhifscv6uILXQdLcX6dpFA/vzGx6qfMvsb8T0BxUMx
grzSTtRP7XBfxBARgTEoRwywMJ/JCebTmPGs5IzIK69Ruub5HizGp1dINKurVaTxzzXD7Xk+Uo8u
C9og/Sh6UWFp0dta3EKiG+yFDFhX7gz5ZQXH+YxQkMQMnI9m7zOHMsJxIGeOq+vifSefbytkA0oS
547ES27gxSi64he3sYl4aD3xLNskJGQOPGMHh7E0nbIdSY2rCstHNGgq2D1F8Klx6KoOQ2vKSo4x
eHs16BOarz3HutSVbIXLdBbBjMohEe5vcLPzucPOra7eSrOd4c+vZCG96FoaGHUGk/RqbyFQ1aum
Yo+CRjwHF2TkxFyy5XI9Qu84ye/1bTbVN/yOzu1SLYz9k9m+CLX/1KS6F/2dF05oWaDI7x+sUugx
dxIFmAxnuF/VMZeYDaQbRiO1YUn+GruoBKIlHNFpppLtNVlgeuu1Vn/pJbMBgKHL/T7JoAObv82N
uoR5zLI+4FQI/NCgpvz9Tfn/TxVAcfgc7PxQzHuzqQe1Dls4u1aHl6wXsoo+MpjnQytKM5R0jc6Y
yUKbnQ4j3KeQz0KNe7RruUNCwgH0Tc0iHqggWbxlB53CvOiP853LHK3DJdbV3hF8gwQjNg2TVQeJ
LxA7VcZofrKuxGXRoQNUbj/WQXhmf4IXkOaeh1oxWYVV1v3XEL4q6MmCSz/d65IfXpvfgzaQA5Wn
W8HnDZ94Pf03bEdnUDDQysEIlyz6rvtmZvLXbB0BGQuy1k14ZPkAoshuXJpV9vdTH9FsQVq/F1pK
szXU9hJAvUSbKNdO2T8bYBvgE1eVndjKu8gPj8m46roUUHmayFzA1cO43DBhq7wZPEIilNhRKzOF
HXHIqyD4hB4sKX2HsidD4p1K11woByfLWd+yMTwtXktdpOAc2wGXp1UYv17hV8K8zgiPghGfL3Tt
kK3JlwDsbLkMJIAW2hUXaQ0S4SzPgLwGNNMd4OSsWFejXV4YK8yMaDFCty3bSKUEViGJ53qMx2Y3
baP59ymHzWnb38auo/xTNC6FA5GuQdzenVrXAdZScrNu3vzaaMd4eWZkxEbpnJ0nIsfBn5dPseIX
gnDQj1NqM06LJ1hyBa9etBcQCbTDVftPsqEiqlJuRA71L8DSOzHYhJZ9tRXq+vwo3U3rqgW8JrsF
X3AmxNWgKEKWTuU/xJMFlQXF/eiynHkhFSXmkXY24qQjvrWLglq+EJyn7M9SJlociv9QWCE/jAPk
MyhTNhAI8rI1FNPT6f+pm2fAe6vFUxPcTtUmYejZ7zc9bzxIfFxHkARv6hEV4JAS/QVwnT5in8pr
kLl87fZh2WAZfkStZM41PP2yJ9ei3w3eFEALEKvpPtIWT5SAylhM0W9vwKzzYFq2gwGSKzJvRg9E
DMaOo1snClGj2jnlstyA98Nq5Rxb35MlAfjRcjuhmQWd4ou6OX9YpRYasO8DjCMMSQ4245ECDFY8
W5MYlvV9pDjlmjez/Es3nxbxXt/icrePJCYBHDiVAliTW8iiL9N2bzGW/tE4A7pt9Eg0iEVVhiIN
m9v1YXdwfFVfvOtztouw3oUdHsx3DfNGQa8CmuePFNUIg0CfFZ3gtQp4x+pCNZcHBB5MPZw2mgEV
Lk1Jrmze8EX72Fe8pZPhq2ekYkjOcgj4++dc+cykPlKwmH0Z6a7UmkG1E9ofmvBGG2KPJXzJO/VP
1t0j+95hoSXlIJeuVFSKHMC09HmDVe0X5I2ryPuyxNQphtXiXhjTEBiyVEO1DyqQPcwYftVnnG6J
1ajjXfMYCSxxiUOkR+PhxmAmcjxdgWF3E7MdjC/5DA7j/VgLcl361jnv+qMz3fdVBjN1LYerkV/t
JaYDwLoPW/vMm3PGaWe0YqItDicAAb+cbzyA+F25kYuV+e4dtVkQO3T6dNfY31KBaMF94ReHgbTU
6pHWWER6Eke3wSYKyPC5V/nDpv3CKNr0ei5p2z9CIP4q4+aiu2SwEV1BQch/KzciB9x7I5pZKx+y
Xrzl1JPkHBJPA/YrU+FrbArCO8QRZ1MMUg/xP7TG2+N9PLyEXwrnQWi2+MTZSwQLk43qGQa/CwcT
RFEzGLUnEvZBIdpMtf6JXKKIOIo/dLrv08nO6uy0L1uepJ8Fbq+wZGTTHI0UvXayih97dQupBNwW
qrvxReLugJG9MUEXpsaFzEdBprQ/kQSMWV9V/cid/Joz3ytehIuQD3Dxb6k3NgZpdtnKfuXDOQiw
VCrpU9WrD/Gg9KxDVw8JMujAl+BYN+4Zg2eBWzr2e2TfP772o9V8tk64YpokPW8ZVOMx/RFSUmqF
zSCcVJboz4MosGza0ezkZ9nZbD3WBtcHChq7bAUaQ8Io9aNq/F+M6yXrWTBllxxbQiqoJ/a8sRBQ
BE9sE7Bkkukxm8oA1rJ0a3rXsfDIKiEFKgPyZtkgsKQunyqU6BPu0lH+dX/C474OzbKNJHCyreTE
A4JFCZCtHMggBvaYOda1+aZ9AWMrlpr6Ye/SKafAZgp/581uSaLHISt9p3mB6d/++vBbJ/9zpl7A
LVTveYXAzvQsc9ICg3PgjiM8NUXIzIz/nykU96XqAaDFRz0nlJcE8G1Vet94ZudAFSJGHyZPje0K
3sxkQMK3tXcj58k74xX8weTbIVLVKKTy6Q+svTRLnj8HZpcbTvJGm7LB1GqYZOyEVyff8NHfeqkM
tQ90+pfcRUWVM6ITLXgZIyXo22x3Rf8kngBEXNBaEAUY7H/l4kBdx1qDvMCC2dRdCmWVP2OYfJi+
6eSkyRfmOTKF7mI+wqcZ7McsCYJRwBDY8mwxIy+PgltToUWLj1HcFGaZVLqc+5TBmbnxSNH+BS1u
bXYAACKEXtCOTWhOcfQYKvm0hOG/dfo3pl1NNIda3/ac+NKUE6ZSeimyW3INd3XM4SIj8ocX9G5X
XlmlzjDEFZPSbX2uG9NQW3f98qTJOBbvbKXMisLCgWTJlnkDn5xE1NLfNSNaB12xDFn9ZQMdSRx0
Dd4fi8zD/tnwCXZcnmlsXN2DdD1ZrP/GdxO0kzhtGTWw/ZyK7qf0Wz3i1w/F9XGdivkJWoUs7EaU
AFMEbkh8SyfzqQIUn2hHBPV0FC4sPgjA2juYjeHpJ0xtMDCnVqVKIbjBvcW0/8k1nc+d/Qj/NSe1
3xPPxuPEsCOW78E90iOyQaXW3XAp1vLbW3pXmYGnkhN/pXGTiZ7t1pARoRAQGDh1tyooj5N+TrLB
aOD+X8TLHlovF0teHxJzldSDGT4owvwKmmyA1No2P5sC4egyZ80hOrMKTGp+xAPJIBeXaYB6OpOp
zdnU/71LiAb0NTzTB2IkLKpSPC0TN8LWAN4IMa8edg3Lf3eU5ANP7CE/vBAdLzSS/yDdQjsH8GS1
mf5Hs8cfteZo7A7wmrATJt5laaLjhfHDfXqrG79mLNMVbkWH49lSYK8+YsqBHf5uBJMs9q9Q7bVt
GPaqSGqbaWFfCeTUgWVdo0Ea/lnnC9bqXoOkbsYZITmwSzY3cGnCWx5cj+ai9IoRmzEr09/neApc
FlOef9Q1b9wFVGJTflYM8fN5l0+WDkXEzf9ySCTL6T8pHdKUvGalSyconlpyyfBs46VkNN09/cmf
DWRNx0fviOfsY7nicDXqTka/1PLxlM3bSck3xOeETUEjTDI7wyn+sR4EtzA592iI1GTxxSRQmvjI
e8NlXArOxKkuU7I+JPf9F/fAqiYbDWh+mm8GHUNQvcLdbOzjsPWg+04+g5O6hPon/NylkE0WcihH
5rnqL+hyJcTjjjWSjYfRy4jz1p0V1YI8HgOvIwKAadYMvC6mqtYXyMXtspFwQ8L0BfSLf9OVdsoV
qCOeAv6nO+nrObpmaxpQFESW0XikjjQvS+Z0cEFa1cXo+WeBfNquFLpZjcDINetuoVaynO5jlIJ1
BGuJiGXc1tbg0Cw9LrFZgpztsijPtRIe6o3zcsDRESLXG+gWKdOQlIOx1guoUd+meio07TYq0j60
BjRJphyMK49gyvWXhudKVW13aai721Ou5Zfb5SF30o1L1+UGfKbhCqQMGTZo0eF/kiz2TW8dNJpC
TiN3oqrLQJALi11WmBcM6EE7b46taw7vplQPivzWh6Yav6J474nvzDoNIwz9xt+bsOF+lTIg5ORX
Df24YNUtQjn6wUB0rIp5l5ntzuuCf+4iTGHTmE4cmtwJy5i5WvQNiogF7fTh7Hwo/1cGO/r/8bAN
aGFC92awp+mUnZWQu8QqgKrHSj8PHo6wt3HjytRVU+9TB2A1omI5BBBDa0wgCljemM0j1jSUxIFI
AI+J4gh6UDn7nMnZXFgO+/LlyuRSxZdzQDdiOfLQyXLADYRPc3FMJgJIqpUhd9TW6uZzebHQN7Mb
lEDnADwEPMdTjITTN+zOdX7M38nk88nmD/lj7zraOHGfFrp0urGAp+bUOCwCws0u+gMNV26XZf8P
j1N7JNYvo019hIqpXPP4cF/K+CpxkEUsdXGbGs+CZOcPOzJKHzz0lJLCiaKpeyJ2vbcxXtHNNILf
iXygWA9MPcAa4G0lv5cF1qsAIwRYdMD4JN4Y6mujopD4kedsm1BsiDnZI8bEPppmtj88f+rF6MyT
ggOUAQ0xdopbhU52yadkNnl6F5zmT8nOpr6tIoFoPTu86KevAfVRv6jLQSzEU4MtkQupPMRow5f/
BO9CSvghCi7mMPqvpzCI+lnUjviHB1MQMKkprq4HaShuVNTENHWFtemFtHpqLolao2FBDiN7D9CW
w18Ugbkc9+IgoXbp7aQK4ns9SKZr3Y/zeRIMrdgs1OhBm09cBcKdwiuvk1mOCHD4eOHHtBCVe6wE
6CaMPjRrEecwWsMbUoxg0LZbCxGs0NXu7Ho8/1Te1rWfG8Qu7yDaT140f/4wI6+OUuMBcNLBlUB7
HPt7b/L1rk/ugfUefUWz+5u/t75w9PoUdJ/D/ZX1BpQiQlU2XL37pDyVHAWtUFLBM9Gx4C4brfgQ
X7HcL529sf45nXrf5io8txhmHNEoVb/We7L0Yg1eV2NEw4UCvZsDYGZ3VurmXBP8iGG1roM76xgY
XMkukqcq9/MqOYUdxRoDZ3DnQE06yAverExVrsPiKWG96FceeRFviQn+nvQWIPxhhjOeTeunfvsF
CtHwquNAQj/NPA2EjInU5j/ArPujFsK6gSPVk1V3Re6mtGOs3CgjbF2EmUCJIwaZJCzDRGynniwG
yOg0V6JaxQEoyZYKsZljQhOXVDou3brko2pebClMdGA8SqebAAixzU2gQIuEjIef9M9eTp35Unwo
ksw8b1SEPOQIwQ5X73/wRkih+WaTOq+R7K5a/vwbabCK6Qr5VOA+EEqfrhVhByxXnpNjgG326cdE
w8Cr+zpUjHQe+VrR75owZ6gJRBOipAOi1Xnm9ji+rBInC+LnMbuzfimf9lMZ+kRyIQUqFUGJOXO6
0fVqQdfX2KI/lohiM62oJ3lGfG1ThH4JoCpAebEzJLg3hmCH/hPaFj1j42mx2U+FHP7s5EXjEoQa
qkqvdBlj0qRPAhuqK5iqOX18zYi91wJYjd3ngxgOf5rm2JQzfgliDc0/4ouOe9OD85v0UvQReGjY
8CJG5Dg3MDUX6mDIb1+z2/s11+rCD4IsOPPDS6p6pLpI/iKCgqNhv3wfnA3DZZoSmCB16e2zg3Se
tJacUo/5SNU/toOtqL7/GuZEE5r91EoxGROtEp7HZ/Vx3xj7dsb04LEPDCWUJDO/0KYKJx/6P276
55Lb1IRVzg7Mdzj72U4v4OIx7pVvz24T5AcExZibHQN7NloHJhT77uPpm6XflzagKD9Lbxxo92wW
SKei8pGtiJSiu334BFy+xWNd6VQ5IVnjW+FjhghC4C0RjZsFO/1zBC9ixuqnWv++CyKdkuIBtVa8
fAp6/plfEKBUkO7LxTokgYG0+XzN+8+iM3yLgY+sUjYItcUZY4MOh6n5O1u25+lsbAMU+Bp9waEb
MpN16ditkDz0wECLEwXqR8wubJoCGmmdYwu+PLAO19dEaYCFf+LfBsU+NouZfs+HUieGuDyQgOBQ
y2eviEj+iMpDgxVFQjDPKGVWlLzjMcFeT6upF6iHQH71BXwSw7HKYlteH9BxDBWCBMKW4HuDE78P
YQmXTDMmg7jfJw1PLjFuKVfVvqF/CmpqV+ip6V1iBu2jh3OezSKPyjb14YdJQW/Vfkm1FYl4jVWS
ZWBCK5WjGFhNzVI8Mxfn86SbTAsaANPXthyOyiRn17/MCiJweVpzMeGAkSZrNxMxw5OIYnkPxLP/
s0bOiQeGiyyJqH10n42NnRozPpoErh7eaCgFXH7cDWZwl8oW9GUhVpVsleEazKOyzpsayopw2Exo
oTaziRJQ3dDxkJNpJlIKP0/vr0G64Gs6SzX1z6bkCB2vkke6LI97p9WZHXRXallXT3BSt8ZfF6yv
cgO82SquYYCLSLQaqKYKiiIHI12GPaStjpRXPF+D6AimbF/bEdk08hohC67WWz57eVlnwiQWOitp
53Kw0h1VSumSU3M+1/1Cqt/Y/qyRsRr0ZJD9Wlc9jQMtivWTz9ij5XKoR6/kBVZhVZgLYuCjC8py
upKTi3gaD/yZ2Ki1sU0fKIJFRxb/BTOpuUgnhoVd/aUwmhSb9mkt/3v5yFwoAfVDxpp7UV2M6c7f
YItgAihtXUeIPeXczUyUnydivDVaFKcz/KPEDFJUut6jO+hs0zPIg4wOnnV7ZEuXuxSKwkOAC1Pj
UNNUnW4tY/rAAStKeJ5FHU9alO0QRq5u9WRCy1jHnAnEaQKmV7r6VEM0srWBMjXo/Ue5VlEunLZb
uksE6cv7wLImFRPBjLOL5FACDgrbIc7RwUTPzkBw0AebB1n29hw1yDmzVSlB0QK2pqdTm487Lz5X
ZMsFN/EysJc7e6vLbnmGdcZPvhJg1j+J8XmV2wtjnxSMUKYTvCDiUuz7iCoOnxd+wv6s/QKlf5VW
OOdGwLNRBMRCtCHSxsc8e1Cz5RynfGIWPcNSH3+ZRuEOz/Q6gHbPyGr/0KWuLYZwy/TIZPKr2myS
YQmy2spNnTRexBYewQfb4q9t1auaW6cRzug508yRY5zBxipdm8PnOiYErYM09zVTI3ROY58JibK5
VQd/bwvvmkYajbmOwRd6GC4e9WYWn1BwrHItvqpjfhyNNH/RLWlI6rN1ACg/j3lC+9sBGHhRs7qY
Eb3i45mniGd9EvaIDp2gwoy+BDF9HJqnHCjLLRKQDN6D1DhRr6vayKt6gEzXF+tms8oUUfDM3Ylx
W7qtVR3G483qgGsIClA9UI6FuRc4KpPeH7e1j6boawdyFSuoaQ+woadIZpRJb7SdofJDd3iEzc0a
jm3X0SkVlqjnYD64tWJ3QxEvOF0sGSajBNv9VZu6nJu7GzVcPvSDuJ81QjrG8LA8zooHjuPgIZFp
AQCNcX/s9n+F4IcB6ZnLw7B7Ch8UH1wiCuQGfUh1hqwe4bke/oPrLnUoMQyFommYIsAMaNFDVTWQ
MrjXCdNTdhyXaOYD5WvYQtjwkLL5EW+shajWI23x2l2bcIi59ixIkZ0VYK76HYH2Vmr2K4tf2UeE
/ymKnWg6cG16iA+/0L12BvLsY9AocAt3hqlqCtJgytzPOCe3j3knTuX5b2weSTjJn8vPsK7iiBwz
Q7sfT81K7zxfuPpQUVAeZF/6VAgxH4IcxDmNkUEeMJLpW0Q4hVhy28hnSAXhQavPc8qWMC4dzU7N
L1PXNYrR3mD13ZQZwup8rkfJUcdEQp2TXsNr5XxnOdQk7B10+dR382swbOHHy1HEQQA6Uz4XXKbu
Y8xBQ779s/IKN+odw3AMVhCT7H6u95+QDtEj5pn+LnXUk6kAIRFIQXdISiY3KTUW1bcJCJHmKo+D
h5t2dM9UrGOwDMvXRWWE1TQ1ESGpLrEGp9SJx0fIG7ctUGdXKzQ1PX7YA5MDXH+GllJ8RLgv64uw
T/OhGBDyLSUXpX8IKrnr7XMaD+oUzYA7yaIB1VL9Qk3MRgkDnISJqkXnEnzLOsGejmo0jEMMOPTv
J0Tcl9WRpHyOUtX4sB3UOod9ub755OkyISoLMu2ghFrkymutezyJ0Q5VgcJTB3QsbVHdpB2uHyuP
JF/52BeTHJI4isjvKasiyNxPqvCmOp6LHypArtIAR14y5CTkbzVfJlY5TyWe9MVPka+8jaxapB3m
MAOEvPQHaLxVVzd220s5C++AbAxc+jFlODD3GeuspJae5nDT/BHMEDzry54SpX98fLy4p4rpVsld
JFmRIODMM69WhjMaF5/v4O0KP3hHs2y12TXlzriZoEYvAJmdoNt1auVNBNK3Lap/FSxyWAPoDkWH
tEV1IzpLYytgk8uSRtK07VjDvCWI9jDwW+5jMkL98x0mKx3SxrkjGtFW7+Aqs6C/8JN4QooXNtTH
xMssnN0BGyEzgfxUBzM4IuvQpnpbUWyC9RThbONSBpIZT29UHVxPSvRYA0VAfF2vFWC5YH39I0tJ
NOCSaE8cqO8V+giw4rwlxWIxq0yrQOL549UjE0hg0yxuJh3nTHvuuDcZrdsjwswEG5JopTKNsS+8
e18swi8QMJ3fnDiCLjVzO+Fbdd1kq/IJ0Z62JV82Oshs/eSJGUmeyfED8oaYUphL3pnJ2P/Rc6nB
Xm7qT48vaPzQ4Momv1TWdI/xYC+yfWX2BU09yiU3NmpmQhwweTn1XRRYTGz4wt239OmxpR5PBwAS
enqaiyXRb+pPKoIlyl/i7LwqlPkfhl2yNMHlEr/RzwhIvhKxr5zi0QNKYSDiOajvo9nemNURTh4/
g3OZneKEQhw1UjaTwiJaAqUG4ZepHrfS4T1B9Yk6pDJphFwaaK8XPOQ3oy9HrzwEb3ufhywHbHt3
JcK+ZZMakZT95jkOjrTAjWkmBnfAsH1oBvSXldYjDrGkSTgVcKTejSQMcGbVS/L3TpXnkszQa9HR
1VK1gVeFz3ctzqube47680dZ9akyqCdn/qTyM1lw3VluRmH1a6HeSR0rW12kxwpGX6akYF/UXeBU
ej9e8PujNxGM59Lcjh2qIoThEMC7aPTh1HMY41e+bFP4+X22DB2oaDmmGlkD0P9MoxhHBCbsxoj4
+5yEXSd+DLW2ShARcCxMBHmmUYyiqtbEz2leI/tLbVuCaRd0exmbC+By7TFICxYTchrO/T/yhtqp
saOHSSS6saxH+8E/ZCobU+G2poVb6z0vExkVk3AHJcYoMPXPZfxyXzx5hQHRvVYbIxbSWOSdUP3h
3WLO4gEtAC/X0Icd76fOA7ysjaZ9KOXfFC9YQulE5uZJInTQfGLY3QjCxw9eAxUCfMfZNlaeVg4x
7qMlOM0qLh4jET+ReKqUIv/avBMDXish/sxeOcKONbRLixLsN5vVYH7wTzJgi6iYWz9Y71J7iq08
M6VP3vTJG/iB6Af61LSo2a630ob0xF6wmmm4T8ERFeMvLnBc1jaZHRDLwWJgq1P+kdk0d37zI3to
zAQpKn+L5zsh3MRuyGXfCb1ByOoINAwKLA0NTwiWhymB1pzG26h+ioYwDabd0qrGarcwSYO6fKwM
0xiKy1BeGqzOn0UhPIWZ9WRcr5BcTcdKvXGV5OSEfZm4XUg6s3mGD+8Yq34uIeutQ7/RhJ68BEkB
0kEBuvFtk5PgN7hf096D3rGFMKDglAQHJSIreFNpE1HOBKgpo9F6RI+krEQnYQHbtIL1D4QupqdL
LPJ9ALdPEAW8xT6nmcB1rq88SK3Uj6FmiVsXMFu2kHicQF+f+41olRc/EJxckM8QYQGF8MG76WV8
ChDawAfKg/vpQpR9bOgYs6YWPDEHcVgWuLPH+tAS8djJU925gZdTz3x9vkDnVE3MsONIzUX7myni
9OS8Sc4+YedOGs1nyVIUtmOv1aSZLImQtWnaI28eXrxkxgvOcClD2p4eheYN3V1I7vJH6EIvKFme
bCQJwb+hhL5P27ZJ6gVQAaykQ0Oi+IOE/8F6miByFqCRyfy2Ima11bgMxgl6VYLiqrz3XyXhNC1Q
HojgePlrltpwxyCHDClmy46C0wcfRmH3nqQosf/f38coyR3NmUDnueQPWXQe8gd4ihO/xkuB5T6P
wbt/B3JTH5FPbZj5HVvhvRG4upEPBwRQhigEjJCVwgwJvsqQjkBe2lIsbauIBr8yXqOiIFRu0jqB
7e8IJ4yFJSQe16DhgdH0eVTThPwYnk8MntNx/UWg1TrZuo2k6IS0ZXmqjDTaaZylxnkaHgM/Ujqx
hHELQA6m55d3L3+ZUNAN5VyiIfoT69YEzuuRcckOjMAPIq4vT3vUIQMIUZgTRbVH/XkoTxaMIhe7
FTHYUIYLlyn4fi2MhjpWqZFxDqLZ2tN8bVje2hMOWMeogfUc+q0oO8PVVos4EU4ibAWjpPM34gTL
N+n0NlTm+D3GhJLzv842vRd29eN1gHlHC8bWIJzcFcV+4ETfExvEdgBv1gaM66IRM1BTKi80Z0OW
oeCj1oYG9XexVwdnTVb4iNpNYQIQj5VPOWx/eNq+5yiaM4p5OQmgPo/g7LtSQHF5lpVjVQIY0ZBn
btU4RUmzy+UUdwA7PpdFaL3XtFQprwSrLPrlwLEN+S88q6ARqUanzgkO03xgaZDGMS3w4wM89p5I
Y3IjPcObQ9tJbCfCBobTGRgAoHhqLfGrVKVOcXiCDwJViNRvGq43CNc0SkdJr2fvO58zKzCpJl2n
nQN9G25hR4D6VsmxLgwh0myGuerWn/GzERqetn7AMr48J7odWZGuyzgiJfnWykUo9uqYPEDALlkJ
cxAO9mdCQjfT7GDagE/oLJStPQL+Dy3z5tgFcNaqfdhVuIYAgXpdpb55DdTPtfLXZO1a1sWlDwVe
vvtJ7Orx6rCsx89H7e+2rvG3IH3pvMKk8ZXH3hKV/rTqyI53zOho/qPbIHUuWL5YHocxP5lyPEii
s8aHokmgLzHgYlrrPLUYtEJGME6jkzYSRSI6exigZAZa2fDl7ECXaRjUGonGTFkgFvcztb0kaJFI
jfLvDceJRJG9t8bIjDhbrWF1P2uz+a3c8oXnBAeA+F8fahjNygBaDl07q3xP9SAcd9ktRsmUX9+J
hZd16hXHEE6rIj7nhWgW6I3vON3h/fMA8StPXKcWn2p+fOcdlhapH6OO8ewGkc7RKAD7QeGcrk6n
8Gs7jD03wNuaLK+8MGH294ddtFHmO44AzDr2EcTsun53qNhKNfIG3aSxpj0+j38zRRfeijEACSxr
WRWg9ZIIRuGcFa92DvQSE7L8TwrhSiWJLxUa5OCRRdPF4kLQSKMw8n+BMX9cWDl/v01r6JVvTjpU
u3LH6qIE6BXjKFlwQPRyll3LUW0BciZEOXOB1rKAE0dDaiNgVrDvMN/evPN3WOeX2HSSJi2Jk6TD
FzqgIFIzIkkBKWsOSilWQUL9uElqrivWftKuDsUqo0wMROPRZ+hvHtC2/wqII+Bxp+fS0CBCnJBQ
irjPjeJ7so7A4yf20qode6DL2sqJJtDh0Zf/faca9wAjI7gjL/ryuX4RlYzYj7StJTbkOoToycBu
G7Nvr+oUWyjNc6JA+LziePpxUBXWMPDxNYrvv1HyJAg5/2FcadhzCC2/HK5qVcGLUes8cH/vKHeL
1cFRylFH9fskAaGT1mDoxnnr0mre5m4Q0ydMtikIjmQU0fi/403r/3sxq3oyZaQJcmklB0xtvnF9
7EemrsdaraJTktOkWegnJbk/dJpeHhhLKqGtL6umcsbvZWpYrJkVljiKTpoJDy8iOLqscQDQIgY6
xSDW8Td6eAGWqDmHns81+QzUe9vMkzeYpOJle0Q9t2ql3NsWTeRZggrXIHSZgzGNGXgGBkTZ+lTd
Ewr49ed3rBoTMkDVv6xbAYmvqkxwQIsQaIOTw4jTJL4JDZjuGoXMxAc3G4D9OyMZxKL3h3wlZqxL
67JRSnzpvEt0hSHjBKk0gr2pE/qujZ02fREeDkRZq303zXS9BU2Wgr4XfX1lCSMVu0kLutNEa7/7
0zQNH6QPE4ZWBXs/ALaxAeZ0/hsPzA6JjJCa06U2wDgme0ft6+KO/wvlNWFAiwPb79+2Xo38PzRH
3dLBsxjNYbjfp/Ssz2Krmny3Sh4AkCvUDod/TNX6omoaMTTTrdurFnoLPnG3yBTfGy5oXMp2J1JF
p0gSTg0aA0I/3JULJrErbwnWRS7bfaMVaKFCUiJ2FGzBELjusbMySPsziaDxcjFiWoocfjNH6r6X
fg7P0U5VCb0WgnLvhsOc/+341WIlBxzxilyMRbGRwxij1fWy9BUDNcY5jpZL+E64CBJsR89ZKnN5
nYDLAdb0Nbv3OO7n8gIn+ENebMveqa/Kh60dMO/JGNNcGcUzofSvQWHOrCsHzVZT9FJvrmBa5XXD
iD+iUOBL264ghR341+HE+cwZ4a5XlY/OMieSfvhW6T2G8or5sweEq5YCTwErnorgIJtqlvCBjcno
cyvpUBmSpBCWwFybAQwVQR9/dp85cV6BiIu5InfrUhSKY0t2EZdgOrkx0bW+zIrN6xnwcgIcPhYQ
mi4lI7+wJhyoZp4hAv4uIZo7H2bgteKckivxYUkkmyOZm4kZFOIJdE8InxbWr0PM7oL2fq+2yoGy
xjwkuJXs0yV9DnMoAU4SKYirsS7jN5HncHJ81dcpQq8Yg6qh+GlP/9twe7leX2XmesL7E+XYAu/v
MWp1NH4CUziPiZaZnSlju7TfJ4BqoJ/lUEkvlK9e7lcwQsb/d8q/gnjF8E99Fd1k1tNner622Dbl
2xHrdTe6AxEo9uTyass/7cliwCjAUQcbEftkX2aC/SH4Jj6ifKPSjz5sEV3zne0aVlVkfdM1BD7A
yG0e0oupHaM0uOS3nIHW/91vIo+Ev6dCqhi54AD7nZFKQA0vYbA9Q4CuWmkYrDAEzcYz0Z5F01tB
p77GeSmGqdBUmPOP6NbPZfXRXES6mvQmi7denYloWMlmb5EuUQCqncxtQFwnqwFu5kA/V0rIp0jh
7dMLRRnwU1YAMPD27COxPOUsHz+r/tcYtwhyVrTwfNdYZALnNIlpRGUHed/i8yHYV2UcdX6LXCLZ
rZl9+0dwMeZ7cOPoAvZh2pN074w4I8/8phy7O928Z1zuLTf2yWdLHLo9krqU3CJsBp5VXAFwdMNk
intyw+EA011isini7HyWYaXOS7McRoj9AOi2aRLE3AUhYF8nFcOD+wlfjFHilkOfEiqNut2TaEGe
Sk0vnghkZDZtqV4sXfD6YfWvZK6++0EA7YX0IJqbhPJf3iaNeQGFdvp9qvJlc0jr/utadp7dBvsA
ES5ffHVL2k45RBBDsL8L9/oIzc2BesiOWAmWVPPxAdEwsvQLgBFk4cvhc0gOq7PG3BCXIUJUSsP6
IvlTpP0+b96Rv6r93wG5dYXiNcEIZFzXP6u2pClG+ZD38sjPvhe4DJ/34zukMSy3RNBNtL8FsGmM
qlva2KXaJungNwXVsDhC4X5n2fmhydPVHcIh0vxk5R6QhpQNTugnyPBQJWBZe8Ydckicl5cI75rK
i1b6XJBGv1WnY6rmXnOJTvAXi/Y8eM6bSKgOACMnI56fFEfTo7ocmfu97732LqXsuxXlKwrVOzY6
dpgTBndyNclvaBkJIwmPu+UyjgLmvhJCB1XPrQEZw8MmKmTvESC92Um42jknYq6NPDnYE7zuiM9K
e8QT71PLmxcCPOF9KhQHbBjwi9o6QQUfuAEAd0m9t5JhMewUZtoURY5hEA82Yq4ci/P5YrTqutAJ
yfiJUwc+8xRx/qPjmwWy21eg+IuVZ3Sf4zp55ZlE8r1dxBxHQhDlBL5jUHtVr+Ipsa93suauZVHL
qZ3dyU5E/DdIM102FRwjQtQX0hMi5BjYDs9QRwI+md/tRo01tfJ0vYeJiSNO9RdYh1c0CFVSeqFb
26CuotyADb1bwt15L0fN5Az3oFZwY/obOcAciYYnE3eNqLXpGf1eB/aQakzjoGfXpcqnQCtJpaEM
QfUgJnI8s/1enb2uThWbYAnya0SRkjUCZY1XSKMSzRF5mBnZyyZ9k8dSi5xX6KaNOAaxzEPf4Ni9
WUXg0Bi8/pHxHVJPhjM01SZavWqnMfx1OzsqDXMvrZ50ArxVc0GeFfeSWC7mlfcR4U6GNppwMak0
uXbH1X1rUKuxOYsERDi3WNBs7RlLtPGfuC+jSY0OLAj1YQvLFLV+j1JocHoGWAGcztA0z9txqMBe
yPUjqRTTkUegmXwRwUX2732QMT3p3jB1O2Mu5VWcRZWT98MqaJvq/UIUzTBRwGalA2UKcZvcQXFh
uA6tml2YjdVueTrmZMYgacWxkjaS5Ru/5+3i+EKHbiyDCScIzKgI3TTrlHndQMwHX1urTLPlMtVr
0HoU0dgIdHwhH4x+DuZIVwNvJQPWlC1m35ROMjtwSS30O8arOhz0wVFwTue3xri0Vsz+YgYPxUaV
RKUOmd5h8r8Z0xXg1Rk5jCq7I7x9kgmS1EBdR5SxQTVAVSuACLxl7Wgxcgi+V5OxozybZVrutzba
JOuZEYg4u79MdEOOAraUnypPKOCpy2gw7JHpM8BFtQPzRwt3596LqlJeIdfU0nuRrSeGWZzvnGza
2qJQcirIap9CaZp3N3cUnRTAw/50PibxYDIZWWZ0uzuz4Wa6Ih1eoasuJQidVqxz4eGQsSwyzSPq
1bxMO0zJ/nMT0ZcvKjKJIBVXr5fWMnG8ZjPXlwhZEpROHsEARd3NuBAxIJ4XNf2l0K6q4fWPGSKf
4Bcpw/JAkK3YyPdksPNejdafj7yj4RfGtqmPGGqb6tlWcJ68jbmZKniBUb7Cgmgzf6RrNyvnOsWQ
yRYNAiS59jRh182/6MamfsccfUK8QFARCS5S1mwoNUS1sAMxOoQn3w6zhmh+quTtLw6Nuckt7cWe
Cs38IDTJ0hLHJnfrYnULhAgHWCM5n9rzRFzDkD+abPRqPUOtrzi31jMKmB1JSE4IddFS5pTvovx2
L2TAEOpbx6HgWBhrHe509drg8EvH/+mCsBjmd6kjOII/Gz29XvR9z6tSSWISP93S3esG09vptpEl
uqMFUPrrYxo75qfo58GzZh2iLpgh4+cWYTPH9QbL981REqBetIW7Owsf95moPlNCoTdUvN2YtUdK
gYo+UW6tX8SxWwrc85LR4ThfHNo1oeAa0f43VCr4KOKa7wyj8F06VAIhmeMqqGvqAj4Qc5tIC9xC
mJjw5ipRQJjmyLxCQnZDT2Rjdxbw2uvyCAASRzGegokITzWs9iCiDyAg2c1V4iFmVWBqiyuBIYst
41X2tq38eBiGKG721Xtrm2O4jvPnVl6v8QGWs0BN0P2f004yD0sn7vNIPvS1OFITw89bYFqADT5F
w2NtBhoI4BW/ROEEALljkgXeEJf5LYg/ZLNTUQgC2jAJL4OA8kMaiudoDTVMeglmm0OonyBC8aX5
MDnxQT8W4W0zR9bDT5xbBUhni1IOlz+dDY63XbRc7tqY9Ry+FWCdHpUvIJVlTf27ugOmID/ZFpkX
0NJWL1b8O7DZ4GGL4Yb8asfRWYmMbuNHjja8Lek+KbzuEXWzI5sdgkwkP+AG3OWLwOBpxwjhyF7v
uXN+NAvAJ+DU1GeryDMOgHBzeCwzbnZ3idt0WKUfudNqJud3LIXNQ/uh1LmThRaN3YjgMXmdBqi1
MHg7j9LDfXTIbXLRArAsO3PBPRVqBvlESyRn+U8790UYe3C4iX9Qx6914b9i6Zx7SNSzhHZ+pgFx
WtCrsmG0uRXH4htrO8inBzIJlYt+iRbTVpUVu3c/p+bfm1FpJML86nwPyhHKZS6JpvZvCpb4qL57
DQxLpXLmeGJRY6r4Wa1EaYq1ALONggsI//NJuPLesLmzSb+wtUfaD8WSuWOfAKrJrSLplwEQUIWW
7lUifD15badkjRln7Byy/jFBaNDY3LaXSxw1x/WJQ0ggEINziwM/mqGn4Hdot/K7Iy/kg5XnmhpT
63aVzP/wajVf19ghjkIrKCM477d65dPX0iIyiVfH6lguACeCtD/IfARs1iwMmi6BrTxdvq1Is2IB
yd9rQYWe/JQJs6tuxj50JDUL6W3jwOQ2LRtj2BuSBHqoHJ6QYTB5ibREYqoWtnm7SDwWxSgs3zXU
c3kIUEzAiC7gM1WGHlFO5zjvajmfWfw/O8L/NsdnAyL/y3nFuzJzUvnPBbriV7KLw3fO4yhUrYJD
dizVTm76YFnxhd2MFWF6BsCUZKVgUsVzYTtQeXn0oNyJe71RRUpud6thQl+Ws9XnVDHet5n9uOMm
HbAQ07YuhpJOzLUgYxmmFpblpDBxDXgcpNQ/IaUV4ZERgw9IhpOwFGvvMMej7imALdQD4QMDxCSW
bO22ybQ2BgW723ZVleqXNkgeHRgqhZsLkw7xi0galF9tFxbgSqpcBrEgaxRx4sJliaKosBxxvTZz
yvdSuGNS14pGmZqoP0giBLPHEGD22seDWhvF584RUj7UtUYNuyuwJvQTp4zwzRz6pKCUj5PZct4V
vUBM9ZES9by/BYbXmQEtgSoVnoj+0VxIiQu+JIGsBeMHDOiJnitYizr15o2fdcZ87AlEpqkrouTc
9Iu0K0eeZDrXV0gBtTazXFk87DCR7M7IUlh6grS1IW0/e+YtApcbLHLzi60guPhnmdEaijh4vq5X
kkCrlyfJ43Og16SJnHCvqz+KrLK8iyqeGqklNxYX1VB67Vlc5OysDEJo/gEPizz09raNBqvJYr6g
7wAI5/BDDYYC4E8cSGe+kaVyhX+JxYZdqLnpki0VnXr6/UNRV7AYdTMOnx4EUdnr3NO+vqWISO2R
ND2/vDEVZ8e+udQiZ8fNOlXrEOTEA/z0IXV6w1acBESrhyO51lkaxNaBvQfUJKC+g65ry/ePCGDH
/h5jdaUHKqzLtPqgnrmqY6cSZ5UfQpjjFy8ce1nnPkmybBh3ZMbNydz+8k0dnB8RxA+s1bfLLQWs
JItnoRiufmUQrSRSRwclm3GS9VQo9A7to02hbtH4AvUhLIQDNX/CUsLtLntqk8/6iTmf7U9zc5tm
+7Ctv29QtmIA16/U87Vd2yo1SZtLSTSJLQQa1RAMCzCbQs4RMKq1fLfJMjJvSBZ9/RvZcH6BEn+j
BWhdlLoblQsmtl/JYzyKk56RQ/DJsYD1RiPeXs1/NIZJtCCZL4KVK8trdqJ2m+ZO3DCSsoqn87wU
UZcPGM2CHLt3ZM6/XzQWEPBxjqu18wyf5TS+FOdG+ySJcoDTSIbFhizlxLyemGQLN6rnALTenMDj
vF1qsy3XNpqcMAY6uk34fWuXnV0QGuObx8ztr3e3x4u3h0c+8QXjBH0SSTFU1UQdiidWeUjVYS9a
p2TrRCcBwd0Zw+omSPOZkVwTCCgbPXup5W3JDgVpnRWKkwSiuG8fFFtCrY7wCB2JFyJL0AkK8oYf
tB3vhSQJjyv5tt7h41vmhIITQmMl6rTs2C8gOoTycmX7NyGOVDkeu2CSWq4gBTR6zfujSxQ0zsdM
eavTkN6JHfjYQWpFaFGKxky1+V6K4MAgBxeMDgUccO2mqrbhp+1UcWTjgZ8wKfjnYxYGWGdxBx6d
MYjIjMcRWkpwO8NR9Hq+PfzeEzSORPj2pSalfDwTZFW6DDstaQyteBQmlLd6nLGe53ZiuzGmYE8e
UohrkKvB/mSBuJ9CBc2fXiJTbrE9+Pke5gh3nzbf7XKJToXK1xIhl2dJPgmJiWmhX4zcl7e/Svqn
Uv07xKen2hKlDHZ3HefOcQLw6f2hiXPPz8aVFY+RIDbKJkC8p056UOaP8J2sGFeTptS237yNlfbX
NDa3qQObsWf8durl22DVZLI8WP0tVA57O9ScqGdE+5tcx98qawffia/5TBZ0lm3qa0D0eGRmS64D
mMpYiw69sZKepz+ehfx7E6TfZD9vfoKGIiI5OClY9P3PpR7/4uA+4x3DewZVwU8/DP93i4/HKV16
odAweESH/RzjjaGdIVXFHNZG9E9LO4IoSKp61q1M+F/eFnikHxCh9i05eGEzg6gQrCSD02ZiqqPL
MY6fZHv/dSoeRwCrNvsrfez+G9ogm7S7NedAiddb2diuEPBlYY7488OTkQZ+xu1FKy7L+l1itmhz
T/bV7Ez8AlZMIYBhvKicoD3Cf8BhJb01l2vNpjTCOqtW/RpSx5cE8Oug2A0Xx7bBGaSx72Lf52be
jQU4NPj9WUYHZ5pIU2X2+IM/PrMkjSl/Ms9lXcxDdYwbYjn3mfKZ8ZaQFiHLYjP6Hb8kAXyTnVFy
iRqpp9JCEytw2/wXKOETtmACRdYHkz+i1DofcG9Qpvy74u6wbClHmSi+MvMujQFXYegC30l+ZREj
OAO/Om0ONyL4Z3ySIbWfclGccN+eh7i+/q+Evm9RIqyZNnSrHsDildq3ecCzUCPwK9Mw+dpmp2Lv
iy6ZrgZX4GYoJqWslrHof9YB24QzdD/C9B6gZ7fuB5XfgawlPosyziORF5gqSPC7UsX9dC+gA8oH
2+WUeCKi1CYva7VUSZh2tNSaK/Z/Gz3r6fEM7KnKK7YKCpfrjUv6zujE+LRghT8oaRTS+1lmW/wc
lavJeB1rjk0mPqp1eSQLbPuA9gT8M7WSmNrBZFT9aU5iFfYJ3Icu2VnonSEuIuLSZg/IgHDwff/7
OXKtLuwyqBSDmGzc8JgmSHJWBexjXqgEjT1zKDk+BAaofokDsJ/vqUWlxryCrKukk7NPJ6jfWPqQ
CVf3v916J8fb8+8UUf9nLA2OBcgJAts+AdnnyLxJDdaBdGG1Yp+iqAxMq9NFCc0xdQEe4d+PUL23
U0WsRJorP0F8i1kTqDbLp0jFC2+R/eHFfACrJoSvnK8hkwMFvQeO8mM8DAaBn3HHWMMQL1oJ3i3s
R69L/i0VS0YxbURy6ECyglQoxVp5ggbswAdi3+4shB4XY2KZ9Zeue/Bnj/x7fzpq4SNplLNVCsgM
bi5PQLIhiY8Vxt/Q7lQG+X94/+dNfr3iZDQOppBchjPzVa9EKiXzq6FB8DrYlZwMiM4sIM/mmQwQ
uVe8cRp7IVR3GpOb79g/tqIBqrZD0ej4+mTe1ucmJSDukyl2sRIC03vdYsi672050Xh1Cc8Dz8Pg
5ol8UK86RtyQq24XTXtoQeYjYd10vi3AxmCrCHDhfpvWiNdK9Ia+fc7x0gr5kKRsOzSHg1vmswi5
SespwPDUvv2sHq0moLiMpE/YUHoSrg9+002av0887hDjYPemalxXn3HT2CKNV+cCEVHhkMyfL377
y+UsrkilgJucS9DZF6MuJu23yBv1tqAXPowH3LTHc83B9eiyAfR2CmGBG/U7fLzCv2rTNijRGotL
RwuQATDoEjeio7XeR9i+jGu9PDApYfWwoQkPGiQtY/SPNA6vTWwox+qNCnMcA/A4ZHP/y5K8dxjO
VTTnUZRlVpvg9Fr1+FENbUIB70HQyXk0L5VvcDx9sQWE+AGfSNb5Ee/d12UWtuxxnbUT+zHc3kgH
hqdPBOTLIRXQCMdxOZV327qGF1N2vdR6xhj8I/f+MmpG2eg30K7ZJzo5opt096J9mB+r1k6RkHdR
s+7jnORfpr/dAWatOL5AQGDdSntRoSS/iMCM8Jj0bu2u38IucWaQ/09EPYlaBDHLcIh+REqbFj5J
suJ1MLy051WbRQW9a7Q1RNYbkx9xceh+E+qeaN6xwxCbzdffyWiMGwWnpWU2lAO7d3xrjzWMgQuA
4EpvpD91AVr+yf7rRzNTH0Vebp02O23R/fEVuNMy4Lovvp//vfO3DEo9RCX2hn7Fe0lrK4JXU7AC
tcCALI537pouo+DGTqb+TNex3ocmzTEneltvTAOwx3st784PWjn84/qxrKmYnu+Q5VL8Och3k58H
Xo6pn8smutNRZwE0ggQslSgViB/FVLj7M1iGO67nVr2+YqU47KkNSDwutF6ol7IQLD29lerQNAWO
dxptyKTi0h5pDJLchlAyxVbXKDYrS0Fyegs9h1WFaueBKlZTlGiF3+4yGoFTWxxk6SDxiSzO8cKN
/lVTLHRFpB3CSvoiaaCVPXKE08Th7lC6Tn//cnqDQ4KXaQYbZcG9lbf4pw1n8rAx2p9U51tsIdXc
bys8M455zeTL51eaq1TKl2IIprY0qWVQKEx+IszsJNo3mY4jmeASlobJmmiIMw95cwS++EvTpqHs
kvdyT5Ny4xgrM2LxJKjttylZ+KAZGptq0o5uK2BCAOqGHvn7RvSefVx4YmxF58kSnd07VSDM57Le
vuZIa/GEZqwZ97zjOr1H1wL4PxTF+Z3OtnQ2C9iJUrc7Yvf1ABFB3Dj+yYME4cphJOiPqH9Ny7ux
1sZKi8cNiG3+tBPc7+xiGBgksaNWip3ASx0uyUoKISFdgRH+GFi0VALDSVn4zjvTXTU9vSHHwYZW
OtEMmCnMRqCyJdaeaV2MPSK3PgOkwDGBYZmogEZthAWzdIp0DR/8qjNTpGL+Xqk243W+/MpnXcsB
9zTmwvvF4M0rYOWIQJ54kOz1Gk+DCVXLjyb32xSIdV8YPu/0ICSNTQNhfMFCZIix37UZEDM/5tHY
CarYIGfVxGVxah8zxpCqBF7qagy5EtdzU5EEs65CzKlyRKk5iSlpYIbQiDX6o77cU5PnsXOehCEH
b8Y0/IjQohKsnEC14ViMhglTRdLcs/UUOC9Mw5JMlkupGlgx4I6ZnGJMlIQRn2QdkMiHfb0hbGt7
VIIxoIjfq6l0smbGffMRxvYSQ4vWD+gWUYsOcMyDpSaqL7Jlq0DqdcatnLOY3SBGqp+2PjjD9KM9
C3bp6BzDzwIbCV+N1xnHxTsVgV1r8rIw7RlnHUuElOGYf7ZLugZnzq3QHWA3TbY7gEFwZkQQ+2lB
mXxlDD46CBvFN7vJVD0m8BrpCUW9LUTUcmBtfuofwz+GcdoFLYvGdBtTVytSFHEK2KbEFueS40Tq
hBQxrwyrvzYZKqJrZPQc+L5sM1bj/csH1bhzJuZEMS0LR7mgDTy6LRMrH2cZg+v3C3RzJRs0cmJD
1sVRpCdb8KmFdyh+XL6e7EOEep4p+j5bES6eqNXKcyjksaMXoC7hHY3E92f6wnmjOdGnKOsyXnpy
kmeJLmFoib1SloxJumqsEIshXwmVWWu8eSWNjhaN922C9gVBS9siwKidEGSorizNLcv5H7Mv8IHT
EuMFR5XeqZXfWbn3IcMX33t/GgKuojRdMBj8AdzafHaX7Ee0Bt8Tad6bp++6TFBcJz/WteksNGdk
7tF+78ptePIM2aZ3NsadvB8ZsnNCnCHpvp5l/z8fFH0QIH8i76IgJ0mbsFNlWrIDQzZybRqll/EX
o1q/YFWAvYVmBGbLHZuo/2OmG0GY1oUeU+rR/ScCLHRIOIurWPJo58+jtuZ6FkVrGMecV63LRNou
TN0igAXQO1ZWXj6rKi6HeY2j9o4BKIDtZD9IsGdR6Hr22rg2NcMEfhSU0MGbauMXLcD9si0MFdTW
9qXL5t+6z6f7FbVqcwwbCCA8fE0nAMJqeVjp0/8ydVRfq0OYsQ7p2rNabvFa8zrszKGlLTcxsAV0
bb3d5BzY4zmZXnwbQLCkHziOVrvBHsxEDD5ULVNcNZdzA3P7SMT11fyLXPGUUS90LZ6vhTm6i/oo
EO/agFgmPknJCQN2/h8cMFDRUWwCvtvMvfClOYu80izoDH/sRfmjVd3psIlu8QNuTEXsDls/upVp
DvFfn5ovqf3WmgOBbEYMlJTnWHP/roxPqJzoJ7bL+37mc96TYIpwWJ9m7pWygjUd/L4uzrq0qQOK
PjhHvyjv0FVkJxcDbxWN8CP0uqgaCY8Q5GcHAXcuTa4Lq4vHsCqlh225eE/ci/GbG4K4AUc0oOt4
FTGcyl/dt1JpXtfH2MCtGoI3vG9Q6jYg/Ui+ter2ukUqfYVrif2Ju8h3YEFC7iNHAiescL3HjqLk
Ezp1GACsjdsYPbQUOl4A4EtysaTxAzR1N7L4jHV4l6hdxdRik0QkKeuyqJk8JzPiiIuprdxlECcy
4k9O3qJBVRYgm8w832dm5s/q7Y/X/YK3txSdYrARzSODuJALf9/hH4mKN7/BO12FvWzT5LXE+trb
795qKemfrt2KGbwBlKqSjK7UvBlZ/iLa79vo8J816P8gIIw/yDSN62e4p4TYu1Ff1tgfG/zfFQ3E
UB4uOov3Z/on5BafuJ9BkFXLdjYRhwc8i/gsIV/33bhOrKnLBti0dpMAB5Jqt+9/G/kIg45L7zji
O7TnYd6QbKVSpaZ8DVKKb1a914XY+tqtR17wEphcy+aEYlijflauFy39cYJ1tgNffkny02CyVJ0F
pWE40nr+qQC9P/sfumV3I03wbrV02bsVsfdzWtwKgemcg2AVMXBeKmcp+iVqKyQ3lP6C2lATDLF2
b4sYaYoGx7vvIfJmovB1NuWZ1Dp9L+aD8ES/P42qpVWt2hONGwRfQE6H6HM/Cds8ubM9EE6Z5Y5U
oKiRFjuiihBAEYA2InHZCvdrqGwzxc13lsVMAJewR0lf0k390xFCelJj7H+8GQViXt3HvkkQGwpo
RvXBwJ7ARoiRtis2xlKFECi1/zA1AHwnjQgYzB36lnjcEBXRou5RTWWLtIqtnmCAywlT9+QyIW5V
ZWcQKFvWPIANMzwJPm+JudRnhX5o9e91s3l0OjCoaGjid3pwE1CI0N2OLTPaWE9c5oVEjkGES1xk
xCdF08KhNunLuOKsdWbIWH9A53eV/p8x5xt+Xdhlby8uwT3s8hXOW5YVob05NivOyimqyVqNU56D
vemH7JjxPovveZzrT20fIMmNx5muM82Sopj7aLhgmQicAcylLN8X3rG8OvPoM2KXNaOL2MA3aoCr
a//CVYPpljYuji+aAUhxbpMeIDIFPgFEc0YMAUIWYl3vEf2Td7cLaLSQh+hND6vb4ZXIerLVtOE3
UfYWkEInR9KgxUqrAJAq7EDMZxsVioqtfVvtg8eSiyCx1XZo1EcMFA1bIKPhQhAuYLoiSdb/++Ga
Tck3Mr68euHN7J4DMjjNhyhOK9Yn8vp07GpT5kHH6YjZ80rQly8WJgCh5D3tByeSx0JcQHWV04Jv
+Cw/1Hs+CvMxt6/qUJewrRvsiSYreX3BmMR41vnzlsDK+ISuzojk7tvrOnP4U0p0cQpunk2BoqzJ
mBOQe/Sa+lcngvBk+98PDQpK9hYjd7/zmZ+NnQs0cxZk2r9PfIAb/a3AoGbGgUkgZLSAPELrt8v3
BTZj1dSLsygzTDa66dfCd6gVb4R+30P46duZ8LW5J52vcTLcfZRlbHQsLRksbzCZizUN5HjL38BT
Tmb7iMEVp+GbR4/gAE7Lv/0XVxamL9PYx6bTfQkb5p2MGeVksahJJ2JNl3kzawoTZC7ZnA328Dho
I+Gen/DmMg5j+d+2/OJteTi+4pQfhBqObviMlih+8hWIgholZEO7lr0mvP39mAvmSSh8+tQnDb5K
sjU2301e0HCc+xUwduO+vl/aajFjWwu9Takcv3Brs725FS0jSG5z4g9cDW9M6VCHmn3mlWPnUe60
M6dnICfHtDGzVYCeth7HPyESCzyFOqe8R01D8v2AyArfEG5oLuNiRwEtd3W1eWsXkrQDmQ5wogev
aqBQM4Z7NZUexL6tkJ73XxLxYF9OQssM0I+FWb9whrzCH8zWIki+sUJOlwXYxvBcDKv7CW3UlG7V
E7Aqq28eOQSAcX3v0E1fX0hYM+r5F/1bpsmTlLJiaJbcsAlu+HW2ayR9FE3evHQpxLn9eT3qjj5T
Hh7T4zdE0I9tQUKWYLRfdm9a/7FEWhfHPzxS90eg38ejbSnBs+u/vklu+7JPwudb5NfWqMCKTrWz
nyfXZP53zAy4WPSph7TtxLybfFZgqONcBqMtFY8gS/ThQA+SdaufK76OpVjMEfFMh88wKgLw1/+T
v7GrSdbd45c7ePceiG5ri7iYT1Sgr7btelsFPSk3FfLVh756Naz78Yehr/z23S5fylx1VfDMJ70V
Ul7euaezxoElXQDxqzdZdIKn6JfoETNFGdP8bVm2d0llY0SpvqxcGF/cxyh9DR5VqJM9UTUhGSd4
31nxHTtqWLYIqMiQ7EGdCln0TYR0CKZWl8KmSBN+0CRmvkbOJVwlhSaMWmsWP188uKYCopWyHsEj
IJ/ZoAb+SQAY8zg20s0ltyCNFBs4C7/CfM/2/Lo82jM6vLnKLv6GxaGiI5pS4OdUl5NV3rN/T5y+
uApwW/lnjr6NQGsgvRRwzUyEiW8YT++E8wTS0tOSFbqU5ek2ESFOhCUinrELNwC1DjzQAMNxtqHw
0HMkIPFIFI42rJOC5RtLvz2qth46Se3674+XLO/zngtLVgauOKIBDBFMNbzNF/uroNsNF+LesDhN
qujEQR1hXt2Rzx4ScD1oDxwvJ8ykxTa4KdhThIZr4mgbo/3xIkJkTFJmTViM6xM0mvYT6KDUVVEe
CARrHPigbHRy3PO06tueVBUOn25UigwpV7Ki1oa9JBzTBIxAMKnVuc5XGGsI46it2CHDzXC/Me3M
aQpyBUQ3MtUzbSyKVZJQZ07l2JX59n8WtUcczop21lZydnryyd5hFYLpXyvdgLzDsW6nxTgjqBcn
XspZO538KH8hSWuiQYQiCMO6RWT1VbM+pdXlOb1LbsRWiV7BaM+2+yhJvPQQZ0LcXCLjNHEdiY2K
hAu00HmseUo+0ZFVrg/3lDHaESuqVfSwytFnqB8kMkm4Jy0NiX5AkHN2Amh2dfAh9ntfcUn45BdP
2M5YeA2tI8hCiZpZyqJWzm1KE47wpcLj+6XxiUvGfOzd/PLQgBlEzsKafGTN3bT/jlIEibOYXzQ8
SLXRG/V6aGE89IWz7bNayOZ0kHU1cW1BPfTjUDbCGtTV99miYYRhMn+whrYP3aXK9+426MclD6VI
FQNxnd9SJNPObZZi7fxy1J3pE5WqzqjW6XRAwN7BZ5+BwSLlC4gqNSATEq5g05UfrNfZI8L0CJMD
o1s82jNSC1nFOFAF+/mO3ZzFNYpRKjbvlCBd0b8ZLtLmoEmJqy4H74cgygoZy5MockVj9mBciqP5
tW+HEcTJ8+1fsnbbz29bw53u2ByhaKp8dsNATrEcDaLI4O5fiYwV4laq5D3b8qEljHB9/B0A3kvb
QTLVHLgdcxN569F+kVpvayOFvnz2K79DZt/T7wfLWF6G+HEQVeUPpX+NgMQjeEhfZHC5WHm1x+/I
xFYK/qT1zamC3uKsd/khJ9Vfb74PbTNZbw0HfW/xEWkGoqIfWTgYzDU7irtKJsr/oNQTMe9yspXK
duoxF5eMy1qxGca7idPP52hk50rHxpJ0GDOI2a/egKGeNcs2L9pCe3qLiEY+wEmpcaUHQ+V8yU0E
uCgXulfC4X5uKyXMo+iimxBMdY9zKIARqsv9RF/2PNCEDRgz68Y+ZwUE9cgEZ0JtXv+yoStjbLPf
veg1w41qXdbbQmEX1hYIM2sb+l3Pk3PPP6HjiQbqQamdcIQSd5Lc906uB1HrtLeJMBw/7jve0BZM
gbNMNGsZNjnOgwcygDuhokHTSdCemQYcRh3xhApYQzqkRzKRhutC0a2OyJxlcw4SX9MoMztD/Yuj
X0yFX2dlUZvSJsb3CDLcVQudfRFSTT6lELEzK5c1Vjf9iC1ur/8K7vA6NFMwj3QW4/VngPH5TQKG
RyEaR8Gyv1AtGRrHj6M00UXOo6Awm0bEGJ5suK+vh1rxJ5fluA88Nh25MXMW92+MVvViU4cYdeai
5WsJOEWlQKVRy8NyKTR0TKl39ZiwDqZQZUGTzk8sDHMHh1wtWkagvitIpNVuTVWUlUu1FbB+tMcf
cOxiRUTztWEJ5QUd+5vxomO07GOAeb/8MtxpU8UuSs/p/pVplre+1aElMyF4ZYdavw4yEa1ITZ7J
SnGYj+UawyyIMvKjmZ10ZBOl0eMZT/Fhf3gMQ4LzuVEvhg0msJfmeD738DDuONAmSNukGqEgxk+a
77igv+riQNp74efb3q9JwLD3dpMCcmDiXY8MoeLJYFtgJi1s/JQaxfqMVBNUS5bNglQ+pm92QC83
3kgC5uBkXWOUXfRZt31xoWXruppHt/r5caphKvdRp+Y40a18nrrdS6GByNcaSX7vwdhICn3PZmpa
fn5BE0MD9sD4aN4rjb6QejNekLTipOhUtswpQR78OW/rI42kCaHe6fPrZmfz2C4IGSyFQHJtnp5H
RgudcZZxsF7PHmQCmzilI3pV6yQX0DtNTE5DVj2NhE00dE/ZQMg/TdYzH7S93bxhWzVsx2ydH+Zw
zuV61iD/YtXaWme/HXrWmX3BqtXfwN/vfGT6qM+YYgSkP1y0PRS2E/UPGvzuQ3GCJikKWJLKLRlr
Enle3iCbe15uqgSpxcHVMqwABFxCCwqsPVFtbFwPxpa3lHhbrcUdoY6yvzvDzGuX6YJ6hu1VlLLW
lW2H8VANVkeLlIlhU3GDGXUyXhY39DQNkafExSbkjTCQrrs2ixi7SSey6jpeBIF5ALPu2lfRqKBz
yo3zvhwWGJhXzc7sK2W5tmCYb84LRsdAK8d3pgh2v2WDDk8A+KYco8nSq+UP8LRBQlcX8T69pjz3
Y5sV30KWALbdP4OM/20SDYiXJZaFEItD4eHAu1iUy1xp8M1K3oKwe03VrGyz8Zv+SDEBYoVTLf2K
cAXIQbQdq76Mi7n4XKsszRSu7mF5avgGYDGuRo5VJAOyhcR59u2s+ZTfVc1R7LMu8Db2r0goT+no
9EiG6YqrVjMohTAAN/mQvVxTxZlLq4VI6YHSp0LmHzDUaHIX0Nz2Yn3KntlcdT4KpOdmXSXY+34t
r5XuB/7DTwHa+OG3xduZua/gSvz7aCzkIVc71BkS1ivV59ns6jfIOG7L5uW21Og1ysiLP15xIfWR
+rX72z7oQrE77iidreIXUmS9BV5cNvtLjXfEkZqnJ0gF+2XhFavyAHkGVkV9ryGVMq8h2j+F0pvB
7mib2pxGfB14lIaL0VIS8zKqsiG5YpTPUjqtjdm23WBjjvwy0d2/Ou1sPtToRUqIFXI0OdP/547H
1251iexFhMhjB06bz3gqHlhC/0JJqC3vQet2QSzDQLSv5H3kuNDLQ0guCvxBTv3+TzCzd7uAOKvs
rPCuaCpXT1OWc5gAXd/IPqWFzNm7snIyE/GQ1aQDC23aYLA5P4Jruk6mbdWkRVg5z7MVHVqtB4m+
51N2Sxa+KlgDFfDgf4zHRYiOJuld/kRvCXtfLsWaX2GaZe9J7cffqIFbP87nM2evLYL9V3VFKarQ
MBMggDOQsv2QKulHw9T/hkc5fEkKrJuFzm5uQE6HC1GLLuomwNlI32bmBikPT7Yd9SXYnD82Ck5H
dumDiOTNkeL4Umdt9nGY507+EtjvBrRIWAjgIvkWp0aVk7VivkXpjJIidm7OMxkCNaaWgC9KLgia
7sdjAhOBiO5X9DbeitwifuCa3DM/4tUGoe7/FF7TgOUwiufkEehgCGdndL1q1DqUoSUL2Sxhb9uD
s0Z+b8IpNloS1Ft7yfxJlDvgfjShwB5VYQR9MYJ9xRsJIs6NOAnS6KWIhUcFkzUjsB87WGANecNB
Y3+osiwBhOju66oLgcO/16H0jwFsaGYLT1Moz+Lq8oGS6iCYldtWPMXqA9+XX7Q6SmDiu+S4ax7K
M72gvIFLkUF4q4zj6EC9sVPhpaXalJbzHEYLor/nIPD9qxyLzY0v5HGhsdJVazifwy5SAsp2d6Le
1OJdjkRDU+yZPro9RY8fN5jO4BdNrnI/87GqBrM9q4kp3Ddmfb6AKu09A44d1TRnAVLuLDkeqQcR
AuEGQ+qlY1nfqyC04xM5Ju2KM2zlF0Cud/6PJbtqQq8HLvX5XcaOCGDvZt1mTxbX701hh551r7EY
wqh3D7SSn63FbrHOxoCe23zztzUUD39IfDaGainP7yq5NbfMI6eh+1tE2NPe1Ane1ugczp9OSD6t
rWovIT+6fObbGrH9soikIWO+kpSgWHanQh4Dbn0ZUOtxjdst3sgPbo9sp1s2GIWlEit8bmCh80Hs
BELTn7Hp0weBq5eR4B+f+yMNzeqFsHjojEN68D34IFrBMJbNNa2682jWtwE3nI/srm6CZ8dGIUPC
C688kZUBh5HqQUKE9Khh8wnel7ugyxU9kYh99rGJoJBQUuHPKVr0O7lvanfQwlRi7bZ7JJgjO7aL
jKyzA0HOd/ATc5Tac/eC2njO2j6Y7RswqgyUDAldknAeooC/gHVp/9FG40es/+k8WQIT1kKQ5ndY
iVV2HrQ2bzIiKudxCg8cRASDhPlcMrmYv1+keE/eU6pvCjVhPYwkPIzg8LPpKtN3Ht8lIMSMXaOv
MfADsSLOnGZ8JbX7XjnhjIwqNv0r/1XiVQXzg9tzVKPmHBPFvSeeXxFfkmxYmikyDqwsUXJwgng8
3JJWPCF7YggW+VWw1C9vtHKwmDJm9SZVXziVt5YV/d/S0LOHit7jPIld85fAYFgzOIByOKbcg6vT
h2aeC5csI+ph2JuZVbIGnTau23O87a85yr8hK3HIPeifQuUHGGlzillzN7OewcUlf9btZiW+GQxU
JuGzKTaQgQgMcX+8kf4wkz8LPtu0G/tTwLrTrxIrzGzcVPoSpcZZ+WPkX+fh+J3nQU1BIUhI1XVJ
uFUwyascZuEQKuxn4qTgBQnP2d8HB3GvGaHAHbKnSfoM/rsz63344i5NCwOahmY7JWT+GUfvbp1G
uw0+2M86dSlNTueOhp7GwcubCxU6p9mfj8McMEIorxM1CKs4p5zCkt/++LrkT44/aiCxeNfhWjb1
FGgh7PoHsVCTMp3/BO9WgN59Yernu/wYE/xw8+/AMOjaG1xH/vlinO4AARpcBxoAUnN8u+T7mnZB
TpiwpHLK+xEFrs2ZyKYKsRQ4XUhFJDau2FiJ65U8hOKy3Njl64q2eT9XBE8gr6T1O6Egjsg+8DbJ
B2d7X4XQw2V+/XvmggIGE4GP1VaL8GMhjugNHVwTSjcZy985JS+yRPPZ5f0WI+T5WZWgolRY1xke
Tv8j0DsBktdwTpYD9RDBvT6j8rlwBVX+LWkwOlgorUU9nDxd/DMkoj3vHW/5eWj1An8A9EvfCcLk
Ek4FTXR+jAvw5RPS24+3lvReDe1bRtQ9wOjs9gkKUeKurcfNrUKlmjkKheGJgI/4k7731lWQ+5+T
uAS+4OeGvye2/tp194FcPGB8V79/TfK5IsoN6CgEDHblzcVLob14TaS6+YifCNVoXWEBxNVxob9R
r6zvORWrfDAXkslw53tZLH4zfbl1LmVKAxSHbqrWqKmKva1sNL130bOMtJ5/A7HN+kxjyN5UISiZ
Xetk/2/t0p/tAJFIrvPI/hlJpbeDefdLLlVfegouB2fQDGHF2z21bP6FTOezVZ3Qon3CDHwv94AK
ANX+MtM2XPu6TNAiQBXY45aPAp21tMacGIXWykSre0AwMMreHPsZ/w0N15lJ33o08/5Pr5UnikoJ
+Fa4XePf8jSjW4lHj8HC7WkFAIEEmVCFkuNLbpQvCBYHVyo1YHXBDENXD1yOZPf7m/yhiiW0fiLB
/sGDB2or0UjVxf2XQWJzd7kCu0JN9hAB/ZnZ1TM472xNuMzKHIGiTudRF2Pdh9Mis1XpZQiNU1hD
gYDi+yDKIRjwP+oi6bvoBGEVfihadmCfTwvTGk/+NXkrRmAhUK4WZh0b505DVjo/oZI1eV39+pIJ
kc9tj5fEG/D3kAttfJawbV9bLJG8S0y+ZpaBn9AFOITqBRDH9eFvaoEt8NVKqtDbs5ORTLaRd1sz
PpdNi83Wiayf7PpbP/a2A5ZIguYHNtneXmEDSDTxGLTeFFptPsMHnhS5iU4TWRnmgvP3k6f8MXFg
A3RHAQMDzjKk2xFOO7DmG84XWt2hphd/LHS3OZY1N6ws3ujaa8qUtiKs/E7iaVi7lhi06xmVJfob
eFRKzvdOhm6KJuZ7zlgs3qJP2pfKPcIB8yIW4PR7ej+a6k6n7HN0kWopETi6tytFSa7oLTgOZmLI
n6HKSTFOUzI8NZ7K/WUJWdeGPrkSzVUoq4iQTbL7kpdi0LWNRDqMdyflsDSVTKx1jHlqDoZNK4yO
TCL1IZNZTHRbqHxQk2wh8gzvIAgseQGLIFmeaR7AfhkS1pG4eIYEv3akWojrU1sond4dTYUmfrXx
izZyQPG7Vjkinruslmg51Hs0OB2AMPb/cqzpDkR+c3J/2gSaDteuLN57JD4oQLd9ner87w9ybXlR
gbxNnC5ga803L7ljRG3B6kX+hwQYVxgK/NSToE7oev2BuPomhKdRfWE0diiFM1rUwhNaPm5Q2iBv
YA8OoTxv3ItVKacGhc6iPC/1YO0CqpE0N54r/VMn0fjoTN+4BTju85MO1NWdgnhFN2bDnxOqTsMm
Cwr+MbojrKihDzU93tHt3d78t+0HyMRltRSw67heXi/+0riQk4Yo3s1JmjfApwfr6rH3rBGwZYuA
o7ODmpTS3ZbjZgtbaEWsIhnL/xouU4E+qo514KJAtXgyqtCVvVUjFoejR0V74uUZRvM2neYI5iMB
eyf9+lhJ6qG8/KdjobbpvEcpWTYrHpvqhYR3w1d52jFWAoBG6Z+K9ytcZ0h6czBddfdHWtdg4fn+
CraW59/6PfKWYyPG14nZV2YP6uepJTH0RVHvIDBp4j0mJlWatQks5SSWdD3H5GSvTrjOJ8Ooi3ww
vkt0xdBioR/f0KtHuzIxnjaNTmXI2KemqKUtiA4mXJS060Avcid5JHmq4FEStTvLOK9LWYXEUEr1
GwR+/3TeO54hCQsYX47KtkFYnfYf57copeSvgpxvS4zFuEnccqR6QdPE7tQxyyY1DeaTXV+Amj1i
A70SIbk49mOdY4LH8YvENQqrHtEvQQkI+S2nnLWHS+M3xCUm0OKdiLhDuKwoYG9sOC+G6YuFzd7P
TMNb4RofLUKxKGQRachaHV7R/smxw46iZivCHKBE419swfacauA+KjaWd8NZehdQ61W9Nw1hs2zT
4hjlEDytzidUfYRYKt9O/mAblr7YTjs9IuSZUpWIYZy4NH2ke7vKOL3UPG4ypNaNzfHyLFfEZtv6
ypLNAb9Z1/vhaCH/3EiwW9wEwI7w8zS3d9+V/s/J0ugm/s+xEE6SdmxY8oI06Me/OqHM9qsAtT+n
g8nKSZH043gp0+c2lneIURCt5njraGH/wwxDmj9SoyquyMhy71kVrTQIvsr6fEtLxpOFFmm+E0p7
nT6Hqm+8xUbVVKY50LC/iuwmDD6h4yS5VtMwMKiGB7FWV+YueLzml8ZT3yJ5VaZoZZzVc1Kt1zA0
rd1zYt70MVlDWwVUpeGUtMwX9LCnzLn0/+UGNVdknII5bNhympK+ZQcG7TI6ZFgpY+IpkeU0hgVN
5rnm8drViXSJjZZlQwSSHxWBPLbQuBQRANTiig/gVbKKCpekK63SKlL7g/KRZiStCaU1boPczwLE
KK5xD0cttooWxNWaB/pzRmrFpdiDp8mhduY+oH/BZEFXVfcGR0AnyqodrE5nV9SQFvBYY/AEcIJx
9DKil4TjFardoQX32QlPKX6EshWdmOqG0wzcM24KyqfmnA07WtkoWnaHcwBWMRZzSfaH/6mnPrwZ
UIfaXkIHtqJlMVWNwB+z2i+ynHeo3D+Kkxen6kRHYZxNUn9LgekmsmFJuTGAqzS/kpiD65mkrmj0
QndO32Vbhmk+Oxq4ijidIEArqjmNen05wAi8vvJLQ5hf5Zdgup0pvetfOyCt1HgDpmOmIRYigoo/
fBkqplJJk3/VvTCt7bbdi2X34RoeAiLbgA3Livxzb3z3LGAhDf9SCLukRahEyKJ/ZWX/zQcaHUSb
RPr/17Rl3Wj4NY8yCXStKUqvV8gpbpUWVTySXetoQaCX86TMRKOja8+nq/AOpV6GfiINwi59cg8F
FFodMcExh5N/zaIeyYJ3G2WT1ZOK1AqLjDmLKzjcGTZCWNBG9ub56oPefomA9NA+R2bdttMaK3Ti
3vGtPsBV/nfIpkeL7tT+wV1EqoPoMiCRGrzMewmzlWVzQOvVIcWiiecn+j9ajUFk2mm2L2WeowRN
FObdqZFfh3A/W6DHBcMzTv538x/7yHxNYkNQVDnfPlwKdJPjOIVGtE+XBji4A4qbdv6rrSX0Ja2z
hRzWKbg07l8+m4U1LkgSpJFqTg2TNRle7wUBuJy0alHD6lGcHWFY2XPIJ/uWBXpavIqxEAGP1glG
wPIGOmvT3xvvu8G7C+Y4w0Sq6WK9wuQo5csXxgVe2dCW9UGZ3X5Jvsd4LvOAu17AQ0WMnmjmVNXF
Kj/6OhAn0oKdpJ9qEH/KbF8Y5X+KUtw1yQonVp/5t9kvm0UUChzi+PabmvWi6QzEYKqKnxq+ub1O
1V5QOZ+5d3JBmfnhqF5/Q/RjqWYlbhv3+1avTNz+dboiG8fqi82TtlUMiRWvhViXOfwuNVMHI303
O6DSmvFXtbkrQ3Be0buGFmP5ZQ/gSCOwkTMKI1LKayazeHS0D3HX2j9hdXznr+j5emSRLHwqOELG
J1nCkE/TFyfVADvkHmsUZwUG283O1dVv8Yz77D+lLyYlA63FL6VkhQrR5n64HcOIJhlAe4ydNqdn
3HIPw/rDjhFOALOLh1rdi8IXguu6FJTGIPTblBwo/f2KGOtwBg9xwMq70RJAuJFDY1q2tkm9m8pM
o4zAwQGy3QDyhAjxP8YE5VdoCjMMCbcKZztuWVbyhJOmu016AxrKm4fc8jLe9PznTpFRS7LQe2fc
yCTut2K7eQF3ekkLzDkPQywuvRjoSwHrHMjiWtutbt0+C0LoQpVtu4fCa1fVv98/EZT9wZaFZwOS
oCzvNA8xj89aC1rAOqbL+EAoJoc1fgEONct2nxZAVC/9aMLtHGxyyks3UEUHHvY4pgGPUJqawIcA
R6FvWVa7HRYQyeZj7XCwVlXAyFtSCrk4AKb3HXW4Qkb3JK3dlAQQfkId+JhFE/ruoF8JwLfktWeP
vGUO1b1BIL+nXWkJjuLKlyUUN6mXBL6rjNlqHHrajzQiIHWbnkJDjE/QwW6eEed9tE262Z28n8aq
Gb5Ud/YRA6JrEFQStrG3D5U22gaXG4kX2FOxewY9hP6nan9Uq+gFpl1QWbFk63sBHnUB1bZMiY5r
/0CqCKif0IhOQSMscnhNgmJM1PFpKN8l4onU/6niQ0Xg9j7/w/Ilo/Hgf2HX52OHuxYnbtR7CPVH
HOtVTV5S22J7XvEeYvE3c6D+4w9EbPdS6Ibq9vAj5jLC+BUTpji0LM9a2Ra7OrEPW+k3L2KpZMCf
bqcW/OSiPrOO6/0tmSPie2CTtaq5aGnKdLpl4EP6RY/YZD+3GNc5Ge3IjrL5OPWunImXd6ZEZ136
2hw6XHZICQLBpRg+JFYlkIjckU4Q+y+QfSu4SEHtE7TLtJgtCrMgOcKKYuCo595CDFyelhV7ndQL
X/4xccyCfQZwrdjxiPtBeZp8n/0EQQP9UWLpZKtce0IybHMJiSgb5Jc243c6OmGUYTeWFdfAZLdI
QOYm6xLNg3h6qJVOMXkb3WYBpma7lFTxxBPO12sZ3qOoENXCJiXMSYVwaB4hCdfU4yripNBciq9i
3GVoeur6/NRpDVyJf74vjLKaaMSpIowRg+4stHLfg48e6Gs0XwxtyYfuNBurIOd7YE6RRbMYTkUY
0oB5p1nVgJ45VFGlZrWBXwGP0FjECmJiOVI+fU3I85uqt/r+O1hKoYAhWo0b5uczGyo41yrj2ce0
ZQnBwFF8zQjPLq1JilR7CU2/E23575278FmwmiKyVqRFFIfAGlGtGQBPUHf1hSwcZHk5utR0C/6+
H2BFHiGkrWBpVv8r/PwVERk7qfAkfciEYaKMsWzlMQJQXki66eMe+Ex+WzoRIhSLAYN6d4Kzp0jE
bpSpTCDyQnUtfQuJsgNyCHQiyUZTXFtG52AgS9AktGUqZb+oFv9TGzh1yWICGTpQkTodKqHT/3qb
WLTkLNH0eMSEzT+JNgsRJtpK5VWzsr92Mrqd4J2/RxaFxTcNiFYSys8FI7F3LLnPXt2HPiCr9XLy
GzaPONAnLFp+J3weU2t4hfJdEpPi339vtwhE/+wN+diebCADiNXs5z1uYnl8TVhJTgLg+B2aVZai
QTQMYUsrf3AZTGizfenbsBEjLQzCrecnjWA634h6AFXJtgFE0GXOOd00GP5L+3Gwr23Yw5cFrakI
nnFCk07T8cVpBLFpVi9K94MqDrgHo9En1FT9lBz/sAJkR2K9SCSPijIXpD31VSfQnLi2i5+bCM2E
XbcwAzz/H5zwJHzUBeId54cTFp0cL3G/4/cphm4Hj6EGLDR7+UBh+U3sc7kgJsvDPqaAVVcysibj
OC60+PlAysleVjVn9SvhCvWXeJB3VL+Ggr1LhJn9Vj+33eZ5jttvsH5MAHtd0pOEjRkurDHFLL5H
QJ/FxHO1V+dQ5XWlfV7pMGlfpDAz2zOUkfrZyXno6HlRXAve+aIVxMtEDAmfkwJSniM661FQGEWq
BbyOKpV6uL9KlLuapQG2+Y0+8tIqtuPLVOG3Vol9R9IjEepe2AjiTzv5s0ij3Jr5KYVlXvXkT5ec
5ZsOW/tiGmrhP9b8kjT2I3NRO0zFjG/iOHD1g61pWU4KFJBsEakQpn4I0iN9IX9AGEZCazAWilfO
EQBM7EokqwDhFlosAjIBi+QZ507biDAu9gFD6blTaGELtgrN9xmQ4wqlvwKKBiITZfTB0TFaf9Ez
+GoH6y6tBR6W7ZTvz+ZQ+srlTD9p/YNiyObFnLIW+lUGiOhh/W6u5oFei+S0Id7nUJzs+o2rXxPJ
/zOlz/NbwjpsTmt8I6A5FewE/mPr3/RXMkSwuEGZGPKcYZIWzJixKLv201ACbp/0iMiC2baPniZL
nLSPV2KnYBxMoM70e9BiZMT4+OGl7p1MydP6EJgyDXe2M/2PPGF1J0OHS06Y1yM5gIdvI0QDW0u+
Ycap2r1o9z+EPIa5uZFOFmy76hio7hMjCtnm928/NJsGsAVdu9x1HvfMm930KxlD5jDoRSDZ1+3X
gvL1r2ArYK7cQTaYqKrk4b4UxhmhjE+kjR7jxtG4Xat1Jj92qEIAhy+Dm8qQQl7CFV+dbdR6yP4o
VX348Xy74qYyzNNih9De3sPxk1UDoUBPZZizY82zgb4cBJNmUkoaKX+RUE8jc99Na7nZmXLPV3Oe
T9KXP9xTebHvIVCDwfSp+bwBeCBdsMtf655+/om+Uv0vmEsTKJT02FMp8obVER8rSzSv9qGwgILx
31WsXdpcEMDk3bKsyU2BmzLHDnkzaHGh/G6KdiSp7E4ipT9IfxHQtEPQLHrRdpgUuD5EjV+qnvl8
WhpF0cePsfbjS2V+Ozhp6bqap8qbrurshz9tBTSh4S+WtPPBjblDagHpMyTia4ecMMEVtz/QR+x+
5FK6DGdWiSUgXcFwEqR/z3tPB3Wm03a9PtJJA3Evx2gSwdxs4f2STFGONeyO3WhxmhnGUzE1Wbnp
3gbN9Ea/dOzHc3JEhYNuSc/HJIoP0sB9SjDQthStgLwABlWJSefDZmoRHdOKZyDMMUpCPCOz0PxT
uf/rDYPVsfVBKoDTnwMofqTLDlTGxf/3ps2bSrsYWgl9RNi89orkpB/MX6U6FUYzywCV+LawRhO2
M2hkdYwUTiLdV1uUa7jqp7FfFzC/ylhraog9RsNPFRAWXhmqgGSKImq7kz/hoT++onyu96EH30d2
4HXQmzU5iM534+8FZNoBJYcmpzS1V5TK8GCUqZnH3f/MFh4tVMC0VIIPwbEEAVSY+TVs+Owh2K47
OTKYZ0fuHR7H52Qf3rwwsj7AjXWg2JmyctnaZ3+CUz3iaRlpDsUWi/C/TMn3ujrRFrczZU/qPrWJ
71SLKe11sB6+y7Y1X4ec1VG58VnqC1fbmAJEyT5RXAsmmBTcnlO91TmoVzmQJencWUycwRohzmI6
99BX2pS0TxC6D/MYXyw+fPgKTXU2weWgFklvRErBNf+8MFimklJRpCGpGH0H3xNkn0d1maY9E1mI
LUx1zgly9HhIhZGFEyROkELEyvUpe/VNiGIgT/q2AnXHRTnyPfhhDE82csl6/qtY1iUQtMZK0wi7
1Dy+j2k9KNrbeJA8yVHXeA9X55tzlZkjizOH8D63SPayKaBNPA3DSy3G1HYbSmypl1EjmaSOXlZh
MqhgdrtzmSc6KvHGb7d/mqyxHHNO2z3b1uajwzYy+VJEv3kEEIRBAKq15wGHqBIOWnphmCCwSg/f
DCDcKS6Ka7HHQSBuIUfL44eIrHVLGAfZfMP8Jl81DOISiDO/FGYg922A8I6B79rxlkQSCZiaBjxj
VQs6GgsEf26KfFZ4hXyu1BcgbFGxNocaLpesLUK68eSjdSjwOe5xc2FtYeVM1GN0Ok0mC0bom50x
iRn8KPBopCFCJx2x/ruXCrM8oGpeynkbKSlncOCq9P76tPgupkUROsA6vYSIUF9wu46NR1yDVpBQ
qRJ0nxaCNeWJA7ZfhYzsUQVDXuTLJmoZquEkwPM/NS23S65wpapRaZWVPvUk/USpUeZy3Fpvx3AX
DPjPiclru7apYeFRqbbSUpSSwrJqDLwcHp6eissEDFpCIsWn5mCOhUl+lsPdWfUk6jrGY6GbDky5
kYGWwp0qTScpJn/9wKCPN6SChI1Oxg0q+k2yk7646BWlBPVDpR+n0sCluzcgKlVilm7vxNN0E8AG
qd8Y+yMWp/QJj8SF13XGnDQwJh2NrM+PEIKEf6dO/OEsTa8tTiGOn0AM85xg7d258Fb6MbqNFAHa
kofSq+rAOSyj+zMCf3zz9itbx6m8AVuqNm+UP5sP+32UMOGBQR/vuNlXJiGSPcm9EYfxVZmkHPDA
K710YOe7EkeMH5x/OeFOx03pE54OXaoH4sMK4O1pbp6GPwG6bOsDJ5Z3uUIaxmVos0qZCVyeYFXH
OD0YIDzeiSqPR3Ws+9SHMqbNw4uuQXPv4aY/QqsC6jPPedI+Vx7WPzGT7wFXwwqMA1KIHl6zTuoz
YEV4u6rC89HGoDvaMWvvyeNbufs2pI723zoPGk8DveIImqi60ayLg5p67oSaX5AK4HJrp+44ECIS
8nYcMZjwVd4bqwwd+V3/NicLk47Ffpdg9jIXRXLVKxqMfWK9BKulG2yxXT4XBzOfdm+Y5khyQZI2
TMgLrtoG2/z3S8RQ3ODHEoLuHitTPG4Zxqx0W3p2C1ld9/9JUFhsZMr6uMUmpYoZXRiaJ1UfHk6e
somqUsUuP5HagQQlwcBWgxogPpTp4eNmaLVb8CELCMt92ME+RlgptEFg6p/yqrJFeIvaoCvCI2uA
gjR5SMi+idnnK7keVb6XqVhnGWLjzn2zMycPm9+6I96ybUashb5VzFGG/LmfLp0G/W8a5XrCf928
VUhB/6tSPNfjQL7NouOlPRYJPN64wLbOTu0Ls0CzJnlxiC8BmfrfU+zVLNIAg5uzMlyDRK/xjM3z
WlbQhN5n+LGCg0X1s6mBC7eup7XIbhHdSq/W3KYfpgyD5kn8+94L/PUXRyuD5tAwTQa7liVSPJOJ
PrsSi6nG0frqF4kSa+4I+uYxyiSc+HfNkaEu2qAdxFW04LuPLt4kV58kC2aH1f26l+L7q/PMj2ke
EK5Ca1IGcXL+aw+sKguq7wLkxAf8tssrZryQpNmdXQguY07i/z5Sry8s5/HWEEYYFpjZBKO9q+1P
987a+fnvLomh8QK/CHsCCQ8QD+/pztWN0KgFIgb90z5/tlZ+RIjydvDus4MRxjnxSGpXwwHqUww1
suG3XCqWtjDwiB3PSCqujfrwRdYMMRTXcYgm0PPOpj6g4xla6i4srN1m1MoQDCJRCLZSV7PBYR/V
LALlbgY1aACkbVcykToSDJA3WPWk+wOxfwlAjU/MvMCz6RY9kr/OVwwBAfSvgIurKArEuqw1+Wbl
jEWQggUyDsfx/wz54QRiUi3uxge7dGAt7TozyoUH3LQpqIYARzTdxGjH0Lrv19/LlLhd857dOLWy
RfvbGF6FB+LxSDH7DiW5ot0KLnbT/jTsXlT0/dVFchDw3NIYEkQrq1Y30/bhO0yDkG93Owihfecw
Lg+/c/labbiu4srUZDFeVlRLfgD6/BSTtlgdOgCe3N35B4OYa0hJYyc6nuEQGeuhPFZVigD5hHQG
7yHYtgvFT6xri0/CQIAMTV7XzEzPJkWU7FZRSfgPAJbvg+4Yk1nw1k8cJZZeqWYrCOYrMd1kq/8T
DVkLnr32sztbE70h+5getXVp2h0AoSFfwP3HMp/VFCgWeJWy33Mv6ee7ahP87FOvBXKXwvP8UsRf
/KMP3e4zl4gcX2CABxq8DO0OMyisOFGQr6pnnljAhDzPvNbBBv+FCTzpaeuHWZQYp/jCw1V6VRPM
XAfDcVQoO5lPeyEKMBuskfyo2WJm0MknUBQD/Lhitxn/8ppzCqf33a4Lgnrkz8h4JHf6QDYgL7uX
nzNXAaZQMfv/THGGlxC5NRnjua7FEe2v3G+Mlugm58tM/3YE8umPXB+J5rvNUC0LXDUD5+Mm4B/C
0PJZjgAclCiBO8RjbuLyLK0kz0sNSDjc4opdHJUnI/saYR3Hp+UTOt4UqoW5EBtNZlPEqqLXERbf
rSezjE8ajj4NeJpd1SR4xx43UZqFPWSsYnqna27bHIbD3JXfOC2ukJC0YahxCuz1kUJForsNIVI6
Y0PH4lFYwWVBFKU15f5V25sRJNjwjzHjaptYEOK0NVzsPrqFcxRXm2kaInJ7olN/go9i2VUfkUrZ
GNRZycoCB1IYcPSmUQAP9s9ifxo56cEGr6sV7w8uU/1nMuZvCSwoZgRMM0kWaynMeirYw1M35zlx
SPzsW6z9+4oA/nKBVl8g7Q1wOz9vI+Fp30q5nwY8zExR8wctOv4z0wnoczmH5ym+99mjFdjR3heG
qR6IxrHZacyigfB5yA/FYw9YpaeENA1qSdvGkS+GXit08lFPf75dXdKlYQvOqEvCr92WJydv805K
Ki17fLYCEjsmqDacxlq/NfPcRQ2aG6nXmqfnulRwwdObjpFfkHJvhk/DxnkT1iHiSEF2PkEAflcb
OaGxVVWqt4jMCpjOf4Ns/sAtrJssI0S9/MEvUpUBGBxDMDERP4mUx3tPSQReUXTzkBf9sfr/uwY6
dvOWFIvejzQgtPbk2VTrGtTHE8BJBRRznKwC1+uKHMU18qBHLoX5lkrwB5cAVnNZgf6ykt46Xn9O
KyA5xcJN0pbz0yrG9R5cAMm8jzH6YckIwqQZpTrUeUNir5pgsEM51FDpfoBflACe/N7v4DW0kghh
c3sRzzMm2dP7Gmz0aVBnzCjfbhvIhnbn5M0KufbE5UTZQNQJfJk2kgPTtCQLJNHzLpP8ya2JEcTv
AxOb++USx2utRaunSdeNEDgIKFCbpP803SfQmHb4TJUN+Z9niPGcFV+ajo3DwH1DgJFHbWDOccwJ
C55I9lILFQPdu+PmupqukGhWL9ko5u+4N/drvbopyzXTnWW/KoCcIl5HsLTpuFEeOfTMgqfoaCX7
7BS/XeyW1PjPMUBKCqBEsBvg4yVRnMfRxgvfOn4utZ9cFdGUjcbiLP9JBcxzGChwu+g2hwf2kPc0
Q/zJcUht47fTWvXNxbZJLW6rAnXUnjZZA4lH+xcPSKb/NzbBODx33E6lb3ZSG9q4IE5BEAR54uGf
Tp5exgRxpviUVXrOcrOWEI540abOffzVSis18Cp/6M/L5RH3w/ef0Cs5R3QU0GGJxttcQnI2YcbL
pbL8FUw6TlTM55+UiylzhxdjR7zsZ31nCrFhpPgxRR/JYYaflkt3f9O5qfb1c+NtVDx4NzWObCYW
q1t0Eo5ljmGbDw30O+c7WPrabaSl+WAqKu/xt5MHqlyQnpy/t+s8V77AWirb7jR4rnhovqf5HJRD
YoMtNTt7nug+uiuZKQJYhKjkyviDilwmvlKCNzVEUh6RPE6gSM0V+wQhr0mlkwtknfUhJiK1kA4Q
j4pu+q6UeRjFCBJZQ/fOVSvPKf9+FRz0Pz4P8ATZoczGLJKaUkOGYipGpkgeGsJL1armtSEHXegs
C1yqOYXR5m1yAF7fkyFo7I8xyqi8if6OlHDjAUiMov1H0QDwvFqpipJRLJk8zs+mvBdQR6YodL3W
xhPoQv2BsslZRxi6vAH/0j48GzwNNQttS4x/w9jtIfAHNgpNJu4M+5TaodMgGaQVTRSdoqN3CVz5
5PliYyi7sCNRnYlEooas34qSZ8HYTZ6VT0Q66xTrj6eX9Gcg255raCvrgRXUdfPhjCff4ZMNvGS0
msqZtR/cCfNRgUrhRUXIyX8Hfjft/kYNfjXuAs8ToMK+UelL/f4jWee1r866U1PZYCIbAtTm0yWv
Cvr9+YP7LK3jeCETu6XBbX8B+14axKbK2u4iPSCIpfcuIUTxEzEoqJ4dee4wB7oB7PY+CU70VLmW
F+WFEl+8/qFa/ChJPAyUOrT5KooSSYDR8QAaeT0YM1UIe2mpVj2kgPStvJqZu9Ky3U+bl24/DbCH
S/M94qa0UauVVHuKJrAqLc9wN05nzZ0K8I8uDeZoDLTDsKIoIAwCfbji8vXrJKdgFe0jly8KEyUk
91qKvaYgiEV/qSkujK2l9sy24jmfBrArXZIypsarx49PbB8cdxYPGE/NCo3N+waAjdzSRptkw88J
wu1BxQEz65x/3BT+63rdr/LKHxZApmKkU09tCDHtNgF68rIExbGVfKUfdavSadMWtENKEsmYzKLf
Hp4IMiOWXKD93s+P5Ne7o6z9X4xf/6Wk5qu5Q96aFgGo8URuPCgamtrGujia9RJYOwLysvCBJIM7
0G4AlEw8spx0jn8wSjXlNH5WnYyu+p0ITonx8e4jJkaZ82/RhAi/kor7V9x+HXj7xQVxWd4BMBGi
MHgB5bQMkYAXndfX5SnBBoahKjpKGlGR0fZt8n7Jkhcn8tb/PQyRioxLfM3S6E8VHgFp6HyY7Eq9
Hq3921UpmtbmbDUik08/9dosHpx9Uy9nZHRkrV5bAccHuMBDOuk4ULnKv2MijiY/GqD0qAyYvaPz
VsDnNjwVcy07ups5TcUhuR2ei+AB63AlHqNI0CGP9rzKXet2Uhr781vYU1dnhahEpl+BcPTpVIq5
Q1Wau6QS3iOYUW3X8miOzecJlgY1psSgC+kz95TQfZfaalWmsCyH6g528D7I4l8VdJfCbCozNKSF
QkfkyX46Zj39RnWYtMG/vllC1oIDBJNBja7zpQZgikq8ZDzcxzRtazTcGYyYXce7G0LpxI3+A7M6
738vA6wKdP929CMnEJIBkc9Kc8pp+HQmF5PX6VewvwWtjRhZzfZLs6WMyCpSORWaEGtpiNf3j7TQ
CAaS4ZrlQyEL5nHhN+BTOuimc2nulPiuRd+yk9OaaXv3CpRUCSEbyWwtQOX/FgnOQ6NL5fkXoSkB
3ZxTVgO8yuWJ0X+C6FkeK68mBYRgHTXo4WdmHhQJc4EPCgKs0CJUAJuhSg/8j3JEoVA36/pzdjIc
yj+erRedERiNGY7BXZpos6U3wvvo5xQwjboay6/5hItTY+FmDt4dTKWO93hCCKpjttNyFadsZSRl
PT6YIwMO5hYJmicmW+cqj/CkqYz1HPzBaA6lxStmjUaacfbaG05zfqna/VUDRgtk1TzNsdGjbadH
QtCFkh5U13j/EQZRsdItPvfjfDgkQE5qkjOBfg7vwKwzNQMFT6CDahWKZ/V8d0kwNUZ9yBGLIUMC
mCWmLOq0ObfO1UUcKOFh7rDkyp008jfSEznQ603IUL782ISQ0bRb1IsZe+4icHGbSBC8PuQ25IfN
Ohags9oqFrKA2muoKJ86ENDMffF41vbvtutHXmi+1gAWOCBNR0TDJ3HcsjQFDipezlWNVLh+iraE
N9dYcXzGq03oWlptw0jBP5EO3dMgGlvqEeSrUcPhE4pohg9IEib6vHJNs9VDi/roal3Ap28d3+oW
2A3AUtJpfFWKQ/mDq6HdLjHOn2qhsUsJJl7FcvIDxvFr4NSr4AlxeJeACT/P7KbUN41ZckvlJIJT
boTrdcKu0907QlfJGt3CKK3Hxr6Sh1zZIK4dJbwSn6fmXYOFwUoUrPUFkSWK7jRhLPiAWPVHsut7
Cpl98HVJYpSLX5kd/v4beC60n8JzAHSouNk11fRSkbhNUBkAD2KIM3x2NV6kg/+iOWdVGy36Hkwy
vEjKPZKsPOjQD3Y/eBeqqU10dQdgGgzyLdyVYwVcfNCj9+VK5iI26+MAWN6ShJ4SylLC+Bh6Ge3h
aQg0dGlNoJHiUZdUhODV5nxYrd8W/9RWvaNTuraOB8qpDbH0iWqJcOxzhfG7+UijcmjPWzOVC5al
y7CilQQU4oih9kIJY5YPDhXDNGipnO/8MOvYwnouItLP5aGgKQiII+BHyy/oVGnROT8tjBNft/hb
1FuAUgkJpW/oIpzdVb2gE//1e6DlgS4gpmxLiBxX7bhrixpt2Ng1skCq0vgf5t1RPEcJqcX7t1y1
kVV1w8J7K1+N/2EYZVikyZJnpJmlnC1C3MZ1eeRku6iK9V3vOs45MBqm17HJaV7dDHW0SbA5cBFd
2Kgi+ey6s4pIywALX2Xein3K6LXFvaqmz43TxLyhf181vDj1kx9QK6+m/9BoGMbJWYcuGlrADfq+
0sUDfnJFGTO57GhEcTbvJaiNc7oxm4gROmNNJKKvEiHnw2aGELn9OXOfV6E3SVyjcAPkEMO8m0Yd
ZGjdYy03CXTjWNS1m+lRbZ3lUftozG5RV5lpop8GfKbn+CBjE4YIGg4/LzhnSq/izOFGpUx7M9J5
LN5nRRM404wZ3ObaxMCva0z5z9WHWqGblrCujuFi13ib5o+lhUrGinnvLIrJzG0JayV8R5dI75Vt
J8P2b73Um1VgWQU+v2zv/+W+HXb5aTAt1QlSwPMZZQrhaXYai1pw+fZRmpEWjmnGkd2zzYLUKCux
VYHJtj+Ga60n2LKvtaB473sbAryg7ca+efPKLZsgULf62RoPHF3Dh6lrt1UVT65qgw4X0j/5OB6h
XXRef8I0oDLepn2s4CLuQz/5/r3zwyPN1H4aoFcKRNgG7samRFF6XbO84SrMl5u4BO5o2a0PakKY
0AJBPcyJmSzT3z4cDMT4XvmCryrxJEGh17YbV5AR9G9IJJCWif8mLwgO7EM6kZAVFC/uhnBhnvZc
WPY6K0unANUcokX/Q3osBN45yjF6tIdcPvuLa7RmwB713jYUkorAgEfaFFZ12smFmPMlCuylNAk9
n/6wV6MB4rbSIfTpsiKU2eiC9AzmrQcl5ElVNUi2trIWUUH3zWbfh6DcVawcqUREm9+WjFF1RZ+o
XoXJE+mpqOe5YstmFzylTdqEKNAo2Mn2CnvZA79r5lzHjoUQ08GJ1WvqdHTFPwVl6j3qGguI26Vq
EIJSIb6ZuMwdBNwEEED0UbW/PPtxaKb7l5F+eMVHGEb/QCgcZPw6jbOZotanvC1yKlm0yYYQSl4O
CpAchJcL6PzWoCo2LEfJ5QKNm2LnwfZSRjoO1+rBzYUoJoBMnsyTBlBTNO0cQ8r30XZw/2Y2Ce4H
D2+Fjj4G2BjfBEA19NUTZeu1Yk4GhOXspstt5U3HE5SZ7bd65tKeHWLSzEF5irtD1b/650LxwmAE
jP/HuvT0LCk9BzIajX+I+cd4hwT6JnenIlyGoG9vIy0RHtDFtmz9+4YkyafqJGxHoMTOECwFlFlh
owttrYQ/UbjO2K9IFJL8gb0utHcWJ2SHlv9lA6OJJG/zg7CUiiANIoE9fpyGdVQmsTOuQ9ax1xIU
dYLTjsz/IOPAHtkMogIxaO42cLgK7xKhlB6QSaHIoOaQ6PiJaeEdWOorEaLgYmyojjiBE00p8B51
tmcX2BjsPWain3jz8IyuVBgQ6tJPt7xJ3eg86N/rIARVuKXj5BZGYcUH4PT63Uw1aF/fg6bTf0dH
F/PLL5G4yuX+phnuSLdFJySSiNcUnKuTQolFNB0ADhkF84EBFM7uJJJhq2KsbKBqn2T4PMMSP75y
Bq6yKtXjyFSRuagxXZ/jSTJPzEqgi95n8AFEEQv3/gBOz9LZ+tB+3g3nU/dodFUBlGLj1F73LgaL
MggI8LKsUflrpuGKiWhThDQ0NfhaJ4NSbr9xLureuSvryc235py0hzlp6H+3hW8eJnd7LEgu+fYg
RqiTz8gkbD/wo4qq2JpBQqo19HNby5wia9NNrJGwubwWCih1rflhlusIwDBz7x+LeEErwt5FLZXB
8xW7ZCJQx2lReKJsJJ6+NVLtZtAkNAEqLb3ebCSd8P9srR+DYGsCKoLBA+V0aLAfmc8QRp5QzkN1
DV6WM8quR2db6dmFCfVe8dPbPvRsEjnXkpr0QIsDfnLIAFTofx/c6YzTYviR5/6rnzvNp1FQpJ9T
m69T8tWtyudL9bQHU6LMFjr1UDH0Ruej3y2Hblf1JqdKkDnfDMp44kbuCcI4yi1BTIGjewzOyvrl
FQTSwseioG/9bv8LIBIlEa0dJagbrx6aPbLM2Pl2OYjzj/sGKESr9HOrbsS7TbNMGux2e9mQ7Y8/
Drzn74HxsbvJ1sh0n7EmfVwvgAoE968KA/w1lqOAmol6Q0MTJu5yulc+jbWCgUzeMozhuxEsBtIW
MtZxMEfotrIm4XLODk1RGRRskJ0hzFsGndWYLWQl0n/wwCodpX6QdcOEckDrMCdRwN2NHN2qoaAi
Mx4KjJXoKNkQu+zwwc7m7Fp/icYVGVfAz8XC/J2LUWGyErZohVE5l3i+i7CNqSDcjc2Z3GgpsEU3
HcTmONBFYaerUfGyN0ItjsRpwlq7CwvKMNLGLGgZIP52bqYtA/aCgy/3RHOsKXB0ZeZz8ebK9wdp
435co/LlKz3KdsQlnbooVcosFg0jCtmeTpjT6KulRas6v+mqQ4auqUXTjxsliUVioXnolb/p7GSB
MWzrPYxylWU0NXNrmhe9fK/ieL3kzoSjWpSgaDG4MIxLtrLD5sMvWuDC53eHQ6V9mc9ZxIELC/yE
6MPu+tYyOcwnLlE7I45xPHi7QUH43EY350DRkhXbzIAcNILjbY6vsdvmkjuDYsf888W29qyFnpyf
ZL4rYxmvA/+oeuJLBDjZlX1VWutCAqcQHrnE9q0eFpxBeelZE6mnhrlnJ9QajkYBUmZxbLK0ECzB
HwLQOpeAMGu0mCUv3G4uQ2jHfKUBI7J205jBuuppyaJNobhP530FQ5dNJ2u5Xeg24EWDreCTqZ6r
IJ76+RRB8KinRXoaY33FcT/GwHJM0AXDirr7MbOe4qf0U5qLw7YuKHBo6GZhtK00KYQgM/wEMJxU
9QgfcTii12ShgY46pGF/X1MH8V40OQKoaGxHyY5/ES1IHBxFqfoXZQJ8Atmnbxh1M6rqIoV5+Ka5
K0Th0KmZ5rqLrg8nzO2z/EKcOLxHYnS+qvrW7OKxALidCQBQjQHytL9CrVIsuq8VqPbKQtVPhOsD
kMJzaQvZ/IvPmp2oxQg/gimHkB3PcPvNX3+cutJYoAn/2HZ7pkmLWobQO6/9zZAlqBGbl2OsiXJ8
JvsreTn9mu16G70IggM9pOii0t1fYH2XxuQWp6kJydguJTRCh3fx19Z72eZwsN/7+jpQ5IpkInBT
nq2MyZnYUT5PxOSVAtmon/fY5ZllWXXKksXmebaquN7+3qBnvTVekMXzOC2OCArAUVLNUxysFmhR
GFEIuOLHz18ykLNB7SAMGtf+TP3QhV+rxm/8Fk3yefiyHd3ESs50YZoUIgEkZUYE2rAR1vbG8OZ9
I6LmXnNFzPc79CVCVxDTv3mSjZY9dopGef5s9G0hEo3zGR6odwAx5G9YuTsjL7Oae6dnLvJAR1yk
3rQdRUE5v3ej1AnH6IA5R8M04uc3Y7O9U2pWPkg1jx6fUR2rw+Q6y9+cDXPyuEW58LbMKpDrnWQ0
2Yvc2CBSPc5PXS+HohxqKb9oFd5ZyfnUkOQFJd2NmRhloe/2YkbKmrrTdttkfLv4CLXJSZf7/kDG
x11d0aW6YFzXFQWPz043XB3WU1mUsl75NKskhh/QgU4N+D9VW45Is3tWxgDrSDlwaYNrgTda1ZWv
xFTLVAgb5GZDKSTKR/Ef6cx28cZ243STjg+LOreGhi+IAsGX7vOd0kl1OKuI6nFfDEa5Hr2M9acu
cHIthyGKc0yNZZ3YZb6FcA1wNxklnLFIMEZeBpZPFfHnHOvRe4fmXlvDpvQ5TI1ltBZrG2m8cuDJ
56X/+ul4U6heNshTVX32IgUFr5fQHclnJWXjSV4gTzt1/qT6i3GTSoh7I0rng1+2d2yvrn9JCNNx
4pQCj6BAZWUFuz54svauHs1rSF9LruVwqDUGDmijM0MDTlnM5BbqPfTLj26seCCot31OFFR4UTf8
BcEwLOJs2AzMaB81FlAxMkQ2jDHwkyeNXps4i6mXulIvBX3nUNDn7YB6joV9l78++/ye+tnIDbL0
SXlCQvHXHDtaAM5x/t4/iQJ2FVuNPWCrCkG1axtCTItZi3o/Rk9jtA4jBLB+ljOXODppqLKustHm
W1kudilm67x+qLOM9nGKSOOaabexNvAG4l//TsBwoAcyA92FqQzWAgQcDXZZAdhn+Fo03P/BSkGD
J0m0m78ZzF1GS9vrW8Ug1EWMoDpU7+CXtoT3Dc1t4wkD1ZdgTbY1bkMe7oDrY0HaI1DhBrugIdMn
9E2/XxgVSGHlLinkZW8FTNxxIEoZlfnMJ8VNab9LktH94XtrpNY09JvfnmyjjtUMOif9oFXHx2qY
Qnqu1GJb6LWtrSWiqANuxITKEfWldaMxXFN5WtdQbAAU2MuxcmlarDdi9wa0x6VXN/cL4UhjAKEi
RgChApRBmt3M+Dh142w3x4A/u2OJkwVYFhcenQqgR3P1w5i6RTQB8xNgbP/XvEC9vDsGh1u54WHb
sudhD/1Af9QCgFvk6oFyv7FHI4j5H/S+ilQc/oW2KfV3JK6noJFsfsXXmYpo4oLC+El71ZsWV4XZ
sN5qoYRrhA+uOcaCnHJXhUSCDEDH1wyxavvuiub22TNxr4IQTSIhO+EloodSMb0p+dAFs+vodOiQ
D1EbyXIqRyMpco81PeK9cGIudjDcZYWgmN/L0LZ/d790HNbonn9jWJaHhTGHCVGszyajNLNbnK2Q
Bn+YNNoPXHftXKsK6QjCnCCugBaLTtKXm7sgnGkwb4Hh1MrNBPcPMiEu2ZDtKun37iBu68ZgcGVx
2V6uS7SCCa4ZzbNO8mAO35rpSavb0sbPmF1dNbv6CKBgX7xNGulc9uFJqJui/iGamFa9W62OQ3sH
pcmMY87br4YHBe2rFPrNFIInbdxkyLTjz1mfoB3BHeUNeGSbtHR6jtwtmqlQ/KtSsQR4yOVSTuor
/lTaBOP+DTSKyU5PxM+0Z19SuUKciIE7O+9G4BZb20auKrimCLq8qoSrw7web2mehka9SuqOvop4
T6RZ9RZb/4WCIRySE5zJm0em2tV7SbhDo9gzB6pQOGfRq7PaHzqUqMAeUKBD5loZyi1LINkeO2xw
gvqJEKmah+jOapO4GQp/qk6U9BB3EuVwX3b6s89j5S3dHCxHtvIsRXmUcaYTvkvTF3qYE03hmyAo
K+FsHslf0Vy5JABYPQwwTm9Jm0gv1NYDzhLMatZ2vp/mrdEEKgdplMI2x1xcoYm+szNFPQcF91n8
Rm5mNZn9mB+3ta4vt1Rrn9uZ24k6B0LlvOAeFhZiURHrOYvIxzJNqrv2CClKt0BY2gK1H7ompG6P
qw4LludBPqbZnUSLBJsVTk91fhrMMgQkeBhruQl8t4ZtGxj1amZRuS1sudqhfLzMACWmsocHFK6F
lYD/ddnY6OAhpvLE6b4rw9GlrGpARA3KM08Cuhg1YK07jiVt/h8eZ/OkiuEkOovc2b342+D28JU2
//ZnMJv0nd/hpJeHgu94UO8IM5mqLmIrbJIOtws6lj2m7xZZqv9ugEBCWSOyJ+ll1QLguhUYF5qA
uVD3Bea0MDkMYIFcdc9PaRpNAPTxxq/Y8qWC5Y57tfXxNtX3sjHZfO0nSyzcapCOIyUhp+zNDwxJ
qhml3AeBczhl7vlHjXIiNc+uP4kN1ixWESzc9CyGTKI55aQBAdPEh5veFeKVetzzlhU3n7pCpkXm
27SLJnU8T6nhhsiIb7VjrpM+u91G5u6bZ/lGorBmv1xDwwPvlW5J3101A+5Tp22WTE+sukTn22z7
k42VBypY9xaSamWqjnjhbqTQG0KS2LizQDCyaDk2h+U7/8la9IU600JGRYYdm/L9AYVp2m8lyUzH
ZIcglb26oFeo6Xu5rZSVY1j24kiXdZD2tmaCVr37NtLB++I3iPgIu+jX5QRrDZ1XaEKhr+IbsKwe
Sgk0ZwKa5vQ+NyZ4L+7mxD9rUsNPJrgSTj/gsOiaUtzzIdI32G7cm+OWhqMmiUVXK8FO9tmdUs1Y
+eNbM3TAZ3HVDPwaUNrkPOgeGjvrnhh7xhMqEXQkWnxHXhoQ4h32gUKGfIsxoTZ+b8kXxvpwimHN
O7M4DEn7bITZqNyi2I9HyvAeQB1lDGIlDVT4yKR6Gm0+8SUDl0rAr2tWtBdCbZ3oWQp6UXfPy+BU
I85W5ifsqozb/gwn8jDPMEjYpDCNnUXuXcW29TkE+vLs44a0gqlnXAL7jGsljrrsLUSZpwvADIl7
IdQLSqkTcLEq7nJNuBvL9d4ZfU+5coqKUA4eYteLxB1xKkavMwfrtFzuWs4KjsDE+wzKNnRsHQjB
WRlXo1rv6/M8S6bz602di5RP3Y3Gb5/9xL8xopskyEfTVfMqTUoQdP6zBybZFJQa8gRLNxmL8Wan
th+fAj1dZ0IKkl+eS48emXZFl+RYt3+qYEnHBf2pp71o/VQazasSCfI7MRuQf/tZ+vpG+69h4MHL
noDdwlYplytlH9T6b7CNYoEgkAXQep5Sx104JlYUL6vhCPbxdITDQ257qUqtL2OyEO9dkkf90kGG
/bnMFx9mwM/h41E0zYxvOfHJ6DqYf+eEoVlE1+DWLXCSMjWcAV3SSX2DdNw3JrYey1zjIlnrwMGe
zpAwR5qjctRwh/bUDxRH8yt1Og8A7bGsIAcPsRWHi/xSunJSfAjj66F+gAsaXOfKOEoHUs4mdwCk
R5R6vho8g0OyeR4Ovv2ECadgVduYHt0MlXOTk+1wm6fKZWuwtxTr+5bHpmgbJ/3uO+ee68wv+0pD
iAMEFsaHYoztEDgBnAvcLaEX1jmatiaJbhwYRelnwG2s4a6v5kIjVSCG20cKqrLycqjtc+I4Aw3F
ciZTppqbQfw50gZgvUcEecJX8zEFW05y/xTgly2g/y3Pj+XZdV4J05ual8A7TIJhh/4NC/Y+hRqw
kaRYPlk0F/Nt5PMxCulJ9Xl6FM1Mcwbk2Apc3m6k3oiGWJfdRUeI1I178/KuPWMo44NwoznFzcl9
T0mt//jG5e4fdRApAaSDwb7XFY3P8IHg2hf4ouesGHM23dwqB4i58hwhxNnh4eV2pb9EQ1Sqglkd
a7itnvzDtv88T0xpLw5FYdvys2m1PSt5v7CTafINNGL08lw9Q7ennJBcpMGaA9J9W701ACCB7BEl
S0LzpT2Jgf/EWUJXA0MM79O99oxtOgT+soGmeKmsRBrKN/9h/NjxnUvABlJMp2wqrD9ZsPXuWYov
Se6TZSivvOH5lygiwOpWxmBOulSO1ZF2AHMQycmIjdP7Wl+35Y9WFzFYTOkkSZICPg0Dhffw/8r2
3ia+QLXAN2hZh3qDtVvuzYCSmoH+plBk8Sox86xZe6Ladxegt7m9nRWvaacJVqLz4VbB7ytelkGY
jRP9F1G6xIM9DVJPz0V+hBClb6wD6b5aOuTtQp65lrTyNXwAsBj3RigTIZmY2hS3JjZAcNIkiYGT
3856LSNeJZXgM2cLixOVjUKFfcCQz9l6fjhHwHGRZMrFLdDMv7RrgDr3s5KjD7AbqoCpbULLEcwS
ZjXMeadTBJQfLArOlUi8+mQc1HdLEeXNoWRnUgU6cTQY8YhgU0sv1u7wsefsQGUFgjtbNcAB88I2
vcTwv3aMlRGwBcSbDk82vgmoR3PN2iZ0PqWpQIt+/TJiO0vTqzYk4quIYh8WNG6+NnAZS74IAAPI
w7WoOZITtrZuuhrziJBBkSu3RQ2oyz9GT72R7QU6vEUndi8lpUBa9/si9jrhPoyFiDMzrG/o1cDn
laMpKGZjY2rM09QP5VZl9oExYEOebO0MIzG1bixliUfxqYTybkMZqi3CVG0vtHME3OopDK5js2LT
YXam+AsBT+luNNcnaQewRimJ0ovw+tm5EbK1xmnDQBgwXo6+nIdgFSGLE2vUdWOKYrPhOWks3eFx
qWXEHjiorhvzmWJlkRFYOYXJjNEf23Jeil4VMt+D19xL1ZfVc/RbyvA+gYEN7ERXTjfRmK/ENgTT
zt0C9JS77K0QlxbfKNviCgWEJwgZK3/VjZYf+DZNRfO8+i2/ekqHKtgZeq8Bk9+mRsaAaOQt6Ge/
XBEL6tqlTioBrtrxypLgkxo6NzUHgHF0s2wRAVO4zZg86jrOr258FaeIhK0znm6WWRK6oBHB2UXG
IcZLruvHSoXqQ2Pg8de1gHTE0sjyahkqxB4uC7WygSYj9iMOAjz0ujryOpQyzuDt9yA5A/TcDHqA
KWAz2uHCU8ny2HNOCtj/JkaFj0t8tmZ2/5Fwp8fgHIiXzvvnS2IrXbQrhDV8TKPu3k6i17fI7i11
zpyK7gqTHtpSdtiRZfOHr2QmWIWabbXLhHUWaqkenoHEIHrn8+4XOIVD3Ir55L0SYIX9Er38MHnh
xpepLhB0pP/IX1yxeZT/1M4Ytttnp5b7ixeCI/GWMMO+ROrFgZGDmnc+3LzceoCBkB38TUQGRDnA
G1pU090gq5unQMsk/RGlXGmej03UNVYfNzG3sewEjuMl+Iyu1aM/ipppOTjJ05KME+uG9nRTb679
QzegMmWWHYZk4KkJQBjoihByydm8R61U+36DLtgxcKGMybc4BFIS+Nj1/SBLc0FCnxNu4s5V8oq8
s+pvgonXnQl9zZdnKTasfjgkSDUHuWf0puQZq1y6P+F/SPpYn9a996EqJTehXgq0K+yToxAPj2aW
QnFA8+z67bKmFyJ8ze2RFcswiqKJI14dK2hklFM1Rle3P6v3ClKBhdtqYUDlsBr0XEY0tBn8nLwU
yslVuHC/+izJ7p5t1Y+vXO4TfU0DVctrCfNuakslQ4lic5yh9ZooXrDE2hUg0hh7GUsRkPcugyyE
T6U4U1cQT9SwE53pVkzwXtjhih5My4dtFmCQh1IXCR3eP/1/FVjxPUjjwiB1QVs+/C9UZhnHMXTU
ivfLkINnrtw8dVckHlLoStufO8u0Ubvs3GRIZsKP1iBtaY5piu4q9maQMRTWktuDbm1RtKuYtSiW
oKkMbKeiBFvCHGwbHt9yuYfmUfiVhQDciUvUubPKxIcAx4bAG3sPnIPDInZkjVCvF/jDv6A4dktH
CYUVTmwHyqxHtqHUQuEUOXTuM5CPz/jIhtI86lRNGBGWnnbeaApLqnn+Edn9JrvZwHJMWowMR269
yZdZZ0JZwVMN7iMvGB+4vI8P9f7rWRr7gPupBi5RNUAElFMMquW9S2IMQ0oSvgdG8P/KMYZyTtxy
WC0wf7g4L+FyYLIv2nWzBJi7rcDa4N5e0tJayi3lv9dcDZ9d1koXf1HbIdqaTbjRr5KKvk4b9l/Z
SPw5eGuI58Kyajm/zWfteApV7MrCt1l7SMpQui5BiITOQ7uNGt+UkzQT3pnmAnOcZ3vrPYQBnfKO
Y6W2cnKFzddVWqgfGUc2eRq1Ymss4I74ctY5nI/Qn5+dUHpQHZCGJnGzMWAxNPGOSt8r9sZq2HNd
vrLCLtP6hsrdtBiHtgBBr62NDfNR4stFo2cScGYr87Hh0WuCJyImAXwUiai22fvRdC4e6nv2hDQS
M8kpy6dvWTNZT5cPWhs+E9m7OPcbF5LdwKD1utjl2kjllQWwp9J971ndfLDcNb+I2uLwBdUgRFZd
ftohpJpebdQdaynnxAIEPkAIxS3E27391VmODjQG3UJZavTPMdF+xqiz92X2LAu+TAap4F9SL1uH
lrsDi+iO+ypnub5Lox/sa5FgReehmexTwZYUNdg88SO7ISuhpgDlPngupJMu2ERHwksbFTUb0Hc4
u87ZdaX6bAcqrjdkxqoh067F2yh9eArdj1wW08RQNBQBD9fUOSBDji8ecMFYATboYig3xOzFvvUO
YjTYhUh8OunhKIOh1+/8Wafy4tluLrK4KMzGVZGsb2ACh2GTwfwsPBUoj3Zrp53y25l9GEvBJCc1
C9HKSI4IwdsGR3zpXErCZKtHqKPpH5pOvpL98DMNFFd9ZOrGZRHkhO6N+PtBJOzZG4sXvqEWS0Ws
10dAKGjuDst4OhThjZBnHxuJHZeaoiziF0MF7Gjb62o4P/f19V+ySFOiLODTb2sk80WL7fB35zEU
RFF2Mac/0PXTTN1LkqBROCcZA8daMAbf/Rfd1aLitXBLPEGH/1IFEltQFMZl8FoDdC54NiM1yoJ6
L8E+bDKTC71SOthcHgFz+8TWy77hjR4fIq6SUSoyum/Bmqa+cU7AKImKUNxhBIx+zR2cGeAtRGrQ
B6v5AirsVCi7xp5KPbW5UhAmWl1/4mxmtF0JBHy1wAIDzDxOCigZILEXn/CqGHxc0JDzeqRZm7cR
9cEgN5K1xz+YUYqy83k6GBuICmGcJNMS5V59j+dg2CHz0xUOmU+Hwd9/GKWetKRW4kmQo8saFtQv
zn/mIKHRiRWVWgciWtEnmtGHiXFs8jB87DujqfBc3/XkT4U3o7JS0HbT0MTdt47r+B7oAQhV4O3+
KSHcmk5ib7WzHZsq+PVfKIZbKGUt5Q3PgnNcnxg9/CjoOXTBbMi39bXgya84r+CHHpqMibYDBupS
GDZ5nEv4aSC2CqYn5xPMWsx9pyJysEuMXjV0n7nZGFzD5d1uZqYqqMslA/7Fq7rOEVAyjUuC0y7H
l/1t5p9Ga2nU80oFYM7wENrvw2hkL85eWHNRNgCOWl6tr8muF2+Dy1XjgXzAzc9H0uTMFcVr3dJ7
3vmPoqnX8dfW9qPlVcaMCkWDgZKAyDipN3/Z38yqMmH5jEiqyrK7t7qbg2eHc9CLF5FA54zi18CD
acBRYRejs9y1xIjJGfW2PDGpr8MGzGmUZB48iaBvJj3iBz50cMhNDRE4BINWYK9gnflBJEMM4koC
5mmBajYoWkvuFRDVnwheWqD9GPAg4zrB670/p5tIkgqixXT0R+agvTwKKpMj0ZxQg4Uw8ZAHGJkT
mcj1FgU/4cI7ZQGhmTax3tY38gsQxV0LgbFeTAeGfumAnuw5M6XUkZ03aPPtb8ZQCKR//LgyJ5UO
dKFolphYo2qAcs/jbZZhqMsUWeSG2lgrS14jXUUECAniEput6vQnWQPBJOjrs4sEX4l0OvZqOB1K
EyEJ3LkGTPDz7hBGNZ8SnmHoRrSBxrlrfGiuUpCFuEQl0hxm8kgW3ajxa+tZMf71K7gTNxoaoII4
odpDp7HSd+QsNSF532ap1+sVJwqMKMZWkqJOnbTXiJvzu19BzVkSVGAqAsmCxxlBrjDsFbt0YAiQ
WEkWp96TQGMGxTWk0PnlTp3zDKzN83SHvNYZHoHFKi6qkJFzPD7PAF9iFTkhx6iVFuuKDK7cGu+U
fMJ2KUNgC6uFvm/ypB4yHzrhjnALr+dKzJ4MEArxKiiaMUAEeDnIzk7oOdj+TL9WepMyu3y1KjM6
Tue2Go143IaZczlDiQR3nB6rk/jXHRP6oIwbonyBDz3EvhDe61tzaaMZvo5ALM4TsgdYh4pEZExc
dDZUUwmhMohBkULk1Lj45dq27UhL6ODMstH7lBjVHNDBP0gLgq+axdhD5ZUksc5zw5//jlVj5c57
vFgifMvQe+Oo4vzfGtfBN/oUs3tf0EW61airUe7daap/gBrNqoZAF9K1C936mRn4F2SpF8PbiN7u
vG/fty/7Ned7UrjUT+SL+Gqobv93tKD6QIS1pf2TOozC6XU0AMafbQreh9omQQ79bUlUQr4efNNA
isIjdjyav82yMxN4KLCExZ+9Yru6infRZOsm2c0/Pe6JYVw2XeJ24SpBM2E14meiCGQOWy3g0AYH
a93thn9VNj2qP2QAeAa1YaA/0uO9xAYNdgesStkvvkt2FRH9xGLZbY36XnI0Cehep/J9cMXqMy90
F+i/q5S0L6KWHfQcdCpuRvc/A0aR1q0uW5Sgeb38/9KvSNsU+6NwSoKxxlmdQ6cxVujJTg//TAov
5PPlnliXbhU2CDc++LvIhDEkAaQ5ALhryVTqQsdTMu4KLwXj6NG9zAqspJs3dZWIJyNGbNyNdnWl
dmF7EeeQl9V8oNZut40vfvmpE2jtVfnlEvvHOSu9yCDKFxT2Bkr/eEuTcr8vZ/JYg844hDn1L3Dc
kDdZLYbQeWOfFqGPqq7EyYky9Q0ulDiMFy4nwnQAa768GFy07i5ySUBYoj+2Bob5NSL1gxEFJU2l
VR3DWygBSG+0v9FAcebYjBvkHC142eMX7+5RiuDJnr0Xymu9DEi90BVFU9BNyi/afTy4wOWCtmdi
CI+QsmUX+fof0LMVVXYTy/9GD7Q2afazZiGcQUucFYRUonhGCZ+76Z8HzAA80P5oaNG0DFN1EXaM
fwjh50pKt7H5DGEVRQAmfRcW7eHtWYKupWNDNEE/rqExjR/Ha56J/IKeUBHQlg+SpkmFRyp4Vm1U
D7x05bhH5bxt+Y+Su/SkWgycoIMD41o42zisd0Qa4DWZEB4REkouVh2pnCmEZGYSXHy4RfGrQVAT
HpFlsJxWiAEHSadoklG/3+HluroLm6rKR/QR3dwthkpZDM8sWSXw8Z/clOJAMpFilTDbMR1gY9Sg
qLgEmQ3u7IoSieWa1wGZxAWO5rGPAiSWzj8rTXEVUI1tB+3Orn39bP5Qw28qmTUaK+n3CYrtY56J
4XgweADl8J02c0gnCLCwFtlzsUQByyfnV380FVuzE4GkM/+AIEZnpX0tgaoVrhAKluFCA3mlQrBA
MOU2IvWe6iJOv0mnPrXSUuuG5q8RTgM7eNSBRuy23CMkmOHUu/s9vB0G9s9vn0Q0uBru1BLqYPKK
3U7I+OQ+TuBuD3LxGnbNfVwAf9Ke5qdJL0rvQQ/nudGANA8UlRLIxVZUcZ9rhtUdl1EtBgUcpF9o
2M8OyHo0+kdkGbxQ28ze5csKt4GrMWAGhg9ee2vuUZUd/FQHKM5Y53XQaFi5BuQqlhywXxVXBVTY
PSeIVF6V3P1UzDGNT39qYCNqNqXKQqpDhgjveBqwb1AN52hGaX0+xKrWOO4SUW5uKwPBrAM5L0Vh
k3PJXqFwnTKHj+7WlF0Rs6qnA8uySCO5ApBDdE4YDYGcRvX+10bGEv1f31gUyB2PNvZvHwbTmXne
n7KJj7w61AZlXfaNfNix6t9x/tVmNlWjgTiPXHQNDqRV5ckcMHkvHswk3pQbLIl7hw8w0HKbiRZQ
GnWSWX67tgzIv5Wr8JFaFpYRMlJ2MBz8CLloA6ZEBnyC99t0YNsJBykG29aOol27ddc749vOTrS7
jdOnmoqO6XUErKd5Me6nraGW2Fy1zM9PS8ml7/Iebn2TyCnx7gSAzgBf/FiDDetsMB7kf6BoqWG5
Bs/P1xDVWTqb9s1gh7W2/bsVEXzdtmi18GeawYHklsQegQTukALIdMhyYKUBjGv+Ag/kqUkEXZgE
ilBRnWuKB3svlJc80KZosNOT7b3DmJzNj6Qe+QcSkb8TzgGMLHXOiCk0dcqAfEErbceyLEs0Ym8v
FCuVt0+42kQXVEMEuQejPATbGYAyNAwmctFxZnXJfdv0TD6X69qCybkVaTQL/2XIhKlzBxPAepL0
gzcP0/6pb5+WM9Vj5uMF0WzkEve5wsRkYIOFCakB2P0K9wQvIdB4O+UTCrgXORxpNPXPMUVQ7QXQ
I0+3jEre0xkkRUf56cGYVishQupj2EvPa6ypGcAf+UaW13pSEG5rZ3xa8aBXAI4PrZ2faifGcIXR
odgIZBxb56xixH/TZlUwnDFrgPa+I+OG2edPrSv89+az//tfRtWPv2UPev+8RiC0bxPF57HHqX7p
3TYcUtq9bzccylJq1TP3oqtYvqhnfoEERMSYnG7UFPwdhhM6iZg72U/YAtGo9JSI9wewYvc7ssPo
H3oWZQV1eifKc4Ww5LuhFlczXvIevezRud+2kUcteW3s/2bXN+VtXyFRUFOkpZiKVJiFt2pa/H35
uNBR9dPFNk/Jt//xS0azUZ9tDNq5nOseJZoVj51OBNv2LTBNbZPUl0EO4sHJ9H6su6X+6hRWANtd
UCOnBnBw+I/sJReLJkqaF0bXNNdSB4zhBhtBgRRlldd6bmP0dYinvjEK7sIaTS8DJND8ddSuxmze
0jYXQmhmR3Z1UJmNRbExWrxWX+dNda5m+v1R2vGnAy8yTQLbOHXpP4ZIUB1pTBXDEP7ATqYbdpmN
hC6hjaUsBgiuzb7mBaPOgAv22hGl5ZCI5x7RsQLYVbG3lOB13yg8Dn4Rca0c+i9PWVUCK0PDjVh7
nvgwLHU7wbSMLo+RBDmayqJEwi4Wd+X5iRy6wI6G7cZZbXVZXCVaNSjwb85LpqEJO6xXAsF5t+Ug
AWn2e2J73S/SMslMGh2YJ+z/0FMDX5C56XUCa3LfhmkE8Fpl7a30Qz583mzqCKLTqWBW+CqsM1ZV
cRYC7nvHX1O44HOxR73BsJJuL+pqIelibppNUks07ezoxC0fzhy8Ipe9dnCcQnMtOfD034Ol3T8q
5zY8SL4OQ8Y8laRHy3GB+AglIsejLLyjdR39fpXadMhK0FcL/E9CNCfO4OwXycxDwwe0vhML+wn1
ZESFTWmqr982FE3aGy6xizDPQ4xoGK1LmtcVAR2aDgtPxh7hbbn/lQBXguE6Ol67zpBQjTIi4oxs
Wt+8hakCueSDBfKEGylp8Y6K/cwv1Z20WWd9wBRt10vkkL+15/lOS+U5YePE5O4X8QtJw2pG2VW1
cqglBeZg1Ylo5FBzz5Z+LHmW6FpTMaEIfbVZye99zobUU/aRZ1Ad3CBGfLRNv+NVehGh08uSK/Dr
y3MJLGn1sD3dmtaehsE2QUQoevWwJhJP8AJsGXCE7cHgK3uj4pcychbTwNMgGdohpU943pOwP76L
ZOFHRYinywKrK0Z6PcRGaJSwY4ijsY5Iqdf2SL3Qnn3Dp+NSHJLYhDwBvDWHfogCdJhY1mU5hVwz
gQJT9PQEeW6H8N+HEAgJJmYBjHdI0TWJE068Tj8KnL7rJNrmoTUinnYj43JnX5UlFPt3bnINlEOy
bGQKPZxmMq2Cn6lvmHsRucWtftqAOrS50rTj15Zp4tWB4CO7GzVxgsxaEyhRqhWaPZcXhDJdlzWs
VFcKTaPkBCvrPpIDlLmEAD7yyDdYMUTtdTV6K0e0+2d7rZLHbb8pAIKzS+d1vGRQlwSbIdyZx1qu
weSZFF/wXrGQ5eWs3HNyXtC8/LNq3BuQ37X31IhZ8uap2gCSUD6W0EUxatmn+aEuybzGpnPKeTyI
9jXUuVFWRSQDA7QqpA72LtriNA3Ira9xPA3LKwGHaazQXL7C+Idf+cOQO2y6LoH1oJB+bZZ5CV31
BuG/c6lJmOyIRiiMhjO/+qnYQaRaxGPc3fJCf6tSnwqyCGc/O/WZEFLaOD9Ow8ptnulxDGM3sxwe
OhKjIkGCvXR0UG35q0is2XxkqVjC/jKL3ac/3BT+8hb8uQ7R+oQGA0OiCjyAgkBCY8SqVXbCK/by
XIBcYuYYYG3ydi8piC9mY19N2UeM9r3QH2qaJWdbNTipnOB+UxFoof3WIRuUAsFcixCno//ss+Oe
AopzL5JSpIbknlTpZvDHayf4OubxCywaEQfYDWyZbv1DaqsPmazHPPLB49Lbz5fCUuEd7xmxYA0s
/0lUnTAAmb9TQnut315QNa6dkEZRhePqDTGUl5NndhDaIRv7JNYfG4QNdZFaiF0tgleebC0Esyq4
XAyeVRjRdA21XPspIMXNbOG2nmVlYwxyTlhQqSZPDrLfkx1bBtfgPx7xOYjJJug8XqxjQ0ZaoMED
+cyhKxIooboAtrBYV4rqmFZnyyCuPGN0vjV52fWYMcrZkVV5yZOSpK4LimhSxmSPhCnlipWZAg4k
Ml6Z5Ow0og4rxP8cZJ1EZRueUxHtnigcdm+9rwojAl8QT8mtvSxgeB909Hn4tWsmGYaqWNpBT+Tx
WwAbmWy80U8ivnkZYr3o4NxpxUK9yq4xwOX2WQHomrIStpdyBcMFKTtPx2FObrxOh/EJhDAzQCL9
HvYJeVPiPQEuatun75OthtTrbDPIb5uIESH8vDS8zR3wfYw2XCHvJxuUCRWqjL6++6xsxvDzfi/a
ss/9sATNXS2I53JM9mgalQgi/Ud36rQm0kyurVUWpVc01mSg1vHsDcOk8G87lo2ANrI5G+wyvA+Z
AbjykjGCQ9DZoEk6tQBwiUL0iIePKqvsMlmCxDwTkETN8s+Ua9QUKOy9jQ1xC0vFnkYCfxtefPEO
fVqGC5oXJSGz2sKudaDaQ72Dn5TqnQFXpUnBr0gM4de4/DCWOzkkwahwgZ4QmJi7/RL+mCWEUFZ0
+u+vgavO/Y129erXlbKJJYYl1L4VObDOeOMODzgqvq+ZXFnaYgAZqO/qCLd2o4ztiTFnQ14+FUCI
6Jv1Oi/NbrDYfoxLz+5a6B2jjeHblwbFrmpJbbrlIWGATosPKPlXpTmIKn0H3sP05er7MvRFFsaB
AC8nITHVM/AeA+PVWmPoXVPEpzSGeDd7aoQRln9BQu/yMLMdO29r12KB3XuCXhx3fyxCohUce9hA
B6eoa3ndnOwtPb69YaiVj2CWtoddEM6MfhFt0/hX4rYhrg0BHeXSdasGffTpnp+8tfh7O6XFOgwz
DeARbnNGVEWruhj8uTi5hHPGvsFgyxKyLVBgA1pMle4pAu6ZXhJVd/tkbl69oF5sL+O4jCTWH7Kq
sT8deFvyeyTB9Mb631DB7mcA1j5oqwbGcuZ05V+AHe1Zu0gAjCNhzy6i84Ko8Px64tSdbnChS1f+
dzRrkEnnL/JgZspXtaBRrRg70W5yJ8lbhD6jIO8hh/A5uzMhKfDaYaQZRgQnj1NOecwgllF1MDvP
za4XBeNxcGmn7CwxNNtYdc75ba75PT3ndECHovr23wYGZZDurV2+pYbgx33oouqLkf8enSPHK+tR
JcF8BDcqnOk5QsSRLyHYVWV7pjnDKZqrU22iOlK5qZ1MR1EZG0BwjYc7Aa9E+fScoQpvk2/mApQA
Nw9hVxkzU8eplcHHtdDHrCC4eMijkQ03i54JPlsS1XJt+116bDuDxHISQqA2Btx9vzi+7u+tVBTB
vryy6b2KX4nReP5hfAKBE1bCB6JGbDUlR9ASGXexqK5IcLCI/eIy+8eepMFd14PmCRlnS0M5IZha
W/WyM47yDtmmIAybt9ikD/LQPfB6wFWqr88Daab/3hSrYxa+4GmYuVbd1T86L4jBi9xgf+K6UNZS
ipEpEQHdCMCnGmh7Gmok4owuirbJaQfM6huDXhNaqRXa4eHnPMsXbtmAUeN+Ex/N6UO+/HXKslXi
dgRzGbOnZWvBTy4BK/2iMCifhfQzQw525NqMJ/GdL+nnyqVEb2JWVYmnHL2wZQHDY9Y1yxFDTpJR
jrkXZlpXuGhue8VSmEbfc5hfqkXUyZlzAO+lDLwI+FeNpZOqgwG0ku+H81LxvjWhcrsm8RI6irp9
7vrgpKMmUKY1PuTznP/trjEoPZp5cZ64hJ+y1yKnW6IrNY0XPYsxmuzwQTAi8FtHO/PZWxa7Uqnw
FUtF+oKEZbTktu4j9Xn1YyDTUIvoHPUM3FkNTeb9SKWPe2wC0yEYcRuhAOKKvnnkQy+sewuI58mB
8/W+sqiHVcP1qs3Qzui4lUjIbli8wA3FST7tHiPjeDPLds/G4i6KOjL+REHTUrV9m19R3QuSiX75
v1apuzJPZFdv7QKnHs7SpuJhyi8DNBmhI0D4hleJyxz9ZifXoklLOtu66DWaAiGsrMQpLp2cZpLj
3fOpoegC6iByBKi6oItXxoqwzOMz7S3hw97GZqajbhdRMMrd/9PjSyvxve1TiHZ3vcVxb4VvDX1D
tj+IGsdvauRzl7A+GSTYzT0x5Voy1U96wA43gnFLU6Nn9ja0v445uVkstACr8WZiLeGWnvYGSJXz
zbGMQJrxKCxSzMZLve1215a+v/YxXA8q937N1mWdSYkGQJmqQOPgzURGGTT+cCVbRVrbSUkvmaGw
IEmt81mtpNNxk7b+LY8K+Z6h1dR2MxdBSXBIOF8FXb58rVMLTHKzbRTmCNxmlTv5GDQHhJ0uobD9
atgqAhWQBkPHYJZHEvm8PY/vl5D6YlWVZyhc+yFIZ+5VQhFw8Cs0XN46jOnw3XenEXDehLFpOnPR
Q6prHYhWA9oROLVhmQJkS1DR2bH1oIWG8LAwmS3NKBiY3QN5t9iKmqIk+/yMqo2pexr7fhRrBiSc
d/RRqz+TeVww+1Q2taMTV0lCrcs+jCQw7hQyHDzaPg/wGJj8DFtEPhU1rGA3HNd21OEm8SGDqIGI
LW6qK+GHMNVdSxGceCVW/eqAEtJk2u4a9anJ0Om5FBdEFPAVlFVxla4/Hp29b/hb4CeNS9pMrE6/
RYJhq+5y2nOW/xg0jkkWg2GaLtrVIEm1h+vZ7JanoYE3TJEH/rj7hAzt3ZusqzLiz4mh59WaWMsk
uyFQ5wVBbQRxBWJxhUC2HtNFZ7s+5ir/jiCwTAnR+MxjEgRVZu/7hXKfUcxZ5pZYAgAxo7TdttFl
xfE+2a1a3Od6JR/JALnv/Qa1eP61gSkdnW9PxAxViZi/mQY9W8ZjdbwQAGBcWShNpNOUyPL3hpo6
jM5tVeQm1cC7wnGd3YUdTtLw6K4w86w9hsbK3j2H8y4EEK+hqelZu/Nwd6gkUEt8c+kGDOv5Y7+h
41XJFNZx8sNScE3jRY5l3Ci1zPwClcpZNiSoloisxd9+U97V9SD4M2mO/utqfDkvPxwBQdV/Gfqr
YwdZRyheN//2Hn9ZtXS5+VJTAmGPZCu+bDiXxT7jvTTOtl51gWvSzoAijhvnyGnQLA3US32h6kHz
vzAA7m9VrDFr1mzA3HcPVRkaSpsmt65ndFuhbPWpwJ+yfGZvAWC+5628n8BHfftI9KCm0FrQp7ra
wnem9ufGKIvQ9R6WSCVCBUO+Ujykw7HT86JcgP61Y0dRTX3gEzwJgKSsauhXAyv5q8d93cjyASre
sV63rvI3HRXCrjlCeGkHNHtTlTCUyuAV+Afa8+uBOCXKZP6EtJ6TXNUy1pllMMxU2+qncf3N4yYy
p4gdCqGolR8zeTUIzqb42n9ebL9F+CrMfQWVEcLDHs5rI7iT4T/53BicMTUMNamdH2qyy2GP7rBQ
aR84U3J2C/OSb6jCHa/MT0JtNN+RfjlCo6dSnyBQ2vmmvexYE7X59gJ3fUz9WiNhT39S8k4dkQXO
y6od0nK3xHQqt7Bxfn9T8tcS5L1BTZ45ItgIteLjtyaxjXZgfYotKa+6aPKukU/9N6M/w1FkHgOr
EW53xlftL38/3+R/bCzEQcm6RDzP6l7YdoJa+J5z9aX9+IcdB8abfEzsUhcI0tx8TaWMrbBxWRJb
swcCn0/YzzFHPDrIxxTegRENxs6LS2Y7SS13Nj51f9B040ExpByvD1B0XZ0i0Dmdp1wAn8G0fmwE
V0ghSCaxMmz6Dze2a7UtYCa9MJy9qlRZmH6SR1usYLgEuTLtVq0JLGVMd2Z2JxsvLagQ8pT+M2IO
z7IbjEBxzRHjWB3CpvoTuaPZmVRLedbPK1GPszrIPClX5hEhb2zdumZ9jMITR9gpX6bz2kJ1jTZS
wSF9vP2IrxipX9n4m6sz/lpX1TI/cwlAFCuaEzi9rmWwVtRdo6hjmdO2ZPSOm0DUIZh7kMLD5DM7
u3Eq/KrDEEnFE5vjlHl/HM/Z4rS+xmNtQVOI1nIwiOZOYaFGtMejxTM43fjCCNw4yCgAPwiHYPad
7qW0oGhGhIOyalDaZuECB1Ytv54XN9ARX9Wa1BHOAVpvDa4KV+AMhHUSoclDdCURWOW8KQb1Gyw6
m80/Df0+I/50Y/Tg/WMWennqntAVanU5+b3nJlHUKadbi+t0i8NChPynTZCxnvTI7213UGeiEaxn
IqagVadFlyMYpfsO1tQTuCk92GhMNHovWomkkzY6SZR5SOf+2hhnvbO+6AXiezvelJNUQPX/F/MV
3svFy549dpTfK96oQTI//KQePuoxCrfAgcQJwVtD+XRO+jNH4mjCa1vOus8Hfj+GeI7bcQP2Lyvq
3BKIIxqg558ZxG6HHb1OtlWnH+qfPIYx/K0hYL2ojY/t1FkXWsBkHl7w1tG413NV7AfDKEPmxgHW
qim67PG3crZbcIWacSYBLoVL2y48tOE30Mc6ojjguk4TQwvCQkMAOPPk4GFkAavp4Q+urHhYPJec
BE6CVM7DQgrvnHoNmc4y85ZOG3LOmJA5gb4Ta3y2yck+ziKIr93mVW74xStPQi9rlJIqikHv/7df
QKRm/1Gt+zHOY18Bxc8k1gJyyjw1Qf59z8m+MtSk5ovjbLkeDG1hK0XEjy+cVixYqhqZyxe8lFKp
BW62ckYOn+D7/sgj0XKB5/uwyqfm/3tcU4s56J4gWWGWW/Kd6tu8NKEq73Smg+1QlMh7u4lvmPVC
s9mN/U+Xvef+MT4bE0Z1V+yt7IIZ3wQl+J2rYBxCI0SGslUls+OjPDWc+XUCSlj/id2FSPzPqTpD
0aJ4nY8SQh8K4tfNJ28W7A81/yUD1wCptj7DRd+tICS0aBI7yKe/pyZvfw9XH6ukhvAnMlMDnAXJ
+TnsayFn7qUfVkt8n3OqkOTXP6HAmW3wiqqqI6KheQiQWkhWx/yCvuDkh0DKkvx3bwmXtu4Zdy85
0mGPwhvFatNrCT3lP6Qc1O+okopfuevLxJn3uuwiu50GqTeuWZqANy1ePEjK6opyDf6hPF0FeP9V
c6AiRbPMi0B6HOrS0k933EUjbuk2dXZnJUX6qpK3FuvK6nCIRGFX7P7nsqi9OT2YxEjFUrftXQ2l
w1n3OO+nm5luaZ4vDAZGODxsUI1oCbBy/eAJbkDtMsMqWCEHD/haRP3BAs19Buimb/TnorqY6jZK
sKOMXihaAk5YdlF0hvDl7qP7ur6C30it0OLNIkQBxg3UEA3V1fnBqSrfJA1+fSn3dZRhtmcsY1Ue
9gXt9l923C7ieco9YngrsxjvxFVU+w/XDknJdyM7sYlXA07UondZvXJfkj1mNWKSgRx9Q3ZreuN1
OTbwsplsQ8mHdKnMHBhZG09OdWvLJKbZtjt+m/qO2ZX8u9QjmcGn2IopWmcyOGzko0q7sAfMJfNx
DnaVn7gqUjYG9rNPn+JUfXrMpRrv8OmqiHJskuchdm2uqnqK07GnmVKJ1nY/rEWyTOfTIrgPNBgx
G3Rm0bSaJdnrvanK3B6SF8eVf6t/Tgi9bUfRsmnmtJy7U6tc7Hsvbu2Lj8wgrzhluztIo1uMa5zm
WPOc72ncWhLpg2y+0I6BN02K+pGea7/Q4L4tnJRQDPrf9lkl723CQH6tIuDTa01O7HWf+WzHY4pK
ubYoB4fMJ8t7ktV0VtJheaXLSlPQPg70kfPEMDHh8aQRL2BS+IblcVJedK3GgNPPM+oeQ0fNUcsQ
erChrw6wm9WQGrK6I+NWulDKOYSwJxaIei4eyGVTDy3/mwaPP1BxzPyXxGuzBpoHPNzmbcrAquAE
FvenkAQhbILAEiTaIdVip9fuCX8QptSnv816a70CbIMlCa/1WBjCDlS37IymKI6tyX0r89iVwpXT
L22e9kNHTYB2lCrZlGVZtXUq9ZQmjqI5d1rUmLt/tUd0BYU1cASLiOuiDuLTObR4hMm/0jfGJRQD
PoKFYpIeHvRjLnCD5rQ+g6gZBU909g8G3TqkRbAJsMWbf2xDSnsHWHNFPYJhfC4algzzoP4ddBNc
Kin1MA6MeScHl1wMS7elWGVjPgedsKyU5lDo9t5Ai4LmJYyX1OHFOebLgWCW/80vmYFl/h/VdAky
iDrsYhj0EoBFCa0zqvb7Mm/QCQdiRecllTORLQu3/+zfrA9jNWVxIhc9FHUgZm86+QGQkQOxxTyt
MlvQ3OXMCj1YNzqbcIgiigJG6NFvkbdHdm8eFM+SKdHf6IP3PPTLKPZW7olRCBm11JpjrgFBCmA5
kUdNa5NY9CNEc6pPqi7PYuXvyp1cbOfBoo8G+NnFzVur/xmMaXnkilbqyI07VHhIlqm068bOtfhj
XOUTbmPGkMG7UwIFoqVa/Eg9FRdjWqPgHo4g9XPFFgCtAU/W52zHtmfdfzlXn7qe5J5sdJpL3nX+
9nB4rgmzTTake9nKy3u+i4jV9L22I/Ky6rJt78s19xJP3MqbXfMEchajhvPBSBvMmP9XZVs4fmui
i6rm4pjyplL2YK15D2zr5o4qiRFYL97tMbLJ/sMgvopzYRv8QJXKIGL5zYCQIfjFaevmFTTQT/w+
O61cPKAZVw8TixdrSWhiBrNNXLWdtK9ayY+4C9ZCHD9WhA9G3KV+br3diJCSi37tFqgn1D1wvrMw
JhVHBG+tLCi6hbTK0KRy2BiQb7hBJKMGGt8gft8SXkeLzvmJPtIv28IQjLT8wKljvcOwncnXsoH9
LGjZlim07AmQu5sYjC3RAmm4YXNc6EiTfOVGSlg3pSVKFj892r4xafCk0RusuviHHHRUJT+uQg1n
HrKUck7jJmsN/A29UWw4E9wZRAEifu1pMABdOaOqd/bw+jDzdyEJdFk6c8DAavBpuZHQx3qzuzch
CdYi3/ecszGQMyuCk7/BI13xJJVvQ4o5UCIZq7rtl8n4hXDEv2DN1CEuiBJqWNlMn6bFa5BbXGdA
7c5Eafwam2BYWtoC40vHNpuXits+mafYGPblQw5iLWTbXy1uwfB7rFbjT9CuMaoJh1kVLdNlvlxV
o4YKPa71z9+YCpXcN60cmWKj6Lke/VXGEbDnm6NYM9791I9nCrVkj7IggBsik1McHRMP2fko6W6r
X72Nse7Y/QVq+acEIpzsmhFuoCy3vbPqO3sT0/PDeqrogMZQUdQUN5LpOUAlIjCJWj2ziy6oy2Vg
TDbQuxJ9DZvGrALCjM6m5EWjAZsPr8Et4tcUwLXKVSZN7kdkcdsZhhvSBNRAfkl6zusOwffdycF6
Am32CNzvK17fi3aMJ7wga0UsE8ON6Vd1M4EbzbYo5ShN2NFa6j6hROhmCA00uZoIRQ4116tcJDcP
DPZjU7c3y3woYqGEvQIQ5KGQDbkyYsMSv35nMl2h/TtYZIDACluVCE8/oo07hanJVc8Bjv0dlk6+
T2jwmJ8ccGcEHGsH3HTIQiDefnSqyr9Fu6UkhmwxFaZsqVnZ/yWm4XrmFcWvbH0EphfFUTzWDBhf
8w4Ml6gstrghlITPmtRBG0rcoAhpTfCcnERUd47LKYtpEp5aoymF/QaH32/VqKTW13MMgdl6JQgs
TEbUtOh5x1yfUIXZFHYMLBym8ABdi6Eek0yiHuNsLtjLcgD3PpVhQqHzGph3Fnhzkz2YdE1buLrZ
jLPdMFi7oSNRA+9AG2yPYp+FkTugX/7gGXrWl/1cZYdbyQrq89fzzlUrbWUb0q21SsT7yurdYvJa
b7QgpAFmzF5z+TfblaDq4nmQWb3T+yeYMrgThoyj2qbicIqcKjhmYH8vMHun9r/MXStBhL9uLdqR
KGEpajyfXgJU96yya+iw8KvPlzR8qjRSsd3KCI7SN0VCApJZOG+18lOWGnLCyA3cJ7AIdYu+flGz
HT+9qwMS45C1iJhT49N2IQNAczMmR4nNvwsLiiyl/JGWBtVmR269SMl6C1cKmfDOBbS1/NtmY8RB
F+O6R+I+TCZCkC+yebNAEVLB44J4LL4fo9u5EgSy4idvt0ShdN/2KO5l16MSiUIRnfsD0qQggkJz
sw9ff7Ak4+ctLm4+OIAQOv3G9+TIqTdZTPPZ75udtMNDEKF6OYvwW4ynD/1DJzf8GRrnltZW8YzJ
dAphentWw3S7gSE/lSNdDmb7Bp3+sUx95mjQiyl7S5DM2TacCSREfUHahqASkhQtm6Iq+J86tkCH
M1QR8atFUzuszs2VahiyIGalAxXmsRlRnkNsKo8tVu9I/IzQZin8AWZYXqmp5whm6elzjWtXS5/F
Y6+61hqZMoh8mVEdMsICV7HCI0R/xP0dYVMOl2LbzrmMuTdXF+fCk8wzEMRPNhg6l6twZx23fB1G
cVclde22hk/GC0GCbdB5lNMgWX3Nk+dqclGCsBjZ9sbmkgHmN9TKVQq1YBMRCBwk9VhycFZAn3M4
A3A/Uk5kXu9gTxMbiBSG18XgsNsdaxy2LGer7ZFs0QATfbrB3eVNtCmhT+wza+XgGEK4hiWYLLOP
mcuqv+IiplL8wDHiorxvj4f4BphR+U3N+JKRCCQXkZQndf/6ni7YXc2VxpRjOgh4txlEGh0Q48IQ
YgdEadHs2cD7bPtod83Ou6EjwpR7af5CjNASoskuVx8Xz1AFIAeJW0z7UhU97nyH/AX4dmEFdnKy
EOPfy2vbHIz1mM5ULeMUJIm8n9n8gzMbZYEwCIEu/xFIWmweUitu5IU3djdUncOO62E23wDGy9qt
n5kyF5dNrtLfZ8xff+hvFbK1EV71/xhfet106GkkbYh5blzynYRyH/hBjsv7AFLCbLpURg25tAjo
ko8qZVxy4NNwT980lwWjoasB11J/cUiN+Rt4l8UZckGMDKzVxSvHbjNMNLMLvimTPTzZSP+C/Nmo
9Y9M76GubPVu4UlaAiklCZE0xTWtb77K57qqRBpp1EOlhdz2rzynDeCbUVG2RzB0N/LYqJ7jc105
G3eqWvndNQcdPkPf6XFuTDynpLDqN68NcbiXhFXQAplvZd4Qp4m/9CcqFmENH88YxM6Ja6Z/20z2
DkIGyo/OGjCiG9VMBp0/5v5yzEL/qOdyWJAskXJGoDuC8qHZlR6IJAvwG16CiyMEwE/n7pkxVNYt
3xouu56xcKNxdsoINgKHqqmZjxDDmmKVr+IwQvlASBaiHOthD9P7ZvrBfzy/3RRTS1IyJ9JSKjZT
GocgzMfxTPFslumWORirI7kl6gSzCGLOKZH7KOnUeJDVEznP1vHHv00fNNU/xvQfLUldHM/uPFN3
LdCvzgGbREHYm9btvpQMYMCv0FBLH5pDUoo2G9CNNcur9oauqwHnOkn+oV52nqi5hrApDAxyTKxW
K2GddpDwGe3WheUvSM4fFwkSVsKhAoh19KjDZN2XynYbWKtU7gtE32YOyDdCGxL+xeYmyCRPndvI
8jfQiVi2yhu8jYu6/kE0GOh3XQbFSKu59h/h0O+BkK41yksGFEiS7Y0WPhCJlsVK4ElDD3E5soip
mBzSfRAT9w1QTVT9vY/z6H1rS+LvAK142xm/8q/w+uo5zHw57NyIByBvekN16h1MV16DRqSQsQVY
9Sj/zEYNMtQ02gBgROjq1/f3X82rdZ6pw0ivTtoIbDxVES/nanKLOzfc0nlWovDKMmZB0vPQIjXa
4qtKkjIp1Ijim8M0OWqNbcvFPQ2ivKwMBHO8ANvTARX9aLBYbAT2HGNUT7kCKC5sd406akoQ4Cn6
prQUhZs6WIUC+/Q+d0LnPlvxybKF8LJUaw9d/H6jDk+QCbx0BOrrznYLIux/+lx2Vn0Du7oPtqM9
rywr4QBLRZdOtGNHdu9lTaF1I8UfDP2a7XIbhs+U2DmPnYz/EGi1UEpgbVhLp0ROCb5Npd+mT2eQ
jCw3/0KW7sFLD3ajPvpBbLa+Dgl9fK6EfP8kT9oG+6hvfZt1T0dq2eg0f3tXhJ4G3mXhF1NuZT2A
0IAn+cmR8iYAIUME8TQG6JcytaqRofNdmjZZeImJUnsS1h7UANaTFD+QYI4wdO/QWvJvZwAarkFw
Po5fEGt/5WKwFjE20zg6QCLBW+76JSdnDfLRal9k/A5Pa74bT2HIEvgDYzNpeOMEgN6/PwDjKzGI
dTIx7SFh2Ta0SwjJ/LANk4Od1/YtjmN1edqYeOzpmNdFrV4LD0iAt5Yis732rRLk4s+sawd0GOCU
/4zCvcyh/OIUX1Oi/zMPZdhu/Y72pNosqvPayWY2Fik9OjhJKcbZxkKm04UMA1/9yIge5L2vVPUL
k6TERI/TAeYM7w3bbEHF598RfCwvG8gHJpCY4eaRB6XxPRIxaVZ2U0QyQoEbI/OzfS6eVSoaGFXb
9wsCYptLowhbSonKOBvm6ZuUWgKi/hyV5T/pffwYRWYl4Eo9Wx+Lo0ajZFVrqCN6kZysRcGRiQR0
3mfDzl0wBdj5uPKcSjoiQ6WxevDSBX/GJN6RjdejWX2dsqJGPVHno8MWlAtwwHEZu+MLY10GUEPh
gDYjnJnUlIqSNWUIzr9NGY5wCaXcCiPYwT7lccEa8DskWABuONfBw2EAEkGLDHA1xoLskfC0t4Nb
tomLdGMvUgq6uqM/Zy1lgf6XIlKpmS0TBI0Ii5P2NNUz+1Fg4m+EL6bF5BfVOf2h66CdADHC4Dp/
LPUH03l6DZpVMYORcMp1zfD809c5ZCwvANOT/w6/KBxN0Q3iH4MTYTV+Vp/Ym+guUf9kFHipXPrU
0h6KUFTEbzKqTKwMYE1lZcTERFowIRw6+Ez6mwQtJoWKGJ/vp4/5m8cfZP4HLtWfEUUc6nzHijTI
qAnri/Z7Cdc/C3Qe9CbT4+yU2KGJBi425GreRDXMaCPlXXsdxCsVOxcQzQx0BGG69ha/9Wrm1Vh5
AI0apKkPh+k6tvrifQt6esDvPrM/1vVtxo6bfecVth9UKcaZYdes7WOhIYxTwIKMMc/bP8clGC0s
WeUe3laXlItQUWHbuaaT5JgFf32Uvx/ZMiUzMlwkOai9nkPBPFh9dfan8+jWEAfgm7tmc27jtXwN
4yAHcAnGGrwV0t61EHOfGJhrTyI6j0WTAvMtgRP59q5NM/BUzEIqkLAildsR1pnSw+F3PHwPxTT6
toiPsJCaoLvwRuG3cKeyLkClHlCfBHt0DcEY6xdgkLgWaE0oFC5UPtuOM9We2aleHLz96mH/KVgn
Wiiw68WbYH9lr+urY7IAOVXon2tZWZIS6YuVVgypxIiVOZMXKIuTcZgdi8FA5zlz6s+Xpgi1NbAn
RaCVh5J3n6YzEODnpYUZjKCEFlbqL00Vy9uPJUgoLteB9tHdrFZAPqhiQP/fcIIzjegzM/0PTqBs
DEs32MUhpEiiDNakFomoJsTtoCjRntx8rdNavZAlDz6TcQFOYKh73H95jVylRPKUptoRWI1R/rMa
JmPG0TJr++uoI5/juP4N96qOGbQzBu8evDEV72MohsBha9yrc6D/AeXFDkJ5RfjZbQunwxJLGBFm
6i0It9m6p7koq+w2bvp4cwRzn9ret/rUr/pCp7fyNkqWlSTWrx5lGJYjCtCI+35sAEq9h0TTHenn
jVnmJIDSpSKztWgoiyDPM4RrRRgzw17OKr3K+5u3NfPrkLN3pDQY6vXp7SaCtcSphPMCpBdbYZeA
3VgjrZy7vCsryuMEqLSdgokz7Flygpv2St+88JK+aI+cc+JI4AxiOAEUqDIRNWG+8fvHPPuZ4/JL
K5NuCHH3aSRledVl0DseYjostSPqE4KP1r7UkLoj0Qcz+xGXy7kQVzHpjVmgkNdxcouwATrgAnUq
MQoH//yXtcjp57LHAct2CEleNvChuSu3z7wbkPdzxT9DgOxNVux+kokpZLsK+EUzuarkgN33qGvT
TRGojAZJodS1S26Ny7Rd3DifMpQwuY74fF+CmczioZA758vDgRJBNfZA2J4J0vKFVeTjKYBql7UY
RT7cxaIhY4O970wD/JrgM1q5588uFoQQglMBImvn4WglhcAd8F11Vau/jLB4lqnhHRJwnkmjAiu7
hvpdOPnWf/hB7rEmXN7aJDqjuVGFDIH1oB8CI6fEy81mw62q44cqdx00uatv336zQXcYzsaOtFxq
BQ4ZTJkRSckfZj0oRLw6yVjbEIYjW39hv5bWFCRYnjNw0jisp+qZ8QjeRqTIuTpY/RiRjvMiNjTQ
RvhHv4QByxNR5BDaKRlII010Xg4b0nv5nN1GxIOh7QG8w+hG8tNsqYiW4B3nFIQ0It+Jl4E2ijMC
lBtYfO5t0UJHm6bT0yzKX36eLcNpIeH/fdGc0raSYuWZGPdUaPW+vW+YohF1nD5PU34vUTCrVmAr
vuozjCDyZN2Vclh7Sxm0npwL/aIwAwuc5mXxvOvkhlkqNZdwawS7fKVJKboWCXciqYnYBZ//NZwK
o+EQF6fkjhj4/2KT9tDxcqaKVp4asIXpvIn7dEkE+ok/urVfRj/ET3mJjj+sUif+huSbbuDELl+X
zXgL3cMBZ+NtUEda5AFWkqvMB/HQ7fEVcXBQKmlFYbwO588vKw9bJI3Y0OlYymfleIv9exP0LuIT
k+akyNkk1JJq5TQ1vp8oVa/PYKqfLFcVZkAqPTH3VLCElvaOKmFHc1hCoSXvPU01z/5XEvZlby4T
MNZBow+oohsVlL6EFYeryP5MVlrM2zbgY1wAmoYu98dtjHwQEq+/WeDrn/UnsSg0jKq9kyE7fN5X
pcc2q2/IMEBRqCF/wHmsfqxLoI7bp8NdvRNOmk3khpRqlil0a6HO6GpCteSvHGa1m8y3vRWt8gy0
dhy3nk/IzaEBbPjvcYlWViHib4ayqSjn/NlUe/bgmbX3ElrsbUq8+wghobWufmF3V4r66hb3gp+Y
mr+YZVqClsfw4fYfN7hnvpwcBBj+ONo1U80mTLDRGEPrwmkWv4C+AKLPfpSPhRfWCVwfD+d0M6ra
5C5UtFvSRPNdpOA8d6LC/xGjBQvTngfGC0ctIXn2YPKF6dMJ1NbGNaNc30QGmilHoUHHq/QMSgt8
xooYSXk8sM0arr0JzQJYkCV7bdY00uinIt2IsjbdbsnM35W1xz7j/jyViHv6ZVIQWbgB4v1yUZ3M
oV++aQwOcxCcqAIwrdunVkXch2YU9Ug6Hqnw5ldTcEI4aUup5DmRCMK27AD2F/g+g2pTGGE++ha8
oaUb8LGfmVFfs5mbs5/VN6QFpQ6x5m6FCfFem3gYL7RK6X8sHJo5ScwX/LZ079iOG3QhIQIplQHQ
bgpIvWFe4l5Y1+3O5eHH20jbJ9GD/DyaeOFTXFTnwUiUF1Oyeh4fp7QT82fqQmiFJi6oGLeVaquV
JX7RREdXSrOUp8omHJHrdmSk+WucxWTwLV5FTRvDtQYKYUYbktYqsZh4jT7QYR1YwDdQGm2XQ1Lb
t1zIDtZsz6dIqNqbcpJiOJE/Eao4bFy9+B4OZq9kOPABQUkOfAu9w0Zyz0ywRZwTc5erup7rCqAQ
9uLN0FI95TGodEPS2jSxczT7ybDuJ6iac50PPH3oKgtBG3fcxuobg3Pxxe77Sfvjo8w2elPOq2FB
sP8+fZeOIsq5Z6GnWrRrYfzm4Jpw6Ejrh0JnzaZXdojkqUdrKXZwdQajyrCcdHMgs5R6cPdO/CUg
385iWc9o/Pg0Ts1lph8T87xEBbSNAW4mHVC3mQ8XQsiT0P1R//iUs/DlJRJvVi75w7eVwX4nLKNC
4k3Wqbt+ebZL5saDt+j6cV7ubrsNVtEObf+LqKm70E4K+JbcXCOL/NlIvognwvJ3LRV4ONpX6Dnt
pHyoxjeTHa3pQh5vKeIhZe4R/ZwxQU8vIL8URh4uNf/uwuOrSrSMCqot4tAvUhC6SNvOlnNTMhvE
RfQv73/E3FSI9+wrkS+H8xA6o5A6ML+Ta8eGJYAYVY1TNYYPFtIBuT3FvhHUCbdTTa7n0U7RvrVs
MQAcnKwPPbTSU27rBSdXxQfeDF+xC2VbZ4wsp1P8OhIuk7Qg4Hf3wVUcuCOiAbRfVMajrWnoRfTQ
aFjo/bKc8NUmNSJ5CnS08T0XxNoxkurLSDxNoVfbzVpwSXQC/bTeGZcHTCZUg60V3/kD2TeSjQ88
cde0zXs9LcT5j6JvY3dEveRRqDLonD7p8Ppp7zdD9yHMKqk0GotoruL39UgJw5iCLD+cJm7cBX2N
sF0dxOgDTJnypxE/wiYcIJnVbPyEu4M8N/xtHZf3XFlrAUnaqqY3bNRaExKYkE0ZlqSUwotsAYCr
plV9vFhF1beQ0WLm5Lf6vZVdRPAmgrJ5MeYcD1+lB/S4OfzLF3CcBR76r31RVTpYjz0YhBgOKsBA
lt8k0rFH7EriPuckGcbkI9qNCCANdVkCQsbVkbpOIK3iqKjNYHgi4P2dGazG13lyuRgO5KV6ClCZ
xJjemfy0afmdvp0+21rmJbyZjVxZD4W4cPhfqgVW1AOV6GhDYdryFt9L/tyZkvsdIRqgzzHkm3k0
zMeZXhYJvzgRtvT3x3rK6VQqz7mdd6BwnelhrtxCx9CKMcmFhgQOO/wYl/sAJkSSoW/02NvK61JK
Q/QCqZ4bHVw9h8BR0PEW1gSLlDWFPLafxCIqmr/tlITFO6nXgTODEJ7jlCwL0D2cIz4ooA39SNQv
DQu2jzW9UNj1YwphOzJZdYiKhRxbA0T5RDJGngn4nUn188ABeFFHFr5GSjoQXZEvBwgmZtYXq6WW
Xr67HDUPu0+UhsruKvcTodp1sIC1u211XiF2nm7tboHfriGdQ2/Yj5/iGOxn/LVXiH5qmQUD4gD8
LSMGM7j73w2HSPa+SsAq9jnVmz/snj3FtnWX/1mvrZzE1jmxfKFazCZXoPDs5X3tZTI11WeSrokn
T960wkrMZiOR8wElWJ+is/l+n+HB6j+TkIQVUaUVoxr5wILYcR0qMiYo9y1QbjoSeVQ06JT9jJm2
Q732Nnz9agfGTNxXm3itBaHsLYe91PslXLWsS8choBokwDZpyOo4XY/jL0JUZlK7kQ7kRlPgGsmV
RSqHU9EFF1sGygkPrSc7Nng4+FcF3gf3KtkdVZph1AQnw4j8fVe3ovpZdXJuwZ+ubXbG2BGFPfBQ
xkjoHQAd1nqlFMF8Eh2SBB8G/iT+lPxqguHddCC9dUliTdlO5vD0BWFdOn0A7yo4i0h6Dyfd1Iu0
ACCzth3IRBTDxXAD12nD1pxYq1dlqDF4LuERoLtZ7bSMkW/+XdWCdWlKuL8OWqbo5vJAQ0YNyFs8
xtpltUwjdsj/y6nQye/ZcJnh1//FEqYp01jJgHCbIbLNprN9XJTd7pmmJHSGFr6dc0NiEbUZCOVJ
wHhlUFeoLZGu704npL54bF3ScU090DHmua2Qg61DTpfc4a4JHJ3rVj3iJVcdyAI/AMDu0tWMa6Ha
GmEf/Bgypn07Ie87hpN+MWLXt9pFPdOLDSjQVbBZfLz3qzfqy96WCsSExQZwE4J6AhZL7B/72H/3
57PUhkZtRRGKNfbLI74B6quhi5KQpdMF7vl6yCMXVMOoKCV8ViDy8wwI2Nd7ZKDQXj2ZrH2drah5
LdtB6bvJLv4vWY5Wr9pBwvGFfjZqqNImLwU57S4nyXw+cUOViSzuUPyTZrEb1IGHJXnns8dQyzRs
hH++mJ36vzG3gkGwc6DCDYKeLop3almYLIhlHvCU3fOr3WYDZMqV40GstEeTECyKcnJAhe38pANj
jGQqezpxnjAESk9FGPye+dgATtGNAkM4XhGqHcFALHIIWv0+Fr1T5I7Z9E2nJC7VTs7He8TwqJDI
KL25No+Be9WiWzdU9ykdghepnQN7iAhsVWDW3JxH7fwGGszHS8OXh1YOMuRBWQOUgiCDDiy5nKix
qTZ4oiuxTzN3NsfQnCNVNgywsNgR/3DmCH6KVBXLWH+t0KIdWu98dYghvKBHsqdyL/DE6aEexcTf
zlwMNVVOR3Ze49ricdQbBkWsRqsikNmGD316vlOjA9tu6W0b0jQY4SiYqMH/ONE+dF/m+AxfsRWO
c0wpbk/TUZHW1C0LSa42bcDA0i7hNWsHqWGpmElCwsTmEIXS4CTrWtCv0COEzfQ7pfYlWDoGeFsO
ThQfTDPBC3SXFysNjvPTHH+Wj/09PI9/A0yIasZ2TPpS8koxVHV6u/0qmiFvrzLjYf6rUfwa8Op/
DxwdmjwLvd4eRZBmHv4rMohctCuCkQi5z1IruVjSTxHo4LZX7JDai6xLhjcRjCKpeXW93LhexvNw
gDs0pVr1V3I6D0uS0UQxmSgNqYwaFvrsVmM/XyzFQvnEvVzbQGaM9H2Bz+xbq+IESGdwIMflhtM6
tflhFXfFn+HDMo814tJVkN+r3KHGWApHmdrJLeYixMj1W9kA4dwZqxNg/gZmFFPQFzT63i7EQAX1
ZGp1dB6cU4Gzj8r6/UPx761O0yhr2OcdhcQNSmDUku/+b8WMVCAO3OjSu16r/tiAGrQu4z9h118S
+xCHcw8AzcPQjlMG1U+kZ8BzW3p26ctpeBygUWh5CFjKfsNd3XFVeyyjjFkTvXRbwKF8Sqgpv6GX
3kX0y682vR3is8B10UBAA4SEd/+dAxiG444dc38u9pLYptdoEqbYpTPxUTS5Rbz2mjk/AtBEGvBH
5af0c3ExPrchKRgNSp/cYudFo3W7+yMCfYNHftJwWoZ+ZBwvClnWeT/sFQsfZbr6wa+qiN0kc+1X
QzuUY2OPLBTBrv1f7uoLVlEIFiG80ZBXksMiXpkRixagBWB8TWgeMxjmk/Sg5WM0CPwcIqgi4G+t
6nDsPglI7hi/gSptFxg5RG4gGXVRpivGXkNlZoXqWGUlfkLHM01lkxWkVKxtmSd9asC6drUByt3a
yBp1XTcRwfTBGMsBbM6fLfz1TDtOa+DakD2NYmO79GP2VVnu7wT+36sOAIxkjZV1y/IMCDStkTko
73AXUql3pcim3CASxtTMF+0GkHtORTfUc4wFV4jG/JtRYpPeifynVtuiRq/5u3cvvEtv7LbkTr45
ml2kzKdzS29vL+2njtD0ORzqpSlOx9mwVQiSCJliAm5hhd4FFN5ah+l0c8NPXgCgeYph2U3ZtzWP
/+uTGYYAXA9L39OE+gSsL0X1aklAB+VhwD8QATN/lWThdtCD7tlPeCT319tRUOMkDupsF4x5/hJt
XVUH9y2ZucWGLbKUHNgCm9sUmaaL0w/Pj8Sjk6zyPpkO5PbgPxdONQq6aYzoU4xtQIHo8beF+GV9
LvBJouYzl/9AgHfmthQYMN1u2wo4VyBiXEB2eFRukhB9zLw3UfB0+iqzuJqFxMZQwnBm2GDje9Bh
L2842zu2vjnDuGlggiBG4fFNy10OVbk0u4D0EgjbeZujib4D2e5oc+4eK6JZjLrj3j2kHMx73p/T
P+3b7sZDJqXJm5OpA85tHp+BGyNt9shtTCapozSjvHPzwlwCz/lFx4QQrK0AG9J4Ma1LCsWw7nBX
CpH933IsHYFTzrB5Ye0QUmFpaWycPiRRYNFCkxfT5aQgxm052E0cITC6Bs6Ue6bxzcO1mNLQ8R9N
d1JIl5p+ahOPr+X++f4CmmFuSIH4TTKeCB7vEnkrmH8TdRTywKxxYrEDEhGS8aaioyBRedghOdhx
80eCq/EEEEDg4GF349hw2ljoQ4itNGp7fwufYNDzxRQpqSssZH2pQp8NqqkmRcn2ZMeByxo0Q45O
7IPUHLGTTrggH97B3XXi1jzoKtHJWrP6swXhAf/7vs0fnJOBMjCot8uGUeBLjzCYiALVn3lwHkXn
fyfDOyPDNHeZgd28zj3xMj+hjRtrppkVytna45tKmf6GpHuE8X58AZBlI3xnria5HN/EdWrdOhLk
98eqhDpz8nhIfE566F4XvsY4L4bkG8p2Cc5iqNtoPH7CM+bf4/6zeEGHgy05CDNpVnbHD5g66/dG
wWNMiKHRww1xEC/gvtvqnWEw7KSyfDjDx/CgN0p7wMU7nVegqr5ozFYjfjnET+UBHnj/sNRM4WOP
+YLjLBv+eUEbmJtu2AaKlZmHcmRlqF/DfdFF+xtzVMHMcicViNkJ6xkiHiLEYebyL6iqhjfW0yUM
Pivn6GxrZ4sqXcFHjjokcwt1OorJewT+vWPThB6WRfRi3jNyKKyLQb3v2AkW0pjn//U7sx+o4CJZ
LhCCzTy4bISRfofXlFR9qlIj8BqP3O0LHWk5qGIGsCHkDzfxc0b9ROBIz8VgiHf+kN5zsJZHYG6A
I0IV1u+hsBn8LE40bhAWvQbxhHr4C6MWMW72u8vWcSD45HdB0X6PJ7BYK4Okrn6frm5EfY1h/vME
V4juP7L//47HfuLn89ThbEO7KcghPeuKFt1lsDHhmXAo6YLRrDIOnb0bODwEcBk3IcOPWvIcqc3X
dAfZ8hSmzQN6wkE1OUWpBb4tmWszF0ghB7tl4fkZW3YaBnT/Ei9pTygq89W3pSmzv2i25VLmBloi
EDt23C2Z2u1PK5rEMmss62s0bYCgs8NKzveKdA9YqBK5sZerpBLmwgYVBd2rbEF9pWd10inRTVw6
Jr/0iUHlRyXIzCnx+si5kPhanwtC/GFIpAKObNHR76tiNiA8CH68bsPIlDY5CG+SbISdT/h3AvFY
kx8Nqu3Hk7aCYHW+PLmrO4VYkov9zV7Ok+PXIpJFXOoagvrQcFGTy5Vmyi8ahiPdEyf5PX3764Z8
BBBq7hDdwvWlFom7fgcev7noQSrfEA3q6R7ic1ToIJYCIn1BN3BWG+McSEz2QahU0NWg28oO2yGs
fvrCgBIRdNewdt7ZUgOH/MU9i8LGrFEhVB/S/wmSsB5AMnFYMCXEl/4kk3j4j420KqgliwZPbkp8
Vfs8Ddny5WAq5ljG+FgCJXKhQ39Xpp0a9kIcVnMt4Ne9QCAfd2zeKC/Nc7SF1iAbaQdBKS9YU1kc
KHVBdKPaoYkwIolj8vPt+KJpwczlc16+FBkElZVW3xqP/cEX6xrvLF9IFclN6wJ8TwP7f4Uk6TSP
h4azb8jttafrVn82pFoej6a8p54NwqdfxZJEXG/pRFJD2VngGH1KI02DukfKXi8sHQeswLI7MQFw
9ZytdjQvPOYmJWMXsr5+CkKAFHwjxTmRSSD/NDABJNYqLNq0YFzkJ9Bdht8SA2yQk9sBRPOCOu96
0W2LSoZx7h8nNsvC9uz113tCfbKkiwQL+1dQb7JCQxU33bZ8i6hH0CzcU1b2yH1fHkQwJGOS5q2W
643P52ogRe06kx9xhqMpM/DZwkxCQ1heBOyRFHvhQwxZK/Q2xMhSoRwEy73EclDDCXm9YeLZtzVw
lf4R+CX7oKRJyPWT4ty1FkdgVzxjGjppzdhCkq/Z79j40yeb7IVvJWxUkiHSJ2WlgqUVIQSPPR1f
jRTQC/zfrHXEtJq+LPTWWT344pYJ/qAnxjbqUfqrT9EC/ruQiFZ1K1B2stIya4XlHz1kZ5CyB71G
IIvNl6ibnL+ce2dTSVnrwAdjYyFtqWwRuXPm8GXCm+3ODGoJEEROioNFTLxcQv7/amhhNSMEHJ9P
lzMqjvc25vItJsh9pTcE4w+7defGfDiodum+5f8QCh3bpmH8JQbXgFz/jiyn6e2+eX8dFWstT1Il
sCBA9QGAC5X5zf/KkXSF1kCW8emTNG1FddD/LO1WBR2FsiksQA0K3nz8WldcZKqNBKYHTSquns/1
J5TYB1bBx05fGYwB9gCy8kBoi4hxQ5Kkuq9ZV/yr4u01h4AAuF+9cYc5n9yQ7GgY7DSDHUlO6NG9
aKnQrgrMYSTsOIrKwC5ikaFlm1FWObCDY16ydVvpXcaBZfIqxQIFt1YuzHO6pyVsnexlT5mbJQzb
xdisrngfd9MGEousZpYXZRfYBO46SAYTcpKX+iFOhwiiLXrd9hpPAM09O6VdZt+JKMfzw1NV5/1/
2DZQ/hWHZd3w43a9fFWa1+uDjKS/AIzG/uZdPOLr+h9m69ODjYaR65bdSRvxgOin56hti02XsfBX
5rjH551cMdHh07xekNzcQSqC1ijEPACvOxutcI0jVIt+rKpAi0O4K+RjRAacvWDpR/1s2vCcIH/r
Rs+laA0Q9oQ54eBCQI/NUo1gjG0VrTHkiCkb15pkUCVNDX3vRhgz3MpkF4AWcGdj3UYHE1Sy4lrx
sms89cvzzoLsFR4W6Gg2oedVbmFJCa9TH3yPQKpM3iBKSa/BHVNqd72HkCwmBCACxgkIjRRxefUP
qofH976UTWrbGmKS1kITLvA11ZcEvbgTLPPeGtD7bYPZW9+/ppqLDQWtCQPxqn9y1EDbRJRfwQen
ebT1rm1VHb5WouL6Z4KvB0hIyi3XAruq3ehJB1g0m9krGGsaFB8yjUGwc2kB6l3WAuoW4hgJiwGP
qXSbnBAE9riQm3R1Z/FfY8j/7n9FlCwKVxJd7enFACvHYFxFm8wFlreNRsObLwCtmsIwYfeukSLA
mYPzjCyZq027tHN7LRa7w/fDvMgstLwICifbc0is0mSU/P/wtdsf3GU7e9Y17g/bo/GV5Ck1UE2I
hdiArT46E7R7PhJlvW7+TDF15KwLOOPcKVyITk9Ft9gzyROd/mmMm/+X5BCgy+aFF7R+MUu/hg43
b8e/iItcJcPXzRspF38RD0Lnw1nzStT1IqaEiiy9rBHkva/VmwnEwvLPjEXbfyYA2/ozeWqMYPdA
VkepXeEwwAJdawqZPlc6kvhE2bMMovNza/iS/zbjS009hS0BOuG1gKzSYX8sSxx1vD8eg09t95NF
+khzUPnv+ftnqPfa8e3fS4+kJRY2fDb5D9Ckz4tmrFycGQUgOmp6/+qqiH4BYn+qAaj3MSq9cqmO
YJ7E8Jt6QjZRay2sumbVbJXQJl7e3ve4EdzdHzz0jxsgFCNVeUrW+ipT+L5KHSuPwt4g1En2pTdz
jAMWLL4zcfR1W/DtM7VTVjruFy91oxsdZfb3+mybmBrcAi79b7ggVfwE53oK89NaRQQdULuw+3Wv
xH5CDuSeDfhZ89zRjjSlPXLrM7VGHjV3P1uqra5IyGJSZBEUetMX2roCffTNuUp26aJu8t/qQwjP
0O9xwlMM9s8WajN2n/CnMCmbZCf3VXj+VMfkHArwl8e0qwT8DVVrNfGCWIQIRfefWeoLZMk1kLoQ
uHBu18jh29iI9ZynXm9+0T8HKvraw3wp2ptm/eeuoEn1GjOtxT96bxAry8kYXnK/iNlXzZ3SvMBq
awgYTgUtbxLoR5a5GCzy+/RzZ655j9oekHpQdL4ZY03ms8S2yCaRWK1KndmcQ1IacaGIhruQkM4z
DUvvxMrD1+/ZauowEqtLGl0LJdoqVnofiO4ypB2vx6egtkd0aO70du8nsP6J81Kq9mUuggBXyjWJ
bYuH3vuMbBRz3DYjUNd8RqEvPWcj03T61hB7eXRdQTAXZYo+8pWZzJYKEjUS49kdA3I/aX/GnUSE
odKzJLVTrmwNwDof7z2Qv3geSiMz+U0Znl5VGNTzaZmLV2x6Vk5i3LUfWp6a5nRD5SVwBSASigW5
kjikCCwn9Br5hoaItjl6ItKfbB/NIBIKuJw2OQSHe0x4iul20r6l1EHXODSht+e0/PBRdqhYsD/Z
50TYOdRu+BD5w+wn+GV6nlMin/0d47pLt1AU3aJP8GU0chOgc/Z6zy2GFxYGJMT26y9y94uZrvpt
vnjiAhqiEf+SiI4gIySAaykitrlm72iwHZXXcPxD2M+AIXE0bnU9awGLtH9A22xdM894S3/0KUkT
7TYaetwqGGk0GphiAokOYIgvKB5LhaxNG1o1P1zdVzaIm5QUIkEBeh74yzqKRd3Z3qwZDuTvpYAL
oWgZzmFUkzddPFt3wFneRYfRwwIxxBFPqf5mdN0QPdyImqMhSdHMDBHpVDltpe/6XASn/XLyupgV
SkrnHUUsArQTNC1uXI9NsJYNJU+OYL1Jv0lj8DVeK9NM2rAto1A/pea7XSlMEig5SQl54fZifonw
9cjdnwv7muZD8ySpjmLy5wDRDFO3TDLs9DW2snXv/g0w4y4eA8QtfT5gZBRHk++53s5cM+v+bA/t
a10nqoAOzwKDATyDDEeptRlLxFPyycX+u18kx0iF97KyjsXmPw2rYJVF7mmWMV5GQScW5cHir5eQ
8lYGJvOLmjgTzO3SGmhl/TR2bWANMDfEdDaFWbepDzNCEcEZEOdc+FaFF9WQq5mSABox8qQP22Yy
p/zPX1b0jBc/e5rPAl8UWCF4iJPO8MICQzIvr2j3xFKARGSIrsj1FoflVTzawn/FNe1EO9024Fw0
wXo/1uOq09TbFmwCH+Ev1UK9krIttxr9p7L5vjCoPZJD7uZnuPKLdaCgLtDvjJYuoAJ1riVPOr65
AIVP3ET/ukwSDyJWy+HWJpNvz4bnKvzU7i/qEprwyoP+0CzMz5x59EYbZ4RFuwR6T2tPhOgPvaXs
TOaUWAAa0xNXzy0i9iFiJ680T//A5Ed5SElAQDrTGLcoQU2Yyl2ViB1k7gPawI5N1Te9Oehpepkw
9tfhKRZlvSK+GFYsQX6tWtzVf+6+qqB7P3nZv2Z68L5xyN5tEYlDusNXEGDBfYADWo20CpXdTCrG
8fKG4zY43H17VvireL5tzgUxJW/TU3UWSa+tApadNN8cRmRI5aXh47GJ/zJdIDkGuK6GY7Q8Cox1
bRmbjyhadfFmOLoZtiOI/ArJWnrtfsseZ2UiCWY961jdMND5/iOIAWCt1jTuhNvtkdRVzaE1cjpE
+NvmssAqD90TWbNkF2ujAKdZm2ZBMU7Hb1GeosFQAKJ8LKEFoyFYlxfRk5zHOsSTzRX+abNlcdIb
tulTz31DV/UKbvQl5gCtVi1tZU7X5w/IQjb0DnmkGSkEEdlzmVKkkS0U0cHqj/PjvVmnc2Th64IV
Rp8SVsdANSsjaIHcvkTCw7mmsPzY3HwlzAthEGpDqRYlkWI9S3NQKMN3tXxNCoO9DrUdlmf6hHOl
CEg2aUyILRM2X5AN08CmqiywN6dHEkR2IyZl56RNfesdDmDK/E3hznqYsLYg3ztjKYMltiqY8DqS
tphuE3Xl/TN/dn4KzfdE1lV2MJ9FKTG3rJLfXM+ZJySrjvo6V9deF6UTmfR990CBUfZdQc/wE2VG
a1luu0AG9F9DYcK9XWvpAH10mnsd9JBa5aaQ8KDgyYgWSitZg0QlFw4cJiinE4P9kAA0+lsontp6
LSmoIQ2Qr7/cgGlHcnCwG3OL0iY8QPn8n3JkK4VNU2yP9VRSDrruXQo6JCSFxHvJ5xQmTynADRnM
KNhWGhNxWG+U2r6rfGUskXPxiRblCSAYL1bgIxiI/1muDgix/S6j+zKlLeQSxs1NlpAgC96Ov3cq
KFrVWnsYAWP+aT0zowommPdvbM86IS/FEgy5Z7QZ/HZhN98MkHcuyrHAZqec733cHCI7LrHqgZDH
WpkMXED1NDnhUlQtkCe5MEDYhowF5HiHVoauVhJwoFq0I6AN2qZ9CP2Tap/vyZYKSa57fJGmMk8d
S0lntUWN1sgK7GXZqKtB+lerDnVhBw6crIWgB/lZs6mqXi96zB75I4zqPRL4Qbr53wtmhn0gVcz/
YQIKOdMnZmJCRplw37pGXJg2YkSI9lPj/q4uvMUOq6NlmOXg0DxBIZrkzMqV1ni8Y/SH+BUupnwe
3NnIBjHzBoqkkxmJqLRJvil53gY5wtDQcDqlzpSjbFbIajhAQ3S8a6o4u9RX4nwoGwZcDEhBOkdx
PR0CjI6C4uyZAOMjBTnkU++AaUy5g8lsCcY70dVAE96JdZURzG7wvxEmbldAGhde55HnfGUav+75
g1OQvJ6tEF579RGSvjadXOzPk8mF3G/Xe4H1YXhorFqp2g8M8NmNJ0DO1ZD90OJZ7gdnjVtXKM6c
nKbAZLXa2EP+nWsM1UlFGNd/ZG8aoSnfEqf1HjNPfZgTRlk0FrUx94SoX+WKda//JB9GAkBQjBNp
I1zr1Q6Y1VWfxqY9/BQqSPkoX5ApINJWcBOYlDA7139SCt4Bn0Iej2XL3yZLIBTgfliMYhMA7nPP
A3I7GRtd2pX02OyuEEiesTR3gAwFkkw578+pxQAXoL56ktexO4oV5xxFiq5Sn+0/NNYg7IGNzHBw
zpWDGclFomWvHrPwHaO0lNLLpcEmT0Q6Gc/HQVLdIBiaK2pNAzB3qJg47A3qL0qw7jKrVP6xqMCx
aiFnjl8j+QCzguuHjb/wq+FYod11Hby1hKiWaGRWy0L1loCb+bSPgZ1ZmP17sAUWLKHohjs0WoU7
dXshMHCDViO+EK/OxqRsevKRPokCMmVH4U8VGvkcrzYiEzb34mB1KJVoQf9JEQgsIRGQkbhflmfQ
wA/Dbu2oM2oVCbKXdrxYoZs9DQEZOuqnG7cjzjsOcJWwFmEtNvV7SE4rBRn84Vz4c9iRS70VKy8M
rZCPw1xBhCnKmsxys3xbwfelc1wSHlZ/kviF6c3D3C8Xsxh3Kp/41kTrB36t0ktQL5OGEAd985XD
tvfrrig3MwLL3fDPwuOROxVTz1637R2OcysH1NmsCOR9E3uvlCrKUqoMU+OZvPfJxZI8gxQxLqBn
pyQAXkIrA0NH8Xoj8dJgk6gG/DU7pcIrg5x6Iec6Ptuv4+I0CrBcLjpT8kP6dY0Dth8K7k/Gnbbk
5WMSVEAiYIwFB1qPo/67UGRgmFkNzKXiQoZ8xs099+CACSLZrWoY4sgbQAtuCNT6RoqOHuhOiXCw
Lo6P1tbeEXXvw9Yu0Us0GeZkmACqWWZ9+5WPCXOCXGolGYQ4pfr3YO2kaGCGNpkV+SfQd4EUkPa4
iLZNt0EYJq6Y6dpmaWvB34CKAA5yQukR6U3PbWcs1LqpKqkVOeMUhR1SfqYE+bIuA7hpHmtff1u2
5uOv21TYUwCfbtgW0pttbaBNeOcQ01vZQ2vOUK5qAo38jf4xhdG8l+Ov5i/Qfcfx6GRARAH3MXW4
TrOo3GUDnpeCKLG1WBAsVO5GPAZ85AnD0AZovZKiQ+VNK2Nw/fKrjE2jgXVgeLpcmkVGPjYzj1up
IYQLTAAWDzOEzju0NP9vgURjj6f5WPcSK4yEhZpbz598kAgBjf5fQquXyL7PR91wlavzqg2XLiHB
YeMZFftYkAEeMwk8eYyri6VanqUlaaCcOrAZOn0Qmb6xezkKZpZfaXk19Vihk347KWyXPSjXf7Bp
s7AWIMQlxwG7cXeegfLcjYuJdEmKWN8wx7iO4N5OEDFhK1bMRnZGX5Yy+UjUPGTqe3VvKdmreGhb
eMhpjK+zGbVV/vXdtcr1ciVvmDYffYbi/wDbGV3JDsvLrdSl2vqxmeOEPA4egPkvzl6hH58mfMw0
mUpveO0zs7D3ddxJfTS/Ojy3bCq+NXrJ3z9MniqJfm19cRgOMURzOAnk6DbWSzK6v0A4VMrzCrJT
8b2y44y6ngYFLaBCxh0m8EFiKQgehNTMBQ8Xm8x+RyOeP5OJwUXCISokAuZCZ/y93FYLSkIQCuos
7PZ7BxkEmh7WWbyWCuqpPn7dRkHObeZw1ISZ6OTNk29MiUSCECVEY4Zv/wq7l0/e7E1zJ6ye79eZ
7AXeu6B9hrcRODI3dFlItt1JtqzTqF2tqpwDKdznKm5WPnRT/vbd3DfNpH/Q4/HDlbOgYkH6tnbz
Noa5zjA80A+Wfl4WGL9QphJHS2mHtcPg85akO6fLM7Q6R8n+KaU9n05seFFeQVBTcsfIKvY8qhNd
nsTUBOwhcDHjODIXpnfv9ySVQA2nhksnSVkbZ+RVvKswh/ob2SIIXwtaelL97aAIRj4TzKgE52rR
78EX+ryldLYyGNoiXDeC7M3aUi8InEZ5WVR20uuJ2aGfUVHDpGXk8OXjJOFTokk9mKJ1hghcDXsa
zcFo0EmfNRdTkUZ5h9Q6oUKAzX29iYgApZ4Fu1RwWPfpjCeKogz8UlKTnlw+9an3s5DI3oMp4C0u
IxMfUN9BFTzQfRkU34d8FTRvlRMzu3m5E2k+igd4CT9MDuVCVOSzfUkz22ZgsS3uJYEb188ZcAVb
V7hqqrA5Rns01EuMPjKn4aGZJG6TxU93izrmKTGb1ZV5/iyWw2poBvpIDdBcMm1yEbLRXt1oyLWN
3YXiYYG9VEF3ZK986YerLxKHf/jQe+HQ3ZXxpIaDr6dT2DCTGVIW8StvXrdYDeqUyz/98+kp/iMZ
aklov9wicFZ6nBvR0tIcGvLKnDsZjoK5hq6d9wa536jxDDHiArtla+a2IFFB2jGwrY2z4S5bt/uI
yvTWGCFG2gssffGzwOB37Q3UnOWwj/ua1jLZjEywlEZjxSPKIt/sVlygD+J1xrXeRUEodOpbPpfp
8z3mqdZ2GjWaS/cDNlOiWtKwaE26a/w9JkxIpqJtaWq7U58QfCWsno2SQuarF7hc1HYY54AsXcLc
vGTrD8r4AVgTvyJMaiIqjDOj2wKXlONRoE2hzuu2c2vtvbeOESnr7ykn/p4RC/K6XqEM63ldn2CY
/2KI7qtrcqbKbr5JVinYlao/9PVnGavh8xzAgWFKNTZVZf5iFz42kZABet9spqea3mwzGbzjoW8N
snZIO/b2hjgkowXyVOcvUnS7JKXvEECytRBUn+79oY3i2FM4OsMsmaRilud1cLofsFg/dpXK4igr
Il4iKAAazs0DJPbX5jw5fW9ALoPN6XjEuFCrJM1y6UZoIkgqz5uccw2S+4LUpSQ3gertXdO4Q/oU
vA3xpN+Z3GniEdzvF33hn96TJURxyWBBRSKo9A0m1DOXKbnDTbG1bctdSqqY4yHQMv+rh8B6W/Uk
XHz8FYzDwJTkK5EFsX/1kGTreqr/EAYdfaICcKYPx2jRBBXHDxNpDtEgIMvwQ+gPIlEcRRtptJ7p
FgwH+x6Cg+BwQ8844wc4SHoRTk4VMZkoIlLtnKxeqiwd6jWxdhlWorZgLDSH3xDbVCpwiiUgzw2J
IQkSjNn9WSzbs6o3NGOLt0PXPMlDysAKHeJtq5k/QzuetLXSWpMWoAMwS3qmH/Rwu2BT07RCUagI
J+BgV3iYMzY7cDveQ1sXYqwIPdFqtXaRHA5thFpXmkfk/ylFrwTnw9cAbZfZ6P6TrqVVXx9wyuHO
AXhdXG/WYfiyKGdSQ/ir7Bx7pqbRNEw1amKXcLTwhYuDMEUuagF17BXmzCoCwLSpHxfo8CkYNJvI
yUf7hHZhTId/wPqoVrFAMfBZ0oJlv7M1EXw66rb7YW+LJ3Oc0DMlBy51rtpnvR3jgpUbCQj+i1Z6
LKG1FA0xywIT/itLSQtf8sjt/Q7nDA+EFnURWdD7PQx2Wys72sx77MstU7xfxY1OQ42VTwnzJvAM
WBZroGxohCLCp282FlFo+bNYQ85UMdyus2ZAHhdiAp9aZg9gnGVqeT/S/wociRYTry6wojjokTfR
+eVEJluc9e9nIY/4AG9T6Dmes/5HqzZ0rYl90Ga36/y52to0WN2cYWvfizGWVwSjjz+tFFKpvNO5
3ryf0yOOJVZmejyCHr+OctoHOe04Uy7RW7HOVWDDrq7lWz6H+0cGoYtE94EdZ/16Ab8Y4+8pElTU
y4Mi8xBL/cN71hoBMLiId1vmWy+Zm2lOGxyeQSpW8aId4J8FzA8XRYBUhNlm3oq6LdtrtQpVim6M
6OpAQhmXxU62ZdCm+TrxItRHoYk+0v0GJi6/lYFcDVp1Td6HISxIqtUV3+golZ3QkHogfWg3jMLC
eomtRod9A/JLFPgDQxTF6UeUFt5dAvNBJVt17m3hE8uhCUkIs3xiJJAvM4i0wAJIWbUwTSReq4wz
EY1AUkSfvPU9dmU30qeCK80eA2ikyoEd+HTw5voLgPHsZIW8nsCPDYcvPkWO8wG7eSWigv/azvPk
W/2q7M558l7cKvMjspxgs2k+Tc0Fsic35499oUp921l5QQFxUPC2sEwYuWHAN6oghRzZUPofddlS
oxUaHA2aYkMCJ6KKbWfKrRsnRxAR0hufa7nBRlwsCunKRblhFptlbPUTJX9sOSk8I5Ma8rdj2nUF
/Gp8IXLbhU7H+tOJHLDTv9+ewiGiL8iGjf9pZPoOOwqI8frtdiHYiYe1wbVAf8jba8tvopdWakwY
sWOL8p4kIPAox4Oi5Uy9Yaejz9d1UDfFc9rYxo+Rwn2EOx3c8dLCZVJzgj1/a4KfnPt7a0/FjmW8
MmzUWQAjepM4NM3xx4rXe3xQXppwGIc/ZZTP5LrCNfG8GJfs//4fbDpUP5qAkukN6602PSm/H1H8
BYgU0aT4OZ6TlKbU0DaEsZwXqcIwbzwNGCoVxMe3uDq0UfVqIk2h+x46CYTlXLnmyMyzorumSiyh
+ZECbNEnUzxBwfHG1PzzVbjHPA76p4axdbzlkqYoq4guO3XjlEs1MLWTJTlJLOex6nPknIrH7RuK
5n+cuJUpJxFzNKlUf7Dg77G1vOEayrjBaPg/MFk/apJUelX8POry/IGOENiPsugA0TSTDhAtYiyO
NOD4JrtgxxACblgCdrUu8mGSygtLDhRzkm84F+xsGWvWw+YxFeihe5NnUMOrSV71dDgOdPz6hjau
ylTsBa6NZrZQiiwDTEQUr9COFVpCchqAHswaO6lKamlQWlTRLR5OzhFcggSvKuludgXqJPKsq2oW
g87+P5jUJBkcVp+WW+iWVndFmpbgFkdTaFGS8/7JQtn7QZWKTPDmIi0yKjwpu5+A0MOmkC7UxTjN
SDy7Ss/Hcmy9cLfhv3vrIcNdOdjHY2Gua45xO+rEf6o9hihjMS+5Aupd+fkhTU+BDMmD1rpV1Kxn
Dh99uOE7H+1qWUkG1OA0Q8mi1DeFB3sRvcYYFzMRuxPdqhzACig5ekkIBSke9+bQAt18PzATyWnh
Y0LmOgTpy4bJ6TKLieqnrCOTz5BIfzNV+nslDpZFzCi34iTseOBW80a6e6sA7b82XKCjWsfClyRN
lDIkb8aiU89jkoGSgZosddqPTd4pKfvM4uatbwy4MQKF6dYVthoJCmuKsSTGzS/X0/obND/OYVtK
q8WZFHzfQ70jBkd3r0Gq3PrPDV6nQ4rHYgMo1mUZqUGMyPJyB3lYg54YkfaMVYS4DKdikpL1bZcZ
I4agLzwQOdHTt09ZLeA35LoPlt2oV62WR2G8/SW4fw75cgXmrjEOC8dtwhyQCr84/UgAMmiz1fQt
g6HkAwzXT22X2rLrlCCGUctBmCZ2pHKVuGczOPq1FD+OR8XgQgUBzEtegykXiTZHLpwbA7JsdP8V
UzVJBVWZrFg6Or0Hj3Ilm4kee5hDMSUpms43WZymVdxG3woWulc2PImbYvRtIcXMXBPt7NsnYoNQ
KSa3jbI97mLP3Ur1tb5oZU0azvK9D37pMwQjUkCWKAI7nhpxuMNuTqNH1hAmYyLv/Wu1qlQyc52i
cc6LMN9rR21p5q78kGCIXSgyWwYQCLcwR4+uSxJHBJQPnFiL4BjL32SbydLldGvF21jt/Hc29QNF
CAG1fvvfIyhjGbAZnfZR+TPpppXDEc8DH/VHizCIESWdaRJMEpeXHzZiXS7IS/A52aCOGTVpR9qZ
nqW/esTsrSHpAafAZRgrag4sGFv7NDo51BdeqPDZ7DkaCJs5mQsKPsrjX882BmVGvXinTDLj+ORy
AzSM6FpA0DapJ/jzVPSmfq4sbOh3K9MM7Mv8WKo0cralYyl5jAFDisQa14rLE8lAr2DKGgFORAR3
ZEmO4+HKw2WxsgRmqHNV+loyw+T/30czvSej209SgHU5eakwTkwCqRu6IZWziKh5Y/nbrxA+gmga
U0fGa/5+zMx8whEJCTFAl68+bMXRrshteO11H1ah2pFYcnG2TuABho+LZpDEMHH2j0N26hamoNKU
bz6y3wcLz6CkYef6sxrTQ/GWbDkBJ4ofSS4CRIK72q4JsjJDc5jTSQ7vNgzhX7aJn1jzi7FB1JiH
xBf2SpcIOKJ0zGS8MySdOHfrZ5QIvU1ofW6on/6xa03Fg9UwQtNtR4Kx3syagyFOlXF2pOEHDrx7
OLxOc5hQHuwbx3s25ouDkpOEW40mvrIsPxT4TXSEeGbuiUbqOcf425EUdcEB/usp9hYZhlHFKe5O
oybth/RiYetL2/JB8I/ROR/yMMm7pKhffZzVKlgaI8bIe0v1PrCMiZTq6OCG5sZ4DgtmDetl/qDH
NE3hbHbNn0MVwaWtABItw85a8kOSiiaV0zsFSH9YvnocLeFusbCkI6Pq1rr/NMl2OVdNw0teenis
LWnh8ebjbApWl34X968yfHjAf9Xl/qvS/MOYtPIPcEcD8BT4UfY1mr/IIgoZ5AiDComc0cNOpp0y
TrX87/xRSKLohdi6z/wjJJuHf4zvXMH4+rZFYKLVTheFXGUUiXsCYZcl331pcT2ZoYXLGc4ahio8
tc0p0F17ITrSexRqdxdjwooGRniIoWAO2uEue8iboHWmFEr8nifGuB++2bpDzqciAc1fvvYfinHZ
fLO9NyhuxhBON6UklotCc8MRkhujMoDmNOFnbB/kMXOBvooFCRRrH+KlqhoUpx1ZKxo46DWyANQG
B85CKT9FAF8YTExjizAAxCSaTDKPL3fdnuCQnaQMTlTkf0JWz5QNq024XGNZUWCCofsXiybDKbZd
38JgL73K0ePu64UZ/5PgHdQQjvX1qUW3rrMAyp5Xk4mu6zwOXe3s8JXIZ372UfXbCRRaIdi0F6gG
h8kexZs6tZMu1mLS5H8mie81MvIOMKAxgMk2+flvQCBmARrwpNYzkb0MTjtSxHX4eWr/+KDml7GL
ake8sLiC3g+wYkN2Rcmr1Wz9mdlPz8LlBG572Nt2K1RE4Z8US7uE1vFMIDBzeVRXfwq4+Am9FkK1
HaMuXp5GVGy2leO1PjDJ8FE8ka14NpAfsJExOhid9INVFxGN82L3SWDn/xhd0d9+3M6S/50+3A7f
WU8s2SlyIsMp3Jfc+mpwpS5A2RVczOkE43VnZWH3yi9g25tAIZc4KfTs2gE4gz5Uol/9s9A/UzhI
3n0raHDEXdPcoa5ru1fWacPrFpfwwEgQ5Z1LNe4ZoFMIl/g/99OtzHUxMPu8u2JkZa+FU52wCVAt
P+lROCwFs/EP/7NjoG4yzY29gJX54n/zCM4FLX0L8nk2QgWOCceW2uQZD6+BTEsEUi5gnuPWz2r2
kOAp6dFrcZI2TC0sFOnN7uWk5sZFkiXyB3zYOA7p9CJfW6XGb4rkCETI1yinpt6sFrXzyBg76C9F
kME8i2Os0476NL9MhrVQv4tZJnkzmz/YqlogP+ZZbFma4tv7tGPLOMt+fYSERBKNdqR0CtuneLmd
qFE6hrruoITUWKHtbBiehWiacuxXrOeqq1ROJ0Ey1414WCa67CQVU5b2isusC9rMCrfX2FaA9iAB
3yXjWdrNrWkviO0Ty4y4KrR4IP8F151NcCSAy7MvYALw19OXpX5hO/2clEorJVX9C7ACirnDv7rc
sXC/pmyB7PBYX4KXnDgLoerC4xHwlyP9JoT8Pi1SKvto7g802WyQdr4HS4a3EVABP8kcqo9YvWAB
Npcqxy7whltpcnFBMaw6VoiiJTXIchj//McIgLNMGoZKcup6O5V/V5BmxTRYLodmYxfRdMFGYm+F
XqlxQO4xjVZm4a/P0O+FIRO78JZLzPvsNgftPtl75QdujjHHD6+D4ZCJZNsDHg2Dwj8uUbPzyFKQ
A9pOaYZBR70cMmbz27ZzNN2OQTClOFWVxo/r/DkzPDlDEPz1Iw1KCpCcdpm+0NFrM0P48AvTRzZT
+oYij4NAigXBAF68DAGCcBSqdwWC8uy6NIMCO4oat30LY4/fevqJYouDsvh2Bxlh5jpE7+RaMXc4
tb2+1sApDnRwUw5dYRwPlhiUJ0Np/YiBB1+IsqOPN35whVzTTpCTAP1LKrVgkYFnmJx/V4ovX2BX
UO+W2Z/TCMfyBrfArDycr+KDVYgwOMmEOYxc8pU70EkU2KZ1m1tNMzjfTf18SJ72VxnCV98lsSyb
rTP9eE1AL/859mWTBSGx6orjBV2lNaBJ97G3Zqx1SPSmNI99wl4yuxCCbMMGfbC7dHSB+NFL/3Jp
NazMq1E+BtRwQd0SzpEUjrUK3AMuG/xrzDkdKhPM/s8OzAAFQA8KDZe2FtNFXEecLurOfXe4JFyi
D3xULWGJcx+5hfmF+TH+6IyStOEH4ouWQpEi/z2ysNlTM1mNiRqyhsjllgoFrIDWL7Mjoi1wwT6a
XA57QiqbdfMjQFHw5TgQXwYVqD8qVuurIJvJJzrrimdBZNVaOHsZNaU2WwltedB5t/JIYsnD0rQC
KrTaWtqTc8wOMPrICUiutn8EUddyYsfS5wABJzdbMrM1x9wDWyGr9pRlRnpQGr/2/6UIg1JdXrNX
LWIXooISXHPPeJMP6XH3c6F+EfZpTqVrdSE3bTioIdKbF+RiAEAUmcSC8Pf8HRyG7Q3E2PNVuVLh
xeRiXZsZndwOEs9NksxXn2U19RZ/gI6EaTjyg1ekT36xj32DJiV/UG71ki2E8y3C0X3guGMVU4WK
Wb1wm/5WIoOWxQfM9ZA4/ITgXkx/lcFHmS6CsGzMYdGZvuFQ+wiCmSBy/nPb+ciFKiF1mYUwixrr
KI+Gp2JHpGV7bh5H2ZYitxerpyqOgUTStsfPRFTLGNAUViCnDcu6zmIIlBBG9KRjPI32yH8h0sW5
idaYcSpvdlkgXfX5/8U02lS88pYa3Fdc4bUAR6NVX7uxcfE2JmnpLuXAW2kO8lxFNlc8ajnKspJ6
/hPF5XW0jzWjE7P/RYDJyRfnnrak9hsuCdsiKs0j9asFbULAqGDNcEokKY69t7wGQCYKXwuKZwJ2
+J9fXOdq+OxPDPw+/fDhx2EbmE+MQMSIfENAv3/0dwEXdkAzpljI96lsvW9H5CQQJUYinqD53q3g
FtCOiSVzkuRadtHsKV1lce12q8ZYjv/hTOklskkM/lGOMEAoNXgO9n2QjG0bDgDQz6Ju+5xwMr1v
eGonZGEwjTIAMOOCnjSNodtSWNz9Yw4juwvlw+lPx8iUNNxAoYfceTKlZMWu9isprGyfhVnSISK2
KiGTXFRsG5L3AL0DqyET9U2i2qAf0H9fI5p9171I3whGVa1HwvG47gE/rUBhq/JEDf2GkT5FjS67
acCzkvYGQSrEsdD8519fKKfRjiO3W5D+eKqwEhOfp3tGFy2TctAAze+Ka+oPHE1h2BBMFdf5NSY7
Hg8WZQGKv7cAKyxo6WNNrWURQRVsawURIi60nBIKH0zT/fMtfNYhM73KAinjh3QWhB+YHHLTSIw1
EKf6huZ6pSrtHFZKvAeMjcILA/7JT8yv96DjyUOLUnPYw4wmuoINpYGrSkQfP0Dm86xr7N41/U1r
irb1ToLJ3/FVs8nieXudkSx/mAV++1sej7vAw2slRZcWQZBWiUS6i2rDWJa97LAhOxLGXxqi0895
Igh45c+gfhttPIa9yr4cMpCib5gHTvbv06Kkl8HLBHyzPdvesD4tDf4q+vzlPNci1PQx5+KFUyCy
bM9dAWaOXye61uaQttKj8zFyHIGSyukcH0loHC2kooIYYOyOY0PiAflD5y4QWGc2D6lmtDeO830E
E9k761WOqnPhmD2new3nzbIa0okX6q7keCO3/Hxvv9JuX+Y2jA7OlcIzI1SxEniCetDQciWGN+Ec
Ry5EO8V7Dx62oUCEWSRK5/ND0LRhZkyVxzcga8vGcdCOq+p4TZQApTHdqTEicYwwHiWAsp9V9ycp
nnVA3lz2G6JfYF4i6hqPxVuAqp7I0qd1OpoMPp0KBKyYNeKVJq22VxjQq9xWWCwxF0BylsfMOeTO
RaPPu45VOftEciLUAOxapfJZY9qP64nxR5oqTeFGJ4YJGM8yWOPLaZXY3GwaIn2YoOTk6qm95TQw
znpbVzi3A83Eq7GOr458j/kkFIbzHagFElvPoVg0YLyAq0mST9CnXcuu0CJ4hAQVeGvt8GBDwk0Q
bme2LSwTk5x4YNX61qWIRVvCrWsd2QhCxgubG0i/hXduwTI8d9LbClFacuSKHFnY3bkJvi/0LDl8
EyYzLpmzGfUzO+jKwu9bqWVVfiOgaCH8rSwiV/Yk2+LVEw/cP5pljIlFVuid1FkVA+4T0GZlLQv5
zf4vlk/wM+2FbD+OdI9k8u8qS6KQ1z56HV5UEp+jFHCV1p57aKgF+sfrrUxMGEty7m5rdvHCSpxC
RtHR3/nx+0jo1xjypOVPA+Au09g1dqBiz6QeLtl1OIA7C4ZsKI7F+x8cWJ/1888PHznj3/tbMSut
60KssunTqkyOPIvAEkAzXjk+Jd3dNSNFMtU2PaTVVsoQGhVstESSd8LoAgPKzGm6EoIx7mG7rccA
ghmZ88lYUA1Pw49sQaZjZN/52YwVx2A3ubgdDwsauZdkE0h/uFu5BRimaKc2C6OLtGhEWyWMVn4C
7d4JW3aQb/Pcmf8Rn4FL+AibkXB+39g4ShemKhNIQv8a+sD15GlTaoIt34bmS/J0EddDrPCQPZot
XmrLC5QbTHy2x2iFtaZaJTO0zMox65ynZnf2W5EmKQzFS30AAGu/mAoewMvpfeicEOiSx0TQOxiK
Rgz6tKkiqTlizujv+M/WasZiiPeyDwIq5p4YkzoiMG1aA4R6yNrujD7uF9pgx5VZrEyKRl5uyo4R
FLMa/Y5484xDRdvqqt9HYzGw3epg4DGA8ySkUFA65dav5fksEINohxqGpPRmFeMdR6hPPPcqqRP3
VPlF6JoCys108e7PNW0oE9cXTnGnVR0braurTJgorSgCJZEmkA5OaNDeoAKczM92IGlS/mMcIhdF
CaKaRzWXh3GywtCr8apkHBs/d5bnbblkKnoA4gt+pZUaDUexrQLOutqZibU9upieU2+zAlRnk33m
GsiECiXz5HWG3UcXiUOM7wU5mTr65k16e90dfkyOT9TJyAQAgxOm7wjwDsxjC5PTaT0VSEDbZeGn
2JwIzmU5RyzCmy8NNjcAk5qJIZIevD67l/QWU3WtiBWpmfaPmhkJuKSIzCTYI8m9tQWI09FOJJ25
WSrP7SmG27+qA7h649IRtYefJdQhJGxZwHPOz/SNc5SPQvVBymbCuj/cg16q83mX6QoXPlJL4J5W
tDrhPyyMVLSjPM0Yspr+vohEjG2FlAPhhk7Id4Q8yxaiUoEjtCcYVVSFTu8rWwf2d+kp7TtZPuYo
7r868ISQRGLx8NzXurJZ9LKZLg5oYglWLWVS+UYpil0ij2olDFR4vDh48pi+DPPnNlfsHeQOGmb3
TXy1/Lz+yI4JpFU+ysgTD/a7RrAAEHGj8IF2aZjNyrRybHq22MDxL43qzu5h5iT2ZVVo1UBDxBSI
HcVpN8YmQyKtkA1RMVua2jTL3NiEErdDduMCsqniKpRzFv6XZh+Pv2k7/4+0HYJJd1uBud29rb2s
JkG91CGtWvK4kddWtaHd7q9roC9dYVXCUhYL/Fka+LYS+POhZldSZNhMG7otbEPp2tLocaY4hhQ4
Vbg3jiKOe4vBbT6MbMpJEY/g5IMK8KL/iHMAAPyOu/BdOJI/pWU0QYrHjUgMxQF87a/zX6C5PxED
WBVi0J1VXV5mla0APADCrM75TvCo4j4vIl/X1KbiPjhjo5QAB7hiuHljzbC+v7QNGL4R8E/g2Z0k
+jUdrz0zeictjtjvnsSDZakdgofx4IGqxe7vOE74l+8om2kEBD1unzhatWAkW6vHbIZNZoYQSqcy
LkS8BXI3a4ClJ7OBzm2wEJFtcU5DDgkl5DNO6uWGu6zd24u95iwwL1ISdNqw+EAaEa12jxE7ag0V
bBjbNl0oT1S0uDBZr053TQuhtBKEqP5JH3cyIskvDnXiVDAVG5CWH09U8xrklWjK7HNzD1juuNxf
9PhrRxKQzxcL0cy6ouOQ5nLfTXKHd/0TIIO1X0AsjCTw40td0zipSY1736FRXu/ZQuESsp4pABvn
TWN/pELAFQHtEoAHIp/H662hjkKhZlHUrWSaF6uONI8oNpU6jUJL9l44AEYpTkhvCT+DP2x+KPnp
gkC+T1ld1kLavCYeAwSmqgKZhyeWES1npj0N6ou+skY40Gt5aP1x0l+GmD+ok4paJwCDqG2/fxV2
dhxTP6PMHS8OpBWRLsOVvn7ZH2oHryA2ZKL7yCvWbt9RMlvWeIGmgRgn1wwAG3QN4n+DdC/02rEP
Sn24dXJG8KXm4pt1r01XNFQf0aHDGtYHjGlRiM9gYGzYunz67RMjrZR2OUNHKRPlQhwkhk5yqRHY
6836IVIwrnR3mMvaH27E+e1+9fun+crpviJFJVnNwvqFQq0HeXHDBR4Tka8nEnOPES6LcYSvP2Ya
sJNrjYUngbXpjvJlNyhr3qpYDkVW4orjUzB6TaXVNlOc0K+sNxOJFsKWZCw3Br8HbNf0Rd7X2wox
RHGKpvcmF9dn5Vcoh3Oi805vodTxL7XcnbsyZVqTsxCFRu35f20v4V0iia+6mrVKUKNZL9uFus/7
cwijsFqk3v4XYR9smHWMV5Kb2zm4byWTsvy/VbvFVwPrF3/6XHcoMefLKVl/fngV98UrB9RT2KMb
gfpJjIfEgrUEKOPB5RjuGW5JcHvXaQ46B5aHgrb+21jWxXWoZOQyAZxbJhkYzNwIEiwrZT7FBNP0
3We8vO/3k7tVY+T8fZGFQXctlA/DpgbdZCSb604H0i6UkCKOJTtYkWvb/4e7Yrl+kMjzUuQakxI4
Ztlo8arnVHOBXfoAuEQ5+2TQB1vzrQkwTc7bWyj8+uKkfXQT1TWS4exJTpynFjdZM9iHUOrKn0K8
x/kDfnNhDAzsZ1vuGwWphsPdAn+cLFuhaON0gy3bDClhMyACN9AzzAmDYVeMN6UjHia7scYCmYd/
Q7hHKP1TuMRnzk0+oyyD0jNoHq4ZsYHazQAv17gH0hWoNZfJdPlVfyqB1veDZTqmdrFWKAsb1/xX
vzKXrCDCceoHGEuCLHiYJF/XadqKwmbq3h+H1+AWIJNeegqrtEitNJbXmNjcMjZMU8Lk6j+ZEfd3
t2l/sMEui4YYw8/uSBVtnlhS+aMmZR4thy4CRK85cqCvRvOElJtYuhI/8Gq4dFz3gp25g2B3eZYo
McJQTrO4dWXBxjlF5pTyYCzRMBAhU7Ou337IeGHrWxq208/81wCh2MMzDjaVnIiE0WQ9zcyveFBC
kwUNYRIIk1aQKdXzQDQYn6UVCJBR9WGcOE6LVFEvTI9DVogr/pBYOrrcLxJMSNFxgXylUr7ivSd4
FeFE8WgovN1zZaqwxLbm6ifIjcjfjrJHG5DAgL/LgFCz4o4Gfuv9nXZJ7bGP/btEZaDNMiNl3pF/
V5jba1VYdPLTqd7bK9H0yw0dzLREnefl1Vi6kY8Y3CgAsWHWryumniJTkJ6AL/YPB+JTHU8JVtdr
07s3DZabJRXwHeFOJ9YXDQ6sWTR1i9m48hk80j06dFZseMwZdhoWP7IcGn2NXXinWwndU/7BYDVF
56+OUB+NB7pxRfwVEOaKDw5fZTAACuBEmnMK8sZZgtTNOuK15HSip6r7HVB11xIZk4OrMnJIqO4D
DGtGRbvGXTs4a0W29SEuPyvf7t+GIiJLE+Nvwq6ogRfPKJi0+rkxUurSkhD1gfbe7h1ki/u1gpOZ
eUlFYxn1KkbsT0NTKnjeID/+68KatV/tpLXL0Bb/OxfbNsaBLLtIERua7+Fh+9lQCCtlteHr8+r3
6qfsM73IsurnNaACO0bmrTyoJsSaomRQ2Tx46lHX2RYm5OkQ8TXNXauMxT2U+z4VP6H432NlAEnc
/weCSqs/We1kfyVQpeNm26n8WNtpWSsgpztJ8mWPv83xxvERPPLWW6moZd+saPyf7kyWxlLKrpd6
vvTF+/4rLX5F+lalKdMDw5x2mJ29Br7hIWHGRHETnwA48UD3CwTJmXWWx3w8LrmDl4rvyt3id8MM
379QjuaCXTDjhwCaJcPTj/9Ah724IaUFcfBr9Ck5D1rSHg1G4uglTZBhOYZLhTAMzX8Y6p9QH7NI
CjAbNooyrgE0g1OfDoGDyHBc38ZfMtn94uWN2SAVvTVun2lVpNAvUcdvP+xGuX116yR2m2OwWTOd
aO6NObY6VqZL627JtsQA9e/qx6KG4+jnB/zdG4OOI0MVAPV51piAYTL88amRnMa7GeCq5RnImLDs
6l5oc/sXQLWql9bVjrgnpo9lNhqnnTCwvqQvYXUYt+najhSu7ambc8X7Ds9dpxWXghqgfzDiFJeh
CY6DGYi/9MasO6NG+Gq4BOZACCG6W3t6fh3739Q6ez35b2JzuHwFOQ8CWIf02JLWIYDC0boBTrDG
QZqdnTgcQowt9M7lHf5wK58Gc8K7TJhYSmxlRxXRdqt7Ym/dqKDcMCCHuoRM6thWr7vi5y8UnjgN
vjEZeLTxcfuVvI4Hr59trMRErbkw1Q2gVUn77cHu1b/wVSOEZknrCi0Fgm31BkMRT75MduCYbtz8
C5tJVJw9Rr7FgyRJuOGZxB/3Nemqee80mv9ayFolt088xlEeUkaUlo6bisGhROaZpHdYKNtFbyLq
tO3uALLhZvawJ68Zj9rPJ1vOKVXTmWpQ7d4CcIUyJ8gulPTbLMUIVEXlIKeeM73SJXRZXXngVIFK
t8armV3vokEviwAxEkNOSaIWINI5tHSNprpJXNTDjjZm20fttoBoPtODrnJGjrT0KOI5TQ+lggif
vGztuX9+9TCUDYK+ui5ghkVUG8NcDeYTd7PunxJQm6jxn+tmly/423EMSNGHM/6Pmuj3P9YLlRfV
oWEHNuH+8tVr+IIdqJd0e0jMrcrbG5BGYaFNS81zbtQdBZWNkq4bTVrh1V9s8M0VVT7nm5d8+koX
+nwksaWgUBsbzh7Oli3zB8d61LVBB9xAyNZN3YsbOy/UfAeP0uok13u9VANJByxX6R2Y1Mw9B1Uf
mfGsrcr+hKEiw9BpuTYWS/t8tWDkq+ANjGAxAf9QA2FXfI2PDnrSb1mEjmglRf3B1U9TFnGhSDxX
HCvD0sq2cYPqXny/vItM9f1bKfG3KU8MLuoz0Hamj6D+TQl+yV13jy/wbejR70Ss091GnRQPzmPX
hoHibejMu11bYKMPiqbQxwrqF5rpw6A+wl/N0qpH9IxW5hzajKcoC9RvM5DzN47ka7YPg20vb+W+
73t6F1WKhS4PCa5wHq/yuXmn+TMR9GGKm4Hw4bZeRNNdnBxXMeecZpvJ8Zgd5/QIWt7ZjjXalbZt
WFvqH2IRJBXrCGFRqggXls/o8VcHBUtVLeYEtWTIqx61d6Und2ACdTDUGR9l7kW4TPVXKTsN8e3V
nPVm/zbPiisjYcBMfQO1u6vTccNA2jH9rY6pnPO9YXKBN7px2jfsjhbc6+1HBsLSiDZ7Y2aZ1gxY
uyTR628FUvCgwNhlodFTe8EjYoXeekPbOU2D9hN4C4ENYYFFSofMU/5XNOguBxEeG3ivKRa1WBJk
soh5gcZbCHgfjbwuLkHRL1xUSQZbrjCBvXZ3JfsEXff72E7gVxBZlweb+rIjQHHNP8NvR7va2Twz
OQQuCTUoLuIClgXpOTCthcwSSgMFPVvegY7119JSoq3ozEHhyRwVGvhjIZWZ+2NrXrdOiXA9KriL
EwcJ082ziXikZhsMc+O3XQi2cK9oRP3rUbq8vglP0M0BkD6l6R9qKw+xV3sUIrarjUZSr1ic2KMc
y211kaktKj6+W+FDtLlohKiTXns9UTgPTUfDMz2ltUkLuJzOUsMk1DY7BAQOgooVJ7cZP62gdKqo
ssqmrZRaq8WhPsqDNvBGd6Men5+0gYu4lfcuG32JnfLVVSlxhgnvP/+Fzp05poLYJAct8EtplSfS
QQDPwrBZ0LnoiGcB2ViycjUz2ciMPY97mD+b6f2c19Tk8nEfNfi1cFscUQWKko+NbhcOsvFdKHuj
KiZZVo3NEm312spVKgVO88iWLZzWqDcKjEWwXrICni254KGsaM3wKxMWSAk7GHzxtV00232o1/Gg
A7UM2K3+X/FTUOFmHHFXghZxBewlJGLZJ8F7fumVX2kXCtV1NehTn6bJew4yKFwNYdsiLbsH+q6B
MTZLiJRzamuXVSDQ/eUxzorm1u1q8GlDOFEKNdi7SpOhAQPP4GhaP3jVFPmF1AcjWZXu+zULJDEP
99sR5RpMCxTjojd1yfkmwHjhwNFIjKT7HYjTRcbgdOe7u8Fx/GSGK3VADzG2GE232KVknF8iyvIw
cleG5WVtw5bYFXmzeM34CEJRqxec7Dpz97CFOiXCyErn86MMj3svvRQSA66gweyHw5d3k+QaAqXr
YJX4XP0ecW+wT2x5h5kjjcwTYky4hDe4EhUokErC8POD0VSKM6UEAlObafHiH5hTWuYr/57hiWKP
dLsirjZoIYeqeVyao3uS9n8koFgFNlraGETGO70eEl0MQoc6emI6rMqqt1FOIyeT82U3cWcUsecm
qEDKP/n9PiFKqjlY+ZcvpP5NIeNeP+3s+PGURaTYfgt05UJ6kg5+ftSlZvqhq83qrl74mCrDe2Li
VsYJCKUzDYdbBcLHXPOveIkwwTxrZ7xiBUsTSvgjwa0schJ2W6SKBA5tDCpZYGMHEoYqZv12+ZDD
oFTqrdRt5Eri5ATHO5vTmkOcVEGgaFRRYWXsOQ6u1r93voUVo8QtzcMr+fV+hRJCLcNv5/Fwxz7z
WMr4kMlhC6MXYdEMnx/17QKrF/QC+rtUEnJRVHBvQ1MQtcoqKOBViqVGIK5eRkSWdj1vBgIqErAj
3pzhGltVbWgNQBIe1dwJDn8pfYYg6Q6YAUmAF0P5lQrAgA6ew5zqcrU9TRbAXB+JbG2AOZ7yJevw
SWrw1A/Lt8KRhPTeWUSpKWgZvgUYCOR+M5RB+zm5H9aoeg77w/RwUujyLSGUX2sIbJza53DDp1bg
yM4Qc4AslkoMnRXbZMA9N5BKnLEX51d7GIoJsaPnaldad60WQlUMiGOTm6Gc4RWFr0964oQ/E26D
5MBRIDuQcmFhNPSMrVTW2L34bZZqQdyepA5HhY9BKRBl81v6V4DIKS8o94d550AGdw4K4r5bXOj2
aN1eKWAdMgJ2ZlZoLt/QIsrTXtxkkASX1xNGswEc8rFGDZyqh/2dhgxsEynESaMK2F5ZeTkwuV+9
mlZXKrKEa7Ygvo738HT+S7spHFNRPKzNoiE5+iIXHf/w+tHLkzUNhnRmJLID4TU5Qdrk+iVoim7G
TL/o0oqLGqMxv/JMNE19jB2jETQlhAm8MGvauf5cUWFeLiQrIQ/+wEibp1ykVpYOCvA3fSwCILWI
DNssZozKf6ZkIiHVvvJgXW1KzsNbkRmhGyWInuB3a+mM9Fzb5cIXG0X3DaqZ6/39uDdeguFyxl+y
00DYDHt8Rh4r1AFfFkuwja5kBjY6Hx12YNmhQhyd4TLJYkNSJqGqlkQ3+Yd2qD09eTiHts1OPaQH
q2U6BlJOcTDbVxrNmnbT6OK0N33Fvya4BzHvwmBah2VctRJrZOXMJsDga3RECqmU9oqAVt4SY8SS
PWrNBcUEs9sqJCCwXgDs6UrafnOnE3cEqwQxcqDCWv/+hoJCutM5mZoXtS8UMok/VfDMdSTm8veN
aRol1zfVZ9j14k3m0v1ohi2EkkuQu6Q1Cy7Qk4i3PQ7x7JRCtNRQSEwL1nLS3xKGsPPiAmLJWs8i
b+ws0XVtxFPGgvrGFOu3Da+hTtTgFkGNDmn8W/ijqCZ7XNEzQBgPvUBx8hZagzteTSrNUA4rd3vq
l+4NPK0T5BNKTPuIt56jgt/frTDjqG12XdfKJo98UFvSVBtIZ54Z1Sc76ocPMosEyjPXx7uvehip
IunwgGfv9hvjqK4gXhhLjQjGQAcE5nrWrPZ5zzl3JVZhM5rhlBdsLQ0Mf8OuHEkgHKgRLVFICsD4
3GWvdRxkq4IxUM3oYdYvVUjlUdiAJpu8dabjeaLtQjL3zDntwxq3a532nKFc58kxfWKHzQw0P9Jd
evf61wG+l7gRchmFwDVbowt+diBxqgddJ4mGMU5gKEQwwdjDxHV69UcisjTP8cKuAfk96168crqG
zxElu31P6csFMVc9CiWs9KscNW+6dW0oC0q5IjvwCZl1MNptw3X7G2bMARkuYMKWwQ9ezJb8pk/s
IW/SZFsj5u2/3vpIWTZ1cJDiz2XNCuCHa2HflZZ0YNN7Qv6vV67O8GYie/v1UK3s6phiIr4KBICH
uywkf5eZQ2/UaDVGAXsE6evXC6wL/AVLS+4lj+6jNHXSLHgcT7E9N/OKPUizCwfBSwEoDih27jVD
vZNlY9+BVygHH+PUo/cJRI9YMQCFzW6U8EVRgGEGvsX80DdndCDkW9IcUytlzWa063H+kaxWjzfL
U2VAQctN6Zllcdd4OjrG1W+0hwFJDmH3sbzRhQvBC0gAGmEgs/LkuOFnaaFUgKItmhofoWxqK3C2
boSA1bpMlh5eCrp2ZulVhJdEYrkvaEi6ulHMn7TXNZtlSN8qs8nlrf7ZDH9EO671zATLZvUh/Mzk
yWwqXVL3azyMMoxN78ML5NNi//tJ+ubNMnTQhe5VFZGFMZ8JurnMS+mAJCvGle/l97MHxIKEYAMl
Zl9iwsXEjSrSUQwfgpRoyUlgiRAiI34eAAm2fHWnYzEQfVIDW1BWPf1n2baXvLdfSvI4lPXYxxLx
eoYG9Xhgxej2KMWrGJg3s8n73qzPE+hM7Cu8ROjMmQIgH5YTy7L+1e/bBMVRDRyo7Luphlb/hIAd
MC/9WyhrA6XBkSYoLFDearaZnAi47OunMrZ/HTDvOmGLooQAM45Ct4NYiVSTGftbmbIYBzWKCVtR
6YN5JsaYtf6UjPMdH4pkLr/LaOC8DZeXqChyxzIC9uNTQD+TTytEVigekWIJHrlIluAncRTyWMcB
DDv504Gj/B+bEqfCXMUrvVoOUBOpQZXgG8c71VVnDUEirNc5Lq9tBM0g8mDdg9HcZBebgpvA2TcT
/7Xc5l9BXrMHrtMiKjz2P6P3w+S9tMeYaxismWPfU9CIWgZHyPdHQUab27QfmPgUWRFgn6Ael8ZG
j2chFJ6VP30KbKFkNGzgJcwa7fuKWLKTDY+Zn6BUxC9LmrMIzWA1a6kID7Jq+bqYnLOO1ua7oACw
SznpE08Wdgj/EzqH9vHp+RBFNScB3ZDNeE97Ftfurc/8ax1prY+0Fkq7N8rOw/4QkW7JaKnjUcNi
V/BAHp7HZqAG8cOSw7u9p2QE2AqGqquLvIz9t8+YgM/d9SyeWtzvu5es0JYCS1k27DNYJd7tGbZH
VJAf+6aMcPi6gVXvoE7h25d0S1Of3PJjfXTsJmrqskqLcqBVgLGGqI0k2tvSmzg52llvq2LGC/5X
/tTXK1LItgS2K+IMUkTs/aiXOyK/VAqF3m8+XfpKho+pkB1Z2ZKQo2gcVkAGCIW9Gm2U9jbK26f+
G01QzS1ywX50qFUSR72GDwPgLCxDsujJoi/n/pbsAE1gT+OJujrb6PhAXAf8MMJtynZBiYFg/SAN
sXcp0/dU6vuFuSm0xJbM7Mx9JTe1hrLRGXozieQ7J/4R+yQPD/JTjRLnoW0bfVNUmJ1/IXc7OfFF
Wb4XAgxMmkFDJHQu7HgxfzPtGAmV3LhC7CxkuvypfX6i+hXbRAbOWGyJVYD85Z4Rcyoj3xvZE/RM
RwYlom2FyrPPDbBOsb1e9eUnj6mGjFh2JL1C/WvG2ScUtw49BWgvxnSgLcU5qg6VNMEMtvQjKQv9
8TS7nj/MKyYfaRgGbUwCjQ6lxrPwuhcSu6Th6B/E/tRwoNWk0Q6IggJW0OA/5x1+o52NFwfzbRP0
Vz7XmMoSLZUzI82Le7kwRXMEM1m6SSBpAizkanxlmdnFnG+FA9FQXPoFuGg6XCS4fxbd/D6hY7ld
0gdcFJWGnJL9AYJOPJgBE9HdECIRxNPXr5AlwZ8e6kSAT4chuEF4jC9P0yns9gQvAqvNdrfPEGSb
fktfkPDreE47MspRE1izWBcrt/5VvjlcJ6tsDERsokf8rlle4nm66QTMJg2gnmeZbPb2Rd2yuvo1
i6qqYkgk9MnfKd+DacbBIyOg3WLhb+DWuWwMsfn8RJIQJ4lqNQB51sdqTZo74lGhGBc2ZIA51bS3
g5iZT/CKshR9x0pEzHVbItugS2njmAYvznq8ZM24LPMWrhSngoprG84g9u3X4lTaJpH/eXlP/4OI
PXOD38BajmTR9kGBWXW8KBdWjC18x5PE7xyar0bw23OiS56ykID5h6I99ZTYEA3zQ2gimel4XhCn
VY23jQroejajlZ4/k8QpdpbCJADOHLMSLNxxesY2XMmp4oGrpefthkfTJxiTyWX4hMz/9UwO2Xbh
4+hevc2OzfuXGXwgGzSxm7SGVr66H6czwiolMEAoo3h4wlcW0RpX/4d/ea3KhzDBRLCOAUzZPIRv
ypz2tchuICdc8mPkZ8RLg71BoPeUGeGFG/D6YUZ4i0TGwBSl2+tEtMPyJRiHxb5fD47H79kdWlGT
nbX5U+GCCFa55aNVjUT5Qn2OB8WsCHTawZgGlNrSgc/YQE8n0+sWXb1R/DVJ51qDCwLnQ9uvL/et
MewO8lzFmRl6TBth3je9+A9EHatfpL9Q1+RHgNqMDqi29WyKCPV7vPWF2aC0/mg44i7oADd/ntmo
BBcq8OLjExPmwFoxWuEuBK9bl1ZylIyqwhvmQdVBsoaVKyT5MuNqYh25y8PljAaEOWtp4vWxgnPP
eXvvQ4yhcfKTKS0Lsy6GDnIb7S9+C22xyJx3NPaOYdta+IYky4Db4NFrmrZ704eEgxHEpl6gzBMt
stkTrck3Sgw8r6G3hUjc9v+KhZkfSBR5LnCz0RQUUZuIl5RHUSAz3sFz2SQGUsioUlH4WGSGmH4T
1cimPNm2GdPAnzfarw7RQkKUZ3uCWVuGduermlDluZllXhEaLMFn2FZYIt7gJRlQG/ZJP+hJJFOA
Nig+/btHpj2e/fbFLo0Dk/n0W4bmTTkqEQ9emVc2AUCsr8Qns0ZKJ6JVJeMNCh6c13TGd1LBZO/D
mvB4NlMO6MCiydxde3Zde3/nfbs6qLUJFZVm8FGSS7beTzglPihc6ZvvDipjH1BDQP9JuF5QV2nL
eGasQRl1zP1jenFT7kTvfgCz7ABvjmKk5lQvVjExMTIWIGlVPwfQop3VWmEdEiBnTSjwVQvVvPDl
Jsg+z1SEOoFTcRKSDZuqjSKgHeA/4IqH95qW0I/pkzEyPP/wSxjpwZCGk3V9YSWXqQbvpK9f6/KB
Hi/NmbUr6mo15rEqjz69WLI/m+8ILlYFtqv2RfvYrDLXAOlj+wDuk/GGOChiadW0Tjlb3BSjZofN
Z+R1mxjQMXZ/QGkoZVGD5O76vZlSGvr+tJQOZZa6eHmXsg2dRP/GA5XyYGRSsOGwAZeoZy8GICLv
/c7hMs9DAe+6Nt1T7wJ+RdODeARpLZ48g/YThdWvMCcy5557/lgDAB9F9TCxbLbh/EtgcqDBPDn8
2yfYp1Xu7WMykBYnTFxaUewEzgMNjBpgYvbG/kS5wwyWxhMQ7u3mwvzYReEADCT84DpMx83Joi+e
9bTPJX7wKLGks5vFjRMKumiNGkebC20GTW78+ekTLB1iTs4X7UKrzD3XiWBOItLOsqj/wu5hdeFv
IdOGDO5A1K9Kuv0oy0NgzJ+zJI0zxeZuel9NSy0EUBrNXoFuNaMrB3cIsQFLp/32vn3YsYFbjhd0
txdp63X0OLl4+G6rl7iyZTF0HiN32ZqTFGl8FgWK3Dbk+LyhdsogbFGBeR8ocjkJoq3Yas9PJCNW
Vn0EnWKRDyf0dJTYBHsIDmONx5f4Vm/2fQ76XM4e/1v9C7YumapEpm8b6pC57rakDTnOPkUgGsC8
hS9NwZNAi5LgggCOu26CR0zHN0jl9w9qS4Lk07kaLRCb0pWYHySQ2LKaFV75tyH0xs2TIJFNJ5xn
0iZd1sJG3saNLHpnkFbAZFfPc1N5wU962uL4j4L3nErbjTfA6Yn4Bblq6hCKlzWZ4uhQtiHVo2dL
ava1gu6yqamvFk9/yThIr6XPN2j/KoKbg7ChWdqDOSS39KX0lnewCJC7aRmfDUAD5xsdoNjCxFAH
f9SAHFXPYaIjTJAs8X7eO5vsv4KhqTMpMc9HVO9mNEm2TyOIWiOKCxuHHgOzC6mr7zb1tGdjR2y5
2FZmqVW/UuF/2D2q6yRG4Cx8Ju1GB0kFklS1/18vmywGUrN1lXUsQ+vSFdlh1qiXVb0SJ+zQhQjn
d6MCjbDhyL6a2U5jfW2rf6WQkGUKhthQFEv4+aw6mESJ/vtJUaiuBR2PPX9gzK+Of1GDJFa+fLOV
dKMS1Ej+4jtnf5ZKZ1/vksfoxtKN0Vu0lpgiXMh5tRAsE6nhNMT7Ea+LzuEs6cI/MYdXxYNuHtRL
4eaSORu97wqXzn77iS0vIHC7QyNXbX5Fj/37FxGsrf6apE2ZXNUPAn+FlkG7xCr9d5gnZG1CjdRI
PzqrZVSIUKjyIzBPs/KobkIL/4Zup7adrJzT7BPK8GN8Qe2xChl8vWFOLxSjm9puDzuOc7sQQfrT
FMU0CElxZ8utCykJl7vB1MRvWhExjvM4LMZLyDve1KSmlzafzMOCG7B7qYGwGpqR6cd+J2ud+6G8
4CpK9us2giVKIisnR5ZTdQTwp4a57ZnStoEVjkFaeUQzi7ouK4ABIejb8yXyfoN//Ybo+PDT7G+Z
puE1Se4bYR4+lPRVeRodo9ZvDLMUTmsVVsez/ogclFWQTvX12HCVdJxjk97j13/v1i+5WCMG3I93
pdL1Ep/NQBVWzu0PNjlx2EUXRKMAujJxhXtEXQNiAsJTnOQSxRdiG0eD1WU6Q/5+/Lj6WJ5hAK19
uBRihqO2Sb1XIYXcoqdE9CEpBpi8+xBN52uygiet8O/QslQDybeF9iMXdK7ZJ0BsKZ1aMkZNxuir
HaP7tTuJkzme02mrZNgR96QSaBUIqa7drQcGIcAEz6DowBNFBaYoP7N3/KgCB90RNVx1i8LFgBuW
KfsakMayHMrRCGsa9coLUiRL24MV078LS2GLQeyj4y9sMWYgxJcZkO1HbKadsGYeZB3z0l25G4lB
0wZNy3bJd5Ia1uKNsjG7n4MN9z9KLaRjJyVkyZmuoS8uPpROS0gxvTp2ArVbgeX+o+YyzRTg5J92
+6cTAWJpjTBQYlGgmYthy12SsuXesrXlSpc5LhqHL1TUrJAnJE9mjd3CKEUkClGM4Ztssytas3Ig
EQsSpRjlTBBDATZI7c/VGo6S3WqnBrLPxqI8fkkk4dfkCkAeBM+P6SUZHUJDXBPccjgk8TJ9ynEq
lcqG3W07qflG2erwgC1J7mm9TLnEI/AG9zz28zTtd+qnQr/3SgBi+uMdGNNVilA5rHndnWrSYx+2
iXU7dZ8+A/qDKdvsHLWXs3hW7S5dDEtAc5tE0f+UtLU0+o0YTs9O7xhzkrdfg1BGJPLGHld7+fR0
Cx2gQp3VQA7AiYtWyJfAzkQjS1L5eGqTwjJpJGsfIusBU5sf2ZX4eGn9eXKJP59UXGoyIdqdwDuJ
zGqNVqKyhgv84ymKbQE1vfVj8l4YyuBp0naMIjUu/Fm/htMp5fufLRhigu39vVA/QEIGwk8kggG5
hrwXHctTdy33+8EoV/SMM5lzRZSCugF+bn7vSZn/TsQJB0RXJs0dcgBif1zoBE9fs8sisKm7UUgT
pC1iXT+HAzjMiujJ/V9Fe23U3HwXAA92xB6BGtpcBFEl+ZZmzMNswcAXD+MUAYS78N/mQp7Qkfs/
xwwu2r4h3baKjzER60g55hR2E9cZ/OhqW93YWXGmK3wrI4t4Qvq09rpDSQ2oxqveI5Eac79jCDP/
FBGpSgMcqmBmzLLSpMYwe1Bna76mQA0C3Z8eRGaX0zhufZHPmjMsFyMy8ukv7o7b/JLWXLX6k4sb
4YFFLUqkWUTzHWLMyXTGowThP6HPBWX7Q/5V/SX+8iZybtc22mZQz7e58DWyuVfFxZGzO2zpCQs1
28OfWhPg9J3Z5SaGGxl/rkwAAyZwQcKjeWf30+Vp7vRwpjfZdPYsl7e4jJQ+nMuMdG29wpFFdw3k
lCrjnHNBCXdhtbW0fEbj0MGmFXvHHWV6BWUNt2cUrolfg0Gj4/4Z5RFPjZB8qw4P2qq+vGDtLcp0
0drdMgOHa1O4v5wIscX1PcpFl9sGg1VCcSP8zlTHJOeT5Hmf6g7JAx0ZR4myCS0wBTis4somEcJR
GNlAQDfm2sktWu+sm70YpxeT3B512vWyZ/u+7+Z/5mjoN6FG5zMYIfGiWjR7vFJtWPnJhAwovjsM
CBL9hw1DfcNIF0u1uP37BEYuZSc1QPoaNRWp26SeGXNbhmXGeCbQqe0DhFefs0xDj8taX5FwcDCO
QyfMsKktisMj66Jq2udI4pcvbjhDez6KGj5tedQ7MGygiKdqUOeftbtUGpJSGIO+I6qdJ7mCwj/9
rFNE63FZqH5owR6RafTxDekCrl2jiPBlnh2hfp6T14MT/vvEVuDYe/4ClADA272NrpoSy+8RPK6u
db7YPy132PVn8xl5BOzsHQIXUwTWq5DuUSLkGNc8jcJFvtlMpmEDE3oKkBE1BBEh37WtGpRTdOQh
i9OIov1/S7nOUjjHxt8OdOARUQyOSgcn5SDixuZJiimJWVxgdPjheKm8ta7jDL+8HAa7qov5OHOc
ndhcv28YTDCpN5fBcFp9CfWwTgtATRh/G435ucczGe2eTggKlKiLtsEvpaplP7qnTJ3S4E4wE3q2
38FC77TtDiiONtnVyCBI6sckUyqjxLBg0MmikDuzTbZm1vD0CFfaK2Mn3zsYXxTZJ/G0zR9bWIIb
MXzuLqNcFTeZ7mbWgvhNazAyjN+Yt7qEJlTwuG0pgFqgIXsqJmcSiatbDBGZQe636Mb3tV3o+A56
ksb2m7qLFAnSdIk8kg7SsoLNs0b4btK2KfW2B7kw33nPA+KnSmiXENZywHN9W7AapMxm/uvsdVIW
eONar2VRJkmJdDbMTTj7II0ZckBdvPUs+dzn7axkTswcHtfcUTj4OSfk9xGaKPLDZkzWONNXvcSW
P0GjbkQjxRpMov17PkQXdY+LIIkNhdEb3CiboTiZr0dwjtQ+A2KdawKWTnGF1QZQJdUoen4knsVl
VBcmWy9A3LONTqdisWF5nzThUMp6Oui/SURF+0/6Z40886LJyjaJD7IFhb+0AbaETjAEe67R9cb6
71pN4MRnigOIqOcqZ1Z5mxdCDHQfUchmRRkmZDvmLaQidPwdjkchS7nuQGcuFFArX/bHlwckfPdB
uW3pYkIGYSU/Upr1oMd8Wxi/GtbvzbHIEG/7vbRQuii8pNsMnG76VUdtiZF9UacmPH/jBkOszzsb
TiLabL9y9jhto2LmFOOvfqXWgCsw+RPx4mFCO2FtpSSU11/FGhR4AB1yY4/BbRzmkfoJZDfSxc9Y
GKxXViIOaO83AyGSC5UfcIBCNWHwa6GTLvumd6/dRW/esPpBuXz2TREBTx2ApH1xslqgn27oXFkT
H5zOQxhgGW5Vp5BcjkW62PF6iBZ69zjjCkk8lVMpEpBGTskiWzX7pAZAlmSX1VW3R+n7AOQo4Ljy
X4am6g+Ny25/eXRtkmu65KaZud8QnyLrTIC07GwveeM8tZzRxqEVtk/cQAk0ixNZFbK+30aasQCI
R6IKmLGMRzdTonir0KWMaD0+EKNhvr5weq0T5uGheli5ec9BFEp2UgGwNBliSYRjxZKndN4+W+b1
YO4jV33xMM6rPFsAE8lpsPy6bUDelWOxQxa7vOIKrP36oKh3eItRgJgVG1b+j5NjJ2ODfjPnY1eq
JbpgJsm5QAo905M3CnUZ7opDNCfmOGfEYqlKv7P/U3BwU87GBEH8jLCzLdhq6GTDiQS1RfnXiKeP
C5eEI7Vg/skjV1gtr614snPe44s8R6O7q7J3J8NNZcyBNgCQJJ5Nx47cLkA4itJleb4+W0UCAkwV
dkt+sIVHq9XSmn4o3EmtRMHLBkmqQbDbPKGN3wjdDzm6oI5FFp798U6Lmmc79LkJSrl22cxzVU4B
dRLwnMggDYcavhnNF+Hf0cCbg9gYdHwCaClz3dQ+H64JtLQl26zhSn3eEWxQ41qt5InPLZFV1+J8
feV5/CtZLf3/o7U4PcoXImR8sQd51rhr9TUu0FrTbEFBv8CMEHNMfYr9B3VDmr1ndJgzZjxrQKHp
vtEJtVnUkaCVDNxYxZTMH9hpuJKy0qezYEWmfKlXO8F1zZ9u20/CCHNGBaMuMuFO67/0GqzIevUY
RydwesFhyhHxZ6gXfu47Dq+hkOEQHCZgfR8sij2WIFMNLmcUY0ixKLZcBJNpbYz8cL6qgHZo0a07
Kimvbbyi9mXYrLb4IcLUS2IhSzkD6DP/TM3ySxg4JHgm51cftIs3nQ6TpkxWczZofw2BmvgUusis
tJclthN1w8+UZG7TEkln+Y4ECx7LHr2hhxe2GiqD0LZANEaGi//qkgx+E+PJpDpmXq9xF3y3gV7G
TGVBQkXIVZQCBFG2PZVeAnsROuDoL/g4ekFehLAl2sUaYFpF9W/SvvmjxCod23vtBR8F2Je1ztxr
NsmCe+pyI5T9Zia4IeplNmX3kpf79pF4NawQmkgi2hQFAaAEmDuLIIEZAsR9tfhsMRahmSl0JtXR
s83gxbEuuxh24iTSbx+P5bM7hjfRrmBELG8fTue6sZa1+BXiaR1FXsHWuN20+9N4I30RaHURP1tj
qF7LsmKdVmBCZVe7q8QidWtGI8QMwFxlQ/YNJ7/LBNZGkWqKDN6qgNP3tFYPX3M2ipNOOt3IORLJ
FrHfnAnx4fir5NQ9JXyM+7phdafZfdF+RQdLjon2Wvma1Sx9+QAGjguMknuO7E34skRj9HW2RUFz
k9EdIyoZlH558vA8AeUNumQAs93A8ErR3QcZAqHy31BLB178kEm99wITsU/0cYRxV4ZkmAF9Hzvj
6hguEGiKhSFK6qYup5yiSTYvSx+NWgt0qx/SSMd30J71uMvgq+ZLi+Dtt63TM3zZBR/hfOcR64ME
AaoR41d4sD52RBMi5JCUObUTMJMPykK9kRG8Sm+FcHnwNXK4EYqdKtGuwoVJHQbJqxm9XBDmf5OA
dppMeJso50DVm4CX72xoE9EciSVYyEksYCz13QGAFHPk0kKLN0ngK8Ej+Z0DunRtGGJeSrP08SzD
MPd1mwOmE/v2VYWQl88NFS14KAnstfXpvPOgzr/pSyH/VWPK3m4k3Fiww+9yM92suVINTiLEhGc2
XIcziyQngfJq/K6E2jvFdOdpAE/cAzQ/dkxAd8/C1ycIhB9TL1EdJB9Q5zR5Bxetojiz0O/oeWyv
HAHtNu6d/MoxUqH0dATt2MVUSTDZf1cz9WY6tBYBFp798rnPiOYDS0Pw8cIKF6arL0Ca5lv2boeI
6OoBESX/5D+rqQKq8jEWvsyXTNid088BqKgctla44okPCcLO2u8YK+4ULCHAO+EF5EL6x3v0dXzk
vnT0wCPqod2ekjy2LUuoOoBM+7fgegk0wMvqcM7qZa4mDc/eZpWUxzgQVewuXJmtOtsZYxhZBrja
wSOEavtoXwRoZvY0scFgAdIOQ187RzYXnxE8lJs2e4pzsDhWR4b2CjyuYk6XjPkiKi0tiP9BQIML
O1v6brW58BpEMH9McKyfZNNAccb9u0wYR8OT5OklrURYJw8DnQ+FLyyf9eJ6zgb5bFLmL3NA34TM
9Po43H8h45oQjGUVupnhL6V5jbtuRURrIwgCYQxeIT8W0xgLGXxFEnifJNBkEwTcX4CZr0yyAjEA
6IQOrkYpXHwpQeHi8XJf1DyHAmxJNzFYIuswtG4jPjMhEUPKvbpT0Zthvll5fPm/XruWoFyZ/OtR
ep1TeUtKnClyFtjObehLFjPNgbFsuaeu53whnadJNplIjzIB8kIBy8vuYiEmB+5rv9PH+ncVjrU5
Qr9q4puJz9UitkPbE/dF2NuqtrB0oHeq0QgIR/9v5Kx6wzjn5DP/O7XvBkhoz4UbxYVWFTckniDf
PIkMdTWJ3jd8gUVCMxfbs10ASpCV2zgFOamXXDRfnscb4tAlH9BolYfmLsMf4s8sRzV/wSu1LWbV
UoQ2pwkH/IhktpCHnkx+0A0HVI3AlIrEr2zfRRFfxEdYsJFNdRsVT+zFRj5Kad7ZNXxJe5MCnCVN
PbcndjVzpFpS5hGdkq++gZ/DBzLSnCqdKRjT/EPfyAD3+TESpFJm9M9LeYaAivvGFuqOs3mj/VVR
EXMNSV80h6sQtnc+7zq6bRut0Wr/WlgKFIz7M0Olh/DtDLft/XYJ66uogDn9vM/ocX0CX6+uOUA3
NJS0dO4gDMILnhAO0NoyxISrl+LAi1sBfFB1zZONe6TY1X9HcYCP8MudLizCCqXYG0aGkH74bHkd
Ck+8JQmOftS4ks9Nzofc4c6w5dtFLPgyLLg8gmavZmWovPDBLQ5I6MzrJPEjklJIG6CeK5Dl9y4+
BHHQL38+1BlXuHpNpkkD4ejhghkCGxYdFCAfKi18bRRjsLTfgMIy/Gfypa7woVOhDnY5/csrfVRM
rjque0A5FsSeo13+1JTQvbsEh21Jf96phXRxTM3vvCpRayLDGgM1eFMDIOH337VZm+wRvR5SNaf9
r86w3td5Die1YHY1emq2ya0EOo87b28u7ywxgp6VawApJ+cRPtCyIKalvuZs0QNlwPECqMPl0r0I
20J+LVf2O1Ur9DUivioqaFxS9VQNECZR01RR54oy4+kxGO5k9RfU9vAwjsSYKzgQ4yyFBDdngNqJ
JFRVtVGzPattFhdc8b9NZ8ynfBbzR7mPKo5Yfq5Qk75ux+h7j0exv1wnZEd+8vbAtdf/N0wjwCtf
bepN5c7vGeoNm5pxzFUTJzBmVkq2rgmJAvfVjGum6NlNUi1+MtlcD2/MverMfVYDBS1shxNPAhEk
OvqwwQDh8O+bu66szRfkNDJKu7BHALFzeNm5uSOOjQtbsvy4uTm8opHJIaQja5kB9gjIjH8Zmv2o
vKtQqSjLaa2TaAUMkgGfmFQftPKtkg2vIl2fgLHKp0U/idb+TifuMp4zlMXqLtL4ikXuMfvt0apP
mioKgNLIz0JfjueCq5m4JrdKl9ADICtvEaI1NC9TOVDJ6fTrLg1744SwbU2pZ3/S/KN3b3pyQkzO
L/5R6hhoO0XjKFPGV40s2acKT34fCnNedEa4VoSeJxnd/0r+5mx24fFUv5P7rMhtKUX0jsgpY4Oi
OZV9fRzfSzbzLXOMWo6FNylsGXt6qlxHvVlleGmk5LooS2EhZ8LbU7Dnc12EZYAWx2SbIuxeVlQa
sAtFLx+o1mSLf+9W1WR2UF5yyX+qLdEF/cydNEw5UTwN+ecAsStqe1yucFXejBvGH0g6xavNYmMC
l1Vj5aBTCIY0y4LKaThhipSdvi9wYX9HHJYmr+NfciRX3zBtO0wOnUct62GATNSo6XzP9b2r1Yd8
Z2Je8Q0JDXD5dGJfv6UVE96gK/sGvcmCXMHVDoM7vYa4SfLxar1SqEco8J9/u/R3M1flK/1jbnyu
NAJ3/dK6D7DmSt9sMo0ae5qsJ9CMkI5qXU4pRNnJbjckSqpJRH9j2MOxa/coCPWA1+fpW67OJZgb
4KSstW2d+hvRDPi/+5KxLtzpe+AI8XZYO5YEP7ad/hijPCqoeIPt0qndjesl30JdsQEBfL4an8fu
uZJZgCkqkYD5axqkqpAFR5DsdtSmq8r7uZhC+ZL+QCjjRldZdPpfxDG39dbRXChln8JXTuBhOphK
7HNzg25EllgsaYIsJQZSN4sL1yddfzPdghZ8C9vIt+jZAPh80eDwRichPBlHKxXmr0vGeDgMRFwG
1EslsE0JDa+ZEV2BGzUAZHWiv+gWfpnWqd3bSXGslsN2zsnuwVXUWJZ2bRgrjf+RbhOrvoj4M2AS
w8lw+wPSBs1bOIOSMVmKJxQPEMgsyDtserKlcS4Ai1f+e07F04tfAvjvEVvFs8++TlGZ/LvpVX34
R+ohm+fjZlfOv8KuyJLl9Wk6LuVh0hLgAnhBY6dvtIzalhwqrLnI1Y5RbhJFBHykbJ03su+0pMZU
39mDT76X7+5Z5mTLHeoLva1pE6xkaVKpOzV/bhOAQHF5O/lwY+BQgaW3yb9c6AuIZKldbZs/lyzV
84z9kxNp83WB9h1nzJrMP7nfUImng+Jn9RV29T+y2Dr81lpoubDUNsBv3EtLUaE/OWMdjd9vKzZ+
zmcx0p5xUrv/15dErUSbCoGiAPLf9ZJkqN0oxVM12E5I2hErl+cxS6ukI2h3i/vT6K/JEWzxsXNe
8/uuIoLp10NSlodYq1TXyHJ8oP/Tp7ySwVR9A4rnqzDguw4/PFctw4Eu/n3rLpthtyyHnNe/x35N
F772At1MOWaNsiCVJONEE4/Mk8kskNHikLWShg6tdkBQRQY5RPJtBMVsAq9V475g8bfZpUHhwhTJ
qaSy1sTnuO2U7N8mPE5b6lhq5XHKEVDiRlwY8a0vpyXUmARTuplZBbn5y841cABhRO6ymqzu40/N
+5CY5hxlnFeMTiQhM0aTjPQ4aSGmx6zHXwenbrirWoD7HuI423QWOlO9RiYfHKekOTB/R/q0r6+M
cmJNUICea056hF07YqFZLFbMmYkzY6hjUHoseoJsPUs28bgcWBSfedwWlXOxW/sAHDPB0OPVV+9v
NbJXTjcMtJ+DktRLaoaJqC+GyAPQybLNAJWHYDA1Ks/0XTNDeRtx1xBCAOcvCZ2SmPj3mogdwoZ4
bH8rjjAHo+f5uoNBA2xsvczCYOwSX/Rh2dfc7ucTYE2b/yno4p/oHQfBxpNEucZULPLN1cpNTmJ8
pdMhliOpVcHE+5A2ZsuzvemL2hSkdzROIB+d/jSPabGwA/eoEVBDwA2u0D6TQFzLBWyf9vgPbCBn
/NZVARvhr7AxWWTDB+l1xDxUHguRTvSRk90bzNwNB1hmldfc1GnF/kC2WxJy7EHiKU1ad9CDfQgX
oRHi9tkpMsyfHtnJnJVWglkDshnkUlAyt58vNUlA+aXDpeTCc+/9yJER/nhakgtXtFjA7Gh/BxXo
Sh58AHfrV0huPQDJlFKmK+1fP2wMP4h1+0FBK4kMl2+gen7Zvn63LIEaUYJa7fzsyh9m4HvEJYgp
hparpRvSwkqDxkBwNcbXw00xZWVLCn4ZFCLwwWP/AvCsyxFjBQtZ/NtoK+DPix8rDDLAkyM83TER
wBXL+Uvb97X/mlvp+q9y7XjTPKSZTIRJE3W4MW36F07j+pbulZYxVnkmEKZw52xlnAEhPRKa12vY
YGgptocXM2IWrTcu6iiKw7DJQMtISScWG9ixX3xEu1Rr8UxnJePDUb2QpRZVGhChNuH/ntdmseLj
qcl8U8qBGCjsVY9zP3c8b5IT+Ji7W1q5+pGsHCMT1iM6DsVxmAEvXKrYZBdNtCCLoqodWCcJG597
od/UrUM/EqjuGaFOY/kOz3aNFphr/J5xEo7bb6E+b580eVhOuaJ4hJGB9TFm8/yNb0UNiDrStpcT
fdyFrfpR9l1XLo59/AYiwNdiiY+KsW+FuhHAKgMXMFvgPT/IHPNFT82h+RbsAMnL0oZtuR0NHR4t
BFrUpU5gkdhKucWwJBi4cD2xRLxsZMkThg2zkoI94MhkWcYhqNbE+cpwAGB8MjJ0wNJGIpcZs2GK
KlyHlO9sWIjWVuuHWiAcYmL8d3F/526m8WMCX8MDLwWYU4z6MNRtIwYUMJx+zDLbcDK699t1kGS0
QLY/F5CvfG89FBitBw0jNyp73tRz+LjeTvLZIXX+c5aV3sHg3J9nQsjmltB5J7oYMcnTnepKkcQn
JNDjkZB6cw3hc0NC8kBVgTa6A3G42V071MhGGw40mMPcK+m7scArT3dnuInSjmFtihOjVKNPodrb
r4VHo868usv6dQWZuOMA/JGgF5o4yD1ZRmEGIiZ5IOm2Ou7zzxJaVJ0311Dr0et+kvkNHztfsggP
yBZcz+uiLTB3UExadftkOjnxUn7AOOwJ7TLC9WfE9oDw80p+FK11x/35JXTzZNB5Vrn/Y1DtItej
jExyYT+7iNrMhSLTsqIMfT+so/txH2GhIIrc/gKt0orwWAWWxV2DsGZLYOn2lcvOCS6qDq/qvqVe
w32T09JZT9/enMo/2OXq9W9vKam9f6ReXB3oTvjDKlgALOPJ3yAqQkr/Pll8/7UZpHoc3Mwge4yE
6a1m1tEd6VaGIox3VZZ6AEKs+zWzGi1bkgA4lDsymrEEGzTuupHy95vdMHWdDm9hX6wTiCgRjRGx
LcqbE9RVcIWnPRQm++vxgckN47dYfzE/Gn3wBdqrxOSTvD/wwiTlhH7AmIX6zu0WsyKP50O8YEV5
Ke5EYayQiRUGa4BAocltluoH86SZNaYeciWAlt9ovMLa/WRdYABQ8mG7D42POdWlRGJaj4s9S/6a
xENkStLnMLffFC+AMnLPlTaNToN0twhsq7HT2D5rOxQlB8OqRfRtMgAFzZtGEkn2yP6WeQt4zQcp
Fdymi1LPVhWsyBwOIEe55y5RMVvYZLsnPSnNZB6MtPtNgVnPuWIZ5h28be6BS45pPjJiamzcv9lT
ExAc7xIiWg+pXxNjQON2yn+8RH4KfdFyRr22XeDstcvDoXyhGDsL2xwHVIbWixhylOn2f6NuAVk9
KE7hJLDek10ocU9TeI6wTNmV2rnvd/5z0mTq28yyZyk9dixDgOXd84V17/2XxfvQD7yp5b1IERzx
6AWj1RHb9RUkTBywBh0sdRbQ5t1C1UUu3CultSvpvSZfSU2NU/IFhNcFo5cCSEu7eMh3BR632Szz
bFN11I0Y+3Xym8z6BIdBONF1Vh4Ai7i+pJZKBnTTc+pmxN43FqXfR3ppCflLq8RXlSnVx63kuTbi
8wsFfSEfLX17nWSnHRULE3WSOq+FHY++rNuWqa5yWEXoUF1lwHwQkhchPyM3hQqcjJ2KsBV827rd
SwIIdO8mGz2voR75Mkbpg4EZdkMHpxFl7acRbLybBtrcljW0gALE5osaB1v5CeJ90o5xCuByaM2p
FlIIoDZ+Sv9M4Io+m1e3n5OdidgEGPRvlrxa9UcEu6iA/5NWZZKIrbDL4jtKKEM7xWwcdhJbm0+D
G2BeN4NONF2jJkVNQBhdcT/GwbzMzSq2KCqCV9KoMH+3eC8s6k169QQvNEV7cCJ9Fis8U7sqd0l5
sGxHNM2k6EP37nrogRGzTocr9KmbfhT7nHsKpSTw9Y4XGTXpDHogb6Yn8y7KUB2ezGmkv2PyIQAg
BdAGpodv2fcokkE1vm8DV8CvJBBx8osWVkMl9CXnjw/RKOtEbXbBUSVBKQbffOiu4J9ZWSDkVCDP
/bluwm28YviC1YnfrSfwX5lt/jYtWvPYKVtHHPwddVKGLVGmd8dEQupL9ZnQyp8VPf6ax6cnrCu7
bDbIQf0f3JaRcWig7ldmd6ZCYlYIl3cEjCvseKddZ/1K2fSy4Fe3sVVSJMdmV20YoHWRfj4Jm4I+
KqUeHx7xF3UmsfgcJovO9gM0/SpsP1OEbXVMwplEC5hO3WZAAzCZGJU6u0DQ42H1kyBg30HCkbty
CdPXUp7qLtzHI1hhBqhR6mHOlabFHD6vbWSSBWLUHUxdY/FIpJrH1UOCFtaGc9zzIHEmNycs+ngw
jm83vJIq6/SpQQMqdNJkd+CL7TatvS6+bccFanyJXDMS86zhhpm4RehDiyCMpZs/m8Q693G23VDk
NoAYTXXwGanzGKb5ifReCAE9LA8+pUce+BvfHTO2Bl4hCauHhXKxrnAKliMce7tsDL57hkmSm6pO
PEfLEeRUjPvuh2Kvk19w/ZEzHlWowEypMKsl9DpPgq0h1EfQm7JlqA/7j29FqzcoT2G4WI0mC9C1
doeQ/91QUnfQ3fcYOCHJPmJVTGyg8DdUYFhaJkAavbFIpMw/FdmJIhVp5Hm5Gq3QlJvv9qxQscZV
d/wfWdfthec1Kin/VSCE3IYGklIafaMO0lQnBKrYJ35gs+BBqTiAUoJRhLOh3Qaw+Joz34+CZM4X
0ufQyoxlncol1AmDpF87rKlafG3+jwXhePsG/rh6FH/vrq7WG8cws08y3O7+i9P1ZEgQX0GICREF
3P13XhUYyBqlmITL2XajxaVpuNTCrZLa9nfJ3K8T58K1f5ZJOjJNKnw3ZvJH45RSGlZmvycAZsgv
QXZ6YZB7Xxbaqb1mmhEV0wQdK7ABpKHDAalKnNRnjQ8F1S+d+ArwBCUhBSboqwh4PNsI9einuGJQ
/xn33G8dvMd4v5q7GjGkakqbCb9O3Ud6faocYUJ4t2ndkvoFPrkbf/PKRU/BInyIrfcVw1+Vn4qF
yxELcIou0Uoezu10v3U2dR8FJabe1c06P10eevzG2L2rMgvXlzFOtdssHyQUShBDuUWKqY0iEknh
0vPdArU8ZJzJENpWHXhFGGVJat8rW/0y9dMaNmwIQemR4sFrC0IJS99c+uG5p9Zz/3P6p4QQORSh
ye4aza7EFMaHh4O55Ky2JzBcuvVaTL37GddClFMTKtUJsLCGSeBjbQ2WO+mMj9jY3rCvowpllsEd
/NWzgdITKTq9IoU82VQggIMi5iAG2Gwty6S/nBmMSSOtn9pEgeEiFWKaD0Q/zZJH0F+h7nTKS/fI
+6gRE3AnJJ1eJBGL6rTi5upZ995tSry4w5Yhjrn2ql5NLQcr/XumNvTMzJXfNjdlGl1vdobQhiy4
86DteSWtK/Rn27cm2VvxBj5LubgXwWyEBCD9LMfIimgDdJ8QtV8k4oAFVw1RF42a6i4xaPhHohHf
MPNMIRZAjjwYdr5ZZ8eQNdQvyqpsIrep5jkHuVPOTjK6SjG/hhLfZ8F6771LP4J9xZXr19+sKesR
B05F2bUPnrtVvFZ7C1t0IsYN9Q0cdGtaJpALD+L5xsKWP51FlNViGqVH+Q9gmy2yQ6ycHlCQzLPF
3g12lIY4S3ZBH2ZuqmOCYSnEozH5RPC98lYUaCzcZdYLwQT5JILvgCZ2hfjC3bwx09KM46JiZNNO
shRlGTsXw0nZ0qdRaIy+ldxpgZ0kdLs1P6gobGpsGxallXSWi2zqstIKCBHdeaX9xGNysmzKMlPJ
NMQH+mZxtHdt0rCV0eAnEdg0h+UVwTAp6hxvyna+ivVZVQ4yrnjzI8O1saPn7Qw8fvGtqwPxSU9B
XbcNo5Qa+8Z89m1u7b/wJXo7tw3ReOMp/caTvY5Zg4wjDuFCmBo4NRNFeLNJwRViiq9abcVLNJiW
/kwoRgIUBTh9E3TO3bpDnT5hUjtRQmKvlqRi4rjKUs7D0BsY+I3Q50XHklGeVZBwNwS++l6epgX+
MhBiYreOm3+0HvtUXViBG+lxQzpJWa3udfyPFJCXp+y1jIeHUNuy9sr9Whi4YgrxKNHBfcEwojIj
kllkIxqSnfqLUgTQ83LQ1Bs1niNmvfKP7pRMdkhhOFI8iw4ZXE3d/tmi7NTsDvpGZozWzRh0NsKG
Pf510ws9Bn6KXWiFxNpHolkX+jLe5stiH4ABRaJ+etvuVTmnZyyqqILwT3NhrSsphPshtyzDQbPh
GE7hdMaKxoq/A3tLnh+bFlhgV0Ls8Hf/Mp3fGbOVUbSRRSk9Ab7cL2SXJlERqWrXsPJxYMEOU30s
SeQpHWgiuqXmFgKQAKtBb2ezrI+gPupQbAeHDEH+7cI51b1uLVvP0sIFwvq0gyiydyT3gB8G6pHV
4g33ZipksMA8pp1MKHfkCClBcldSni5QFxtqV8v7iCInXBsDFVsZWM7kIR81oVH6FTLbgz23jZyQ
/aBYhmohim2HzuXkIQshKxxRHK7igawWvmYsE3nLDg0BvB4lhRUPypav0NTkXL6XqcBLpvwZF9IA
7ymc0wbh15/rcJx5Xc/zkMY4P7uciDoARqeVvydVoJiVnNQD7ryFI4IvRjZkS5kFmMW1Tm0lU+Z3
YLgIdg1ZENHgyRssTD7NhiUWMlNTVQa2gqIGyELaZdgxzjgkefWrcHg5UYPgUAixi/2NMJJio50S
XUb2hx6ZpIVYAnPdFoiuduTGq85wyMe9287b1nz/2oR2rDf83cEYoWzVt/fAqnw92mRpR0D8zVu1
z42wxcTKWhuYQhb24rXrkuulcQeTp1c8TKqfkd8NcYw7FLtLEJe+FAVmRcGXt/5YSEfRXspRgBuH
xhw0mgyRIBMXierBhp4UztuF/6aTj+4usC3lubWUQcLMOgGqXGtxpJyauH6HiSFo0W6rUtWxjOY2
NgL8wBxsbvaiRB32rZL5N+7O+0kIus3vqCgcqlB0dBc2v90pRT89MYvQUxjxrhbLswkA/2dF+Rhk
n2e1AfFK4s4grTsFfKYFUZtlXQh6XKJmxKezhV3ftqyYxTXnXP2pDltDyF3cLE3VSCWaFW+K/Rmt
Wb1foCfZhQAfeoVBT6Y2AwBkJfBL52lRUI7Vl/aMilYD9eei76Ap7skk83k2o5VzbtqfGUUNbB6N
t3BGa7EU96MXDtucmctMzPqJgaDOUbJHp15yB/+umWBLqLCckTH3rTxu5F54+77HTV09MDG3LRij
i/cDzNTb/ARHiZG8JjLmBZYewOGL0ni8DHwNnMznmTwcl1RL3C9WVRjWLa+dcprf7dF+nVf1YSpj
zC8JGBHCukJNx0Hk9QgxmAhvxiNdvOBgnXsuWxRN5FRS6cpghcFZaU1zbwqV6qWW4m97wVdJWefb
NYbkPyMC2mce7Obw7/EfN/nR6NtyL9thu74+vMOpHX1epJB9suCYCLRj8eJJXlYW8Fns3HIrkhVD
4x/076RVCkiX2WHJ8QBLVCOw5Mc6kAoNT/reJz21x8d9A9aQwbTRrWeam9sY+l6s8+XV0yK6Nmlc
JHyIhYf2bE9k2DEpXFx/fHiK24ZdcqXoWVuMXXKoGUaoG12HxsyGmnIM1oWTbhC2Aiq//pbuRPGZ
qXeKjFSmv+n/cOIfmzM/p90LBaqx3+S3Wi5tf3DaOLD4zH2AUG4gHy2knjL1P6Ih0TRYLnpq2zrV
WMfRgWzGaPxkQ2ylOlnpSOIgaRRBTt3tj9T9kDYt4ERn30mejjZg+NYI9WrOAIZmJuTLtEAf7LmQ
IuP2xIF6+1d1NH92SWzrJc36x1CQSFXzR6yw84TBYsaqNiyt3SnsAgSUyL8WCvKTNCBSGfhlV80I
kg+OZiI/FdqLt1QWTxQ4QG5cCDPJvyF2yvtLaDUmhL2AWzwBbLIHtQ2bVzF77urJxnaVI3xH8SnY
25WeSihx23/V+61d5UZLgupVvq2Oxq8OggpR8V+RX7b5z226xRctQTRiZcfNo8fUT+BoA0TL3FFD
kIJsgdOzHoo6W4mc9yOu00Tj1nzMuLhf6CRxkM9dNtmtaVCznaDw35uBJbOJUDtSmuUzk53ENH+I
3kcX6hi/DV0FsAbsF5KypobI2JUOO0gLo19EvpPEt96F73D5ZrJ+TLStv4celf8p7GsDUpTRh6Uv
BzmONJ89xBxJVr3bFyiGleI9Ept/8i2+bO30O2WPXQvlPQrhiezkAD3PJoSZSP+60Jk5NvXjVcfK
W5OlGFRRsseVsOCjwcgIq17IpnhEuzmiyQi7FktLl/WYxRNZbmRTMrPVTOvROEN2Rlp5XpiXgyZK
mJVlm0pI2RqlolAsX3B6sI6sHVp9IAzsm1xx0c32aWWiKkJjLu6vh8iCQls37MhkyXoYg4VjzSZZ
tD6ZDHcvLR6Yzh+GlyNzaOcU2nM0K6oHm7f71gLsxz8wGVSQOH4j8/2fl8ecmn+4hzOjwKFbznOf
41z2n3+QCS4n9mO6C4zr7Go4ViF9EzRDJ5XOzxR12CeGCv4DQcDIP7MwXw8syHt2DDG7Gs/LFfri
4goAlAKz8v860CU2qi2xvkPRZn6uxAd49M1s5TU2U9KYW9GDdCQ5ByT9igtBOBKqfcvROSEYiedd
P9XZ3NqnE61y+kRBIuBetjheyIJBk69He9FJdTE1ZNOX2yeoJAs6vvrBO2aZk1suB8F2FNW9PH9W
2lLY0PJVUjiQz47mgXwDkP8y0Tvt+eNf5OBUEq872qjc9bGf2dxa9AGCIJeyWvQslGIiDGCu3+oe
IQNxMLRDLGs018yu1ldCMbEudBaesZPjV5XmdXr+rU6Mn5a9rII/8K+o1ko9M1kHgVLL6OcuQJGk
Tv6weJYCJoSPFJn9gyLw9YQWGP80ibEDUqa7lCSSwgu1jU79paHBf+PTKKTCJ7nUwwuLIETlUi2U
lJhKMuaxj3y2BcASOqo990pt7oGr0DadCRyf3ySnJSk6zKKO/Y3rV1eG3jZQKacd1ElXTV8Pjd/Q
TeVce2o5G5m7dwT3L4gR3TGIVc/Aefq4roBIaURTJcLK/UA4H1vJkHBcNd5ZJOXFGhHGCyg4HG15
I+8+5BcQWhkKb3fy2gC1kxAIERAt6uFllEjTbMvxIADK5mfQemS3fYmHJ7c00GFdugTo8SLSciKy
W6XBqMQfZgMRyRN8zw3mT8YPRrJwEJk5izzkrNTEIy1ljt7etg5BGtrIGYRRoMckekLMWK/aWF/N
YWQkMBpqZ37iY33B/iq85Mjnr59Ivx9FvuCXDc1jp2KSht2ycqsgUGYENxe2iYHPXlOJGMRrAoAZ
fHRzHSUEZK8E/nKtE+EkPyPqvUDm0mKUp45kAqN93mEZOkxNx6zpZhXciR2FOcXkq9cQKo2CXNJJ
vWUhscR6vgXF0AU6u15H0D1jViqIOpVfDpKoE6kaaXA0CkmG6wR0WoghlMOa+YHxwcHcgNatPnQ+
mUtTanhsuMIY43nZpXcd1V4UTLe+KzIQ+fOW/0QpAbit989S/X/aSxXY4F+Sa5368aUOP+4bpUVW
slZyDNpIJzLQN1vHlRYS5EOZJQQZC87feYU+5UQqghut4DMATxb8q+gwAViz/62FR4NwOyq1HmU0
XFyYx+ouj3qq6gEt5CIqb4a811DdeHPieDwBlOemnyQf35vTEi4HYIAovCnz1zpH1i3AhKyvmnhn
hP8CHISJwkZ1qXN0nHI434HGtYuyUn+Zm9XEoafTwQN2WYMsNw7l2rGzPlZVCeHq4xNTX0lBvr5t
woQbKq4tknh6s3IU4ABzHngpxZVvuZvwSeo6faU2PSXXJkIkdhr8fLjKF12Y1UZdQfvuR1geo1XF
RMDAtr4ii7KU2tcR/vOcZ6cNX4qMyJ6/s2goWlxgteVDTLddKOdcTaD/5Y4X9KiGsQ/JlmBB9NFR
bU82c5V3DbhewLCNJNfdS4ay48iva5NSE+ubt+6K1xfiXtCsiCT8U4nXoFsH9A8zku+5bJKbljEQ
st2OcBFzW+7DjpqcX1Xs5VWLEhpJnlSQs89SXwwonN45UHg8/456AJTXgT95VXwnqx+AtGcS/MSo
AHJQ2CQPIo/eEmDCH2lUiloY1xO+vlbZAtbViKkQjCA552LA7RDEoP90gDhxdoLaiblzg7CmMlaI
pMmxJYo3u7WnCrRn4bAGa9myxfTEQnbJBpgHQnpmzyArNqsWJEc2wb25EQdf5995KSxvrILNP5WZ
SZwTQWWHbfUgJ4FD/RvV1h6TiTWeVPl6fos5BKbfy3xp1UwZd9OViZch7kIOC7COmblBYpKPb+bE
nvXCJrq4wXnbydv4ZCdHRJ70/c8g75xhwfJas3Y4gzuCBSC7aKRv3CH1f7juf2KNh8vZ7zj2p9EH
ymgSP1A7Q2bdFLg4O3o5YZsOh0M57UkjMxnNt4CF5dIObM5N1r9o/RMv1Hzh4PvxIMPNvtcxrW59
xtMhs+AGzyhBL/Rn677ySRuOOVODU2v+mqUIGuZToR+3ozL26RE2NsAF9Dd2bCabob1ye8HoPRQF
zalwDWGrBJ9+XFp0Ni4n7gWZqLW+gfRabVTdeicFwI9cyLzoSz4v86AFNnIlByi65gkbEMKcSg04
FWubxnmIRnJmF/wldOq+WoenPjL63ueE6+sqF6bLXoXd5NtRp52mV0pIrPw0GH0h+3w5aMwPWNXT
wEQLlOlG8jruo4az6OB+thblZi+xpDuFzI49oNym0DT+76hYIhlsQTOX/treA5LmkxkWuKlCSJ1J
BeplfvZhsLAkBPxp8fUculm66fG9eAIoofot/FEVtQmrWH4JeXaiHgXlQjEJ2SqKxMU39D2oP9md
3X732VW9staenLBS0RTdL7aHiCR+MhOjIFiLiLR4B4jBWp86LUCwb9l6Qb+ik/amlNN8l9DyKINb
taw6EF3LWNTIJVmgI7GeSlqBu/6wt29oVjuRcJGcdzKBIFxeLNk2KxnhGOFwRmZY23fskTancziy
dKbjHjjOzEQFJDQbceHjjUa2VE1yE1ZX3PWE+hGaQvwAwc0D1JhbckoskSuPRoaWheYK8juGL5eY
s+1ve1UBe+wbfdeLH/fQu3iZlzzAtZc8c98oYsiI8tSJlkB9wn5Ko/7/jjOF5hNbcmvoD8xfUkwW
Fitc/mP58BqaLUP2DBLJpBKSIlRsgU2HnZnmp/hn+kwRiezbbPvNlvvHeqiMVxV2RPOIQJ8lDohH
+FPkynh4hoV/phnNfi5I4GW3Rtgy7hvpSNobNNWQcizxhwfgGxLG6EoZZqgbxgYouUCdJRuWUPPe
26yC8M/JXA8ig429QxMEKsZw5SeFiKqvJAW0ByocDop4a49paPZH6ED7AIm3gB92RgCiswUQyLkC
b0ZebhrEgD9ZX6aNXW2kNFuZ0VfEJmzaltB29yg4pV8IiMGrmBnrUV/U063N8Mbup7MMyyo80mIK
nxi458O4er5LhytwQuxQWBKfgY/HxHMHGw/n+XcsW6/ceCYy2KytTJOr057nWnyBY7RZMu9LnF8N
E4eGelAIj7mfMuDK4ju8Tv11a5OmbnbbOO/XS2I35MOIScvSDW/IzD8cU5JDxbkrMtUP7RjZ7NR8
p2NXzjCrMxcAfWC5tYzyaEF4ZUCPo38E9iymtHYgxyuHx5PO/vURW0ZsOA3Cg1mO0Z5Z8htUlEXm
R3VESvSMVrY0KsB/KddAeLCIGb4OzqgMh0PoeIT8p6G6+NAoHNM4LhtSiIaMQMvcoeQ0DyQZE5X9
LmPn7SVWUoGY3xYJG7q0oeTaW9990Lm7yG6ES9f1CuIP3Bj7dAQ+b0x9+/+4YVKI71WfpQ/0I8aB
EFcZzGD9GZOFR7OXEh9Ie7/viqJenjMLNX8IfSB7FYA+u6sCrlQ4+vow3R0bi39q+48xHb7pB3+0
H1L/ByGBDecbdHLHC4V8K7TxIwlE8cHJMaS9Kja/ZUsu7JLP7LCq+xyg2ynsGw/k+x2oQ0O/N1N/
OdPScujsAUu/63r2g7XSuz2eSnfuW4QFoSj9j4mFs06nvkO+cusbTn0YMDn8kv84xbstBEYkkSX4
Jp7vtUhAWVYJOrLi4dXnBNuMNkgdSWeReARM5AnOBW2xxe+tfmgnamGwhlHWEAqdIg6D5SfibTcS
j2HD3ho90Jk2DCfleIj9ws5vf3C3D6HWRN+ii6kPczeUdYNMjlQ45wuc+LlkqSd1s5ZBIe7nuAV7
Rl0SSiEQNTsa5XDGiR8lXuKyGiRDD5tg2ibvmYMVRprEGCKfYXJ3ZyIdQYSQ7SQ8pJvL6WMbYH/J
+ACRuRSOFL1I5wkaywR3ZT4Sc0GJejWVVOLZfdoLxtuoamvzjIp+Qnn7ZJtrWPSy6GrEF2JDiIf+
NtZz3h/2JOo8J9i0kbm/JdMBjoqjT+ziSlx6tnh2RymkdfVCfrvb9kIhkjQTsZqZ2B3CtYEIxuZx
1MMAj1IhlZ/gxijbwKalI5J6aD0mZaQAX7x1ABijdr3o+McfGU3awkDW1sGlkV6HDnyAPAWCPBUg
bImzbC/7ESSzY4AT7y2DwM/PY+uCJB3E9PKq6As5O5G7Flam2ZTWUkeErqqPjl6U7tXyw4YYBunz
a3RwxxSJlrNDMXdkgow/m8PesI8XxtNOk0mLh+WuLtGNEzlb3Iz1XjfblMNB8oWC53Fnyooho42D
M+cIMc++qWMLs7EdnPzZ6PNfYspSa8FbWP1lrFNmX2lp0LYlpLm133veaTssI4jQ6puFa+3Fe6eL
2yBm9HTPrIHsMrYd6xOhmUqkrQyMW+ry3Cu3TDmPvIhhhwwx7ShaQRHUhqhuhO1bQm+u5N6ALS90
+tB7QDN3f8AX5b4RPmnLKliMIYMO5aPHYyLPTE219wBJDXoiftiMXy1vEFGK8j2uQKLrUI+TvjA3
GdinKP2sRQcrWHb2bYxYDACZ/RddVzZ66QrcH21Z0PD3946ZEmyy/esH8PGMr45iLVU8jkUETd7M
uTPnQH42Xt0yiJeMf9zhyKkBzBF+c+NtaW03FaZ30OjfgaBoED6BlanpvSEoxXuRZzjFcz43Sx6e
Zet1q4yMKkmK7N8B/Oens0VzqukwvoZs3gQdsV3NMVeyS2zqeCiEFChvGr6xVuSOHlE3fbWcd/W7
leP148VRCAHGFsZN+j7oIeorCkrGFwVuvauyC5bSnfJzQVnVcMW6IQg++LEmaBoFXK+u0WhEBvD5
vHpoeUVFany94NfAs0iwDB8oWR7+Eaf08Q3nSIgxJdeZwTuKfNiEaiecUIQ+u5eXB+hZZDZTTyAD
GEu70kGcadBSJRqdHJu9IrybRoDsxKdToYSDrPXO8rmXiXiXwL1EprBwPvVfio74UWb1qdqX8BJd
6ajuEjFKhdmFetdTqOBWrK8taAMmI9syqPkex3Kz0i6SOGA6PJVbk6MDWeGK4XCCIVLEgPJftrrz
ltjA5naHEAiD+56w/cgw97CHFdtz3z/E64c3i67A1fxVCdTKOMH3DmR7qpnuQYBRxjTcO+OuEtKF
Dy7xW2rsFsF2WGhOwDvY0yrbnBI3DgqpNwg88CECKrFZ/Mw1FG7bK1VKZxgyvuGYcMRnu1mT8Ln9
4nBtsDnw1G47Cu0W0r1WPeAeLv2DQVidB5hFO5fofu8uS7PfR+ewBLw6GxWy7iUv0InVD7ANREjL
bOPUgSbD2w0rI9i9tuktehBw8IKd5VF9zOUNNn4AjYZGoSnv8ujhnjlghxL2RbrYoMVgKz/7qN36
zU3XekPtFkW/kj0Hb2kmQMv//NE+yT91L+448lquqCA0oYe7daC7uCeKfOzirQo/httBDtmMnlaZ
VdleGp0Ec8DpwdSDROkApxEmQ7jN7gSw8MST94d9AEeJslIh+kMo/ZpmvbVUrFAo2nJd2pR02cAE
4R46KfBP2Oqizxd+0lo0nFr6d7y/ep75wwiYkSJiJ9SnXPYLsZVXk+/sy2JI/t+WqabltVNoGHg7
ztt+E5fJDIRu5XI6J1eFHqcZ2vusKB5yxpQmmDFDMI0GljMMlB3JyFapvvNkveT/fe8HQJoYS4pW
C7GO97pDeEjKPgNie2ONd19NZEVogyQDvH8waPIPhYjkE6nGlFbJvPGN/DyNEW56758MXQJ64WNq
wDvswtbvcayM89IWbKlwuMAMh3ycyHAfNmzScAGmwW4MTGKxJb1mgdlSJMgmTwt99Hu5TDx5qMKY
iPkNgredCldV6VOSTkuyAD6Nutz0IG9hy7iWcwm7b0nycmGmLqiI2aNhGcBqyHZ39Jx+g8nHCdFE
+EtHTw2HqBI6b2NfkgC1VNnP3WYCVo8gTiU6nqvUY7L0KEK0fdGCZPznu6AbLLzdoY2vPUXkuK3K
OCoK+weXEGRR3MHFPBkSugQFCk/qd9jRUKFxblLbs/5U6tXxC6sAuCvPdbz2gfrR/VrMEFTLHGJ6
dfnHkEb7Un39hfUhaYeI5MojutJqx1ONHqbxdFvd/73Y0MfhoRSRBsU4f3CZYIvG1mCxr3qeo6++
j26swTgsh9Zs+Mv0GFEoZZo4gv8rR/lVMuqdy+A48OVVBm7yVbD9ajcaFznfWmSagiZjoFbGKIrC
P9K7+icvQx/WzDOiuXVora6FEx5c//sW6w2UmpEEJb2ATKM5sX9/PbuMHfWa9IdHK5sXZxOXOJfE
5Mp4D/im6d62wMGlgzFvDpyebgF1zp3AQEFNNzscwL/gTG+HLUYDUD2m9I3kKj19bqaN39UE6Tbv
IO/USj759SIq1NDpqAN/RxlZwdw4x7hMka7lZLsqVGlBAW1uV9WJ7iQoZmGK9GLRjGaOkRIJxM/W
/lGhLMgtoaQGQcURdbgHhvWBeMYapO4B7XOU6usG6Y3wZ669bDFyVDSZprw5Prowkp2Gyy8ahBQU
m2XzHVInuexz+l2f6fz4E/C+/PkTLX/641VjwGn29Ke7PgoGR1mRasAMrBSpD+I/ujOvG7b3ExUt
AVAE26SV3NjeUzO14JuBxVfntygY259ZGPep7n1CDhYq4+V9MBlu5U6MREW/yZ2NjjIUSer1QNSN
XvUW03ds0aqgP8IxTG0yVv9OxN8o+8hHC1WeOQA9zd1kRdjXy53lotHitRkPpxyRtF8i0SC12CM+
ae44tCHFugeaoiWwafS0qe3CEL+SvYhUoFUPibp1K55shPfaySqXXn0f9e9oUcHeQ9IXnCuNqnXS
lKKMGBAIebA5u36m/lGmEzQwuX+2w9Raib6zgn6Ur1qL5pXjA/BWegsYbyJrU+ywqRP5m3YCyMa1
VzB1BWRPmrA5PD1FZfB5tvjXECT7RCV8U1eszT8Yv//cUdTQXOoaK9lqaLFqJshZ7xxRgzFfX2uQ
CT4AGRUv4QD9gx0lkrkcwH52YSi+h+WuUIcJpnRjSH61RG0ltCOwdKliC7nQ6ND4dS9pqDJduj/h
GgyK0wY1g3SE6/BXyIIglmQm3KP0BPU20aAX6H64XK+tMeo/p42FPSvrv3sOyTV7bA3KVjBHY2jr
IlBo735/NO61aF4xu/67p+fdyAMmOL9IyyJO6ceBhkuU7CeWpjbV/Ffegs5TXj1pJcBNIKmDyfGC
k1i/TKfdD4i4J9JeR1dYlGxgjpuVf+s8ijGil46h5xYr4DHcAUkD2nLS9xptEd/jCKD9868kNgfP
MoscMQyY6iEx6vDHEYo1pDPXsRkt8l9I1d7xY5IgvjgteqTnv99FyHtLxifSsMR6If4T72wDMJOP
tfqdzgQJPgFEbLFKyEkyONteH61W3jswRsZ+z7bQ5weJNh8f6LnMgVb5HbSA03HuHDfOG2RNmreD
CvgVk2COSlBWhOyeFfb3Yu77GpjyYBR8SyYIBW4lIAhYgUZNWXEkSprMENKzrb2z7LOF7mdcDEDZ
Yvftuyudku14XzvnJi2b3bZsbkzHF+aVEzGP7NeoFbHPOK2UtBFEbxlUIhmvrsPabjhS4B/sqLbt
p1Gb+depfmp6IeX2vueDVXnFD5T5mYkmfRE7lBUV5TGiJFlvQ2SLONt0R39Rnf0M7GFltDoVj3jb
Fq2pzh4AR+VKlSq3q8YJZurIXLDZSomnEcx8bKEQi8Idc2fRbvVfe1EDrFAfHcjZFq+Ixr0elLoA
bCbx40XvYGarT2h4WPhZsdBgMom6wrkGOZe6slGXVWbiK+jqok0tL9jk9QFYVhlVQi7vHGSjUy3K
Wdc50s1sRiEsaMuKLBeSDqM6e5hdcvewCOdiSzr/M83BF4JfNMnM9FWjdLjRQw/W8MDXrtaELrhN
NLa5ZKzYR1+9XAI8vMAUJ9ZoQWMmkjAFsduujJZJl/Xu4qDePLo4ZcIR5+tRRILNnkqfWUzecSaI
IUFl6GZH5MMpNYoGUs7Khk9kLf725+lQUvk1mZJQeQQ7i2PXRotAFay+8eO+pPpJY5BDkHqiUZVe
LbQs8vekYkBG6u8kN3cYUS0zM/msOPDQr5zd4n210p/hOjy/TuyXbl7XKT2Hid2rUUGXAjDvdRHC
6O6NxJXqp8YJ0ukbWpRohsBBPLsSb0W8XMKRGVyfGt6xxm9+aaY5b7ri/3mne3elycKZ+jbdi7H8
wfeMzwzipq4uY6KuMo4wNb26ftOJaBVvWzzeNVyEdSDbvZ1nTPXlZb6mycfh5PdSBGloiuJeLc6l
O/NMVTZhsOpsrFww5LO8J0xVVKXutDhIZBDVGy6ilADw1EwyOqgx9uLUaA3nwUtBQlj2082UobjS
GfmjOSAlDOCbO44F3nTy5MX0G1a5KU8NGTLvRuVkdD/7vf+D3JEsxTaHCvkMlvY191RFKALVp817
+nrff18R0Kb1yCLw7uRku55JMHH4D3gHV3YZq5B9nF9dCRdMlYTOXVv3MpQuAueA2qGxlYV+Hmvg
w63pBKaIcANvrhpa5RrtQaWOoLi9HeRBf1CojtsU86K7Jkg/Q4neUmjthgXTngI7vzRETIR3fpA5
Dz7SXz66lGd5IUeK5QK0zPvgYBMze20krI6sYNiz+QPb5WDHHqSKKUWKrcEqBAgIUU6OwTJWcWH5
ajtrfvKbLzJK9qTdaxX6Py9IjyTTqUc0emqzrvq49ntui/j4mFtHEGku43Lsj+07XlB2o4VnG/il
GVyBtdd1BSAmaj165rdJvU/QeJ0O16IEzuJ67jFTQl3yhHjCd3ulWETli1is8d+92mDc/ExkTA8z
SXbrErcve2TtqCr4DQjmd9TTOs7FkKsGQw4I45ZJVaGtGuvld083LHLPeSl+jdH7ML8LrBqLE9rZ
AVU6GLnvEVwI7YsUDZs/sMvP6wIYECuX/56USbYeCl2CR4FrGJ6mEyqeAERC+Z1thoFCS37TTjWW
zEnbPT8vfRgJj+iFid7L7XQ62azgEf9JonXdFXKoGIrUB4WSTMvJSMraKTGR3YqteG/0x+6+L7uS
07C68ne7D26FCvNBC2J1qBo6UdNn0ENVCgzja+3AmVeo5jua6v/3Kw38LL9IE4Xr8VQR5RX7YTZV
d/suQCcBM5ttgMN7+nePrmwJlOYp6hIvBrrZo5I8eu5sYCWkbuZ75zjUH1hTLVPXmeAV7767n5i/
y0lLWliCRoJo/Tnok0AkO+ndpVSzJvfh6xCUT4i2tjfNnZ12FQgT02FX8wgRs1KBbsV9D0OCMent
Fr9SclHXxSO2nC1j/6GFBSNtIUFBaVXOL7gfe97DoF/SY2SVYxYGLrv1fTvI0jxBG7v4dBcv6/Bf
J1Cn/vNnjoBhjerIHnAWsWQ5STcHX07BCp4KfZR6pWfSfVY4SwlQvJDkqcDTUeu3inEYKlU1ixol
TsT53pDn2jyh+8isEMy+t0+cApH/rgK6hpV8zPBigD3sQyl4eqq4l4SfFC0p5/SQ0znXX0PIXfsm
7ySEKPeBggNa6qry5lPOSP9jbcI2wFskXT15tqfvPmfoHDKDSTY1sXnGUicrwbENGkr1AqWa/H5r
A0eU6SVQNNKWypehIsb+pUo2c6ErweKJVwjzQu4697DKmJ+9NFQaccLjKEbIHq9QIolBdaKuPVru
+z33eu9/6aBuiOi6Bq+488WNnQHGVT2KFdRkdoryJLgW3UASdumTMKPacdZjdtHGWYLhyPlm5Qng
ec92MySrUeKAQtXREVGZVmguoJ1A69EukGR0+EXqmvCoGcy/qFhZGwc8vucwrqKNvjclHURazXrt
KF0Y6EgYxxh8UH2SLttVn+hTu0k1htXDe0R4HK4I0x1ZLcFuCJyo8L1IX5CVX0Takctv1564cMqc
n55L6vHjMfXkOuoLbLV45LHUTVcCix5dzePp3KrNABTRfXtmQ+YNcAddMfTIKDKe6nXJ8fHUA96E
VGzv8j2TeYFBbTPyRePUk32Kp6oK0DN1DiY6OeiLERq4tnamK1dITUe4MAtVUZWTjs5QHxsmjgrt
kRFO8pEfMgK5HQq643YciB9x1CeOmTP9j4nYZn5uYGTjMVb4G9+MDvEu61vqglPbKlXtFDFSrW5t
t/sgvXgtVQIl9SitwLuxgUXZphvyaE2e1DMr56fxG3gd31bov6W1DAJ99cbIRzW4zgVO/i+WIF6x
/fI/zycBSDg75XcdIYnxRHI53GP6E6y8uhCkUaOgNNT7XE1P8wzMHIwhmE6kvNtWNSKIrRT1adN6
0qD+oUcLRoerSC9d25uCRo8T3X1OIrDqB9uJ14vziGxRvPLP9P6pf/cUziK+hpDSWWd0sFrXGk7m
aMF8mRk9NKcXBkiAj5xLBsRIxmNp9Gv5Ocd0q0TqcMjmiKd2J8PG7GiU2aiy4oH82YlF/cnF9dEy
f047z6ibkguBFz1+0mBVl1XYsFmXAg5navIv/qhN0RUVi/izVX+MvGaEOU6bbgTxDIaOxQtT7/20
oPaMlUKl28DWrSGQDHoKiPZCyftP+fUdWLOvpFIq/dtCjbHFNgccv93/r5kCpMheb3sqh/8/trCo
wFEPdzGU7gY+Q2NyUZMVQIfWOAkav+jIDkRweq2cQZ2QKiUmn2SVLqoOrgFZRZa/Lu9ur3YZyMCu
JjFFyFMCvjWdxnqmjNjXu9mWTnusDXvfYBViYeiCI5H7io+q5+flQu0eSEpOEo/nZynSgV81SlFU
Tgk63zkMxkxx9MSpBFWf5teh88FecQlMcQbmiykhv39mRrErVMZSuFC1RlYzZJV2FJCPV4I678RK
Mh9DGlUiUZFd8CjuloYpfgJzv6WjXcUJe4M9mvmEZ3UAgZ80SARfdC1ka9xHUuf+ue6fcSbD987H
ChcPEPLYf1g7RLFtg4/cytC6V7cUe0WaDL5A/0ZbGn0LX012FdlLhISK11zawxfxopED7DKh7fhq
JrM3CaY1P7a8NRN9OWHaRxZ7NpEr6NE6ep9OVRnymrSl39yxmMsnd5ndKbQC+Gya2ICAdglN09qO
/zlrRewl2LAOFMiKUKW7IVCN+Tuynu6i8FMYGUcbtLNGIBcD/KEJIClCQfn7wfBmiUVmYySV0gwJ
ZHVro8sOttYloTJxPBEqGYK3o3N4xzR2Kfsk45wVt8KPZwki2Y9HC70D229xMl0F7MiI9vck8k2R
IetY14ZuOJUyahccoWrOeiR4MiUD4KoWCe5eunhFNHDwhF7jF3WKA5hBm6tVaLP1rWzgYOWD2Uk2
Kz16hlz1s+WYLHM9o3FvIFNVhmfU3YTObUaIEq5E+q6a2a/FrpVF2LEKO1kzXBg5udHiKw6sCvd9
2w9RZfh4dHIMTF2mbW2JF0ldovwikAaeQRBPKM69icbSz7VNcXH5mjWU1OTCVc3r8CtCqWPvM/pN
8jxq6BHIQkmZ3eqa5xJoRnPIedtDDGs+BFPTktaMNramzoOCR2eTwAdZwQDS+Ee0hpCiqhq3wOOi
0KcWkrJhwtVJRwc3kbAQjuktl69dbRx8dMwTU/z4R51izLz99AyNcxMHGWci8d6couvQY8EY89nL
V+cOu9VJx1pY0gT1nHMMqd4GSkyN4/PXjjh872rzOUG5c0FoCy+HzUm8suTNu+Hn7FMgStxAth7d
MJ7mFaZqTepiHsWD5wNw2nNnDzVHGc0igsEpuq+f55UG08a94Ho57uMeIjyOcfiCaKJ52Ffh1yil
yzkPjpLVotqC+dX2TjZcdxxPfx97+aN2yZrPlNbZ/uXPfUPPOcnzB+XgdHwM/Z0PGUk8dmRuFnLH
DDjMW/9Cy+gLWsLaLhHuGU8XiwStiw/WPtq1mVKjZsqpNMErHN1tCHc+s3d4iDXY2sE+COb4+l+R
V+uHdQ0CYkpwqQd52HJkYqO6qMSxzyiyDUVKJsM8fropz5ZD6N8FUjO6yJV9xuFNQxmphG3GgbCs
bX1qXY5fxt9btLP1PRrBxB2+jWfg4G2+0RaTIR0x6ih41gV42nhz2L7+Ti1+O0pOzo7Q2H+JIZ7I
+8OOyzyNRjC6SxL40+cZEvrZHhX9etf+hRrDR89FugRv4oh8tAGbMipCSp0zn6BT9GgM6VX3bRH7
L/epLgqV5jLW/rfPtac65tjcTJS2nj3XX7jqsiauJUHYQE7sCzJSZ64Qep8zlyI6QSrgN7lsUuZf
FgcHSs45r/BeqLY4LA9Jydm+OD7gQmhjiA1XMyBAk+Z12I5npODUU1I86DryddqIpZzSPYSFxLHJ
GZ3N1gr/1/T7vlFvvfzmCL/W7bYkxZm0thiEx+astOlaxFZJZLz1v4lxcJ4YgME3pq8sVtDWOCMg
jJl8NuIcaCUPfxnxdmNF/HCgqwUAuI6wi7JHwxxzR+hFy3SoR5KKRKcaQt14UpuPLcDxKTZ/zsZx
zYLo1KjmQSE4FBu+oswcEjIMxC/5rXvWKMCal5+CVFcs3DOZ2qg7Nd4q9rhAn+2qSAo5Dp1Rtmu9
jU3pFB4JhMu7vUV7N0sHvQP6jVFnDkXZcMqsJC73wXoNrWO1lL+CiMZNsqga5Ey02wVUx/416FfN
g20ywsC9aIbkqwbSYWTSwJPQDxB6kjbc2GwGryBzAYw2wXC2DPOFbmBjUgpVSGETki24nZhMWKvA
egrjFHsfLkiUgrdgVCVDBp/dFr8mFSTjf3MwFScx94FxFdpiy1/p3NrP/zVBLkRBqgsVqqxb73xG
iFiLPb/kTWirFiGxrVwzffgV0jftQGp+Pi8AG3LJSjrLiKVOilXloRjjnhemj6WjhqWZD7UrUyGu
CSMzFv6KeG6VPX/foXyy7yBTfUSjL55GEnRwDdQQOj364uEi/66qpQfjDwnSXwIHRY0mu3/9+ZAZ
wISfO0gMAzSvWXA9CQLl6HZcTqubbfO3ksdv1dKshD0g46QjkwZOqYh7kBRVzKzeQYjdkp1o/YvO
bGUX2SUFD0SpfzPWmt9Lk5IZHpO0UgBfDVv01mUkqF77lM8bfIKjLMryjACq9LawqUoo6SE4HHuu
Q403yVhVVCcvDblEjPxw6jwHB+j7aDXcG+Q2eHFjaPJkzK/s/X3QaPl4yRgnHZYJMG0GqL2Ddc+/
RbccP8X5AYHX5TuvfPuGJtvxyutXcjwgA0INGBgKLS1sf86tb12103ZYPHk5SexhStu0PsKszgEX
lMvNU6J61TOYSCWE2oY0yC5Mxoahc4VsG9eyQmyK7NcNk21YaLZ/AAb7kQqqLvSYIDrbGUe6KVE1
2GmsLNdeVW3dMJp9kFcM6BWLQ9ilGw0Kcg8HmEuHmwLJsFjIkzmUle5p6WYEH/KNWYUc5oKPmKHu
653Y+sFUvT5dPtU+SRjPxR8d/ZWZgYGsRejNipz/Hx6K4eAAw5DcFi8T+JVtXMvQQQQZTPHHRega
uKHn/TjWzd10/5WAV/4uNvTkwB+6Cg0+IJsXU+CsRRXACRi5+SudF2C1J+59aQFzP0Ej5U8z3Zq6
7m5/OAscQ+7RilT/RHST0xRXbMTHH+syM4l7sgD1etiB1LWEj6MgAPfb35eQ+qxlieDlRGEUFbhq
m7IRHpLN34ONXS3moAnRKTA1Tm+hTpBiPfRbCRao2Dd5dHAizjFHukjQxf66H4+qEl0ycHXBXU5T
O7Q2+uoxkkvK36tsUI0P6R2b8S/jT71Uk18/8HmvfL8cocdFkGWTQfez9rpEY05th/Z4TIDWjGIT
5dIO+oczst9T8QogE8JNEgBWSjZ1+FIddBTMwZUrg0VrQ+8pwmoQ5ptHqrlMYVMibVaqHGej28lP
2dGLN6vLASJzP3yv2jYeFqgkNEfr2AfOS4QYNfVAcolsgRJW4fVrFuoj4bh7YeTkaIeEejpl/Ull
N+kmrQkx91+lETCt5bqdVp8Ra94ZRHrn1nmBz4NpWWw7hpzyC+0O11q5qrtqcpsFMESbSH+hsVOW
W9vHqTh/UT9azBWQKjzOEYg7wGvESH3lLWM20i5X4UjCyodXvt8LhZeXJOrhXSRKFvvqT5YLtOMK
KxbyZgrjBu2j9mGVwu75CSFUF84NYzWN8V5sT2AFuq9tl6y1TI0GOgIlX5i27dW3Vb3LLyrRG/PS
iaGF9gDUdeU3D6bMXni8wO10oZSJexqCM+ds5nMLpWfSQOgJF8Kgy7++Y1Scx922A9rL1di8eVR2
AhfhgeeZ2ZuZDldpnBqMFHUoJtuimBxfkgV/5VUrdq9lvqlfheZPnYKvX3P5z2Q7JKKFPtI7t6/0
vEmPJNQ6/jQgKF6I5818P49D/5YrquAZVqdEyw3qdOXVrf83fZhtJAGTbC2kTX0faNC8G9V+50lU
AR60gSwVIu2N/5Tnbp0qTB1HJ6Q6dQPsq+GbEtrAZAX6o++GNyzpiGTik0JAa00LTDj/my2ceDHc
whwp0iJjuKZkwrdCgJ5jY9GEfBe4oBb44TKPGdoPwzM61DL52IEElt6IKFkp4dpO9S7DISlOsi7e
9k/Obol6C9YWzoirpqbBrwCpXeoRjzOW/+X36zVDHt0yJFi9vP6Sk+F/77/bH8I+lKhIQNhDlmh9
1jfGvUZ0tQgSC/LjeD7ICgSoGSNynreA04qKNN8/2BLrbbKA1x7twqgwsw8YBbdyCodXN+tHreh7
z2F+/W3v3/j8vGgyW6J+c0AFD83xS2HCRpSbT0M/noTp4c4jma85RItUHT/89pNqo9EznY7laXeW
yXuHLJUdmO0ONFZW862yAD8WLAOIFpk5YNP8FebufF6/002UxAQ1lYoGBDZrgu93nXrqlsDB8M5g
IGvvqhrlmJap1iBBUcwQlJL3kirqSPTe+B/WvhVixLrNVN5xLGOd1OS3RUsXoKuoy7DU2c3WMY5O
sreO+IjIT1ve5jaxST8/UKGMbw75WWXEz7o8+r84rdedbV2h3dLQyktyZKbf7niv2GeZhlgMyE3V
dFQDptafQNMC+EHKO/5MQrrg6hc72UTYxds38SOtCubfL5ZTxDKBw8fNMefwOnj4F3sApzLZd3pW
bvEbe4skSYhwudzEqXtY2JlTUcQXvQ9JMZLJ9/rKAZPQ7ih1km5CDnixV8aEwMKYWn0JDhHwJTsc
q6/AT8XllUhJPVdrwTg65C/4K3BoLDUhr5strtC2kQ/xz+N3Xv8J3uCLXI361LiiSN1neT3xYxxT
iF6JjquzxV91PcFae9TzCUMUFlAtoEY2O3J4OMquyCxk7qkkCZBeBbXtUac/Mmq+hmnCEtbzoU4F
Sf7Uj9r8J1cfp7SHKg0K++KyqI+2PqTE6AssB+I/06mPC0bgYWmx9EYG2pKeuOU78w6ylK8PcNAL
p8InEnYvs6r4NY2lofkMaPSNsnEAXyZ0QpS3OUDSN4k0qdc6zHGRVDpu5E84U5w69tOxp3YjJEZq
OpaK1HfqpmKg4pqHt4RG1l2E/dNu3X0rsPLN7EoEIwBpqStT0GMOKDDbruxUQaN7gyXeUhViTLlx
P05L2dWF4U62ZDpal1zI130puF8LXDlg5bC8t7XiI2q+Rn8h/Rmw+ka6jdjfFFlWzFw7IbTirwm5
3uuXFWgKsye04VIxMNnaH+Qpb4slWz40FiAeVkw3XCG5UlySCjvcUk1oSxcncQjfZByS/bwXg9gL
GibOM39AIcvcCEcIS0W86lrpsBhkmxLn/WM1gBuZKLInZZ2eRb4Z2sh9DRtfeomjthNU9BWEK/Ry
95CtWLQzGKhPDW5alhPA0EyrKjQ+ge0dJNBXdQohUW+f6P0UDLiaNk/8CeRB+0f1HhVFjIBUom80
zF1CaLlricqtadaplepvC06zh4vMQibZpxdgoRaeEtyxJuls6ptDUzdqwleIlIdbRLVV9kmVjZiG
VofAb1VVfAtP/PZjp2R6IZEhkqHOpxMr74NGvbOsbii7+M18XfsFThr/Ru4vLpKRVagDQrwa+HhK
t4z8uBBdjxryBiMQgAx+0xgpHLTJQ0YkY2ISPdDqGeZ9JdcbwzJbXE8nlgg+6rxkicVNzWY0oGdp
3jF1VoEN2KC5ZFoSMeifM7+kJNDETMN8dY1Pu33NqA/F61ZvwAtVnn1dJzufbX7Dim1mM39dU5kO
aXxeFvtV7AzIOJdermqtpGsDxAu7ZHaZIrhnxPGIQ5lppdG4n9okJpNRlC2BGDUMK0NEIaTbeIKQ
0kE6lZYll+2JmuQHA7ppZ/s8/ky9B6Y4k4zhNvqpxsz5D2/ZFxkmQCOEEeYBOnQdykq+TwLv+PQu
ov0lnFQaySuwORgZypLfADBs2pyW43RCjYMKf5TTkF9wJgFsf6Zdmlv2FLDgxeax5JCQLDBzrpaU
dEwXQ6W4c0lN+Y14GLhMPi4/pJSnPruWs7HH2T7KJE+57w0P6m+bOu4kRuo7+kyw08WPVSCQmyxt
BGJmwcE6T5kx9f+HHMwJaDy96W9FAtYaQV8Fth4SzFfu/zc5h29lCT5bhj1JmYLYrxgp7V628Rm9
O94rWdWocD4ZpyMXwJ140pAmZK6Sj1IRNqX8+xg1kFZm6j0WqiWixMWdwuSrU6o/e1DG7tOHZ3/b
yHvA80kIAXIkpbFchkczqmVCu0Mv7XNMrBa4azMYZnLY6SgaT74OAlypPAcG3y3oej7NcnDf5SNn
W37kCAU+KzMl6mZDHMGjvXAqj7e5kSSafJ+S7Laxa8QyVOX9C4MdvjMUsetoIR+JcG3nMMiiTHRW
PjgKFAZufOeiWw+a9XsasrMHrJCp1JK5Z4Rscmjh9MbFEKLYdTWV4x5kutFWiHoOVjGWt64INqVY
T2lG442NhAmY0J5wdrrgBSVLhWQfn9iUEJD09KmMBlkmGH25CNbJLDTFcPD3UEvquGbIwDbWp+bi
uGcs5E5wQ3HW+mQasZNhIBfvPbpQYb+A5z3Al+IFBZwaRuucH3l7PmYT8bvXdvXv4TLZVuMaViHG
OFm5JBbVJIYVptdEvj4ooUysviR87gdAVNCdjjAsqJiqnJR6Hx6WXFT0PuoWPdnUG/JiDUNZNDkI
PjaVseJ7SQi7bIPP7S+hhEe6jqI7p/NxvwhqSN2CUM1e+bEBQD1l6EQmNWmHd8KI6LKzWzwFYI7s
0ckTetuS4vU7v8SALQp+MVS6IToKwZUkgVvV/cBewLF8xYSGVF14syu5MWzR7i7CYdvFHT1uGt2T
3yKjFfPTMbEGj//ywnQWSkyjalZIRtPUmVHgalmLhB37qYiVR5CLqn2YplE3enoN5Jt3XjLXzas8
Xgf5DSWuxTlpi2H8gVtFLsnczlUvtzpSnxzjGshwnsH7IiMgR2+06QyubSbA2V5JHBl7gwAu5WA4
CU6Ees0QDcQGX5bD3aN9pU92evN8h0/OOjc+LlIx5PZVAeFTjHuIq7dfYCJCnkhH9zf05NqV1Kdi
eOvV/5X49FO7omi/SmsofBV01BtN9YTlZYy9D5g9qxLkn5ph+NDZHcR/GmpBo1zXDIMCYMUSpffE
h1TDtM4jZyU2VBFlX2drELE1ZilZAm41twmTV1WYNXiJb2LnOFuZJzh1aSyDCi5SZHrsf1IzTMSL
ORBUUAx0aGrV5tVK/VSpa9a3QmXamE0fpvUcuzegNdNB8/divCNqi1rkLrcJmrJN2u6+Z8uDwGWV
/bJcRtxdJgYs+EZZY7gyqY4q4btmL9JUQcT8LweMiuYbLYyAB2f53ScN+3ahdZsjHC0kwPxsdsTo
c48/w/vQuj9fJIro2k8jqPGbOFg1BA8ExrTxEDfvt/ejdSkJ2x/vpcxgSAnJLOSQHKTqkL89UYc6
ucbZfkFOj4OCGNv+nYEGRSmMsV0GgDKM5W85SL7tfUN/IDhp2KuwLKrdPbUjbRVl3UauPSvNeFJL
hF7mUFLDbBcDff+YIY/3kaM8dllV7t8T972XTTrEokZGkcEe94jQB/LJEa/Qvf2WfKhyN0p4NwlO
8NThCBZzzo+j21RWQUnHaO6WqkLrh1s9RJjiiMQ0K8UTJ53gbAA+W1wz09xJvn7LaWxqSqc3u1GE
Q8A5BDcvXzWw59hBBUjOS+kjNgE2UqDmK+AnH309Opp9YHnuQ46cnLBT89XACVMnh/bCmCfX8C7L
Hkc3/L4ayOHibt0e13JxAT12/I8dTQRgWXT8Nszp3Sf8WvvOBlvmwVOb61I9gHrnWJo397BJ8vxQ
KMHaZWO+FrBPB2kByZPluUOv2/c5o+iX1y6TVyC3K6vbJiy1lNuq53SATP28XUvKLVK3VB8IEaQx
wtmidmrUlPx6qzndm0YDp4uFh+8nV7n96OhutCTzEfqfR064xesXDBq+wEi3A3QdbEGZWnPIuesi
8l9nKiQ864Nt46P0e9lwJ0qcCvBcofx0YBMopZekafQeknnHExRrFHnYofBnDcXjiwhN9fphN6YP
hrFwt3NBY1CgLtWntvOxajxBiO9x4A3ZS3KSmOmVfXOxJbkjMz6DHIziKTS4uoG3yR66IJpui8a/
An/mkC+agq7AxeAet/G1BUIZtFI26S5KpMlem/AYyZELYVFu3sjxPRuSDYtz15z+3OkfKBkhH5sN
4/QvUm97yjOD70RoRGi56dLvJB8fKoTilU10XDbRNtrsEiVfWm6bkuW+MEuNNkjQ+EHhpBAMs0oz
gLJCgDovdSyDRj0IR8L5N3ExAfCJxBZ1RBqyBNeRZb7Ymwj3U7rPz4sZHTiGXmnpAiAepLRuBIbH
+KBMy4EXHvPa4jUYbxCBH7fWTaBcOcM1h8/nZ9W1mADGrmsb/DizU16KcJqhu+I//98h01p/OznY
BtClduuhEXRG/OfErkrEkO9kMmHZIqFz8sLh0S3ynzpaQYN7B9uZZcQ8lw5jJNNtc0e0BZI+9Yto
HNwNCZ62NyA8SgFaSvJkUlHIYfgw+KNmtC/LB9DpLM/sX98OPdC/JHym3HvwIA8Ffa7VlnGYtKqe
PZQoSBrvopGWXdE5FpCUGeD/wjtXws419zCAVZAzKzeHGhMyBSFwYmHiH72YQ/PMsHE5bDMbpBZN
l71SnhpojOM7hosrjePtu3h+xJI34XHHJArkDUbScQKSoLNtBPijfSSxHhhwA9c8Tj1EWB1LLGA/
+dbVZIuDcBKDdmbFWOI7wCj/cR6V86pBle8B9tOUK85tiZoOHnePBZIDoYG355JumrHtNeEPdBn6
7V3tAAQffBtIGnnONoO6Xu6yzNEU7rvgycyURlPRxv2K0hZh0W8ev388aeX+Vwu29l7xqyq7iSRS
TuuimXApaXmMFJ28x2n4XRG9HrNxfWM0wUsjKQaH0ZOQG4TMlednX7g34UzaeRKahqbxiNy4wVP1
BUT8s38rk53hxtR+F3jpWGWeOgIMKP4UbMSVQYDKG5854Bccf7mDJnqa6fC7bX2jx6CSoy/ROqf9
VJ3QaJwS7wb9nwRrzmaK0lXysDtphPzkQsjRc8dkoizqd+JcLmDAye7CZWgGM/zKLW0mak6XGqmt
gCr8j1rlWPp4WlBK9RPOcPFNf6T2gZpzOTVAW7ADEL61uUs025UZLNzUtb7jPcoie4rXG9JpjzSx
H06GTE6Q2i44UDdf8Gi5hga34mR7afAKnf+z39/rbJvyV6E36tmtFkPElSTg8BDsl4QAw+mGxw+p
+HZeFNmp3htotoPFjxAdihkVPJccsh0MTglrgBXEOU0Xi6D3sFPrwEm9Q9tyL0X35bCvOT7KVPdg
2qEhZk/9U9ayUsuekMAzGKZvb7Sik0+e6UUgiThYpBK8eyOaItlApKv/xUvFnL+U2zyjjV/QElw6
MvVAe/VC5C3myAODQ6nMfHZaz8i99jH8QC+b/DW3QlV0ZO1sVuX9WdPuUGze8mPaxHC90qIulT0m
W1WRYimsxIX6WZwYxQQwxAKkBgL2qv7N2neMvRyrjJzXNcjdN3AYhuesBuJt+xDeR7IqUUSAC+Oz
gbllp8wmY2nrJL1iJC9QwGgZyeXyIACY0ouXrtseGA40a5cPlnogSKm/HjS1qGaCgSlH/r9jU4Cc
zKXeh5beEMM+y5/FlGrg6RJjkoKJScRgZ6hf+fs87Ug4n5PvgQdkVwinSskxww0O7pMoV7G5BAP1
zFpem2RuaeSt+4BSb3fGpqmcexLaJQgvklaZqJowAPXpw9ZNqjq9o/xv2q6W416s4JjqSkxJxCFR
JDZiqnU5HjskdvSAn/+qZgKLHtsuog36TntOAEo2GcDCe/i+TZIJYIPs0B98qOA5VB8BDRY80sTX
mG0bkNRXYBjkYdu/a+B4EeVHIceLDp3WTAPIMimvVDK/TY7ga/JNhSXtWVcCQxJt5pyLzQiOPCc/
33/Jo2Qf/laV6y25yTpBq4S3IuX31UNft95m/aIQIcZ2cZx++obNgXDwwi6eIyCS6pach6WXtFWC
9ux100HaI3LGNqyd63tPaMIcviCFoSQhiXb/g81tZAA+wC1w54PNfqTGo24aO4k+ZCkW7bC6ewRI
UXR6KaIbQ6DQBs7ogt/zvGN2oYCrAP9swKnIFpOj0FvpD7YtbETtz8Mf41iUb9meRHh7tLelSE3w
CRK2usIjnwqyKbwe2+Wxz0czTqoHHa6W//PYwfi+6vAliKEoj88/ikSJ9SR+qOzVcMe+Dbfb5OPm
H9Folru2wXViJ8guC+f7jH6V0tfVT0OlJKV1sVDleXoZaokSrZkkwg9Gxw4Xlb9MCJSFZyP7JHnu
MnBdHDpSGJQgiZ1Yzg8dDMbv3kRFntOkgFKgWMFtyo976UFjGOCJ/8LCijf99GuzS1WmOFskn56n
IBmraKmtvjzPdlXEvUjXdMXD5I3TBr0vG7aoHG+OaptWn6GBI8T4vxjGRPhCFt+IC60LNkSBEwVE
27tpdIT1VXvUzvFgdnMzYXVyHkRVbKiBBuqk1HnDmiCSU6QKFBdVFlz/h6NNfQNnkcmoBm70Ixjs
ITzJKiDL87RGoXvtdJOAIRxDVn+iC174kzct95GbmbhbTTaeUU2nKiH0caREe/8b6ZP7EIspeAAM
5T+xsJreJo3y9zmaZvU02CRBxUzJtx41JsMYJ38+rAHWGvZOqXYIyxUFfDwDjN4SeSMiHuAtJjQF
dx42KBWjdYViiUV9YQUY6kY8kDsxW12fNJ4F+skbiRyAEuuRB6wlDtwz5A2B+71y7WJaWVumE9aG
qpBTdn7R8uik6JpLshpDU7F9gTW0ZeWe40wOmC/xypOiJO3FBfhx3nbyeWHCTw57SMOiLIZ+gjwP
aBK6foiwUQluDSA4cjLtstfxQ52SULsx7aVRHhNMyzROZz0eHhPJ9iSqXBgjf7Db61OgAoeQ9/5k
TbZTSnSHnn+UxgGlgO9gZdlQ/5Qa6uXvYOKbmxD7F7sj+Dq4wwN1vSgA2AO6in673E8vIuHbQwLj
VXgiROh9MWQNOl0WqxWflQoNqnEVXdGy2nZn+UH+WQ16RZIe+O69PoezpJKKeCBH1A5+KvMpASiX
UWGu2AjpXY4Q7oNwi8SZqsznjynxkqqPSFg8+lkokL01i7fYgoe4nhavAZilYSY9LuT1mzyHjZ7z
O6NIuNRoI+hSlEca+iXRgIasraofJHvjXzW56miEIcR6wF+42mszmyS8DPRt2yYmRnSGnINfor2x
uLSVd9pD0PTuC5sI+paiYtHUxnpnsp7d0Un6DXH3V8CV+uAiOm4dE8XXG7FPuuFzzXc61gNyIwOy
d8kguXfOLjFVbSNhoI9ZbsZgIeOKMOFUUa/jQ2R//l9ae9rkC6gEq5nMF7cXi03ixDNPVYqkM+8V
PryOVpaTCz9uFz8EdwOuPRu1FUpOPip+PgLvddqNQEGhIimSKAVjOcxPRMQRo3hAIgIjywwIp1sE
0b+OmkSZcicPbqhiiyuUMX5E+RLkiACjKJgfdQXuSXQASXp3LmyGQbKtwZzImLZmwGafrmf5U2XC
6hAGffrpfy9lSKFbuDtBL34msUtFyixhg0gl1cOUq3ySl9tr699MLB8Fso6A6LZp0PmW9tiaacv2
VrXlMUkavNSM5ZUW3PL5WoHXtDi6eC8W5g//g/brrSeUACaVsIkD5GhdZag8MfFvZVaZNrGfFuW9
cZgbPKOO5rkd+P5KejJOzpfctWLzhmGWEgLftbf27blxOMzAYUJ+7E43Jw9iEWApfxfXZEeR1DAS
f7AzTVshrQ9Eesw1hCZXbrG3gaKJUONKIPmTH17cYECKGojpwOi/LVAr7AgH2+e2NMwHA4VC3i/A
imfgPXRKcc+RhseXs3SUFPBUypvSAatftpjXfddTRhf9JmzHOzVJrzZF+NFqd2B5XLStwOd9BNK8
Z1r//hF+o61Az0Wu7B1ZvaBQJJXEnP4zJyuJOn7awodXqyeGMWvql4W/222HrhmX2HY7ZSvLEZMy
nzHbeOyrBzzhXIbasgRO56+E8s8/n/Fhm+RfEttbIFct6gNQD6A44n9O0JaO4GifBje6+eIwXJGT
YqzyBu76y13hr8sYgYheJBIzfL+419GPM6Nn86fl9JN08KIKnlFRKjjQ5sM3K4pU9fmKxVFYQocR
RPXhNl7k12b7qXaeO9QyPlFilg1UfjpkjRnx6iJUzJFirpqeTigem4T0rm9JSsD2FfVnZg1F4iv0
v4dBFARAcxKFhe4mtL0inhwnOtpnrlnpGO/ZVlTUdjhUCdFBwUZYEBY0mx+jnnUIY/c43sOaW2+u
SGm2RHHZLf/p4E8/Kaz6opyF5Z4kRWEmYm3cswXrOdc/+lWfa1lXU7jtE3m0vojDvsRbL0M3oWXf
IcdIMklHRLZ3SZhRC4o8N+hLmcz1qUFomPkWOpayia/GisCMh6poQoT5JBNxCpKf7fVX5Xnbet5g
qaeAdaoNgNWUgsDxsrYmKnpXI1m1CEH52cuTw2bOlgeERFJpxt6THtxilronstmFdiZzJk+Nr/uz
qyeKS1dYNCTBiZ7V5HKznYzLiGAKaI2tVVrkRcntxCrBtbJrAqtSWdNMUjJ6A4fzyPSx65h2zMz9
Y0w1J3otoHMxY23CnEZqEPv+R3XwB9fGycZAIAxSkVJEOT8bk2TkOc57bv9dDtHvllfJytNE/QGA
K9aB4Uo/RwjgY3TxxrYD0dWEh+5cWQ8nfl6B7+47HyST5Bd+nACBOk8uY2KDRIh90OOfmLpZuMJk
/OMXxZ+Cc0eNsvYsJWrTGzncKXaSCxAxvpElXiyMwTqUFQIa6nSUNfNynhA6v8D3UhoP6hiWI6QO
ZkYlGTazLzgWPkQyw4bMZZVi3zASMPSyOVW+mnehBwjwLxFoyKvHoGIEvD2cogsdBEFh5e+8D+3u
z6q3K2lzmXrhXkMSfa93NiLTbqYU8/3jZOMXPsrLYsV8UZqEikDKmlQ+h3YbciNaBdQ8//YgIEqT
pxwD85ZA0OwBLVepZoQiesGU8zGtrGurptMP2gQRCZCgv7HMb9IoWSH+9VvgELCLzrmds7uWPt+A
F0iLimXfQnd0PP2T6V5BKojgSnZlvZWDZEa0dBqxueIGYrZhGt3qyUQoOIA7JUs8cbp1PF/oYSi6
tMRwjoLit5cqsFvuJKEkgNOHg923wVjs1G+jdwqH03nxNhTyYOS2tM+b3EdKasr8ui6AhP2K3e44
R3IRoNnkmEhKzCjiL6JTv3+yG7gLdjquRTZFAxi9XNFdYeBkmAfsjD1efSVcGZQLBaNmAr3JCFEn
P8/9qv2rLHujB7YOpFXkmojh+8GrJYKilaUc76Br/KsT5kCnKkGNJ9yKLrDavPPjNeVqDOnkzT7q
z0ZH715FMHUPUQHJlpFMJdxx9DGbnB+eO8SdnXecmD8zcfGJQV/FFLK/Uf/u8A57RiT02fIrWTBO
s06QNrh6YUBBTp1dEvE/FkupYSuvXzB2GwC6cR4x0/3H2S4tU87HprBZa66Z+5fK1iLM7nWjppJB
b0gzmgDx2dvW+/0PxAvYzko4w++G0gcKGoZyuD2p271OP9X0tIlPZb8uDfwZNs+LqOKRdaf58Ypd
RZsnCY5Hp850DXTGu+GfmJPIIzfUF/OZ7GPAnAKcZT0LYpmj3WW/VXfla6zrsIO6fD70docuQTUm
w0kN75Ji5h1Ss209Mafme0IPUwo4xRSpVAiFWPiUIIvBmCVePD8sv0zD05zM8VUdrAmSqFfDQM9H
zK1YS10B5Li0EuGaiFQJYFSZ7p2blPFr8ZFqaRmfdi2SoPAcPiclLaaxGJaAwZvdQX4yzBzEGr4l
d67TS3of8eQB4RU8SXqoSN6xOymoPATH1JSr+QewKdtuc/64vLS8+FEZzwc6ErP+HQoXJ/j4QYud
tYSwtuaKIHLNpxuwOLbztX/pijBbBh4vZ2fC8iqRgczU0culitOVUhVXXtPL57xa/mh4homFJpgy
BkmCfsjQslmnfSm+N8FNM5+6ZwvpQD02v0qpA7T7WCI6y8tcF00sp3A9emUNI8orqMqTbjbV6uPe
pNvT3GT5WJDGYRjNAsj1LQ1Sf5PcbFk/YUjKhA2PkYXm15+NPt5L3ULOigMPhca7IETIWS6I39f5
ITlD8PY7ST2Inku7naA4L68FmZxy9yezqW3C7yC+9ZrMuN84g0sWQfp6GHBpg4L+Iu1D+BbLw4qa
8N68b/g2RTdBx9jcZ8TFvaUs+2EdvKy5XU+9C1SU+JXDE4ptDsGqcD/0v5GY1Cnvq7TlqHbQGBvs
REFThvaPlcOs9YhKsdntyfVIFK23ZcfDXETObOPKW1KTSalsNTD9B/iSQiKrOxpYxm+TcXoiiAtG
G0tgjJBN3fwlw/EMkykpkiHqeJj+tz3cmE+fc0oNb52VDzGtnAA0/45ZU4u+SouFlgfFLRojxTYW
Bm/Znlk6p2VoZpJNrATAFHCt292z892spJ8VFVZlXNFpl4D8voOslRfAJS3h3oWxnEE23/OUv6Yv
jRN9Z7+cuGFbyHQzJBLHX+7c1wrO/yBcvD0PwDCvItevReNqKt2DxGosvRetiVhfcw67jdy0rpG4
t0COiWFAM3vqi9B6XE0yIz8NWFCnF1uz1Whxt+AwgYY+lnIwzY+qcsWFT3IHvcgWwe0F+PqGTPzm
z4g4yYSvQ0xWFU+4gd58HWmkMAGafQ6IyYb0mwEcez7fPQ/qbdgwjw9nOh+kXf8NmPJI3FWYk52b
tp36/tYivUdNPxnm9tEjkx72uF17SDuBqVOos3E/DZBpdORiD3sglPYwhHFrPdJdoXvhFtI3mktW
B/ogFCMGHSGyafRo4dqSOLpAoPUw85RsdLBNtLIMHx2Zahrn30CCrFph1bbxQ/k2vtSzaAz6bCRh
7RZXZ9a9v8U2+gclNmLIFWQWkz9pJifBDJ+4n6xQIeKfYUZA7wyVzXSIg4UgTKlgenspFoSDWRuF
NrhqkgfWtwusICZpPoIuvMpP0w6MIz0lChspTEw7BdQZu8HX89G8vGX0OJwRy7b0bkxor8OFZ+dC
9dfvE4gFXFVEh9T5aARWFeAp0GLnBfcE2cHI34KWAPe5ec3EM88nkXeAgDcc1GGMLiJBE44Yy3lr
YOp6BLV5UlsPvd7uYwwaTXlu1E6tDC47SiXFftpEYzsbdGyBk9jRRH05WIrSc5GrxH83YLfjeP1+
HNmRV9ixx4oyEZhhgWjUnYF36xmsjzJqPV9xueH7yM1aUrDN8DT1AaeTG6DWGNUSfklKPV2EO0ay
l+1FPhnhqXxlFXdoXAtvUdxYWxA9F7lbE0ab7VQh3aJQ2YPpJiXoQJFrJeb/ioxeOhpTm3uJIE8X
ZwS2I0KbgrCrU9RxoApEVxNAO6TbxROuDaJiRnU+p0MPaU2yu0q6L5idy04CJCMNUZANFqbtIUaX
7Bpu3alnLYrWzgI6Gx5tgXGIQ9vuYLeZc/RO4f/hz3cfIZu584v+xKDpS7qMl5PWpjbT+bmWumVa
lk03Xkh8feO9C882JeJ8oT+DnbBMXqKS+upvJKvw14yzGRs3IgOWEqglq5vhupA8YNuGfW7NjZhb
vKVT5WwVXGUZ6ggLgiu5tjPllo3PnBdYismDsomypIsdXYoB39JTfM/9gX59wZtBA7gb+8XRjTom
EmoA0awFL+yFZzPGbnOTD0f4n5YGGrcMoggZz1Fg5PVp4OlTna383LWqXq+wEP79lsxEH76ENUDw
EPtniIUAUsqkx/+UeNZgBK89RVBYDfpj9n/g7bCvgFy1fkUMXdIYiuCwNWHAKxQ7dge8pE12OK/r
N8lYnVLh3BAmqO3hX3EnDrkpIG14GWD4iLO9KWedXmR6DuxIPhDZ8fzTABI/ALvCJtmTnv5H4j8R
jv0gBPpQG3X1X/OuKrzxKzUtlB9tkqVUGvACqjm/krzJzkYKZTtRtH20+ubPGk8rW6p/GEEqRQal
RPsgA4K1WZsMGQkRqNQBAa1+YvwiiegP9sI1kByzOBTGwznkOwDGOXWD4uhHD7jYyDaqrhijuFYf
OzTpHaOWHg2vob21lFc61+DJMp8D/XG5wozs4II3ka748PM+IhY/jdyIa+coiJlI8tez78Spa16L
39suJDNL7uMNBgufZq/IHu8QxPbwhNJuD9CMn+QpF7uNcfRKYcpr3+niZnFNNiieSdU1bEkIuvR6
tiUoHuiXISf3nlEhwuNEDFLTUq6pzkjjDcQlWszvmGYbfiz7aljcd7SlfbwjtWIlqSM2ng9LSDfI
HCz/xjkFG6Nxla41/r+e8IwwS2PLPDHJyDmnka0jlmzvPFMh1CmPcXEEDPKKawhvs36HantfyZDT
yg5m5xzWmGI7bzW9KwztVUWLB/5CWmYCslmhHj3LlFqSCIgSr+/hmZEViMCO5o2kFP/abRYElpQG
lwzluioohNTGtPNrJ4SlMK9j+0i8HPKaxrl0IGbxv9Q1FRSLXvm2PLTKw03tHujolQw1HGKVx7mc
TVszWTqGdnAu21QQzUTUxN+e5oGTalYmYlg60K43E05uBniukQrY6Rhhd09KHfWY8JwG0qMsNmLl
uhIKAhclHbtAzccSXtZmaXgvUXRt3Lpo73QBlAvz+Uf50DLY9vYSlJ4Zknkt5lYr0KtPSQPN3n6S
vwxKa6hcoAkiqLHaAbAVbIkwgB5pC3ByQm3uDds0px0DwJbJy0psObM8wCHOj3sGkSL/k+vy/nLL
ys2/WQyhJkiJvzUCPsNRLa1kLJLec/FpRDzu0YWEGS51m1EFuk3d5rEbOYcHRGm04Tntu9h5S3jP
zNfXCIse5mm3R/QZ9Qzo3RrlCRX14/eDaiBt2NdsegWjTCBYaIeuqX2gX/Dw0pUb6MNpDBiScyfI
drskpbTyQmiAdsEJ72WnJqkG6eH0dC7B6z571hd/DXq80qO0dkDlvfNsMR1spverlJQu8GTYWrxJ
92Fuyo70oMT1mAmVHFyd0qIC5bnGvTSfo+HU02mf3gmGKXBjd9IwJt0C8HJc4CBIZfNhQlDyB/KR
7j5lUksyvUQTTyTNyzOu6e1l1OD31k0wqjhvhdPAoZJPiqYGzPu29FCXG4TdwXVd9WvUCLDZubO2
Ky9QhWzXcFiwGvylq0DMsqwiEyjmKWC4k7HRsJDptdG62ySv+tRPNG+vzVrOjDNYDNUP4jKvPqX5
BkLLZR+ucJtC5ThHKVYmp2WdUQci5ZOBjZpjazv1+xzvIoL4CV3aQ3l4cODVfnzYlWBCym824vAo
B+RvQ/M66tiJUQ+xebRG0oHRgvUZByTAthHQek3r04okWXhQoBwHSuk0EyQ6Oc3mFLPUBuuC1pIe
/GqR3/Fe4C9rGWSyTCVbTJ/EcA3Wgy4PjIARYW7H0GJ8t2bEctQFnsd82IumHUH7NYvZb3Xm6ydj
Hnguft4eEjfbJydYUtOScEUExnSko7SmzqdE2dqPzkURXzpjbdxZPQvSOfSwoNSCwKGRqdMIF6k5
2jaStq1NkK/CwKeZnvJ+DFlUBs02ZHOt7fZoNQKQwthA7bs8warc3DhlNquG4N0YY3Fa5D9vcWh4
8IM40vAO5X0ngvCK3Gpgln90w1nzJprGdg+FEmUyXgRBLAPSkFQrvVbytuuWS0OmNa3xMJaAkcXV
8Nkhe1TdI2nxJDvqdkXP1qS6e47VpkGK2/u90D+anYvl1/gzkSHh6NIQtTyki34gmUwpBZ8+GElu
vAxh8jQKmuROR3dA+D+H8ln1GS1Qv7peZlDGR28rTmDUMVaT/TXIu8SUtyYndfiqbzevHb8HdZd7
vEPZ7PGFMpdlz7cJnyXNSKiIpIPM4MvDNsL5Rnz1FXBVcvDHlUxce+m050loZAZqjbJal4aHaFh4
YyxqkhfyHU8rEV0Qs3L2+LBWrkxE76M+yjEe2A/bJ9tYdSkoWf+YtUtLLHMHXkrN7gWZSZ/P2kNx
LhsrVa7jDoBgFj/fYascDc0nN7g6Roh0eZM3ostyrbsAPNHWQrV/MAyKfKDw0Qjinbwudc4d+I0f
9DZhpg1y869JgwW0nviRDuw8IW39hY9FMsGbyCyR3f/sxBMU9mcmMrXG8XjJ1yTAvj7eWSCyps0x
5gbaFIECtxBckqjvo3l78k1CxqDShVWQ15pWugWi6X0fpX+PjixgDtTGUk3jV6jMHjXfWwD3hRCY
SLD/H8aepwdp8deN9Dpz5M4UZgennHozI8Z4YHrfnp5G4PSQxtLiKqkksouyU3PhVsRsIemLcldH
bIYwv2Zo2yAjrinXgHOpDv7Kybs3MeJ95ZJ9dVm3zi4m8aNmUPKhPmQVAjSS/k8LIQ6N+hckcoSF
rYtAl3gvZY07NSH1LI/BjQgkYxsvQc3f1/fqsRrn58qSHtJyDEbJP70jRIg3e6BNMZQJhMmfG/0B
K0b7ckADskg6LYEYGsmuY9hOcOT7Pqyz8Anr9qsyp3xMMTMYtIqNxGvGFGlz1Px4WmHkp8fSynJ5
5iSRdo3xnk/BZ/lGZz5mEvGj2ubzTSxPRSwO2Ft4NbE3YYT6T7EQrMVXuL+LgjpzcWca8Ot6Itty
jvDpr5uJDUnyD2KOOAuYgWlo6/T8u+NsuqCA9IAVgaJctsjWBWf7qAkL3tnB1GtnCZuprmAefB8v
8bC/J/ZONnPkm7SJhf9T+IEeOiF2xEehUsaQikKz6JDd5+7zr2+12PPSj5YNt6nPNCjuZQCKysS5
DSHSZQx8FNnUPm+s2eoy5gjDIma+RtGlQvpDAeWpDQC9ihLIPxUAGaB7LApAIu9ZKj82JdOt6qLY
pYxIDqNi+Gqx+yXVjNU9jWEbYt3z1EBkDZ8IB8R4JBboVqOgoUCXxf+xWQTwIj+CJyeKDgvjz/SV
OnrTCBrm/pr2TGblYUAPQUYHFKu+4hbRV8ObrCyX1sc1a75gge4TtSfMEcxEodF/rSwuDH6sAhfV
wVvo6th543tnCYz1ZTxHgC603rcSM7QVx3aR41gToegD2qtY3ukYUkuJI05k9pP0V4nEu8vYRbWd
8mILK2Lq1Bi/5TDzrTUB3OxUGjJjhEUFoSus6+SfelUuXmgoP+atOP+9J308bhLdUOdiOiYMpLDE
Unn6/bd5hUSPj+8FNN16aOElnFWPkmKOV703+YVQpCyvXHMOa58WOJxlCW0OaOtm6mdB07uki8pC
Slf5avrkQYt8xvAfqYUMuFG0cyQ5PTMVFhm9ao33pFFTRQvKfB6/54ASY3KaANHCe1GJq1y8zKyp
il4wu0SjfeNMLztAhwaP9kCoDS+BwtG14FeyEKQzxZO/X1nZ0bgRFEdQfs7vpLuXcm+q+a45FNFQ
jya5w1ji9YXtafWTRgdVy5fQK+wcE1huQ0immITUtNP0RJ97KJ8qUphBR/CA1w7rdBsJbsU3mcUr
Y7/om6IIs4bshuye6/tOXGIQaXC/Ya/XiZtLdH9o4rlSQsAR+pLfarrXm2LojL7IFrxlknALccqv
wngyHhu7YEcksa7WznlptddY0XWewXorHkI0fgrasyKKPul6Bw54lCRgkpKW2Y1IvoqLPGm2x9EL
xh2cTKcidzolmQh3SLnGI05QW2H2/KHQvjWUaIQUGTvwQGTziXg8yhcAdShtbI3M/bOhtiwnfLlb
B0KB8FPyNd0xWCHoxcinF/poQlZVsniOnQmIryoHIIbWMRzArDaDKSOzD8Nu0eXEabnp/7OAuT1M
Y55rJbKBjFiTJf4r6ktqMlZOfhumG3Y+GKY3Ljdc1ngxfqGsaa2Vpuu+dSDriQ3fQ4RRGSiQXhwk
+1NRTBRvonk9gXLiCIdbcb1qng/2M7JwhD1CDjoVneHNv4QF5ae41ZQh4Xv35Xu2pQKsPKI8AA/F
T7yJbtxwssHRb/+SWwxzbIRdBirevJ3JIlOWvE8yfLj+rcmie0+yb+tORTfjqeN4duHEYmh9dvJ8
CP97fZ6+AzW17zOnbozQKFANkrlVT+O6GwMZ54V8yaPLHZ6Gvqlp4iMg/KTwEXGu1ooW9+jgKXDT
E5YBrZgWzxfm8LUPIiQpitC3Vv1lq8ZiLy7xpRIErScdM5Al0rJ6RY1RCdrSLmVYN56V28qa72g+
2Ch32vpiRacpNp3rD2XqGNc4dqd5x0CvRKfqeyOw3/wYAYjYHaCPdMKL9N5gdRJyZ8nNgTI+VjqI
hOVRnmwUgEkoDNzUQCjINTalfvtvHUtZvno0Ck+tD3tc79csm719/MYz2Kc1EjhSnJFkvGiGiNtx
mlVWRz5ZAwAjNREhOE7KPdAR9vemO99F0OF1BYSwBOAfW80PYDQ8fp9pjMzAfMDOCUNcjZn+UyX7
7U+AaWNnSjfcosWlDe/EOCyVkS6c8oORVt0kitdef0t9Ncyjfa7JLhMi5ht8qsP7tVE3yvbG/nH1
bWDbf2PTVkW5BKrmVSr1eZam6H5RusKcUxkG5P0dwTtXU7EsMciGok6M1pUXX+rEfO6J5ozdr8bQ
9PZvfnNTcfqnVzjeQlmthpeLztyrIbv7+1EbWPknwVnlnm0Q95URDHBPmihzBbsg9+OEEiKH4URs
IZe0LqBCUqpaPQJwSW3s0loOGrn2kBT27qoW7T2/cgewPtTRHYAqo/DSt7IZx3tI8MB4VNS8BgQu
r1BgGFaOz/xT2bqX4e1ESdjknwlfoozHQZ9rZK4TEFlASBjxr/FKMiOxl8B69hDlqtVYF/xuJ4HN
1f0r4lC2E922Z+Pa9Cygs+KgzDaqqCNskHcGg0hu8UCrKlBhfpWrduj9pDGKheahJza65AiSDgIB
jm0VgSEFhn166Bj8rTSjjCHXmwQeYz2DPw0qdaCeb5SrkKnxIddnVJa2zJHYVimLJuBiUNkKdgA8
yfPODd8HupmIJlQirQ3jUPHX9EiyWFpShMV0iyk5bVFi9n7mrBY9AnJct1Q9hGW1e0MPsI+t8uhm
wO9kUpPiAEcx476YYG5Cd64+dRJKmyMjZ2FI2aw2XFRJfPQOXtNhd68mnEohKL98um9lDM7XUFAC
UBwO5L/snVSvZaQwDx5i9SJ05X/Gy8QmRJuqwtRiPoGfDRBtg8/DfjmNsdcCKNEJLw4hpb5XDqMo
Qe/sDAbVK1xwrSjiYvwzDbKAsQYtAjNVGWVZVp7nlwgljNd/jo/Wu8I0+gt+v5UXPg2dBAeAMbAh
Enaezczz+SJtZ5T2JphqUYf2ggy5fQ+vFQhuGhKDpCfnultaJtblvgZtdfCv01g9j5N2nS8oBD3f
Hya42q/CSJvKN07qnzUjQCj6eiBmAbh6CncIPIWqHPEm/RGqgeo7yqHW4TCvQGbTQCtI+rW5wVnk
nYHI/bMTDsuSkgd6xoHaH6yYWoFhkL3ClMRc3uMSnBgTko8DnO6Z9GxRNsJqYX9daVG9xaKnpndG
nTaspOzk2555g+o159f80Ej8pT0+IW5u2In+irW349/0/pF5f5t4pJganohhtSHAIU0AEPDT9uvl
yTH+OI7Wvms3kXuCUUWGj7w8wqY7lohElM6GKouZTX3EIpGyyl/EIDjIDL/GuE5VS9vNXLBxbd8R
t+xzOS/3u7vh5/BmRllEluMkP0iEBykOPQawRNTNMv++CFGiYOwFvBl+DON9UTLe71uFYHptnjPC
N1b3H0Un0/PPIF8ysmoxsim/PjcXpordznk9Evk+NR2V8IrrD52Ey1h5ZXXVdTlxbiWE0jMWqa6o
0e/vmvo0+1TUZWn4NU/fdtGyPiuWsj21szS6A7jzwso7HPhLCNAZd/NyOQrSq1lXwmTvmjPmZtVt
JRg8XQ9fqeYADuSPFm7cdEMQplGx9cq7VFIYyAWqoS0wgyq3WRbZ/X4ZZG8Ry0qcAhZSyPXMZtsS
ptdHraQg584EthZpP2zBc01S6s1fd8qECnn0x7Z3BX+w71Vpg6mnMBBjCXLb22Fnr21bdbLj9Us6
pwnO/inIEDy1sPvfBHhMwQgeJxiXsFacOUhxnd0Wu6ZxR9ViRPMN6WLlCIGd4USsi/igXQbg+HXx
QRbhbpqNIsF/F3atiBGZ05LnlMUZXCP9HIU9p1Lad9XFH91x+7bo8mFST2p9R+y9cH0EmlmvQiII
ASO59BrXK8SeAG0dkWHlTu2fZujh8Xzzgnc+r3CM75aCfL9GsH2HZSMKuMXm/9fhWbBv2Gu83ZTI
7EQZzbUiW4oHBbwWy1nSSafAix2FIzf/j4WvVL6ebiCSltBgxxu54oWh19/EwMbozlHj26Bik0KU
1YoGhqNk2OL0RnolExOEKI/kpHXDo9n7nmuKHfMYjvwOR2Fri/DeXjnyDGq+GzVCFHV0b970ZOT7
z8qLf2H/I/4dtQCZJue5vNTBfRMZIOJd/Ak/kTsdX3w582Irr9DW1S3xGtzoYlpt+VwV7KLRl0ge
0vkRVMYnd58bedVNz0HwmNJuMQrDItAdCGj4t3Tm7v4NEe30xZLWEvWTd2KiG9FkXg9zRWMbhc/6
3Q/hffVH3JozZgOVcPMA3nBsFHoeHZgwiWfGXIdwIw1GPbdUHTxdsdq2f7NFsBRsEJkGHMef20v5
qlAkm8RPcHFQ8h3BFVS5ldR4+fylfsw8BoDYhHEgLRWXUfF3XiaHcu104v2YGR7I8/cdd1MwEJAI
WMA8J8BvXUOedPx24joZUi2kED3qK0Hohcy/FkDLVxEUapdVZzn1sN1UjpByXRU1d4N8xP3Y1/LS
cLa54X2ioLH8GluUsG03jfe/B5oB0mOVAp3CSmB2jaAYT3QrPmD8loqDFXWcWTvJ8AQR9BGkMu0l
jfzge9Y47a8tPf7M9rJag3MZnPg8da8ohHlAHvfqCRlULYscIQm6xhYsKw9CRZX0XE2NKxt1hXwK
6LZrtqZCgb1TA96jtIrguWEHL8LSJYGTZ86BhUR1uLGQWHJRsVDFkOa372kI9PtNQCVpL6u9O7t0
4IHZru/F0LljlFlKgYSp4e8pnnpHAOM9cIIx0dTnJ9w2gjxd98rsd+bdyxwRwP63vJ7HCtgQdwXp
PC7ofFlFm/LfOEXDhZwRr5fcWgXVSbdKdyZKKnwQjkxzyojmLPXy0X+UNNA3FFSBLl+WDZQZY8H+
/J4LfpkrO2ijzgarSVa6LPwfcPfSpMlbQikeYC+TpP3hMRzedB+VNaSDCgbgbaKYjfTYVMhEtAFj
nZHlq92NsdmsMNjO6o+Rw8K3KthftdXF7bM3+v2gaio7Vi3MBB7KjjyIH/K1l7MCicKLnYm+H0Rr
//cQb/yRKDJ3OAIImGDmH35XiRWhvkkSgBcrWk9JULtnU6PbTYtmRM+MUI/PMW2t6bReP/A/tt89
vhq9vhHWvTP8yrTgx+oU5bpVtRoYwc1/Q8kZMD4KEnFMVK7IJ7HEAq56sHRCUYDfABd1/9B9/C/m
CZ92mDMKEXEU5/UTrXcSm5K6Ll9oAbbP7RQHkpxG45oOzbEbWdoRNeYKuHLaAPMJlvSZo6aoPgz5
O4sHKFU5PN4aFahoqrBjW2+0lkX/fbuV8hiu+YD+PW6Y04/UGupldawGDx86R7ABj+pCyidS5R6R
Dqj1HTMZr4EbAtlRS2R41j+0B58mk/sbqa6ahljOAMrRPxE+06dBfoqFkGb6XbHswj+5lFH+92Z+
7Yb/4a9GzlDJwtscz0RPZJpS14Oywp+/Y9/d8gDHoNYAvXLx8wwpy6Qsu6KwGhEOuSzSAE6Bc139
eQz2IDo5c5nmbGtE6fC15U78Zbbzi3DHTeO2A49qI0jHhofcK78W4H/COM+90aHQs2WwV8ZlxrqP
O2TmUOZGr+KvjAyMi2UW6P5Xo0UGgBA+CVvyLAzcZqqIt0283+5VGI5IUpiD1i12NST2TeXe9A8r
hc6o2aLnFSvP9wDsBKdGH3AJ6Oz8NpdIA9X6/7/wLIeak70rr6v8Tm3dtHegxOmdKb3/0jGgVH/C
dmzuDoljFj/aVBa66K6hRZzxtOSU1LY3KOQqIvstmr4+Ugua3U3nIQtAY/HiCkUMbuyK5WOj7qx1
0gJe/4FkkNvWf3b2AqhlJ1ohJck7X2D8Ja+FrGx8OrF1auSBeKPREC7//G5bxjz4P7DjiMkf+Mlx
jl1XzUG6TtESgGNZgcvKEUDaQZxAaSoTY7sJAXCqrrfKIO7Ia003yroECRqQHl4vOBmRmYQgwKOU
2jp6rnAMRunA9HEIA7T3VfSa0DTMAyiqyLmugwiLaiTR9z7B9gevPxrq56mFO1ueQ1Sj5a8FiKax
vcoxkZ2Ce4IgSdzQlKjv2Fg4o2CRb0B2/L3BmVkTK+xrB75kOtRrOnLBfnNlu/a96poJq1qgVz/8
YDsbV+XhgAwqvbAxhotCL87DJTRnfn0GFuyKTHkLp5NAs/qxXORwd1lWnw3wphZeG33RE3NuaVx/
HKXfVH2RAfDXnP7sTEHuUxOvbrPXB/l3mCEcU62Tfbu+6sqOyzWmOs+gkMh9+dGS1WQ6HbARk//F
EifUwPoNF+0zyqA/jFNumoxG9Ln0atE2A9CUM7lk/eQpCCvfs4yOU/qdZ1F/1wZ7LoSCWGlmH6D6
tbG/CF9wLvvbWmmJN7zGGk3cpNo9R9/zL22MbW+y6SU9Dmidr85OUTAGELibxCbnmSYqBGu4rQ5h
GwByy/JsI2zRPfhendaWSliu9s7U45JtX6zKuich0EogzH0BKnOntE4EVopiu7FdvPSWBWYZKgrL
QamoNBoESOdm98bytEYDn9CRs4/MD/6GAu3UqGvpav0/UzhMElf66fe1aUJuRj7EB0McEWDOEOde
SzQmGluKYKeNzJtRu+QqqG6ldk+UJsyvC/iRcLtAcE9yf3nBe1bIXO9wqNlRKLYfwZL6rpTx5jG6
4NsBMu8DYRalYD8Sk7ery8CIBp8Z2c9Lk+aaxx9hCs+LpN4v9UXgpDBTGwW9EUeef4/npXImBVgu
fr0L6/Q4mJEhF2tXHwga7vNYMwCMGWHNapKtB2BEV+bEOeYNY8Beja4oKz35gTTSSDEFcHnCnc5I
aoCT2Y3mkuSMJ3ikocukq0QIlvFcXzEM0xdTnBxkWk5gEGkwc+Ps+psVr9gbmc45T+u6tO365i2I
3c4a/Z0MD6woQxor0ZwNhg3L51GJ7qKPGI738O3x1Txmex8sUchlGD6AjF7xT9bHVi0mFb09/rcW
sTuYR684cfjqHS/AIBT/2zHJiz9mQtGNCxIGu09UV9r9YHmyynVvu8ZY4ES8Yz20qHz0XDDTT8vz
njOvbe7F4V87mlAKd31wIGRBBybbGkrLX7qd4NxCYGh7OeuiCXU0P15MwzNyske+hMZVQqNqjR20
ewth2HeZJVB+GuPoLJ3LKDIZKLaY1KCOqdi1eDfOByYIZE90SHo5ErsM9WH058ToKv0SulhFiP2G
lAULKQzmhA51iyUQxXMfv2pUZwtSevOr6mLTX8MjB58kF9EYdMZXdXRUjG9cg8tuoJwipoHtt9E3
1tCq7fmngfRXAAi8SSw4NUG+6x0K97A88+uhGd5ALClV8LPw78xFSBdh5mBNvDPte13EnfZuYXcP
DwH4Bmwz3pdBVs03u6d7NwkUrfOdOeeYTOR8R03mQlTp4tSAS7/ZN3KsWkzhReFLqkubNKpXVdTS
3gcNHWhYoS1ZBiUBxS+ahXY97Ts8MoPSPlwut6PnTx5MSCf1QqV4wQ/TaY1gyiB/UzM+ve5n7ULv
W2Ni+ne1fSfGHcJCcHsQxvhz5gj5rriA0w7uiIC7MYUKGjJC6pKg2joP6q5QxhljPTZppmHnOjBg
UmT98T07eWMvUEBoLYg0+hsztHxDEmG0kMY+M/4EbTXFnOAzVp1fGe70REJB5PW8GMbZa8/zi7N5
aPXWJUWkgMFqyON/bKEHqps3JFX4lDsHK2PIaMe4oj13BWirqfI2XKnbV3X8/+NKr8ZBNiMlzR9B
aJZXt8ntmXuSAnYoFolgjGbWctff0cHB15GDwk3EYJbadW22slh8utTjGTVIkkjo8Fy3CZkN+zOU
wyyYB7/2ZtPXMBQJbVLC5/8Htg3qzLLavaCyaWh1qv86HXMhOJuAfX/IweGEj56eX6KBpK5Y3AUS
ya0IekhxM83Yr+INNNHuKg92YxAM88jsu3OO8rYMfJWFcd4fGjgX0CyOnEaLHEuITDmHocH19/cY
oIqZK39+jM4QVVxnTp4iMYcaZKfU0TU2CnxqGIE3GJ4kfp7iIP7eXyQHgKmJSlOR/mSxx3lx76yx
odH3PCICxJ3RqY6PfyAclmCLSZHcdUl3/sh+dquqS6xDKAXCygT9GzarBh66sHe+5d6iOw92qC53
DJtbmmeVyepG48dtWkSYT9yEdMAyirB6g0RAUwkEb5O1/UZgIghngej7XCcEXnYE/B94ISVcjr56
EBAtlTI2sJgbT4N/TVjNaoG9KcftJEgswo9tPRi6LHF7UxDy4IPevo1RE1/U2U6W/TDNuDWFyb65
CKHedRnG8XDTWDGy/oEvedC0yppW4+R9eyD2h8vLfuISc94gWEVyaem5CZ4L6+lUZVLmVvnN9OIl
uAKEWhHtCxdS+vVKvqQCFxPUTPbkgjnrbSP+UGRnB4g10sM1WEkRAWEVzhrCXi7GrBcftjz870ud
/L6wWoXq/cGqNtS1Uu7pyjE0PXHIyJ/6YnNaE1s9QWjGXMjlXKf9aXdH2xLDfh4fmm+HgAjdNCVD
atek7AsuZ1NSDMdfNIpcbisDG/NzRxrIKCT/Nw6zVxhTmv49w7Vt/kBovYQHbLuMak7euObdURAo
7Svai7gfvApCxrTg7rlAekk0IS9ufLOCx+hcJhwVHFERXYizbmKffL8Va+9gkXgI0krpDOCI2RUf
QgPkc4CnRrrRkE9HR9a8z3Kk/HyfEeUdHUE+yJPFFK+IK3nAMvSOH8pooFIfJYMG3IGKgIi5kqRn
deD51+9d4mwucOk7W378QcjSKDWch6CfXf+ZAVWkqJCN9fLw1PW6f+DATcRCEMpCAV8sIsyujZLP
GKwWs9yR0HU81QNkFmNaEA/XyZx+zZjeZeX7u+SNsO9gdZD69qRDTOZJC6SC7ZEL7Yu8meDuqgdP
FfcfEcxVNHm9Pnswm74iO8OU3/dOMOxSsgMu5LzFs9f3+kaQOWBsJzXPx4wZqEm60JvjdUq0XzyH
cWaXkLs2ZD5UqgwV030fudz1+frJsMOK/n0ErzN3qS35pSnswR4X37pyN+saW0cP9SEpzW+jhqyj
rcQQ3bVmQZCa4wBxtqZn16y6NcnHQ607Y7r5Gm/KLue9Z+qmqvw+S7rBt/E0US5/U2nKpczXSfdM
yONXK1tz2xTxA5CehCW9dUlVlVmDZLtljVaWwTuSKOEZGCIUSwPHZVtKjqfSC4D3Xd+kuTPRQN+K
raQa5yZ7YwBPqwHjmOdHxn5YlZwvp0Qms86J5gpID92RieKneDGufH09gwoLK07hpHGJeGG5iXz1
5zPiUvqAZODpexPqKjQ64sk333nGvb9tLNx5kq151FzJMZYI4TaKJYWZUWx+n9nhm2sUdMq8V2L4
3Tyi6MrO9ASwGQkTWDRY3JGLGEG+pDslM8isu8b3r9s/G4XOSO0nqs5BHbVlZ8vWzydtS+06eOsj
D7FVnFvUCRMcSmmK+aeDhZQlqCGDp2hzW2aMzASs2UEB9kZqwUponla4uFloXGngXyZt1KA2tpgq
yre5dsUtwqZqkA8Yjy2qqyGpycVOmkZWq2FQaYplAl6PoffTyr/lf47DRC+VspWIAS28LxpL8cdK
XPf0j3wDI6L1EEjau0P9gnU9DhbC7T2GLKwCCY6yIJdKH+byLpZm8gnrhukVHLtrJi73hKdW2A9y
wxOeGC20UcnO9pcOPZy5oEws3eFtrE8X7nIiVYH/ZhZn+H/KgsWmtI+ALGOFNmgqV5ZzDimu1Itv
KT/TLzDUmh/DjMOlnokdNAuh3fw3e7lr+TzlIQB4ZUNBt7Fm90OhY1/YIu2VMM0BkB26jn6Wv9Pb
eJsqBq5S4jnjsUnNPbe+krURYK7IIO19W6W7mQ+w2SwXfS1puYIlG/BajnNxSsI9vEg3TKo1scDa
+r2otS/CWNSGDn9TbEf+tlXYQc4nZNVHKXW+dHtYB/rOGNzSEqKZG0zg4cv88UTdvYK2N1wMSgo7
thkpJ/6mTEK4yxBKjcTI/v5nBdQjC4iFHgx+MN77R88gdT4q3omgOW0gzQCepEMptvnGzhZ2fuiX
UtTpgaBZoUxWRU2JVwNEy6H1AxSInHg/LlRJHNhj9zvG5AlHWqs6s7D7K0rko3teF6fs+QxqNOe9
DPZZ+EHJsQef78gASruT+qd2OQhn9HDSY3yV/Ykot/aFwj/GZIkzbqW+f1O2ryoRZEY4YlQEF81N
AYZvdw480FZnZSDR8+1nsSsPeAvMfrquesla5pUkurJjnf9AUl6+y29sdtqUl0Nu/lBUEIuu/wAc
Tfyx3M2OinPIvioqfr0VvdI8FK+NEzHkKMfMcZTZk8KXkLFeLUpXui74JiqqlLyDM8lRxv7bb7ux
uvEdg4Y/qsg7bu0By8tuYMKsL+VRINIgVcz81+4+QYuphJfAtavbdXGzcdZyYvts/e6rdxypgktl
aMofanMlIholFuc973ULS9XPdm7rqfc/hm4m1TQ62IBh2BABesOnF9KpoDPaiGEZqOkZtSIfaJmK
QGvgXGaEoo+uEUNYwJ7wk989UuxHiUJLq8UJtpH37AZPS1RW9poowjWfHqU5jQmDOWCGwlbg5otE
oKwi7V1UyzBn4C+WjwYqzzR1TSmCvd8pJjDWu9x6GdYgfiPrweae7x8puV6cF8nxqL29nxst0fZH
N/tvyUMkpxXmpisCVaJqiMha99uvJjjbJ0a0H+AzaBf54wmbuXubhvnSz5LMRG0amU+VF9aS+xdc
msD2NQL4gfPzpB8fgcv+nfGdzpHEXJ/Hp1a9Sk30lSM9RNtstPR/Ota+RRCLvZwlUvm26DJOeRqN
nhH7WjwkqoDgfwgi48b11jXnzgFsEpLHI0n10UKZB9eqQYUn55dc4Suvx8qgYGQl975kczrYYgUK
zHVm9Dv86MInaQiR2AQ8Rxn596A32KfZR0kJbEPdPZj3OmIMpsHNK3E3OBl9ozNTI7KTCS7mWO77
T7OBSdnKJUeGoTuTmxn3WQTxr7OVZHh4bY9p7aChUQzd9Vmkf6yRC1glKfwSN65vfsLjrN1/AvuQ
sGiQtkebrEgAabXuMOXrqBlguCiSGMLLReNH9mB7BDHNM7O95YkoJe+G7pZpJ6ryorybP4dmqLP0
+Zx6eELpfzpcD259ir4TTMCmL9anzHX+s3eef6QMuTtIeHZOmMcPe0WyQm8JkARt1XEQ50gARIWc
O4ME6phs2z0OVyqtt0XRZEW7ZJVR6Rdt+i4TndotDjSUdmpvekcAtHNSCBpE7gN4U2FCDp56yKcy
+FzRZy9Wdq1zhRT0Ys9/glxvwiW4p+FMKybra8pxpuWbMx8p1kwKIxuwgETWlontT09mkS6+iyMj
DMEJ+668/aIsycVpFU7GL9Wye7he1msfZ7eo5k5T/BaU8K9Jwf/EKA9xVa8nVPo39YO5N33WrrRY
AvsuOmh6/s9OfoV9/g2AZyVdLa9vV13to3kVWEsUOjK9r0BiYQC7uTF1ykRvZ5pccra6Aq9i1Hsg
qcsJllDxQM/G53Jpn/CK1Uv1q5BqHdNz0g8ni2Nt3fGJboyXbyMSDBF87KiF38nmwGEV51sLz2/G
cR2LLzcBw7SBXcRWBC84FiLGbaTrC/FTomNChhxWuELFwOAmbpRH6WofZhZKSTfSatoSRRkD4F79
laRas5+ftAny0HYMlwdgPoDWYOrk5UdTTe1F+v5nh3IctrN+ImP4ZT8PByb52Nx+h+5CZlX0Ht56
CABb+KnvBJ23DghxASfYMAKITvmsQsR+MNKhn/1OpQ//aiFzQMYxgNbXWAJk+gdH3YLlt0tKUqR4
ldmdC5s9Prt7Qr0qhAyOMsPPDoEl6gK7Slf5R3KfW/jNq2ivls0cTdaXOUGo2T2Wq/+bL2J2t/Qg
5RfemBqBikuHMGPmYTcnS5gfAC63XkP8u+HjNc/47ET/hO0kxWhT5f154rAFzOZdbsQvW+xFcL/2
0SmWBq0VmjyU48KB5LcDWVobM3uViJPuY55UA//+bBecY2rtyF3q1TJmFY/6LmNeyMgUIBmAA966
DZoofHjd2mX2Z0cLg2hcjdglR3+r21OwbtKBszpZmKoVSqCmTMwu8DAxm2LnlL0pJZwSRIcBNPfr
ASS6qa+5itEPl6EDhIvJMgvujO3NFQibbn5oiTT7iQKW5UcDGZowp0imcaZlEch5lgED8zcMeqH7
dMsxtgT8Z++HYjAeihbt/wrTyt/AJOB25/uk9XbDqaQVD/RShH8jMYqi+Wgbx6FnaAW9n7Q5YDkE
aHipwKMGF/VPnTlKEYPqlKZ0MVxhMx0iNYJYcHINtA20GLHuR5yVT64B1FGyl94SP4b+9APgzmgH
AgFNSs1mCyILhRIyQ+7kbpoN214wTpLPy6UdOIS+lsJqEBISZDsKDvsAXqfJsGVEu4hltHn4iBAX
vq+CrvPL1KBMHgVoxrahbbfyfc7zd7YC6gpUV0oISJ9EqnDqcZzzZuqjqaqgmyaT8h0TpRzap1xk
O1MnrVqeXo7+TJS1ZcEC9HEiVRDN4rff2BIk8QhjEW0puHH07xkacqCp60Ys+qBJkmzZvPE5swBU
pPBEQ/JV3sQ46JkxS4vY5FAWuoh6X1F5gSgwI1BJgXKcEuuysMOd3JTjPxVwX5ObEoD2wAK8pqPB
TM+Ocb490xq3W+1aOVZ+/QoQ8qDW/TQL+W+t5lvKvPpV2CJ72dXNr4zYS2GfVKxu0/K3jWC7m+8p
4ZuEu+Y3paFc87ra6LxzyyEat9H527UmejaD9wSTnqrZxZk9Nktd8QrLiRkPDPq91MtU1FqvDfWW
5SSAWsUSqBq2DdKHEHbV91i9oz59ml4Yl7gcMaSSUAfM2mNhk5D3fkQCmnBb9qE0fLA0wKDEqImj
kWrJi07fm7S69kGqO9qD8KEAVAqHlD4kdki5BjHOukQ1OILMKUdwQeZaCYtQ7HOa425Iyt5YpnoD
nKE3rP1+aAJEr0pbKEzw6pnk9CO707jBj31mxSwNl0jYajiSE4f82tXBbnsgCo6WRgXiMZeQZHSn
yezC8xscLDuUN4JxeU/bOtEPCXIBxvFojxpzL1FMi/xuZiWMhQWSK/IT+k5Qdoy0JjXSwhPXwCz0
AVFQ8IPNZCjQCfyAmUhjUTsUzA6nXpnIFCNTIg+Tg4/l4Hcd15DHH5Wd6v0hfgwxaEAQnstwwlm0
Ftm2XkENDmKaFVKgJygMSMEinuOcsqJ7QG/9Xl1d/BR3wAdilkS3EqDFHEwY2CoELGdYhIDE+b0v
9VAyB15F06CuB4QsKspvnwLH1xGobkKEqrg6JOUraxu5BTHMWFP12sZtKRdZTXNxJdgnIx8TZUMz
R6vJjTUA+SMseRD+DYzDvrChR98iqFdeMpq8Odqrb4ElbQ179d8YPATpY7JO9RSSbYWcV1NNBE13
reltBm9+o17FHvkrkwVwwTDpag7MibYiEL2RLbTDM41LVI7cn68fJbHNflMcJpQgEhcS7hsWfcbK
O65Q8GJfGRtp4HBTVg9bBWTnGff0FAWOxNjzl3SpBYBAkuZgW09TI5L22EOX3LOzBmVFQjgPfkXQ
2Ku/wawQVPHand4bt3DqtTx977mZEp7W+/18CvRT1XiBR78WNEP6toLMNg68MV4lW7HTsUqbrvyl
hgY7QB2N1nzJcLckYRm/wbFJTNp3FoNRdI19HxnLmqchyfz/bVTL1qloEVH3es2cpDjofUjaL0+m
XvQr/XM4OfJnWFQVMDyx+/5flUxetJSZVoMkZMsXCXBV9WcUlYNkMQIgni33dwo3eBdQu2g+qYSU
ksAshdSaD9zfhxWy0gzLATHc7OmNCe/Iy5tO9JYVXZnSpXswKjydB6MoSVoK3kc0n6UbAs5ID2Ws
Y+si7KIZXBfTovNQgF24cWWVV12224VN0pZYorSGWtpZHCV+cryO0HD29Z4ECjuDQ8pAKMR2QxA7
nsFa+wh2vvtGAjuQXO8jViHzUFGInncoUgDE8sjwe2chSBFH2AeRQx6M21089Foiz37OqLNy7QfR
qpt/B9b0kJ2V4sVw5hcgJI45tAshHrx1l86PhKFZQs8nF0VvxTigwJoFI8jzsrfHPTISkwFvrgpM
wGZrkv91zosAUZHld5IisHXh52aKmiLaUvuYKOEQ5O1v9FbMX4tf/wyGEWFiAgnkmkeUuPn+kHrt
23M0bYDpC2wevchpJso/qIODsZT3GTfGmnQUKAwhUdQqwMWiN0bzydGBYrhfIf0MbZRBlefjkBQ8
wTY1WWhxX0yDYuyDPUO4sEElEoWx+/UNrUtMtFgaMTAt7KOHzfeurQcZ7de1BeT+YE89Jhe7Ckm/
26Y7suvxumtI3UnCkq2WcOpJa6vfmbGmW7tfnHg99QG3s6/P/wSbmAA95MEEZei66Kj9vT5nIfIb
7/rv2xPy+pv/tK2BGbH60Ct9zqP99kpOufTT8S1j1EqhxAAQ0sOuBIe7qPRfv46H39X0C/C+M1sM
KIMwVUNVUw/400DNDIDNjnupJUvD0sMSLc8KhPP7LsyrI84Ak8a47iT78djawIRlbcrsIE3jBdgs
nAkVOGDB6MuMwVhlcoGTCri8TAhA5wdRFjplT3rZjv+Ma0VvSH7h/XSt03tgB0U4zkQoHmR6EqTi
8TJWc8XN/V6UGG72zXNQPMzW2GV3G2YqPYGUCt/KA6OMhNmBDWvBfoOSSqtGsWIZVtJkH8h+25Ac
fmcQutGDbRyyJ4yvnz3obbPJ4iB/ZGBAfOqv0QZHAYuQFbwnwUauxXbINpeQUv9K3IUdQjbLvKtJ
vXaQ8cSkutAbHi4vEW2dOEtpsiTsmDllT/XAmjlTx0c1Zr2Eq1XKwUrwIv9LH1BIGn4b/gGbl5Gr
AY/25hGmWd2hzPBHLLKsqukRsZYQ3FZpEZv8kRU/7SU9XvQMomMtNR0dBW4sT2xjwuGPBsKyxIXD
J7dsGTdChzb68PU2t/7wu6apVeuBCJRRV2GpHbDPc72ngEJuXdXwcRvK631wDvudhWKsZqeCOyJO
hAYBqv8+RAe+SrIFdx6/jFHJA+LD12lb3L7ePHiFh3LpcBlSMixcqP7NXzLDcN9T6qaoS2lGsGam
CxTDSLXlHeYdj0CyrXPhxi1fKDuNRGb5CxpPOkE1sX1W7auybYVF4M7r8E/1s3Ha61Yb36+4wEi1
T+VlYGLCqn5rjQPHCQMI6FQrtlCojx6wSgZBuk67DyNyBvsNSZl3RbJPKfVNsIaAnwAhd7+gRrZ9
toImnlRvDU+Gi9LMBjXJlpZF9HqO4G1ZfrSYGQUqjMnjeM4nT4A38X2mj9BtY6yZU/SE08RPWy8N
sl5YAEWfYPEs5yQv/blg/2ZjxiJo3lM8B+G307EsvVHYTHWlW29u77vAKN9tc8p+R/a5XoAgQrxU
7Azuam7L2FYlOkO+1r4L0ScY/hHHH3gtlUkDPtNjsq2PRfiHC2wjUHgp1FB/3Jf6j4DCcT402FRt
+SDLMUYvZnfRAJZmrpESkJD4GQ85OyrExe8PU4tyoUZNESxTWUevmFUNfUyHxZNy2x8HFtKRzAWP
TCT0O8/EXPT0DmtOWRlTgwqLyBYq01NvFMiJSd4DkXFsMbVAx9pj+dUdC3p21E6dRMbOCBt8NcFy
cOLnA1EP2y3yhL1JANFqvp4DznO1qKUIbW2O5/hFq4AN078o5B0ZeVAUimO6AULdc+8Y74ce/Y7y
WlC0rH4DoRwnYyF1ZYIXkDG93fqoATuX0BHNQEOVMFJW6mssoCXOknW4ZwcbbpchNxspm/0UInEP
pB/AyRSLRVwCT2yUyMZKFH0LA4XLrQb9mZtdf5bDbtjLP+zH0+tGJ/xlA5gOSx8LtosbYQ1W/otk
p84QHSqmQnuJIkatdO9U1rQSt6lp2zX2CQoF8OOgRJ604XOWQNgSHARAY0gOWgwjFouDcj15kHqB
oFqMtF4lSj3KOE9nrbNvmDGyRBUuT0RQ6qNjjoXXBLRgijLhhFMn7jYSsJYSsIrUhHkavZTvtIvD
hFCu5wi5pwBoudziMHrpDUhO8NCYXzMNPnXeq0xOVSMzdeVPx6AelWCm6XnwGcAaYTY7C3XVN7lM
qR6ifvDvnXCm2nj27w9e/knElQuaa6rznElM69Av9ej39TWPL/oZ7ngTXHvqKD0arKgSMQoJu/m7
hxdiWQODtkKqiGPLWPaRJL2lMHfqWn4mmYuAIBDTjzgV7/DpAIGBZYTQxLDwm+XdYr4KaiSANTLg
nwzKNdtKxYTbnQJUX1Jye+9ua9lZcwhAtJSlQgcNFXVqWtyoxm65N6Qh3/1MYjovfI1rFemCPCSQ
wG5XnePxmiVsH1YEeQ/D3LCyMvE6mEq4jGZXmBTxTM/JOEUhW68i46CqVSqyvYHMlNq6+jkd+vEn
PULd0Du79Z1SO1YjXA9V0XoA6s7mRYsjOYyZREZkAr+RG8Ru2g5eLdiawmqsh099FIM6eg/qM5K3
448TEK/dmmfUeLwG6zgo4dh/bdIocSUwN8O3lmEue+CDwzRR6W4JLJVWTWgYxlKvr7EFJEDtOuRa
U2ALqFZO4AjnJUMaZdKEJcuHPUseEtn5Iv1bSvuj1AX2N2xJBexIF7JB2GABTttb4Iid7ckkucfc
UW0s25oW8HLA+af28/UUn14HQarNiPJlBpXO3D0WhV3gIXpa4iV+1LAUok682iQb5psKTrdzOJfs
SiBj4WtvEshOzUmReXr6nOuDnKc13xUdyqr9wCpaanbTES8ne8PhyadylZLCjLda2ATjOADk+Hbs
7S3zS7avSf3RYFXWJFoQdiMhvu8jO+sOcu0x7wkg7EUZlAEZIUdKqWJ8QHVyMASbomoqa348ijR6
kmD517cnOQE7MT2lTz0aDfQSWOx3HtxrbzR98EsTMOx1QtpONgH7BKxtfPg2eyiufBFCfqitOYkN
M8XP3AoRth5LR9h0ec6OeOB6kt5rPXpaFuaYyeAQej4Y+yoYoatMGwS2pTcdS9a8WCeXI8QwMyDd
Ih+1SC/+8OSn786rXYUKUmE3G8pedN6znR8PasZcf7dbU6a9YXlh3usDC6mBQenJ53SGTVhA4R2Z
mg2HeMZB8yGUjVQMRmJHpn3bF3dOlMmsiyQLQABuom/SwK/kv7FVBYtaVXj/SwwlfbGAW85PUrX+
sEzQYbnzWK6tVZstAy4SLtFGmUY08izhit6M3wvJzW7hYIQDE8k33WD2+ACt/4J1AuUgGLKPhcei
G2zGdHyg7K7gdvf8KcRfYrwoBeiahzOVGcJ2EQ8hGnUrFC3KNKKQrFKh7j5EhLdbKxoX6zCcQaAv
uCS/lDUj3bKxhfPzRztBIgGwuH1sit1WCLVGFES3RjIH1r/ng8XkFKG5V61UdW0PZbHWo5BvrX+B
tgV9Ek7NP8knS3b6i0K9p8yklq/3vO7CcCkw7mNwEPCxApt+8eGexaQyPXmZaBV6KE/Wh3eAQWdN
lqJZ1GL5IsrFajHxhX70o8b77VYuC+UYIM2RR+kfAUKrUU75Q4KdXqAVa6uZMNMbP1farOEuyVxn
PpKtuL4MXWXuQ56JBphqc+bKn/I7sA7rEZ6Xs0Gr66q1ybjQFPVpSa1gLfHRjn6pOIMU3tYaBYDe
xFG3cmuORDD8eTmw21ZGaGCN1yPF2R3klP1lZyZeuWu0ftM0z6x4DrSqMFrJgy6GIQd8vJixnyjn
JheKlZPzBfrwzBq7kiwkQrD6qrJNrZVr2PjdSK65pA3BasQUcAV9BR1lWzc41JE5cFzJpYu4n96P
Sqil7a7zR0GYunby/4UjBcxc+jmHRCqZhW4+9I65WSdngkxkCBXvSyh0m4Gy12RJSG5ZCLgO1imB
KZzbj6eZ9pPxwXzckGjq9a+5opCu2frzw6fyAj+HNa1snbYekibT4lIBJxYGFY3bral7idtWhQgm
7SIl8Y2xG6OJkS6SgR/JuH1GZFPSqlcgBYB0cDwjTnbTnQTCz7aNkhPntKSZutCnMVEtwwJ574QI
yWeuIpcWpxbIDsR0vlgsuLiNNEd7srBA78cJ5vKegNH7/FDs0aXLS11Zi86xZRiFQY4hCHjJSiXr
a5cvG5ZApZ767IBBcjaarTHdjdBJlqLGuQlhxLOchpFCJxA48zpQ2XQIXE9Y5s+i+ZU1+Asw+zdP
YTQ3eq6ujoaGJlpe8tgMqluydGmyr1EJ7Zy6E4AhqneHFw4ooef+GLF7pGNDAqar4rZ0LfHTEvnq
+xnOp1AFQCpZ74Ua1rFEf3+JSHjFc8RnaxFYCJ8se2uZjjzY4xoVFEOrUV8hjO1fvp+u2GTdMAfU
63P87VdnvNX8/0nNxroskLQCfaEMYbviXzplEhV3EH7J+rlszcQH5mzzcLFY2thvDOkn+Ecd1P6A
IA85dhCd33CCR8xVbYO1J1G81gyWqKE3Ye5eFtGbxAYaFU+NwfaQ/9Sx8Uxr4ZdAxW/hQzo4Oa+W
1Fr4v4KuE+kEnYJefTKhRWoBD34kZjpUmuA03THbudAI00i5UOm2sySEDUV7sGP46aSmPPFdmWaF
s7Yo7jcSabksJ7zB55QZY+Oc5hZHo9xY61K8HzYaQSeTfAVYVsTkBTxOc4EPxhD5hCjBR6bpHXpf
iBUGnK+W7+OCfJ+scGQVOcp7gnSuDmH2gXVEkBiBQi6W+e/qIgsEZ7zwQFwnb78ZEiOxa9PJORv3
X+2jL5EL4O2VLaDdmrYUy096faqKFXe4axgQT22I5NewblymNLe/z0mDpBfqcKU1Zjfgxud6zWbw
8+XFFgEqi9RgNgoQ99joYKPPZy3+Y1VKXi9+QeiPugaZxBab6L2c4fXNZ0/K80anzi75EtJ1Hxcf
1VXVW/aMW/FTxNKgrrfTlib8qrkBb5bY4zk0fdm7TQxEstJYesfe1uraqyQpcMH4A6ILyl25l84K
2JBgj09dtSbr9OLzKu8mMRVmIeJBqqiZk61YNZCxhGN8QVowdwsrVnJysPSFV0Efad0fzHwrgWGM
orEDQWjKRRwkQXK06f6CbkNkSHiGQtf+VmRvI2dQoxtxjDHYdkFumndYcWrSyfXOoRWdSxvdxLgd
vAe74HwH2XEumZUPOCNPEBv8SnMl0y/689u1BogHDXtz2bkayo4gY+yDNERR2zrG0FjvFPKTokuR
SXr/B38ZChB0hbStLuOLxvVNfKk5kvz3q5k5/cqsbD50IetKgkH/j76h46/319Xuxg30IjwyQQa6
0wkuxlH/Y74BL5F0zkxAhLGqkP0dfYjsH40MyE5jyZtyMpp5JLS0H2FiM9Y1IKHxYp0GzOM7qCLS
JLcSkGFLjc/0InhdAqS+EI/hifpK4hHP6q1rv6KKCaIOjphNKtZuZfZ4ZgUskRAlB5qNsFzZez8X
2cdSj9LaJDuTcHI+3QPoX6+X4BH8PCpkOqB1gT9X7E/WBW0Lt6Bi+2YnU/GSwa3F/JuxoJWpr7l5
N2zffjrfC5D5RnLWPng6OlM6KpMsIxuChMTaRloyH5OaagtAuzNCx2893gUgw84cY8i57ysvV8u3
fXVKa/JqYegN3iOnikzmcBTUdLcNEXoRCDXWrJoOugssV2SRXP1lKUMeIKpzkibYg/Jt8g98ZEu6
QrWj4bSyYxYIPhr4z1FXZ+7Yqv5Co+SwrAhVAunc9pGWXnFaeC/cSexidvufK7tB30c6PcNNOFU6
zmTvh/c85+mxinldcuvVT0Wfa4jmWbzwXBfEFGkdifm1/zokU3Umhc7GQ87epFKywXrWIZCp+6YC
zT/i/LDuozROiIraDI+7KiJFWLn83uI+8RsDJimdf3TZN5nvhDVt1BJHozYY8d0oNDP36eYAtsby
tEBDWi6JinH7tQIdhBZJ8Wc81fSQ5qXp6T++XctBQQEjPPQIYIx9/LyS6PnBnBssOWW7AuLHPt9k
UWlRMiPKf0kH5kFcIlLSQTR5R5Al3tM4Ykz5rfzgjov4+9EbFIb+2V1iIOOd24rxyh3d8T3z+ot2
oM9su92F35DaIIFcQ5IEBM3v6UVCSDBUQ6B9aeRodTp5bxTREA6gop6XD8xewqfkUBNPKM/k7jCX
30+mlpRMgZZdcYHLw9mC6uJ/SH9rC18k6HkHswNBws8DK3l6qQi4UB8pquzyqYCuAqo6xlTRkb0b
wg4vLljpU15bCgpTKxv2oDLaQt8QDO7/5Lhkao4K/PC3va5EBMYV7AGUZcfCKcqE67IX3ezD+X2C
lmsa7eFWFaL4izC78hGYhNMr4hjVg66mm44COIxTM2kO9uDavHC59WjURYAgGVeMptglrv0EzVRy
PbTFqxlIAu7X263WBi0FS9bZ98AoC8AD9p7LWMtqj3DsXvnd5SfRW4BKqCnCGk0tG1HZz+4QPeKZ
/6oD+CxdkxdG92KFdcIxM45iyoR+xbw9bgA8zo30jdspV60q01UqFhPIyR3k3YLU2WYPIlHFCmwZ
PAQZTJN3NkrQWl+4aNr9f4UOdCtJ4Yhu7tgYzQo0RYPlMOGdb/oSPTK0um3fq8bbok8JEQafExVv
FEs0Ebh1oQtXMhWwn7PNe14E8fYBi4hmOdrb4sJEf+/TlG1E9H42XCBUGRNylSwYMjKVl1R/U/DX
ZMgYNgfsFe+hvkgHqsj78HbXl4ljVXJbMUixyOhmOg6CDyocFy61nMeByyIwuIO3YU9uYEcvFRuU
oSjAvN3NzyrjgZFEl04rYloijAnAOGOZELVOu7Ht3x372A9OQOEpkI+eApDBb91pESsmvnrBsahC
XwZZX6iTBgFE4LsgYeJfnOZQonMbihdAzr9Iobfw3K1icDymhXHtLhYQ2PHve0Tft7bH3FyDQueU
EeCBYPHir5knW+uf5kNzRVsGF4SZe6/ZNPPUnqRxSiy18afvFM7wvwaAeLEaBmIX05f/UXktZvhF
mVo1RRYxngnzvFCgyl2lMO9jcpY5PGJ6xmRPsvkHA1bYd+/kx6VsO21uPQBmLz/7kfp8PVA5ANof
qYgellRsrYVExtZTIsAW7BtvTdIeAqvFE28L8vCf5U0lpWMfMA+JbfRh042nJliqldh8MEA9GBDk
r4KA6UXVO0H/yC5OVIHkZQEardRkrs9x5MhUZxwCpmdCMMA08h2H9i35czLXvBY5+9m8un7D1nlW
mJng8eiR3HIHw0xPG5yJx0KuMP9/WS3B9OpbKSS13GSDzImlZE/OkEvHULNBRYeTwQEGOD8CMdu5
WdB72S5rBc1MyA9+1gNPf+igjA+Oeu1iSDn+4J+Du3yl0f9kbydqBQ5URtVVZP+PySDrKjLHlAJ8
ZBbdokF9BL6UkAXMvQQIdfVtJnploOX3JHIdmEaS6Bgez4v5bA2GvnLOrELpJQux5ZdUensJHV7e
BpwLa/1XfI8+//d9OVpH18Ea6HKQI9t/jef7bPoJP2c4/B+SwQ8yfiFDBL9ukNsDeP6JDcSARj3E
OwkBNZgz9QUyJLg582QueknU/RPDYsIfCKM6GJtdjWqOiuFfUsRSC4s6pe5sLTABMVb7lkXe5h0H
goJfggtsYiBZRtugwaNsLjI/D1bd7yn6r8NswINwbc7SEmre3zsU9RvWhngQtNae8wDZb4sfHzyz
qMkXf+9G1NEp6ONATO2jzI8XZVyXP4k9W/8xLEy8KuiaHCbo5Afk2T1Jt3xZC82awR3T3vd/vbJq
2uZF1XArVDzn+eo4NYa6DMHd9rYkwI8xZQzOFjHXs5xY3evplVTI0pQqt8dh5WmQjO+Z/nqiXGrt
WXUTOZPQemC+lkWM9WRpD+GePJcR+aOObbDBdUbnBGxnhQdr7yg1BowDCR1PMwmo1ua4Q6UZhoDY
bHwSIkEY+l/krwLHNbQuopKwTr0/WtVeixI2q1Af2UNmXXV0WbvnVOghJMXAu5ANkL+Oi1o1tLsE
ZBAinb7nU54ld41sad3NxPcOQwGHeQmGzplKZbbNmscQEIed5x+7zbWX3Eoq83vZNYaCZeW4AgWz
+kbIaecO1ucMHx1zTe5NmSw6Ok3+Suzp00E5XiqNlWbdhJ1/6Roknz4anjQaKyW2x55RuRQNIpfJ
I3fajOXx0+spxdGxz1sFFNzg6m7WvrMr82dnGvdAH0VFk+2DiXCy45A+3pt0p2qFMS79rAhoejUi
WPTB1Qia5fYyDgEgMbr99Osm/XnZCZPvXZXRP8xKOzocuanjN8Z+i9LZeZATKN0AMnXmuvy25ReV
hP21dEFYP/Q/5s+YBx7IkzgtdpvkJ2z0vWQGzjpBHewgr29wjKm0PFus4Qg4aUzzMx7TVT9KNR/q
PSivpGAg+pkZVjj4hNzl/m1ADRVoJ0nqLlnU94vwTO2J321btTbKo6l1Kn9EZVDwHArO3OwlOneP
FGTBOkR7oJTfin1c4yu7De4wOQdobkHZVGQx3hqH7Gg6LURqyQQDZt41snBLZqPT8myiJgaWt9Wn
nLpeDKvOe0j1pLe3mvuUX0Cf+PCidxv6M1nchxglgaM5g/5qc6Am9sKNm+43/tCILTVwXlF13G89
5xUCiRKtCOjD6XSPyoGGBjVfWWeraHH5n4PWPSfkGZFRlM+4+JFkk7dudzpY5phrpdtNa9Y9PKwO
gP/K8Gl31B8I2EEXoKc6DzNC3ki5lBlWKzIaM1tt4jFrJcudMzdU0Db7DTinc8CEyg579TOxsYsl
qBhM1F/6kumnSVvvkmIXYxz1RBzsys99zi+V6L6qBv7ZoWVEERn1Mk0CLlBJ9e6DrP765nfNrAV9
M8CaEsgrjsujKQonZT/ZzpKsuud+rvvlkZCeFfRY3b+J6xrDAkxuuCvnTRIbh342Dq293PIa8X08
y4CiDTqshH5BPpdO1jCXzCUapPXb13qxdsUT2AGtRPEjEwLXbtHR18nkqjhAkF1rmJT+14ABltL3
CLK4XUdpb09ofRFUWZfn80sQmeY3GiKU8Fk8Hvr8K/sQD+jcCx8j9s9EzSiW9dUa5Pg8AvkaOO1p
fe/ihKDWOtMr3fPMjWwJtwDRc0WTvrb/giFulAp+bvXkdHDmp/bNi1UXc+b1h0cxGNPE8WLG/MYt
Y30vdSkGCRo38XkrI8olq1QVZ+kpTCExiDLiCQJySB5Tx3zXFAk9UamdDOEgZI6sN5NlbN52GwSx
XQjGOcVPwmJN184Po62xxcPgC4LihE//3OBejMDYw9paWJskJ4E46PqTaUhM3RZ/Zo5DnvbHyf6d
eTE/7XCxMG8IyfuvLTRgpgBS/DwWd1U/Qn/CGgtQ4UWR/TST035InkNOkJ6xv2iSdSn2d4vmjzEv
hyctYVYaN7/HZAqNVlRdMkANrJUv3IbTgasA6F1SA/JzjsdN5O4HBl9VVpLwI/ZaShq41VtcSfFx
keBlW7AWwva8R+VGcXzvSyUIg/Wfthc6pSYVxNG5EniuKdlvLp5Tgcxt3lo0LvIt8RbX+m6WaIXG
Eg2SXfWXJA000w2fqii69ikI8CplZVCLZ8olSaYhS3NpeoTcm243urCHa4/ieGq30R7PoU9dNnCv
Pk0ZxVy3My/aLFZy6T68fiz7eRPf8URBi3uUyFuicLrTcNRGZ6JU47rmcrXugAn8u1NvVLVT1ZqH
h2ho1Q9iMt9jcCC58J9p1ptD0TBaFxj5CLgbk3k3v4KMCodh8dlgo4zRBMtRNd5PdsbueHUoePeF
XRB25/IWaE0erq/3W8VARURTjhY9q9ikr8ZTR02Ju/Jzm6T1Ab62jbDYbmR6unvMbKO2cTwRqi2l
LJF/rAbdAgMcyLcXHQofoIVi4Np5Lpp013usEhweNqXOFc5I3XByH7y9oCoD1cu4uBWuVjr58EK3
WJZg9DIOBePk/WVTVKGIIatc0NQxOxXnhvlgQZUl5ev0WaSLK56ChZLxuTi1VcymaSUjhypsoSOU
3bpwOj/OF0afZsYo1WJWOpmWK5pO1qBQpQf8UezByXcvxSKEXmraquD4Kl0E8JmfFlquaTP7FhLw
vfENPLnJNI+UAXEohwmwiP+lbRT73WE3ouowGEvXWpLYiYfNQw7HO7QjzsMniJPlGQPC9QGryGMv
qauKGCeMrkRM3Nar0uZsNLAok0dY9sS9RvZDm2CChDOCHOkaaZRNn6wxkraX/iGK9iw1t7iuMKX/
a2DMGefP+m6TH0F6TglkfbcHbcL5wavP3RmimN6FKkSY2fhDPU5bXhV44h36MGb0FMzEPzDPCeuh
/IrBv6aGb49r3psrsgcW3OP8cIE6gj5DnCAihx2TgHQM4bPCWX/OtBJ/pjV8etBKBgVNrNhGU3ch
p4HFt3nWZD9285NOH/H1F6cUG+UqxbSVmfjqUkju9gi7w0qpsX+mb1pR/5nNj1LGnJg5RGEVJynT
uwaOjEquJLeW2xDGYa4tOtdIQpjpZZ4WJHsw0wthR2DnUpLbFDblsI7NIuQtudwVLCkRsSZdu1pz
8sFhTsToST07ajvSRPIfCHRdZD93DTpAM5awCJdoe6vU/mJ8TgxPctZuyCIlgjzDNCpbdkCBKzlD
ws3pvpRyj1LPyOVJ4Adz4JXiOednKk8lu1I6iYBDvPjO7ktyS0ryVbYSzGcg37ATsZx7AIAindXG
8tKo3kAYkZoinlSmuJZ8TwmjnP5tH1FIRqkjCHZf3gJ3SiL8KqfsYuI1uilKMYDSfcUS2CNkbgcr
d7Aexfyc+0O9CqAdD+3ap99toU26ZaR/V5CLD+QK+ZSCQRMh1cBA8CN9osnqEy+b15Z6qcILN+n/
L2LWSMTOxmZ0bzv70T82olegBhea5qjCFqD5qSkyOivvJVvh6wMq4OKbldgHak6jkyhS+BZUWjYg
vsSESCw2OsUsOOm5DstsuOj/ZrqyVE4XQ4Rroex2VvgVk21fR8D756NOWjtAYhPf9e53OXk1g6uM
YlPnP1ds6oXh//ssSNzu1/GcBu5jecZb/nTLvrO5GjMQVn7E7zeiwlq9DFPM6KX2wbLI2EjblB67
RSZCbgUDgacZF557GUPlq3JRi/W64LhnQz4o3K49F3uS0Lx1D2ef9PBhXhw/IeEMcMPAW9NLFhVy
J6F2tG3KubASnQrGk8nz4a0d+gkEYOEIbwMuS34lW5xZG3tCUBGSFgTMlxvrgim+cob+zxfdqD3U
DO0qTzbg2z44l6qq5kgxgpSnT2YE8HNrFXjuFqcaMAR1Q6KGRIGeT2lhcUirGWn8NIdBJTkRmOMA
UB9Tw38CTC58fDQx7Fr+mM4SrF0iBbuPpJTHfo31YI84dV0ft+lg7H0yRtfuSdAMZIteDRc2yfSe
CPI4Evsv9ZzZZRSVtvgr7A3LfdWhCwBWDn1hCXnVomtgjyZXqlmpGIu/S9qq8SMgqjsoQeI0FjgY
yEtpHf39bGCo5LoK5JNm7/1AFf4ac5sS/CFopsuywPFYf+oi3uhfCrRuMJpkpE0SQl9m774kY6kY
H9ebEYwbUTB6RdzaVD/moUnq7wU37rLb6E+ALrK/Lsqye9mAw4WS6OJcE9Y9MmprKmcNNxMbG5lX
KBIseurH0F8gMb0K+sAEorksjfyD9SgIBKiq3QoErIkbFyi5SJoW7rT+pqNA5ncn4ybq0n5Axoux
uSla0I3bLEp3zxg3Ho47skWtUvmuUa9ArOq18HQLDwsZHKHuOmg9v+zF4gO5le++HoLWgZcrmcdv
woMdBDGkYzNeR3d35DdcU7YZ3g3qlubTmQLM4fxsfN+pe7y9ilvYqB9HRvVB3lp9G+tdTXVvBovQ
RsE4jCOgHxkyuMTDth6G4JszqDO6Z/m3Mak8rO84llofosyhm3lGhMdU2unCuI2GM9mHRiFhk1I4
LkmsX9wb8lzVjmr919sWzl1qFQPY2VC1nBzjGlebk7MhP272PqKU7JgBvuUY4d+mqpTLbqJhcrBa
UB/KdYYHxJCTEt41DYcCNYDm3AzzHqhtQOTJFPnZkSoR1W2kI+SXPP6wf1pwIWKchapA80gd+NIx
q2eyjNWAuzG+PPam9QbIkTJwTCttcDWN1tLFMkkTD3A4aBXgmOWEoxqsrqp4xY7Mn4uqvVFaSw/W
eslaOHuRAeBQzaCRPQ7LEY9Gj9+Ck7KrwNiiaEmMcjxEv0FTWPE14aZRsIZJsHebW9GrrQC5fDv6
2N64xErX32RCbHgqf3PYwQ4oMmJxKAy1YQucVgboRp7H57lGPSBFfXB17FT5Sxp7bJo42UINKjA6
RUPeUxBltKxScjO4Q6bmd6QjtNB8A05bYUuiokw8CojxPatW9cKNGSXpH2JTUFv/1mi3GOmzouyY
ot07pRkPfOJ8AQzjVvudOllEmHZdFH+BySzFHxHoOdcGKtsZgIk0jWebniREBfxn8YR4cKDEfP+k
3KSz3UQPD0N0Pc//1QV5TJCCk3bzvX70yK3fJwRBAL/kXpTk9IVxOJZaNXKrx+4aQW/Ac5ScPNCl
o3x3oIuU3sv6alRymm+04kT3glVWegE07uYgMuYY1jWodgNNnxML88fbsUihADD5kG1QtJ+ivz5G
Ca10YeSifMze4o8tYui2Mf2pnjHE4ZEYLlTl39HcK3ALniWevKJnUbGTjcUnkhkcw2ANM8pyShZQ
l05050+Jb4b+cfexm4p5yj4+EPQoGvOS0cljV5JGAywnW1HI4niBTcAgldhdHSzaDajJjQviRB3y
q+doJ3Uija1HePSsjUZtzcyPgg/UsPr0WykBDoyAJXYMbTizMhlqkzi+eRMMer624lmELKadhqdM
iISVucj5vvI1bQv7LCVQ+9OrZ+73dWWI6ah4XN9XX2a651WwJmh31VTduVX62VH7xNfcyUkU/2zW
I8kqoAWobWN5VdcKmPeVvXWrkEj1myxz1RYzoa+zonKf8cE8b4zPJjX7U1T6VX/vteQrp4P8pnWv
efJUDucoAGChKaM0Yh3bEN7gQtzSjNUbGANj1XZLoW+Qg2iUT+pgrPcJBkTj8BUFLF4q49KfLJWA
kszPD6pnF6d7gAiL9OtLTeCAmCs/sQM1GJKrdkIWSc/WCnVELG1G4Sdzt+5gdeD0avZqMXj58ZbD
kADmJRmnJXdPgIhgHGsb+20MKAQ4r9sKqbVlmKKvImn0zQWGDTgxBF2Bwl2ciaR8Fwxt/hw76A2l
meFuJtLLfM7FsgQcUEIqRt2bkTBS29swJIk04o/X0gvEb+4X6DDUZtrTaxJzx53AEL6YcHLoIDPe
dT948ajoR/Jn0cDR73CBICt5ymsLfXbWwOaPeoVfWNoDx3I2CmnJPVYGrGQmA2u2Jnq05K57SwrL
cToMjzVEFTAkCdFgaQoCWqi3WsCMsH6O1UdVrCdqI/gcN5cbVB7NYD/muocbNh2/4oxD02bXhTdh
Hj8OfwgvRNe1vzznNchmXTogisSxqnf5Z+eOMi5svAsKLrs2WujHTcnbPbY01c+y4vz0Qdm8Jmio
gvk32VBeJ+y/eDEz9NAL/QOtKIK5HQMbRzjlrLAJhZpkMBnjFpuvTnyizIuVAL8VxpRMDutj7cuo
5AnXB4fWuL5RYdNvRhX+6I9B4Dt/DMQ+6n2Vzi+TJ6eYGU1UV+8+hdsMEa4oi5L/pC1k3uhxDCwy
k3NQ4Km+YyQ6AUKdg/ybQLG1/7127zNgyrVcirp3zf9RmqwmokWbywcXonNgnvY3pmMXnoQwapUL
2YZCNcwdQNbzsnrXAtIxIcyxX5r4Jj0Dl1g8O/IG8BXkDhm6hxTATmdvlIX5sDQYOOhRw1h3FmgE
B2M2Z5OS3KAjZZKbOHEhkqKZEBAjjPa0Ko9eNm5gHC2mFMMlv3ifAmqkVQjgwvLdk6kT/IHijn1m
sZ32RyGMRk9jEPcnAbAa95nczOAjVkw8Jh3WdL4/UGUYE5z5rpJ75rpXvPUUGGDrfoDrQWBIB8wM
SsPC2GwqiYu/Bs3jnFF9wzuGYnv6G2Eitv++400Elf71X8phCd54uYUotCsjuyEy7a22pbuEg15A
cqEo03CD92ixBW03TC2178ER5WrxdQolhrqnYlRoA58P5pkZ7oV1Ng22Z1ZzxsLmmODH90+iT8qH
+PsSFPDvS1xl0SUUZOk6FSchf/wmB6m22lpSoiczEvw63X3HIo0/NXUklDMIJlJN5xdo9DeYoZ3+
9xqgBj40e4gQVJ83ztQKMMdud3EHlF5U4D4ldjh3XFLLv135XvNGnqe2axZPifoFD2MXBgopmLM/
ivTCy/xonwrZqUZI32ORBZT7ok+KOo21//XX+GNe9UuGFYtRyEAGZQd4rdkhpEl0C9J4bX+NyCoy
dRsBVTOlw9lvPmxf+Z5jVy9VOwrzA5yHNi7Ea5qLvAWZ9rNb2WI7aCna1fHKVXqMALg8eyJK0pBp
UF04HswNNOkm15yWz56Yf2MIpr2ulf0WKhD5b/8oX5KGfrG+iSzURlKU6SqKHc6kKdWiEQnjDLym
L/OKCE3ZpLRyadnBtgaUoTo49Wn/nuj0boJ8NJNUq70yX9UCMhRaLNIahkrzMasL63WfqKQxuJIK
zwBIGLVziUzoopk72iai87Y1vY9fABZkZtEN7vr6xSTVpOGGs1JvdlYfYc+aSj7dG0Kowz+yIJT4
Ta2pUYxbt5jEiTBjDiKt9gwg76JrgYkfKt7WtAbB1okXfi1Uh/SrSFAv2rr0VvK3mnY1xE4nvq2M
eD9aqShy0mpTBB/9OvARr0nCk3Y2pBgBqWLpQzhnVLFvWnPjw00fLUSzRRse4iKKm1UvImJL9ZX1
SkZyoQBQy+/lDYB30WO4OPbxrb0aprmQaIjkBWC6nvWLQKi0MfhXPv33Rfwn9yokLqgsti3b9dkg
TRMzvkJVZPczCm3640dxbL2P79marFqdUX4mH3jr2nUYVGnEZa3Z1RurN2WU8ekUwAtn71E1BEn4
+oZXNOshsxKto1xPBN7O+xPw2jp0DDD54GdtrHtEUjU1H2KAOJ9ylxFQmkmy7+o4Vp2yuKmdM21V
O006G/O6yrAbFRC8XxLL9j50ARVC2Ag6QycMBrFBGZBqVehbB/Y7RGOTP2kpaiUaABb8zdEeibwx
x6c37BH0HgvUIw8Yw8pIZqnTlIbT8dQWWVcoILGMDzdoHjnRtzTBfY8Ar4VwOFpyM49FQwaIbJmb
ImjZoj4/pCPFkt7mPYxY/dv5GKLNa5CsMUFFrI4me88tMCW0fQU+5mY0UZn3sSvVbnozOZ5DUoGc
dyK+D3+jiEbiCwCS0xwmBL9sRZClkow5pRfZeqqtLFW27kalz8oRGbzR8SvsWR45NEmr7Ztv9l7H
RRLb8JSlGnXs6rL2yCrJ8qeIR2TV6b8ylMmD+7ps7aXGYaY7yS83OpuVMPVhvV92KV1GF07o7AS8
qtqpeJw3fIOYmp5RqfwhlDG9tnhhahhcd7DWIVjapwZOpEFiF4ruiI1G8CNoei3MLrAMjKLhQXne
1VyaxJQidFA2wQ9Hb/S46+nYtNLXVHSr3Lk16+oPe0xyP+ZmcgubKEo1/I593ZvyfHW9NZACbQ/G
Klv48gHILmth693LYaHtHFQ14XG0CB7wyc20lTrMiOfpdgF3Ko90n9TljhbGgfkE/a81fqTEATPe
xW7zv3bKt/OU5yE9Pt4EFFtM/NjM2BDl7xfqSrkoE+weCwlFqQqLwMTVDDzLndL7jonYzV9lJMYi
kyImAqt9XEFUk+D7pHjwQCVB0VVDCv4IDsrXn3yJ40U5T29b+3n+4EBsNvCwO82tIEt1cCWyugJx
bshCS3PgUXfSlFFmfDZC5QKKOQleIhAAAAFwcHKxvTZMp3jVPPGOqbINStEO2R4DQBGEt3GF6PVc
HN8N32tvlNRMeQQGeGwS3AM+NaF1SQxlFnGD46K/iV++EFO6T30ztLS/+zzNcBu/oAt0S1KVM0xs
PPwC+swDf9+53ZmfV39RoxKVCrQESvgjCuQ7ToNCIxaDTaq6i3shhPAzQeoul3ftLib3lIXQXQ0/
WcGTYGHYL9/o7s2J5tP/Heegwtb9oDtrsNh9Zjh+hOntYD/CpXEv8CbuFgDZNkM5W2BV/l+z7/Uk
RFfQ+pslESkcKcNQS0pdcFfh/HBqyvn2BXzRD4YsZJyb8CCRk6S7OnYlWK24r6ALnPl7Zh9iCmBF
Rwd9FNt29ygJRMmAue7nSTu1YuIsDvQ51Sc4eY3uU106IVBHNx+cyDF5qU7pDMZ0sK2o7qo8Rq3Y
VnvxiM2r+E9BbRIMS06c9ebSgK16pLp/WG0O2+wMkSAJyDpw0SzYyjwwSZqSF1qilTRVG8cHJ3do
dxcTBDgOkV3O8uTQA/RzNybKhGxpq7FDB9NTjwB0/SOsA7b6d5wl4UNZyvyWWLqz3JYVN6+1rRJV
w0uYdzAbT6W2yD/9PHITX92skMP6FP510Rt2deoaUM6ofaZwLb9chh0JnV7qqle341VmA0YV84v7
MmHIbAWmwZ6n7dcjlYAmpq8IQb0DZoSRJSVB/YU7uGNScXxgmRNs7olj4H0tnxCPInx4728+cRS6
qKFWkHZQ4Xl5E53wlfSXpadFTmKbb662pPjzyVCiSJWQrfDbvKGiV1frnMT1VcQpo9CgJUrrtnNG
A9BRyEP+dM49XzgZt96jQPiU4x7KytPeFCCVhvXo1tVIrRBUgLVSC2nfbWJkZqWrCHRW93VqS55O
HZA3/4VznO4eSb/2T4j2uprTZ7sTdbdurxn1BmjivttHiybKddZc/oVhIjBqjF0uPTZKvlZPfJMO
7etUneTIrR6VJ8BIcvVnUMdyLQQHVy/wt2iWPFz96XRlV3TXej4lDlT439vKIPHOV0WKLQ5mlJAB
UzwW84xOgRHwjdehAKKFkRw10kXaW8aOVoR/z10WGoULNzcxgP2hmDirwKHP9YSgtw5gw+NRWLvQ
hv+KfJKh3/NeoJ+EJV2zZGIOL3IBl4hWDcs0/rTgmdJYH1ibtokYTXDXtQXLRNn1lKvmBljZBRDM
HxEQxa7e1Kxqb/xDs/zoC7raOQOtIx/L+Uoz3xJL0H1dkI4XP/FcfWBqp1q2lWU7kpuC47piaEu6
kAZT5y/GpMk8DU+oj1ioKS09U2c6o/32B75qmAoVWFCUby+oYTIL6Z0V+1gWnDtm6yxIsGDm6A2p
TUi0W2AgnkOgnnF5aIb87hotGP2sEWFgo+uBZ0aMPjNyWKpu1bmlZjH3OVciQWX+8tASxWENOgTQ
e+e11qulXT1TUgus6DsTt0p3K+bcKiLTD/byW7Fy7Nb5ynUFqYtE9Pgrxf0wgzxScyOCaCfRnH+V
6QTz+VhgXap664NxlJ0zl7D/zw+ZLIOR29aS5NZmTBAYslb9fn02yp4D5Xf6BRAgrbJ9Mr0B9sey
4G8cl/zclTtxAelFqHysF1SYIqCJsF6FY/5SvFJZ2e/051SwwWSO55GSB6ObogxmIVSLE/ONlr2g
4tWFB/zJmqWsVOGlvfKpsnE59otb0D4hHrnQ9eKCxYtI7yx8KpKy3fIRJ7+x4YxcSebv4RX9gZnt
CozEDsUJRiwUsB1jQ46+Gs9sJBkVPCBqCI2urYV98TytGUvq2e5TABgSS+vZI7KEAaw1I2vzmObL
GY4pak2ZnAW9rnLklpwFszkn1eWGmdEVp2z3/L9aTlPR+QieFGvbA0/Mj1I+xVJa20S/LcXuUjgt
kdz8lm44hcQlQ7eaWhbPX1T+Uf3656ubuV5PuQoN2CtU4PsZfqIIOOdg4OgdvkBWMXAQW8QOY8D9
wRbUftwkqZYUwLqOEaN8/PPjc+0W7jpSYlYSCy7b6UV6U/qMlBvX6cfciyPU6RH2ep1KAEnHyiIn
puD8axrYo/zcv8PdYtErwIxDK83RgDj+nO+YalM4HZK6ou/vgw4HF5thrP7hjMqedrNwVe3lOAxl
T64B4VrEdXcDDIvJzgtidnUeW6Pi7ZGcdp1oihw0/9+8CMhFZxRrD25qOqF+58PyjgzCcSjDith+
Dn5kv9CUO4KOeLwBsqvoyY7Kr47VYSMbZCqn5xDqNIsyK+QFVwLk/7hdJKzvODygsRuqRs0fxymF
32Ku39DEWqVHYyL5gX75wWRpSaFCIysYnctnwItKXUzPgLrZN5Sp3If4T8DJpLOHAe+dq6v8zssl
cGuThFPaLnPU8S4kmLzTI45RO2YTPCvitJkgi+bidiDyTdmn3g5XOh6s62Qah+uzNmRsxcTAOKKY
SE7U1U9bQl1SDtkAeJz1uimNLFjsy2UkFW8JYJ+kLRQnwAmE9IVazxZnuNGshII2rCnWrPi6NY7d
RBs7+E/IzaUQWBud/1ZN8tg9PIH/bmBgoxS+qmg5s0ZMWfxavWtnynhuVU+h4Lwm6wWZRinBHdrM
DDsNqnF+cgS4wGBpoIKz7VLTbdTzm51nt1f0WhksTheT9vj1xCJ78EfZPi4KeLRl0ug9lr0rOKjm
mVxMOhWlH+7WnWsaqJfX4B/Vy5oinSJ1y5Fr/pOxeseYD1tl+3LxyH6H2MBJWQ4cSDWvfdp3cODh
ifB3Mn8zPqUIVr9dLFP3Jzal3glX2fclPbpS7YqX3pY6fXhUvkWMKIVDwLwUXoIMGmGN6ttHfVmX
17ZHoJoT/2y45+4+Wb/PrswXCaeAo20VTvhQhU2Uv6Hcy2iR9/NqRLhgSb5dMhBJa29bjJwss0W8
rVE3G3XqxC8Czb00ocY8kE6FcKwg3pTnUFNNR+4duJ9UacJWjlmOwW16rvXm4aKCkkirZMGc81a8
gZ5hgpOBLAFLsD+p+RDXvkzsLBPAfuevyVmA0CJeu9xsu4QYBybWS7d3LzOdP/8umGdspNCpU6ls
tUkhxFeT4WGcr3ojn6EPQ+6LVcFiSt/luKb1DD2QQ6JvkgJyilGTvrmS6Indhv0BiI2bK+mQMtGm
Le2MXfAS8ohMcvbQma1Sn4Iw1KxBvgKydt05jdbHx08FFgIe4QB3rsYYs+x1fxj/25a8e6cneTKg
uAo6xaeVij1sth0zhthDSPZi2u/azErDUH723Suin7RcavHfMkXkccHmLq3bBIsAQjkIOQTK9gbV
Uq4WUFbszz9KZXSh3fhxg0FJtVM73QQo/zW05HGbQDNv6Nlw7JIoRVLu+M9L8b/Qoof039GgeVPk
03EEpt7unREaXHCR+lFB6/c+UV4Xy+LOrO/GjCZtI9JeyhyyidaP0ZEIeOCxtYuQbXJC7a2GfBC0
UvVo+soJf00mkgZRVoUIuV6beN+EMX0rVAh5/g3vYkFYfHTfUYu52zLTIwvUDEnaoo4vDsXzIenC
9jLkLwcpPXz3YEreLN2tQkJ492yRKCENQS0H+Lrppd1RIF5WsNSvqLBg0j7ee84cxmbr9Fwi4qSq
+tgRc1+5i3+a3Uwn+v8kG/hBzFOSoEWVVikcpqz5tsaMX1GXUGKGaCasqsZ6KZgAawH2BHJnb9h1
eka2TrW/7CMYyEOIv5b7EoHX7bUTzo8Jc73+cvU++Bg+bH1Xc4j859SpHvOV9NyzykwfDMgdenaj
ALmkBB6FGwb3Ub/lZ9C93DEtKEULt1/xudyyW450FT+NiMCNxy2k1hvBUhibmA/6rrMgInR+vhV+
NqKIiP5p5UAyXaiEhfbuLKvvriwbCNuZm9Z0+b8DxuhXY8/3tbPdloilwgiJsZwui9E+RZO3DYLG
/Bo1tA+3SzdUDgDtuLb/Ui3EgF7fzfcf36VnkCsmu8X99iFPwyOcYp823M0BR+9C7dSF1upaIbnz
K3Jt9A09TjRd1GDWcRVwGBMdtLstToMCpUaf5/uyHFkM//e46rJ536Ohdrx17upySW2gpV5fD2zJ
zBk7y6Qe5En3MYpBN0+FokLvc6NS+AQUGLKqImkKU4uE/+HuW2tagqBdrxYY6t7GPb9QZbImFzMW
KdW43ccxytwjd5n6BBIiWeZH39jB1Wc6ERoCnfGLLg/urONPIldmBRzZozdTPiytA7wPssSPjIoq
cRsM5bDGz4W29mDljqNbAJTLGI0Q+bmPpCcx6gPkUXBX9kGw2wi8w32/B8hkpceAplJyAHWD0jAX
boAoVR1VUkJBJIw/mo9NbGObWSl9nYYS32B5AyvHkXWRK9dTZMnandbr9RzxVx/Sm91v4UAWq6NF
RhoUJdgpGLBSLOdZOA8vvoVqi1F+kBMEBHHvfVn0ovN3t3Yrwz5t3iTUdO7PffAefuO8qKk8wTNl
Dt+LrUZOha1QEyt+Q8r4MSwy0LxuxdlPx2CAANOaWu0Y2pqmQz2MIafjxw+RXL8pRgfzqH6blvn5
qve+1j3eowszN9XFsblO+jU4EdT7d6gZRnu//JWd9FRkxZ+pjsWfS3SSWtWlvIvAQZQybpTDX5xB
iB9ly5JiQoL85ksvW5PzL/v6Knyodwxv9V1QG37oX/2AGDqndj2RJvOOou+2LU6jgBikUcOb65Rl
45CpiK9RHHynG0K3OB8akXg0WaOYIu7XhiM5R5OuyjoYQgrTalkN4VpBFs8xAs+1nr5ZfUzh8/wy
1BoUTyQqyYENAVX64Uqo00sNngygvDQxKma0E3GyotXqJZffnzsMmHY9kOU5IjAvxhPp2dB8I6o0
SOvkEvcCQSu6KfAvL8gBMoPl/G5a4l+7YvpkHvS2zm4Ppuc/BcfHGKd6iEwOChadhZXgEIF69krY
NUgZ4EFRsWqToAyAAOBf50cV8LqsHvF+xc90gdeAOt8dbeZe7wDNHKej8CrJynGw+XovBRj+yHWz
axCZe/VneLW8NTGm5UG6gzxEpocRrqm/acUiLA2yrAXRAzCmKMUaMrWiYOxzUoXQOQb5ScLIF6ek
4me78yvRJC/1DhVsLwWiMmgwxbx74yGdwoFH2W1imSL2ovdLk3MM1CWAmuk2PP3WKcN1Me32EHYx
1OufUlImwQeTFs14h1DZZJjFh3xY55g9J6ThXMLkzryslTWE9XVovE6SbXz3GODAdU1wuS0vVVDR
QpXmLNoyGaqewLtyvokktaMPLLHCGdiF/mONY3FoDveuPzI8r/UP0VBaCsN0maP/zYA6RfrhatQX
SVV3BlqnkslBU8pHzD5qXd8WrN6YRQRcDgxFhgxmRVPsMU62eh3YDrFURS13Mtfn8GlBnQwOvN8w
u2aBKvHX+ObsjPauJnZIQx3kgdp3dDqNIocmMiDQD91RP0IuvZjsmRtunE/qhe04UbQTQxOA5U3M
LE5ZXM5nCv1DUwD4pEPvkzKfTqU/P865fH2CEaOkSallNfKUTa+6W0F7ni4/COtOcg3VBoVbe/g6
LOPa8zFU1hXr3ovuHPgJk8AIjrt2O+2SSTvDD/mPsK7usj6J9Ls2HU0v4FtXYuTxBe36GeHzZHEg
hAIGcabhCtpDSYd1Gq5cnbhRK4Iw04Nk9Te5R6lZ7r0ahmes6L5NFlcCAAZtV80VYuZlCdQHZa3K
Yp/WCJ7XWXPTxWelSH+Il2gpsVo//hCydrdFmSeLqHHx1bQnIhUHSLIu28kXsxe4QTYzwdXHnx43
3Mtnq8lGC5oxNKWhBSbkH8wuxSqnnn6krlW4IZ5Z98oPIyJmaNaTmANNQz5mK5OrnM+zYgT6M/LZ
ovVgW8P0IKiwg7F/xBq1krwbfbv/vcOK1db9RUFlOD453x9hb67zJyKQP2SWVDDX0h25dIRnSbxb
FJgoXDxtuveHNbR91mf49bC8a2ic8530M9MGXCgAc05X+7CSG7npYC5KM3dWPEMEIsZyIjZ6LRaX
7aDrboUfr4GbmtedhwJBQk07eNJNcAnJCXvq8rIeqgd33pgr4LRQVtEbbOP8VMcjI6I8gOiTg7vC
pDdIAX2ZhxRVF9DzOF55ZBG+YwtWKnPz4OUGxoU9Gcp6/LSXMP39pRkrNT2WP6mZYtuB6Gh0oTVq
ydnQoJq2KADxa9+3lPCbeFBeVEvBG5YJiEoURNy/z3dfya9HXYuuZu2GiLYlrzTkT4UNljUn0O7n
eQcfMbr3LGLInBI9dnKLZjVr4VDrRbeGF6gOhaJ4QS28SzbyG3iVMH5Ap3sIEnu8duR+/tFOOGeO
QnhA/vYVI3OVjgEuzf7S8O1T+ym/xTNbujK1vqiP7Go5HBnGLhfBoSRXuSvhgb5kFvmpf0v8qDbE
YoEFwLV2fvw4zfLNo81vOHilwRRnm67Pl2IhhsSelBZJwtDWXd9Jpr9oZybVfqXkbshFWpB1RLYQ
0zUi959qpujXXhnlhchAf1t3clQskLzeb2OuM9ep4fVT0N7SNy6mioT3Sg36kshE4Gi6do8/XaLs
fVBOq0rii6dCXme9zc7kho6dhfOkdg8OnVAJRm92FgpRWdfA8KbWQRC3+6C0MFBJcVksg92Ic07G
z3RAysV80LHC/KfpfpLyj8fK3u7NkjForvD5pEChRiruvrgxesw9zN2iqLE2lG0iYZvWo37BouBb
gtXgs/djL1Dp6Uu0UAEklo9Pzh1ktpHskQ9eyf7OWNtxjzNmbZ0GCIxvpcOYukYdwbFo6AgxlIls
iRh5Tn+b0vb3N+8+8R4gMRTh+v5tpCX+/w0WThgpLmWfEUfji9lDAaQxp+t6oGT/JB1O19YLK5lT
ep1XZwkMEu5JW7J4HGJz9lTlxSh2YhOwiiQeQfLsNoNbBGsUuNFsF3mQ8UsF0JP2zsFGwB6duj22
lglLx+cvk59wSB60bSqodHXdGrBUHr2HgzitdSjIGFaG4DfNJ9S4oeTFFw2TMS9ZR8WBtem4kkqF
ESfYF38FUjlwK7yPTh38+OmggJz7Rmc1TQEUxhQa6sxX75gvGaeORqXAy+Oi4jgSeUmplHuKPn+c
sEaDcdnHzvSHwoO/W0urF5hGvRr37TUjxy/4u4t8o/nibtSHbj48/XTImTonBrMzMnplq1My6i70
gBjPn7lLEl1pZv3xkbIw4Lqj8u9dV6fQ6Zlnn4NRpoGhI8/d+lgR7keX0/O9jz6fmlCT1XYG4YTr
BJriB2uZkjTyTXPqpoWjfrx8Gd6tqg5seCIL82gEgNO4B/clecW6jXBY4Ye1PLx1UxvNj/Zo89ql
s1wMIxkjoy46k619Y8PTz7g3VHFxkKqLfuB9foL5dZVD3z0fwlHiBzLgJWumfH+KzHSAOLr6hl4f
QWlx0e7ggki6ya+FcHtkriBZvE+8UfiO4CIlczJRx8FcdgocpjfjsbXomiLxXqeIIsv4Ba8Xjf7D
ZEj881mIBm5YPtqn77oqEbqm8uMZekHviB5K76sgWPiaut5YqeSnCIqM0bDHAPNZfvVC5upxjnaQ
YqsAIOsOhPm3Qlrwbazdi4J1/yZcvP4sra02moCPVhDSJ9J4l2CKVuzp6SEYkWjLd0jVSSdjilix
qzb/3NGlQahaN6OtXZkE9Innb+EYAVyy/r56kMmUPBsEMQC2ijfyKWHPTLZkiG2R8h8bOmudr4gw
i3Bin4bsCZlbkNvM2Ij/CpvFPcLMJJJ58Oht9Js7o/vc4JIS7yUwHAsGhU13MnmFYQdTHTW+pqt2
0J5GjME0ewrrQ/GvYxQtV0fJrIVP6+W+aOpI2LTSh8LNsE4UvfTPb6FYuCCmb0piNz/4g94+Unef
6bolIiF51smGrdG+WMo77mvezFk7BlOmYHIthKB+sLXjKUtLPMrtvq5ac05h7HUSzJYIeG+BRDkg
artHCaEPzjtENS1M6ZrchnlmfTGZHqQoFQG2stwfZIEPqRt/vvM1S7Gil2YwsIL6X0kiTat0UEkE
tHaK0JY69vCfPHhj7AmD/VEllTmYn6GVmAoU5a73hZWpoinb/YI/APwFNGCZN0wR9zXrbyFMzzBf
AMetCpKlEzZg6Y9xYZXwdOEIhaFTYWf+soGJNgT4FX2fwCcIuNoxpm5GcKm9OU7GFGoCiFLCsl62
nTjexH2EJ6FaWaRBjSEZCEx/x2AURCrkB9dv5nnLD1ZiMy0s60PimUbzZeba0ZQsTc5vtEya/63q
dOyhkaXr/kw9FKTgZQj9muvC53ySxuZvcm2ofgTHYg8/tQkFiANrRuHaKu39ldr5YvTrqv8Plspf
QGhoY5M4ZryOmRPi8TdiMkf/A9MvmFXWJenGJTqUhLgHSMKFl6vr5XxdJPI+6MDQORq0bJWN/RVR
bIY/bc5mxqMkvqcmMDOoI5NkvQs+AmVUsAeg11NUMRNoKb62NRDZ59d2rAxeeHcUzbB4kECxPWHk
TV3P7JsHElB6V4eJ1K3zIKMK3yR8yct/tALbLv17wXOvRojerbvjM1lQ3Dd4bFOKsqiCa3aanyqb
ES9hLUjf9hZOLQ6pQRLcO7ZHBZROwXtAzNscpuNAh3LkmBgYLXxc2u6/ZD9rT/2ZcmMMQdqZE/8E
yGo03zA635QeX3nxt282HNRUFjeTXxML21guMoHvNzbnquRVPAsG8Hzalp0kMh8Qvimj54lNFD6f
fn4eTj6WEjKBsvi9QcDBH2dWeVn0wAwxACoHE7Jd2pet2ztfaQENjtEpm2EYH8bPS1y/W4oCBoEm
mnXpMa81sw0fBpIGw62qJ/9y6mBhlThq1sEOvddYhft6e8Xlq0KXXT0TAnPFz1kbtBUMMbyXVL4I
ufUpQoDJG+K+gUIE803ZfwUZbr++XmkKE+1C/ddz9c8BfpUC6jGL4m7XjzSMH1E+wtGSBbey4LH/
EX1OIOx24lx0J6YjMnb2uuiL8T1kknr0qGnwGjzSheu6oSLtmPXCSfpR3+PXqkjODkTz4BKBSOZ7
WqqodDHXocztT2/DzWeu7IkQ+GwskVF5nbt+EmPV/Wk2oHPXviUrfvhQE5tF/jgqrz+P9YO4yKnn
5YuueIeZOpintsNhyeUAGyp+3gEPUCDRCVsfXqop6xuxuzhfPYP++0DwYhXMTcsQt+Vhby8FnUZN
vXJAEskK8Jpyis6LleREaHVvQbS65K/oJxhY2gIhspSSvbaygcDwDgdccLYYPUfN3qRyvCuPHw4N
urWezXTty+3C9kYnG5KI3KBSdVFnsKMwkScE8xatugil4q5v8shL06ZD06DxUiDW+DOWGFMaZ9kR
WFDKVX8BSoauP6UAQkPunVW7QicHcaa39ZhPvT9dBtjEs+cBuqD1E2YFDMgw5ZkT3XY5rJBnSy6C
nOL9h0Hm73c597a/Lz3YvCHsj7x1cgpJOqDKBKS1sBlw2jPl28+1XMiP3d3BHlynBDg3CzctfDVO
7X2b1wj8hGVRspQqV9T7c/DeixRnXoQl/CPCYTS0m+AKpA1pkxapFKtMmQmSVtf/GunyAXGKUBP1
L9xsE87s4PuODgqBo2cmOyMwUSuNvGiXzHaMBU8IXrrFgG1A+YVKP0NHefF+1hSojlRTQLeNxBNH
TfT1f3aA+2GlhEkwVv04RlpBbLIRu9AogQegO9iL8eUKTRFTeBBGT37A+wToYCzBA5aEIWDpfTj3
iMiYUzJrX4+C2JFd79Do2bqU5Q4LaCl/ItbAwLrfa7YcXHByKeCElUceGvU5Nn+hFSekfXULyYGt
B6Jy0G61Dokzrhy0l7nU7Cji/Wb2GUXH63dVip08w37BPprKmyYf8S2ARGRnAG4QtM4N3XlAJsfE
2dU+5GwtohPAKOmoTGA70RH6X0uCYnCPlZPZEPgEMlNatmUnuH+D1OBqLyhI7pHUcutpkIDv2/ep
8ByEuddvYkxFyUaZnCG1F4QqWX54/pNYIf1Bq7rj50owG77sTJ9glFDecfwUuaXOCnVvMOqpsMBk
fxM/lDhdY7IHUdwoSOkoHXCXOebz92wsHSUO5O/suihkVdfk55WX6Vj4YBddUi7oDjlbR0I+n+u4
mYBWGajzc1jChkz819f5NyJ6YqB1TzbgSbzidpDBzYmIb+XoYa8zDhz+bCNrkFIKQEAHi2o/tzlE
jETmo76S5K02crlnBc5B/Yt6MR5kuN65audW4yrGtewHvhLeloJreyDqd/6qmHZFq04iDsetPSpN
ArKXYX3PzH8MFSqsDEPucxzyesPfEvWq/+zgs5S5U1xgAHn5D6qeK3DM74kztfl3iZrpS/KYj1dY
71X1OThSJsw0eqdQ3DFPSF8Jhc0YDbZe/ueQC8STAq11Z+QnI1JrTDnHeESHt/ZHTkhfZUH/M6mU
ljVTMWyRr6JjIJfGt1sD31FpgZbXMHwY9cxSIWclHCHS/Bxl5suzf7wpfJNg99zHnYaKZx0d80IJ
r587wVmIJYQQOkQHMGCAFYiA0s4x0y04oeMit7W9d9rDjCF9qO13qBkG7weAG/YRRR9XAm+TnS4b
qXZ6/mqxZfnXG7mF1VUW0JuaK8Ke2T0e1oyHxffoeuR/JXtiAh0uN9uPkv4wa5og7gnYJoiB/07p
8m8sVkE3fvJwqkjP5bMbNh0oOfuQYIHl+wMQLnVswsKhds6lMVQroMwURjwXGtERsujmHipqCf5b
PojKYSp1AgLJcZdyEBEBikscZUzGG90LCIiPszGS46+wz3dNbdJqot9+dxV1aDSJfU77tx5ydNf/
Io9DlnQjUouR/o7K3UevcPvtXx5T7rQwaiBCtbQ3SPQ7wEaOk4DVYSxcr9OGlLArjxwH6sjFKAJv
O2RzEoUlwHjyP2dh5feHIQOXC9900POSPwPmrVoF5LWlXV2bBFlUR7Sbgcc7RfBDMWcCABsmd985
8UbTFhORcIa2iiN/viZSXmnV2kuFzlxm92fiX8ymHXlN2G/I4bwJ/Rt47JwUWlmxTI6wFrdcSEik
ns99EA+wkhGOLGp9v+s+vGDpfu/Px9m/tBGfN86kH5nLf+BMLOdOD3jQMKxcezRaSpMXJ1PNx5tV
KoDdlc/vSBROIimBFrFHlFARdPX1413IKi2ccUtkoVVeYzgxf6uaC16ZTwyj10b4t+zYTo+bWAMj
nIYSQqiCHOWOjiV3zixTRzjgdekc3p6edL5UnKesltqpeBeL+MD93OswVOjkb3DwLxBHef9KTIiU
qNjccH/ND2HnkcwXyzm014X4DNJ/7qfAM8Gf5KvLbvSl5YIqMzv45CpIbVPtTpbg/NIq970deZo9
T581HttLiouTk7VZ6LYvpZCzuKWspB4AEcT3figXOX515e0rewCnDTK50cA8yIK+wGuQi0XgTdDn
1BuHSTsfhDnGOusZB4dfQrOSeGUAGfVcEiQx4/lnAtFDu4yb2c5ICR6SfYUj6ooN1sj1+x0p/sAt
FkOnMqMGZN8Y0j+YG3QrzLIJtXxON1vjLYLJwERHnzozJnKU8/yC1+UygTa2fzhTLik2f2tUmJgq
kx/hNvfUl4QHWFMzbk52tlu9cN/B4G968zETVEPjhSLmwiI/3fKpdRyBdIVbBNJxc+DBN660JhV7
1ce+t/SG9Am3GEdkKK6VNlLkgUs3StLGpoNrqkWStN9kgOvWZfNgNyfaHtPHa5ebGEgfbF/FOfRs
gTFefGgcH+EQKOPbA7fJ21c8OTvl9UOZuHecqvGBdvU3xziQxwAMMXuNf/Q7bcux0uSR+r8IlVUW
1FC0gElqa1o5V+YbmEDkZ5LfW5wz0mjN3Pb+ZbojJ81uJxRTUTv34zBqHjJ1vTZm4/9P8SMpOfjI
soFwJ7hb80QoiqGrKwkdz2z1Ys+KsfhrlFCftGxdOLuzt0RiKCXDWSmenGkGAnf1iQTu5zuLbOk0
sqFEimmnvEdoFhHNHdvxZLMEMGOSqBXO1ubsL2QFgwYmEoQ5sPundL0qza/5G8HVzD70mLioUuvU
/64im5ARcKV6fQN8BeIyuyEeSmBKZgv9siRMawA1Zot4EN7Dntvya6ZpMP0lHm9MTpxjddAGzTji
1VW1PjrWTal+hxPOYC+seelMwy6f5CDb7BFwPupW9xS2VfGU9INypBw8J9Nz8o1jnQgTnw1p6/4C
UWtK3dCRl6OdJrcIFf0/r6w1ekidCp9Ns+jNmWH4qnMe4Dme0AMmoBpuiw2WnAVtLo/FXm7MH3OF
U+13iw3aJ2Uu8gsJr/QNgZW4jDeRGQWdhBuVCDgkUM1seP26CSsc6jz2HbEgoInwuOxHwrnVd3U/
MWFZHfNvnFGI97nBkKk4HKXTpRIUuoDwz3pXtg1FHdbO0RlQ5AWvaApiBVyF9cdGwly1wI5nN0yO
iZuexO8UY5fRZVXKjvn1I7kYTEy6XXay5T02hqTj/JMKf49p2afnVYkZ98389r0f5nS/UkE3Wrpf
ReanFC5ZxXwKgA3zLjzmKr8y1tckqMqVxU18BQA7ERXfdtxgAOP1Yb/CxxltnTmnh1KnRmZZjS+S
Me6xHVsHnpMa5pVU9hwxZCX0MfAbTAgGm4TAtaR1IOlT3ypHCKEeEhG2+rVCpAqFTAb6G4ItR1C8
Mxm6V4dRvIw7Imbd0kW5lIck1K0KHjFGHY9geEWr5xmCK3UCOVrMN95cM7htXcPt2kQSijnEaTgd
KAWaqFt2Drk4ddoYzptIt3CIdoF+YwGYvP55Dt16bdBZfN78xzhB7jtB6MwnCNURfgujCF4dt/SP
NXHf/ZnowBCjM6gg5ydF1s8yuI2thVreniTdk3eM1hjVVFY4H1QFNx2sndotLYozV9EP7/rb86VJ
dAJ7tDbPJIOX1yTJN2kvyxh2FNnuCupTl4RGq9o1EuJffu9ZkdYAkfQvOiPskz4i6/oH9ml+XKIj
0jgwprJX8DPrNiiPh0McKj2Rk/laLPZmb2FI541SC/ZqNfCucEmsE06Q6JMUdWYH5sOlW2YisNXo
J+S4o9GBNA1IxVhL/VTAtn0QBtGZ41X8syjSlLwqbko8/NFQs6rB5DXJL/zecqdVVnuK6dJJX5aP
pu3hU+ejQO7pcHmoMUHEUmAwD9GvkiRn1LTAST7LAzVNcDY4NOmhiAbLBxtvmLTAKvT834CMsNyQ
ul8NArN3vQWnI8O120s/O9HUKT9zfCK65gH9tj2+oWdlXOQXf2u28AFy0rkkdCqw4H+pOUzg9g2N
BxvpqP8J1scmR3a2Xt9N0EeGJue143ZKxNEkm9zQ4LGFvwHNYR/7+6ZiswgKJ5rlm2KGibPVxd7F
JjioFyzAE7O8QBqoUldg5yi/5w54bWqzT7EGLUwcdDnwXb/VBoEiZyZzEkcV8eQVu8gjn37D0GW0
rGY5bL9clge2SxScScTZ0aN8Dvp1aY/mT5FXGDlGY1eZY1lC09vsd0lJi2i2iD29FRqawGwtktKL
v0jMvbvWimfVKY94QoztcZIVBAYX9rzADURJ9mAzzGCbw1WHrAE91Ithvob9/Twn8fo6NsrQxFxF
3gIswKvBKyAVmvFoWHS8FbkgI0m8dNKHOE49fQ5vuROxISebWBZJNMYJihgfPGTzvEJoIAu9AVMO
yezbNFeMs8EPRydRWgVNV9GpMCcIjLHsGSLdnkOfoCuIZD7XfHZx57a0Aq9UcK3IO0LNBE+ZdJuV
hV8Ourynn64RFnnDvRR8rFBRQLqZ2Ba6iWmwOzOo5DR/PeecDmy3bHRlP2Z2pQgNmEHBXnGlsUi4
bBTMaNqzVFDq7Mf5KUmsF/Lo+TLeAWn3FZPfKvKBfywAusxYUcjW7iNroYisXIw49zcHNBP9y9bF
7CM1YqchCqDnlEKj7cmRwcQJdUvwH8NyQCJrIvfpovG8iYoOOQM1GhKq2VmwPTzwBtsaM8mEReXK
WakWqV66qIBXNvoWX1hZ7L7FGiwJjHtHxgqkTZvYa2XK4JqIsSFb1kFqnbI3jk0W5sehLtS+Q9pe
KUFssfKY/JApEgHbQvEhMge2qg01UeynqUHypw6auVun1O6tCKQRTRMlY6cPX5y1bu0hP19XfgtX
Umpyg0sW4Wi0hGZn4qN82MuKVSiTNQ42E2PpeBEGU2R8ciG8zB4obtAuxadxv8/aK7xT8F44CTwS
eaRgCIKNqT9uRHapRJTVmoySaLLVREKseCL8r7Zjg32vnjDBluQ8bHnoWX/eZqAFotpMTzPixUtO
v1S9yidmeNxaf0N6J934o/8czRQTUw84297FboKpGQpQve0bkBvrCZJqlI8J+FsXFBqIa92G/ynr
nJPDKl9//7QlKWhQuUtD4CuF+sDu1G7sx4G1fdK9vKxl0i24JA74xCOuaStl4003DzBs9kL/W5sr
p/nlR0RP+YBWmjEra0B0yv+qkdkp2N8wf+O53ggJfkEjFkPdG+it3dMDQuzirpc3z48azie+vZCO
eN3DT3o2uLUDTsqqsrUDgK1JbvTuFqT4VW6BC+Z7LTh9ub21lHxgApD4sw9pZJ7jpGnhfH0ii5IC
MHXk3CWiOIDOIFphLtNS6haO0S1TSRwAam/912DgB4nKzl1BjlFjR3NsHETZr4LutseFogyaGp0U
W2CgJMuz/8Z+HYAOMYTB7w2DGjKM3pa6328cZJKq2syQsF2aI4T+GbLXUdTmy3REvo/cXOtu3Lsw
obRDseUOC8LhHRgTJalGxzLTR26W1rECN8v1VAzhD3OPU6JOSSPRKkKyRy+kOBvSBiD88RKKA4LM
DjFUoZIsl4ty2cMpoukwZhsGcfvR849V5sAa4DujPMUWYTVZjbf39nTfPJi3bNtWCYf7Bc46N5Xg
aEGBAz5TTx9JuuEKUyulbwV4Hj0uDU/psmQdS8/vIcQvKGnxDMJ6po5Fk0cN5JuiJYkcvLvIncWc
yV714NLoI2LiJcFjNsD3NfysS4BMvSXSSbdrDbW3l1x8/EfeVso4D1sTi24YyCH7KACTjw0sdp9N
Z9EE9NJddvLDBDPpXFUGWNykX68wA02kGF7bUHGba1kOj9VOgkSFc0cCYjoEjjYiJHwhXziRHQMh
qyZZasa098EsdWCrnMmCbAijJx7pM4p+VZM7Gy1IEVtwn8TpZKvFU2cfFDYN1co7NTlymMSoRoS6
UEvlV14ttCzDlkCbcJNbJBdlrWgG6WtbQSY2FB6LMDkSEGYb6pSuCBRYX7wlSWjDITtpEgbubzly
OQYeH78TBRxjV+la2blZMqvnphzjPic1fFiI70eenxnqJP4Zz3WPmzGceIodKdWQLgu+psibh1Y8
C7BfT370GIJXebCdQXftFnWSsiXKb7EvcY/mDJ0XT15QQEnRCn1t0zKvqI6rBZBgr/wx3QPJchqC
dGqF9AMI29TCK5kthFqo029PoNJXr6xJP+eskkGpuUp7Ird+by6uS3oPTfJczhlCLIrTzvAY4CKa
TDQqLo4Wcojw/JBumNse5JXRutKKfOaQCH7sfYWZde+n+5qTQ3RaldIm/yxTeZLKmSKKQYUxPWcH
Q6iK2VKG1IffkBNVQeSdaYH/YksEtpOn0t2dL1FWcasxIUAwzhu0kAVwT0YVeOfLYMLxxAHcp6k1
fyTEsYN2dVPOkAJtF53vB/0p7lFBUTPBNkdV78vPNGACU5TT1qILxXXYyX5Vhs98mIPqVhiNl3V6
s121Kegmbra9KwO/QJqYOqSKOvpIyMjKonSSthAc8/4aMPT+2hwiuYAtaZlo+pAQepx4+nLFvwvO
WkZWUNs8S+v34iq1pOhTP18r0rXU6iQoO6GrjRhgSjs8at8daHiX0NA6JJ3v3wVh1Fp2rFc7UjUo
L3vUhaPm6ZpmvvZ1lGPpP1N16jkr2EyHmTT2UMu4mBsT1jUn1G23rJkTUwrlHg9zEo5Uffi/IcsN
HuJrASl71nDPlfR8WV6KnBUBf+aOmUKsBAsAkdbCgfgJbutGzNMUiDpszqy5xJtiW3r8xQoJwx5i
LJHgeXEvL9xaSQk07z0A8J9j/JQD0HLkacpqtI/JD9r6c/PtFrI+I/1UukSUXSLlb53T3tK3lhUi
FZ0VOeWay4G+O8Rsvh6xU77vQbPAJPJQ11sZ09/OE/ukQ4ZJGJMDRbF3MGdMn0OZGJcNY3NE3cK1
xXn5Gjc5CjYCM0yB3gcY3Y+p56RpOmsonyii2KAxyYbV+2YPo4A3mDq+iXJylteaqJrQ2BnrbXtr
Gg3sOF8t7C1H1RDTz8ucYtYNYhx5/+znh6dezO76ghR8H+FHtcIfrF6wuUAw2v7FQpRQ1lRwJ5kd
wclr9/oJ7f0LKIEiKqIbM/Caesf8vCHk5SK00KFeuBGHb831ZydrSy4bHTpF02hs+YemmjzEWwvh
k7VMKUArm4NQuI8W8vbpSNtvFVrse59t2+X39ZBzwuksloSbkDy1gI/9kPSxyAr6D+gH+OqyxGrW
ghoHuRDJGbCsTsPqjq9s2G56r2BQIVRtr7mdX1YtD/Np2DLyZa4mT/pDuDiTj/XaeuYlbBy+y7D8
2CZOFTzYDlTOlSACZMWddQ7256Ox0BUWykb/0qHbFsxlLtYhPRJdk3EpTEl0Ljzcwqil3KcGtnF1
IX3SLg7eiSbiqu9oVhAQ/d4lHlI+nfuFwNSB7tWUea4mJDh4emoCDQkYYIBvXVYReRPV5p/YIOEY
OBbu8Ib8VnXpnr//bV2o4Ron60ZbwwMGGbZziA0NmmOOPCAxTrGn79h1Y4e1inkgNgxrKn8hJ8/K
c2xzHYktEY9N+43UCrxi3xjY11ZdMf8fCHY+HhPU20TfIfd4Y949aIc2u1YRz2i/PjZ/+EWlc6jl
qAh3OEgkg/2Ww+1BqWlX+Rzualav2IXj12evEIox+2x236fQOkR8MhOc9U8mvlir3BCeJmuthulG
bpiv++AmIVTaX9Vft61H2vC7V0fIG2FZpLGj5HRpIuP4w1Y1Vh1JhdECiui3e6it9KYmFQ9fZMML
mHvf4mr4glpUT6m2J6t6KWfL53tZ+fGluYq8RBtXQ1jBZ5wXLAjg5TKsX3CqQonwK/Ib7kJrbJ37
noBqmDPMC8SoQPCYjAleHp/tHJ0Rh+M7dzfYdle70uxehJUX1i2d52lIYID6fBjjVymek/Z1obZo
EKTBrNDSNQFIIFLC51EJHtlApZfR7UmqvDwKZEwTBM3hoJKGecLu/SbWrZCUZbitYLiPwwD+4KGH
ugJCKt168k993yYAIBflXMwf/iUM4bk26h287aC5a2Wv+xaLWT0PcRQT6SRPJ9UC4anrKAwGau4L
yD5G2DVNbWvgm6P9/r4iiTzIaJ2oEoPkvdc669+7vjjOQRod57cFT3Qk1boFlQhfEqBvOq4ooxEV
Y/oAJuyqVZv29mvq5pxK4UbifZPQJu/i6C6/A+xFctx1NK69YSox9Hsx47ncaJWIMZ8KhspK2TDH
b/MuiN/yDsW/2mt2vMgtWyv0FMY2DVqtyHNIrkKn4AnrZxbKz9hCHXgM8No/IwKYJrdIk4j6aRg2
76nRyl9uptVbqcadLkIG/QNaR+w9fpBMRUhCIBk39dA4x3gXdb9wThR2wc7eDc5jXgGVGqmCR4yJ
syk86K2WgGqXUaBjWNh1KvVyTHxynumJGgeNtGBOa7YnQ0MbLr03nhWFMipNjxhogFFQ9fkH0m2E
R9ZWWxhIauvPtjzhGYokAiVjkNRB7cTFyxFMcO+nzu+hLHYRYedMEOvQ91AWbqvYd1bMmaFXxAQu
EBn979XMcsDUo148i1XCleV06SjVIJ30qY3nS0g+wVfGRvqU6iTBZRPbQPJddHxY8H+YTzOKrTBg
oI3lmZHq4eE0rzbBbRUBSVIPKlGn/Qz+7l5e86bh0vYuoWpRyHrrMSDs1yVeukmLl1O5Vl1wGr+E
p3kFOnO3DUrITZFIjtxsMGRz5ItyDBr0CB7DDgT1m0JC4tRlVVu2yN36PUucCWHDG7BhybVhx+5i
c8lz+f3YbkOu2guSMAKY6ZWr+MmefFpsvV55PeEp056nNegd1MV2k/4v8cg+B/ty/Czg3oDINyyn
LtfEzLFqeFrYjoaUolKBdEsSHEIhyP10Nh3RH17J2MwEqgqx7rw3JDDhZg4MS/HtZdL9qb6WhRqK
dxYAtzxeOA7NjPdSYBiVAIINJMx4f6fA11COb4tul+nFDTP3AMAx+KwEeyiMeSu0yBI9Qfh0qjF0
wJz9NaJeyXMmk+cMsGTZZf5SHkpERuRD4xXh/PDjDvTUGAg9gUCuOqNxWXDwmoWOXcR0SHrh6eoE
i/1ivM7OqmVjl5RyLWSeLgO4ACG7uBupLmpgzQsMwmHaeSN1T0hZ8O5SHXdra0QSLqsHeFU2ZL6N
dvKV9LnKXoQkxCCP/82A5T3a15MHiX1wjxRPmsHpQLGLZK4mrMqh6Ej48g0eT/P3iTC0XQRFYJuN
qNEqbEzrrfxdXqJKXIp0pM0zsZnYIkcFhpwiQ9V9kmxdtuTfszhnYoGUeN4C4Zaxf7mR7BepJr83
jwHLl5gqmyxX4QSRpfQVcrQ0/5HcHI75Xp6gCyRefhBAPEJk31yOmntHI8Vw5fsJED6WaWEFyEnV
ZbOmz5QDOyarENJiiMi6v22cH1sQTmFm0bTEQkRSaN/k46KenAlx4Jenx39XqSMFifYScQdD0LB0
kOYQjD9vXmdjhQdb1gZM6SHuAnIgnP/vOd8OjK9Ol5rPJnHxQEJANvg8DU15bQNhVXka/eWTP6SZ
jReNfuRlcbk/BnRzOv6dnBBAWrDfOh3PfCpL+v/4Xf2lpbNkDMUzQTl0ET4lo7W0O3sApRu+LDXY
cBDuQ2Xn74ZrlJonOQhh5SUG0iHkBYVz+OIx9M5nn21TwX9eUCVmsddEKuK5sgMfbxNaPvSEX8tP
ytDlnzv0Aufi98Nk89nfPToxVHrzyorgpTjx3QRJ5XhYCmk9E+x4rquNoln6QWw0iFNah1F5GIxw
R2iINGe3rx0qXRXhsxg/2Tih7Uek4fvK10oOosMK8PhmeTW/MrAdb3IqzQ9S2dxIopwm2sxJVOiy
QoyFz52tLWWQVZl5R2zsFexdja7+sOBmCufTEZc0WTib96jm+YLvO5EQ2i6n7KvN9fsyEQskmJl/
UHPAdaSqC+WAjYZLpQO8zbWFduE3DIpxVjSvFXQAxp0LDoNlCfiWFNwSvi/QrjNaJDkyn/63pimp
b4ilqrpe4Kev5fkqOxUTHECuV/dNfELpKA3LJUXKT2CjBZ/qdz0H+KxOSu3WozTDFV+DTcQIJevW
Z0a7GbGyhvosEcQWPEs+mfKhE8zkCCdZRVdUcNcnler6XGeXX3mrxtOH6R2pPn3dyN0rIjuPcMsf
WnrpBaEDnFs6gxt5ICsv3Cr/5dtV3iy1ibkHyiWqRiofn+DxHu6pakRfhrrNNTc9Z358xiihaffJ
5jzeU1xh2X4EK0OVPgRzmWRRC5qHUnloqeNJgyTcTZJeNqbsMhWh5/qxFxGIKJ8bCZHOE5rOG11L
6FmCP1+R/0+lTcVgqQXSYSRHEGrsQ5cWP10SmB8xn3J6Vbp4Gy8WXuyYMAc/VuWKWPEW6gt+28f4
EyMtXFHkajIeG3q9/RlIpdgD9sewXDqYbpQVFgDpvFqCxO5D2+BFPo1NSGNzP3TE2l68WW1PCNAo
3hALFigzae9VtDaA7o0/ybEjl+mxXMcnR73ODhrGfJ09yxkCEwSco4PVGVKiwapOlgQQoXZySKI9
eKj2GhnZTu8RQD1o2qBR3qZo2uQACZmn6dJJgHSqImLcfalFY5oPbPnaUO6YqwIRNfwDHeButcHG
hiT5lW2d6RtV62e9Ky2iY/GnYeUPdEAdz427C/YvrLljkWxMdL8xSBY2oDWsiLiiiZfVBqHXRJ8K
D7xqx+cB/98vopVZNO4yfmXLA2/gvKgF3zC5m5MHVOE6WkWnU/tX2MCtHgQEe6lK4FNmMwhfPEZp
NBc9ZTWCFf2ItMIKoE6tgNO7UND2AT1W4tNvTVQRsSN9YtiNWI5umuj6p5dLg4om36YC3EuPwZ0m
ZdyYNeyeDj3sy1AOauv1JJ0c4rKq40snZN2olwV+M954U9A4i6FknZk1Qvdygv7Q7uTYbQ0V45q9
Y0EeBVOetUTzxT88sc00k3VyEmHt0laMRYpE3zvDP/mHFCgoqccXdBDLSw/2exAAdKEud6hv2O1n
qIlxuj2Zdg/pjUWodOdTNQ/Dq0GJOivQBWDA2qxVKFDPVOorgRxvH8bXXKgD4rD7pJRIxn2T7hb7
Pa6SAj/DTxkJCltFxzU++5BaeUr0sUiW5LHJEiNAFrOxNCc/3cCsi3oLyHElkodOvEXEIfFfoLZk
wdOH6PhExaJ+V0UiJjxZfIJrJf6YDHf8Z8L1XMi9/vlhwGHu7ip1YRFy3zoTrdKQv9qgyvm0tXn2
ZTN7ttvLuESlv0rW3ROZSiofJ8QFAd0gJ3XShAw6edF1vmsxkYVxKYb/Aa4dedCSOBbOiYfWW6Cj
Vo4Pt8mEQWyPb9aVjeGwr7XIi8djveTfBmFazFg6rpH0Vi1BmRtfrqTofKyK2sqiTr1SSWNIevAD
xdcXpbpcIalT0bIkWyaaccxpuyQXgcMz9o2tXqFk/iNzPxpnE8c5thzw+9ZRXfHV4SpVZo05KKY/
nZR1wJohXpmpu3u3+wkmpBKU2HE8HEBIZIYw16+fi2KcsSXFHDy6TbS44vSXRBGovC+hhR4WIQHa
/ayr0CKYPiP41v5BPiOlHEomn2XAVppO3NnRh/ZDSuFfnASUvCxMFzL78vLkg555pO3JGwnqu7Hu
ncsj87eLoIDXbJQvOWEEDm99pIBGnFRdCu41zl5otnIpGXjuN3XFmHrDbSuJ1JUYBad4xtROzTVu
u8pFPFMRuzKl9X9R4W4PDRcC847TDB6DPKyVBMe7Qe5PUnqwaNbiyVzfuMzTDBY0oqgWutPIjLSl
y+UnrPt3mSsxFRqyGLsUmriu0O+LKA5zP8YEXrE7P9BV/RFiBz1mt9Zv3fkHKFM+vQltnkx3R4rQ
NwEWfd4suT3VfrUnX8JHq+53qii4fmnOmD905v0zYF1mveGl2lfxatgzUVgZFK6h93jvf/WP6EXK
4zCJPVxF9wv1GVt6tM0bdTYRmQFd7tMC5w8VvPMPLkCJyAo83LNyyH2wwp4En0ghj0M0iwtgnIPg
k2LTwAoOfv3zPS2tpKizmVUF9mao4wiBkYL9RN1CdjmaSXj9bZK0uRWo81HuX+Gx47SVm4Hc/w10
j1BtW0kCu1Qm7AynTdqvXMonKmfcRVezSb6+eTKnX4bDhgIjoEBE0Exy4g/H12MGhBRtIKivnqIS
7fx8Hju0AgncyndPaWePWfyG9Q+bzjT/+tWu88HdQdFqkP2KJ5yYMIAfSFPGUKpHzAR60+Y/PLgs
3hpoZg3CUQTNymQxMWTam90kx9Mh7F9C08qg766yHfGB+ARNmB/e17ycwWjw7SlX4lMKs1/pS8Am
NO6a9iHhFHd3LaEZzyjhxm7DGD+p4q2Mx0BUdHGIqR8n3RAc0hbP7MkocnH3XVH71kmJCT+fAoDp
BMaPQM623U2flCmXkxhIRzGHTYKKDqR5tmygm8cNAgTvc1Jvk26saC8aNLWEyot+7EnXezGpijmK
ZnJi8bIHznBNmy37UxkioX3EaI7YAzjpZ8KVgkDOBk7O+MZwmMjMIieX+vkdLAs3rlpfwlYO8ebe
LITzvjhOXJYQobTOJUpFWHHn2FFSxkzBY4N4mnxqKOpN56vkSZxvKaNsKM8+MmxqVdYTdjSHqXDQ
cqQ4RrjGWm6MHHVsfFXp1Q7D1LWTO/i2rJlBoH1ZsEvoS0Pcv5Ro7cS8nRsCwKaRfJiKJjY9X1VO
Poz0JXohjORm7mVptX/FvTarWTLIgus5cRW9XSN5Vgyh5jUv5CHun8MHIcwdvSmoCNTVFY6g/x5f
sXe6YflEiVInxBEZPNbMaMlhHBmmbZerMWROGLuL5PcrLe39GV1Cp0PpZZ4jwnhEK5igeanyKodf
aC8qYV9m8TLif3bmLQCfpdtlJSSTQrVbSorhhxNrs/b7BoW2lD81q53/9laKtR/eaIzxoPXKUmue
l5kDUH7+Y0FVKhFSc35z/MXfiqoHy78F5IM77zGFJ1f4LvG/Uhb71VNjcIw/ubkkY702ibpWJeVW
KxMAY/MFJH6urrXQo6ii1+j1g/J/1ff8IwgOWwzfy3CWFSmIRQDs8pWSw4X/7tXy9tUwdokDUnB0
9SZZgXJWaiNqDmxy2JsfyMTDrCtQ97HCU6xWzA9esjA/1cfUJT0AMFWWZ5rJ8lOyxZExyscSjd1d
q2txnbJBDXYlQkmA11Qhlz9srXjytmufggkzMBqVQWq+zjU7ho5kdHBDiTLmPNFrIURjjYm7BrD5
D2OyqZrwzebakRvrzzcjFm/ylQ8HCHTr9vi7G2sgTdkUOWGdK458h20hYm2ZjFeIEBSrhRjBAxsx
N2d2ZUPXXcUrmrptTeJUig7gaj+c+ZhqyqTBWF/7tkOq6i59lgQ4Yyb2owv8vFgaWK6Wlh2Q6YA7
XMrI1IiQGznO8JxcSbXyxLcaG+YoU8rsuNSn8xUyD+dLb8FmWH7lUPdS68JIUZNq3i0/hK66wdxC
erNKs9ff93WRmZhyeCrfwmPmfrVhjAwKTtkUAUjavbNyNeEe3eup7eWpS9fMN5qY+E2RIuEBVaTJ
/+Q+Wn9Ng4Yzubnkz/9M2TKKtrSdHf7PG+vfhSCSU8jUCBlD747yxb8Hr+s9YnXpDICRUs0iwjqS
2U2F/j6Y4jwXY7pZptuDK9t3ESJKuP36UAZb2lS83uH7prH9xRmS3A4TzwzOgDVbrRp+k5w6EJDq
ClPqd/IpvnPEAmdEri1C09Blefb8MKzX7feqFZ6DCNXlLO2yr4pyq5jHUJ3FjiOyOsRmnohLFVOp
ezikXqBN7CwmgktH5bv01Jj2A08XsKOxdMNEk3A+OnexK1pM52ZKHE16K6D/S8vZPNGNQrn2+E1S
GvIpFaxCoGTD4cVFPPGUndrpvTfXSVjSOEbJpFXuOxKkVmc2h8KDbUO+G9kTE1CUKeyfFTm0gmM8
/pzO0xxxxDamTReEWDDIjsCBuXmuEXlHadzI3E0N8H0m2AolKX9TQxw+94p3beaYxro4DVjfc1kO
PyHxfVlTsS+nKTiJ+qu57ea8x6HMRa0niTtcgiMgyWBDslQydPt0jtsYIgS0Mz6BTc/5GbXAQK5b
a/Xvieh/iYccxNnbmxs6qYtLn0FVUcXFGKwtE3JAYNL7qDlOp4UF9eeuZs87+mbY261Nvlqy4C6X
lLfqoUmMJ+OUXnH0Y+0jVtXf1rJ2PdiObN2Hto/dQ/SQCFBbalbgMPQhS1KVD18ltiZ//JemSCsR
CyitWlRGUZMTB0JZco2ktp3/udJRop9C2EXGxgxZLvJKQMgypJ3FSE8keNTaXj5GvvjdN4GJWu2j
xLTGmaapcYPejiqBJRD0QE6N8soMY1ZzSOlZpXtrSRfTZLau677OmdRNxX/lG6Ixm6R4j84X5C+/
4nBqPH6TBqPF9AA/QGaaZPap+a3GmmiD3FFhPPaB+WHD5zaQiiUmHs8jujxk3pQgGSpeL2NPbpgL
308L9RvVkFxUaeIztbGtoAVZRH2hqBCfimSfID1B6nHC0l9SRLcEwtR4y6uvkcZR7v8WsWKxBNo2
gYomH89dgyZFfWFEPO2Sr4liOPZfhP58QT+gQpMgeVjEfJSTR8NIsDPagCvkzoZY7P/NBLlr/1hg
K/s1iqJAZub14UQVzkoA6QwGOb8iDmfiLwluf3RI2gRBAzv93uRS5JrfYw2cE56kb3YXqFfsNlmk
mjxBxmY20ydw/pkryjQcDCeRGPh0upvL6IzUTdSJvXTqSTkGnUKH9IvpFZrvksbiWq4HstG2SqHh
1YkcWc+vJ9Nr/rrbihIVTQ43nMB1gxMcR0JoTvGGFESrxXvx1ZPFEtWvILEm7RhWxyvZo4zoP2t8
XRdO7UxuJiwKJBjc4abwFpuI3fsWBdo6kKJoNnZagy5Z8S1Nt9lCC36nFV1B9xnBCI6HVoAQ6233
0F0qMtQkehSgZU0uZs4PH6xg4gK6n/wuhCGeseA0ZNrqkHW09VspEw5VImwrwLA5sM7JN1sbtkgM
Nbio6ROlEXUfXct6eIzLxZiCP5/8ULiGmRBRlr9MndDO0wwqT9xtdcSQkfogGcFiajT+zKTIOnii
ho0Z1RmPP1EktX8GY8CDwwuy7IZbcXuH/xeEir0EGDhC7bF+0Wh7v7xqCDOiAKcYx6jsp2hNUTbJ
tD7z2hLdBpm7wsMjAFx06kle9fN8KLPUHLs+TwqeIdiNK5VH67IKPB74HQ713QwOvmiMh1JN1Px8
n+0/9I4AX2N/15i9iX+SagDywsxSVYD/2qrDcS54Y4s184uK48ZR0l1dfIW55+Dcp8lhFHPIb6wp
OZVQA/urZoybQOIKeEb+2j2yQ+ZbbO/dtxG412Ji22uy5Io+eHyW9PaT9R5OalZDV1yZvM+nn6eg
YAnQEnHWGv/ReqWvW5itAjEJiD1LGGrd+uaAbp+nSlCRihbVyc/BpiqWoERj2itsK0WSQW7KqaOG
TCf0n0U6imACNfchYzTqX3pQbZTGMI6vQV13XBeM3lDDUX7CD6WvZ7a9Pg6Krq+ISaDG2bLc+Ycz
9ORgZMSUr0zj5XjmDa6bdb7phdefFkN2ApBAYTLudw3XeXVsfjJpUPxuHP7KXb1FuOsCqKaWp2rA
nz8DQtS8tqtc+dJi2Pl0lPKTfGafyYsxdDg4l0vlsC3ktr0Y6QFoM1AqAb3/a5nRS5Mi1uc5wdyx
2piNOY44j2KzdPLL7tLAu97tRqvMudDoM0iWtt68FC7FQPS9elC23Ep9mteI0hrVBxViYoxrf7P+
Ao4q1+43B/f5ArWwCC7J4CKzP8aPiJiGvqgbhMXV8yrOgfS0Hv9bBTY8S1zGqu1e/tSfqiYdTex7
Z335GFTuRpR/g6C26Avd058Vgu6PeJNYjpf+XXIT/P8ZiS/IJ/UP5VDdP+prL2hlDsu/OUnDGtRa
Ok+/TtOiCs6cYLvDR8DgIeARfzm5yZRSvxJYs1JW1/2d4+XahuES2i9FjMppMnaQ7rDb+xAkgLE6
K30AKV3RkCC+5Yw7TDzwI5aqt3/Dl0nYexA498vFOgNWWR5IGUr7asKy/axcBB5PvEFLah75O9D/
HnIgwbaeeYOkiv0X3ly9rkHIZxpR2OKh4E/lUafKvDCDbHYJLCmymTUVH7y+lGL3W5vmrEcrQogQ
7QSSx62M5yqpngy5U3oIF/L2WCT00VKwFRg+wft5nVJ81Tgrbh9PQIrFfodNjpQaV3YkGibIuiQu
qtJfS+lvX3qfXWN0VSy9cppUQ+vqRUAtGjhZ1ufuFw1p0r8BhJaugd6hPAudAl3KnW1KHL3rxiXx
GI9RoVc+1vC5lTRlYOP+RF5bwKNqCNbf3hG9aPY+mPjDMgbxRbYC4lLqLt6/WFntfHTVUlpOP08x
fbg/j09HPZOLMR+a13Ixi3O88ShfUbqVZUUj6hE8my3UvQ/GjWrRvL2MPtqu7GnulBQkMZfHHA6s
/725kvgcoriycxKB/zItJojgim4VcmXV3HcZdqrsChNlC8iA3dPRiG0gseAwXqZ4i/8LWt9u2FkK
7OGlKClueV8sywKwzfbskuIjXqrV4V/RoXNwc9pJBnU4Wis5LoqQItAPlbK0nB5PQ1EtUIOpIFc3
iaDQcYvE+pZizKg+GG3y807ffqQG6KpycoGtKENtMjqE9CtML9F1XhrbTWHkATsrgLQKuAeLkSMf
L6ZlVYrAu2whufgwTXeYk8R3WTdsIRHMcDIwOq0VDuxhbtOFVyd2NG4loAT1Fc0PKtmm8Dce3Dh/
mvIWwIhctepirPpputZRj0wOUjDQyUGcV30Ezp4ESp4Hw4csf3VCixLyBoLPBrvyKe607mTJpm/G
M2xcWvGbolTQANt2PKfLmFIb1Lai0TvlWk8BQR+AgLpczlevVYq4O+x9YCBxh5dUTcM0Bprm/QGJ
PO926to8ElQZ/2/HuhCCg6++gX37u6ogyJubA9b9T9AysuIhErX4E0SGctO8pUJ4CMAxdlXigZn/
/sLCum1xLbj3u5XWf+e1mtVQnqiuxhkKROfZonIK/Ix6/ljeJ9Vxgka2GC2VzmZJ2lq0IY2FAtQb
72WfDhsqZvPPFaLfeyFrT+JBR/lfWBMuDG/2DJHWhpH8aFeSnYi0iSDUrtDpzECO8FUDfFmW2gJY
dAqpNf65sWnHJri+2sZFTITP+JHHersZzNHgA5Ez0IKGZ1BkGzAMKOzu74H1yp7TmKvEHTzq0hM4
SYtzv/lwc0Fr4Oh5h6xOGKx4ukp1PnLULDIlrE7vqyOjFs3zOHIvbolyMwhMegoZ3XE54Njhs0kr
URpicWf+UQCNAWQJAigRUJWE6LtGSEpo9gyOMdgUIx98W2yJyiYwGQAhZ75SyVlRBjEg0rArxygu
VF7WJ1wuBOITwFYjPUe2ARTEGhqL1m7cud+PTg68szxStwuVmXj0pCvl5h/hebjGoYbatKxtsDAN
nmI9HNzY9HETtyh4Hu198MS7Ewp7QerIVfi6/ZsQwValUCuTuGFogVq5uCeDRoXb1VaWWDIle/s2
eJEwKxVwPdvkbpGCXnoqyp4X8MktGbFzknCDvfIzrsOOz2EqySTmfIyi4Dh6SYO1toJu9aVplibP
yWGtLzu7NHl8360KLKYLJGIlIBB2crGqoeG/gTkOq5crFF9LyXxGgpIxEHJCYinchX4R1tgDHzmM
IoMDN7cs7mcNrGReCaJlAjgJlorqDRtHzD4/EOq8tgDofyl1JPCxxFhiNKsI6cG6gOhPOfG14KQs
8TrGz4WdWGDgItPpU2+3BsTAAOR6uANB+KU+ssQur3JJoKB5/Sa9jRAeWse8ERV6xKW/gwZhIxfX
M261298e5o6G+9woAvUGCifasvM8bSAEdVEu7itBr41Jjpl0GCBZv6XbMaDW/GMQEMNXUF35L2aV
KAWUPPLMR/s9duz+rqirc4V75Qv71+zlbajPtRKPMSF4hzb6Jlh23eXhJ8BJ5zEDDV6N+65YSXlP
mPmviW5bIQuoXWkDtZM6/gHu/v59dXmk5/AN1KKkyWJrdfZ1ldMwOIHAOM+8fagu0YgbG6bGLpzu
hAaKb1VUkSr2pL2WFzuaalkm+EZxT3ompeNORC/xnDMLf6qp6oCTBRw+CZX9DcEhcm3PqI+K6v0e
xksvHJxRvOXH4dLgWauaV1XrRZMgMpmJX6Wf07sUxU01bYg8AST3eQO1rOK8Pn4i+dtItV8WppyY
jL2fG6LENIpBv9J3OoBzuPbwDmmf37B6z2JJPyE6IP8JYhmTRs/3e4Nh4r2k39QwXwZ2uKu68LZO
Wr6Be0aupKW9bdsc3Fpg0oeZZFY6aUDvLXvO58HbCr9si+AA6BMEy8MTkIio+OJJP/3PnLeIaylC
hTxVxFgJbgx1XpmUeNCrKF1WvYFPSxetV1DJG4ngmZHgTB3XA+TslzUSe68DiXnkIb6cNQbp+cqG
MyCNn/gdHqw29uaeWxS5u8PxLvqVV/pGcNLLJvf9XFAae+bSvWuyV64UIiX5RK6iTfm41/4qclws
ZXzzEIgsBIiuHm0ZPCxrRj7ZgZmtDbq3+NngpeVa7pVY4f3H4YlqTo7YqfBLIPk2cZi5yAYQ9NPC
KgYy/5IXGF0SLXlvRqc0qXLHX93PUMNp4tOU4j6T3kSr/hfqs8MDQVYnufHTrs+7WyeLNbudIjnp
iAExY0awVM4XjmiACD9JTyD8oLegEYdYI3i/dZwiVoN9JQN7BYAZFcIr/qSuEwrpFcYLG/7m5UTe
rmNUKmxcsaK69cqi7twy2Sd7zNAOECB/NScPtz5J8IAsG1dvX0JF+H18gP6YZbEClgnAskRRRvY1
XglH0NGzk9CKHyqj2KdPqRY0QuPoq4ERYXZFuIsV3OK+YD8RfHOy/KVX0k6q8X+9/UYGs4eq/8oI
9DQJSgl22XWwlgsQvW8CGxPcxL4de9JrlrUwIx9mGeXuP0yJ6Y0+ro4xeg6G6EzwqGnBr45KXq9Q
mE+Cxjx1BmYyB3WFo9Z2SuGg6G/Fq0rWv2i4sYVrqZb1UPn/rTofiXd8GYQ8zwKX4Ns7bQrI3Qdk
uy6KSU+ahJ7yoaFS3M5tbyYvPK8j0zeX7/FIBJ0SlgFzdKeAs0c1SLG7w1n76FENcjKeTdu2GYuu
wJaES2Vn+W1Ph2kIcuvBezbOJSQ+ula1UscnOnXB+hO8L54ESopYTcmelwuT3BZMAzapnzO8JKTj
+EGe9ALRMCUdieeGtrGzn4Z7LiDtS4u02hn4mjWDAlSyEDjUJGgTPwusU/QY1HSksW8d2TrRNK1m
JRImuEJtzmhLx+tkOSzJnRwZW0FWreVRd5EAZrg97CM7Xk1rWcWPcgHdLee+UGIo7z8SKqzKVxy/
GxmI4HOcXmxXExZwOMS2OaEPz9EzoaIQP5JjS8IY4TSHCzoTdLR2nsXpQ5sIT9B4vImNHh4p7JlV
cBouyauPaxGrUxo15OQZE9x4XQWc0WrUSdIuzu+innhPDPxntjcwTCkPx9F8RXFF4uOEamuWEPqu
qDWKsEmZsfNstOLhdYYZ9IoIfp4npVTPhAZvIz6X4+dXy5o5e+kKfEcnXt+6TKgM+U6/Z1Ogn7yJ
5Es8lfWv8btJ//MIb7xmupuQhnuvZLwGXbnZw1ogC4rBS5B6KNcaB1wPOEFhKb9MLdKHU2Ahcqu0
gfBKplie9qjPU7biCzRL3X76M5IFoYkbQjlp56VVy4i+xi4lNgWQr/wd69TqHfxQSIJgwIuAsnzu
uuZ4WQyZ4nCP3QWK5IHnaJi5Gt1WL7p9WDJ9dKmva5v18fDVJPshl5NhU2sxVKcD2K1/jzoJjzqD
diqnXNMQ87PEe4pKaNtci9dl8JUIF7Djr7Rz54FI0W1hggxeJFymNdW9HVfmiK1Ytmx7tcuwgU19
+g4O26FYP5QxAzmQXI8zxNOOPuIG1bPN0q55oRhPX+6gio6DwN9qwdVNJ9QVhvQ4794iu5XJr1oR
KTvkECuf2V91TJs6W9kqJ4GAKeHM7yKW+o78mt0pNvUXqK41a7h5g3zbndUpxrQ5/2Qre0hnSMAC
ZKb+liv45hFwr2AocCjkSZQ2HTTlXTWXC4vTMneo5IH+JnAggytkJHh6T4ORPo93kGD0LHkwheck
OAwZB1bWuT+RF2CGTVYrUBf07Xfw24UgkKkcAb35bJB71oNTG+EdC1MgEtZrs0/xJvwv5mW1DZAI
pEvtLFjtegCqtfX1yb/Xeez4YY7F+UKmNvyENBLXpGv1DuE6NFEXm3lf09L/fmetlszk5I7HrwvN
MPRSN0DSsJlJgvkx3kM2pFmAUNSOIYQbY4KDmVj4Ej39qezdsQE2R1+cWp+oH7GSJKcyqD08Ur8B
y7qelWXBnmjwutq0KhJK/tllGI3tl2LDG/wGO58dq7Wpnb/LddtOydP8qcj+Jt3OPMPAPBnD34ug
psSQT6whozW6bua7GuuA+dOt34O9ztgvGiYWdof7qUWv5PvtOsX3UQnuPIXlUWsXoc7+K6ia7Kto
srOoCPiS/qP1BWF7EjtBeQs+TraCctePfbgW5javT/hRni+2J1yxIySNCDMLXhE31kd5EiYrLtGx
B3eOlMfyH+dektW0XaXBXyX97a5nLOalYHN24HRGBt0dZBxfwS0m/SL9Ynj4co7ZuLZ46AbZTINL
uE677hbjleKiVwNEVtjv8CGLZkkLp7Yg4Xwql26RqSRA+we6qNqOev8Zf+KdPsHcnbqlTvuTuioh
lxsB2Tf0eounQk2r8xN1OpP8TouEcRcaKoWQ0zJXlojnpYyctsFe200eA6oNyoQeQUb+F/yar5BB
8bndCuYCtN3opAXp1DUI6VZ4uGTXwvsDpkSx5XyMnJkQ2MsjqqbkEW+citSdmXvfCVbqkoUoCguU
qZX2+MwbwGQ1u7DC9SbJbR5MY7z/QGjsQ00Z92iK03mg5wwFkeEjcyM1zpS/6UJSRP1h95isOKkQ
aaawOzAyb52SSG7k3OUKS7I2yxOPu+UmfBpgKC8g3qjmkOzzArq/53UGv3pavdcrarNl6VFtDChT
eKi61Br0ktwSW6va/0nKuHWEuE2N/eVMOZNPxbchHlNikaXUvNBzMmuL5oQY5BZW9R3yuXer9CzE
PZ1xbqFiBZTgjuDVmqgJDeK6/ofZ3iWa4OZ3zV950R83HJegF92Jgh8WzXGWbONmPxUTzlkaUDcc
LZIF+C+RWgxx7wtIR0s3sAxhfuk4gIsljyOUVaVC6rKx2T8DjU801vrTUnyT4N3YZRJHGnuXL7wH
cQXMYTy1sMSDkHkct83qi2GHFWwaoOxtlNNAb8vFj0cIDWoxdE4asDjj3YYzJewgiaZ5U/5JV3i5
4DwUGf0TJAkMkhJOVlOoQPLCeseVC+lTRNjFu0y/HDI8PC4nOfGyDO31TL441SqtGlR9ywHPRPrR
0RJboHl1cSdDUJw+hHzY7Z85QWa49LAc43m/hnUjnCkExfCqs9l69TSt9Pwb7IT7l1AAMd3Pc7lW
leDLFUlWcZp7bNzPsX4IbI3CdLieQ45KFBi6NNsLqsa2HgY15jOV3d+wrqgef/bIZZQN48jZFN3n
PMFZZl5m6ZijOre7reR7mXegX8kmmpOGnBY+SYkXDfhfxWMsieTJDF5mrbm7QrsuCtVnMSgIyKrG
HDiB9iOuvmBwVJ6I9q+nX3Hg/DscqeQDyTWQvK9bb7jL1xa4b0147WX/9S5mtrNO24Y+yh6S1e2T
r8Kvmgpar5fs/iqv8GR23W0zzsXoB62Ol9B4v3yy2iyxV87d0Dyip3fqBfMG7VbFnPatPfP3K6KM
XSPJV0BK/7A1ZZgET/T8os3n7AUIXR9pfJzuBmtG9k5gIybjGfEisUWjGVPesVuLssYkFP45XSMP
0K9/1bv7qZcXYKWZ0Fe45+AL4hAnDWWax1b63xFwDwwAIy/oYAze+47bsosHJrFmXVMPFejXh6oj
ldnqrciFsiu3Mvx0zJBvWEonDJjLfGcAsusQfuIsdqxKFEmXJDZfRf7WMPN4i7ttz+uOO1IvXZjT
SjhvUasQhSjG70HrP0O7EVumH7k3leU5kRUxjp5ayRDK7rqMzsswBNXgyohVZ9FpvARyEYFtRC6K
yX8e1hO4fdLb97tx7Fg7hZe9nwB1Mn6g2SuJEur11pkVPlBlCOzM0INPmolHjxW5yAl98tJTZHdx
NUWD8waifJ5vEzEgyJ7Iw3C1tEDizyPPRgSCxlVULsRv3yO3fLgRuSGd99+S2+Maf4q0yaS+iBAs
d6edYSCqNwLFuvVuJqeDkDkv35e50XJVF21RPRS1hRwZ0BUkjIlCcYlLRUDlNwe/Cyp/kQQCNfpr
w6lh0yiI9M4DgRlRKocArgk38Qu6+nvwncAv3g/R9wlayUJ3dBL0z4BRzeCqCgNwQr/cOupQbaEQ
fCbnnYCWOXseuJ0HZhXSY/JQnTM0rwqKkL6FF27d+kYSj/8dP969RNZjJud2XG50oeV83Q6GpU40
27fc9GNPzJpnIpYnAf471I4mHTcao3Vn7fzzRrFw9GGf5n2JDfltj4OmzxHCh8hC89JQp5xLQFJw
y0/7ajUDVVKeSCaUcE0rPAkyesKn97DioHTIbQlrxTxoQul6Tm3rYB7qoPT5jiOT/ZrdLsmSdtDj
Ri4EZAxiygqYrBDTm1pgtXt2rpYCKGaousC6rzE9j31Wg3BnzdnxL9NFy80XxvcBgyzX7T6bCyHE
kQRo9kDQjWDSaXHQZJtM7cdxoEOXQ27fCcvNMIeCDRwwqnP6BjUbdIjhw8I+/cEOOZCFKxxTEVMr
HIGypfx0CzxG2dkTVaXa+lE45qbh0NyjRFZJbOGKiMT54+/XTN/2W1LKxu1C1QGoadoZ6dYBb1vf
lcTUivgTMkkcWUVPbU2abIc2NKphnrW0vljse3vAyDdx407kRlxcyiK3NMgBjgg1XaKTztOfTBJF
3li/oXCZknX7miNS3hYQ134jz3AzJ8Kms+Jj7JitdUWD/Fzgb8viBxvwU3SeChTEcLBG8apv8F3c
3hsSH9n2l/Lfyd3jA0kreuuOg3G2Mac0YvgOQx76otGZRxSnEidhwir4HzPkHzayHABlepwx99XN
vsNR+MKrVQewSbDmynw2gplWnXtUnkVfOjiy1fSDzGtXFdtn77q3ONaNvHV7rAHdmg6ksEslrF01
HhfGvM6jQdCrbvNjmdC+KE0yWje9Q0sgQ0sBHLnHANCVuOz0sU3xP0aVEKU5BLWB8tAB8QeZ4Hlu
P1CeBQGzc+ELdchKWooDDBkXw9I3sO3tnbqvms5BEmHeuehgbuEIdvQwepHjVw1vU4VVHEXAQUML
rwj4sg856S+7pHZRnIuZKRxyBBWzk2licW47aTtdpNoacYeIKOBmNb0cgf8P0S+OJmrteXEFS+cA
uQELHx3QcslMxz4WbkvemVubFfr6OIf2VGfoaXZlJZPKUKOfrk3r4vFfrpuEq5vBvpHV8csfVUlx
mAwk5XseJNYFE5mQEazo/lJ18GcIB/7HkMWgZBc4QSJsIvCVgRUzqQmIpQEoc/8Kb1Yy5ED+/Lg8
yrWR+FjcfaccMfOLdrM89tSOBf4O9nZKz2e+FVAJZjFTfuRtafzLFFjwMO42grAEX9yJGlOOWALu
WpsJDEpLZcY/UFBVb1ppC16HU3wqbLKrz1KGku1oxt0EiF9LXeqw90KPXXYrT0g4gaZ1Ts+tTiN1
+Xpa5jkABuG5K3wmuSQchQWzguXG8ertWzNUI6y4rr/9+abk0wk7oWy9LHJwfo8KFqV+JR4u1Vz2
6jJyM1uRJOXHCkw+TtRVFGDxBRSEYi/KJZyjJTWLI/8bQ2alTuRge36V9v5/USVqRN7cVM4wzFf1
S4uXH6+3co760cfsX87lGFDewAo/eWmBIfgMb3/Rw6R6xs2sE2SnKviRDuqHztUtlUMdr+OZF1zk
0owfarzF8j+BRAnMFJxspZTeeyPamHu2DNiyFah5+0/roPk+BF48XsFedmuxuZMpB6LS/eCcEmvg
woXVamlpD509l/5jetwbgcZZq1iIUMqG9QrjWed/u5pHuxje04DnU9Wy6nYon6T1BYMciQ+J8o3/
i1dGmxGpoCbOQLn5f0WxT7q7qvricbvNvxYCvcD+gcBOrEfdRTBwkPUisnYk+gXLzw5P9NUEu6a9
zRZPxr/c9QX1eUOyEaNq7ijpphiKuvtBh/c9JbhZsE38g8bv+H4SWaPKroue+EBfzOARtvasaxBh
NrU+uwEd4pR/XNPAco10dgSW//9T0SIAaDZTxkjxvuSO8SkhNkwJUkIeB2rX6ySWeXdSR+7bAF1s
2mDC0wwktMKL5yPnBxkFvNbeDE0FVaapSrdqZ/6kjylNeYTh+p6wFX6rYWne2naqMZEWJT6KVtX7
ISg9cRyIg5fg1hI2Cb1Rjxc2QBLipIkY8XemFLEHBx4b5mzgw34hlg1OVk5G/CwSm91qssdetQo/
fflZFHuyJbW57QWBG0aD0IiCnTzyHx8G/+Pdf8UYWTZj8gJ+cNftys8ZLbQwttARVhDcSTOJr4vf
t4lK67gzuPkcqmiDRZ4+OvnwA64amMr+K3vdvWwcSwSvCJCg5ROiwzDy6mFu34kMNBYEcQhPUo3G
sq2+4vgOEF/ygkHmxx0Amj+5cyXjl4bWD5Zl6RYKfcAs1uZZKzDTS5PI3uHpO7/Bekqxw1PyrxX7
ZuY1umFJOYAortLDFCIIPR45rx3xxOsIGiAsakgxHBftqPZ8SKo0BOnza4mdDAX7t+EbnktEqsnj
E73SMk+TaMMSDP+lWely5lwPmi4hzdCcQLyNdjYj1Gv/799TQ3xjoF2mDGHSd1hrOHVrtYGfzSN3
peJQXIJL6Iu/aD7CtSsPOwZUIQsIVe6Z20AR7k8voTMR2fDVUm/z/33rgx105GUqk5LmiiLbHrSM
JfYTZ8N4GqnDm+Mt8tIVFdM5jEHKbQgGxFAitI9NzM+pDvkDyJtkRySYxL4Is0UNjBzEgfWbUzmB
+K//5RKYnYCZadARCCFWBg4cDtc6sjbK/+UJhLvPn5nLYZiu+JZBpi9g3uwwxHzBS84yQVKIpf2Y
YJrdDxoJpAjFcfVt/9bnlD87ovCdW2VtBzgF6yk1oSHOuEqXLzGLjdvhhgn1VfBqAcGNv2iluVdi
Tn+DmRZ31oeFHrtAnm3YZ9RMXSKdjhiaoWx9tBN/BkQREghHryVhLB7LsY6ynJywzlg0sy3W7xMC
JbRdH+EId93azFTDxpeHX5Fn2S0JqZp3uJ95otKnxvPKZqyxV3g7xCgv6AS1vyQBYKAbf2Y8KLRQ
CfKMifhH4ulSW1k3JPUJU3ORlVXLQPyoI7qybz1vrwCuXgR4RZpv1bEeXrrWy0boWJRlT1JLqSZq
Mdp38rTWgBmhOOTzwKYipkVRGtDRtQITJtW7rFiXvciuQTU+77D/PUzsmBKf2s3l/D8OpSjH/BmL
aYq7+D2l07BHzPbQgSLmmwbyWxadQn1PUR+7BKG/pqC1Lv1m6+3t7wdP1VfTUGJVZVStagU2CKKK
Hg2bbMLHbdg3GxL3T2xuIG4TqcwHXDx3t6hH675+gwxTnOy6yK/zZd0fti/T1PLKVbjyw4d+YHZ3
XCyuHEXNSuilTWKhFHkON75U8Xh4h6pDw99pBAbvFgvcpC3/mmSOznw8oppUNb6acwDcLjUscOdL
E3r/fiWPzABOTeawJhcIPKDl3EJoNOK/LZtez7+NJH3+3LMnpsg5fvZDzMtDvI5ahF/F+s4SS3BS
hO38lN5j6RzmqgKCALml3Tcvqfwn/rgidiiQu/TwoF/Opt4AVDSaJxjB1cVUlECylmvrFfchu+43
pWDK+ZrqfAMsQ2OZTg+aDV2hBTOpIQ9EUJxgxo5DfIh1jwvKJVZQUtOs+2aTa362AqhEb1hYARu/
SAZz0Cky9HY2ErXs+n8y+z1kFCbbn60PrJk4u3drBi0eGmb2+NAxVX9QJ1eb/SdOwr4c0KhDdA8X
a3qPncHJ24bkbJYs+Ymm5T23WhcSrujntlo8ZchWig+VXta8yulE8ouvSZmIkVGbW84gnt4ADOHV
p2HBmxw1j6kmyZVjOnyMOA846mAM/tJx7LAcaJa67ePmVj4cOGrlxK2fC43kJrkqTj0r1RAh6AZ2
0sW+nMfWvbcw0qxc29j324PaY1DqzZsde9mQkhu4akJIh906c1Xyyy5C79Me8fmPKwwioycAK2pT
9eIehr6fkK51IfISVjrLoiryDDztTDbZrAwdyLKzDHHik4WZjg9tWuckKIp3x95b4bKrZpfZluUe
ujvyPzJvZkHO2s3aQsctVxUSVBOq4mgeXG5qTSw2YFp0l6qIeQxuVLqDf566PFNSmqQbiV/PvN1Y
nmozbFZj0qdNVM+ksrT0fBREITb8cBXCxIGUV2u/J0rBd5ADjq/4xQ4VqzdKAgUAI9xje9csG0cX
Wu8ktol3kp20n282yCvVFW6wbT21VpZA2wEevshM2BOmZfDtmwHIL+KBmFsZebLyAcRIbt5563/e
ty2okfxPIT6cSGvQdkqa4tUytVTlIMmi5S+19a7FvB+TrqQg3wEYjEs/eRlQSUzyOZxgXp93Lzt+
vh1KqlECgZbTOfjnbH+lJeuXcfmkeOiEwRl5NTU1EHBcFY7OtieUseMSo8Y3b3FY4viLuVADiXGS
Ou+XEaTXhphB9i9PjToY0zeTvvTBjHW2d9AF0k3mbCjDQFXA+nsq2YBMvNFVpIuBxGxhMsfDNf30
jYjy9/o+V91SuVyoKxYTgJ+ycCnH1hB+qspnwnP979EACzMWQOqirrJ0i18d2zaK/a9lmegPNpct
8z+ArsGCb2XCnhimqVcf0/VpG0q/vD1/yjZ9ATTPyi5qIWSxhCEYx4v1J64QZql7+dYZkDOPR3kc
A89a0ixB5sCNnFyhorTOF0+5betsUx2tfHk9J17Oc9Lg8HYrCB5dLxhE9RVD5g+GY3LSv86mR2/2
DAb15CRBMuAZA81lKT+jP5qqzAxeOW8efN1M9VqhZdkN2/Ml8lvCSqkMYpKt9HqCpdfcoajdyN/K
GSb8WyhlPw8Kh7bMjwHnn2SfOhlyXuMpxl0+HLAm4HlDkX3ZsJfD0ilzmcDAvBfSgH+uhtEptnIa
kWq857OAz3fhsHYu0N9ORHNBQ5ojs12bmc6PAhGXapc2MpDXsFDm0QvoF/bHyVmbgDiWKmWAUEWt
RcH4I+40YZvSXEUL6GdxfAnfCiJsU3UR/S91I7QWJwqO3MlvNaEYcTxSwR5508F9Bmjn1KXKSgqr
qX+Srkzn6Hq1Fnfb16k3c88H4C8SaNmeSjDgS+nL7VBryIeS0EtnIv3D9RGIJw9iLA9tKy2pzwev
+UIoH23ma8flqnR1NF28lt+BLZ2b8LhBZdAc2TYFnQjjph1lGI2l4TqzWSkYMM5ssUQ5mJGWmh2b
r/mPN1Vstgs+h71jG/GDjWShEJubHrd0/KK06d4d5pEYI7PBs2kfQuTA6d1q3Yyytgrs7ZdYLABy
GwQu8Lsg8jEtfAlkMhL8s1pUX7cmO1MdhhJGMUmhmjMThfjBQ3732kvbhn0gDlb29zyF/XO/QlZG
nFmpOku6JNOpae4gYblJjpUNYL4zs0xhP7wLhZonE+JwvAyxzcZYQmXgsFWoYJQtId40XoEFJ2dw
jGLwGr0qUsNU1l5C6cS+DuGvSLXtX6g/9n3u54iSxH9QKKvDYsyKgQUOIW+jUzcaSLABJWUW4v5h
bLlk3tEY8y6c0hS4N843f1R/SAbnI/cU+mVrNWasI9Dr/6p9SEAp2FqrbXwSZe1u5bkfxlTQG5Z8
cz3so6y7Ws9xJnTIdIls+C+7vblCC6bCu3sxVffqU8fCojPKb+EZZ8eO0rBH5bKzmW3LcuA9wJoO
538kSQC5ZDT1+VC8fPFMxv4sZs9/BT5N/jsYoVk0i7rO0pEfMnfoAqQg/sM4ZHnfyFiEignW484E
/RRHuj2P/5qTddrz5+IfrCduiXSckcDEdgELLThOgac/rHlC+X/gBujItcnqU+XrqbVHm6MvLMLn
Uii5W+7RnlEUr4eMGMPW+PV55RCrB8KuPrxSWKuhX3rM8xkEcrLo7CuPf9Gj37wnIpbeS7Ixp6Uj
jvLoZu9E5oTUTlnxwFsuy0qAIIsqaQkIIbwowiIBuXMCtE1SqgPkTaBJ1puo14GUbOcp8u/vme32
Wzzt6S79t9RrU55kZaPv6hfPBVHvvmTmb6yzDi5Xtbnk3OWGLlMBC0fPjvnFIjV6gRuOb3JLnSOf
V6PmZ4gclf+6M6vETPriCTCsNmEKKXZtI6P3GJDR3iO0BEEszbxJjCZegK07VoXgAikXJaZ8ugVT
Hw2xKOtoPypIa5XZJx47IoGynhWLBGoqJitCuciLC+O8LY+vLSMQ70yYd1McxmFFl8OVES934sh6
3nO4ydp9TwHBYaS+vTr0/vQY1eS9dGUPm1x+5GfBcWssPNetmLXf438fMkxUv0IFqFWad45iRONN
ee80UJw6qIdEh2S4M7PEdABcT6hFQW0hPb1xyDqHgI7MJtoM6Hu5aaqUSWwN+ycpqzUj4henrmLR
LOKeMk+BtYLIRGP9uMLIchpHI1ygzgSfspQUedmTRgP4kTiFToszRoDSdsjo+fXy4itiVNQJzswH
kPBFH0bH7qOFO0jciR4ZBj+FgOuJQbMigTWzax4z/nTgdz24tkJUbOwV8b5dZd5qdPnkdD9YLJp1
b0gf/7rJzQmw28teO7siVXaf7muN8VqBuey7jLNqlvOJtuCwYaWU77Z6t62ofw8MbBMNkuTzdRkG
MiwdFutPFOGSoQM7Q75KFf4uci0xbqMBQzwZ30YXKhN+B+oJx4Cgsb5Tsb9yfNvlqIXzMrscLrew
jHzn2dgnEBIKGMGj6+p4Tr/zscuViMGNXLCgWMb9DNmjB5qNgmXL/VEQAi+wE1lhSkNDilOspcWC
Nbhytzi3GqffRYZo+4REqguaLjbBJlS65phi68OP89FNAEnsaC2IMviF4uKCEakus6IO6rzfCdEC
Uuj+a1MFd7X0VOitn3jlJkSnMT2p7piSmM30jEe/fMSZVHRCcz0Jt0y58ovaxZWs4+MDErJ3Alyb
q9gkqrjss3m5Lb/qgv80kkeKLMQ/3HU8iOfcZDf2Fvj0/vjoueekM4qNF/5a4z7VINKRJ9j/UD7z
WxIfdF10OA/1RHpET/No44GYUCHM2MtYltOfLHabMnr5WkIRxvJ/z3WHUahhgyaolixIHsfE9HeV
QLV71FL8RX/62/T4z6+p0sAym65g5gd531yzYKZsbmz8fLexg3EUe26tbpCgq9bN86kiF45VPBo4
5HqLBe+1RWNsz3/hzvHpPT1vJpTDLzlQf1RPFLDFoT47fonyYiF5znRNN5qjXN3iikwfWxiDXmiU
OLfshBSj6ozlZuhtuK7Ico6OLZiho4gwHkM5L4xanQp5RyMHC5wXv0T9geazsQa7JEU5bRM5MxSb
hJGSHN4mCrn27/USbhiOKThOgeYF0oIkwrM0sA0gA/qnlSKCl8UzaeOw71vG3BTCa/OEhTGe6bbh
qjotIDgZBDYSEde62wjtTx/XZI90z6jXoSfn8e3wGUbm1tJRx8R3Ze2UfqvqlCTvunDzJf8T5z39
FXfeIfTXxL4rKEf7A/AYXsliQXYkk98V0uxxbcoS0O8RLq+RxOqy8eQkUXhpFeLX5XiZbFe7dPrl
ZcDMq7QxEJ6dEcO1kBa5FD2jYXdrE6VPGUKBDBz5zN0xTTrN7l7qp13clYpskZiKtsSSzdF3Gx8l
JYzdLbVGArOCqd7UZfOekLutWAg0WhCFQmEGBzNFDBKXqC3cRmimSCGfTfpawGKROqA9+m9SBq/6
s4ZR30egYYioWbXEnj7HbJd1D/9wlb3oGwhL/wYn1ie1fY3NgYUk0kTobM6jTDnNKg2hWQhTn4n0
JS6M6i3MYAxoe3zlNbHO8LeBwba+UV+sVy/tCBx2yjn+ZSD/JHPuocUKDS7pg4q2/1GlKvegniK6
Eh9WemNo1ytvEPS9tTCA1DxlrLzSUMtFKLc1+DkY5TVHR8u4osduk471YzUMSVApa7AOBj7eCbOk
B0XfZyPHgHvlubfJh0F8or1vjl9RL7mNSDVCmn3UL6UUVn7SAq0jedjkOjxNCMdIm/2ovHvHPFeO
9Qkr3Aau89BXWjSp9aMoGavMfNrIVRW3qU7E5qRMeystUuBGdGQPZ4wQvxvMv/Qwfspu8mxxTNYl
S+18Tk9PaCercA6mV+LMa4A9xNt+cNb9sJqnRUSl12XRE1zJIWoaOYTblLV0NmdIQp0nGqXetEko
Z82HtqoShW1N+nOiZ3hJopEsLXkxLAL5/MOkHuy0v/SwAK1q3Ztmv7LmvM5EVkNL/XzkJnK0ZMsv
QrTvHgYcJ1zBKbajDX0bTROgQiwQY4uuDWm9gx4jcK+ReDEyAct7YH4AmZ4qBxIXV0xW0ocHCUnv
qdIg7tOVUb2sWcEZFmOtWak0I4ex+U7K7hRI5/uUUD5vnZ2rm4ltKbasJqiOjRqgz6tqs7sBNERt
pPRMW+gBFYiA6xGve2vygTGODbe7I7sC2sD932fp6PObJPE5yMVcmLQZmMv0IEAYrFTpO0dyy+go
PpHxaesiCeSbtTYGtnoeNF22SN2IPrVc9mJUR8Ai3jZTwavpBYgEh43OUqiKQO8VfNRmkFV2mMq8
LHabQM1kfu3avUBsvwUep8oJ9TwzLCj0p8apzafZO1dZNUFv/iUceUDGabRsn/FFUWeRLhqWOyel
16PiTL60u6KQ0LMHOaz/T84Vy8I3Hp31t8Po4EGn5WdW/cPar9MjY6fBPsU7L/LFi/XwYyj+vYFK
hM2elhdmfYgjUbikSuTTvF2axVA4lPITDzt9POBcG4hjjLiOPGMp1bE4K4wHJ9R9iDUs8EleVsIP
Q9h0CcJ/qhsIu+RwdpmcZgGwKvfisZ/HI4VjTIpW1wgqe+jr09zBbv2z3sO/NFO52DgebIzz5Mee
9DrtaklPnlxKOHh7wXW0d1NOQuq6q6E/Qg8CyUaSh9PlpRoUvp3tjes87krszA3KVdBgdji4Lh+8
qSsp9Y7APKiOYqEhYM1RdpNo2xIWmjvgoGz5AQ6McHrd/PcTujV4NLYTuppc1bJJNt2Y3ktdusBn
He/s3+ZGLrTnHlWP8sMWSZNLujjbVT4QKLWuTFPeZmdkz8jYvhFP0TZkM2O1i+dpwZZeWNeF9KWs
oZzcSUFCRvuWal8Ye8x+2TNMWwd6Q3urXvnOYWTMbe82IpzjQYOAMsh+3KIYNEvk1AqIj0ghBTE1
69OjDwzeeL2PI18N03UaLOZ1zkl0FF7EXaL5Rn4uwwnZZ6+lKuA/9LivJt4lHumHaA4vcQ+tX746
WpfeVSOSG4erz+cuSSia1gABhvcuODZlruB321BmJ2F18gBEgt2Ekr1d68YGoE1CFDGvg7cZQv7o
pC9F0NdoTL2ckemyOeKlR6pbleDvm7AyaVgBdB2DxLi1N6YiemuIbFdLCqQB9QKnk6uquH8hoq2F
EIC2w542VoBOBVWpjHwo9XbpzfnotysJ26YktTmTUyPuMGaGAlhw5/lmJjh1ikzOl0KCD/Az4lnI
sDvocX8U3uHYjfP+I4kLnDWO8n/B2C1R2q8cKXBqR20hfwTu3lfb65yHDCuC4dhTA/V0NUVZpsTT
plOBD79P1IHbaTUpe/6h9x5Q8KAGLm1xDlsKx8c42/Max/otRCUQu1I7vyolNmiBair3ofZLEZt7
CYGbk7sPVipdutYOvcrOlwQ19w++bCe+f8cTWoAUPF7KhiXnTf87jA+8HGa6folxRN7SF3zTBE7r
6lqNQPu7IgPWMds97uemGq4/TliKYAteHrevVOLNbZP7ii4BkT02BhHAqvRKPCYdJHn8UkX1UMzY
BYdw2bi7P4xE48UDQo1bHm2lazgk38uLL6mWiX/tgQBvZmZHXY7SYkbK27rw4w2StLwXy6RTLMBa
xKsHU2RksyF8bCWFqOAmDNFDIPa1rtj7SwBsDizSPM3ucYiVCad1/KY5R1Eu1SaswdGyxisGQHx9
wOj43PBpGcHl39lYQl2jeTWcWf+dlWBzMnDmkQpX8XadKHlR3i+lByCwcGBSsp0Tt6ybYYNxb0QP
S01jtS/zE7Jw3QzXiFzw1VrzLOgdT1cPAGuj1Q9gIIb3Gem76yvX6dNnqfXCxhpYN+pQ3NBSLPNB
leZZ+0qCRY1ZY1ZHQ2wcrQx4xXxvnsuBooVgylsLGQ9bYD0dpVZasAaCEo5BoAxHinEhrSRX5OcU
UP4YzMnVync02lvXF3Pju8uNVuxYIP+a93Gh7AGh7pEHQzkrxipQzB/LnOVh5kvISm9upItxLdEJ
W57AQDfVXdLHS8GxkkWH2upZN8ZIAypCJJwpl9FNfuZOFYM9B/PvcfxjY4JqBxfHUAoAdSP4yEb8
DRIGE40wTsxF1c8s5wLXpP55/c/bm368jOUU3q6ipF7WDnyuVkhjQVZeDzx9txjsuqAfXjgJwoZ8
/21x/37FdkD3YoTuXLyoTs0j0GoeXKlCCHGQxthE3rHvNV9xAIlwNlAf4gEG5V77kDDsS+m10rTt
uyl0aItYNZB3KLSYcfWwQLgVgVYK18xGhwe9RsZ8qCoISIo2k4KXy//HrLVHabHPYkJgF5G9xfx2
Nk4bpnQf2DR7AMWDiefeVT5voazgPxQq548nGIY7zgsJO0p1coW2GbX7S3kuPxJKU9qXMBvhNDoA
7I90KW/W2ef/lAeu91e6WjniFNOZUKJbgzqcy2HzTByPc+jwxrmMOmVtOri8ilJWDuIcI+OZHLeN
QAaltOXHzt75AFjZFzWBLH4LjYdSOT/C+V+m/OJY9ypzwod8KVt+FkCLR2HIQZnvHK2L4eKxv6TL
p727XIQiKxTkngtyCMTXrQNSLH23+Q03FOlj8UIVQZhNkLbqaSiKRCryhYAifVLaxvAsFHfhqGsl
LnpYvdneUSSz80epmFUTfE5U//HU/H+GMyRPFOkeXsVweHCL3/ZPJMjUClBt8pqh3y1i0mbxbYmB
JbO5LvqBJ3XTFi/nloWnVFfJ59XOYO7vFv8G6yyCuHChjeLVn3LBRwjFlRuWbZOle1nckmfpS6bz
19tBf/ZZWdIHdlfqOVwkUwNxfa26zgCUQ3wo52mZhlymM3nvSSn8OxFzuFbK/dlVgmBYj7/b087s
Yk3DgjrrALQdpkqswLLb2muomX4OrLmr36KJQCnyTmop0crUX+LzMZaS4PAa1kBYNEIx9YUTOi1Q
iy7Wz4HeGRx8jZLSMey1tmDVoncW7DHPLAk7QabxG52Jmx5tCdwmu48K/b7H08NAntGWCSLCeiiy
h1VrxqYzD9oOA9RzN3T2+oM1FUIrz7eSjODZksyPAa+lyieghJfN/t/1tZ906jvDaCtNBYWbqQSj
qoZCO22GC9mWuo3WJHyCErS5/0W/xgkVFW+phzQc+nDGJiwF0Hx5x/Lw9cyvcvMfcj6gjp0OTtqb
ZpoGA9AoJx3jQT7asvwdCBt104DVzlItwTx/L5sr67GEIp1Ux8DGTNYbu63kRzIQ/npIENCBgF/X
OFiU/RM9GAhoxQyF9ayrRa+yDH2Y406hAlCxUHmKfcAmrBtrwqHi3Oyy0iyNTrdYPW4glOTdjYTX
VqU707kd7/3rVgbtRlhwvxxsvgSvpwKibLW6AxGHpb+LeYXOpKorGtlMnSBjCQ9xe1WumpFbdP2m
QGQmgsDcIAbyPTSdlzkqzldway6/piQcFfNqd5djcxSdW6pshAFSD8qLlqD80DfsmHzct3OsEtxR
urrBYaTAUbEWKV3GumN7sVRukD7rv0jhrBMbyOPo/Vk1hsj2fh7Mg6hMeUobhua8TFrDpYIOWI6q
z1nE5I2PzB2IJXiyqm9A1NrpE4ruj/7AvBjd3prEbk/vfF11FWQmU/q2IosWqKr17/l1YhH1tz6E
wgY8MzTYWDaOH1VVGoij2PPn58AIijBSaxkOjgDnSX24/eLYHPemZ4zumddBVsUhtR9n7g0tErw9
Bvw3KA2zRvLmZZ7nmw72JKGCljX+yoAraRWoa6gikABRWUO9Nh9eOhJZsU39ncGnwTpco/8gAlPL
B1xMlugsXrn+hOiF6UYNhD7q+aokWFo0Q6lLafxo6mo8SrByPvLL0tapR5Q9aycTd7Us63WmKT5w
qBNYZNZkWVZBVMYfJp3q7seBUPUuvCULJcCNsZR6/OA/DhB5QlefGEA5SU82FNyh0RMNxxKY7YgJ
U2Eyb9EsPcevBe12HV0bF/WUUVTIDPTv2Xi1IRqra7/Ax9Wfguib0P936N7/5CUWzVsPG7M5DBn9
SOCrdDZeiXjBSuBSZi+No5QFyk9k3qEevTxM9KXWdbuO/g18Qvg0oXC47b6DJRDQQRu+0LKUO+XA
Hde2tDfGz5yEkTdurOxwr7aGMqeT70knl9lN8II72vpYKbVoqExWQgR4OM4xGdyNn03T3kijVgDK
a3wiAAQN+8WHo1WsFN8RGPJoqS4s3RMEvGB/AdxuwkQ0pl6MocQeaJgnm+XT8b4XUYo1pMPyGxt3
fMiqlZOP/hDe4ii2V6E0V6Rrgp65Kdyd6J4zukqLHfGl3Y3YXlhGKX4eriIc6eMTa2d2fX8zIDJE
oVBXKeMLz8E8MKfaAliePahf8LjP0xkBsVq9dmAbpDYCA2nWdB6Qg+1Wf5yesRJjVSdk1zc7JBGM
MQpEz4z9aAnuhvyoGu6tHZaQbgGK9vnsNTHzTO2KLCOvThSL84rDhosQeQghYBFR+op/lzBJAJSI
SpPtsw4D6RNCEW79GpIJ4QwNn48SN4HjCE6yIAyv8/tSwen60aPTtMRhdvSZ1QI6N2tony22MH09
DseYBnBJ6NBf0H5rOAtLkkskDYE2jAG686F+PwSv/aXWlpZ8lXYV/DRW17Bs7YpiuwMCcyu3yjLm
HwwFpDtgSVuLqciGycpUTKVJDCTzqe8nfFIQnF/0drI8A9q6lrXWkw2jt517ugWw4MdzM3wNIki+
UZYTklDOYGkrn/LbxqPw8M+fX3WBPZtGN2GpiM4T7Dtvn+3j2xIrDQHAaxmufw8MxudxdrZRQwu1
nc2zcxyDsEy/aDvx/swbi8OmKn8DIafNP8rsCBSxJO1fv8bT1S0CL0lVJ/rmlgj50AEfd2B33796
o3gFkfgHcJ7cn8uHklatWQqtZaDFlwsmFGp5kvT2bNOg80tJofpcR0/NZ9dGmbaI0/JyJyH56qUe
HPi3dLEWvpCkJJKI+BAJVOpde+BAgqYV/epBmrlns8c4m60mTV47vi9NBbTUkgzmOy48/+DnZO43
dCEJSTDr2LOHr8JddymfN6JtjFiTc7ECkkAi6/QvCC/g9sCBaohJLAQYTCe57tpCe5+I6bsnMvCg
jbpdQsSUJ+eq5uZO7kQtk9NBaUqFkm2qHB+NDfkfUxFY+MrHkDV2Xn1jcBd3+aHR+dC/8RRpULfC
9UtUAIkRBSLBJAcRqGVrEgoj5a4eAJ8OGm/7L+lXRlfXkB19HpANeXb1GVjUyW9dPARt58nqROj9
+2i8Kbt0Z6AagiA++p0D1r9CX4xD339gGNFKRXk7oItCn3FeiWW/cJAIAkMn5yg6JkF/aSfVUsZl
2w795rI0+0OIygmLLihFtyVC6Hw/CnSxuzpkKTSSIlIfrm7/y53OToknDcOzG0X3jVyr+2WMGsQD
tQ0ya7QX4H+J0stbxvLjNaZWrqntmAct873vRTd1nDT39WioKnPVhSQSjnAs4o81sBjE8iBv+V3r
p+Mgp0bAIHZyq/Kz93UE4VSh5zV/SWGtJa/8jACAFN5UMGxogljwNjd3O7nFUPGwsJHP/VblLpHP
mXo5/dlalo5IEO9+gl2XKuHWHYnm7dkNqlWP1WPSiHJPFGjiHj35c+8gLr7y2G0cl+bZBwzVdWWD
ymsnieM8uTNnwvzSU35R56dwVreB+pYMB8ZlUsMgHSS0+yXRVCvuFZYTAh3Iu6aITj8KGKaGLjJg
4KPY1/l0LS+KM/fDcJ9S/GHNa4UcB3hYi5h7C0zIresvCaamx+Ee5hAAgLO5OnsOimvwKxQkBM7b
47FuSfBqWm2RwQ7ed+fO/JvjUDIqRY7xt9mAaUDQx0wPx8PRJ+0RjNFnOUztvF9rMfGKzweP92Uw
/hZAYaYNw7zDX+PZJSgqMWRvN+qI5Fa5/FSGcztbwxilBrzSaumywYjsCYxPPendTaKZd19zy3Wx
TMjv52A9egqHzHyZThld/foGttIlYffcY8wJ9HIDw058YbaHP2dbqaTvcy4phARNOZnAy3iPtmIe
SASvOOLyMgmEu2Tdq2/PGFyFVw2+Uzm2uZo3zRRqQMA9j/vhlzXOCBVT04P9v/+8JDpDphJl1asO
m6Ce4P3iA3mbAbLvheT89A2YAEMWB8H5+WlNih1JqIB1KMhfnsXNBHl4yrSqJE0Z1fFpCEnfXeyP
DBVIou/Y5QSLu2UyI8SHWi3Hi3hVLqM56cTj3+xKUdzl4gN9rg8ffcA9qb/FFawhrTDj759QuX/l
SdiEgehSTqcNnuiW5fEcSBkki79Wwjv4ibQzVfDbTXvLW7AUMZPDoBd5xn4wJyCFw6APuBKNiDIe
8RpezrT6dtcMEYAp3Y8P/n27k5pIS+iV8qW/uGLrHXVkaSQv6XKhNmrCVTOLFCwmb7RKn8eMl5AH
z0P5OiNiz5eYg6LBJySFLuAwQ63vQaKJnb8CGozgoKEBrNUG9f01O1Q6fWNweZTjSeqEVqNds/+m
Kz8ig2wBiS4y4WkxB96sPXEpgcjDH5nUHMUZCrqJt7BgfqWCRY7K3w4NEDg8EnWowbGYox+Q5W+p
ql9WuPtnVLCDq4RKhnE8puC4WwaXxmq7sSGIlUIo+HaT8NUv1WB6z6OfCLF7quf8R4oSXtl9atqq
QjoOoSxOzJNCY3kAfsojt1sKnpPcfiLDT8XSJC1+swMVaxbau5p6c/UruHCuXY1sWhlThN9rzG5T
UzynakN8i6AwD54bAr4y4z1PsmOP+theywhU8cZdMGYpTfXCPHO1zRfAbmd6SBWkbCgTjtXm1qwo
phJy8j8k63ODxGFJLSxN+f1IXoyQmpOf17vp7+1+sJlUW6Xf6LhHF4vchN2OAKuPaTxFTTcAZ4H8
dNAlq8ApSFH1hHpt9vcvmH/ZGiH+RqaWLeTHhTr/Xi3YpOtQVfxmx0i8SBkWnmI6C0iK6IUMOquL
jCYOlXmZnCxW+627Y32eMo7VSDnq2/swcWWIr1uha3IiYh3bzWSWtYj1cnAPYs4mRHDifxFA/pMK
B+z1q4mZ1lY9gmxQ0TgsoARLKpTmyp3VClc3RS0D/AF6miIK5XapT2H+HadAVGx9iOT7oT4s33+C
bc6H8G9Pih53NOQwgUKVs71Xaly/p8Z2fUNV9e+SV7PbdGY55d7XvvbnfnIOK6LlxJkkQJAdTPvp
+QSOy0AmcV0EUAom8SxhLWKZ0/8hPz0cBmMm7+Hxbx5qatbq26pqDYI4zAgAXcXJDLCJW82MEuTj
kaWXXVaWwjgO1kd2TEJyLGTcHDQtA1w5YGeTSBOi9Kxu5B92KZIyhlo9rK0YVXhJk7dtacTwHluM
J6bkaY6+Tp9Cxp11E7hWA4wDVmWBnhdqxqYSh8iocj7vSO7feHUmEU0NEM7dNi69qi3CeSHQVxSs
YTYIYs1XLCHrVf6JPQ5nHQIGtXBAVS+slQftuV7YsiEcYhl+vHoG7ikBLKYmUo9fwhtC9DFfbyiZ
+4o7EFvIVGHKUOtuU271E82vd87Gl1Lp7yAnxafzWYuAGTF2d45nnlGvZmiR50b7+3zpOsQbCTlp
9yUoLL6rzoZWX4XMiq4L+s0+ajlBMGptNKnPY7pmiwFKijqbR0AFjtc4RZgdiQYSe2DdLXyeCmIZ
Kv63Vqtaq4PUp5zF02DNFRLTz5N6w1TjNPjF+oFq5Oi4XOerwI7Maa4E7/N9pc7mkfffmuoC1oM6
WegweXdKEGHVTC3XFho2XNJVkcbpYYk1CIa4n4Zgl00RPGG8NyM72HcFIF+erUO7fm8RpqQURy8k
JkFcxVMwBQ55ZZNSigaBOvZw7sv4IyTKct1P3v+RYcUHbbMGaaXqkq/Nof9Px6CgbevDn/sf3i58
d7QgyQ9R/GU05Zc73Q6ULGC3hvPv8eS5w10PpIuuie64QHurM72WvJH0YB45iJn6ZeyFZMuHyGqI
oMjCLaCBGZSIYe2BT2DxvGySUlJs7oQuzYEJVbI95oN0bs7dnVTQlpVmwIm4Bq9K+e2ilzrraod8
jwRXVfI8G9DR9iloUMQ9+RpjB1I7rN2Pl+c8ViyF7mQwz/++r/si07PI8sCl4qc3QxNhBnBtm593
t9FZgAkdeigrP9WnIONIxOqgalS/xOiGkkuA+g+BtKb1FNR1DWhLufiWvHAMWenxHfhYIqHxn3WV
cE7x0gRla3ISOw2RlY7Pns3jmS0U0OW3gIPBmxvubVaNrTK9dTRwEIRy0Sv6qfjovqgSCcPo4axL
j0q2qkOh3SY3ZbTGZAablf+HgdQ0mh1bQR6vjSNsYy4/suQYxpsCS+KwzSTGeHKOQV/IK1e/NFQA
SeeKi6/A7nIqZNyhSXvH+tS0Lpn/bjRk3EaO/mX3DhU1yfW4k77VwCwnnB8M8uvvHep+keA+60zE
axPtuxAJyuxJj8JDmajJ8oaZUa3XTA+7dsPwD3V8ks5ElsUzJvQpo8DzfZ8rTlouzyIoliceFMJG
zcBQ7AYIsrSmqv7rInILSI8UF3xSaD9mO6Q8p4Mbioo+MN1icc7QXuh+Wv2CubmuUva7dxDv04sP
EFJnfGqBso1iQ1LnULvKrwf3wIDXxgvYtB/eQYol+nB8an07fN0m7P18mUf7wn5vc/yya9Fi0oj4
OHDQZo3Eje3ADQGK+hKCplHS5I4GU/OsxrD3p77H7yKWPLY9N80hJzwSH/wCxF4uHPiZE8nvE24y
pI2W/ZNogWojgT7PQcUji+9wXjc8msLFFwpBq+VVTRvuUoKZ1CXc1MCvo9+Xc0NYMvw/svfB/dGN
7EOV9WWp/fs9bqPaitzHmakKKXOGx9+XcyGNzS5/cmBb9l7CdiN96nYWkgVH1j9s13+saAVsRuuu
1ilnYV+BqXGDo4EY05SBAZgKhdDENnOeTdiOSJL4Xqk+4Hq2gUR6Gu03zH3vUDQtU5iF64oLPCwY
OH2dSFVTF3oN2hoYD+dTQ67fns7wlvVBAd2iWWMcLreBOwsi4JIlNNdqrPn0FcnArDsHWQwyEbu0
3fsHPbhAr526G+Mc/TWGEFiDs00vrFq1JqJTqHlN1GjVqI5N9JEJiALavAoFNxU/Daf9SX7v9RSr
flpDBqe80LHyeomZrUPB1/gLRnUXpaz7NNS9ydbOWxMvsG9XLPq+d+bjkigMBXochqAFj8tJu1eG
/1tVJ+ZQnb55aEJEg8+Fe1shzB0graDO+dd2RVU0cB9EBw58PNLeQH+4mWXa51378n9z4wLX/OBx
RaYDrPkJ97jjdJi6EaemsBa1kfDoFZyi9Hr/i34OY8mPURm2Y9HRvumo0f/PwAXgsy2WZwwi/3DX
b+3lEMsMb954nOEEjPMGmcTTHXq8On+3RltMAQ33ISfnObuA4qprRilPbAOVFargptWe23UK4QPo
R0ffOCFF6+o6ab9KjQiCPGkbsdKBmJyi8A2+n/bFy36ZPuEte5uBVznFVLsJa/IY13FDGZqM3Kvk
8zspC+M7XcGCYmxtkVzAgQ3g89HCHDnc4PGhtIcUN2v/vlPg3REYQFy/TKhtrP5caL+bEFkO6F6V
id3qjdrAvEVoQYqgIcvdcTDY9IAZRKU5GMCEsOTdBPnYwlJtw5ZuVCl4JHfNBn36muSsONAogn99
5WTMxDLgLtrKXuW62EJRRAbfNc1LQWNh4gYfl2h6lzl2g7p5VZ+eL6Lh76cI8cpanBUKeBT6YPLa
Y9+vdaJyFnNQvncJjIAj3Q6F1aJOnmuf01Dd7qonTNBfdadvYe2ja5gM715decqFVXzoOTxDa2JN
fg4P/LZac+6pEpaKOGzGSlOQhhYH3FsLGViCaOgPLHBtsY0fpRKRAmX2wExJvpOpLMMrgTnmPJef
I50swx88KzaQ/Brbyb8Nfg+MBEfdaMLbY2vjCL5jZsUw/DQbj1dqeidkQDdsnyIsBIqtyUscUWfi
eOYgjj5tXTkafzgM4UXmL9un99EAjURvB5w8SvlRlYoATIBpgRl2cdWpjDa6mgM2GS61eu1HFUDZ
3mdJ0VbYk3cFCAE8SZuP3QHc72hPPd7+pgZwVbeI/lw0FlbVyD3vT3j2z8E/4tlLCVLlS70Mi+sP
GtGKErWsZ74pjjLQIJWrbZuHo8ASpxNyht0H7cqDclVnZaLRn10COBeFmEppN/lNWw5B5RY8549b
xK1Ar9/GeH7bMCtoK6PneR22ec8AGFiqEPk2KvGbL+328jigHqdKKqPeFCjzLo/v61bwr3nddVxj
7tK8dI+4QM59JF6idICfdyH+GpFKx4j3v5byBajItyljNfUlKN1hPHxLjTTnW+HQw8T8yK/H81jB
HKQbNbk3X2/YNCQnKxEMt7Rf8CsefRZAjs3YNZh4t00x2C+c1KcGhNIHlKpuVqI74IhDUA+nOXY8
7u2PMEZACK0RCFOIXiM28/9e2bVt7b/Ur1L7RBmnb2Zxz/2DEs0E6PGP6R5/BwZzjkqK+Da70rNL
XUy/G9tgvaAaU1L2SYX5/LXuwHs+aYZ+z1pY9W8uP9giK4XRDUrzXDMuFOFnqjQ2mCmCGH/eMlgO
ULlXuAZkcZ4FPQEezsJN8GLRK46K+o5qzsM/V2XG2Rvt2OlrGa5SmErHKNWAhCyTY25cTrkHwzkT
fLiSslWIV/M1tmB1Kbr7zH7W6nt8A0nD/MHx9f+MryQVJLj4CKCJlb2av1cZ39hBq0+miStCVOTd
bKPqSW2YsArAy4aAjohJD6Ke/gYAApKuJ+ALAi662ffJ9FPRuN6QVV0bAds1Ff0AxUHokrD0gSpo
VGO5FtKtZi0Lyp+oSUSEIRRYrB/btlrvdFLod4S4ptubW7/Z9g/PwtjYsQV7hCjTaLBUl2KO5orR
vOvVwd22EEQdNB81h116SLCYB714CCpXGp32wXPqNUQ+c2mJxniw6HHuzQS/2KmMhI1SYjc7CyvO
vthYaKsLOJOmdt3PqJRkGoUNPGNa6OouJMEgj90mJgidb9C1EbDJ6N1gWub7iqSzbI1LSvPacSjc
owtm28WSY4Jd5LqGkSfAT5r6DOdvSH8GawdAedy+7EQR8+WX8lEtt5oc+KNMyYFuswPniUWnUQlX
zCXRgVHZmB0rNTnNIJsvQBf/nvkc+5K1kJW65h2rkNi34LxZdfNqSiCQ+fB04C9gJa+kPC5zBjxR
+KsO5okjka67yGjgNIWG+b2DvsYWYuO8R4hJcGWoDjWZ512ZleFYFRnpha/Jo8/USTe0Sp6YvNut
JtU/PFf8L3YmFcPRa7QEGjXEqjAbbFfDicJ3EutvtHbUO7gqrvt2ci3Dv893GGA3n5PwDtcVgJrM
XVNzrIDKHJfYHgm3pw5i1gjBScVQSkhdOTnTaaA79cXs1zuIqaObSfMTMLVg1iDrfFtLdVtFKWY5
rZzMGH/aDH2G6NXgN9BLq1Rz0MwBnKVOTzT77gE371kVIsd83tHcIDD7AIwioWVHOru687OE7wOm
NPeo/gNLQ99kjjuhnAh7quQHSh8naJkB+/Q7vYoWO9gRIhm6NiBhkX6LREhHcPb7ow0BAnWv0z1z
00lCyhUHoql8UrwRtOf+VmlSY+xv0yHw7rERnoF3jwA+8TUi/Wk8xmJIh7QLmar7TpqONSzaoIRh
Cfa6H+Bf73pNV8TcACfdv+UHMEMRXzdzaM/xohVZ4dsF5oX3BOrA1GmxlZdffLymVa7Ldu09ezco
sRY88HDF6QpQHHrsOykEhrreAAJl6Z0OAWLvgs+LUh8tyoApsz0n25JZ8Ulp1wsnasutB1fOcnSm
ySEe+SoGse2rmLlWIDHpoPyxNHuwLfVZQQHztkVTEZ+Oen763PWP63UOIVxjbYGqBFAgH/MCpkPG
uBaoUVd5vmUae1OO1p6lKAoLXgQh4XA/kcfopUGb+JG0ehcgEKPUcZABkaFBiXdmp645m9gVGhvQ
0nqHmSRggFoIppUdxqwdqZaKeVsvm7wwDwZ/5zrh5awaigCqQtmvX9RsnuW7ssfTOoZ3E7ynkxwQ
/HiOajaaudJevrx4Wd5oZwTPowkA50Vkajrs3EqCNyNMZDrTQrDyZ0idzUXsdK/D+FEUj6xkDT7q
h4EjHSM86MU7fa0+90sedWNbblkTG2pO6Lp4IJNO9wtVJsEHHDohnD3maEAvEUIBpV9X1C/7JOzV
7z8ph6pe6V334YT0urzLqHlsxmfbsc6SvD6Nx317R8LGJn/0pqzI1OZLt0rU6rDAhRKSKHyWBLRF
7ZXacvV3C6f1DpCZEez6qZ6/U+qQ98TkzYwr+ZZKklIUAkAvl35i0P8ENJ+9PIB06Roe+qUbHJ3E
kMKdBodY8CdSajTbswuyGb0KR8q6u7cpBS7ZUXgYzs+x9VwS4cya2gaGgQJuIOLHaqVfhyqtDU+u
/KxHzYbWepY4MZRs91wyWblohNBkv+7YQal9BFthOiIE8a0FyBnzF0EOx+z8nPjLCQoMKtI+cZqj
gtl4IV9rEXUWV5kSMAjKySn7FYwWUpzWWJzgPTj7qHG4IbMz0f/xj80Ly4y7zjbzeobXjO9K4h1L
CTO13gU1Oj18ejieoDibBDevt2CkKnziaGPaPJBV4n2yQWYSlfrFLo2Xr2JMWJz/jQE/QQOFK+V/
6k1fsRyhh7UQ48ucgp2cidwh9+2AgjDQsK7kDHdi/wRv7hqtc+f+YVbVzAN13C0YSCZurnmGyuA4
BTqWAqrJ36RpNHqRY0kKw7dHAloYIEChyrqVUHXEgtSLqA/HmCs5zqaqtXO6nhXG9sXO9DsBf90v
sLUekwOrzdAIqlyzys7mS0gO2Z/juK5CUnyKCUH4x5JYZ+EpIzsRUieay1t+XMZjRpmJQTx6ypxu
KEIV4EDCjqebA2WPuM0OEilDfA6dAbbuTe+nUacR/yt39heN+KXV3kFtj7AWUnOhaGVzFXGex8Oq
M5Nsec23IrPQbcJ3XJ1GE/bvQlNWDjYlskiEcCpfvXiUutIwZY0fL/MfW/5J2mmPO81IcecfVpgO
lLOaN/lkMnUhaC0aCUendZOwLRpnKWVJ5ICMITzEFfFnsKM0DRYmhwUJ9am5b+clcF0x+mV2eNdc
/EDLnWIVDf32CNJOxaxOHV+r1xJtu/4hqp0LH0uydwRlbnWZSnu78CEqc/mjSAgj8mKu+iY8ssOs
guM9RDdtcGu4O5Vokk+Uwlpg3mTMMtSU7maQm+dZFMsV0+FQu+LJ6AfkqpCB7ZUR0ghp4iUL41MB
iNZ243BlmKXmrY7leVHp29YraZyEOTHk64sB7XKFkNz2aP9EF9gN+JbSEbZbprQ5RtybxZ8JirFz
Yhphebg1vea46Qkue+4G4e/2afoLUcvUVBbwBuRkdYrovnzNoLUyFbpIYli7djD68p2Ju8nAJkSq
plPZV6qEbIkDUJzr9GPCLPkkigGoEjkR6Lm+aamKI1s8a19AWwZim3gsNQb6nkRtW3Uzvm2nPYxK
juKI033yp9oMnFYN/3WtFC+CDsTO7mDOweg5hdA101XypVfrDhwfOPM3dYPabcuu2pydhiaCBMB8
yd6GpuGL1PI+VqeQyii8PnEHwW93Kvfz4dCGr++Ucd0ZI78NgUXpEPACIiDuHcEQVwB1JQUJoIq6
QA2IOfaCWbNeTeQ1e18H8o6OyOogxCJECzZB6X9O/oQ28cYMRF0TktKzz++lgMlkf2TXDNNKBt8N
Mx3OkEHWA5Zva3Mtcck2jkySyB8DbpLfTRVCBd6EFQUDCPwjM9oppeUb9vAp2Gczc3PCoyLlT+lZ
/4v4IVOzqAnchwNkz9crH95G6+g6PtvE9xSBMKSwzp/P1Xf3r5jpG5ylzhoM3IZ7BxzHxS1fGFTS
76/8fDlml0CMs8rHyetN1LWRBu3pmXR1PHQSoW+e/M9ZUR7wXx/LuzBCYsqVxCy+gvEgwXlVguVw
BxO7TeGnY2wtswk32rYLfZ/6/b3oYKl0bQdIMADBdwGSMksDENCPlPcT8clUJIG0jfPeF9U64Ut9
eatOdebQJIume6gUa+eoJVnza3hvlFrkg9GeVkhKDlwbeyLwb7/lBI7vbrWFaRda1sFdF08IVBig
n5b5oZCHhhIfwI6GmWm1Q81icF/ccqkyfYMiQcumXYpTA8OhnM4Ksba59ECmtISjSdqNmIkwtIoV
btwnMSeaY7/ml+PE7movV7LSN25Xobw3/1M5/CcVQjn5/QOo8pMdQ7ZFWfQQvDn5ejoqHafSXEgH
V5jTQtYXSVQ/gyJQnjA1uuIO+M/Mkgtmuj0+pIlCLEWo0x3VJCELcb9N1Oj19mOtQ0scJXaW18ag
JPbUM/7Obt57g0CJbqxzBMqPiKgk0iNhMoCJJeXifs6WZcpSxfmI1h/dI0B9k9ZSchcE97SBcy9F
Q2csTyByQPpb07bWH99eq9wZSrf5F6nFW8Gov9BqyWi5FkEJgby3VtiQivy2t2GUzQqHrBHVREfA
D/zppkPaEMl4R7x3hf/5BfMTy9vy8v/e2eRdmUnxD0U4bIoKfszp9B3OV2CZxDPi1VJI49yFUPYr
6RygGpD4//zl4Ed6O0c5T1PGdcVO+yPWJAAwh3OLPMcuontxGYcoNAP0M7Hz0tvgz1qe6v1onUZg
yVnwjJiBaPMKR7QM6/yEP9gbltHKtGan7BlBoeflvieeYGC+C64K9ojUoeDehvYkX6389w0YnkO3
3jlhVQKwYtqof74lScJF4VrLedo+Rm3S8dvO+H/cB1k0OQIeDxAvBdY6G9CXMagJx1g0NmuRNnFf
1s3+nXIssz2j+TCdj9p/OxwCn/etJ0wROmyPsNrTdgTTmhl5QZ3f3WKPl7SK/t8eIIUNA0GjiTb8
lyAIPpJteXQ9PvJMmemsrMs2xkpypAtqjthzaNLXlIE8QrkQDbje3zL7smOu/v3TqcTQ8qcdevXz
KDp50ZlNBrikwjRXy6VqPZowRxy+TF5we6Ty031+RbObjDHGIF5IvSmrDz+p5HxMwI7TUKtQQT/2
DnoiHsIz/ZUU//4VsSyGoOwsMg+IKRCldIN4c4LdvO3KZ6ApGoAfFk7wPjQHXT0bdmcVreuhaHRU
VAwLZEErqPn+i3IFbp2tzLG+Ng8lBiOgbv23cFRUIl3bZvM+2RkmR6fWfcieoNzXme/hwOVPuWA9
LGOj2/vYO3sZcojht3OvBn0NqohEik9EPwKAGzuNV516QZC12mNs0Pt6HlEf1nQNSFZXI/oJotNf
eiS33gw5sdKkCemWSWc0kKvez+f8McV5/4W4rN/Aq8dEgBFxT+KWxZJa5vRpnsUATwSIfrC3LRUU
V6U6HQ7hfTDiX7d3tsSyQyQpNxW/Cg30T5FvgJr6IrC4+98bEtE2Hsk4CASgyDy1KsqeEuLswzFO
j9tx6eLyL2TsR/qvYRyjgm6W5sdrZztKO6B59UDQtwjq0IC9KURUvB1Hvi1SyuW0wzXJFupwUpm4
trjt8RIDVcmUl/6i3w0yMMdmys3I9s1810O/vy4RCa1BnLIaWNmJIeRKrXZbs9MCvHlewXef6tF3
5c8H7JZrBR5KgJICsFHG5BQrg+K+NiZviNRslrVwzcd0Ld6Hdc+8/WtaayKebs4KgsXY25Dj8//6
0kcQVGr5FLSteuHR0dCSXzVrJDVXZzMC8TxZoifGGMmsNdAcl1igaVmDq5XIbyUneyoyxyzW0znA
J1i8P42Ud31Wo1jyU6zsjAvEmtz0DdzwA9nAa0qPvoQRDSPBEMfYPY8ZxbH5TiaR0E1cHOPvWTHn
PU1vXpFeOa5QFTx4lfnEMkYAeHl4z7uOSDGp+FfhoJmt9wfLM/D1wYs0VzdDY14LYYCBZySKyBRC
VnfV6Xp7GpX/5A7UpWMQuFemtLBDR6TnyKwr6jcRSLCHgO2MVCAmCnKxchtusOUEdsVnK86Ce8qN
VlyAZiVmNCBizO774xgqtiE0z0Kufl9uPL2tVKMt2xctcQLudOAQfQnCC6hNGBGbA/iofMQSRYqa
BkDHvOBZPD5lSeQ4YQZh3hYvdvFytnf46BwqbZ5CpeeDl5H8EwPXCWHwDp9nBvH5morxVfVInH4J
qHPccN/dsmB9EZ4jMR/BP7fqupR7syj7p0rIDZQgnxQsoppd1HfEVmvvGAkzD1JTNzXnuJa2ultN
xUWN/UC6K/MNc944eCPE1FU0BeK5FHIvetkwbcJbnKSnQBB28TYvEOxHjqdUBC+fjF62JkdEE9nl
NPbJBSOCMsygMpV006ZT2Ws/aAnJsYTUTHIbdNOQv4EdTT/PaJt/ZpkZja+Oed66sU17e8XT2wnp
WFewLtwpyFx84E6OYp0/+FT9wWGuo8xWOkZcNa8uVJzZNNXwE8fHFa117cxP8mZEKG6F/6JbMUup
q6vfgKpA1ga1nTVBMpnxXAV/spUtCZqap5cx/hBR+4LAssZYzPksJDoQ5AtvZiBijKmGlEGzFGA5
xsRFgQhvgkM6Px1H0DtvG+U5140sIGkl7Ay5NZ+odlCCZNrdZLX5+bm+RjG5pkQQlRruuDF6qCik
LGbYvHTA7MXvGmitwygAZMZpXxNClrrw9vafqoAWKMvXDi11IutdxjzUI44v9l/WscuMDslhUgVv
VqPEBBBTN7jh15DQVYGsALXrYaaR6IM800x3lE+zj4PermPlR6XvtpDYs/7Iyz1veeChcudsvzVg
wJueYW3ZUO4pWbL0HrPfswCcyvKuTOecrTCMZiMh6oSG9Zl9YQpGjYrHpSLXoTWThEhGGW99jA4n
EZmgIQRBgrVglupyxCoWjEXwxvPdOCBZHn2YhHmp0+EFWbdsxkgSVOV8LSPjLGFBmhAVHAk6wCdj
EDMjopdLcZqnE6oNIcCw8dl/qcXqEADbCmWPvYIjcqI1ak69S5iZsVO994QK746cBq2P6i2vMwM2
dkiDTLVT698QWUtMGKJeT0ToNBbG2KOF5rRN8dukCkQPHsjrWQTbMPN5v6Ac0RigXF6iLZw3otr8
65MqoVmHAKP7fHUkp24dGuXKwaR12onMhBwl4TVSO3zv3YsUHMm4NxspxAvbizNQvBe713aFwJUY
xclZqoo8f5/CWmOuPKbPlzAg6WxCyKym50n8z1WwojzK00B0id+j2LgbD6hPEYJpAljYoCOFcwdt
tkhSsUhosQVvW/sXS07ZuHnwAXuetNOEubJQx89X9OyHav15qzzzbWGo0pumEBKiym6ZyW4GRrKT
aXfXP1rl2+mys+s1/Dha7D1bw2OiBEqf6eLr/yvGW1t0X58NlLd2xyEl67bUI96Wf4JJ5lIpN1G1
f+YcjDFqONZmuzGV/8Zb/Ik7z72aFD7w94XFmuSyzzbQaBj9sjPeRsf+o2f6BLlmotmjhXTNTXaD
wFwIifCg1hzXiGX3bCYxvsH4g1MnDZqJ9PJG0WSndyc/Gn2n1aGbQqaUun5LADCwsQ1GK3rezkwd
TZtbUWe6ydP1dC65Nuxf3djw6yrhlnE3oSFPiiaIyrhGJKvtnnkX/a654hAMu+WwICCTLZbcd6a8
d84O4aaq/h1gGOoUNBQ93Fnz5v5x0Izo0GAzOS16/RRcf7Jqge3wYvno2dWfvfqygGh7l3kUpiln
ytWpjQ+zQ9fye50HKY1T5DF1Aln2EBaSNyK+3yysT0IRNFPV8ou58xNDKR6gVaX6CHBPtj7pC0+3
VW0diGMjB5wxJVa1Xadd3gWAXY8kTH/1j9yJiO2/J9j/5M+Rg4Kdz3YvAuCv9aQJ3rEMJ/MqAfQf
X47swGQ5qq97JiYLN+zyGW5ANAGDe1/dQ3DIIB+6+3CoUwsn73ugBSDwde6FtSJ+LXBRIBMPl83P
fbZaEgVVrIxPDxAS/TPPEFEOEOEHyc++/UKE1maDivIVFbW8m0B+O5WoHf/GE8t908cSGC0dq90S
NVFfZ4Om3fl13rjy5X6rXxP5Qs068CcOGxCPtoY5Ega/sJe3ssBUvrfBtREtSfhu/eZAfKxNi4y4
aeHbubSLlUvkj0AZ0wFoNYupjYO1rLApWliW87K3Eiz9PLSg1AI21n3JWvP0/FMRvaN/2XRJHmty
7HdUkKX46SJ3RUHJt3lEOM1VdZ/ERIBEmDX+1GMHR8TftpIjNreXw5u6B+a5g30b/OYQQ4h3ksD2
kVI0E7UNxn58eJRNX8UeaDv9n9ii39Y6XYbyekdp+ZkDPuLqflc12vbhM5LCNURsMFXeQaLi92Rw
wlyOjJCmmahnnDIP7MBIfNGmM20zKC1OTLS8F2eU1I+VvTE6TCcikIEwacK9xBNSfL95lusfC+95
+Dh/Bq59DlkPxKiwME/thmI987m0Pf3nY11LIMkuxu9Ex1tHBzcBYKDINfjTnxWqsK06lXN2S82w
6emSRR0byG7+5AvyIpzt/2p+DzKWMfl1YRqMcCqaMH8JCIZtmlJr+BkUjh4xeEnv9/GNHZn49JPZ
JFSqbsewZCMVbA5yIrMUiHIzUZwyYhvuw5q6jphwj1rwmjcl+fe7IzdcOWKixpYZtHdRZ2aWjs82
sPL2GcX1Ev02Zyomwzi1T8/TWU+lpwVWWTvWJ9Nb4P72cTJgeAB4wmHNl548/W3mAzDAUtE8KVfI
7wzlxU5aLk19e8wlKW9iOEMzPYHAn+gQCIdiy2HdB7YoBZpQm2HoY0AqXzYCSiLOT+z0MVSmv89R
gBNiR6QwTSfuH2HR4I/RP5po6ySD4brPvi4EKOrzSW5fivnpUsJWwuaWX+noGCfXlTxVGShTVk87
wxkvw5JjUaNzIzEkPCV0i01N3J33qxikhXiwaQEojGlK3mCQiTBrVBGKiYcbgEuYRPg92bh0SLyI
BfbjxxnUlVldNjRkfrU90K+wUyILQ+X3Evkmdcg3BbTp+OmWPzRmHWgZdkXByQYj2pe/3zZvX6EP
OTTMhqs37nFBWESBntor+Mgh6Bo4XxOuNwo8Yssetc1y6eHE0VbQ/ppIug4OKyaE9ASmMR9yHmXk
6eR5m5PLXzTARMsOWjG7SHHp+dOeKSEATpsMyjS3/a2hg7UzLOKbJq+kAl7XdH7/v8j63Rl/8MSD
xdFGdow4s7+w4glTfvlBlORsFgendLV8jrS0aKEwpzVOimatSueZ0i5aFj/8Y36zvFziaDtEE3xg
N/DrJ1f449Gc26iEXlvKbRtzIgZV2oBMBrYoHZ72Od+TZc17pBtIcwOzWQpQYqpvchmLZpltJhq4
2Rhrk8J+FI3dYsDSVQHA0j8ubZbrQq6YpnvdsgpgjVT0KUs7ChT1rDeu0HQlt8VeF2Xrb9EqA3B+
bjaJVtbdYKckkkkCaAIo3TFBQw6462paqEDD2vccyim/zzirHrpp7CG+Xe3Ge3VUm6E/F969usbn
JDFLKp0XDVNaFNUv3fnpla7MqHVw/EFm62O2ZmSCFNqkCBiujY4MIxX4o4oIq6zBKuay7gq38ONu
qSoep+RaRVCNdM0I+nt6vKp4wV+jXJKP+1njZTnnh+lywTk+32hbM7ADfDY1YIcIgzE36ipryKa8
5WsqBjEEW91Ads9z+92ubbRENibNWHwzxtJKA8xTuQq/M1sQq1YfGAG311jpwXl6RCuetAhf7Knf
pp17tn/53ggDzcBGbtSgSEERGTU7m5YlnZvtTV7mVumU8CMb9p3Ic2SVBnoqqsyI4lMOiehkMYDU
k+PoZ4SoXduVf87lOi3yFtucQLZTLTm04l1cuBaee1GP5fnkq8OuZcdWZTw69JdptaUUA3fYxzmp
4KAZw6URHAHchv7nSfB+1aobBEDoxHsySVkQKbcp9o/VfESelakA6n9jHcvvWSYdzIxZF4Vn4C9J
WsTWDXrlGbTeSkz8SptBix8Nnywim9Y35PypBx7HddE46fQEIQozD2fIXWJGlSHDQ2keViE+lWM1
hthkMQQvGRFBmD+arM9ty8Pw3jpUqQQfMighMZXdCORZfRqhV9s9X0NSPYYEGrarKhOg4oNkIYOQ
C7VqPs+j7ihTPAd8AYJ2lprHCo7viNSl+GFplGrTLuxlLM0ejRxw8kno1aA2zhiqgU+lUmWdJOHE
2mRhI1WUAI1zCADZ8734c9hCqAT7J7olSq5f0tZmWaJ8OlgPdJyjB/2UFHb5eRgFjOArq/eIeqE+
dY21ZKaR650ptMq4sCz0O8Bl9lbVF4v+uvwnCDd72+s1Ff4PsW8fFUcOCHxjCY8U64Y8bAYx7Xf5
S+SFQSqZc9BeNn3gdxpUreMtObuQiu3W/0KjC8k0r8wJXQPTooTC5dzSNSfUgeEr+XCJ/a9/iiv8
rYRVa6HdD1tZ7MJodTkyt94ltl1ROtGIgd24j8dIQH2/ao0muF0SLYrPgIaRFceBb6kj2U/E/5Y6
tbNxO63KeVjEEF8CW2GHsGIWI0+TEPHJ/Kg6AhGWDhITtqHWbE83FQDUP7UVRDmJxy4Hhi9RXY+6
tDG/dezV8oTKd3v85yXdetM7znHuja8JnGSl13wMorWeoPwTYO1uDZDY4SDbXklD9uzg1c6EM937
ntPpf+uGPb58m5yiEIuakR6KNJpmHvbGEiRtqUpR+ny+4/FZJpu6hg/jukiaMui0aY9bEGsAL/M6
HTkrAKjlsteFR+RFajd8EQDLNNTT1MeevpOwWO1pLm5bh1GguzcEa1RUWp3FdXtUzxArFZxWEW6v
+paCAkLOeBnpqzJd6TBnfyYm6mS4t5UpQkkCh0fEMxeWtjtjgayQwsD+fEA+pwwe1kJvDHJs6o5J
aS4frAsE69055SmaGKCcglNE7kYH0P92Py/giVcs7F3OStMxnBLxeBvYTmGok0pOyW9J3ehTYBoR
GL7RF8wQBqKuLkJSbeWTQIibxEKOskoSr8gL+zYOgpErEF1BCvH0ikklgQax/lv/kfstogkJcKi5
cOp6Yp9ovgyaif9N6b+woD3aKimq0HLDvR6C1HNnxJQxxHVjEvz1cIqVR0YUrAg6Pfm1Ls8FWiy7
iUVU1+8W7MJqr1K9ByqgqF/Jt9+VWehrKWtYyW3xMgMrDONNmdHmRFIOCi8/tuICKVw5CZs0oJEM
pMQ+zUh4ptmhVy/ZcKzs9W068G3igrtxygvHUq7PkY6Z5TCGiq8pUjZoj7IxRMqD9fMiouM1klHP
ey4WXZW4yt23coMmUPJQFOLvOB2dwvKpodmW1Tmw4DDIgTKGZyH7ECgqeG8QKluiS8sXPWHUD7do
R/yeO4qMHGDHC8+wW7yH+fwvbzADlNtv/3n7R3ATGcgSpMvZcWTm87QKE5goKhtWOqc6I4x3ibAJ
JHMi+jHZcA/He/CRTXtyo3cMLyl2D8WW/CL6l9o5qtAat7moO4vN1ADgmkKgMAx+/Unf57C0lbc0
CDSwKO5a73SImAxmGj/G2UdhRp3+6n/Ax+qkvWHZiLN+wm2VGvk2ekHLXwjzeLcjvATCL7DZ3OEU
jyZ8wVMHIvxyqqlT8c0euTiKe/cHwU+uMrQG3ItzS52gRZitJD6f2nkJgr9CHIsLlW0Otm2yM2Nh
teVXg5EUHsbnS9k9SJlu0EtPjDXszeDQ9D28dPu0CHhxLCdGviflDb52VPiIZQrK/TWfAIml6ulo
JYLkK+VXgjPXqsuO18oqymDqI2GjDxDSHlXL/wwnY5Cki3Cv1zM0GXX69SH/TyvEchK4ZWffN4ZI
qnPcjnbLeBeW2Vup2En3kZFLMWLt5iZA/Rx0tFv+CciSKFT8P+rJwdyC3XT3Ke40bHd1GLpW2yK4
+INwzHvQg+lM2lNxAFVhfOKlMnHhMUZ5YTYZ0IEFENGFbc8lCy3VHjTFWbVqnCfuk/W04yno3zzV
j4sU1M9TJVa/NvxlEPxtsl6JjSwowX9Rc16uTXQcCDihkkogXZMh8KMeNvv/q0iZGHsUcC2obGUk
uNFrj+2N2tvf2mKYOh8bcBbNnEoV5tgGhbEJMS2qaznN6jj0KJW+6hlKpSOnLFM08vND7DfpdM68
gjIWV0aI5eXKWU5KaRKlAO12WwoVpdl+MBsCSFBxrSBBpJXWme7u+HnevNqjDWJBMYIYGzk7gMPH
dbte2dZtkrlza7Np0ByojOwRXsLFXBnGEX41G8KGiiiBdWb/BXnmqu9dJhiwP3sJ9wqRVSlTSUKy
5YPPFth+6r5OE8uxrRi4HjLdBpzvPMcpBlBjtCAvakwU/yvPzpt9+lbyJWNESWjbo2qx25qWSbjJ
0PHOWPRWX/CPG0NdMuJnoaRgV/QfyWxXpOnVlvHEzzvHXpvv1mElRQlOBXro9t6T+04inx3WFPyI
LWvu6wAr0Rqiu/SjqKr/eWagh7dpGl09qNUCfMVFK9/GY87MxxH6axZeu9GkX6KylO/jh46gbn5C
jwxwq5Q9AIr5aDHI16OT9IiBqv64LJOqQBiI/KtJypmXpgA9/l3iSlv+/w789TE5IfngLtw8avlk
Etj9TOJwl2DLBjJJg89RHk2yJLrgB9F1rit6PAMsHCb3g1PJ4BSKYVr4uSAeFf2bjt/tlpDKbh7C
YAXhyD5tEeWDbn8zn3+Vczf15ovmXviZZ6Qw8LLLu8QD8kzoNMqYMU2m76QbcgRzUEK9tp1TLa68
YS8IXlxfT4dV2u+5lwWCaKsZGHstQDoE1k/5cNOEl5Sy20BOJbDbqbSi2ccNRl/v3tbQzA0BlYdz
MPJpodRuGGupV7SSnGNXnIkRziW+rEY0NES1qtb2+Gy+2UrOFKkopdW8/v4K6SbQwhTkGGWbMGwG
aGZfdvQQ5mMSUa4DDGQquKjreIybcZF6sqrwGZUEhsu4YmEHc45f1WVOKV+z2VXw/U1aRAMP9uoX
jv4BN9U1vg8v9SPPQTUg9E3UDuXZDuKc9Q3sd2v45faOuTeudTMIpX5t+rmxc2QpHj+oCUFDGku7
FBW89hNn6Uswk4vkF0ENtk33SC8919p7ae5xsUdiX0FYeI4EI45y9Hpci+bW2YaZMviiyVsMPpg4
P6s2FEe1lm2sSdNjEwggoY5eMzicxLjHpAjOOcsVnc0NOIh54Nb45fIMfbLcfk2NWd2pd5mUceIb
IGKMdFr/3CYb4U7iv7zzbCFTaqf1Juf8DECdIUkI0sJkU/MtXCH0Jyf1g87DPQJRy8TzvEdQIAOF
fLKJBEZptWetGH+PAJzOE/5WpkzSwbW3XMLVdpeHA7NcZjCUjSApmF1lLXZF+eShatwzTcofhnKn
+uBQA/LKCDM6HgZsiYKvXAwM0GynEAPFsvDxST9yAUCWYZHjHJod5EAT0HUjqVEcgZAlngzUFtge
PztWozORwErPw4YPaLMePG7NUyYoaAwI4XqS86TFALVhq7OcACKydvx7vUAd0j2j61Fmj4ErsaiU
cWcR7m+cOmjUNEp3n9kzYaupZVW42o/ot0T7Hadg5LBOkxPD2qXdG0JYrKWxUXfxMLdm5dwfNQCp
v0qEEWFlciMgdddXfDlgCgUMtnOsDFUS1IOvs/0kizJC8/ttXlKAcB5N7zXr/bGHNAsPb4INci4t
qLaMefl8worv99zYEzkgPreDxcvhNNkMnAeGYUrX7h3qaXTlMjQZuE4Jc5/sWSeyWIgFn69Lnyg1
lgOPVg8sWKgCA+8N0a/dOY1gex/lkczFL83QL8fcVAdI+k/cufYglzDxhDLSqqXPRPflyd2pt7Qx
6iGza/iU8pY4Adhyg6XM1Ml0gdF63RHzf+9EhfMPt2WEcxcBt4gPZO5EHikdsNVzvscaqRy6R4O9
eT2JIDNYH+tAvgwMbTcoiiO02OBjWYtDXG2KcYmn15g/R38uWdCxJvt/pMRuHE9LeQn87JsXgNYi
oevzNEphofEBV8LkBWO5RV+apmyDSpaYgL0ueU7xW/7cFVlvBz7fU50V6zeIXVar/oEG5W4mVh/X
l9LCq92wkSgdUFsOR6PlPlZgDXSQ5cUnVchY7xzkefmig+k36dtiQy3erGzdaDGfJSSpmfSjQX4f
EyIvKKghF56lhHaC7+109ryvDThoxhIBg9MT4GanPdqYAGkJO55OGia4SYRNM7kPcyPvRh8F+wS3
kYFZix5rSOnCe3D2txL3NVosyMJsrrmjs+/HEBWpUaSdd683V6ylhNF1D9/Y4sKt3HEVVNrfmHOK
1hICKFiYpMxIj4BUoffdD1cMaGQOKuFdKyd0cx2Shd1WRU3+jOG16KkYR5YZu6OnDd9xYA/p2uVL
1ZWgmFd0LtWBsnUoHNOpexQz+2/La6d+VIGW3GE2M8yTrkuiz+CmXYUmd3DJlASGc64nI0bZtEfk
XJZDS8MNa0PJGRnOdXLBJNC2F+d45zAtht3ovntmz9rrNvfaF20qICXlclJrZvlLA+JryOvlMiaq
gR+qH/m/i21v8E4wQnp985jt73pWNQfn3RUJb4Vx4tQ7TyLgCJ5DMTanyRzKCpCK7kWWypLZvF5+
B+U3zco9uHioptwxDQIkxNgqEje4UOOH8gVyue6WTKQWBsjZCvq0P8pVLE/PuBbXlb1uB7QPZPog
8xUTH9iNSlhmtezfP/jIcSvXsc26VmS2Y6UkqyGO0OiK8PND23nz5c+gePWVtD0es7tK5TAdIOBd
r98+zVpQF8vPJ9hygltRc5jzZ89Z73E9fgAZThBN+TlrpCRhcRE6AwqnZB18fGlGnNCpsFuWUFd3
01a8aD3kxXlGRtjsLzpZxbzRNstwNHOKt195772A3vHkDX17aq9oztPKC0+0KQmo5v7DMyEzCtbx
G7yhT1RM7FsJLKG5VtVLWFkwPeQXs72YyQtRlZCKqxwC7K9/Sg9PNTJ/mMx686jGFJYnvB33Tugj
FLvu07DSqZlbIceGlXS9YTKPNT9tNLVjlpxmN4/FWFHMaB/yxH/Opc/08VS0Muc8g4D85J3WqQka
bStSaXgCwnbl8+4Kl3cHo54Z6lSGBAreeO5cLH88WCCs6U1G9EIzY21cz0+IoDve6Yy/NPjDDZFo
TIm/0cAwybHvDAtj0oOuEg4uo829HABqimymvzDXtYFwmdPKk5z6BO7LqyFuZW2WlvQ4Pw71ptv6
lWEODfl9RzdLE+Kw+D18W+DvLYRZjvMfyUoFZWenLBKLSQ8ZNcN0UYsu3xaDnIJx6l+st8sUzRYd
KbhFzIe8LiWMKNSWyZ8zlDAUw/nHK2bESjhhQ8QK+AaG0Q1qIbtD0+hY/LqZuLYyBVYfiy2kXW6F
JFvhfNe9G7zAQvGgYewsY+6Qf4obhPFmNqbpZfziQ7BW2jVodr+MxVSgoUFJLF+i/zP6RDhxb/nO
v1b4CETrn/5QWaMvGNvalhFVxln6jS+QwKSnpwrinmOPImghEdBj+kkl6hYzM1pLyPoeEy5EuNwa
Rr8qWefBsx311Pmc1xtb/oo8Z8cEHHcmS2fvQH1UXLdK0Dl453o+5K7juocn2nH3annQTXChHDr9
WYVX99ldv8RrqCFOGPljlqWHUyXytyQrl/G3BuZcjMRVjJCGO21lYd6MA8gImWu8l4c8+zWlm3hY
4FPo4PRLjzQf6x2unhYNO4QZe7cSYEe6md/xW/wp5vVoCXQqKbh7En6N4DtttpYaNlls4dqo1zH0
Gy0pDIBfHxqxqDYrpo92e89Woz/oLf9lE0XdQJkSxhGUhIfduvWYoiXDMgouonLFc8B6qD57cLJW
UOO1OoT9akBHRF9hmvTHPgysMBkqmfleXWVh83zNbIeaLUvkAqJWYjOSrjtiCZTjrR9n7TCTeRak
JNVi78bOBaFXewhquJWB351S3Tth7S2Xj40r3Rjq1kjooLLVlYLxmMRjo9ymMpXzXoo4O90O+C3X
Oldeey6FMpJbujGoIQwZnZj8F9LTWsZDQdm8ddhowPp0WXFt9G6v53GwZTyyrmpEGXyIZ/wLS+lS
kfR/YtpZdkjQR7L9kfpeRW2fdWiz1pEbMPfL8IfgIuGc3FDSfiMRNBGZTERDxsqSeTMlfii+xwZ8
D8nm08uy/8UP0voCdclvr2LHpZveEK161zn2+KLQfGFdRFqQkHGhWmdKPwuo7f8UsEo3AiWdxe4H
JW8RohMl1kDsvbxNTlmvSBaU9RRA2cXZmIHKRB6FRU0hnjRws3A+EC9geTloS56AVwUjTEzzYsyQ
tCy2bNyBZIDXK0lfA9ue8IBcGspnugr4siIclC+5JYWQQS/IXemRy2wxWBLkVX2kuWhmsQcEXtZd
9+n4Ak8kj6qM8k2CLNN17e1jD+8CbuklC0+VfMpUjpWnwrx2+zuIUOuRNabNyVhycaAF4+kp3TuQ
a2APsfRNO+2F2MSSxiqlTQnA6gcztdWlOQL7PSFsaA/wK97CHwAhifxaWOVvacRd0vdis/z9cBfh
YCsKA8SO3a+t9rELRs5vh2Jqgg/E/jiZootbYm3PcJdInekqjxc2kvcF5m17LKMRFji74mjnduPc
CLG8i0w1L0DUMrHsKJMa3kJRm2ru5kRJvpmsxTK2wxdxPGV8Exo7LY1beYXLP0yfwp/qKoTXohhj
PohqL9tQMLg3rlPhu/GEPy9Bb2kJgnW8+86gzi07WAsNkfPEhVHxJw5+ahZe57Ti4futnAZoki3r
26UcxVJxBGVm0EvmZgdSvFUnw2LzyZwTkaBA3qgqW+GGPKAc5/q2ewFT/rvY7OKeAUMnvPyhJ0UD
EUag1qYElKfFiAK3k82cyL3CmBdrAmRImSRyyoP1B/8d2D4NIQkx/71j/8sG6ZtiHGEz4UXwRa4Q
0tKncTFXiBzyEzMQLWhSH7HpFa9Y+h0clv5VgsZbUSjdDcj7s6i3oHsB23c21RtOwVxpjlURjLhq
+antjFZQg3t8C+VvKwbn23cFZIiRdXWJ2ugq7ohEXE0bXd1iR4blhnoEYRlrJWN+JWktCfFHUkxP
zoAE7+LouRqHIQpymI/ux6HlQo0H988o8lOWKTfnQn6Nd/ReU+T9xuUTrVOkJi+iyK348zeiODVO
gIohRXOcW3tZYw6UngtwYVyUFDjke3Bnhh4VgUIUmlV56ErMYndLsMpztOWXBu97WifHYM0/BwMx
yrYaUvzPc7urqg6wcqVjM3AsQBZ0UEja7B5sYJlwJSaDvyUzi548f3SI05+z4EMHQmosPgATthw7
x6Y4gd07XUYopNGMfUptVypS5EYWGcRbvXeapF/Zxf/p6xf7OlU1wie8BCQocqjNg9I/rlX/viKB
qRa437mddIPMEjqBVLDx3irCi+0fp/1Ug6XVurEUd5gC/Rd1L7YVf7OL2XWSzBqTw2dwmofbW3Qr
XHDmaEapvLa60PT3K/DeILkYBVB+bTihoovPjdgsQatoHxAro0buTMjq8a3KJiAig5gQC4LwJ/ZH
jl3x/QaVSwHuA1JKrYqHif+GZwDTX6Ub1TJsqtucf8/Ro9xZzIYaEyHehDNfxD9SRBIfa2Yqu0wT
3EngwmuP6NRL2Pb3pIzThIhgghpZ/59NII7lylH1iX3nNWMljYfKPrQl046bttrsfFnkJ+1DV8OU
kO1bPHpVeJFgYrMLkj8Y03HrtFcJIrjOrhDwC/ybS9hDBZqChA12W4/wzkz6k4TZia7piXYd82nR
gGYd+b3mTJwGgd60CXfy+iqTS3wZrTnWpCwUJkS59jeFuwq1FwdApy/vSuVLF+BNt7V8kqw3JD9P
zReeicvnN6Hvw0NbmMrKiMY9Q+9hTMSIzz2+fo+MteHmC0ttEsj/grBhK9UbwdKEmNmdG0bxG7Cn
w/uJx0/yQZznlzsxN4kPvb7T3HFGYpLw6rs1zutuSbEf6Tc3m41DdSnhfzM7RiCUMt3Jn3wgNJWu
k5K6f2y0cQ96gJxW9q8jIVIYKznV8gWdHaYVl6WxtBj2GVz/bbmzXQwD4A0u3So0d6prYw+KYozY
H3RKJe7yRPPHI7FQr1jGhuUzupf9Pz11pfPTDtAaCbNy1DaWQdrcLHrMXUJrcw+cu6GQ2em81okh
tHdPjOa9tRPNqloRgEP3afEt09AkpvszslEvsMWMxkvo1YKSGEZIsAOOn3ZxY61BvbahA5Srb0Un
B5t6IVc0r3t/qM6ij5s+33ahUQjH9J4N+zenkuQd211RXyh/Nho/Ny/laYM0W1WYEgr8bvRgBgIJ
qKZydw8a4ZooJ4ChDBQ0VrLRPlS7jCI0ZO+aX41nGxsZs7B7Vh2rV+U007eeEbSw/ixcUZhYSQ22
NIbvIKGo08xUIHdXPEPL71rezHcZUsurhw/ikjcofxgBmR4xzMn87GEyEdcictidiBpnCg7YfPq/
I66NrJpt75xOe32p7VFycQwOnhyWVJu2LfXpH8+ghLpBwieZQaWr+02IV24kbxkqDBKRI+Thvqqw
DtIN3DZknYrE6crgxL2Txku8OEViexPjgkosSgLycX1Y+LZIf9IjD6RPCSLEJ5f40yhbmttSffge
NonBC8nlJ98IcAEIIUwzVpqgNjrvtEGrB24WA3nA22JnMuobf4WjdrbslLGNpELp35rypqh0k2zI
21LG1o9cSs+dVH3Z0xEZ5ak3foN4JmX8wTSkej5kArejxBurG1K6DnSvcKqjy3pOHg7FHiqP4Pbb
6urWoOGtZOdUQf2N/itu++TOyNeI3qsZONjtQyk+HrL4JPwxcNPULemQlzo1mDPyHK+qHsP1urhe
fzbVvnksOnAzGdcku3lVfJiIWPlUkItjaVnYnTKk+yS03+6wKaA5fVKvHhlbUEqnvDhzOE/LCk0a
ecmpRvLw1UWfxz736JnWpkJpqri8DMq6s+SoIR0zxz+if14ZbTK9ZYk95xfFk3m2cDsVgIW/KNIv
xfVh3/ZG4nTocufD6Jnc8auj/emUUBb+p5aaaYad+eXqSsEWuh3PTSlhn3zOQu6rrMH7tPEgWvIN
kkp+3HjtgEdOadzF8JHMDrjkVUyUvMkYgvTXT+GlbJZhbc8974Ph34EleU/mmkBOJanLWCSMYlHL
wVXb6M6SWAruGxyYHUbKAbO+kZIXwJOjXEfL14/O9I6/RGZN0oNRY0l+nRoxl9NKUPV7tvanEqE1
hCEDr/trWr7FFzkahTDuKxYqoMc39c49fOoZ1rdqruEHjtqFnuRI6mYaPaW/qNqlYI0ePQaCfvwy
007w7aBidTsS+YeKJEaWy4z2+Ilq02RZbyJ+y3tVfqXXwjElRrij7+x5EVSWmG2Zxvrk9zdi6dIK
CNN8ZIMUxR6tHpZlfXMVQOQxlMXl2Dve+ZI2bq/FI2ijJe309Od+CM7XYYJeH/etakb6sAOQYY/y
KO9SMhOiAVJhetbgBhueA9aqi+04xCvvU9saLgY9HosYj/71N8+FcdL/jKfYV30dC5tDDY+GYcHz
KYNdu78EDEflzpF6e4kb/cZtLI8fZstoGzNy2mmZpZ3ckxJmH7+2rWhf9HPTWqDJMyfXACYmD4i9
4qlSXMx0CQi0fESiuo3/J07zu/Ag744OrgcCpVYj1bu5I//FHnR6SC+RlWMd3g3phSpy4CF8iUJv
UD+RPHso4RvTjUWfekG4Q1mWbDyntASb5tK/2oAoOq5CgAJz+A0VCXHj1hz8yvBHNsXbVb/LKVqC
BC+5g4cncrZAKmRdi/KeqxsdCP78QULNPxPutY87AWsX6Hz5A8WQ04Sz+2DT0Sx5+hO5UfiAx87y
B6/HRnIClYOttycSU8DNRH2fFE7+TsgkoMnbF/nYrQpJlf56ZpcUSMt4i3oW+eFzKZ2CDubCLLk0
Kb3MK4fFsaWL1g8jPdfxy/0motswxBNxggQSvx5hSve11EKRRyxcCJNGPt8tizOx9f+nLoYLslvT
ix0hiVyytDDJcpfTy8UdAEk1dFlTJlOcOl7I4mUvI02+uXuoW/6Nxw5jvOLDdCwgFtL6IPos8T0y
8qr7ZfxgG/E7IYXhchhh9Z3l5JfUL4xG9WiqNN64t6yD+7nXbA4cHtFuqbElmsfT7l0J2P5eHoD6
bGJABswYYkjSrNwPL0m66XM0wax93zhyqyohWGy4qO+hqMoGBruaXYEtGtN/Rf6I3QH3+jq4+PXb
WpYsJcU5luBlyQb2GFKXxmiOmEeWGY8aF2M083qojLihArR7gltlsGy0PbnNzFIKfl7b7GUedyaj
DGIvM9GgNtcyA0Z2mVVv4ZTpEbmoZjZcBqOSQm8/FG3t0J417syPiqGCn83cDAy869vLsFQayZhM
QNnpUmY2BBxx82Lt3lkNlfwwenXQu+lAE1ahHvkx/VIMnxmtrhUeNdT/EmuSrwW8EHHWWqef5GSd
B6aossVAT91R2zdvOxuKCljlV0hSRdUZWfklg75nbZ5IobVsu7AS/jnriZ4UqtroEpo052/GicxB
M8c2UWVfrIJ8YAGyApTp5nC9DA8BNFtj3udwGv3VFPhFtYwNpKzNdIhzQCNwofRBdMOSzdqFHihi
HYVzk+IiihG7GwQ/kLcGh8XsbhZH96B/njSubWFrRoY2XoQuxyGAp03u7ycTFfFbtA41qmpJTbUM
u2TZHB4wbS+hKuE0KyRwcN4ZoHpB+/SRoqZO7BotWbpNQwVs9zaIn6oBqne1A6Kq/h4YinTzEPk1
s5OSFgCUTK7CbutKFX8CD1m4EO2+i9xCViBd22RdWPlIdw8pQBHBtdJafPYJ84KELvu10v3CMw0a
+wukKIplUFUTlzCjd94F3XyO1Mx10Pfj3UHX6o+VxntpBMDRh8l00U52nYgq2UNltXuVeYQYBlYX
/KkjKS+nHAYm177zpTbWq3C7wHpBN7vh15MXzCAGE2lxFW75seDUnQG/OxKNN164zS2BGdAQSRg5
3VaA4Tzrx5BMjynA6MemzGa+in3Qhsms9qRlBf+bu6bFXTv7n03K9jb1o+OguerIZ9BBnSnVzSa+
d4m37Dms20HmBOMTo5QNvE9hCUDBbQ1P368oDUG1ib+BWpiyhAh8SJQRJgXISo5Sc7q7DLPhvS0S
tMM3U/KUEplS1ELLX4FMpmnoCUUI0YqwaR+6Df4ySAo43yb6nKQfA5hi1e9D8lWKBIV1nQgogclR
Cv/FzTN8QmefptFy4UiAIEMWcGNhMRzKKQKTXUbNpQlM4iBly5N+CY+tUUeMrj+4AWnTswvMAOif
8SS/2cm+j3u9G1gPZWLigtj+qxFnKVARFFCxIf17snZ3oWSUjCTivgQe/qIaHRa/SMfOfnzp8xYi
NhE2iEsqXwOqggawTpRfVFTuS6L8EM7ptsCI2aJ9mff+bPRJ/ikIzqfoTFnlG+qH0uiEi5Xkoaad
tJxDG86Z6QqLMYZ0jdozvUcrllp7pdcmb2bTgq2Grk8YTj3rAJkEMlS7qNDeTDvYmnnympV2L9Wo
iCbaWhUvnau6qS5NFszXrml23M3W1CXc782nMHqInVrrMCEuu+0ZrgqwtM+9o5T4XCh+FbJGvktW
E6rloU1aCx5tJoR/f+tDsTLWmVuq3A5KK8AuoznM+E0A3/AqjcAyfMNGJt1R3thTip4voF9kr/xD
lldQ2m4ORCnVSkwr4Ily47XuffwCJWB3EsXfuJSBAPZJ8QXJK7rpFqmCCJcpw0fIbioDS1Mo9KH2
Sqa7tvcjayN+OO+fqVLWKoUCWXDkmT8xBIm9MdApgOb3+Nel4xrJtdkSA/1et91i5MckmZOemUlM
I2/igt6nGJIhMfKhNP0AQi4+X+RuqXvZSyLYG95RojTNZ2z7u8RaKqj6zjJl6oUAeu6E41WOcG0s
FNsoK57K4wYz4m+zTLVvGBySMMNj04lXseZ03P2A9mzh70TEHNcDplK0Gn5eJMePSj2XbgastqPA
x2xkl2KC1fb7T9zmbalx1qg+XPOfW4KwOWSX+dvkCU0wXov+ljRMHGJ/OyCQrVd0vHP/g4mN9IU+
1dcl0l7LKLwx/KLaKF7nw0h5pDFNQC2RRMv09Pxcr77LI3oXTk5GFmdcJPNNkx4lU26ITsPzdFtY
lEPbMHT18aeelvB/XDQy5wfadGJIdqP8PjGNl/jrOl0xWRyjuX6GBkG2OK1ut2xbjJHud4UmHAYV
pjkK5HjYbU/y/Y1vIFIt5nC+N0MxmudemWGMmFVZ22SlWezdGEmoX3TaM+o7rHq3C6aEKsrQnwwN
ZKHkxXX4viiwCM8PzTF/5vc5uaE4RSCfXkw6AOvK+ZXnlHjzNDuNT7gRMdCFk3lyzu5uWLECdEX5
HZll9Lsy4eojlAx5OZWMicpb+k56WY2l/CeMKxhOH9WbjEVlBaIWUTCCzBFdWXvvT8DhJDjvAsY1
HgEc+rtwGy8TeG6egF2ohQINKmb2iXwpya0IhRDJPTHgk64WAQoKGGHGsZd/2iDO4c3ZJQk0K+36
JRR60+/kSgOptiDNEBnam42ePV5Ff5nIQw9wNdCIYXd/OezCAt5LgckPlntq22Cm2evy7xObR08y
FmH8Tjw2tboQHvASDOBgBKvD8YeSb515FWQpvPgZjWtk8DU2yiBVdSr4Uq5SkLISDMdsmHshmSAZ
KZvJZyNbO/YuuF2cjj+nQrMvJyx3rMffq3CQdrOPUOvvANXIp+ZXUxrJbGbqQkdQno7uEs4ekON0
h6tpiwaBXyGAb4KFPfgGDizOihwkSpO/bniB8yxAeTedkXROYx75rgIZgw6Fm5zf9Nisuzaz9Ruj
Td4+TKZw5mYPla0VczhDaUlMWHBP8HNYqLP5sbQRu9G5lrkpKLKNREScOtb+TpOJPPm+L6KdIGAG
X3i2YaoTd2RtqTCGNGrQP5AzFMm7lINNsp/pmwTmj5Oz1pkUyXuyBt0yLgtlWByhmsMC34DeL8cp
bybCduuAXSSI0hcm2faUC3IQvKMjvbw6ahXbfxTBXUW+go9J242AhqJV7nWMeMpcPFsim+qJ6m1T
s2014bHuupQyA9ZfYJx5NPjQaeK2Kla4KqLVGH2uYKJPTDPirWx4AlxrLb7UMe82YJ+wDujOflyL
pybObO4z6MUhyXh+UN2q0/Ook8VzZX9pUIoUG9hVWSx7DDPAtejj4217DE35tDvzziBqaF5tEmrF
aJ4bKYUE5GSAkn/ECDawoVEWrfab4o+AnX1Yu0lKp7CpWeU+Dx4UXrrL9PfaUeC+18nDFBFULGJE
jyoRe6giX62YyRki9GL+kSXFOMZ18NVB8/+/aET1c4OcmifBU/2FEEvIgPr9qTzn1WFSxO2Aj5gj
ZNY0tHdkYeE569dVMpPhmFQYl5YD3CGxrlA3A7cptBa5h6XNx+vfWxMnuciqNS/HZSZM4TW0obLs
JgAWX1LKXlbMO5scaT9EK36XBknndGDGlfOd5VwEBao9Dj4mlEboSiFiiVr82U+mO5fAt86I23YX
mBBH8w1QazSQ2QHY0ZxoOodSPWMiVhsrhAEauhXapUZcHOlD/s3nypJz79s8Dykeo2dQbHefZzj7
2VhkgJUUAdDoIEZv+AfSV5c1bq16AD0urDulYK/ry1U8qRqhRg26KS75ue8QaDeN4RU4Hc/ItXOk
bXDyDupTWfPWd4LIIvgIseOe5YmMbbdJvnlg83HQ56DjGxhhR/xLL0hYh0P/k1btfSipRK2aZcKc
D+blny+Hs0g3jlGZcQnkywWBy2R14PVGgqJaDAk/JiP7vs8Xx5xyJVNoURHMp6TWzfvhn70jSbjV
/R1N04m6cwsmjbzLMolzexQe3sevNwXCfpL81DA+q9YGOsznxqpqhhBRPseiDe+hi1JsmztvRD0d
2tfb67zefl8dtUU8ve80HiLINyOaLEgufRsxAcKdyKPMjBPESkm8Q8Nxg6GOoE9A2W0gUTos+um6
6KrLLByJDa/jYmEIuQJ/raDSnajSZxGQrSFrQg837g66LBTdkmZk1oVVgUTGkRJl6EHvdTtWlk/l
4nqEa0dKb45LcJitkI0GMKJlyHYG9hcrTQyv3dhC86zlig5wj72t8TrmMbuvTQ6F112sVtcSwQ6P
PcyIv4Mxg+7NkPbN0L6f4twwdZkiuULFA64Q1AuNjCRLMGmv3PZckfKN2FQzaXUIIzGW4db3okY0
PUuV3pd0brbEG89VbUI4YkKIK3AmCQZmwkUIB4t3vj8yOC/gHKNajdshn2pYHamGRjh6sSq71kTH
Mbi682Rf/MPu7rqbGMYxsttPMBhdfqo53sEiXEla//5gZ6R+oEzbyjSiWYkYAGAHKUnduM212bRq
0A4d/61u6WlNk+/n+In6VZZMRAEduTgXzHXWjCgpv5k/VVtWJGkRCgwXWVbO8+eeu4wwxatXcE7p
K2i7pGw3fTMhceLXCxkf4V6RzVdbbPif8/x3YUqrW9HJmoqppPF/ycowA5w5Pm+F9Xvvl/Ur97+G
RaH8tiUaYJ9XB8rmsIQ0zVzVi01L5iIc76uWo/aToHnu/qStYWsSkmXD8lvpoAN9t5IJ7ac5s/Bd
/sA6x+g2Pd3nz0ZsqS4pXyK6E/P0j1l5GM65f9dczbo/1UnWygyS0sh6NFmVcwj3jGSQjU86e6Aw
mKDS709cy96ftlWvkxrC4VqZlyZ53481bOuZsqkFFFsfyyaQPSe/R9M+nPbX2zS5odpyY/EQa2IS
eWFgEW9O5h0WZA3/aPh1p+IBYxLEJ+TQ316Cv1CenKKhqZTgUKiMp19hpjJzqHU1IGOUzCA0neNB
2hkzH0xAKY9Qw+i/p/au1K/5czQLpnIpAnYrFnCebK6xzsNaCrO3I/Cix8eBlcA6tH9L6KrinfLU
XtOmU99r//95tefd8YzRhcNuqvnZTHcVXVEnUKQgAtVBvZyXNag2yEWl+8KuGruZlGo/VFQy2EDK
FsmL+ctcrMqGI+Amz3GqVxBswOmpV/znUIoPRCTdNeIbu0T6kEWgRq4igQgzeRkkA7j2+x0Dytyj
211Kn502BO/FOzXmRKtP4I4YijgoUmKWN8q5S2ZsOfuh2Xla9DI4yQRGOCCEqc/6bFAKNCUOqTo7
kMhQOhjmMSVrbSkTtSlng9+lHLZ0Fg1wsOuTfmw/UZl6X5HBgtituFW2SMMyW/2oxQrPMyei7GlX
4BuuegETaMmc0QHEHcArdZh4Sd7/EZDsXjJLWfpcL9k7/hYobAibjcJ+TWjMZu5JzDoNqb++RZSS
YgeWq6SM5VR1jYRq3zJRnXl0f5CqOBNhQOVOGmSAKgJ56mTZQw9gjA2d5x7Cuz/ROuFiqRLUM/qY
K1ouJpo41NcV4Z9mPDTZWdoKT/w/jPMb7YMHQ/ZpnCyPQvMtCY/pwDvGf6NFF8MoPXGKxyJLPx4a
4tKzmnAcHReKurLVZN7tsVCCFI/z3KCG4LbLELE6fPivNQOHqk2s3FTF6V2PDsXsqTsrQy8XlmJa
GrXxPb3Hir1/VBIVRmlZW+mRNvg0vuPPC3JfpDHcBR2IV3mT6Jooh06u0MR+ZmP2iPn+E7JQI4XU
hpCjYt17tLI1SOUqUfYStvJuzr+WUwH9XdXPYa/XHFSwJETQJUymNbqz4yi4OLFqrTu+/0OM9tFd
/bGjnbE3JqJDhNVh1TjVclBIX7Xm5kLR4qEvwFjy32seYH97CLfN1TgwkY2LvHR+oEm2O/cjCCMA
TWyOeo1UWoHOdnjJ53uRpsGRuhm1Wck7T8qx06nGDmbENVQUqmL4jWjg5cYCTPAzRs8fIm0goeZ3
B+0rLrKa8RJvcdY7N4upnj8OEwSX2iIFDpfBVu2R1pTyWbNhiFbhEreGf6lPTVNLwrY/Gl1iH1jP
Ia8OUoNu+Od4Uf/sUgnrtcampgFVA+SKiSP9PNodKCyzc5mNX8pK+V0/KxrVqU+TTbbcm5pB6Dm1
02uBWKu1PCUkha360Htfjo+8rXNeVzNZ4LbbORm3UIiXE60o1FFl3ZcCC9/mkAzpPbG4D7gYMyI7
O4Li1fd4hmhINCTiUHoA2SNH033ifFCHPOrsUFtfXoE8+ZhklmiFczO1J9ccURGxXsPrGLBjUxxB
SAScq/Y8engKCIj9IFxj6mqD3Dx07B3/4dOtbqFwY7DS1J8uBH4RKffqriNWDAOirwf2MDE+C/KD
2hL32VX9NUD2/vNzlzUmZY8Lfvxswif/Mrv0iu5jrnQQ3zuULr9eyIur5vAJrRBqw7HcY56gjvju
Udsic6XQy5qiMeONWgk85In7hcbBu1sy3T2vNGP96XVTzwAD2TNRM0BkwR76zsK4VsAWspBmC6V+
ooH1je4nMsJ5i12+JplTwRiN8mDTsgSxHLcZhVoR7krR8gkaQD5yA5Ivi9XWlTZZSZWHe2ZkbQh2
eL1b/gTFV/gs72ty/fwTz2r+XG7WlhlYsjVikJuP2dtPHIvoqq2OhchDTBSwf+3kEk4LPktMkIQA
3p8wpUpiL9AOCuDQt1IoUYSRyi/e1Abl7hmDEaCPOqa6HipYNwQaSiv5fPS15kGzTSib0b9rQ8AR
FoMiIrGMkJ57k0h7OzvBoPMGFAp0yjV1ybEF9lqp4W8dTpMnqu0AEHZloKcoGIly7iK/0EO6zWvh
4j7JVZ8hMQQJEaDATQOoO7J+RLeLvrpRGUFbd0zqIVq1aiuvM54ixH6F81g4oKTmBiKpb0p1nhoF
NzNT47matEKQGjVgvQ4EnC9Gkd1xZdOLx1uoLFgqp6hMYXxyQtPnT0w/gpBaizkc/jdLfdN7xQpP
2uA7lWNOHayMAWazbuqkjO+f+r/+EEIHByrtNNyUg9D07Bde18XK/slvBAth9g3a22NjRjG3govI
vJjehC2P/jNLmJ8SGFvJuc9tQl5gYrvAaSbUE3tMQQpKi6ld9mV9QKrQwbvF9EobBBsgAKAB+2hL
6k2A5nbeeM4gT/Dsyyjq4QP87nB359BdGhHtk9avZmV0dtddY4Lp4z+Mm4Y864ZV1QepbHD80ef5
J1A41lvYMo+gAjpbgA/mDMYGQQ0Jm+opDXhS6hCFYJvvbGYYWt4kuR1vJCzVdlAjHk8tb0p1pys3
fiWp6ZzA4UrqJjDBiGiQIIZ5LLJxx4OwpVVi3L7WVRHA8fEoWxujUUDOLVCTLj4KV/PUWbwC+/6K
N+1vAqLEF0Cm4+IobYOxd/e3NYhzucxxH5N798Gu6cqVLjC0sc19BvD41jZbbtGMsBdgFYF/mkCh
3vJR2PkqEbGz8jgKvV9l4co4qqE69xJTJu3WuDf8E1TtRrdyltZHE/0nXYYGWmbnN45GG0uYsa0x
FBlJBCagOPSX1/HhVW3t69CNjfTGrmQ1LDzPWXmFDapz+c7vwC9tsAWJOGcVcf7G8mmSH0TDsVMH
2nVI2XNxBVbgchJ1p4UO2bwhdnFqFrXMx2GLSDIIqmgHmDCHAVPTeT7F5Pc4MrX3lE2I4PBi5Kd9
rBve6kEddGzdAPUyCW4uN1GNjlra3n4P+OD7ktyrB2nWLOi2AOauBxpx4qWGqhcJiZP5g/Q58w3E
PrSb6b1SFENtbsbJ7pcFylcjxUJInYvu/j0J2aHfhXdOE6v/8iIivnJ4bhQJkmP6opwzbMWcDLKq
LdHGNk80UNQcbWtGyiV3Ex+l+NdWWD/EUigLSJm17b0bR7sM8d6AkeqJ8JfZlFvr4Dxbs6JRU8Wj
EaRAb9eK57Sc9rNJSSiFSdVclfk9bRhaWvFEFvkUcyDgSqj6+hsf0ZOsaHzait/yRSgy7a2Kz6kE
zwXA3MdzfeE+w7UELYh9Xtq1BiTm9sVmudDjr4tK+FW6xNynBGqupuz1qTh5q9tHcbLlitZQ7jvs
q4hT/IgrMgl8W1JG2Xoqnb9vC9gmzLQfVX2+AbcsfGZ7wJcHN9npQBgQRLOI4T0KgOFnvjjgjVHp
faDXRgClF8u9GWcO6EYL2Ky16+6IUExrxc5K4LXdwbGfaSwX7GT/g6+7VCBg3JQcdtXaFtxTr44u
IDbLJPQkyRhpn1lPLiW13R5g8PehVt0iuySwWwA6UqcU8Yj+zKHqdWcuFtNg93E4Amhu6doGL3Gn
G0PHwTq8H24FP8175zGlxo24/zt2CAegUdVkTfN8HhOoJNhkVXkGuh+3MdntabTk7ui8vBS6LVbG
snDiaKxUHkXaSDBg2aOSmOFq4yLv7+/KdndjXeg7ttibNkbN7exvrsn5a0881c8E9DIR7i6o/xuA
JgPnjcqPjrmte8PIFpCKb9hhiszBGOSbxWO9CapXnhu1bV74HKgH9Cvqnnfv2YEn427Q/5C/w9Kc
jfdtbdMjDvoaWj0SEHqiljxXhVtE7QbtCv45LIoEMLMxqX9eSYgVrWqUijJE8zsvTWH4madxRVxG
em7rh0XMgxTTu2WnZJzprGSd+eBUvpLKfJeZ4tFqyNNxxA0XFMwfBnlwCFsoMglnWfPRRFPx3dtE
Jq2I53vOC/c2uhUPqDBBl1qaC4Phm4itP4ihSzXzxFAvhbXOmj2zq/NaNYOc5zRN6YDVdtQE43Eh
vdgxj76lPoIz7DF93yr+CjJbbbrZ7SYpryQnK9ZGWW52zbRYZnwo56mrpADeoTgqwnBFZZ8W4xZt
/yScZh2tfGcuhxlaPdPAGWXI+ve8+TtEZ/YHQhIwR/fZw/tJHXfia/AXhKdc/BMGndVRp+fKME+B
u4X3lUa3m05D7raqy/Aw7sk5zxM1gYa3bXcuwErWjwlyzqClnDkR7IxGO1fto8G+5flK00WPfudn
mOSVfgV67+4BkVmj3pgOqgXdUE4VFhiiMx6xByXnw9K+DshpKYap5Qs44RTomfrJv2mgzmkpM2wS
/DdffdYfrW7cEtmj3EJQOVMetJ5Lgwv1EOe3fbz8glh9nRYG1e5rsCYE2ULa6R6ypZBdYMyd79GT
0oImoszmz3JysH50KWLepP6tS4QJ4JiAopCVqNZ46BmS7fSwIdWzpE6BT5iNthtV9U/eWlok7clP
IsIhQ/pqJZt2JDTEdZagR8Y4iHVSkVhsn9aGDVp/7y0fb5Dr6yDzLXGfzE3QKFjc84mGf/Nr2sEP
v9eL2mawxokrDa4+dkwHUCsIyvPIk36Trn8lAyx+shDtHeJpvhWn3Ah1kWLMp1HappifhmOsEO12
OZigAddzMkCwwcO/HAeZYnEGXePIpmc8da3ntV+OpdRESctCh9nG+slJ5xXU+Kg/U5zD43qj6cDV
FIbwmfFBhiC2iCa6GnjHbIwmfDmEgRmh6wVj4yNWRRJ2YPkJHwrkj+JVOTuXP6GFvNxtcqOS+WhV
zHsqUnYZTiqpMoeXmgpFhf8QzdqytOrI5jATZG3ilBZYb3XLF1euXay/HatbQp/wmhsmHRzTyxSA
Au2duaO4n1eqI2AusE/o+XrOAZmEHDss7oXa6rpgadGGyDlvbM1qfNoSipaknu3KLAZ9/x3OJiNN
ygingSKyFW31ezu2ZZtuE20VvVCMqu4CSO3tFKPJhYy9TOLFrB9ccNrt4xncsy4oOUfKIGeslvTC
zDeo9vRV/52YZjzmKpKXmhtifm+R60+Yjpx2Oy9V3jOcGD+fpmLsMYD7K9uNAH8SpN9aYmjSLpm6
oEJaq2H+B8hV5WVh73t/iAAvZ9MvPnhkqbBcDImFWXCs8mZC+jb7tZ/yy6VPRqIZ85hlg0NplCAs
ZEROyExu9ZHHq6S1CKnm566J8RTgJFGZcvsP7+MXVK7J3yBrPR0DkrqbOY5LvhFHU4jc2keXVqK8
0k0QS9Dl8SAZtlK7My4V/gS+eFVjVL3iPJ696ZNJYSFPa+4YhJH9ko14+NHa0rf64c99jsRQcNkt
/47BrELcV1iGxxDpLUe7FnxMhIQoQ87PknlPlJIzHfcXBMYqW9NPlGA5ysIunRRtxFYhS0iN/K//
9oDg2d7smxWO8qsNKX/9JqaSPGbkgqSDff3bVqjHJdFNeUnUoZ1RkxqIR2UUgjiK7W1f6gS+WDI6
1CgrJtcJqogPWB8d6A/CYvHynvRQgXjGXGsSZKj/TD3XG/CP/1N9u/Q8Yg8RyL5chk08/UaKrB7I
2wMBFkeugeONHyFAstPxGpxalsiADtemFDQG5xQhTi0jgggSYUHLAcr+sLQcnd1EfMpVoUbT3DcM
h91Y9Y6d3pXGyz62Qgrt/ocv8mpnQPUbXsjguMpG0uDgbeyIvhrnJL9ZMxCmBKH+HeUxXwZY4Dl1
OBdrqUVQOEaAeKiC/ra+Muhgbf6Pv3DlgYRNb3A0/5VS9r3una7lDs/sdIwAkYNxyJMvfs2yo2Cx
X2Fn4nXzW6K+L5fwgyeMNm+/4BWUUyrYx3E4UzIXA9oU2PtQwAu+e/bM2oTr0O10WA5hCrc3nPue
BbkODzaH4p/mtxSn2MGSLXrxupNvrUrcSomhvB4ucYlc5E/7XSV62TGvtHsyjpMA81TXz6zxhXEm
9UIYifAQnJf93l4D3cAh0ewRFPEHn7Yqr3cC+rieYr9Ow6m5PszhalBTIIzgsugoSKJLb9opS4ws
VrIinYItHe4LkCFbM8PoywgpZ6KD6VSnCRCW+9m1WiVns9/CslcliUWlrUCc9Ez4H8FGGdIA6Azi
2n1ZV/nu6OCPxntHp5AnC1ByQStmV/EW5RHON6OUDxrLmWlWFGSh8gzq9J/mgyEgeIvI6iOIMwtJ
BUO5OT2NoujXBCtx7rRwGHVbAhxMyv+nRaPRCUdgBGXWboQh7/iG7YT4FQFyYgfsgVre6nF4bWSE
REUf4brW0Np6Lbj7LVYPhoL+lv9NzkQHPamR9a2D+MuHI1M+zQccr+w7NgWOiseL72Nk+A64vpqX
5YcsAAzKUR+WdN+eeOenaBewoN1OjIpHQY+FMwFZkD87OG+mtWnFOgBhLvn8cCRuEhLfLKeKjDYh
r7u8ZIhNkpwo26RBKkAoG2d16wJeR5uc9ginF7cdweDZn/9VE6D5puQaNKkvHGbp8U8bVtAaTgXL
tPJRM3lpK/+PUZK8I+ScdFw0YL0RVcumluPoJPVnHPcyGW4kLvgLpeVWBEBXsUYD6EG92BvkHqgN
0kDami7jBhy2zVzfSeXYKZDvKJVG5SIy9VoS6TLSvJEDRx02+0HcjFP63y+jQg7tSZjOXSajTOoV
pJfYqN6ktY8hJkQ3XuVfBkkxsO+atyejNehIU2tBrfQ4X4uwjP/CQFWQuY53JvN9VuALpelGtdVM
I38ROOifEBZTt76Ewhqj/FO4q+XChmppjpy5m3/3b02XjK3a1rdOaIUhS+KrY4Bmief2/pnEl5y/
eKBz/wWKGxA1u4BxSpGe7sbkuzTlS0SYo1rdkMRx4fgRQNTsdWYQYrWrucLlC7oONwn+cpNDsfOf
QaimefUKoT0eifk7JkhqLKUc+eMx5QiV9xR/AiL0EYWqsl/dKM32OUP2ALT7ioezjLu0Pa3ZEIZg
umX0pFBwBeClzx+KhLFp3dNv+jkBPn/G98vSczj3WYZPkqs+VRk3paf0lYDGtNCdswBlIg3958CG
lWIDnSEG0WDkyBuAYK3l6+7O0weJXSMbKtnJ/LKtko1kDVMP+qo0zgBohu0pLC3tSF9Yw54Mll6f
f5+zma3z/qv1m4Z1UqrIripUeEQgOZPiGz91hX1lJH2OPtHCO+2W1U5F8vtHAop676tc8AHwZjeF
b6bnSrxc5ePkACVlHLnMhyel4zsCFxVXACBGG9i2sBqKrpSISOVqLx40G0ArcEeyiKJuEOGGMxQy
pWm3QvUSoLcJiMiOHkEfwvC0qOsW8U8HYE/+nbRjmoo3lJd3Cway8OphTiNrRpyZ9afiL2Ni8nXL
Q6Pze9Yq9YF+8+uRiOClQa4xsAlNkRbWHLM6w2UKz0gi3rEcIrzvcVHnKibA4sjaKuEB/ren+tFq
d4t2IfsqUkiBC2DixDxxzigiJLtSPfDXLltHDGfNVG6LvayFFw4Mtb9rL60ZDLqoQDosqRrjiQdK
e2Fq8oIeVKtOmQMwGsgO61wFMQ0S33Dcrm/olKexOCMEaGodPNiovtiQDip3JhKQ6liCxkykq+yI
HDVvz9G8XFX8vz0zEkUUY3ZUYikVtfBc8De+Z5pfq/63oy/PWGczXpxy5JiVycBJUAJH27ZeTw5N
oOQ1h0hlVI45mGUJlmQ2pVFxiqgUU4JF46ivASeKXBKSc1rOGSml3/85P1xoHyzFx5wy6jLMY9Vz
SIJzB0CC2OEb9sryidbrfTPL0+FQsA3i9U2pzqZXJHVGK+hJb1EcnCxqk43Gm3OxFBNXMCzHva4N
KxuWnZyk5NYfnc7pegWYt0hDam4S3Pf06kE9LtH3H7e6XmDxW1TpvCB0yH9mgtAPgBeARZBLqhpH
+mYkJ9QAnpe/PsefYtoARi/Wpfkb3TtcoiLQJxj8wJxSx3lxofih5uuuoZwHcXDNHZG2oz6iuy0X
hPNkjulKzkMmFgecMu8fYbwvmQKwEPN54LF7k+nuuvY2QqK20rE2rgZTgsuYtbEP4HaLwb+moCfA
92lvgtXLpG7zTCaaSBS+yHjd7VcWYGCNbMP1fPnQU93N5NgsXjMHuUAureQiWeFyvRlkZ8l8i2Le
ga+Uo5e2C8MWnLH0ngVfYlG5FPg89uV1fcgzuNBChmjlC8HaUiG4XKmNrwEbIiVPsZVQZ9h6rI4d
5k8eyUZFA6pIA20VQBaN3CzM0zwvgU9Qwy6ODH7XrbJMds+s2vP5NJI5Byej/lU+qjK2d8+8C4zZ
ti/oa1C6iL0NZL80EFI8Hnl987E5wpZSWKHE+rJJRWHKSUmMdFalHfv6Zpn0eqOKN2SoLyYkeQTA
RJ81hEF1KEqV3Ngfn5LlFuMu293pqJ84qBMT1c3jGjN5CW/yEhQCKY4o/jRY7kmxjpBN7RpnNfd+
17o4H9p/DnG+ZbrtACOvafgCURBkIMdkUGPAx+WbfioIp9UELpvPZGFZUMFf2tv5ht6infT++Fi7
Yjh8/FOeWP0VjfNahOmc8AxPTA/D9bIz4wrDfOBr343ID2WlDmKTjqjZlZxghhEYrAar2mBcG6R5
VV9mCWaAcueEFWCCwIqLCf5SUx62ZXbMJfdWiUIg7IruSNYxGfypvOB25YMx593FJJeun3DqYl1y
op+fmDqzcfleIAuBvl0a8JtVabeGQDuUfcg6eOZEPUi/Dxgli+vidO6TmxV+NZ12y1g+Jiq/NXLJ
9V0UbzVZYRrD4hG7GYrzhpNk88z/MvOp4/iqPYcoVY6yDty/XjpGmz3Y/9QDK3GjOO4PTK/sRCza
eTh1WQPS6gIU2NJ8TifP0mmrvFRp/8S3Sp2k/m2vrP+cDCqsxIXtOx2mHuqNNWkgalRVUhJwmZzs
qpouO7VRiGb7QfoXu9tab/P3lMUAvjyAPYR+kidnQh2mgR83D5c7LvX+jEiA00OPj9Rw4pya1IPL
BVyovP3MrUzCguTll2zcl0UfMIxS5SNFAf5BbevMokB8lcTwqvmDlwn9qsRStLhR7WLXlUd7gI6D
eCjy47Awacdo/TUTNnFlhpBXtvNFXAzVQZtrw4n2fuCZZDRn2dst9vNTtITHchDC+WvgLRePwbmW
s1u+wMg5+LCfGp7jDlTl9g5MbYEXxrC6MztCMeZ94CdIX3FcWALfCXtL0AY/PL4lSf+hkZt/7cHu
XriIBSGeRg9C69nD9/h00xoT8ES2dCO8daUwW20/oRBQVtyDXakvSJu6gcaYh45Xv+IrVN5/415x
WvRJ9E7MjPSZpS4C78Rie6BDB3NEEMbVaqsnvsFw94Hz8Kdfm6guoBGHikyZ83hioxLGlbeD5/9k
krhUC9vKVKRXFHHtNcJmUgfh+OFkT3TCi+l6VLHREWcN7N/0HljzxrXMIBiM2p58xW2wgYbJqwbc
ddkaSLK3Do91bUJokPMMhW9IXLMcI1nRbYMg8ArEkz1fcrOKXxB4viFHuJ8PgsRI9gkrYKL9mM9a
m2eqAro0fCPgJru99MIUI5Pe5VFiFW/2/s6wMw+/mZv36qcU5hXoeDLsIubIN87ZEnFhCQ7jUTDi
CnFUI0O9OxH+ecoRzJybkOh8RF4iqE4+G69OgsYUTLCThj+B9OPB9XNIckz6efC6HNMXIM5yp5p6
byTer6WBjG14LCbl3V2YrcYYCVsuzBBx30qJ0FAJrMx40syt330BDJEbt+CW2Sb+EIjH7jJCz7qu
ZZvQZ7QzPvnf1CDniRFIefKBFZgid1brS7ipmt/ApBs4fi+jJRyH2+fH474lkwKeSDral7yb/7+0
JPmCBlGkoh2z0csf0EG29WFxMJ3nOnXA9kxdEr+X5X5qms2cvuEtfSwfKw8DltQoHXRxAPcCQhLP
IQ58u135/huNEPkyOjGxCF5b9YYVmPMuDoTLRx5ilAQB9LEId1TXGS9UXsqF+2A7rxFPUcfVPr0B
t/QXnzUO7yBNevl1dBL+u0uV2X+e3pWpv6bUes50HkQ6QRjE3PSOPYhkWeoyEAqZhnKEQgxXJKla
Q5hbCoMrSkhJFU4r66Fwt28f8Ua/OYhHLEvuk7cKY+S0rolwljogt/vejHT7nQvn3BghT4O8nCX0
QHEYoi29vJczHsPhNHwama8Y3HOCi6xw6No0fUwRoRrPqBRKppl+rSkWR9tZhugC88925FrSN7gL
B/2ypmIa0tBhGOP0qGkt4nDvKtlN8eLRFHFk7dniVY551qc7RCHqgaXt7V88e+6Q2/j+aRpE7tB+
e8CTYbHyuEOwufdmQhjS8c/MQiOYtTsNFZdldp02Mv96snS14pHl5eczvKuXcT15RxFjfay55/r/
jhnpMTCLJVVewZ3fh2kZN0/cy4Vel/tAfFOjQDQCFfykIV3PT+xz97KqSUq6GQYZ9JusXnyn53Fq
7EVZgPw6lrlCKyGCJ2MB2qog9yzeYWaw7n1L82csSgb+gDGn/yeP4iXQeak2kWk2ynILT2VgNxRU
8hGsBOi3Rr8aMdNqyP6vNwi0OFRxdiz0WvpavuevxJgMj8bb+MbXk075OrKK5qjU7JamBOrO0ZQb
0qUx7CcHEEWYcOZ6TpRH/mZIvvnH90VJj0Det78r1UsmI6AvQe9ixlyZIWwdzMYvn3DYnLnvl0Ks
VbV3p9LHZvJmttP7Qm6Zac2a0PaDTr2ut/DSjE42fnEKsb8KSDxF0nph1FktOjBbiwAc+RCWkc25
ccgwbMZETEeWCmRWSwnnSJWl6I9WAMObqfKjDMmaGNP/EiujibjMlMFuVasBTb1qu7XDJw1/6QQv
41Ij/WehJOGqqZIXBOtL4chCSG3Ae4xlw6scaWz/1gHkWd+9s9MduPIEai4TKh2zdp2iTWo2aeoH
u5z5MS5J66Fuh5qlh3CkWaEsoSRu/OXQy/WJv/3viWSPux0OdKvHVz2Y7NqMzejzVT8lwvM4xrKP
FZV3WoOaQLrVCkL9dtHktQhMCiCMEGBypFTCCOD7hvWAIpY9Dik9yspJhucDRB4Vmjn2pDidiI7O
YZGT0l4a87FqD/FRDDWsGeA9DyAmU0PyBjpdp/GoiXGt0aBRULjjGO7h9eg9PtrYtjbcG7KihItE
AcD4lCfpXM49y7XgOH53zui8A7f/W37LphprFPHpPTRGofTLVpGeEOwP7AX7YSjd8ZZccE9a3Lly
57yWn81DF8ATiBxV7C6eoTzEe87d9XG1+B5jeWR1j9XlkjBLkEDJZuyCNNOObHN+NF9RgmDLsIc3
crJiOwS7STXm5U7mCI8vdrzSaG4mbm/fzM/b9Jo+rAbnJ3Dy6EXTyGlUdHf6Fazgs/NLJgpxCMlb
exBG2xGkcg6Ud5ENA2XE3rWvkXJGin3YnUNTcsn/Z8cFtMpaQha7Vqc4We/ugWDxYv0Hlb1qLpWw
541AFNU7agS0Wg0XtUNvwsVsnx0pPRsFgY+NJpt9I3Lo0ZEnDKW94fFRCyE4Z1UrulxM/hpb+nVs
jIdQFeUr7e+PTUCvl9LgEnVLgCWz22kk+Fy2WgdmnmXaSDYuKmF/ZSbcu4MJ+JWher7CDogdtTMq
G4K/6r78JixxhabRFJZR9aLBuI8ce8RtZlSFrYJcbnJqYOzLaBJRThjtlUBuWNbUk/EkWO9xpFA3
iXuHpbHiFa1PjPgad/bx0KgivvnxSUnoXZZgCwNIw635Bwk2B7ZL9YlfWSrMUHaNsBHq9oMFRGB3
rD/s5Xg+yhaLY8KwTGCwzvBJHl+/xT/RwZkTOlTKUJS7w8NYvUTT/LbqbdIL3xNgwART8KlHC2dr
hRkL0MB0IT/YxFPzeh57IfnKo1OamForABYLZlM5ECsvs3Du1kfKsbyPy+RpBKKdNFk8D7iJVWyU
easVKY/9RhiiYEEdVC+xs6Nn9OTl6dX3+tMuu5ThjUMJpWJhoNLWPGPNcFBcjrHqhjiU5NLBtd2N
887DjewinXHBQir9mXFuKiOSEW2WhNIcMDf/61bxnohZZR0FKw5Eg5+6zlVmN66Yj5yH2xTq5/BL
/9xXKO8d3o/arMtBRfjCwK1ibL6wKNUzlNEKduunTfu1oZ1Spf99edcX+7aJ75jtKF8LPi1GE3iB
i1c3j/lcuF+MH9NnHOj5sPXnHnRiLHSvEYvCgnytoFftW+prRL/w7r0tsQ+viw9rVMOvsc37754x
4KDnIE7s91EkzySbPBKwmAB36uhXkqNJt6c76SQYdSxGhP8Si6prTJILiYHcRz5NLsjgCBjt5UwY
4bAJdHni8p68xupCGBVCBJIXjg6TZlmvCHbpHmmMvzQG2e4vcLNF0Eks8uPbtpKJ91FtcOfXzlRA
mimWV8GLOCAYSA1QP1m8HSJkEYOQZWXKOau/t5GJtk6ELJ9gH6C2tkUeLMLxaA7o6+EL1V8bKzE/
hc1x1FexvulcWrs6yNhFoTYaEKkIlq243zrQGRCot1jXpt8RtLcxaCxbnbQomz0sCIMAiI1HHJXN
u4QJ0JfaWfM5tlj1Pt65NCLl1EhKapNHBCQ+mQDZ/JGx3K0xPLgSt/DbKw5NCfxsWHdZSnmyseLH
NLI2jIah1U9DacAHEK7xFovYlvEFsKOt7qeuxXKYZBxsRrcvx+S5ezuprRniSs0dX1+XKhi4MQtx
gVSIfaHVrbg8/gTVs63U5awXtyU4FcOQMm0eOmhg4dvhPaTgBjsdm0C7K8/3XdeCd/EBO5GIF2o5
7+2QsVqMgzakA3HNRs97QD5DExb3zOSz4PcyXY7/SW9BAU13V6iFCcwhlM+ZLnBnzjLVZAJuzIBG
Fye2S34lD8DXqkllO81iCo7TwHbH3BkuC35BJibsEh5OQaFFD2xvuS4jiD9LYdzj18lpZo5NMEv+
drN7+DcJINrnWhJj/WnTXGJri1OEhJXdiTYQHLB+yIIvVhEG4MQJqueYv/wTvs9/Qfvhv/WgcutM
HJUGjqlDiC9LbXWfrXvwbbajzULNGN4Bpl5XpMoZmjiy+pO8XsZaf8evwSRrByarQsMjbwoTKUyx
kyCXQWkgRFlIAU9FU42eLCG7N23v1tuvtFooZBi2i/C0ls67aVTHEkxKj7MMGb8LSxjzK6we0u18
3zdxLnmk8/r1s0Ry39ofre48LzvmjONjOCDN0SJNj8NbHutxyi8GnxyTpvd8GOCCCiiltRbcCDkY
zG/ZN6VAoHJSjra1ykrtzAdP/TxWLQnvHjiXY3OxcEb+U9R3z8k6j/qexHhPQXlQHyqZc4s3kjNu
Svyo1slzPJvlfkCLYJhMPeioGWKL3wOmQOhLwgaT8VBkQ2phdqkFUVP9svZvRITM5FSD7WmJPB+2
AzG8xwQtLE9EW9f9KIZpYBKCE/jmuTSfu9XIwB/nnDvrPEQwlO6+88GEKKuqgTODkXVBhvUdgLZt
1wGThsuR+FBcVGQrYdgRF3vDtufXB686sPRI4+fKbhRJxAdVixis6fuboe/CVyctS2YyiD5TqB+j
g0aoX8i/sSPgAvvp6ZDPUT7AT7EOt/NSiFjVQ3rJ+OwbW32rYeow/xMUShL4FhwR17mKsyWCzeei
SVVnw8Qq/I9YI6aQRd105ajduaxrzEKX+r6u245Ua9MOyMQBGft1yqtTFXNQFnL51PGyD5BHZ+v6
M7e4EGrLVsL+VXbygbVxXA0bbHzdI6K/BA5T22EXMHzlAxIe1SlnSd+cGZFB7Gk+pIgcYm9QNj4v
sbJK/FXmeKxLxZqoMa3GxWqyBWM7OHHWMQA6OCtY4T/tTCrwf1KwROuL3iU1Ck1mOqDKJh0OK2JB
26qvJcZKTBHCNFcuGm8DlTZ2Gng5jOoLsn6xkdM+Fr4QK601/vC+x+HEg1SYPBLMBp/OXuKeqcMs
VWz1rWrmgkH+oWkBPsH4yIE5ic6Mz+wPvalJxIRB4z9WSX3oaqb10HmuH1JV/Fo0TEiIvFm7u6ZK
MZ0Cn4LrCcA4buuh+qQBYNUFgxfaCt4MWUrVBTL5TU+vrg06BZdLCm5+rOMBpR2WcsbSYW0QOEaW
vxiQF/8CUxLUYpUpu3Ca/WogZEwMfmLdtrHGohJadQL8sDCXL04/mAdgED+tH1ako416eDcK3/rO
Wl7TE0RRxUKdacDkIVT8H2Lb2kcY6MY9TZALgrih2tDilD3uskNKViJbe+Z1Z95hd1MoimZrZORk
Rvwq0NtiPy+O+uG2w/RjSXfbDmCsICNRF6ddfJnjkCsCb0hCT6agR04Lld7wKNvooLov6JT2UrSd
1aAtTey80FB+7fI56pr6KPMnohxeTqfh1czueX7jXZcUcriCYHHSM1ri2h5PEZfFhMwQpkuGFfHK
dfs+R20T0Racf+HJauYlguADcKGQiOVQte6i5KMRCOVjfeHysy9sOStmjYUbZlioKzrUEI30uzb/
DzaMnOXGlFZNv+LNGzJC4VL1K5M86k9dldJHkQ33O49JELT7wVrlPfKpIlpnBJZf4VIhyCqBVtcT
3dOgW/3Zfk4VU8ZsEIC6Unl2b3G/P9OylXCMaYC6om19LyanVYJlbQEvUAJ750mcptvohldyY39G
GMkVs8puoYLzwXPaDoXI02oJs1orFAZgNE02hUUBHKFLzvgW1OqlvimRZvfyjRA1zH+g0inFt2Ia
PySWNPcayzEWEjf0rNyL1xqhYhPqmc4KuZB+4J3GBx6oVLkPwUCaUWJwjAx2ji470kj1S5omuNby
MPIEm93u69ha7ImugDV0vXxBywrwgK1ZEw9HO/ABMhnG2ocdWfG7Oz/l/UFRnCNktoj1G+VKweFE
65uXjbYnn4ZNq+u7aDOFM8QbccfTR6p9ExN3qBKIn1IcU3BRRBpij/ACcaCdWE86EhiDjWA/MQU2
XrW/96GZaF3on0DFbANbZWzH6Z45jwKbP6trhYQdEALbRqYHih8Kol+W1uPKTO7I/6wsPE+MdWxj
hfx5jdd9BhJpovPHxm20HoIVyzMzBl/mA+zhSVjMOCBjYWyMZ28iftEiZnbXUqxgUUmO1CzJOyIG
0n/NpadKBieO4XJJ1p7cix/ZUlTUUvCtxghNMoQP3CcYTZmo/GSC8/VKAZ5ursiL5yXDPAETBJVp
PpY5ds7n6o0BQCu9fwi3GNTFEFgwP7QszzQh5THOFMCK9u/lOcXy1Iq6rpvsf6+9okuI/DTsvyRW
3WFT4u2cfgMWbTST0jDCy5gKA6fGJwTnCo0sfSAALz2T0SgcrcUn5WddIHBrmWhf6sGqb66Z2BUZ
ip271PnypWwaDeegQJTrH8k58Ro3kJjlu6ryw/stikXuHY45bTiCRP98As1aGVfKuBxgiFAfH81f
DcyaeAMs0HmMTmfUkKjEDS/2kkBP4lWGXxntv4T2iWvfNMHW5RM5Ivl+PPj5S+BEsBhTY0J2DzHf
hCw9AcFUuu3AM2CZdSJ5KZr5RYuBI/H67yNtnPta+1nLAkOhzRAXmeoeCTG/j7xC5TyMlW42MuHT
8c1aG0wFv/qDGQB4W3ofefTSdjgSGEUmOb9fO6MgfsnkWaNoQYHrWUTUPNS2Z40mNUYNCNzHDcyP
eRGq49qeQ/9ZPQK6w0hfMW2MS3SIF1DhAhUvUU95ah63ET1SEW7+vbMtIPJkTSLk9QtvgSgt/kl+
dWWzyNRify46psOkB/2GRlEoeCwUadeUr0zP458/kucnC8pBF/KAkib4dTDJnHb/6yszAXLcmyic
44z3rSR8lE8+xwPqJCnNa9ICC2k4AlMAXx1fsMGBSomTK40WLwVyDACNR4xeNFC+ECVOKkobe2tR
5fPZ2W4cUuneiLlnRXkjo1ucrsHfek85XMAwb2Hl04/UQnifpfIqtJwyrIGohl+dptmOfIaf8Vzw
mwpmv2QP0uObw6I8L1/OmUXFkM7tDZKJMXfCtJGN2bbHVc0XFopinI9D98X/rWCBUuILoE5/BRph
g2GUjn878LIuTayLlhVCWd3/V0loP/Stqcr3Ix3n6lyxrXcETppD+vK00bxCL9lW4DBbfcXz7xF8
J9fPTLr5fXq170a/4r47FPAHBBJ+U7xevhmH1RWtdQQF7R6XvK8+N8vkuRDovnYtEz7rZwqvXd0u
3eB7U6RFZvFxPrhKzY9bQzurz621o+z/uavt7NXYl3Wjl828s6DmoEKe2rAvRy7qdCSj01lgOtBV
KSvB5j3LQg4ZACU47Fq+2SAgj6fu2Gm3McmOXsleXURc99P5IfKzimR4aK2XQuVGuf4SKNG5/InO
ROx2uFEU3SrE3I1m33RFlSSSZY1/k2GOrze8RhtsAjhcZvbiOtwM/ShSE58GH330bTFX2yLNF+ds
N3SDOA6SUKxmjlYBXAlvnBbr1nYDibmmKvs6DDOaNFPkxWtwSgePv09iCQJxSeUFdQqkiUo7hJ1t
hg9jbKVKHgyi2E9kSOy9OM7MiB/xGxtfE0by4z7d0vP+xd0xQKomPIWnCqxYIpPuADzeWEVbhZ5C
oaOTGi13xxbTHuYPQKq/WwCzAb5NtQ/ioEjTXiKwGM3rvff9DQBBgfK/kMeXEuBuQEb7pOVBtSsN
x/UxT1dErxK4Ny9wMQicZsMw2hXhkrCd/px1/kXnLnnPEoVtwuH8lj9GBav3bz9XOmk7saSGD0nA
Wg/JzJW8hp1JVnbVvXVQZPoFtW/UamerpWlpHaM0zGnQrrzzdVkTIIars5zrBNas8PBIxvQ4iXFN
9ay6UmCeHWGR1p4hNHMt/oM0H0KZ7YARdjeivmneDSEJ/AwayFB6OeIo4UTb1q1BCvGy7/Ml90OK
f/q02kStSkM1qS5aWkgA0P4Xx5eh4pVLOgB+3qVWR5FGrpW1PZxUoWRek9hQWbFW/MUmrkkhOmao
Uw3yR56WvvbtxqpWkNS5qFA9Cgir2OYQDvO9+Aju9LLmxH2XPCGsp26g1KKehdE+oPfmZjMyysjv
YGoYJYpQXghA4pSfdryCGFQqe0omAMrXogvtMLVXsvnsJbyuASr538HUwXxXeONhEr9PE2nqoSOZ
ZmOM46165vV9Ndx8fhEyd+vKgk9lGrDALQbP7pLCyOeAri2EwFKrHS/ZNaiibKxgGH9UCcaNhMiI
qSEFpE/jR/R7XHHs7lp4wiaxahSDfw8fkU8jmyTOc2UIBiIdwOcTTm9TWYhLJQxdHs/LxKZ9ZpyU
+0Fd7Mo9ofWlEvdbuoH1sfWuVLQ+ZoQQRidLihTQvT49E/N2jdbcWC4rY0d5Xhc9eJ75uPnXrbJc
t4dIGzoBjT/i2HLjz/RTWGc7zmPTNMI7iTqSUKyESMaNG8RcUt+l3mrieNW4padCpStF+ce1/AZK
S0d/qwMEx5PEkbQZJb/gfIPpt2QcSPjnmolRzAjwaMUFi5RO5WqLl98WXhP0wWXKC2KeMLCLg4SD
8SuR86DAJXfNckBoQFzLdNblVg2NP1h7Uhv8BXP+X8Oz8lSoGhtPWKxwOuIKb7eWr3jDR1NHFMoW
SU0+g/MYuZXLZieG0FlPyMs0RGpa9DmPVXRmDO6QoPMqQL3pUmEwJch37rmax+gc1gp6Ih/vMfj8
NPS2yfF96XbkgI3KLNF01p03hBCx0z74S5RxrN4fLXzSv093CExyAvnRAj9tm0BFD/jea6RoxEKW
XXikQqQIlTyQTlJaGNv1g05zTMnrCPcULFt97rJCb67HhFl1xT9dqW/2SY/4UHYKb6Uw+/cp22ie
nK3+TGHZiXRiU6VDyG/beCKs2/buPZx8CkTC0kK00QwEX7EFHa+UIb/bh0ScVyN6AOiOlMEnXPPB
3EHuJzlgS2ZdivMtCyXm3vxxRB2UnC8nESvUqMDCufthsdKbdUqWwB67c1ThOpwpA2CVixKbnbcc
2Gp+YjPsve1OxccCRydc7j4lyDl/aWzxdsqDGfR2+28IurjhRJzvCibiJmulvzrPrElO9bGlaved
+OPngOuwrMPZH7+JLgR04MSn2ADbFTfv6CX+wpbqfHbmK8sYBp9y/JnNQNmy2QX0LlnQM0Q4vy1y
lAR0D5IuBWe4ihdwb/0Bxajqp7BWTzDfoPPs8PgXA1m0swsvRRJBME7LvIyToZ701ing3h7yC5HJ
4VCDCPmtB9STePZn3JIE1OCrhQ1BaUS950B660GI//jKcbyWByPEfpBTrM4ozRUl4EFGfFi0CiRr
jemjgdaY0scvJ+jSwKDCnzIxelihIsBBJbk8KQw2M66ELOEy4WkjP0Byk5bl9AN9ZU1DxeSn2dMO
ehT3h7jf8s51oXPfvfEb1wZ5tTE4Inu8vNWMgawseeoSTSY1pe+Ll9qa9pirZWoK7fmFkWgtlcqj
C/HJjrvWo1LauyRD2lnIQDBUyC/lswluENJ5BH7wImaNpE0pe3xDSNZZvwq6xagDOXGQh5WJGbnb
2g/xcQMpYc7HNSpZtR+O1K3tXS5lfuiG5CCnE0GswRJZ5Oh+Ovgvyiei86i+Chp3c8oPgBFnoXC+
N0HSXSZIOYctkr0cA+FEkE9x26OfGSnfDCmoEly6FeARiIJhyOsfAHn5A1CCKII5o4b7zciblyi1
FxJLQKBoBV5Wd3/64qG2AFFQaxlYnjpVXSQKXc2lGeokHRv4lOTL7+GeiUVV90LWZAaGpWOkMYW1
tUSyUTMnN2+FbN/Q7yVC2+HKzk8UAjHFZqhD1UxkedjHr1gr+u7ygCG96K9VNvX0szuNhFXQ9ba2
GIileIRWoNm3K/HG0RJIbhd4gVxsElxRSLNUIirheJE1voFfByeG9u2Hxs5xTM4pMsmEtmOHfuan
TVJJvmvs+wbcSYV9/HjyAdvaCqtQVXLxHVeYRRQV046qz1Wb3dOfhJ63pxiWUnyqaOGE4rrcqgfE
etNHpH549Fi5dGBLmr8AmHg7xO/4tB6p1LUnDB50Fk2azzRoG01357naigYyv+9KVOlW12FgAVUF
PoKrP76a7rlq40UnDoOYAFzj66sSfrOzJPG2qrkea7neQdbWvt5Ni+JV8Gry9UrfspEeMGUpN+zA
DQSJf6j/xrG1tQT5MTVgfzOkEPuJAY3YvqA4NQxL/qvVhcBbhk2HlL/Ed/kY30tg05Q2juROysea
0CaaeOaxM3WZS2dN9ZMQg7jVnChjPoVMDikf5kL8yYmOp60p+irS3c6NzYKG1TRa+PADPwzW0xri
lwNy5Pq5CO5NpHd/a6klK1dkk64KvJSvFEgInuJQp4rtMDGXm5jw2uVOCEplOKd8jvqkP7m8TF2X
kw6VO0Y0MWkw5EC2o2qJnMm7GYYCfo/6DvkPXk8aoL4dSeE7RVTjz+RUob11mn+K8P1yOc5lM6ts
XfYjYMHNY6hksBN4NzTf7b8I1KIf21kuEzJVZJxrL4iuHoxEuX6Rc3mcJhiaXOzd9KWCase2GvE9
e8EAzP8YiP6PEaZXMTZ3JvzZW+jvFYOW6WhJaP2GLBTzXLXSw8TwAQxTKd3QfrSbbIAv+210mVb5
IpJN5Ut4bnKXH3igJPtUd6en66NMqGfwrzsGoIwikPY314lq65fc4RrWDkVggcPNxLw4FYKbetaP
K3vTn60/6OrP/T8GS//Si/haPzg9pHT6g84s9vcro24N/h7tUwi65h/vzQ2VKx+zwAF36PjqhWY2
pl1+OceLuoBL8kBo5LvbJWlSB80oVrxqQVmFq6D35n1EjQOwth95vSFDguk3GDlI0fxYY8zgfFTe
4Dt0OqbwKYWxEXnOfwpQQk7Eev+2X8wXuKE7YiRu7nfvNtJkinYYRtm7xLCrIkHy0qPF37LOxdlA
eD/TmhssYkaad6D0onW0wahqtqXuJuqjueZCHrtr0DWDc7bOePzNZLfUoMjioDpGslLZSZVOyp6t
NsdLVASsZQvn8b1dVmuW+lLOrUQgA8e8iNKSx/lhQzDxh/Uv/Tnj1CbqyPvaMwdNUsdzPQrSqQon
rgT6U2j3eOZG1azRQJJ2E0StA6lqSGgxvbDlJtDkAm5tmv9QthOMelOHZB1IPuNWU2IJJgtfhiI8
xCLT8UKFSLoqguZQWZF+j2k8qCzs76Q6yNnfdApLDZoBJqxBdd06m84wAsXfj4GLYryLrHlLvDfp
LtwG0OCXFiJTGl1LJAT4c8v3oes5S1PV7b6wocXK94x9dQJLSwK2ohh0dnRvD1GyVEOigHLH0b6i
LGfJTKpMfC/uZeSprZH4P8KwX1HjGbhPkI2sLRbnXPdE4MfcUqEas/TBuzhU9GmQ6Eg2IdtZFz07
o25WoyODSOAbpqCCZ1c0asgzeIkUPbU7aCo/RSD7kE0P742fLXqA1XhfEi1QBenA9YOkUaox6VpD
M2oQmWl7bkLGW1WEdyt16GR7/Vx0ei3w4lxCKPc3OruL6LuONZwCVfJ6idU73vZRJ/JvMRFiW9wU
++GE011/dt4oerGr+ZRwUYCTpR8cnRy88q5RNqaQVujC21yw5+Z4kEQHWapTI4EkeL/mxIS77bgM
JFtoxTZDIjDCdf/UE7J3q6d6y2kPs/vvyYVV2kResuVQxiZABasbSSe2u8bf8FDNLKXom6Svcsnh
2OW3PDOcUw2bVgISdor2FUY+H9bGW4zQyMIiJksRZ/lhJ34hi7yzTMPHgmAiEkyiaqc2jjvnjbMu
ksXaczY1Yh6SfCFJX6DIKvdXDprldUwutLyLSwWYd8nAO59hJdQBilbWrRfvtNrFlsyCkX8ocwtg
HqbqUyyFafdiQ35Ex12CVQwBrw45lRUHg9v1cuHoC2wi8Aqz+Lz6U3UqqvcBqRfx9AkLTpexRcup
BAR6L0+Ky452LbOp8CLfxZDNkHHPLeuZqee5ZguFo6I5gsT7D7zAQ66Fj9aJOTi51Oarp6zc9ELZ
1qFbEgxd5dW1Bf6pG+6s34FX7hWUyj9RphTQSUGywU4F7loh3W/6v75g8o90V4QWi+VxTgnIB/4w
l+E8E3avCE3IOVWIoNhTWTTpye6oQgRbrCZndl+OuQIzWVvgdea73qjeKI4mVN8HqXWqmULYT4oA
ft6C6toI7RGbxldWkNu3BOUX7QP0Hs5EgFWoIGiULc0hIgNwnkKQiVvGM5g440CmBVLhIPein6m4
ngUm1to1r9Vm9lkOtO7D2SzHNqfV6gF5lbNA+XAIiX+NXLQ676euOH84pKLBxWusu/HqA3YM7ZAs
+/Q1KqIVau/bRGDI7TxdfPHE4aHRSpE2fWhyAmqlzD5eYnTx4yR+WqijMNBpUpdXyGejcMe1pc9H
0zBfr2egJmat6g7e3EFi0Jdi8q+MJ2DkUx7H6nvwXUBGyuVHpiMAxKwj4ZX1LjrxOWULcO9RTn3+
EAAmHRgAMYIZ5GjuU7QnKJ+idfjvRYcfGbkaL5LfuNKGCibWqYQ4ku16lKSzAEcALY9xcU/wmfCp
Hhtv2Kz5JiwZUThskcfyPhPYjh0CB9rzLyoA3BpVcqRGA68vBKyI0pWVLcXToiTySrlqTpXE4hJY
eYZb9ACD0WjGQiPZ8+kN8i+FzOwF1JhknPJ4IRuD8ImoZiblCDtTZYdLS7fwpP+FJoUo3EI1KBqh
we9uqhuNbv+ZJ5854R73KfDUBTglbMbtbvtB/AmgJpI9CwT6+VklAtu7vbx6q+tiCcjk2oU6sDYr
DbKi6kPPRL5cTPX6ExZ6z0aXgtRZ4Xfgv1l5TfMIooQ+QN+7IdtCiUy7wFUmacDkXSZd3X69xq/h
20YbU2w5mZTS3FXy8rewjaq+8GaS5lmjBENsYjYFU/4xcBdj223aweAPmojHs3qNE5CR/cXbM3v+
WM03Hsp9euMWlTrdyoCKPd2OmNqkq9hy0yytSiSz5+Jcq704Ea4wIHDF/cSRAZ6OmZM3Oqj7HmFm
W7hlxI4gREd7b+Z/SL8aE++iR0M/LwhI1ir9hbcDAj3cOVl5DXLOc9qvmRgUOpDA3KVcmh1pYLQ/
iVdZYvZw79PQqoz3R0qihoVVMWHJYfZrwQk3gVRN42YNrIhaNxcvaB44RuS4N5n9hG14oEEe4Lc5
R3+kUScR8g4hRxm4SBswQVNcCoPCIcdCB7eno5oUipDaWeThFVeLHVAPcaQGZEYLIsFSbW8XHasv
ZYLT5mJWeU5ZB5hTZf48/Kx+U1yn+K2lZbFBEFMwK2qQew+ouRlZOS8hjvRIs1iaNlqWI5xAltHS
5zDelivVjweEt48rKs39hs5q7OhqSukT6rh0omf7XV3jD/+IqrvvM/+doiNDYKmZjJ/0xcW7S46G
gtXNN9VhXax1DmYREJ13QSR4SuRgk/U/33GPiqF6KM9kCu0kIU7YliklygGH6LtjBjUE/i7eGM6/
9iwDXFZEOyk38iS/BwktTxg07fzyysxji5hfQ6KetSo7qlggB9L1509yt3a7dnyycMTZ5MDXv8dH
cJQ+461G2zM5o7r4qFBT373woXpUX0IYNeQDizIqAsNk0Pugu+kXFbdZOOnqyFhiHgI+OBIzAYn7
ykWhHAhtKMyVlLHF0URQcAU4RpAlC6X5UbiX+/J5OGzzubBVTcns5p+XvATHOK2Jb3LdGq4qVcU6
49LHnMa8eanJFrOraKkUuinzYjycUWE8Xm8EsLeINpMeN1KA57672+gyeodzZ287/mkkiHMNOEHM
8lPu9TmW111YcogTel35uBVN+FTDGxQVZZz324Jq3thHpbTtAtyltzM0lsgs1TleQ66YuLaEMwSM
sohj7o3ZnCfqFQwyZ8NLI7L4D8JnboaB7hLmQDF7XnUG96gewMGPxbYp6nE6W54h9IkP+VvEVKGY
eOnnadV0vKeNkZJrrtGG3JaE4COArVji1i0URYnsetrjAj5SQG4sriW9Uz/dCg96/2/cq3UxUyTK
foQAZqE2/HhEoYWKDLu744HOmvBQJvkV62Bxsu8LXKilMgzLFGVqUPllfcvQtw8+D29E/DBhBY5o
uueH6LPrcbC82dOiabDWXagKvPbgIMwTLtoltZzjAXeEMD+lGW2l78OeTu6/V22JsEzrbfLrxGzZ
xNy+/59PWz6SoZyU8PDk5tKobPzLYBmIRGlX+d2/yhdgVsekrj6vOK4hVLEkvpW7ztnmTfCt7nke
rAuiHDuY9sBqa9Oq8tDwkdrItm5d9Gg4m76T2tSSWzZd3GwFY59jgUytmEJfSKdsPGOMDXL1EuKm
Qf2Aav7JRX2KSL2hpDikZCcNBdrVZu9rJsA0YkVAAM2jUMJawu/r/dwnm+E8Agr6Ik1uYKTKXWqk
1W4nFJAjpWVb1/sCEHmi0WaLvD1TpabepZmzfoEKKp5ib/J0jcypCxm/mp1VOXJWIkYEtljnrH1r
0rd7g+GvHZ1PO0EVgANmVK6tG8jCj6L0gZlD5iSBbh5bKZy4LBWklluYShG3mJMCwplAkeNgSGST
5d6s03gqLQAuD68vL/CN+8IMC2CYW5FJ8HYLpA/CPipwibaRjS/Dr33J1yG6+ufanCZ91udAZNil
di0mCN1duxXajcV8M5EgYyd9ln9IdOBmxoLEDnK+CPS96b2zoXSUTfQx6avKtyE3+B89aszz3FXk
9EJTr+ZGN7PmE8+Jhi4sPQALAx6zUNQQj44cZAYaO94yST9LJWaHIPggl3WL2CI2sZE5CHWROr6c
hGd9BrWb+e+c/39kF4CrRjTQxqhWug5QErpARAE4P+U2G4uj7DS3rDX5NvDeoxtf7tYaeONZpwCo
8I8mAhhjIXu4rcWc7uU0eocFSjnpn4UeJ6gHdU6R4JLOVQCrrYBx6VqzJ0Io26Hgo2Xr3V1a1rCg
rpbDoO//AiRDGi6A8+cgddz4Ot2n75RQJpH4/nNT3EQttbWiHsMWt1VDltCmiAkHIaHIMhmFRuv+
ZS2BBHnfURUMuH0yFo39a8vH4/YMzoCHlLaVCOIXqA8ZB0oFUxfWNVTumg0S/SNgy9yHBl9hycoK
+kOCcCzAj38QaUezvP6O7H7LcErLeJ4cGxqrAFOcpVlqPRmnzOx0YwrhPr5XOK7JcBaRdFEEuJhy
xHS0vZCNfZgg5vk39g29YqkKZBGrLVkhYNWvP8u84LEvwvAsrHPaToYndC1pJBF9Ea7VWM6PxdYu
71nk4nJuWsh72+sMw4MKftXMVzx9n4H0qfYy40dgo7vZb4Y96XyvvRZrz/UGI7JH7aeXNcSjFLFJ
KSDIXcmaIfyWxZ1O2ssrqFva2JWEsT9J7CVw4OegVuQUUvbKxL37J/sEWiT8sBtwoycqpe7jhK7B
dkF+AMU/xmJ5jDKbvXOoHoRKc2CytBm1HrxWk+kTgxdmkRXCgZ5k9bCuxlmI21EDHf0YcmY/zQNQ
zZcNtLcrpOqAHNjPx5XyM2nEomk3V1Q6/eJYYuZ1SxRxR5bN7BlaWo+wvFHrXtl1b94WnJFbLjEG
dgGYeFpiPCWRF34LSxM5A9ZzaMEHmAX4dCzgTRw0kPqz67Y+KFbn2xhql0t0ld9K37SKxUrzu3nm
I9SIAupjcjhV3Ab5LwslOTcsSC9U/hGKakRTVeWOqALC4zkar6n8TF8/ucduGhqYJ7y5houg2Atx
RG+kiwdrQ4E2lIzVP98yxGUkMsfcsLsJdSrP3UYVgmKKYL4VKO9xiouKBTXxsahuM/sFaeHvoheE
alyM5M05skzsxQAgI2k2KUnx/ePZx2lUnHfzknrVHmYHi0xcwmjloe/Ox1euW08kDZWCrZBqQnxr
do+/4SCfEMew1v3Ie/hqyuyAM/xNwOv1BdeIWjmmoqtp6eud+PEF1jxRftN5naeyfx2EeRJ7dYp2
/BD6vatKa19XGNwPvs9B5flKCFDJumoObGsNaRd/iBN4C7PnWhtRP9CR5N6lEpDBRAaCF6Jb9DmP
n0m0N5ahkwDwmchGSkBhuzKzaJmupDQ7kL1H085n0fIOQfEka/tCK4aRbOlchP3bdiCL7iyjKizK
LKGSdZE94PHd0iwpx113P58ZgiSAZhVCiCRWWausJy9t6fP23yh0dq4hw+CwxA1ZhQRaCGp+++16
XXsE1JikxVmJUyDCxgUelqkJRWTbnmDkOJNBQmJSxSQsrYCFrHS4Tv3kSCAsMaoZ17YFBWOQmjxA
26sYOrhJZ2e/HPqukiylTWZI1xGzj8EyC24gi3keSRnXw/jPJhhqtacYibZfAjS+sXpdqwG4SMWY
ddSrORvtM+OizSYLjFZDpRXGZJTgRxKfjBUY1NTLzFscn0xdBi1CB7o3+Idblh4Ds3uCznvMtGeK
Q0RJxCTb5TluC5IzCOKf7gcwhNFixjrj9DnXJhbBGQ6I12DMMPd39SO0AvL+xXtGzj1dMuasMoMn
CsgMhEoWBY0nQS9C86wLfWAFJe/TwIpUiJlXBumGmvmn3IkYgoyM8EY5oJwXDpzb0s+AQU4QwfZ9
UrSy9/iEliqonrL0z6EQr/PKYrLJrkzrrdsMGrgt84LfHAgZZWdugrAYxaa05PYRIxKwetco8suA
9eRmAV6NjUGF59IBgk7kS+QX+c6ndP98tbjr6QWRzoXoqenkc7YiEzW2g85DiFjn/G0Cxjm/BaTe
qkV7M8/iTbWsOId+o8bc/LFSnyh3d9AJ+JAWS24Bt/zsxUMFLa3bXUwMEIThEWdwaZ3JBu7b2eDT
qpGxQnyxVDQGa8H5doG9pvjTbCwcu7eFoAmicCpFS2AxtG1Bbie3RL+VSXmeCgdV7CO7h6mHP5J7
VVtJzDInwKqAGbPgBkbZ95BzCOfruLmJ2bhYQp+pg8WuZWYGfN5RzyCbWKE3O4YUpaq4a9Y1MTUP
AThiuvOon3h3wMiVi4sVmX/qfcTd/KmVxx57EK5qR9mZdl224pHF9ofdMus0XOl/iqXnRGyYSmQf
bCbSC819/xew0OuZVSQp23ZlBQuduOY7caxTPIB7MtI8npI2u8enm5cCZ++I8jEC2uj9Lb986EZE
4h98yNgXMl6IiQSEToc4DP5fSh0LNqttoTNb+sQhxoWjLni05su7RXuot8ebQq2eYuwkp9aRqOKz
1sMlWZeBx17QY3twO1bJicFz8gyByafzcRc6Q8bTiOwkTPyddCdV/G8A2ZTrdtadW+RCTgZ+pGUB
2cdiSjS6UE/Kljp5+12//faqr+78wl+L7mTaVYcc1ht/fG2MG34y+ORrHdIQvQ48JiPJwltB8sCw
uAXyk2+BGEZz0l154KLO4JUe9yl92fc/LyhjZIgzkCnfF4udFfkCOw1O9RL/DFzCHIg/R22Kwj+T
i9w7okwPjIX7MQLS5rL1nMGJ9FHFgW15QkedBIGsTgcpWZ1IjHwSbQqg6MlyV7RqcUy0tZXrZzbS
LSX7ji/Dk7CYN6RI4g+2ntRxqXb6edCrVxwLkU0vu6TcA3JPz8VcRtv7TytC4stL7OIJenBjlmye
xdfZVkv+uq4RHpCQ5obvN2i9WZgSu48T3kmeUvt2Huaz1ESQ1sTQahwhAgMZQAS6HYbf2u7bcMmS
N09fA5cZ+Ei26SvVpo/fFhJ4J+A/eLpwgfmBTQQ3up0FHzUNCJzh7muwXHbt+m1PFZX7Ncwn/cSF
GtHC+TeKUCV1TrXkHwWVFiGbFxRVdMzn4/FCTsdSFcuEb96T6cSJJxxNItj08q6fy0smLoj4xVhA
JynbSVFQ2ELy4GiDR6hGUAT/moFZ8oiAesdrWvxwgVyRzdwXVpjD95+T9Kc8fhAZ1ZW8Vl2PYNTl
1WMOMGQzecM1Ufxz8Q5K8ur5vJJkj2wRpj9D/J1yAygE19FddFItPicYOYq/obNThojoNM219rWs
tD6Bzs6yjLvzsoBtjnvrRSDI0zZCoWVyhI79K6SkcaSH4vv8xzOHiLm27AJwZaJde+v+FSWyNZjw
y6IofxO2XV6kiW2Sk0sWcKslvaAzdhUnt9RF+/G6PJ+s8oR9AByE8DIkOqbHmaW6+5hRGwBpSp04
X94cPYYf2jYNi65Vj942aju+sCA0Xa7AKMb9nBbcH6mVbzUAkh8O4TgHtCPVukmy6xbGzgTjEqrD
BYooEvSVUcPr7jAu+ws/joeDuGnniqcEphv8G2pbnozOETvjIj0HN/uQXDuffxDI67SjGRzn75xJ
6MLxLSt3GaaU7daCcB52jlD23/7YMNZf0aYkyHjyfXNMEblyXDG98Nzz97rfcqFWd++WNoeHvS/n
kQsIqPacQVNHiF/QabQEyS4DY80jesrtqmIOVi+ptQ4I+7C8XtWuCfI0HAMstlxU2FMKCMlkwDrd
Qb0o9INFEQ3gSS2rEr6DJpHrrKgIwIMrKpSAzKiYCVXcIx1+rqHiF7meY1zbX8afBrArTmcQRmCn
TGC9faIsO/3AJOncs58KVe49OXZBiuDSxp+5h4Z6ARFV8HOA0KOScdaOAoh8TlXlig0SrDW6PlTV
pBRAKF1lgqVx/iMCmlkpX/80d7voJUZSU8+hpbDkIwiBpP1AsEQVInetpB3gncvjlz6AixubOXjE
sVUIslCDq0XWrBfYp8Rd5wDOwq4LftRPFF4dF0EOxtL4K5knR3zQx46LHMPQvEIPuOq5HqN4cd1a
qQZe4tev2ld6qU4h5OYr7sElXIBI44Pth0jICcTshFpEHgvxgRG23Z8ZscLFBkvw0liEAaI96PUm
rfio3GH1YKCBeb2ItOfqLUBsnaYgPQJidcZrBcZizYWDDmPTLeC0Yad2plu2qvxyB5iMy4fmm4X0
viDvLebCaWjDZpEgd0HUOn6lQp+Fos9Rx5VtU0K8Q4s1VJROccN6jfE603aqgmULS9zy2h8chOl5
JHIxRLIz3tFKAaI9pxLeshYnRJweNrmiV1ct8u9jN1JKgt17ntoaZlEhwtNHfrqXRGiEGKdgu343
cLfWiF6Nq9y/3XEUw7R7wkxKcPbs5FUx+xTksa/jA5EM7ojovGlff4XvGpakT+NPHxtJwQWTjipd
R0s5oJFZXRyiAwsP7rPVUAl+6C/KjTkitS8FF4G7x7RlLXohTKyyQ8b/br1RwPwpcCU6u8gW8Oqt
mH4+by/3n8rMkYOyDyuZHeUyLFu1HjrhBfqzYbJJrL2EeLe95PnGAtXoa4XTYh2pXQKFQ3A79jRE
G1wa9UV2OZ/YZxKye/33YUWPKxkhdpNzTB4KWDaXsHH7/NTUVSi+Sza5ZfSCo+hFHyZdKROEEeqZ
rlbUe+AUndnHtt9S2BJOlpmGrA4+P0zNTDc1pBFEoax6V4Xn8T8CN8Bv6BWiLwieSPCq9KVOAdDi
Q7ISC/YL5SoPkdv3RgtfsajaCxMgcqknJnGvnWkONjnA3sVEh9uoEpibbjRKX/8dz4bTSI0XIYZ9
bVyfp65VDDpF8KOpyLlrno0p9QwoovMGzR5r33L786k+aiX+ZXHtDmeqoo/ufgHu9K30+TV2yJ80
DLed2uxbcQsV4f9Z4ORZ488aCHoYnuu7EtGhxqzJraBTd+M5TR5qxAF09F3+khZuaeBuyuEucLVe
++ghYCF+x6PMcApp1U/JuyOlV19oVPsebGEC3uu5yyGtryP9Ccfepnm1fiwDR58bIeWJ7I7bLgRm
o4FquD17ywRDLNWov+n9DqmB5XzLVDooXyHHPJLE3zS0xUea3F8Y5gCG4kNwdcgK+jTwZmymkK2+
UWg0ifiFH2BIcInC3b3xfkKKHUzCL/64878kx0yUlrTDYj+xmSWAcGdOmkUY00K3qoPLP4ZuyPIz
DSiiwZ3fG/ta59YxF+j/Icn/9hjsyA4/NsOyOMjfG+KYsVSWnSRZpSWbfuO6POalIseMxTN73pLk
NDch3cajCUAFszoJ9muIbscwAr/zd7mkzlQO84m9B6qZ1J+oCfi89VGyQ41wxNNBNo08J2idTwr6
97ZNisBq43sFakKgLykSUvZ3i7NfZqpntbxQJd2YfPwHFKV00jpv5w3F61dbVlQbdyLW4Z7H6yKa
zvglZKXXcDX5RqVCOU3rS++gWT+FoVGfIjC+t1fvjVlH3dqB0kxahYvUtnMXz2+Gs7cGVLmSbJcV
5WO38UjFy6ZSaWFempwwjD/tnvhwvZWOx/g1KStZ1jKHLLI1la4+fh5UWz/NkCPS4d7phlZcUlhi
7ey7Lq7xL4RRxcUt5IFzUyHscyTYgWSLLtzxPhla9AGAegy52MB3DPInW76BWLNknBaKBdaTc0Hi
h3oJ6bkM8tI4e2+LgOoXlDNkCtqjKA6aYz6pDYyVx+u7h1XSF5VWv8WA4MjX4RaC9HN++T5Bjs0l
5PJmy5XXw4uBgk68x4O4JYzlRnqpKzlc7LPTo1umT5ovB6/+7I/kw3VNP7zSh2gPh1rhwizGe1m8
sQnxCveNqZGTM2Mm+sm7+XX1qovtmSHOQSpf64NT0q1VYPd68OhfYwTSNToKr1bhaor6BMGslV6Y
0dD+/NxejMxwrS6oME70KSQ7FRJg3PLfPwFusnA2Lbd3y+fEsFw+h4isq22Q7xtU7YHoWM3U1k9k
4jCGVeHRCbKUMKQ4yCxoc5PCSax78Q7j1aeLbodOiUs4sUxFB+nB7J8fEb2uSXK1MgGxf2n4lf6p
ej6mwzfDr0KmtbiQdnAsIGZXjRNKHuBa/+iyPwTDXcMg6WbYFngsC6vYqB1byuqhDnINIs8994uw
9kYjR3iWDoQboG1LcK8w8K8AQ0ycECPq2Nbjebg1KfdbMUoXgDZFXKn0/tM5HVA88obc4CUWBGEc
Z8c0VTSKTqAXMdKOrUvlKCf1bvuYrhyKrpYH5l8CsMP50JZbTgaT4xxEhl/TsI5BtzWxqIEdaYJh
i6FFwMkLZeSvsJBu52N+VKvGHWZ0GCukJ4U+5gUpSKwWD5qwQs6YH4ij1K0PLp8gsC6H9xASyrFi
DQcUujh+IV/DThbaUeOHYA0x4PH/e4UniLocfKtqicUezlDnXqRerLHOKqJYeda/Adjf1qqbgJZC
BUjuE0OpxvedgnvXmaHMbeqIAZV9ramtVBMQ2bAgmfwfaIPPnKYB0mkQtWsuL7oOW129Ylu52ePh
uSUnE3w3laAB1ehoXVAz6aPM0/fZpFehks0Rnm5tJF4blQrrkct10bbtLKEIMHt/dm0CbWBNa9ys
V2go7jk8uugXg8JopO3zEMZp4HxBs67poED3CAaHHcPZHyoixiweoaILFJwqCKQV5K/DtBHznBEa
lEFKh0LY6z7FhuVqxSJp019Y5B1gxrSJKrXhaSmnkOJpMebOoGJGIjJ4U2n97DmXbXLerVTVf0bk
k+QNcn9qINIJWXxC4uu6M6h/TCtbcUR42AUqkB3xjk6vlNgj1WI392xTQHkQD+Fe9P9Atm/At/W8
IJlADjz1LKLAcgGV/ky5RkVuK54p0K5SZhjXSUPHH8YCp0HHgYK4QEx8st9c/+mYhrgVDGlC/3N2
j+zi8YphvQZSRi1jg+Kd2/xv2ZKGyRwy5D+OKgYV54NmIWuJApJwxbXNhErQmHOkAqq5miw6fjyN
jXpAz8VKRz8NgdPEv2vxg4c4tT2pc+b8B9cskmVg4zkQdvH/NwsDACnXk6CBl8le4jWjjFEW2Y0v
SckIPGdmIjcC4tpiSZS20Q73lpamP7SAL7izcvU+SfA9J2vWzFhz+nawg31Ih09zEf2Gjb4PRGrZ
bouzmNjNNxkz8U9ayaD/MVQDmZg8fdatKPpBVHA4h3xGybWuo4uewGpApGuBuhasNo3r86BbfEhd
yegCceOd/U6+a/Fp40z6pHC4hbbdyQk63p3ckVV4fwHCaOxyqdt9ec+z2NHjcyxiX5jQGxLoJ7S/
fn1vzwMioj5lA1NnEr1h1UxERox02P5Jg4hrrLum2JTnXgAEkdA20IuLnkD3IYlUrBBBqQwxhdyv
QJHSogQUz3usBIDQb69sVUR9lYaMlHwJoEEKQE+2Ett3c/3SwzjAYsqbIZEx9b4aS9rxZJWaNvJp
ARuFjjdj4/4leZZctK6sJ2D0a3q89Uhn6cE+GffS32UPixPEHxgoVIVZMfynnyPi+ZZEJNh3ik03
FsL6k30Ew9U71HWqgR4YAa1X5aDCGbzAPg+Ty4mwp6nxQfyaB1VVMFC+MUm53I6g/f0kFbdlnShE
u+wkfXsywM6Sc1EC+BgaUu5lrBwZqCugWHorqoVe4OrHlDtcDzdLoYjB9ZVbfUxDx7VjNQoGeagH
QXBzg4/lfWkQnK98cbWo2BZp6p5ZGssCncCdcItJloPMMX8PsUmn1z8yUTfAxKdfo64FgZhRmUup
oNSwiPgNoli45cE+rblIqM5K3n7/gpe6uf5zJqta8MRN6mOtl9FK3QSDheOWGDAJTz61qVQ9QH3t
5MmtXWAp2vu2oikySKQ/vL7mGp0MtNmbyzUEo4DiIZjlB+DfR2s0LUG8/ZpkVwK6UJTkPSJEoAVl
mM2wa0pO2pwcte5bgzzYPjzTP7UToZ7YW/Cw0yWHk/AvivIyQViyWvz2V/r77/aUyRKQUJM0KJYF
HZYwYsymvveMTZFdRbjI/wlerHey42hCzq8lW4JYR4PKtNS0W0rkqWzB0TIt2fJRii+p678z0w7+
owQ8QSIvqxc70ViFiBhFZbAH1CUrhmdba3icxePuCDRRkqkFyVjryVY/Mw8tTlXR/SdpCNWiKW8c
VM8P7/J3rLFxbqdABuY2Y3yGsuqAqc4hDbhB/FGwyk2Vi1FtdcXiDPala7lz/D73l8UcP/agdkBv
UW67wOjXu/wKSno/r7b9uiLZMkynlWhMcNwIqJqPzvM8xqDCWecxirusH8kechzFIZyUwcLZfCws
JDk+1fjnKQR5yxKJmTAYwNuBoYR2MXZaTGnzbQtpvunzih440EN8YJcuCcZQoWZbOgteRqboRDHI
+byyXmzkLgs/yOL3XRpIZoIivX4JMnpFSU0bJcLylrfoIAtUuFrbRsR6j1wgkJvmM3gIuP67iBAM
DzNvWDKLVEy+6u9C2U8WfGvtpM81EegVaYJxN0mdGqrzeZK5sdUIj3sdyD4V9xiAPJLMmkIFYGv8
VmIfME/uKCrQ5pfGWQ4kamD/EkaGi/OT7SiuPWZWpoaqaiANXifjMpWuTTBz0weAtx5rYf30IQuv
VYg5f5gBhZYUfTZ/nUFPrr7QvjE9CCWbv5atv/kKxllIYyyioATbUQK1lHxYCD3CJVDD4CbSnuM6
PZoRP3PjjvF5xcACjWVpO98KWYrnG5DMtXG/Dcr21eg3/fhRjtjOJVu999Q8I0oO/YjonOUcZgeV
DvVnorYXmUNNmWc1xUHVuVwBC4DKuNsXyAA6c+V7ymy2UUZmpPPZuy/y5ysh1qDoIdQ0HccFX2+z
KdpMXVPFz4MeADaXODW2kiQW6DSKre0vlV+/R+FLutuHssb5Lf87+uUk44dj5rMoKqcZL0QHg2jv
LozIqT0Mjju0wfReSNh0pkjrQ8bbODxsZLid9HoDFxS7R7mWyC1Ue7OLwhILv13IAvuKUbAegjZD
vBNjYcMkR04qkLIGO8lJKZqjdXBoMMJ/OhThGZStcjDbjMvqtpveSTtj2RsVct4D+e9IQk3WRmM3
+Ose619J602Hdy3+SzEwBPTNakOehHkYNWZgmu8+uSDgjEFHGBEUAwbKCR4SGSggZChkgT1IGi5z
ZLObA4WqkmRv7M9ZjF8IYj3NQiY0pg25wYTir+Oviu03a/Wgu5Fkr6qWyy/f+fFZ0qeTe9rWKjJK
Ihjd0FS67wZ/A6cQ0chfjF1apAPfg1RwtEud8UuSiCKjiWhNZu7Mq1WfFd0EZExHjkuvb1dVeHKf
pb4M15YCW1swuxrOe3WNAPOGLOyt7eWzUN1nNFH5RXE45BVgIIFFo7HI0UoPZcoIfPtn0fFOjDG0
bgdX8PvC1uLr5xv5Ugl9u5dADwq0FeoSWHQ2BCJdH2+m1Vrkdle3I5DB2LWdkhsOdCrGUcYmq7RN
rRgkELf7QA4H3QtOMMagbbvwiKP/pQfx3gDatWpKLN7oiQdWgCRZ/3fCPPipUiiysSUMhWyR0dKm
A4EERWBWrbBMtuhTVe5xIc+JrHggGphmOG6IvaIIf/ZPX94FtMOOxBFVL/VojJQ18QcsGrngWr2p
gAqzL63x18LTA1TqwqH4aiBKRJw4RGl1lz+amX3mI28Jf2TCXV9DBasbcH5sg+PDjRpNSijHu+f4
njcO/BygqpDzrM6+wAkTqP4F+GCHMxyZ8YhEtxoxHmpSv6aS3KOThuJjmgjGtO2QaGG975XSEgJT
OLcoODKPxo5rBp7jrDxDoj9j4szPx+lQiTX2J3YOldGvkouqvzSP1KDyRTzObRh3mG2Ck3Tx9CNu
gHaF50M6olDuigp3STlt8vKqWNT4PG2slmLzPNEBilUB6pP/Zzuf2DA2mpSLmSRWLm0JirRW/7NA
iYBMdLpL+a4YtTCvf1yTVfzMW4TOwVr1QfxWCyOXmnF52vAiinIVyJQq6iBkVvzBisJAK2GKdS7I
qPFVSJc3zuWe0Qfw48eHaPlLAgXkzKUXxEW+as+mENfdn1FUFMon7EywwX+wkSdGQPsbbxl7XzDc
iRZh8MGfUIDu5RFGDyYFMbIXQwpnffMnDwkZjPrQMvrtYXw7Z6cYdy1wLz0FFjiH+HREotAFFVgq
g/zCVYIVcCHudgpGXzPSM1iOdDijc1i7rkpJRk+TBY5uMD6fUrX1AUz1bTDjA6Dx3RLD2Djag0jo
7mLzFBRj5D3+yvk4SNdRc8OV/EkN03kSc3RrPAyefl6BdIQ8EH1APx/I7lnw0hAr6D3iDLb2HQwc
EIODAOmkR8Ro3dBc4Jv8WSVXfNZaR/PJ2jqsoGYh868lWuYRkYCxn9i864sfk+h/51CZ3nAJCNVE
OLm3q8mWCz3g9WdZXMat6mLtcXclRKU92Ex4vazIeOmwf8Bs5G4uWaPRzAzClOxFwpFSS31wEIXI
uCoYWJx/2CKYWE5+wAUQ+Z60RzputFxicoQdVmIcMW5IRYm7M3EB1WLWknih91MIhK2IihcutYA5
UaPtEb1OA0fw4tyNupTrzyVPfDhHXBZPeDphCly+3E3+8Jm4DpffpUvyj9tQAa6GqIRI96o5ae/v
jd9k9MOIRnL/hpHFrsMp3Xe8ZZXxNssXQ/8FkzNZUfYXGzONvRU4e4w3PMLLO2USLYYSJoOgMd0q
DaCyMj3ddYuqxdinqIcWgF4oy5QY+xG9D6tq5OTEoQtcnGtNhVocQ/6TLHVE2MJ3XPj6MW7zP6RR
A6LiEBshGGRfTuDDALOlNuPxJuxcIPLJ78szg6Ro2p0UZSYrNZSUsXYvhqT0GMbr1IgQWYleATNL
2DGfcHZRiQ5zXUKqCmEelpbJKDEMo1awWLKndUqHAtpUtynXf/sUIUlTofWEJyfLe8NMnOaquBdq
s63WL7zhYnoOgbEliu+3TjyEo4WKHYd1LQooOcswRyTeXvFL7Ts9XSuXdvrxHGH8DUXUzhdloHeh
R9Zcl9GgzHIYDpNhoqRpwf46mra0Pq1hOSpKEetnW4Ti7bJSj30buTd+ZYL3g+3JVkL/we3b1bam
U7yguBE86WDYuoUZaHBNPQ6gYAmNsTt3FMT9O5zNC7tdiJU8mqIbi8lc9KNbW2lbG7MTcS7Qu8Iv
jwBLniWREWgm+FwbDv8G0olICeJO331LOvbzEEo2oXBRrlegn5jzwO+xhI5rutcc+regwvr8v9Py
JYlYi8mRoGZJn9y4X0dycsMr0oY4FSlUwCIblPyyX5+iT14DncpJLoMM9f9H6RJXQ9W50i554LkG
uu58Z5nAkUh/1HzA/fA1YTHcXP0udvSm5fywxa/tgxfaPNDTmbRpM6ubFWl2+cRbD5dsrDRh10mh
Yclx01IwbB5GtO6p/wXI6WQfCfrdF5hPl786wiaWioQkAAZV96r3eCxukHPbB9ivT8hCrEVdpDfG
RZY2Nbi2N40Elak4QzHFIJQIccgOcYuXz5YHqCpzF0wP0GlRKEa6TaR4wHfGILmgKD67dHKHgc3J
jILtb+AGw/5wmYPX4gar2ZK9fWtBJYRzVBZwiHvtbzUj/iCuan26bzwRaasU6h8d3h7C2MQ+SsS6
8Djls/sQfflLQxOCwGyepG+v9vypS70G74Bc/Cln7ymUfQCp6kNL9WZs3L5VAO4wUL8DiB8ezD+I
Gdq4ynj5uChf30sBcdBDkO1cB0iZ4V9/NVYGX+O+Vo4RHxkbsqCAiZl2h647qwFvw5sFs5S/dQZc
j5Is9wNmvKOktVZko5ri6kWpC1T56YB60OjkAmFAsAyb4y6NglwXtQitsqlSdGyjYb4887rdrvh6
midabOe3p1l8iKB4V2epK9+WeDa2GRXtYsjITZhSyvtgJIBeZzh8Z7vyLx/PG8Qa1amviG7Da+K4
bvblvYinILcTSajF/yGPxoi2ivPRlBOPc7uco29IGK0Yq8fqAEE2xAiFjD74y6JHXyeNXqavO9V3
fAX7HHEFqqoXzEhVse4L1JAif9Ts7Kl3KF0vJQEtgsU0fQZN2A/6ONITbmlJY5PI/JCuTBvhHdeg
Z/UX4Ovt7fGah1Nv024KeFzS1oyAhAP549SY0l+WeuxZIva48EhoWCHaQrdHRWSl45wSat4SFR1h
miTIoImqeQ2cmQPVvURyW3k1IU2/Dz0f1GBQ9de5ySa+bwYLQhlxxYCun1PljQp+awQ4xQgBnSc6
UqghloUVM8cqAFCV4Kygjq8xZzDveet419Uik6WjV0rUg+VsTBZJXPNT+us4SBK04Nhg1JQTYAJ1
gDXumAu+YrNvUl/TQW1umbeV6awzbx7pkF7NtIln94yQ5C3HHPWlits9uDdFf0SCIz8k1AGLYRFt
2LcDutsahLbRJI/acFg0zgl08MYU8SzIfrV+YJ9Ha1KB5SnFWl+nJJo8+d2xVm8NiW0r9HFyVpCk
sgru9CX5ZIHC8jf5tS86DetCgcwqL00zOTATEBPnJaO9QNROqdzBfC6iKhgK2hD5CH9mnv/QVCqe
hQd+IjmCej/GxJttlR9rquDhWH9xxBp7Mww7HzFbTaZMEMzLiGlV2nJRxTy4XjhyOk5UO4hBcOV3
4GqXcZX+L8W1Xw++1l+MHqhCeIRsVip74fvWCWxQ6P5r3GjPvfVaQur3I9i597dbjDHe0I0XVOuB
a7X6FqZ8qlkXHJVxNcMjr7PTpUjWk6DGT4ce3T9ZF/EL4BT2DGP1d2eeL5DVSnxE07rIiXG49Nv8
j84nsarg7oLohc4Z9DRyjn62aalFjcM5btIe3H3xNKjrskp+SvlhD0WSwTQrnBDBqosymfPC8mLQ
wbikDc4Z5kVTR5EOp8hGvu6NBcm1IXXf2yevUG+MY2pDD2WKaQf+vtLaHfwaf9bRdcL6tKiTElo5
CRCoTD/Ihed/aqyXtLj4F8cgOnSG6j1SQzh9jerIK2OFKUgfsjXjc8r7wsg1oRE1JBGwIfwSkMW4
RVuvwPJEB7EbAq07dIPBBoLKzqDKns3w51FsKm/fqpvSIMc5gE3KeOP8foRxDuBzIvDeIwlp8eQA
0jsW56/Q7X/p2M1yX9QKXTb6TDnW7Z0Kk+DmH0KRvWwRXCgX8NURShVfHv0NFs0vHYHprUwMRXRm
4dCasQmKwuK3Vj8bzfL4ZtYWODDdd4dRTewu0d5C9UqhkVzA4sELHltxSIYKFHCMJzMbTSBM13Yc
Qh6Qah8wQRY/aXtfQDyg9GpuGsgCVfyS20BJo/ozkiVNBcNsUiyodYCuKo9508UiCcfoLZej2AVL
PWzRkjCAMyOxqLtDWg2gA5T9JeLhmgs3ZY0+1Ykh5awLhfLEuouzdmClksI/cu1Fof4JjysazmdT
vZPishWfb9IKRZ0S+TVJYaLiliVoaC141D/RTgvtqrZ8lQIV4Hfvzy/mjKeDBkZLtvXtHv5qXzHD
rEcPuhC5renNXcIbFP7Tk9NND530hN0REoRH8dpcNJZjGvxDfVjj8Hi5U3NeWGE74rEbpeYhw7S9
eSX+T0JmZ/HsavF7qhj1H+xSxBBYYdc0fUErBzDxoqq8LddsCems1SSDOpPyoFRh6xkfJ/TfxzD8
ekNjwGehwEJWBKgSSr8BgSCZxyfT5sKktCGC6Au+AZ4JWpdyf3e1NW1oZVPkOX8fP9V79HbfEGbM
/RBv0g8LuyrB4TN6MAr78l2HBIR3hNz7Vuwm78g49tdnvAvly/STA+tDx4RPVPZSzt3867ACHSZt
RSqso1AODtOcliBJ6b1xaOBoRRXSj1C1UuqXQIEcUj2N06JAlwIcZ7dFWtqoWFIEyY6MA67I8iiG
g9Z9WxoWQriXR1lQRIqMD5QoOvY2Y09xJZg/5gD2gJ5cjG04kykMwl6X0bnxKVZGW0opHIO9kM8n
INrLoViQEeTouXDjlyUU36RDpL6aR3u9FLWgT+1OQ5g+u+vMmDBWXhTSMyWuQcc/9rZ8ahyT2SWj
u3LyXQO2IaogJME3gdVTORWWWtQQgbLexysup9YBPdIjlWiUwzJZEm0CWSdJ2jg0cy/RCL4pbEXv
gbxSIkyT3EqgLof1kFoYYK4esJmXNC885u5n8tCzr4n8Nz52lCyUZFFrjxJv1Rx9yzklSOlgu86D
+bP7dMQ9XGU+D9El7kn/dGmPs8Z2Tgm8poJCMVmKBJxg4PxBSil9q+t3p2qb4Yw9V9hD9XK8WJmH
b0D1HRuYaAKhhbs8cgNCmZsHkPYsCAukBlS1oJXFKdiz8EBZTGdHvi2UqooLdBU5qNzUcxbX540P
T77yR6R/xic/mZbB1I3DuIuctRb/PhPqtRuFi/lbWa5T7GQQlScugSGDkLGK8hjR+pvz3r5dC82o
/3QvaNJg2/rbXbUyk3J6GdxMW5Lr5x7epMairYXUCzWH2589WrFWKuHmtPAOcYBMOjIjPgd/Et+D
6i1J9HpPsJR6UqaEi+mDdD8hlV8P51qoQkhaTucnPMRD4S01sRlOLNOWKpfYGUQyaOo++0VbXT3L
BzC2CtSiXaE5AHDvQ/y2txYz2oYsdZJ50pR0TIKnjDu7KtHS+kaA7afa2CalLHz4ZqWZ0cqpjr+t
7A8vQVI1iQO90vHW02CCSNPlzvp/cUvPPZtU/De2djg1EmjQ/5bMdyVSPWGPnJzubjx2aFnjZ0oa
abKdsvYE61X2BNBPDTdDC1KsoGxYuMUqGB2PAvrk95TJMjSpVHu/Rt0pR7fI1OLbXhEWhy4qjGzD
jUGyfyt3cSPkF5ldpjksLmpVpXDoqactf2fDxkcCPylpqrrk4TvygaNQx0xqfeMC0WmSv0HezJuk
Yxu7Oy4963GHz7vKdmbHeMKRM53S4d0/uvv2LKHMrq7Md2zMRQaQf/CWxGGfGVgdPyBdPiHu15Me
v1PMsEFZsEBAYkCfhFP7CGnyIxnLbITvEzUUIXcLMkwAKm73GXPtom4fYYv7hhzpcVAkLioAuOuX
YqDHUl4SylxypLcVjrryqRdOF1g+RS2MYxW6H0SwXpEwCqCWX8szRbAFKFePEC6ceulxd+PLp+Ns
18+Idx3f8/v19cr7PJK8oAiX4bhMua5ogXCWVTZ8Z2SuuUHiOXdbWtKHhfldRHfCY5EdOBXQ53DF
VkEvXKfoVry2EJ/opaNdcMYAXmHF5TkQvdsE8u2AkikMEkR5Ld/IY/DdqC3xtJdwM7HdOlaZmdOU
yvOdtwmx5eTsFQfYcnA6ueJ0K/jPduhxPRCyE7BysRjfG7+KijCDwvILmKYifExnPHUM0M1//xOt
iM6wi6yH6d/EzPcsuXp4C+GoZu7/VOQV5gnr1n5ldW5dNUg8IC5COuMGWNuNk/gkd69yQlKfBnxY
oaZI5abWUmcIXv7QrfLzG2V8Pu/ynd4tB4CsDnxsJud4AhTz+0ELWQjnaRN8hpkGUrhgkvvoSwZh
K7BZ/V2Y5ZB2IdWyETVG/8/TuWyAB2QQBACH4i9XKUJQUy6Lt0TmP8aGg3qYDYX4B3Yoj6P9Q5C+
akWnNQeQX0y3W5mRkXJzU2CFSBC/hVgO23ZHWfYqUULq4G623CzpP1EtlS2I7vurcnxJ2QfO6naM
y1xyidV/aEO0SsKGN6CoRevjyAbqrerh2ha7LYpMczSpU+U7gZPsmM90kmFJTwR0wRXuA+dAGELC
LI5MBIXw+W3eL91ayc5C8ItVE3QDeNM/lx2gzivG2MA5e709qvB+g/+PbjDaGJ4F/uhLq9cq9BdD
PPF6LZ01s1v4UB/NXdIeMdtMdPU9L0x8SNmZnAQe9q1ZC+LCxUfJi2vvhZ6XCAbbh/AGpCi8/D1N
COKwFrxbZWkXbgov7WJrWh3r9eosOhQemg0cP19gC2AiRKKfSDQjpKxPoIAdIBL8J54VEHX2GlZn
+xnA3mDaWdGJ8BeGBFg24LYk+CmLouucGMSx2qWjl/vGgSovHErkPmPBNt7/sstrCkV0qEFw65k5
iBxiDOa2F5WN3Z1Mg4YOAxJZI6/kCWnYNKhlrr891jUWGAlf8zHKeaB8lOMubY/oI/cENwgQfHE6
jOcU+xtxDQln4uDL2H7Q4h8s0h1WJyqOZFZUqHSKv9Kq2+V51VIF/h6d+UEUmDxr7uuFpnb6CeaC
tYHXLWwtgUB5ox/8ko9Ja6SdxESHyqLLwZpl58z4RQ61SY++buYmGVEPe57Ez0AgRRlgHlQQIFRV
XVpM0wfbfZg10LcuopqszxHCI2O/JF0tVcuE2y8vTMnskDuU7NAFox/8MwnbWWhY03W5qSzfaxDv
+2C3gBk6sncgzdfPJnBJTMBO2Dg0ovsx1BooCFR4DY8aevQUgQI9eAAdGPvxKk8+Lr0FhmO2fBKq
Edj/FkOQ5iaHObU+OYdLalEITuXA5cXZXJViq3nXOv5HCoDZ0IqCOLf0wFDBJDbEJVq+te+8TA00
G2oTjKY8nRoU3LgQSHalA+qyNQ6uYkL7OUffH8K8U5WkStGN6aBauV1/MijWybg6PCJ2JlDTX9dM
EdTd+yS5VBi7kDQkZLImSvY/UellW3/8SHE6gO81RYYFMFojrcmVqVKWNvbPsaKt5cPf2icWJvtW
1v2uqnrsrXF/qJE+yR7d4ENX29NPLcPdoe32n2ugA8bR2UkKr+kJRSmaGQ+sHzsOfpyr3F/hJTAt
Z/13ycehFlVCaZX0RChzxr3TznC0u+wWGEAZoyb8LJlMvI6VzzvF7hccpmMOdpEMYT1vhBMC355k
6AmDIMtrULOxy7BISooRv1mzv5nvXyTLw+7xXjwoUHm1EPOQ9VOzSqNFJ+GJ3QfqTULMz65OzmNh
fCTCy/vxV/tDUxS+Gm01C/p+YM9ZTPebD/GctvV3r1jy0KDCfJ/O4SmpiQj30P6kOG06s0lK7FsK
9z3iyUm5sJF/8NEUvALI6kS33UMJ6ZpKL270LHElcFRmjgZT6uUlFg6IoCbdOWZ+81vD7Iu/sDDD
GUNEpW289BXC7BvXD6pwOyTR0JUKDu20y4gsjct0SbLe9aZ3jf9nclGztIHfYEehOaV+Xmk/2fbl
tPzcWpX+Cl6hyAv6yBWnq3LH1gpAD3ML0Zkqxz/vQD1ABQaHaXSwug31MQSHsaf65C+gWo1mw0j/
ojnhFhS6c94veDlc2dlJepJiz3h5KXBTIXnLqhrXc7nCOVcXj+zNYLBSiyEZY3+3AnKrbmXefwN0
2KtTSs6p7Ccf7GGVj68g5oLETX87JUR7/bMZIhk15/kzfS8VGUZ68ZqtFaiE25/XJFpTk9GFk2kc
ElKJQQMaWqPTXSAqIIPx5iTyzkxncXFe8cF+Evg2ZUWDjGIlV+quLfiH4jClHlLbB5rKqU6bP1Ei
HQlRQyECpa+dlAI9qw4l1PSGNpAPuB0KHp1aOb7Cinl65BN6zIuHVf/yhHj249B9lh2IDU9Q7nJ/
1AWR8zYJ9r369MpV92F7j1Mqw0FFJiSIKUwS+yxbwUwIRYyW/ITm2LLZIZHoJvCbNHAxKZW3GSr8
rGQtNJQx+Ir3lLpclCIaa41iR4lZQ+h2NVCHXexShSLM6dgxstQfp8LwshDx9augiJ85xoZIG/yL
jEVe2wMUIt/6z7l+Rl/pt1KJSMyzloJESeqOITpYtpucKkU14n7Xq/pz3X6E4KSWs1PFB/fj5Dvu
yb1j0AcuXnAxR4g65afQNkHBx1VlvvUf5XmAkh90xQ9I29oQx8EYRhPlIQ3vQrF2/Xvq4v9oTNVl
zIAPCGw9fcf1AlHjiHU2maOEErx6MLf1bdHKQZ6dGsn6nOlWbleDgDu9WpgJou7bTkdSqw4rwRL3
bkTAJlcraCgdXzud6hY/JjBoZVPhBcfqGuyFHZpU8fkCGkITo7CCMAQhcuc53wUoDhNn3EZbvgrN
5RKXBaiIWrL6u6PXpKh6Qs5FnJwM8WVvDgPt3rR0Zf8d0qgXx8+wGwv4rScX/iQnE9U2UMox5D7y
JM66F4+qARtTeEy36rIK8cSqmwRgvVVc4FmeKjKREO4SC5WJcQr6zdZqetb3hbd5HDcSUtIxFP4t
15MjMXsLT5SrmXEAhReYyJ65V8hC9yzKtwyMX5x0ssBfsUsISNkEVrkzvSH+y6Sg93CgNLgHgHJ6
DtrjvT6kPkRJeTGwnTa4fJeuFMUN0f42qmAnndtyn1G1BWOHaV1rs4gYxCC0nXX8juckehYd40NA
JQpkHZroofmETDebMn/DCedWvHXq+5JXYltKJ+RiUVkB/1I7y3a5JbbFPh72Kza75Q+/Rn3N6d2E
y6fCwRQ8bDscyeuhJTWnnXx74BpYJDiuUYCjBxfsNK2Eam/aRPJIi1bCB7m4H8WmfuOGLJdJ8x6+
HMVQizP+5ono7Kb0mpTF4B6be/TwLT9QptKnCrUyETKMkXoke0uwf02xZ/ITM4sWji8KMD2Bm+YA
KsCZMmQx0JjKD2B7gBENKB/sRBJOufSjpELXQiYZfCt+sEDDWCSzYIXmqGKNvTKIT17UBvr/SdoP
6ZvvXyqydCkMxFpEWf327gQVjzkvv/J1fnMdxnfrKF+dzvs/7T0r0Nx1LCQR7Y+AvygdWqkIhOcd
m2HrtFSmxGcY5a8PZjl+Kgy8rWGEb00+2SgsEaXL1Pu0O6q1NmGjHUZrrtmQwStDYdRRftzEWx7X
GPHEuWuHtTMa0Qlq0SaY/24OPiuP8QARNYPKmFX2AzBxttCkIWSioOQGLknryvqY2oc7KwPIFMOc
N8m9JIvKAwMncwoN+bj9+ZZvm/E16IkAChhSM4IwZY5rnOvek3XC05V4FHtR4L/zG3vYLin6S8wn
/qi0DusBK6D8HT4OQx6BHledN0wlwAMvAn4XWIMHRQ4ndm9bxBJc8HxwMwKzFuBFVWEGdsiKKxMG
ZlNaG7Hofk2Qu3Sd4dfZuY2Jh/AOY0VQBVHK4wrkXSP+Mz1IrhqnHRIlIVdQ/9MMALjZmacaPrfG
sN+UPzYTqM0HB36mOMzX0jC8ZmBg8baa6GNekjKgl9MzWerhc9rsbUnDROa8aExsiWji+DkDc9u/
RHGI74Fyps+30PG8rwCSWhUu84Lqiq9E+2X1jXFPa6QCS6CBlD5w5YwZZoSHhhz9elAuSlN01Jxp
Gs0gUMRouA371ilh8S5PabWzAqOk5CClD9KPvSwe+H25am8i29dh7KYJekBKaRYeVNFlWImdD9WX
SSDO7H4SkpPyka9w2R4e8q88fbpEtknt+k4CpFaFqI17GiC21aaot1q4u7jdpwx8wk60G7vAw6Y1
wIULqFgpdLmxa0fC3vDfKNVJLI/hQMkONbxGtLmxf7oKXVB30Oe096GBm2EB/AoYSDYvE+o/643T
iDcVeqtZeGVSEVGkHrDg+yRrcmcZhGg/JUEjz2eKTQKeUEuzbpxMRkoH8804O8s5evg8z/A2h33v
2nd7SjMihX4H2zQ8WdOcCSqd+zggwL6czSAVABjVUz703GVIsED2sCs8hzGhcBs1tofOhm0bzj1F
bt/gVC2gPqIY0M8KWRqabL3kfYHBumsyL9uqouwSFd0OmaFfPNxZxlXIqcKeLrcgogwLLb/kxOZm
CEIHMlvcVcBo/fzwQJ+FjjInfUcDIIDEAIOB+aWXl3YDjdhsJisj3kpOBkAnqqq3NQG0pSflrOXJ
ScXtSAHswjDoEuu0HFU5ORj02dwJgONL+zQozxMUP7CjUtttJeEyIHhen8FyeAQ94MucW307/qqG
vrCWu4XfOn0r1aIU9RqHl2Kzdi1j8mk4FnsrUbAtf89Y/+gCyTAEJ474ttQkPpaVbjuCHmigHNwB
MUCdGpl22WdY70tP7rSxJvlPBr4zo07/s5fIzCcdgoJdEvPR3vSQmSpFEOeCEZkqxtiWOP6mk4fY
WzlE1O7fBaFK5rshtWTuVx6cgyBj24Ns0cspVdzg5ghxNBKl7jwLP8B6G9iBiNZ7ytJx3mQdSfqt
3Ldzs0mDRBBZKPLE+mHahvDCFYIR5NSSvL2ZBOY0c6tPGaSaSSN6164dOO+scIToFpbCY08DvshC
o9D9NLkiUkQO2MQa4o3LqORskA9oEBFVzrFlA0bZyt4RI/o1IYbQ+L4LhZn2cGqCLzdB/yi4k2Y8
tGufDtefQQGGgLAjPzxm+3fxsG4PR2GtICh6R0Hui2fHkcN6/1P263ivBxJMFG7sV8DqSYSkSjXA
0/rWVh3diZR425n750qgncMeyg6tC9c6B+xM9bYpTM31BVG/lVEBcfYkbtl2AbmBiWKZN7I8iuvD
mOL45PWqw4ewTCwCUzDnTR3/3X3SJK1FLoHIfgZm0XA65wGEy/jA2UdF28llPPdUatIZGtjTCBaM
rM13z/hER7NIdZxeZ6PUzP02H9FI73Y8IlspgaD9BYH9vs0YOPL/RB7YCffN8x4KAvScFV7BoNec
vLgLcJvq1RXn5rRhohYi9HIZoY6mtzzXZA1lRZNO/mDg6hyjC4ppK5llYYyNgtTor8u4sCkZr/Ik
c/M1ve4+cmUTmPRH6EqnxlF5ozafH6cSQIt5dgxMa2yafgD2EOYKH5CMrnRPQYvDVO6Je2LkK4Fb
fhQWhHEZ3wQhf7TaRQ2SYsPCIdaErUX3DYgAkEsGBe2+UDcQsh2rDVJNAK4cqisAg7Vl98YRW6jL
Qr04EuDN/vW8qPubkuWiXECkEhHqgbRgmtJm5IOm2lRDE4CdFZ7YpJofGPJLKD4Am/No5SsxYml+
y5dpeAMpLFYYPH6knHDvIX2x1AIAVnb4/LhbqZyXf7arBgbtg9Kfa+SIqyLw228MgDMVA+NKmz9N
N+RXFLGA9V0fr7XM1x7jzKAoXCnOa82oU1CYVULuNACaYdO+DN+ftVa0r/icz1gzhbE3OI23F4m4
CjeChTc+BrWovQMmFmzxNMyr82mPlVmlovZ9U95o5KZjrsEGy12kz+mqLQypf61PQiNX3MUruWuP
okMnSLt85DSIrp0BWaiztj61wYLFafdEAEEoOA2Akor3iKIPdohBiW/kW7LEhpIEEzkKRzkD0Ad1
CeK+kNwRIrsRDTma1+QaJJ9APsRpq+FZwUu2eorsvUWGGbYL9bzatvVM21j+d70++y3iWuOGNFJ1
nf9JBAjr2EpDniANzlP3EgYxPm8qLNgjkxlSAHiGg2rBfmqpSjAJWzyqJnwtaRX5XaZxjLUMqqXg
ZTl3sn7gWy2jzEMWOejtJFup5amokKUGoECCabw6nOFFDTJYLM9GFX0bbynIHzbTr5NDwM6fNBqb
/QM0Q0Br5vHCnLfMkru8/wyBv6zi8vWpm2TmN4K3+dYG5HnF8+vXk9EufQ2iYGAUol7NcNgm+Byz
+W9zHP2lPzoI+xCgSLzOE8Xzoa0kO73UHrfsV2tIvG3rIZoouayOI+mE7+i29DVv9rWuAzOZkZ2H
Xf7lb7QpjgRHEtthYqbNlpg8CRsSIiZr9T7KYW1xZhgW5upd1+FnVJQ/UQxKkLPxW5gV8vb+mkfi
0XFJ9LqSuvowNcRILG7BID1TUJvNVmmDG9aXOIihd37PqTD9SPOtuPhD8dpx0NQLodPLijsTmqaZ
a3CFBDUzfHc3hbE3QuT35VoVZAFzBrHYhHs+v+vJGEGfXgQRl/odUKBMKRQ5MvOaQIQ58vyQdn2U
Vm0oTiMSnLvC6pNoNxd5l6XZPLeyuwhzXFX5ilQ/Fg1Xlvxc1fNPtYK06Z5Yw5oVDK85SVApWWRJ
f/kVvABWH/Pd2qCddD6rate1tkYoBSJAkInz4Ac0JinKVLSnEDl4Ac+0KvDyJnlEw30DMSHJ5f2r
bEU4/UrrvS2pZB8cdzxhtIpyAy0VGmcB0IvsGKPVgORMZyhBPbn+gKlMKDOBzfmV5wZ0XRRBBTHv
dggGcCDXpeNEGRcjMQ5c1rNjwdB+D0xSku5mP08QiH32GKoWnYwQQQNB+U8UwoWmdELUUJ4K05W+
BQJMer3pNOF9aaeFd+UbDU0zinqBGYCO/7VgeKPMtgQl7Gg6CszP3zUegGrBbVEOIKgmQrUGCJOs
fMAodaiCsTvvTVgW/pL4BLEQ4hjVAvZTPFFwy77a5ct2jeKZ6mlQ9eats73MqvJ4WGN5fpK7zj94
dZG4YmQluE+iFNnRXMp9sDH7fTPNk7SlZMPN3YVL17S1ka4prW/oR3FtXnbP+SRoRKZ8MFkHeLQT
wtGdS8fPasNaB6rh0h8gDxVc/iGS5FM+7/FHfT61SUdJ3Dzx7S8sgouDAC0bEB2IXpH6WNgBBycp
2vwv4VeqFZpHuVjWysg+8Mr7tJMlDwpjf/7lKtt961uC9KkfN8tyXjtX1oWIUNdn2uPxpN0blkR8
ha8Yqbr9CWm6Bbfbwm8TsUWZeqfP5BzVOnpgc/TN3ap9kokXylCqJyzWxDoLqsDTt2OOKBgGqZmG
m7KVjDiEnaRupwlarZn/1et2Kb8gjcWEVL0qVGnKKW4fB8Rnd7FF7GCg5Cd+6w87ui6ivma39OQS
Y6yGD0L6v775KIH5CqG8bMElRpABddgY97KTyqEXWkXOSVzC2WwoxVIbhMH6gc5P4nP7iiJ74gW1
6aOUR5I20Bm8ws4volVoF63qgAu6cGZvY3/zBSvUrcY2pyPgvSy6gysU+25kI5rR9tHA8VGZwQ4/
X5tpD8XBMG5AY76AbUoagLYPePZbbPJIZplPeieOjuDtlvAn0fV+75dzpzZ9vJx2LcYvSSD8oYx8
wa6lJ1Is6995INRG2d+MEdcsRfYUv7IJvXnw1/PX6j0FAo1X1F3aqXQpQcrBoOd89sQmULqCQ8Gt
HrrPZzXPQW0dOYqlw55q3FfZ9tWHMR+EgPTuzDdsTU83TxS6pD/El7+pOfXZE0M3VW2H5yrMum4t
yAEVJD3LcQVVicv+eAsHRbFpUa6VO1YTw9+TzKH+DUJXzUNuJPVhOvgcCnzhqryJu9KtjbolVvVR
6YBOmD649d2u0z5sAflLohKzfQqWsFt00EGjJZHFQ+kp6KiAdwj0MAodADUFk9t8nITk39ODqRby
ppd3SQHNxn5lsLb081QGA+xexYlmm6Q6jDT/7SlOCCw7nGDzz3yitXjtWNHnWkzGgwsMYRPJuAgo
M18pV1/rMv0vfWIMjyICXbI9XjtsONBMngnTjgiATLl0A3sahBsGYsDr8W+qkvccYLVRLWJ+w7GK
LNN/tenIBsfnoiwvNqxK2ukqCT8lW9f0+9qiuvQsaqfjLjBBQDXOIjx73jN0vdJFX+d/2bbUj9E/
9uPAN/vXdTJfFpxIqf7ixPMCt4XdgUFI86+ZPou8QG/uxhsaSnM1Zneog7EjQDvpbsymQnAySO3/
Jp0hjJWnu/jkCSxX4LausY34J+w2PL4GI0Ejuuew4ef0a1/2cgX5/wMp8ZKlGvOaIsklasfudZhm
rH9h+YihQAAbBE+NyNWGK2q6HOm2Sk4Srngk4Del5sb/VGAewJhWP/Zf6gtU714j2lmU9hni5bXi
7G17f5oqwdjQcES/YJQrzMfanl+bN8G7ov4k46rOokf3v2Qb+SuG3clZCvWzf3qGNemFcyQtq2wt
vykexaowRiILRpW8wnCRtoG/O9kkm75kt5bc2Q6HABVejueeKZj+H01g8uJQ3Ahxgd5XoR8QE72u
7w/8FkKkMgtJAAO9kEYhoL6y5HniOpNZWJHwK/HsesoNPcW2iDcaD7rQJbkKA9ibYql2nVRVAhRr
WZhJkHvQgDxvifno89UJ0K7GSBTw+EyO4eWFs54tSNTAK/5/Kq4PUdh9nlmDKmYBz6QYshLI/4Xp
7zsB1nviVy+RxVdK1P/i19HO/WA2AFY6qlXo2I3yoUBpt9+qWpmUOc1iVik7O4qVdePwtIWcHdXT
Kdn5TGZO72hbZu35E6B6rBNzXQ4KXwlNXt02ZSSnmomq82+dDYWOKRW0P92vNSMzuf7PIkypkypp
ACmwYFBUvrs8C1On1eT2fdLd7J6RTDMi4t8af0UHALgmhWbxRcd5S5D10Lg4cVsDUN/rWYxwIlcv
lGvijj1s1GZfMixTeoMS4p7LbQfiOKvYfTJrj6oVcyFgLbxB8AvggelfUPDZq5UqZ5wVGzJ0x6Bs
v5MnOi7XjnxzQTk9wFCAeZ6wYHRxr4gdRhFuCo+VTqJo+H9vnWxaHB4WfwO3wkFSTCu2nSXpoGAQ
s+6qiIFc0sxsghpJUp4BdACCo9etU8rzLQ+7QgGHLT9GFYqjSSBNRK/YnuL3Wkqv9QVeO+EUICdU
XOd0vH99V89oTcSk0dE0hhmCnBj5OlCKUbePHBGzXw8Xf7YbQ15x4A7I5ZCiJ+vWTmq7YeicKs3q
BGWLOCCmFqWGMH5qaVaeFGk+KK7/OGakh0LX+kjMOIczOPEz+nyg9AxDxIOMfoumv6dSP7Om6sk2
3vc23WwQ3IhVPbDp1TXUXqq4Bjrg0fGwnaaUWGbTdefKuIrfnd6ZdslyTGxl6hkYyzA30/4umEGs
EZjjRk0u6UsrMXKOgNJZy6aoyqjTXFskcccPAe+QwNPOPrYurYrUuhHsMcgMiupxzqRJrcY5Z4zM
m2xndl2ETESMqVQF0HrJbfwirsKVexxBABGyrTrjcJtm83pzu5WVnRMjLxaLA7K+NxAhAmWEesKo
tv8ad4J8TlO0krFGWoVDYeBpOC1j6MfDLgt1yCMvGg3CNKBBA3xBFTkXyv7Kr8UpdLwfRSI5JJn+
Py/73bRuNSq+5Q6i/2PpCbCGmIjcKoyQikBbi7jSLNGONgPWHL8CeHV0Aok2j1ptZzk6d1RkVTYJ
qcOgMkD13iJOl3axu7AY55xs6geFbKfEK52Gbdv0jaYULPbHt3tGZslTIxQ/JxgKT6GBOAakDSM9
bkeR3hdXto1w9bExAxJFrgONeUUUjHSjKxQe6GFZU1b4OXynbhAKkFghWCQOkv6LZQM72rn29B/Q
N59x8KH/Om3qg8fx1YtlVEO76CTUiwHdfSoRati0xk++4gAnSUWbeU9fzB+7klSXk4ByJKShiRh+
BjioKf8n02RXa6OQR4tLSG7ptw5k9DQuSYYH8W2lQgApiIxzD0iuuncB57iNp1uk2i2XTXbF2IaB
aPGsEtm+sBjclOFq7AKkpbhIAr0EH5wrbex6z3SZDANjtt6f17GEu0nuUdsJidLFur2nfj+4b9Cd
6rZt89SMCJWcQ9DJpfC/gwhpfseYACOH1nuBQKevAS17Ej+X6omLmnW8GhaGMmKA5Nxl6Y3UTMAI
Vmk+9kDjqAeeufidqgfWi9yHwS6Wk5olGlV0ZDBEyKrdeoLysYdpqN7r2stTvSNNPFF5/M6mVP1j
4L/PDWRtFvtAQeI3onBCLc75E9ytTWhaMYfSCF3RtUlfNvXF+Nsh0e4FgB1CWLixPLT9v1zfgMak
HuXM7vYGbw7gff37698m5wC2wou3znjdNjVgXGUignqZMNWxOK3aLKfX52yACW/0fFLOzGC2fWM/
ZnS1gEhTx7jo6w3JLq/NMJlXGtr5ZFoyV+TWZkl8uP5pC0deKHCFCVMRKYnO0Lf+5+Jxjz2lm0DU
urw9zglviS5A5ToYaEdP/mZIIDRUvGWrktYRYpywcpiR2Khdo/CJccvpuSP24J441TnPO2cBy/A7
WQCxMMl8xMs2zhQdcPZrjyAqKeoEGe6yJbbJVFKRdoJAALZ/K6N2qs8QJqG0FwyQJbm7FBDQOQjb
Du9k7KhBdko8X1bFINjNcMcmuv1YBmkHKrQhTWEpIl8nNK8NKUZ+PbqP/Dtkjvf4L3RMIv2Wsoag
BzoiZD5XvTNINd3j1rMtzRggO7HqnFCF6In3Op8pI3tHEM8j1fYxplNKxtrHwAWOiH5mBjPRb/LR
Nc52g06Ctg3DvPsnFxXx9dhM1P6PHOsH93gTqR1DoBKvmP3WNj2NBjPYa32885eE+NdPrLC7m3xJ
EmjHWCpuoYSGRkHWO/wH1ZUC89jo/VfyDN+uo6ea6TVucERnr74C+82HvBE/MhlT3qhmlVcXOD96
YW6l8qD77fLt+sRUSqZYuRcHvw34/oaRUoQ4VjCeXZoSRzslwE1FqWYZGptQ5M8aU6HphSUUN30S
paMRX2wWQN6/PPF+OW4qU8ZJQoVs96/sATVchbXuiffxs0h6tr4cozFoY31GVJo2BaJJRiHOXBpJ
gmCsG4PkX2OdsGSayCuVk2ar/uexv3r+NZl4MgjB2d3LQZ0jNfyrA3voPVoyE+IiB/NahyOZrA2c
ECTQPDh3EGnvIVXjdtcaZha4eYScISeGw6Eqtqsndb9vjUV4/RoOa1U7T+UpC5VyzAIsvswOIsfj
PV8BnU+YRNTlf/B6/d470sZGqk6AX23njqIrerKkaP2Akt27o7HbI5h02P/2UOEb9s+7UJ52xJAL
heNVsOBnCF3b3gX2OF1Ft9l3xNKcgDhjEG8PGuGqut5p9dg7q9kXKM3mfh1keHOS/IGQcGVJDFFx
JVzGJFCoklxytkTbdq4xwvqkijc414hHlNAop8tCY5xz/R/fug15db0tBhLq/FgfWbwcdvdqcwoh
+/oHqw5fmDlEIVFEYLKe5Wsz1I010q4skzL7qijfupeyWJqcM8Ng2PlKg7SQwmAWZE5FjyFOx2aB
wfoZd2y4XsmdFLcZgqTHHSF6CxRwM9vg7AcEDFR7ox6PxaftiMiXRsfZe/e/IO6UCUvd1Ds329n8
jTYnp8gIekug630UPAGAXl9f8gRJ0JsTB6ZwfC0xDMl4s2QBUgaBMuwk61tabTQELPVPNDHzgrDo
6rzq6C4XxBoAmKnWqo21BPFlyrs07kAA0Bx5AY70Eluoy+iL0JBRNgRbXZOsEWqW6g1rRa0nLO1p
bc15uJfFfBpGd/hz7iwX+1ohbX+YKXWqJBrBepio+iBunIxgvcvKBQCp02f99a2gehj69rSpm7+P
RlXPgNr60Xr0Eq97qflrMPuktKds1ui8SabWyR5sw4eDdx/D+EbMP2/Yg7RyhJ/31IfzPhtjOj6b
pW4EnBRp+AQWW0AWlCU5b32qY61pc2x/st5KZM6/4tX0TBpT+mdC/IyC7IshTSEBijvnWhAr+vJU
B7/25MdCShFR7cktuODAdJ75NCl+tElAwZrGkig/5l52h94xxinFkVjVn378nMyuYGgKjh9znE8G
jcgknGBwYCz1ZI7W0NC6B43l2dxhBJlOfmoZFI39dUAYsIr5sspGw7JA4bTrflvmE5qNe0TQqkIm
gM5Qxr3y4Yb5rgje0mP9ZafmLJI5qVMpoLemGe7vNt1AZjBXs371wmeO2auTlrpFtB+EVdlL+dHa
pLujrhR7+MlcIiuiEfA0Ibjfynmwzt6MTOoF6KLDFrCLdDhVG2Ph/CB/20UKPc5m2MCH5XLzIMFE
3EiOfcJR1ez0VFiILz/X6WfOlAGjo4uJfDxi/wiDIOjVLmFdiuDGRXTnuEGcKuUs1jg1AOfoqQ9V
dZvU8fMw2IV2hmFhtLviPUnvRFU+9UYzrXOu8PINjeZk4jkRSdLn5k3rIt2ujZ3k9TbRl+y+m7Y0
nSPjVh6OQCB0L1t7WjbBA8E6T4xaMHHRG1+JmHHzGfdYFDfQNn/slUcGe2dMGbwuS4KOBBaykn0P
mZhZjsCMq2vdtvmG4EUZqzejvPuvDKAU6eFLMqdMzVqYBPPwiqw+bOQxiiFZAyhxUfQMpRcoyM7O
zTS7OFUjIklcoBhXA318iftEJWWlKJEH9TzYcq1x2u+WwGnsSuMhIhpfQ54sxKXDlO3HVWaz4i5W
RT1ycS+9X8sSTUKLMgJRZD0QVDCFSucZDTI0U+VwE2v+6xEXrdnKKIEAi/4Dd6HK7cBKlD6CldQv
KotEuChiLwjMYd9aAR1mlmOUepc6r071+OliLa0sl2NxSTxPnc8QrS+kdYDeYW8BMDcxIBLQNH/V
kbP/R9dp+/Si6/Xn9ixliy1N6MOG1maukNEm8QcYta4B1o1lTs/8hJZ6DqJHD1oQmJOGd20V3fXZ
WEaAylxc68+MSacY5a6XL8Dgd5H2f4vqZzwx/RLG85RFDt3ZIcelITbAaBvKFIH/1+FvPwZGMyiN
j4RoIIgxikL/HIVCPjoojYmUF85QDB5NNIutI7WUOo9VZl0AaPL4caUkAXRhs6WSJLBti82Tsr3g
jtaWgc7EAbUTge53MKI5Hj8UNp5R/+5aLMuDCnfpxO5g7mo0BPmCcGb38OiIyZuWqpjSv6Aay/yb
2qnLzSML8lnJNytyUaMLaZyLuUXLxb4VFtRqGAZSGvEx3JzUjFVh5z0wkshedoLzUcNA7ywUNbiO
UU2nqlg3ffAGMyh9j5SDXG7d549/ft6JIcExjlHzXArI+Mn8FUGwoVbZEhtkHVfcMnF8eivNs3+m
gFy7EkJGevXsHsJcdDkr6cdHO/QfEbUai4q4SJQZXhep/gR6E99Lei87Cybnc/FZrlKL1vM4CGR9
9jP4Cjg4RChhW7CMmV/ODESYwIDjTStQea5rjIxIS7QliODZ8P5iXg7MkAh+FllXyNPuGhg5MVpB
J+e4m4t+7W/OLMRQhNt7miiOPe/OR4bHTPfzSlVO5LcOZT+IL8sTb9TpF2zy/5X4+wsuM7o37mKe
BdOhPyF6lrvLdoVWjsXNjGqy2k3WrjYCKpBr1TDiXvNY6GNpgaQkyoVUXDEayDCmPjryoGQdkwuN
2bXKIynScYl6YR/dRz8tUgNwIR025nzmvzfylj6OfCPkILJ60g9WWB/uoWpdNAm7Qn6m1UXoEcAf
XtpeeunElZWdREf2acCe1nseJs+ZvOvfzp+aChBRnepmJysCah8wzy/hXaugAQEhHrjMQy7ZpGHD
2A4hQwLVG9w35fHuNULHRQJl2RvbWujcY46DXBWBj1XnIWtjorOo9Kxhr/Ar8NQn7MylYZ5XBe4T
6Bec3+aVksn2TpPHQk68yMvtb2m/b64p1SlU4+zDUwie9hlb2CEzNfwANvxTdAT8gy588+ommQP4
nQaxd/gnK1HwZO0ZFMT5aa9cAYAb+5R936Rs4uQDGvbfcAdz5xo+7vjRWDGzdjbMhoe93nm++YRk
6F92NV22NolzY5MwwlqaIJuE4HRIi9bI2BLO7rkNJDX2zizIFKjj6dcL80x30sEAsZr1UdfhPvie
xqygHswcBLOBcdMkDPxQFJ9yU/GAfdNKkvnn12wgUq80APEvhaNgVL62ij5JWC6+dBDepmCks+SK
Q/t9MPffGYVrbyei4FKgzYbFxipSRSSTMpDtsBHJLzwD/KQZsKNBaRkVjv8C8EqOuQQj45wUiyTm
PVvy+ZGvB13LdFF8ElD6U37WJk6+KJ/wlm/k4sDm7TgxjZW8XQKaiN3+L9rn7xcVvgYcTP3tqOnd
tc9Q5iS2yYdkv7vrv0k6YzgTQG3bEBmM6JBeN5+pWhsjwRC1tvh6lyiGFAGCQZdeT5hBUZhGNLB6
NXCxmh9AEzuG1Iu1P8uNUhtKL8pwuGhdSk8XnjX1xRRxZXuTc1+EnJNWzY19Ycvg7gPKsnjiBXdZ
NDjyBzH4zfpZ4Hb/xBqHMgFCWiCXFYwL2eadp3vPyvYj6FqxKdloLkJASZSbdBia36X1/Xh1CTLI
LBbqAardGi0X//6Rz6zLKwnmI0qcCXer98dr/JI/shiuJP6iIEZ8FvCBv8W0nQExSW+HjkfsHvvA
IzvvVj6OuBMhZKPgL1DNcuxQnOc9p33a+E+2KpveONS2rZ/uCqeUARpl1mI6MCGjp3yGi1mF/ZK9
Mod5AzmGIY4mhzsbhWoVSzFoXWT0L2aTWmS5YTTU8fBe3hY19EgwjqYjTiFynL2QyAZKDpWApsQY
kqw2IU7Eg9XlZnIUZg+EFGqJTx+GaP6EPp1o73ZW59Cc32PYXX07fEhY8+iGGb5arUltA91bYrs0
Qk0ICO9G69cOKv6aIfL9cc8EMhtI4lHudWOZ1UlbNYg5yev4bqbFD10gfzP657y7my232pqljwZv
7xlmLmKkXSsEAhGrvlDfDixpH6FgPwgUo6ZY+plUe6MO+U+hT60zpWjZeFUTNoXNTQ+ef2I/XGPa
UTXIpdmEiZrz9rhpa/RK8gLCDULUAq2lDvQMfVBbaTo5I+BL0nawJTsUuN+2EWsEA4Ej4EphOIti
GjbbmF2uAz3/fVkFUWaWFgjgoPbHXJWaTtkEVbyRXV0/86RZzkpAlym7OxavJC6HPDaVZrUc0aON
LLMeN0rqVKhfxLyDwYpHqSUxJREC2foPtFCRrml8e8cK6CfGJfJErQD9RAfwDr3W6uKhPdp6kPxY
iWtdB5h6cwd3zXnvWADd0stDyDRlRUXKiDFZWwC9fDRwDjewuafgYVvHBXQ+t4rXz9VuGrd4rxne
AqvcSYuAIrSNaeri8krKaO49JJLfQZpSiG+EmizXVr8deOlxE4uOtL55GBFOFHjL/L8gCTh0fjH1
g+deI/G4BHn2wR1o+ojd4PCVO1FGaf7/sDSs9fUDmhOz+hoHbjI6zzisTxGTQ+XP7kk06nc94cuZ
ozOFfAX1oMS4DLs6U5wKemH+6wrlX7rf8Dw6SCBFpyoRgfaMpq3SsDnAngxzKmAJYlWdb2tkwmUt
GpTjqUDwFKFKZcas3Afvukutsa6Nyw24MPvaVJU1JrfLtxWMwfYZ+mTxs7F9viEdj+hKcPv5DHKW
0k8TqlB9n3Vdl0iq5LRTLd8kt1lSLsPApY9nCNapdr3DSBj06ZaaJRX5+xN50G4eBcvXdkQ7QVW6
lbOhs9rwI2GhEhrusdkyQ03FHYJmvjs/6E99ZABrVcxllBUX3tg54f7fkt9OTS0deLtGLuaOsP/A
/za8z/YJQm0hRLRU5zNP1w2OCwErYS+367+7ZUnycxUQKgh+AY2x8tLwskgxXvlDEa42Gu3saPVF
UTJFbC7Wk1GR78Sdx/X0zwL9EkZ7/yLWr4ux5Qfe1MWHDdCldmaZ73n5aQeMXGPdSVqoj48twksq
NVh8+Z6kHJfrxhwlxgjdvUw9ew/LmZBf9oXnfTOXp+veQiiPgMVmleWj0dcnTZZ0Ia7S4mq8UuRg
c5nKSPURXIMv59ZImItqLipSKlOwJDpA7fwQa2EUXwHjNYW5iEGb87UncJXwzCwFuCxtj7vC1H38
YdpsgWI+IZ7L7VfR0J9MQU0fXDtCXWJTbSsghP/9zx/KvX2kUNXneRzos+n89piXsE7M8NiMoEE3
5bvqNl7zOoPEopO/LvoUoODdE2q9HKPbiFovwTe2i6/5aOIbSKqP3rrPIIZZiO12JPzzifzYtxp+
ZYpV7tXvMilQRr7Efa0CyV9Z06bqR/Q3kJ1yPKKueuZxFvTXLLeXRG7VQi5wJFaTJMHO0CnBSf9d
8pK4/Ppz+5sgvp/TWfLh1G4n2PSKiYzWgjIusFsS8TMnEpxvj6ovYhjBOroMFaSGZKpz1LyPowVg
vH5zQikRzhU91l+eXwTb/hZ8279OEHLXha6h3v1xh8o7Nfdc6oZ9VoQKulYhKRa0sqI9uxfrRkza
w/43NnyoWtsepsncZQQqsoFngF7sNuHEoizcsVEncFB2TAn9g8JwPjxRHIBE6E5OZdpacRr6xoOw
Jc/oeONWu8iiAGU4cSMOptlNBiR5zf2JET96ecRDKXtoyOAp1Cj5DelBWsnwUnbdW6m83EBn4L8G
x0C+4ZFYX5Anj+B7RRn0Wgj1EjlFxFMJEROm9o++Cl7wpkp7PG9sCNscfmtR4YZ9nnABpj29gqmS
nmT4PUCaMWbMnz1OJCoXzJTQIXMHs9f8O1+BVnF4nrBwRj+ZHgLHqaNh0UTmFAJ7w/tqU2RS/t5C
x4TbySRD/r1piHF3mk8QRRmrnRWc8SSFvkpMomW/rAE7HUtSkxt7yOyRcfrBGTadpiNna/jmPu8u
DupaUXSdyxh+jlXabbJfc5+icJZ/IMsXElrw8uSJh1O9rrFARLEfktZmXUySO8nOL2RNNj+KI76i
7DBJe+loLC7AggQuZPMdCrM9xJo8O7DVZjz3ZDXytuNqkoxFnL/nqWascIrGHgLJTeuvD8FkDN4e
GEXtiVgXPDBI5EH0gIiCE5/iVMQ4aalbDBKm1OiFL28uRTsUBk2T9H72y0YDnLVcr2HSBFB+i0UZ
TP8Zbuigcncmrlvo3rGVa5038AYhJ1Kvhy3GV8eAXh28dETdQgnSCTcfq1OIdwME6NOc8gs9Crgc
TgDgHfBagnI//BHpQLgcADFiEBnlMwOzyiMxd1W6MPtymi5fJhinZLYaJ9OpEH2XX8Ma3PvdqpvO
WmwYx+rIrIUFXISYYKlKFw7/vKncL7c7pStvcKUR9+dyc61aXzXRevNCea5BHGnCnHAtfS4vfxOS
BDPI75BUwMLtC5Id+DC+0RxngLAER1Mr73uGVsH4Xe2uYJQd1AZXODJap5A7F4d/zD2OLWCjjuUD
HUImdgqE/sMZ6PvQxdyStVmtRbH2EVmJqU3JyGt4iJO3TQbzm6wIo8ofHWMJ9pINcGlF0I++KEUM
H/Fwj68Q6kHbCBFQLo8CAUVmYuMsTATHt53Qaur53pppLcUuhFR/mng5ObYjK1YFmDyvASiI1BZe
w6TrCBW9pleXZiz5fgLPtOdNgju5G2cvVDHJqtt260xY/mx9CkFQT/JieqdGmiPHhKMHQ0Od1oFx
UfNhoCWHQXpcOg7ZjN/7MLtzvAT4CPNgLoW1/cWmVChioRaiE21F9UBesyq1H7BPm7yk6QGw5vBd
A5sElsKowAZP7pMPgXYdtgktJtzxAT5yfkIv+jCkhiL9KGbJGJN+6OQs34SAT6WV108drG1iMyuN
1/tRopCAJ//uw436k/KMX6YrFaqLx51Jvmo47XuDQYYn29GeUtCFanKTDDTxgbfLfbDn/XgaIoAj
8S35PSTHeWJOUOzDADAkTlcFuR+poom1MwNfEj5SbAxNar8diolRTSeXd89fXp5wHA1cYb3YtytX
24BmR++QSS2WkEiXhhob9FpxBp9XCm0gqwbY8IRmrPJ9uM1gSOPnOdA1PsYr1qHgFKLCUEQ43gTt
Z2vPr506avcyDlHVcJvaSiq181UHNj6iRNiV1x4JCqBpJj50/XH/LMB+j+TT39o/ODr1vqofiIRH
ubiyxPgqBx19JJsMeaKI9iYUtdl3niw19Yap859R2VQqfjN56FaG4corm5i+jn86aJ+JF4h173wP
t4gaw0qjXeqJ/q+07trzfmw8GrLF1ZCdKA9XF9fPsMMNeH+U/iMWhoD0VNzpjQwKi1kh3rV7VZfW
9wIx1tE8IiifZU+4jlYBv7KSkRwrveuN13e3EFCQI+SNc4FJ+daBc+OaolrQQVjZJcHHp+6cxiGZ
C5RjQx394mV5TJtSjRDmnkiSHoWNUI0WGuCRrbfPWwBbkfs8jTQrc3pihrS/ZqcIFcvkadroCTMX
Q8mnIFmR6dSNCJegbd+rBj0gjYIyCwIifrgH15LHorvEN5W82luBA2g4vMTGYalf0oPiTSy4cTue
cdcxWtz6xK1nvYfBVhDDPu/wiEpuJ6iNigrXPv8g25/wLlJmW1rbtv1dnw1kPvkPgZv5uFtOj0ve
zxPJnI3gDKnRdom+MMxU7CNg90uPtbAnmZ5sAQG9y7H/s7i52d8JglMZeY2YcG74eWdqFMN8M4TE
H4iTe0JAS4gk3ClVG/WH3QcULqJDmmjr28yWZyoJsX3I5iQlFn7343JR+JlKIlhPAi0Aa1R/FT0U
GCbQUr4NYYpLZnA5p4nk8GhiY0oT6JCdmLg+QMBTP/KPCvC/fBHeUNvfeSeBYXN0upZG8CpSp4DP
90S29nPOxtZbrPAaj2RE8+ZNqxkQBsbCMDTi258WSGJc1Rr+hYoXcnyYDuOvch3bTZ0YQ1mJ7lE+
wyS8w39NvShLYt/dMU4Tx4EqWEt7ha0OfYKzO/qYjRRpY9kpQLiaqiA3vy+Qrl2VtgRp7apBZjd9
4gtafm8FKnIr04nPoQfUTOMHduRIJmppe4I6fDTgPdilbRM4+K6yYpOKVCEneDsZV6pjs+zvMla3
Kef067r1yJAdo8rYC/JCVkiTw2iZbL0VD2GK4d7pxHWNsDjxcGP4RnjsR9499sik0bRJK1LDLc7m
3jIbAYJLiXZldkMEVJms4XJxN6rHTkXqOp/392q4pPgQ48AXFzN4Ng5JEVPbfqNbVazA/BgPWGVq
5wZj4YbHCXvKj4sce1g8P1IvzqpksZwCcPanN/ryCjwP5Gk0cQXv8pBbt5Eyj3KHl1sbvhfMPMQq
bO46Ji/ICTT8QnhiUwA44NNq9Ta3bzgHmbjjUVJ1T1+p4K0kWlfYDEIHDMS6DztXM6spvIhpzRDt
AYzdhCkdOBhsaukXBsBvdH+bLkB6J3sXSHLJGtlGTftV+UPxY05GSYbVZ5wWCmbANO3R4PIXY8jL
8vXKJH+j+C5+RaYSAL1Xht806MtHPjNqr1jZr6RUWVFgrlqeNNDkCJSUA13hhUuiONoaxoncy7pE
Dsbva45V1ZZalE+h2QCQl1pQ1zKYi1xGZYTtgDfwQ/8emos2t57RZ41zK0MC6WQiK6pH+ZX9+N8G
rWcSUCH68JER7VHA/ZZ2MAoaVLJTuM/7cdE91bOhNWBOBirYp+DNcDXNksinZoEMCFruiq/8CG62
sLNBn3ZzeR5XN2t/H33mTR7MYlQSDNRUbEfeMqERd1WKD14TUKnDdcudf1ISD/iiQ17EyMbXBTR7
os78SqUICpdYNjuKE5iTMMNpmQYTY7iCmNtc1xFKZc9X94qGm3s/oIdZMQnf/8P8ePz4BkgORNqK
9Vn1oZSPL6KZdfKvIp1Y4ttFn8RykddbslEMYj7m/XSNrEHkokR54wIPXidfw3IhOruRnGbjop4A
ryDk6T1he9pZM1plrZWaykAql66vU08aE8XnSOOh5A3J4mLY++ge801M7jov3XrsOZTTQuBo9exX
SrhHotw5Zal+zCkltPRw4jrpK9orlIXInB7v0aRBWhXwTtCHrsJDnJ3uzsSr3BvcdHW57wps1lPO
lIXA7K5C5nURNW9Q+O4bMy/kBRQIvZQNBz+D/V+Wuxr0u4RT74N/lhv9glENje5w5kfdKRN891LQ
GDmdRuMrbkkAUrKlqxSW/2ExrUwkwCoeoA7d9cehxZfbMiRks59eOfBk/vHobYAI3zIIt1FKpYk7
ZPZVNSD9tUyI3KcZ8vHTDyfxVrGTix83vvzSbbiNFVzRzbHNrCIzSDHkePbRyKyqdpwcEOjXW/xD
cZApjjwB/lyNvDlAUqPd/XpeN9ErbA2jee+yXAkTMq3uU+RQnyX+i1DXSARD5O5Pzk5Q9B5TGbMm
UCmrP411bj2V/YSuw5cDoBGj11LfMq1X7Zq/rEXc5uBuHhBIBhzBZlWlWibQYJgk6JdGBSAT8XTA
GPKJItRT+K2nCRdQVRy4YT4XvCBSCKRt+7zIuC6gpM/b3k0USw2mt3ql2FpsFVCQ3tzj43/+eEp/
UB28sCT8CvrkFBteNZHngI8Oh7ZF2st/BZle+D6CylScfOEckWB/yw1y4mdLks+hKqrmEEsgByGS
wyiwiUrrBkyud3Yx813uesMxMhdsqglEjMCbQPe1C53+grNZ9Blyh+qdYXJtCF77nL5i4I08RQ4l
Xr2xIq7q2dN4ylzz9p5R9NWySgcBS9BceVAkDjO/675038aHZuIUPfFSyDb1gm8uI5++JAStxNDW
Oi70s5eQCORo5grF+wgWREkH07/Pq0NWhuowf9WBSeSO0/dLphm9JYIWoePLf8IQlgUI5VdwE+ci
NLykDh0DzwSGMpvi10EgTbsrBla8jdgNQ/vrLh8mRE84b+oHvVJZN7TqGpaIn+B7hGzPF+Y6YJQi
kPUW1oQU5+mxIXQwFC4VojFQV5uYJ8bMddq7vIXLff4TakJwpnmDkqw00XK9NodChcwK6nQffx9w
Oq2EgG6Cq3H/97CugWfprHKDCb3rUUgVWwVSY0DxkIbz3wBEuUAfoFsC3dnrYaeX/sIoBs/K1KAl
iCCZEdIBDCsOU8jwzauLlzoZoKo0qB0WI/fm34cm/T8g+tSGDFuvRula3uaBrUa0RkYcCEseLK27
n7f4XARlhzehbK0rJUuBOgOv8S/gblJJgPtKFrgbMiqUeyb4nyXY/jEynVP2aQ7QXP42pYbOSGto
fKicFuJe2QO4p7Tuu+8Es0ItXMFXW/auW7ZXVBlVAeha6JManqPc1N+czoUQHWhT2nR70RUku6GY
qk0jCAMomyk/0C1OU783dBeWuISq9erb/RGIdSOeuPzxiqE3+mM8L0qIIX70k/T50yruJtnrdAtI
U8yfkkcPNPrsvHyQHL0b12vRt4Fnwmyl9swXUGvbvdaiIALyN99KZI7PCNHFgZioRrodN8TLH8Lx
JckCWCidq2YhTEInWy5ZM6Wqk3m2uIvj9o7mMbxhxHs457ueb5H+86bOmsMfrNfktsDOG+nDKdG2
5WsD69sjcW6mtGMBtqq2thbxcI0nZN22E3lUfLrHChMUYLwcVhMOy09IDhOmTNPyhzMKtmij89Ln
KsWszLE8zLVJQRbQ6PJfhIS64ByS6DW/AmOZrZEQvHtS7ZnzUhcX3pD2MPxnTLokiyYwbgvYopPY
qk+eB0CVjKi50wXdCg5iOw+hiLJ/NqHDbzo914cKTuBa7msQjPAR2VT6ugFfLeyNVD+3UsFdY5UI
K5n8ke4zb5vC9HzjQQltYvJMf3eu1B9h8MmXQuMY9bGjYZXHDRYXVma//EKA+9VVqTLWdgnl8aWC
RN/LA5R6ObRqqs4ONVX700Metwz/Xyav8WnNaKU680kY5uTF01dClKCzU0IE8t0Qj9jFbwePtq5a
ypdu7n8QYjOmsdrDx0DxQdr9xNtOlcm3q11UozssJw0w3YVXW7Dw9979MDDJJGF9oDbZUsnvqyBE
pKm7rBsOCPER0rKhE0DSKBV9PRW22cfaSIJg+C/iCwHn6MTEZAgiME36M7K/Zh6tjSCBFvs9MTMo
qnuo6Xy0ycreFt/idDFAnWjiyrBaA6lb+kmFwjuAd9bkxh5uJy/Ss6ybiTlg9lKQwVoNpb6tl7Vp
SnL5DsOyRSmx3oTqlCKKT47yOq5wFlICX02o1EbFtUza4iyn1SNuINviPzXF1Azj3wAyyIkSvmkI
VpfFGoXo9OHNi7uhqiBBbGcJ3S4VLwJ0omCMF4cCD2Ti6A1bXtJO6m0+nI+Cay6Am0s37VongRq9
+gfLLHK3nJNYZD2YlByUYBbTfn6fIofrDkBxNSGtU04Q2+6gTknEAwk61o+tKgezeBF2H3CqFLKq
rDOX3lzjWxgMITy1D08l2zpDDGSgfbcL8JE2ZolZSaLwMdfFh19SpltW5a9dpgfnxlelTyCFT2YC
Sbld5/+kHMMO8CrqbkRuq9kedi2qJSd/pQZHvN7Jm5V72A1tIZUlbQ9PRJuSeRa5w7SJT1GH4TsO
efuVEYndG3bFLQEV6jzXZOkQ8oZ83/Ehg273cLi49Q3+Ko4hHS/u74RhkwgfR+TjqnAcxELNIgB4
64ID7tbttRQOJxO4P5hULF197N79jhmNMu+1zJ+5uTIo0snLZziuX0aBAyfBPH7IM6SrDwfmR0sB
knHNlEf4/V3yJ96bBhm+M5erVBmdQyYwzUy+P2R5zB/4BYNTqv9pIAPwnXqDqPq4aIerAD7Jywev
jczduS+Seec3+iNiEf9eCiGo/mqYp2anyeROofm2UzmVx7eAGmbrxkTDJK2QWoNro0x3p9JXV1kU
bLMwau6C0xy80MV31zJbJGPjuD0mRsY2VmEO/vsJFrHwe7qOZLm3P+45HoaSNN0dM9+yqVGPit7+
0vFlOCqZGPqYRE+nBPx2T1gfiowNKA/VRgNwKiwq2pyLY17yjv/I7dJSQE6IAKzX9A1sE2jUC2qZ
rjCpUDMycxJOlPlkN3RrkdFz6F7XtwCGXesQrq38Ay5Ru5RJ55C/9R8yQc1oBQcEqLjUw0zbZQ+e
+eosYmLPMIjOaxMUCgJTJRPCp7DLhw1NMFeUpcWCRPodyeRPY9uJKkXY+eJif4HS+Hhp7LCUs2wl
lGOaCCs28ErU2kVo4Hg5Z3HTGI1e3fOAJnvJHGs/zbqTUz63WSrx9K5OWWfxl+BGqYJitCiyTQs+
qcyaZ/x6bLFWrnlQ8LSslriOj4PER35j7nctWeVe1OpOX7mDLemUA4+qeJXqIiKCheWDoBsPiSYk
7poyC/kTq1u7tqrpSuCrs8JDJZ/R6xkw/39R3iCiygmf/KBcOn+rR5rYDvUG+B+32Xzu3K/73TOK
yVlh3MjNgyxt6Kil3G/gC7vEZATTii1zR7N9GyBgdO6DIrHp0F7mBCqFHdBa760r0AWdQh8nQG4z
raDaPXeKjoY/e7B0FsAr0fUZkwxGWd5vJK2vRX55jAOTGbLSzTZv874veHBNjNHI1+n7TyfSTcSY
8ZgcAlfWmLZ0ZZnLj21uU59uBju7jHtbkislqLgkdx1IJVO07LoPAHFaiHLqAUwJOmLELJTjkd9i
jGy3GTTd1NFp0WNE2Sv2JAijZ/5U044sIp4uaRcx2aqM2Chx++skUjUG9LJP/42Nxvy9yUP0bOzS
tlQ0bLSdXJ+gECGlGNXwfj/xSJHzCS5dU2aJqNXdEtVOSuY9gwOPA569srC7ESpqYf7dJU/D6OC2
fZynyq9nlALkUkabVX8Ydl4TzanUYNb04Xetpx61bLpARlhaUcR9BGPc6PVJZ4Vk0X/LEzqwdauv
P4RMK08xkhx2Ckz6Lquees4XmZgjlanK507gwRxmocbLJnyk11PPvzLZJAbQljlNMrwpOFyGphSf
58YWYm2oMv0mj0td0/vWlLzjqhrLknl51VLQ2zQPLcfC0F8h7dI6Nu3GMv0XUjpg7rpzjACIg8Vj
V0vSyTDIU2ATimtUVr8f/FQwRMwHjk1OSbs+2ERnMKL3ZqCNihRC43Xqumc/O9DJrmZaZMCWZfP1
PWsmk6P5p/z9WlqcCum6dhwczptGQCaasjczjpOLmxcMjVdZpDkITZPdhfhslFyKFeIozxWHcD7v
o+OqRenChFGs5IrME3l5PCtNXsPOmKIrr0FXIa5QYFy+WwOFEtADAPjgM8341wWTggRAY2PDeu9a
X7TScKrsGRgTnl/HeFndF5aow2R7j6xMl29Ot7LvrmM6h0HCZvjOu/Fjkr4b9gW8cF2DlPDLN2zl
FmDhu2oR3x4ntAjGZtt+q/CioM0ARGwBjOF8zW0z+HcTXTXSVNl2WN0o+5hG7lNakKQkd3PPTWsL
knMIsPhxyM31ys0M6a8NHO4X+2/375/cGNY9A5ZGByn1rROoqRmzMTkxEvQ+OqaobHMQUYDuUzO8
H40PMhaHAwnsn1oMCR+6DdQJDoSuYrgcxhruuGwZr0u11Mg6EiCy+HV0vX//uTkaZUNY8xy0pN1F
FAEuzu16H6bp6EoXcElcGvkhVCuwvfIddi14HTmhPObqfweXc52ppC+QqoEzx5ABbN1X5c1wYf6d
G3g4B9FbmqQsH7u3rNVEhrSGZjwZ/O6J+wIIyi68r3nV2430N7Zd1NFROSFPCmRi1a5vEJixDWWL
XBGLqVA+9nsHsHl+kldIkpjJgRmeO+dSiDTRSkOwlZf7kFPDUrAYRgmfs4u+AWPM0EIca6/xtUvB
8egptir2zDvsA0lov2e+TshRFbkXpCbuqjg2xgNGNzEWjev264Iw81G5jUOveMWoEeQn9WjG4S3c
o+zl5QuT9/DBwhpISJ1Xf/SKhjMdMk66AW6QJ2OnvJnhTbvASFuxBt3Zd1RPazYcChK5+VE1WhL3
XexD4AVbNAb0+24DSMDccEW8lYfnT2oLtVlQPr1AM0UQp8R1erxQWNT6jvmrhrVUDs5Cw1UfXyIT
GhimzDkxpIdjv9h4GDvt7/qPXParPyVveb7INrpyYZ8TqRtTNX5e+KnP3Z8A1khRW5wYd2t22RAu
g0/d4PJGS0vnR0QFPaO94S/C4NlL5Bv/VlkrTB5Gm71zjUxXer4dBiIAbrPNI5yZ+wf2AUIDUaTt
k6h2trbvMfp7zNC7MYgzVSm2Z8UiB3BWicVrXMdCUc8yX0lpmql4u1rDp3kJaMvtIbfS/Tfa/C9f
lnVKy3ihIzwD6r6okkIQ1J77SY7ev6ErvHSLw90OPXSnq6FUhl+MfiFkvg3NQLMNoM+dXuG0TUWx
iljvAT9tcyHiviz+on4dPXPm+Szk375ttD6epL/EDBZTeqmtQ25PZqZx1vMxvmMSRKXLhbg7PWod
eVDDC3LVUkgIsC7Q248sDgjW0dn4l4+H/GMZ+YzSt+0tqa4tsu6XAHZUBxg11UTKevlL6DCU/YEz
Z8eqENCZB9/jEDLNy8vcPnFh3z+BgiDhaAUING1P9AoX1XE1yGpytt87p+Tq7SzIGRRQzedwEIB9
rS97k0KZpIye+WnCFvMziaTZREXkxPuMAmiOhtPn7ATE7tJknDewJ7U8G0w4AUyJj2xwqD3YHuUS
o0b4O5amVMaVeLNQx6ncQtyqv9DYWVpF9Rsg13QxxWOrBeib8+0oZ10RoGW7dIVU3ZsDYQv+6tIV
MZSTh/9OqVMJGiM2gK38orY6hCzIOVXLQ+GOsbZ78Tmk/M8iCYfAGHkUZMqJlmuDSxcQ5hmcJ/n3
w0xYRKRZTu1hbO7Cwgb5eOGvUKC01zeSpGWlYbLuMTSCRjsDmO+8kwpp9Hp61Veux0ghS9ErGuuD
vFpLB6lLD1Undfe+62yi4a/9eaNNz2c3ChPrHZRGDF2tIdfm/Fd0VE72GHA/a3AD2ebet9MkH2G3
TeCG5kLEqAYLrrgnPjgD6KpxCAZSsiwicQcBov2k8QXxxc5lWnRfGLlJdzyBe3bO/VT5YBGeckWr
gWQs9KABItFIs9DrLVvdZmTXYT3Kds5Gbe4CQBrQF8vvbYv19u+ZDarjNFAxpMPxsRQVLF6nQgIH
Oa1mo4vF/1WvEt+YtWVRv67StuYlH9G5+XXdqtCCGNpCs6uavMaxkNegxdVShhfMImQXXNp7Plwu
hmo7lTcj79x8so7MTvRfPPjL7RorReqRtCi2zn2qgQFfzj2U6LEZbwNsHxtVIdI+tPZqojqeVNPX
rKCMmhP29HRAENZS9pim4wMhQPbhwWRbq4TJQPd9z4Hf7jiXFRZZ9fj3XCnpfP6M6vHJCvp2/qY3
XCwjrEQoy3HfEcLhQFGb8MNvx3qKk0I2EsyUlekZZw2LeY8Gw3wIMD/NW4z3kujSpTkWLJr71Zpj
CA+rFW1V0OXiyeHX6YUNd8txM8iK1HEKvPOB0PlHidSnSoLFZJBU4gLweIMHChGkrp9iSt7NJQet
uJKSsBUUruVaT/2wtm5Iqor622egRvc56LXjsT/Ag0IitBCKOVKn6J43LMdQjuN0FmI21Jqh+ZN5
uEdMWQYXMtuwTCZKPmlBwHHL8OFsPQvzeCrT0yhawoeHEOVBBJwMdSy7mD3M7P1PKNtHH8CXAEfA
T6pI7gtKpfcjcqDgeWW6foifEqwmcGw4gTi9GGhCVtpXQ1JNs156ksZshUOsnzrc7OinJ3+jIlyb
m7OiR702/QJPLwdx7ZzqhsMkjkvJYmflR0eFH9N8wUyBD0wBmBaMBZ5tkQw3dX41cTz9hpmEvbbm
AZMTg6+V8YUyzwGWXKc/rZS89SoglnJdKE/W81chmYclK7Y5X291vqVFdt1Wnt3AtBFbWI1FQHfK
jNW5JXPK1LoEUOVKLVXK6hqh+lHCqNKrda6TPUx4yPBbJqlyJoVe3MhyfEtE2VufodAaPSx1BgAz
0jfAZ/Pt8iRaLpa70yIZk8QkIilUhog3d9uedq6tQkm+WlAxprcZKOh0AbiLhUYZoCQZekqkSEPf
vHw90RLQQIVTjO/RHbx5T7wpQKcn/wvmAMCVHjMxbKX38KVJGWXarc1JZd3vvGnFKc1YTAguN/JE
9gh4pvqm2lijZSyT66GvjydODvFxPxiCgS5ndRdgN2DHq9j81E2MsRQVlxB9ooqLyYQzrh+mDP9H
V9bWJLCHqGEmvZR2dWRTmZ74t1YbTa+lCz/sw2u0mrrMt9OPWWHZEKWTfnsMwLPmTZyqRJpZTIyb
MSh489d8SBqX/nnlw+E9d3ZwCn8oP0vB+LJDZIsx6W8+zpf4nuAewvxuZF4ZMmd1hEV3nAXwNiQx
h7YjP9SUZE3y/nU1lCSn7/5MZHbDYusBnwsCM5wP0VE92xThfW04ew9IOfmpiWgdBDZPvAtaTERy
txubaizXnw0I7ULvF/3xtdhPnBS2XO0K+mt5YDhCwjVk2Ek5bpmk2iFGqreRgcNjH4DrV/dnifI4
m++/LPNyv2+/IZMVzIYSIXUO7XMPpX92oO3N6QnkOjZP3yQJlrPNgy4H/AXrj6onf68KRMOcO4jf
Mm+c9JbP6aqggs4aYctgk67dChjI7ZrZFGWkL8oJhhOnb+YQ1jRsrP3pugsK7Oqrdy8PbCGYP5ab
BxPqnpMpwBsr/B5LQIDs3RcAbsQoJ5BScnmGGkjnN0FKKLb22VnnmYl0GZ/0vx3pDEJ/GYPMJpgL
ojKC3YMb1YLWmK23xjjzZ/4zrnHuJEAcIgiMXKEVePPAda7wIdL+dTg0oh0LhHj3y/Xo+wtEP8rJ
aTXDYxrQI5cgvGNUO+Apch92CSs6oU0Zwdzn88Qo+TNCs5nopg6vy+1RPZUvBNvKisfyJJdVmnEW
OOimxZgR9qISbz4NL2u9D6XZi66th/+2pFEadcpPWw+zw0EJxKBO5/EB/j9CA2Mi9sABQ+ePX/jZ
+aKUiPOv7p9daGGV4oWdpxWbUJNmm96Ls64z3Nl/TikHwEPUc6kC6XY70c0ahLqwkSebB8VCB0z9
k9BspKZI36QYlhn3SjyuGa4x9h8ldDJPu6wd2qKeySJIFghX5HkxXRLMQgoxXjhbS+k9WugfiGho
9YvGz6Xi6dyJsf3CGmo6Te+fB/+Zn5seGuR0/IqdjK9H/i1zmCM129yAsPbNMxfhSSapNLBvgEFw
ML7miLr68v2kmTU61lx8ErJUKRVuAk7q1hfDk3CxFRW/0QULJg/QyjfutNL4u+5bqywzWfxjw/OQ
PdBSWJ1WhKUa4+Y4YgmyJpF15I3NmryKGOk6H/VRe3PojGXYbvGQwv6h9t1YZcFx7rdG4UVyr0yD
8vsTL1uGuS87L3d56tbhpBFcehg+Ptkq7EeDzzqLetZw11ffTdBqgsggpJhfqWd2GZ/wKxlk1h86
megrWSEqvy87GCnEd6+BFoobJfbpTdhaUeCvkrwX1+ydVzxC/Thqrt1H5NichKlJqzz+Hbw5T6EK
12f7OdIMa6quNRKQEEuPo6FLCZCT4RyGEP+5nOa3MO2aUf8jhmfL1I6Pm1WJ3/8ChDmIwzPUJK0p
KnPKWzqxc83Q+xlComp1/ImNDEXCD0DhoOrN3Y875jTfxhrCXist4pOFmvSUggs9kN+YrpxRcOdd
HrN/UjlNH6tTlQiUhya8yyQMdER6LB/XWaHLxG3qYtlgiaXNi6b/m2lISZc7M0/2ON+NKv7ediKj
MoGFeL0y99U/nMGRTqUNrQZvyqK9YRUsg2OHVM1zrcDT4g40MX3LAiHuK/Q+XvmMkWt9xc6N7HRU
strdev/PhNt+bDRyUlgcbfOzXxFLFxwOgkCKfwhO5/kTcUFbper6NyV1q9Xd3LZcEIye8evOrdfy
34m5lWL8CxGyD4qJl6EA2+qm2vhBSf2EgrmOO8xVpsWhKgaqdEW5ES8ZTiakABf7jGODHGXIqrPW
ZBmoPI/775uBD5BEm0UXNIHsro6h71QvQviAtc5HFWNhYjzVWWbGiRCJMD8c1E7fFlItcjooCs+a
OXRRCIjd9AE+MvDLUMArY8IEpYEHgkNSkhq0FMfXAKJzfpZkJNIy7VgGaTGyC9GKaqFk5fbjH8vK
64ylZJBDBvLTXugyWVLNwYxl/ns5ET8KTmB5qsSDLHREbnDiQWOpRwSHBST0T7a3knq80J2z4aNP
qkMg5KYbTfb22BkohzXOrOwS14025TyIBrwTs+uvqroR0eAlb0bXgWUVwJDmmP81aHI+MMQW2cGA
3dGaQG0rw07EaDPum9FKToemdOm7B3Jf1GZiGMT6kUd/S+mZMI9Oo4mjw6MBeDDaLbsEDZtCDZR6
YrpxOh53HyFin24cr2MDHcHtFyKE7tvjm+/u3/zwjgczuMbJdri1ruIzjg2JukcYIHJaJXWZbI3C
u/0eWLJvdCiGd+L0knMAsRONcd04Oh0o3QjwTGgvjxdVpYhXhTD9+PXS10e3tcnB+NcWdb9QJveU
9ouZy9VN6hY6+kgzAC6+0TFwpzlY8jeDobmNSR1jgayQfiqCGR9GgRotxOAz11wnktgeUpEqEjz1
5x2/blVIuL7Np47SQcvbMWgjJTwD6szEdbEfnaXoQ74hicjF4xJzvyPbUojxYbCXjsKZCyz7m1+h
IZ7oqvCxzpnVMwcsB2aO+Q3WVhZt2hETGz8g84NSs4XtizpOCldDQErfEO6jZFsM4EmiKjjyJ09P
S0JJbQNegSr5soMsr9n45ia7G6QbyGFDrabc2hPthEig+qHvlSypeDKaYYDHnODh83oz4Q9Qj1Aw
wZvZB83KZTnk6idLUTx0OXUqsDPa0x4BRNSDfTJjY7hHz2beytvIDVtzbJ3Yf2250FMPCSRFngMd
sS5T5m3461kRr+rwV4UqbHwbSGRFNKOhI8KAzimi2G33p7hTccRmosbArP8vHqum3Hnh9CO2J7+i
cm0Y2x4fugo4r9Qzlmxqo/1F5cVFj7u00s0SW7/O0Z/uP3sqdpyzl/HyCD2topqTsZvCW3g33/dU
lTnCK/etiX5LzhuVWDN+BoulaOL92Idc5l2SDnbdme5FG9jzdg1AotqGqsleSAU7qsBw5v/+0T/P
9+LBqiyA2hej5KZwieTPNjuOb+K2XO7uHMN0x7uxpcMLS1ijT4UgiKgiYfb3pWRwrqXU/shw55Br
JiyqxTLD9CoAWXahOQ/Nthpd4njk29QPD7x2iHJC3+zSTnWK1bzkOsVtvyVilMWmSry8tnTctm4M
DXyJ2GiL2/0Z+7w0RGSnlO2lKfFIMd4u9+ECiowE/54TxpF068zHznXqaoCk70VHe/ZFk9vTNPaB
LpIvtm9binRAiEwQkoBfVOzTCgSLPTGeSLX/8Ih6F0QpOVaD9YD2zDT9VfA82+OOWqDr/R4vnoYL
y1Fkj5MSZru2sfR45cIHsf71DYBVxgqdlEeBUpIjHFqZqjaRpoHB467d+ZCQc3gV01cVm5TTkOi5
3MlrIgi4H4ig+C7NW4wuj+qobx3ZrhiyB4+r8Y7VuHmFJnmnDrEPMBU4hJv1XXQcsA6iqct5qwQz
R+yS3+f+Tr6uVjvfjAGBf/Vedn62YZmwJW4RcZZuyOhrggAX/VtgGp+/PUE/b0eCGnJK+xQEPW8H
zae+jWPimRnLf7dSR1u/kyhNskLQ7RqTtU28pZTdd+RE1Ao/w692sJOp+sd+5E3EG6EoeEu59noc
tWMckrBG5g4bSdfVBS5U/+8d94XxhbCyM5uP9LTwzBqEl0Mxd9hIfVJVEY8RVoISbsv/on3it3He
2jP5lZcHQe5xY9PohJxxz5W8zEorqCLItqJs9Ff0evj7tywD/IHmd/EzH38LrzCfHyaicrWOnhuf
woBGW7b7D5pBRGMIhd5XwUxSg+MNbp3sZmUyRt/h841xjF9x3qczFJd+z80weey3JSa6gqhvXT+/
jNP9h+N1gRhZq1ai4j64UGsu/ak09W9d10JHVWbQD0mtSJS5NcjVKe+DnMMM9r6TSW30+GRq0wpm
1DfvuPCZMsBlnrsUV9H+7+F1jn/VgAZYXM64+QZE0OFlzFf+klkrAo0Db7abU8GL6P7Z6v3qeNZG
3bG7jmJC3eiLH3/Awfk1iCz08GHqd3LCgkgHPDbbD9d3N+cNsGfmeID5bvL7FpcYec36lQl0Dyfq
hS/GokKeQcDd/RzFWI5UGV2kYEbk4oS6tRX9KJc3rQfnowZ07wEdlRDhtGiY1mZjBuX4Y1yemAPR
dSfuc5DSuD5sO/HXvoH/0jLiKybFgUwn+BubBZhYbmoO68Jer5orQvKl48ZP6qTH+meafeckxC5T
iJK1T0oxmI9xrowMUynmPl+PqpC/61WFhaEL5sxVlAGEPD7zeeXHaH97alab/fC0zs3S97/7A5E1
y3EB/Iua/+Q5w1aegczYDdEOgxiOJGd4tLE/iJWlXLEijkHaUw0apqjhcXklicHzK0uwgW5z9B36
f+sBe3wz/I99G8uNPh7n7v2ylGeKzXb0Pj1lXoYU9p1VVX8gPGesaUyGisG45jKVHthARwB4GWVq
nyZ1TZb/DTD1iJhx7PaKSGpntV1GIAuXWptaRexHAgwUOKg5RfhMf7kl+XXBauclGrKt5aIDnsMi
lmyeQrr2nMiVK+4fw5DrR5b/6OaSotBcfLmwPcwiZGHPlrVJnxv7yh0WL68/PGJRr8Wh3fc6D5n5
wi7b7O4pzW0Ofv8zI43kb6yY55jnw6EPLJmuZS7aJLvFtFm/keJLCNbtmky//Swl16N2WP7lEoly
AO2YVkzvB105PhN5dQU0mVf+U8nkaF/Yl4VDKEWic8NtyFtfgDy93vWOuR9q34ywbSVv2xJdUeM9
SBfhQbQoLVIIpAh7VM1+yDwOYZIEmEmO178Xs6hmd2hQeDJT+/CK1OOibml90Be5FIcdFA5Mbh8R
D2DhTwqnqE1JC8mFbInvZRqnzah7ynBCoJyzEtYfoicgJBEW3maGidlPktTXynFcyHoNaJ31XxJt
urH2wm0PyjMWIEVIvq7jGBHFtWvl+y04OmMEsTjI9fYyas8zZU6WDdIm53duzNM8ydTKGsSMrAAe
jUVxG2TJshiXXbFql+FvBTVTFxmiQYQeYsDybypJ/Z1ix/Bx2w11mjDT++q4hWgl9Ml9ZaYuqcSI
2s9jzWu5PLIIH42lvI0UINxM4+6jk9/145j01pXdMgHVAxU2qPB6TWbA2SiF5sQxuVYxItpnL9dz
wc/Oc9lEOCVzPgNkYx7mvIvD0NwQBEawK0rdFNRuYZq11O+A8+C48qavvfeoLAx83shF35TgLIye
8jUpblnbKNhEAuA+RxgpWV9UrGNbl+KFo+ZGLbkjX+PK7weWt2NxsaNi+DnkEtDKj5NzyFpzy/kl
XmASMYeNc0zaWeFGjt+Ulsxez22LKWUMzNiY9EDXJdBYsgpMvAGADMBE8EWzux7jZXw33K/VrC2X
BPH8oHnp6WsdGKD+DDOhlIkzYApx+5n7vRB1mD73Upw3bbxzd/L4Jk6aEKyDUR0+KIRPOpbHMYW+
XwgogKB9NyUN7o5CZBzIFsdmErR/ZmQDKDCmNIzCHTGaWsbXFiAjmCvOppY/EHRN0zRR0Ciz2L0K
VnWcXNlngA9HqxZZFkjsgl8tSAGiHRnYIdQ8yBhUSBwpuQuhk+1AysdKY0zTffSY5SWJbpgN+0iz
+dWxRdFuhD8iCMEacrQ9WuzxuF1x1weVBLzgHDEhpE7O3f/zeRM6G4D8Wo9+1gdF0dEeyVqoAtSe
heQ5PiQwk39/K4w4tTYNF2M/u2L/WQ4Fdy88tUp+T4dA3X1H+zi1OnHrIgVzpSS1XXdRHpR0P1LF
aG/9OGVBwcgE+wYcFG/wY/j6yymjT9+IrqHpZzffFK/xNQNhBblVQoA7O+CpcXyTbc7ABNm+Hb+F
EmYf8ThP8+ryfK92SGeZbXMvXqFP1XniAH+52lLbcSeBma3lz2qH2OSTqn7AQ09Rmc51HcDdkywB
fLWvGqvwZSoWfmRAtoOZAu1D0zLoW0RZKE1H8D/IRkBXxpxEUEnJn2xsz+0xWTWmP8FBrv7aD5Wh
1vJuoAN6Y2rBi/5QYt+OIlGnVJHJfCzuSWcDEqQPkk3aC5pTL4+AXBUs1CA19KYGuzpaqNR1Mac7
TNr5IMQdhLWdMzhVOgqDkA4oe5gbXDVOs6UOXMsEUzaa6Y5DvY52oj+9jkJ0n6oHlwbDb1IN46LO
oUU9zm1TFsnFK62ilH9cBnN8HS40IrmUziZFkRqp/jSbg4ejepRB54NUYE+ks0KLQcU1xfialEcr
ZJsliS4rzaSIODC5cJ+9nWqKB+dtY2pf4s0O6wirQQIf+ikFdUrvicUJU4jm5Xaz/uWCcWnvVhpg
PFg6oYR6D3NRTkBmu6CvBZdVGed0SJZh2+KS1n0r77VDsI2VexJMzReP0/0CmcvRMCjYZWixNMkC
NrFBKMc7jm4tbePgPtbgSRbj42wDF2ypA7dVcfkXqR8ppL61Nh3lbQNVIxyoVzHt2nsxFIgmqGyC
h1sIM9UkPZl6YZCXC8wgecqXT2wXllybK2Ft+BJYHg2MdQ9UA0IWDVERyAZAjd4UYoKQzm9OyLOd
WvcgX+C7K2Q1g26GnvglaYW3+6111I0cy9iQtsYnPVY2ipiMK7FV4GRRN8U4WYrUguuQxrGsyESk
btlwpdHqg49W0UgFB0WrDKaHI6beRgUuPyBa1D7iacZPPdzQIpT41XZhymdsFXcArGyvtWnkcAgd
QtB9rZFJMhzMlgCb0g5gSAoASfhR3z1eqkLkEKJkK+yN3eMQyA9SxLxO95UK1qUDOn9lvdL+3l3V
FzkfKp+UYzm7q1L0Gekz7VlzQOrvn99tI5XxI5Hu/c4+WgI+wcaAKzDGUw9gkR+pkWBRwypYsA3x
mc4iudpFf8D46h1OE91TTZuiTjJ3wPb2Xn5RtCtd33DW1MyNPxzNvq4YuZMaeoSv8b6Mge9sUGy0
2RlImaQJiXX/GnAO7+PhzjtHazXKCJSP6NnQkxS5TeoceU6H58/+ddehqngZTkjb2SW/kxJfFYZ2
uw6NmrV6SF/jQt/3tdik1gmeBKycOukf17yItQcm0gzW8/wMGGYQ3xKoZBFS3IfgX5Ryg9fII8mr
xKkgqL863JeXzAuQ6JDXaSA5mHmgAuDISWHduEkfpZz1YE+YkLMx/MWrh3ZcWkKHUcTsozprtr2d
wV5k3gTyfs8x3j1em8yY5Sx8tXNaoj1mlc+otadHWCXq8Z/zMpJy6sPxVFFmbWNZDqrZrWF6M5XS
z8DjdT2mbWkEM+4sOWedW3PHSsJIatDrjtpkmMm72PJNegrEHCSQDMVOJRkJxnZN66c2pH+7psbx
Ipn/wfUd9ETqPlT+qFZB3d55XJ4kDzKy/zMLbgVcosueSpY+RMHi6M7uJlWVoy4HnnLoaLgGCDR5
ksaaAeGbLBVgL/YBsHwqB9+S+Ifw/2UWVTk6+dSDjFruAiU4nQMBgcEx8pmzRONOZdnhfZaHejFZ
GZefdXh+j/1LTSpH4+OLFZTXVcPhhcfAPpU0CmZtMDPafjic78mcq4LvVDatYJJoUHKAsZeXslkM
s3Xevw38HFp9X//9twmejVZGcTi9qFxMsAezI1rWTxc2rtu9CaRokMtM4wFHR2aLKmnEZJQ40Yzl
FmrCsFValemqGz7bRxiBU66I9sf+T2zeDrGtYHsAEPVwq3wXCPvbkStBmF19eDhrQMS9THeWFuvn
jzDA5i6nXuoWJgyhkMBDwWmELYmIHA9IINlGnswTzbpr8gpRBbxkvTC6OSjdW+m56DVTyrlG+hOz
nQC9K6eVr0RnjiOwivd51UERgHPrUe6MNbKAlpciK+RQL40KwOTZHnP9Y8zbG0GT4qhXmF0yDoOC
v9d2/H2bJI1bOMugoNwndEmAUdGDaOQFGC8++fUSQMU5GPc4fsx27MrDZNdYiFPYuHj64LhHHqmj
twaqtkPGciP3bPPlyohENbYc3oV125zf/A7yslGHyAKOT0TzPEmTIOJilRk7caQ7UH/qx4FuhfSX
bT0R5IiYvzd3hWgrMSWyQfLGqnkvXZ37Qq6TNdMTShxI8r+b0HUH6yWMsFAYi3zjDxoWIgFzcNjw
FLBqdZJuR0h6IdpsY0qIkr+EBYIPFi+mIieyEG+zBNV+KNzuN9Vr9D4l4vUEmaimS/tgQdow5nYq
uAJbjq0kFej/Ke+pp6C6LIkZ24LJ/IHicNNCl2Tj8zocZYAPRTPGLV8XYsbP2CZ6Kc218GcGJWWU
dQEtCzh5PrJZtanwcI5nvKtBZXgaGzpRw/CiCNPnwzkRZ9mTdusOP/UIOMUnfHvC8XXmUpMOkXhE
iHP/B9IB1vgF9N3w66qhod2yLoaXkKXcrcOvPhZtjE+kLKGrBjBVTxJGb8+kt4mWSeoEqh16Bma5
fEPOc75aHrcJ70vfJnzD+jnb9l5HzvRPkzQ8FfLxO1uZUfp2b9SlHsSF748FkSm2n92Kpn3aj+wL
c8YKyatiF/Muv27fLIj+fKiWPp2pDggqob5ATHqLU22xzTRjGV0RbXcs/quxmYE/fTdtqVK/FHjJ
myBGcLZM4JhtvgD1dQw95s/qjiLSFjogVgd1GaeVbajh6VZjqAVifNj+hNPUPSOg5y+1CyLXDTZY
dCh6Falx6Yh2lcAvsphus8EEzo9LXvwHAHnxox/BKazTvQmPQ00eqICawG/KUK98YhW9fNNGPkFh
jeanQQ2riG0d0lbOEAOJt0Ipec0usc9f0yRJszJ1AUFN7XIOFnr4qy2kGJcoBNp7HejJByttYnlx
HpatwR8O+Xo2rZvf/IFMzHSVsvipUEjQ6VfgL202h2XyEbMFl8ckA2xooB3C7rSuM4VAIu95x2ti
znecJeGmZMeI9YWwMOOh/8vz9KxxtxmlSVQwEGYtWiTx59tCW7K1/gynLjyYvnkpxU2LqDxCmghu
CSdY/lshNlpVzBzb3/520YQzuGvHnjUjSddzyR5ZzImZ/yPj7Y/MKqRJ/vgvTOyoNW+SSoUAtmZT
dY/l2+EUxC87C99xtf3a+LGyjG6ptzSTQ9Vl6s09Lim9GnZSRzUDqs0QAdxLHWUcxFzxcwM8e+jQ
ywiCX5EnVP4s2ez5BVcwYMzLJVIaOrEmSsIcyzlEBIZ+NEEA5dM/e3AfpuiabeRogaQG/MvOdn4t
Vs6uACzuHVYRtFVCMSNHUVTojqj97MQUIfxBsfqZZefjzYqm/JsHb+Lr51H2020D8kxVW5/f0si8
rE35F2eX474W9Y8Pkm7gizyUBB3Adjfk+9R121bcu5UWx4ByMWIColnjbenj+l1QZjQ2qzD9zZKR
WHHqm2T41oScqsSD0u3dcMx821OxUOHhJZM4aF7VeY0CIYXbaf7U5CtQFGpna31MBYNj0+8BuFjz
DafdaD8rq1sTli6qscUntOmmVKI77c8mP6UxIlj4jiO4DAVGB53qW+5Lm0n0hhFmb6zi5UDL8vv9
NWUv+V2TEBLutQm2oKM1r91u/fMhbPxZ3yrGBvxCtBAN9AYimMwjvs9mxFphhoIzvkqX3Gmh+vyL
YARJ+CAzEd+JYV7Tkb8RCrGwVU1ml22zcgjJeKUnQ4jXhUSP5Ek3u1TYY8kF4FkXoU43/zIgXcSN
mFOGM5AVyNFwZ8+aX4C8Jg2GFXRn1pyA1Tv8ocVEoxvdN5cVezCpO9xV+m6ejiOuqkrAzQgFwuX0
yVgwX87PaKk02fjcYx8UEMSygHCt5s4TrPjEpWV4IA7H41slUxuj6Rx/PavQGNXXyOSut6e8TTtT
HgkfJhiyj/FRtzYm8x9ULCv/d1E8hw3a3CiyN8NRlrEOKaBkmhmdWi8BGddRjitaA5xBBJZAT99u
2cytbcqTpgVhtyvxtbzM9GPCQj7SoL18bawsMz1wD3xHYsF8F2dyJ28y8w5V5Uoeu0+WP7zs4hie
zRvN7d1pzw15QVnSE2UpjwAxUmb5WRyRpjX1ucH0RyakKtnULZBJibZAP73WdSH6Mg1oG4UVBGJE
0Vda1p1jcfWd4lQGYHWzUHu63WpzjRqvG/SiAFTn8VBjH3usYc7q59coFbjTya3B0r/ktSD6orF4
GyglW9WpeP4VAFhUAj0N+VZK28kftroCBCnOeDv9GGyiXEdAV9qusTWYkBzwfQW9LHiQdxyNE5sS
k5p3ocqwRRInRKx4w6kGl3lHP72dNlHP32ZaJlytBLtKoNWKfNGU99yLD75GVSW9dEnQfICWKsY2
GaLBgzQLBRaOZI17vVgb5PpZd7Gea+Ib2B1Izrbb/9TzwHqtsPyFCt/kncYTykGxobwZZo3JSKbT
oQfXFhb66ymha2DRd/oX2Cca8yehfEtR4VL9vtrHMnbnQu4vLeG0x+Fu9ByGLF/+xFTf7dONTGQY
DLNp917MAOBWuqTUvIlDcaS6u2r279ctV3naWZFcP+kmvu9cUsfuaqYapl49ydeguKJ23Atrv6HF
sSiFo/v0vo+4lS4/78R5zaycATnQ+1wy9Uae1VRefu9RTbqRYL/2Dd+hBEfszR4TAybPwM8r1rJ1
b6oqyi1N2+75vHG0SxDvFvahZbyv9VD6hgrFIWvuOUphCQYXGmAWcxpO0TYKG+jTjWVEeroOo0YD
MNVtbqXNUlmJhJP+BAPHluAcLmlxJuQEm9a652nkC0n2Ky2n8GWG2mOY3trN7v/HYHmFq2RtzhDp
DtABRZr6Ak/eeZ+DT1XxUcEkYGvKfRT3tvUaC8HYr7doC3lfqaOtDvv5aCynBJ5mKh+i0UNb2/0D
bv1iifmpbEDqIhQmt38uZvUo2gEuinLgPY+XXdoeGal0ublVrGq9XKOtRLmmNlREHxX1QEAoTlkd
qMPriSJQ8QsB8O8iEqEZIj7HYROMg/8L+rA2LwXXhValLnVaZqhlt7DOKw4Uu2IP1PQXMp2/wC6Q
1it6bQ0D+AHK+Oa4wNssUFPI1yQCcs80LG/DxMvM/SGXbNYMedOFymcBK9I1dJRgM1oWKZ5Y0z9H
6Q3SPYuQyehgj4CU80pnN4xJfs5Ydp+27kCFwMArZCG5ShSK8NUIxrBSY+d72MF98l7S3rMjdjOg
rHsFXvGlDvAODj2lWaEBnsf26lPP8HVREBqXZWoeSL0gAix3tAR7Bo5t9e5ooXrX76rDMt97r907
4hFZ/j5kFxwsopZh3Hs/39qfcc+EN0q0CYJMNzaEHkyvy3HfGezLQGD3jWiUcJBdU+ooedWzkufV
KzLQrY9nznwILU/Owog3qq3IZltprKxzBa+Q2D3h6oFmPaw3mAJFDURRr3XYMHRsLmmsZxD/FOti
MewyeKtsiisP/ZbKnA7P0zBFpFUhIkL09xVN8VhnDgONEmgs1LY1OHwOQlbOdL2kJeBiuexmrlcz
NddFaAPdR5vtGVWerqIIjeT9Gs+Uq449gcFNcIu9pEDjvWKgAb9XppVtYVdxB7GT/oYu5DnlAOSr
pyujf1rRzxteDS+Xd5a/yY68cYH0acOU4JkmmxCdYhbHVjOf8QHp14MtsSfMVe1m0pipHGueArnF
0VL/ZOwyS+OfbyR50hvWuRzXKgySObe8Bx7nTLoQC9B1oHaieMWNIVqeh5vJDVI3/nDLwW19sg5Q
vjcfht4cHozUQq4uE1LPDshpdFNQz+Gh7srVqS4TPwx/a4RiTIuu0w9Zgwpl6PLqRjmeNo8IDBHg
e5SvP7L761ecN3edM8/E2X3weIcaVqcpikNonkU51tNG/ewY8GWCavZK+LbiZ8cdxA1E6vAC7hEb
0sV1RKUdwEgmJa41kaJmskB4ghuTy+5s7WUeAT+XZgAb4leDpe2wqJS4eazF02813hssEeStlRf+
ng8DylhSq7HFfBLqHmyLwdiqpTO+x0/Ny8mFaOZq6SuTJsyCNKHTeOPTG09x5oZNxXKe+tWKLjOF
XkaLMM+8CNVStQLDbAG8lIp1sW+UiV4r+vqYZlXwIiU3bMzqiQjddj6g+aH0PpYD+pChCKdGqxqD
4aVTID8sLpDIqdfrsZku4pa+r1yCbNQv8QSJy9rbJ/76zKcBESjpMgDBwYCyeQgccDcyRxjsSSdn
c4s5M+iM9n8P+H018JUfbeIKMJ9wRoxuJc5QuQjoRe11HJMVnlI+AHYzDn0gRoNIc6HPnI92xX7r
olj3HAghGTlcuJhQ4REMT3sug2YoPbUJvcA6NLqGckFpBNLBvgr52jig8G1vAQ3vXIFW4CL+YPJb
KdA3WfjeyW1OCF7SQFVhs2L3ZXA4/JWETeewwSSHptIk0EKaaIEYFgbAAieFUmApWPybEBC5ja9I
OqJEweyRvhsmd/5dHOb2dT7IeE2tUVr+abQ9Ye4ZPt4gh8DO80e2Gt6d57pNx6RqEH3X3g5LImcn
wPFl/sirA6blir28h9bxXKdwLg+E9A/ojGDtBkVFI8hyPLYwh5JHNShMFok91hNJ70AZk1hWvTL3
s/KL48do/PH+kQ2xSxyh9VzAEzKP+49o7Yc+Dqi40wOmfBfGC6BqxlRiGUqI3O1YSSvc1EkztbaZ
0Tunq++YcW/lfreSFl9WtmkH7hC4hbAxmopzghk4dkABXZxlq/svIj6hZye1wtZ6VTwPXgRz+/nz
7Z0997SQuXyBc4IvCAISpIcxIcdMyNkXlx0y0ARpCoZkBz+ZaP+sjciWcRzhPd7QVbZXWC9czqF7
DEcJgwuZsVAPDAfC1yhZ+W2tF96w8sRddPmzAhOmv+Hlr/RhGYUGkP3i3cpfhmaeub0uqhFA0jTH
usIzdb1O9SUINMimPcaBJFaJn3wuYscJoQUgW9eZlbAr8ENSDrbixweGQv4KUh6f9aeGQhecWNKI
y6dUlZe2aG6PYmNsKVewAkSwaK2bBtXOtv8lWxgE4G4DBgLeyFfm6fkKK4KFffXqxOTiZcH97Kcc
hGEhDs7KyP9+MNWCWx64S478E/MFKBR/DaERrAJb5QWl4znIKFIHmYkZePLeHVQ6zgMcFokY0WKm
xdYMSTUs5L0Oc/mRtgB5Q1Club71fA65oDksqdeccfd7+RodP20jHK99PUSYuRbLDyu3IFeOMiYu
fuqNFOj/sw+BljVSTNVDut1PL+f03QWKm84IfE8xTCyPzWo0L8lpG8lNPKt92X90V0WvqUmYAp4i
F2gz/1e0PTQdGppGYcHQzJzCtkHwpUVzQ2WqymQlf6ixnRUMyXoJJTfZSlCyzqlhm+X9Q0GTFw8G
kyV4eCOk8tGnCnMl8FRNbWkReEIv8ySeUwmUV4DHGofCeFUHTrRY9Ktrl8vRUxea92t40gYrA1nk
F+UJK/ktD2e/bQJ3jK5lbc2pA49XiOq64Rl4Ax6Jp/Zoqj6nCFWEUMGgkfZl2VWe+hW05hGoeJW+
mG095y4QuWPSPdaceIvFSrHL5XIFWMEJ0FdvzfUH4cZkA+dmUufLJzTHmjCkQqjN9FRqAR+WPYGk
Wqrezttp5+yfoW8962bzbN1sBoiNLvKB4J1PwvRKoINn67EJytXzKQFKqvhzw9mwRJfG8f1efoNo
CGA5H7MeHgluyy6fcE6sdTmp6Kfzm3AebYYet70ChPF192aLI6SoyZJS3gsAVlvpPY/fTBV5Xvlb
OMjJJn9h6h5/g86YP3k1pAYMudkB6X19Z5pgVuBKVjj7i3bktB436I6YxgGtArZZKv0zRLbJuBsC
pnHgca0EOYNeUNyvuvyw5yB+XonagsEGYUgBRRFEKIL5rOKUFEnr3xh5s/0ph174rs9aj6CHG5Sw
AgW+byZ0TZirqecRlDTNM+pLX9NH90OYljYXtGVM6qjLwUI+6xWW+Gj+slIUOxwrF0U36Xsv2yiF
2D4a9/wx+iy0Li3QWspLT1+ynIOWtLIDOA8u0YAVjYPME16v10iVa070/83A9apXV5Q2YH+WznBb
HM2ldcC1wW06MjTMeWMK0k8rgQhXnkb2CLbQtwdkKNrHcnLCLNHb0FgKUR/Cg80bvlHMxVtdZ/QG
lzb5Q+/rq1ku+GF7/PiYHNASD6I4FH36HC0oWe0zh82uIVKdv0a8CXTnU7VZVklRh5AZsBcANYeI
o9Gd4AbjDxqdn4u2QawfewhpwPsZdGO3J+J28Y9QqYLUnGns/AxuuWhZEB+qfKQ46WRXC5O4nM7i
paBpTvVzYywO+gGpvmgr3fRAukYyKVvdQxR2hkY0sroGCmqNtN1oS9KmJeMFgPRz/0VTofE9V3Li
TaUgOkDkPYPFxsDt3c8FynCTiOCJvfF1oRpY8lO5hXu+IyPmRsAq7m5DaQ6axlAx/7cWvdvIcRCx
/hs6XNPylNjza1+6DFpcC5tlxDn3AruYOXm90HIaVnn8CxpNarH5sW7PPiAXxOj7x28HVov9Y/7F
A+I8OF8t5oC4M9+a1l3RBVL6A9V7R0LCKBJgk5pJ9krNMLzkYHI/gXYOlt9obvWR8qT5/H5uU9PW
j3PTtbLo8t3/VHD5NGiJ1KY6vLVPNr+hLmspe/ALfK7HQwlI71vToVMvoQMrPkLaxVM0xoP2sj0j
8yKuDwI2Cdlq8Y2XXwxaRKTkJpd5bgYRSXitdAwcfBLdFa2veSMlqfB7vv0JRCSAOpQQa/zDgjyZ
5hAVfBvilvBOEqGGa1/wiA/b5O9aymDk4gPH5apbzkbiTW0ow3eVpWbKDqv8ou0pSVzpRg7nsuEY
wz2bw0TAVmgXW4iSkl7h/sEsSXbqQZsmEgFKZ5jgaJRbJ4HAbSf/XUNUHn1LHAzreu1AVoFq2vHV
8TWyaM35HQ00dxTYaqRrcrI1sdlMPwzW3FP54HDN1xcdbJWzVYiHuyMcPS/lGoOj6VyYoyjZ9B+Z
XLuvLXjLtXu77IEk42l770vKlVa4Hv8wzIchBsfZpEB8Ld4/6xGJnNxd8uQFq6ijUgojYT79gaqn
sXFlX+PEL0dz84XEfucdXhxkbuaabqKl/WyMS2FwlJi6JfvDPGkatTJWWAYM6+yvim/jaWds4JL/
0jdtfMur/gm/hgOz6OikPzE+DCw0BocbJ2uywj6RvZpCvg2wVRlpUq7uWOFXPn4fqM2lflzZDb3x
3VQ1X/CwRZihHrT3LxcA27D7FzML2g/HwJLxvAcGlX+BH5HNfCNzOOszyQirCzfGHvFkqcQkrxNG
xk/8gBXU0KjWwxC8uIZmjW8rLGQYIaRSiD9hQGASvoV5bxheNyRiP1kNRLoTABgGqsH8TW2+umOm
hNBOfuVpRXYZTAK3CI/lHR9mqOflYVrvEcmNX+MPQWnw96bn1VlW8wD9KSK9wmWFzTt994vl0z65
VIJpuQwlqnRxoblzN0VCquzEEDdmL8F3kxJGbbk7JlQENIaeK1ACkdDBwe6s2u65okIMHnUO29fu
eW4mPcroSHMCOJe9Z4mNFsdw3uEd2yR2/lbZcams05KcjYuQ4QrFjmijPGEpzboqJMNDL626taQF
y4cm8JusZmrJ9FQdHpr8N0UGbcsyO7t5oCsXwa9zmeuiXtGn/cWGpH/A9N3AUeMWI62pVGLVFmSw
W4RLKFOQ3K+VabDKLaJUtlCt4hp2CMSk95frkDX61x4Ka/JtbRjL5rRWF9X7DdzsYVJw1mMufNsD
5mfdDgECvHEqi+sFsVFFZi57LXPD0wDHaFC9u6yIO4reiA16goOBe0IYxT60Ui4fdzsfndYKq0OJ
jH54VNUf+prCIG2OjNb97xY42tNqQ2vFkgs4mvlqltY9iL31A2SG+ETlxEY7gGOZrx3hhz6KbO9y
NFRMOL3TEpWUqvYqok0O/gKKejXGryVqydfcdYUUfcNsAcXVTAy/xFXf1mOZom1w3nxhryAwqg2F
J+qM43DJ0rmHFoV0vuGuGncNaBMhQ+9rPu2drxOxifK3WgrSM10wYSFaCSN0yBZ7Wf86Fr/lSsEu
YcnuNEfx/riUcH+O8/vqo7s6tVXxQyH0VnSc+gAfQMpQByst/WYRw1ERxzIodUy+xYWjT/VmRWpV
CcCSorjtUetAOkSmTdSZ+hoRAHbU6aezi8MQuoyEeA3v9rz77HQH74f1LWqR/U9XUJDfWu0plHRj
LtSJAM4PgpNH4VMrCe7ygs200E6ruTYORtIy4nudKVgqaEj5M7/GHG3qwzi1eunYzNvp3g8PxWen
FDPBUuar8FrK5TB6DXPTZNhLMeUR46fpTfJjwX2MVr1lO4owQwM9tj/CdoLFiKiquoAkaGNQY9Kb
J1EB+bc/tfD9q/XjlN8umt8ZZ7vyUSsDOK2gQ7NCezs7zGEOAe8iwWcwLFutqUCirqzV4wDc4ui2
a9+0lhVggnFuzDi4FFLk39GcWMvHHGbR9k75z3mEmAjzB03LuilbM5yTNLc1YSI4AUE6Z5ze4KdL
5dEh7+87cprGv0Bt3fsFxWYyPzZ6LnRf2zfXFJsRsbQg7nUII1sv2W2ib8poA7gPgtWcFeY9LyPE
e3zisbbUTnQVXtfA/Y4QmhJI7aSv4j5ybcOCHRSYNnjz6p1INMTcLNkiuwkS/Pzwg9uEkJAkCxYi
clp03r7tPTiXcv0XvzlTXcfuXC0o6NrbL5H93tB+97P2WR7WMPjzU+XOeNbA6ZFgsxdE/3znQBMP
MhR9x0SHoZV+Zfu2TNatn8bf1yXxCi06IW0xQHOj+u7zPDfk+wAe4M4V/+v9uCBhI7ElJh+KxRnk
hbmKmHoqgP9aqUSg67oRSyvPE9oNAkWZQGWZDy+pmzwR3lCxcsfUpnqeAsE2sCgfIj7uybMffgvr
FL5UH8lS9hRbY7BNpM6JOUya5XeqDME57qzEFZvun/CjlmqHyht/qkPYG9Q3aFqoqhsqZNc0Yumr
p5fHmpiYFUAgv9hzV1/Cmimk8kKhbRm1EVP6PlDzlAygmMQD0n3jSfwcnPblUov5hGJZf41UYIZp
8f5yg0P6R+JLbwrifNPhxzTaNYoo28gS8Wl9TGy73PSkuF4baQGku2A06tEwrKVTDGct0JJg2TgY
2+aeJ6LirYt31/So1izEIQZJoifm1IQo4mqNcTbI4AIaoHQE6xqkhaaqsODlo8eplhjqcpTqVRss
d51CBEXcSBNItcPUvvKpnaJf43g+HzOBIvQ+gZLMah8ar6eF2qa1QlQmdSscN/WbJKmPCh5Qq5ij
dBPhd/n85jyWxGZBv7grg/PXgUKbl85yQCPDt0JvkB8wlwKvkJ/XKwp+fGElrzZSacOGDwdlYQBx
/wqvffbU5f0evw3olm6Sf/7hfWsU4NP/d/up/S6Eqv3CheH3GLbOW1WxXmo7Y48smhz1bUcz+auo
8HXKvBYz/q4gAYZVIEZeGPDJ5rS9Y3J5+1RQHZs/pkOWrvt8Qe/gYJb1CZAX16Q/h1ZSZ/unYbAF
+d6KFabtb9iI21d5URPwyyxMeHf4tNUTCCyLUyifXRqV82ko9ZRVZQtxGCzteEeDhHqe0Tin4+gJ
D4InrGxFZpX6RCDtx2d6VSNJpzGCg0AHujXwfwkBoRf5172ydB2z/EANRnPGkSpNAMRr++cGI321
qMgtCyZQ212SZ3TISpg/WvaskHSjVqaiF94dcg1XOtkf8wWBqM4ZapJYfNIi4rCIMK/ap2zMYNmp
pHlZX7WJHFqPhptIdUC/hyhiFofcmcXs05L8f1zkhywYUvT5YpVj7A9hHse/GTH5lhMJ51SlWoJn
YNWnoZGf/fpUDVeuWROGiyegoAFffkdWdQYVlqCcza1JBAiMi2SBzz/nV7FQ67lgMr1ZBtVfgo6M
89QgEIh/Yb7VoIao7mLIm14d5zTh7jQSI+vnwEyiT/SIcxb7JlG3Lp/bGMeKc04L7CvGSDeMZE8j
hZq61Tkt+SEPZSBC/Xaqio3LlZ3tMSzHs/qiIEotRxZEQAgRqzE2+Hi+oLt1mUSGeDBQzwNmrpwB
AzddQPlopEHGJDgB2rjn/a7e32+oFylFZXYICyOeIYXFf21GewAydLFbDGHlyp3/KCggmBdf/sxX
4ttabAqUCYcLW8ObEpHmJ0/oni0ehgYp7PBmq40jy18ghkXV40XCuV9vfO+pPcSNPMeAw5PMMKZn
LMtzTO3c6c5IAI209COcLcH9fSqZToXMr40HF6LlVbjRqsmw7Lxa7qB9J7G9raRycQxo7XVWaHP4
/TOXaELDjUgJktfnBrmeXKHTQomk0EEC17uGqyWdYv/a97bOYOeA9fx7Cv8sGXiKGD3RIJZN+Reg
xkpJZIk92gcTcWY6IgnfXLj+mKicjN6mRZSaOleQ6C6CkVYiLN/3bDAQu6jx029u99scXUDbMav0
5anG23oDS3c6PPM5T8CfUd3c3i1jZ1cDhf9eyRP6k2fEjPr7zjAFvzHpVAQCPXwT0GKJyrZ34dS2
Q8TEJc7ZalK6X5ePUA0zKZCYoqHNbzucPOUV9k1MKb2xU0P+NeknzrwbRJw/eXjqjE4eQlhghqha
F9hcwlqJzl4PLIohkq0nDchItQAePU67J8LQifjonLeTcDvsiFhUQM5G2/mijpTGMUM4IFv5sfbo
Jkx5lAU2ownZ45egD5MD3Q5bWnfqJCZ8WgEmkp7MCq3dovwc73t9jGWSSNzYbZ/acKRkG+tC0yvY
bMfQb54fDXX3v98s12y93lq6ojhTbHRlnzdt+Wt03050Augx8WDg4nwcVPN2bNOqIUZ9RCNLnfJD
6tlv1mUe27VzxyWtzXo9zNK7wtiqdR8FEWlbSAoTXehcCOz3Gjv5YRmY1MlQbD9VJdXPZvmjHP9D
hWcuCMCgv6vUKHqB5d/BEIQWHuLlYrLSwloL4QX/PM8qAzKyrTES5GFeti1C6vqwyRRx1wU2z1hw
FKHyiuD9WpcvFwfzNkYavq2344r4ft0D2dRTn+7paVcnE4hFlJKTWVjPJZCxLtrf1L2DoE5+68L6
jiAZMuokdS0YRyWNmbM8W/l+QX39w6BZIEsdrNNqrWMZ5lGdUBhPAOL5WoYeG6E6L0B50TxkjP7O
KD3i73jCwpUnOXezZkdDi6vDzF/oNrl4rcbUbiyOsVRb8PhGeonFN56Qw78G63J1ZHDypZj6G4lR
3IHMbX11QMSLjYHy6mFUFGVTZDmC9t6ej0Fuxc1dqQ7fFzscJBUaoe0R/QqJYHmFsCTN3PD1gcTw
6ttkPEasHFkiVBe5DasFPOX1B2yqVHkkPQ9OyxHQQNGx2Q6wBrPAAHiFnFLXNsHnn1HFJY7H58bb
CKXY5clYoZAWeQjzFE2F3xT7LpKAPAacPsjm7exiJl98dQSBuEV7xVpiRvDAs2ERQyinD7YzInVn
4uU+1w10wFfwk6Zq34OOMdVEch5RDHM6wdbWvMgSYI6ns9fWEKeIwDgLxJIQYMEe1UbA2L7log+/
yVFgQv2BPetOT5tTFuDdAzhbaCqRzdFyT4LiqLSWVX44kV4zvU5Dz06DrPqowRaTQAMILx3ndM8c
KF6Y+sxsH/tKMdO4op1q2OvMasAFDCqySg2ZDblTp6wL+5FwAy07GdcA0HZZ3xoYgMtxLKYlASMh
OezTO+ho2vZPyRxDvq3RKI3Y01pu1Ss3gtngKGOPKqtnCYlcKfV2DJXt9bRtrRm8uw20xasnwJYN
HGKIVyFAUCfOF69jkt6OF/CtrPu4MTyVU8o23cMLdLanzRzLL2o92LWTSJVmkD9/LiB/4UMGeR7F
FbHFMBrNIOtqJArl/nZunA3A+x4bGNGx3wlXCwrEmDBUbDtl+dBap3Z+DKYB3DrHA58HPSPjdSzV
lb0FHC2E6Tkz39tTmJqVkAJrpnd30UojuK19Juwc+C1MclZAgLZA3abG4AlZGvSfrSox+j6sdlBZ
qqa6YMH0SO+KGLzh2G67PLk+hbLgJ9GXozPBkggUiScY4lTe7OaKREU2QCt007N5zjQ13mYaxXeR
fmztcdoSg1cRC3YHv81N3XlZ8Jw2M4WsA4gt5HKiXW9QtUp3zLFWIFLmBPH5tkyok97wxA7ebfTt
YDmEtA24VTXXMJDZXYHCvZXPjkOM/7tW9ToUobTNzDb/VByx/WaAYttZCPQ4Y4yryr3tR+jAXg9C
8Mq+WDxC1iRRO2rtjv6Vst5yZmiZPmhvRffFv1D/s2hupJZica+ejB4wHe4CWMNLWN26t3TrEeYk
lsXZeIiTJs2n0ge0jrCVb+XZRr9O4W92pAhB1QnxDvoeDG0lNaunTkJoin4hApRJH+q/wrIEcnws
GLllYjZi1+mIdO57TzMsDjFqcYfzS+5vkyetKtQoxSSz92FB+Uc7JqnTvSoA1RC3n8zSS57VtMXt
8u8Ux/PdD2MpeUUxxoknxHQI8iqgSKIEsM49FcCSRisY7q87JKDc0ipRd75MpQL4ZV8ZJpvLsIZb
82ShZIyUP27MBlATSPNE2Psnfbm3MAMUzYlzsBFRaQ9UUv+L5iyJv7IxmlwOE2WQNjalWcSzYsYV
lh295h3KuKUIxrqozYROLMow0iKvDPhFiKi9XfxO7R1pWt8bU/kyL5aOjYZ50/augdKFJ6gVR4fT
U1CH27QWmKj12lg4w1nzmKHJY77+96QRjEhGkyD8AfutxOs8ncmuALC43so4wE1GUUarYb4KJye7
8GroirOnboP1pOf8us2+JB1D8dPDDELfRmIl2aI4uhLEKk7O+6MM+QBRRwD5mEf2bSOmUTeaX90w
MGn+8ypNBlPVgEkZmf1S/gfYN098PB2Fq0QR09GzsZffJuK09bnQvBzjDc/u15iUn9R6aBkam1v9
6Jw3g9FBWTUnO4Ycf0H4YgNhhxH/rhZaBupqE4F65Xg8WAtxOnXRR4uuH/SYWzGowVSe8D5WP9Ll
IJ+oTxV7Ve0GGcXGz1DgOYSZEtBgRQPtvGfVZfZ4rF5b8d6MaXZfB1JashNpOqueXVCf/vIYmGnr
agWarPMNxCl/UDrlto8APBbkdLssWSZyE8Bl2ovJQCeiy6a7aRjaTUc7EWyFYNMrYj+BExySXq+I
E08G43KAaeJlsY5AFQCbLf076mB/IQABhlhxvwhQrlXxhsPwe0bnU6EAKmoPe4B9Ww4aRdFIk5RA
hMNs+bQOnSwSM38UtgXfmroG2hWjibKYgr2f3p5YSdrExQ4UopeVUvK4AKObrjRmYmkCDPr0yUkO
i3PZAgr8QturHLvKLZsIht1irrJ9cU72WAHWofDvl8Wh7PtPwm4XJp5IcEkJrGDEJueIMaWm/Wjl
9RkTzherEv20a5bCVsmbRohx12gXcK5MDDKVjsnErUvst1Th5IhJGoAuiQBu4ICm4CnjVhEBTycf
YjLuqYwcna/IJKDI7EpDU8ajj14Ais6ElOjhuySvg2XjWIvsGmM/WVqNjpFCaCGcr05EWlUj7yd/
Lgdeop6WMXDieQQ6HsmakdXoaIgGCNlk0lRGrx56qZ5H8IvgvBbh5eqdxCmrpeI4hTyHIRuV4oSa
Hx6MYlZNAgyr47bRCYXNC7a4nYoXfvMgrj2NCpoQM/XOiC6beSnGxQr0w0UbTwcAWd1BJGdFMj4y
XdsskEcMR//ihAuIreuK0kuW1udvlmLf7z1feekNGfg5Y/GkFhhofRg7fCyPW4tLS0sVwC1XssK6
aUfCneowSnCM8ad2pFn8IZRSNcCPSGvhn5o2BaK8ik0WzXbmn00jeHpYOn0u/EUtPoxrd/mjs9Dp
Wu7/u3jt4an/zRaxs7/pfkxCPNHVHBWaQauO8bJSVMuSYTz6CVfDlPo5fB8K8LgKoUiO3OGGPwbR
ZMYWPLazBZgh5rmKVFEZwz2g1zH1ICWDL+H6Bz0YxOGH7mFfX/OSDvc/r4hW3zjn+CZSnKSvaiY8
oqilXr1wnBi8QSA7GW8tk4pU8c1oLPXLYOAm/1YYlnKQz/UeocBCILGIw2BXIEMwVyL4Uvzhbpqi
nzpJ3hVm2LikwNBAMNaH9sVPoWgWHD2K99o48i78AfiL0rta9OUuWVpCrExro/L4LroA7S9O+gUW
XOX/CVOFE8GqdZoXu8uWPbs3OjwOiHK61HXzz1l1jsR45ThVHN7jobjhSqFZnmxGuP7CUUCcSnzb
K8ps74/HAsqSOgqePJpm7KerZDUvk3NXc1c/O7/DVNURnNq88atXepcoObOfOGEn65V/S1iTDP5e
YMS7difzZxzBp5e1Zb8kE3QbcvOj/+uP8VKF3c3zKWrrbnQeeTIzaF3tBfk0d6o7jJB/bJnSD3TH
abJYwvXircBe7rrZ/flAPCSatE5Tv1JIzyD3R4mUbFhy3JdiQBt4UvR9gcOqn/jNyHKb+y2NdTzo
4GEZfUOM5sFNOh7smR60cdX7gQYNIR44IPeh3KJoU27LXEdm5PQB46xuZnhGurbEIXLMxNmXw8l8
IShebAwA+KCfI3lOuMmHdC+MWXTrCy0ZzpG+DqCahiKhqMK4HeClz6JBS8qiGMQCv5k2NM132mNP
7KkZyemzFAEhO7VErZwO6IzVnhuuKC42zUQYDG57NmmWQL/NVr8BEWr3AuuAGA/i7oMIYyh4AD7Q
fitchh3s5cePwJ5ua39vFFf3rG3pOaxPREgWjxxkdtdHZIOszsm96RFtK3MVzlVPFCHua+C8wxrG
uMUvmmhcXK/2SedFHXNKshQ8yx85p3wrwzonkq65M4MdvpdhGijJJ/Ou74sSuaCpSgi6JHtEOLY0
1ffx6LNQPIe3k/9/9fB4rfQK6HFWzx3UzV/jHH4iAEQdHGoL+MoCaprrK1LY4PSef0yCRScEn1YU
muFMIadeK0VC/K5+ME/5mAinwYG7YYRLxgHCIl5BZgZ1jXKDmGn8Whoz/ffiVkORZuOIvDUnElm1
rtQ0OtqoDCV4LVQTN5rHA/W21k8eywCKeao5CXu/cNtVjR+9AlNk4/zgCOVxelw3AyFUsVyQU4wk
cnDpJ4JIKcGaWY2HU+v3heLpaCFomwuwumQputZeCC1RXtzhvayMtetKLejYyjBfRJIEWsWhd25F
4mcVpSZewYSTAz25A5+3WfAEkO/NaXzD4yegPsDmscWHjOaUtI5dJ9pbFzYB+9MMibdlcNwYvUFP
ZWfPFD73UUcPpb6a54KeqUi4hE5QxRCMGKaPUNCMCP/DCbJjw4Adb66g+I9PquMHYUQDaNrj2Wlx
ZowYqvZIeKy+sm6lw2z4CXvy9mcnA1g7/SXWyhkZuwYrsNNtX4EJYWH0hLiLKZBBHSeRta9iirmF
SD6/oNqm7AHTaZ7/oQqapYJzvsJTgp0/YLa2Zcfzo08qO/uDFNqWuPkkjxVN4qgIU/+NSKvbv3/E
IL2hg7WrXa5lm8ifrQ2+MeAOTDfmZFp6BQ1htY42MdPuhKnyxAvyd2YVP+T4K8fi1Q+BVvkaEt+s
G/0zkV3a0Mb2nJtMlEHud+mZPeB1uZx1j1ed0y0uM5W/kCkKkpuTfl9/HFkFJ/7Vpi38YZkjS4Av
4Za6pmcuXUo4GoGKqF2gzxBvZXbKks/iUasyWaabi1sjFjcd9xV56YVZ7lmH4IjEFzAqWfV4Ws1v
HpImEt+HyGe+F+z4jtO0hW3RDlAzSjTnqGwB4xUMVkFJWdHxxaQCXsHl79gzaJ6Q2L6Bjs5RFWZV
QUIXBaBDoYZrCu6cL2UoN+ckimU+SdymoIGiX8R+AlVweCGrih5bL0bM55kvJlXlY2BkQlvRxtrD
x4NB9CXx/j8jNrgfJohD4MKYsCPX15/BFE2JuwzAG+pIYZA2wx8CorBf+8+4XqMogp/eXp50MN4y
hx1BmWWdzDw2hZJ/gKDeXxk0qsRhyBORCbLpuEGxgAjh/p2I+U3VaG/rLq1+F3u1EnjCo4NPwyn1
x+lUzvTUuX4OzYE7QLk9wS0FN8G/MFGlKAG1SfH6swrS6ufKQ6U86mUWe4P3eT9d4SfQOg8ByUXz
wwuTkEhmimj8YyFOE2xWWVyvg76hGfdlR2FteKsAknB0qMjxvTR23GdF67bONkfaVMyBWILlXZj1
nPBIqdhUXj3AeoOJF2EMhYojIDErVUkYF95rd2MCyZ7xyU9rD4S2snm6U8kdna/J1lLDN+I3HPqU
kmIJXbWlPQln0uFCwyDJxVWsogKzGc4DXwcnXQS5zVaGa8EkIT2Qgk0oXA4QVF76vW/Bb9qtoFKP
IOMxssE/y0U9OKRUZFz1Pzcay07+Qtk4hgjbwsskS5JjktYDawCJzpKFmwnrV7x5UF8lpJuuZnpo
L04DQbf5NWSD+suLnJHF/0rtipwk8Kn0gQi/64QkXQNV5DiTdcXEqbHqjFK1NBp/eOsN5Yi3c3Ep
NmDukEvpNW9YyP6SZ/FSrq3eQ3SSJjUykmgLhZivdZEj5bCHq68/lEXTlnpvhCg1ozUPkZbS1DZm
S86+7srMmw4RvGTCedMLNoEaoSEmTjpwXGJnW+0xFv8snpy5OU++5U7X11gP89c23/HqvDLtO1G+
Ig2kT1GZXssM/6H0FAXbls1MkEcOFaAVMbKqSBTU0PpbCPcf6pveoHDzRQuCzFEoKH3XrtWa9Ihj
tVUkQURL+VXnPHNNsmd2WYoVtvZRHJs1U6ASilkwMm7sLc9GdzaEUydm9+rAstohBVnT+sOUfkB1
M+PJfieXN7j2Wa2st0UNwh+X5agYu6tmVwq7c2shNviEok4iIOXo5jbSj+J246fV0MSlyRpKpLsV
aneZaTBhmxqUVz5n71pz7Hu3+FJQum8WFuOVjXMI1iSJbV1QzSqZY8881KfAB4Uai/yMxbJm8Cbu
QwMoqg8mG6rOalpRoBLjkgHa91uyH9FUqQZlNYw+DTrPVPEi3fB/6PePI6ghk5XLZHL0K+gJnaG2
j7sJEj7w7Uqf9pKvl5pZLBQCFe836r4S3F1UCpIRELuEHgsFjcjwzyy3T5yhyJrh7U5sQ04SAZaT
kUvNRS4359fkS03CA/kpujwcjqr73kzfbEwpU5TI4W2kC4Bu6QWzHm2OD7I3V7f7JdSXRx4/K9e+
AUscLnUU+KYy2RtlOX3rbqcUADKZuKZ/RHOqX3oaQv2zQB0/QGyl+wkWsjeHCsU4RraJxFClKm3F
lmOD8JF1tSJxm4oJGUmsLv/Yrue/uNaCkyghBVyqQXuoNYANk18pzyX6NvXOeh6gm00FirjY+Pc2
Hpe6RXh/wDXx8BeHdr50otdoJ+2gIn54G1kuJ0e292HyrsTdU3MGmUgsre6kdtMssoYHYVmvTmbc
qhfh0AK3USJUyJrUgWeLMrfcgjgDcWsSYQi4vvQZlF/YDEFLnm+tjgn0cLuYMhNZUHI/QFLsO+sN
dLmeISGmCoja3f9vv0/adW35Fr1FYk7xtHjqPCjGMDNITnNeALJyfRu1UPfOoNsNrPtpIdwAiqQZ
sbO9muYq0IOzkrbzlcXeELxlFqxjkM4BJCMsWNT3oHde5YLmsRTq2NYv2gBEaRYnhvOrifHJCbHj
usRydbsfMfNdJH/4XWQwpgFc8te5rUuZ/4DMzCtAoECa9/Tf40isMCuyCR2Nh7TEOK1V3tabBFnT
Qt38kSkFBw880qYxtRz+9CDubgZ+NSDAk0wz5T6Z+8SwcrYyD9Y27OV119okWZ/3sYG3djiQHMxi
MtWEHKBb6nmtjp7vngerdcrihc67+Zet+i07bwK8NTF92swDCnItxkvUfS4nrfekJo3/E/xNAmhr
s4s3smqKg00KQvnmQ7pe5XqDjxvXuqq0haqtMNlI2NjVQx9rNu76X/YS0nRmrPDyvcFjbfriZnnB
d/4UU49nOcx65Cpl3FS1mVkrZePexL0py5g7I382rq0yHD5h39uTuhupPIZ2AZtd8Hocum7ejtAt
VwlgwctWw0zFnD4Df1qx45xEfZapUixVeIA95mMC5jaqWJMj82lAA8sCEwyZI9V3C339IzwiC0PO
98vS1N7YmxVw1oyVPO2Z2gVP0pWao1BOelAzm997G7FDB4Tlm1jqM3tW6J5jJX8ZYppbTUqBjEBz
4hchBws/viZNa3DU9lK/L4tg1VfufNx49XvVkhz+hZuuMN3bM0y0rYb7ijona4q8UaeJB8O3ASHq
CswtWseewCigPwr+4dC7Oq0WE/Qr+kogOvsurmCdjEIr+9BtWcW2PnVXg378qgfcnIQi9RtkqeAE
2YnextD1ObLvzkqOwYzIvgzoMKHZsK8Gwkr+iy9CQQuTrjLTWBWQkn24+DSCTa/uZzUpg/yQXUtl
3QnTo4ne9flU5v96EMmdqE2xKiibgh8oZvlg5NFAg5/lCHNSWLPY02K6/HaZn7gb3s4LBSDgJ4/5
jh/Q//K7/0khFuSnyHYaksNowmn7ev70qoHpmyvKYXeF4uAQo0gEsMzdJikPgLTp4gAV06z97myF
o4NHd/bUs/Wh5Wsv+1AzNtzfU/Av26pWmhN2I598TvF9dcpBEzzVnZkbGeu0/oVljjKHoorjvNCK
7Bt/CCWk7KD43M8e2gflCewKdkOKB5GqcmUZ38SGVGaBvtyGYXi/reBqsuaY46yOpSV5rWXw/+RY
uMdVQKqjAEHVSnRC6u8M5owbodgjmk7Y/ApOtUcbCTO9QdrdYKAIpQp+FZwnWsCN+HyekNYG5FBL
2TNmKhBmbvm+f2ho9C3kD3uIgFuqBifWhywnrfCQoR5Hg1Eic9Wq8pv5sDn18oRzySUoDjydOvMj
4kDsQbuoFex8+XIwgPpNP4t23A3uHGXyh6dRJbWBVvgwNgW+LtY7bjle5IPtrMSG9LVPK7FEY4y8
CzjrlItE8M7AAkoEaAjV7BgAFRZtc7qKylQiUS2QdPopXSs2StdpQVFQarkYQfJ3mTMzKBdyyT97
kO4LrmPcR28jRleLLqMRTEJ4PFDap8mol8/z/EgxAM6y0/nCGfm1q8c6ThOrOjfaSRJJCPuEfIwd
qBt0kTIPF3KpA+xM5EFL0SRhszc8Bcwl42d9KwpTwf/BIW49H6MZ6CpokEY8E0V8zudVzRQ3khW7
zEULn9wAoCQfy751RZ+zGxerBn3CvdEWx5/bXCoqzc7ARh0NSl/DhPJCetNSfHgXCgzpKdtlBMeW
yCy1DIZykKppQz1x7PYYqLakDojuhdvYZ6zy60bPe54ZLYJTFeEICCunn1vIJ8KAnXEF2eg8KLvb
c61Ljq1BiVV8BvWeDizqBlk5q2hQj0zq9GuZ4f3/tmdifYxIqBt+9iDJ+GWNiDlQ7S+3mAXYJZHx
zFLpM4xSPCE+EeB52bcH/s8aSAcmZELzhjbFCi/uBAdluctE28OoNHAY2L6GcxEvEAN/puZ7BWIz
T/4HQ+vcj3CdtHxEqU9VVSO9NARMNzbRXArz5TSSDLgNnqpxaDgHlTUJyqD1XE7asqLAzQXPKKWV
j8c0pAW7tNDfsl4nHU4n0f6FZwCRV5GYY85Fu9ghnxeYX3HzJAZ5cCA2UNiQrGz5XdOH4/pUTrT3
ChPuvASFkjm8i1d7aPLFM7spCn1I3Wn/rMTRikamtfjujzSUmwE0vtiyzNxv5q9WPb0Spqn0yxz9
IQwDb5ISG92GF667DZAS+TI32HNP8dYZ/P+EVDom2uQFf8QQxr8hho+eAIKzrwhNdCX1++vLfldy
GYZdQwdZX+AJtTdSslKvOcIrT0SYijENPDt4pW7862MkYwGDZjxl0zFwdsNslEA2iloaq+JVt37j
6o3RPY2X/5zKCRAU8KzE0sYXspM48nUfh0XByloyuSRlL+7XPRjGUAc2ovJz6eWiq+PJwd22ZhnY
EhX5OC4VKU+9j0SP0IJMQCYhnlYb6ocnZ3VT8gBUSXBofW4WpsAbn0qJpyDaoxd1Hq08F1lv9QDQ
5QcukMglejC8KD7dG7nLJIL47NIaizgiRb0NVpxc5pkWuRpQy8rzysGWndligf/eL4usV0Ukx3gB
McGUrmJ0UqItnAV74r0zdIRrrhYOh+ugDhBH7eg0ytVE3xzN4d0h4+abdyS/xbOwt7FIcEW+lLXU
NlXOPNb07JwL0xMzqYjA5Jgr75EXVhkHh7J++IS3QIHxYWFF6fXF5pp9MMti4hrRLdJeZb/dGjqQ
1NRmLI9k3tLaLOYjmVNj7deqwU4WrC3yAm0LxvkT746uQMCimO4rtWoYuIgl9h/h+zRdQRvo4GTr
dPdGpr7kzXY92Q/rCNbnHEp8/GHKm4n0uGtG+FLk/QQSnfKi9/nFtdYdmbDZUet6uq9DrXMefBCG
AwdAuzGXTHYN7YoaYymnVWB09AjpYY5vLl1ONTttyAbzYbuk8E35imCKmHa1Jy4TzJx7yfKfuIWf
5ITPVT1xAlKS6qY6RdpdPgsYaNIg6xmcDNe/9Ybf9F1QYaK088Sf4ZVMQyTdZIuyLJS3fl5QFTz6
6vUYOI45uPHH28O3QUSwl4t3o+CtRFV/SX4OGveAA+RDmD0NXiBdM18duLvKMeOz2dzr/7HMctTi
7/hNJMaus0xak2B73h+ONQrDCokLhyb3EDhxB+fN9I2eeGRFitf4F2T2bzWOiRwCo14TdgZrFmFv
2cWmrcOjN63jr84NhguSvFqTjtK6SoeuIdWX7/1BkPaEqyBvH+K4v9d/wdDUtI1v/LzUg8tjpyhT
qntvuKa+Lln02Z7qUCOA7USY7J9jV7o2osm+JzIB4c3a/EdIS6uadjo3Crm8mwT5bwCCnA5oRV5j
AQuIF9hNUROMgclUGd+f8CNRl+D/ihQJeKPji1AmOIraoQ+y70kA7s4zR8dUO9U7FrmlIZb/2HiE
R5VryV0kiAeMHvB35ysNYzJ7aPIrA/DpRbDczisUi4fj5z/9HZC0n2uDzDyMHGOzDiKj3Qwf71Qp
wBc0LnzcjQCXDDCLpaiFsngWEcDSRPpazf14oomIaXzxAvJInHpiK4bXRXJ+5QGY6nua/hW1w+Ir
LqCBPLV+DE0C+wzrQg3DpTOvLp5D0fV19vAPP0qFoHR01LQjQKLgoBGYMpnJkwkHWs7JwUqVuLd6
oZZUxaZFJuDzBny9/z/QT5jE6jeXdQZpkMSMrLJQEBUXsoXsnT/uIMdO8BYs3qxjRtx4RhfJXIlN
p6M84wT3jr2nC0A/n2zVhuYdCrBbj6Aoz5qvYa6DtR4OyTrVO5645GfgDIglGveoPJsRbR79NjKs
mMahlgciLEUZlGSFtIGfd5RKdqSHXB5qOLip+nuJ6IjQToMz367P1frym1jMUiOhsFC+oKPQWNac
oKFp+EDsx2VdH+XNQjYYVdXHtjdQHW6bghAGUXqoGGYuZn0Ml3/YnAfygOnO+uXX3Wg7QIMRMIOT
/YSOLoPSJ5YQX/Zb9g8vQwqDQ0tKVxTBFIia3M/ctA3xnnjeXXmvQaHiCKKMYQwKVV+uAzP7alRU
dWV0DlCPOUrk/P4vmbJauf9UGa8o2NY4c9IYcKP1wBDHVgr28UiE4+7iYky3kHKIQq1AFNqXuQe/
RI6EfWNq4cIOY9j7la33yZxAtaL5iZ2QMUU+cAA/Qz2Xyd4t1UeiXc1gECnkkPG3MsLLpDT4YLCC
0o0YHyqhgxrpcW3MGBhAV6RVJNRwocXGGu/4txYeo8D6jO/ch6CWEq5QM/Mj0lVMqjq8xeMgVTyP
45h5VM5fECZzxZSAb8aKmud4RJoQ5kjGrlkyTS/RQ8taqXQMe5lwWTkyq4bEXsyCsir7nJGeWPRg
P0YU0Y6VtaY6Bkbgfu8cuVAk1vYVslxclfiTMGUrtv8WqzCAX0j4z99CdkTtlrz5g5SDNViTdd0k
9+3EaIBf1LazlyYnPBEjjk9iSuDCi0Ovqh8AklWrmWt+magj+/ztA2AT9S3DxqmO7tchaQDy3S56
b1tV102SW6k+f2F5ZYZPnAZrKmydSIUCqXopltqLLbHZIc8ho1VzsiqMlCErjqH2X989CC218nNI
eGOCTkYQ4zvsJ1V8q1jJafwxAdDbFV2LLNzhy8SP22zQ/Kvpud0jLMWGLqZgXwgiJA5EFR2kZM4j
WiLrA/B3PzU8L2XLjFwCj/veYVX3nlZoXb3y12dsa48G22KTcHn4uAFXM7uKdXsXAXJUGED6NNjf
MKvxJNj8cV4eweJL1bkUkNUqxOLzOZHutoRg3WxR2VHanNvLepg+nOVjRuIrfk5944B3l5YpzJ59
II3W+NgqBd5VLwXlqxC8FQ7E9kAqY3b4CsDQYkajgWrCkQVfIU7EbTA7NpxBKQk6/B8R1ZS/j6TV
fi5xViLvJcr2Okk/T5H00Q/Q1LLUcWpuM1ikl9U4hnddOiARww5u87e1QB1hwye0sxviZutl5mlI
8HvqxPjEfw1+8U3dUfPHG4yUcz2+npyGVvrcInzLVSrdtM4IaF825AT5Msv4bR6pC7jYJ16TyWvb
oVYnOqBnpewDJ81hEfDPrtUoySqIdYKtxIrX6EOb2DkALLMROizbSc54cM0bUt8r6vTU1N0aweiP
PeHw21b5ofwm8rjj6GjFWLV1xkTEJHv9iZlvm0Vh3SnvwRIa7pcpASWNehqTt0a3RR+tQXtvNqSB
vcLCQAtS8VYvvagKQMxDg3YICUfGiYLyvD1edMKkW91Cyse9ojr7ZLfqSz+3zlQhqp9sSu6k53El
HIRzo4eE9syspqUC/VNKlu4ViuUaeJD1quHRcYCm+fFthmjH22KAgg14J6TLJPlUNrBHz+PsDIOr
m30UpSYgkOPf0h+jsTdEmHeJihFdNGZVus8rvif344kxf83Z8r15gNNkf5aSZl9DoO/2ZYWDYYs8
R3Ir7J4LuPyUV8fpAyMFamSUOnbgak/5CEUZJjltdyFxvQueF7R4paCAGm0goAUG2Z6trAAd8dqL
4nwbYAc4X/1pVQQTT2WyiLC2+HLAPkaPcNMHI8+LWAKsl0RHj/w3WeRu2KXanGn3JHgZ9wNuWkyJ
A9dmdkClnzX6aC7wgSSUe9KID6omjicLHRT4vWUSsoqWtHlY7n003dSwPaizELnjjJpkfvYHDek2
A7mQ5Gu/rEPQcrNXyEUy0viwRL4mpf3Hzsx88aO6CDf7YQIP58YJoLSaaILCt+dual0sHJZjxYIP
uutck+uioxT1aZZ0ovUpJCBaJeTTLoKMq8yAeSVnkRhObjDxbBAzf645zYYW8M5b91MDfBZF9pzs
7VxgWlI7z9HmkV5ay/JGOZ0nQEYyK/K3xRFX6gci6khJim+rXUAFPBquUNbXyq7L2P+TsCxwR4/a
GAsZ/MZJdC2W1/RbXw88cFbeIshNR0z7stUFjjY03N4b15ls9WLF4z0YrsXrheVhEuCoXCmeYD1O
uV9RsocDPhBcktQnWa7rOMZ2SxUqBhmT/o1SZlbdJ9WX2kcy6LhvVfo3Ojwbgy6dtwgZeFp4JAD/
KY5INIqAo1GzNzjzREePQsqTwbcA84y9OGYIHdbdBheDY50Puz8VfLkSIdFoLKDRpUlkIMUaY7U2
UPNlavVuuPcyKgjb5qRU6TPG91VCS7PHdiCq1qHnBdxWPpSeW5F+UX3mdXdyIRoQ9VT96+sZw/lA
lqfwmxQfEcq7QdpOUg+s+Qxp1XYLw57Vc+b2tfohsY7nXas2Jg8WGURNVufT2d5EBs1pcpaEwrh0
xflegHrs+BmfMY6XSZSW6kTqPD0qQj6ni4EwYBkdFojrhLkkE8BUWosuhktaXpp4BKaep7xxs03m
KJsc7+sRFza8F7eoP7qqv3f9WWjRS/aAtrxxiD7/NakohjViLHBiYHBkDsN9gTFhoqqIvp6vsul1
mo45EyDquRaU8lY6urHkDLPp2B3S6Iky9uazzaQEWvdXEtdTnJFfteWST/4hK6dzvlubhFuZqIVi
2i9Y7/FN1Zbma5TuJZhCCthuPe84Bdkt2ZX4/bOLQgkKzoD+zKMFWES2opbLGTFShNFITc5PAlrK
uxVBeADz4dpoCvZvYDE6wY0a4RfhIJjxRE+0I5w2T3CrVUuFJGIxnQ76x1VU2bhTePeW2Xrr5YWl
zzfU80dOvYGfVAdRzWAgY1BLVYJZJVXWz2GDB6yyAIwS0NgSeVpS/DjPwJPUHFuv/zGRMCtp34qT
qpqstzNjjTpT//puva3iDIuC7EuurkQcB4H2qWCY0kyzMTl0KeDDQL3Crwb+E+LQWaGaFBKkEDDn
sCHlE3m+2XlgvejCxAOcIyLYK4EbtOJ53cI3PN0UfjigZmJ3XRwavRT6pbYWivirtgtx0cPvGUQW
yrh9aBgEDmXgbaOFkJuDtlSWMOqHIgzxiYtpZcZxKSFJrZCCel9YRNQ5e6P7W7Gh3kFNA5gKO4zY
ayBhk+BHPdzw0ZKhtBd27E0R9/R83TsBhPJubqwAoTHkEo5XHg0Dlq82Ha1BB9yX9xBvP5YKmu+N
5EBer4Dc3vyp3/96LbdCLu2+B67D0ydmV6xG0x8iGoNda7R1UZJ9FxHS5TGN5VkL45C/ETyausUZ
EAiSwTLTAyIvGbbd6honlEc5HeaY1Kh1xdHWEkzrdRSQ7sFFz2aT9rVHEwI85W6khucTZppZAT5Q
juhp6gVGxoHwrFuNWFRAOUG83ilrOBi+w0NoCOg6VKC3hs7Wpt8vprX7ovTHxaQgr618/RkSDmba
v4THot7hxgwnbZ6rWiQvrjMRQA/AWts+C6ihIDIcZKCHUu0gg0UPZrSv9O/1B66Rp+EhnVWOScCT
b3a+qAOBJ2eA+edKfGaKtoiAYuJ8At2szlh+kft23AkeOD+i8E0xWVa9l8xPb4SH+GGbzLd+/HuM
LW3yWEq3KjYZSzhbpnpSlQ/3ObJvkrHBxOMexPWaCrnrt1W/HGk28WKLYbyavhzM3NVQLait5uNp
NHyhQPg/95COG06wjPe2xixDx/Ob3XlJ9iPW4UtleM9bYN31h9liljE3mg64HABjzGwF07HSaZlX
8l6qyqRWIjdOIP1BdbeRhZLh/vi7/ZCeAKaBknZf4pkaRGSQBxTyut4yG41GmnrASty1DCQ0fK1j
BVAC1z9qPg92Eed2/n/s19MccdYzZo74KZ1t6Muh5+cXfuzIA5BOV7v61kZM1XvILlnLyF+kxx07
V5OIWHvQuVhMQW8T/q8JEwRHQhhZjwXAH6SnpviNaqpWrp5n3Kmq9DiAjSZf3vmjJbdR4S7u9kZ0
87m/tE+4hpaepyr0Hhoh2K/vyX5fqcMp3DDGF5WkX1vJqBznsNB4tuToRG8bXt8XeMGl+4O7P7xT
QYcXqRIvlWiVycBWXlJoqXzPobvPFk7AmL2VYsgwtwbhwTsqFiyFUx+pMsPF8jS9XxCb+vCJMUaD
xjJAEPe/r7FgxlzuQGfdwKE7JhfoGuk5qe/CiM0EUPlixO45WeohBeVNKeplOIX1C4gvteAeT4el
wsaUvm1tLa48DKzR3GUaxiBMGNLZJITj+iyocPpno309RHqnBsccdaFFUYlN2OUwnYA8a8CEuuOb
P01qeslpnX5Ce7gwrestMR88rDq9Vv9Yk6f7gh/yoe2uPQtnicVTgzl82Las7GZ8+8g7HAdzHuME
O7bJmfwNHVsXJygXz148Aa8IsZt+L814TtGFXWxoqptmy1dsaJ7jXhM/TYwd+gTh/RDZc0FOrlRr
E0Pzr62mSo1Z5V8QuzGlgCYPZIBawq1mxOPxOE5go20UMKvDLET72DDtwTcAQlRVOj16d6izg8aJ
tMi25JYz8DD+A0L3ZDuNqUVnUcGRlBXWxEJ+fAEVs/i0nUEmWI7tiq/+lTdEdEN0tmNfDVngiSwL
zVUWYto0iBRpIukfNp+7dxxyWNC3tkNTFX7Y7FRPojqgoHQ438pu6bX6U+rGbMYim4IO9irmt1gu
YiQ6pVQXfs+Yb1/4eiqD53oEgvTyhk0tK5WBB092pOzQLDodRIMzdZFqjlPGKDDGhYZuI18qO/C2
9peul+Lw+P6U8B4XLopSEwkxlWDD4jGldzkefNNPSv7XYeEK4r0Y6EOpog8IKBEzdPjzRuF6OOTj
znz8aYTC0sWXJsPP1rSUbkblK+teKgqMZHm7WH7mKRzMTeqGgTkSD3bevNb0N7Q+HOMCmNofRW+9
0I180bZf2Yp3n/DWWwWrvx1Z6+aeQy4dQrIW06qzmLBfTt/ep3I1BKB0plxbAXipiQz9ouVo9ESP
ksPolvqwjJHgVfdhGfUDbhF8DimZ4+tQ11Y9QnBpFmwlo8VY4gA1c+463jRgf5mEpx22IcN9G2Bp
LipVYElx70Vbrcoiv/yKCgUWAJ4MIeG9X5bKypCC2qH7DbsZbGLEI2dyn2Xf3+vBla/o3W79Arph
Bz0PCOdJfptnDquaLojgrlUuXN/o+9wW1b5I//xqlNf8Aun3JwskKX5IPRQawtOHAd4U/Xz+0Nib
8eHCOuhn6oyU/A4ptqg/7gMtysB8ypOGcPuaI+WEZF0vPN244DkFGZ4j/G/Sl+LS9jGxV6FCkRdn
QTt2avpSRdtxos7syc8txM1lHz4NXAvrgmiUH1lsscYRB/3YdgLwIJLb9ZteUZr0PSV4ImWDGSxW
FX7T7gABUXUYFOgP5uzI3lddgX0wT9gbOa8SsN7nqGPJNaoE1U84ToXwaPULjSEiLWYwUnz01/jb
JzQ1n0ssEsm5EHztXHMxEgwW2Src8z7ZEO/oPw6nVdy+ysC1kpbyxjEsFnHT7p3rZ+7bgQDNSuEa
7tWrvoqOr+L3JNWQNRyViKuMvPIUGxRH4dCs9dwTYkqU6knFQzi7HO3armuosqe5Hv25ti/FlsnR
c8/LsDgh1EH3xqp+jzrw6K0/MljbsbBNOIKneS3+rlQnOJHQGtgv8Lt+oETWjFKQbuTWW03gAaKJ
A1ccn6jbAKERLydaWd/BMO+MkxVmwMNSDmSlD4XS2XxlltCOzZJ0qgQL6nIqAjx3vBYDVDgqKy1N
xIXeos7AyKrdCTzaU+LI5kB3C9kkAXzm+YsSp2Gclca/VTUhcFt2aUmvqYE38OPZLFKZ8cDm3X4p
87tB7J2L3uR+9XNiBWMbIy+cGmzzmB7qskm0W9RvAnPmawxpzRHRw6ZqxoOk05g/UWw+mGBv0wMZ
Xkdn4CMaw+j9kdpDM5RNFkZBsitKx+UBAtE2YJtlraX3OvJPlWvSNsmcfHu/YQRMqcAh7kMa8gC2
W9EF/Rep1+22lbF7p8DvDUWL1gW0Wwb7LpahahUwXBXpU7DfKr+sixpx0cw6X3qLwFcStIYBqJ9f
MZhfXj8a5eil9rb0MHRLSBiXPT7VDJtWrcxawueA766pw+FaHKSyDVNPq8EDEOcaauI7yG15tXlP
IGFYR1DfBkK1k3B+XNeRycqoP3uO/6e7uuWFOy6gk6bAo72ZW2HmJcjs3hDbRLrvJUvIugXnYkvI
jdjS9huBFxYtigkOmvUmiVTfetjnyQdlS6tXyHvxwN/Xbkvb3iZv3gxcEU9RTBiWShhAAL0gyhS7
BImWykk9LwGTyBzZ5sfpJdhEihg7XSoFp1QxXoJiDgk/TjvWX4thlCE7iDxRn/fBhrf1oc9fYG7z
oF3XV9A7gidAGh6yCCd7DgNLfJZflAsjexkusjXytsuymvVECSl07eSbWgke4HzgclKOD2NRW6jn
aWYwA+YASHR3rqgmFacrbnQK3GVe/Aic5V/YK39JxoJlQYUDsjSreSp7gn+ENF0XS/X9cUY2Q5Yz
QIDdQNbKXRWKLCy0r2JV75e0fCKhQpfda9XB0ehsAjs6vazt06d9xRI1sjFHssM7chYas7MuclRv
YCP4DMzhTCqENj5Fj/phXHK80wPepDGiKXIdqzAbJWa4lH6Wm/+luhRmvPLM2U6VermO979TGy8q
INcl5eVbK5B4LNAV269bU2cGkNEkdQMAYrijVf2tJsAj7mZ8J+mHr4j8O3vDGut0zCztB5eSwZWM
4qdEmAjpuGh+glnf+5fpc8iqGia4KFxr9qhhv03jr5/UgOaR71nXxfmOofJ22+H6Y40k3Ek/HQdW
ctQunrtjjlp/QkZGFLCxlH6jQ5hKaYRQntAmsJzPsexbsr7gLSo86O3/jxs6sHB9cVDgJ5axiITl
0rBlHiPgP5GPv7Vko3PGk4MZZ+xad8JgW8txd1wGwtZ3f8hiH3FDnVck6lNYj4UTYX2r9XvQXMpN
+199M45Z5iZlEiCbDmNqzRccpmXp0b4lzGDuwtpU0tkNwXwDcUHYZkKQm6v/6RM+MUjhu9YdoPZz
cf6ejOkZCgRKnHm4jD80s/O3rU41GPt2ESHJnfa04nsU9l5W+uAAfdY04mJ5MXEaweBswhIsoSYS
nNNMejaHdF3x0IhYkJo/UrEu8HSsKwnG1OaiqlMVZnIs+6upwiiDxEklvHpgNuu/ynkEe4MhJz9P
KYdSmiBP3ZJQiIUC7TrVkstCinxAZnuKHj0R7ZxLzOwxqpuNR+frLyjylbetFCsP5lkC4ccNCTMD
C8SUnogDO+bW191qBu7kio+mDKqnbw+DiKTdFPDAORl7hIAsutaZCm624+W9KHdY5xMC2VsPqhlO
fkVZPHSvTPG1cQ5RcSk5XUCSv88vLl+UCjrjJcc5jbaZT79zAsLVtdfV4l3Bv6rHMQbFgq40eAQZ
S+9L3U3VyFO9VzaT4uGg876MeQsjnMi+6J2fd2n06jA/w4YU1vGCroSiCNoLNnAV6KbGAPHFAnnq
7FfL01yb1v6ejsVrKDksDn6NmvciEfTSJf+wrEyuBqJRUnZtJ6Zh2SMiH8mzmKwvPaypEitSqWIz
dV4R3yc4NtkUnfDkdK9lLfWftRIQ66UIqkS/03I5wAWz17GC7VhqzUS3NW8EXoZL5aOEVnyWhwX6
iOUSXcz0gXXTkm2gTiJoTocyisol1NFye3frT6Aqi/Gc6THkbAkzOfFfbQZtoOJKkkbXU0kwhzLt
O4WFDsVpacj2LsxtCivIz91N+Eeus3ZBJwkuYj1P6rr/WzXJ9fxj+x//UVbhYyFNMMCtYOMzV0gC
Tfugl2HB97Vibg5HsGKQt7XK9vVh/x9TdG22jDjDhQ0U2+bSrwc/Fmx2f0ID7lkb2+aoEoAMd23j
SZQJ8hJljspjrZY77Zrj5pokmBZil8quRyMx/Tg0wAHMq6w9mFjfxca6imQeJzT5O+ZB73Q9AHBf
CNGZG5hxUnsrFAs4o3twjctgfmLWdpOTfKP2LTXR04MXpyZStpAXH+hDRVItaFjMftDUpxdv0xwb
VaTNKebmlA9TC8C57cZLSkiIuNhvVCqGXlnJ+qzoiaR/GOR97nh4u1i4wzuDdJA2WTwcgl4K3ynJ
yDgmF15H/kK0bbX71K6tN52MijZPXGYO9H5n6bHMQepTJ+bu8E66XVVUm+ukgMHi9BhbySk2nzUp
x2qAop63SUB6n3QI6dbZC+HzzoB1H4WkI+N92pQ1y8MZ+p2+KU6eBIrLGLIxM/7tkwVY2k9F+6cP
QPjaGRhokH2f+OAjlBiQs4MtqM2SYm+y8dZe1SJHHXoTk8F0q4USlalqm9WKz8f+y+xct6vcyFR7
12+aN343C4zGudDlmGKUaSxgMow5wD+5WHkijuTQSz0Lwjrj82uIhw8nANneQ9jbdxHFqBZ7uiqS
z7Kb+czZmSRkFwqGkpexGnf0WSiGqdLQaECZakdcmkPzpUv+e01lqqTG/xWzedeBKtk0zawwcOjE
v422ugeLYS0c86lU1dPzCkK4LZfUrX4XOXhBr9eC4Jpmw+7aHdXcw2pESEVBvX9peRXu39UboKzA
iavU6fOFzM9vokTMZ3Pt5BmlmLckgPwc+Owl3UgG0w9mcPmWLOnCNOQ+HcvSdAxmZ5yg1HzNl6yX
CTpSruVKlh1uO8dyOlEIx/4EotB8ObAPREc0lGHF+OstLp4iUD6lRAA/Lhmxoe97qZ7cEoXfn57p
DgiVy8SFUqXS5VvkLxnytmkv+EFYNTOxEySm+NUAGTMXyigXMegTyZ/OCHEveIgi3dk5Sreu448P
3aDM7xqO8JTDuYxJQQYC4/ZvsdGb9CaliY3kOCdojLD7u3JGPuSFhEpeyq5RoMO7raSC2aesnaJo
X8szEC8S/Ftx2VC2RR16Bc6A0f50HbnWSYnW6bLb/krmxEonclr4GRmxmrAGm1JiZ4/z6tSOF71u
xq0JVdOk7HIY7s88zbsG0X4EI6S6xX4l8NpkcJSxT9R03FezvQBMt3hH/VbbL3bq7eohL9pKiYFS
nzFSV89lbdVvEoUXd2RQXuLE7zB9wfN3c5nnsx0PYD7wrBHY6tSi4MzKnD4ZSo1A8eVKK8yLM3IG
x/D8y9tyxxBpCkdQR8DgzZLjlhonTuP5JFYGjb4xWvjxDDVVz1x/JePtquO5SB/n3xQ3hOWSeXmz
VzXM3Ims5SZoMWDAx9+0Nzv2H/KBJd4fVH5yEZ771BuQJhXjFPX9ELKW3QSOCZsH6JcUVwYe1ag/
NBH36Ss8tptXUDmHEbIfmCeDi5N7+sOH9TAx9Y/DJObhVAlGF/CMYjDDwO5+f6vNSFF1NO9E1npw
6cUR3BrrVpkcXtiAlbwg03OzAVRrws0gCzAS1ZPQ6dOFnk/H2qC4Qf+mJDcABIrlpLZ3vjpFBGa3
I1bkC2PnYnh5nWy8m8c9bvf6cKadXwQI3GB3+GvCaaFJ3Fk/7wPrq+bE0vCkAvmZ6TaAdR6aE7mY
FpmPp0m6RcoTpJCWayGKa0D0hpZxgEfg15913WO6sNHJZENwrw60oKRpSTvmfHxWAe/Ajs9CCiro
pSwZYL4c9ETXb0XBsAXcd0YfSAHqfqwHb/wh++UpFLE3tDZBB33NU5ztwkPepJfSClJZqslVWAIW
DUOUnHZYBMeScFPmf5YSJfKvfmJsnBEPUrsidq/zm/sQ2BoWv7Aju+c1j97t3kcs+lmFrEYZcJyI
FQ/G5uT9bpOsc7ukkWijtJtzq+fij7IjNs74AjgAgf7sjD9oCBhXXSiWnRoIHP8pIncQt0xdcKkl
ujSzRqju8DL1w+i4kwFUT+MpaozRrrbgI1MZfwFT5jPFpVyyYippUzMqtQv5tnSQCxiljCuPo1qE
p1PTkFWj1J/XnD6DA4k0ZeXtcfhDZGeseczFvQNQ4QcRV9H4XA2TtQmo1+OvqbRqAS/ID9ToRNOt
mW8zuGJ3cRVh73dsh6sFkSGo/Q9lorF1DnupDICaRvMNOhy0a/wSthMlO4W6sfSI8kGAKM+5/mt9
bekHwpJzWt+pczmYtftQsr4vwCBXS0arwm6k8sONvcCE/b+vPZ7msKnwqilKFKkEwbg33Wqs9ZuR
hiww6WssQsWsSGeACoDbuuq8IKjl2jcMgzikCR8Jg1tyDdiwQHRU/EMNMnFh3Cp7ebH1Jv59f6+Z
l0gd9ivi9YDtwhBCAwQm6ViAsOGR+cOtVhKqPqkhEIMbMaWGBH6BjJBHcK4NXUyatF8aRpFOxnXX
n2qFfNWq6XwOoxnKtKAB8g7ryHlHCdmtZljKLHkkhVZYh9DHeucx6N7eqC5mUXBzPSYW3642JKyg
qfEQQ+TjW8n+9ci8W8klnu3cDPo/POE6FewXez0Kax41LpvCMbP95r/P/lhDKgguJ8+GgtVU0tnh
lkIHjLuarbIpC7Gvs1duOWmzVReH7ATBTLH7uatAwzdz/2R60ex226Uk4H6Anrx0HmBlAbUmKiAO
lSfbGIpNHPe9/63et7FhoIIj56MrA+en+D7yOCvEK/3PHPUL3zx1KYb9jyFvLI1O3ok6Qpw7ENe3
bPrR/qtzbHbFK7SUy0j4td7ltQVOSmx4KRJYUjuB9yJ0xBSe7uyLPT4vdho+LWDv/V/MUKsaKc3t
2wbyBCOj8moJ6siYssWiCVdCPydmsq6okWIS3RiyRM6BO3OFW5JAgs47sorL1WdUnzhlBLOQqc1U
ZoCJQlKYrD3HAuMnTCJzP/p4z4dMXGznNSOrqZN45H8wPTE1f2nIQ+P2b9jjoaevMjlKXO8c18Wk
INjoSO/X4/O+X+6PeF3DNG4i1+nntom9iErGvbRr2zZdKdjCZvDOV9N7xqyKbgVFyX/5UPj6pA0R
FkAAiSpHi/WGuskI2QzVbQuQRTnmuzscbTVvaGTJdNhUMntoqIlTMHo6dsm72581PGOpJYPbffC5
WRstpE5nm2hs09xYOEBnIpqbhInlELfkvBlL0EncVilzJ3JX/X4lLlKzWKzK8pZJG3XOP6zXWqPm
VA4CNWlflkGMyIB1ml7QPHxGCmERbJgQv6Ge+VB+co5Jp6c7YWshxgrJIzN4/VZzYpIKCLcdHVK9
JiAk4VbvecJhtjEyK3uP5Q6k9rnpkqZnWQBxTypdNuXP8TUjMQ1FkzxcxgNd5uev8WGfTRqRUmC2
gMqAsV0/an4pKaAJQTtjDYLqGEP397BjIDLwCArJXrYjJz/1Q7bjWgBMDPL1GRfQ8W0q7B4cI9q1
yzIyUAj2pWZhtlIQLl8ijwTyv5GuS/LA4HzYkA9GnF7RPgbhAPgBPoO5I30AQitkTgLjFe+xzjDo
RkCZ0Ts5kPV5L0feUbEhvolNuYzl1vc90pw9LE9+8elNRlAGHY0iz+oG1/+WfDMZHeuwJCPy+0CK
0z19rhpU3h8Gvk4UX0axlbhGhJUcEey4dXIP5pvt+NM6Rx4mqxcAMwHgWC7yRmF4AgptZxr02tox
uneh1lu3eF0UROSWMRCP6DKKlm/vdlvVvsRXQq51T1BBG3Qx7MEoCkChsO61GvQSUbiYi8TX2urh
tI3rkHvp93UvCC1qAeYkxR5R+kT0Iw2YueBIOPIdPpOel0bl6F4QhHK0ybbv0vBAgxCwONtU0VTg
bTyQ3XDE6kqCA82Q11BWywkizYDYvc6knNZf47QblyifIXefiuxs5bj6QydGzl90SRPXuGfe1ckU
fM27t+FaqbtthyOVx7lsx1S9+bIg6TEkZkAmJPlCz51JLKYXGafG0l2GFdoPcmm109H0S2iiBdFc
8797ERyND60vBY9Sb/V/FGzrQSVQDtHOdj8UttrfB4Twu6ujDFy/BjM2Ekih7KBDcu0RbYHNCtjQ
tEg2aTwD/8Mg26Rq+3hs5+YFc/liMmA9WZE9hnVacMAlMG4EIZfRj+fHktQ8+RPV4jNcAcXlNBnv
s/qsXS+booo9i1F+N2iGPWKmRjGV9cDka4TKnjypCsZntdYenavrzYvbRFM6rzP7ba/6mBNQsSqa
p7/XbF4gVFgm2hmW6eYyj1XQYSD7EMIdtczd2e4jFtHL7hG55f8xf9/l79yfJTbc+EWcF3fsDAaW
LSFHZ2gnHUAs1Ami16U8UTwOpKtHyYhBlURWOk5azk4Tx9tyxtXajw1u9io7gnD89zsvINxX2fi8
TM+pz3c8NcIHuaZ2rOrT3rg3tqvEzVTmo9N9S/TLenSBGF2WfefN97riSSQxpMpPeyhRDqK0VKNy
KkA1KPcYOv9me4K7ubVonNgDm9+aGTygnoIqmJXVOtR2IgoyydMQYTaTI5CFpZzP7E4Cb+3L7PuK
8jmqxySxrw4t4IsrjcedAxKVvdVpa8AoE8OvheBLfxG30FKCsVt9l+6ns5tgSBGhysngDKTzR+oS
Bkj7KTYrwSYgeUQJwXSdfd3B6Xs/+9IvoBiR6iHuVH4AHgo3ibEjPQaqUj6RO2ZxxvTRP9TShHJs
+PeFbnbugcJBiTx3lflXrnrxBxONkRmPWsEX3sEbYCC0AbPRKmzrgQ6Wed0jiWU2Eg0+oopG0ol+
vHhzMY5Mqzb56+TbLqnu2dn0nBuEt29i5PROWlsbD9rNIO8JtVS59Q6kweKmdkUdzzyyOhZMFDTz
0j5xgiP5vgADDyCTozoPnBGMPawP7eRmuXL/RiCiiXoJCR/RhpQTaz5gb4SgbVzbX4QMwXCIcjgC
R0lpRP52UWW++a7a7tuuD4VulgvjLnzrukybIaxicrkw6u7XV08JWAUDXRmIU68Zc5DIaSfTBnHh
wVYUpEvuKPH8x+KK/JUvfOcmizKUvQdhQMvexjVN1U2kSgkoQocp1xH2DRw4Hj/SFubL4zwbCHAD
VRZuO0cCllzSAMgzlbBhz0gqd4CJQqMmvtlhgLPeliD9V64pwqm9Dw1u7OzUewM/FwpCYbtqEsam
6y1GkbO+NONO0zgpNi+z8E/6kJ+ee2szx1rTi3Dgvo6xyUmhWWUjPfQVAa8yi+6b+IDh/enMCHuD
oKJ64uf5XiYRRAkzxBnBUhOTD/S6douOSrV0tqH+4JcPv9gXPjTAWX2vSh613QHqXeF27rgdPEVu
MjffT1TUdNINfkgcymXRgDaUCPsBPTJ3nX5OPhRKqvr+mpodM7IdL1qXXw+dx7HKNkEdPXp3mJDd
w3wVD5fE3x/4CjH33LvoYv/WmzUeon1gNvjzjnzAWzO/4/CkU/TrTLL/TmUVQWqX7oUj0SaHpNLN
FnRBlNLIWA3A+nBgrKPe6CQAABbCzmi1Gwl/VxrdMTRkvz1zIvWtZRTc8R30cHptz3dhpSLWouSh
PkmUWvcEuVu4xtq1/AbqkfAkrVrodY+73c8q/pI+Z5GECWiHU8A+eMz6DwFY3WOq95Pxg2V/bBde
WaYTswOx8TUQN58coxO9tmVxWr/V11FcfYANJ9yWRzYJd1YyYPXeJIA4/2VQl9MSRZ1d5uu56U+P
F+jBy/u0SPQIkhmg5wm4xFIX6FVGtBJbkfqIVO5cxcNQ31DRDfyObNezq2eoe+cm98RsGCsq6ABf
15TwXtpCBDnGn24n2I8Csmrlh9/y7JzUN9c7jIsm2pbpZGQwb6sqtNuDCTW0q7NOtI61va+Xp+Zc
AwKZH4TDhJkKWSYRbrtWQkYwL+avKjDg4F44evNznPRgqx5Uqe23Xwk2kbA3aGwVAojPHDmXJyz0
T3lfmiJwYkgVXUnLwHnv4jOQFC7vh+k71ldgr+BNDZRKHpX2PrrlcsdaDKm5DOkJIb3RD5bOOe7U
xXJ/H/YA+sSmgXQOB/2QGhgbu0E8P1ytrl2VPIsSTF0secEuZHn6mG3dOizv3YpwYQAya6S3kBAl
VyvqOyfHnih4CKPmIsYpUz+ERl0JLoR0VMUH71vdRdz4qCkCuSPwCYszNDeXP9PKB+VMgXqlnUYt
wnOBempyGcJBdqjUE2pawpwsBrVTKmOki4LoRmdBym+DCaInKCzixYJxRd3Q9OIwadVnvQW7T2wL
aAyOuyu57iu9+GQVynfTxFx29kclOtwFrVxcn9lNIKtW4y7BlRIUiCA5DsxlswEPcEXTLKelVHaX
8vxk4m+LOLQztoCFogif7gv15XCYSQW12CVe5dwcIdARCto2ej33GOqjXFrRpa9Ws3P3G1QrunVp
8pcn+op4H0UzOpGCKEFbnemPVeEFL0oQx+SvTDYPp0JHLCWVF51dc/Cu8XeGvvgUx+Js8X9R/skp
QDfgNJoRIJOCU6QRtLmyfZXCMN7C99nl8omkDNF+8sEXhpM1aVXnz71NTtZA9cYPE2Nxka6TfUn+
yg/AnL3F79XOW0nK+sgKrRDSWmXJkqTRSvI7AGEwHxUYbYb1s+tN9+YoluOttoqlYrcNarnEKmac
1ZOeKcRfvz0aPagsgmte5gesjvghvHsoZQaxnFdcp9AzUoUZRNNWoU+woNKyWbo+2ORTjQfy6kAC
F+QyLlHxZwX8pjM9qBQtn8YVp8nI1BGJTzazFCX+3E93t8W6d0lTsbVFc6yL40J0bDKyeK4ZIHUp
WZXWRJ/ZQfkcGUVwCeIPjHAQIL4MXwNUAGJqFB1POuVtN2ZgUSwBM0NwVt01oi2hcd9MS63shE4L
4SDNhgyzzwTV4a8thIL7qAI4yFZ50355pFrZX7GmaWiCzyBiMKXuPGxcT274Ca9Jma/D3IPWljmB
uupE7Mt30vg+q3aLdkfZyFq0tIKfQggXLZdBT6pFIs/yM5VLC+23CEp2GDjbj+TQE2hDDiBoWDja
ImLuBJj1VXWCFluGtRAU8MFR9/zqiw5zRt76KAkgSbts+2XxUuP3XJMDhUwPYzIBgEN/c6MVe4/D
U0RyBk1IdL5iAYBbtAXuzCz4TJduhauU0ROvjCczxR6mM4eMO7kga3Wibtz1r7XKyqW4i9hlt2zj
5mMFe+Ta7x2n/bGsODckaaa8pOCtlF4pRflidFRP2JzVc1t23y+auEgVrwV0RrsUYXyFO0DWZ/FG
L7mtCvCMwB0P2UMuvIFLewvTVt35Uxfaksn90QKnEHd1pwImtwDjvmWBGm2YaneaTq7kcsg0XY+0
iVgcoxua2IQcT/0xmA+s3Xa4JSZu3KPFwVM9VCo/BNrQ+Fz3yN8D9fbYNgEblRcl8IGyfLtkURfw
mPiwunUL2WLDEXsm0nCP6YWjPv0wW6/mKNC90fvB0+O3+7JR7aKg8cc5R9fwjKwar1yH7aCBKpz+
tCK655caYiX6a2s+JvpwI5tvDW9B4g8FwLoQ4h7Jbku8g5propDuHMftcriEIi3IP/993LOgpLwJ
KXh0uoNc0GDSlI25aNEY8zTpVqv1fQ2N3LfWA0EP4gSKi9NjcecSzGVOWSCORF8QJYwiSlRTqmuB
7Y4p8mE7fOL1+yMoBjSaH8vHh6gpMTqeuC9KxG22t35wlkKL8NkM0hiCbeDr448CSrLNvXibhugT
D3YuVL/5Id3MInELKoDOqOBHV22njFHTYlV7YY6UPe9Vo3lF6mWnOXOTbxE+6lqad8IK+R2gBQXe
OE6IYDlRt30Gih8rmDugCzNnYnz5wWCQCBdhuGuWRSktlOm8oOcef6ApqDsUBmU6s9O5+EBw4+26
V9AnppMABAGR90dB6mmu31kgFlzb6gxHVbQoZZ07N5LwyZAygy3M0j8YDNe1jbkFl84LaRbpkudY
Qt7zGXPGEP6oggtaeyYxJzx9g7ZlK0N1CVGmeFofODcsrhwMICr1T8dcQy+f6gWjGWGVljZ0OHTz
Wb74ZD2X4oU92gFHA9ODH4ZP5s7P3xvBVaY4OjZI8HBrm20mbT8Lb7HcFUMPTfFnjm3A0UU3QI3P
qv6JjoV4iHzQNGkQdbV6iuvzd6YDw01Q+QsLSxmW+kcQXv3BAjWy4LwyWiKSJ8KXH5kgeJbR/Inu
AghinP19cBW0DPIYCY41QCcg9uBJfw9FkUG2UBDZBcMZ58t5O/jskC4/KtMWp/43jUb2a6LpQ4eT
+ZOHmufx5lhAsT27tNf1G/iL0SpYS2Lzh4XCUJIu2sTnB7c4CTfgD4+1beweiQdWvXOm9N8mJxqx
Y0BeezROMgoID2ZkSsBswAKK7hy6EwsbYleoWMLDsgED34RtskPPC9HP9f4c9chQS0aOu/A6p6s2
34kd1tc5xWUk3hblvE6xcJfb+4uaMf6d+NHpOiA5GN7yMzGkTEQZqHZgI4BQ5+Ok32N5cN4PovrU
zPXlLUocYFh2IlcKyTfxeqKkmI2zfeLwev6ok8vYYdScCylsdXag/yEhfK/47x2dtAZdka+sQHKV
vTfDZf2pTa5ZwhbUMQlr7sXZwmaZFiRn6t3Piv1UJJHeP59jvEJP6qZ3L8rbS3asKoyIFr5FeurD
JweqTaWFtquRINEvt6/uBBKhzf0XvhQ8rqW9AH7zOOORoNhkqA+pKJFbvVviMgDTKtc3zvsvNhgF
l2iBOxl+gASYpxN3uuqSJbSKg1Z0FaEQvoOFoNEaPyhLpx9XP68LNgXZawEg2aRiCt17PvVol4RR
I4SDowmmGa922QoLjbVxvVG8zwDzfGNvkNfvK1O/+lRg1UMkA5Bv8RPYwru0PeiAqzHRwGIABfj4
De5asNQa0NAuIz135H8bEWbNBkiGfOfv8yNAnGNg7/RZ3+mQGORWG6JwQ6Xx0EnTH+Bj14kl+qBX
VEimWZjcGSPIQm4ioGCURz6IYutNwko+lH3To2jTsUYsCwr/sqXxAUKhdfeqscFKoWeWgTJI1pZe
FaYjNngjXHcnyDZIbdNIepUoa0MerxUUvDmOkw9nG+b0QD9hNefehn/nXSNEukioqXgFZ1hdkzmu
eSCS75gOVH4ii4dTf+JnFu5zug9SCVoCxYtdzmgDCtzaKMZjIVYbYYqr3FlxAYX0Sv7oXvF9Ze12
eMeeQ3GZpTiGN3x02GPtAAplIUvuSRZ0RomrELM+vKsVjlPM/WvsBxd2c1bQjt1+jxsnWbXeiTv1
cBUIyZa9ccZ6wQK665493lnsV8U9v7H9y1qPYuBhq9fKy/2TQffrzJkibWRVyFB2nx/BefsANN87
jmkqRgGiSKbtH/iMH6kGqkZ2DP96TdFJB93fAx7fjdCUCmzsMnmbeVE2XNaOIM0Xu0oGzwaUIPYt
lGWLrGYzChaMOc4AunTy9n6yjaa7yVoXpp5f3kNbrupmpBNDB+JqpGhubkwG13o7Z+x5bBkcZNQq
NkyAOpvN8Jkz/9JevRFEnQAyDOC5nGT4mBdXdmiDphOgXqk8sb3aFIF662yrDSgf3uE2eAKUwptU
sc0jSa4bErKtkn8j6MRUNMQ8sDH157jCSL5Mucu87SbG4fC0MCivh+BVP53UsDFcTjpmDiVd4H7J
w1qKq+xjfhu6fXKk4AoZdJodXAG1AJWXijLog+5DLnvn0hHx+zq6looT12OpGW/woNPNBrS76lCg
Ew7z/uyOOmUqhX8QpFJvHAZqx6RNMZVYHC9A4RdnR7EbURFhfPev98QeDz14Ms7xgNG7c4QUB30Z
jqjPtreccRWze+jULRTfxtzvEtrbieb22lspPl/7ukDcmves5wg8661INj/ljXyOkLTkTpQFwqAU
1Owinh1Mnflx7DF2MaVDpeszrqKNmB3j5KsYjMkDL0mRUJaC1GzrD/+3PdG49Hwxo9HxWjOrHfsJ
dNOohriphZGnkwNR2961pl8ju17CP27b4voplTuezv8qDDoHpM6WDlfZhJ8dg4w4RG2OOvot4fZ0
eYiEmi+ecwc38tbCiS4gJ6KKq/MeM/4yAAkpsd9Xvjf+G7Mu6DXfVAEj+7vmUT1vHyssXrBMJ+Wj
dbrUvKgClpabemU4QOkzwLssrqYkbMCqnLnfa6lVfKG3F9N1EoPzCHB0g0AgEmF9DNOinN1ViPjp
5Toej4gAcpTF84OqgEwh1ifNZtbFOm+CkZuB0gCQrZAPJLwQmHtpNv36mW0CZ6fbThaPcpgNUXeH
TfliThskasqjwnDV2UrcIDC5GNe0nI8yeROhPyxXt19AzW/nrCPEQEx2mFhZP6dOHbmkbEoMCt7A
6q3JMNqkWoWxwS0bYWE8T7R17VDC/tN0Kw1cSuVo502g4UDwuqph9eZ/JxeOh2oWB8dH8EDS4Z+E
+epLwFYiQJtyaQC2i7ITbjeUFXMhdw/wbtBJRV9eOpZT/6e59Cni6jS9r7n+b1r6ttIrHv9d948/
QDVTQM71RDvo+/jdRFRS2BRq7YJDZZBtqPeOJ1Wzp9aP7fO+NkxdBlixfLW8KIgpe/2lRSYAWbt5
3CYGkFdBHPUA/Byu/GJfGjtTe+6rpBFmntMwXHjAPEUzR8UZu+NJ8BWhEp4lWuuBKRw/3ADjWWgL
NVCxoaRHomeTe35wcR7QZGWSFdTnjo4Prq7e8yLXKgVnUqUNi+as53BDvfvhDiBbC51uxI8XKiRG
TT4BwOUnxCh3D2ZkD2jCxH0/HY662DKrSeiMBNAOnIXdqWoxxTC2+HC324gQqVVNHWMBIRQZy1u8
O0tGfaQQlm8zfqMbERVNRHryWCaAk438+4cWM6Pkf5ZZiFBQ7eO2XH+5IwXyOD/nM6EcCrnEGGTD
xwLoJaSDoQsFir9lMcZ5OorDh5QvUC2r5YAmAChPa8Rj6xkXbJAU9DPMC7C11c1OWJWQ0esVeps9
l7mh3fa3kIOGbgClMW+XcTzXeUuqODf4RbzPy8ps5yKVH3fSTXeHjG+fB84p7CZFjfrqdsa03NNx
koK8vj5Fd/L/wnQH4Jn9KSGm5sTvKD1zFQjko46Lfg+gHpnV5qDMxasL0g44Cvu2HszwqLDKuCfg
Kpri+jbNhjAEveyKV/pC7EacHFnoZXT6IYkoHZ6WLmwCeueC8WmjSyF05+muYhVFA8ehF6tj1bM0
mThz2Pc7N/NSZaUpONtRLEG7qYwvwEFp4jdOgz70wWehtu6lzHgWEdfCN3lGPffXoEvov+ufEM8j
EzzGWr762YAal/Zb9XXqL/9pwnAqCM/7Rmr/GJS+TDTlyD+WeDGGEdMTnmfrH1bPYdtebaRLYuQ7
O8BB1AXY0GMZDSHi2EAZICpBBdOQZQo3grIg81EL3KV8QWdWd/KDGzTvi9e5fjW4kF5z3wVxwJy2
a5IKmBJjOfVO6ctPCMLKoeCeVIW1FpqIKb7RAq/gANgEYX0wOwiFT/9KO9cNnMFVVWDjgdNFfJ9G
GfFDT1nH+lSI1Mcu9QLY5BMTmAi8Mxpum+pQCwLYlacDg+pdioK3jN8U6B3ELtGF4u63M59305Xx
vKYxkIxMdu4I5DBEgmDpA3Uv4dJULpSgiAuq12lyLoqnMidmRagN4IJhOlCj/5MCGj5AacmGllhz
XLvLBd4mJXNbkKeI5BHLccuk1a5AMrs3LkYNVUhNkKSpfWpgv1THo6n1OLv3oCGzspARYVuY3ZkL
F7zGlMI4kyK6JB/ALLri2Ufx6gdR+RU1emDV20uA8roZ1zHMM2tDHg38tJimsOZ/YH68n/FLdcgw
IWBh1Jryz+4DD7pCcquYzjtaCFWbNx7hPXU4TLpwAM2AeWXF901m6lImOOhBpQJrGCwpu6k1k2Cn
/pDuFqyhQfQPi97rK1iMnss+btCBnjEYb3y9wVj7coEdJa5CbkhPl7kRWjlmiKn/apRuESSf1u8/
kA3laR5GtkCSztA0qJjW8uzBZTinLKR5yNil1p2H7KkXTCcYOg8AhIaYGOZcuMKVB0ssMYteGuYW
ZwVc8IVNdNonSw/e7IUDX6EYJjyK9KkRfNMa8mTLTXl1q1cljOzK34XRpOk99ftWQBhkE1YAdLf7
1/rJECOfWrn8KJp+QuC+G71Mod/KxEwsVeqKNgp7olNcgiy5Dz7z6h96kOumb/o9LxMTbhlkem84
Hl6P5LDWbXuL/wr6jepMgsr7zfAz7rkEjJRWI2yt44/6OPO0OVrcDRCH9xrYuLvkd5a6qSWiHhYC
ajN6Yo5TibC1Z09afemeUd1Z7+GTgULQ69qSquik+4jNwNw/dLXXnkj185d2zoSZltBm/BbaYmxN
SxEiFuZqu+stM3m+pNHtF9w6cuKCkHLL6kXSNK3ubBggioqCFd/s3h4+W/1m5xpgE7Qv2GMdXZKa
jQm/GIbuWpzRNbfJf/+WkHkr2jq3VwT+Ohh8U+wac6waLbegzUK4ExFfXjHsPV0NN/dK1zPw1uRT
ykB1HFoh9arv+LuhUu2Jn3QrCzhJvSmVYd0E7IpSS4fubt0JONXiFTMJtex4+QCNhDX4zZUELOtq
xK8JgZdBeYrelJnxjLiRJd1auRoAbcUaMz+rQkcv/7R1l8+pWo7tniZLVLK+N6K7PfDS68dYPRZy
E+ElNZMTs0BAhlOyFvhTHuC4hOX/y0Rot2DEeyIavaBn3rw6ghfqZikjdBEI48opphtrmtlL7509
4kQb2t1s1jqGy2nN8DHwajEcxZoC/3ZLpqwm1zk6gOB12vyR9yIKm0q/pfd+uTdwaNMRpViaoxxu
7alSHQZOvkYv/wKMAdV3zfSA4BsZJEylVZjQtd9OMsqTZysES1XOw6DzgFWk0XNd045TrjSj4YL7
HAlvglT65BB4EOgMroLO8fUONG7TyV6eNsLnM9alyMCuooZM1EhNrAcf+UfrH8BGeKlrpi3zzAyh
E3pXkmJBNJoCBAD/kcZO9g/m+Yyz8MVuEEED/UFE3Qw0fQA8d256N0IhymK73o0mpN975mBUVHDZ
u3uUNPl0jrrD1hqAkBTwWgksP5gPXV6cKQdxkyoYs9QyjpxU+4HFK9AaSY1iNG/2RhlcvUH8wcNJ
FuVFeouLA/juwm3l2gQ8M0j2H921PaJA9VzRD9PHcZ5Xy1sz/IHmUkkbcR3W8wLRPP+8F/1HMpSr
KvgngGWLyw1ejL0x04/RQ2eQ6fQWKznEBax8gwz06xMyc0/+Hs+ipOOimEln1gwb9omnHRUDBjWl
TeEu2df3gAXffLOc+PV0Gr/cfsLpd74/eCRTVpDZNib19umhc6omEtPQHjGPvQN7m5wb0XbmHs0t
zM9ghstbE63StCCha6y8wWbFq4cxb03EL8XJsfEXG8P+zmNSxtmAH6Jlw/qfvhCgLwMcfzJYP9kX
IGtyp+wAVpyAFLtLiLvRAH+WYG3hC62Pt8kIk8LKjwPxtVempwM2tW4NH+c3LXjyC1b7+x4LowJK
SO69dRJOYsuFnGAPPepJ2UiAUUpaFdDukr7RvGQyub/1hG/1pGO1bWUlNuBCaPvQADd/Vy9nZGPh
+oYlraU3a41fXjLmzpyyhUCVbRcfXL52WiSukD6WViYsjqumVIWXfXxpniJf2Eh3h4AD2SKA9OR7
a/YJAAWoOmSULXgVYVUHWoF3uv+YSgOvL6w1KigZzqdVztQJuvXOV3xcjYcvtsMgBJWqVGWwodlI
6EEyzZqoRYYBZ0DTtW3SM+lA5+yW9U12t8qrclEyfkwOu+YZa4+65WISdLdgZ0mu84fieN8paMpY
aWeJPQAPVXIziuOuxNHATs7CyYI4Z+ifxg6OGW3RAGxRcJ0egYRuX6p15gP6ozrpzMK76QoSBK2F
XOjbzNKBYETnK1xwIczTAk39lyUfIJJsFfRFfAWhoEowcZWCmYRGSr5j/5Hx7XZFthYN4VOqvUDp
f/dvj529ctiSKbI6mqaYx86LVyje8c0K6cRdlKGDdSzLYzA8agX8FdVamImWZfrgSHhQZnPcvr5S
W4jKbrKzEW+vdkH4nLFxPSsN9oavcToR9SZdqhZaVxUlbskbhj4xE5DnJYbnZ1fXYb6wdPga9ZU7
Vzm7wTtBSSBdDjMI7fN32Jn6GfXJhRC6nuS5oEpEU1MIesyo7peJoT327nn6PBN20EA2uOWqQkZJ
/a2ugJO6hECcQ2cB55OQEClZj7O6Ue1jTA+qqK5sLP5QqSj42o0+YRa9qp0RC8ARv4ux2B8yJsvS
xk7d+/col9myaXFVErOBpYz60quIFjjL1CgRPUFjljX2L1n+nV4i4SudeK04FPBD3lUK3R0T8kPK
SUYyLJnNkG47uuA3WW5Keh3oZNVMVlXLas10g95Ze2iDHycMTQDtfwEUzRYAzmOcano/hCkKkvrX
mXHlXmG5GJPKQdE+NCVPFdnrqVOcUijGgw1LC9jol111Ennp1ztgw4a1Eq+nEMuIAcl3YTTYc5Ea
vKm0IR+uG9TaqsmEBpOsXkXefgUcrRo0p3Mh5bk9L3usGwAbMeFLbp0rHPM8RR5kqcLw1evU/rOn
q0MkL5SKgF8Cla1xtX+95DA9EUafWUUI2KBJE+b9Mqv+ijBEyfQ184M+z9M4tY7Zg2QqvFDptBQL
FLjdo7keMdYcPNVvgFKgFjyazsbq4Mzqzjdf0G2ux+5duEEjZLMjjdhsR1U9Pg51oXPexmBducOj
ph8P9Ive4kwsg8WXCYfRa5jmt9YDaq2pML/c9A8TxGkrUdu2rBV1TzIE2P7eO7AhAa9mJX8QWZGG
LDMFk6+gjHVe0M4teKRPOT9wKBQUc3JSmIoQRTAqvAAjmtx9FnE7VrNZuMZ/9v/FzjC1Jngv9Nn6
wvhAwu8j0XnROyCbaQYruXcRdlDono9AdpAwxKaecbAgppsiH9w3RpH0gD87rmGQsRQH7IzNSo0H
es2zYg3HrzeqctcbTblEFz83fKu3mr7iPJ/tQfmoztprCbnC1sxlqdFAxeiw5nQTaZ7p7dFyqJGG
HtxBQLgUMT6Avv34ldFvaDsOLWZb7lqFFznFmfpsw5CLZwmnYIx16MC4IWQRXXU6Mod5U95Xw2au
HdtrvqhuLYXvVk9cVhx/tCX4wnG4gZuB2oOS18aq9a4Cdn2g/4mWaxJVlYE7Ax6RK4NNzvwmX/Kz
a7AwwlGE4E1HtHHF9A5OURQUHbCmu4ROCtrpUHunPnuJn4M5yJXK+UmMZwfcat7bXKhcr6V6zIjm
JcKvu7O9o0PeN56x7xHH66TwVVIqSAbU4opmxTj8JY1ske1UldaZGbiS9CcVfw1dHeUBBrMqtAwW
lkPrFtt9f8ycKbc8NVke932X8Mp2ziKhnx9PtVV7ecw6AXO91DfUaH1BqKOABzRZt8/EXGjuegCD
qYqRwf5ebTgtpbJKn9Zg2+Ajo8No+WtX+7YRbAr4Jijih9my0OlRk1wPPujedXeMSLw4m8XUKPfK
qXCUvW9k579Q/EIrCR+RrpxlhNGpWhzO7a/hrbOfGz1oXXME3IQuHZX/u8p4NVFpwLaO7leznxVz
BygPNGnN1RlW91gKO/vN7flVO81Tt/66j9uLbnQ+No4qCQxtdFo9CpFiMGM7JpXipAudLGucFT/T
i2sHM2p2G2+Yn8+24gkjukghYouetAddfOCxcxoh9CbEhASqZDCyT/kGszczArG05C/g6AP68i3J
BLY9NP3cN2Pnt0MQyWIliVOTSKLInEVlc1G4S9+q/zdGOsWK6Hal2kAd083VTh8TBR1ipm7FZogL
S+uzXFKoESNMmpIUobTOHMhmVycroGMLwlZDzL5GsDg76wqN7Vdbp88VApe39sFUT7TH0BCoepla
mVinu1GSR26AvYAlnkyQ9RUay24TFXr/0IxN2PMbKpyiLYeQmiCKDnONMN/Epo1UglD6DNJeUFr2
HITKCAEdyJfyLdDo8hCcJn1Za3aGJhbJ9NofWWgOwNJ2InvjWCMBIluHZVY291YxJj7NBtf33WzH
B7ft9qnzkrpwoXlPSPgXh17we3ubICNgunpclwMQN2FlkRTLjTWOssPpNUbjEZGD/eNLSPGmzzZl
xQB48rGr8/h3HL5MZ8U11gdsPlW1Npfe9AAk/8fnK5rLnNqNDLGjcud37Losfq7SmiqKTeceeITc
fmRtn+BOHR6QacpFaEk4C4PYqfsQeL7m5MXoViWAfR69Wx0irJ6y2WuWu3Ymnc+v+vq5o1iKdgGk
Dwzyw77FvGi8i/rFR1baQAA2Eno1KlieEmTdB1U05oOvZ+Y+lsyHFxunU2XtpHqSbGdcGKSg8kQQ
KYWKqXJ2DgLiw7cOD90rUZYzB8HP9aLzZiazscAfsmWiwuJWJ+0kulVgeiwLMw2R+vGrbqIJBvfU
YzUqHuUWXRR0bwHK3LJgmOJWYTBx6FjDKiB0tKsI2fQLSphPNSwUzh3dNkzYrjqhWmFtHzPG8n5K
3HK5Gjs6jRTjy/cv5KTlnvW4X8AviDRCGb5d0QCmKtahS2G2ABt3iIbZLzib1s+0+ZBVfKzJ7BL6
rC2erpxs7tUYmtsBhw06HKzBMR8YmsT/gsdRhzvzx9Noq+eKr82OnYNLG1V01giv3Ov56eg+VBV9
N4hKH+xTMjUPuhk6szZYmjMlbQ+0weTOme9wTsBJTVyNz/1QfJSbHqkPadLCUvDga9ksf3VyjAUl
q1av/7tVngp96c6IiIoVyKr4B0DHRq98K1bhVPJI5FtP+FqjJEhD8LF0PryHozK+Ho0oiMe6vcgu
cnMKF9BPHZJW27czeRf+KsQoAiddSll+d3bmIN7upbJ5F3LIRm7DYkBrxletTzBqlh+TIFagEsqv
TFa/SaI081PxrE4dhSLsbAy8Wc0KDcPKdlh/RkrLsRd/KG43kOkql7ejU7XczgqrEJzbTZSzxw0w
F5lwH1+pBtS0VdJrZFaTCBGLMNYDCIuBeSk+wEDpeefl9EojVjQEyBHjmie1T6M7samDRYkN3LFZ
tnS7hZyhBTnYcQzelvdfOCfuS8tIUrDnYcDfIKEJ7IGQxSWA8j/PCv2U6rjtDpQ1VobAR6hMBM1f
lEyeAvtiziReoS/KtzuR9pydHZahUiFXi44rOW0FmDnjsE0aVE9WWeNp9ZJJ4BHy/tQMjxBTbxfJ
6/XN4BKb2dDgquIyBbH/eOkIMD/OROC2DZ2GMEvMFDHNZ3AgxWo7WG5XBfuIvvyTdJT4kwTl+GJr
ymX1FC6ZcmXVz4HRaNKQnWx9TsAytvzxt+Lt2HJNx2rjJeSclLdp99JdfHJYjR+5yFzpZcn+y70Z
BjuivL0z+bVkZXdHz2N7euPfrM2X9Qy71J0mZ25jGfegBkQ0oKKkYLP/MsoOvRR5kQz/iAqo0KYj
NxWsp2uTWgZfMFpwUtPFPh1NtWYR+QkzXBalaRzM/QhSPsTxbatySHf8MkWk6vKvAyiQwATpS/rv
w70Io+h7Zz6geCCBa6SwV1vVEHN7eiHhW4oqs2rmjvkatnkQNfk4rCqzG7hkGaSXQJAn2Qo41WTv
KYOTk4xHVhDAsEzZ3m4XH+8shft7PSNtu38fq5iwcv6cwkmPFRJpGTd1CX87blw0AVHddTj12YZZ
xBlCR4jKcW0Wh2cor+P2D3w7i5NOzNTwTVQrgkGrVYwPtyjUSCp1GkRumMDG4ZabCHTxn7iV3cMR
FOLVSlLrCpsFdyNuTlbg18/eE3H1Ev7Mf8XGyGcyLxEjI1fUrxJC8L8KBqiTExU/YVyS6wu9DyNH
Lx1V4S//syxg7HFDPDUskOe4/OBxhzIbCzBqBZ8BCXZVSci0i85c8FqZy+eNtVHI3hZ4nfEmkRmW
ND7GYmrzbwObXHOaLc+NhFZiYj7clqGBIXiw5wIiTQ0h/YSHiynEXc0sxl7NbCVMYgZO1i9ZwPxn
eUyZwbKCjq99bRl4mqXsP+Zt9JzCGObvT4Nzf/vaTsC3B7G4Tr3KiOlDDOH3ZaEhk/b4KyR50kJt
FmaNkaO+bvVzG6DkRhgHOIqhyNVwvA9vdpPKBym+LTJz56ARyB31NfDlRgWp6gq3GTN8YmdxX450
7xEcCkHCptuOJiCZ4iAy5yVPdMpFxMiBoSd0Aq/OG58jvdL08j1NT0GMaPQYGTD8mhvskikrz7Ma
LXgOZzvG3kE23RsAEEeLUQP9k/G5iVZOZ0KVMvvwtryQwE+GtORJTMyuNZ6eTK9nx0Bh6vEGg97y
me0GAsFTkxh4QUJ4d2TueXEOiX9yHx2ZAIrReAfex4/eoLWQRZwgVn8yA2WWnVWjpwRZSbz5GtMv
nQ7ZWcNzWstEja2SSkF7R5WP9Ge657B/OGBiI6OU85an9AbNV/1XvloTInkiIYY+3SQ5MZ1XCjRr
k22FmN+10cDOSRprMohZECVS6YFBLUwAMkYIg5D1TI/IOd17q0cfdhW8lD+cWj5jHE15E/zTayEn
fHtUZEv/e3v/yPEcYgLzIczHJcD/vUFElPHEwhvPLC9FzWpPfMDQEY2AGcWTaDblRI3momBjT6gO
xx9UYm+DrEKo4QvAmr4wC/aJhFRuPIoD7MT/XbsME+64TY4g5kyKA0p4m7cKp3x+ImmkRD252YPj
u7QKO4Btbgp1YCkBG4j/ImsC/Ak3PaoqhDCHXYYNecoQ/XGxaUORP+XVVjlU9NzDmh6FmgppS7nQ
44GxvgbylgObYz80yGPCWyg1BTrQhe++AsJZVY+k0TExpjeveSQC7swFXTm02+QcZdb4RJSBYOyI
HcQmr/7uHmbghchmmpq/evm/GEPYoXnsiA0ImJxGGNu6EsV6DWsFfpobL0U1bvtEof+jHxjyQPkJ
NVVDNU5m21LwIEY3Bf7YxYTENYs/2rzQqor7j+Wihyeilp9i6+9UMY1rPqgiq5xG/FIgXX3agitv
uRiyZabZWlG2knmPUV8MSAhJ2oYtOTHErPE/KHy7qATNvjQ7Qv3QtVC9im5bxhgyHG81V4JiYAQA
seCnSMQbKXVNa/4tkH1/LS3k56Pi/AMfW9Hjk9XkibV1WNFo4hpz6rIcpLapJaAHDWyt4bFaZRi/
USzOiknD0Nzo7DIW9hWrQ5q2gyjuyNaaFBCcJa06aQxAyLPWhCiRlS4aek54mOJtWDsIWnNdPYUv
iSfHm0RM6ZE26gp70nTkdCfHj+N7zrTm3YqRKsKX0mxYBYCr+E+ftedQb/dlSWZaQIxfuKNrTxRf
+vEK/1vAarfTA4RaBYvgNdciAk0GnBNUC1sn3SWN+TF+VDT4w3hR3JbQeEL1qYjp9nB0yULMWJaJ
vxuPa89M+yqCn+x65/qvH3beyBMtdOyXFT4K1cA36Osy8TYr6PwGgG2qXBidA3TS+jBsDJVqAzYB
QZq4JLMV0bx8NTCmlNky69dwYSNf0wWxjNzN+HbrRZqt2pa2WBr30ono/eTDVnPernl4B8AfS5h1
Uumy/3nX8h0TEw4vMp3NVXt/neQtn8BXhws7MFEPqzX1E1kBj+UmSG2e1AHC8o/LsYkToQ3HLJeG
m67GTCbDFkH5PkFFRVbn9FvwX2xaWAicQFgXVPDnEt+Amwwe6YlwXtRp9bow8bY+qSV83NPDA0AA
FAZvswGSB2ghV2KYMrs0QBZ24ZbKX4iaG6v3hkO2KgK0UuI4CyQene3XA7oQoZx8yRLno2ODtPSD
hZ9hNHDDlGV9/fe9mXe1FsouokODSjDCWJLNndTf3bT68wgj7s6NvlfciI/7pDC9+o4QbkaH67aK
W5OEr84v5mYf+Bp/PYNKiz64DJWOsgc3gAsjNb3DVedQ0+S0Nh1Yhy8L5zBqIuRRGhYx3hZmFl3g
/jn5V5WMWy22y+w++Y5wW85O8jJ2GJl6XOfmdrEU5I8bTI9nsKGM670V/jdnYOzQXGT2e2zuNROZ
hiKZdOqyRV+YcbcO63eblQnUQLs2nyFgm3C9Mo4ywHfK/REnETH8R9/2ZYSyRiFZyljw8F3dKf6V
fHledoji2OstTHIG2jRQdeMNU8oB6Do33g0hYWvoxztIiIQ+CwaFA7ZrayZOYHuZg4Ky0DufvInO
jJNK5AI7txJ2XbX5npzf+pOfX991QxrFqbJnyNLvvNb7sBJW09NNX0SwBatqwbpsPc0fTv9s6KZF
iHqVKDs8SXtGko8RwD+KpuwuxqTiGoiakgTAvIk877+qXIDmg9eyXS8xyMlvEL2LHEy0EQS/MsWy
z7/aLOHsgxbsWZhEIjk1FnMIOXIhlWQyN/YDZ/hLrO4sk5HC2p087oz+IQCCmh6bQUl7cfMTd+a7
O/TTkXzupwLt9y108qFNIMP6IoGiuo4R9t7E8xRF2/QZLEQBTdLxEne8wyj+G73kHpJ4nOptooty
SqwsRTRoQrrND+33gkf+ou6oyli89iTSwaHje80QHKzUE8RASkg62BCfdUzQQN7XCXRcej4gUGJ9
5fZe6vmEokcs7iEi8y/AHEO/41c2sj45mtlXKN0ogWLC+vPEIVyJv4cefG93MXAFZLZw1xGzztsV
dfadoAuD+CCUQHbWxuvEJ8pV4krYoeUPb3CGCdyQBDxcPKmymep4M+P6CmBRUUEc9nZNV2kN3MQf
nmF3s7Lqm0lNVR9AvpAZrW3RZheyx9Q417wQg6U/ItyPheGQvLuCgujipYbquBlOD1d9rFcvGW1S
cRRZS5r1S/LGHL1wAFnoMgJdCbAIDtRaWJF+3S5/c/KtndYo7yriaERHRiYmQe99RFfxRbvG+lhJ
n+pFhqRRkEVvtyRzl1MjJQ69O33VPw2NnFcK31EgZbYbJZJoiAjDPrUBD/2RSOFBhKDWnd0Dmkug
OR24nerIbUqB2pWwWNJDsdRk60JiK3GjF1Gijou5fb6qVuBkaV//ruWI2pu97LbItYXCfpeCnA2r
n4sgjqVkAXUn68R6x4RvHQ9Dy1uaqm+skQnSHMcMJN1DkFAyDKZrybXCvD92pKiGBkju/C/R+0gh
K7pTxfZxIP0K2OuI9YvrudH1OOG/bRF/uiZJjROjVJgY+0PtOD3itOJ1a84wzNJjlh4Vq2a54RTb
le930FLautXuI+lkkdRxo8Xy18ZZQbYoF6kvdH86hLsDQ+QVjBQ+RAXyXWvogpMfy1myBXYZW9Jn
fVx54viTb7ofJ0+lhOuqTyK66XuWvLxQlariCkECxb2dgZKG3EFWMp7+to14psmkPzfu2XB/15GO
BCamFO898+h1pAm3HEaeu/0O5DuFvson6HRgBj+WCNwS2PAIyUwdR3MjG0M4kPpaCGaYbBcf7spw
7D57tLCvsTT9sh9AnI95C1zL575jtig9JP/Tcy7YA+zMgII+y0JmXgkXg+tib1Wqr4sOk8q4Xa3y
EzBif0we4uT8ajUZ2Ok531RZpIwaPyjHm7pe7rD3MNexd35S5a0nPGZBxGu6aIxspum/wDfKLGBD
h/SbU71KrL28CP3rm3yW9Jq/+UbOmyOEZ21rLRhrUowOTkskiUQnIp+pUthr+FfcVOOziDQtQYuM
Bp6mkagGFjI6S5kaV9MlzlcIxZKwAJSIhRLBhDBPd1fUpUkW8K3NBrqhl45u75xch9hlknD/rwB7
ctOQjmg6QYTjwrZtfbk9rm5ZPu1bRPd1K+AAmxDzSC+/Hq3GIj40pYTeWWAS1quMb9Bpvs6n4tk+
C4sC6e170FQDfpmYmw/hIzCmRSCJ0+veNJW7OGdi9dBbQ9I/10Bo5GL6OHpxAtBgxmfbokV5KqFT
Rs7OjHH8asGOldyI3IkBQEXd1eqDy5GC4dkj75HgcLlSlLbHOtuiuF7kut2AvCg4G+rZ4BlLyywt
SYOZ+MDPMaKo1D7aSwUBlIJSj1GK654UW7jrc4lY/XsNAy8aeP/HDSHeC4LnbgsBxMCQ88j1ekRs
QTyYzzXVsbXUfoUOKXM0WORihbwqs0NripEbgzrKZDkIqvuSt+2AvJAPWyD2BCtoEQFNo+ngVNqZ
Q0j8RaDceL8kJufMQPK81Mqnp3tfgmt+X4Lb6eT8DsVQsMTDlT4VJooh4f9HDZCbYCnJ7+DerNab
BzJp2p2fA1cd9dZvd4xN6zvqkK9cAQcf12lWFoC6++iUpVWjYvNFBXf3Qi02pynga2qEciq9shQS
Ulf/dTxr3V9jeSY09YLGF51zP3x27d8e0qZKjDPz/LOP4vxrysoOQWYLOtQUi4N7u24YUPv41Cxs
DpgGwBiZzHWhAEC/4xV5kAh23corq+nkOt9zfgO7PKr/gFibL0GmT0i9q7lRwPtE1bz3C7lULO+b
Ie9jTXW+2hRhtPDl33bHQ9pZGR4/sKgXwI2PgW2HTppzgoA1qFORBHKoiN/lJLdTz4lnsBpeLaZD
3F4/X7Uonf4ifNKevoN1h/fwf6bf6yGqn7VuLEHVK2zuPMvPtSsC8j615TSrU12bg3O4i83y5Gwk
x6qvsqcbZ1k3d+ql0lP10SJlVr0/MIS4TxajstILoMX1HmMvURwDoiXz0Hfpq0YW6zeRDQoXPVQb
NP05zGujtmHMSr5hPFUb930szRAiCJC8kPNXeNpV1igqFfoIQQ4qivSvulD/1vf/T234MLGpfibD
sOFCFCms2aowr7LRhrtsgDnEbu8jh9CFLl63KpxjXQXX1UV8lbs7FZxfNTntuwG1lG6I2Hf0DQ0F
TPzfO4o5ROVuXthetqI7zEwF5sMNJDR7hAOtQEQFl9NJTBAxjMlppXTLHCgUIspord1khiHOKS3R
TmLxFZvKHJGmV6OBUsywR8tOXroDa7tNuiIJBuCpVyB3ralL2ih3KvO7W2KjR4KxiV7nhRY/kRfa
3YxXoHbJeL2EpF9tnUBxYlyzYBCIdtgV3EqzBrmg9RpNPmbmqljmlO0sAY69ZTj09x3r1qlt3rep
HeYKXrQHMucLXn4onRriYQYqVtw/9eGTCcXhI821K35CcMOXog99IY5v8bT9IuhJBYa9HjxnmqYf
GQDXubmckWZM0YqgTbm5cIeuGOLwUYqKhAKccaHo1iV3B14eUgWUlZba9g1Z7PCZCRjI5erL+a4E
G0f32PoFyj9fuTri7ewPuufPBkzvWwHjJV42gA/ADIOpRObwT6IJWyfNFtbRjLH0AaVuPrN6jfi6
z7CVV+gi/UppZ/XFNrqvGVC4pFhXvz9PkNkSAUkRj5qBN05I6ZIW12mX0J42BXeGi/5gdAyd2ZrQ
ZIVDKL++l00KnBIry3fRrBcUakQBPeTKse4R1/mXX0fy2W01IqmdS6UUcHzag389VJTztp3zsts+
Xi6NY29BsXxz18VDEVjTpJQIuQs9Xnk4aE/gfM+8sAmUHumIj078IA3l/1a7fBGHAZCI4uZEV677
X6zdBeGaO5kye2Nn/AsTzz086E+IbcTIYCOTvqGoP5H0FnQGDKSGItOZLCECxpEdMC6weaBe8Obc
E87ERE1HtpLBcylShAyuL8exAVu0/IRKz4mhAELouzr5hdgyNp++CcvDCFwZnJzLDCmxX9s8y6QL
x/3SdBn5cuKUj7f1f4j/kkB3SMbvhtJ6CMzcS1AE9FW07rtzQdO5oBPBspPiwgNL5/ZuAGAlFgNi
1CGYpEJSuYoounFdHfxlD6MP7VgMIMkiHqWNjQpPoBxQZyTtPWK5neclIIeRuM41rACOaPMdHJNG
JSCB9yigJA/zc3foctS2TJvdKUiX3S8G8PdLOjl6X3nDqz+mJPZ8tsbAlqYZa/hOoPwD+A9GHDE/
7QUcO07sOTt0scENLP7bT0dhI71HEujyXQ2H3ngkqBiHKiRuYdUBv2E0v0OjcidxwiePrWrDxFau
ScD3n2PTXOzO7q5dWWZx+RK2yGfdfJLrSC/2ko0URGBrFcXu+JD9Pgb7z/WCGgrhUl1OM2VLdKtY
aO/6Dk1rtrpiLlBR0dSI0MJmtVBISW6H89URKLF7BHJHXxtDa78nZPPzCJo1i4GLDWQe5YG8BHDL
zNFAwCDLxo8q2fklM9FO9d+mxnntsZy5k4Va7TFsKxE33DLPbRlArZVMZrwvyygzp0KQt2LCRYIa
vdFbzUw5MnwfI/I+GVJHBUSO2nUi7Po4GVtfUYdyNgZUoSRZzHBjUUXg9u7iSuT8sb341qeR4wAu
UXGIdD004e3I8Wa8Yg57ZpHnZBj/OdqmJuwqS6qgCeQLlptQkOYcEv/U2rpqus9xs7rqlBtiduGg
46gIPxjx8TAhwz0wZJOc3UVUApO0xJaj+v0ALVVlohlf69HJYJAE0UhjP7WdGGyCZ69TOVIE5UeE
o4+UEpUiRT6PqruiMVWxd4Me82V96fIYLIwuxyp0UUeQ+smVZLUR1Ah1djPRB1dWnK36DYnGUYcR
gNWi7x/CfZCF4muJyt+0sqv144GB1n00gyatXHOBObYQgo9l2uMqo3bVw64b2CyGOlGf0Y+Itxl3
jOn4K/6sbdVP0jME4BZNMHXXyA1Z2fWoSwbB4CHEAyjDQC21OCftfgny7KZCnQ9ZVimkXbPQE5y4
7lpgSuYKEVMPPlgdOcXrxIWKAoi/e3qjmeQreGbLMrSNje1m/eP93WuY1boP8HiNDp1FQKu7Wd1O
ZgKf280SrF+kdDZB8moCjmA9zPX93IiCTMJLoqxvMTWWoK7TWPNgFUVQcqwa8WXWaIFX5RGUK3b1
jHL3wOmu6OOhs9PJ/ez0G3EqNtJxKnilbdHVm4vs5NDjfRJEpnZkPAI25bvFwDe0gz2UbTMiSx41
uQ/Jo/DV7mX2a1JZdF28oFZZ7s5OH8u/jDu8MQflGOOVi00dsXa4AsmNdNdMbyRWdkUDizbBGeQj
3+lDfXagpkWo2iC6hFrBL2kmatqOt8sX2DAJtSugSsKgaL/TRzCnDxszsLnh0HoYNi/6Gm5/Td1b
pK+X36GMzZM49AJi99wR7Vwx5v9tu1jOD1xTvX34TlJIh9wZZgGqZa2IWxP8ypxH7pJRhFskEunb
Z+2TWABzX9OTovO2CkzQtqVN9fAK/EtQe/WRR886ORIEUOOmkI59+4xl6bPvDKBFyQ4ftWBmwDBy
AF/GkVc+HKcM3cRnC1TntO4Meb3lFaJrVO0DhHyxvdvsT9DgYEka4C+UqeqWWmsGjjMa4uhs73+l
s5I0NmrxtvUZ4D9fzJB7zg0FUSpKJfmag5ozTli4FpNi1eUv+UxVdYiFZjKcsAuVL2b5+yfUBOlD
1/fM/EwYzXn9P6fNBvqLnN+CZrah+57KhR4x9qWXm280O1nwSaojWK/JbcBJt6TUsknh8noQhNSh
3ts1r7uzxs1lEKZkTczWgwcnS7jdkII3cWh19vprDNh+8ZF2w31USCKxp7JbtnE1o0VFa40t+Lrx
5eY3VbgW/bvUoPMwXEZlanczXGWXNpHsBh+KqNx1YTK5YXNYr9u+rbKQJMgXEF5wrO6LPU0fdG0h
D9xMXvoqHzscpCbToXlLluLeoBByOKsBaENacqA4jGJLxTmAWbXNolqz23p4blpRU7uo2pQVmFO3
vklzh3booEEvYItGAXmlrdW9zUAk5Xt4flSvYZkUJSIRG2GiSAqwL5W2zQnIqeaUDEcEE/j3tNj8
j6/aaSiqtIECsmoKEutwpYn6ViAjuE7sZbpMjx42z8bnV95o7CcJMCFCpwxqdpt2/rxxqTpfnsti
pWZdwU4aDUMkdCja9ByK9HNh0omwkoJ9cvxRUDbSmGi1rnfOvgscCsDFH2xyyOe+lXYZlqSYAgLf
4/UtR1xY5wJfoaS2sqlrl4FFJ1jmRjHLuagvL1U3l2tllPKYDVbGc6DG1XPvelbt/2UPPj85KTkG
8sunNnRQ5kStJdT5zm46bEmPQXdZU9WB7Nmsy6XrjZqVHkzqd5sSoxzs9+reYlZoeXRYeIJ1aoAA
nU8JwHdd9Np3r9wKiy6tis1vsEgXllA5nOZ5UOR5GTqRiGp3aCjv66VBVnsOWXqJmfujYmWDsKOg
8ktjPCSAmiCpRvajL3T5Ay86WkeFysS5eMNl9OzwyhqIzGTdzJn8ud6rAxd/S6wlKeZgiP45ZvfE
DqTd9ITFDSM9d8MkRNzSIxO2Zy8prQN93F4KE3dW7oCeAQ4RNLWT97cDJVTXXfDsVrc5jV1BCGDI
EW4GZlIOYr5j2zfi4CRWMWSzmICiWwkOskpTJeB3rkHVhglRIk8nR4zBwzQOrKvLVJebc+o4SHNN
/aZEhalASVsJ0Tpa77z6tqcoU0lhC+f9ZFZe3Tjj0hAIm4imN5dNItjR5bHtAyZ0fxlFQq1fJlAO
MzFBRAbiTWy6M1z8MEN2I7rvC90fp3C6sMDEqIKwsLHpjRtpr1nfDScLJ64GGXkuFzEslgsRR2pW
+lvXwgEqBtlwfkn5z5EREieMRmrP8efB4KGbR6SrOAcH7TCTzuoQXVxUid1rjtWYs6ji7TmVHlzu
le3E3RQj0u/zjCvZxc871xmUNwo1DrijABhMhsXwnlX3+BDWDgNRC58BfFCakPQdmyRgazHNuVEU
vsI1Vxa0ETjnNYusqLK3rc2sXPVvia0Hm7weDjaGdjHC23Lii+eWx7bcFKs1A1DKY3ahUS63OF3I
kwfEbQFvpZGIqVJn175/nOpuvEgy0egmw+4FnB8j5M7SgsVR/2/pYU7pa18NgZDppIUR5jWdxW0O
s7zcqKb1HlBZ8aaaJilU9FRwpwBkkiVQKk/m+J57ekXGbLGr3K7N9gJgZ5eYXW5yYhv+oD4hHsWx
x/zwpKvjbu++uUv6FeaM3G87sjt5MR1ufJzbBOeKdhBCo8mAZPo66NkChSX/DJ8klc4zYKzoI/9M
b2dMz5wFAXc3GJfyaYHwDuxNAigwx97E0rrXo1TQk58y06Gge4u1MaQINBSqTTiKI0swspgdoc30
kCoHTvC3XCkewM0dt7YRHA7ocjOZJnIGcgy0TdxXzZ+xAzaI1RdCFnH5JINW5LVirr9ERqFhdAgQ
uXDEr/46zBptDY62k2NxBz3384oXPArEpFl5c0gFuYMo9xfvEjBEsjjRcUamXKmtjKoReKVT3oAR
fwilaK4C+ohuMBXXIgBt/XNwC0XXty+R7TBrGxe2E6lOtbKg18tpDLSGS3FqIWpeY34VRUdlb1VV
FRg01R/0rRX1mjfvWJEi0imM7hXCwLV8CvpQwXHgQX5s4s9t/HFNqoND7SDTSe3XQX7WHlvF2ev8
izsltNzuHMJu5zaXB4a7N/MC/BI09himVNjHI9BcqUZDyyZosSLR0iK37AuguVHOZDcoRqfWsRe3
6LFizj/xJzt5p1ofqM3OVzMF4S+zx8y2yqjX4Slg+kPx9E511+pURv/m37ywoRXFzBmocMfqsd9t
UCQirK1TbkuXROP/vAuSILocNKvmMUC0pX7SSzMPZhWipmq5pmmIX6XCNC41LOFk05uCqIl8tf19
v5Xzg1WuS/ezxUL1g/DGn1/hzJ2z0EGldRYqxgWyq65JAPzL9i2OI/fkXfHMDOcoNH4gKfh0B2Qu
DsITvuHyUtPVSaV3nmoD7NYO5b44m5xICHa2QX0KCmPfJgczM849gu4HfMBSZUZPzhDzi4pCheTx
G0glIkhDltRY8VQ9rVdUEZXOyG4nWIYNhXMLNmkw2CGAQAP84zOn+5lZU7rQhxJKS+QtjDm1bDDJ
2mUVorclrmukkfpGwitwq0bkO935A9rhmBWw55o5BUN2n8W2I4OMPfSht8+bTVKIbzpB9VO+j5lI
yf/GWFovhG/QwDhKSBE7n/ms7d5LgAObkKJaR8+x/lBNWe1ujZljxj4CFHd8T2TN34hV2wfRLnru
Q1VTmGTZByC06pFRXZC3KFn7Z1umkosYe/z7R/Y0SaSvefYNxcc4YyjQX8F7/Wm1yqxhYZJS67kw
2DcEwCTmkWu0WNq4IZDApQGYIHcPbbTy3mQUrzCd9F1BFa+V40PdMDM/i3a4/Cju/AVJJaiVm7op
QCZ61/s+IRwVbfrFBlb91S/WiDCkNXWwk+D/n27z42FyVeWD7rwLr3PU11Vt3vFlQZG7K4enQyGj
8dPn6/YfWdXUigi1oGT34KIP8jfuSG4WiqnEx741BaqesD80jmN5r4mP+/SBshdM6aX6HD4ZBToV
4iI+has8rkU/j2AgX4QFm0h/CTPMlgdNiq6JGkoprFXTjxxbThTUJDnWTB/E9Q6DBIH2XIp/p5AI
2lSwhvTz9N0yp+2HKhLjDvEwMym5gZmsZKIPTHZ3ztjlEcp7al2JaRD5lOR13BEMPjOmbU6Shppi
B8T4zVJCcmTnRN04zYzpTMntrmaGNV/JhPubjmV8EudA/dmM6YZIjp2ojLjmOhqb+LRX/nmEEFZq
/DXGLgIk27vjuW0haiD2c+UQzaR1rnRAQjiQeIB8zk3v4PWUMEzgqe+GThkDlGiOJw+d4oYxrBo4
rou/KbHAa4Sff1O87Vf74jyhsqcdcOPnfjTrREKhfX2EPOGvWbz3USR+Quv4ErZOmj6yXp9JAFD1
EUnoyVjPNUk75vDhLiyNA8BZHmSujR5lacgmdQ5Cb+keLKFuKdJSRyBsOh+GWZNr9jP5SBHuZcyM
eyukrdtHeL3GA47wRxhI8u7Zbl9a3LPlgnNbO4t1Qd2+N8x63so5N1QqGneo9lujkQY/hfqnFYQI
xq64AHg1GRVhpvGrI0U31fIkypt9OaxaW3Hn4oA+9QbnpBcxhI6SylyOtMvcZcSc6fYgYX7OuRgt
2rz8RISmu0Qb+dqnz6UIOsUyRkIB680b2yip1z/YAsfFPk2x2MPWzrGqXyHCE7ZyBwwGxSOiNm+R
dwfB++/WBJrsTfbxxnV01ZM/3apIPACXvY62m9AM6lKfxT2BJo4+cBE7/pviaWRXJwE1ZyOiYkWx
oBXB1S1CwmZUpUMIsIPjv/jEphVw7dMkq4kNoPJbPCW4+g+/WHNnj3AIvjDHH/bKGLxxWgh0OHzH
tmySAlzF0zymudkyoL575s6Vzsn4P0sNB1aPFuhJYjZVF63R0u8YcOvXo59gFAVFhcoeITdTJvOk
txOmrgpXF4XNCJgqigeleUVa1K4xiC/xqKRsVEdkt9XHtV6aj/u1V2GEn7n9gvsxGkn9nNj8xU2x
ln37hWWiHBFoLFJid+HXGQozUVRR+/K+5P9prAg9BhjRerccN5zwyA8HVUTQNTabzyMWiybhxYsq
JsuNhziR1/2JA4kMN2yMyhXjTEUyb7s3wplj5ghwcrBFwtqyBZ9cPfEOqbCvGp2UrrFViG+7HsCZ
ObtwNx10byYJMAkeqz7GPm+6pbc9DiiVz44bFR38kwh8RHMTCFJDXu4kPuwuPfG7mZV7B5Pqq/IL
gwdRmaqQ2nx2svf2EKikK0zpTY0TYdGT0r3oZtNeALTg8ecaZdd8hFzH1A2a/mDDsrOU8qHjE6dr
zMbHRE4kXEHb6otdLyVXdEkT9+3GMX3lX/5G9uVG8mVeEj2603vKTB+5ckIZtfNBcuxrAEd7fnB3
Qc/CzqdE1huxZPIPWP+wZZwTAVGurmoJ0BbiFnj7yEIqqykTQH9w59HENYCfJVh/q2mvqdXh/+vr
RVY7wKIEm2f+VeW68JpzKLfJHaEK4Lyr8rQ0uHChwftwk4uwNaLxW4kdppc6D7+ZxCsxSz+nD+rZ
DNOCMPv0xdDZAlxXPdUavg73xYJlkp4bbRIlTswgIOvesuIasB/RNAnsxNeKUzA2UNCu9xt7fJf/
m9t2eyo6KcGmO304rtOIub35jhiPqunZUPlDLI1txvFw/KmUqAClu9szE7CYTMFFJYbfPhJoYFll
7EjRIoeCYXV8xQ0A7xz4R34TPQAPdRbEY2ecUFdWXFbztlR17oIFWRAOLCvDDIcrukjnc5bE4NjH
Q4hqdwoyB5nC7xJNHY5EXZ/Y/nwG+OvBOoWA7zDz9DNlcd7jSnZyRRotDEEPqSKDxmyV3TOL3dHh
ZbjKTqTVKzSmuZ7yd7S6I0y5Hg6atm+nzYJXcp/fXLVZ1B769jcHKWo3pdmiFzTADb0T5ivJ4gZg
BYhFkSInkxAQig5opoHrfKRlk/lK/Il8vOXm0oh3deniRUHt7OIs1wJe3Y5KpKb3Ydfo4lvxcRA8
L9LBc2A4CTTOwsKEZCpy5skDv9LXYATS0QO+uVZmEYaWp6jWK2pP3hBXtggrWXL1UOUf8v1pLxSy
4DYHxBZ1RRXmKkoqWwn40eQGyoDza+ZNjgD4fonZ0PFqFaczXHEItvhRay62WaYr2Z0u6MVchqv2
LPkm8wL2V8elxcKDgUXs4VDD+9ARiJpdrQfAqWc6zU2w0LjsA+R8ZyT9H/HfUbJu0ZWryJeqwaYP
P+s5/JSMxgrQn3J1ByQdl715Jpl1L6AZ3dQDTvLEWXlgOJx8StNEHHn+bUlj+MkjZjZXOgxQ9iqP
/9IIeeU2MXU0KzcqJlCMOu+I63DC90HDJgobKRlMgwHGGM+MQFG81jimXIn7rqFXIhM4DoZriMKF
vLbR+vA26YgMQ2ug4rFqmUIHe7UwzgXLDstsLTB51aMGL9lejxdPxtW7zU+7w9HxqmJn+kKeCxEF
uEuQ/g2XXnvkf/MX1bVHQ6hG1zaE2ahgCpBUvMk6vdpgtx+EeZmbwkBwWrXDY2j2VGmGLyeFABzL
2MsIlE7coW/cPCX7v3WtTNaGpLViqEN70jkLURXckHNmgK3gt7twQ0keYkfY0uUmDzMkGH3iiKI+
rnX5FEvSH5Q6H2uQkA9uOpo6mtVf5UP1M3sID00g6bRfrcVoHeU83bdrsHgDQo+KUsWRveVQE0tg
UHcOpha0KIiR0r8x24kIgdOK8sD7Z7tKXum5gTuWoVjcAhu3mxEi4zHyFB8ADCWCN4n/OmWOzayA
CkT+HIsvMYF7UTmG6PZXOgHJ+OT5Tiit7fAM0ir4+5SvahFFZUmiYy4L6B75bfg0wLAwAUpRaOsd
jo2MsYVDl4af6pO9ahnTb8WAkSz1MUwWGRq9uKP8OcNXbaLraJ7JKbbAY0HtZND1NKUQK7R7dW2c
dOA/Ce5yh/okJhgdO7eWU0gQwnBgDIBX5pp6HhFA3/Lz7+0NXUG6tqUiZndxHKSPYkOnzs3TtGbz
BcPEmfJq7FJoTkQvOtJRSAxhTi+NECerjamtBUNG/idLGGOQx5OjHPrmFArY4SelQfYVkkrYiSRk
8xI6CCMqgKXgRtcvga3x9/AIFisVDWNTNm4oLcI/RZPlmO3YDzXzO2c9f5mVDO2K/2Zgzpe6twd5
/uHjHpaUccJIqd3sr6oaFUYRVykkQbLyj4csxMQCfTb5XNrNuRbsHsla3tTZ6m3ahY61q7JG66jz
jFCcnmG1cdU8vHh3MfVMshN/R+/Y77csvTPnRedu2BF2EtEpfB4Zq2TOV5yJkzE3nlWZqYc4iuQ9
zLY7YuLaD7Poxh2eOlv2axsPD/CsnJ1j1YdHyUwUhss9wdsHq78M+gaenT7045H4gqtFiEy8zBJX
rEJQOVppvpNczVAXxXTcgOvfCCYRvkouTkjFb/jI3i5uR2PSKiwf+6f4KtFsYm61yGJ8a3Kz5bX2
B9MNNzlWCF3jAuqGD3ZvLFZJDI6Jw2XVYjzt2ejynFDPMjunbwKlB/vu27KoTeVE7/DmqAcGMI4S
flX0q+nOqLeTT0JRO6oc7WmqF+zUHuSdWjaA4Bivt9uaPNzedv8U8gfwjpHILW0u81hgqy7I+5hb
wtt8Kz7U6NVqPXMaQrKyu1zJbOyKN38ef7eGIxfPERPN73q/IAxpAb1JJ3R+RuyXXCs3TDeIiyqZ
aJeVv382JhbgtQuQSBV2JtnQzyVsddVpxJO5m8RjR2PPRc1UcVLsOGDeuy51lWZ8oBtKAE3icR8u
bflQl5HLuLXnYYOP5ki/7QMhrGVswTZMJsif8JoZD60nUoRsWm4bo4xv1XZCWQkWuLQkc5Ix6Knd
RLw4LpvUTObgKjqLKv9dZ732joxL3fMBdwIEN5i7dJ/Tetz7t8uWStQZW5W6v62MWmFYgfE7+UNf
vK8y7a/ifQBusLnu6tr5lxxzQ23MLFhgqdJBX67+XMK6KVEr5osfJp61wY/vJFmarAaxEsYnnO5c
Yje0kQPAcV1CmfZ7125uaDIO9NuWMMwaNnU/TnFeuiZ+G6+DD2ApKs/h+XwqP7ieIA2EYg0LN2xO
JTSjifFOr7dRE/+SYFPopPye6+fBPGgtBwEro2z0zu4OJbQ5CQJKq0U8CvScqAL/AVOuPSsKVVYk
79oZtDZgPVLlu2d3En9D9Vv1RFw3HtX9+F5blpsTCLZkzjHPKLw+l8sr51WGn7hfrWcLv8td6QGK
Uu62BnDxrQw5BLGwpZ/uX/xKaM+3z8Ft2180zIkBk/62PToSeR9jNr8S6GJdorZllXAWHunGE6CX
qM6xGiE8kWoh0gOOBFe1eh1o+Y6daoEIWbhnH2ckXe1eGBwvw7mWLx0GKZ13ILC5VyHnkK/+rWSF
19rOuDowi1eTO7/2dKi9tIMZ+ZEXrFX1I3B50zTjrHHXq8WKB50SJHf71OHwDbN4iwe5nGDEa8KU
rflSFcmjSzotKhXXXkgz+lLpZfxHN8rjSqfP0nmhtt8BqozUIVtwEScyQc5hEP4VUL0wWDvtD3AP
sBiQ8gRKZ1fe3aKlh6jGo6rX8pOeKeNUxhjDFLr97w+qb5Rhfnsag40tK4Mgk5PFiA3IJEtccwVf
hLEwa+Ua81jVSbP0eMDN5JEDuCedUr0Xu7L1/r2Jfr0N8CrGz8t5Kfaxf2z4D/uCZbv78Jsr0kG3
la8DzJMMMaz898FJsv7/Wwato3NKitiDyFh2226ImQtA2F7GFFp6FbtBgo+15Q13N2l8LW7Koofz
qAIz3M7bFFVc+cQDnWJE5ZDHIEhgA5F7EFNkvDupJv/V9PFy8denVDG2BXOnHMATBaYTBd0neve1
h8KmV7WqAo2lc0gg++8u+7x/OkrK/ocoo1C8CvBT1l8DSXlgrqfE4RiYGDHKENaUfKXYxMl74+WN
x+aEQL62EBl9Q0BTg2m0xM0uYCWfuL+rUh9AQHKV2XxZ2aPY/tAkeOVTE9E4BPl95BnhwOrFEtFz
sw8neH9msvpJr9JBAr1kndwGhbo5GOTYSw69u69HjaXOHhrAbd56g7pOaegVD2crr6gfTMsX6NKL
ro40iO0gf8j06YXNE5C7XUXtAFOpVnl0tQkOuZvXcNyzWWyXoFrhpdu5xhJWjsq9LACZgSd2TVGl
XDmvItf1wkQPTdAFlKVhKUxv0RKGUHWE5NlUAGfu1EJOpxUcVkdSntanoBwhkNhrJDDGxIOVNUQd
SiWbd7fZmHbzPDkU23TpxA4HCyA8i1ZKo8KnKlWtUq2Mr3LvefLv6sBHFftPGnBwGLBxcwOR8PjR
FF2m+iwnqDurnt8XxUa+N7sDWn9MhCMV1cWfbbh5Rcz6bc6NmzI69JpYq+Q7L+p33qbvaQS0U/ZI
3aKmzW8FnklsXeMm125skGBCa5qE2aHhvDbObIKqNIuwSnsswfXkXHNmseSM572imQdS1HaspKCd
S3umO2KANPuRrF+Xun99UkfebSaHF6Rh3A1nIF7IkVXq9to7MflJo2bmXlHce8VvA13H6E6Ab1QX
6MFFLqJAS8/AB6n0OJ24eOWNjQIGpz12uLxNJQOLTiIHTLaDSlkXoF16w88wtZP+1F6ebyIKUyoZ
1m+5iedjYcjj4foVyDjU6ZcTnRcy05XM7c5mn3oykkeNmZhn6Y+pTKveV8YFuqhu7u7x01fE0r1U
y6y1fKAE4UUjMknV1KcaU9JaDSyzdKZISlIOITjlqxZDVZvmewdu3C4KxB1+FMaUVlqQdxHZ43cK
gCIXP1+Zrwghi5NQX4qfnxXe/2+TKVpFVK6tpvBuSxFVDt6mjF6m3Jg/Jcs/ynGks/OML53wkJyK
m2MCN5K15NZKNymJueNBTs0ZMIt7RzSEwY6+3JmlwUv5c7rlBccX3msYUQDNvZNvkX/t4Lh4ouB4
jn1RMBP2t7UGVnGbQ/oBCNctdGpzxxEqD3Bc6hzDWixttZts6fWUNTZ1j85zY3M3UyWbq2Gi22sa
ziN1HfpBPvqB2/YCZs5ReX0ri6upMVo37agaJdtJiq1Y7mubb0R/ImegmpZVrrKyKYanMqrRumJ0
9te+zJaBIl2Wu607+iv6IlpVspZtNqyFu8BaRBfmoLPjMcuAHDT3surTvOHudpylku1wu4lXPNoE
7kykc7xTudyoK0QQmF3RS2iTn7So2MOSCK+/I+dNQLydAIx8TFRPhqnpVvtnZJ4afzQ8SA2ECKGx
ZniYuFe3s3FZCEuXwMB1EhqOhP4vyVrw9dHXeoezBHX+hwCnRSrrBZZZiTn6u8qXb6lmncUpAgWj
kgF+/RWnlI353HZhmJAcLPcWO1FzSf1Pfp6JrSfquzIaJzma9wLff4L8u83ElJ5DICvXMpDoUxXB
UJj6TmMU8ThaL+mcUiusjpJ4osgnZuhopYyHXvhr0m+JJq2MD3AzueJe3U9kdB8zTKfPlS6zm06I
ubabyoCJLET2K8fqShRwafZ+5BpXnIpfKR7eQDyWAEFzMibAvmpllciSeJxnMlMBcghr322Ayt2j
qJzdvoIPAmr/H0vZ5tjCm7FkisZaY9vDzQsUj99bUGp2/L5PsSqBOFEChWSN4OiIvqQiOLRUuX2X
px2bXS1Aw6d8qhAk1CpUufQmp8/6wm75oK44PyGK9QYnUg31z8t2onedgkYW3PRO15SXVabInS3n
Z/JDQ6ZDDHMC51wpwK75aaJuJjbAMS/RQy0+4aVJn1OLh+hPQffmE2CDDCWowtv5JxRq86PRDxVa
5HNALPYO/cTvqwQOGBQTStvfw5V6nEcij37sbSIM2sRUc89Hs9OKw1mu4uatb+6Ou5Ru+8fN5edJ
WnaYkeFUjnevTThGbr++AuPKq+CWQZdict8biGckZAr7C9qfdaS/Av0ya76a6dQDhcNUJcGkGepk
+qGMu1oelhRZmlGrcap8dYCAwyIUgT0M0tSpX9t1ORD+vBkknFApg9tQyodRdNC0vfqCl2PMDqP5
dVVevDPD0Yn2KjO8KAAwyGMLbr5F8kMPMMOtt7ksTBysyluLhPzHOKlLHWA1JpMq/3qU42RsbZu9
8Qn5ZygjHc6y6PddgkOomwO0UrpeeBaai1QS80ivBjye1o5FxnxTwcubc2MxGKk2nFr6y5BGAyV4
bhSiho1aARnKYAedtlFFGJm0tRO+iV8lfzirT4ZD5/PFcVAiP/qiACofNE4hxvUKXkEvediHvb5N
ruyQ8za+oRddBZETL8nOm0lOIZ1NmNBKRDtEe5xzwa9ZJWNV8viQ8BVjuEVXqeW86TAhO/KHbFgP
s6AySWrflUvFHYR9SGx6V+OUlFX+jg8cSWaUsyg8fIEzBuERHg026wKSSwHgX1dQ7y/RLAz78ZWa
49g9149MGjsoTbsi8KpR7GVtFVVb44PNjxKvT1wPmIdJ1c02jDZOIQjO4LI4HJflirJ9tCQHfNuM
m7euRRQ+SuKcNeW6nf6esK02KQr/hKRcnYU51znR8M0IwkJ6Mr718D7t+iLjWvsKi35RMJHTAH/e
1bAtg0xMZOSn1W3gfFUyN61zCIVfbwpghvZwBOYI2yhBUb1G+lTCFxciPZEFqf8YQxX9A2IZXqb3
Vu7LbnqBdX3Yg9vnrZZ0OUlEJ1G6DcP/PNIF3dAzSAly8j27yOGo8N6DnMzC65DrhCcoUqe3YxJB
HcceXFvrAbb1ZICbEX1iHak95pIWqA7e2kBwm9B963fz2kx1yl2DkbkYA4xRxagaA5lcTwoFX33A
mCAv2C1kQNKBij5+gjQx2ZQLAZPbDmMSyY2lX4ND3epr/LLYspilhqIz8o/cRBqHFR9B0ApX1KYu
EvhcV2pNKtCY5AZUukIyvv3/Dd5IoHnSnz9j/F6kWRGqzKMzeMhK9FrZN6gLtEOGoXB484MrKVK4
VnU2ihB+ZBjIt+TimA2phKYYHUxpFuC8UPN4A/PnrzbsiRxRUWz+yuEVwXzzxYwelLccSw5WAfOS
e4VC/wuX4yGlXqVsuihGZj2nudgmcyC+ja93J4FSa5HCvwns55LJIc/vcrjvN2q2Y16+bioUU2eV
i4BqTnTpfh4bXrQa/pm/ne4B30KKUBpB41U2LyBnRRd1ObWKShaA6d9NfpuuJjHX5xqrmhx5uQIc
NBHMgUwS9IkxtfWkoP/A5mapGu5hZKl9X6SRBgBiYC2MzrCi07sDQIW2aHFYMGxC1thGvYrtMXON
lsnCtFB/LNSGysnzySeocbcFL2Qwcgekm4ZAxQnZRFe8JzeVlZk2CuNisknLkX1cTAQJGy95+1Y3
AbmIrXUEz8vqywUcPn8OsBSOOgRfLXbrOqJ0tu5pq3mBpPMtj0/NrULwOERIPQ8relFBopR2yiJ1
AeTgPXnuhercOZJVG9KIJ1sfXTr1URE+KxOAky470YKsU456xGSeF1vNeIfHaTOrHDYiYQbO/mdg
1u+CkQ9qnCJYFKUGZiVJLtBG8CzGQqL+bUf///ay3HE1kbiT8u9Fu7WFUqyFwCt5JF9Tbjz4OFwL
eLydvB2l0J2ft8Vh0cje07JyLMLyKnp4iTrgdBNIh3L7iJAj2zNnL2A/q+jO3ymijJov3K4S9Hkh
4Tpsvd0TJvW8AjTN9NkoYFOFBckwVfyp0hUKrhRfJhgpwyYHPMVhSLxUaLSP0ezw9tfAc8JIyIp8
rUYeV3UGHuV2l+77h1j+/mTvOEiy64N788r43FXxpmiUlx5PYivjeHDGcTkI5/vOr1l90OcWsiZd
9cG7y7WySmLzqE08rpUXOGMDtezyjyJQMG4A+nJx2YGdfgHcFflHBJuRwJP9JDk9t9jkUFGKdneg
2rrtBq0/FKk8o5Km99p0mIlq5RcF09d2lXzB8tvnKpbSFBVv3xauBHrMbs7touAIaT6kVzmpT9CX
guHtnNiNwqkWm23edZjUSb4wq26wVxjIr4NQfB/rk3N360O95W0mwzqQ+KT/Jq7cg5N2wESX0z8D
M/EoISR2LqZxieYx36PB7p1wP2t724qswE77VvVDn27E55EH/tOSm48cG0YBk6suYr0nVw94pEk7
LR0BY07tNR2bxaKvwPzcJh3xx/0rjO/kkZz1IyY9uYMgkTctf2Uo5vRnEZrWEBh1zG0KTXOlYnVs
Zb/ih3HtDL50mz2EVcKgRwI/rNH6dmtb81Z6Mii20votESYw3Z+nMJimW/+ztG5FFHOK7wQ8OV9N
2zA8jGM2ZHtH0Gyoh1bbRj+g9V7/D3qEr1Ksq1ogIQbdzBOAZWM3z8p3v+LCsh11yKaKRAQNmfvR
02jhpnw6B6P4GS5kpD7wOGReqXmanZYHvng57j+Mj0zAtRqXn3nzzraJhARvFv5nbMAux3jfT4Ew
bcCxAwhMr9UoPwLgeyAE3+LgGcgHg6b+xQVglZmgQ53wIEpXc1V5dHjAoHqb3VWMSedHzvzzRiev
EXH4SlhRggDEVti5v64SG2TAZBvo5OJoYQJ2xH7IqSdoEx5B8Yn6+dnbwhj8IdeH3hr5qja2w+u1
w/lmV/AHqbb8oO2v1Lov1TVbxrEld9z/9WXc3EdybfP8MJ26JHtoT+E3iB0CMtWuF8HBN5P9N2sE
JyrhWowrlH53V7IGgnLgcnxNrfUKF31tRHzC7Fy2ZBWhGlhyd5PK58Q6V751sYprX1r0/MS5WgMf
J9SCe/TiAoEjgcpUhvehNDFJGh8fzOJkh03xM8++NsUCKP94JRKvLymSbzU6hGscQS4IQMsWS+pA
hFCt7tXe6SFnJsO4Ce4fZF6adlJz+T53SmMOLjCtJFfyybEmFtOGWUDwVaG+wESWz/DaHFFooT5t
P7dU8D5pNNGwgETxPTK5Rg/S7F4gffTxR5DIWcfK3B04FYeKpViVr7cGoT+OCsjNUT4TuCEPZWYo
85G0+yqsKYilFpM/2HCuPtyeiTQnps8UHcvepe+iqmactLeBZ39xePT0FP/rz1YWdDNxIGNZnWBf
DMT2Nr9RVVAJYegy29FPUW9sUvnpaZNBenNcy9Iio5H94ChjDe9C6ktv3b9JWjZ5BcGnnnt8RsXt
YObAS9qrHBBRqc+j6SBYNH7bUdK+bDJaH4m3xIMALzS7Y83tXOAZeVzyskdu5bO8vJcLqquEMZvb
csmVdC0kmIrrzPLkOekLU8o7Mk7EA3fXpiyAozMCqDsB6vACNzlYVM+i6jTgEUdTnr6dQfJZFrWL
xNcB94fIoYVKhL3rXMc1tnRsX8IpT/oISQaHIKAJKeYUTA9TLj0GOnXf5Qp5nDGOQheNEs2VW3kX
gPJKwOyMEgEAyw54jRhpGJByld8WqrKlkb/60QtIupSqbv3T0bmPLl2OzcnZAMYCmAhhKb+AkXhZ
pIlpUHPSv5dCwH96r61OdFrL/KZIfiGFORBnOCl4qZyOgj1wqjBf9Hn91hnyKRWWLZ2pMTv7d+qR
6E5VIiY18uM/Az+bsKYhhyvsPFnykHnBhX+oTkXK8JQPe5L6BDa2BisaehfU9wC5eyzg9PgPfp8m
j+H8IlZJHGE9nyWnu7uQB2um2vz6nRLJ9OWUjWv3diWwII3g4UJp8z556hlnisIWlXcx2BWeNN5s
SIEilkYA23jThM9OGxi8koTaQPBBVzaYq17NdC0LTWZFJ6E2CnSUCUSOlzG3QR7MTjsAku5SoWJ1
ftiRlxl/PfxdmU/saDFagJRfcLRNyl6pXE1uXJXCAFuZTlF0wOMQAS/hWfa0WlmUAiR23TPKy4m7
+61PMxh8+IzKqkwBrar97fRJGW8p+6vsEGxMQ/yduybmt6I2/2+Z5qVHaLMw1SgEGo6lq26sDiEj
KX4MngmDzkMZcY05LolF267rTI+cs9SqBiCpw4TXPNcWlAgOdroNsiKV9AtB9U9kqIF1Lob1+v8P
C8recxOsBNIJsMR/ctf10nsW4ZZhxufrzF5AF7Y/lXB4RU/5H8FTI6XHIAltR/8JkEDJepYYpmEQ
L2QNV+mC2GUtOLAywgWBFyKu+oAnq6NAPlsn/egF1tts1BygjBObyJcbDAdVq8MBfED+n82/XmRW
75oA60vUGxiYEzrs8QPIZXvf9av4w6JrO6t2+HIf0ULP27chUZhMhknCFxAB9zwJUzYrK0Lzesgv
8QbyFVEuRsyG27MyymLnj+yUpBkAez96DXUgqxrh0VuH4GaF+OoZXr0P+CVoDhTQwQOcA2L+AU64
NZEbVlRN7nvGc4CDoK1tvIJcth1XIeSpg4CSkIo2iYvWpsfYXUerYwOkqW2RFKtZHgPs7E9Y+/uM
s55TFYAPK8WSvpMJRai3mBwAqXoMlYUWplKPXXNIYaThLANZqey3nNZANGQcEAFWGjk0I9RAPmSO
r8KXwmIryEgoFA88d+9+XPOzCPqaTr22gfMAFVW9o2HZFQiQ3K0jwskuYMNUBfj39dAYFSlV4ngd
ERKKcbzWd3hTh4VBS/i3okFKj1eckgdlrBgIWXnS4BL6NOLUx6XNhqBoHys/LMHjdusCDXvjiYi3
A0bog0C1svHbBlno3J/xZr0vkqGvjbTuA9wsZZWPPAmDEbkThjGlWmN8yQRMU3/2dfozL0KASCXI
kmDUu00Lb1+nOusKbFuUVy7dR0a250gZvXN85Dm4SwOsuHIFaZBD79nY6ok9JfIAxG7HkI6UqqrX
CnWvK1mmHIYnmmSwMOA5RI0hC3aUC7nvG+ra9DYhrmmbAxodMcJLKXf98y3Sa0bXeEeVFUNm9PSd
ggpIVzsmBoWmrUqf+FQyx5ClfPqeD4wHlbtVLigk3K9IhD5J/YxvU+fRaExxVTf20xnxv/KxOZ3y
H7ceqKfnbhaOa8tceNCdsyKqXpLCKSHaeStRFcRvgxz4+LXI1IUJ42MZDVxQZar9jiLve/DSVh2J
D6xLCJXlye+CNsmjHTAUgWfpwshMlECB+7axWtU3kQsH5/c3eS0FI+QPHKJBpis8zq7zoWFzD5p5
s7tl+k9p50SyACMorqJ1ywh4sRz52lvc8fvts6Fdq5D27zbVQiKs88PndOQNaXAENOaDYiy5TJc+
zrcYkY+peWLvGF3oXlZ+8PpyL3rRfmHvjeTH9yryfeziTkaSWqJXTl3Mkm2/UWypoIYIwMHOmKVJ
pLRc8suM/2UZGjnpp0Kg2qD6jqe8I4I1aXA6tuDCENF3HQcfu4P197rb4JTjLrevEd7CW0YI909n
R8pmTbiLyu0KhkkAGnzW6WqaOVBy1KSjnS/Dy1gGBlOmipfiyoWL5HS1vZDJXuBLKvp4js3k9fOb
uJoJF9Sgdd0qrObDGymyDUr4p3R6ongWZV5J39OuCdpp227ipGrTXJinASvyvrTxKQ8ckaM5MgSD
qRJzDhYXAbQXNZzB8INLAc3alvxRsbsPPKgDl2OrY9l/84b8kZkjyeeuk6DCNDD000mtMQXzm7sc
AR4fG9C5RUeoQAQInVkBlSXF6h9hToGaR3O+VavIWYQ9mgefawmcT32twCfbAL4n8X+fInGkeW+U
jS0D90dOWgIBmByCsQczlgVY/N0VyVGPVlkG8+zXwCso+vmTo+DWcHj3C50/hSqg4eFP1JpAyY9m
0zVU68SHlkzsFgrUgqQdu0B7X5y4mWGUVbGlYOYtc0RObrDbuXiS7ZF2+oalsvpPatY1h7FIvHL/
WkHmC61nbejgsZTkARnlYw+tJLH4GYStZEMXdebNhsJqyPFbo4ODO6lrdc/9SPc9qsKMqT0AszKu
ALieVq1KpnocbgWKjLL4RFv0CntY4v7aBWDma5pXDgDhJgDbMmn3pdDg3+PY5FYVh+AjgA2Mb2Ae
9A+VRE8GxWhl6F2cETJOA2jhaKXfr45R8kaMY1Sv69x0qfqY2SVJlB2P+VrRf4puSljbgnzVWmzG
qcdkR7Y5hQpbmgcbkBrXql3piN82TLzQqy4Swf2vtSsagCbXwpC+W74D50XdTI5HaeCmOZ5Fb6gG
O/G9bIzcQI0FQGBp3aJatiVUzpRyb52rBrUc3muERcjaAtx3wtLPAjkWRLY+WWNa5GClcskWgEuF
GROKNGRI50rc8Z5Aqz2+kY/e9+6x4oDqE7ySqwoZDgRFLUP1O9s/a+1UtXpMBcAxXq6EBITHMLXO
8ssBeXQhNajYgIJsRfZvVSBkzGZfkG6Fo5tMQgXUJCDGJ2FzCN7Neib+Mv8+ywc6o2cyz4xkXkvg
dqkxvm88MDzS3iDPU8WCLsUWardQ5jRqpuxexllO1SwAQme6N5esTpS+69ZZnLJmFAATT6kfTPpy
KTgGDthIamsU7XtnFZ3w3G8rIZL98gsJ6yOqXm04BcSJcaTgexgD+/sFlogbEFZqfIGW6JcZALqk
1dTVP15U9vitGCNwF4axfI+FNxH9Fen41OleJAaNzoulNDQtNmhZBHuCIkyJ0fZ4WzHFrSHifgt7
+7gVc4lFdmo4D+WgLVFSDGY01rpF2wMA46OtA8rhnAb9KwWyG7KLMa7ffOOq6v8CJDK3ow3FF0Yu
x8nQOwsiYLH5DkwxepaXkiV2YzJ805ENV1zmHZPIZEPT2Ar9tdVRVji8Hym32EgDxv4hlihLjgyH
b+pTzFyzJRihlnjseOWee0emnSg64WVtWUhVGOVuYszmuV3aEHbXGuROwzDTdtmzHV2m+YXQM6MV
biE/GxpOA0rJDdi1ezMoxJVRgVECUGWsAS/N87KRZGd8VHafQA+13/Rl03Vwn7eP0Iqb7q9TwHOl
DD3Mlm23dIn4+mykUbWcli9QKImHB4Ttd4oZSoAZ6vmdnfwusi6g6bT9awWvf10NHlZolMkDIS+J
VPUqP6DWtunpIndsWIqHJFfRtMmJ5VIU3oMOlWe6UN5Ms4baBCHQintX/OacRGjgpGOV9RB8zaWF
sKbK/sUhGrV6dfNt9WNvh56WkGSNBBnevGW8JDSQhy0Lm2TzYrnOSkXBQw19ukXIsh9aq1iFPZFQ
xuZaqXtnERlFaRj1a/5lxYAf4ellOPi7cS2JFVvvbfH0F40UyL+Go1bzw795okrtRSsrBnf9BbYd
mUWj4DL4kRPG6LjWDtKnaiQ7WhxvzYF0WQVryz0Nvggip5agHVOU2/DVc7rcXyvpMrZX2zQEtPLI
rd1zuJLpAdENJGl/N6nNMCQwIspbLcgTH0Ahg1S9/Oxyq6Xs+GjVQDhRLGqWraUTwuOsaRg4Z/ve
M/7l8cAT0vNZewWePkcHvB9WTjU9AshnypQM93ptkHkgRDNVQPKN4RpAEOt+R7C67XeD2t1dy8Oj
apP/w6gIWsFDXaf6c6Bh1HrZiaaIpudHiaWLVK7el6mHiTtkHn/hAb9N5Fu1L4stNLTBvxZztTxX
9CR74g0Vje9BWxpME/TCaxOBFa1Hh5WhQ7K2vIApcBvoMWDheYsFprRmvmz5/b3kRqEvFcAmBBIt
elTF8xDP/D1knpSw3g3b4p3EML6ovVCO12r0VxOD2l4YHeIcFcVRRPSPg8hP5QH+R5wlpCuRXERw
j9s9UXJmfQCGVqV5jES8Q6eklM+FTlUKZDzQitnnjetrw/8GTIw+bl0lj8S0lv797Liy49fMzOTj
kSrpm0lmINF2mbWPQ9vALK4Ke8e5jwOfBBSOoSQa89QbawxBKjVugy31wAapcaQwaBpuDDr2YsW2
LTgxEReITQQ3daGRrS150hAW290Ob6fV1sJvYIZjk6W1xDSnPkGkMZ91hB3y5nLozVFLHqRkmlu0
xhGRHggyYWXk/vjR0zjY0BvPPleSYRVXEb6gSXs4/qV0dzPCyvMKQVti3hsTfwciMUoR/k+UxlFe
7j/SbWNNan6SGokfJanRLpeMDGGJWHjsjSZQTViuMGC0vLZGezGNNWLosienWgLHb+0BdhPSUgwY
AL3RrmNkHbwJQxt9zM6Cz6X50a/OPeMBrb2eD10xiX5PaWBAz87tkzgiE8IF5F/BRg7+OmOtRWd6
wz1eY4oRZnKMar6W/J5Sg9pWCr2f689AaZAlmuDWlvzbDkwqnSOJnDEStsxpUTvmy7xJJccSCIzu
icjZmKX09QLTJkIzs8tOi/0b7CDXfMeqO/4SLBs3Teh8YSCFw+NVvaQ+NJ4bzCdGrIBHwNmzKZ8r
2j8PRg7PBJchKQKNBCpCJo07uYNSzb9YqVAp9CXOYnEQ7eIsDYt2TYWv3Wgf0gyniDpIquPthq4R
PyzuZQMJE0VnKoAsU/6PhaH0vIMu8kO6KMdDeThM9VTBuq9cmZpx/NCfxx0OQFdJy6NumambbDxY
DKxdq+j24t3Fi+gPICyAk897VJ6lapz2lfmuzG1etzsaRT6JPoRqgCFMBZxTx7tO1fE0FFyQGyRD
7vqlZZrM/4SQdKra/LrDoWNnhi5zpl4FZs86KlcEXe5V5HXkX1FTaWtskWq2DmFj4GPYMan/UxzI
0nj0ID0LJJD6GYZJxY/nFCsdyzfWeZDQLh8J7ginFVrwl4uOedF7po11H3ESDBZPiWc2iq5XNsp0
GvSASyi33PVB0Hk0t6aUTWhGzOxVCHjOGfXr8/t3zKJrrZ39lpPXYnbSiCNAfaMlGgkHUI8ZYccF
qschpGIQms84phEsPHwhyUYdWQ2IrO9jW5NWS1ZyICZQzIdAbSqLEFqUL5AOx4hnnRyi0DNXMfdv
vUGyBsv/xAyeyKgiEXsFfN35Eni0OKbcBiGnZtVVBj/YkA1XovCykaAr/YVQbiSbtkCQnQi5twq5
MG/rsxRBYv87Tq1HdOW658r+Q42TDgmFQee/4o2nTxU2hfzJcOczk7rQLAHprWoiK6tYm3+eALOe
khYyPxghnBvNllTGPwNTqMX1keudCIp4i3zCpV6qVyo/m3eVbRakGn6vLQKKLxZlGkF66PgzpLwJ
VkdhMMlmt7LYK2suZ5c+zFDyixtnvtPdc0+lcvpj+YLvTh7ZQDUSAC6KeJOS8Z0X4Og8LFuVvajS
g1gSYEMnQBVQUAMAtBp5mqWpIVdL/au5eygCiXKFOI/s2mVzEW/OVqyQa1qPjiK0JZEaV7zfFZtb
gzthKXYGTQurnAWYl4cP6XhwqjM+CT0/UxAWPO68EtySFevnGiGHQbY5rnek/MyRI725x3v6o5/7
R1OOuKJ6c2xarVoAOEJngvYUi1h0f291LMe+10uJkHpYi9z9TUhmHk6ooR+WFyTKruuhNx1JTua1
Luruj4OZLXw3ouYCwFqVsD9knexgTBXH7vQYjCEICFU7UEz2NERUTR275v5Yfgy+Xc4mlMOLqm8X
X145FMLZRRdL2QhNFBpXDQ+m1iM3BahYtb7mm6LPS8igLRuBiPxkWt+8n7BdlvqRDXtUwDVs4L98
ML5C6fZjApSaMMUvIucePLnqSsa31++oKrRbuObF0yFH+6VFP4zRxDpBF2U1N8DB1Xa88LvhMd+G
VTaIbVA0xxurR44UjEHxluA0HBblHKb3YuulbhbL89AhCUwoPywNoDyJIcYCoozuCxz/HwbC16Lt
UlD9ye/5r8or1TISge12eWafqwImH5DVtbuM0NWzseeL3aqdZmfjvnc/M2PQismJYmJkD5COMwCr
W1RyW5iksxR/tZec9ZnZBSKrtvCiWzfucmkji/7g2kT8lZR3a6S6BJ1holTGlQ1sHrNqFLPdE2UK
GnMOdA4SNhQcTdpvo1PstqzSVm21dQ7FbsSRiYN7YDeB6XQ9mCiUdKIL5GNck67lkyuLOTlFpHPx
VwxwAi6OHXDLAGWxKg18JPrL1eCXzKyFiDdXZipZWlYoaft520rTL3PNwE71iM8mBLUvl/wcPmtF
DnMhEfwyhe2z1I7hDk53hE4u76qr4NDdFTRClpybyWMh82a6BkOtX0DrD2ZYLxbWka/7LkCXqVR8
Fb8FgCmzukw3jPfnL5CGn3rhXfBGUaXN6IyxVSJabxo/cbyeulq1NGaD6Wi7N6W4a6pSrJbrxODt
ypn6hvhUGmdZp7YG3GSaRoBHHIj4n1sMf2lM/c4g2+yFcs9th56wOPBmxH/hqbQ27zTe5DqLlRGN
3H25D629aDXEDvODrTlcwhiLbq26N1btG9GPCpVGYIW5tJdOFRJyHZsBeoXmMnmWEBqjCSOlVNrs
0xwQyH/YJBPUoYv/ZyDpO2vNC1ulsvKYGkyqqpOBmJAznzehZePfk279RhpuxvxK/CGFD2ftv+GA
I4OJ0MjLCA+qdt1mxuzTGhxPGLjZ0SP85ct/m4IJym/cXXy3mrPRZtyAumjU1+EZ90iA5IzIY1CI
B1p0xkBwlPSzdsvBF9pcnknmC2s6+B55r5UQYHpQb/7a7X4q5ZrZ05Cn/dJBLchh3yDu8+eX7Tmk
yU/WDJ4YeVWufAY33xv6CzoremTWpKZiAFG0ismldEZkXVVPc3R6qW8eV3c5JRsQ+odTnfYl6SpK
IyvZ0FTcG0Uym/HXMgyI2zVkFmv9MW6bFEvltMa9wUeQCeLw92LgFQcIzncZ2rfajRP+8IchPIQQ
quVbVTHnjTzUB4XSeG8292IZR625jIeHSJzIaolNdJmerbC6o58JsxOmglqUy4o/CP8hzPOSPAvA
JTh961e48i7RZ4P3wZ23+o7Ek0YKEqSOvq+Ia5Z7DjfECnz0hWxJ74HJUmyJNCSoUGQeHAlAhMjW
q4c08jxuYMT+p45BKLPxAKXYpP95EEn4nLJyWyEwhKIDGifFkF7AJNNZ5yeSeUdhki5kYtW5p6bT
LjfKMbtmaV21Sk7EX75Fa1b+7JZ+HJtn4BSHq0lj8nrlzstEHyfEp6DzpNxtVu6knTMzjxO8aypu
5D4zwxh69Kgjdhu2AmAAOQbOQHe39D6/ZdMp90fKQUeFl8rKXZUKqRkOctfiLZ/duTZRCUHsVCg6
rhGmxEIEvNlawEurhlCRb3+HtfakhFfHRLmF/FYGPxssYqM9kPIw2bxWBsBcr9AzCgytPEYK0Djb
F4GvL40bVR/FmvdVzKrbc6f4a8pNBsbPC8wele0PwNn7FCXqgkvCUgERJRDeZ9OOTX44e/S64/hD
qdUdIQyZmSVMzwUC+OrSiLsRHW0EXoXLi3EX5Ge2mh1ymaU23dRw1iJAMHw3rW8cZed8jREf0KYD
VGWRZHj9FauXbRUENr9rz2HTaI6eeoP34zzT/TwN3iEnj9XRtAwEjFtYiNDx4etaaEj/3FwJ79H5
cJruL81nQLm/w2yiRbOn0L4Q6NwAmxcTaSFJzm/FLfJYSTTkbSQ0JxQv/2c8GQz0WtS9WZlrN733
PPHNIhrojrvxXzHbLKtlaT1xf7M+GzfOpYOyFER5GfZcaP3KvYXncAYfyYuPmBpZBZNF9CXoZ7GY
5xrvoGFvLTIoRN3R9wjazQmPIQ0qjZ89RBHc9CvGWyLADmJoa8PAvSQV04UV/+HQdIWrBaBwtU+m
qGVMVXQKIledxA1Ycgl3aWc3Ec2b2pB2cdD8dYyXmzD0JI1d6St1/octn0ZHujswUXPN8lkxal8H
1IsTSKRKUBqai5MmoSjFP/dGhy+0HzWPTRaNNBZR4o/fZ+TBZrz+d2mE1QqH5KE7RwZC0Sdua7s7
gW1Qy9t29iY34TUFwRK8bKE1GGJii7vG9cYr7IGaXRPgCdWPAcTWgPcYoS3Loe6+U/x745HyaQUs
iRKkyY+zHoGA6t55PXiGesxnn0zhILXAwyc5VAyMr1wY3gbCBDUNKmg6i/cFsnBOYKqncYnogfLf
x13Gh3Tavto2/pORkB8qQpwMiy6raTMPQjdT4xooS0dUCFfRGEboaic9SqjpHGAoCO68xfjVLWFo
aUoP1s5cx17EOcwwWuuSSq199p4MszWpHQmAAqxY+YrG8ueJ27RpVMnw8ZDLPAju/6eU0OZ6+q0t
eewQhzf/ZTudMPHk5x2YobBmP7L5Qxt4QTTKYKaG9iWHB91y5/zxjmEdHDT3J8OO2xSQah8YfIAG
Tb0gNy0sIrkUM5bVO0MZ2iLe2ROdCG1CmKR4qUP2sGBoPeW+hO4VaE5KxsBQCo5nt8d/R+a1a7sp
ogAWZ50lEgzOfcXCaxv9whWsSkGR5zdEKYNtbM/YUjK46lzSmLukDb1ZAYCAiPOjg6OYTvUc2+2d
1P1HihZNUGlj/kM6dp3Y2vsGCTb6yfg85ZEeJ/bZDox/DqfdUP1ZJqtRzZUcjsMhf3/E6v02InMy
uXA/ZBibgvpoG52MyK9nXojf2rRK07zwiZCVHtpHw8gNtdwS3Sv96BzTWzzcFT0S4Q1xGk9/wVNX
8VVPR8HwSK0DQAM4PbrL63vUBf4eSmwlG0Nupmd4RfLbFHzPogPUiwSDOIKH8gtu53VItwikGkId
b8X3Hz9cR/x1opGf0kk+rFzCYUtYgq6+/JuXQNAbAvXv0h6AomeEC+6TIb+cKtZvjJlD6Xhk2F4y
YovqotKVrYeF4ccmjY4szp0AjXsdCzxZN0usgru/fQQ6SZ0ExAMX9kNKCpTl9HJYmFmxxBSsxF8T
YL6NkOQ8HusC4SXCPpH9KQ2i88HmjTPBQWuyivitD75q5rT88S3503JwjLm853gAYIH+A7C7Rc3f
aR6LbQm0mGzw5igAaeNEpOzHIhdDrFXFmrHuBh/EUFzjimXzVvj7EZOXJfPgjVENn5CiEtmgeriA
br+9np2Nj7pxjAwM84YVYJBdxpgsOj0zyvI3I7oQBkLCz+j2I4vM9ps26rWVnR/m6fQwMQ2MCoeu
ikwUCxHB5KCtROU/F2Lh0wjA2ouOMltRK82yKAG81umeuRNyFsP76A0l7CuO1Mn5CmYcpOSdhH19
U7DFJMfT5hi39HpYTKWC1I6N0S3uAZY4jERfI/DTpO/x8CdtmgxJ4LP2Q2313hOvdXrFrtnFL9Ot
vub8s4xiMsSU1pv5/Zhg1XkjE9hmZ8kRa0CH606CY/i/9WZa5f2Gy64aOQrmEUd8nC4GWf/hooLz
kUVBfP4CdgtxwS17uYQo57lbZisrvD9jEhEMpPCBH+6jMid17eDMRb6GCRUb610MshtsvSifsVsH
TG28nou71RBLRFFHtv8ro7pQ4cCiijRn8LWnRVIi3FEdksCQrvLfgCMWInqI8r/a6XJI5SFwlhJH
uBt+pyek1kmA2y31OB3lKYTqpl94zBdm0owQwN5CJp79Qv1mXBmrKJqgGxyMorLLYtrwTIm3oT/a
2b+h5q2NjfkkDVE4dvViW4KpODyhLAMsnjUIl65QA5MbKvXC9hKPzYxPruKVv6zjn1pkCSFJYO+D
Fh2m2l/1HVmEJjWlL09S5QLGHEhR9OjL57CW05DhHbQLvXjQky7k9atm0dbYvgY94wmOtTFFaUH+
onkIbpIBGsvfrujLHODfBFIGAli6tdI3ULc5/7vK7mFbyK93Kb5+LQxcTXKqs5CnLi8BPfVuBhVk
o/nXwTJy3Ci4LPP54tP563r43rpLr3Q2NbtH5W+5TSF8FCGF2dTElEqaE/ViepNpjNSh8cqsTJla
khEOExls2q6t5b/2/aFirGjYJ5Mu9cwp/XX+HD/RouzS3l0S+CXp4nl63oL5mZtdav726QpTnUwG
zXgnAYCEpWoJHAkB2ZokU+DPZHYY1iJuzPml25x7SougEDs+DF9rXy3J1RfZ7Lq23JzXnyl41oK/
+0U7n9eYb4kc/JIp/hV7n2QxE7zjc2hTKsqcS5E8LBK3yRXKoFqe+uyNZhyCAMvnDjOSHHHtvHPj
5s2TAFBdnOcR7GrSaii5e2NEoZvV5AO3sR6ZabieK2ZuYszPv5NEd0Sumy0Bqel4Qi8YeKYsW8Kl
SGkQ/uM+auUZwAmHfnUcSkDJLM24P/ZwfhwO/OEPFjkWX8O5ZUx8lFJ0iQu+Qm2J/2bjsdwGoVhq
rRc8S3D3tXvKF8qxI8z32OhbK+JSpJsIxGLfcBDzPzQgmelZF1nuvXWhniEthZYaLo8zfZAyVata
5MtlxRKbwZXRhqFF059AyxByTFatXroQsjvtfHZdXgPSplZ+fLaMrIJlpBhiy/gX7IprMGF2ipuX
pzREppv2VNsP7IcvHEwB9wIAbIKqOR528U6+qLLqIXDKlsn0GbN4THZSMm59iiCUC7KqfWEA+Djr
QQYh4sCKOuQugHS0Aq815FotgLoqlrOD+grVUCDPvkafHebo/X1m94oxPKLh3lhaR+bwNgJsDbUI
heVcdf9xgjzBXU1J8NII/1kV7jQ+zXPD7cUcqh0N01Ks53kXLhPgcmbnLu6itfywEHDufzQ+5yln
W4l6H0C2WpeChoAfI8SXqEggUCIRXZE+Add2uhHRsx7Dq4LqLSK1Og1SzNnuDBH+A+tba7XjBxtw
eZ2es8Yl9tWSYGYDvSYw7H47IGLxqbJ7JNntPfRH2JBtscB5oPtyGv4hr4pWrQf00wxE51bP17Zn
4HylnCPoeZEUf5kx5Q2vcR+wkYmYGKsxUZn9+ZwiT/OGdqObuq2hqtAq10a4eGPCR+j0GnHB4eRX
wItM0DFsUAs+bBGLvf5ITAkwXsExRMAgpQuzc58Z8q0lfaSW8kKsu7ZGwcwUWDeYJLkLT5uKfmOY
pCpFRlBVurwdYV7510cwGW8GohibgVxG6tLsri9GyPkI3QokM/hAymgigEF6tlTn9uaK0JHMNlsW
5CZlwLIXm4qblB29Qh/2dMpCyU06mdaXGx119hRZhNz334MPBJMo//rHflUWDRqGKgLZUCBpFBVj
qZGHM6ktJb2QWg8F4HyYQ2i6hauLoZKUIXL9lMBMQAi6Mo+Vc3CptJyRx1K5XWVW1IRFf8nqGOs8
w96tfORVjDQ5cgSP+aW4+tHSPc3j8rpM87GdLIQ6N9YFZWNmuBlgof97tuAIcHuQiPVMGNfu6Clg
yf2bq6NBjDzdYu4ppOkP3HfGejrp/ztnraf6FB36kvT/Uz2Xf1K9jhdFa/iQ4Pgn4zCq0lTUS8yC
3XzFvuQILYnhx+jCzYjsoCZLfzMOyi9rvD9m3dY+MebkvNdbWwYv+o0yssSUOWqqE89sezBOKpWE
Om3abfwbfkAW8iXC8q6oZMUYwk1M4SC12yqI57yJIRBI34Z29UzTZdAC1ygYFK0dxEzi+taox9wp
53gC5Ew/YR1yoTDOd3gUYA8/4LKyQ1/DcZb+GGD1lcySjLtkpFpLgh9R9jin/ZdDJleD6V7ZmLBq
lQO/fAuVdSkKt+z4TD3h6nCtD+W/B5ihQbHtSQnLkxLaOBrrjcFO0cuQCRUFKLg/3oussihRefQf
DBB4pgTCBBSp4nF7+J2fJ9d4SoqPcQuyWuts8uIZgLIl0d3KCqsoHvJHVRCSJHV4jl/w/tbKKINq
H759AiQfsWvWCbWEjvgJJpvoMSwSu9owa29A8BPjnINznlqlAOdnxgbFbf/Gh/B0AmRKtRgT+pPw
ApkusaZgJP9sBcDhsXiN8rmh+XMn2C+PoC2TA3qMX0wzvzDG0iT+hJ5O0ku66qSioMmtWag/yPIh
rcnUMfjN8Sx6SVlya9iS//TmCdrrDGwvjIOAFovuxhZRaHmAAID7Jfy7gQc+AVWgSogLmPjbYq+8
u8VZZivKkg3Kf3B5Qef3mOs2v58Et1JscB2oaD/o3mBlCz5FUPgkEYKmytZsd3TXW89roYd5zFto
ZAspqzrnsYMzvc225NjkWTRYDfKgayGPu46lkceRgSQ0xEtLLFSS4mCUzqLLLqtuz1jhwDEuC8Qo
FNiNSGNX/5O4JEuLlfij0jlrSsLF5dHadWvhKtzIQ3mRMh9V/PX+rNr0ATAgyc9jZuZJdZjbCFtb
B8RxaLI+YCAfKrf7Br+hfVhzAPzniMzHQRRTulScaLFvPB7hELyIG56oYZYXLSGZnVydgEQSmOoj
TKEHwskL4kQzGwnnDYAig/zzDALp97V9YQwHCm4G2rW1jvquQYQCSAkgYmohHo6kwKrjEi4/Xoch
dRcS9nKZIdtzCYzAFlIH+4TyFcZBv8MHOSMKzMdmA2f0gPqICNs3PVpfzaUikYuhQ36YJHoKpBj8
g53XljyTjHjANn9de5VfDg3XGLfTf/vQlqsXsgfCu1eIjxxjeu4aXAGHx2xyX5AeJUg382AJuYQ1
1ZMyURjtuuGjIXFixFZ8Y3vQMRavf41ZDN/LOSSunIjLHRyK2brlEqQnBTRPLTzvsEfLttcbxvHz
D3P5uQmxwg1B6dBwtZy3n6quML/VVkQmrnLRe7+/p4zR8+dnHLxr8gTLzdOAkjojxlsVfYc8QyiF
gk4/B5S3gTdQqeND8KWvH8eInPVmOoSnmqyUqooqSlASskLU3kG1MOHr2VLohUAG9QohVwdVSgI8
OkK8pxUeKsBYsAzEp4gc643tP/A+72ptUtfoc+cx/+np8xdrfIErzVey5cJHNvJTHzm9c1fjFDWx
NhONT9OAAmJAGaJJwoANYusFl57E6ncVvAP1koVCg9/TwtkXCHFlMyEonY8YPdhZp4TR3UdsmiT7
6r26e3KCp2MKs3cSkGfBc08w1JIjt6rl9X7v4c/JQj6SB2sw2Y74Jo2IGfxPvWX4rav8eg+/GR8i
qFURvEtmfJjSK/oXVKlrw5dLsBAXMheAzksWmgkfTP89fJ8PzJQsiorOIh+Tsl4qLLRUOqzKevhE
0+oRZOqqVzx5fap8LcYsVfqGCijiv6gDBt1+KGWOESQNa5nbaYHGioJNgqHNLtVGWMup0xLOODu2
VW4ilFaRAlon/E006h9VqY+7mo0jH75Up2g9Jw43Zq+Q79205OVHgVqBlvPdRDTjlPDrmKYSd7xe
gc+2WCQIGeamy553MWtSkcesjXg29nxGjFfGHqvUIA5s5OJmSuwaaX2c778Y/VsX2bB6hdZPRmBO
78M0k/eXDupUYZiLA6OvUUjhlsbMjVUohtpZfjgY1mNywi8z1ozNnmrkFKs+Ny1mp4OmiINxK7zi
/N52qMFxjyblubrrlvOxxdj0W5I83yPzXwQvcGM/bzyUzY0tBzP/l4PNWGynvOadPwNMuNN0chjQ
WaUY40kmyub9HbfzpcRsf0dFY7gq2mP4wFi2l87XWefuR9uPqKUqG6BN/dTvURaFaliYB8jjbXO7
rfeZ+WcVRdSaB2NBjm/PYeMt+mxR/Hs00eWzJQ2k/j/YyotcVgqKrCFM3KCMbL6GN1ssDqk5ZCBu
XQj/ArT4ARAhhlWlAhLkPrTt6FYUMZyvZN1J6J/44/m966S8xclPC5UlwVdOFxWO/ISHcnfaSacr
WgK0sRgQWKo1A/JA4TGP135Xfyty3njTKcHodOu5qBfYXWu6fTl+C0gwtbVS0p1PqsCVBONJp8Fw
QL/gtk7bbjIy42VS36KQBQsJt+Ozvy/TuMIk2OAzbeJR5KcSbhQyN6Z3xmTVKZr89S8z+BtrlL3Y
RWp9IRYN3R/u1JQkLhaFKojWwKBNMvnPX4YNwjxaD6F2uLAUQ13gT86q6v0NfS5IdPD+tVT9CSyL
ZFzdY7EHsl5a2XALFu6YaXZsFde2lFoXc5ZhSOXol14ENtbeJarJ6mnzS+EIa1drQVYWyqeSOBzF
iy7+SVIoI4F/tVNrnWEwv87RZxNl/FHEvmaPRiqIzwzoJZ3HEYo6ASFf2C2E/pnejpJ9lVhRUHhQ
4M5g9E8IkgwPLJiZVShbP6OquYDZdBr8JORTKlNMbH8LVkhkAT3T9tEn9umSbMTP2V93QRz4316Z
x9lNi6uKsogBi+/tAFeKbYkxJerpBRNkZcrzKVAm4bGwGIK7OP014kLygl1SwzVSqpNurJapv+fO
qQssLvTuF+DeU2FTLOqPM6v/E8218cmIIQ/sPa44WK3sIjxGvahBAj1ztTWi+QzlAvND9+DNja2X
gCmCt0cM9uVq9N2U7VnTQA61DOqUnqTiT0YKqqvcdyGvKLEPVLaRidw7BACBYUv6TOyYtTeRJb2z
OML1oCNiTwOslWs24QozHSdeOS+zljlloxJvxISXg4J4xUkQ4C5RlFgA1Or40O5FUxfz8jxiFw1E
TP0RVXJw5x4mABVZg5soq8CvI5jv6O/9d/JCyPm7prqmI4euYj0TLaygIwV7AsRK17DP0VVVTjaI
Q8DtKWTLnmNl9vFrrebm2yvVtFhMZ7mdB7pwBAVLvxtGWacRHGnmF7W+0wDf2dviLLNEB78SwbQ8
KVHpFo7BqS9Y9GEjxRLwcGw2NyjqCK7UEGJ6NeIJS830PD8raWlk61eDEyS2HxaV8fZuvQf5bvpO
bpzzvmlxEGxlXjbXr8Rz4sGODYAQ9+5q7RqKSr0tXiHRBSFwNSnzIQJHBhvfED+5yeKvNEzZPhjh
GEWvkPmQLz6qDhCFM1HVGWBp2xbATbIXT07pNXTL1rX+78Eg3xjxlky28iWnxA4QbW8TZ8Tswv7c
g/1OC+Xak91k4Ijs14Mnffld4kVNzKhNd7J9O7DDQ8JYwqXXv37PjuHaFrhtIVkPYDECH5p4s63p
QBLmlK3tb9iDrtjDXGw4tEaKROSllX72SFzCGdTHm/t8SKMGNRwIkPfeQu0ZUTK9vUFcuvCcFSdJ
WXkZnb8gjITl4/VTqcBMa11UUUc6ORHiNF747SRczFWItmEg/KlRjK6HyqjzwBWTrVZ7Ps0856B9
42eKrAtaoqG7hujctwlO9SMcoEHYwrATR0DUxDzuiJn5TVcpV676bRnymExazo49D8Ykiq+DpBnX
cI3Q764QyaSXB+/wtDkSstKcWqTSJ6hM/Pi6orFXXLci9J39RhR4mnwoORCxvnhfjINwmkcXJJMQ
v/zGk5rE77Ip9g92pM8dJrXDs1wTrf8Ka491RvHH0l/VRTauoWiIbinDKaqIKp3uQM/blwZict+u
FKvKtnN22bu8Dq/IxGu3xjIWDJHApREffSAQZfG3p4dNBgndb8BlRhYfG3HbaxsWa9zUgW0jNkhb
KGndaAyhgcj+aiRLpVR9aYLoOpz/13DsYP/X/8yLK28GUgoX8ZTuV2o7U5OAnGVgzW0PGvj/vnSi
RjcHoj7TAXmeY765oRaCQ96w4r1UkxI9xGtgDes847CvpXDVLi4Tl2iFTA/4ToOie0XVWjP3Ha6k
eD7HLALkSHym6W5sh3ea9mzWNwJZHjfBtFV5aGLa5Ejsy0vwtd68Cv1ZIqdzbytILij4ojQFL0RS
Wt7fpX9ZLA97zotltWhpFm1ffsCTXgt9zKEd9E44Jj9+KNVwaHUD4UERdhk+Vq5jrds4syEt+E3R
UNlYyTr0uwcG9kMWlesfTCzq1VrMcXkfmwV4PpHhwxPtfbZeFX0TsAWGnIcWNlhCjfb5XZlJfxZI
p6TgunjXGD2J9xHHi8FMjCVSePf5qphDmoDgPPhMr9Tt5JMP3CnIbumyEKA8/Xz5A6fm17Kp0wzn
ZBtbuVk4T0YGvE/TL3fXozHt2qWw4/seHxCurnH5MLaH1XXxKaYzbAOK6/9g5m4GxIaZB0cm1Wh4
rIPMaxdfm+5ly1LuVaBec2LDF38Re+JLSTtW6b/Puedrolyr1utdL/aVgeOPKS14+uR8hVIMeS1i
bDMzeMO0s1/tRKselL2OEMk8xiuQlgXiEn6XqQQ8pJZmnCr6025yHDRPKnX74cW/SNS1A0ILR7ao
1RD/fo06KPMvLo4es++GFsetZXbgcxHoScC2r8itA6/iF81HCDxrX8HhDpTgvT725NxpCAAxgc0e
E9fg260wPyZMpSJNF2tOoamOVrJpx3dl30IcyREA8BV/mnPGyqcHN4jYkPd36oCke88L0I5Ttey2
nyNrP9LJ1o/UQX/HSAFWz6EHAmC8ibNqr5JRFzRzJCRm72NrpaloCtAScJcnJlbhOS//UBadOn5e
ICwaqXX75vrK7xrwuWYARoiMdi/jm5j+umwPMWJdfHv6a8XTVCHdRKOKpS4irtKgoO5W8asPjlJa
z9ZSWSt4S2XKrt03Nbv4Cm/BXAb1zCqDFMXSEaWmFaPv4CEKf/CvGljTV8bSl9jeybvnLQksh4VT
Bs+gF7r9f4oasgdmC29w4rSXyFzHA9g9mLmd4bWSFJ8VN4fYC0pQj4NorNntqEyRcZ6Rsn7LuC3M
+yopujEqLLRzuYI33Qon7C7qZRS659vcOm15RTrN5nDof+LIvB+eu1HQktEHVgNat2R86w4RQM6C
KK6YgJhZs5qi1a2OKgdiEqfKDPviNZIx9pkZeo99umInw0ieC/KRg1y28Eut9zXbpIfjc1+AqUqZ
xOA9Kc3/CajoJNQhWAstj+HmypZoudyswxMYjYyKKx5ibY70sSUt8gfWBOZ8Jz2xU0UDK4adZP5e
8jtn/FZl90mvtItOiDFUwv7LNl5uzLKI5h86aLdnBwPlPbh34EqISvTTQuCWW9i+mLTg3mJG02t0
sdoWbEGMq0xne8IJfh8uAspWOzGQKn5r/kwPVhTgD1pjv54hQ6Cq/jBTiABRbKd4AdUfpPT6vq38
Sqc2szeCcySJG9qbVSchklrkxpU9v0din1lzjGoIBL9+h49lbvxHR5YJhVfAZHEboqlC+ldiVa75
0aFIqizbe1cr2sH5nGYPMfBFAm69oa3ZQsiTb5UQBFICrn57NTDs6/GI1ucEfu0KkntSRrvwGU0w
6BRepMwQOcYzCVrfoRVl+ss4cg03EMdnpE3WpjAXoMFDolJgWI5NFN+ht5IZph3uZbilooXOyFsy
7TINRivPXgvM9stS7kkrs5rNCEDUIuXwUAkVkviabp8KaPeUXKZVC661WHpeQSq/n5kXZf5T86oH
EKPkd0lW0CgZYHa2QirkaPttiLsuAcUOxGtiBq+o8R1cqtCddUvhyaLkAbYBwKvvgfw5rSoe+7Di
0omeUKdGQkHrhMvkHiEOOuuy/IYfYaj97YO1nAfJQZHkAorH3NptSC1/fFZn1cId0DdD8oTpx/t+
aR/hDnL/vXXzjFiKbDz4IO5d6qWqHmXOiIdP0Lwtt8htzkViB+PdANcfkxj4EXigMQW/Xcnm+KaU
FskGFi4DKklsmkv0WcwJt3HdHrrvCXL+IUzERgpYbMJs+O1nIZQYYlJmDT+RIAXBJy/9U6V48sbz
BZPXVh9fVWoGLpRN1Qpni1Jcmk3TJGkPuDKt3LX41yoUXswtJn/dO4rExE0uOAH8wLrT8wdS+sCV
71a7uVighCEPYqIVVUCesIOEitzbrH8/m3PevNHMZYVNlk8zuIRAc0i7bZ8Vkospd1xVyer+P1mz
cW2hQrBCjHxII1wBMxQkbbVNgZt+9G8rU3y2WPCT0rL2Wojo7AwL4NPWI4vmIggBm6nFc8uGMz+f
vH1nbWMAv+CI8sd7pPHnbKjZeAt1Yc7oYZHtePHNn/zOj0IjXkDqAHOE//SfmFIx2xBwvP0cGepb
o1hEApD21TCBkdXnW8DySo/wROXnsnii+yASMVg3ZLLrunG5NNQM/CUAsuK7Q4oQPrK6TQQB+jvi
smjPaZDHOrK8FFFWXTv8IH1bADzcgawBxemc52zt0nAOixH81XEvWxKaVnO2W/2ePs0/H4ud9oKw
F8DIr1mxPAmfQ2mrFLblyZLWACjlAUrhm3S2Czgu4ZWSVfrtTkG9Ay9gKw2eNggtE2VvvzujJcbH
NUHEF6wHxvZ4tLGtLqXbBEsbXe5qyc36bpskyw8QTr2dOtD54k23ZylsU/hb7sm0U2XhArWMWKs/
Hpk0iq1gAfPfUCL9YRKc/o/Nio3ntMEIY25H9ZVED3JMuKZk5sNJizGqgDUkf0uYW47cDbMbyuVa
haAtWEOZp5tBDnjkSAflDEHreyHApbVn21bcgyzPnIaghPVJn4tz+uqjl4sAHto+GEAx67X22aFm
KEhHiLzI6UekJZRc36p7hAWC74bvLVVkCwWon43fOswXPbMrKsWdDjpDD/ap9ClLBai0LGdclJm1
uI7Du5e8Rw9CAVW13o39SGcQQCKuW/d1BLXIV1k8+6inX+l9rqYwIvKv4aFvrmPz9gEZndXiqmqH
2m2bKAvuIl6HihUaI9hI5eTnMW3wr2csu3CpYrHlvj0NjYK6tfAfyvw+iRWv2zkaP3MGKruI3t4J
FF4K2O2szOlEKV7jw5fze7RiOvn2jtXCKoexqqfd4x6aDVZoMdupat1d4gYvlruJLE4P22Hqb394
kvEXxNl/Vr/8AoEQmEg6X532ApnjyvTJEcc5feAV1OuEF95vXpZwywOOn/1nDB30Jg9XcLTYIsUz
VEAqoXI7T2jTC8HDrj9EZxj6d7QwJvKL7WRjjzhwDGFmva2tP3iJ3jCYGlqEahrE0tkHveMe+syL
W5EJXUwtSO+l5/iYzqpeB2Co+MiurhHLUEtu5ubHVwAF2MMs8K2iRKS/9SL+JLEtvdP8LmFMcNe+
JKCQBRlNro6d4pI8EBwslF27xI29BFYAY1IiNo2trcYetlMPpExmapRW0IozrDtv/iVTgIFyVaFs
rZ212uqbL2iXODJfJLL5+1lpJqu/pUmvqLK7RwbGD4y5mClGS3yih8G3Zgn3fjQ8ySfT4kDfrH1y
3DQLliuveOOR5S5GUMPKG06pBWRKBt5NS/Xz26ShMrfGDBWo0FCWj7ANZswHOJfiz0WfTCzuPaCG
RoWrfZx6O5cZdmOztZRwF2gWn/MvnW5V/WRk3c3m+00/mMSoXk19l1KUK05UgwjLMtCO3YUak7Yf
KIpozmyrOFel3Xl3wFO3wzNBLZKwr6BL08ByvnHWjX+frJTCDNMxVLMpTbCXuT6BolFBFUobz3lp
ED5mtzlrcfA6SWwQ0OPU4znm5H5KrUexHsnBsaEKfANdRQ5/rHs/QL/ZDE5btBEAcikbMF+acC1R
A5jQ7rM6rzbYEsM6m0aVOixp+2soXmotppWeD86gimd0Ox4PijziqJfd0pFk2/JZx4lDqOTIhYHt
yn8JvmVJLyh+BYnO5umXSMNopgHdpyBeV2oKyk4iEot3vy4qyBVdcadvT29svJkA6S37QaKI5BUP
Yltp5OrOSiLVyFxumx8UCNe5gBjGlSEXf2e6Ur1K/T7agNVUfH+3f+Y6nVUpucnNUMlQGUQuaOMv
KI4B/Z696lxa6esHh+4oJWuwVbTOBnta58VDPMhGLsbohKKNIlna3tBYNPkNBRetaU2XWr42w0tp
I25s+mQ+EX8EMbLkw/AlbKvDzA+rKSCwkwnuNWvh+a1eKeeW19NxlpEFW+h01DqC1We7qwbMHKMF
JIc18EFuWc3ec6bKDaTnkdHlvfajPCK5RvcZscwNb+tsaadWgviYL0D9sXedaaR1Gzys0pM79ps6
bWM8BeDThiUIOZSyIHBiZ4aJ/I+0evXV2E91cqMG/wvv4lHeXvpYP2Mr0lEWZaDT85sBab6Pt68s
FqthJCyZvRY5AdGx/DH+Lj756bWzsjEca3pHRZ62K2GOxIXEBAx/WJCVgzsVHs3viPnXaMOMuhBG
/tOc9Y0CRvolTtzu99Ngc6LIvSbv1Ifcy7REBtOaB2fP7V/n8xCWOp/Hy7qtLTxUSoSuEXOSTsQu
R4+ayC8nVJVWC8XCs7HWQscwLzGxjivmPkQ0qAiwi2hAD/2dRRJGlhUHGFeDYgzT3QvRYeoH3IN8
igyBkASwH5O6DRgJB8va1j5M7WPrb/W5LGMFBBSyDMWUexrnA1EW16djwjQK2ovw/f3iXYXigDvn
SieaS7+GKtDXleoir5XuHujU75Bb58b98fsLEqV0Aq6/oFyxBPvy22/CfjsO1axlxvVkcFayKzjI
pXFv4KvfQfRJx4KuDITsWOVQij60UFuuFmswjigL+X6xv7UTmKEy43vL8zLfp/Op5rWE//Hzzqp4
vkl2wrbq4NhnGJJBOxZS2RVnqAuPfK+o9IVo9cnoEhfj7qpUfFLLiikYdpKFJNie1Crs0as0lRPu
u3+XamebJliyMdQjiLV9wrDBnEEmCcHhnjI8JKsP+nssqfl1z8SXKPPdHa6tip4reHl1l7+dS5x6
ENsN87aKucUfS55yXuK7kzJCvEb6QdzpFVQNHwipkjkvmBSJD3t7nDFjRMt0cDj+is1m8rYgxWSw
Gd83jZUsFdgW2lwrT3VeIbreT3uaCqOJRJPvXxCbuymoRX8zHl/CswNgpevGZvp9mi2TABZ8Mf1c
Pos1h1KYlelfwCiCBCpTwDIqixi6L8qYnkjhwVohXJPDGCOHuwHXMmpJNGSBo4nAt9T86FIKLYxc
Pg32g02FNXTllOXrNNIRl3oetv3wMBiPj5C8Na9UDrQntBHwvw4HoaDpDQVbR/7c2RLnhrGaKmV9
QU5hjEryBzQN5ndNiS+Fw6ytvPPuGjwDHEnH/yKhMLBewoqnt3X4qfDKQxLGwGrJUA2GsNoRoohh
cb/0TSsR+258Oa0juP5Qi0lW+4DOUKnmvTW+j8xTY3qayOStKWF+A97xUWwt91KFRpaxKgbIcztW
bBSvLsv0gO6GbWRtvUYGhtowk4kVS2QPA0oCPww8oJEPSJ1EKjQ0xqux9Yn2Hv4tFZAjHtTKKpT/
bbgcYdRufuFWwbN4V9mVf6TDELA3yVkOKXNEsKwvx4fp4sesGH71UpchZFdhgfzHMeTxkKFX9N0B
5aCm1CrlXor5CbEyWLm0B9P0OUsPpxvyRj+qQqOjII6AxF6RvBVxr+xwOrsostruw84GVjRUGuRO
ZPx7yBNW88teO+oCcmPhq11lGPHqEeYZ71HVnNw0HnTcrRs9NfgBvEMPsBjO3vRO2y2Wo11pR2yZ
jPSK49ErIvPF+Ev2Hklpq3JuFZrdXMeRjUe0ei/+zmhlFFIHMyNEI2tzWjP2Kob3SFPZIhwhIaMN
52zMw++V4/glcaFI14znTkpx9O2OQDOXn2ugu25XTE5ZOADgDuhEXtFEaXToLN1ZgW9SPvWnygZG
VsRF1ZTsd3SwAouaEUVbkXX0dEdtKLjmqv61nFco1Lmz+93QKTY96ofbARyOE2KyAZEE4SRkLKNC
Keb2RRu8rffay/jJdnhVmGSxfOxb5zoS98/wcw4HlVO4L+lIQVHnZ4YU447YZgjPvoF5IDOJ85nO
yYhBmbPQS+Tigf4td6Ad+Bv1QPWiUb25mslhPtxQueyrnfzPBbOQEEzF1tARk4oKKD2RVZeKkZ4J
W0iOlXnAsiRbXge9hoSladu6SRnBpt14y6/QwM/ANpl8XDcDNS2mEZNgxMCZcSkyMmKvrf2o5fSi
VnxCmuW4dLjmq9lmhNZdvGbyr8ca6prMivFpqls4wdx4YrVKRh6669+bBQbKbdm6IBIFJDRHk7CE
bwRH1Im/+uxGDrMtAZV0b7/4Ff4kciI2jzel9M+05SVVbSb6PJZfPQq7GfIxKdGk+y03DOMK0jXx
rbVV2v0eSEkxSIPJac8w3FzvfOzhFLuilBgixA+O/EEuii4GMHLC4WBoyQN7jpSqeMfoJxJZq/EL
hmBPgoXRVVNqFJDGvwaHCHWO7JJcA4FVau1f4P+GgMDY8bbllL+KXGWF/H9QDZSH1Tnx8R9QrjzS
ISaCpHPSPFfsHOy5dE6MnU+eeu1eIjzoZso7Nk8fAmSe3no394FquaO1CLjjcmpTB7MICaKg6z+P
27M1kesYupy5arEAd/EVk8tNzSEtNA5IwZSgtsVxxvgyj95LQLTRTSo3w8s/iQ0YpD+G5WIJGO1s
9ytVsLCYOLgGS4Wwi1Ov8Zo2XSKs1klOY7DcZYlq4AEkcJy55kc+fx4qun6BRDrb5mmojtvoPEda
keIAD1/CxN3x3DsWL3uls6Vp0o2ijuBd6CQeJjrRa8cZfbz+g8DZfZrOg+GwHV0tOCx/z0liUCG+
XsfWo6XRCGDZ7D/xwt3urZcSyJEmPljQ6Z4xetPpgs9jXtzx4Toecpb4iree7NmuwR4iKrMqW/TP
piVaQBdD7aZtUuYid9LtDMQdFotrrUrjvmr6wupOmCK+A3fzJuFYIZH0bRPy9ZFxGK0yP0CmTdOk
CsLw54GpacsxE2YATDEX8BMuo+mCdVLw5Y//GR9pDJ7f9DK2xpgn4gbXU7ut2qntKDYSZZ7Hegpp
5Qh/fYzJvaIB4/fntai5Yq0qIdMjcaFZxfrMCDnph35Q6WV/3L0xyyy+xvv9he2G39rOqv5yXEhX
QOgekcHBjZkdtlvt/YqTY2vhWuyWOnvmim6eJQGSPzOpegtTvdj6UvdH0zhMlaEUc0rqCdfjaGEe
Ykxvhe0mRu+WiN0ydqUVDIUmpIFqUAtK4ryV8N5Y+CspgpzVNwXb+gYdWxHpd057kWIqncmv15pt
maIwYTHRCOHqUYKVrv1pPfUYvRea+lZ9ZkGdg8IS5Hf8wRDc1VFyUmdo04kHSo+bbj/sVkNSVUsD
um4PD1oQmMkev7Gxd92lwAV9r+nbb8fOq/n9MHviblhvmkRrmIGeeq8XgwloYOoCR2XLXDdnXr0J
+mS+3msHeEug1SE7sv79yaKh2XADMgxAailXCSOa5ZJAwAfP2EdtNIayUlcB4N9pRr4iaS9Lz6HE
r7NnI4L1WQi7OZMGwfg8L6CDFQbuEpJb8jLwC1FY3bp6SnpD+PWVZRKYCO5Z47Yv5WdD1mcT0ziA
wEIpFEHqBOLMqAeO6wEHocnmRwR1ZGny4XABdvWHFPHzqngnhWCvH5TKrZQkyCEZYXqdPk09vTud
yhsa+S/U1ceSsWPfLtHwjUg5v3NS5rTH3MjDj1mW63fWZBIP/+bLh4/GSA2wIg0IrUkHsMUW4qqU
V9av9TFSem8HlboHaZZ/eaA2akZwPQQ3tNCAvS/xybACQdY4qxrohVhx9h/0YUTQbpR0Zdgjwpr5
Auv5RcwuWcZq7QxkfeQRpQecv8MlurvNX2K7a8UcF9tAwpWVkb3Vw2yvV9wRlI+R0rLY8yszL9Sy
/HIWf2laAfk71pVnYboHHRgWNsGQtOl32/tJwntYtQVA9u4Atd7OT5N03L2g15As4uZEWUDCHm+T
QplRYCwxf5zPYgkhJJ/8z5aOn8bz5IHNd0RsEvILjesiUNnGxBhwL4bOXO9a3Cy9A5VyXITH2Qy2
zAuysb1MmbSd+cwLwjCtjK5k+jaB201FmQPJL0NLfZo5kNb37pl0akT681TEFRtwFnA8m+jsjiOX
LUF1qw0xKgnyO5dZOrYpZBc8HnpLxIYOlqZ88PO1BHCAbZx/+NfiE7+Qo1lKxVvVemnDSegvPpp3
JUPOE87lZQZSDCnHQDQJUAAyFiqSUXWxAG2FKEvyWPv2LEPHsUZXLVUZMVMV/akDJ1/UTy3ZgjNK
ZCgZFpcUNmV6u2FWGtCiRlF0WvWSNZxhh/x4rbYpvjfLfBSc55jASgpACHX3smsNeH36yjqyfSnQ
HtWJhhfqNpSIKLtop51STWgPTq5wkgt5SB07TScEY39JIXi761B1mbilVg3K8M+eB2m0DdMa7yAo
QFV09bg2+wiENzaRpp/9V9uK6vqt8zu72zxwxP0mTFkBNt1J75UVbBVRXGs/tuuMt/TFICsJmwdT
b7xGnyCUH+CtQI+lJ1Zt50IzUQhzOW2FNQr0/VYTOwPSHHRRW7QubeWEuMHx4pI3lPXphmLq+ISr
LhLpXeukqWHWyKD25FtqnDHKts2lNnzqHEIl5TfR2WrkszUGD9IdsWUGtqnttqdJrA8/QLdapylz
QUBVF/uyzCJLdiNtz8VfJJUwLaEggbc7N3k1TT09veZV16zjGcZaqkBoOJFfz2o5EB8Ns6NvAemT
RpTDBAsq6aKp9/L/2P2VWuLI/Jco527Yqmm8jSVwpifSCziwCW+j2SvIH9HGKijzkztNoSL4v/u1
/Pym4vVmnahov0URC2s1pfaBcAbxIhYlz7MzqNeqrfDS/E73hMSAyj6hWYNEUSbEsGFdwARyTnjZ
34kj/etj/uEHgbycDzm+XJppoSU8gmvyI6Orh5e7zctFHomOlJ8QnXbLkBAvjTNdpIXYaan+bSlG
ZFuJLi3b7IHbquv5eua91YRJhXaK34y6mIpjhBESkGSHDz7yAuaPY7bHm2rEHtDeNpgzuiUWcgbl
N6TUKm3pY112jWnC5Tu9ikHgOxbXBtZaMTcv/ypQFPukYTUvezGlsIX6qYYFf9o/ybK9XJJLCeAb
UzV638FSbVdFXeY88MoP5LKTUOPwada3/Bad2ht+L3UNiRzx7e1rMcXzsPkAuFuqd2YnowBPHL33
csUdkbK0f6QYaYHmRTlzw4XsnixVBUFlzr6a/YUxN7LlUUJxLPq4UuRtJKHT6gIZkWjDmBvp955n
tCyP4YUhMUjsFwtzbKa7TXfyRyYfMeCLGFG3DEXuMG67UmRc1KB1IdhHtBT2okWSF+W+cb8OkTVi
lRMVJ3sz18C+VvTtKCH6ah3h8+3U3rAUot9Vg4SjxozIL1bjH7wK4k1HZjc8hPUbgiuZhWZjMKji
bYYUTMTJ7ekSDfZktSpeNBGQSF/8TvfLQzSLdz3D258fZcPqP80351IyQO+L43RfqvfTMJySuoXy
azg27CzYBj+MaOQLQOl0tAgbBlNnTll+AtFXVQiSzeAQY2M2gCnDGBJ1RX8qLcgeniZsElZNr0n8
thsvh2y9XoVwy8D+ds3vvDZ2r+Tae1w+YT8EPrsRHr884mrQX2u8/r5tZL250Fs+J91iOSjCjJOM
ByJNXHuG3S4Q7EsKbc7YYaHAcUiFxC9xkCYUi0s1zyRQqeBrBgw9CT3RvrL83zR8KSrvQhqJyGM0
mNmZC658dzXM98iDS93gHA8CyuYN7XSNXJogTjzYw8gPNZJZjsryVAUO9ve4RBtm9tA4qHjjsvsb
aMk6rmj4dTO/9rqAR0j6CbpbzisIyymjiFasVX+N4/EFk3kH8osNebKKpw12KNZGg3uq1begodzO
BaIOls2wLWtcA4Bt6JXqA8XEQ5E4NOYBFabOskRyyTxBlfbK9nA3hosVcA/f0IVRjo2vdogddgrf
aveWgznY7cMLoxB8UGFs2SMRXfwpB3ZmG7igIdhEhYf6utSxw8hY998nAOpBJxTxssrE4B/xjmGt
vVd44xqzFEOdIol+ptnAdt3CWa0SY6WaTgwyrhftHTQhdSH8ZvyRwf3P9+9HMKx9NNn7qIF9LoFb
qW8d+cPLTlsY55pigAuHOiX3i6sTU4ZFYBCDktcy6oGDoUKTZPMJe7qtczWq1fyfjw+L8QPMrseb
vxl4dINbxfzKLZGN8EcOVZLxP21F6dyPlgbKr1cDCr0I3gms0+JGQAX912DkQK8k2M1lPmyUOgSV
cSPt+gwnu7lL6dmvX6Lbq7P7X8cplXJaVwC0y3fvp38wHuy1ia2GV96T5XIimDwt+PPW8TYphlUO
XQBiTEvEyZXwgP3BbPuFQlCw+KfpXS3vZPtaECYm8R8c0qWrVQYnMO5DKwcTbq1RAVhYZvywPVJ0
i730vNMqdb1KSHmYoq3NWLZyDFRYZi7/bj0h2y34/AdMvyvsLhjRuFpSQk7fdFk833nIXjuwoW2S
ZA7AGe0fUqcxGZZgZI0ohdDxOBOWO2aTqT3jkRGRFQH6pW/wWuunRcw/Ynxi2tqpoU1dXPWsZXSz
SKQ9+Ax9O39F/2vi7NyH5PjWjVnKKV2GDVDztB6ZhoKsPZRmmY811EeoTvYFVeShbqmhyxC+9AxP
UY3o+fo3L7ns1DJNZPsf2EfNZl/VoJ+cD8vUr/WZKV6kH2FnsM9r5weR/Z/SvzHqOnNHPehGf5Bw
O3tPhwyJqyvOmPVCKQWou7fZY++kx5IIaTabzKJv0tTAvJmaEHPMqIfeL6tQOVU9CfLll+lXRbp9
fi8Huqea85CgxmiPTbKqx5axP3U5+YXfhafEnilpcGY3txhLKEtLrINoaUtisvMieNixxRwdLPFV
DwxVxMG5g+3lLYuXPiFBGsCr21r7E0IYoDTBlaD8o3MfU/Nc3kmewyvYveNd+00CDeNobouJp/b6
C13YYgdIfhpPLseegac/3sKRmtMArwEn3+gFLkzV00N2bDtClzm6kXAlAIrcdrO7vpAgj4wy+CZk
TJP+q9fj14jOf11x0WanbgMYuEY4xYgPz9lEt++475TXjOylRpE1bw4BIz753Pkxq5wt4h95sVMl
xCa2oQ+Ox5IQeLkSUz7eXgUBJEPXrGozyeleWsFr/CKj1nNrb+e/ORiZlKvyE24VJGUpTaB33Ys2
SCG1ERCpMZ0RdNQF32Vk4h/ovi45Bwltp0p2OGQOj1yq/Qr67LGcUTWU1P3fRHrZJxOxCXer00AG
ZDO85n+eN9vOwFwc5I3fgM4HHH8xQB7jga98ZE3Ztiy6UIIfDh6YQNUgRblQGBytxs5KJo0P+DBO
OWpEzFu6HIwqyDfKAmlqe6p3JC0sm4BdNLjo8uvgJSo4Rx3KUnCLyy7IBdAkE0hCcD0tBLi2DTqU
KYMQxK4zsKYk7jUB94Ecl82hAWx9U/Rj6Cl4hww9Vc40OWLr8AiGQ2hWcrj/jfj+6T4Um5y3Pk61
b4AfC6PZPLdUSwsmOm9ni4Y8lHXi7a9ElSRCFe4S/J9MDti82nYaOPM19rYebLL7aLcZKc31oElE
aow5ten2M/4t8XB1c3dBw3GW8VEHPCUsdxlkSkM+tK5msHvTxsYkHqe4mCZVRKhes60QbtCo8QP4
e2nL4nOLFp1dXypil6KpDGv4TpCKwl1HcOXcV7wVazOP0pueU1E5tSXz6RVnshvCxSoteRPqizmk
E73e/Hzul3UfeMPflaUnaDHoL8DtVuOz7Cz2QhaCWmsL/+fJS8wR+bk0NrfYQD/OgMCz+QAckggF
QJMTDtlgrGe5fMsO0B6dE0pRq5b82n21f7xv8GCi70pnIVSrAYgL341+nLA8oSNQfejkURABTYHr
mt0/eUAD9B2UPQJHvRPLXWplLj3sbn0gZX7tPHSJBN4WhrUWRi3676oZjtxBxVBJ3AltDmj6Eh7P
RpMjmBJ0UnmcyvlzCc/acgXNd2upqRRs+zjBztWuRAOYk6+mDGy0JQl7A8B9O5UhX4RIKHyqQWHC
Bfah6modvSWQre8tc/M4TA5aGuLncAfqFNTMKHhWWGzCGUZOsEDQdmG+ZU0Q8Pub8qpvVjIPEMJy
T6xlOvGA+YNimAGQM2CnhpTVPinGRHUJfsYDt1k0Wgvrg2ZY5DORS9CINM+pHBNDFic7RhvMLPUe
h4PAjvPv9bbU9m2cnDBz0x4AskNVeA/SKEkdaHIdmaFvvu5teWteiHALVKR4iSBXsC6WXeDxreEt
h7+sj+/FGGrJs5b/yeq8e7y1jJH7chC0kyNh/+QxTZCfVb5IvVPcDz52D8+dqAorH+vyZyG6FRRW
+a33lUO/XzMF3+unjKv+67Ijn4iIrD1E6Dbf0eT/rueQe0hJSZg1L1ArhSkTYbG0a4qnp5Vl5egN
1EESQKcYUTBI8xN2vuwXJORmYzIe4FE6k+LxAfWrs23D4IzcMg6A2VSAa9kq/jhyvLCgRYowel9C
6zdnkrB/33WJaENFzFXnvNY9AQD7P6NrcAZvBaC1wU6tUzJFj6ZCa6ctgfgEZmc/U5piEuYmqGjH
0vgyxoaOB71HSnoNm1gKejgMOWxFZC652gHmjYyHC7dAb5XCNsj/jg1dbRoRp00qJzkHqTMJcK5F
Qbmkj1T+38O0gkSjVXRPQlUb1cANbwfE0X0zcPsWpXXCfo5Jw6NF+dbIb7qxalJqFnHPaBlEKiw3
HtOxtYuEoYvxiCusf+o+muiFhj3X3iEeEUCptDePhyFGAAWrwXLf30Y9zbDS96/Jor9mDoChRFCZ
3enfF9GDPC/RuQYksOXtrVbmzTO15XE23tBJN4kQEyW8VdqwfsDEIIrU527MBVF1mY1dGHFKOZZx
Xc1RicZMAu7AcQxd5nfMKHBkcwOaQGtT9ZfYm21SYlInpxsN8e5Pxyw3Zdn51Q9a+kFDVK5YJBJv
GeWZ4apY4d6eYG4dnQm1OHmMIvR12drGi7qGw2IjfHxoRsy5pQfaqMNEEBUrnmU9R0qPi0QoQcwc
5NVFFMlQFhrnpRCBeTQ8AN7xHG6gP4fARCucxtozsd4vn+Dy1FpB+Sg0YqHcuuc42XOGJnAs7w9I
rrPz3lu8rPhI41utLb0W+pAmS8EFeAebrUrgxIjlTe4ZabkRUvnGNXti0GA8Te7L5+Nku4J8N+Yw
xzKbeU2XSDRPHdB4pCMRBb7i3ikom2simREJ0Tng30v5rVVIV6CenrQPgurOfVMj3+NdB635C6tO
qfUlfJaJ9hzzIg/kFX3v2uBoSlUnCJfaOtRoLbQXFRQBj+tAxKI/XZIdDTuwNLOJtw2QpmGxrx+h
5ohv8Ehv3fpW2d8vWDW7A2o9LqzD9xqkHRNHxz4wgc1WJT16xVDUetfgMJsa3S+fGEK7+zecCAKH
+nAgs0mjsc1bz95GepDzRqjOGrrm6xuVSt0LcEFtDr681GAGH3FiZz+wBODEcF/ZLhJ8KtMcgRSY
3qacZHsssud4IFtbvetJLJsLif3T0C2S6KOToJbsav74oSJcz7klgcKIvyxOCWJpKK4p80DCrAnR
8Qcdf9HJEuc434FWWKygzH5+B/sh4oDM0ML9ZxhFIYNztTDxDyQHq7a6rD/NzuHGevaetwJGlBmL
7a77dcfyeFm2qTCRW5gbsYwnRMEI0Rmplmz6aqhjIU5Jew7FOB4q2YuRevNReopBCoTCFdKuNTcu
Ell4eN+rv/WX5FOMU/kJEO77dUOyUaK6Mfzxl+6tDTC2zXh5fFeU0TJK0rC3+jCCVJSnkn637V8p
TCX+ojoruMYRiFArwVOfxKLJ8+Ks6UCuTYuEXj2kLSQqT1WwTdBSc8liwahTDUH0eVdvcxXZ5TWl
TzOugl2gUQ/FUk/vVBMV7RklNpn1N8OI8MbPOgAbTWrl7Ha0nL1oDoj3ATCNF30JOPN5fAUDjw8s
RN4GBcksCaZybFrbhUi51p/BR4KSuHheNP2s7lGAiHMDMEKQFpS1KY7ik70PV3qH4rqknz5t9VYp
gTR2cYJnNhGo+ySbHWaWwoANuFDvVhUjbV59nNinX9lKBRkIgPLYxPmrmJB6g+xpM2xQAaGlYty/
i3FX8Ue/pNUEICa0TF2ChJM18fW/vXaskPahgjx7Jcg93Mt7QOVwXx9K7mlB9fDl7tMl26Ufy63N
EYUeSAMjSMA7jHukT0lSt65xh35+i6W7cAN9pAEYx8ib16Wyc5bL9CFh28MHbXCL6g9oXch7EHfx
e77W7dbGrYOlQ/6YjqZnCSyswGu4Hs87Hx2tQ8HX9E/zKkBDZI/T8VYH9KwfD5CPzndnqW2EiR5C
x+a79ixOes3XBU+VBLYXegB5DXtJoXGJ5MK+tB6V5w9irtIdYKLPxJKDTUN3Or1L5pQZz3QCClfo
ZiLicaTqwPDrdH47KawuXdyLryJ/Qkslc6Ddrtc4DgcAjfjiG/T4Nvk7LHPwKBpG6bRA5oOliJk8
cTyHhP2gBNkhxzDek9a5z2bZiMEK6v5T20jpkxn5iAtnWBsFOtGtUMRzThVRVviItv6QABA+3W9D
ySZ9jjB/taZvQb47LEwFUvP1TzlUnuXEvxi68FVU4MZ3RAdNj9aAgq7ptXYLQ4+vCgoK751+crl4
8/tRaaOYPjxh4nu/OKJfmS65lgXZvFqBOnCQpaBDC3vlMQW67ZCrDsLWlcssiMB8yO8j/EDswmNF
VNouV0hOqdZwYlzjZZe/UpSE0Us3c+BiLmBsAex/Wt397hlYs+QPB7R6uQY6QR97HoQtpvRu5yer
w5fQeM3Rkrm83K6nRDZV2idzL0aAf90b8kJ3eFcXtZJGcOCJBPHUyF1Bg949+8n72eib6bsBYOk8
ZooJkvmqwwhzpvzvFvBCwaNpLjftP7hoqxsTEjpLmoAmZGszQKbJJs7b4dX/035SDlfS7VHRkkCy
dBqGSbVaUT9veuu69/18Bf0rvPYgXySZUKu2yZOHfB2R+wsMWiigotl+ZCucG4lgnJKLik8qhpY3
Q7psyk4JDqUI4vE5WKdQlmNz/uhaMCnTYGXObP1Z+ZPhpYUlYuwyQ24IaCIYOA4ByKf+DMuclmFQ
/4GVgXALREu2TWJ+dt8IAchOMdf4E4Ik0PGqBL2RCMP6VnfDiYU1+71YpyrJAJVHDWIs5/wjU1iV
uug/QDiP/hcGDhgeXFviMo1Y27bUwfK/yD48Fgmqqjw9zr4Q302NDnqhDhcCsTZlxc9qtne8uvb2
mQK4lMGqpo3NnyoBO8jUR1vzqQDPtii+UuQZy974scftxhKJbcbKnfpfNUuDVaJ5vD237wyKzyj1
zM6p0YeDdwJjU9jFu5l7DsY8he+QsrbF5sEYKLjl+40IAEGO8R/nZ/zfbd1nFNuz8fTUkTNepQtU
vsVTGMeu0kf/G6irEWF3x//03ZvCs8urGtfkw7ddG/3CIo7d8BCGBgKeNOUVy4uKICXzdrMUcZEg
7AYFkeZIpfsuYA4utX4wd36uDCIskSoyYNattXiDHsAeiir8A02je1JiHztM+7EdOZi4xGqSjaPN
7qnDu39KQ/UmFdTKVbGSNqXw3Z0F3ozuyLS7TPLhXLn2sisi6NjER/Ef8Ivhr2o7YoSWrbHsEqDb
GWTUH2AKoHy8DfZS4/g0nRrY6k6/cXVjmZVAlVDklVF4dVX+6JcEyS1+IRvQAV26ejgKL8VXsT2h
FA2vhlm6B6aIjaiZ6+REMsxWpKTVtceAdQJ8wvgCTbuooq81uWBI5l6JSa9sJ14kgE7xTVg4u5EX
QNOQNSTDubkc98dCggPBU8nP9WtgZ5xoKRo6S6L0H4f6MI88bNBcHCZ+PgmZHzJT1a6xLBnS1oWp
aXx8LY5xm76aMRmUjV/n+I5wDO31sUyqMEHISSgkx4cc9X2e87txS+tFnLt+LzySSz2ZWh8gzK8b
NOuNqq8NFgXo4WiZp5jWjV6KqxiYe8wNFIBHEQJhFOb7bV0k1L3eEJmtY1uH3PpttTmy07Z6XABb
comw5tXayn0quiQiPTO3KgFlJ8ulp4WiQY87Dl2yvlcBOHqntZjEY/Y6XaWqKdREK99wBscIsL3G
bxS+IqON5HGFsCGSvxKX1CfLxA2+JAAfo2Psx/UUWahzLS2k9LnVMazSYyXWs2Tdki2KJvfLtG7h
0aaGPF7P9PzFaqqy8gHED1mRUxhRSVnatr9s/XDml0uVp3WJtA36L7NLLZZBXuZUUZkyDG9xtDxZ
bnrM52F54H7PiQ4AuJM2mRhTkHSj+iCteptC3qwvjYWWuukhhOffeEzHSloelqLKDiMV6zB+kPqz
JcYO4av8BynSCXQoH2TyVjijuSI3Uq12pHgUcFilXzjI8noidxB//BomKoKoWfLz8M7YwNsjPqKW
pZJlv/v5tCF6OSV5U+T8m3b+mf0/uWz/oy7wMk+gIrwTRhD6XiVJa1xph/fK/+hYjh02sdcgwrME
3MGYhosN0nIgxlkF0wBwIbuuxBstE1lNKa6pOVBMa5btj9GOcB6wx+oXcSoQPVJDBYvY3nr5WkCc
l0Gzd3b3ilob0d69N7rI0zHs5NOsjWGgqcwas0iefBzrBGfWc1C4kYxYlaVz4TyFO9wo4OmDSE05
rMnU19yQKXWpolhIqHHHupAj99KUzfroL5Kh3B2bhVMwWwL35UtYZk2bVPjeVJJYDY9BwLnvkYZi
97KVPcqd8aiEPfyGZDnYA2HDYGMGyxD8WUTzRbQaQp4b3I3Lgi7dX/Uc1908tbbaSQ5RhTY7tkZW
siSQCWKdC8hFOSHuATjKyLUSOmPrL/L/b1It8L8K8JPonJ6oZzk3sHiYuGg8h6k3JIQPSMCGT8v5
7Own/TG8bPaTFUSoeJo8+rvijwIFjtXu2wItijh4naLQMyXwD0Q63Y7abuOsRLB/spCKAYN9Uw2B
1IRwFrYIzPlOusn7VGZN//6f2dQcFhQysspClDsJVFoJJvXK6mb+OIjOEAJnu79eLP4y1ug3bJiu
bdnl0K9nIURnItgWMESe46EMIaBx8oQjXmVgXHJbZpaWMEYMOZdI4SptE5sB+50pYlW4RftOLvGT
+f5R3PAD/Fqu2jit5pzqY1AivEDPYs2qTrrY0hnCbufeP6ACVom+KoyONN9l5vANMXB/9tLJ7rtd
Y3K5iilQA0INca2siVBIQkrLuF1n1ejkn7G32Ebnc4+XYqURm2h/49N/ofKNIou2JlQPK95L/9m6
x/tv+vH1GcDJM2y+K3VA215demdPZrNWs1QCFKVavXtOPrLnuoPujRtYRaBMdnrggHmE/2dgBdBm
A6EfnyMiJIdMCL2tc/bFJgq7sDWljVaCzIJ4N7VqO4zhASq/G/38GrOTkvpK2mHu6MaEzCbads72
qrKCy9R0EvWME/V3Rx7+OOl/s3/anILARDFLtY2XEl8fi6xikKKi1yhfsaDGlYKWeEcljK0t5tsV
vCc2qotVn35K0lsdbpes0nSSjdhanrlpBV5vsG/J3nwEyIUMDfY6Rg59p3aYoLCrB8TI6d1ZsbKi
+46/2AvYVMY0aVbSj/G/7+60tDen76grd0N2yYMa0egx+uPt0crhTa4c7Q4cCQxlG4ooUBC3Oz02
MwPtEnmY7RZyWamfOcbvQQeJluggskSdY4zi1kuqKFdQhamYM9nWECAic9OZcEwgviOayWhG5b+A
p8u+JDdrxMXrmf4vfGQCy2SFbRG1bjhQIXXiJu64XZxXFMqCND2NML0q9C8AhAqrjmAhiGtKSy8x
1IqbV4LO2bSxOyJwPG4xFPCHf7pMbDCIeiocjVULJBvekmX6P9Tfs3ZWwmSmusAN7Ziz9f7IK+Fv
BJmzfqzLo0dPLvp0II5qIZyfMxdY77ACaTNMFnVucyhYgapFFE798L7SHjPhUaQRdOH71WmWYlN5
wdPQxgKX1+ZETCoM4pFmFqANMAK1PuBQlCczMEI5ZQVl2YK5bF02XM2ff9uaG6f8hHzHxEjEXfcJ
lkUJvG6Cdja7PDLR4wwes3o4cTWs2pXxKzLZx6TRMAsiTkhaymdePKeC9AvuGO+F2OlFK34rRofq
sFArGrSRsZ0VtnEDb83PR+5B8QuMp1AgetetoF/6TglxKS8IBjkJI7C6rgx5J1B7D9shW7KFCKef
ohXWdsX/ndRcemKuTafZOsdKn7z0U6QUITro0kmtjkdDVTGm39qd/Ra7Avd7dyGgv5GnqTys2klv
h90dL1z4mbViJf2+5wjSfJNV1WC+w9jCsZ75ugXjbqwYahUyjseVfpomTxRMP6ORtVSEymGDTizM
fTOuzK3+me3wh13ssw+Xi9wSAJ6hyWAuH0afYk26M4/ZMKbR+idaPkEyib4Vj2LhQhlBUWYnyLxV
1xqoPHiIwUwOMTNCHiJfqHYzLEUJSGucRFvo1W+9fXD8vIjKoShrMJVvAM77XqVPYBVruZfUQHpu
yFk3fvXZZ6sK+KOdqwXiWGXherbrYeYjPle5/LOisomywjtOWzC3uy7967yby3m/ARPooSahggNj
aoB+T+1z0oUuXqyIahI3xiLXjqGtEAhTdRJOpTflZWQiWXDYvlpvQ3r0yR03mp6AKYTf7x6e6O7/
3nCzpwCSKek/wzxnHYkxG+5vwSRH1DXxlUqaknrSdcRCSThvIRhYTjmeMUHNBFdr7XUXiG3kuOsg
l+q+LXVi9k1+OVhqtQsYitqBk6pHQFQXa9xVfoFsmaduMQWaDeW21IVLjDWOQVKittSE/F8+K0sj
6mwprPs8r42cZpT6Ie/uO8PmPWZ+Ko9FkNYdhK8m28SOuVztuPdStXKspxOk9egLDORW9iItLL+i
51HBur6WgEBlZD6HiuP5YiUsY5oO69LzRLeeJuZbXtgwVXVqMfS7QbPlvP8uEJcpguAYo47obln6
0mcO+LO864eIifkx+aA3dHSOxJRmHz7dGl0OXYWD6hnm+rA3ol/idNd7I3iSxiu2YxstwvQEHL9Q
PD3+KBO/6NsQAiVSwku7sGjQewtIPvFDvd+YCceXvNEDKiy8iZgsYqzqJYv1zTfLQ6x7Uo+emPI9
9ghfIeZ6eKNYT2oU1D5VUjqClEXnWVHaHu07Ffeqy4e5Qj2Gswl3tRNfbb+0MrIWryoko5MsMV/Y
Z83P+GAzTymxlh635YW5XCw9gC1QkLDBgyMINZqJ1e+J1RXMqEWvbHvqFA0kSFFzlBV9RWCN+g18
pP1ih/odsI8WQd5Ap4lePNZTe8w5M1AQl4m2+ayNwzBwCnywEJkV7qV6yo/bohtm8ixwHVpu5XTq
oOG7UMC7mjDoGoswSHEkSG33fvrnSQaEinCNI+zv/GajEvc44/OjbFWcd8Beq89D5teJO8REceTp
G3cYK65ZRO/RJFfVGup0bGFKhdEMkNujoaJMj3vI+WbQ2KKytOn60DqPzHIldEadSxqpn02+1Sqe
aQvued/PyOYCsm2SSmX7O+3J/xtd4GUWjM50OLhsgSlXBcDlrQ6hzK20CHSC77/zLc0c97GHFvth
heVhcptPNToSCdolwEq2knN0CMMJPPPnuOVXDdEbz9UwSdgChyZKEviCXfLib+WgklTKEBTnSUyq
rOXnbYbgYfj76gIVOInsgPGJTbEwsQCR8N8bdDD6koxo2DpVD+5IpBg7b2dNpgEmA/5CMirHM+rA
p+m2VMASNiJzD4gvHC4k37m3jSz7yyWpY5eEAtDfAY0s8+b8HJ1z1ugS0ahoZNAmwMImmPDKyrnk
oAoaX83jvN/I00N8dCNvG/pcShJ12AfVlClB2F2ovrEje0NE+lMo+um6YSgpDVh0G1AJQA4bw8Ec
S1NCgskQBzNwb8qKmttGYwWA6q7ewj/LcTJqPICIsg01pWOdE5rOvBJgraF5IIRzmx57qIhSHLqJ
tuw1/7haZERMlX19p9eLU1fSATz6kJ4CwdjrwoPicRRSUddZ6RuXdmq+FCws4VokxXTs59ZHXs83
52biEIztR3zXvZULJt2oQAp3MUnmn94zMVwe04OziHxqXQSdBizI+BUVrhyqyYQfH2VRkTuo9Tk+
GlVixW24s9z/a6Msj3kgbU+jJ3iq7nhpqfD/c1dvFwYxjm3aKGsbYtq1nwgB4mVSTFcGtFa/r7iB
QoK+XsM4sIaC5iSJuI10AxkHnGDPj8S67fMYur4mKPLHwQoOrLPWxRBmV6L1USrfUNkXy64+bhaq
RPH7bgyrgWpMdqad0wcRqRRq20BCslhpAIsf6ug3Ys268MOzFCtFKSZWgcNYpRpNxlD28b0BqMW0
I9GMHN0PHSMPyTmON7K5Cwkh+T3B+yuWOWtTU25gMtPNgQ7Ag3aB7PFOcn4Quky7msIkPJ3p1PCY
a3YvDye/OhFtnzARn5dIzomYqExY/x8UjGifMz2wYwaZPhIYQsidtvbm6gi0QaaWvgs6SDSyKwTB
A5KvgiXvwwS/XltIQScQXtcGqI9vsko0vuqByPjCMzW4jpdNivUzBi/xaakKOx/kKNOp6EcCqvBE
fQGrO9FmJlhFeQTx2OSLOf9vCQCkxJlvVRLF3tZ+QAc28sZTFYAu6IWiWkYvZ01DhMHLQ6/DvymF
zhgAw6CRgN9Hv/7MjYrtjBnkp7P29cwDvYLPuwjoTn5PuSou7emFPAk7hB4mWR9A1DWpuRNDv+Gm
Ge2BWUL9UqErrED0AJCMivV/CYGUO/uon23VOi6VEBuTCf6CdRODeauDuRnWZyU5E90BKEJ3DZDq
0Hm0zL2tj2b1H5QJ/pVCQI532mpRtzBfNU4EQvl/2iipfIi4qJhNev0LbCfXlL9AXGtpJZ9ViWuu
tdPvxMlAVSns91l18x8ptrCA7FOKcMNL6WJ+tVTgrwQUEpOXkLRNbrcNyzsr7Jcv0BWlCL37fWqL
t+XDFHWBtkc/+IEW/RIuJkeXJiFv2Kndi/Ky+IFg75+LqTCEh03AqOlI1Wk3PCiRD3RJg0bKpMgs
4z4k11R6dckVCqy1udM0oPCgmj/1D+xnPmfTRcyDerASgTx4F4lPhnbt6qgdLAa9nGa0zOjs5XEi
4KYRW4m/a/1Hw+hwE9KK0zNupCoOcnZCQY2X3XsP85apRtx/dOGcegEvx+HhwI9C8Wf5L1Qwlx6o
tcoJSv0WmyA3izhgWfuM/0lLm8SS8BdFGhVVcKVoR6QF5X7v0ayqtRagaIqnIH1idlbfjaLKGEd4
9f/VkIViu6kJkaZMJhnQ6PJXcvXhZ2DE/nM9ZB0wlPzY2BKueEGWXdO4NLUYx5+CwsVGBJCdAFaO
WP8vk/pIolX+fhRZ48DgF4i2AS8PTvshr6s4QPLMXwSyd6DnkixG9ocoTFHwSojl9x2cjwWCp95D
hSisU3nJEdQb/H7Z/t+WRMn9xfPbtzL6vxzM0xRWhvR96ZJyt18QbqkWiRAkUQzIgG3i3GWRg5K5
a1igLHUbfxfbMTxANWe/LeIj/h1BqodNdvOA338sDogQGxGoo8RdD2E1sBF6ikByYWzWQQPZ9v5D
6HzrlYub0+SSfyMxmpvp1Q9hYrtqg+hu4e39ZCXd/2l6AR24qZeqWgbBZFbHS29iBi/CmwVn2tiG
dTcwUQc9n/mWVwutYRF7DRh0bI48nosIlQJCCVtjdnT8pkQEYlFzWkLDhwdLlIaG7nl+fcgVu1bu
1cO+RkhmgQ2wvQLqg1R9wEijZZe8yo5ZEgxz6yYOghMEBF5V+8stXwF9DDf6f/igPHndZwD+WDy9
noVGAB3zibCXavArrfTX+iuug5v5uI5/j5S9QXeW6US2NRMdw9qxHLS5288Cq6+SOf7AcqJqD+kc
imDkGOZtMtCj4B6c4I1R/Acb7KGgHeuQrU47xxdaD2T2c8nyVfyqREqxhRZPeIR4eU07xZrUHtQ1
443+ngnVvMeJUVI6eUWxW3haL5WBtY3NnaLY4EVgQppSOb0Luj9V+oBt15EjPBBpIZxHHMrc9oGN
9f2D5MuoXS5/ZcxMlpUy5ivI3QbfwWn+TclSASpCcPTTA7MhjGzqgr967c9SNLSPgzw81Xv8rnv+
4TotCOj22k2M8swECGmnz/KW+yz4xCtDK1xpYGebGo5Z+5mzY1GuZ3s8QmgCZXFiVuDbCU/P+eLP
g8qCETr02+aqT2ARnRHeP/gg3nEdloRTiI7OmSEESqx4ER/rBdLOKsWEiNJ7tEpbwJxKsrPgLymg
ZevjB3V8qqL4XEjR6AvzQoWUeyX7+qpQO1sPlxEnMJlnF5VRLgG20hMVOdVqHIwkdKaXCcMbXK6c
wOM7D6Mepcgsbm358HTGheL4yQajyHnl8AIth8fE5llwtJOqcqp+D+4QvwdZJ89siQOk44t3F7aU
2obW0u9PJDst02k1TEkD6aN2LbFVw2oGM7TGZgB/uW9ITNGIejlTJmh+vATuDeAqd8gyV8q5ntxF
JQoahqev6rdyzUrRi3PShniX0n+D8/aVvmHhvIgE/DZTmJrsaoV0wZTUkmNwgMUXefvG2ADSRfxH
cP2YXg6SeeYz8TEX7QLnMzQTtgntG+tjHuqePi94zoLXrhd4lqynPekpZudilMNoxcy0SHtPzhak
QrhoXuD1hHJlb5io5+As1u6plBvkNjTKUdxlsyL7HictOAIiLdVz9lLsQV1j0s/S8iCbxUV34LhJ
PmDMcp/BPYZLqrxGcswUCHbwr4PTRiQL0BDJsF5okFtVhSHOOmRbsKmR/AkmyA38PD8niCW5rYtA
N95UqTf63nRnT1BJNvnXIh7lY98lWXcYhbkjgYOZdSLaDsxNMguxPc33XzyHsNRBGlL/HNCqt+6o
71vkLuLrMWYKahcXyRl15skoL/9rHY0lsUeO6G2Nxx4lzqRwdaQ2YdhUo7EcwU0rWCQElF+Ron3G
g6OGIigtl8l3shWwYNDHJvm5lIE/186nRDgBJoLpKEIfgTAa2NpPTWgXY5GSV9L69JERR4pLk4HQ
FAkdqwg9htP6nSkWAL5pssElEJ/zZbb4d/nbhBQZRXW793vmncxPSFE464QNX+21eiwBDzYPu8PV
Y8jFFsWDFkKdeZgRWGYamRCmqYTjsAurhHpRcDff+PjxOZICcHFdesrwnRLNXfPYlBtOLROFqMMO
a/tvULVXqFGsTIOxtvlRHHXlsreGsnrk2M8FIhB4ruLetBD6WaLFQfavSdkUO/qiCq0a84p/MA4L
PCqJD2cJd7EeS6f64FO6wMOqtJJY507MhqY5V3fXkB2rc4F5YhEbPKX9M2TimW/mPo4Xdwdk+BjT
9Oe+wDxQ80p4tsM+GgrIjib7JYOz2EmoTzp3SX5AvUA2coV5KNnUKvWwB84Yxb2zQLFC1HS5vZnQ
rqvJljdhh+/2q20HCEI0yn2yCN/dxp5es0oIhmUZP+2O541FzQ3iea5A9DvEHDeJbjVH1ORNLFZI
tyZTAAsCb5yK7Ek6PlQXX99pHzE/UXiSFjulAIdWJqHi96LNQjpEtnqX6wAHMdxFmJTmv37WuyLo
1IBp6w9IDUWY/R1qRuwUTqdeI8q53n6uDKHWGhlcuOPJOC/s3CamFdsnBVkb8SWqJJhk5fBHTaoi
Kgg1/Yd1cyLYYJHdb6yVkwD5F3obgo4U8m/v8elkA4ig913ux2pSm6aCsnvxk4kvJ4hquhIwomj9
jXhROKIEgl+OtI0pDBpq5BPZqrLWc5MJF9DRUjYYz6gsj8arVETpOBiqkwu/IO7Hy8K5SXkJZLzR
F0BMcnZgElRfY/p88yf1/9qP2k/RoXIO1EXHnstkzwdFO0LrttIK56K8/gbyIwKpvRa7I3FXbj/I
G0EEk6Ya4x8MMR7FiJ2MAGigpyo7g60bai42xhDopzmmH2diaFW6LkGJ9I2hbroJkJTx5Y6Avyfe
uZWXZEz3QSF14XJ4Wl4xhihUcxxxN12qtKieU1JL+Pn3pZcby55o9zvL3EXS/KKtzC75fwr7sAfB
OXhu55Xjqpw/UBNmYGMo2HKV/KOmIoiil7GjYHOQuAHWsZBbmTkehvyZgsL9YqyD2i/lBenh+QZR
CnY6OwuAs2MgWWaq8WhK8cjE8y4lw+34wx/69D7Z1f+zNseTA9mJbcqCSu0CJKgnKWPQazENxssZ
48cFAWwTEnKJqU2ASyS46CJExoKy5WkW2pZiZGzEkdbbkkl/XvnIvK5glTjt7Ale5/gfG+yoXowb
RPBBMo9dacnerRER7oVBMpRdj+ZXcmtXuDXdJ2fwGD4L1Zm0WKenTRowtE1E53gwn0irQIhPE2hx
z+kCRerRN3HgLMpRzsb1WOpNWoY3/VMoF8Rh0sbjBuU7yqhjXB+sti8qMaCiMA2OG38SsYygx2Rj
oZcl/hClMQac6IjOYgj4HGZtkKKyEby7fw0i/I7+m9NqvNRNOSaBItmJDrG9J9JRnlhGttmLizCY
oXVGNc4WtrgiInYhav4PY/hF+FmRLiMdXGqncQlAFGsKRUYe4HqmRCPeA5l22fBuXLIkPGstv4Au
ihEHLeBwYCZFR7z2rvHd7NYPc10WP9vsnG8tRygUVuaEQiCi03JU0V6I7LdL+n/Z7Sry6MHD2Nrt
da32YmNE/yrRTyQ33lCC2UoldlZkZ7w72oyHh6UF2cbYDR3Ihqx/fvTYH1sYorzvFrTHhZhvfUu7
7cCPIYLbH/H1oGHfkuqX3pwivFEcztTh2eAAWUk9z7NrnGzgkkPHPGSwJXcEwD/VlMTNvG7Dz4CT
6MMmTtLYGvnIa80yBc/IGMJOGFZyRV/QXCsCE2ICAXmRqYsug8pjiaCTQoGm/Zw+BCVcg8W0YTEJ
3tox/rtDT8/JxwzkptvN5PsQoPiat3pdpfglzq0GHFwf12iWzu1hNLheKMtJiXJ+dzkP98ogfxAY
SXmZ90Yjx3spSZZeLdxkCuekzD6YwcRXxy1C8hxITa0/Z9UKzN5oc/vm81BARgHqQjdf0LduRCYX
1iGe/dwPy4y8ao9//47Ow+oOH0eBKB7S/nNaersofH2LRt+adAf4/G5rYO+KhvVT9wAUSke+Q9cK
4KJOdlDlbWoIruxXpCphp0J9MOqoNuD2hhrEHb2FtYAj4qhoRhF5LPmakJetTp2fAqygdQw1sLmv
tcZacl+uO+DIyzetkYWM570VNQ2HJXdeY2sb6VDjCfXQVlM1s/gk2ubiN6nuP5Ja7hhEnvaDxfeP
x2BBRY+96dx7PEc4Cm7vWvGEs9PH/6tOFA98DMTrlp9o5lrp/2qQMKDC20UNZ/Cy/RPhsXQdtuxW
GOWWcElsfqZ4xDDcW5PR8GcV06r8TfEYebswJDk3ogW5/l7TgzLmEOnQK30mBnhwru3Z/ukiibCh
sqJ6CsGzGGihmpNBDSUeKW7UKjxdqsvrtauYo0DJSwQOeMHQQglABUzcccovL1WiB0Bzh8qkXgqR
IbNkym7otUH6x1QpHZIT8L2bIeVl+kNV9AqhlsBzlZDNxL2ZB4+cpjDM3mHztmABhIV/mo1H1+ik
3o+ZUl+gVWYPnEMeVayasBqx95ZNu4mb9z+c4odnGcMXOb9PEZVEvfMZvwM4vgCQUOy55e3SFN2w
SIgZ2OBd4JkPla0QB+NVM6ZjJULZoDmNZN6t2P1d4Rp09z82EzFvESSNakDxKDk5q6FtF4LIddzq
6ZiHeUgVbFHcnhMjsDAGQiyobZdL8FTEwu5s293xlLVhz8P4bHUhx26WupxO7EsjUM4hEnEGjmcn
mMac/aXHgsiLN08u6FNOGyFqVpBciufQRupuuzGgdvRAJPJ8bT6aLcd1zxA3uFioLZavri6o7/ln
kLaW8K8G9vnjV1NX9nSqhqToFQm5Ar94Xm6AajR+UPR4zHnDh5bbccZjJXtQHbc0+qYJEbiGIMEn
NYorOLwnAxr+DO/eM1FdfL9aNJ0Ua3blYnzzvbNHSCU8sVCx799sr+/RNAAkSAYtAUrme5iSV5xN
DQ6a21iheEDS+W0cMbxPi93QgSPndjNpqPwC56PlGdte3p5awJCEmK1RlguQE7Tl/epxzzR8PNz8
5Zhi6uU+4dr4V0z52L0U0a2U05HsiyxrCPwITWgVSCyamNal4f8o/ZBPRwsd/Qzkw/FAM9VyqL3V
ihBi/mdfto+zwsMNyWKNM3LE+rlto9DZUZgnqnwEkvtrMcd+2gu/ZaHYPczl5Llwy7CKmmmjT7N2
hm0OFg5CDl0r93B3YvOTGHHK3YTK3ART/WZ57cuNyceo7ufkcheH6bUcCyV0Fb0YEPGDXJ3mSZtr
+TgeZnsx0RCGtA5qO1kxgA5JoYSYYPlWQOnq5EpNbErETZcmDFmV+5nJPVHuZApMYs3XFf9N6Bda
XjSafho7a1Lhz12ISBOj56MvZi+/sCRY5o/b0/qC5tGH2c8xHyTUxzgughGSqR/1Eq/jmZUGnGwU
J+op2jQSvHP1cXn2sVrHo4+9DOq5n1Bs+odpS+bkAmQ9Eqhby8Cx5HQXz2yYZeef1XILVN2PglEE
jPg2EWLg6cHV16mPpQdDu0FG3xMyatWYEAqwcNDhjLRxbqkQEuQXYRGXXHzKXDb8fqkuzYTbdOdm
2ncI+oSQQoRcDK9Z19yRtKGKTsE/ip8+3yxTG59RRLacWwd7n1jsZk2BNPMgaiWW5ysd6v37KZtz
SBBPuxt5/hx/n9G6G7cjZiZFTvEIceePcMb6LL6ockT+fDttdYj+amWg527DaD1phR9/dyoH8Fu6
TDhurmr3E646XONkDLh5HL2EGudyl5hv2dLvyeXtC4FnJZ8mNEqgRlGXxqEorYPeP+oeCH6vhqjj
Js6/gChOQ5iG/OArc4QTouINvFyC/HZ9JhWFmzNdEchY2by4rGPEmw1AtY5DwBPx/a7HE1K1N1C+
W5+FZJHjVo3a06NLK5FzK4Zso4/O8Qp+LtBx934+kKdUp2cK5f7wZOzsvx0idmZZvCU3M4Vyrv1X
Ifo2iUs7n2M13Uv1A3nvd98too58UWuge/OmLgeuJfT2KD+JUoQbGBtPvXmQl+taQfTYwGolbklD
SKHu54w8TmNnOiwvY4qCwBkRLlWQepYp+14bskk17IwJvqRqAmlvvkGjjsI5iwyDPqW8KqH6tzfE
tFjqCHSPyUoG6aqwAJMEKBRlG47SbetEiP0Z4Dim689YpRYD2GfqYln3oQbw4yuHAXimWDSZmBWK
9sv71x7zljw47akigLqgtKwzMM5YdchHJ7aZI3y6svY9qK8f7rypyAAi5JfvWqzP8PSLRlE0PMg/
9UNItmAzYNw2MkYMyAX288ANfBLLDYlCanxcUn2BcNTtwk8YFIL40oF4VG214ZABkx7xWzt7N0T4
xQ7pjSZOKpVOE5/F68oO6UgAtEkxsCdqaM4PepOxyk/zq/xUm9XnCD1tU77+WW2r/ZdHirI/W2wE
V5irk7w/un/BeQKTx4EjrIdPNLmXoYMZ9RPF17BUjCTaD7VxK8KOfxhkGvSRNzDcTCwBNZ4MZyvM
VeT6FR/IyhAvmXvHfVTtpWVdAidIuCXIRlwj5zL4a9wjFWF+vt+22aIjqJadk2VkJdrV7am5yhEF
O9lDOeHnAfA8n4qCZKYMNeCwtTrySQ42nFmWf7Xxmxkp0WuTTnSboNnEV7cjNvIDiQmr8JqZjrMV
KW+tkW2yk3S3QiprlfOnOqYz9gh26tnbK4J7mg0bnQZWazIjbx9Mx07TpK5gZN/nimF0Hr701+fd
Cd8isv2eW1zuTae1pSTMa50RLxUH+GuaUYelbyWocTR4FhNnYdBxofE2cNGiwxeVkfHFXtHx2RlV
sXqLerwCCUpW3vd+AdN2e8GWvfnWMB9sYTZoJVa8OVfhg4dNA6eB+9j6lBRfRtiX/4x6lWha+zO1
JVHQ9sxN8kBGY6GaKDgq5owbLxORpRLoy21i2B+glGSXPv7IliGhwfnKLabNEIiMR57qz5+MDbxC
2HFF9REVZFyx0DD51K5A06NKYplbjakvjH7UFeuOD0sWuRDi9YIqyhgp9ap14vblgGGnECLwyeFw
Ti3VQKkqpqlzXTnCsENw16vMXMOgzM/SrHRG5Ycu6i3COyGAPJxg1IRfw9fnGSZ2jBIg/Hkfmpdy
AX1WejC61ANZm9Ah1obdgs1i4l/s41NrQsinOB+YmhZwAqqzMgcViAFVvRN8ta2Ebp6UHrtjSdUA
JD+YYEEV1wlhffBCoSPcxUTwP3RN4I0bvJebabw7V3/FM1NphRB/DqRv+758uNLFsdoMa2gfEeyO
fw/sJTilwbmB0gx/tWvOlbT1vjybFVfuPeLT+vUlswb8YZjN8al/cTk8AwT5qX5mmj+1lnoDGqdr
+KGOZnLr+bqhYPuo3pPho3wAFg+AY1orDXZE1fS7cBWR6oUglK+0N4NqXpL1n1lSTRJVtGxdr3tj
BAZVhA9X0tj7WF42/1zM+Ssk/jZqKnoqJlCjiG1WieQX4mtHO2F1Grqg+4NEG4z5i3Ev5BuA8gpU
woMGV5v56CHy0SRdUkn7vPeoyniv26SqHLCh53lKlC7eOTvquI8/izzWwWwUSnGDCzHYbju5j1GX
9BPp/JVnUTHNrpV6TGuV8bCyKJRwue/ICM5h4yPpwG6kpzYjYo7NhEYxDsY9SzG33jEBA9a/ajUw
cfFogDYp9/HTJ6b8a93ZDRysXNZWmXAwb8bJ3P32TzHlhzqpcej/c4MPCNh+OmiLcokZ/LpeaH1N
++6TGhh03tsKR09Lo9c5RjB5xR9lXvVrG/WOV5TE+tCFCF+j6SoUTP3XgcgciYSmI/D9P+UZX0h/
OOzVcjZRqwZXcu17H2z6X+teZktPLajSVklAv+8Zr5SLi+fxJtEjHjMu/wn9/nnvrlHGyE+S5U/Y
izbHiV1blmY/aeac3HJHv8VnAFqSmEJFnqjWYgbRH0MWmI7R8H2nJmHnYvqeOpyiHKPcPDymiLgv
chn1nb4i2c6SFYm6gf2JPMpJzwmaooB/R19O7Uuvjut/0ToZEq1+Q7Rk7DpKjjWxmMGEP2fayhsG
UINA4GxXh+ENESRiIkCHLhEhQrdUjiLqa+lVTsFJXd236+8g1Icz6Vs55XlMZC+SxqvPaDZ7IvX1
Gxz+9D3R14LRBHl/9idFjm/J2ZM1/Uz0OVZOx05/anqC+6uDlJmuJggAr8kr0ZjxaBjjKAMqu15u
t5jQEaOyKpN/0F14Jf7aCqQaRhQWPPMG40Qglks59G6T1tvF4EoyBiiqJtfGtR6FgJ/iFHvxbvJ/
XvKYkEY6Ku3+KaThJvT3zZbb/XdLtxbI918CwtHRFF/O6XHGEHl0WtAOGYABFs/EcPqjcO/0BpTG
4mWbnHqDvrNObgDI9nlBxb8aLnJa6AHthhGc7gqeHhg0G4uuWFJ0c8ch/PQ0smDHHY5D0RmhjN1t
sprjG5Am2ORGCDczZhsmyY+ssemEUZwhj7sipd7ZHfdA78BBc6HQWDdH+/UMVRnNoT7qfNp/aw9Z
Bc8AHhbXvgpjWNmB1ip096eEIQVn93ztSYlSHvm54h9vtkIVTLVuVKkb+rL9WOSUe5+bOizt34Ix
mhiDmzfjC/Mu4JoA8wuOYz1Y5FQR+oKT+XRbH1uEpoF8FWYkYd0ma9ukG/MzIxL6a8SLXrL5FUiP
kzv8UQf7qca36AWi5NdPdWroTzsmLZ4a1UMR82wNl4G/E7R3b6P9Y8KaEVn+9GpPbC9GP4312au5
kOCjLI1ecfc8qlk55H7+jsahhqq01BGojkANJyz10jEHOG8OyUwTb4bSSpMHG/2DCtPU2RTmFdpo
GABgujXDM8xvek+tPfadeGoAzqYxnsMiJatCUOLSKBS6eED/ZLkYNDqTQ5V37xrmR9YRmS2Be3uC
3f+rGfnEMgt8Eo9SwJJMIWzTCQsPPkem8VxnJ9yQW+bN6Kn40/LFjQ6UHTA8xcnEGtCska41kfLy
wWgDAHv32blUlMNnuAEPJF026VFxjqsfgkK95VhsheydunH3aAasgWvd60p1LTrQBpDY068dfriZ
lwb7GAIPqpD9UbeYPVQMDt3PDZ44hRknhms5cPap34nfK09VoXnqAgy7gq5Ngc9Wlj4IZxKgcLVe
KoeVrssWHqqcpJvtp4B/Sf4Ta9bq3vxilwX4HMpz3NV5RV0m6s2VPTGnNDpUKFGs/02QoREzs4/2
NJNByMIzIrRn8dd/NRqQinhvj82gbHwbiM3mMtzPnXy8YltPIoZRzYxQbPMVU2hNk1GHiZOoa7qw
+blvOGXkq7T0UgIbUXxG9LS9zdyvvtZRxazAdxILaJlD/NRFNzbzIWOlorj4HVgBpG+S3eh1eHUh
jX0ufOnAPl3QPBwY6GQ+/k4Eq+x2Vfv9GkPw8thHK8Xg+YEkq1mM4T5zU7PAyPnfYBWIuYY6Y5Bb
MD+gAdDQC1Ny02avbw6Zsa8agt3ONx4bSZ9Qq89X3TuZEXfA4l21U7bAmu3BkyaahU8+N3IzDziC
LvDi8v6LzXmkWOwSRm1WAlKR2Ozf2p4WOSOR5I9uYcfa22fKLVyqS49boiA2Xw5+HDnOjbe/1CqI
thqoKtTozJhfA9AbRR6tAgT3Nk9uNk6oujwvw3xobGf1C6JDac1dSsfyA4WCtO5d0lGG0qT2GT34
PUT743ApR4/Mp9/9v0vPXweMFwkQfdGz8kKm2l+3SPMA/ZRH28PNbJL3mYLvyta9GvNHyTMEGtNq
AYasryPhsb5XQ7NThyIci/9VeUzsdV5jbRrZbrGwBrCz9RviYj50ki17BDH5R5deAxetG0pFFrl5
Ca9kcl350guQ4Ob4aqoBHPq/S+/vV8hKf/xhlkyLD7HGou/ECyIMqEfVgwlia2mkmYhCjvx1M2Kk
qPX3pUhATnX3sHySp1snwyXgRhWrOSoVgWUi5WaVBi5fUd4sL6r0UgnBxZN4ncqzRHiqiwZGo1es
sSVNOl/GfG6TYvE0hEM5vS/G/ZLw5sxGAf6OTL+7OhC9hB2QmJCZqBsoDchrs6SDWvWzAldNBQMc
eVpVAXPdy10wLBwzPOykfelDeoQhOGEKsHOPYzP2nrOhNQtkGUxAWge8emGsiEh8aLaJGaej7D+L
+CpFbHCl7LqdxY2xEzyKPA6NBVyeZ9bGy51UzKbmMBB5nSaqCX3/U8y9Byf3VoLuJojNxmmPNUAB
YAkFeDcSZJ2Ekcdr54dgbgaT5F9Lti9gNY/1nSIPJ87+oXUngDN+c36TdH7Gcb612VU4v3uFg/sN
5CT9B9a5HjAfbusvXKI3twnfUW+uWmSBCSmArMbxv6t/vazq7L0oyr6QASDwIwSl0LKBpscFVfxA
7cwBT8jPTNgVLqfJHbfQ40R2aKEMAq2WtwhSrzlGPaz4hcdFKNIUlVa1Oz7a2MXwJcrg1kckmUMH
04SkvlmTo6mWuOsS1v1h62GIwh8UlHTECUD9prD57Fja8fuJjuHEZOJAzvjQbmeCp3ZhAybeK9M0
MhNyqhhP2DfcrHAeviBIa7VP5M/CVwPXxxZY9CudweTlqf7oICP2lEJkQ97h/35B+iCLrkfRThPU
FzmJU6VBuZsFL4cLd+4O05Ej0riYbZTc/IFg5K4jC5OGD/gyjSAQfGccH/kvjggib+5SGT0JaIvs
uJml+BFRePV4m3cgpKn70/lMV7ZkSeXYmqvn05dPU/0LzaFEx44Ck7513dR+PCpLJkEZl2Iv4Lqt
eD3NydwciqEsJYpRhvGAy38Yo3wePsNOgGcde1z5gu3nofj+JnyAD+C13RM8EGRF01nMwFLbEA27
xg3QZ/JjC5bYsPEqBzOAqeiPezrYCxf+a6YMfs9U+qLjeLbWxLDvtn8MIN7lbEfJnly/jdhSqCjE
biJdcpJU2fhAqObJeVLnfTJrYXCGSiIQwdVvRt2bQtyASa1avp0CPUKKfN7uERcQDroq03bxFF7I
A5g9maevVlD+sMYEsAlzUkTUK73SXFQg+owyGWVFAoWz13L56k1T/NkbVKpLkrweEGUpg3o1JwjT
yBCTqVYdjWxpnnhOmkt2YlX1idYuRzC1VAtqKGT05Ft5zfWECrXdrHJoDhBSqWzCD/wCT/fhAw2u
IYjxW8D9PrSw5G6hGcg+ngFkMSFSQxy5vDtPF/yUOmfuIAQW/MbvrQlqvVPRRpLm41w58JPAV8Wa
QgxJoQoCFFqbvfnA7ijgf1UE4XD1KM/LA1wTox40ewICB/KQDxwmbYKawq8g0oFZwC88QHH7R12O
dp520VwsONY2NJlzYzqHczOmfTdCoRV3dpsKhx3N/MMKQlR5u3CfA8c0pa5eyIkiQTN2rZc6DlWw
mY5kzsZIB41fXGS9YGcF7j8IMkQdpoqrLWM6ajACAPIcNdPCMpL8ZLLEqo1vrQpb/GrNG9/LXV6r
G1Kl1Nyr7yh+9IqUjcNB25uyg/rjEIdFMxyiiaphfmIxrGQmdEV4LUgzzn78DWJEjUcOom9Mhf/n
52mKfOGVPpzqprVcsb+Q5+mcr/PkVw1fueeKgf5F6PD9qa8T1S3e0za5RS4Z86JzKOyUrJ8vCiTk
+u4epLTMkXelP/rJa/ParoDWWVUIiaFwsst6ojl1GEWKybE/uvOhoLo50BNEP3wjwvPS3xm2qqCK
GQHjUH/hBz8P0E3xRkDkJc5EZbXmwT65a2GuCzwx4XXcWPRUI5c1/U/QkAQ2VnBxElnv+mmyKiTB
vFfvBwcYxuS98rATET3LejxTU+uCw+dETPgoOsZsGtSegCro+/zTggrLRArgMdgViqUxaVRV2sQv
xO8U0oyD03Ln3FGnrHbNhVEov0l77e4b4lCRHNDaI9E7t/e1OkL0YVZxRe3b2cpwLBOd8lhbBaUN
EL99kGN4FKPtpRNIFpDuLkD5a+u2lOxrTHf/1+uehh8LVRCYH6RGH/rxpRHU792RXjyVyFIhdVgp
nnCHXynAoHdpBAM60V8hzdVyBQkVN7JSejayVl9c1v5VN1chKVo/9RN9KTf/svsdhJHFVYEflS5f
XR73MGuxG5zT9aHJSM/n//4WpExDUqzWJ0AAcJMlO8TCvuP+tvg16zUWK0sOfOXDs4Xe8DYjLYFt
Qa+sG6ydL/meEMqqqXx/nZpZCP/M+ViFdmLsc1mzNOOvIn+eaEoh0mgcxU+IcaCIMtkI1I1+GXVG
3tPpqNu5vT9aV/QCCY0k30FjrIiQHksPyApGxM6EzPHuNuzllqjQEkYTr8OBXHo9PVZxGdgLg+SH
eZg26+X6qmLiLdwOZo8oCwH4vPnWt3cCEIsHXG28Ydz91mD1mvbqgs2RIIPX4EzW64E4gR5bnTBz
bhBZLj9/crdkNX4r0PSKNEfCg2pxCkn0Hv8nZfcYgE5otcCGL4cwcLlM6PWyA8OGCj2dqd+87SGr
StrR0iGbD67rM5cYuJfAtacA6Wak4qavS8VlZL76w//MsJqNUVxkddMK/UGRl1Qppt4NCHCfUYGW
X4JGlPlvyySd82utjz2CkGTnBaJEoTCXEykBfaeTCI0kpR293VZ38ewcR0vCaHEOKHTIsKa6D8I+
CEAMZlnTMPKXca80m+MClqc+k/Mc2+hSeQ58Z3c2bOJGRuv6+KwEU+wVB2q0wXbB1flOUazIHjBl
D5hdct3AURDp2NYzNOFrJPSglAg1FV6EOWXIePjUoLENFvAD6yhy96gK2SwTP9SxInytPtYqKycj
zJYiyRXl7inyiQ2W/C71QhUJ4gCnfOCXFk7pwplCFRhl/WfRPkNAQvRZfZPq4n+bjPlxvfkXoU4T
TJHeGPLeMyVcH1ZzvrcMBW/d9I0ecsfaYsfFt9N+s9VzacIehvroy7grDgDojcqHbajqUEpuAYv3
jRVBhDZbDJYzVRropHqLJnhr945XXk7/JRU/VnsYDNzYNkNT6gXtVKj7b5Cg7zkmNN9LkBqJMye6
5RMPuap8JCTzoTKK3tEUNXGHeVa2GSJfc4LQP0ntS8WD6TIlApasREaEElf9P7q+vVBTq83wMb2d
fBgpA+8vdosgF+tQofc+tPjYWhaDQrfHm6seGwKZaxczUyXuY8TLMgC31HfEZ/UCGFTpd8yq+04N
OPxiHUSQWafbvYnpouwHu42/tcXedR4bLECQMWsZcei6VK1/i1DT/TrsrpJ9x/iKG86znbQJsKav
h0Gj/HS69g7jBoj+7FMKLp14+sJffJHZrUsXrrWQyBpMqAXToAd7sALKiR8TFsRr0JYwcn3yqVx9
0QgzvE5EZx27pbvq5Z354mNTy/n569Q73+djS2lHRzKIsCKYKIcacyl8l+erJkcXArC3CJUVLAuJ
CrmwpTAreuj9BHzpCy+XJmb+3SFK7mfKgrdYsmT0gU3pA2fk79UoGXjLOfVE9KIChvBXcEPn0mCP
D15Ua04At5W1r+jtC5M7dfeHJGosql/xDibB825QOIqtMzEjwQDSFCSQP3gTfezHmEEmhzmIsP/3
Q8rWy4eyBucbLfRzgRDj2rIl99f7cLUn6fdCavfhzLTnqnlQJmWda4nUoGKHFXNYnp3r9sLqPKWH
dofOSpR1ldsYH9xsvH7l32EbwBKMbDjJb1wc0NmmXc8L3C7OnEcRiX3ibmNmGi0hEoa27wZyPr59
3C2VD9nGT9jyONNqDdUCly7Ee3yFZRduFGMfFaRYccG4mfhuBfCJZm9ZjxZmcMw+9DYc7HHC5rLQ
At3QypKdRiKXywy4WDjxwxwRJBtKD/IO3P9DTxHlOHRHhLb9Wa1gowwuOm7g9G9dX0WxqEqOPo6U
ND6wuDwKl8HdJBmKWtHc8Wz571kxe94RyxHwAGzsBawL1u9P3tPyZ+BMqfxQvi4+dKve4wfhPOec
X6PrjC+YG71BHlAm6I5m+9SmU73JEiwtFLj5E/8dSshfDqhrZKI/H9LcNqr24tXIsh8CX5kSpFhC
w9LJGd27ynYjcDD38MKTDYOHP19PFzjvMgXqrJ1UiWosykSf6OiVW2rriXHgRakkgvIWhbmk2HGn
+DtdR3neYbUG/2P5gJmYO3dl/tpoJhHeABNSwL7USDQRAJygLSJYF4/csSMJDU9kQ4vwLYuBMAxy
HRKHH0Mb1q0RJXN8UZi5nrNpfSjNOI2mx2/q53V0IUsTWoFTwLbeNz1m8/Uw86XX0IwycVKT6kPB
t/LyajMMrjrn5LmuGUcrxaqMkpaaQGYq6srrjLyiTjqDvs8fF2l9sTq9gEVLLZ99mQaQrlGM6+bN
UNx7fqHAi5tM4Fhd3TqTqEL4cT+uLwhYDBEs/mLNzxk35C1orDnkrvMgV9yNTa9J+yNbs/2FUg8H
/P/grpsg1B+6AHuami+Mocjk+XO8f4T7JJMNkBeIz/laRwyE2zTE5KvjViLTVgOgXUcp9uuRh8wm
PVKsayTLeXS9N1VWTcF+0GlQ4fBhljJqIr8LUfVfzKSekyZfIhGyyRxpYjnHqwlxKRH8WQSNQ3nM
KSkAQSh3C2yzbTqz+BmUgRl0MuxqlCuSBjpTt5Mdzn04xWMxnK/J8Or6WxjFTwzovN+Do4qw0amC
jv+yalY3dRrccFRReMnvL1MJs68rRV7GsVMNTDPd2Me0wU12phz8nJ8zFE6FFlB00XOCZM6YgSxW
04xnUdWNd0i5qOxdYB1jWy/0QeVlrf2H+q83v9vpvnfE9gsoID+vJK4IJt1/q4JXXW4ukQj8eVv5
F3PzR4yeJyJ4T3drqtRhWzW0iK8ZOz6/2DPE0EPELCVnP/ZEFYk1LuzkFjG9AoD9NrmVtezC4/R2
LQnyY70wJz6Q+0BUyPlYYJ4D38JcmAMyKKlD+ZXt8Mbc7lH7WhYSvZ085rZ1p7smNb0h6lF8or5f
JxmMC+YG16OvhT8cT9QM+PsFdmZPDHjyVlYGGHIImn8TL1d491SKThfPEDyDBrUbnNYQYKEh67bi
gn1RRsjP2bI9sTnRdBrEmm4psdYYWyOfP8TDBNt3rfjeVXPkYV13ZhrsYweRE1BUl69rOoq4Nhzw
gau4H9mR3wEYdHB6iFaxir2YI1UYCAx0mC3p7YqKYRmqEyeYiG3QaQvibeowkr6RHsccUBKGlByC
1kNGtev8kqmz7T//1jz508/G7Jk1tckXbWJeESkfR2R7V+TV5+IlDIGn0Sy/7NNVto74lMwb1RFa
e9WkMT4Mww/5gMTLNiyhU7wQguI5+eB8IUTf/ZB9d1YxIeUkbbBpKUDXb0qWvhgCUv3r+pwsUNJV
n1CMu+DpPlDSE/q29Hx6xQyKpr7nK86GK4R/Hm9gO/fMDySMOlSHHdW/1/IGgFc8JrXksIWb9SkN
ETrlJq0/dt+hEb3j7SuR4DJoi0c7kRSCblE4i7LhRYT75NM9ILs/h59bCV4ZYZSVxsmtu2Sb2BOR
mVkaaadTERqcqw/w+jz5i+Wr1neaxIBYfnyCckQHcebLOI3ZADX8LiK1xbMvNnqCwddTPDt7VOBM
+isIu14LSPTyZW+ih0SAtt6bewUF4xQDlzlOhCLeNgkJvLleq77nxPHln3MYA+ovtfyY+xvPe44z
uno1QLK2wyaVyklFh29IRCIFM3acKsQxnbEiIiDLgY/cG1dWzykMto3VjaZkqFov0jxjySXBMSAR
mk7twL1JPqwacI4sUrRHyyumGyJpc/cM9PZVygJIol1G65oaPpeLxVWU7nlFd0l8ELlEBAECD9Uk
/eoCJAbdiIjphOG1YFWWbuQerPkN8h8AHNoXj5AXZWcgJWvkpknsCnMkfm8JeruqMablRO9NR6gN
nHx539wpMKp3eVTiPOe+bf5Q+dQHTPKQ4fcho2CNdgPqxIs3fShXeS4x5ZyuKLYU0I/GL4LwTHE/
nxUNi0wFI5BLA6lgibHWDyTaoTYIcZGFZZg5mn58M6ibIfk9P8KeQ/YBdbBlsgdjV4C/QyQxhAK3
lAyacpiqA+fo3Wow3usBGatQgEDZajCdLwWsaBtQ/1hRYNIUPxGVMBpT9WU8mJ4eE68p7h2umuQa
oZWlf8m1RBFj0smYesBz8SpWWH77V65P3m2Bzx8A65WeFNJvUDMEAxHrbGY3hZRfKl2T6hQwz8of
lBLGavEKghPvCGKwpQ2s4DkVjGGHE4rnqDUhHByCHWzA6evlid+xAaNd/2zH76+O+MjyB7E1p92A
oOJ/yLNzt3LyY9BhJkBSLKQlQN8SDiWzQ5p3Rm/jtp79Fc2whUUmq+EepETjhUA2aONoRr+jluUr
zVgrBCGtXzwiYQCWi7f5nbPkHLSshrAEu39R9lRzWf1G+w7NNw9+ObAofUfqgJe/H/FMtMs4LYvt
2jQ+jW7yQNHIVfKDWEapH72AqAqbJRDbRso+Kfi+IAsYSeKGQM2FW5zFvGoQ38aTvCyCLVwC3UfM
0vnJBihwNew0mu/GDSANogQ4Qw/i+rqaEupx8Kp1uIpcxyUcF45fsE85aQDWVgLQrW4lRlbIN15N
2EqVswT92vRYtvq27I3qNXry3sRtAA9mmXy7WLkHSh1Ui9NLgZraCKnBZTWOokUaLlhqMizvfJmJ
yUwkKFHGUcT1OcjjdYJfciwTv8omMNMjzSQ1Nj2bJ1Tcmmokw8jGH51tX+XwCJEEpDMH8nkeWFEX
ZuaN2rzMA4UEbfZfxn+RWR5vwBpzkFccEnagUG5wS20kQ0+Mxy44uHBY5szor6DwuYeV3aVJVGV9
Kr/jHVmUOcU6J4cOOk6b2a4DaGI3netOBLccRwRhnlqFN7bNCjXVGaXwyY0ruePckLKHN7dSL2J4
aQl7xiD1aQAfAwBB67LZTpvtjX+oDOWAcXviAQ1Wv25StKxsqw28V9+mjmvd0oGOT6Ye+dLCiiub
egmy5ZyEuA9Aoamp/7MTUXPx3NCO6NPAFFfZvujfXUavPk3SiRLDpVk1yqiqXCB0S3TvmVmnu6Nz
iiY/NoML1c6lAO8cLCvNad1vrY3p3OIB/ozbRkdpqw/I8bY1J0paMMVyRO7bHGiTlKltkuvae6dE
AXkIZvElSbe1X93Eipa8weEa3lsk84lusJ41G+5V+6JIKkrVlRZjVmt/DxTggeMRHcbsX+EVElv1
/sp3wgDbCDM2e7aegSiFRKoQpBmh2AkZ8Z3Iyml0YpvS9JpuZ82NrNpz4+P6eUDJwkY6RQrfPPN6
MCGk7KSC2nfJdLTIcZ+6nvrEigtKgSwiltHN88g6/pm2MnQ1FFFOizVqUsfbH4JeU4yJmotYdY9k
zWhsIDg8/jhxwoeMs4Vdmu4M019oeZ6fruoflqU52Ysoqg4sNN0BTuRB0OJ5EWABmnWjkCUSdfAf
4y5zmAlartKseu4KDhgAhispSscq1xE7N+ZIuXM0U9325MMVagUhSDkqOnaEmWrQ6+1fM+6FQ6zU
SGOz7gDAQjKJgj1h+TZPpwCSuJ9PgcOoKlADSW7LSNAtPt8cKk+tfLUVFgjoefNj1cQNu2IRhPfT
4oreIGodqnZeti1Cf9kw4ktDWRT3PszlB1aNZJLEdSFLpK2YRHNoCfkY+Me4zXsIMtTtsp+AgbLV
G9wcZZoF5oOy+F6afWCZ/oOOSuIvmDNOdnUS9N3Jvs2dJ5BrqMA+fiX9uYXNp+PdqR+YaSE6egQu
SBHDZiLqcuRX5frsrbsaK62cNPuiQ8kQHpQZjNchp6UYZWsQOFu8hUNIWw12FaPiodCQQ++F9TNL
HH3FlHOkjVBcULtsG5r8rg5dO9IGoieui+P3Q4yhQWLX+tEE+q1uxbBQdo3caQr3xdYqgLuCOgrp
NXEwcvAxjYGXvHCjcpjz4ucptZBYpfNnHF1VwybRaRPEBOuB4oSqN8dDOeyNPPOi5RHwT5Jb0+sm
8Lyyz/oyPi9kq8CuokbIQWQ0KIXRd6LeGgUrI6ULDuCq2Wkr8SDJwf2wYmkTN0laOXgyBAU5c3xx
t57BZDHf7jgIbhZFFs98xi/QF/7SlQY9rgL44yKurBGCSNjE6kXcM9BSZ+ryaDJJTttg/Mb2/cn+
/gaFl79eVEo+GFz3Tqym+s30u9KhhZ7fCZl1fO584DV8b+A5Uw6iGK8S8ldWaNM9s6798+4G8Vac
1hioqip25hGMog7GrV7TjK0sQgHJw4RRZHaSxiIAddcdXiyg6aP7ntmWscxlyDAxq01AU4bezIVN
M34AAECOG8ZJpA2A7vP3YIdaz9mOYPiF1gxFtRs4fkqIQAZXdMc2IPjdoSQL8I4r4sSXIhV77bj+
vqr1GZ3rM3zKntrUYawQHXEfZOLwmxIQ/regA+u+DtmKlXRxoMxPI3LnZzKf2I7+DMMvdIPnk4+T
VT75Yo+mMAZZRcC2dTc0+qzhpUt01cVNpdn287bswpuaHx3XcECmuqjbXuBl6n5ncPg7Xj4hRx9l
6C71ov4fr8MzM1SX9VA7knH+M6dXb1a6eKYjhF6fm4i+32xjAW+XLmE1jIXZBWLk0d+ia00lnaPh
wQzZupCzUiSa5VVQqg/DcELV9FvfPxcv9+ty26KXZ8UPhWS0ICam2m0v1MhsYlJeYF/TwLcGnhUV
6EoE+ExzGw9Mh/M74cL6+g3h/+l+x27YqFJEw6M1fIyb/W/3lbJLbiSGz7Ge39KA5jXtMaGdTZvT
Q6F90M5osHHanKS/q5+92W7MQNLZxfU2CMmV7l3FQrJo+lRjgdpKyT3liifD9n2AMe00SZlTMxw8
k63cHtPR7VsAJyQH/4xHiWoJ/f3153F7fuvSjgj0m2738XGL41GaDbn+JDXfs3gmIGabHJgd15jP
Wn0yTUHkl/CQNL9insDjMuNJAbScvjimWkP14r44Gzah79vxZ09qPE4MjE9eGXHD2nV4n+KoUoRg
y4QYsvE6114VPYl0dDSZkHHQNd2DS2aGVSuxCRZ2rP6MQWBcW9TS+EF+k/YLw6RMeMMpZfxqC0x3
JP0LorfC0Cp3JcKhwdXM7orcS6dIahSmafZYV13yXk7P5vrkwv2gXGZ6IAz8ZVAq8RkamWJGVHyS
87XNqwIivhJdjnGKuNh5mUzJwuLpkNRFb9mg1zC2RBXeNHMaW4zcx5KPxcpZRTVs36OWDxFdcBKG
9TqChQykAmXRYAm2pY4mo9TuPpb/Axda6snMk5JNNOwx1X9dE+QzQuL/JWRq5HeOt3KPSRimhVV1
wleGBPV8fR7/tdjk57IUwkDJSIUvvrNOmfgwQREKVcFESqEGgb5uNE/srhVObK2Yhig2GYBc59/Q
LpiIT8N3ik31IJxRkwHvaVhvNKN0bkG/te/i8rHOa91PJkHtYkY/PDxIbXBlj1Wo7y8V6CPeJOeV
lNTvtlfGTH2S2PslN0fviZNxPfHNTBayKw2ctwOmWSxqTMkXhQNthE1FozeeAmWOPnHD1UYqErTb
efEbeKV6z43fkjF+PQo2V0cMnKhc6RiDrW3yxQZWSBNpbPG4ObNI7njRgYeEE2+xLmTwq5DQ2/lO
WafzPnulESP6vaRL2mWRipVxVMrbMIYxp+Ygt+9UkJ+w/EC6ssfs1AQx4lyvwVkaqLf/w75EsRO+
2B33yeU8s5e1T17qrAusC23sVCjBkVbl3MfdYi8oGzFDstTm8vCl/VpzKQVlivPazBfUshEFUq+q
/fQZCMpTvU4wqzUTCrHp5TB0LWjewRQJaZMu+7T1+pWGtkFBU0p7n6oRCNRHKgrSW0HF7qVRq1MA
0WR3RhQVnh+cZIGjJeiltwltY+ZeuCbgsmokpXU2GNuPEM+/W7Q2RbKbG/NNx29cvpIIvv6XpaeT
jsz1nzdA1mMVLv+afRQgekDolZSbFqo30qKnwj5zwKma9HaCVHV2tByOUklscEhCB0iDdwW9DXUk
PvQOSA9fvpeRHJ+PyHSVO5HXgyu3MS1je1+BHT3vbWRuvYZ7lVdwvOree+ycKKEP33yi272KDwy9
8anjRCmcgpUDNdFwjv1VEkwdHdLzrANDEq9DbzZP72f8DTfKO/3Gjt0uMUtkSRwAlVVCvv2WSz2s
VmPTzcttsRTVJXG5g1tbAIaswgK+88oXoIGxzQ+u8OVvC+xkUhf+EKk1HQh5C7cm0nY2xhtW40uk
vEru+ruq/ytYIY7TnXpoX51fbZcnQuTiV8PhTZtp9dHX/JfDo9lKU83iKuom79tRszWZbspzpknP
rqkEENhTuUxE66x79VdaKGEC+nVnl+tMp0/z7GvSAqexmqQusvbIttKBX5xnVdT1PR7wPKfOenSe
DmE993PDFYYe73gtcNcVtuC9SxB9nk9QFthFIAbQdkryvw8V3p84gPSM5/OrMeY4cnaHdsdUpSDk
qg1375F+K3bUbVbOlnLGpnTeKWNdX262ucejq3/MSJZeu5pOU/ZOl6OTyhwYG6lH1uK3MJQdXQt/
q35INzqHqyZXrkxrMbV5Cixzobw9KIqtar73q4b3ilYASNSoYEd0uHon0MggDpskEFHYwePJk3sM
szk3DT1hjRIUlMByCMnwB3u29IPyTUJjKkEUZybmDmFLX5km/7jsWtxhIj9u6ZIhc7i9l/phZDha
m0ijk58ShbgRQ51AnSjskAGCfitII2gu35epn9Ger+myHxAONMB7wZN0V5eI89gfsPGdNQfZPwLA
X4Tpgcy92SsDzr7pxMAWm+uoR+g0j881BEL/pT+ff+FryymufwBoidaA5Bckghog8FqAIoIiocS6
c34Nq9kISGs93i3d3GrUcyOKbNu3LzQQcShBrBO+P5Qwi5a88Mrlj30DtG7D23YFVIoZLQNciAE3
CDiJMqNf9J6wcNOVUeTxe58lUiTAyOmurj4/z2ljyrZke/KsTALVJpDRVVvVL4Ebsniy+JqqU0zD
Ob8fezeSCj4LoybdvgX2T0hiQLU8Y2tN2xICR0ZLwUXJMfWXyLVCf1vquNh8NChVb2/7nnzlRfRv
eOUVnCpjRoxbHNaAwkW7RlvLC36ZcVLJTTnYnRlbp4XDEZUn4DmXB3k75W2f2wLJROPap1iyP6AI
SG39LNZJ5hdYFBZW9V+YOfBJfvfEKrJZN977Q0CLCs+PpTXSPjI8LXvthXqA0CmtEH9k3nqEn2xj
zXNgPcCUvn/sp0aWWIugfloIvufjsuIvdAQxNOWPn2Wx3m/rdk4tsJyEJN/G51v+135EZ6ZI4kSw
zZcjPIgnL5mGog112UTv0Ckq8MITowUnhtHhJ4FvSyNKRMbPVXNeIRA+WvsNgsGr5NfG9ExSONW9
WaX7Ib3943wGawNtgAKL5Y/uwfZSFuCEIdgx5YjtGRFKaaiCtL1f+8jBIOu61VOm2YEwaHIAZ1ij
09o0KBrDSnVPttjTa0VzUepkVqj3iKFSdOy3UM2gcy83Y6B0q0kJTnR+FGdRAYfo+3WyVCA3ByRO
PiVS8emu132SVwy/LPNzXDVKQ3zvtE259tfl4j25K/6Y7ClYs0c8sElf23MgprVg8tll5KpCD8Rq
KL708n6YGEoDU2D7u4bVaufKrFL97QLCuP0g2nA/JB60Pj+UNOuNskB0neCZLkGHiBrEFYf5BhbQ
vinNL4LoOgFRy711C1T7/4DDD7yXYowsfgmDgA76IAWsXqTjD0CVJHXjpuHUVvp63hSxWmABsceW
Onge7XFMzru1WvDZ+5dGHmdBxPz77wf92c37TvuR+SKxw8CtVlz1DBRNgugMDlCuY5Z6fls/6mID
KsLq/RRP6ffHoq+kRh1H3/6ieuscXuAkL9cVb2e/rrCgVoN/XasQpL/FtIj1GljavRHbAxQX+6I5
+LG4cgpoREzFDblJi/W0qyTNqCWoQE8W8NDarDPFQrXU2sgoom0pDo4LreMtHIQEHj2fIBS7ER0I
ODD9b0vwEYbReh+KadfjFvOCB3fNF7SwZDZy3E61bP8zyDa37ZlfzF7fqwNiysBNZWmIRayy48XB
G67xWBMuFvvDGBgj3QyktDS5HIbWKSC4xxiGZFwJL2M7DGbjo0gUkwCRcbU4lGfr2dI3054L4aNZ
KMTc4vI12OflhL6wcKerqxuCwKksIR3zJD7Znwn9PtftekvowozOiCQNd08WHBHKqqIZEdkRBjKp
yDIOIunCxOY7AcneT7tlYsgCeNG2c/vAwE7IkeVmAh5uSUtaHL0+oboDwosauA6/ftvJr8xbxrFN
u5e9dYb6mv7Ct4SzHW0WPJ/bMZQ2MV4w8mx27TeOPUe3mGauyW3JFLMf5qZHtN1Dahcon3t/W/r5
nK5XSshw0duy5bwej0AggW8HzUaCqwedx6AH6SUUVNh97fRxY7SwaNYjY54DzdHKuMzNrHctr+Kv
N7UlLodlg0zEJzAh/l6ocnSM9w3/kZAqB2hcD2SL2PzrKXpc2CsDZhTWvKKn8dsIT7w05T0cz4KW
czwrdebzYnVECiICaREvCh8H7EU9VRJh4j8XC+z6zkbpdJ8btJAoWS2Us5vy+g6t6H91AxjUdNDF
CR9xcg4uIHE+1cj7hoB+ENlqKZJdlNFnbfxslXqqhhoS1w37wTLJsD1rM7enMXwlabFwTr/vq4me
Z4uWdrpUZAc+1VP9mD+L9fdPXKRz2L2vfVhLLoS7M4wG8nYsDxwxVaHo9Wbs4vszk0VHZp/nQPLL
TmWmSgXTNiupZ8ZU85oM18IgxY8LiwFFBqlcA7kavhDwwLWwG0Bv6Ya8lUIiFlGw4p1efszZgevU
sYh4yak+2hVz6j0hmulqFmBgAm9Uz4Um+X0TnTobOEHxWMFME7zX+BmlYyfqVXnLE8FAXnOzxB/f
Mi2gW1ZGNEgJVZ7rPTOHWoeTwPa805xCHEnZ9K0ZORRDEZDmhKW5aLQNixKCKl2usN4VCtbexzPh
HIfl9vifkPkql3vWBSH/eT91mUDsbuubjQqDw6xjLbKLt0qzA5rmPO0MrjFUg5kepvkix+f+I/pS
tp3G9jJUigPTr650tdkM/loNt8rpUIfBIg9m6G4bjBdPd3iY2GeUtCBMhdTPN/4pkkkWXKBS2OdY
fjW6FBnhH3158fZ7cgzNkZAJU5GmhcW15AcFAbjOLCqs0qKlDFjMmG4pEeP1wGRfmNlK+OoHEeHS
AGwfEXaAk/fdBDybEfEpqPVoD67fRItCtiylYYB3lsOT7qha1ry3QYcHWxqs2k3cHCM5oW3QUaKy
9Drpf2sOHrnrA7Bmg1arEkXaXQCEHVlJHfEBR+rQ98NEzF0O1RqyDotGwrk485NcBbcMuDzTU4/o
d2kBbfQmg1R9F1WRIY6NxpzX6LcjWqG6SAjfB3CFq+Uiuhm4ZIzpx5FBJ5M1faZA4xXxGR6I/gbL
nx/lsrrrrP8QltiNIkx15RXdO06KAn6Kct2StdWnKgNXQJp/eoSZPLA/AEkHzGwHsTyGZYKKyY2W
/LgVOssgB0oLFqJnduZGjj4Dsp3k61DWjBp6ZtqFpBrXIhe6s+r5F3v8CrT9D41M+Z1T47VO9Jwi
wAp4PfCpkbgXNRp/QjL8aHCmKC0RYDLTAiLsoT7YtUnI7k86u1RdZ1r38Nu2ZKvZiyrVMRmwycrS
fKY5onGCskoLcCosAUWbobqGSOuEaNW3HzOvqB1JUjveOA/T/GWuH5KYcKDjriLq2R9z+1lcIpzT
qyTKtfhfQhRc9MqMJeYiiNJ65VmBALgXtE1x74ZJ+LtC0z3OerESips2P+q6CLjAYvcgwsDYY7oh
rJkOnRD8r2O6wKsW6776ZqGfChCvf+SL6usB9yqkpFtp6768qEKt1k4YeNNXpETamykJYoCoMpN2
/gtSGXUsWIB0J0VKqpHV1vgWzSqahHzI8IorV06U8e4a655EgbO8BA9BWcCPwJwFCXp0bYCb2a0f
fqVRnT1JcIl2xAcmO1OUo7rrKuzc9jB6N5QvxG+Bn2E5c6hoYe1z/BgXl629ioo2t+scC6VXdPNf
UdK9mo00obJ1YJr20MeYx278TnazByMfLAi0c7Qr3of4OEKW9JRuYE9NIUa8X/tBjX5DzbJtnCls
KpcwP9JqjqAc2Ln5mzN1PvY14CcBfsnJyO0NiJtIOUbGjdX7CEOiA/mslKa2Ir6TwcrPRnMqsSCT
II+rGGKl4dqeBRc+fLnUboZ7v8fsf9Q5qwYF2BS5pbbZ8MMwjQkCJIz/P2+ZIMmLc+xEVlKhLqBJ
SOzpdH9A5kQQSjKzNSeFS0IfAl3ORPG5SsF2HX/Ac/LanioD3EL5yMRDS+/+NCx4emmvo8oFNVu3
GoNgMScAQULmedo5PYuz6TsN3olqUVoW0x+rjZNIoZxDr1tHqBUUv1bAQj0omKRsVdlYS9UIgEw/
rhqc6T/HAZKl4sma8MxwA49JHqeLUoGUcvvbfNU+M4C1Kuj6xgJp3PSe8WDSfFjNd+FseL7ZY5W2
cEASsxYQsDleVY17gjcFnnNuvQILQbH3a00JORrBZ7qgW7ZoBNXo1GnIsVx+jbdlSI0Swf8D4Wxc
CSXmXOTX0XHgF32V1LN5sajMULrBYgN0CkPtQ9mvW2Asy1naUO7h96Uaj2UCtDGEPuwv96fruPT4
MRnGj/Qi1sCzkLjpA8GdABFqvwXR1l1ru2sslYZ9CgQoZMGrnurqKPh0EsT5KbBaNnC2Uq6p8gQG
vsTP2IGNei7L0ybiy1uOWCZkSJ+KBZPu6oDCH9Rs0aRMf6ugF7cgWS74+0pXGLNDKnKQ5Nr0cprz
RjdNtfV0KOPOODMFG6wO7CPEHSHsSp/bx47ncO6uq3kbtW0sVViTwI8JedIV9vbCWE9VXcpX/XUP
8ygVpgelTeEYue3wlvkPmUQgz3dC4FW+/yPgO2mlych4fEVz4ZVrVwImDimpH99ZkNxGQPsb3wu8
LfU6MERj7WiRhjQeCdL4AxUVi3qhp7z+XLAVFmFTcSGYj5AheagW+We1m5WMU1KBSuILZoo93/wr
p5hsqRyCIKalxJh/6mUa49WyeLHirnZnUzm/6lzDaSeOBIVochIQHQI2d4TTeQfdUIn0oN+wxbHJ
hlXNznADFfMNjesfNbSNjAYVRBm4V8uX3UFYEkIq2MZbNTp8WR4oIzu//xAfoiMYcif7GSL8QX2Y
JNHbijLiG9d39sdDecM2scqCI+YTaA1NAEnAQvX52b0hNEBmIW4481jrmglU3+Y06hGPyLT+0FNX
C+h8dDd7oPr+rAZz376eVsgN3EwDq8X64bNVbYPc8i1YKKeXpAtgVX8U6VkIZPYTRGjLXfs1SwEh
MNKV88k0a82MK+FvlQ0ULs3IiY0urzop/kCCnEbD1yP5QTZ3vHsYBuyStnduQ0G7QR8RmM7thjET
u4TYwuWrsfFJFD7ijMwTzmbw2bg9yCrWF1UxZKOHvxCCJntmaoKbepe5iTfD873YhtM9deVGi0/r
E3HvrjkL1h7H0WH+mfSP/0jA4Tynha2RiIRBJJYVWic6XuQ5J+C0+qHzNq7kF++v9XK95XqBE5mv
/SZFHa5E5w0dvpQmLHolv47v+onq0C4Igb/RHtL/f5ndVN4PusI2pD/0dAnzM97XXYLak0r8i25M
hOIrzuqonfLJJTJHwIHN8Xk56zBoZmb89kI9RPetculecp3T040J9ZiHlbna1OmXb5anAZmj88jt
KO9zJ4GFzx0IxuR6NVTzH62tbGzIV2IGb/zKQ4sQS8Lr/fdruT1GGU6vPFP8IbXaT4ANXlgQl8Rc
kuYn5Yw4P6LcFbLDwzO7lBULHEDY0GjkEQ6l0Xv0+1I41hbCpzcQstAUTin5lJU3sMov3hWPQDlF
xtQ7qcCuXDZk8CZKkG68sGXCuNTiewDzjM0R+X37ubskvxkNIkQCxoc5Lj571Vc+vFJpLPAO+WpU
qoBXx5fDC/XVkk2dmxw6ouoqjWGoycsxJrgInkiorD6od151NiS9pqOephdVCTGTt1v2m0U1eYP/
OQOFfYipGtB2dZYCFAWH7Lqb8pAfl5ZkiNlLuRBOAkpnVc5UaflOgr5vFfRNMyZK8uw9gTNZ9W+s
QoIyFDG13bIHlWgq2fiBGlTCL1vZeWAn21K1Zgt0fxJibs186I6+Jzmki2y+vkRQZiuXIpPHV9Zr
ivVe3noTTeOh35n+LS/ag1r2jRJ0yQ0poe2FD5wlLLTA4boOAfqoJHXX67pBx6JQB6N71psvkBFT
JbiKEOHNY9F+Q6ccEoHOz+XuDGpqPuaaHuda5S9uc3AO9Q13Kp0qPT5y+eGfIj/sriiEsYuQKglc
fm55gwmIrM04UVOBqucIwb/n5OFGzVBlA5v2leMchX4Arm3FSK4HJRPZOeQqAbZopbqyNtCNxs4D
hwdyNgF1nTPeKkeTmrSOhNt2HAp98Tm1BxRaJGOYasfGwR9XNZ235VX4biepbrtW/O9V1plx79ZL
kEKKxGl2qorjiwOA1NSs34eFiRmcEmhn1y2CXTS8DH7jmxKUZTbfcA6uQjU0ERV7FSrU1mYNmMEZ
SxEQ4+IiuVIvOX2tpPPlxEsleqjfsxGWXCeKH9jnGeb5a4JLe692uHzGqlOzCn9YEQ7O+dv8c5Vu
Y7KSFN6gqBVrgFUWDkCXvnettQLoRUAzYg7XtcmbyyeiOf6FDVRmleMlkUNZM5GwwhiHqHiegnoJ
F8TtnylP1ugGbINWtu6/AbCgMkxVym6ArMR7t7NYz0yFqabtkQFv8mSc/2KYKX03JCvrBFc3LMpV
C69ayekW09+2+srhiJXIZTOGkjXxeeaCGe590qktK3UCvchxlLyJs6lOTw6V8F0IlaA8Bk7uYoZ5
iBmEiIUt8AHwlRs6yYWZryw/iLX0p6eKTWub63tzFqoaTFE5rh9LVgOB5JCf790UZ1eZuySiQDHe
OW60C4vnV+fBPdXnozewyoyGrks2u0ec+t/ffwaGs38sLVdgMNTTOxLGgPspT1z1C4OS3jWa+C86
0Ql6wHCL3ilaVuXAHUgzfK0zF6gHx6q1eOfgQy6IwRyPgNmhZBpQn2z+EwwBlt8zc+Q/d53sPFBH
kAXfCH8UCT2g9fvanhaiJHvJuGLUmx6YlmQw0bzoi899lQJeg6gVprzMnRerGMHgZZNysqgUbHA1
TqE3oWV9gtBFnCk9/FHL7yzIF/Kpmn4E7BNvEgO+yM3/Ag+Hh67lrF5AshyG8Lm7cGDEZsamZuin
sK3vOZ8GC64scUrha6POjdo4gdqRVJ0YYl1P5M2JfWXtW4GdchqYKZFBwoxV0OtrrTk7r38fFxMD
ypk87d0iotBMsWZ2VAnpw9OjTCTTvUAS3KsSkKMZY//I5D2A4OBlO+IP/POqjw5yhDPt7jbi2Zsj
oCWlUINMQeu7JpwfaZDJdV99ETHeUJO3ua+uMG+HeY31WYYgdHuHk8Yv76/gJmux5QsNbc8JxwLY
LbQxjypCZrZzSqWwx91KMk4QGCcE5t4iJyazioLvNZ8xpjIReZdkHxepGhIK9THtqpkz9f5bNSkf
lgx4UmzGbdy0AAEzzQoF5GhpBdGk5i2y3CSE/Yok+OcXeBrggtE/tPvT1Ap5QdIwFpTSq484bcEy
i5DqO8eczFqxuJBPwyTNq02ldI/cndhV+xEgNWB+6Oaj+B2lgkEABFL+SVjA35Z6XPPi+yBRg8MC
7yrUwjU8TJpbG62ah6N0sz9389vBQ6ZAGkjvsEhN8tsxJTRte3tx5oZATaO2ARsmRm+c0V0v2hOd
eydC7ckDQciquNWKPaX7Q/O4IY5KivKao5DpaACzt9Xv6X5jRaJuqFcSfvmq3ryaXJD+KLIVI7dz
mWveLb5KV65LaTXtO+hCACj3EnhKnFP8LN45De6QToaqqWM4D1SHUfGCrQPugxaO6ZyYj+lwN7Ck
j8hpL/3KvLsuK/ILB3Liqngq97VfXl6iJjdeV0ZHZUQR1OiIL2OFO8v4K98Zqg71z5hU/zdSfHtz
N7Ya0IvLylmFt75TdtFI49V5Aua6OLNus6MH31mdr+T+QOP38aWQrux4rwKd/30ZqFfiNTvePB+S
b4PG+G+7U5OgHl+3vGOq+9CXYuAJojTxQ5mD+mA66VMxAkW9OjdGjD4XUgE9fCZyr3cL6B0TDdbL
81Zm/3ES2Fb9dx+c2N8LOjN7qa7vMClIEiKiZwPeagpmV0XHulsTdjSsSCs3b8ZZw76My9vk2b/C
EaGBFTHl2XTyUteYPj0p+zVd2nc9IKE6/pME+dB7A7l94e7ClzwRlmkmJdF9PFRRmGgXKW59kcSK
uVPBb29+7hNeE5XhywGckgdyfZmNG+zUSHgQ5dUN7qQu4eMHCbHCrndxvc8mkJWvPwSiLkEptQoS
o0Voh4U+vl2ARa3Eh6SNBjccFPGB0QqEkallMlWTRzIxWiGMpaCTf/xXR0L54znFQQaSZHktCEZI
uRvyXxQ3qUZRbsNCPLHkuQ1QCB6jmm3o7HF7Erm6OKiZ4RygVaH6ZQrf5GMH7px9leQcnzqhYkPO
IGjOU+vES+sURXhslkN0Vn6YGWxnkgmWK/hNRrxEJTV31Ul7DqH8kPr8ZB6z/Hq140eXhq8Yl6q4
jb6vWuSsKTjtBhPxArpPQXZMM1Cclr/9DUajQklQG6DeL3CmBDzOgc+7sj5ZnLWztbZtWYDf531O
yoX4SGzDYURvb45PEgTYUFOpKwGOm9h7HxHCdALxe4a1HNKwMZ38ScvAJxoDu9xPMGZM9JaHuq3Z
BfUM2Yw2mUeE3TlXepEzYZgAZy2F7GS5yobvZgTXVU8m+8+elG7j62VG/W+QGVEG3z+nl7YAnFCt
zLnjqUmLdnBWq736gpmScV2I9xhofu1Fqytn/oijoBCGLezwMosKWgI5aUfnMzkz1NWrGAUnzLvG
ak8bc3YVb+r/aL0JbqrUlRihkgjH0DeuWT4i9Sv60DHC1KUpJUavvR5QI0ULS+2C5D4exa5aIELy
Pe+9b1qzLL+TI2OSLCwMrPP1T1r9CeNKHqkzFqrms4PVD95oUiP0QhE4uVd0wwuODFm9QN8Bpkq7
G5Z7DAN9ib0HwP8UhXagQUDYM1qo4fh34+1RJKydXmJ4dJAMQ4oQLi1WujGMXrabMP5TgOXjLqkG
FtZRANSIt2kVSzYK88Bq57bZISiTrO2y57gTpZN1rn0Ys2V4s1X07unafkcrGeCBeQ2dw/0qwJBh
qr4BxJ+mrq/yvlJBTenDrlueovsUWI/xxeIHATgXZp1pbGbViQSDLe0Dofvlu7OCb6dQriqSEAc1
g7BTQuEfKSfrqLWsS3WGDl5onKnZ/GNDS+Jv1mHWsLtnXsdujEiRGrxzmfmOdBKg39TP5SRp5KUp
f95LZUMXU0DdNeAtf6kImbjVuncCjYLLe/3Xu+I6HPGmAM8SRbn5+WIJGcnVSsttUsHDcXwHEnqU
yJSTLYIiYfqaYU+bClckuggnShY7/yb3lDvQmiyZtrZOfJvyuprWV5g2pI671mRyJOUMOj8GMLCN
h3yvvXLGiC3dUP9qyy/QE+C0a5cLipcYYtcCBFVF4zP3GCc1HZRKPXDvPoMkA3loPojkAcF4OvAA
RuzktQsHN7Lm5WnWOPkBNvxfz7NfOWGXtKScqGKf3cGkc1n9JLHPaqddRCyGzAo5n+pW+GUtNGYB
pmQKzb746VAjdDWQcPhahflfBCuinZUDrZEiYsNB0O7aey7Mv4BMKK1Ozu8EgtRj+rRNuWS73CrF
0gz9y9eNDVBw76+vq2WOXSyntT/ASxzDYDO7AO9f355Ajt8daEIgmg5CKL7iBqAQcWV1T1LRZULs
xDDdxOBkuvFoOvE6g8fOLk8d+seZSJpEs/H4WztbEIEtxEsLaqbqEPHl0BSVO2blLstJOVFu5w50
JC+A2ejIE+uoqjHCYRDD3V4dGoDOKkWxPCMVeuk6gNlILZljsI+QE14V7TNWm6U+UBHvD3j2GNax
XmHp0gQpJz/jvh7PwsuUQvDrAgaonkpy6hL6T5R/D/EyLaxPdjKJrsHTKeT0x9z8x/vr1jW5l3k5
JRPKjbMLIy8eYENFhI0jAzVrZMu86At5YTma8NIZ8U+xzu4R5VNrm+btee7GnIqHJX5KNuLpnWKT
mePe2An4hf4THByPPGGcwFHZ4+2vkxhMEuyPVdluot2zFF9q2S0w12QIAfGPbslImlvsLQvI3D3b
dCxgz9qYmDVBF3MUGKAFvAyzYzb5S7YNyO3yut3zUUYgyiDLhTH5elxzXcnjL7tbWWGaW6swRWYu
uK/vbE8jM5dtaJBRBqbQT9BuGl+qVfFUbwbcuJcQyLqpibVb4aqCsTGfHSSSnk/rBfsI1Ln3qae2
+Zcx+Jg3g6YlyylRUntmNcYHk2bJPVC9yOijtBOIT96ezIaRZezawvScpQiAp/NCeImVM2jzCu9r
gL48/co5MoREYvkg92c/i3Y5D9yTWn7V2iZdYjOSmHtw49yAKrk3y5aZVfhEtwu+ug3EM2Nfjqhx
WuFJy04Nb9ZJ7/s/Cw9ODs2ASEkUoIR8+fcva/4t94QGSoluKxR0xEZEhqfMz0JYNbn/SDVW9Wi+
OlafQretbaBeWbXSU57YpRq0u53xT1er2ApcWu8mCAWTHXYWoL9nUUbNdOwA7cRIo/e6Hcjy43TM
ZvPZ8HEzX4Vxe3IqCqtTYQlAlUmgk6bWzhoo614YidM3IX/quPnw1WcqdwNO4EX2RqpXDihHGDDU
IpOhQ+4xb3tCPeOozM8EWOL66y3nGIx4auMZlKHvMyBiP52yHbp7Sqxf1/KpQjGYifIe8WQ/lGTd
HsOs4XNoBhI4wmsa/cHDzAZAvQaAGDJUN/RKR4nx7JleiY37HGC0hasGICq0upm+TJjSe77T4B9l
U0BlK4t3133BaFjZgsVwCIWanJKHXfA8phgnq8B7CLiYJ1dzcRF0/LfQSjrth2ibw1o+EmGaWDX+
FmMW8Uw6MSxYPghBkRUMv+g9rSaFIyH8IZXu8AyN/4Bct8Q2ipBKiEuhzHvGMNhSMwjBUnKVIVT0
wjlbZVjbxbJDqrU3FbSFiACyg4BzEqC/krSXHDcq79VTXZWvLk8D/1NiLS5sljMx9SYn/DyM58j6
auTogQD/ahRgPVuHQxbuzqFtgD4XjbiFvVqLKS8FGfKm8rCnh+G/MV4jrbh/935ca9CGTuacDxdE
nai2aHm3sviIS3DCmnnlxYFzAsSWEMbm/hip4Y8cvTUmScuzNtN9bO36hl7nm7EIFFfDa651eaZK
NmLM6zRbQmYDNadcgthzT4RfKueHfIA6npk32DNF5oTFHdlpj0nwvpVWhGAJs6EZ7sYxxtgap1kn
1HB7q6ORTRnrSzM5mMMcQPMu6OIY/mYIiZ1QkbQdSwiE1rz+0WMu81CcXWbWDXk3+pUMizwaojUy
qFBMRQvzPmdFopKBOP4GGxc9CNVqavxe88E27GrU+bL4hf6MtezmRfPPcDXSrzrCDzAra4X+BgD/
uL/vsf5UGfX3qu7QrZ9bMX0mPRWRPIyKznZPvjKvBp8HOnOZdDPsd7Al1AiwadqV9GJ/3OW6JA1A
Ecc9RP1lxXer1Yt23z4ETyb1Dvii3Ck/cU/wtH2H60iveEAeK+HsMzNKYeizGLf7sMUvL5GsijS5
45djTgU27TDpuN9Nx3DCTgIER5CI0J2C08d3fCLAKkj/nhbLNh7bp5ovh6DDcmBBdvAWfUs+gwdm
lA80/XGK1bf7BGEFWXtBBRMcgiHlm/EcOI35f2r19bDdRs9lRvMMTw0xmFJQuvLF9vA6hsCRYGtG
dzXTfM9fnvxwp/EB1HUCYfWeERj1gf+M3qF+i8fRsXq9HaYoXvzN8e2wu4T5PBQBgGQ1Q+b090S6
dgnlHNS+MIG9a/oryKSE2+rH8xg3Y2Pm2j6WpZ6cxyRjOkDqTIG+TvydvKoMCY6DttskYB9/XECO
HBrPH8gubro+O1Rj9IYgUeySfe9aOY2qF8cE7a6qpnWMuHa5YgN65DED+97w6fJ/6e+t6cKNWamc
8NEPtJQ7Xhs/5ExQMG3Py/x4Nnqv365iE9YC8HCvz9DApEruxfXlVeEtNF8L+HXWYAQTWIhu6Ae3
mg72u24tCJVrVWrB29OlHvPd9rJ7XBWqPDuPRGYhDHFDNghWvZuH4ieHUUe6e0lP8HVsOaUy0+XW
wr+Bq1Pt958xBUtn7aP1ikSeHsksHHQbaI6Io8sKShgRRncy04HlKk36zMBNbA0CTzhJRj7wrkWS
rmOuCEZtJRHjfXZ0wMn3S6W1gCRHd20v/dcr0cFlmfntBAmkx6ghse85HiaT7Zi+S2DijaipVCII
WBwyurPjPjllVSVjf227DerBpmuXIIE58fYFfbLGNawCV5RlGox1sm7S3r/tAnyZCW5Sa+knG9Ny
idaPp9mSLcmDPl89rVsSJMBxL1Kydx2W1lPruuLJDedrqu21sFTsjYiJSbK1s6ElWJi16Qcn0MT/
QVPEQduee/WefxdEZwRf+Kj5XapKpiNDyPAvNd7g9XKSNQH9NAHTGf1ekrTMEq3n9Y1B8MwPR5rB
XRSMaLf0YX7Ve5yBoVmjzP6YV2MRmiEPQsB4CkcnTd6xLQJeSQcXzIr/nl/dYQG9rplR9Zn4jmlc
aY7BqBV7+hfLJV5C8UxQzPgpW8cX889KX+YyRG3JDievc6GmNqsfPIMWskCyrosR+Kbaqypgt4sI
K4zsD1OGA+qW3Z/XArQOd1/sODXmoXt765MXSJbPzthvWFunPkBwbatGt02epelrZWCtdSWi3r8p
wXZufdEg6i2UD3TkwHFC97JxxGLJPAnfaEUKJp7BM4xCSe5nz94j5vGlzeHOzSSypopz+h5D9epn
X5jQQFEQoIRy0wEX1ODFBAuVOy6xJSmvM3qP1kRKg8cdujgvBvP3yXZi6ufbqdDOXQ09l1FB2Ckm
xyIivtwrgtV/48SCx0R/LYP0y8hAez04c4avzLW39VutVG5dMdnTZ5dH5fzVyQgWSyTqc5GR4Xoz
6SdTr7ZPydqqI8htLePTFLr55AUmRtprZ9EA1Knn1xfTRKyo7EQNWrf1Ffid5P/Aw6plwJ3BF4pX
b+0EwUqhZwBrHIsJQCRYtLxnxLdgFU3LFwEZt568s19BOkv8mS84ok4JMdsbtcTC6VK9mUPZXwof
aHSiCu1v3uUZPjkdgx38U+Ha9ZQCs/h/w/TFBRb5y9kLPZp5rv2HHuN9kxU5xpAqYuBQQnI+5H7v
2OiijZA8ukNFgNI6hXmHf5eaE3e04dP99xPpTVVz9ymG+EZ1QNmf9zX66yIgo5pFAuUhfvwxzn5Y
r6JO/8wm0li4JpiLgdqM/nEJ2eIekEVcFfnnUN97p3R+0YkQ0b3mcOuJ4Jbtv7Jt72WWgKmxDpVt
WDl9rnauLHSLkLE/SvHVwjEIeLH+0tQDfEZY9BTO6/zLILHP5OG+uFFt25M4Hg8pOdDDwJ8EeMHC
zFVhzwMwuNHagfT1HfoSpdPwx6y0LXE6IuTqPtuNI8YtzA11sVzwCuSmH3WBwt6DuPaYi1qRqonD
lH8kTw+3c9PV3qV1+Td8ssNhkyFkaKd0Jb5XfoO1A6ramWGpCnA1nrTDMx5VAXmOy9nR/t3dK+sp
OwvIjlTjPXa6js8KnoVQS0pN4P6KR4SzhkSjbxWEaympZBhyLWhepnhfZ2pqHBZWb25ad+RHr1Aw
uUSNUNh/jPo2fNXYXhFnQSmGeTP3tEtSNxiwkcfTS1ypzaqRoLqjTNPufSqTPf5K+aHRatBeTtzf
iZy5vRpcizC7nKFdkFWDNNQZRt2vY2bzXdegkAG74xflNPHQ9P/iUp/5pdgSvcCyxZulOTFeLlf7
oHxz9MvdxYkjPXbxYdJysrhvcpToufxxqAvvVoWOd6IYQS/RXT1OA37mxsIHoZ0zowyUbohMZmXF
73KTc14P+jA8RTLe0yxZ0iy7xoT9YJkX2b8dQ13CmVvq0AlRqAMVMuRqIg1w+owbTdVzrO9F5339
M+EXcmlEN4ITDOMx0TeZW+La/ku5b5ptYA9Joa5WUf/7cC7AMPdmf0mmVckfDY9alpoAGD20drWh
f6uPwGWUc5c6VIt09ZZe5dTmDZVyEwUDxX08UtaXE14hkeC6RmaBps10MCIdzU7v0kObAiRihljf
3Hx/MCxcVzLyAaT8q5Q3eJZ0Wgq7Fh9+rJL+XQrqbo5tJZuV7jyMGOtUplmeuJMq+SM1h5/XBCV1
YAoIVtit6AZw+YQTlza4qFFY3mRL+3rgWTY4LKQVt4yCpRgDStTb0TSD2tkTBIYp9a4uckPBpvUZ
m9m4KWO97APrTbN8XRmWssGN1AH1vhVjrznYXb/D0JO/DwhsoIyMdV3nueHjFmslpZJirFiGctp7
JDua3yt1OAU5k6O+UrJCH9jdEtOQVyhcVch308lmy5k7DTKh0dqotT0yNRXtF6a298VBCHkd7Yvz
RFpvYuAElFqA47v1PJ8tpoJWlBXzxe1Oi6wViCeJ6VjIFcatebt7fqmTpxx/qjevH4lHSD8aPSUP
QnBcVbzZEB1c9XqHGPpH6zWJpouckPPJUCs+hKNl0YiE4cv8NRvIajI/fV5Yn9VL8xxQLI6ZJf8S
7Q1uNlfs8Y+144EUz6fHkk7z4KH5lG8MxJ3lsFRhq1AcaQxST6V4p1uifK8MW/Y/SQtWWkU4YE7u
lYdFPuyST62Lv5rUyoPOwfrpfyQ6r/9GZUB2RZuozrw5XaNSkxFBj/ExVBiB0492FbX1OpraZaMq
q0+jUaI0GtlN97cLzOs4EBYtszlqcRr4CoXl1pGmOwHSK/TUyLpIFfA+/G52+sWK7r1m8qJ3o2NJ
JirmcmRVL057vlRZTK5O7CXGFhzomQZAxCTZ2ka4/+3Ta+SkhvmY53yx+G8ERmgL5f4w7hTinUI0
v71mYDSsx7RfcAoUNP5CdPnTh4awSyw95f/hqjn9QDV7iWfS9sn+28NsODpK+CRVnnjXy7RRvnAr
mwNIBL59ZtUfb0xJIhnuF3Y9Kc9KmX2Jx6KkfucNMl6OBpjhZjGnz/R5qVAlzi3viBxuwTj1yoJS
ol61CnYqyyCkye1GCDHC9qWZ4dY9ajqk0OAImo/Ofb659LUj0MDyLo2ZJlEiKk8mB5YQ3xQPvvrW
685t62A0+zjnLD1uUrmIySWt0oqYDoxBpE+7vBqMDPcTtsbSDWiz72l93nUxl7BvMh8cNhAIJB3M
pbJDH/5Dzvp3gmiLyia8AroNh8xLDKksDvk/ntMK2ulc0kzu7vNmvPGOjwjELNljra7r7Eg0l/xl
xlPNAkUBCZox5jwuc4C4yQAAasMvSfNE+wrMGYTYxN4rrk3y292k0TOjy/qYjN9toCNb2CBGh2Si
Xoe/ZAOam8DBh6ljfK+RIcKI+yzOmzroVB9ZKrLRPhv0ZMA/wbjzIHxNC3VnbmsPQpQXLZJLJkLx
sty1NUDQHt4J47eqsM185HKYUELWj1DGiFEqOhqNUnvCEb/n3GW6g2nHdJTS5VhNnLBlPbzWd8uO
H3hlJJ4+7PdxPRrubruAsB5ECMkeNSFv1XvTjLHjikVx4MjIU1O3UVV+F8QC+UxmjgN/3W39347d
B7tKS0DvAUNOc+9eb3CQkrKFAO77i+GXqm679ZK840OBbzisiat0hMWqvoSBfUsOrIehA/6POfi+
kiKNTX7ZqFqZP/fgKDbRmv5yOYybECCihnKAayZm69Lq1wOzMRfBztv67qeV4mbX0BYuG2ozutJz
xmvIhJBca4mFUIah04LHl2Q0GyxNLrzNlPkEHWeVwt6HFpw5zP+3wFFH1JkA74Lr3mJX5bcZii1q
2fZdzXik4W0d/FWozSs/QMsevVsqzIob/ko2U6pGri0WVih3ogNcmxmsHUuZ5PX+3uQjx2leAqQc
SzFHDkSmGhtMO4ow6CPKK9mjeGjaXuRGr2V7asOpTpQ0Qtzy+Q5fLKyb6GLZakLzLD16IrEx9Zo8
AOdPV/gVqn9o3gyX2W3SsC7wspx8ckGYwSvSu575ZBLDkwWCLWzkkMAoAcPD+nRIqLS+iuboySfC
i6ExRoRi59bmQA4FPC37p4lwodw1srU/J6ej4+OmpY99PAdEM48SuNnAiDurzKxcLOeL6d1IOROp
EwJ66EtZFsTxCeG5DYjV/Z/XwXvsMchYFB2IQrPJG75yXYiruKAtJ3BRo6q9Ff8F7fR+297EHHfw
s5wbtQ6RZ2AJglazXiUMgdUNvFXCkxwhv75At71RYDLjvS+uotgRaaGsJ02mSEr3q9ZmgfLWeX1F
+jcd2PbIIzgoDY+Nf10mOKDutNDf2kVywq7XP76w7aULGL+ZyCtnCK6yPMu+s+sxVuhnZW2WzNAi
UPX62u+4ksRDnov+BYhjnnGfyLr5xE28QxpIzh1Nq27G9YI2Gxsi/BMepfFqTXBLE4Z+mNquoM23
FeW+Ia1FrxqMTZgM89BAsl89jej0Ul3VHWU40HTCffGp22aEHWlJrIFyomEdmlq+CjblViKjGxpz
YFEv0yjQChKUloDWNCyPqkxubbJjgiYkfIt5ihTkVKMvjC5976B7BT51vtZj7+4Jxo3ImLAIMQtv
8QuLL8U3smniRnF42ncGlxUFsBRV4j1SRLV5W/rBMfBAOHwVjde3RdjKH86iug0THP+5Irlle3ix
h5XMIniApAb/cmP3WEf8MdKevw4NJ37J+KNir0cJXNtyIc4VSUnuAroqkwlV+Sqwb8no/eZCBL/U
6OYM9khVC/og0F47i8icfcr72k+zD1SuhkmLWwVxk1fen5RRFKzIVSDMqJB4+Qc64RPO5YTpCuf8
yBtVCbAOq6l9UEj2VRfuRYParcJ3fP8FiyMvXVlFoUjB3bHnHpNB9CvwZBjWuscmPbYgLv5Ofyc+
FXpyfJ/Nh+et1Z+Rr7gBnruTbfmi/kCvSXPfzYRrwXkfTN27aBHysk3ozfEXCQL2ETvYl8BYZmIQ
WhWj3Spp/BgpRRndy2nEK5qahbxknPRc8roQVdRC4FPLMgS0ckp/F4DwF7s5Mw3EB74S9lpASkqu
oH4xVvVPtjIPuflvfhqerVTypOXxzsmDbjbeX1+jVqoti5cNyfgPqV6rz80ZVrS8UOrjdasyGLCc
esRY2oob1q7w15kNT9gYAGusKPL30LTiL4fMo9PFD9/GPv58/6b5hWgpDvrEE05icB4ndsfiltQf
06YP8wNNlQlasM6f/YJLM8rEomkw9tbJOpgMsvBaYLoNeqyB9cqX+DOlpJt7TB/IW9zBE01pJrFL
OVU+zuGPdtR4iMl1ykSte+rLsfcmym73u1V1yYHux4JzFYNfbBp+Swp7QprL8Eelxr6iSPKwLJ6m
WUSnKq5BI5KnhlINzDq+PTX6zUK6ykSaGeMqL3IcyL3HD+GdshDqnrhdT1lkHly+VQOKoWzxtlwN
CIX1HrZz6q2erBHBt8HmwS6yLFi7XwrMt86VeqA/pJRkMSsLO1zcv40Edg+rMxO3mprISh0UwjCw
vA+c+T8fACdFSUjKU2D6w7VLuu9OnHZ/fmXzc/cu9u/7b8UQih9MPnklsZ4KYcr0mMabf5SXW+7x
lbfQKxPIjJ75s+0HVnkewhfQZFxvQvFfVHqITvYvds69IWFI3Tn5aiLkfHoz7X4FAdOZ/eAV9s8B
T1039jIg3S7PJcASSYFgxBRxgbfPnP3tkB4gLvQQRKdlCLTNzBIT6QqOzMl8tjo9wD/LB0tTVP62
axuvZnSKD8/X17AzyohFOztFK6n8Ob3cW9cZDRaDOGv+koArdmecK5CivCdvektpkzO2tVgQHMNl
Cl5gAHDPUj3Npk/lVvAF8cZHSrUxmJYAzQbvT5xOSfdxELwpXWO4oGw9HnMVVJL+q5rXQ7jLC7ri
ScfhWxbwpO+wccfOEIQAR56+d6fXqxgMW9zNc7LCLeQi8iNQixw3Rr4yWF742J+ohXRhyv0QGBSV
bZ24TrdUnGw9Gqz/N1npj6XiX+1QvBGBHb8Gae52aHjPVVIY4cuX2rCOKidG8yx8MxF2z/BPgcAh
X5ZSSLCnbj1xSbXq0y0oL32Zx2qMy2Hx4X/dXQV0rTQAxSH3ervgtWPGMYmEgZ3sCZ7Q41QKJuc6
C1UYbpSnFkna9XXHJ7QhExzm28q/be8rTjJaMlSV9llTnu1p5/kF1hbthnAieJa5B9PbTiRqm4Re
/LOQ12ajOTAh5s6nUlK+hO/EhaNi/TNA0jsggJ0l28FTHlduEIyemcpcvfh7NEAQs/uL6o7m2mGj
9FFgI4wcf7xO3SAmEXyCFMYI8OZdYAXklJKFnkldogvZ9EhIKxf7uvxhKa2oQ8bJwy3AqNzJiyzd
PNa05FFUtxPao4FSOQlr7LJ1WXtYySfeyC3ZVYg7WKHij7ORP21COszvAyBoHuVDhaBCrgQSXxvy
5eusnEDhqXv63+wuP9UWnv9XhMh+muCRWnKPIgBFRP+QtZB5vIYgeTmFp1NQsagk3rzgQFtsgR4Q
1mTmVHadtzDT5sDH4C86pdN9WpVFrXccBee5UXyBW5/ek8wrMXZaPX+b3tGTrD/PKXeHdV97A8F1
l3+qGKldB3UXdldeUzlkZmmD6pEyjVjkd/2w5a/60JltEfbrt4OZNhyI6tkIswToeppi8wghZ1xu
WSS+ZEqJOssgJJlgdXrifYtCjhq9da9Sauc+kcu9hnyPIbku+GBLSUrsdlo7j5Yl2Ys9btNBnj92
lwapgD3cpAXtFLoSjKBc5aikCeQB0l8kSBumBemNX1AsIm1x0Naw6R32Zpu3QxwvCScQwDRbHXpB
8BUuz3UMjZzPjYahyopMWCpHR1DYJlnrKLMiVKI8QtyNhv5vYRbzOhpHVFUva3vDWnzQSv3LEE5t
/lWAHrCpzGWcO7D4iG9T6pUGGuoRf75BpxO48qqHXwGq9IgkVf5jYVruXGVQOpcmMDaHulSO4rVC
hkxFxrctP6B8CeO4wQeHqlv8u+Dg6e21XkJaHGmFyBlIYeyV2pzjvucOqTmXdCAfYOaoHei5SKoy
O/wYyUwHoP5sdEnD/0bEs+FQaqUrIGKvyUNybKnPaxxqvrCCVFI98xqpXl/Y2PwXaMo/ZVhP72JL
bKULoaaeuBuBOvTaR4TKhW12Hs2Lln1DCtztoOax4n+QJtgVUb6GA5C8zS0c4E3tChBd5bbGLHpR
e3y13CSpv+QvgJtxAOXOdR4p7yPs6lp1WRbkr+w+EZpBlIUx6vHY3i5ERMJ0MO1dGqYw4c8/8yMb
ZwALrc3RGSA1vBXI2siYO1ZkTr0vPLBBhwiB8fr8n71vrB7iUPYeG+3rVO3SaD4euQoY5NwAbJCp
AHa2ZgTBUJvA0xcqzsEpFOULT9RUMsxwCvcwFjov5bstGiC5eFMYnT0NFzDkEB6gaPzBRWkGl7Yz
beLxQA1iI0WM+YFU+UM8hikT9GaHGtTfJy/zA8lOD6rLQlmM5tNUsxO4teERTJ3QVLx91jVuTuRv
6fMlH1ZbBo/s8Ef9oW3m1Q11UgUH+qdAum+CmV2PymxStQw+ZYwoXHqgnbWT5WuOjHTG8Oj2c5gg
DiVrLVNckQvGctCajbZo8dTpClKge6qfdkZhH5hkA0nRHg+1oCN+E5OzOFfibqw6p9cHVg3j5VGO
dp2VCXLDzoUr2KYqOKUR20dxgZC4H/mWoilqVvdbM6tGaTc7q1N6SvXzdgmfNT1ohcV0CfNhVC3j
P5REZzopbZKlirzDbdJtjxeplJY0E1zugUQOnTrh/Sm0xM73dBlJf8kYAq4OCAnlih0oYcGx83Ci
Tsy8u8grdsCw5s79z4sS0l6yhExvAthHeJwIaHgA67T7I7RkAqNnKu4cmSeqDPLWBd+dxx5YTiVp
3DUuQoBMxqdlbvzCc6so/yYCNYI2v1m0KW7ZngdrW588wf++PoyYcsA3EmbxmS81rtm734f9lbsP
51amGLNlHnJWNxl0wufd6gKmHX8iUSIkA6NIdirgiRkxhNhOvtW1kee/W1ocBykZuzzM7zHFP8GD
bffrg43o5K4pRynKHuYSbCVQE7w38U/NhOnblCmMEvyeVoeibJ2I59XMEwj7DborzU+OWZsE52mc
YWCAvoeQeo4txtirwlNhuEbo0BSn6sma4RHF7w9aOAgSFRsViulRdu7pL1XPnk22mu1L0PYFbdtg
1ct04056ANqGc9pdJwcI0wTqCXQ+lgZMDRrUePW2hooNXsDBhzy7kv879VuWK5W8TWS1S1W6imDI
2WwtXB6o0vd+d7EEziIgwtT9Pb9ti0WuAD0/HE/Le8UNy7MC6ebAPSUDRqjJtFyz0drtUJhfiD/8
oIDFXStC6lmPnidlRc+SxoTJqX3ezWO2H5V3uHJd7EeCsFChbUe7JMH+wDaxuoQup8ejtgCo3sHv
OsL/MomMNofrcJZrzqGfcSpl5LYMVy9/DYSliwC7Nz52dvsF4ohEs+duyz2tANBdzgOJI1Khlm4i
WwSzk+UGFfZtlcbVVfC3WeTf0E9AvWGg+gKZQZL0AbYwr6N5HvwSeJfjUX+Fjq3OYYdzFzS8XFXZ
82vXexlzhVwh2GFk4+u7rYmWLgUlLy8nEHV//CUROTgZJXBW/98oLjAbwWPq5UkHnSG8CEZp/UpW
Z9W2pWx2gWc235LhNI/RuKXX9Z+u8m+Hll2ANsj9/q2jFm3QaOCZiDkFnUOZC+bu8hAXJ8Mvqb78
3/5IqO57q97kV5IcymUKOyUz0jphx6AZ9NiMBjzweRUy0Hs3gRMoA6kRcYGPwseZ71TZMppHNUnR
2GH8l+bnrB+Z+Ht2Qm3hD9gs+dPM60U5UiPLw7Oy8zwWaC5YnYTNjzJBKvxKCX/4/Yghe83beUN1
3/tfp7pNw494zdPcetKQyvmtcKOgWHOYHHDXs9dfVaWTlpL31e+UZgsYEX4X0bFP1XaUefm/jeAm
NuY2dJ/qGs/Nxk7zkpl2YQ0wDmy25x/8r8k630WjHfB3VlB6b8uXTbhf0xjWcIhrUQDAqVHfgEpe
AYCXsmkZoEgJzPcaxxhsgnag1iaBBrvO3j6Qf7b+PigxYPZizadDkOAzM41D06pFdLzaUvfKeEmj
DzWKM66NB1ltmeCAMj1aEkZF+EPAvv3M9I1dxbqE8/sCWg5x1ZQhoz88kevvdEJz/6rnxEMUXvfM
TuZCeZbkLXE1itXy1Jc2Aduqnw+8kr4GdHSB4X040KHoia2ZMut7cWhKhZRUzWySCnKR/+D2NBod
Oxz6FrNk4/GxZ59BRIC0XfiFVHf17l0w+J11puuqV0WlOggWb7Y0U3Ke92kWlnInhw/LH47h0w/7
TAWlhtE25/1oNLYuNZhUxwyqDpWJja5gygU5+U4B57giddyO6imfdVt+D74suHyx38NGboSPm8GB
h25pnlBDSVmEGjn/TBB7vOviWvX41mg9lZhtt+SUmYPeTTlk4eJ7bIPCchd0do5UTEHE5Pm1UWYt
W9+ulHVArqsZX8it85WzC/bPeD6ok3QTiNJY3Rfq1oSNL9KWgL1NRqa1kLXDOEpXgSO9M7cJpinJ
5Z77BCUT8jkW0dhvMs38L6DQd03tzyZNNqLxy6XetPvVCuNK3Y4khzRSARni8XxmI9ck1p1X0//L
sIlY3IjGm3uYD3jIh8G8RrI1q8T8wBnua0TiPLsRYEf1xLWq4iSlNoi72BIsXGAMJtcDlpR1pefC
KHqKIdbBj4bs2l8iimHd7hA1vn++8r7boDGzb/pGjlHaA7fm9tdU4OAgiaHqUdypv2CRQeJv4CAN
/wscywyBWTELGbD5nG83J4rPxNVXNWfxtKgsISA1j+hNOUvw4djPcqMw6xZjXIwAnb5a0SH0C7kI
TNkbVYPg3MKmdO+C7QBZB7y77eTEw9kA8FL3+t3OdHUuBokLuiCpSLVK9GzJ5GfuNsburYplPUa7
4NSUKn+qDRPzOVTOKCi478+u7MUgawVnEs0oxl39XGvZO2hjcqhkRtl4Vp2wVVcJ2NhWoMEGvaf4
+K+ch/sgiMzMWinqaVQP44dmwGTJ0+alCi8ihhC3lCF6OMFNUSvJEU2AponMZTv26juOka+XMWjy
gjsfZSFAuin/d0EmQGhfN4kt5khYvvRK9Qiooh+1/n0emDvYnvdHYV7LO6RSX2ezZysyRQ6ZudyH
hjrF9G0kOHAXKh37dFHdwPiKIVoqJI44knt9QoagUZs+T0shXjyxcVngv3GqBJuRnSPSy9ItdS7s
zZfUuWQ+JE79vf+4v3sxN6saQfwQGWB1GgTKzDT+0veFFULAHZIuQtPPfGUFLk70Q1sbnxaTvUZ2
XCVmgVdZig46Sj0J1gny2nYtoGdYdDEpRSbLVaDnGVEnrmHs3tglSCptth1kvZtK2JvM0kCnIr9S
eTLE5dJYxzGmhKiulGa6EtVQ9762+upXRlHDmpU+vWzKADKU2+q1CzqvxK1mKgM8PXq9nya1N2z/
myLLVFnSeOG52ABKGo84In1r2DGe4hG2axTsI2aFIXlXAATmIuC1WHlaSFfEYphmDzmez4Fk1RIL
hx3+TBAozu4pvoLZPMiCf2DrFhwGDsBPdFW+NUOLEXPiY3HiWht1UIjIh4NURZG4BS/5Kkb0G1D+
QFLeQwfAiE1EcSAufv2VbCRAk6km59CLf5o+RHByHvbHdbCnmxW0YjmRGxRIv28svFOp31EXzllQ
stEXOSHICVwRzffRIy0+2b94GL8lj6i0ozw0IEDzC0MAm848fYjpvtqoFBnS6F5rHkjMF61BHAOi
XpTzLpDd9aJLotpXpFBDXKKQjQl5PCvUZ4MRDrZWZyDWRJgm6Lw7kRnsUYzjmsFKjvEWuIoyfBzq
2ZZsCRvCu2gKRZjz1gV3D/RKmwk19S5KdRQrTQcbwWcjCncnGnVjZbTduGG6QcEVp0vVCyrPQOeh
aPPdYwusZAxWmBX4mqKp2wxijmJNl7ICL9SfvIqCbhpPfabVvlqWtAV+JL6d6Dbo5qWL3PX8etVx
WhHxG11BtBgbyItmfITkBZF4b6kr2SjGEFnk8w/1zFpZrMARPoxaA6lJeVVLOUU6E3j8yGhUCzbe
w1byxHYlCWBkXLJ5xI7xS05jLUbcZsWpjun6SKtgCOLYgcQa8ySexnPx7F4UUDdqGnOnttq2zSrs
iCpDGleI4dQU3FQVGBMJnGK9/+hsOIB4pWPAilQUaQ/9QyGXbQnzyWXn/K9Bezn7VR9/pfoHLSGc
luM24ejesbs7scpri+E3gvwa+gug/mDXacTWRGIEpnRXVWkUns5oflZvM075OGCeRUSQuURnVspD
sFUggf+KjWmde2qPzpMgUiBHwwVlTrFQ99R+SLuy8GtcuMMMzOINyugKckoO3hCH+ztXRGtTSNR6
OhZJOTSnfqexag24pFvmak5otUykaNpTEhuYbUHgqH6izS9ewZAO3n5drYj9u+MvKtJ2VVWKRAko
MUCIplF7X3SXazT8HmHlKvLgu/ZocD6egMxCEj2oM1EmMmJDeX7UNjLEYOM9TXAgJ5bRzlVH/LsS
6QWdYOSVr1CzwbU4fJwkKvSYzVOUe/amNFXNjTXiC6IOVH7mAKHR4M2U/Wa0u80edrcZcB5eOI6h
Z0tPEVGzRM6v0d4npTFwgAOSohoAI2nE/w3aZKb69GKD9+B+ht9zX/SDEhJjPcDP7aWX4KgmRuAN
E0ThNw8LSTvVvOjfcG0bZTDfbWMX/TE13FAR6EQJMYVG5sG5BvrY5YMb4i8UEugyZtBB54++HYSL
ejYiTF55TUS4yCtm4LB9eB+Mwdsh8i6bxREQgXztD8t14SgI9UuRIEpEcDTKuz0tdie4viqMukNV
rrDqtpUdQZgDYBJfvi5944z66X7hTBr7GdtFbx3q9Ujl7l/YpS0t17ap9XkrQ4bhrfVsyRqZkt/g
aBsWW+l8xJAbTryxkoOQNziKEoJvLEUQia4Qu2QpSziheFsLdEaRVbK4De1H5Mo3p3WxADA6EmXy
MVlXrdmb9uveHqYHsBRFlm9QRp5Y+PQBwl2N8zdyf7TyYfb0YIyb9TyIQuHbuZLn4q7CPvoFsx44
WuyUxgCAGtYl5/+veZclcCXv8+zKBy+i8ORo2BnHWEfaBQXTOI2Nj7FuIPflPTHOf76tEjNUvOwx
u2jtcVuue5lgymxtqxGzRALaK2bEf8gSW6OWD1X0eAzxkE6eo+vC1lgrSTTwRM3pBbZCUGQnnACq
PUVULrKvhl+vyzymoqZiWpjKhEWTathM+5nY/IyuFpBVM0Cy98KV01JcaPHY+kg5ntjHHYl8QVmm
ln2uCUmnu87kGfmFPewIf2oOgwImJSxmpu2bKMdEByzeBM8DXnu+xmKmd18DHfpJSVZm8dpbyE2Z
gC0UlbFZ+yDnOEVTG+kxCfDJXU5zJInofkfOYbuGRlaslkQ9HcRxXiRNL7hHTTQJa/Ejb5tH5jWU
L736uAX6ELDzD0SkEDlHeNNmmcFM6vyM0vYVaWWsvHzveoN1w/3681A7Ho7fb7wPIlqsUc2AlpH0
b/Ot+242etL3uDCoeWhyf5cJOAbr5J5BLGj5lu1/n4WkBJLvK/7D9ro3LntApHM6CK9C+kqmGw/V
SwZL5C6NeKZplo7wYzvK6gFndZgAU84IwZ5dgcLm2vkYA7Yzl9JtsYPIMSywt+PisbQdOZphQjWd
9q0NW4cS9iHS2rxYq/EckYNVmMPl5GtV0hWn9hWQthBXspzxMsX1AXBYr9ANWPltayb5vxJNQqUy
uXDaCXEn9LnMqsKtEWf55YKITsvWk6Ra4kGj2WOTR6VTp6/uGqxrdAu/KfOUK7lX555bt9psN5xL
X16upA63h/uXPerH7SR3FsBzorZonPyoV3GUh0mkecNpyfC31zqFY9/5c2oMMlzS3j7G1I8rX3Zd
Kl5AQmDQwf66xDU9U6C3pLs3x7YHEQ9NQiXfD+4aI9YMfgOUkzSd3qkhBmw2AJeNIiEsszqC3rV3
A7mbPPAggOQSi+rvzG+EcybIDpS2X6RyOX+4gETvb5ITqT7HjlLkRwpUN54Mfx0iEcxc0pWLoNrR
KA88IoGhwR6qzcCTFKd4XN5MIIDmPwSvhMUf3RiBMoE0YH8agUalGt1sxqDZt8fzwyW336tI7Xjr
W7tpMZsphLbkgNBr7evz19Wyq16dfMpQ7nSQjBErmQiLT0riatqZ6Gvfp9pGCmzwYHx+Yn6KAEoF
wHuA+87yyjlPsL8cAM7S+8rWrRnuqFKs4dgtMoD96xBRtGsuP4g6RnH1H6mYChb4A835ASUbz/ON
GncZDlMfGmwHOLYlr7uvNYuQBt0HC/PP96qADPaRTuO2Le2gCblM9jq3UHHXnoc68mzQrM1EVFIi
COEpyXsgPT0TvxHGKWUmQvF4UyQcAeBg0vXp/gw20DlFCSwwszKWZnYpl+M567vz45Jb0ciOl2+8
qnO8E/+Kr1kSz/wQqre3WOzbxUbIFBujEawm4DlDYLUjpUW4W9fK5paQu14/0gNzwQl65BuzBoXO
DLA7lvFYT8w6aiHukwcSfnuoPLYMtZYTi9DjJk55WgSEi2E7oFPzN6nP2phN4XkWuMrgZq35cM/s
g0MjpGaNmhSPrjAcIqajUwsQCNgtnBF3p10pZzO8yiuBbKG6E8D4OTv2e9Go5mjN3sW9g+CH2l6v
lpmeP1/c6NUahNtpUzaZ0dm+MWOh0zVQGm8ZSQAoWBeq8z5D5vZgY4MwPnQPNrBUzZ5zTziozUVa
2euQFeO+IGspJtjgP5lMrIkdy6K9jC7BEREGjpWg6Tc/tsTn2OsbnrotYQBTjf6/4CND0RZ/yKm9
pktuNP4DgVLZOgWD7Aa3UQWlHw9j/8pc9JNRZud9dIb5M9l44+6ryFpaGx1ATsmxSeUs/6156rBR
tpl3nE4WsNRPAY424EMsweAncUgB/QiuKFQAWxxFRP0EhwdMMmf02UwKXspdx8W55SxXvYaeq/xC
7urL1CkwwFvIzVyBslAwvTUCqKu1Uimp50pI8stqxyeV/d/aIpbNSoUKV4hOaHoiwJJfIxuoctTL
QQKtiDIsWfBrZ/8B/79y3SKwamObDxx6BZpp7YQYZ6FO0IZxTwT3kpf4ygbjAy/+We6n1COuZb6D
qe1H5mOtusgckE7p/w3Zp9Z2Fiyyy+1GtDq4l2XxSDI0EZ++AQLztdkIcn57FV+2929EqssPCim9
gg+kRcJ9txzYEl9+8x9H3HMtIudiirSXp2bf9BtYzUWwoLFPLjSOYn6agLg6uoru4nn+n3uymJ+b
DT8mxJDsVtTHjYEAPcn9wHgeBdvE3u/AoJlZmpsBval1Ad4yU/8V+hAZbd6ahXM82YWhobg49N0+
UThaWEqyUYI1BurETKzPVwrhLdzyHStMppG78BG0JXi96D0jn+4jzYncjHvhAtxwui8XfRTfuqde
DuX+Eyf9mM4PDBEGsjoxkdkK51Oa99VsEIJc52V1SjbliiKu4l1T2ZAP6R/Rrjvux7d2L72DQDbw
XCLHKWzIdrIVaI/auQVfoih7ceNsubMtzqMIJWrVbuX6QJCdNKO3z6NduuAORaBa8T58TVipLcZb
E8rU8nekY4lhYcfnweNHWBWUA4qsDKmy4hCRAwJO0TopczXzbkgE44lTG2uqKIZoqqhKNgcmX+CC
yA9FIkYpjyBsnuyNaoIh4LttN9G1wnjqM4Z0y0HhrfqjngCilF+FZIVFAyBUDEaRjgiWIWzoei3J
gaJhgQl+VnqyPHWy4aDcr1M0shX80TW2I0M5OUmInc7cT+1RJkUEYMv4UurGdZZz5ikgNlkhX/QA
ZL5Y1P/+97iLilvyQlisGBBI1kx3AdgtE7MtFLAJTE2MjtZCBs9uKUEo61TNQPmeVvgsu48rfLae
wCYuPMVrrlIEONkbTcVxoUSArLPCzkFQM/d3OCJTvcGkkCod8JBQprV/x9XY/vLKqd5Gp0XF4af/
V+5ODsWfUXZQvZSgL+L03qHszfBQ1SLvVm/IVu/rVODnrGECFfRW67HslyGTfGzf4XuK+MsI0wQ9
U12bVp2mMIjrrUTvOqE30X9iDJQappxNZX4Qzqi61dyel5YXTrUOHziXU3QB5JeMFn1zJhMcMXT1
d0P7QNJLOv+3lJX/tReCQ4ZobAD5lJzgiovYmbVc8ZQQ2IBgdhcbREc9n0yLHJU4kP+017cbNmYF
n0SAyB1l0YDR0B8bn8XplPGVv6nbY9p6hTzWiOcA+imgDuVbhtwcx5bkEvKIOUNmLNl23qvRZYK3
qCD/S9thfIMcx+SbjRK94XT706eTRumygyakylTmKlUFZiwrRGBgMUZ+jMf6V/oyDOdC/u+rezDb
qHAga4kUjSxEtB6ZeIBtD+gpdhMa/8jADUauJh2BEYCHzXyfM35oIbxD0jNzlYNbPCcbIzI3yI1a
dIGUGJTaXGaAOJa/oieES+BNehdEY3VbAsdbRL4Vv0aC5zBQLRq3LGibqBu4SZwbrDVAyna1izwx
ETQCzLKrLWH3Oh1ZVy9YqjC21KfJ6/42kEg1k25kKsUzzwr70cvAtAY+Ewsv6T92vovl2g5BFzrC
saDSv5g9qCLDFEguFxtIb91SkhN1wtxoY3raC8WYrhtdose2HOik+ZFEN26KxUTvOAhMXjFyM8xG
5250vrV2sN05GFuOX7T38Lu5/pAYuFLrpK7k4cs3QJBjRIkWsT3WrM8uRGefuqwm+xkAn0L7tbYN
HXVjXuat9LFVFXJMKJPfaCX3b/6isufYrC0/yTW28RkWL77CRC0XfaNFAe+CJmpBk9faBiJxttDa
uUnV+9pMFbkeh7fD5/P2l3aGGbA49KyF62Bv+u+LOIkum9jJ7HvSd0sLzJQqZYMNjG8KDwa1Mtdj
dFPqAQj62PNkcOIe0wOrlqzkmZDrsc6ibeN+Fi09GzirbFh+Cj4pRRguAtkvaRNLkAquSdmpIHGN
FN5VyW0MPincwWy4/lLO4DlneiHwDx0tN/nCejY915nSo1a3ZKfIn9y1wrpL3O80YIUZa+BYazwF
mC3LmIy28jNAws3dbFV6qqbCfr424QeeWSdYyprFUCoiv3UrtBNsLvmE9DxbYHC1240oalNrR6Bg
q6iVr6J0gcohKz+pOIxFUwXL2LQvzMd6Z5SpoX18lF8bNEsbu7mkIJ8AAn8UpgexdeqtNQiLTlJ8
ll4WFDUJ6L3e9WvxDLJIOBK/vDzRHKc2+Y7fg0okOm01N4AfkKDME2jZ+hmcT7WWrqdffRjnPvUT
uCjQgkGhu+mVwN89oOk5niBwr0U6CtJ5sBKnKlvmTC2hFAGu/8YFyX8ELngQVvfQ5fCLXmo4C0J/
9zjpDZb0V9PXhhSoir7PrxhjbvZzoBqtzY9pTy4/TkA6lLj9MPc5VIkSov1+EMKDxyvYbfXYrreq
4RKXMocOvoCtyQZkUuNL8//yhNicsiusUENhbmxvbXKAB/kyeacedb2qMIzc9vrx24+fFxzH61TQ
NppoAfdvGg8yehtsEFNRwtkN9OrkmIaNbr6erppPzyFQKRZiKMFQKu9r+PMTXBkPkk6AHxGzxK25
D2e14MeHZiKinD2/eCB00qxvDe2Gl7Gwx3UCW0XK9chvhhLQUbpEv4L5OueGgfpgKSUEE9WZgjfE
sYRp1lh570CR2ocxWAwwJqeYIO3yeTYeYL2+T+XHdiMkSbM6VmalJjplzD8pPXg8Mh23AGoUEfWt
EWL9rixTCPJY7lfCTZuuWkn8OdCFQhpxTdlDv6bLkii5bAn4NS/SQeR2fAq03eCcbXvBvrbP81xi
vl+EnbxQczNTX/SM75qsqs6MYGd7K1tmfxnAMxDdwx5CJ4Xe0Myqpgu3F8TFwWTXOb2Xgpep8Hnp
LDuhySyxplghTeEq4WYd+40tlzg9iMM4tTrle5TnUVlmNV26V/6KJmXn+RBTMsB+yjyHbXUArb4A
okl+kWQqrJL/dHUgb/mGtwPabQuLcM4b1xRE548Slz03JVleULyZi3BJkfN9C6mTlntBT4gUJEc1
7GNDN8QWrZ+XslzlKfkqR3o+KO6noP+IV+q9uV+uqRF5aHgwrIKixos+KpE+E4eUjdTWw6NP4kUI
KLo8eH/EJfm+ZSLlY6QtxPAa/pnyuwKtKsegPq/tkVaxBEblhNLsMOHxv1aNKIlMKGjzF1S+q8zP
u9avzkKCvcCqGBE8dyoNL6AeTdD5vHZul5+xiACUYZXacEdSYuzMgYDppKcb+y/1LbWoQtASPS5l
cdmKa6aU1pQs284VvdhBZMiFK7Xfoj02WBgtAMNsP0vARSWBoeBBTkSsbRRse5eqLHBcgT8xxETU
JDO6YjjpYOWyeX2IDU5hH4uUrKaCmK/y68gLYFidhnGTM8iMKV+yFT3+mOQ2GgQXDgHZzCRvr486
FfpyxHzkQWNACpxUB6jIPvOvA9tvoIhVq6nSeGe7D3V1/k6qK0awNbaWR5fLfRan2Ampk6vxPSmb
3GgkayhIV+DOmjVUmuUTZYNfMdmuMcfyGlZJ3PCqfcnA04JGzzqs8ye2BhV/8iQvflorZOUi2GlC
hZqecSZFItAGTrh6C3qix/2xhLZ8kRIQnseXYRTJHro0aeegUoYXbss1k/gu1vAaH1dDyMjJbLPj
/q1l6ceXlJunon9y06ijTyoJGvE4xoABT48MF3TyS2nacqstwwtItc9F/ahqMrM4IhNB41kmsgIc
NVPesacmm959rsvt20ve8KpjYHt271son7UPUYHB01YwdyXJwc+o3t5bnt24dUdKsh8kOFw8bZtA
CzCQ3R+R8056pPlp5T29aZOrM6htRKd4kRsuOaTP/S0hVQHMO5PEc55L1tjtSDGFRW9y+zmuEXAc
mm14wqJhlkb6mwVL07zBWUj9daIfujr+xNSVdYoRqqP0TnlTFxkpXbNPd8nSCyn1NfXvBRuUU9JU
UUkbLWas83SKD0p4hzs9Ym4vshoSBOVFsKoRHdJBv1SJXsuN5iIOjRm81NznNRRAsBF7MueqJVtA
6HCkq8fZjqosFGNHT1kumBLjJbSbHfOnZC8Wy1hA8ETZ6Z1IECigy22BXoDRYbNFkiI/M0EtClWX
rC0+BErSooqLRTzFfKEdpRkdUbqrfgP4KSMOvBMnSJEpS2efkO1MN32qOVoqK+3dL6xs3VtSh+ZC
99tzsOjBo8uHWYz+jX8cpbr33nfIaahH8ThotR1SOVGYetEI2eKydjNAcs1nNF7cJKemfdsapjx2
LCHHDg+kZ4L101FHppasbkEQD7GhseHGTMAGlhbkbMnq1Ukzntn6Jx7OAxJaVirwmSqbZ4Uh6arN
woG5ehTP8ZTckhu/O65kg/LJpNiC6XLvsqJJuWcH3VcKZ74QUClhDjANET9DussKFof8wX8eiqlY
c9Snq7CBxyEpka3N+7tpuBQmGnFTgy8VYqotVG1UV8qC6O5Y3mUZmwt81SXBGxXaC6zFj9vBj7Pv
I4U7lOdVTRzfpU9ly3qU24qUHhuPxrFab+ODol8arWdhSYUQtEh1o0MEAWyomGz0UOlUy7ttzcHN
3TD3/tOLL9CHT/XNVr3UqaF297agpgFw/BmjHzISeqvgcKpTsnGfgiTH9UN726G69BjQSKwzrBSW
3qgCTHmGAafrVK8wsnSbOSxIwTXNgmYKvqmvJ62IfvqboaY+jQS1xpYsCtQ5W6G7ZyC4PaIZjHgC
LGjaA3AQM+FpJqrfx0HcOFLy/0lOAJdgkx9IiUgFTZYA2XvlDGZ7eHruZOKg7B1FN9ZywaARS8A0
Q+rb9wkUyEjkX3gF4n9v1LdQVBHfmxQb9O0uZc8HpVdFTx58RagIM9XSbFBvTLt9NLiCGWF3e6kH
5ze74OB8OIb359fKWWlwvxLClkDy1ao6PSbrlpKiwGhYR2buK+AnjSng5IDjhfuCLLdA7j9vPvPQ
EObAYICrZj8zKd+5YNobKcr2GUhOEdrzqJN0dB/JHqfenFZhuETLNFfyycbcRaaUoeP5KWrjjlir
+yU1NQDj0T50sYD1ag14Cy3mk3DJZuaZ+KbVu7MJwAj0l0SYCmSRF/8mSypEXTE4+BcnZhh1QxGi
OHXGnrrriaSZPErcY/mDw+v/ameRuJP4ktHf+QaIaJafwn0GDks+QYAO9nzjQDnQL0VzgU5OPZ20
INQLfecrf3JAGHOJGG8t7HY8frVCfRGFKO5dk22dQxywFFJBXpxkyW0FnTHBXSP0L2df18JK4KsM
4e7cT5I8qXTuhLB6rDDJ6i4FwFFWTQbmTjian560zsSZ8ksrGR+W1je8KFTGPhynhFeny/04qJtV
JESTTA3TnPBZJr7+zI2fnOR/OCXIfz0fa7+BVlDeY6gyAULrHbKm8y1ZYCBKrfB1sApNaOjfEkIi
ij1Yby0sI/ewqGh4dfsQBv9wWtcrZc/qKPcX07OjkcGY4CUsX3i3XY7ySE6FImQmZW7RNK2wUqRX
ZGChQhrmY4Q5KKHlCwRxaqHdgiZUBaJg8/8ZgCMBGgQkOR9jzUdFHBnyZDnNj62lpjzPX5LjDr8I
5eTIjMxpxAmVKFkmPUR/7pjcpybb/ieKR1PWP7qX+3sKhlcjPzIoqwZkfNFdmhiYj6hTkYr19npO
anTiN1xfk/hxVMq6Ls8us/r6YhSZ5zTAnXSfrZ+z6YBWybt0ubGokpt2VzKf0S4fiaIOq4CSYbuc
+7u47fhgOaOp2Z8VRg57KQ/GgidshoDXdnDKgjfDsQ3UeAhi6amkiYa6TTHqx5sdo8ieOzFR5Y7L
/0iwxnsX+aYI3hfwvrKLKKhJpgpRew/5v8Bf1CrMQlHFfXgWuEHJgTqIJgO6nOMxR5JMUdHHsU9X
6hBte8TLYEpWyH8xJqI3Lcd95lrVAybEvj3QAkCfsN1tqFKy6ISJL3y8OO99XpoEHFeMOwLrTUj0
B6q/FNsorN8868RVzRHIVM1ABSnlF5C7fiodbyPgnpw1tTAuC1/hz0nBIMwxIO2kvr6adETdYOSu
ggrbnnKokIrDeHxCtZzhM1JjcspqVl/Uaor+LVr/8JDrXOqZW+99CfCounuwL/pN42/KFj7U/+zs
GkrgDE4yI6KonwK/iILuSOY6uFF88OHOsLapHcfhTqpgR10+y5K0Wf3U89qT5+4UYQY1lRVvWmt7
Io/cfegX7uDVIGMItWfWVyM+3n1z+JCz61IoTTFJmMO2OVLVyUDJCuWaphYmdQsFZN8Oexb0bNbS
FrRTFM6g/M1cSqdEzg3VH+wW4LEn0enN0tCh1wdlkCWTFt+dUgGJRascEVjVSkmQt5elDzL1ZZeS
s6I+vg9CSLm8k5IGGaolMtORZYpRVUdtQWIzbqtCJC1we02yjBCz6GKa/0WECVFEXWdAR0fogcWg
OtAP8qV7uhqEly9lb+f6a9DbeTrZcrtOuHuZsXmTAUVtMdnidh8CWfls0jO4Y0pYDaQxVtYADW5e
XFsrTX09xRPK8bCDInx4ApttyemR7kRIljrzSFC3pfl4vbVkvt1wBjh5mMoqqI1ghrETCLY3fi7a
xflXTEoRUNvCvu4AUH9pmxKutnTIGRn6PTFOYWTlNM7uUGeTWSKIAEI6cqjEzq35mwTtWis/a6ee
w5q/sfvbsjrH5LmvYg1JKV3S5d1vUNcw4wu3gqfla5FvxKqD2DwGYOqw6GQc5dJSUecWw5IKLPdb
dEwgHCaDoYu+3W0xlN/AsC83c+KNNZMGvGzOs6DXUoT8q3bDHa1aUXhMDibbrpfIfZA1mt7gIxXY
udgtuWVr75fIMfo/LQ4lOQEHw2Zr/BG7Nlk4uiNigbrjxgKxer7s2uVGQaGpkEmpX1h26rPCWYrI
tjXWLMAktaUOjiMdlrXCi04s9uQb42IR3jGqUkJzkpczNt2cOIdbOkY69vHHcZRGiE+XFgPbFZBR
23Nb1EE2a6Pl4iABq+5JaVxBp48UBHyuc8SB3AEWB95+VXZEEg5CfbdTWSiF8kz+E6kekt3ROewc
vV/GP+/b79GD7wq6dRzzbJ0bbGfB9fS9y/BTM9fj74XSkTVWPYJ3m5aYt15TfhluFwn8V+IkbMO+
IfcGUFfvcI2EgUuVpzd3SZ71ryVMU+DIhZHSDGHCFXctmZQ+7zqPtm5iqn3PlyyT3ngl/6JEWfG0
LZdLMJRDgWRgAtHn116WbmPIsF27zys4KjzkStm0QPgFEcSwxTFCkAbLhqJh8qV7Uv+pjdtpWmv+
zCCYxO3yOHOClenI11defOruO45hJBFwQc3S3oPBj3zAGt4Aeu95goTWI2ZahseijxdHn0DbKcL3
9XFmeHNPlnU2esvrzq+XSyWL0mO3vqoygAPZmOgzGo8UnYeRJ7d5BAwk837mDLi5oj85Z69qu1cS
4SBDJfZkVTGFkbx17e+4BbjeBMVADwrCu0MHPetsCiDYdYzu2okgO/CtB7SpSUVTUGSe9wyJz3I3
H1CfiXVcht0qVJYtY9WKYqd7NH5lDKcR8zqIFtevZBaqsn8Pt2a9zmqh/Lo+1U26R1ncW+py06I8
UXzEjW6dq0EUjZZAk2BdWkjjeQhZcdxOxaEOTq8Xj2JJBy0kBr2uhevQbxTbSeMWUVwaUARbxB+s
ghspuWmYxzjKT6oC14af36gE45kOE9QB2J/b7W8vnCYYEqHrqJQvA5gS843C20ss4OF1AVyh0bow
wgictjzkgoTlVIBNmOdXajncI46YZSs8i6OmjYiW7ilZ2YizlZM1fpfGnTG3beaFzqEBHj25uBh6
CI77NGn4szXiHa2cU0bqewoJouYGkwT64r8uSs4ggkq1TAyxh2//ELqx5xMgtgKpN8yRQWA3eiOU
JuPhuJvAd9nnjvpgemnRldm0BUNEeDPEMqU7x/sP9bZXgMAsHCz4pF4u02REZzX/TlwMv1bZVzxh
dRcozxrHx7NXb6tPUQyyaZKoaV7w18jUHaiCLK7T5bxjcCkznhLoAi0PeLZ/bRwgmFYqmzrnWerH
CsiOO0Z09q1aksnsWtE3vp2uTN/ya5hEERAz4aBfvkDD3vYNLwJAzycLu+L9JCq6ALI6MVzdB3JM
UAKb8efq0b3iwyE08BAQN36AaaFPMhCtZ8JN64TVkeO2TFQ1PQ323wRMSMKDhUGvTdJDdt/CMbop
7EskWcPYCTbsOiD3p2hVx1pzBP3Dkj9aiWQVn5N40BKiJHMrPNLiYkaC+a6DWqmDBtcqCQwJviTl
2AhnED9CpxjCpniinAIgALO4+9DMXMElrX4N4iFLDXIoWCDFl1AtLtefu2+9ToBS12p3XZy4O0fg
iaKhKdXR/LGuLBmlrtugugKW5AKXMC6wmApWZWmk+ItHBSBRIDncgpX9ffFH/zrqIUucoE5hmcu2
VniI7E5+ex0ickQi0MEp606h3/ejR6U2XSUmF4F07snV04eU8nRIky9RghVK3oE6U0YiYvWhsDo/
NmEB16h4YPGNlxiJnXFue0P+GgkkFuMgiqhyzUOLjq1AQCkCX+a26EJ6PuqmUZloPhx0Ej6DqRXc
MKsAas4xTXjSCZ6nrTTYRSckS/Kbw0oTChTzvK7Zb/2kpm4BqwegZkTWlo0De6GMF07YrS9nFrn5
ltUsitcuaVL+0deSYWrD+mkPXZ7GK0KA9TmcUEe5Gdf8diUAKWIyl0Y2kWCe2j1L9FDF7S28fd5A
2xw27j7j1+bCH+xlGTqp58B9Iroyjf1Vc+GywPLAAI0n/UnAub1RS3a0KQb3tmGAbR3DdJ+G0T0f
0lQlWs0ID4lRuGZtI2goaoPeZoCpdpR13kjV39Ti/KuXonjWq99jZQR09Plb9dVrd+W059ABRZXI
9PdUeN9KFaGcVYYgQksWrpRDiZeA28vIu5F36Z1kLBHDT5LVOHl3FmkCfeXoJbUdtgum3yYhC33Q
d/jTx9UjfWsMkAJNTRrFOE6w1pl9d/m9LXSATaNiKqsEAwVM6nKhE5C7NjMil262nAogfgiZYlAR
AHxyWoK5vUV6Uczn8rNgy9gIds/BEyizuyZuIR20jeJMH4os7blKoRERiY6NK9cjPoOB2fYA1feG
6+dIyXqY5KkkUrFkCs9M8GDvtMyvicM3A5T3ifdj54Z5sNkwUDn5LInASdTeuN0KnWaIvpOET+yd
HFCSKwSfs4ydR1w9nedechFz2ZCLSFaNeHto/JL206lnjljEvPJTpRb883SP5Ewe5Z02UGGSK4/B
HWRVt1ExgXCIk9uQ+Abh4iJtIsBKfjyQ9ujhqiSibNhWwvCxee5Ng2GEl8hOvBpi12RTxA+vm3S6
Wht1PEkkPYznHtDfalIut+df5WLox0tn/QdVSFyIzptsaRSnAAQtKLCNSug/MmQfuClymDfyBpvn
az4X3R9Y9KzhsCqqhjOpMUseRINDVjF4jd9nOQYjZhtHeHEzXRX9aUKXm4sfB8y+KRoejtSIwARO
3R+Yf33tfBsoemUWNLgjp1b41aGRZJjHjCGWbMLkMv3wRpn+Q7Nra5pujQ2nm5Jv9qgvg7AW92ff
1PBy8SiUSfN7ezvjw/T3100Te8fjqSdddFZUuS4sDCz35ik8KY6xhwntVp4G2fHWu9TSFRT+83P3
RDMQTdfL7qjxV/26/mQpyQC0mk/qi914a4Keq7Tc8nwlqCfTqkS4ZYhVxXtvjTfVLSdA+80MPy5q
HV7sQ6trdNU/GiqFTeAMZt79ZHlbeAPknSft/+5LRWSg7M1m7ocQB/ll6kRkhJImviyVXfzsEInv
fbr69xCpvG4fPr0rNuABIXMbwf/a1LlMbrH73iCuJLkYP2/sObQHgxWEK3RLXVlzBhTW183JCx9E
VjZEEbAk6KTuuLt2WPdY4BooeBjpugDFoAwwckX4yF9CvCYlMONMAsaNU0/48B4OhscFSdfG9rzs
XLXU+J0YiLO6na6aA18pzGJW6SY6ljgi6oN68wJPdog5jOoDyqLowq9pbQHZdB9h9yaCOq+MmNcr
uJ0ppKUvfplQDRk4IcjYaN/RKNMGnGliDd6sLlOEXEZ4nBgYl23Vyr3cIgFqcAoda/8MtRNBDeH+
sEwAtAWvT4HlQpKoVyg1bvqOZ/H3ixva4nyCgHxb6sst51pWaVCfmU/aNwBFzWe6BYmsgjwm8zZr
cmfFpIPcMmtVcWuscQJbgICCLEUAcE9s9Sw1bPCxQg5ts3IADcpG3HzvPluXo4rLauNBLOGvrZ6h
REdpMjajk9isKjd7RgY0VLcg9CJALcu3n/iyG/aVqP8I+MNFBpJcav1aRNcQkpUvLqLtAiOoWwkG
lqFrxu68GkntVF7wdNZuj+qzPXVAhC7hSmSsaQeOm9pLTgriE3sK96EoD3VwpKRaVP1/4Z/J/W1G
P2gyJL8m+5TpqrHfqahXoglgbZhqIi06nzcURotaHR+dxIBoJAcrLvWjFV5Mw3EBo030FqZCo0gu
2TvqFPTYY6DCEouXebMfEnCvRyw26LyJFpiPg7x+XoZh7evr6FUaJ/J0IL0YEWszu7NDv2GJmRrd
6dEbe7C280HFWqRqis8Yw6WaW0IizAB9Np8RBMoahLsoAp/+ZwFj7az4YdwEnY3yX20tvJB1cedA
MhUSoe0dMyszkHy212ovtFHZsSrXfo2FF0QrxINoEdq0C0sL56CZ76N/+ar8n8poQRgeSokXHma+
0HOjgwkIR8jDYEVhb2YA4Fh/5dBRCfxxCCZA2pDkDIgWuHKVXIj4qG1g8VbvX4HukqVAL5O3/0yi
uQWBVoRZojksj+faUHxWgDDcUJbGXIH4d1tyHHykD9E6wosVzRE2w2j0h9+aGlE0cSYamukiUMJY
xT0s4P1LT5PwlH3TRxfMend+jFT3xkLqFpvBxFpjA0CG8ot3BrfU/LF4bgQgf098VJJDrIVogdb5
ltraI+FatJO021yWbtwv5VORL4BBdsVpJZF221iLo11ohrmBOeLrmyF4DcZ63rdeNVMWl1IGJw+3
aD21S7ncHo/skycBiMSF+JRFhLLzaoCHIbK2GzWTRS0Jd4Q6+Cf75HWQZfTnpOn/BCZHa2lyGjHn
6ushwOtjABpy/BXuayWE77i8rGoIv+z+1+lSDa8qWsVQBNRKrMqNeXt1p5yCCHn93xlEBtcW1chT
C5U58z/0zK01jMb6+Jz/2oA6+H8jCeaIR320iWujHH9PCPpP6WbWYoy3E1b2Q/BKjLs+hjmY5fLY
pAjLe6tVq5ysITw/MzxzP0WvmUkov5RT3fA/uVSsDTiWH1TwvtjrBGCG4E/imYzZ93ZCnMj9/LjS
L+SnUH1988FTTdKSEHAPIQsqcr3IK1EHGl7SiW08v7BcHvsRQkqlFD06epL+leQTUdP+I+D9tshz
dFWi9TO9me7dkxRZ52eg9BaYn/RmaaF+ooXNIjcNsZjFaICDOujH8wIus1KONpa1EQ6Ajw2chKfC
NzKkLO4H+GvVU+Fb3yN7oq+PCF1aF46eJ/qTYWD1gczhqfWuBzpOjUtVRm5F5GnlnqO5638Ge7OG
wYwpbKBR8rNOT9vr6k7CAgsaq3A+MWihTjTYPwwleAtr+OxYdwP+rjK7qAJ3ixFY4hhQTT8twGQT
SWkP9wr2qPtxCU3TkjDdQKozMDPpxipesMpiSMM6EnU7U8aDJJZoWCvEVd2Jx0m6xpC/T34S2N72
j4InZ2shJ0XQcoMxnN3oF4OLoPnpxKUwmzdkHl5AYglTcsCi69CKcnhy+DoyTMtQ0kox6ysm9PYf
aEMrv8KwyOWzaRTkOiYvS538AbeEgkDrPzw6ql1SAkSY/iH05BSbdHFrELeSG3UodnYLgKomkdqs
EuGiUl7Otb1+XAxyjaXm446Qn4B/C9IDGxU9/dMHjYAMqymwT4TZu6mCsIs7fSmqTXFhwo7DFwlG
4U5qC8Acyx/4IIm0Zfoz7x2XdxjlCUZIdZ0FeXQhu68UhIVTyTw4KVNRX/XnFPqsxkh7BJ6S2Z8p
ANvriSKamrznZiQ1UFzo1Iycjn0vSR52xFcjcx5YWfWWxbo61Lo9Lhn3BSMK3bWG5U1rM5RAk8yh
JLAtxrKelys+/KZJ3u3th5b2eEyEoVdlU2IS9cKs0dxSIGoccEn7NMpQzKm8HUU5px5IYJ936kFA
r3twOfPk9fKbb0GyUhzawwBOMAsWx4vP0wueUg406C4zFSERBnCAdBxcoztW6oyO0ajEFosmME98
4kimkTfHgnIGAutVGLaR9AKXIWuruOWTC1xPZOddFvYNG8Ns5kVMfP5z5Wc1bg+WKeCXWZWF7vBI
jM4zpaAH4ILy7i79AeM/Tu2gUULh02pLyjBqzjJqunGvenqcgQOL1sDwxYuJBpZ2etx2or62VMng
H+vZZn+Hnb7fewR5CDq0M1QNjmELV5aYZAh1c21qHiQtMHUTQlWe0SbZtYii61fV5kJw1K+Ph4ub
DqUL386XTv/vsB7Mr+v1NHFobJQ+M1zzPv9Scb0hErRE3L60HibmXO9Ezx6JcgvEB8+iNYSUwvbv
zmFfcMvhXxVvUdiEi0z7fk+k9efJmj5699ICuNujUZBCCH08f45jSLc9cmDiz9zkkt5Qiddl6IN0
/Ms+pFdFyS9HBEQn/tAEZEnpG9EowmwFt4RNbjMQ12212X8VD8Qkgxq1EZAuS8HN9DjdJ8BJ1YjG
V1iQkK1jOq60I7NLGQ77naOROsnJIBRyyCjyGVToger5SCt07zXky5pmgfZagUi9L/I0lhD9snvn
sIcR9nOxhmZrlDri+i3yi+jQwbSrUSp5tDlLpz0+hyMQFFSs6iNfcEIJ/SxMTjPyzPTluY9p79qb
2uw0mV0wou5t6KImpVGXgfJ1fiaNMBlfECSojaI8KR3h5p9HvVMO9Kh5n93qddWinxQJ2/f1IEww
wqHifFc+aQcJRiuqKLC0CHm/N3BjkAzK++PrSDYcFgocp1lB4QEuJ6UQiibCLgjoiTOiQZATlnaK
z2IyFabBUbr+v6Q2Y/CKHQeGJlN28yxOpjlbygfg4TZ/RJs87o5vK0AxEhU/MrInuCRy3lqj7teO
TBTIYwgQEk0n9fxSPu6F/76z90Ib2PD+l00Ngb7WP2jlOkIaMwiH3BKkd3FjqfjpyFYHGcoDDn2Q
o5ANYf/cx8s6k/7i3+qRkLgqcfaoODjto/V6PUF/KnkN5GolrmvBbEUgNGslxB2CROPascICt6jS
ggSD+xZWNymd/T4VMToydscoiCgkhk3wjRx2aQsbpQYIvsrdE+ZwTJedP131q09nA/vI/cn9IRX4
f5+KAc6O4LRlu7Ob6nfnsGNrg441D2wF1l4cStnLXRzWKrmQ1BBOtQ2LFul+fFRkVFtVydR8HeAx
qY15Dwyz5exhiya7V/baXJ2NSQM0LeMsfLSm9m2I8fDCOqpg5xxW7JwguBvblTeFgoUeJx9e8z3b
cb/t8mMin3q5z27ZNm/u/sey7d+UJc/tlCZbidyO0OnSzJnRCUW7Vz+eogejTLydXtDBTT4z6H2G
YNMcTAekkdSeaiGjPTGFP/g/Yr+u6EOJX3+jpw4ogWFDlaGK1B/KrVhY4W7ONn+AdqLPWnw/fFsG
myIKVssJy2hdLUiXQ77RPAx0W3NNzJ4kNhJZJXX+/JqbuylVk7WX7ZvAUs1vF2XGZpo5SZskcVjD
FVUeENx+3LU9jSY82GoK8iH0Zx8dQlOThCbYsOCYEoCnYwnt1OHsUnkWRspAq3FkhAox8hVLKhtA
WSncbxh6UNnRFBZIBOZlONIZJcPWaJzvXg2mdF8CR7mkxJkYLJdNHac0NK9VtrgKxrYOwosLF369
TU6Sp1Q516QKjy8Ouxr9SvoOdzH3IvQ8MDFF+gzRCeJ8pT/lpphWlVlsGCgKG5FHMfSWsGJzB34M
hJMaMiHJrWu+e05/5+xNAykJqB82M3VB8VEEztWzikCzxH0MxpEq0A8U/xn6UFQ8HdyRihaHB5HI
DIPF445HchSOL57nOB0El+J7NEpwCJ//ODvHx42HN87JVlz2fu0GPQ0vrWePxyuW1AA2N3rb3QRr
LiAXykDvQnyoV4Ubo/W70kg+YmXwqUwD+Af+xUKV3fcCGc5kDx6l8yBf+4gxxPPqf6AIguCI62kr
uv1wLBUNP+kWsL3QrSkIJ2cCHtESc+U6v0xqOV2XFUY4NtHPw7EwEEg8rFqXjPFNiLLr6E8oKMQP
yPYF9qY6eDfojvBxey1Ssuvzx0+NjFB+4CAF9AMbCoQOqkQzIYbY4z+UG68u4GNCdiOpkxq6ZEma
n0TUagBzpWoVlxZ4rAmicke1/c9DtpGdkdJ90fyJDgDl2YNGHOlP8wlkdVn20EBf6wZqd1ExTiOw
sihSpmH8Z+Xxf7Vi8PDnpNyPcqcAdWPZNhNAGGm4GCbN9s1gjdlUBl58fDx5/CaDC1/5UpPb5pNc
fQWkOEHpd+mkBEzEUrwvHy6Ff0ItmuATzg/aJY5I44fcM1lCk4DY7vxWQK6Nfb1RFmvzQ6NMSMKo
QTVDnmAjsalyKFlkdT+MUb/UDCmV5s3vFoxAlUW/KDtUmqTH4ihgj2+Kj7uVXER6jb488O9vDoNC
1eo6QY5FzBHuehLG0gcQsfFLISMTD6dGB9HIDQQw9HGu8BP/66b1K58bzZDM2DWClb/Jj+YdVtGq
KRBYk59ZmvSsbvdQgLHw1V7bULPYZfCt62ASMgPgPNcijpnaLJn0i7/3mkF4xg2mpp2sgf5vrK09
iryLRqHMKZvIo2KCmhbY0lc9tnbZE86Lr7aef3Nqy/uO7KtDJ62qUdXRRm7xZMtZC9TEw95EXaIM
glbCt7q9ZoXNsbtAM4f7h+f3t4kPqV7FvJZj+iPDb6MRFw6N5nbJZP2HIMJjR63j2d58DkYkIxgl
PxieUp+UwYQGEgNJ5MdSMz5U4ZR/IeM2gf7ZM2L6NBXMvEdCBHx0rooNb6Bj9X4vQQ0cbjwSwCeU
25PxZC0zTaxri5mE4QB0VKirH3rV+cWSFXQ1/5EteJjvlPSveWJlIMJ13QlCkjqETQ2dObWoagpp
xmRFWEvXj9zYYXgPlt/zipw+UTfxXt9kkw0ohjOhLCvX5Ja3SIRx1CLph7cURqaxjmnUNlhblDhc
Fcly8gBzmQ2pVHDVQXWNfDFZNGk0l3Cr8WGFFEYeGcISdE243HJsqHdyXi28kQpqEHHyQVuuZmS7
T9VTK9HrHEyHrP1Osu4DN7k4+/tiHNfdKRuKLSlD3AY1Q81+Va0FfYnfP2h4EPIVKEaH4uZFQz2E
hptU1oGAF+AL2yorzdVAURmBPe0ObGXVNYIsgMDIljB39LUM4JPDiXBosdSGYS4tr0zxfgdcZ7Q3
Y19S0G0PSqTigCGes5KWYIrrtTkMampGZTh4+r3lMf8qzqke2OMl1p7P0Ty3tUa+hGlynlZGgZx5
six9XvwvfneKFNAkYmuKtBXMQD4trFNL6UFp67SmjMudrYTjwbnDgR1tZb3RciPwHAqdJ0DA2lIT
Xz+sM/0E04nv5aCh5WXk4hdRAgHc3xdbOMrT+kj3MJo6ByBW6g60uAhIEUPLvvkxX94JkK+6vEBA
jjEAEcTKJsV5ZZM7fjNrKh8nyBIDErx+H4qvJDrusHVqI6ReqielOYPW7GruDZ7l3TOctDC9/W4Y
ak8YfunM55SznjUr25ND5ppCnOCAZlsOii+JchRN4LhRIFERe2bHnBBUsJvJHQ+bsYE6pDuWAXTX
lg16sIVWOiN/gXQYaxR6pG7+73KT1mXT99JKO6r9X9aqtO9OoBKF8o+MQbQp6/SAmtDCMFSbdU/v
/OBNfkgeNwqqeoRnXKkKHgg1RwHHC35WVOb40mnQS1AsBSVeIe1HeAd9esXNdChuPlkbUzRmKLNS
MAxBpHkdPtKvFpRgdRjcuaaqcI9aMcgrPNRp5eQdTt+JobDm3hAEWfMpbC8MGY2QNwv3JMlmK037
q405Hlyhdqr0SSj0Nyz5FAX10MNH+YVySvXXJ3alWkihhp29+q98em4Y010TKc+D18YPy3di5YUe
ARpb5vMqMbdQ9hZ4J+t0JH4OEeu3QeRS/x2fEm42Tj8gX9Ma/gsOAL0dpRte32r1yw8MkPSKFmE3
sI0c6NXISLFeaPc8ch/qOXnHlGSR3qoDVt+jD7QV3YFpfk1WTnUlIE4G7M4VxWRT9eiM4phdjwQf
Ta+lKMMOEzE7e7zFn3f7RtP8kN2r73eDYF/bEFBeT5aVdk0Hb2MSH6pPfKLpZylN2G9eWU6lLrnZ
vvMMYztJdLD7sey2LMpX4UWn53OzJmRrY7iRWkZSUtAazcbRQ0bzzUMsVqqeFprKTgZymOZL6Qc4
7UobIb96+UAegHFQBI2CVoktZ1iYWPmqdTEUk6DtJ9dy2cmDf13GgOODJRIt7/zIvLK+yd7lb/xU
EHIAIaZ+g+RKaBC5mfpoKyL8p6ufX2Y8y8sTMrXkQYhPlwiF94dV9JBoaF5BTYm+FzJFfjAPdsJ4
eofYrjadj9SksWpSoBM7uXa6jn/CM+q47prIO2b0JjKMKpskgeH0z6ZhsAXnQef5UHZLf9TrzY3E
kOFlwUxNqSjm/8ezF4AK/o6O0WxwKXGKJflaL4LDWWD5xUmW5dcZs+ZafxYKdTPq2MJkM7JBA9wr
mUpD2cZ61CSFiscSoINuezZoVSE+GIQ5HsaZJaDcjEnQrkh2fD/a38kz/bONDc97vHOgLc2doMwo
h10e7W9H2Ax7fy4dcUwgP13NqKDtzEYkyGwjHk8ZBs/VeOZadewPU2woGduZDaVEO0iyrZfJ0gTY
x+duXg9ZkeEmhLO0iSIeyF4rt82fsfFz3/KuUmlDRGx3kBnx8xw82EHARUKkvRZAeHm22Er2kcah
qIP9e02OnptwQf2ZjrH41xuRhNfUPer+p/V+2HIZqeXDwRyp1Lv5kYZFRKUVToOhLWWW5AT/Ce9C
5U3LfSbZqu5jXR0tbcWMhj0UZKnZvhpBRCxQYiupBxNJlDkcs1ODm75rlP0fnekOLQORvc+q2Vue
r7n0sYiG6t6tHeRgsrl1tRhIL70EN+K16FobwdHSq+yP7Y5MrVUS3Xj0aiZmzi6dkG7wSZjY3bpI
pc5p35/j93i+nHClpgSlvoFa7MKmJqp6G4NsIFVshnNQDn+t2DB2SGhHmvRp0b2TQ3t44M5FgtjR
lcfa4gA9u5U7KOK5C8y9Fyp0dT5wi7nbxYHvwtwPQdo42ToY48WnuQ3H20zliOHek7YLnFjcXpMJ
hCOXIHVxtCXg2xa8f7piz5aG9aBLRGxwYMw7GNZXVCwrDfWoliR425kngVdBDBUPEDKVRavLMjsP
kpv5ZuovlQ6whIH77ENPNLZCFtCzOFBVLjoRzY+1s3yzbtxxp1LymFNl8A11Eg3g2xe3U8CzCd8U
v1K/mdFoHI/ukIFeddUnsDVaFErPBhg0ckdsII9D3CJjaxfSJSKUO6zcZLpC6kLoZkbzmnVFc9M6
M9CpdIPfoIXZfMT0UlmhpIJmrgZ9EdUs1otS4rZ2P3f2cpKALldE0pVmFWVYTjOiOGkWqjvlwoZB
CpJsHJVaAWnsjNsSihQ/s4gBP0YaD3YWyxd9enJLMDyIoknd02llcE8KmFfvuioM2MV9v1yste9e
wYYaosdi9d/hRMgy61j9R6EGtFiILT80wS1KiysIfCxkaw2FbQwNxVOvU1FCZpfJkFa13Waz5MUM
dtk3NsAHu+nfuRRDwc9tREvHyt5OsDPm6k+ABaj8xHQ5wG3A4uzf4+GuHRzyw7f2jzacCikV8kA7
W9jn3mn6aO/2E1n++bf9s/SqXDRV1pBR4PVf1aVC9ZbzuKMCj44Gh1ORV0Jj6R2Lt4AkMthmWr7U
Lj/X6vspTuirb0dJ/bSthAXcuSe3ysy6W7KpWJzSTMHd1O2JQivKrvDhQnOK8vLgmw0XaIAODabL
pU+2H8iFotWo1aC0GK3oO9TnMELWStM0i+c/GR9tTCoin42bQO8aP/ySQIcJmjFwmIraPMScT8cn
4cqaqRRa4ZecFFJCGeiDbsvZtV9TKwe/kSrP7hLRXAXYimnj8ZjVp9R+J20AXJPdEj9Da7mowsGg
GFFFzplcQb9tk0Qkp85jsQaRE0g0qRMyCwJm8YklBoObe9Yum6mncRZOrho5XgFC9jnrjxUv1r9n
FS1WMs1jrpMWGGcYICY3Ahg1OMr5lUtpzE5jVKr2NiEjwl8o+RdpI6Zzt1APUZ/xnHEq0T0W9drJ
ih0Taf7FTlMS66TWPIjoUvQO3/aNHCw7hAQ85kEaPRck+HkM4bQBvOm4ByTAJaZfJ+fDl0tBGnZK
WT5PV3Allk9aSoS3LnHyz2uqHIQAMKr5DjhZUIUbsj7FhO9hZgsAGi/tSsmBX9BIUy1oWH+5E221
xowuWkevqeM0T+tk9gWnpQ+vM8WybpeCHZeu5RxkiTe4svp9OEWc7gyKiLHjYBtbnyosYzisSXkN
KWk/hAI0Mr92FYxgeS1RIa2Dduh7+iWToaHAGLdD4YAmIDoyHuGw5SWHjMJmVif+XPz19h/wCYjy
2xeeOHYLdzB72I4D+CRnlT8YQxkhResNicwr8/tA/LaKifRT3mt8qd6BVV2PrOXXEYSrEbBG/BfS
DlSReyLyFw4VG9BaHebv3NlUCu7+7j0v+G32zFl+6UGQUqOmVUMuHiVCkHYxQc8gCDWweIQ7qG0c
8Mnxm672+gapVXybqCb0jJgrxepW4CI2kfywjFBrgId6K3k24dpxxD3TiNRAge0PjcNjMtNC9D8F
AgvTGpSGV5DVU8GhUj9ModtPWYI8bEDKFpVF2ichhhRCKRLxnG60UqKDB5WXmffJiwGj2L0mFIas
2YKVRcugM6N4pr+NW0KcxU0YSJmUHSCUs5Ap5JDurQsbIEtFPMHwURZLRG1O0iewK3BDKjqUoSFp
/VIDIA2dLg58QyrK7qdRr0UoCdWX3jmzqsbKynimFZykXZtCMIrt5dfj9bhhxzcio+1aVB2qjyJk
QsiRsVGWhYP8JECywNRzbv10ghfT8iV7QdstIk2G1ILA9FRW2rB4rL15im3RCUoPwcOd57O//DKr
SzTfu/jqG/g/7MBZ+c/wwWbOFLwFHPYc9GqykJstAjIInWAWIL/EQUbBYvl8k3LaYxGPNZqP/fvP
oSS4CFfELM8PJM7KkBU75wl/BkxjHPZm8Zj0P+Slytbx5MPna0Q1oa58Pxc+NtEOLj5HW8uZ65RK
dLS5dWwnQR2w3JUVXF1j2UbC4k7A6Q0pSl0nx2SSP7lq8diGsicyAGtywpxvKkxbRAZ1e0uc0JoC
P7wL7ytmYpFbSJFB94j8oxYDVFyncFszeMJPODpiSaoyKeD0z113vahv94iVcq/TdPCLCwxLcbBZ
nmHXB14kfBo2fXoFohDbwG/3cEcD0FpTE5XZREGYBzNYuINCAtiJoXTrDehmV1RkrIdT2GufQDSz
YUorhHX0wMf2y8LzYwjz8AB2NoXsav18Erk/tBg8sCyfAV49S51oGJhkMqbeMXbDHUht8WeSrK5Y
eI19BnGAPOiBw/r+fmAQy1RASalfu6I+SxZ6YwDxqyYNnK/g9oUJNIk7Bp/67uPncxXv12G60XEf
noi+O88RMTq6QPj5mqcLrmDuzcT9CP/l3yPrY20/xz9ql+ZR1QubQyil6L1yOY4/vfUW+wbctmGB
HNjNterr88g0B/kyerz7KmPHLwQ3O2CbVmXXvsFSc1Wv07t8ux+ciYIQDsBcAr2xunB5JSB0BGtP
FqxzWtb2TCxg5K4QWGNEnxk6l6Id3JPR7scIHM4eRQaMpsk9VC577gKbI2KJd6S1XKwYwrawI5DO
pDISb8KAm0bOpos7vM2R8a2V+lXCAr/P9p9yb8nEzvqx0rD6rNY1TEY3JwUiMNGJXv218KIcdgN5
i62DnQholkKjd3yostnoRvG5xg85IM28+pfmf3TsEYbs21GKWRo+wHl8gSlayxIPHfVdcKblI7DJ
+6jKF1SPFce4zSVfiP108umJv7fHN1xRdqLNTDcbyGJUjmD9ye5hGReLYJEJa5yIbxB3QHEcYdSB
1QIP/NyItC7wTeYeIZdKKO+ccjJObSsBft4WTwVAOYhTl8IIwehFFB4IxgqDv5d2LCzzoUtmoqKM
mvXQfLp5XVELb9ylFY9easazFJNz5bSc8YIwYg2ICz7jqvKyspg3FK8lFy6TBRoj8Y/yu37tdiGA
XlSXm1zouZYvWShiTSRcykPURNRBrtpevDrQ5IoFO4Ewn4/2fA/N9YQ+bQ77OQnt3gnNr2kWx+wH
jX5HEzfNDdGRgvdfGCyrENtJ1D+is4ZuRPdmU6dc/WhhaV61mUVxyV2t9/yUmsabwF/6KynTdUHJ
w6UHr/HIMqn1BSahwoOynzpJDz01xL+c11ueLc9Mk8RkDiZMv1D7LW2mn8Ezdyg3M7o9HDwXXU7g
3uQ/GXMqHa0lkbY/lXsBymhwbK8a5UKEJ3/uhwlitiubPEBf/jy/iKOklPa+SHOTtSoNYGRfbthx
ZqDklMtBV5AdDH4yumqeThar8xB2G0XMhJ0bqcfcUriulNgqqLbi0xcxxj1klN0QSZkFWk0cc153
jjNzLbJXsme7qcIIictu2CXw5pyB5TfS5ypguPMcMkaKNKaotvykbx5SpNZ5dZj17Bx4vkzqfoAU
ZDa1fvDvvoTe1pYBkzg88An6THQsgZ8h1KBbNdKAvOJ3SJHhg40uP2DtOZip+o3XFtEP1+8+80RB
vOjCo8cXAB3gncTRUVWKSD4nrLq90SBgliVDCYMOEcQG7JLKcSeErXIVqf/vPR/md764rVW+3tW4
iI4OlvtSzHQ8OrTlZPTU/bnZuGKxJvNYpk1yGCKTuuFGfuSo3rawXTa5Q8sSHI+fwLuxhZRH27Pj
+LkrtiITVMZFAXXInh7/lQom2MX1KUM4cMoKlWMSidzcEtq07TCtXrxcdLGbF3Qxpm8hEYZG3Bqh
uKIumt9t8+sXNGZcb7zNnCDFrRK2F1mUHa5FQityALdTNpRwzSQaw/PP/8JXZ+72L11aOVAFQYRT
Co/k1r2T3XfjDoUBoJHREFYU/4i1EUWU/VkEnjHYzF5ua+0DibCELfQMVsvoUpgbm41VOA8ycyjY
Zku8edTPDo7Uum7IzpsczLD3EjRMABKB1f2Ouws8zQ3gQAs4S0oOUtwOULc2YgW6zIDTDYuh1TkX
8ISHuLVLcxsJ7bxbqwnDJUYfnwNuce8sqr9HEswhgi3Djlkp3tirsXZFqmKADJcflBqS74arXOQr
r6b1UzmoAk17qjEAtRQ7H96XiAvlDPmtjO59TcDL8Dh0xHkTSXrw+P8kFXbMru+7e7IPCEmfbc6y
wCtXtliF1gjQQKOqF4eJET2WtAsv6pHIlumYSM956OSSnHjYBSoVukc12uI8uYO6maRDlDqAdXGT
NUnhCyCKwLSscTcpw4ygEzYz+Z59t4MaSDWC5ZSqFjvpCLSXJjnGeY649U62sBAiX24ygZnZgdan
KTV6D6+dQuBFcdnwg1nj0Io9NsrR0FqohTGp4BDLgyfi7khB4EDYfltw/VCXdvVBPYrWZG94f8bw
qTNh0M8SFxxIPUnaZLV/6dB26d3EGQ4CPY0jsCKUptvzyTX+EkGM3Ez+rG/pyf/+DvBAu1zLOHgH
RkV9Gt5rsKEtDAsO2IqytNqTQemMPa2Zt88L67HEawLICPij5VzzkJkba/OmMum4VMxVlsJYakAe
wSj6sYiW8mB9FzZ/halL3XmFYRXPgeS8EUcGLu9enl4JtX9EJwGxKHK2svLHpCs4kBw9cBIbhtnX
0J8BQmiMVExljZ125EBmu7B+jz/XwXCAKYCyborfkiwgrbvrEZCWM5rTIGbPpcZBKpvooE79I6MH
Wlbf+YvZbxkkaxzIQfC0AMY976bkfqNQYz4YJVjmoqTO+BQEgjDLXv7HlC8Uqs030wAw1E2JuCtz
mUdtfSPPil6Iv4waTQRx7AZlssBRYQlzlq58PfmhLGrKApBZ4bc0q17uOfEdC2crC8fxCBOy72NC
wtrwsAknVHjiCeMD8rCNWJusLKbsThZTV6myMks2Naq/5qqOEco8EJIu0aFPcrmRAzUTFzAnb8SY
42FIW65QUJDVOT2nRwNn/cMy5GcWRhHgemckQxSxxXj0bMGm8XX4HvfsQrK1Cor7/nIDrWgGy7P/
iiIsZ+1oRkEJxtLvC8ZPKVnaplUwR3flboRRhsThnKiI61sG2SX1vnKn57BzyQ5r+s4hqeXG7F7P
RzUmZIntRZQ8S+oI6sRFRh5LqKtg+cPBfdzVtd7YMDkjdfBjLLI6PiEvpsA3W0V8GcITe+i3q4Tw
uG9luo5jmOacMhH7raGydJYJk6Yt2sRc03sE24HTfiJbnlpb8DUd4HoAMEx5PmJH80wlNTQlI9Jg
935gti2qIwrrT19sej0gg1vkQuWYrDjlJO41gN7ZELr0BDTHXZ/Ls8RxMsoI+MwRG72+z8vpCV4N
oSiIN0ZdXq2ucsyno2uRJ/0ugTKhVWenrlOLydWywcWhL5AHHwiV4s3GwGm0Q3PPzaL3UEKm3D4Z
y4wEDSbiy546zvMXBFB3VsKOtM+oqLypDHPCXVGTLPGWjUiJW9f/gkRzMeiCIxYcP9cgShZvdk/0
PPiJ2lr2qt3+XDyjEhLnFFgZMzYMlAeCys80qoKqfZZNaTgMSIbuW+7EfbXMaMPyczmd5QzS8Fcy
ojgvJk6CkKZpYE5ZX/KgZdDxtHzoZGUvFHqm5TIU3ng3+Xj+q3v4kf8uEouAjYidCc7xExrtM666
QFgS+9/WAApjXpaYXyBMD41clVe1F5M563Jcj9R2tRmqFS8Ibm+mvSRdfkg+Q0/I698paNoBFPHt
STPOJcmz/L8Z8PSH4J5NXWI6tkFUJmfSGUx4Zjl2Pr9UQ/31A3EhmnA6P1WJQr75+oKmur5EXKRk
pPPSJGDnw488KeEvXkA8KZKi31AIyhDLDDlFRpA1tUTHXeVgalCscEX15c9GW93TNBBhVGi9LyX6
tNZNGCNivwccvTzmtIs39nskGKqkrDOem2wWNnLN4bbKRtp+XgkX3QNsvcDLd5IE6af7nIrOLaGw
af3jGfjvEn7UqO7kaLUdZq6fCPHWi1l4PYWBStrTyGawq6M3Zisn1rjWN0nk/PZAutk9eA9KQHTg
w0Iv7OHB90ih0pFtitgnqLY/c1a8JAVNmXHxnzwlfHBqbjmzNtkuYgxaK+5+CE7+AtvJ+5DBKaGk
wR5hC9/e8dIoMPp841zcDUM9eIYODyFirFdQRQFZ5QzH9vC86Ec8QXTiq3S3qhHU+lhBmTNp4OeX
yjnq26AdbO26ezfPW6KU9SCSdb/5tiJuM9z01Onr+onwGCqvuHJTxTjg4DlcPzIbNCCqrMWChUwG
qjZ1JOgN72C1uXTs/xkrXpUG4FCF8RV2Z6z3+hwh82u6ju/tZLiUtY+pyoRtNTAYp1ZcLPgNQWVq
lMgwCCRNH2RIzJXSf7zZ8yivYLtxd3qXku3ks4eutQVdSk1esh7BfZbVWZgVZ/J5etGgFwVVxOVS
eFzPuZvHx7bsGs+UYf2Y/qBG98QipbKa0+IxPfJTEXLWq4FgslpmyCCmAqLnynoS9qg0hf8LJChP
U5psAjCus2jBpayMdc/+ZnB+T/ARuSUPbWARmszY8R0tTc1onCDQk1PhRjBb1PH3KLW0auZqUjsG
JcnR3neReX3kOqk4pSOftup5wCJo1AjM9f9NumYWaLlyUyAhwtC8k1t22yZksHGAvk0NijXzQsyb
wWDf8ZmK6MCTdM6erClms/jHvG9rEyXrZlVKwG6b1yjJzEqHFuwjomA0UD4TFug49lJlWvv4v5J3
+7LpkoY1jGWEP9eALI9u/x3zWZ8JgYNb+Ibf0hpRtEmfDRs33Of209zeYTag7zU1d/Va3+fnBkeD
749MVhqEmAnQhUefG1j/J7hRWULvOlT1MIegviB9S94dh8lD5RFa7ipJ2AaPFEG184/hZu5iVMMi
y061/quiSqfcBORqGlS4miBBKxCjjzSkXtJRwI53zohPICP3/6Hbue+EB+DFpbvviCpCQLs+4AvT
60i4f8OQQT0n3oodlZrA8Th/i4Mrd2EvnZfCUA/tn3zRR9c3Ij6mg+7EH0BBFmzqwjRxB6wukzRk
rLyhVuG7PjnkvIpnGg+jWY1sen935zVgy1dHIP2XXI8w0OiZC4IdjfRX23jAJmmbSNzgY9P7mpu7
H4aopqg06Ez6XUyawFENUR1WU0QbR9a8ivuGidmk2ABaNUhtFfdMm1Vt+XejORM9uc0lim3bSVHm
+ZFXtZXZukohON3Xg7luAQkXc+Oi7Q3Q7pdo7OphNoMvOAngwlGIzGfdBHHo202plJMOJDzAsmhR
yIsLJVo91TxE3DLy7q+VGa9KZnG6rq8K97uV/w/cDYUcusU01roLaQHFJf3x7837rJLl+MPRO7C3
YIj0aU0iXmbDvsT4ODztGeuTWXiGsEXZzfO6WAczIxSQOMqQQA5/cyyzSZVoKrrLFB4lvlEcoIkh
YCe0JPdKGIE27bzA26ns+juVI/OtOy4ZCq1M7pVEAmXbcIEjUBHHd+e9ZsTzC8Pm+pJcU+C4Fkn5
mkzoCb65WCm9E8GuZJKb/8oUCaEoGrR8hfagj8+5zTfKwoavg/wWxn4YHfh47ddQI7xqPYMbNUDk
284DYgjGE4aHPiR7gOoPlANT6J/MU+ZG23nqNIXF2SzaoFn2CxiUTKF60xf7P5xfR4oUkUz+msmd
N7m4GzF6x25KhrmWUw8jLjgVfcXW2ERUoj5reGvjpADsrrzSZUNZp09+LMO8dfVuKb19lLW3+lez
lmbI58GzYuYrANBCaUjLIIhDwbF2xB+GmUdjuk1lwJn4rPti5F3FgPdMf/m+viGfAqHM5hEYOZIv
jAE+APdF0UAidcW/H3KPAQ5d36o4y7gQg77Njq9cOiXUs0NjBSNwh5dcJWoJeZbgb0L3RtBaR+29
SJJA2CfEyb5bDuXe4PSK527nx5ToypLIpNZyXjs+IG35UdbjfZLFImR+fKv/tmCDih89vonaQRs7
9xTlmao+Ev4qvDFOrAvraSNerknFWBrHDCUdI0D6xXda5Bsg3mf7lTE+YP3WeqOKGEtcusBd8e6q
ZyixUURZJxLg58qD4dvpArn2dWCPP7ulGH8PzP4UCyCOTEhCoqWZaMclj+z1RVYvsnminx6+FjqY
lRaTxb/qfgThT2u7tVuA/TMH9RsXwGHrWbdVRUurIaVDM1WDH1UW12Ve3QwXDtZ8IADwUf9aP9iG
AX2Z0rqogAztFCJot3uR9meNobXhe8x0+etjaQI61mCYI/5r+tKvxnmInbP5ixBNZSR3F6stw8ud
OaGYdgPjsuOMaqcqHTqqC6bCjQ3fgi70obtIwlkaqdKEEfkyMRSadEmdQBLSPI7IQvjsa2G8pvln
jcAxple5O2YPiqJtSWDhq0s+6J4gZz8GAg/svSRhYSk4wHFF2hcvWqhL3TXEoPLdhN6kBijOb+cD
8YyDb8dyj0QbQWYtd6kobNxOxsSVmRtx2sDw9fY1IUrK45Lfr/Tq7xJTNF46UZI1Tm2uvZFA6G33
wqeooffUVsjei/hXqIAPsNoEIYcQNCPRZrnADM4Fb/CtPJeDbmzcAT271DetwVkziMbEeBNA183p
rI8o+eNuy7MqyfHMgzIRT/LW5F9c+HrocFeuJhBmozTan64R6eOMzUID4hnN3NdO2X3EeXN5jUq8
l68rZIeqm1yZZtLeOV3IU/X/PHqdRISVZQ6iVtZs6nKp/8Vbxd29/QXHMIxvXgXEvj6BZyhrz2Dj
WGB61RLTOMska6kyGvBuPtRzjeebDPcRYNeEnYygvA/vTRfxVd3G1rHG6R4AnBzbgnA5aXh6yQ/S
cg4k5th4nMXL+202txxW6i9TvQgGPSdTSemBXjij26hT5bHU+CulUZD9tObcSpkF22nOpoF0GSV4
HZ2xMQMHb0l0Dw1ECP5cXShvgVMOQXk/hTD//A+9PUDGuvSJ9kXjZtuj7iz+mG+rNaNnPzXs3AJv
3KwxJ/nRFfiMfWyotD2xOfd3ZkSViYVruXDBR4YuJ/5REcI8JF90p+AAq3oU3KLG9P2lYDMozA8h
9nqoNf53PWjW3liaZWPxL/7tKwR8Mha+xY9UoAzqaovxezbtj2hR4rYtHTPmcWsVZyMNfccr0EG0
JOIVM6CIh+g7Wt/xhehGDAiUiBJupjAMeSrPk72EToMPQ9LugFNO/T9JEXy2VDeVUE9ETwQ/xLW5
XaYpG1a/p+jzIaIz/JQQDjTF5MRcMPcP9JzPLyKUQpKO+MFU4KFmZ12FSNq4JkSJevcZVzHeUXaC
aZZyoeok++3c5JOSbPiXIkq5ug0inFhz71F4sRRHCGUOU2I5+zDHTC7LNWnFdsUWjrArQ/JlhOhX
V9EV5KnAsK3a36H0kfFTL/xwh6L7mJl9r+QjfzkG48KuH7fplLwYiLzTDqy2LCcuV0YZPuyfm6Oc
7jy9JhofXJB4bTK3FB+NpeWO9Qr8fA5UybHOGm4C4ODRlO+GUJjZZspD6LsAA3luTLJptx6r/T2O
rFr/0UEj0b4U6Nloj1oiG9/fyCba2y4cxfZ4ogvzyiP4ZQsRg04uh5WuEUowWyenc8IKNmy+dZ9n
M4iypaUC5sR8kvAEgGxR6fs44u7xveHd+qhf3+M/IBodTd2FxxkFBseqFHdUN8tqMJxnSEunjCrJ
OHp6YNVnI9DPSwF45+zv+AJmAWPhFDTnWlHNOKdusRIc8LBYsrtC8F7M5AWM/bOkPj1XTzcB9c5o
Wlj7uq6BnqlYdFUBBOTw34nE2WOaZCF3l40aeQaHaCD7XbtQFv7clnxWC10m6nMYpamoGSTBnzug
r8bQxfVd1tKUzSjZGVbB0J515bsoVHmz+YdrApovyQHdNadDPteGVcEoeV6sUUQpuAq6dOnGtVut
KsaItBL8Qig4ngwWPQyRdSGlpmZC/Yv0GNHrvVoPInjXSRbkZAFUXa5qYZT4N2qDZ7lfzAuFfQJo
LDkOCA67RtewZgEF7QWRaZ5AQ5CnHwqjhnB70mUw0eACa5e4GDYz7f1xBB2v14hh1IPJmPwWFxrT
jtefHVf6LRc802V4Adofu5NATzXcwxzj4ZfB+zx19KQK133LpyZYnAv4LsYBEqHlBg2AJDAiv7t3
n22WVLJElNN0iqrAW6nirMQZ9sm+crxS36y7xLzFc5vI6puxTe//Oic54RHdoX2oC3aabE6XlC4V
tQ92E2KTzGO4w/8nsACZmtq3QqaRwOTQ6KMNHKO7iOp+omhYMVgY3W1LanXI3I0lzf8xBvrUGIWI
JG5HbenER50IX0qW42h2mcx6GwXwvQ9+lXybBd7GcIZOk6ARakOFy7kGHnS1auTBBQtXRJUy7fWT
iZgc2q3nQskMy0mR013VyNOg1SdYWLm9LuLSyizx6VXAFoqzeYfy3Lz5FbGdkDbAwwR7a4j7Vyqt
W/RDhITT0wqWXnpKnFyC165SHXWKDsDSNgRjDwlmIlqjjRMU6/an2Cetec6qsX5wXaHXRloWkTnX
qzKSHr93Pt0gwdm/qCzqlfXTOnCx48Nm5eiRbuSVScVK6tb7bsrvuWPnGovAsg2iCmKmSFPIQ/AZ
J9Yb5SngJHLQ8nBq9UQH+Mrk30wVOZgfjRywJSWLxM4H+kg3ncB06H+LSme/C8WYQ7SfY+JGGfRL
SBannHh+bm9lzTwilApFfTpNfO9oxa6t36G5em9DcmR1caZGjwBEx8PsW4Ggs4Kx6/jInqV68Cad
51vP4mMT7whARXQa3RW3JtKAJHzd2qvQLrtPuC1hGI47Hro9BO9lVDV/ib53VrC8r3aF+RrQnAXh
6vZMCWD1JcydMuDWghJD4jDe1gNdFD6L96sAzJJ6SPIMHpQD8q+MXF9EkFjolTIFrqRZMh3+wFmg
a0phPqblshLxvUN+T3d4hUP9sTrwKig7q3F9wTNK1eaARQBafLrShMTqd6xVZErsoiOxQ81cAqqy
LeuM9aeeOk3sKAuiZeGxeSTc6+qpKexYezAMBQn+Z1O5ct9kOEwwRv2jDYz2b8PmgXj+pltzQG0N
Ma1DArs6QfjF8dbQnh+/6tBXjXm8C8XuH6/W1zTuHUcz8stiCBF6+AUtSgwLMZ6kh78B3JX7JGWD
A8dTFwQnTzDuAO+IHrxl3Nba5ZBDKNUkx3jRm/KRvSyhPhsNxx1BaZLaaAkOF4ctjVsj9J78ZkKz
2bFRgc5krRiFIpSGN5dtJIsHwg8PQv/pspIeZxdt+2k2FceE0GSB2gRkFHud7V21MzzIEJQIp+xa
r+QfW3do5ScuRJsqxgK0m1PoKoBBa70IqluUbvtWCfxqpYMuFSZtw9rB4UFP3KDA9RsQaZXYJwqr
XebR4f/6Sh63x3NqjqBwiB4yDWYZhY9z3TIOBgdzRbx5N34W5QIniBkfHwjUMAZYGNWLARE8vspl
XA0/xRFwtVonjxW9wJW1kFP5UMs5W/UMRWyWYlwUuASc705qpT1bziytn74CCg5CP7/Fen5zUCEK
frQdzDOsN2sAqiwgeMbIgpaV4TOOpV3s7IBNUquyqVJ9E0eMKXCs31pIfNdFWWBQf8SgKZ+EVo9o
HaHJuRb+bNinXiYGavyC2OZFTZUlxN8/SfhFsSiD8oAWi6qpp1tJHMLqV8yOqy3bXzCjNhp67ZwZ
4lFEPKx+XlYsmB8eAuiwEh37sGmhVdnWZQux8RNTGJ/k/AenwJnX9Wn7tH7yg0/VYQo8h6y96g6G
phFqvHMblXwaUl2wZyHHcPbMEq9taQ6yGiDO/x1+73BW7OTeMA7r0PA0OXKfyI2NrLNFInmxs+Fb
Jqg9PRNjIL1rWkGX7/8ApvzesmMpJLWX2uh2clza1xvqmAkHDvmeLctV7g7EDbC+1UVeGhgNUVrN
QB+sBeTVCZ4Q8N9BR7VbnYbh+ttRWlkQi17qfIws+52rSGN1VjuFWbwfn965hN1TQvECXc0OnGEu
4Lf2yebZvvQNS2NYZ9vLtG8a+bFivxMy45w9iNjM7jHNkbyXo1s/RRXv+M1JmEgW2UGPB6iwoxAp
UOc3WB9AnXxeHJT2pEeVmw85VdznxmIbiilFQwum5bBXFvMAL/XKyDrtyUMMfvia5Na+Bj5h9Ay1
KwyxuBBqLmdhX+9eq7vWjeHIFIhoJSLyglKtxOq4n+QvBA0wvalLyICk2g8YXkLJMWXjj3ZJOMq5
uByt8KGB+PZFk7N1OqatqnsMB8cP73dyT/mXDK72R7qBDuZXuVK1SuoFO/1QrZRaf9btNnHlhZyd
8/jG/LlQhZO0VklTGI+ljEWJDJ89hy2tN0P0wwDFVzDEa7bOdA/afShgj1UQvPyWdp7j3+xGZjel
vnDCVPWVUsoUVzvRN2b8BLfuXW+U1ChWnFkTK+KFAb1YhCkDWNMS8rEa6olP/IWaVjUM1Pp8dVQF
orxKE7IuHruZBfc1e0vdL79NPcE7GGCXa4/2+OQIgazrDcottUa3hDYumW+LjzYaKQ1iLHqSk+Kt
rBSTzJJ72HKFqlr4hlzR4uaLY9YJgII0As+JIG52zXEmnzlRabCq01GMSP/e1IOIgyryUmkjsWSG
be7bk556kSOngXgLncBdVwMrXBo6AD4xvjIWHdLfaT+UESWztrrrbkQjbisqrEoDV0rvoR4TJWYw
OLsU5peEdTp9smbkeAuu0WSXvmsL8yzz32L/OIPi1U+6SCFZvSTMSYvz2WGYQukCSqiSuPayNarB
zn6KzgLmiuf32FrLZysSRmixdSiitL6lR/9O4S9P4w+ng07TghIsz1ocU891ME1r3m/fneKpBL7u
+ueQ4/uclZoMdD7SnKG1sFOOxPrwP22Z/K1v5xTCW8iE+iTVzJsXAbMJdW4eNddYWj2tjBwrXcsC
ESt/c9xzYjAM359yYK2or4Av/4YkdE7adY0vC/0GOmaHxPCeLao3jPQBf74l/rpHW44Iky2+FHDx
fPpd/4dr7flfaawdOc/+f/IzXz5YGrzNaJ1tf/7q1rRgMfc9sfcJbrsLxzoeyo687bQypOF3+xzG
yoVgOYXqbnsh7aVMEwD3yN+OxrXx4rk/1cREJZzytAPyyLeDnfb9EoDsDiFdSmgNLTl3dPkLlpIx
pfHh/J8odi9tS3Q+LIHiNhPHtN2SUio+B1k5LbYbvTv3LLVo8FOH/qwFUrSdTTVMgKE6n11usDG/
d6M/07mYRlmb4taGCu2kz/d6IBpmUuW3jY+1/RQzaDXFsUJDEBX0RTSmYiTgkdlXzFDQMzG+vMBV
T3wX68sd+0U+4QInBktF7DaMqifqbCL2X2wT24ToDAfPqJx67Gj5cHbOwFSbqF7lqfFlWbC8exQv
pbA3z/5qCA1gcNHqWX7KqYfHdeMK3soqs2DZXPx6OZi1PbC7xAZVETys++NLDm1BChj/DqjHL/pq
YTprcwMqYMGbWg6+kRFZFvyHaGjEmmJUPHuKXsnFE4YkhRFVvVWhwnKZb7NZZipLMXGwy7nGaZZp
bsABu2WtvSgW8JZiXWhQUADcL9WvJ0yFp7W0m0LZLmyFwsKqrE0ohtcfMxewnMbnPT1UJobAN+sg
0qzEBPz+fbgniGUGZKncMbgWAn9o6+vAX9jQPc8vKG8HihK5oNcjXdHswJgco1lLtCvpq7LCJ731
dh5ISeslTM3tXFKozNZWvqeImLqzHVR6urOhlcUYcVdV+A1yw+lqR1kyVcE3tXNMNQI7Pk3yU7eN
iuT6cQNxJ6wyzSDkYWrDk0htH+awgkc8aggQOG4HZZOUTEx5HYrEiJ38kqw4HsPFYjSNad0LvtsU
rxZ8CjbNZipy5BohWzYZv7EMEE/j7uyMaaVOuxaETlB7/GqoLc7rHOwCB+RHYuYwbfyFpKQVi0Uo
/MqBX4B4tbrTQu+JFnhQsdAkaQfBwCn+3JxQkRl2j8UjqJGFTlr2n/m9l8q+B3rcC7NFXKMYrz6v
8992OjKSNZhyTFCIz6vp2553aSAND8Q7I6PGzqsOj3HdPtnyFaMgbkUZUwg015iJcfKWB5oQqBAk
tXvz+B89srSu5Tn/psPOGseMm1hkgKOdrrCBeHnkrHT0vZjvy7yIaB/k/1xjf04SXBiy6u2clC6D
0Okgmn/Xqqisnbb78aVpikDlp9ZfSDL08bE2MbVNFXZlvxAViMa880AJUnVsgHZDGmPoZLi2MCew
/T8jS8Tc8eQBsg05dU2eR9gXxLF5RF7GTxShH9kGuwougd08f2kuWd62VqykAmLG2Ds0b8/VwIcA
aHcyihmCE8oMw0KObOZRLsA6TjLKCwZQZmfpKOMy33SnVHo0Dh6ndW7rmYosJLy/wckpOQl5O5yu
qj8VY+UD3Ntlz1YmfufzJ7hQW6vZ/jOT21/UUsQFuudLNITSD+gTKOyvrFmwaqMnPOm2HOxMMO/P
jopTpfvudzdRTrtMbMrcTonG2d2hok2CVyQOgA7bL6QHfQpI+YMnv3Z8DFRh0cyfjMGI+qaFk9/T
7iRh2Z+D+UMY9avzE7dNqDfjeL3b89cnssT1o+nPFulOH+wy7tb8RHJuJ3bjY7rXZR8oiAtcwHxy
2eP8z2poapnR49SYo+JgCboycbLuf7otvVO5XVSND6ypJrUxs8asew4fTlVUyuIgMCR8wKPubaQI
UGsdojvHPLr/VckrHb3a9Z8nz5g/iExlRtwirVcnpUzgaCTVLLmEns0GtHJDgSwF2TZyaZeQL7My
UKaTglkm8bdBAPMo7CtiHfxuXhzPZBpETqzgB9XY7067Em5bldGcFLiNsyGSm+OPdfDz77VjBFaQ
fkhYR3V+kocTWN1N/PigIWv9bGySnWihabCoYmkddcuuap7iFSN+zx9rE5jIMqTrzDBDkqUM13h0
IhiXpbudUPHeDz0EcEWrsO4x+j6m5PzOV3lGpzazhrPlJJxs94NKz+8hG4ZbqFI2Vg+bXG31l47O
QDZI2UxuoSD5fAmsD79nwAYsCDV3YJXbsDPTRfVxGfZnGCcqWiHvsZxbhuOI25BbAWvs/CyRgqmd
9H3dXqSlNJmb5nxlsMqL/eL9gB74Ce2YwPUYt5n6tCk1prN2VLD1aVNIaajeuAa5mqDVRCsRC8E1
49abKv05CXVCs+xZOlluDwBFdWGJj4+y9xbXkylBhNcT9j10h6SFkmoXBus6W8Rrhq7YAr2uhXgr
ivrjNXQZ5/Uy3mQSiRTBfxkq6cfd5gMXRJh6Nf2/00igyXTbEIX0uGkMYSPuJHWzN6kxT/O574Qg
ppR/IPTymOCH5USoXm/Gln3AwyuoAcoa8lykIKztD2nI5q5+KaEuUZ94woaaPfyB82yZlSIudv7P
QJmbmhky1ftZ2vNvwnqJPEFxGHGi68mrY8wXQ88bLXn8V64qK4u5HSgkKm53O4odbG9u+EYVYFdZ
L8b5zQVW9H8wjx9aZtY08FLeMMnQJEaEtVsSRDF0neyOkyThLM5AJN9S2ONZED0vhHsRUHc5Gp72
jV2qzT8esz3B+jrt7T3IxPI07QiLL+Nndaelik/EFPGvvi2Yeh5fcflvnc0hPN6R6awvR0CA9jEu
zJsRcjtvvoaHMOY7HkW99IrB7WjKNu2KUrrFIv6mDdt4ZyhM4aakJ7+pTHGVgftlbWNu2ZC+qPfz
6YHKy+8OH2eo5TsFLOUMrvxY6Ts7t+XCg8aXsvZnN7PUDvk/Ndi/2CVaEBVIG/pdPGa5WzfRxGoK
q5UqT2q3LD60b5tmTfSXIumI3VvmfQDslBtZRmfVZC7J56lI1zr7Z+rN/6o5raJT8eoHr130g8n3
eNvZZucRnnaUrtz6n9gCcL0CzAUHA6zVZMXGX7mkGKS8Fy3uEVpVt7UI7qU5vcTtdxjHSJfRUBy0
VDMp/J0E5JTxm4fKTjZf4Rq7bvjzYzQfxRHo6fcxMQi285+FjFt6kV3/0Y00UymCb2r91MLzpwHL
+J/Gpo2417Ryhgrvw+tiYMhnNQFTgE9503KZ2zLmI4PR9prA4ObR1azo+p7jwPXxA8KcN/a16mrD
0ZNfadg0Rzvwq5/4qu5aSTipKGgcllqUc64+7gMxIXC9r7oK3p2JSMu0mRThmKVEmnw8kR8taQAB
xWI9vG9zRKOdmQei+0cwaTIAbQfgHYtbyTiHfHlyjE5APZvI72Cv1ccm9bV12PAa6oIdm36AyasR
aVdxD96lMjHj8VCZhkf9yMvIPtRusO2PQRA7MsV1EfrCPZJtPRR3I2uJVsKps9jRquFn49sBqvpS
EQKtXli+ekoMwnubg1snLRL0h+6dpg6b1pSOIdl5FgbQlacyLD+AnMrMZuGJXohDlbyj31ow8oMx
M7fXj4wcIi+go14qGexbSrrAt0eGtZEKRfdF/P0iJynTJC/cgz85VT2s/8EY5HC5j+9Y6J/JtgrP
oqhqp3dgnDKh8BXfsfYrD5u8+O687F8JDIndpeJ7pfd7tTRNDAfTfCt/EGWk5DMUyNMvTSPnFWs5
LWEAEBu6kqyA+KrbazRmBuprak5vtyYvE0tNnDkJtOerhpjZuWKFerTW6aLT13ZtXLIZgeeKQV8K
rkKDYmvj9FgQyIK7cnyDVBKdXClnN/ktNDgOliSnZhrFJiAFm+h4EUx4VbxuGNurvFQdD2hLFkcM
DUisa3qpQsYCHRdbMrXJ7AmR7AKKr+5nryrG3REovHPfkoYXHVXg0If+zY+EjhEnaPIbYPgr4R/T
UeqT8mCUh3DdaFNjI5wxU0JUYq62LAIzkxBz1uiKyt77mCGd3eKaAnMQu1U7HEsLS8sGSSLzUYIn
g2BHhwH6Ivc5kvP19vZhw5VxEmJJMAXCw2EmziQYUj09IFCj2YArAlt78O+gpK5S/fgQdR1FRmI2
JqxaaF8iLGQWIfpMDKyAETRXaV+MYd+KqeCfyvf/Wz/0LP+NP3iTDczWDuilBGeePDLPnZuHBeOI
WKD9UY20YAZYLq5nwcixQGqQjNmwJQAvrMGP4QSd04t4OT1ZlyKFSLci1X4DtkXcrUSTgoFLNjwG
OnJ8pTgawFk+LGvPDKsxJvjPhtnMp0cO6jE6TaFXAWq3NH9G2TcV8fekOKR9/rDPFoPCYEyXkT3n
0aNhmF0+VlTQoXIfrT6fJkBHVUExqTZD19j3D5g/1M5p4hSm+SlApQUwD+A5g7TUio0pbAr329qd
zpruJyo5ozuWdfQD6wHQd4PZsTvfq/tgtvVd45tsLUYlu7biW59vArTzzNc85jhLECZ40NDvAJeZ
7WGv7XOkPhbdGct8tPOqzG/+UUG+aJUBTQ7EVSt4VuQiOUEDo+KpY/nC2EQlkaZtRcHh/AStKjKP
FiFUGw8C611rQHrIxp3vBXs8TL3CwTskhdy9Oj0TRL7IhBKkjiIqBrKUAyV6DPDAAi3BXN/fOcuZ
G68yOJ/LPYkE7yOK7pf8mYT0lRWxQ8KsRSnJ5S5/P+Qul7k5h22MeT1/qf9dEp01NKxxgfHUdibU
AYZWMvvkhkGSbA3rFrGPMiiz8n0qOoJ3+SzCt+GauuctayaKmkERn81YhEHVhKFrjtpiUX30bwku
0hwt2QDpChcdwQcIpQqpVqAmPTRYLzE3keQR8JHO15qRu12D7oqWOZzlZqPJ40SPBMVuavyp1fsr
CjmwCFTWCYrPvYrh6FQaCMI0xIDwhNGCmG5RkKjYF39VdGb3XVpcNRLFnvqibUBiHGI8IL3D+Rvf
3pOHYaZ+vYc0eRhD5n+FdaC06QfX+tvrL+19oVyNbPh9dYHv5+/3YyfwQZWeLq5oqnUzMYCAZBdF
LXoLCEtk6vRH4Or2AybFFBQrtU3VwvfCJQoqD3lG/6h0Umy73Nqccuu+n9H9Fgg9MlxF3yf4luDd
udd9OZrdVto5Y6sFZmix0Nf6z1C5jycPJfZQcG+8MXteR60xlLFcjyEbLn+BbuQmchBMpDChbHEO
olMKdO7gtqz88ZuBO8/WOBtYN5af4r0Ej+5zWvqCdO6dZoAEd7O07bjgpDJFthFbcHWXiZ0DLt6z
+qd6A3zRzPViyOKve8Fif4cGEOrrH/bVWUXV8iDz4O4alMfOesrzSHYJz1eGXTG9dHRgKNm/4A10
twSzJXJuRNL26LjXVJMt7FHBM+4trDCTU0tT0OnWLPN+o13iDpHn2u3HwOd2LdRt8eXiSsZK2FRZ
IYZxTHtqTsWytcvTSw24OPiFTSCFfaFrr2j86HjFIIXIYGo4O+2w7gHIC0PSCt2a0B68eN2JjSpK
akO579jp79WL2L8WnjNnfod1UC+E1Bxeru81PftsYlT+27wF4OXG+rzajUQsDLYYHSDBasvw5b6q
k4qjCKc1TZDqwwFMKOvARrBgABRF8jfAc4Ze7hNtxqvYxnKV89q4urc7EYCkFQ4XbTz2vwU0qEAn
OavOCs9X6GaUPXmXMKkD+RqWkbjvIT24uDrqqHpu8DYdxSxtzZVb5RndrT+pvw6nQVhYBXX/600M
s45cidw719acnFidzzMTle+6E4hOXjOwt4gWwkwc1bXtB6Q7Vq6J+9oRqX5jNZhbhQVMS6GJEuCy
TnSR0gKgGY/9Z7SrTCtl47jW2qlCVcSM6mRqc6Yh+/gHUFkCIpM0yQax4o1tXJw/dWP53vq3VcTs
pEmzOISjT3CvOVUVssXjRCOYKEYjTnQYuBVEC+udS+vZ/0Xi4idtV+utARidv8EHBtI/tE7pmLc4
Ngh8jk8QlLpUt9u+Ui/Vdno/Eu8RagmY5Pm4CxuSLjQZLx7ayJ+fogmMgnkTMCkqGyVCgJgm6h87
U5DLDhWF1A9DcqS7MBfUcSGww02gBmu+dXacipsz6qPiMAgpqAoKo2WV0jttmg+LUv6TJZ3OCxMZ
SjcC2OjBNm+zog0GaAWfvM9fvaUgLIHzw94Ugeu71Xn3Hg0lX2KRuKrEOPhdypQVKA6b7kYggu62
hKCoP2mVe7u5cot3JxEmKd6fgrJh/z22OG2L9tyJs6HjfZKKWLJ/QiBGCZB/TJBVvGhNCXUsxLq8
+0SHpizOUID6gwjq2+kG7THIJFZWXrfn5mSNr6FqrWqiHRFFHhe/AS3Qeg4F3KvOyblvi/3mKev+
R1F7tuQ1JhdURcVBqNwJL/cyjDBaNS6IFLA54SjUPup7qqn2GM3hHLXiNxmbx7kdOXMrGBNMliQs
69Ih9uEDVx6IIKD9ISDLMSPL2WBPefrB4MNxpSiVraj575R/Ki/DQ4pelb2KRuxL0cXJUUuzHo79
vcTiaTcWU4KR8FQB2O/doYoTE+dBxbyZCo48KW+0nyRQ9joJNKYOdo4+kpM9NF3jwshhd6Jy0KjJ
VI25ha+EoUPZL+ug/94ujMXcx+Yn+e1xvyJGX9Ars2n2Plog6pp9DlwDRyr6ujHtkpqtHCKouv/O
yfWPzutFhyRj5kol3cTa131RDVvy4cfDpnYd5RSg5PC7JgQOQNovLtNX3nUOECltPjQpRaBY1CEW
QiQRyfesHF5LfnCueianlClHsgsIpjH3zuOh4MkGWRM1aO2MpoSjLwEe3ezF0FFEu3IJy+L8LyeD
gEZEJGF4cuT9rYlNIwRydA8CNaM1HtldeBy50xPS1A786PCAQnO8y4ojfilmaSqmhI0R+cW329Dr
pjtJGiAUPG2SlENr5kLTZkHr3Uf3rnT5i2evHGB6MT1y+tTA7/mp6G86o/yPmYAYHQeiPRdLil/w
+rZ/QDXrpOtTpP6NJBuYk8pwzBVrNW0MwyLKfSTwxS3k0N8HOJavVlTpCKVtlKwxlrs25XaK9UQ4
C57xyMvK7Q5RwTL4zMid+god6x7zX4azHRzf4KRJjhwmavhdjaz/6GkatT5my+jBqXBgnWj2V1g6
zLvR2n7wNMzMBXvpD3YfpMKNl4vzEBSCmHLK9HbAlv0iqzc6ksTQAP5nDDxLJKJ680w436wy3We4
plQQNDJgcEWC/wYswG26D7VXKWSR03jau7Cw1G3OyHwVbMN5TncluasHMkk2vvLpiPI4B7gt5mmL
dpUNiwVfbJNi7M4X7v88il1DuQY9TPhGrnVgFQjiIQ2Ecu6BQmMWbEyzsEBMdwlW4tMJrjDMSsrw
NVc7KBzfcgxv9ZICiSc38eOpEbYMtb5ZZ07F6OCN16jcSmkf8MRpY0jPCFYWrKmz3AoM4IW8xH46
I7Ea5IFEmxChWBojRW9Mfa/11cwUVIrfyXZ+lvJOFox3Epy6LhOE84sgOZOtlbXE3VXsLlYw7Ic3
/x9Q4kjfUaly1M6zOjFNzJ62IXWGDDuUIQ9CPahQKt2M1iXtjof4QlcaEBpXh/eqZLHYGOOBiqnj
KbBZqqncTA5wx2dTl9UIJo7gICRjkUhpeJte1CbXuzcn3FuWtIXeaD5tbF7frPrCai+zcAab/uEm
DHZ4Y/AYtDWXGz0PTfFQEhENbgnijM4IHIfGlB2jONz11y/EXEqn1w5EFdG0lzN9H3YoAjNwhrO9
ZimZORIRdmtUdVYOI1doRs5/GwWrS9OGyu8vwLrhMKDmJhO36tAq6wXvYdWMisGQDe3bHtCDdAos
FBOZlWmg1Rzv9KSk6Sd1REUJG6RyYVcuovoRMl2PxpaHvvzHj+jzZOY8NyZ48u92scpuEjJ7CwGc
uytl0YaZcW2mOZY0sswd/2aE9UAzfMBMyqr4RXIf3X4EZYUJUtg5oR867bPYLUvTnA7f4PSGN9qA
H5g0jdW2smGck2SyqQu/dIaFQh41ZnIkuvASIfcmCCkY8MuOwQDOERaKo1+J2XM9dYF8lBsBxa0Z
SzwKyhzB/oCKXvvh1nMozagGEREMJLfFPtdJO43mbVFcj9lTf2oPFpfqGWmrAosbBOZgT9nC+KiQ
B75bt7fVpoT5dAXsOcnxl1JyON+39QwKrBDX0wHF5Q6zPHkCGB1gqUuz4ccTN5kB6tttCXH+hdgm
NbLYnvwTsWttj3oj7AD7+6Oi4Ft6oRoY/LstW7kLkwa+ouvD2cNg5pQR9FXDZPPivQjpK7F8481E
H2nIP3vEJU5J60fyimq4mGFmHgLizu3jKqREluY92eNS1s8YILdqtDMtt1hD/hOMstduFVmK3nCk
IY7TNLY8O8zvNeEXElj6hlA4JTjp6bSq5p2J1oooemqWr5ALjvI1GJubSiYXecXJ6u3MRRiYb7Wc
gm04isu38LF3pf4FtIOoFht0/Ph47+mmy3JnqfILN9JKmk1QvjvuIRzZV1C+7fyR9AJWuZ9pXV4f
M5PJwSX9DeWJOBeKce9BgoEbWXkunWGF6Avy9yWXQHAnHECzTG8jVpEutLS6qNwTs//6HLMoNSgo
4/KsgwnnwZu6et1MuQFQLyn2cyebkCnpauK6mO+Kyhc3WE17gIW0xArZ42rBaNHKzyysEfGoPOAc
Kxf9LxUkzVSjixxOf/e2lp2IlEvJBshov0hepl2qw11wQCMjh/9GArvm/I/0KEU3reaVMfRLTxmL
TqxwMjRFgXH6BGM3qDiNxTTHOxj5Su6MhQs9OSyjd4P+SokBsTkmU4ePk61Fz3jrfRKvK1jlvwq5
LaIkHkZytdxkX3BCxljXg3whRIKmWls/PBGk3SSstqjQN/xexz74jQ41qgAXaa4Rgr+xmEN0uGiN
wDT/II77DzOTgiUOvEVmA7ErC/u2F5idLIZm13lyunZKGVLlDMSbo8wHjldd+V5d+z2349uO7Q7U
xQOnaInk4yHCXMfVwOoKRBsFy1489sbE8d3u2ZaVfLyyzpT4zPexTiN+vbK39fYTplTzuBoQ5afK
oUSb8lUbn16utGxh4nSRaCZrVBdnuDatthNeSl7e9lLHi+tVShc9UC1eVnf88QrRfMRsA5slSWA9
bM/WYEFnVl9nUV8tJ7IbNYwP4bVDYnNhwK7ui+XUjkhi46XZHlsPSjG1LRBFppDsX8eRcRBPeGUW
3ROlefI0rMXhMGClrDb/0ejarnti6u60/JyM2i+1pa7ur9W49nbYdXjzQ8VDo331oFsQ+/Yv8Qk1
bB7PqvS9VeQqRQej8Sf5WGXrbYuRMAFsPfmLJi62AHj00o5kAdUbAFNWPZ8MfAHhknXiiSsXpr6B
jNKzItMCQ1DPcFgrhhQJEin/jOPG88wYmjRUxG8o1smetTch1xFOsKye4r9M5Ge9wjtutRg06216
vszrPeFg/7jriMIZlbisp6rXKNOCRT/NQ885eP9vJ7AcOUc4X8+Y/JRp2EhG0VMsaSDBUrDPgmQf
BMPAi0CWRpxmkhgQ4ppwsvFySbZP+gDJOp46h4Q+4HiOLCTHgsDS/15x00frvNMREDSWv8Hrhp6S
1MVjKZfHSpQ4xhHrfPMT5Yrv7EUnyKsl4+zxU9bGZTRswmBrHd5XDuw0JsBmF0HPSqcW41z378k4
OD1FKmp0+rIuagbHATmWpdUGuxg50K/Vu2SRymOLEnxxTMg1XLolGlINDA7BDCQtA6wsaYj58Cjn
/FPCqjiZYXZMim3cCvU20IKSCVbaHpfPU+IFbRSXOOXvL54fUI9y2zQYglHluyMssZptDV2DnSdn
uVO1W9svOTiVCJf0p1R5MZuljczUDL8+uItNPrQMcdASufce2LiWEDconbgU31PkY1Moe7iPRy8S
YNJjbGG/RnZocVzDA43ImEB0B+916qYDb5bPNlLX0HEqRgKIiqXIOinWPA5dAfpM8J9LCrUUgeA5
AmPdWndaUN5GeXVtv6IFnWfitVz0gGl9YNxmIzbpxWOA5Cr1JXK0iYt9uCaqfMQYhmxKjDLc79eR
U+dbRisifPpc6emQCAl/INmiLT/6HEYtCGlp1iTcfCdrzgGRExDQ57LRF4gNFeHYpCpykwgM/3tC
Li4szmDh3AvtUF0YaHCMmPKuyTFDBDzBG09XACSfyDnb6xx60LALFdJe1mUz3kmg8PCRLPzzQn6h
fCfTrLtxurQmw/lg2+NPlxIhyeeFnWlHWt7eLwZ/fjntGYruZm6tZT7XZK5LRbnzFz5JC58NF/D6
T+PjvmgxJCqRAS+g9OsZzQMUkSLqlTRpUx+l5XS+9rzzbYsZrFG5twG0o445pxYNOH65cdVTj+BL
tnYounwQItW1/5XyLBdWGpQi7UxuRLMoRlpN9/sd096cOINA17+Q19Ll4qvTn/vCccva9YZhAnbh
kGeIm/RgAWh/aFHl6t0JiKT2g7H8vHqNjZSY1hSDEXVzZdnZD1W7KPzbjQ1DDlNVsbWH11zOZSwX
ILZ160UWVS3rdX2oWeARWmhMhogtimOBLvNnXKHEHyZNNCn8kaun+BCw1EDJj8QyQSDLyWQmobd8
Ww45dNPzrwJcYCUQBKzvHwA4pQv9FGsCy0IczFcY/JD/pkttOPWGho8FImUIUsvJcJTn5QwuIEc9
RwniMorIv5CpZ632NTlLUovnmVWB0fvz2IqIp8Nw7boe+rVEucWmnusSlFCboIwqN7hcqxWrTXnv
ro1Xjhs1Jy5H2H5c8fXa4a7X0icWpZyBnlaGU0kRYr8ejkozUdYpnAe97d0UND2C4DXkE1UiMISR
8XBIkBGTXw3gzyvKIrVxaOULAQFhckm3ZFz22hq8M4zDp0QjpReshXqqC3x+Opq5TCdFfflWPpz9
bfNvx4KkB5fmw90oqlOacGUFZeiiiNS0YkPil2qoSkEsLv5ASFYdfrc3WZV/ldit+ligV40nEdqp
mwGOBajQYHb3mYeu/pQ6BqcTpHOleeXoL55MvumRot26RaulWkHIGBkm1S2OHtQC8vaDFKmUUt6q
P9c1B2rq/YbYS9DGJQojGbOqSoMHOAzaPcTkVH8DhyWilixuAuPvfN2bd7to6OH6kHbpNC5WROCY
KeDxmio0dJuWuAZaX69NSnHNbICa6DZvk1sFgdpZK1AuYYOL0BvdWl9q4H6wmBUwuTgEsngJUwlQ
SaYWlMg5sKMAuvnF1i70mSPytmNfqK/E9mlaY0sDYFtEn1r45KD7VkyiiySnoLyIDIdHXnptSIyt
0SfkgVGxMRxQvt0g5HV6phtnMK6udJrNglz4g5JmJ2bXvxwPME92bT1BEcJ8/gLJWFoONKe4uRoi
qxDxAFibxhUMo4zzMnUIdWmjcSuwtJiewgUmOZdfrVKc0DDn/Nn1y4FK9aXHHB1JLw6L2/e9Ast6
4bu8IvL28Hb2poVLEu2MOEuhGDwvDRu00AufzKRqHZxC1dKRIdd7VVH5yghOg802oRfMsCNfgZ0m
FOFJ+S1MYevTQFyoigRS8IL+siHeUlJZFgxlVsG9uuRAuJpXuRtvAyPKpSyvEE26GUn7DCcm5GWV
Yiw4Dyw/YzoMdYU936mZMhMclz28nx8yExwOu5NKJcXmcIZIiXszMXjqA9xYfPoCu3RUuK31+YZ4
Hct9gy5KO7F7oDqp4zE4fG/AW2vdMTdzPCm0+d8HV49ur0L5VBqQmknzNtzQYOAAhUAn/MVSwfQT
dzfBAc89VPjf/R1sG04EaE0IDOanRDAajQZkiOmOk1zbZMl6C0K4yx2scuMXazdQF5phkSF9Y1Bf
iJrfsqFSccK9dndzKB6m1uUCNJW3CySY+6IXlHGg/ysNj7ineBrm270HAi6aXv0vJDRw7YmQBXMK
pm6OvmYrRy+x55HWwEe99wumnVyzGwmtAoFHMjSy9GLu7aSVGqIUkoE1URttPV6EKINc/suAQbVb
F8GHjidFojTsWCjIzaEr7QnzQnntQkliwWcPyHpLtQKPHOa+SxUwq5WujrbGz3xKyfd7wQIyQjur
MgtHHtkSBImeqJPW+c6b86G21ngaCcPt1DRU3gTCRksEWyZFEQO22xdxjHhdpMURanw5tGSa1DsE
kWScCyp0esgKuMS7J8hq+MVI5t9tkdk5BxYsA/jc2D3ZMADvnUR0bqLlvzgAGq2UNzoVJnMnKqgm
wmq0U3AGKJ3oLIG/bjJz6xHHFzlC1+IBOWRwXpMdGBf8DYCxjyF3tIWW4gcJNUvITseMKcYH40dE
SmrQzwe7ji58LwNGA0keGm/XBfZ0cqou4hH9NjGovzdRZMLVKQCu+Qv7fIumEdEFh8J2rPfYDx8p
5yVr5NMHJgZNNsFTiAUblyB7m4aGQLz/6WJgifNmZuSApFlxMViPbjZnYjJ0MIEqdc/lKKYZNZtf
ZtKTegRw+pKnS9v7FIo2EFgr5P2cKO027i6anPUrM5qHfXg9cUXrEQGhLBwZufVVr/YVHj0QidPG
4R+pkOQ4trC3nRxVm3vHrjiJ4ONBHUVJrS4ytblzoGbeSpzEfdPY4tXzBdvqHPaubqVJUG7J6rSt
irXNI+nG5iltSuxnxc/fOFBPzrBqfz6+P9VU9d7t0k4XTPjH7hEgm+rOeKjrkFMPWnxG5kXqT2Rv
ECWZzrKH/SAHRpn1lVVNJarkIFFuX3H3//LeIYZVW/ch/oOf3lr3MiZEiMeb4AS/Ybk1Cr0DQvHT
ZsY/YYSgcSRmWK7KAmXy+nSNAwDfc/xJNprBIhpZ0WadJpbqJ6mXBXogY2dQpwxDTtqOmcluyjLM
YZfMM6SgQafEmHH0ejEtVzacAyLSp8H1x4RtOMWqqqF2V8JMQO0mneYnjL548tYky/k/pTAof6u4
dAsaQubFX1m+Z61iSCcRyjbLQoQYSpMrtuvlO5C7V6XziiiyJFADOJ49wlZwqqU5g4ejHBp5zu53
CohCpYlLa5WF9xnhj7LWvJLYTmMCC24xsjX+8yiRUdJ2/8iBhDTjKLUJZVWDhOHRklE1aag4Bnz1
1TtBh+uAP8g9FLK8/KuNqb0xLdSwNvBRjzo7zJvTeE0zW7JsHFGYVXOgvK2N23ItxxEkm+FBQMWo
SHGKRo/D0HYuSvEQPpfb/aeWJ/mLKT5aKqMQXgr2Ea2UmcAZfZGcEB6Lw5Mz3cw+3fSITguVTJB2
4dhO23MzXIASrBSXyfKDVFvkgADuqHGeAYo1me7wRYtXOj/tdh9KjM5SXWr98ebVn1ktY19M4wvA
Ud2kNdWaO8SjcTyNfAAuOZlOy401d1WU4BjwYlSn3vULpeMjZlQF1HScu5XyBTZJeX7TOMflGPmC
J4wwkD3qwQc1cNp8LilLETQ/gBHzubBchXtJlAhIxwB38J85/inLsD+ff//z9QyFK8a8p+OtF2JW
2xpP7kZPNjXu9/UBo/a4F+jrh2PQ13n1D5xr8PS7P6Jpa4s+eQarxW/mIdAgM/aNGh9p+OGkyuvh
2zO1YleD0kLL+v5suysBaR4J5t1Xmno0+wOgi86Jb51KvAFrCvFjj8nefn0Iicn5SRxf569+O/OF
sBRHGiFtKrLVj2R3TdbzHMd7eo5cHBc5Fq9IqJUtWDeKwUcSCbY81ScioAxGFmnzaqE/6x4n8UZG
HahlJ/GfbpbXfkHu8PNug0Eo2pa3UB4ocQJWN613eFzIVINE6wtcHbEucSFzGXqV52BD1+O3B3M7
Sm37HuMinS8Pe/JojMxfKE6FMoloHRPXr5Jqaz92gWlDK+BV2T3sCZzWK0Nx/fmkaQXDRrPOZBqj
5jHFkQJ/bjGiyXtzMPPebe1R6FpSeqMfggdYvB0JL46KCagq9EjZprOPMVag/kAx5fqmL/u7Euz6
4SgWby9t9vHVl81RU+MgV8tBOaMJfy8Da7xxPUwhp8XVFZDF8V13iKufVPkPo/6XUrR/HbGI7IQ9
+vCalv8GFdQdFQ+Jbl/kxsL125gN+L2PRxeNsd4i+drBSPgnbMFbATNQcoiUqEv8rHURlcWPXVZN
EJ488DaAG9ShAsZt6+dgeohMezfL1WcbZMGNZ2V9oTYRdufASZ/2sNhwEbDNc7MYfp89K/i3abaU
SW4JXJolBFdgVN2JDLxYSOWyRMfq5Jo8Asp4+qY+2I2A4cNpww0Ii+3HNBClC3d4OWc1cBIb/DKV
4C7m8d7LCQFj/x8h1PSR62H4gWYe+R5mlRTYbcOhmMI4CR4FDm45pOrQ+bKMGfBbxR75G965xEMS
IQG8ObVII8cwoKLfx6g9Aay8jtEaNoELxD67YjHbgoFrM+ALEpDvCsXXkelZjPew9MxakGToxuig
uHGVoSNtYbyRcirPX7axcZM30Ohrm2D0hzOedTHmNSYyioLqtCyaDjS92EK622/xYJOZiUJURuFS
EPs5R2C4Rdp7BnJZwq09vCjVL04HO22M6qy7pU0eQYCmrdaSgnWNYs811S8eKrxnTNU251qwoIEZ
JnPftT2Tmd4sLvpc4VDFLWztoWLifU2py7pOoeECF5B+Av8I/i1uivZSzD3nHVfqICnL0FV5cQQ6
jHd4YGnkLRMXalGFGxY3pEchLZrcYBw2LHM+FFroBJoFbRx9n7wWn4zMtlbVvFfmr8CJjM00JmSL
3pBdtuZCCU2y2Zi8Iu3az7B56ReMehJNdik+9Ooq8vWV8oN0z23J70SV2baUcgxzxZJ3UInRkLFB
4KKw3LETmQcsZgRDg8Jy0fcTypOU3s43OUMFvoxsgq8+MwSATaoamppcpbJIY05PEHCZt7UaBmOs
wnWbeNfrXcc2ahoblduvW2U3mT1hdNemSlG7CYdlP2YuyzYJHANjUFm5QttKU+BUKv43UWnqtRtQ
cPxZc10Wf8xhTfggAvm+vBzyVeRwVgLX78VWVhnuGIWIYKO4oroe6GN60ugZ53vLveCz2AzuS0ol
5I4Ege17OY+JSBMrfpIz+SgHuGrarFZ28nY6Rmni+xhalWdmPCQkdefzMVdpW69xST0i1kYxaExD
mge9kDiPF0HRFi8NM4G9vuSh6uzUq5Ivvq5KqZhplTUqYwFxA/AK1o+m9HnjWXI45YCsWFE/EyRx
XkajnWKrRCr5wpStXnFibO6oZ0fZWhdrKWMgo5fhrJKW7hUzKGSeDXrT1sZ5qniex1c/WmETrVXL
a7/4quFeXgHg4fY7clCt/xjpcObW26OpIRKWHV9bC1eSTukaFhRrBmNSxrnFyU2D/+SHrr2gr31V
ntXRNdvAg43QUTmgkXMWAJ6RsKSA2DfRJydGqICN6eDKdevxTZavCWZ/ElOPB+nlaU2G1qfApAxp
Y7L8Sd9XjeM8WCEFuzLuYvFDAW0uqGof64j4jsqokrP47YI+Uv2nI0+QqvbGzkPcqWMO0uQeNedo
ygewFNLLOrNpNkM/52mxC+c0iCwWdYIK1LUfK/e0RFkan60gCuHGjc76CQsmsQ4SLPCFcsw4rE0/
OTx1tMQhCaZOBR4/y9SuS+9zVwuap9cGx207KQFz7DtUkf+/WzQq7xPPW41bYdjRTQfEUbImE1Bz
PsMp0osabY4hpHO8QhfP9kJB74BKLVv+VzRUrhjB7JPIOoK09xkUTji43esDAsal3Jka15pblNcB
6tE7JwrdjQb6STGOU8fXu8yQYcI73UPHpg06bigk4HaIyYFBNwqD5rkzZE9b5LuxvxwT9p14OHYX
hdIcPWCgpQu/UXzntGNwrB60ehPkSDR5KwES2sV0bgK07vVw6n6EsGGLZiBTvn/zdjsj2Y5tiM9+
omFHqq2ASIXOZJXexRlNdyTvAj7+MXMAYTMHPbEUgJNeDroXIYsIylcbJSMIUekH56ieWxpULSsH
NCrtDkO2QfEqE273QzY8beLNMz/jm4GLrGQKfyoBAX2XqsQ/fGg/7PC8joDzS2QVVJTgZF0lKjGS
wYwSTurIJBst3y3BmyuwQMtac7Egdq1WgEfg2fwnMTFZ5sLyUeRLcbTO76AgyHbsZEhv2WbO+cG6
HFxXIlD+sq9L0DtodTtcGtw9JhDHa+FPNhOMDexfY9Zrzn+BsC8+D4/x6tkbMPsKKvydUCUMY8fd
Li/d3RD8NIi95ERfjgWEP9HZDozwbivoG5vuf+iE7tSHVwmoJy9kDYkkUzj7kP2BV7Q6y/c/T9Ts
3o6PthGvZMGEBHYF7LRh/KqCZu73GQOuS+ku+0GT+cNQ+Ga3rrZ9Kb/Li59nZ0++m3k/skcEl0NF
LmZUbMVqgByuzNMT8PsZxFBJhC20J8mhVskSz1k2byuBQW9KP1iRizp/2OX8vNNMwpQgUBH420wS
RaBea5VJEcUC8lEftCyx1z/rPCUYs8di7b2r1GJM4yRjKLavqFjLNZeJ/7xL/bxVEW+MJBvjC1t1
jww5l3IkaLqrZPR+jWT8aiXkyL7K58cPpeNRdhfSqUZS0oMl0RQPltzB3yYakK58x7srFizimvO3
Kl1nJBIlDT3nxdmNv5lmD7z2PCUOBc9jnUHWxwvMEYUiN3XOwqF/9jAVHg5uxz+uhUMzSZk3JUZc
gI312Z5iR+tTUDcd8/sBIMsR0fd9fdF6KpWk3zrqYyyl3tnEiZVKJOeqfIkAt0HcDIPZWE3ooGIV
I6+OTkEqgThKhER6IMbD4LbkJhUXNloGzsjI7yySPdeqwlxRLjIPtYFwxo9D/w5TavVaxj22jc0V
k/nIwR1ViW286JEy+ew/9WqtrQED3OGw9ijC5HWULzTJbdGIUBLOTWI6XFKK5CC9lkv5c05+dr95
I1qOfW0DMj0R10wDtHaIswR3alpZUGiOOd5xPVlH4ZMQ7w+Hu7x7KjJmFbNRDovCi8rnHlRXe3K3
idPmxIgWWMbNRNfmUzaVbVLwxNONqt/UoPy2pc1Sp0NlGQu+nds86OnRhy1a+o0MS7o7B3Mzuus3
B+NT6xbQ6XlOiU4nEWu748WjUabnJ+t7IAKaZUmEpADYByBm4flxhuaZ+0vIr+VThFqRGRt2eNB1
l7LyJgziNRSOXqb5iO7LX5X+oyzKK8uk7saAGLIt9sIa7q8VG6q/AD+MguUC0WOXyV3By30TYqYe
IJ+LDJE8yA1lmyEz7gPSfQs1MaSidT0JH5joZ2IAfgw9GaS1JZuZbxU9b1kH+PoEkh1h7U7Q9tzO
1wVNuW1xUwCBbR0dMmqJ36IyumggTHI+ex67dBZcT+JuboR0E/ywGBVWSaiJFN9GrDprtO1gxsvM
TYmFIV/UJgdRKc3ouOrPsBiS+EbsALZL/XlKnbEhqTxoaY1WHRWSKLGHRqN3Q3yHBPqiDD7ymnVH
UIwX0s8OcE3xb8WPbdS87a4A3agsAgKgiXwQcBLl1ajhlitcVReCrh5JcVMUQ2EgTJ3iQ7SqFWy+
XtDqRdMwAhsPiy9uGYh4CnWM6XwkvmHi1mBsLPirCe45ZVW7+4NW9E1lIviS92Obf92o3mmQyHl2
3o4XfRicqm33TpxUFRzaG9TnF4H/swhxZ7da+4X1j+nRUCJuAJMcECmeFtBfsmdl1Tz/LCJEGPF4
d88DWyZsGZFGYu1xiAHvXSzRCwl07qonrlqg2tWhUSRDcOxh60yEa9COKBCDSW6nRviFTgpNzHwH
Ub4PfQO8h8WYutBsQSnaIFLRc6SLnxUtu876ESXfkwrUzsxyMeO2xYJy8kdMLHdNKHnFqFKlETcq
K6hT0PZWTFxa/v4gj7tjhccxb4skr1H95jmIBPCzTXYdjmEplVKdEchJPvUh+WYev79eYRqOXUBs
t/gTEC0xa1gs1I6Kyg6aE+QmKRzYeJjzYLeTyK9GEaLnmTJD4H/5FUtA26IzSLx7AtlJfdrNZven
KfBR9XZU0dYy5uiiPE5ieFq+NynEXBTLOAmR8whVFZBxMFPOyeq15SQwHmsb4FTYTyWsC4X+KH6J
FWRE7gZr1EjgAfkxKh/CKfetbo3PkCC1ae3ZpwlZaGi0SW7xHEkpD70nQgPSuJQCXhKbrDW4XW0L
q50X3BNWGxnkNyzHyhvtCANVCAbjkrlwchAbZHZflEojw5FPer9A6dVoOrMGOvxqfHk/xuVQmGkv
d9uuvz8CtMgXkOWFrAtPX9RXL8Q08FAhtgUJ557+RmDXojtMqvUMH1Tt1TXNGCY6d03AewcW6AUO
XtA5sk0wy3Oa72Zziyx+flYiOcPJXD7YvPE7PY1p982CUrVuIfcDS2H9pjSj6TFVi7qDZysrl7F2
NCkfX/B2hGkVGW9GImxl00Ji5gmYsGNHGYK4asKHEGrRcY74j8OQzO/jUIeI8oyDq2zd3mYbg0Ab
34vWXS5TaRUZpPJl1YWksffJb7SAbixBq1W7YoEOrA8KNU/cWE9Gi82XBfxw8DetZPX+HnmR1+3a
CRqEg2zl6nkMnfEe+xNU32WvG5yg4c98djoRlGkONOtQmycP49DLrv/HTFiK/fly9zfi2bMD7NMJ
Sh9njew0bP0jR9PtFtX/7S4gXgnRDpom0quMo9XKbk6H841g4x/fjIvp0mbR845mQo9zEemJJcpc
BF7wyJ1E04MiGdt3O+wWYH6b9JnnwquJofIoW8Xgv4aLFXsEaFIPrpvhEqRfkriUKv+L+LqZBbwq
J2w9H7u7bMRIQfowEDalhitJs5noZVRADB9gars0VTLXZ80POAI0FJSmO2wtOtMFFxRhibm0o7o+
NgQQQrhmvfy5TD+mznzPccIECIQTdDMpS6ctmL8AKZtqJpoagtVdSgtyxjCvQ/zlnDHUh0vDBX+d
OmDZ43oF5TknRVmygCSG5GcGGIiP/Uhdl1nQjGxeW1ix0cvMqErjaiZqmVyr5wc135iEdJ/Ppv3/
UToqqAjGg7QV7JjkvbtqsPUU55ygZw6A2QSG8OLnYKfpdyCKwFsUuBGmm+N+UymtTqhCTGMiLUgL
QsF3GeINQx5htIsbdJgsksqPwqgB0aEeaKIQSMaD57gF5VMWDANdG6zZeZ88ws4jiiVhO1buRdYH
omRqF6qfjVcR0WzC/i8Dmk62NEFuq+JY2Bph1+tYSqeBZdnovIQizLwDp3nRW2kArY4SnbvvjgHG
N9xsPFdDlzMWmDNq5ij567ISCxDemi7kq4vsZO8zwOmwDsdHMQm0A9CdijtLXe8KzTiOMNj/PHd5
Zv7z1zOm/YLG0L/c3hgEkpnyEqQBzBVhxptEy5BrjHN+vwqXfqESLaBRfaij3jultm0Dih+ShGex
BGYgw8nmAe2KQrGGqhifMLn0hRt2umFTcZTflcuv2yM8mGbb4QZ/re+jpTWIO34MaVqb7JNC7Xdk
1V4KPZ+oMqiHRVmSqnrtHQH2ebaA07acXh+GVTzg/KdNOPQ2Cn+W7YKzm72yhbqb0uvdSkSZ6m+c
xF5yLYEthtc951NdeA5Cr+VyhSW5Tf2MQCwbg14ITiWhV2LLrgp5d82eW1XsSquOZBCikxxUgzp9
WjGMjO7o5tEZrcZiOckCzLo3a7LbE1/q9Y4eJ1cSoZF9fBeHJ+Mrhb8swEe363lgnZusXj3qDkeK
7N7+QJU3k6powx4YB+FGgDIkZAZiGan/FDw8li3sM1OrivXrc32/vVEnReksUADyiHC9Sfcpou6y
yeszr39K+Q0NgFmfnn6YaMaKGDk/KC4Dp6hzpu2eazyTIur0pDIT+o0cMLjhLqo6EwX4AHbrOR2n
w3TLW/I9Ax3SsuuMrBOu0AAZ0g27zH1jXSpqNrjIdQtYB4P1ZLZ1OLePV1/EssBdrRrCegUzNLhp
ZeVbEdvzBzqGusnDxAspBaoZiIevsDZiWGfKGj2PnHSMA7+D3I0REddnWWCvEZgoPrmUVqKAx1mU
J4wipXZHUaOPIZ6xULmsdCmrfmLkk5m9BsPGaLbVj4Lkg5qY7dPTYaLDqZwF70nu7Sjp9M/byemS
Zs0LMTa1nsljKYpqZC3auxdxq6zM5tJK7+yL2OiqOxBw8xj711VwXGIY0pIXAqZGJuP4r4zs9SnN
JHgq3xF6I9ok+H8PVLE/wKQ/SQVqtKQaz3Gz3cGz6aDLkcHIppTJPa939VyNz2zVjC8ITCPD+2D+
+mMgCaSSXI5So8XFgQFQwkZ5WRPhI1g+zRwVmnHbDyYlNQFilTurJUtxfZIW2T6yisvt3NbpWv/W
4hKXeWcBcXCBgOE0FbwJkOQWLKQZ4HY46jhB6fkp9LlqunZBuL16jGGQJjUTxTkiL0kGExoJ2J20
mu3/VJQZuggtbFFNZqZF+7b4s/UEGboq34QQ64aEClwzpV583GOCG7bvCvYe1TMjs8EoNGNBm3Xv
jHGKWKRqsJNwbJ7m1dg1cQc4onRmdRvC2RpnQ63Anxt6pj4gblDneTueoQQamAozA2vDKaPam06P
LV6SDZKNTreXAST0jCXYM/lRCa90hkpZjnAH1aedfR0IxjqZds6pB7w5OA6UcIaFVR9aC2Ezg2DF
699rjtzdC6c1q4Fr+17tViCzT/A0zlHZlRrzuvPmecLVxkVX8wkBBoQpuA4uTIwxYOkLnHN1+VOv
rgHmMb1ZfQ4NxVDFQUCMlBO5EMYElk4mViXZyGqJvL9cIHQdZ3Kh7qyDuKnpVNy4DEO7TrldFj+z
VNSYC7dFvGbRr+FCGPKwJQjZHcDTtLWR2SdfhhxqhPOfT5TyIS+uoakie5wdD/1HCK+vGqwl0DVD
eczytwqIC82GD0KX3Zkrvo5zwMw1evJPyCaBWejDEvvwlHNzRRCR4CPCTwRAIHKBi1DDGi5SAUjD
my4TkjiY+ljCy/BmJJ7Ul16DkTlqM4iVutsKuzXgwMMd96uFAWVOIl5p2pSvA4xNKZPZgaQ/UhCc
zakuuu6pnn/BaySyZ+VCVTZ2oldQUKIOHlgK5Mo+DHTQpHjWmoJ0QmBqFeMJho9F2fBt+kMAIany
kDgbemeINNhlorer7KiaNS2yQ/FrBxoG4n0hlmNUVYv8ZfvcfACbCj2ZqpGYuUp7P8aw+I3mnxz1
UG7fcCJGqcnUTg9e2D4MINOE0bo8NE61eIBHrwgzp4NpeI0qpKfi2Vwt/3kIqoRJdzX4/zQZvyyQ
rZ2JUNe2jesHGCvSi7a0IIY6NH2iM8YsoZ0jqJCowik1jylQDj10DqnkF5O0WadR44UTm7tkLEnq
d+Ta7T6uVyp1/+pEM4rz/79Sn9qxl9WtmAyWwn1IxMq6nhn2bUGq1bMk3IRd+rfUrYnpq/GhLAIe
HUwFlt4iwxLrDf1FqkrbDEQwHiC+6OKtJJy1V33+/RNarUrsRB2Xdbl4xDVJWNTuBoR0AJtNZGtX
1zjpQpPBsognOpVNuZqZ9faXt7I3o/3ztFX/xEAiQ81PYcmp9MAXLGEsrE1L50RwFTuAFMWX+n1p
utMkLaGoeoLupEQ5iWY/35bi55mQz4Pu4wF9YGXDPoXQ8Mf9uM8C8V5NK7mGVe17N33WwXvjl7BJ
KJt7JtWHORuM2QFQLUEiQ2FfFXPYd0t/VWHyobHVja7VrsWXwhUYXoTDiKhNo3zw+8bMrVhlWesu
tWhXn5sYR0kUP2vQMAPO4z7lKuxklxr9EGEAiIqWz2yETk0Pakp4IsV9yUGOIX8ttRXyzbr9Hb2t
5UaupRoD9iL32yHY1IKqDEHh2UtJPSoJI1Z+S7aA4jCwsn9KSmNDpPcW/RzY1hfP5WbtWcsjW63a
EPSgE6BfG/1F/3sW5/mcLm1rEF0H/HMSk11fbAjuSMEV+XE+SqlkhIOpfc7C6gvLetmPpPRn2E4A
7a5virHNYSVd6Fy7A0XtkK9AYZGB9Q3DVYhLDp0BbFjFE7yIuzOv5zsjm+X/iBN1JMnQixQLc81P
Wrtb/s/yVXHPocwJ5bCg1BIb+ZMIvMUF7N7c6oFgz0r6BLzKF2AuGy0MDWn41qCSt3QlrTZkAe7i
C7jGH44rUxnRdOTalbYSJCz3yyCIwqWTCrN4uSJ2fnua5x2mSJcOanRIyb3wTfthYxS/mPL1rgnp
wUc7nnUAPo4O2wuUpHGtxTVx/zP0NtrK4JfeDYydpgxEdVmTF5ai+krXkzYLiGF4X9qU771QAvuu
GuOj6QRK7dYKc9XygFT41NMR6azk3n77p8EMQ9tQyIsSsJxBykpguiTcn4Q79BToRG1TFVQ6iSKF
RQ2bxnG8GoZwpQYzg+rgz2W/uMZUnTf8wCTJu4PQ6WHJBc2JQvwHzDDoyUwIk3xrxXbaQbe+FrEz
IUYgoX8wB6jTCqOvdzaMwc6/GuyS1aBj9CAXz6g+eh+3MmkCFm9DWKf1bL1ZrCsTrfMWn/duRI9L
bmAy9ui6P9KAf4u1vBUzu2NPFwAEOA2JbbNhu0OQk307K04cCLChOzL+kLkjw0hdT/O+xsVeuQcP
sQ7UvUnCSK0ANx8B4XbhKoPOy0OxMaPAjGDIXk28AqB8e3cW06WGkkgopkO2/BzwUO07qTJ7JsTX
71lSEeg+O2cQ0KDMOFBbw4GIik0PU+XHQ49fmdfmkUnsYl10KGEXi6B5osM3v5GphSl/c+f+6/Lg
Vz0wHrcdOlyQcVMPGgRIXqTepTpMzjxZlzW/YDpyJRtNLQT4d4htglcK5zWYL+LL6NbNMG7h00v1
G0nUMKfLFXtoToWQTazkYsBKJhhu7T89aWQmfFsi+lIOX6a3AGX4y4m7TgRly6ynPvvlOQM6rOok
USVoEv95eVuhDqjkqdt6ZWrZIGqrLPriK9r6IoIjflEiUKOHdei0MSzEDksDIAl70e2c4AHCbHMB
so3XbGPE+GC3l85O+zXHB+QPBEBQOaeMq1m0Jq0NRXYN05DX2WtaEe5h1eKAzF7C2RlGH6z/+3vS
wWhWGN92rzmAVf9Mq5vQNELWpfi17gE+306tSPSgsXI3RS5B4GsuGij/Ii8ycU1QkZEN5wEFWWi0
EC+MfsUvcR3/4UDryQXIG988W5xsAsqmvuvnVLn8l2VJhfF2BfBEnfbavOko0jgVGG+Et4PX5w7l
H3+CbPfe22nREXw7LKsrO5Xg3APIphvNIfg4IXXpkxjhHqbAvqqZZJpVCcZAWNYmSIP1xc/IKMjU
GaUQYNz/K/oimgwTSr0QDaaPoJTUQmM1XRX7fovV3+VreVuHLzgkOge8ZTbr7ouswbSt3C+ExVi3
n2uhjJJz0t3OaUK6wO1wR3DldKvREocgc3pQ9UpxLFOHsfuDWzTch/Cg44/0Eee67H55mCpk49yp
N/g2I/gabq5lVh96Y6eNnjElFi5MQcU64LrjjAJmXQLTILtjIZqnrGjgb/+doHtkMGgL+UfmbokC
oApjDY6k+76wwdEwFnmezSeHEA41rSg6lfJki1QyYhPWAYl6DGvkim2lQMTaeAtLkrZRUf4pvRb8
eRsRAdSfKUy9HWKZvoy4ufOQ/tJjFSqKS8u0jiwF5DoGUXmvpWQCNxcsKP7ASYgFJANFn3y+QAY8
4NN8hTakfm3jbxJnQ/Ao4SC8UYjQPIHt5qcBsNrSEJ9Cs8hycIMqi9p+mu96qBexRUBCsgEGtCNz
H59JbgchUq0Cp7gRVEpl3NViooTzN/zh59rZ0xUitEnn0osnCbkpLtL5aSl9ibmUAnGKzeC8P3ip
HwHnaI62lnKZPYrxrwgIu9J4FUc/b1qKzfAMlM9q0ERcYpB0hhUujWUafNdwq9RtTpa1TeFR2a4l
QWtH7SBngKfF5mR+QvMkyBq4Y9UXqCb1XuLmUuK0jyGxUhOi1smH0VADEMJ1170ut63TjR8EbYDR
xOfjLbDZs8C7jCbEs4r+WHejAvYkYVmtW3us0yQ+unBYEDznSdariHlvAoFsApLQG5sRp5uyOWY9
cb+yzoYgKA0nZBhY51HFggElstaIDt3+bj2QJE20Tvlgo6h7LQRUpq5WH9OmsutHSe0y8DkffbH9
uoH3I6k4rOyPnysajzfc9As1ROMbVFFBxy47igwyTsfFfodCLCMuzG3hFaA+aGcu3xV7lIM54EH5
P4br9GMKeV0l0Gl8Hz/J61og9bSGNnglhppjs3euKR83pwvXK+40kTfduYsmlkr51M3Zjn+DsMpV
wPMjrNjG9jShZWXbDlLzUM3kLp0VN1vdxfzExUkvx3H6aeuy99ELaF9kBxkF2slD/o+5ppO3okru
DKZyOMCoU5TFCeV5B3S449f4yBexge6WEGlvIcfQGqQGPIvEkUPFA4Q7fEQP6kn+3BoaRgnp4K4G
xo9Dstrh1sOLqqbpRMUz8azyxYlrWARV3/anckwnLAzQcToqV3nOECRelFBxQTAr8BwKyBHllMU4
SArH1nmbAJvyUsBBmQ9Y1A7U17aPSTGAgLXu3Poprqy50TwZFbys+ylMjiKvOBLLGOlSR7xcCtim
sxfzyrB0r4PJKIeBgKgoDGganA+7Ws1vEj7s4sQw7R7JI/niloSVRX6E4mMY1ndbU764gnJq4Uaf
jGBEo0LmO8dEN8nPYtSTwMXAx2z2lu70r5cqqX8e8f0wYjVg1qE2QFW58Bw6xKr3SfjKIArst6j5
2MbTsMUPaV/5ZFWXRlA1N1vkjbqJKhQMTOZ/7WjXS/7BJltUgUQTCx9bI4cIdT5cYl2vXuUouYz2
bZvsWpAFa52bOOwFtKMGuWZ6z/Z9u93xd/xSpv+JuSQE8WvebO7//tbzo8qn/RoiteAEyyLa/lpJ
9uwcvnoq05OXwcC9p0FiO5yxhfhEhaB2RQFuNTWNz21vpeymQD6Gc8i8whzF8vZlrtZzp+cPQ75J
nuxb8NvrHHiRzWaoQwyx9NzZCb8Sfazdjh5R7hX1+edsI7ldlgAzetKqeWaYtcJafJD4lnWH2Wea
coBEVXH4TLpXAkMdLAFsAzLQrhZ3SVx96I8lo1oOuliB86nFd5T/q/06YxqPyaFPH8/YQONrlERJ
VSKp2LWeXp3k583pC7nMNMUqib37E0frR4rC2inPF+cJqOgPf85PYVeTUAr1Q3qju9bKKOvGzcGw
qZbpqKXk+fC7G7NwRRPT49grPEd7esB72nSY8dyKK1Ynsz+hobdHSfSjnVS9RfYhAbtFctE4VFAZ
0ntN6pOYTVh2PGF/SG+MeaFDGg3f/TtnTo3WUv0Reko6JlnutkDiFHaZ3r6GJcM8IEdrDC1U1/oj
0debrk+N7T0Rl1i7JQKIY6rJzWIdSVbfl95KDcGOE5MhWQPJXNWDRGgZoVdzvvfp4THSS2+hS6M5
Hw7JDvrCyGt13aoZg22ngLlMmW2A/6BwvLAiovrWwDlqtt1D/o7PwYPw7dZqFuWtfVeD96DW+W/Q
qNX9kWt5wlzZvJBKq9DZLFwwWzudwK/VPGJjneZMSFojDsTKHRld/WLoZKtSrDcOM61+4E3gVrAd
KY/UP34hsSjunhUQCeRWw52cBNqdsE/Pc7qy1q9fjw2bij8gqunC2tGugj4K+OnQ0qnno8DT/I6I
CEANUV12fBUS4YLzqGANaeCAdYK6r4mJmchQZc8T0nTNrJk6kMV0wbhgwoNN19y8CXukBS61nmYo
BBluRgJ0MUa/s1HIuSHEY8US0o99TLnjiZgT9O8Bc+zWvYwolGZpHl6zQSfDINRn/NkH1FCCC8Px
6mpWc2rkCNCeCg1oTX4f2v/2J0fHqLDi4gZ0EGedvmrlZU4eZQhvaFj0A4WSYQX1sIHNkRNSQ/FV
eGcGC+DmFUd9PN237gIQgr1FRqUAuYoO9ZTwVF2ut0my3SFbOR/67fOLmyJKudhX6VBm5UC8dOWk
tBbytg8v8j1j61LNOjFhoKPgN+xsLzL7AbCez8qUG3N/EBthTKVd/NA6B0nFCQIDp+gQ7Z98RJal
kIWtI+mEbbbLrrVFNv9MCJwP0Jokoo3VcTxdhECGm8tYcrn0Tr+4Bov8wjS4CF1cEocsaI9IXQrI
DWw0pgg0IcbuAEtOp4+NdGgvyOmRX5ropsMWzqL0EQJ9LNvFPuQXdFMGbFsCVEkGLNTlhvvMimd3
SckCkNrRsqFrLxgQxDE94qWTqQMETLkeq6C0mmYX5XjupEc0xwgEldeABO5F4qclS3rNRNMTu3QT
hDMA6OWcgqinOUipOxLRgRNr3JYmhv8dBHcDaMUOs1R34XjGtsYhq4moUdnwoXgRjFcYq5wI07uD
jdmz+v3DGWBph380bQ5Z+kAYyHd4nzT3R6yhC0W/EcYtXnIFO+usqeaYvIWfAJVllEwoHhAdhXcm
16ygK7J3lwIscri8wswq5A3dG692p6j/ZzSl2JK/iEmcuAGwmSTHuU6XsgrSdm79sg6p42IJdZ2H
T98EqXvpNWrrCPWCzYtWhPXW84P2BfjCIHvCTIiKStgcxvepDe0AaCxEZmRvZH8+uOBl7bItXlpF
Qd76UfUsuZGO+dKJJlWE9v/hzwqQeT7F//qClP49fC8iuaTxn0PRU2ZuzdddpZ4RT30OkpMfq4zn
k0X9cydAQ3cppcoWpDPWseJqOzlKrW822QM45cw5xrIXXr9kxZdVG3MfPL4vYU1z5cY5nbZ1Vi0y
en/oEN5krnuD2lc2f3T4OuBTJzR5Xln6KZJi3E8SE5QZqXerDP9//Y5s6TTfBHa3PWB061qFTw2G
uTV4yWcfwTA0+49P6bnyvnqnJZTD0Ti9gcZ3gI1e6JejfuZAC4t8i8ZJOiomDlyhuRSxORJE++rN
qhGLP+tQMjmkiUCcLtlz6GfCQKIWCJTAqOFqCVbV68jzKCoeHQ3lbo8PmZNtPVqcnRQv5Dv4Y1Fb
sbexmo2WzVW/XABSIXR3/gzVbhuxHeixuN+xql5Vy9pwnk8oXZLNGqkRvesV/LgPnmAiakqe1zhE
p00bzaibDAZoM6fOXPlIO++67CF28JDxYmPeLAuOvNLYLyj4KdMKUOidjYSBsUrpdjGE6I7vJDxX
RYzqfqa3GwkYxKEmb/M2YUAGn3g/058Dpjj73EEeMZ07HMsPdXMuCvePzGDWbB49zkIwrJbZdyvK
G+izsZezeR5Rf89jZpP1iPlCJ3MtflydLRTtSbRivrRfbI/m06kNBR4UUIAMRtSeDn7yrW91IuxP
tUOkozqUwuqjLj2Xe5tXUdWbxGMmZoQ8/dxnCQ0C2aDQA3Ed/bnmd/vQ0NLuTfKEx+5tZOLq5xe1
ODWij++1G10QSoCJeRNyxZLRt2L6Du8qH75QJlRT2IPdCjJHqH8Lk5W+Zouca42Fqg+6sl8Ubyg0
/fVuYCZI3iai253FBTSgg393y3uSuWZBb6tVTlszDl98hNpBkGNAyqMuNtcSy5jgHFZPwf3iyKt7
2PYE93DHgUTMtSF8n8icY0XRlTN80PTlGBECWyj/8wxQQhQb212Bnkv4F9LF+FMDESCp+7FJEIlV
l9ajK7irOheitxcFSJl7gAEDhqyHSMD56SN7uFyoK/9BHxWFJO9qwkPelxItugnurM/9DYhysnL2
rTD01cXn3mFTzlk9mjqQT1lSe/kXTnydQdLwO9n8xpO6PmHMrLo8+Osft9YeHLcsX+tyOFXl7gy2
cFIg++kb+VCxkFIDFONP6mTaqhCXp0IEpv/V5CUGt7NdJZkcPXyuh54HQWZHexggZtt2WzdYzm2J
l5OoSHH8ChQdptz9xdO8A+K8YdrP9ncJnCkgJj1N6MYVHiw/rjDTmpQuqe6nvTNqHkwG+Dnfqpl9
oTbQS2K+LAY9BTg4GaJlP1gLXPK6yEpRH6I/n4MlTn3kiXX2/xCeABxsY21iB4xkCKrgq0Z2CAVP
xKcwEChSCNmr9INUWULusLXG572eZzRKErWLlZbwbs3MIRtHG8TimECBphfDzjGTKEevZkc4o9MB
ii09Dh9L/4ACMSXyd2Dc/C65by82jFdrnWNE+egJDQpIldJ+/pMuZuooeLuaX3+QisOoUXLgczT4
Om5VyRbxM8wQbcrGJ7w8PpuCX4y37Gu8Qr5BVp5jsDKMT6W5cGnGm6M1jbPeJqkxIerxjqMkKid6
YTV8lLrWVwXLAPgAK4w456ZExoECHK2U/8rUzqDsI4J9lnK2JUWQzVDu+aIKHnSCITnF8oop8ZUc
vUhNezeV04ub9J2RZNx0iZR5uLBn5pFVrW/SJ4F0I7tSOtWt3dd09SihS/gqaCeF0RqtYilzKGll
huPyInx82t3YZ6R3dVJLrr5QfkOCwpIK2C5x5BRezi+sMwKr27xjVufje1L9bTMMsptZz2XqL7i7
Ebr6LyYYIDVZqfyIhgeNW/piObkkByPfLICd3jRqd00Q5kUDC2J6C4iXhqVZShKMqHsxPBqfg6KL
QcgnoQK73H6XOJqi+kgLQt6h570MyYkp14RzkDjUdBQ/EQH0k1DvZKcc1w2MGFkqQtBfT7MUCFnM
OP3xvRmO/tZO2aGZwQaHrW3S50opxOLjGiVA4yOZoEsvCX4u2i9KuSMb9NPDPp+ZFaGXhAzCNVfm
Cn9qpasGm6JdbN9tJ5npL5O5mXt1UQoRAivbKcusoq+X5K3iavl2Bii9Qr1FWG9POsAuaRLT3xJs
oQjKeZBbHV2me0ZbeiV9aXTfH8iEcB/Jgj2RcWuApb6Q6Vyc/JcIqTWmpWlrrsBX8z8/nU4Hs0wi
VHPDmZnser+1/LEpD1U0UqEyi5p6c/e/WTq2GVpJ3L5gbBAJriPDH8aaZi4GNTQs8dWanMT1OM3J
7i5t4OYcNC0jJIv63LXsz+I2fCQ+KhrWNkifaf20OdkBAR1sQiU2uijN6knlJIkh+8s0jA57BnJ8
Uol77e33JnYJDsgbinvLPoe/WvUu+q6kaAUG/rgBqlFCaTrAltc7eHOwl0HPoNz+9XNMM+6vBd6d
ZLN6vFI9il/kF/CsFni8hzlGQxupAJheNuB9QlAhsTm5nlOQ0i4K9Ypzerp9s/XFZFzrjoNZ0512
Q6raJaNSoh7722c5Z+MvcgxPaDnml+7VYHxD5vrmi3+2I3v+bVI1R+JQS+pYn+iuUoZsiZsZjzwH
z22jiGfELM1piYOiIR+MbQpUQmW6sfV3ie3oyB2Wais2NUf02xrNzmi1eYOP7DfLWdYZQqrasTQ8
fVl5BqsGZqwHHSDm4qcdP0Ami/DryqdjpclOjHXrV89qDOW0xff73cbJONgs6sfQkN4iXbUKFemz
acZQ4gU5316DaXKYKWQ1Kilvd6uFJFVLN7qSCauELbiI5VrLGFdfLxadHGmGTpH+5wgr9mRN0pwn
ZiUbmHBwTcic7hoPWTlssEVM52/6glkvaER/U1xgewBv2cXVJwz94/ZZqnPpkjFcmbt/g20XOJft
87bF8Kumr+ilysZOv8NjpPT2OO2TUZ8HUdg0z/t1sgPA/QuCIz21JzzjvfeJ+rA59msu2ToqSSm7
bSR2HE8sEgWc+RJz1P877k2Li9D524tzh7h9QBx3FMtWjKX6CbkRYEEeThWkppBOZhWYcPAIlaGf
7550uRPgQpZzbUqFHIpcSTf/+IyxIKEVeYnaUhyHhjycXCb7mj74fBw2PR5XhwOPii61rUXKR/G9
mAXJq/6opnVss+ze3l/XW5jKcTJwDWncXB9ZpuDl7fhbRYj+ZnCCAucEgK28iY/6HFrAK/hJDE5g
JJaa1YD919+9GFRfTDVLmoT8P5eNvMZ1lLUTAhvGzTGSPCrvyeudB3SjN2V+steRK3OSIQvxmHCO
L/z7uvT2ZJHaGgej7VtQjM4SWUnKtV6G0vDnujfpfBI7QfGEKxQEqMqS9goPPeTNhrldCUeK2HVg
Rg5xYUTu9UY2H/TWU+q4V39cRiZRvDHmJw2AoBeRZ+vUO616ITFc3iojvfrnuX505tLQ8cqh/qlp
kL0yHbqrh5VpHNOGjT5eNdgjCA7RPmCsuvDj6ghqNkRMo/Zmqasp7GfmJIPA5N7RkMG+euzBIxzJ
neUhNYVecb4GtlkyJ6Gh7iYpNgQ3G5q2UvBnqXfizg9Mjc6afxK1+BkKo28HByI0QaX5Tf5PkBkr
+lUsKTZTzDpvnOvQsOn4GozIpoe2Gz8BzyqZ5c0OeGqBfevXn71eh62ryYgl33BRwsy5F/UWP0cf
nFdOJ2JLx55QJQkg2BScFgY9xhJlySDzBvkr3lz8reJgiPOJPmRLnSh6hMGxaIGQIxQLAk8cXcum
whx3rGZfWxCtXpYQwGqkNdhw6BAJM4KQHCtQSiDRPkQb20D9wueHZ66VqdXD8CeYy79vTv9d3Xaq
s4BVrtsFqMhpUL7nlvSbwZQ6PrhSIUjdG+dZGfvkvOZcUjdKcTF7O3kZ7JterxSISqxr8sGNfXlW
YkMqebPiWzXO0GjFtMH0lo8dO97X5flAsPoWo07/LNscxkWyoI9fTZIVQUC+76n9GIKC+M2m61CE
/RFipFnCgy5YdLIz5C0D9HlCuNqTapkq77LOiuojN68AUD6qevPwycExd0w8tLpeKZCnsVOb8yCu
SLWlu599wXxSpIZ6BnkQeuA7fTLEvLpMJAa6Xs3tZqOR/dzboVLG+z7LdKJUFAD2NDLHBvH1jos6
CyZN+dzft9oDkeHE/Jvuej1LgunoZlZ9TVq5TLOAGyYXjVtEobr0LL642gES9n3Jdu1+Wpd4nPkW
QIIs4uUR//2Psl9blv+C9jo0y/FAxtl14Lg+6wEPHADynQOZ6lyQMk21nqq8sM/Z1e5mDl8+j7cg
Lm8Dzt/ATCD9gqqhPHO2YJC48wOw8c8XEpWVaGtn3iOeDknyIP9CMPWWQJOBtcuvLi/+Si2l2moX
ZUM1eEHTgg+YnHd9lWr02adzNeOYl0SfPD91X/r8RKTajkwBrtQJRDzo79942WBcsjf5NQPEInjw
tBLWfeW3YC9M7BJrqQ/aXvydtEfR0nJPmFw+1I+BScGQ7haQaSxOe1opzgLen/i+7gJSa7jgHqai
HazvkjLk10zIDIQlRZl2DB5JvSxFYWAnmgqMPjPKtBpfoy2H3oM6pVg/e+ZYkHkGDSD4ed4ABNjy
xWYkim+HfSitXxLKkI/OUGS8ZCw8h1BaW6dlkuAe6Aczpq71xJO3hyWSh7utzvE0kdLVsy2AHwSo
zliY0AiGt9EH+MMmTiDB4yK7pJPm7+sd79IlTy8dJgCm9btFtSCoEdzmv0fRyFGKTh5F5Gyg6QTz
1xjBv5i8PMy2iAC+aVQ1B5NAXH2wKQK3Heacabc+c2LxDlV70Q9yETr0oZUYosH2kZZ9SFHutYvY
53D7ZCBn19BTN+zoOQsObpwMjMlNKFlgRT6dJSdtkBN1euQL3/x5v3U0TzSb4wy14bVNd5i9W/oh
8E1eua2zuKhLVdRrYoEjclwf6ZeHsZ2NLA2bVRhE/mqECj34anJGJwwkHz7pDVmYUwnc1wdR0ZvG
0KF54JPDlK9HTLnuru2Lm2h4fU2JDIsKvY3bheELkPE3Cm+A6OI7SIEm2teEGzCmxqFlAhfQ3gCc
IC3k0Zr7p72Rq3aiLFaE628HkL2V09CMq3jx8pw2IQ+aUs+dNn0S9X6cYcN4EiyHyaOrCcv0UFRm
evxztToN+2swUhJEcm2C1eemX8LVb4ofRn9tGAFaSvAy+nqhJRiPgBuz4v0jogu/fDCWiHJx3ppg
jT1Ym4mhYgS+lsZHqcodxBKmVoUI3+3ud5pUlm32V9bywtEUqAEJsOEgO6UShlKK/TNWzIXVXkLs
AYAGwOQOpAsUfOaTi4qGhV5QSoYv6rw7Z8eF6RUah+FQ1RJj7UYoY61FPBztuyQsIdXRHYw09xVw
jOnkLPsD/wG74+/SXXmKn5AGUCUAeOvHGAUdA6YGmCDTPqZaWO1weE7F1ZEUCXzndQ+KQEmWxL1+
Rge2N8qmSIs85kJRSCyD859WuB1gcZQ/uskEXNJebK/FAyYqYD+yeAjquwLFMUqTEsTyjimG2yTA
LrkXXRHVTxHIk+nSuHC52sDgcS5l6Jc6Z2ASH5zH/fDOlj9ssY+VGm5cw2nSeZ9vucHfRS2RPsl0
i6krGJBYBqO+eFjKP1m6wFiilKHib9Z5VtLoBnJFAgRi66evPkYaiGb8Mt2y4YF3CeHyntn7LDBc
uaIjqHgS1aAJTsKaVdzDBzTcNPVfxSdg6kZcoJpq27NmWmPEPn/cyXIj7JovYsP2g8yjGeY1SFLU
2bgodbBimvi7FQ3grFMI41A0/j7jJLoPd4DJfNS1k5S1Ci5Gc8a1/jujiUAkRZnrC3nkRMr+ZAl/
QzeNWpBqPBHb7jZGLGBsYZWAhVuh+srix9z/d5vkATWY6n7ugTSV4NRHcd8XMz+Nav3leBrjM8hb
JLSE4OrC5POdeR85hm5/C+r9Dsdid/bRJ9LaQt/7oLKCHQargCkTfIOnjw1vRL8I20tRwoBtvsC1
D+JqI89mgkdJdHTLcQglEXTgSivISg+KemBFtJZgDBjZpv0OLARekdnt+jPg83c5sZtjV5QlVZuY
oM+SEBXEeb5IrZZFfavd2srDSJpVsgpiFiqsPWYDc7BVVuZ2OCXPVRH+KEKqCFNX7PpO3eWC4iU4
yrk3JbM5DcPMC6/k5tYZirXKz9TKIC7glnu6ULewqSNu1J4YmRaXDnpMDj7779fKxyi+6CzdGdfj
3RrCG/uoICFBKolfUwcy03gsHsYU7FTNwMUels5iCqofwMZMZuNlnIvPtg9S1rCa6wbQyo2gisZt
BLxY7MwPu2hhTuzxUAI5/a8nXUNT4YPejyiNNxreWb93/mxY3cuuc064Pc0ew1OytctDtCD7yrrO
znjDZFiOYN8bm+TITp53v3EPvM2tfhYz29emicEEb5qDj4Rd7iJtaofpEHKnvJr7St0BBfH/00PE
dy6v85UnPA3NW+vl+eIvE5iL/t4oKPYUjrL8+7Q3B5qlDzHao+hQmwIst3HLZFKAqHEyjMciK0ie
I1eUdPsbzCAz5yvmXXj9aaJTkD1MYAh2+piiPHB+4uMY9AFu5PciE0eLO4+ta3Fai5UgA2D6RBuD
TdM8Pj+9UGuQkjkNfrRsAdUZg5uzV+G4+JdBuZyMC2u7kiXaCu1sew555AIxnB79eZFPqxw30rCc
VUd2+FMAax42CKXnB2x9OuuWECN0X0V9zz7RburjBFw0jOojj+a5Y+KuTlux6LWXkmCTq6EXfno7
46x3p3ssqK4bqSVybEy9H9k+rpeoP5aBsvNDZ6vKSthZIKn94hSDq/dIuPNXwd6BJM9G8GmJKkX7
hmCTablII7kEgWfj2XhB8lkTIN8pf6BOM8+IZAOLqRIBINEe7/Z2LKQ2YCO79IHiGd+y37V7ODS8
IJaFsgMxHQisgDltgvbOS8PsQ3I9DJcgdUTcRyjLxdFAfCVryp00TB+YEbyikxtDUyFRGOWIT2h1
ND+A+TBdhHXLGISld1xI5kivKaENT6N0lXxlRaSwYcK6W0pwe42S7MTzcBrOPyG6jmitBXY6Cx0d
IKg0r9ZWbPbwhMqwGvKc32ki8IxZB1MrdOcU1h/LBvf2Th+/1qPzfSIDGbBV4qrq+UOq5O0wzrAF
e53XFedyO8DzYxqwQsnAvQffyh+sxKWpcUvyx5cWd2XedhWoLPairiBX/1rxsulfYMxpL/WblFC2
9nMlhWIMIhzVrFFVz19m3AeY4l1m/mol4OOuZjjO4LnpH+Jv+t7vznBMtz1DAO7IPff74pryPUO5
ib51nBQuW8V3zJog9pG1+tojV0DCV0zkWWsjfUW02msDMvyvBQVXVWxa7kI4a3tp87NQNpojNalm
de9BSkP2CIWnwZ4LeP+5x2c1cWIMVeyzxy03K3zW91SnC6q3mjgjIMcLe+uFmABt6qgVaFu8D0GD
isTviZWL+AceLLR7hz76QbuAfeSH7gD5qB7UZuzu4dqIxsLV+f0V5lHo4/NbbVBeT9ZxHIwRHrBo
nGDICPDK1hABqlefkITmXeSgJst0BGU9JzauXvoIvGQJpMSPl2hC9B3wWyu+iX+V/sEzzs808J/P
muebcpN8RkokphzbsxH9Yb5b/RZx4MTNZiRBAuV7a1B7dgKQzw8Ux3ia8VDg9IryTBTFQgDh+v9A
rhabb1iPMbIq4jPyc4uXisHg8we6uqlBl4NpemsqPpYXqOmpOX7SIR4xPuC9Nk4GsKEC8S3hxEsx
wSyyl3yNVszAdJwZYcMO7b6+daftrJs49xEONVevIWW4kJsHim2LvJLUh54qu2GCAKbDBx2enrVX
1FLoqqe2VCGY8/ia7ya0P8hFhK8yx0xbo4VOOv3/tVKbdHlzISl3KNWuYp5uN2aldfaJPD5bJi6L
GZbnjjkr8cnNpsQsWWH1J3pOTNxdhoPPsL6Bpsmvge4xQBLZgmFzKqGXn9kTMYUeLC08hl0kYc0Y
jMB90Cuyy1e4iAkXfVqlFR7uAOouwLyCN0BfCIbH9XQSgphSXhiRqJLpjjT7D8v2zWiIqhLQYLrr
5EcY1IakTmWleWHHND1/aguDvhsaMjUxtDJy5FLpW5KzMAUj1OvzbmEN/xuADMrUtYAGlkROgm+O
3FwbEqdWFzcNUO03oRb+zGrw3oBuuVnCMFANPKGDUPxrgmVXGIvF3lmTVyiEvCmwDzGGeRtYG8uU
aJ0oZRO4oQAZk+6n4Qm90TnDDdiNdmDayufXTw9V0tey4oz1U8xhKm3PvkC7KBzUK/8M1nrf5NRe
bkvr/+d83cNNXpN36DRinwxrtNr2R/nDBhk6lyEMy6kwVKaJ1YgjEFpwTCk6Lagbih/rslY88dN8
iJuhCegz7HZYh8/zsIY3Yudj0XqH2JJux0skqAb3nNcusAvg5zUlVgfcd8JLusa3N3tXDUbSKE9x
DbtRZ57ok1CnD3Ijc66IXah4JL9xjQ17VwdMCXG7TGVpIWPOXTYBH5NKSIN7Y5hxvO7QSPhnRTNQ
JDKTpbnpyXh4TC4aM2u6Z3pUkXTIFbcCb+FVB9o0QI+KEQCsOzgsSgPjPWZjEYjFad07kNYiT7qH
BVIDHeCN5u/fllW0MT5rBtZbCDb2+7B0t71agTxCGwrufLSBfqBMGjYaRPUdBSWuBqTg1mhc/EVl
mY/086sBj66L0HMGVdfYnKnc27MgEY/5298uZu7o2DdFX1LpGY9GITXASBIkZ73Q05M+yxjeNzqP
Ea0iRGqN834umI3JwC5zswEuogaQCImIMipgg14NaGa9Mf3Q0bSmsoULhQ3GrS9Y6Xon0MzFKC9m
yVMIsCCILFvzfqMWuaUj6rvQm0SylZoYehhnUicCWIQ1UWFtiViVF5tkZKyDALZoC4lUW6Nczkah
OJTsvWR6SWppWzRW+J4Wxm4Yvsm4OFScpfYjQ56ymYqhd6aJ3Eos+Fm3A2YOWTD/CQ2NvSapwYm/
yeW5SylPq98HPpKirw9qMQe4Frs6163vRsP/r/t3ha11sRIm2bxYJlMqsZEp3sLMPaj68Pt89q70
gxRHCaT1DkJMvLOyWuiGuxl5B9i96g+dU7M8kFInLHq29GpSr3w8yOiytN15fCsXguweikc+Tn4i
u06jpuI2ytkEQoOR0DtEZKPzwjn/PJcsImC3TYOK5P+3xR2efJfD/xKLvSPDjohh5d6k9Fg2D+Pd
L9dIpQuq3fJBmT8kHlTZVCDW1H0d3V5e9tPGksTIgcyy9+3nQ+qq1A0H72BiIJHVLj6h4ECSXSxQ
GSFviJaEnz1PVxdAT87OMSqjc+4UVEKsdt8HUzZ0iVD/gzL4d+JWbqURjfZn3L5/umnL+E2uVGRm
v3/CgZZdmqDlpDQ0S6Ye3zOzTargO3zTYKpIttWy/79dkD2+T+PXsIf/o44M5463RUVjwKuyhtIW
0ntphFouCScg3iPXjPcQFQ0DlYZB4QS3VEnMonSVhvYZ7XjQWogjZs2IU+pm1mH5QnWVRfAs5OwC
CqyX1zmAG5uwS9DVDV7yK8hl0eAMqQZZqOcL4Vvly0MuiiBV9pNwO3FP2vz9hx6znrQUclMxN6bQ
dW/jif69ALmoAI9qZaLbmwFUlwwGySETuxkSNbDsX0Q6qJkffbx+SJfl5Z5LxGCbq8r1tBeRXmfL
ZbLjrKT6kkKmlL1VipcDCz2mhEghbLzW14VByKUb+bOrfkt6gGub2uzyNzQmWzEbNgWuBl8zywtq
S08GG8r5lfjeJu64YCKhFO2ENQE9JEuBMaxyDqFEoFhitQ1Lz4Pzd3W2bfaRj1LBlBKyC8CZtX5j
iB3+q66BYzAzYgIJ+uDInhsLE5zHWR9OZT1LMBVL9PkMbnkEx6dmJwXrGIV1k2JkO4Lg4Q6N7mLY
XGBXvDT4mCBeygtUd6M/9LmWQEu01taCSYBSIfu2geMojbB4y1JSDXmY6u8abqtmLbnAQusqv4L/
KqSkT0cAFN19j2Bt4LyP3PLFwwJx9hhA2G3pW/n2t9atRUA4JXf2u9QOh8vMdd4c7oIJY+SRgcbH
a5M6sV01Z/pQNoufmrnvpyss1QFKnB+NMRPHgJ5tADhO3qdYA1y0YpQZw09ok8iSFa3AbJKe/TM6
j8SuSBA0BTK/bnf+8m3I+f1Wj/u/qvdEdfDWBEON3UjKC9RJbjQqWboWXEa7/4NuKYBgprBrumCc
dsEJTw7D+d3+YpiWqAyHWiYuwMD6m+l9mTcbQxfp5zVZhVwS87T4fP4TbaAdh08rllWMLJ8O9LZc
m3ewY1AuzIc8dHklg7BMjNJ3k1p2Hz5i2MV3ZYOKO07bk9CM9RZ/s+bfTt7tzJ/2zvLiAlhLD1mX
uQeB+2nu8VhinhVXxyBhOWFVQOgzlCWc3XSKVen80qKw9v7JvBgLD7vZs44T0/Ei8cOHxKsgte3x
21dlqFxrwp5XYsDfdcPuHwYjn8mgbKEAOOc4YxDZtqLEm58CpkB3JKUGLUSMUlnZ5vZxK6iKSGId
sVuaivtxUnGLFjgPZ66mxy1q7umwrmohmiYJrLXnQmvP/Noomlb+5mB50RDZyKa+NGXEOOFVV+4k
F1jjXYffjKKi3u6C8tUPoOKHk5umuX4ZjoFsTNKmU/INyegW/wTuv4oL3oRuEC7kmwmFBSvCG5pt
RJHoCSkKFR1s8s2vuBA4lrGQ2/sladdq0pOQESESZQntivijjgJCfio5NT1MzoUjDWDLSEoRGTbw
Mthhhif5tISYu918fwHoTPp3RmNHQuGUJnrKTLNpondWSqYC4KorsBj3/v5Biw/ci51j7J9DEdZs
QNsKsrgu2i+fKeghsAekB4WpKyP3BQIDriyQx6GH+r1Yhb/XnvGjPrHPoEECE3MAnXYO1D03hX+/
QJpvKQd4MpchwRUQUaLt3oOtyE40jToK/QPSrsGOUPwYhXOz7jYjZPzyzWfz0Mttdwl6iNg0hnZj
1Ylyyh+znfnbyoLj3TNNC531N9YUXaEq2wj9OMPj1Lx40XFTjo0ieHGbJFz0Ut80WLQZ7k03vQdG
X0YykVHu3W4gh86w57YxnbpCmPufRdPuYfvSwL70V46sFYd7WkJY9rT7/hUTo5ryHM7uIOgpZQdZ
bOm4c5qdoXujtwBiyXbM6xeIpyxThuTkisqqQXHt1HVAxmtwqLkgc9VmbzgksfrCojNAz8nc/ihY
tmyJwoWRXwvYUnPiwWGLROxZA0M+7N8qknsvOqKUv3dm2onysfvrHdb8n7qh4Wx+8Olno5Rom4+v
fj+OAIhGI+z6EqaquVA6+4N7mjPcah9Le5h6hTnUpthGVWbUhSFCDApvotE1nYoAoDIjUNndMenB
HUntpi497fKLK6JoSxNM7rw1btxj15WqafjTHVr9mwCN6yeWkaVi7HCR2PBRdalFxzfGCm84GkQ0
FSZNOCyknuNcFBEaPq+AHf84bLWQJV5uITcgVcWK3mM70DEtfcAaJ+c3B8FSe7P3SWfUhCwp7OQg
cDS52DtzkPXKFDLvWBYlDBp0Q3/E3OEfuNTBLKzRgzQtYwCMbn888C27ZfA/UxYCO1VxuXKzunjf
vkpA78O1pYZXer7yFXlpt6pOxisXf4g1avdbkjVLd2AK1yOq6HZGwQ2RKQZGoHhVlHQCgCw++0qA
Sz2605jQGhXtAivWuiV37cy6qkjb0fW6yCkqy3XJudCyw0ikIvSVjhma/3a3dQi5dLCUI4yjDmdz
ftLH77MObhJDaPJzaZJMgJg3zDEpkxDSI0SpBpS725hq6k9RNrvypSU5wGZhRthCm+L7xmE2tz32
5dM+GYWfdAP5FPVyWguNak4jJY40u5bXAlezE5K/4qh9eHVezSIb5hnsdonh7nH8NYSwKM9JLX8i
fwrFUTvZ222pUz6hrT1o9CuVuqcnVc5Hq7D55M6qnaFhDyMlriKNMy/tVl4ZV8Q2smScaP7/pqCQ
EYSTUMsHSqp6o3GHSb3JJzHcDj1dqeXbyV7g8RH4qoAwJ5uS+lGJj9vVHeBCRl7oR0TSp7EbjQyr
XK5wTWYHDPbTpZnr2bkET1/Seqwd+tyIb5gm3n++dHwV4S149cfBPI4QSdt0JdBTtUVFQjsrupvJ
rgc67dhsMBG3a0KWxuCNRd2/D3parb7mhDbCmTdll/yULaKKNOgIhP1VabIxcKG+d92wcIaZHCAc
H1pPG3QyO5NjeBlB6MxoOOB2VZ1QzD8JuyESrWT6MzupffGufml5dyjAr9J3a46IMCtFTGNtGenx
vLLCyt+Ad3mEM89jL3luUxrwG3abVUngAWdcj6lsd7elmfQI0bnrstkRse2pVMvQHuMc6TNgn7N2
H1qGgxsfD21NLvYtkFBMsr2BDzb0okEnV9EGwYnMqT2+3X3+20B9MiEzA+RXeWqHlDTKjk7nNjHS
AVKGhWYLzOFudV09zoyYK0mXhl8p6sc7gtotZJCqwDE7YPNEPBxFPjQKyPNX4kWaIEbjykLC1W2Q
0QaUbzcEjKh48QSHx0WUj0C428/rwI0XKFzTHoyMl7h1bOfnJ4vSau6MUD5O3TmO3ouaRdNEwQNX
rVnnoI+t0rB6zqM2ZWQKwCV13lZeKUjyWb3Ty5kvUESeWJoKFHBNX1Y6GCTPme9pZW35tMhDElkS
uStGYzokWLY8O9iF7HUNtIxRfxsQUf2rgL5g0mdIKEHQhuHj2S7T1HLkVrIAnkY4MJUVPgO83KTm
pU9V07QC2QlgTLO0sqHF/5I2pdRLDqg8vw2LysfwEidrlfjrtYn9obDKJQYry4V4gWSrnl94PxDE
e2ZAgXQcdXrX9+bdLBjDk57Oy2NfhtomdJ+uOVmQEm/ZILJaYBqyGFeQlZNhu0OfcYA+b51t2Rla
S4ZYorRf5ThATAp/GRUNWh0S/sIQHH8azx/eFfWWyyssyCBOPvqb/0RWO5dqf4mvAtAD5KyUo2cK
tWcm0GrfK1VRPMQkBisBCTeP0qF13JSWRVPAuFXW3hEK9FNm2TisWetekUxxo0thAo0fcEnQZsds
LjB+6vyCb/0kT1HYnKnn54uc5Snf3yMJBz/uNg6oUML31npnDbP0rfWpra/atsPmXzgd0VQSLUIO
UFcWlDxv5lBFu4CJHaWNjqjN6qNOKYRlblely616OPKXG9dH2I6hpx/sFfhyzVQCNd+WEyNHSLqt
7iv/mCT8MZ0+8gdoj9gnM8BbokhszUI2f2koJZty/mzDXYgdlslGdjKAgDUJgpW9UJMn7c+hCOEi
gpvyJM33fVsWswLvIa8BPUhz45vRgtL+mXkFp2HNxFqpd92vAsnOFMOM1Yyq3jt57Cxueh2y5bjc
SPW6Y7Iqu3601aHgUTgxO/GHVpr2BfmKrtyDR6R21YMQg5WFxLo/gGtqGNwlXnkNg5ZFCeSEWHxc
3mkla/KYXk1sUd9VqlC6Z+IP8NLg3YNL1Iu0FeWrjnOvVEtoOHAlDPjKyq5ifASANG5w3wAGzR5n
11qEKOj9ume0U2gukWeV3oXbMBk3dYDMnjkm8egu8by5kbS+0dgkC4+NvSYXTeRSdQZ8I/eIUFbU
2tP986x85xfdztRHPmXZOiMUpW/RQbhRbS5edE9cy+/kw18OL6YuOY/G2VFWe4Chj30R3bz5PJEF
xQuIivLn0MYDCjqFXej1rhpvcd4jBS5oB1hXam6yRGa+Q/YcB+yQoaHmwX8inQ2cOuiTZr3bWs5Y
q1GmVXq06Vn6mrWvDLtOEasFCEuAiw3wKcgphz+7HaFTO2u5hilefWJ1Y0fK18M0SqHKxp534H9f
vdiLb5dsE8JlElRImpb+TkedVh/3R4eemOtXIUO+vgADsiIdtWS1MoiqQBYRwSP/1VULTraDXSGr
9ZYErgBWtBcBFR9rvheeiS4PDmMx9BB2eR9oXC0Zb/kFghakNghzBvfUJ4xxrvnKXvb4XWojSjh/
sVLC3uy+TznLc8RfZQn+heoDg4n11ADy9bJ+1J6ZZ6NIvShBPsxf6YPJ6TLM80L5X3iCT+hFGKGP
yBymBR/Z2lhz2A62LP9GurW+/JvcJRZejc09+5trqs/OxjTwYpyu0CclpWOAzRcHrzuvdoZROPpZ
IgFkt2DvJFAkvt08LJqutIZ8m1auc/3AOEcvaUJ/Rg+dCe7HycZ1eiHrPDVWiCjwr0tNW+Lc2+VC
0M6p2A8GPcdn5rL+jcJpKkXx4uXkCFFUBWmnI981eWGJChGalEFTZ/8/aKj6xNTuO2LFk67tkgid
Ylv4Smcpi548c70wJw+ukIrVUlOHqREADclFKg2UnhqcipemJ48dk5MP6/QKh1emNa0tVNnVIkrY
Ex0YtKPbuTA5770zi90W3T/vbMGH/KbigW0VeldOshs3h+oak9zuJ15fMbDFOt/+lPw5ksXAmzCA
gsyaw0S4PKRytkPa4qpS9LmMxZ3XhSARqn43YKx3rpLaNsXPqqSybPa2QTn5Itli1zAe/nVX/nom
679eXvSuuqFwI02BbgwvCZ2f+uIDCfivKPpnust8ur1bc4XIf1DWjshfz5O1uMWgQ9kgLWY0EhEv
0yPUkVerS31iyxT8x1SUJjONX1+gDyoL/6K0jkNezyPLm03EaymgwJDuin3lkTvn1EB/HKrh1Ism
5v4ZcLDAoU1Z1uziVJEWCLCE3UX4zIgTwE9d766Z0/Xy5qJU6kyeJBIMh2I4+JXBQawmci8kbfSF
m+gBx4d7INlwrq311snhiBclNqUOmom4PRCreMWQ8zeGEheM8yr+OrC1c7JTa6H4ne3cIduxnu/y
LGFXozBPKxAfkllSSdsip9nO1iqXd2ozWLQ3AVGJ8WFbEoaubuNjgDmLvj16yEYVHQ3QD+RInY6H
bsRXamJNvdplyFA3Qwg1mzRlE/qZXGI9tAllkToP8GFVmhCVMg5lxMENaugB3g6Xd/ol2KQ901Qc
KScXh0SdovrZGSMIgRMM8mWJ1BTYMHuVHBvhehKDsj1p1uKFXwB1bojGpbedHDWX1QuQNnQEKlMd
lIRFzr/xXWjxCPy5IyZo0buy9IzsFlCK5eZDKm7gad0ep1lxghY954Ap/VE5EscPNNHDv+XPebVh
D4TtLFoWKyLk8Klc21guXJ/l0CFHPXh77essxVCAesVL0LrN+ASE/CWgIIfdwdRziX6A7Fi7iqZJ
qNFBFQ9zfb44YG2CsRXkexP9HYdPr/4UooblkgjPj+GH3/I8IiP5trLhpOjOAfdcITXV2w3Q092j
uoG1gzv4ZT8anmWJDiHQG91Lch0W1bz6ACqA/E7Hxer9pYEex6Aqb0IUnvxYgYLe0VLu7CmqaWtx
8lr5PjRPwCEhOxHFDKf++bydl9tPugVtMcevzwe2+7XpUt0S6n7h8nl3rfj5x5J+q9E18JZLzCgX
imuBRfLn+t1p9MvNgypgYoVeEj/cbsYlsYmF05zf5nm2GqKkwZpGuqfQso8JMrBtyht+obXfJP9h
t2Hywtaf6Qt60knY6hJV5ayhWBvLrWF9GY3bBxxdlCYW0sLyBQz5FbiMAqbONFkFlT/ssdBXac/D
BiIPsQDqNrvC++QaD2aeRcs5oSrwhR9tOCWmERUyak82SSpFdWtIV1N9Np45f8cxAa0i308vHP+y
Qp8IyA0odt4Cj7H8N+xQIOBezz1NW6y4M9cY96qzOMMhrc9O9QEGpHSTUBlR/TVWOmDkkA0bpSEI
iCb323aHegJWYY/b0rxJg8igxwsiHUEXhmCi4kWLHroam89oO95RKcSaIDBAAXvFylFaZwTFfdR2
rVrFuUZIOoWos2yLI3H3R+HQAV430YGAIE80sUqVm7RH9uGGNMeqmkwPfzPR4vV6IHeqWa+6w1IU
Nv+GIZ4JTc0Fu+RGTOppbv2MtWCE0I/dfsrQubtouxIqXVnMPJLzI6MKHb3KgYsGWMQoJ2P4d+XX
7osnnHeJh2mDSSiyxt9dzLm8FjIgW+/w1YbMvLvkoTmJG3Y62aDguTlw5KuD3anEw+lVrKbO8dSy
Tvm7EBurIKujQjbYqGDu91m4s/9sii04Rh94zsMqgrpZAyQCR/z+ve/jY7y4vUca3vDj6pNhxOgQ
5nUYRS6hPUa5PSG02KVLwlmqzZsimv7HCwkMVmihRHFkAqsM6BaKZmbB8Lz0SA7BO6jtVF1oOr4x
zsxpQ+k4+RL91KgL32/96QQLEkUhWhSPRLkiGdPkhIJ8PinBjwjGKzoHzP5v0jmATZHFDsc8uFFM
u4KF5jO1UiTllSzgyiOfEvpm8iWMQp1oFhMOvGViWCu+vFXz7MNvKv2+OtDbCRDcLOflNqnaRhdn
QwWlSz2p9jQyJQxM3Qg0Y0rf5exXGOoiUMgqVVeSBOVEJA+8BdYEY4+sRb/wKOTFijsjeMVgc5TP
Y5qlmtqiaILKiTsZhZFvFLOA4tDuDpLiq2Bl6K/gHvXEwleFB3GjODvBPTRGKHtKAgh80L307Eu1
kukfzWuE1j2zj+j3RXMMKg1Uw5PyNJgxnOt5pMmtvPOpx8FCDo6Qamk6A2PPtY5e0zWanRbRlYhJ
9Uf3qqBMoffKJWF2KiXEo1u2fNCZMZOsD6r4eMy4q2B3+5+SdTEEFIICjyQeqKENPiG9jMKgPtsz
T6laSKGskHShgYf6DlhI4+WqLQbym99I5KbejueIXHNX/F1yVnhF/aJ0LUT6x+HBwjuvSnL1j37V
9GN0gRBpRl4zfI/YHKuThmw6O8zkb9467iEy1c0usgWwrzglbP90cbFV3af+Ngf/FNpxE4zw2Pr1
6zXWavNNCdePq2VAMjZlwyU+3UVB76+YcKoRrvzwIV79abF7eSTIRr5AfzWfCRGBHwIKfFIErkbm
8Wd8Qxvmk3pG7owqj8G47Y1e9dVP/YwCRHxI3ehRoQXmetb2pzhqjbzsX2SkZ6Z61cOXjaOkMXav
tQOstE/3GZFEaJO9DW8lBEjjrM+DywD4VJfOrvx1qY/6RWyLhlGN6QY49elJAnb7OHJHJ+oIEFD0
icn3PrNr4mcRDYCsFIU506i+qt09QuzEN0JYd1rDXempr02JFdhrdGTkJNdlA3wOaJqb3Nqud6cv
+1mAHuUaeAsiKmPx3xjxg8ZowMe6qscLIjvAqX+cBN4bUS60tUXPtbW9I26YtGK/GJ4aKngx1uXb
9eKg6TtRHRb1Z5hnBebYkY9IkDx4QIrUBLV/TyLosN9/ZKBBf3PUDK+PG8CiZwVToSXgwlOFDAze
75EIEwCBOLt1JQc7pRTVik3ZWtpP/uYoYEhWtKIEMcPSTB+MylNcvWEqIwxPhLKZeDkHkGhyGDr+
rmfkDogVP2VaUf1c3XjzNYvw9kVxWVCtQDQ//lYC6FmFCAVcyw04T5c7IUSqMerMLYdn4txEdnNo
R8tywylWVuOUpOb9piPdsUKbS+hQvm4IZmVwMdhoDjd+UnluY96151DS3RVZ1sxQBZd9G2NmEy9a
sxBosGUmyCgLPDGG787kumribe+C/d3Vr6Ri78H97o+9yf3eYI+wTAfDGSCdkGt3WLNfgijwwt9p
uCr2SitvEa4oZGI9moyteZNkHAvXMS5bORtq5hy9x8c29Pvbrd66IbdsbA+WFLGo4bwfoiAK0W5k
yvh+CwwTu6dWrWt6mfB0UEeVZjHjtt1VWAYLVfkLO0DxenUCaQOEikPP3VAbzknZArzrA2+H9eSL
AqJi6DHYjaucOoSb5ZCA1KoS9z/iXg0wEvZGVZppdxo9Zfdngc3/PvD20CBgcqqo5EVgmiJUu0+T
g5dZJWTdYfTKQpuID37Gnk5f4p2NQiETXdmlanbl0gGZS6aJJ53KX/M2E5yB7M9WSoQZER/G2qnR
DGzHusGxpo1eyxyWJ9EnpSgMLY/HrLpSvN85APPWYe/94f2SSG0AQw8Cp0w8sPIwoSrlwT/O3u6i
wxXjG2pvH+W+y+FikMc8PsEyKDoivZKwPtgdyz50e5PRR6FRgBsxFmNpwpQ3VkAjf2YxC/k3LktX
22TODkAWUeKHxYG1MoSQmyeBzI7fQ/2agtUAbQtzQsl1widVoXeT0EFXrwGkHSSu3UgBCRxAMhnB
z7p1YBapkicUUj7OoeHk2gV2bddV73q/AlyCY6a71abjOcWforu40B1WN7Majn1h134OR0vvHtSC
PThJ5QZaJoC3gZSySIa/wI51Q1MB72jfHMfdAo6APUZNR+VsNjlwxkQUs2aAAjJmWGG5exz3Kb7R
4qy2rb0BZBvlbPQ7GPtAcdL/xQEAj5lk7d7EykL9a4YKYv3HpNAVKct3XG8666YKLVqsUdIVwLTH
ouxGiWCz6maNQC+Ejusph/HC93PjH4d2limAzmhFJ7ZJFeJrW4pgMhybIrkzjcH7giYyI+y+XADi
Bl66K4LauasLYryJtAfr6rMLgQKIxLDGJijuHOA8JY09/3DP/EWllXaduM6YYWcAexpCUBxRA7+A
je+gQI2YBAFQQJi8dw7F8KNU6yNmq5IQNRHkKJ3ukzuFkmEoCtjP0VMa1jPPW1TNDQ2aK8Tup2BP
MdTrqjKqJbmyhBCjgojli6lb3D++6B0FqPVs7K1x3vnq+7etbdcOFJnYKXpPsYJw8dv1YcB0b7uR
bnXIUntA5SfImlJWEJT2hVUqEu2exASygnFAMYgQpA4wcGcTITW6rX3DBJitG6x5+dJe93r3+wKA
wIiyI6fo1JzwYE4ABoVukta1Y1qZ2hyh+qmBfx2PCRMpaCQ8XxRPpy9UsPB5lAiH+J38QGZIrLlB
lMXbEcQs1/1gHVz1AL4XYd+VDc0FZGRbCEXAWekY+emTxJiGAQkuvF6M2B7MuFQZyewvLNWR64Ll
CMolwF3oT+og4zD/zVLj3HOnXACIsdcocgFhtjAbSJVVVfxNzT0A7nY28Zl9KU3epJFZaRo7tkpY
3ar2GsAS7X1gVKy0AEfIC4rwlLFK9SgNSv/KOyD3ZWRTb7ko0eGntmk5ffIQjKfx29eyE9/WWgA+
0bUwtwDKI8EZ/7vaf/zeEQhKZLfrd0ovdgx3ZCQeKeXlcmTGPS/rjZA8ZRMPagxH+5QawlXqR3qI
Dcr/6o4uF3VCC126GSHbvszwiNDuXA8R8GINQj5Tumwze1SCXitMu/a+7EcGiBVGkCKyY50ToeHp
IZvj4AXCJS5jCHC2+uUmWtrYLPyqTkAi8YP9q4lEpNcFDSDTu9nCVYIieNjqgTrwjQYQoVBjWQ6u
R3M0j84Y840okyRUZqeJEl6cS9XJgPIaLg+surh/isSV0T2vL1nCuK7TZO1VzJfFSLpYsmV9wUq8
iOFjiDuldY1t3jcbWl7SAk8m5C92isDU8qFYyxu/DB9Eugl1ltdZzdY2LMaJdAldrEmn99a8Xgwq
ZLk27KaBu3swF2ck6EgAtxhkIE+Mu37je/TKHiKA8cAJi3O1GP8hpbdmcU4hsv9ZbVnRjpEBGgOW
Ea4pxrA0/6qbtoYGMHbNsOPoWQpubOV5At5bDuGRpHRN+rpUvbGPFmATXC/pZuGfRbvy/xnZol7c
vKlL+gv18FRGekihwLZUSIIxOCStOUkSWHIz8u1ikN0B1X5CI2iO4mWKloAsnJ4Lyr5ExruPLpkJ
GDCUHwpkPJEjPps+CKNFFyGlKzXi8vQZzvUYnekjcgeK3pwDhcsXtRI//sACy7kDvM3Xj1VFsQiU
zTRwg/z3jJ0OjSHFLVlr8sNVdeFp2HMqzKWtnu1Vw2IpN4FBrTJKBW0xXWXNYtxVWjkR8gCln3kJ
QVDiMDX74yP2rut7e8sXSnoGRhSpuKVuG5Kq2C7kCn2fYcUq3wV5EYejJqOo9pbOaSPxPLbXdMuh
3rIPjfIMdlQkB06tDEBGJDWEqyqQT3ihHZ/AlslT8zqsq3wxdTb1OtNhlYAF5nv68/ljfCMCu3dS
6vvwteJMdynU3RMncMs2dQY9aWS/KGVyPFuVCuReAUCG70v6+oueTUl/sOEp8wPm/nUFjmfcikRM
MisIoi9Yp17MFD+A+Q4Gs+9ctlYejwoUH5ZsQSOIZhZm43TfxB/tsz7ejJyirfjyCUMX1AUcwsPB
HJHyhVzc4lxqZpzX8rrdypXOH93nXbTAHbVDDsQHU/qMdyno0xePR0yS+LA2lB0+zlUIR3IdyOll
oeYof1q1i6D1lP0aT0Tx8YSWif7RN3GwGsoJG+Jh4sT/P0cSKGF/58qUMFRif3HMudNXK2pBoH4G
IqtsO5RbesTZw61KoCrUhmS8zb3SZnKowb41YGZhu3pqpJ+WjYiDta6smMOQbpbdpT2WQR47jIX0
8JGNCGMzXb/b94dgOEJA9BY5gX9/1dQ3cjGnRh2EFyjI/ovKExcVppVNLnRdtCxas59aB5tBOl8p
tff/HRye1c6JQ2IyXoVhuRiHPIc45iQF6FVZuzcEK6fwWSrkbz1cdSaAk9+f/xyosD7vZWBUPOKt
acrYxVzaH9DGlbNATAqRrAOskBoyJVuyizd+EN+tSIpzWvpjTmAgzC5miYZ5dwplzB75Gok7MrDc
GHkIMCaglxkEXjsvOiRNCh85SZUCwhIq9gKcAs/35d6sa27ZaNeVwaA0uhnAJRNViRTA35dsO4IJ
Iy+FvTGKJe5+xTbebx/kUntw5v/3JNzhgtdcyjNs91NmXYU0bkylN06K08NZoTOQZnzrdDDu+Wt0
eXovFi3LOsBSCpIbZ2epIaf+JmFD+NeutMaQH1YsfbnUs0lmUXKmViCTJqiy4M5nDfOI3Bzu9ikV
2P8Pg5ii1Ght//3C2fpOSipLDLPOxLEHwKWTPhK4MNAx5+UdU9W7u7HwLb1ZVTtlVD7C2HJxUfxd
EzVAyNmF2iQMAkVLHCnXhWfgvhSp3xSVT4/gznLE93CmjNdDtdo40ZgX7msYeQuruYkXufD2lD1w
4dW6PDBCxGMnYiLwdPRvM0SbJqkZwdJOnloDHWAoxeShPpYrEey6VVUSetJbdEWr6DmUwzckwtGT
jZ2DlJUGuluSZgqNqzWVdyPTsy7kYmbcY6Vym/nDZmOvyoOXbq1gv/3NdmyK2Ji/hHCZKXYHTCYw
dlZvpAYXjYumSiDfM/AsKKKU200GRhIhhq8HJSkGYLoh+hsLWNg0mVtQlf5qwQrKvaF5CmDEmmUH
OTGnrhBwEwaFJF+FWRhradTrOGjxXwXsyClW6Giw3wj4xkweG1lGKrNc+cIVGRqdunehn4GNKlmw
FC+ptQuo12iohIluLm1gWUHsEZ/DQDK60T6qa+Yu4qoDp9k2SeR0HgJDIYn+P29Kh8OFGVyFdvxU
ALd0d6UiVxVkpwdv1Hl5qYv91ZMV+4sVteh9AhbZvA8ZGjMojJQIYMu9KTxR9FxR6v07gnosJOtD
+BIHIH6CMtv1vHovP6ExKDDGOdo21EvW+RQNUd7u1DZGL/MsFQl/9YXqBBLkI9ZYNnl0Oc/8pV44
uaFZs8cujxQMHJwosWs0wEy5iYa/eoiveLHNVwZBMgS7j4MfUeeo8hiqo++0NBhlKJfBsjRqSPrO
5H9sex8iHRLv0xYu2LzWjpPkA/igkhrpzWgg6t54dEjH+bpUtT8Iqu526RqBvpWlfqtA81zi8u05
dKdfk345VwLjSkZHIEbrFQ5pb/dG5Hr049LiVtI0sGbDO0HxuD1f8VIkeydqBpPYEfronsh3Uf7p
+kvPyLUotZDmHGx/Qj9cHpCXEdEghezqfoIo0rdTvDnMRv33X0TdcbbFW1GCTGtsjABE7eGQDeGW
YueTtRi2Q0ija/gGlmOkh0UKm/iv+u4LqviY0XVSIVD7RlyTF7hvAKKxyftXE2WASzm8H17zIe8h
cFDNcLPnbJUlqAfqbfiXpKNS79R44Srk2XzXarjvkBQJP93SHGpUKTV5LTCWMHiHzEsY4k4crLJ4
FWgpaBxfzhuIs7qyuxFfPxODCOCyLt+qdgL2IK0Fl0ddlj/65eUwnpdd7h6Un+ON5j/Mxde0j22F
VjUUNabA9TdmORL3TBxa6oRS3vQ9zs4PtFayfKFWfoE2J2itvngeuJ+GfrAkBmmMORM69nEnlLwC
NAVSSbz0V++8Ey3wvsS7fwzdBe1/BErqX8qIHNZd9aIrUJQu82SWOgs5ViDZIAbbIKeEVYe7MPWh
sy6bHlphlJKh4Cot5io5zhb4XpcFXZHjoub23X1CwbcelomRJSOyk/jjhIYutfmhL0ldyB0id0YB
wsQvH/jI9YZlufCnuNkc5kqLBnqyAruQZg1/4ab4BOp7ZDq+WK+pPwfpAjJl1MVexPghNg4opCC9
xl08OdZMVcp83wcChNusPXpiSthka03ZWsf1kJaYCa0Rs3DA8PBg3qQ7qdmrlUZavlJceNsvE2xj
mjzzD4itp05mvpgQeSeDuJ7pUvJwLrWbgL1xLr3cg5DBbFwrrqCefyJEfcR4Ls5J/ujk7NG0blch
vGbAl6JEpCWaGns5wp3I8KTjaHAnvKSY+u25jQp/v3hyiuMza94R7cGzsuJkJwNpSpcxZ7DZBMlI
LGGj2DQS4lU5lLWjQm7CsJ0XllrnezZ86zHEPCmQFju7USQuarvGkC8Fh7E5FQZ+V+2Jhc6xMr+0
+RLnfTJqjnjlCZnfedlskOJdWFYxspRFKF94jSvAWJfD/xiRCWVxvuKd+6VCldrQ+GyGmd9gcBvB
t8BhX4Z8lQl53BiELOtA8gPLLZ8B9vtCin34duJ0OWC+TaQZaxUsv8EcKCfcpjOErQS6poR6EifS
V/i9Ood264ce7b5EB6fRZgrZdrrGGXB3AvzieVyV1+WxpaUxxj0SEittJ4hy+nDc2pcv++RVZcDh
M6XMhcHkpdUnU3uG6nco5lXiFTIU1ayIfC8BuDvFXbxHwKAGZn4PmJPKHCCSUgICqHBA+3QQHP0c
Wjw/OARGsiMO5R0tn4QA5Zq46SMoHiu0yp1d7G5ef130TrNgn7kb/0yahSTSBuPUEdHjJgzqD2vP
OqswjFp+EV3GkR2bt2F9Judjh4UMFSDygVk7t71AuWX2lYyD07+lI3Ba0G5dqmSVSIDh2aOSApWs
Q4tNvEac5TDoAIDHlrCFUmhHQKrBR49mVfCJoWod6VpwJr3MdateNfgBRx0GHQu7UNH8yQwgF59y
5xowVPRmQS96B3/V00ysJRDvrYWStxEax2OGLVHyIKI9qqkX1sW5DkT6G1AiSyAmH4Aad9Xz32NJ
s/LxdXJgis1P0q4gda2xSPoYpbmuzjFlbIpyL/e2TYb/Xs9ObZ7n3RJ1ppcCN53GO7na8npjaaKn
l8wc2RdfNOttvVv1eDyvGhAdrbYeuJQ963R512q/VUl+dKNEjXy8FiyxqdxABA3Lzb66VJHdWHi/
qQPG2wHHylUovPG6s23r3srFyozWRjHCV0S071S/kIn0MT8ZbIN0ttzW6hHTsQvggeYce3nKGUeH
umGQ8Je8vyl40xQkPhelJj7OOiYChIzqmXZg/hFIKcP/SEv72jUBzAQJMTJUGhNge1b/qHJ62mu8
v61bSnc0iTaFBZxeP0rAKjmYmKZVMUHUpo9vf+nTYwH/S9WhYHTh+DG9GdvXRCDPu8EguN28uk54
wb3vnUklyujoh1CNp9f3Ibvvx5QfCwumQRtRqrQYf992STj/NaZdidSZguM3+u3BbHaAdDWM05eq
v8YMOr1EBlbqnhlLHe+Hl5D2ZFBCiJFEPVzSr9QTdycLxzOvHsUl1Oa5py6QMx5OurA9XtYtaQDh
/5zBmR+0bOZKwn9Oi/XcyYOS0SlyMa/P++RcQdUYY+2BjKchOpNJDfm1lSbwmT2/huhw0RTwGolL
w3gIcxNm0YZs+jv8KpqUew65sfi8/bRthNFN4LSqsDD+0FUXkZsLuCdjo2fd8Px8bsfB77PpKuSY
fUqJvXbXRby63rRG102vcxk4bocRNIe9wn7H2vi5nTA3aW8JQxG1+B4WIZjscd37ND/4yhhHmhKT
IPiiMsX4f97qL98CPyMb5hoDLpvs/5ODb7ckhK0GeKSOcKY5x8ESZ3D9jEuIrGMAVrlLve6Qnzi4
RhX4Jhq0PbEa1LyY9pax9dwpvQZKfgWxqvDa5f+RySDsRcFtH7HnO7qi/xlxtiQ3lamxpvOVIz+T
iig//WGkxcJ6ZnCclVkDymgRQye/N3cXAypSOMhb13pxCBNh7OEM1a8eGSAAR6xy5uLUWBhcFjKx
pIWkf0WCh+OM82171GD4rVRgezBYSsnOKaw9KiZ79A7NK0y+y6i77CSrmAx5FywyoOdxaoKg17Bo
afHP7Th5HJVrTpMD67ZiOMry4kcb8z3oDMwFsSupB7zykZzoVpiwMIkvbIhMIw2mq4d4xwEkp3QR
dvZhYLI4GeGQwYW+IvBaVoVAt5KDs2AwxzaVjoesfzxB2bAMAnsOSIYYVeBEgQUcGEAc+X3Skeuq
h00NJq3E+oJpEpnBf+ZiZaD78CePXAwmTWFNWwfAjzhXANKIrzx1e9wjOr6KXiVPYCWzjERRtf21
8wMTsIaBsJd302tnDiUalJncixvGsT+SJ8R1mR0cNi9sh0o7ULC1MGcwduwmzavEQAaq23x4xAQO
Lx1Uq5qEHkgIT9Q+03yR4CdsDYczoL0225Zi0W+h4RMy841Oodo18bHkdDk/6tasgw05rWgnizRq
wAm9NnSZjf/TC53AM3+q+wkoIWLNh18EvIRZpggrxXMVFOK6uM/Qp33X5KN9MuntTGM+lU+7m7FW
L7nos9wSy6YftdLLTLJ/OjuX7fbkKc/dpZoHXgPe+XK33BqeYk4UopTXO+Cs8YxJRyI/XdhuIV77
J5xwuZ6Jfn+z6WwyLxiVepku6qQt4xLXvnJx/lDmnk3hVEbrMCTgs84jW9ZL/aDH8MeymzkfGhHH
6c1/5qeS2Qi21ATZ0h/jAKZT5EQf3vDQ3FPCiA/3VyPYd5Pc45/Bk9h0oNUsxenRup0Cvy9gpB8x
S6cP1PZ3MWap4UG3cWqsEMRCoxQZaztWWY1d6DPby/ryA1+ycNOdIQ1f0nikxhBAS9e4HRGwtOuu
8eTCpGPY3A/+fSlMMp4BqealwsemD4Hr85fLIjk4tchj+dW/4JOBCPfGtE/PQSxG50GM23+clBjP
jRz0ZLeVZwrImGurrftI7dGZQOA/T0yKJFI8wzynG3ggFNgAVVhEldi7xF09Kli77/ITNFUt3l6G
1S+5PnoCe9puskU21o4JR/t67VzbC5lHLEpNMYY313OCKGM2+Y25yEmTqR5+6izMDCJrOmCsoPql
wDru8OckgCaKv5zdJYWxwrLeen0Gyj4G3MQFhsPZdx2vZkq+dY04kgWU0qEvtg5I2eWZUVRrUrsN
Z44mB6hn0DPszDcEMT0iyLVS2SizaX9e0eAfNFKHVETZ9x6Wtz4PWmUV/k9hfFIUHBqgFHcNfo0C
LbULjLLlDGPZ4Ulol2XJ2d3BiDsXRKhr3vr4DYYo+W1xq8RzMXGKao/KU7a5pgFOYR0b3uN9t0Bg
sJ1fEaWgVmELftVk3cNeuSXbi+OxPmcXF0S6ml6Vwu1xQHVD87lra4L1yIHuEJNaHPKcSx3sQ1WT
AiRcn83gO0iKHlMn+oRRrfHLg1ps95mevU4Zpi2SccggD9qjg7gd1LLFbtcBZZZznnytQB+1Pt/T
mY2JWlnvwilT8n9A2jwl+UgknsdqNm8B038hBFtJfcUdPGCh9HRDzY2sD0W4+6no5dHE/q0R9dt2
GQwATB8ATWM+BJuDXDCZw+/NoZHHSZBAo4Wzog5hTLBBAlei0rLrheVG+Pcrc2HNJd2fn3pUgy5w
0A13XFz/yzTbcQ/eTQ71DGe6a7Xm3PMcp0MirnOw+D0VWUSCHLEZrX72XtS4GMZDCdwiXHsbeYpc
skQgjrq0LUxBc6UOuMR9LlF5Cd/srftdQ0Yl5ZJwl5n0r5DwAYkKq+pt0JrzN2/7Uwyh7F8CSsPP
blOnymCO+8ldoOT8yVoZcxB3Oibsb+GdIlxwoerwbog0ffPEuVq4ky9PXFeIW/iJPCzhSZkoivZH
v56Cxqxwnq6gFYPBP29zTLwP5PApyOERuRz2S7asxc5CuZIzvxLI6TALtl8ipX7Jspyd5DUJnZzZ
47+39ZtR3hfmfM08a+8PdXGwyQBs2A3dmmutKFXq9hWFei2aDwTLrH54DTkL23ZDtk29WDsuBmnh
7+yakj+g2h6xhIwgkTwKmIAn0WOQWckqIZxwn/wue+0kZiZMMUpQ1zRlqudoJyH6SiEVt5mli2/c
i1O4Ga8fhYoPQ8d4QX2THQ6q6tyZMXHgrJ8ufBOcb9XUieiIcUGce9PZnDcPq0yPPGVltYvem1nL
RqrLwVEo0y8Q0FJke/yS9sIscdsj12SquzkG8iBCPT/HIbGxu2AJCmdTt7nWdgtAU5s1KSLdVYV8
SXbESi3DrCtw3f89KLkeU+6gLqzU74TSz9XXouJ4P0LYLMhUTBZtGOTnEcm6pz5hw13+YXZ0+RMv
KIlYxj26ic052nqxFv9kU4COgR0W/ICpp3B4jX4qzAYm7q+FjuhD9QYKzt4h55YWfXyNdMu2PNSo
BP8dNARWvYQU5abyDRAygl2BAN2hQYqXtjHbyVxkXf5qVrDh6WMQwV2ldttcgd4xGHM/p6PI7iOH
RefYALcFdPrCJHLe1NIZB7ITYcj7iyWJUcLgDK4//IBbMwzYMYI371Bc9VcHAhRiz2SWGTwcX/PE
1jKM/R0YY2Kn5OzRpyNLOuVApSDk+H6d2/BiDZiy3NeNT2VdKkgurM+u0xQRiBFUcS7eqbXxrJp5
A9+PcyoRTkqDBlrU4uBKO7EA46XkP3hxxE7zB8FCH4Ff+PCYoBd2Y/+Bli1XVhBwtdKIi/Ews2DX
4omLwqwTBDBa2xORuLO/AJOtPYMsROTDjJSXr67duRhCAE1WI3ajq684Vcv40FT2l6jqJ7bOF1Jb
56Z1ibjm2nR80s5tQ7jUIyfx/wjdAFR06JzCetCbrep/3a3HRuJ6WOBTfNajLcy/7FMLvDjA7gUl
W9ajhMpLCSJDcpAKrgsU1hLhInjonO8KECP5AtBiQjcq9UUWgyCqi91wJu7QUuLkPyviRdMJUFln
3/tdj35HfERTbRZQMM/XgP+qgkHSXgOCQr4oFerx+aNl8IndWwG2cSQA9yvZqovM9s3eb6Rh/dfR
onlwOxu+XzXsjeY4R1p0qgf72u3rFxftEfxxaitHvpTwhg4H4vsAryoNGNoyR8rMi3Bx6ML+G1Zj
uDqeB9dzNR/cTkOfKtajXKSoN9S0B4rXTSifcTNBJMRDycZlXlw70YFptHNZTFLVV61OQhixYENQ
M59wVtNE70xSmlIhdGd6ucbOQFq0JOR6d3nI8nvWWUsIu8kzUeWnfkuAiRqpui7orIKZokD60zfu
HgXund1N4aroD6mhr1FcHXbMrIzGgnNSZv6Pz+cPpPcXP+8WORYI1oKVcbIrRGIELKSDtj/XSwrz
04fWQn1LI2K83swjJoioYbeLAfYP7s7meHKzszLZbVRsT8kretcdlRZvEJSFbtbFZAiS68C3c4v8
jLeOZZn+tTF0HNd6UJoxB1+mtU5qH+aHCRj2B0vxxfur2QRlQBx6n66gQjTU3VOIhI/tYyuMzYUb
iZAGn4eUoqYlqRdhG/fXWXhQEZrs8lK4diYU7YNjvwPCuoqgzBNDCgSVtEtvwvwhppQoDwIZoqF6
0nrurA7fq9QAcpxQAIn4LvzWADg21ssWfBXOuLv54mgBiARxRKcTI2oka/3+lrDvXmIv5Y2EnsK1
IZIs+ZIc3hpSOi0nu4j9Yr0Ug5UhY2/XRBrwNcMCflc8MQLQ+kd7EEeVx5Hjl8uZkSqTBCB7CPvS
mXEyVBI7k6gj0LrRqApEgH3rBIQJx46YBGdJ32L++04R/pC5OsMqyQSWY/6E67kq6uaA2TdkrC2v
AbUUZpqX4C6NiEnsA4UVZPcF02NOA1OWDgk9j+U7vM7x6/jraoC0tyBcqItlicYuQZ0m8FinAmAB
26kVhQEkUSPX9VjR7FucKVOjtI3eGpEYqANRcHvhAb+KQC/50kEjmaLMpMGuDMenFnarE6wn+i0L
iKX6MmDwYLSoIlrrE9QuexkKpwLfhSjw6k/mGY3j7+oHhX5EdsO87uAkGMMofEoe5uD6zLzIsMPk
c/56FxNEbOP3FndadS4uP/R6OfB92a5vQ0CzFl61scOx4KfiNFQf5nxBfKXL9AQvC9/n4UXQscwN
fIDyc9oxYoh0B4zE9xcxOf3Bgxp9dCBvQ5PXaPLdkP0ubaBFbNDMO5q01RYlf4nx/UVSlcTF7d5/
M1x0ZX1z4RSzZWSNi3PjctnVhRm2Tl3Unn8xXkcCs4Y0okFIFdJI0cteTyDQzPxOYZi1GMckiN5C
WjIxzNJe6UF7IHNpwGAYwJSJMoJ2hBO0AbsnTm+kqlL78ULj8G2zY620FU0EiYxfSgUcB6sd+//s
6VbQi/HuiCghGNtpOHTRVGfJLqd6FzT1p5s1NVG4DU8TcDxXjW8lKEJH/4xzAklt1P6AeWGvNfW5
xcLbL7+tdy/wZe+9LlUVRvNPf33wNqQIJrNhWjTMlZFiZ2Ah3IE7Uqr5fWdBX9RihgOTx+kR4tWe
gHwh/sTV9hTX6ceKcyfCPnoz2DI6qbOs41JliL8P+RQf4h+Up887RFVAUUveMo7KBQwUqEnIN+gp
yzfneyxJEdRbtc+fXmVlMxoCLpId4u6s2YnWNaGE30/miZRHkDsc5G3iloRlFalWEsIGudiAx/3F
+JBz3lvrGy3SZ8sfJWyvzTkfY2nOdaWHA9ILtQLDw9B9/QsMCCu1f1kpd3FmK8oN1dgCh+0m7+Fq
QbsNG1ui6U+TT3giWmU5h/Og1osMbmFxG290VGTb8GvkQOCRcGD0FaXlWcedx0ywqckTjY4mzXzi
bs4M7ZbKceb0HmMOTY2DWzX2JoUG0Jb+IKdhvYrKj7CTunmzjjnICM7j23SVRKCuCTRlitunEei9
PfPsJ9+F/o5OkXi/HwlEok3v56sBvytEs/09ZXeIc8lKsH18VIptmXfsgbQX3cU0lUrZMyOYl9Qp
b1Wiw9KA/S3g5XKI70B0QXQIFzrPoRhZnx0nBt0/c/ZJTz3bvXy0byYwyAuiFFNrHqaXQJ0GYPwS
1fafEjB/O89/AqPj2A0Sabso+wekXNxR+ExLSZFn5MM6gqWiiJeA7ez+SMabUOaB0L9uf3VWxB52
VIvT0faWBFrHEw4R+vGdntPZqxLZrdGMp7PL3trkOXgUv7tD2RA9VYgCvyT9j47mUeHTRLdvVmS1
QHdii7Fbbn5m6edb3pNFpMjvlnAvN9oOtyNq9pcZgRWfk+m1LWhfmYYJFDx3LDsM4CNQy8vphlU/
Leek5NN8sVkxhJ+FcTKXECGfm0zSSqQG/HYy9YMRUXOAAbPhaKAaJj0BGdxE735UJNAz2de6pAx5
GVkjVePOSmElzZKoqqaze1HxFV2VoTQD4oTiI0KKb1b1KE59btLDL+O9H2pzguORsDaZzurwB36Q
3Vr8sDHvEe5Y/avMLviMD401SA0rB5sv3+qLly+La+IgfHNagPNFwJ1f3W9iYL7HOYkVkguCgP5W
bbCSrCAv91OCxyoKV9ItwvWp5b6RQbpc9MPNEKYXMhFD2FYtS/UCnC78o0jUFs6zVvB8nbKU0vp1
nV8Ah5OZSKXLn6xfRF8mSq/whmvGaf0w8KE+cWRByeGJTuouQUo2hQnOPd2mxejr4VVBpmrX8ew0
V7hJRolsQLvBYhnwx8oHzU6++K/1t+N8WQhhmdLTnZ4k4Y8FVI9cnUb1P5Q4iA1KClQaTBqTSdmi
CRhoejtzr9V4oNkahUrFOqMdsuJ8Ng8FR0RHvJBcTsv1HEV1789JOZVYxnj10vYfA+XjsWM05YQD
79mWpKWdXHfcDLNOJwVmrGtsfM5kqpXb+JCG5jAxyRBadwd0ZbaZSOgAyJ19LMd4BPlQTRsQDXle
PEY8rJFiNFTbKmnj8Vn7a58PlhepqN6Rw5IbQEkYboSDBN/p629n6IqHwngFAonZWa+KB6lihvlw
IwLNs76wxuFAmdX0tSJxHOXPiuuFUCWCfhJCoNqSSufb6MOu+BB2qELWTOyxeh9nDFpbM+dWfxDS
x/s6/RcmUv3xSdMUhvlxMxqI/etR5tnCfRVz+uktVoIJZMafdHSV8i+2IMxGEqLQ2FNCJLBKo+hh
RmFN/0PHQllLEHfEGJX/BZFw7QvWqO9LNlL0r5lrDFxhKLgcuegpqQPYvqpBHPNipCK7DMhFEwRP
Ofh2PHqMWwy3RcULht0auNIH/QmeqY5EXhErqR7tp+OylVVNPi/6E84ek85g73+opeZ703VwCi14
g9CPef01dNEnUOT9cpTcxkS8hMce59uUIm24uiswJFmqfHbEmc+Nem9855smpXjs+vHS61LoGErq
pCvcdn3Z9k3v+aVRYVQ+NNvNGbAPn3xEBmx5ymncIOnElorej7lN1JTLgYP5ZrNdCCE3IYb+oMCX
VQbkZkJ/oY42LmHY1+0dqtqttz9PwGkg0f7OlxmemIvNKXxbrX/UfivJ/WASl0Qdc1NwgeakRmau
DFfLTBAhzaAK1VdRQH2MS4v39EFkeJdcFPvvMnCu4NrS1APnxUtneqXgaqTMExnRRazDi9/5IeXj
cWyo3o2fxPCNsn97X1p+ygNW9sWeJFow6wtJtlyCYJZHX9znnu0HsNc6YHX+fXQAWiJ6jZCfMcFA
p+efeG5uSCG62xeNWtS7tv2n4I2WG0rBT41I1A43o33OKXk8UgTy31kr5C+mdKvVQBtGj2+apSmE
OUkjj9FTyRAvcDwgsZnpQNQzWYjebQ4AUQ2msUQImL34c08UKS8aqw381cuQxjZ1BAwjfPUkvuU/
lJFW3h8l5HwXrNPkYtI/XWuwX1kRTbmqXx+xAzbxx153aCNQmHBOwmiJHiZiSPK8P7Z0P9Iboqae
+5KZlibQeVk2QZsLnJmFmfQgXxJ89I+PChRl6nFuZjZ/9H2mBsfGquF8MTUnR0QKZ8ZICNrI6hOD
cuf5DniJJMUUr8mIJdmJnxsHuzJXvQkC4eIKHy2pUbTjWHlhXMyPQlv7VR/v93aCleN5a5lDjRSl
IHI7NuJYZQVsQa79kE/Fd05+WPNWSDtEo28dRYsuXsf5zYtNXF2McsGJ9+2JCJbYfqtj7k3PIFGI
XViQA6Bj77aRTvR3GSei7lMBFimxYMHUGLy/1RG2Ufi0rI636ulFZDCIFgnzvQI7sJFjnKDn0ULv
rAdta4i64/oFXP5aZPrhV3aH7X7tLZfOmvaBIGhAtLQvwb0IqpZtgyjmDNaq6hCnVpfIM/olfVii
8//dz8kNbQBOV5Snet91cFLNlzrKD+DYnSredMF3VIKDQfoocqVt2uQYi1joVNUa+nMAAPJCmAdn
dpawypy+ETZJy5VG0khnSQmAFiXeCAtj/Es+vj+RAyxGTuD9E1YQwuSQvnx/4vqCSTRmP0SHya8H
ndZJ2AnNXvvlPWOVLX62EsAmsgvOuYMxWZpkT+Pfhj0p6BDT6k3HHiCnOxN/8w7lnvNeA9fy6Vv0
9ZiguMDjG3s+PxPcKe3zBhQylSV4a3YheKsJTXj2BtS2sPxkLUNN0S4nZrXrbnfYOQvqbPKdLj4i
wCz4tgLz5tiC/kwhT6GjKc2KxrdizSlY9OGouasRD2LFL7B6Q06jy8SyFLWZfmK1mLfXzJFD5WGm
wxcGKGcXUSK6aUtOGUuOSmq7n298p4ASFtfWHvWHp8iJbw+IYs427C/Sti0KU9QHhOojOwweNTSi
mLq7Y3RX3kHf98fRgKlLn8/PwXuJWhHlZR4NpNZZ0QLSjdW66CHD5OTw3OoqIFMkh/teCOSVoQen
TzwoIqBOCYTGAJYDRB3KxUVqACWLAk9twJVkQmi2QkHdnBF3BRniv3+VwTTq3oeufXJu2oGtrufF
pT4Ksur8UywhfDMddh11FupCNukHxW/3CAKuwId1Y9bvWFw9pkXVB7DeR7AxvADZjTtEPy5ANswa
b0u5FNX6cHxOdAFKytIpYmbfkiDMf2dzuGMzxKuoqGdjtN6uTytL6UZNchrfSR3brW2UrEhmF7B+
xaOxtOOijMrxwFxRU9A7XghyDVGlfKNnjGkl8pGEHL+BPz+FAH7EH8na7VT7ixYaIob6hlJl2fPg
ZNGhMEjOOKvRU0fkBgCOvSoewfCNmCtQB0JJAqEhqIaGIVyUADARrOLspOz9Q4ZGtXS6Bbs7DO+T
HGTBiiBOQgWaaWMBD3hyRQzqg1ArI0tS7rqYxqV4DmmcDeuyWJSdk9LI/18qushLk8g6++BAoJPS
jjuJ2WzCRumUbdb+7hS7fm4HSoCwxtynfsyG95k8TWnAgIv/YM84mF4C4FpUcaYo6zOQ4pvraqY9
lbLdNUvz4FhHOCVFmcQVwxNel/ow+nTm7AVwBEEQwm3rpUfJDUX942blKZFqNmUDXH5YzTMWx9bZ
aTHWnt2RcBhVOTPzF/PGKVDmaziHbd7xxxDlUuEHwTzg+ahY8mIvNOOy2LwiuY0SN/g4FVq9wGaq
U0dcojGjN9LUQ2qHsoJAQ8CYCfmXVR6kkwWRXDGVQymAZWAIpCkuasBWzMbHAP/F1lG7ZUqzsvTK
qdAUVKjwfkf2g8o4XdlbY54QInRab0KoMDwiU5P3s5+0XGW2MR3C5XDve4kz07nKHj1asm+bk0Vm
QEmEUJQYnI37u41sIzlV9ZxuxCikcMHL78UTOZTf4nb4hOevRYT0tmS+a16zKgpgUqHyy2vrwTCZ
wzBuN1qS3XjfLkoch9saDHuYCfJdC91W1AS7nTC8S2lqr95FeFlAg/tqKc+PaPKqa4CxiikoIz3P
AaKrIsT55Xzqi30KPBTAo65sAZ7XmOnEGscdHfmdXMhNWKSsl1Q3AfHzQ6jckMZtcwVKGVFtTVgt
LU1F1yIk2E/SwwMeWHv/oKjCZW5f6mv9m+JUromsdAtpoRylNJ9//7hdSdD4fl49ApMFTk5YdoqB
yC5203J0zPaXL6bwMJd5bkrypLlMUIuiaWb+P1lY7+OQoncCTDvcsn9i4N5ESrvgD+vztwd4fJkC
sLHdE3hEw7+Gkuc2uFjATkiN65Bp405nZ7+ek2EHlomcGROL5k5euocZaVZfT5raG/8sHAXzgZ2j
ArHFKA2XmwUiwbWau+HtYWH0vBQANnjSamhWsFGPxT1Tb2C4lCoNnJSB83TjUicIpsIKfSimTdUx
ur8lAMn5II/n8W2k4WlxzMLZdH+XztI7yXbaymRmHbot5T2e5PGvQTjvv/RAuIuKOonCZLBJsQ43
5OgSuohmAoKzpK+b6OuvmT/mq0ZjEIsiCIIizSGCoFZM7QkIZObVGoKOdZCYiKltYtvsWaXVsIjr
aryqXCYGxeCox2Rh2BYSyqdrS3eg/O1SGrBjGvkAD7NYLeI5XSiUe3KLbSCEUBPzwXGi6JgkOmJf
tSODJHbqLXeTDsdKq55vZT7ryeaow5Ekq8iVlSUrm7Z25slZvdpMTJx/0eBQ1kBh25KPTTRTfEZd
xn0+NvU5G36ZbM1bkf9k80p1zJlMrsd3l92XJyPMp+284t7V+mzHDXHX9fShiLa3iBLQr9imah0F
NdCwKYFXCUe1V8RoVaayM4ACcH5tgeP9ZWQ8aD/W49i7HNdqua5Q9x+0AZIBqgYVBSXuKcvN5cvg
2YokNPMzY47cQMAgP8x548/Hx7tBvXrranCBif0tBQFO5O5n9/N/khNIdgi6Hzno68o2wYBjYioT
EE64kD7PW2YIvlKAr963JAKtcaP64dVbIQIBIgVwBQjrUYPEMaN//OdRY9RqUYrEiHBEkpParJfA
X9mQERWaGNDevIlwYakVfnO7aLzhK6nbPHZEuPvAmugYT7pyR55tHsSCBsKb/5dhHSEimpfP0xib
0LEFjUUArjkDnJHKiYiOUU71+1XhVV4VnralBxP7H9LSLcFZ9NDGaN4+D6yNJCBwtT4WUYU8bO0t
NRfixeVXhjGkVPdaoOIIiZ89RjmSUJKub3YU0bGCJBqCjjnwd0jL6rm2AgatOG4ECproYDLvs2rr
3VT/RDAKAnmXSsJkdpdZCBblPAVdjWYM1IcdVUr0y5RhCNdOzo7l+bTcfWFnNVpMc2wamU/4hIHU
xco4cQNz4czEXxAi9Yp1MPo7FWXorOwT0/KM4K1RtUBUagH8i/gnIDQd45yLwHhNh4T3gNbut4o6
s6NdK4UAe637s/r6N0uyiWypN/WoT6RLu4cnn6Xgn/QD/HMKxIIqb3i4eSkymDaX8IJghrjvq/Ju
eBO7Ajh7c61ihMMz7eERUOT1VnqGoq/UrMQMHl5RNZpBNX9m7UWzp50gCtwWkmfbljNDwc+spWM6
f2SsCnIP/IoA4N77s8fs6it+Je+5Bf24JqUUKZRP2u7gV+l1eICtylguBzfye3fpE2syPC14mt9d
8Khujr0nMw4oJm6hzxAQ69+vZ+D3cV4cxmXGEgMHmKPjsR2Xmx+fwRbochGIyXv4ByxqkzVbpH5p
Gehr7ayZ7mzc/h0U76oA1cf7lTdoYDPEOAHsiTtfVUWM5XxM2SZegUZ7YvQWjI6o7285KR+bm8PU
8gYhU8D885y180zxEe2E3I8UIcIY7gTXPu4mceJApuSvji0xX2ZjcAwU3AbyrUTwR0W+b4QXcG+p
9MT1ORo/Z6Nxm8Byh3+Fpyml51izf5ngtlqIRWo3JUyOeneCxQu1r3hL0D279ehPVxAQzgpNm7wn
Wy4G1WXYZ/De6ST4Po/xbl9eR4f40gJ9G45woPqPb/Cu15D5ll5IPhmeHkBo0stRQuNRxKTmHqlI
Wh3SjOBHFPylHqAE3cs3Xk2P6rzTKjpxJxqG3Z8kDqBbR2ayYRMSCEDBGU5sG7tQaW06lIdMAnUY
LbhT47hd9tOLmTI/gugbONyEmcVd9fQCytLNhgIiBHpm/RVdc+84ZkFDLTjod0D8jv5NqtBcdX43
1O5Afk/hIccBei/nrChaXV39N9RqM7kVYh4U4s0vOdPiMQryi2nOr14fXgnOaW8l2sagRNaRU75m
d8E5s0y6j4WDLGTaK8N19SGbUhEK/3TseOvYVtyfaxkZFvMMNLbLDydsl4QiAeoKKQe2Rx/K3NOn
Ps6XNVhTSUer9I1sUkJjEwLWhHEKa/rdjrMSt86DYLtzjzfp68wgQqzEtcIJphxri/XQmTeNbmex
NlhuYv1qO0Yk/a7Xfh4P8KpYiSKDDa4cAWo23dWJSxNAMlgsQmSPJ/Ogj7zkjhuQpbrn+m8fy89U
IsWVcKBzqo7F/pdnHfOV7kyLddKH8Ku0Ob+WvaFR7Oe7eaRx54di/SKddPMR/FJsN5Vgjxqa6PSE
PqxEZ9v5NPPhkKiZn3mXMwGWtvXQSezQ0X06t31E616AQM2qu+nMHyOsGxtgFh7rBIE3jUZqij/o
GzstlCTKFigeyeARra+fky+VgywSLj6UMaGPDg0OkG6uzHbiNibxvMykSCNJpf6TKi3Z+lKY1iGD
nIdhvoo3hj1EP8wu/YkQyPR0XEBwO46xejNd70nLVi5VUYQ79X6tZKLl8O2d9++270VIRdyYpWGO
mONdOPflAjrL9KPbVGREpPsJTwCHGaSmh2BzEvtjQTHoj31fmoBlfr0+t9KdzmN+i/pIwHY1fmId
NuyicX4sCgjFWO2ED2yNWESXQ4ftkSjE1azE6g3Hw7NGTHtc29QYb2N/x2WvXx4ULVtoPOOJlMCQ
HG/qay4Vj3DVqhbCzKauwaWl806Ar+YU7ZCaGtSYVOIZDq8aVoYu2HmrBJOGtjJO5YZtrIzfn8iG
NG1Sis8FR9S9H0cwXBvK8c8MnR/ONN5QqdQ2v9PWBi1Y1sEV3RVUvQWU8bo3DS2NDd3VWjvVQjs9
v7v6m5xr7T0iZPVDl2AHJcuBMTIOptAml7ZmwIH+ezX8ci0xBx7LWRmGQHXIqgXlNU6TF/1oEmuJ
g8iGa/8gXUKbEJhINBSvSFMX+kjFlGv6hxAQjAFRHA7VuDeapqoTtkiA7WWcf7Xot6txfzOt4oZy
n1pMFMuO4AUCmQl9S7yKa/sKAWT/mbd6tYirbG4l9LNqBDBWh2SbDxSZH1i+2uCZPGxNj1eHr9rk
UGvr+cjxYRFUc8bUnUU3rMbwY8KjfRLcbP5QPq4SjiWMJU2HdhL7L/aDEt4VzGYMNhzWRUSEv92P
7G4loi7VVyI+k9Y+cpnzMjYNPIHg1zymdqD8t7ivFU2AKcJY3391OjWGbU4fvwXZT5PKauv/C/1g
fKLcSngBa/OvBRBmK7ujzcv6HhdRkfcWRHSXS1vXuWFyw7tqevzugTbrtWSS3WIoXCs7BM9qbfrj
tGZvcIiW6DaiwH55P2U12NboeydWSYjYzD7g7/abOAdUrA5TdHBzee5YtpIBomf7WZj1OAd5AQ+C
YrJdFt5ixXegAF8+tmxzfIvw/yhKLPd4vhe1vtNQC/GEHvTHJaIcfgAVXAG1wdW51NAGmcVvweif
aPQEi+GvHo7qtnWH+PO0jcbkJw7SxTxY/3XyQqWadmjo0U6iP6z/enSsbkj/xZABLAR9g/Ic6y3a
z73CdQMCoHdK6M+vRwtNqyHL8Qogje3BhuGOznG5wiOx1Uhj3LFAfaW8XymmMi7WgCTnEt1XOJeh
2noax7U4GNq4n9QgH5vFPm9PaMBSTeKj4zJoZ5cuXvxBbmGB4A2JhJKU8cHjdPkjO4nqHnDC6rYw
7dHs0si0yywZ6ubglibKV5GuJinnjlcFLQ4aKqfASIO4VISNey41X2kjcxTkKWOgOdxBKLJygdNN
sf8L//VzY3F3hMvVs5f0V2i+bar0ttsYU693lY3bouQA3v4gmGxduFAz/rbp3h4fbk+RuxC9nlbK
YUTAH23SrCU+7ND9v8uzlRBkkuApVSam9Brfht5QQAttCAmaLygbG3qMeUTiDnLliuMotiGD53QG
h1gcsQmcmm+2TitfdjaF20iSLPHq7oHMt3P/r9+Qs7dcqWKmS4DhbYJj3NEKDIaKxZS0nt/4KCKP
uNUe4uu/nAxVgsQMbfy0EddXmeY1Qa8/Opx3Aca1F4kPRYLEx35srVxHWge+CzahXtS5fZ+YRrrv
eAujxVt5VYLwxmfmiV6DB6ACtmaEUGwb/yAyp2LuLcjekMFbOXNZ80AtETM917O3MHaqCWf75Epk
MrLohOuimosYAVXEgBv86nLG2JuTGU5Y2WJRu34AZ88Fk0D24ImMXJUAf5wycBykdOAoNfvQwNBj
Rj+oOFSu/Hdyw9awY6EgHwtgZlQCO/X0y9HBl6gBV6iqIAlWcFW7ee9Kgf1aj393u0TPiID/ZLK5
5hx/WDHAi9V5ckswzfV0XOpS6TqN3IDcOWtEIzeVJyBMViJziyPG7n+8lY9SEd5A4rHijC7TTPPW
Xz2/SolW/dlu3ifGoQminPhy4ZVKIWNEMkgfm3WLVC+AscvNXcQrhyXYuGpBcY9zqGnJzjRA92y8
gvmzIQhtEfYg4yc6+Iu6pe2b7e0x8DBB2Cgyo6miFvCOI2O+QyojKRO8GX1ERC5XJzKhXqozcxcl
NeztCFK7n6lDe7pNR41G2pqrcp7Jv25Q/E2oS5rXuJogPXD0gyVE+YxiPKtomgK1haOpLRF0thVT
zRCDBz5opsf/f3Phpao6UDi/3YX5oHxZsITnMFbctfm3LhqG846kQhMquCbhE41fVf/tWZfClU8P
ruwpRKxYYqKvfs1Y0xDPsrOZDLIakUUvYRyZkdN/nhWwUhJW7jzDPb+6psnRg1+vBJLDXMqephHS
9ncQHpBnwUwqAvNfW1/YN0oZG8TbrdwENdsKPrlVvf2zzdiRWSjP5POooA2SaGjY6pudQwc6evvf
3GCi2l0Y98KQpr1pSk8h8xgb/3yfblxEHP0Wwnm3gZtp3zqC3TQ25eulmxIPYHqd9rYlnDQoLoY6
D5HVNMQ47j1U/oVcBmC7g+auInkWovBx0AAi+MnvsQWudyv/oso386tA/BRnWVMm2xQ8ky6x82li
gdFhWHlxNhYhZUHKnMw66Osj4Jf1ASDL+IzcuVoWZN/Abt6oVM/zq7QWKK0aaKTN6UJ1eXBAv98s
/5GDItzgpFZjO5no5ETcEZ8tpmhpn2Haln67tzB+oH0bRSHsoJGNfOHR+OFWhIOVlAn+knxSp/oY
gpyl9nc19MGxtGQ+tLSCnpn8eV2PViqhzSHz/bcEU7+LgL4hT8ZYpysIAg7Op8RqYPBrPjSz0Ads
74zYYBMLVg5i+L2pi6lY5EaMloS9gLszJsboHT9G3/6cmsyYveGFmuUvznhxUbnf/iiBEV3rIU0p
lQotEGiI15CyAGpirdVsue2ItTSx5rgUZMaEQyh8J04KgBJxJ72Zxz6GzdXIopm8wfdmxuuxP06q
YF8IwJqUWBKUFgM9XR661hS3xvNHPyrp2uX5pEa286q3Ex+OWjtow1jmXsnPtEhrOHxQS/9M5fIc
vUgdr9scc6fLmnWlZAIpHja7X9X1C20h0PKCjQy4m9PvcPxt6GTUsFkRjpO6tjFAmdT2RpGAgGqL
bCOeL2PrPLdgXwYB0X7PrBLDrhZlmkL48D5LuklatwwbtBazIUWYVKyByanReiDUGMb3ofRv6LVA
PD4PtUuya3XFO22QcpV7B5Xug+a316/ALx9IRoNO5yMUYsR/ilo/eTfTuMlT6Q6MVO1h6nNJalPR
MKifP3WVk8F3CVfBV4ux9B3AdsCiSKxbyAXz274kQGJ0rSgdMKowHYHOR+liHgIb5cT78m+vRUU6
ttPeD8pSM35FKbUeEj8HAO+6Dwp539Z6LlwKszyT/HjzUuVXzkDCInbC9j5olgYNDyiLaNJoUTKj
EHyOW1WLz3J+3hm2tPuvj2Pb9i7AtWDcgTN8zip1pxv6Q7vt69k71/ZzivhdvhZJWr0tw853m7FX
wK5nDOMLTNHFnSI3q+vPpQGZQa+N477QwefzNMVe2RuXCGAaHvBkYyLnY3iFlJa+wY0endO3P5NU
zQC2Bo5KjD3fUKDNEmdlhe+A0cdQQnRFuwzZ5XIcpuX1geJn+mZ3LT+ABa8+TliuHeowpsPl7Ymg
R/vfdQDvfwoGOeR5ngQqFheIoKx12his5thGBhMbbShlhvVp/Wu6KIHVxebRI4QAp7hCrstou74L
jjV/wFn0jh345StTasd6DVDUItAbxKslNcxxpmP3JXq//Gdk+I69uj1CxES/UiFY9DCAGuLcsZY5
SZFGEgSCcvAbt2PfIPqQPR3oUO6Bh3RoK+l8MFOb8qdextKvRbmKtWY1bjCxi7XFPN1lmLN6CTql
lWK6ZTFV9WglJ/m8zaIKVPSFSnslAzsP4js7QN+oXPtKOVCInnoIb6A9YnzCM/WUR3mX7i3LrA14
vW4i0bLSUTio0yCLpK1p4FuFEGbS8xFVZLjHc5V46DaYYidexR122NTSz+Xmq9F/fwzwIvgASD+5
sXAkvwXdkM4bLD5TKFUqn5c0NlFDd8BPPBPn/+XChOfZaDwXWEM59bFDcM31tzaDQXTYWp73cQpu
XObEIyTgZGXGzSW8lA+JimCnT0AXFtz+IrX5SuqusH/IYhJSEa6MvEDIWk7z4VnJzoAZEANgKXKs
myEGsG6je++o7FrENo3NIlTsRO34TrrF5W1JSwY+adGZB6AafclBzdDnyu+QwsaKth++R9+Se2Gw
x4iCByHabDuAuiyQuhaO+NAXfOFB61Yp6RvFF92TBB1OfxRzYVTgBZnyzJQFulmp8IX1QJzbq8M6
6gypVUJDNTgeg56w1sAG9EEyYL2k4cR0VKJCmeltP3e0qNooeQHK61ZvebWio/UbFZN74+mDMZwW
HioiUzCFX71uL8R6BZAYFwQzpmFl6wdUzRUH+tdz2vCKkSA7Wluhzt3LIfBFXVLu8e/HyFDMiNQF
DDTokDZGhOegJnvX5ny52jEgaJFPk0tJy4Anm0PsHih4T8kJx4SlAe/ze6HCmitAusW1V0NmTNEl
FMy+ZXTuEaVsYfoBV+uhLtkcmaeaEgmJa8YxeDA10tjINu/SvHgOn2hF0UwHva3z0pou1iwlNuvo
v8R+j9NmS6RXl+enZ1rrGOSFn7GKH3lSmxFhCLVWVvPdYoaoBkMvaKwlqeTSw1yTAvWPAzCXU6IV
kQYWcxskLkIysOapnO1htXiXc+ezPh3tmWCnJMGzlxVhL1OuFHmGzNs45AEL6xYzHtadYeEYuHZ5
D09Gw/KZr/Mri/wkgD56houzFzeVm+6jNSxdtHXHPTbrzwNfB473v5rUhT0dqzYI1WvWYP44dU4k
EG5XixOCPGwbtBJUIZP5Lk+pMTGtMjI/quhLbrPPOYTiaWIqxxFoj3sGzshbA/RAH6t9kPBe4w6g
U0J6EwbcxL12H3Wuyr7HXvd3Z0PToKUC2b0796xUmdZ7+wpC7KjKYPo9wtoQvJEexyXF1xjpQl+F
/eeNraFECDDYvAKjLKDxU1GU7Q/HxZvyXdBl27XKq8hSqZ6KFKETVsFTqqgqZEUZ50ktL5leBz4Z
3I8r34RS3328OPA2UJxPTosFDvMTd4b1V/EAhynTpThIaZw4vbPshYrZh7+76V0PvORRLWwpFj1t
pHLwwA5sn4HxwNmDS7XMi+v6L32asHkpFLcBVeSCIJIosfAJOKVMW0Wm2NiSO++COhPbAnk5K+YB
VKeg1Y4MOl37JAVOI6QivS/cnjroMkiWs4frXALGe+JLwbnJw4meTxCD4Db4gzNB/wLaw1ZA+F7J
4PghP+yu4RTBkDvTLkfPCtgY2JV4FwzNpAgaDzL4+yUohgGEpkaYYdRvXvW1k72z2czrjgU+errm
qJ/ISYFZz1ykIFfDMFf/IdOr2XbMC5GJOmxPqBLt0lme0P441SzWI41zl63jWFoAA8F6zQggP7ND
8q6m7mHjocqjp7MQceYTP/mc+RJ/1f4HQTua8o2ANgiLC0wFNGM3XDsvRsHW+51F5qxAQUu4cr64
VUpnFa6/XzbTRmPrsHq4EFlTqRVdovuf1HKNtm8Pb4XNlY0Q15+d7u4IFozLK7FoX7Pq7XJlO3HG
B0xq4sRAlSAUt6MsnSxTfJTpnljGaTlRKo/D/TeCfazQCdKExRv+rZyaqkP+CIn0SiR1AWkwRSjM
zQOXeCRfc9iVp+MAWg2zlK9DAD9bYxIoJ7r8CZJp58vTOd+/hF7jGuDudrHU/mCI/I842bVvRdFz
cIvxAzwy7w3v/0QudtN9bCULWJDcF/4x3iQcT82Bj9Ve2tlbzQAfrjlN8NPTbW5eWdY3aVlBtxNq
qC5vco5zKz35Am6ffacFuOehdhmvDwfzai9tVdeVvUaNf03sRqaeLEC+Rz3tmgrnYoXCWTtxGXNA
BY97gmqHyC7NA3g/L+2yZUvt1da0bLGWUyTNk1SdLUIHWkWcXyPRqMOk7SWFu5LTyNV2MzeTGS7Z
+Uvno5eDrQlhIuu0Cw7LGTn1QKalhoKQp1tOlTLSw7kX7596a66hgySL1ZAqhyPNPu0HaOHJOwKo
xyeCPmk0dJ2duF7T/KcjwiXMEetUizyFtrehozOsicbB/6zPVm+EAR4jMTZQEcHIVAFrr8isi543
IWsM8pD1bHteZA+X7t6Mu0gWSO5FmqR90CD9oL3qndTw61A9LnABDnFrf0xJ51rIUKkrJoaVDhLU
fAxKRHZ6CPoAMhco5Qt73HcOW7ZjBaJoMPjKM+vDRnA5yIF7sKHkA2hbxFcs4TpkOxuFMvlJeYAh
xti9zHlIteZQlDsFkrBkU4d8M9LJoOAxXqykNdl07DHEE4umg9NNoCcJqgxp6rVscblzNjKquUSj
aA+gkaddFjuzXHXl+QN14dZU+0XTe8TDxx4W+RBnv20rEdyDSDJGBFabFARqZDw3KD18SdldnsOk
FLqLc6hKAQwnVsp6sSMf2x8s/a8ka4erVrg6i2sb15ONwNLXQs8Q/X0DFD5UL4bsW+D3s99zrzFm
WdodBEDd0JtQ5sCmrjVDNj0PZUUgRc17L0eVmRTikJlLP8BW0ACiNBW3DLnI/NIpbTFF6ZFx+5tt
OsssnfwUBiX5PKHz6OJsue34vAhFN+i7uKaKr3RZ/xSOIBVd2tE9jL+fSMRwdssZKcIZ/MKGbqs1
t6ltXeDcCApqQV8u4GPbqMy0nhAIO/IG/adIJvVq/gRw9/9mlo1BUSqqr30OC1/olEJX+3aXcTZg
xb/v4h5i1TQTqYCf4hyeYiO2Om9ihP3CXRTQWTsDwRaJi03X4LCZy9yBa1OTZlcC3Tx9ahwcD72E
Wr0IJDAMfl+Cn55zlTPjoW8DBaz0enMJuz57/AvG86FTht9OQr+G9+Asyh7LWFAyTvscDdwWBLmN
f2TfjVxG6vCEG69JLB4WqbqMdNsZ+mfdkjkgPWcLtISoGHAkvZWRZb7MynqeTS9skPQDkBAbNUkc
QYJsmDtWrpF5hoBRdHDSEeBLlG35Oin7NguhbixAb4f/TjoPEFV8zYCWyaVIaNSrF6V1tSVYdAcQ
8qjFw8gS5Z8OEIiHYKrK+mF2ERiBnCK6doDRh9eq6hffYWZJawRbf8zZNd0vRxls1JKap+dpNgBD
VTEijNbB0hC69L0ml70IZvZ+MCzaDKf1kAV9cqIc5RF+8xiEzK1Ttq47MWVpKacSv8bek71wnCVA
y6af/+ntIpcEC/D9D4XJjbglWtTKUaizYfPFlid6PEjC76eGFu8Ew6TKMsImstdQJ0vmDDyePMo6
YR7TttxJVyPNjCdnPakdJavtY/NMFf35rnzDHo/a8JoqywvbABcioh/Sn1ZVknbJYLWa3kc87j5P
WtIcutzf7B1IBYHlLNBW1i3EoJzuIkoSqkp06Hhq6VEE0/1AB4bpZM2WwHKUPsrA64sYJmuX8Ppl
a2u3ii8PeJ4eLE8Cw3xyC41BqqlmWxSmcnSakeieR/2H9LL52X5SntU0o9SDQwhTnRtsxydxS+iN
OMzf4cXA6SpnJtq3FJSjqq53n32Q4Nd8F3YouQW5VVRcwTQ+tBXW7UVCtSVaVmUmXUv0gu2d/RPU
d3v2d6G1QvPj360L805jSsOejgynlHfy3xW01IxSDHawbd3GzL7E0zDXvVnnrqnjSqQD7+5FMV2l
S549vp/DuOvzL3DtI2+6eyDdK4zo4uVIypPURbu3mcPidrDRUnL63IvZtkbttb8WI+9hDNCJ6mVr
1gtJninGW6PD7QZJUU0HMWcX2w2OoS+jbu7Uep9yVKCppTGnHclbBr4/inmZux8CIphz0eiVgwA1
NXMKa1nRMPgBZ9C5P5XCe2QuCTH2q3lSQUzTwUPLYg7Y3dQmyUfQjzkyOHFqLJCjjbdDWMlYYMVY
/l6BoVRNzzsg1+HeRje2VjD6VkaEmKJbaoG6riEWAgrp7/mt5+J1+vgPDcoDo+gQmvjwvZBVaCVn
o9aeF82o6yT7qbnYK+bHpbHh8FsORQfv4gRTDeqg6LOLoEgDPwO8qbmJXlAyGxqX5fJZiyLakbC2
oHLz80NvcnwaTagPHfarEqEm81PwibwA2DeuNj4KLgp3+3YmARJcmaJ3XJJQW1bU9H1m6mcLXlAm
TyOk4JVbJuqcnQn4OltR92GWSK8yu+wuNcD7D/GQlaAJWN3JY1j0QRNw2qLWwHuDdlEYQW14vUuI
wkWyaVa+MpGwxPWY9SqyS5/WoEisdH5jGRdsFOLQQAvqd+z0EPuEuRaweQg8iXhu76jL4V8dsvgM
y/kZMm7cO6woMB02qDyUsdQ2+HNKjzJoT9U+fvlebXuCZdijQiHKU9nDVbu/yTxXlJJwvpzmvo7w
Qsyk6/ookwNTdulea1On/VNJBms9H2phwpPPYQNH0Fun9GMqLa2Fx0rEdVFUjNlAccTtVwgpNMxJ
lRbwgEw3CXNmVr9rVODuAxDCyF6J5/wULhyK7ae3qjoAFlI0kyEQMDjYogV+qalCIWe9CUGw7ins
FbrECRtnz86tALJZZxcAcpxxRLMKzIVeAd1bbYEnjiK+rmYXuEIDWOBwUsxqk/hTWLD+QUCnj5X2
gHHwIyo+9ZbfM1mJpJMY1lv3d3GsVF2M7R0mp5KyfaDcJpBdEduy662cuVZMu1XWfrOwtNn3xx2W
Fub/rjhAuojHsfOq6TCe7tKG3aG+W7M/eYHqgolL8c9ihaL+rLZtIJm6H3Vq0dERBN1en0Cvu8qh
QQRcYuY4sXoH0KtyIFJX5Q+5CsrSnsWk07CBDb9dUS5R5tWxzt/9xYapC6l/7rpCwmLeUHJTyQej
G1/SR220ue4tr0Ru4LV3KIJcHixohryvji9MtAEy+FN6TqoLb3k4NRL7D4iWSYWXT+SWaGFw6omr
SH0RZFwlQ+C9isT0AkpAXI1QhYY9QWKHuyFFkOQt931TcCmPxL9QbSY+H0u9jVzvHoMocSkAXiDD
hevYGlPurcE14tPMTU5c403kwihpm5+HrnrwGkZTQnU0zUlNKpZOT0MIDZpqzMk3isZrcAAyokVj
QCh3fhoS46ShRaDyRbky/OXjIkRWwpNcd4EZmHGqrhR/eJ9wbBDWLOUZ3Bnnbkqofx5p28gJak6j
s+Gg7MHyo5VaPoqYEhsQ1+a8I1Mx2a/uvcSNnXCyH8IE3pnUH8zteq6lz8xCL3pziEwhPATqkY4A
jQif/8evTznYT8pPy0uwQP234aGZKsXwbObwtAz3x7Z9SpZYFDaeGEtvrCM1mxYKuC6wbuRhAUXn
Vx7XyeEZkzFBkC9LHa8Ccf8FhXpOSQNRCDtPpvqst+Ix+RAPY38FkuxxmHtcQufRXomR0B9PMozE
cOsShruYtMVa5WZgwSby/nSGKlZnTN80tRCJWiPn4Kw8OBVUZqWc5Chi5ENwuAWpgin4jszcblNA
Fj1CsR6MhzbewjyPFX1jMHYyy7CJ3ZqS84hJdyhWWeROfSFLVgKnj6NzjJ8K09uV11rrbfpXlHSE
Z8CkRSsj0YzfNJ8Zcsbt5u24EgLt7AVrEe5B4faT7tBQ37u3a8FKiDm85mPC4ZzH86SN54IEdILr
5ucoXNPkrEWpCcckra5/rtSPpxYDrhCgn8vM+KtSwzlS+ueUtlgsIyXk6o4iVzuWrv/r/tR/Z7yg
IMEWPDwSVZNI+iq5tPzZETCWpNs3EdNR5HVTe0BNX0ovhHzlOk/lM0d7dOpLg8ukCsALk9jyub+s
BLAf13A3+QK6Am7wp9VSyOAaNbgOhCHScWtDR+eP6UvZWM4cM+WwOaibYwopMYn2sOVwnGXkbcwG
jVYXl7A7O6jnQPo0vXUtt0PyOzJQQClyD+9Kr/J6EkYceEMncuR5rQGKXD/zMRt6sjcEe5/3QsL5
Eh2LjVIf5M4QXVmlzPIOKzZoFN0ifuH3wWg4QtRll/1mFrH/C90jSchhigDsw+afcTJzWQkkS0n2
ZicrlIk9dA40+HZ/XwXcBckmOYTqO+PAO/Jn5ycMEeuDoZedfD8/XzWwXtrzG4ZlGgfEDMi4Zuz2
Wjzbd5KjPAiSDMynMWOxG7tmlUzjpyRCkOsSSJQ+0g6dWYQ6OKnvzMhu/3qQJ3mXM8orjgrDnsWb
nnXgDOA9hdUoBd3o/Duy7NRklkhaJC96ihiSXdtlWIfT3P4p4nqyN2knYZw2eQAcXs+kv3GQUTWo
DheU3i1W2p7w7i6gZ1kwDLMbnsUVouQP1yHiwG32tkqDEe3IW+0j1T48V+UBU2Fu5BgIpN6NGFW0
Ec9b8phALfNyPanMkPC1YuElppBMmL2ULKbBiI1R4KHVeSbOHCLkj75ZDQosU/utNPqRJlT7vK4H
lXtcTi+sKLOrseNSWCtOoPwZZpb7N+kpovPbuJJDLOaW5OZOz7dtaLBlGNDTI+zg8mIDdh4fdWjx
ju7fKOp7ItLyCIK0QWR2IVCHM0hlZzhwwLYXpHZ9cQ2YVSnmFn9lqDiU8ZwFgGOA2c91ktPDO6RY
AnZwlSpwWMhg1XkhxsiNiHRMLdmapd/9eGYEIYh9bxHihltGmcrbG+Sm3X+dVaqjhcnGww+PUv1w
0WjV5faZ7Uv0kIaprpSZxZ2pw7+zMiIh6gl3328ZvWxscAtIAv31qbtzW8pXv7+Fqk5oNgP8tb3s
nf+XeReRpMggVR2sY1TQqECRY7m9Vk9ygcNpwD2M3qRBPBwcOOu/+43NYogkAAzBmqgeF9Ll12+v
TbujywEmuwj0OyydkxVKdJcofZs8f1Wx4meTFNEmhPTmEUEEh1pvjnxFK6c8wVmrfxnfEIcMjggp
3ihrJws8q3Rzvr95+Esii2ChRhYmqJEjZ2BBDDnAKYUzk7aaLZlnIO/Dflzo8q5VWvoIXx1cXbgU
Hxy5NtH/QtHpl6ujYuFG8Q0Px0YjS4ejB0NVjcjMYAp/nXzxoQcRFS4E6ADMDWLehYo01rxghqKS
SdiqpuXu258e/YlwlyNFodUyRABivjRhxuldyKt43X0G23kGrZHq6bXyAN9urs9lScCsKHTR96Rx
7ycEXwNiFsCsQQ7B9pXujeXhOMmgcoeKM8pK0bOEuAqSsfbXM0GNubu+lFCfNgOtI557G0CAUqCD
EGFhnG+y5aBdYv8bVNIdAyXrxPgDkcLtupLhmkAyzVSgowZacA+HcNd75Qgl2dMzEBZZmLsmuPZ2
0nxedl0Z0kvn/4Vy2Y9X/9nSpIw4VzC0kMcGVbbgv7Auq9tP62kmaRSs2DZtJ9IqjzdTYKBt0IaS
ONICifC9Ur/eG7duzZUWmQMuzQW3mGB4r4M9i66mTpeXM06dU0cobiPajMp6WVQ7u3Ew5LMW1pmx
1B1K1EPe3qoywTr/iIS7wIB32xfqLX60sljCct6uGwNoIiFEyBkAAHC0qcqiWJugbDmKkQCZto46
LuYAlLOV5vyq8QvUL6nEKP4xm0Qn2Y87gqq2Ec74zM2i6i7cLH5amC8Xa8VjbgPI9iYeddjbJc6t
vWL/r7RkrBI0PBZ1HWgG21TtJdhnnw82gUM0arvWDle5f/xt9SZVla2RGcnQNAQlM1zmTizPe56T
fnAf3+ptbNBppndYOU0JT9ZF+ykib8S1NehsOxRTHw5DsDM/hX+BSwZ30LVOJ7Fld4WZR37DtI5m
qPECBwEjORTCoab2bMofXMHErLabPntE80drhN7LpTJ2kmUnL5iFX7rHD3kmlSDJKH2lBKNKiRHL
vGSSRojBQQjx6HGd6TeN2kmLQpXcCsN4rO5GMKYJVFcnwnU/5/xAEIIfemY9OcYjAaFDksWXNpuX
8sU3lZHHzKyz0irzWF1mf2VeuZUNoqlXUZVs1UOZMfdYlJWd9Wzx363TIX8R9waXOdqCTcgfnLEy
QSXGlWYqigJyYvplaAzlYuUftQUNxRzzfc7P+6GpWvBuz1I6JbjtgT/9EPSoaot4etasIBKFrnuA
xNyC3/W83n0/YkwFlkgMFb4Zig4QcopZEWnBStwqEMXgeDE2yqdFRs+fifhhW+xqDizyMilc4HBC
6q6f/hZQY7DbfZuq+/Vq7JuZyaQbQ//lBSapVJamj8WZnFbDK9LXMCftAIgVIaYE+AOGCvxJ+MWb
ihQE1i1nnB0t4u1KTRwnC/iKmAxTpo4TeizfjxBh7glLGhZqm0GHVJUqnUwPp58oRZQHObK07ivV
nU4Prfu4rYRT4rVK7v9RqfC9In7gH/gzBzJmmqSFS0G/+jaKPESR09VyfIyAbUkElHk8F6LPXezm
yevO9QquyPRIyhRfOzhdF09++50BQXD1Ac+mqTSFXRiB1nK6AzNLQV3mcr5s9acf2Ib43+f9Szuv
TmUp9TbF63u+9ZiuVQeGTp9jstcE+PUCRxO+aqaEocmPYobCEpXTHx+nHKWFja1C0axbkFyvIfwz
QjYE0c0UJYiDZSN5dE+vnsgPQcIIFJkDFkz71BId4xps34o1FDjZXSwGAZIrjnvCfBvWpoL6we1z
YizhBWkvZf+xv9VGXv4paydukbBNRYkbk/ln7tmLL7gOAz3r4eg03Wi/zJUf/6/uMqeGcEBU0ozc
OQypeFEcJy6rGzt7LeUU/4X8wKlLe6eNRpztQoS09UMbzy2v/lp2pZ8LVJU50lnJlK5UZK+gDh5J
U5Xwc3uQNR2lk4QyB4lTcLadZeukRGrOV6JfAovWz+XUKRBUUh3SXvAJnLpqSBeJWxatYsJx4/h7
yoG6aoabT3QE5VGYxWZqdg5GBOMqlO+7ptYMoCdmkNlB8artGzsSRw8upbkec7LwlE5bLzQcFnbm
ALI2qkE0R5kLetO7t+e1SZLdSlAdei5Mc/rH8lCdzJx+KePXhwrN3lfw8P2cqWa/T7DVUU2yNPo0
joil2B7ZgdD9g8nORLb766s5rXOdbh0rwlR8p4JqpHwdUJOsaHXqMv+viGJCvtyfWScI1O6TlGzt
KBtss7V6y4Ps9GgvhsIqaOIdIGjDBQVFrNsLC5Zz4Zw1UWgLblxTrCWjLLHCtxjL9pXdPAcgTKFW
f3RRbT6Ok2DF1+opE33h+j/mmKNtOZk0a6Pco0A/udl0ZopKvm3/wNJDJ2eyuYgwjEWO6B2gZ5YJ
rgdPVwaQishpQr8/R9muv33WgmGiu3Bzth8JyxCXqk3vwI+rXyd0zvl+GFsJjsqhHWO+4EaK0hFR
e6HKFsXAlWB9Hq/OkBkkVygyOebOOJdire5Uy/fuEXNC3rrt34P4A5xGyB+TEo+UZwBZEmhNxPEi
MDd2lxgwJ2zhdXtX/Rvle2vdy5+OEA38GQXl8V/DXGDDbni78FMQOy7UyVB9ENM9J9uBxrHL20+V
vDvl3VXY9P+I+N7HZ/lze55qFywKnDMRqNAOm5hxdlkWoDTbeOAykmTn6sM8TWUITbI0OWdMwjv4
xPOU6yb4Jfk75mbpqFc5a/hNNdTRrPWTMCkA+WH49sw7neesgPHl4LeX0/NBC4y987z4clqSSU/m
4rHl3SaPNHSXettwV0g0rzubJydqvaPS+2LuJfztksXSs7XsIjdyFvFOZXuPF7JJJYg2sjgZPgCv
PFGzugo2/zUJKY0nfh7vRjrsE8uywhHfraLacyAqT8IPUuWMcwR8rW8bl7J3Sl/O7J6UZarrQ8hm
QtWuj4AfZIiwlX6fFnEaUN3b8QP71iGH7TB+xlJbs9Tuv37/G4X8acirOZlqb8zukh7UPugXfLyr
+QIWA39OkyjA6bEaM94mvobBiS2Ynvr0oPGcs201MaeNJViN6Cn8PBrGalDh+wCk5SPMf1KE9fyz
KxMir1WDj89aopAQgVSXvCQ54zHCUQbIE7C5zj3zo1LT2YAjcSRmasTiyW1Ftw1I6sK0BY6L2zOr
3KN4wfK4KKOwxky8fD88eWNloEkh38vrsvqtiEqycGqrqRl2meiG6NVdjQS1AlgSMhZIPAJJJ5+h
5vRDHVZu/ELeHntV1QMwkXC1zLV006h5EnkT+1lrg+bhfpH4THbr3Xq36nFO6FEeE2BENHhLq8P1
U/PWwo88ywkVEQMPe9JAbop6vMGQQM8cnqUKnW/Bf3AJzwaOfbiBtUhwS91IHrI9c23thXVQpuLa
0DgiwaoeyZBu603RvjJTi5Y5U+uytBBcftG/RPo/5/7DharwvMF+KyX8twYrnq06TLzibfcYmevy
W544R2wvloyHaEp2Bjt48tK+lKSqJbtm2qkRwW8QJpXe8VM6L7WCuwjTl7bvNHMLwuFlFxX6gYbh
lMghfhhEEY3O/eGlTOfJjMFJ0KPwFnBV6MEmtY1veAWGtrrBUv8kqwSZU8Ev1vbRwc8LgIuDqjIS
6t48X+XyPVq0D/RR2KZGjXGcfaDvb7e7500ugS+RXGzo1VEwHy6Ac2CE3QA96uTpys6rcaFaPTwU
rFP3KPgFRb9DDHrb3Jq8vrP33NUkJV2QFiBzy8ejmMzqw/RupydFmh8Tb5kyTuvD8ZXGhZd2/bMc
5UuSyJZj0KImPLGU8hvmjpotZtwrSRA0SYw1ACqE37Rqka55i1bojsYpZS5uNB7BvpTHnH7N4CXs
LPB0d156jlYC1reBq3aDY1zMceBxWZP8TzPS+DzPBl2SwDZWgrAyEjuonN3kJN+DxQenFhcZjj3G
SdgDYBz6dndbK1QNI1CK3T1qXWGlpC4uSA4Khpyw6YalyN4OtbHRrFwQ6DW58kuz3n/n1rUVLa/T
aNy2UQPK4PiYgK1n56S0N4qqjezIcCCJo/EkPM8k3H/UoxusMj5sRK0xjwlbvrwE1077vzfElSRS
wRVU+cspSxipxWpzvwz2PKy1GhHkJ84z9fkTzjKyREs05nYmi6geidkenImY38L8twaJo8XO+dH/
BUK5CGNzIKXFN2yandOXYXuJjG+Fu+foGpxbl/J4hORPh0pk6n5zOxXNaPIGU8t1XJAwUbIobMKM
OJwaZhgMzONqzbPt1NIoG7QThJKdNXSTTkM5mgMYAiZ11zHws5tsKIC7QWooEN6a71z6TWUFBy0J
Elr4D9aeGLF2oUgmrNscxF3W4aaE70mbjXdHawtglyjH9K9tNxZbwJ3+LO/5p6yqhLVMhXPzAdpL
AQlBH9UWmuFVniEkdiLMSBtuEVyC5/BAjyi8oPEQxbt4fMjrTyruZQBJ2j1OvypJtBrsVB4RPbqT
VfGkrriA+yNBRVtF272PILbMm8mGv7zsxsObSTS9inY9Ynur9tyQXYSSLqlsxoTpIasA1rzAmYW3
wnk/wuJZypwWG8xiiTh5rJQSqirL9TDyZhIVquwLQbEkBjUp+EF54Tz4Xo83FybKeGZ6pmF2vPDb
MHgRa+xq4nj/RIF/Ay1In8MZ5aK8t2ULIt+XOobIbI/vJtQEukQ0nA57uTJOSBZuk1w9xU/M6PYi
6CmOB2HHKBY6VNa4OeDuD6+lXwT7X+Zk5LwEq/flDWGUQ8rAGtci782hNZIwQz4Aum+kAW96UsG+
s3ui7hj1wNHy7ACxPbfu1vSlrfkPxSHlQ3ZxYZLSHM2AqKHaT008L/WuL7KBzonxcBoR/RrG6C9G
+UkV28IAGW8GLQPcgcQyPsRaQH8zR7Y0rWH5hOHKLlW5qyjhxi1gTwpGam4ICbTSJCjnMiKKUafA
bYKNsfp/EMaUA6qoE7luHIl9nlT5nH6VVuEdWJwQfKiwaUs+yMIxT2Y5QSL4ttqBtIUCFR5FaF2K
ybjiJpufK4r6smqrIIC0cN6HFD7EBQTmGatAm2z06tgrKm0Q65+IDs26qTUlSK+oq1MEY6FT4od/
LmpibSdCdIktFt4Sij61eje38YB7ijmFVW94bzgqF5iCYG+uHcyTRQE6mB7DvETZmv2/5gLmPMeF
lySGP2UiGMNVxqs5fkGL1PksinjbNL6eBeQAjXCILteBExucbCCRh/GR1j+SzAPR9/Yes0nPZ9sU
xB18kkpY4dTWg9H/49fIqx1gSSC4tCZNz5tT6vryFevV2WfejN2uxFQ52dPiZNZ249CHNVqBtJEE
O3B6dtgDhF6G5DdhmWzKPVKDsNUw7H0K53HnZc0DER99Hc8BDZOKNcNXYlbLorNPG4BdksJ3r/0I
qmCTe8WDm5J5AL03E1JPXpWJDLg0t3eg44S50Dx2LJKOtQu8s91j3SQqDtqpL/pa8bZyvr0FdV5q
cQb2M/7c9FBEadsBsJkKv67H3YGlmtOR4jo5xaDERU/8e284HSXbcINRMpRiBsGst8tmY1VtILCK
8Kc++yBHy1nk7VJNV/wTlOcoGaQJ4aYrM4nxNB0jKcoRfZuvPgCQTNwDvCFJBXD7SPi3Y0KFqwRm
g/+kVtXKMJS7Nx36yujf6JJ1JXokwQ6ZNiowPi+xw8600VrACMTj1YjVpm9+050pt/Ylj4XgbTTD
qEVqaSbJUP84fqrjlOVF/qqn34kR3BV/a2V1OfPaT4P69He7ptF6fFp0U2of9Kaj6YvzzLdigXuZ
o5/CqN8NevZdYq5zYukWt1b8zG5D+z0MTQp4FXdCfx+9E0kkm691OpS5F9Zv8JkSYUcilJ996lJz
Rdwu8sRq23yd9KLnGfunZ4Kc2AuaGoY49yfqsPHtiO0/wFii1ex5C2oC8HQojD3En4xh1rvfjnku
fsoIaPB/Lt7/gPZnLOF+pyVUj7Vt69FKZvfuMSDWZpUU4K41OfBNunT13O6q+p+WdsdUkMKvAiFN
/yh5+9iEY8+oMryZzSJJWwsWxF6aJpojJNpg710T5OYR3NPIrpr8anLKcsw8/Gol5A5AhKKV62Pq
9+CoMgd0sUaFtJOkeIdzRJGpOwJZTU982kv73H0ckB2oLmFXtUqPdqmrwhtoRFu+u4cRZSnFmkdZ
fBvhgxD3yB3v0k/S2/cRCBPo97kRUhFl6T82iWYtucrsE+8uCsImAF7B4LDFc1LO7EhrqncIYQZ2
UnvPRb7sRjtndCiXZweSvfQGoiZ1fsU8QrN2dwECzH+4mpEt1z2hkAgQmfXaaOfvDCrcnbCAqC0k
46KFqNQW2ANd/gGQzA4BSjG4ZNnsyN1vXMMv65mvifnAVpSSeoOgwjlpnRQgjbRMVOfypfvnOv0o
Tb8zjhq6SDb3qnEvKESu9lzPxBA+QkpVHElqaqK9YDbVSIgIa3o1bj5RTyx+yddeRuLkX8mbkel7
xLj7C0O09SVjwTuA4eut1LYZzJXYJ9VUCSK7dj5849Yl/+7rF2xzNmOVR8EUa3bGOABvj9hmUPHl
hmi94kOwnqhwoACfK8d+lCS/rxCuLrO3oqiG8V7kFUNeEh00l89KzT3vkm+Doh5ZwQomp1BaZDz0
OpOp6oTq8kx0vuxlP5C/dIImolr/+IUlR7FTcmmWy4wqxb5hF453owokbVQycLYwOl5vk+hqNQWK
4Cu1iVpn4IQHOqBCPBtwlD8lpWg/c037rDClnNqugJSnopGHutN4nDCYGMo/ACRj88W6r4lKSL+H
1i+fZ0Ob/NoJpi+ZCj093xVsB8Z0n+DYcZ/j68FiJqHvDG4iBxGEZ/LuN8yBYEDlBaxcsOlJNJEC
mhRUhNeGVnDTDhJ4RMeGfnFiLh4jSI2fSiE3MbVv9t8zU8l5ai0MCyOemFHNg5RbSowQh6kum97U
ZyIGdhFgGcQQFs0rSINbIgEwz7ZT6AaykodiLqrcSrFmkmG5k5bH5vx0qA4NeShD7zh47rFRZ/yN
3qAHCCYJJgC7VYV5XhnPktfmslvhe5Iu+Z4PaWKn0oLYCjuEbvgBhMbI/qJ+CrqS+jEikDUbUl1T
2GyQagLJlvb+5IcrHqLEX0Eu/5y50uUzQLESulhJvk1w5uPWb5GmSN4dCUP19xNPd2uo3FmMLoOa
DBnreM+hNZXIEDCzYIRZQ2WM2me4l/OXdWx9KLFf8vog/47f+7mfmHZo6OsKhnMEDIHol43uVcMQ
WemZRoqfyNRsdzKc8INmTqtNjb4an24kHFf6QecaTbrMKelpK6PBU/cOeh5LP2QZqHSM2Kmph35O
fij5r37GHLeD+tgoI/6X9tmXizO9eDmXj02aQ17vO4fAF18GqH4/qMyC6YpUS+wllOJ8omMVBYE4
0DLHYRcqvnhjdLCBRD2KBWVD+wSTkRqv5/T58dczRavfq4K0vT+x1R1o6B0POE/yrw0RZwTsOcan
vzTt8EuTJUkQCObyK6/5JVUuZ7F6PPs7aGiGW8J4xvpOIuw5EAdQSLRd+dCme8gws/+X+EUhqrRh
ywbNKS68Zhqaf+aats6nfZpnME/DTdqfVopyLf2c2Kk4gJKnU5bytCh3HjKI78NsKRZQXJskd9CE
eZqHYtWZWn4FxYBmHVv+b280Af6XwD7PB0WAdxQ/PgJEmDqQ+XTxngCINOCen4XwZv1UvNrL8EDk
QAX0BnTpy5r9UOPPr3eW5t4ArqtFbdL9n8yEkdRoeEdaH5odV7DnAkIKW90hqDgEX6n3yrjaDTI3
jgVsO+FmxCURKXHdh44XEeN93Q2QlyHbjoTFBXhBBoXHfbLd6xON28PxhGD9r1aNNWw3i8WzxKlZ
BTien9wP0n5jWvlvgEdpj8/MlaFTwhd6SxtPZN3RvaSpJDWu7wN2/CkseDV29lbkkNcMGihAFPyd
jrEovy+8ysqyhQAlXNNR4FLH77JrZRBvIZk/BzDlLOksTLLZ0ODY822RmFOrPdwsUCJe7GG4wmLs
TWPtSBfL7DSZ+EXN3p3jtVAyM3j/vhH9U5w85j147vwmc2jMf6iLtXKZrDuui5zp5v5IpYmeQ4NQ
2wxG4Aznjrt45oIpcZPLn8Q/pjC+3xBdL65l8NqFGNFH150j0uArzA2qQhx0cskk+yhhLONCmf95
5LSdnGnROCjnm+GXNGNgcOW/5aTDRW7qCQqjz3e5Mq5182rw38HnDpthRto6hyK9r/2Tb1EaBHZB
jwXHNrnC+k1uvzhEzoj7eUXzU1YGsme89/gocsW8UZ2x7BvjtaBjUiaY7F0Eb7+2RaF44oPrS6Q2
XEakdp1mNpzwiDaiU0abrtUB0kJdKtTN8pycuQ8lXTL2f6v6KR3r7g5Z6go6l4BG96MQMh+e1fY+
QbkMlrh96F0Rj8R3xa/J71x6F7wD7BSvTYi5IZFygYJ7g3w9qm+2It4rsrmUUwUvlBw+xbTn3zUf
DAlluZZvLxIAQuwuDA0gG/wHPSB+pLwASgE+hctm2nNYz4Kuwq6LLr0KFLGudQw8tdTyGcwEqc0h
9zqqrUPYxk2Ze0K5L8Zu8UNItE4ah3mTMa9tVGzIkC7Svx+JsbriV+dFPfYO8SucfFrWThIyUviH
bdStu+NJ6rygptJeu8jMOcWAhYkJRqDhY63acEsL5IX+FRp1bdgv7sQ9eZi/km69I8ccYd7yc1T1
d/nm6Gh+7YcB14lEjNOwjyhKoO5SAWU/44IdafzOpwyCOPWapY+E8PeXPJcisYJMLqaPhjCiUl8g
dJNdA2eiGR06A7xqPTPWYZapQE1HrjriacQr+e7RN0HwMhZd+ganyUMLwf56Saif2pCK299/jqfW
s1JoV0W4K5HxdDUFdJMAi8tm05AJdj7PeakXHdL9iC+KndDmsu5NKMx4y0syOxZDehImzGOIH8Oq
N4ZVGpqmpxSEIulqYgpjSqGPKmFmJxFX97dx59h9+Du79gRz+Z5cM/L917vr1rWFB8y+eGEt6Q25
6VvfVgmmNVGekyzFjdGhnq6R8BYLZo96yP/ZhLzt+rbULld25ptrTG59JLnTX+RsaVRgxESzoMdS
UWqhxYbCvI/TFS0/O1jjEPvh9e6lulp/AG3ivCtTjl0NWeR4xDdUFF1ySO6BJk4YsZglhMHByKrf
NIVtNxGz+pqzf29UyaU7XoX5oH7uHT9UObGzxST2MjOCCXWltEn6tf+N3b3LrtWZZFSXAzZk3OIB
qYGsVtuhQTLSVqOZaw3HoAqvw6a8SZyouPlgVCBI6hdpJRf8yWQFg0d7LcPZZXiQZ+fd1bcz9snv
7hx4X56Q7dtKKlcmch0g3cgvvHVI8+1+rqdIVOYxtXPvv16adh15KVXNiEPyYsJz3N/Y65dkz02t
CYbBMIvpfq06kivJF3R20xDJDPugAA5gJuTGWSJlvFzPTiA8dzCDHdOKUJrp0FGIuayk7rQz2qBC
Whfp+/KnNN/w9lLDEFDmLv3PgrLZ2xXS2I48OfSzeYyjU0aDbDZtXUjQWlqKNoifLA9j+WFCXaHs
VUkOvuMd2NAnxwBsp9bT/ZofHdywJqfnh1vx1n+es6clQOl9qf4nrXc+zJ2LBUgdj5sR4whkm48I
PGxuXgHsw+r2XHFCY4czgm2Ej1BwAxDPZHyk/gs6BZFqaKj0UTMTZv8h/TM7d5HIdAYAw/XGp8Up
OxqXNR+IFUYB9nk6pWLUoKGv8tWSonrW+fY0XG7h0qwaM338pdkCBM4NzCfk6Z1ksvpDyZpsr7mH
YXMKSCG8KsShOATvFeKZZ0YUNpksb6062j/zeBuqTckLnEocC6BMT1e1C1ARuFkgoBGwltbTNjtA
Oh7vodhK3t7ZtHj5EtHEZPU72EBWJye9ORj106rJTuAV6TS7OWkm633O4P3fappopgPY7RhDuKrq
4+eT7YloOOoaSMjgRebXpCztSNqvOF3APRj4kSF7+nQPNSZ/vX670DDbfGmNpEfax3XMpeMTO9jR
mWG4k1XvmEB/FiyJvUWebp20iOzFBo+jYgTm0/3dC45TnbS08xikrbadJw1i+uw9YmyBvyFEePlN
43SWGC9/TK99dBfdmJyy2+XHs4mloW5Vkx71D7Tn292/VEjwXRFmvTdzcX5zhwJ+AQoUB+XL4vbW
L14ELvq1axGANYk8Taocx7sK8hssEL0LAzEJgt0WDIe5Seit1mmHMtg4dB4htw635s8mDZbNcT23
8CRA/O5LS2f7tmlHCTPg+adL23fkrnRX9RzNdRU6+CSx6iBwJbfPxQ845DdnL2ZhMaVIYNdTlI12
7zAtQT9KXUQk1yoZoTHnG5rgdKR+xNnnY36TMEO6SWWfokHQLcoOrDxMMnBbSJfeS3oL9c9twhCS
tkA0Yr+Plt4InV5yf304JEA26InjVHFtK916O5xcmWdSB/oWDislCHTeFzFHl9UI4XTQcq0rL5fZ
alIpCquDCMKKPyYZTEbYDaDAWMiz3sKWzkjVFeQh3G2+9LgNWmJROFAd2o2x6K0/cZG3vRylTbpr
P5RnbzJe2mCTGX/dhJYb7kBdQkYOFvlipD07ksf0UlWZvFRY/QXcesj5t99CPUFbgqg6BE7J/CeP
AA8m7ldOAVo/7A0jUlUibsittEvmCzdn2LamUZYG/PdJ3Xwlaa8vF/Q0VvNxFplTngktELKdbQpK
e8JJqJtoN5GZH8g5K0cOfftY/jNBKQrTyX2YFlaaTbUBQEDkY2w3knWYJ5rg8lTioKhm670uCL32
zCLREkaGX6lEBvcum989Wd4dsTzm22LTDK2UVizcnJHcdy+vd+K2f1VymjKgZNL6OEhK+1V0B+VI
LdT7d1vb8yQm4qzYJ9pIVBECIfZWIFaGgqpscvXLjqJA5/h/POem6tKqCofNKiR6ELvch+tk6Okd
hnk4Cr/yOkcxADNH20CsyKESOVi03LrjDmBnPyEZQVwhYQUjT67GXUMDnQU0he/+auTzgahehy21
fRzm4K2zxznZnmFLJyxn/46VhRi6jisPFlvDdwyKzaw3V7JM04HONiqYdVrcb7yvddsazIuGlu1i
ijZDZ1CLg5oW6udSSkLrZcNQTASobfB3WZOzLZ7qEBjHUUhdvYDs97An1xRvqLaoOJrt9KEzIaqh
JrAWPhgtMNmj+TRJwTVYdVSy0OuXJtGFJ9HVB6YiQdQK7I2SLOrjB8ddkD5s1KLvAuJYtYeTEpah
KMtEPSdr4fS30S4Iy+CbCidY40CiDBXya73CMBNwNLt7cstA9iQh5DNk5czl4Z5r9fIxk1c9mdA6
GVLwMrsy+GGvYQgqXK7tFOnYRUJlts+A8RIu5x3wjubJoVhRcQJCIuf9YhVH3Njn5y/d7Fh+JX7v
PHhWObBVWjRX5omN5sM/hYurqqknNOVWVhMAwfs9GfExSqm3//Ls6WPHFWlZZsH9LujyHXMJq+Bf
8+sI0gYln8WmuePr/p/VBNQUj+vFLkEIAR6lZ6C/r0IqmXxmmSNzP07AqBDSmdvJX5XJC1nTi7Gu
IAoWRWMUuwBkM4bqzOeq+0a4YpWFTR9sCh3T2U9JtTwot/Z6iDAgDW2mPQd7wYgCi4GGnAX9/yvI
gP8j8p2yIsYort3fEHPyNIP0Pyg7x8p/Dy42PKx8umaWu49sLSvq5bI0vOokShV1qAuOkAn0nQZO
fK1NuI/54hNgyIq5xTgn9+AQYPRYDn07WrzO6NuWwfypH/lWPzGS0Ljbqi6I8jv35GXuoVJSHg/x
X3DXzQ2Dk2lWeYoNuaiMgE4NOSIoWcBXJwcJGcuRY24y8lx3CSAXcwdfEs17MTfS9UWkmJSye82Y
ux2R0R7nl0xblek495Ucj2pxTJIAABrPWEhSBnrLmweUZHF73yqbMuZzHCMFiV91hwFqxYSH2ip4
zGgRtQ8H+QE5cHLvzbLGPnJYdM024NHnIKmxsazGV4osxbqUoUKRLUA26ts+W3hLbo7H//TIkDPT
LoKyEw/jIM8IwGno47xI33wIwQLKxj9bkcyJkI53K6cHLKw3ixF3EC7XyYK3DX1J4G+QrjtOiRw4
foomoPsjrOu9SEFIOqEk6cBvaelV/C9G+YGBvzuXldWweRYf+WamcxdkRQj+EPd6EMXYA8sKWP+i
vi66RhLLVuUoaT7JcdZ7y4RwamCjXQM4GIFNGuqQNRcpOW4UxVTegHS6Ydyuu7w36HEzPDuYzeU8
7OPcGRtNGMhYKS1xjePcQIpw2Tc2sKh6deNyEGMmFjABjFAm4EG97kpuccQjrQRUMtUbNaYJqNsl
Twva7rM1NdjTn+UDnRB9At0bGskvcbugf/ZdV1lVKaU3I331FaU2DyIgfhaEO8juHnu1duz/aOwx
crHqFcdv0NBnyH8r4sIaRrp9STcQ1TqSG8b+DEF0/z6tX/dxzoSYrfPLEGyoHEePITgITLo1tIjv
cdxxCwN3QvmswlD9mO9JLbX0PhU2JHp3gJQC39+Gqa5ocKj9frpSBvzRmrn8ULrxs9qaI++Lbang
q9AntOxkgh6j5FyUTkS5NzvxSbp//SUNrfIjRIOfzQ1YELe46MvuHmB4iEy3+pemSgYds/5dp/Si
jVvTMdKu3iRzUHhFzh2nONfN5pA0k7wZgghKFDFQEzNNYVDqyzxe+6FJYRTUXBPiC+WLFXLSsnIC
y2qAdWmdgN+0Kr5f/qD0RKfXR9x++yKp86oCmL5NZHQv9S+DLygono2wSQfODSdiiAJkAAAlE6aI
nsfKplo2Kq9uE0pTkBlaD51UMusFDl+7B4Lil8xfb5/HVdu6nf+DNc8Bo/M9VJNyamtQTDUctlWG
HTM1hExAR9jZ4cl3g6Ff3XGj54GLT2zykdVG541J4k+1cz48/nkMVoqI2polpKpYDQtS6zl8Cycj
OQR4m91pXZhlCfzAqCFdXMI++tru0E1V6Ong+4sUukPGweOy+034tmGsc7qtoV+iwdrvf9/vKSbv
SYifXIrgqD1VBl9v1GwsbsC34e1+7nTjckrDVf80vZiJ9fWMXM1Tr2zIWrz1RVCPaAArghIfDLtr
Gbh8ZHu6Dxkb+/fkeqBmy2OFloULsz2GT+8GZ16FJFJK+puwo4qYkUEoCmRC3lRDqrfY2wbIDxjX
r9vHcfpzmvgxPI44kfIO8R/Ng0c4PwL2A+xV03j4qN48UEsJwIfu0fQlqZWPU+Nv4udgao64VPv5
g26PNV1eP3HOJrfiN9IfwlhgmpeHCIzXTa4xJ3tEaZONau3RyriuEQQnfPmevuwbY7M20C2NAQqz
SK624LsegnyDlO83bN3N9TjAT/H5lguVKBiGWcwHTiPZo4v9/F/uUNAZ+hKUZr6tiuF46KJhB/bX
GbsIhcObN0wDGBHSVCvck7lL1c2l1fIHVVo7GM158P0N85gOs4GXjWKgUM1mL+Kvv9jw3us5MO6t
Vtj6TwjOiRr9b109fp3x5reLkN8JQdenV5CYe5BTULH6+hSjyb3hQxYbLPRZ+AxeIIobmQHDxS0Y
zmaYqsgZPzvo2BbsFYkDxJ2LRnIXdqgAhaZw91g9zbSQ/7b50zV/Rsr8YwIV2ZIdwUj+k/7kiUCc
gPpT9Tdj8srx/8oJId8WpECU6V+9j02xIdcqv1wSLGqRG6XN8Z9bxuN70qN2lfxL3u8z4dnltzXK
lXV+z7WWOE5pky0qeKyWejlKmTG2svtaVC1Dn59juVquZ3yugajY/euG+OECQWms5+KGTSbs4mBi
R5n6ch2BWffmKflvBJuZc756oV4CqVkYyip3PEkC63d4P86Tpz0oGW/xgZMQnf/xwTKsytkgkBDV
H3gymgILB8Xz8v9k1b/00AzRXwvwIIiRpEt5MQiCMXct7AJeMjf47s/FHiUQQ5WNYsYpIWi5eAgM
7XT7CYX9H8GpY7az3C8IC0b7c0kcZy27fh0qfzNBkRDWhGmMVWTFAyYIuTeVxLJnPvqWJ0s2W533
buM2UBOFFwm8rUU5Sfy7uphYTUCGVClHEqBVL914zaAllCsJvy8WlAH/V0NsQCeAkMaTjX9h1ybB
15tTcHphYHg2d9FHr9scOzDQOOX82ccGgwcP/Jth+Q7B3mOyYfzLfk2BTOuLMr0P8lyinbZcW5tc
TGg2ek6WQ1a2PE/51X6H8CljeIHUCTLYq8zK4ZX0KL6KB0fLJ3DO6VOrQHMICdeA9rQ4S9Po/uxW
A2Mfkx/Yv6T4dW8LvdzzrkcJThPZpfn7Gr31LjOlS34jwBSBvyI5RaNR6FpAYbNsRZso5RyNgFaB
A30s427scEg05TIOdIHndKf93sKayJqFEg77kWiiBzc8yNGTp+yLYA9LfzAkSWHOkjHqlh4ZQi/1
C4aHUMU7+RoaBVu2YpK34NB+owzQJqwmxzWe3qpAi3rTLnLrmdlT8WGXcE9blN/EjGFi8Qqe9lev
FsLNl0GSmtHX3/pQxeTPtBp45Giol21Gg6Xld8PRkAaNKzvbUbrXHLkomiQi0KdsZxWK3tKDHbt0
tOtPa/50jXU54xf++O9OZ6kW119QWSohzngndK6IjWr/7pba0JZmBn4bAtdUMZLafopRQr/EjVh+
rGpa1X70KoZUikZ2F22ux0P4sIVu8TGFuT0OaHk1a0S73Yx63t7qNeuwLOPslQxc3RH5IRch1J2g
ttwz1b8WKxTdabhjs94OrC9ObJjBX5HOjV/91sWKYJUoGVYuVWij8SVvILFLHAN6YqR58wKfGTsq
WHHz6x0jnVoLePwbR5TUtiYg96aK8i1qBd2ddV6WHY5XBxMikGc5cprPKbG62TLFuAG9TZ/Ne0K7
EmFq7VN8IyvB5n6xbW+6koNnPK4TI3xH2U4fILjadEcof+I0KluIq/MroPAsZMDjJSVgMt6Xv5e7
KyjKYM5dhTh8qKEijW65PbWkEqn8c1ymtsRhIGWjb9c4n+n11dmt3543aEQCDVj2ox/jZphhetKv
8i9MOZgvhG85w2k54zJcjqqMrhUNTyCaV5TjyDiJUDzAoi6KwBb1paP2PAO81Wwu5Q1eeMslkgS6
oUS6lfjvz6zNe1HXgUUUP2SXK0NQQLjO7B1V6StYYQAZBXsWW58FGfMHIVZdQfM9SpJtbelxOlDh
F0IRyW+f1lrgHGCRbHt4ElJjFTVOCIeetO2vzWqlS7TSVisPbJZ+c4qjiEz4KGjUl46g4GBC56fJ
uPnMS8kN+cEL9fGtBI0rTmtFKZL/WJ2wD/Pm42n3H3bGBquLE9Z6pNAuAer5uAK99xVBw7MzoQGE
W3uxrzp2S3+yhzfq56acd0A/uFvAbRis7QlSrjsBVLSFO4oh9WxyHgF7tnwJqyZpGy1rKvw4D84D
/Sg/YRL57z7QoPMOrOZ8Fon4dZzSN1LYcyFEQ3mJOdBw9DmopxISgU1iwMLFZdE1KfCU5Cu4aXYY
GtnLmSjhEUwlZFbnFXqnaqs4xiasqxSKXQHKlggQtFOywPnXeS/ovQeK/hlNrusM3lMqU/GO+NGO
r6z7XtstGls8LVPLhrPFd89z+trm8Rf0JIfG2brPK9gyy/gQaUIgSqq+nRaU/4cB0bwCkhootfnr
a4Z8irbxC+W/tcsHOarp+6sgC+3gB5WpubTcuaj1zalMnpq9UezNKZggRrZPizo/DYiZqrBXOZrJ
MF6ev/f9BgNYvHXfk1ca7Sg37WGxMD5leWCgyO1BaEBwdAXa2jwfyvjxUWJ6cd0eVfqjvgfCcsY5
zMMAvQeHoDGweBqzLJy23tXNpxAsowG8UT1AiiGBWHsenv5xAi5PPQxl0YKh8EFNVRzYSPFJsNyR
whNYeItV6kz5ac4uShKCFwiHXwTm/wMWiDCzbyHxptltmcDVru+Zxgia938J67RfqWVRBQWzeIu3
5OorgpzNDcbWwemF3Lx0UDHu/fTiNn2wVBmBnhVVbOzHNDse7K/8c52azzQyGJW55F8GDlLzFHuD
+0yIeqbeo5/kSFcSa+qqC1xWcJc/En1BWlk8agJEiQ+vF6qLBHyBP3S7XRDEONL0QHavrhHzAxBP
Dxd31xZmNcYhA1TEUiyTTSYaydz+qOFBvxeKOWThHQIk6DRO6vG+Qlt32qKVxqMzIbAua3g1duQx
ZSnfsPMiG6Gdwbbrsrp1UEovATERq62cmBt6EVk/Gr+/X71lv7d7a8yvzxeIMCJtRzzYjEjsr8K+
dOwmfVoisKR4WJ62qpuHYplUsUrBARUE1YIvWp/gbsXd0NFfZ3mpH9epHxuBom9ct48sd1CR3r6V
/Is9YcY4KoFcKVmBEdYobbOjNmoLmKzSLT0MYuR/4I+fG212MJVPb9T9SGAjl9OgCB3cwr7dG+YJ
Qinmg5c/JmeKjpdm0I9+oo7YBGcL0YJPw3Lg9tz3URonLGnKSTnetF6KdIzx0s7hhLxQQD+UeEqA
0oQHXy9pSOfx7/ZsZpDit6PKS/F2el7U0nIcvQgsgwmK+KLgT+idLQIAUS11sxTSuy4ibeocIe3E
EscmtX8cd3YycXMwN4EtsKm47Th6t+1OjpVlCruMgBudA2Jg/oxRmW67kVZLwdx9Y8a0e80jrUkT
ijLlKcOLYLjrOcnmCsYOx6MABofeATEa7/reX+1/Xy+uJMY6/notzdrkmzZcZ1SSDX7zUQFQer76
isSS/qzhHS+WqtPAO4mBov28xx4qLAqDlf7v8ICN7zZ6L1zTufV9EPzHoWZbn/zZw9pT3E46+niH
cpkV6tMuJaZvcw2zrjaYKath6Akcay0wWvRSOmpExNuTNJHvaBurEE46ucL3cAs5da+oJx4A7nDH
k1Qak5IpIGdZHRxcK2FwgLt10/9VC5RIzmt9vJdwrYtzEAdSukeGxtOvDMWzXpq/PGJ9wW112yXt
vzAKqus+wsqLh5Q/32KdYlm/Q2NO8gYLcOxQIJqxF7ES03kdEvTFqYr05lMulzL3FeV1OBDWY8j4
/kPk5wfGYBbEFiGrPCavWOsPILJ3rLwn+U8NgmBXcZ2ZZkTiujGQdVIrVvwpFuPulOCx4ROqzeY/
4XKgEM4e/vtvTSAKM/2pCX/JmWqbFkHMgwy7K21eN/kLIP+0QbuWm5oy9A5OtmShx2b2kLA/GKfp
0BN5nxbZUATxKWnu+cbX6tRllG4Cz1QMZIWQyanXKpDV0wsvVvWxxsxfjgyRNKs04FYGGhmWgHmR
ThGrg/VCJm5Bt51HnAk28HRQHjGf4zITGFGdE9r9cdmLzUP3QvjcVAs/QFTvyU7n2FWyiH2oGO86
G7eqk7V9iJp/jY7VefI1A3EBpMvR0ymFQrOAHr7NvG1UApzHlMkLAtyLksL3LkbDewy/tCJohUAQ
6dWbvXFpaXBbynW/eSACSy5ChU2sS7UAJTmwMKOkbPNgDt7otRit8d9F4WS2RzvtCFucMqkeuzvB
QbnCNgEAmLxJbPSNjP3R9NcHCgr4Owl3xAQ4mTaDcpOrg693owWPWakGh5PYgWFKTADFuxpdgO74
Unvt43PyYkdKQ/INqV9gMhduPciJRotqw4WDpoioceeTfLKuLnX1U+wVsDXd26ZzJ1ka6UHBhSwo
cDuTfJ8wPaYokmTYZQLZnSiwF24nO1jHnTQd6pJ8OZpduA7P0apLgU+23xin8yw7yeKuPthNbTos
r/tcjTZGoFH5zq+0ToCW/yr9paqqcwG7pI6kE0yYoswKRm3BsCA+dcTt2xYDC0ejmCoCespqHdUG
oJOnj1JHaeOvwWe4fq9QX9j+qzk+6ElFY5p3y8Uirs7c+KGOdNVJIkvY7gvXy3YOkiKnLdUHXTg5
nYWUT7tTiRKaEIfnDteklw+uztZjrYipvKbjEJ6C64FYAmyQ0iQTlHIq4VdMD0AiGfht2o2jqffm
1ZWZo0Mrly86wrEVZOJDlKwQGFTJDIC0Hoemdw880HZxsc94vD6A8XmYbsPwfWLtV0lQSpu0PQN8
gfx9T1bZheOiSw+dtXt22JGYV4OLqF7uFM6urIg++2GkHnj19VqSnkb5r6tl4qDkJucbfZTm4knC
XApJPzBV90UqwJg1k+tyVerYh+sro6WDErjimFi68E8FrrNZJj09fOcT0crJIPCLNUEAJpC5RYqF
cplWhBpF0sLCJTKnTi7y9fdeffcdkDkF+pG15ufFxC4dmILI0Qhd2OVHvQjVsQtFjvlzfzT+RjYo
yAaHBcQDD+r7/Xf1PX7tim6tOpYb0lWw4L7bEov/r0tL5PIIrx3EvO8g7UwN5hwPf8o445ue2Pmc
s0dpO6TK9xRcdg1x1t+yeVq9ePBG4ZRkgD8vL8okduPrsfzdBEYt+Vs6szXaLInb6CygOiWn5C6o
Qcfwa6qDVRPU19+EGvhQc6zit1e+dLGFP8q4N7KGaDynidHcavbRPAQqbqVnq0NRZkqQgP2G/bfm
hiZwbFqTeN0jh3VE2mauVYxwhVEk2L1TvPiAvbkF53VZC83L8aV3ZFFKBEA4/DF/rbYqglqd11NB
YQrvjEujGk9naYQj7Op5qRtZY12j2PsmkgvL3s7eIzGv/ZxMfaHCkimyx6mZOPdGy74yWZYulceg
ei4nkarXzTYrGVO6dkCdTr+25pY1Gnpskrj6S5DwQmuJM6Lw6vZ28o9tc0Ap0B/pUrQOcPiInhhr
SzjQTbSYP50RonJL6IIcWe5jqyERUrKeegThaKvc+JzQ0Mt5JZQDlQG0Y4KxkZdWGhREmN2hwX84
ufvWXepuIOg3q4+ZVOdmyPROlyMkeZNeXhp4olrnHYb8zTE/BouPI39BezBvS6NKhxkAxQVLSSAI
jSvpwhme6f9X9Qbc4JVAf//kfgWGdyL8zjwTbvmqk1r0HxvlgV8MmxBnhMaPYHDnuohjK6ogfCJ+
R1IaCispMOxy78fQXyuVn9f6L+6rJAW0QIzXGJu58uIhlAOHm2Mhdq83yqJzMVxig2xfIEoUJAQU
a8jXJ2J8ORqQ8MYw0OLZqBtNaGUDn/6vfdn2tXaEGp6gYMTH5EFSuBZ4E8mtAYxaVIMJkuvXojd2
BIGnePrFWhjG1sREPejRwXSfrwznVoig8bQdXKPzBaFVFN/cxr721/wpS5CTALJOPuK9G5AvhQpN
wsAv/pVQkUAdOCT9Ar5IEU2m8e4YEILiGSCwZZ6PJODMlY0mMz05W8oYKaUDj1x+dINbkwVF4+du
ntqM17I0K91OSydOmohAB7PzgCQf6uI5XHLAo10MbpHb8KFwGHK0OzekccNvMa6Xi0y3mK9f7bEm
0pkrQBsA6EDe/BkweZANyDRFMVdSFELgp9NP9l3DHn/9m+9LZOon3mxNwzESKGxYzszZRIQXe044
8x5Y2oNYcU2WUjc9f8iIuM8r3c9NNyp6OnDimf67g/iK6641pyFkUJE57E0PDT1dKikqQqhoPA23
Vitiau92ryYeGcEfnCIN1KzpsaiFB9CnKSfAWOALlQEpfZ3In12IRv4VfQWIJeMKeIq5j/ZCmOVi
IxmaxLJSOrJuic09LtV2PonwdRkZg1P6KeGH9blsLk7LXSjhExykW4GB/xz3FY3LGqZutkNGvdlL
H1UN6+NDPJBRKIOiy0sJoA0TWylXw/TSOnQtDvS3hpNkUkk2gvoy/qgPdSV7Uy0VsOEEXrkrTWI6
0ewYI+CqD7Wa89A0k4ilusZLGjqa/180Ww+qnTJPzS/1gdj2DWDQ7QQzzjUXt88Bt/NaV/6oLp8y
VFOMdJ3tXBy8gzUXaIbfKtAOiV9T5j6mQh/UEyn/X5MWgACFRBr6Xi7odh7uEQ6+IuouHbCv1Gor
uW/4FitO84QEFpSeV5ssPFULCZkPUaNbI7ygQVx/N531jAfyufDcNm0dDaaQcQU91jq9qwNpzlrU
JLh/jCT3cVDM46xwC9TVTviuMQwMpqJlYo+bjXDCBvVQdx/KcLIHHG3oTUmHPX8gFqPttJGi3j9X
45la7SSPiMGECj70sAf5hhM4obEjPs3Z1MiIDZqaeGOocG75/9Jw+Gwfo5OPuhLwJfTgWSozPkjk
jLNKdD9BY1CA5OU1JnTcvsTHxdfocfoX00CBzBHQ4CP/9Y2+mBcj1/P2nliC2SEHJ9ROgo7Im5ua
BQMrx6qzhgIRQEp3v+ErbeBIvT6R00juGA8cwGpctKzRSqqtp6n0/f8JCASglU6EUt9uXD2Dc8sY
cnpSQA8ZSgd7qys35XLg2nBYdP8HP/tV+xg3fdJI0M7zmFCJCqkQwWPJBVcCiG8Rk6J2i0C6mPws
enyyw/0pMSqrae+wiAohE7qcGf+8LVeysW4/FKAvQv4dByUHnVavUWcDsqzc4iapIKATLPEjTS7V
EjnOHmNmZof2yJIqIDLuHI+4pV03Cb3CJnVJm1cZLnJQ+Eq2kSvaNDK0DCVGzAf/NNmyiNn/JHK6
4bdSuQsaXdQlFlPyw13fGk2KurQ3haYmziFE8TU0oY6jQhoVb1bvm8w+5ori98/8qfooYyETQVp/
1FXVz3WhH9/H0dbskk+3qeaVZPYqsz74iV236cI02EWUAX/SsGoUn4hqXKhJXLfESpiDIL7DgtRQ
dBUYxpZdLLaqbkXRY41kKF+hTfrcWBBd2KRNsOtgIWhIvhGzv+nioJVO4+R+jcoCKYXJVOYIOLYC
Lfj0mLmh5WT7CJGeqD6R8a1E6m4SVIBsgR2QvrS3zMKKu4cfd//du4z+4tMJoc23qpfW6Hsi1yb3
uDzhHa4htNesYRIGerBoJfGML4hMQtWIit6EsUNkavB7bI6Ceh7Sn1wvJYAiMkowgsSJntl4RwU3
dJVDRDR8wbKJoN0oywKsSYwMggXj+YElerhwYUmeauq1GLD5bd4wWQT15W0HDzbi3wy7Y39tgRjV
pMUwtVAQD488iGYWdsTa4j9hknb9B44JRwsJw4ukDPYndUgU4C1subLEHF8rOYbnkmOgYvKiaUVF
hfs6HveUGTm7NNW+lLvbTu0GCMgIVG8f6H9UKK5JgKeeve4oAETC2FdwP1uJVxhzbi2xnMJjSqVg
y0DWw32lnKW4nP6FVfM39p0TILGKIsvzwGXK9mVRKuDPl4XgvptD05ZRYCLzcFtg4uNtDoimWwoI
7gpwl7aNd9aD9PNgA9EtUV0oUIjmbcmfWZrhcY5is8BKfy/k0o9eKPJ8JG/9ybYBZmIUfjyTYTOw
OzUm2rY8KXfhA5a9ZWwsSrmrXB1Stpq09PmZCFDGNSCYJVy5/f9BiNeICoDmPxpHINvvdsWZUHG9
PMeV8dRiAh/Evk0d1afjjbwArNoJwNj3dC5pAgDMi2128H5AtsaTzVxecyCI2yPM2QTl/zjpUqzH
BtonnGoOFfLJlay/c2mGPveVuiLhRxQ1JH5Its1UBWvoeUVNQr0i0unmyK1vK9eyT7VABs4scmKO
YqGUv4yTqIRvFcd5EJGGraDbi4xGu4EZq1JK5AoBQ/KTtU0PZAM2au+8vUsBHQ0hpMGYVTbHHOZV
4OWOK+NwShPBBZf/qGWYszNpXBsiIWkvRR65NhoPlHAXhlly3zdHn4T/7R2Ny+mTjMfUIefLb+4w
uI2HT7ukJRq9Uq4tDGrtIwHXBSxij608A5aey/QomGDtW66QaCxz4FXQyL74EqhZFkMbs6pla4Xh
jHPUMzVRzAmk+x8nP2la0k0tW68jaO4YRYPfofT98UyTwi3QPHzhVQnI0KSBbVpqL3NpXUBtgq4b
knBqzXQLiN02O3kKiaPa9+7qtYiXabLBgSIfTQ0DAjeWfioZt9kCDWi5xGh+6/rNa2zvHiWJMZr0
LTY4jUbhI1oxZGHcl6ujMJd9r5VeJhkp3BU2IHnDKMV6EhIMNcDZi6vulYJyll5cw3f6Fa9zsrVa
FWD4BXJ0m4KH5kw5rIo9OAiYk5npIlyZSB3uQOIOsHT768ZRZgLvS+xgywga68bxN/EgysMetwNY
A5qFcFdxLHdnB4PjcXqd5m+f7DI/Z+rCrsWL7+TsiRRCC9viE0b40LBIpShsSIhNzldkMy9WPPbw
1RC4CqCCPJ3K1BU6iI9lrTLb3Vu6yFZEoaJim1eWr5b9jk8XmdcRpCSiL0hStX3pg0y/znkkeryk
vYLwvoyuYALac2Klvx9bLDfsopKaTDUCHmKETXs2xYUXPpTfxMjZR+auFsbrap59lgp55BlzA2G4
4JVEJVjhdwqFrm/OtRvlc+ubqLPgp7KDrooqFbJsFpi12T0MASQfl9+gzZV4atTYUBCmjabhVxbr
6tGZF1W6+i0LnESADFTfr3ucGkww3WXrKcqfQEz2Wgm38YQQEbJnY6prriskv66iWPeCfnPF4YuX
9IZrvmZmsORz26VmB1gA4dLQSnYiRQTcPAtpvFTtTqH/zNJsm+c6NzWF0XjahpSAfy1XxFmYq7dn
femNynmVuqM/xmpRNwdAygSfEeW9VuHAD2Ow+3T65inzlnDzTUaisrOMaj4ukb0yR9B4soqwhLLw
UdeG5UKjrEq6zv6vJROgaGRkuzqQ5O9/zweOjH06tNpInLmD8FACt6SV49GY/zGuqNS1NUANke4l
ivowmd2cEbtceHOH3mcemH9Bt9Y/dUE4+fYHGiiW5WBdE1XsWWrwJrR1df8eGAQynHlcwKUh898Z
4JQUCFf5E7RJ3hNGm3bdxJQzLmowhqb+8hSYfSmJsk0ULwCxYbRICoFUYCVP6VIV6weLRS1xi29n
os7DQQwjYUdCIqCMochqzLA37N4xz6dLaupqlNb0YoVJmWdwKC22ZaG59RDY7tTqALwhoz9bbOeF
OVFsRbkI8vw6kIwlUq4wNRXQqc+SILPhC5K8npUoMNMnIcxERLtcwXQvJOO+g4OpundOX8mIq9IF
Zz5lrWu1rPnssx5Rj6mKxJdWC/c7DOCTPUon37Z1ftKwTbdB0CslHeQngLVwcj6UC+R1END9LDaa
J0OLulBhe3p2SRA54+oromFdSyq0Tofa2IOPhJQrTxTPhTEqSdGvHM/KIi3OagYr8sWdF/ru2xcu
E5Psg/fpeplhtuUV8XtXDDHt3bqi72eypUmBP6T/N84I9oYxHr+kbnABvcxyB/2Ju56eqj6TO5l6
A/VDeuCrC0auCrVHk/I6muU0uxQ5VoGCee3nbeT2gzzo2Sa+sqFEVGO39QhiiCtCXXfDkYd74HMu
Ns+plCkDAW1Msp/6lXdyqk3eh5hAqH55HZ2ts/joLtXcZCnb2weGOpic988wl9YsUMrAGHtGIOPe
3Q0xqsd1FAmLI11bJE0pYWgtvxn79pCvIeQfC5/JkwJrZTMCYPaUrL6CUT2JpbKT+AHTBWl+mBBu
luk6Qd7lYsmIyXt4w0y+NsH+6DyOqpK/UoC2ETWEcAxjpasvPzgnC2ErlH3gTgM4FDCqWDi67Cvj
DwkgAc4HtNQqjFkb0aJfzLJVY4A3qTADE1FFa0FAQOmbec+qzZogxBoVOlUyHILTx3G/eA+c30YS
jF9yhSufAmCHuvWLfxTmWwalFLJ79GTx34RaBo5+11Z/aR7hBnyp/3ReSG7+F+KdeQhkKv5IgUl5
9hj0Y8yDnZLDCFqlHJdmR//haULtTF+3ylFkkcfJ/UuXHMnwgE7Y7pQ6pwzmEz5aTuZ2WcTdHkm7
STjzSqVGROXRtP8A9Yt3+jIb0SshIyLhVMOLoq/3qp9vNAY9xpSpeNvwyB2cNw4m1g9y5z4753Ct
YvaIbQ5rNcmI6goMBuDijmmktO05mD+Mlp9cYVtF4kg/uNqY0Q7HVmps010j35d4/xmFvjCtCwTR
lxKu5B5B/dpYSCaxMcuAreAjKYA5PPcTDHIs2g7gC+oDNfCF8o79yHdXyxnwlaWbuoXL/WhV/Swq
a1tC3Rf09Kc/pl6v3b/2EODCVblWWXZ8Onp/+hp4Y5wKvI9NCrxrUO60UZdN3GGGfJ/px+tNRhDj
j3dBZ6zxM87LoR+THjEncNX6xMLL1vS7CuGhZ7QfxeUR8zldlNdunFRk5M8rXjB0i0U4C4+qxx02
dT5PIUjHMvh1reXaybGckraBAJti1CnJ2Ur13qAM1fL/GFiu4BzUcabCPK/1JaQpmpTI3Sa7i28I
+HnOE1xVsSB57fmEZEDH0ntdA1zYHorT8fcRr7J9xGvp561sLNXzbu14QLQorR4YRYRciDTT2MsE
0esyrmBLrjgsgAMSiI2Jc+hv8t72Nee2Wy24iNFQ2kShX+MiL1lyJtzYA0q7JwTNMW4Nv7UtZqYl
iJqvF54Ck4itTBEG6W1N/eo/NwSq1lxbjEnsXRVDyO1Dw+on0YJBGGQ1BhkwmBWQq3J2weqmJOmx
ygsImpHzYPnVP+wPqOn8H4gz7A/w9DGScGa6lvwfVdKx8Ibd6DlB2m0ixnADfBACMlNoh+h335iV
bdpqxJsQhehZuVYbvJ4aOD6W6XlTGxgV5brLciIkDrbx0FfJ9JrvhRm4S5f0rHvKTTW/wY6sWba0
JMXdyP/szPmPbL3LTDSegl5BcOHrhGtw7AVz/OZZVWFlawhAenEfAHxNRiIqp4SA1QNQPJhMdEGl
A2YpOT5zbuQ2CqCr/AfLYWD3pOE3mvFby9a7Q8ygp2sD4PfhaxbKsEnUM01BW+/xq2/xjadZgSHA
Tiq5H8PcQiYiidtC6xVIvYbW5F6L14nlR+cNAlH5M9xZSgtxCd2FIsoeOOmWOzAcB75l13H9+YV2
b12L65UfM5oCZVJQxpGjbdpWMFR+bxzieLNZHQ+ppSEVvHkKn36rOKKridT3n9sGPoVpSQuu0v05
GSZz+ORlOTrHQKykOCj6nKbZ69nIwsUNnb1rCKbikAGHIsfOW4IGnQ7ZaaMcGddblkelvPuBLjK+
QD0ewu/WW1ksj7uilZre5viUo7pEMEupLMtzQZsRxklHEyj6oUtKF2YfihsSUMrFe3PrrlG0KSEz
08EKHMV7+z370oVvjPUrtZ/AxKKbuwx+pgGlfXIWB9rSusv1kwqE6f9fZE2+pst6cwO/b70+zfDM
/Frf+ePKzzClWYLU4iVTXzYaVxcZW5O/hlMFz02GxcJHAs9wZmG00Wh7FmyYc/VE0S0vd1hCNpZD
7j/ghRfMJMC5lccRlqVrWxmvhi8ihWlXYL14JZuKsy9Ltf9iYZyfWGsqdv3Rte/j/zy78ikkROWX
95WGZd4NkARatTMJK+O7Ihe9C0GpAjD55IR6Xm+z5u7N4TlhmJyJsyulcK9ih0yLN+xCLzY8MGi8
C1fU9spbjAkvfjrqr45BGBmej/0IZyfO2auovPXaNUZy4SqxaxjxQ44E59PRG+ub5HvCdqEdpjaW
3ujVe8yr5WNs5y/pFP7PXbEy4u9NKYS9dZnO/bzYYPsGNG9a58YRgIFF2DsCUu1JAQ7ZLoXyzGt/
lAGxYj8prOlTubl7QQlWNNTo0K8WkLFf7kkEavnk8WtA7+sDWi20XCMxdyMiBZUU+yEQClPjKk4I
Ic4l3e7/V8wc3nGf80ciH2VPnLmzzOEI8pwCRloGl6JiAMPW8IxK8fRUoqowqLSx6kcGkSvG4Ux9
tLBXzdtjeogsBVD6xN2HFUUi7aKHbn8L+qEU8TNr91b2cmtYf0bdZJeBOcsJ+u7m0yurSuLHQsvi
B43nmcxn1pT21uSz78Uw0V1S6OET9dTwvB8kwhyIfPWHr2fgA7GmEU9+zbOrUC27hvQfz5+QJrNS
uZv0hXfyMs29Tqk0Lu4ldyjc7Sigwv95OyXDAo6iu9dgo1FSEuThYW/9wA9x+Kwh2cAw+tNXRk7H
URfTyFL1rWQHuVdr8fUIpB9OPvnyVFnGPkV37/zewruThUltnSmbjNTAcoPTCfGazF2b50tcQ8ai
8n1wy3T0Lt1HCCnXAWxQDstBwzBHguc9ODMctpPQWdS/QNLzRAakC/qEvj4tIE1zFhwgjtuwSgIi
xdhKm2kc0HliGyh8ZGe5phDcYRCk5uAoNJHLdCoM+2Hs/6eiKRSxtWLD88CcCZGE9Lk+IqyxFwam
sc2NYz/6kgYQlkSutl/zJL5jeeZWXDX44u2CLF/TQhHHsmUYWdHHsFGZnEwId1lj2NlSuvh11sXO
qLsTZBSJArUdwzZuh8/i3YAqc+S3LMHGs+TzlNEKZVqVhVkxPLzkt+subSsKnoU3dKKGi+EMVK2j
tFhKcmmuAfEc6ILf+mlMoNH2CidehQfqF0wWX9xcuZ8eOPR58f6Oc7Q3uov8ioPOEyTzpL0VBvZQ
Y5VfBiPBoXeqMz3pGbdV66twz5bIgOgbX6RnOGihyLdltBisdTdebXSAPuc/VE5W7r+MmTEw2uJQ
rY3ooxRdc6yNtav5Bp0vz+3LcWX98+hxaiaxoVbIRuMAapCLm3ZCdgbxYePqlvoUyZpEQbuuq0cn
Z2FBYlCvcF1xcjor7sgA1zcPX80MXlnY8xUGpV9JY+XxzzQOnVUBnRCX4IweepuztKrsJk6vUPL4
NLoytKvDMDLsdJOByetiGksuvRuARPmh0WyfbUH0vwH43JUITzkPAEmNRnfhr3OttO23OpNnsUws
pL5ja4iZC3Biy/e79MGPXGmylVRJLetS2zY0PKyFbHAHpk5i9sx2+JGDVHSzcfbgitOMlOLyo6F4
JcYwhbmqV0AzIb18NFMxOk3L/Z4giAyCAIpEL/tqF7j0BOBOZgftsaSQyOpvQdQJbBPip9fCIno2
xC3H5gVV1zrQ2AiagtFZDwJ5ItWPvrVOUky1Yt2ZelkmKlux8Uxvnoy1mKGZTqwCUmwtHRGfqt94
UiBIDSFExQhHtvWurnHUf3gI9F89NdissUqwGhvibv/FD//Y1kaeua2er/Wq31qWE5Bv8afCul/R
lvAKK54LFg7MzsyNR8oMbxkygvTVYtb/mBORwvsphpQs9CmccQfmpxL+C2EnhEGlEAtmUbqmHKBj
xOOToXe9dKxzcz/Ta7IB2Rl29ub6v54PoJ0e8GaCHj0OFDBeG96DC4FB+wJ4ee129MRGx6B8Q0nI
03cLM74mO8rVH6gthO9jhHtExMA/9tPy/3aEDYY4tbpw0qxJ5+hL7RDO24xlhAPPUO2yVzj2n202
9u3KM6FS/zlSCtrkAZ8Ce+j6rcnfY6edkynRqa+3DGq17XMVyPQlBFgpU7AJBGLckydeEsZ2bLr8
WCv8tEoPDgocPL3gz1tJwskW28a0H1EYJCFN0HLXOId3yIQCJoeJDZjuKt9LPpXTtVHk0n/0oo+Y
w7EVcw8t++wLJyE3YwWf0vrP8e156kkMqEJexIW45ORP0Y93snRMQAVmadZCMcXbW/z+xPnrx87Z
dlk/lmjw+2uzc6hWUQleYCHO89luy+E/4w7w6VKlBNLr7U5uaTTD6InaGvv4UQCEY5ca0KepMU3H
7j3VpenYCbfdyvyebAkkAQagm83XZdLskztwt0ZkMNBiF2LeWuU69765Rhz6/Q9qxYPRU2MkeS4c
CbVzM3mQEC8evfFcp6IYtIMn8xLic9EhUyudK+8Q2wfRto/fUU86w8zdWSz48NB2uUzeI1pOp4vj
9eH8Af5fa74Bf2H6TfEjiUUDR2rstwXmjQ+n5UFu6AeuRWAhLgthGTxYsPhwypljYwqRzG6EU9Cn
dgnIiOXHRqlTSTFEsJHjzQtCnQ541vr9eRfnw3PaIwCYD7dS1Nf0KFw8/OsWK02jwYeZWjBaD416
hK1/hOVo8R85CTYl73jqSq3NO1rUTayu1jviUQwoyLG9Dha2+WEzTJw9rp0yBLVZ+9sW+J90U1Gr
BieyupMIoVMUeR454cKMILaufa5vnkKAN6qX36zO0l5B/RqxHor3VY5zQNVDB5eb8VuhrseOq0RO
hKSLW3D0yk4Vm1H+zgXbpa5fgr5FGs4m8wsPZLMClg7REtBoBHbu2fKO1g7m6vQBlXJKkxSuCkzc
b73xI1I+DSPYxPNefXXavFREsPuwhRSrY424ouJJnpFSgWx8uItsk18KfI5lhqF5XpGO0Tganq7f
u1vCCgDKn9UhtU8DzgNSJBPJnLVou7iw/K7EYcJTjtY+A3YXBPN6h2rfGzKNIoCxslE47i+hg5as
C0pVjwEdLZp0TXkBa4cgYNcsJ7f5mv6PqEBVWOGBFfsBwGKtMWp5YWOqUaYQ0Pa7F7mRbSPv67Bk
PBKnqJIro+x87RQgXRtO9KriJKH6+6Bcg74wkVfjz5AThu1NT6VzGmG1Akcj3yOkDnbXjXDrd0Lw
Rx+WZ7l2M6/cuSdpwxTUf627Qi6TtktcipqvA3mapxgTXqMv1jlCDedXdEUB+9HRPXVLFrsqRtGv
HTMoS95KactRIl/pnsLWn336Zw7GDIjjp7MiYo/t6dRxu/tZevcHdlmNWGiadKdcocAsvGSuyYQF
XqMHUFBtYD1zp0Ku8FK2hggL+jq21QYszHeB+2nGwNdMN8lZ0Yy9UJQ9V2QdYgeABEarlyNHWVQK
TBRj3UPkL8ffexH+KeK6I2O6jxHgINhE2wUUQky4hYGP61k+bg+UfweQcRsx56FcZ3ceNTY0XqKC
1bmxLEoASwA+7klaP67xjNqIxU9mgiX+Aus9xjyQWbx1LUN0m9UwSA3eBN0VI/cjJiGk69bRrNg1
NNs3NXBTuG6QC2T3ri26XZGyCfioT3QPgTftfwdhpNltBlbArpaUcULJWBuInmpzirgKlfOvO+eU
74h9QmACTOybpQErTQ3zLcagp9VfPmBzK3Pwi164zXci5a/MDj58tLDE0a3oT/eYZgEuEPz/UD7q
bF0EslXh5YKoX0rVJHZFti90xxGCUtqcFOgP1KJ9Jv/oCBy3gjjYTIUmiLpopganxRxGkCVjzSFp
VJsjmZt0izongCYy/O4N4CuyFCeYLdic7y/pivp8XYB+SkXPBn3fwM3Mgpsi+vWfj/RpX+jeMK8S
HaZ9hPvdWQDJ7+4FGGMNrM9MPmJkCX7YCeiFca+EHX6dvxsUQZKF4NSpg1QIuHo6T511mdI4x4jw
0brO0SkhFbvICZ9ng/LkyNonsoj6eKczXSukNgiCldZpIY+U3Srj6lPWSTfv7Vo7fLnn8GZ6hQA/
uAQzcOO9mTeDDT3ZRiPbvOIe1bhaEWjgYbyRm0ue4hiFu64vJ0lZzPKTyFn29wKPkdiuvu489vah
rWhQmmelrC9K+Bv5uuFE7GuwnyqYIZLDOygLmfQ0nEsQk1/Xn++JRSuSqwuQ4E8GD1PQSK3lRhxS
k4ODXffgojXtvs2PQ1wSzSboC93qx+RfdUjVOJg1cw5b9sKrOvwe4hYrAUON5OHHSdNWy92KGbiG
WpH8O9zo1bY8BCGsMxi/nsf3raCfcMhwt0Q7su9B3Y8PVH9fEgNpCgEcbXRNhG2Rmj4M0JI58Y7x
XqeWKHGJ5zu9igi3clV3KlaVwsqvjdSFE6aEwCQIV2QZayFPDUBstzbNe8Q8u1Rhm1i9pI5kbO/w
7xybm4Pq9nbAT2JHoGHFd+/yLwSv8Y5P7rRuXQsHAv4GR4haEpqWyYwRb5BXy058FAmTFhD+qdCb
Q9erROXKtObDH6oqmZgjgxaq8alg6kEMB4J8QJ1sDQUSbwwhgAPdGbgnu/qifWAGanH+MFxwnrB7
HtlSp5m+rPaPh/u81BQGQYgBrvYhIvgSsExObnS7xHgOLbnGcoF7NK2mN0ynZDckFwEBKRWtwT5Y
Y6yFLnZhS+OlP4i0IXVF6Jr34Q8G8UkZK+9PiddV/Z/nqtCpBZt+pfSRWdvxtaS1ze1LT22y1w0A
cg29Ii+3+B6JHft1foYzzOCefVNvsFWz6EAJd39AsBfr9Vofa/sf35NhISC8Fw7Up/CgQHFD6suQ
biJjWQkZuZY/iHRw/sKGeOtqKZemNyxCVhtijVdo9NcP9mm4woE18hLiTncX9HPyM8eRxe3rKGF+
7KSUdLkz2c7ODgmmk5/mcLt8JHVxUvrCg6CtLAtr9jY2m/jxD37WwPntSLoyPvBvHJaRXIpMhsFq
cZgl1SfHenIb0xXA4qxKLcC2+tLNmf6/QPXAzZvdPqhHHBjGzEFfR7f01U5hLoe04rgE+nADddEq
MFlI7NrkYPgOcuQNMfx3v7n9jV7uQQflr0Tj/XA93VipXsGv+QW3N5/ncHR48u6B82Pa0cZw9GaY
gLEasAAy7gPjCmNg+3WL71obmQsfns0lRg9XLVbjqavTwa3UtjySdJl2bxYkkW58GV7IiLcHR0qG
w+PfkBAcQVOHUvGZ1iAVqzzoLoVftuxMWiVFuifUqRFKMUDt6AEaFMduoPbDuDA675gZW8QKSG0U
6+bF5TQz52elT9+ODWcNRqFEQRTglH6EAVD2o8y7iXrQYAfyCGw9t4k6VsFEqO3GgBcN6IklhVCN
jZ8kb5iAksxHkcNluW01slH3vWdszaHuwNwyjg29Ii15r3y0epOgOH6hD15GPL+NHE3vatvOxra9
kIxMTTcN426zBMyg8UICAwK65HQO7KIeGyA2SZtbQtDhfJuELY7512MYLnqdD9B6UAE+E4Fea9s4
jFUgOoeuTF3RmH0qMgxaA6FOKH9nksMBaYnqDRFsPrc2unAj3OnqKAVYz1nWGvY8alKUanU8aIXR
R5KEtA7rUIFdXpD8uIcdWKiYhvp1TYhVL2Iq6DeJeQohb2eaJcjLZNoBJy6YdYyFzwDsjqODzuAP
pS4/84e5MfJPwx87J1blZGW1UGPSSGt7u9m/L1Nmz1ZIjlJAx1ArIv31VfDVPFU3iucYEhxFG9jp
bvTJUgsNbAzBAaiwljZ3vjsVJ3m7hMQJZ4oOW+elq5v3lA+uCkO+zh2Udkx+w9Sr1095UGjiLOuv
lsAypiWpLyFb6/vgP8I3CuyKuj9sBj8coVGlU4yek+5wZ6HlL2Q60eALAFbmnL845TV4WWKzgdbh
lAiQJ96UUOGI6rq3LaRpwcE7ogep5N34xtVFyCvW/8Ixf6LAXbab2CFdbZ7Uzru5Q1yQskb5e8Zs
Mq7oEkzrCre/bs9DKQJpNO9U80OzwzEJz9GxN5ad8QjgeLsRjr86us8/1oJ4ZcohjqBKm8JQOn3b
A7a3bzpSVDFBz/xZA70QH6YQUeNdaF3EM4sfmCodxuk4noAjWiRu/K1NexNDPFGRYF4Wr0EB4h9j
HXdHVatfnWsufY+HuIkoQKscwTEH/TYdi74HZ5pYjTj8C4+CT0y2lQOrkra2U1xT7XEp4Fn+D7br
R60mZGvtSsBeMpfMwt0vWkQB86XYPlsVnQF5OoMGTiJPkdIuHyZc1sVYwFsbZQDTdLYMuDClkfFs
VYj9SOHm2397CcMCkJs6RDzjBaSGAk3MGybfghXEV8/uyRHNNEXkt0f2bvKpEPiamBreg+7Q4hpg
97Y7SVtynLCh+qkjayo/olawuCmhbVDwNqm+PuzKbOrzIomAkButJvR9zfzs2Mbmxx6+ETDt9Euw
AMvnDqKaO0hv1JUKZE5a/CtG/hSCHnTBUDGe8dmo1nHXPtmhpYuKU2ow/j3M4htu3hYyiBUaV3WO
0/mZGOL8jChTbmiI4uQMOv1ICc4dqCqJxtbfiK1NzEvhupGvhRiEynl6BgW2LGqfxHrJ4amvAKD2
hqKJ62dhu/5xpm1rjDR5bQByfUJWHArbQGwU26lmIbAUh4HSNBRKIyLck8TbtHzSM5mn9g08CjsD
YiNxGDNJXUu1P6y5dU8pEZKaXCUKuhSZNxe/bH0oiab3V9oYWLYbfdPiybNQU28ZBcfGL9VQ6zbv
3lYMnbUCHqmIPiterut63I2twIh8hlX7dhHgIyxBF1FCY9tO77lKFE9vEV2hU2R3igq/nexVQkN4
oyTV/xaMx3QgSTtZxCm3qwVTshiBRe2Aqm1BWwdJzFmu9/GuukmoJ9VyHchY+kyl1dk1qvxlNGX+
hfLq2rwHPMujoOB/Bi4pDG9cB/IemtY9Xkzxn6U+32QjeryF+uZEFYOIi3U3wZ6wuE+hiQSTNVf+
ejlzfYQkoEv8EqM0DBadkL8/TBl61jIt5gn32wEMq5hm7u2B+JhP+A1XQlb6Re2OWVpdL74cjr+Z
oBdY1XI6HDdHdczaZ4R+TU1OpipbLVQNX4Xxztt0XotL4RhDo4SycXojjBCRZ8jb+r5DyxuSxYr5
Gb9YIK01CbQ9bn2ZyBqs8w9LPpabq4Vy+j7sIkVL7jBHi9D3tYcPWtKoSzFaxpcmHoB4p9ZqjIX5
YM/ykSKztoZUj4tPlOXwVMxa9BcK1ShV/2PRjy7XihcyKxRXHytFRxfTDJ33mjvC8/zA8jo1TA17
lqt8+BcTOhjuuirLH5EDCNC2NZWSMH9TPLeJdPSbzmAwtsz8gzKDEfhvwLo0OfPZl4oCJdJAO+lI
i1W63h1oJPa9Q5sqb6R1BZeGt+/Inebn23QGbaWefyij2KEsN7slS8/sc/RL2+6nNmMPuWmu35HS
KhnmdH7helJ52XVfY9DciQxn7DQAsDrs9Qa63aB8QwmcViNWzX7fvDGC7gcoQqziCpyA4AZZ+MTY
bnLEZMuwZMsMf4uAmcwUcl25LLfegVW6/xYTc5sednviODYlnF3/jMQl4x2vzbZT/bvZeoUgitmC
okbUSfpz3t5RThkCm+V2YyLEfFmWpvdd1Li/ApkUwkI6G9N6rxUDVClAF+uoF2OKg5T+cG+f07iO
g7WH3heaQV7Utm9cCOv22/Mh4tWyKbdcO7uDOZovfPdsFHLXLzMDJTwbJOURKeto28mKQ9AaMeWK
cWHbbAKlNtwGmmKODtGuP0mkSRbjvWUA9uGDiwGvIiwXO8xeTjo62oLPMfyDC6ruai6ZKTgO99ED
jVm3cDHWJSQqgJz64d8MWl40rrr1qHk5cmT1uNxesNqjmCA1w3avKNw656kIejUW9nVutXztD3UT
qBwqMxQaqo8fC3TeLu29usHAF8BrmxqsXQUZvIl3skFCfZab72a/rkNo1KyT3kbsKpx1MQBT2g/o
oXMrtPCCmVAwbVzrXA75JNPNTu0NOqi59rR6F+RNvCaF/XBFonh1A1fA2fTt7p9JfW6rpPZYRdfy
ZW8UrkUgWqJIyY/drXRks+2MFFir5lXc9K8Hq1WI3vTvGWoi3rPHp8MaFJdS62pJj0jNleb3zCTo
wUrFwwxHxXn6rpai7ticgGBFdbTF+YRw7zkvT7RrG+mhQII0bDyJ8bFQarcEz7QvdDSlpmIpFjNO
Saz1Tw6jyjC9q4BOlDKzZKhTqjlhh/Mrh8TeYWA12CL81Jv7FYzv5KOY9959sqRLpfn++oqN7YnK
/mQnJXarqT34JyXUW7ShCsA4rYHWuLIfg6MpL7bJWh9lLbj+wTHYADPWaL/zLggvSF8ONXhML2YG
hKlEOKCLX6GqTh/HFyf881dUrQ/ewdRxkBWwpjKYuoxlF0x2IK/MSBEBUKJK/wh73+tD+Ch+Sw1L
Zomjek0KXIerZ2QNi0JxxVBvbi4OykalqwVEBMPX4bMNRZ5ne7Wkd/TbBGeBT6jb3CBBkiBlGM2k
ts5zISd3MXKe9WzfYPuQwuK88m0BzSbrYDBoSpBJnG6CrSVoILLRcF8x6EjdB9g3kc4/E8X8x7kr
88+d/4xoejspcNJR6+ROXRTfaveS7t+td70zXFznPPerJRvjGwkh8AYvEEZt9KOibleuTJkOLyz4
NvA6Vflh/5TOXwMkXUr6NDhR7CqqdLvJ13+jkQu5THgozJboTyubZQWbGoqtY55bjJ7uQVfePXGI
vmBk5zTIVTiYkmebWi7fbjESem5UHcy4MjlSvwoX6EKOaTAZs2+vwX7VM3wt1pbHrE1j/iwlDmvV
Q5DO5tQVB9ho/zTj60bL+2QrFYxzRtPhQw/4i0c7ZSrB1ZqMugCclJUM5Rcdsf6r7e1EBmNgce4Y
7Kvuj5w4d6P6b6yZRCfHcihdXJ72Jq6iOIDUQMnJbMQHgAu5BDOo/DcGbWzaeoglFw6Xmhv+gvUR
LUh1c0WdvfhsHPiEvXQVW173NYWOfZTENSQQY8OdodUxnWEyiTKGbqznDcnNMVz1VhnG/DKYGrUJ
buGXfCRuj6js3FdIE+e3oqsZy4+hiXL/iqn4kFYWGEIPEZ+eg64HCuUJgt2d5fJZx9A2GRjsqm4f
EPnJha9COT2RKaZ1MvUSFjA9y09xspiUVhaLfLUQlbXJFW+3H3P7uWr6ahkvVpHsGLXvCgceiAxD
PF8muwOpbP8W9S2vcSjFIJaub26YLBRm1yXb1tWp8eCrpKzdzUcZK+zZHqIaTSkDj2ob9eWnLk4M
2DYvd3gk4Kn/+N5ICconE94lCt40g6Uv6lKlPahPn2sdZ0IoWLcplHe8tzyVPnRvzlnQjKXQgdYl
kjBPSSfaUhOCOguicorSpdiU6CD2E549CfqkcPWBiKNGsk2Vp0SqB1sD1Is4YuXpbXSxrlP0dxaR
ngHFweYYbjBBFVXgMS+cFTdyPOjPeJsNBjlqJbE+pGrIb4A3Jktrnp7jD2M+vHtghSwhTeaRQPhf
pc82ZhPfCIbnK8qc4YCDTkPq5Xvlvf7p3t66R4TBIgwS/aO2rG7sK7jv4GqAkg6nzJ6Rgr+1ZzL6
BG0svweuclUGA/guITZguZrNWgi0iV1yK+xvCSN/L7n5PJxBjwNl86fDvhMVfheZS8MgSDRzVc/m
ubMZ+NrO13+zqvtuEFjhrIDTpXHCpbUa/VItVM+giRPH7uEQrgXGGXurgqNLKNS7RCe97wKE2Z+a
kfS+1jOpsZ4xW1t4RAIWP17wCg3DQkgKNTs3KgKzHNj/haOSA+6aqjsz3kKeZqIEK8L77/UCkr8F
z461vgnViK4bL1h5WQ1X5ZeJwIdRvfxh8MMOHGNrSNWCS+cluECPQFIlPgkjRKPaT0KO4MItENHt
36q4NSogfyh1o3pNX2FWtjlbfnKM39w0WH1BO6fanoLGzj8h1scLri0Vylv+wKijRhv7mxOMnOPr
Gh1BldgiMf96m5Qg/i5iT9c2jFAGxhISpPTRxGexEukTHcrgjnVoo1OaFhOwKH1LZHUhg56rDDvc
agxGUxaZxL+MjWcwNACDLtVimbbIRvMxiG3INwJHFkTvtSQX/0GM0gLTl8uelJ4HBQG5RtKva0nU
duVXPJAQoxni0lBiRynckYwJcpk63w3QYN6btCggAO6n1uUWWyaWytXWWHZWRbMoe5HMXNV0nJ+v
jKoy0P0Q6j8FPGNqN+G/U+hO9UMtu34ZpCqd2eMuQwbg0UnIS4QESFW2Tczm7tJv6lE0LmpPGUHU
LvRSuou7tmtjyMa82T3TMzvM4hS5VYjV1B7P9X1JZpPk00UXshbeAHooSGB/JrNTCj/P/KowQsfS
M0x23C/JttHBlppmWMSOgS6yXaOxLQBgT09p2+JGsEVklR4EQYo6zpsqgMXljRL7kE0YiN8ARuOL
Ur2vnIcRSUL7kEaVTtx072qXSZWCHuuDLxvKOcwMqEnT3WFENyfuvBeBQROxB3fhnNCvWwEUCR7k
VaelOBY6g4DgfGbLFL1zQo4N4O+1MyjQZ0/edOhFBsI0EeDu7WMXgVL65SiBcrRehXW2tWzjpGNT
Xzo3T7qRpoaAzA13RP2kQ+36i987uB5I3Wtfbt0hUDp9JJcUFgPBr4FvuoUFNYzoxraN22s7uqq6
dn2YhLPVI5Qnv2Rz6lKdIeYtwH20RIUtGmADV9YxFUXUatRYriY0XedwJqB8hlClhApMk8nhqLsZ
18rYqypy0YSQWN5gP6TZNzuBXwgSI9syHW1dQPlXUpLpAgGtHcpXuHl7kqz0/lqiRY9O/5ox8jGu
EJ6Mx2WDYaJ4y6U50R3mwKjAIL2WCYgEuLImiDyEJ8UP+39JZ8/mbAIyH+KJVTpYObfHEkebC3ix
O6TffgEZQSbujmzI9O+n12nrqudOqjQBmd+iGRR+MD/RcB0JK2zzFaRetc7zZM0MoSva6AfhPZ2/
1+h/9YwBqKU3ynPl6uLyDBk6A8sczvKSlFDiBH8H209yDDlTiv86ivZlKyPSWZ7KoWz3ucUA2u0b
gdaoSCKHeYx1XK2D5ZHIXg8n5NAHfXeT6R+0Y1sYWWv/Ts7ffNJZDV9EFUXF6PijloBZClPOzKqN
PW0eh/IMR+zh4kZKtdpeYW0Ndp+FW+G8LEYn+o13Jmtu2tmBX7/tT4AcepTuDzi2HeBL8ssNhdgJ
Hysh/WdjJrl/ccKpNF4UyVk6ePgYScqjBFkY0V/1/dMLYFzk1a4U2GSqEPe5lcO0RUx69Z3g6yFt
ckxwacOs3jZ18FjoE6WAiAaHj/CqvH0mXAG+QwQcbGvU3/KmX4O9INwVi1C8qK9vIMALngDQaoyD
vdeKG7kibCqrRdCr4ACB4Z7iGRJOiK2KIPVHjeAj4oHDDvq7HFlGY1ymCA6s+tNGK9umG02k+4+g
j/pCoUYRzEwhzyqEe5SSgqJqcmdzo9hrtX2CjKi2KgZVtQJTmOzIuWgHvd4BZ0IgdqQKlxB77pcy
vDLp8ul/9ToQK9h1mobXc5IFITYtkpsYW46JGdggD3UOzHh/t5OHptjTWoWyRWTFO2O/sE9ii1fF
VkwitqU2JSRpw+y1tfeLjRbp41mMv1vbfp0ImuZq4gabsWijKt036gcovFw28JJ5jDIPeIJ+OS8+
gMgCj5vPYAy8zM22J5lKskGve+fPETjK6jKj/EJA1lzlXnpn2o2ShcC+uXdR68Da5d/4Cj4XYn9K
6Gb0ogJd38VvXB3R03ghG48z4ElbMVM/a4kgqGgYPBQiP1NSaNDIjHi2U7Df3/s6kWjr4UE7JAAA
/ANGM/9V2V6Pfxu2pnwOE7b1C8GXCCLwsQ84vIuL2mtU9rmpmkprzMF1H+yn+ygS4RnBmAaewIKt
nf46noX20bruAGHcdF4+QAkn/gd/tFEOMbaTGCZ7M7vuRpflFHFgtS++ycBcUO6JcvzBRcJJhZnJ
DH8kUQ1ri6T1ApR5L7eMu1hGE7MmBmF4wVphQ0avHo21CCEUufIlU9g+GuS7K+/02voYvK/8ghCl
0Ook/UbL0paJTDvwSgD7TSunsjV3752czk1NAdugutErGm3gefDsIe8yfu6XO3krUDu3at+Y00uG
aMixG62Y0tqkYF8FMdzc7e4GuC8rCaCR1oeZdXxpP10aJnuNL5SrI8UAtJ4h8/YDBDjHRCVXrmCr
s1G8rU90zQd1rHRAUnGvUKmOfQztg+pN+ihuTX4DU6NcUFOvkeqDQNEywdZwKofaxbZaA8B7+Yj5
wSF59p/AMorIfqoZfEMkPP5Xagt5WTOdnmV3MMNoW1fOk2OVOBMpzv2KsnipEFjfj769HAj6ikxE
t+rt68XgB5eIKv0TLuCw4FWRzpZekCbBqv/J7g3Z92y/hmLAT0frMpFitdNWYuC4cqYp/ffeqVJp
INHytuhqf5oqfNQSiqC5nd5ZB6TV42Risftu+Uf6WecFCQNVMVtZmZjag5bFbJzYs9CzLcD5Nhqv
Lg98ww8m6Wuhl6sfuj2/Z3rTbMa/o8BESDusMruVbbhW2VJP4D17rIjhE/FYKxFCQeIfItQPPKcd
QEVlShTMUAfnCMp7kxXR+UVTy03aQ/Tp9O2KI494bukmRgebIG8+HVql3jGrDlI2dEcNhlrL1ILM
KrfwbkHxmojauSXR4ZgigW/tMcPfihdtNFtJ2o4n6O7EfsNeTWUL3SOZ5QhmxjmjZ2gzD+WQ/+Y4
QDnb7TfSVGvAqRr03vkrLdMdv6Y2st5lGb9YigT8nFjlJJ1CminN8vL574VXi7p0lATaS+2G4je1
qw1Hh0hYy2AYUM7BxRlGF2BqoLdihzeE8FqHZlpiHCvl6PVpclmrX9vD935NyY0yif3meHkjnCoC
3OHjhnr+dYVMy49363HctLhNPPOg7GaVDN4wc69Q0kflvnDj7OlwmHOt4tQoiwk4DcxCPgjEFvs0
KEW9iuMPzJN8HlLIYf+XEY6XaaO8wegMnNAX5uPFE0iqrWFY1rMPz9ZfKYZ04AdlrZEE/CVdJB5J
NJgPlb0Z4a6SJp167OkLotROcWpwqA5Nmf9VKwGjNSQ9HqLmL7hk+iZZ8s5LzFAQSHzk40bOUxZU
ao4pO0MC56LJGDCnaZAIRoeAlixDEVDMrOOeEzq48WZMcBfFqZXYulkr3PwPNvI00gtTu2vzb05W
a2WVASAx+LfIrdkzoX2cJ55Cey+BvLiwi+PwcNP7WlawoPp59ZSZr+vAyXPocmfiRCbqkTxYSrzj
23IOUH9zBBCvRYTZA5kpj3PAIu5SWyNagBNgsJDZdsAkshDDmVsi4kGo1iawuwCeogK0A63cnxFm
oWSTFZXehUqoE+HaFnTANaHcYacO9wNbxRfNs6nhcRsZieTSH1sZv8uaUZS9Aho+/hiMVi8VwitK
sezc7akzi3xxSLm/GIpHd2/vnzJ5paokf17wtbz6L83PJWOnkKaZTXA2xYh8Oailz22Rq8OMM3fh
jExrvDk7Ed42u99B4G2HdkGgx9DHBqf5uYHXClnCyz1ZnIbk+Lnpejm58sUTtGx8EW4IfvMpxh55
K3LinzSfJ/lkDf10Kx8RcaVKDv7Amr4vqmJTpc0c/BA2rkpQcI7DKGc27Dw+kQ1ulD4phlSdLFjT
0MUHPcC/7bZAGy8LzEtHSMKJ5pZW5pMYIHzSgelpeqePYj6yQT4f+VhGnov0CYkVmrZHSW5XAZ5V
vN4Md3nwCUuswUiRlz4/b7J7SIObxwROcwDsJCE+Sc0F/2E4RtJjAGEdGlmQ+UlXB0rTmmtNp9v1
9VOk1NLCYL7glOUZ7d7um/ArVbknQf33+0ufbj9t2HUTpF48hGwLZkFRMe1aDWjCtbUR5vEjsQbi
PaG50QLGBLpA6d565Pz/WJLqe16YpudcNv762x3PEERogd+09KLlNxSFtFY0ZzbprwCZRvfreYJ3
YP0uxI93SDl327LEvOmLyWQUZ7j6H3zs4jSXJV/OU73nz5DIn3x0LJqlmb+AkDs/XSugnIVu3fo1
BKTWtqKjPVlt548LTrnUIUAai9k7P/Yyt4xo5z6D20CTCyOB2/7uJ1pKBAeL6BTbRXtwhEG0z+lS
MzbIjGoFg36qq8zVXfOeiZCP16iYo9ewWzc4r8YSXoBDdlMvNUfTjKs4rDIMXfHQFvXucgaXR+MM
tzRXomB+T0sxitL3EJiDATjJiVv3h4eIz5uFdpu6nMnXQuOhbscdV3ZWLhxSjbZFXDYhKb+a5NtQ
NXKHCLERj8PfDYp1PmjQ8g2sm88hnfEMvrgMgOqG8z7g1atl0guFzM9crqtNft3MEJG1BO0ydRRH
8Jav/q/bqYei8Bo7VIUfGe5z74f1FuCW2OcCGrM9mCYOnc3W8u+xzWrvJc/mJ1WIF2d+t6otYr/q
SKLLInPUHM5Jjyh0FKscpNsX21aF0/4hyillLsjfdYJkM/59sp4KnkFMfRBEeZ+SCaRCPRA1EmUj
dC0yUy+KDpEJEMn2SYkWyScq3JSymfe18P+UQBEvckLxGw2toKosygVxM28OzftjgfRNO3tZVEzw
INxVkycRSZAAq8DZZ//hGxruSl7oj6HuF4F51OZ13AP9zWsrJ2BmnvqiU2/uFgn9Nnp7R0ukNCus
jjaN/w8hrN/JV91JYtLfoATDI1y+B7jrooMIPIBrcnYZhu1UH3x0ja/1o7cu3JbAsDW1XYve6ar6
ox1+UUthZ3od3wnrydzzO5tXm3npKb9ftM82mNaoC50HbHOX9CH6FZRly802ETnPJJW9gmpckqQ8
FIq/y9WlTythnoN+EgCcsYHfdVvxG/gTpMlu1I/LJ12WalChCBRnnjkS96TbBoyyLHDr1GGLFZwJ
roVe1izi9Mc++HBDU4MY8R9zwVpbsG+1566HdfiJ0nTvVy5Zw91Muh5OjCLJwIyTgYwDWJz3Y1Y9
juoFwQFimnkocBsCRFttzNAjp3TbM7ao/yB3nBlNy3lscifGy06epbDbuVwGDPAQwXV+jwySMD8p
eIkLnWkIFySoQa+WBx8InrM2EjfwEGfVA+l6yycJT42AXit3AuCjUIlKpG8X9PpSe63B6wHu0+Ia
0cJ0sHPrFVNLgbxcR4SIMED2i9vYhCF9Y/kJJLmc4q0qmq9Hs85aokNg8dF4rDVtkrS+w1ksk0JF
zJzUNiYxVnWjaL3HNrZfjBn9yhw/fDTmn6eRTRx+pLw3lgOI2R8ClO0ydaUg7FhuYhURFydgoa5P
MoneM6HQkPjv6pHNUdrL4pT9snXrUBi2u/wAOnK0F4zRgdrPL9xQ/gsWxxtZ/Tn2ZIPewJaeZeyB
s3dbIRtp0nmmj5PCh9REYeLdwmuZOCVC3JMZ9YvqdkaAM4HPv+Ql9IN7bXsBG1cjoPPV0bLViWVD
PwnWPYWRidmJlPCTL/rfbbR8f7r3i1FHsfUlf1DJ6QF1gtyZfsy551a/SGKxlzOkGmc+Dx1sIHzA
haZk8tC5Rlidz/IsLG/xHd3o2uQk+yS5kuil6ZNVKy9iViJgyTmiyI309lAguciN1UOAtaM19PHn
c8MfOzal47ZmFgw43UKT7fUCi0sth3q73WyR9PxV5jwEvG3te5o9TuKoPeKHWwPt+ZwV790CvQ6Q
slXrS/a7gFF9tqqX6nw+XjT0pGb+CxH6blaVuJ3bdyvycEBnl6q2PH9RtLiRISJedj8RXCxM2+Gs
QX58xk9Qvi0Yj3brJNz5UvPtgKP/KMErRhmT/pQsmWbQgO1drk+pY+xelwbJ5yXz1YA62nrvFQJF
VAGWnZ/pL6bm+S9ViARYU86/cJag06VHSfuTb/UotEFjMcMp7R2exorBz2mS77lFJ5kSB+UOlzou
4d8AFCphJHBZQo1ZSpMrq5V6fRVe61KnKJeILWSV40urKM9xICu8Prpt/4TA48Cl+HXiaMN+PFST
4Yk2as0hl4LgYsznlt2QXJ4P2+laYq/zSHmjzyCO6o98Q8qQzRv4TrQ6yiFom68l2Ux6GIVSYim5
6aaTZZbRqo88830RjwzsgL9tGxOZ9OPXFGTzRUQX5kxleRHCQcNVDTWq83kDlDQsqn2qY6qH/op0
QU1/dFLm45RJG+xwQhWKanzRhD4IS+Xi5PC14Z7Gus45MOKBtqig0OcrXNarh6X7VZeoZUXSepM5
TTbQo2VRNWsKtiiQ2xQ9Hg6PVoJe+4YlL+MCqY9DcMbTEDXfV8Ww2us0wkw5pACGjSuaenG+U6Xk
XJ3tEccdHlAfnn8tX+LvGGiOQkCb99Sxib2hAm1OSEP5zhJ3zd2UMd5GJtUkljffOuEsZlmD9mL2
GhbexcHzckhqgLqsnsPobDysHS/csJYRwnVdzr8gl0sHyVnAYF3C5MGgwbaYJXSVoDeqDzQ2Mk96
hcjNLp2FM7WhmyhGurynoh35FLa9h69mH7I5LffDd6PAVl2OD8KjVVnKS49wTQh+JxU2dx8zuBc+
n5VSvXM3PB5X1l2DjMVfz+tXKKQZViZr6BCCNP0EAqkWEcfYsrjJ7wbkC+unO4Qj8C057pj58Hbk
gu9p2cyEj5hZbGlTAjNlQXAtDB6PaDXWErkmanMPr4wMJfUmSbD0bWs/ntby8vxnQdwprwV1ewxw
Riz6Oriea/sPGpyLbMMJvkSIM3Ui6XOJ3FA4O1kdlFM707nPglbkFSRdYl+cR+PxpjeSs1KWtHKL
XmAXstndHgOjGHC6FoqmuhEew9ALPbKhDg+ea4ioOHqmbyKGLt1LKFoFXmVYg5dzZ+zarL34CuJZ
Jk2D9BONs0TCYv06xpBC+TWkqQ+hv4YPqorORYYOkntkj+goVe6SPYwnXNjwMX3xiOOfCT0DonH/
DEK4EDVMdDsrVR3nwbyjZ6i/AuMny+K3UaZs7mlxW6vnaXjmDNibM1PTSuQnfa3WU0q6SqsxAXKE
KRyhBz/LIO6B0xxQ6hdpF7EHcx3FfnNGMXvht8e3yAy1X+sO4mGA/jUL5UI9BumyoCeuvLh2FM11
NKuNzBwJvsBpeshQKRy/al3I+kzj1UBG+tOS9B5+5R6fAVhMVHOQEYCTfAl7nHJNJcuVpq91j4m2
B3icfAwWkpBlfd8uz3fvGERE/zEMBc1XWAR0ePQq/rX+9H2ieWNT8LlpUP1ZjSO3K1XVj5z5fN4Q
FuffEhbAINHA/+KeFvfR0DVh0DnxJRQE63zk1mQw29JRLXBuqvgU3ys5UrBINiG6TBKF2b0CIykd
v8btwscs5JhhoFE+9MOsuWhjNbAwUp3ei5oIz9Q6VX0P118yTbWHpS+RktD4bAL3f+8vrsdW7Xuw
jhdm8j1ZNVVuXRJXQyUip4Va1P+SG6XmTCSIDcEHzj2KKzxvEoKi3RRYqDsogxNAZl4CpVbLBwNP
nKh36FGiHVlw2GarumMiuIlr1aAf/vVLGhqHTPla00+pR70fplflhJfHdAT8Q/tzcf0/Z35d6kM0
U8huJfVhy5NDX0wtlIHXfyhBnJKXsGv9II5UtuKGmnCPH7FzVZzw+CvcKwV7MF1pNsd5JSnYimPB
spS1JiBAftzUL6BmoRRvsM5NlaKpfJ4FoyQphC9TdhZHZK5aVy5BSig/X6fFkEqfFCxAujwGOW94
IPe7D9g9u/UV8Jsi4nU4f8jTY/FVwWFgyXX8+wYL7XvZdkdaWOOn/0aDg/8JickXfIrr2aiZC0j4
Kzl2AwL9o2Fdh+WQkK4h/3MWkd3A40S9a+R8o7MpcOhePbybCWVIX8EIxaLTxEUVQ3ReCPTdZVbp
iurumrwo9HX0fDxsWaLwslvXnyEufn0FQQQckIstmAh33lo4V2sTlPTvOQnskImOfTc/UuEO7ijb
Umg1/krcukXY98C1h/ipKbmjhXs4+ZU+8dojFO8KaJkzan3TAtIZQf2OhvJB3tT3qtlblQL5ZKTp
uqojfkvn8rEVIyWmP2DqZZgZft4b9ijBdBgF46NFmQn8HdaFGk+brf9A+KA9apoUENbGAvi3qy8R
ARU39D8I1ccqMEQpX+GotSDmJCn9tzQWnxtfS/5ADWn/YhsRkUrIc1qAY2D4k/h0VJts6QPru1ii
xuHiaGGIU96XhnEWIfpHvhAaYezIwsxwbBASgY5a5j/m2c7PpiT3YeBW4e1O8Ex20DHwU0ePpg5v
uLGL851q54U794eRjiwmmJT/QempSlihVnwhqeQZt7HkLS8Qdh5DHohfwGC0vV0QJ2iLa23H9tZj
+3SAblAqlmiyE3Oq6T0tZ31iOZdA8umpX4B87E9XDN2x/hvoM9QEqymb2Y5lpyYo7olcgKCydVc9
nIKZOgRb1DSbJgYGTX8YR+XPtrT979VAzvknuenvxykl6/1Bj/tPB/9wj89ZScunDjFq0PMnHTca
j7+A7eW4BLK3e43im3Fza7HAjcPg1QAzz3vyhBfesHC6onv+tVcBAQq6Qx0ef49/vl9EBeJ5fpa4
W5EM5+4Sdt5dFJj79HrZWpuu1CHTPnUQ+xVjVD4fOqSitdXwXV4Tv7eIkazI1c4N1TS+AjRnHocO
o+LmIebzGMXQ9/dCbUNWUz5M5PjMVDZDcqERA1TevXvE4+O5cdDsrXMdy5tMk0NXhS6cHxg3EpEb
Dx/zyEzfEjFTcIMDdavY31P6i6Naxmr8bfr+B3d8z6fvsQNNg9/uhKSRgJW5dcWtdD01trETd7gb
D9qkv8ZXYF7qFcQK4FCuVdkRt7KasivPJPQzDoq43nEeC/25isG2eeX1xF9pC+UadguoZ4k1NqyP
sR34k1LHw1RBzLVIVQe+ghZxNoIathc5aPbm26ZbtEQ2rv8odSte4bMEim+q7GWaOYWbrUz5cbjG
tePkv1HwpsnhLvODz/7HA96uVZjzGDvy8ZL7ecl/1pcgErf818BozflF36IgqhwxmPMEJFcUkDBX
1ZRljG5nWag5bnyJFHM+F0JSW14Fcc6N2bAnSTzIYvTPXoh+MWs4VRqd41Ne4XkqgbiBNj9qgA9y
JjOdhfKQA6GxAdYd9KVNmjGPPUfNEcUeqbPsFA41vMenxUeYxjFrP5Q2zmsrAFrI9vz993Qg069X
dasItXEwrI8OOnULkimyOHM8xKvUj34EiyN8BmaRYsXYg7Uq0PCKZzbhdGPcJOeQ/9yrVxZa+BMK
fWqP+uQxbB1KrvJ9NoHbmxeFBP3usxYJmsfxkHce3iZUAMaAEgwo7OtaDugsH+6L+wyyHSM+PfB4
XVbrDZCEOqIEQG+/1JiBvDlHXChdEiTRvxYngKJ6xwFNm1mpWo3goOXM0NwOGSVPgWjA8DeuOeBL
4s9SSM7l09Y1h3yRnbVZSV3gt46/oqE3mH9CxwZhuiAIkLPVs9qvWgxwBaTmCKR1vP5Fxs0WwwXs
vtqR/g/n4HU7FDa7mkhzj4DwPCgiQdDP/X4RUaoqD6VkVUBWRiSWeXijyX/kHNgJOQQafJIXW1ep
/IWfTJES0fbTvVbz9vsIZHBSVyzvNE0OSa/rMfTeGm4/z4nVAbjidaXEaB/ZzQCFDweadwgCDOns
mHfBp8CQgYo3Vpbq738Pf6KtYpoZc8vRB0GezErFXocfz3/UbcYiay05zgqUBkzDO+/m2/yql8XV
iR8Tksa534dJoxKg2IzFzrFwM+DrtzlElctiFAllHnHLFgdqU8cVQyF9ruHOAE1iEPgc8irKrOqx
BmwkoNddlWY3KHYFT9CJXnszlZyYIUY7lxM1IRSP34Klf92LQWyolifQNcve88TRaWFMrXpCf06X
6ygtH3RFPnKonmQf2nHa8FdP/D4PCMre0GBx7lWJDzOe+dxYLMtqyN4g3Ga2d3nwKotdS5HYUCog
yiYrHGgGfK1jNig9XReeLdLpSxr+d7VpMo1YmTM/+LpJAki157kAeCg9eE1zPYCxDOpUme/EoRtq
hfsTn00UojmfdLbIxbeTctnwNF//Et1wKevmCgmnx70WlkD4nJM35uY9jfrUyjPKuQ/DwKUlCJhc
5u5YzHwA69AHVToDHlN3xIwtM/Q63VANpoVQdzXUN9PpiinFCHCD0qvqklj1Yt6PzEn539IqlnW7
YkUBz8NHmTY0+2g1C/ObFrXBkpdva3T2+cwJAhKKr4HnRICy9C2XsJKwdHMUjgUdVEWXiAVN1iB1
81+BuWLYUU5mpkQnr7lIZe9flVh2od58cABMGQxXmD3mUdzm4HyzPWtToAbjQzX+4FQlmQBWfDSe
K77v+lOaH5cDaP9rXjvuv5yE3+1xk27nv0vHkJfoRn6AurKznIn2ZkPTh9olFAaZ5ihSnflxMA3R
kKcC/PQv6fn4EYh7TQmH9r1F0qJna4q3pZ94ZW8/pwsNBolXzVcMAzx+bOGBjuS8QkSycyB8m9Gq
IwB+kyEXibihmJAzyT48gAmKjpYEcZ5hOi3VH+ZJaNsbRPWauuLLXpNl/oWP5NfJsQsEPiQRfaCe
CtGl3fGQonJ+4sDanMEgRBAF+Ebc/xTstsNxwO7JZ4iRfFCDz2EkrMVJUzFi5EQVr/llN99BecTJ
Yruc4iwmL6Aqy2xf3P865nqnAX3vs+Z7QiZmcJZ1f2QWql/wo1VOAsN5E7Ta256kSFz99CEO7KK5
vY/tXjB09fSmtXDFmC6b8KyYfIISwpe0wWVBasRsfOpe79sboysSeF8a127XyLUWG9f1vjkvjCr7
zKJHFbVOdSWB9mFWP3r6gl0wxmJW7+t48CMtRTsu/gs4qy4H7v0ZuEJJfjjmtVQkVJaSna6VMhaq
FJklobKBwIV94AfZCJKSx/9afIWS+g8TkjquKyjO6dce8kzkQqskWDxEPkYWTrs4gBgHKTWL7KZg
xnwtm06NQEEMg4YLY1XL+PmIaPUZs9Igu5gg8Zq9zK6/5uh7BYZsldijweTnIob+K5GBPhMlEDUI
zHTLveciVq6+u7+gzEB6B2uCx5VjiHwJOu2yc+kg1eNflxg3Zv8TDgWfURSrGhyXE1nDdovIVLwQ
QZHXFJSfbImAhb4LjeDftrQO7Rbt8r/pUhD342P5aP3AgA3bWKydkvxGf9KJ/oATjr2CnAktnc3q
JChzxQVtO+Qo3nk4aFVI4b2UGNRhXp1CZFXX0CzVhcHMr6W7002SJiHeQEcAkjDnSchhNdwDeMaX
2JPUryb9zJt8OeMeltnWB4+Uune9ewSq1vhtyU8Vnx60jO5CFhvZh5fm3NrriqyimkMdjkbGD8z5
GDTMymuip1wZ4vAxd2+peH+LbEyZ0zEdzeFDoJhcPqPb52qIkgt0ouuMrUy7786bOArYK/f6Ufe1
9JlBt3o3CnBQgxrfkm7nwgspzZ3G6ggecz2rLTh8DXJ7yKPrfhLa/ATPFKH40VZ0Z/AzWNDoRUaC
D0S4mrmy9GXv0U7E6YwjgwS2IQGNsrjyn90f5RoFZnsctFByKSGprRbx2f/86qcUCzDDnPjcBhUK
p4FXIr3+bfyK6UZd6AUlYzyz54iHJwTtb6184DWwvl11wBxmVPsSDu5gQ6rCW8C3tAO3jRxk5rF4
3IXuVSLSK2tQYj2j3HZHBx37F1LgWfUVob8PgmmBI9bFRQNMEOQcwNDooqiu2It2UekRJ5AJ96mr
ie/0ge/DYoKpN7EJIubIneS8KC/pej60oUYf2VAkMJYrdeh3+FmYo/fpXMRXrlzawiGOXHX89RJH
soygafUjhwx645Ytk+qROBhiR2ibIbp4DxMYLh5OX5+laO+Xt45UB6AEjio1v6ZxGG4Ppj2Ye/JL
6u7PVkRbCG3QJs+ltEzK4gY5D+NNEmjX4NWxd9zk1B2an1yy9sn4XP1mQeXjSa1d/++L0Qdd3nyM
NEHuc3D4IkAgnHIOfglZktsXM7G6+2SANqiEnYd+6hdjzEtPsLUbjULdfnv/8m/7VmdzQORvM64l
C5WIEMTafgGHhVIOJitF7XVt6koOK6W20OUdhh1Se1IdumA0MFQQ5Pj8LH2r5VlL64ahKdMssjSk
qiA7HN/UZxnNRRU3s7H3wIhKotejJ33oBQ1mQ0/OicYg3G29K0OSwSXlK4kEv2XGrEYhit2zDDIT
Ga83L3Hz1wjSg4bd2d2n+sPG6iaOwM07YJts0MqaC/+hX3ldpgIVogcVSmE13rJl+ZEB7snEgYAa
tpq/ysEN8NHwzfEONVDyxP75fFsCB/llA+fcDeGqjh2sv7wF/4uhDbwxceNvcj1N4blwEYDS2WBt
qigJnUsvXNEvg+8mCN8l59Ebo7DKr9wOdQ7Ki6qiEesDd+wttbfeuH/WIBSXJRGtzr/oDKtl8H1h
Pb6iYo2TxAbTgz0JvhwmUeUzOeZmBeE8DGriIt30PL704FlurUCwpLNaq0Gh4lGDwLC2IzslsKhD
CUQ+/fLNnXv8STTw85u86+u3DbeAMiwiyRg0qYA1mCw/wYeyZ+3NxKE41+s1X/nb6M3y01bUltL8
oTXKILcwkr5wlgJ/16gwW5NZuXUfhTwwM5VYQmACxN6CiCoDM3cHTHtQ35knOO3ivUDi1EiMaWi9
gKmrbkELKBXa7GB/MfjlH0DqrL0AyEeUNZXqumqSjNkmwNy7+HMw0uMhAWCI/+Yg6xJ+9OSUMIBK
qdIXQJvh52oNIX5LAEN7RT7pARq1Wnzo3/0iXrQN4CQZX73CCx68lsq2B28R6OGxjiiZ3QWQ00PV
Zu46IN0EVI1t70nQ9k0kE9XLSvolDcLMZUgVRdsoZv8pHgZgchsaX2kfYout5XNmty1gOodNdbLm
JhDapS3qm3hLPUxbIQzKgIK4OWV/z6rpfMW1ntdoaCDT1R+GT5EZws8nTQcw6+K6r7Te9r17OWzx
uBEK1zAYr6jZ0umOGelsetdaLPlpEowOU+lJF+X7PqjU1yCM34hliGKnjjCfr8lfu+PnXt2xwTuK
p8P8XChMeKDhJrh2UxDzp56dS1FtjmKHSQ9flxJCht8c9nHVPaSJGF8LdSq4lsFNR6/qLsceKqlD
J0gwha8VIm+qkeDDqRIrdqG3LsHv5/km3W63nv27KwMxjGMq7FNBQyF8axF22Hn1wz2V8WzgBtWD
EiP7SKlWdzREomh+/bm6MIcYhllqJKAds4JrQat8Yu04UgCBZvga62EXRbxczK0UaExdZ4oesiuF
M7SKxdQZ4PWKkx7+zZ6SMPdfcQlYIdCVLo0tAKLl1u2pjGVuIAUMXWN3aKh7uyTime0QqHAZ7F0d
xvQSqJ1u17CLYVGQqQgjXAky2eHlVO1igcyZlofDA4MqEHFPCT2ctludsHnkW68GLm/HiP/BHHtA
3Wm+YzKmML6aRtwZxEJwXyW8YS/q72O1eN0F2nJ0CaCYVSk01InOzipk75CyGdM2bWovP/uIjSAG
qRDjI71vGiFTuCk7vQ2pUWd2SL2jDCG6ftWsX/HQtKO8L3FJMidzCKrnxm4j0jKeWlNoQvEqnzOI
PfAjPM8cPkGp6ezyr4dx2dzT1o10guQ5guGfpM8Ez077G5EJdt2fi6bo+LvITY4ECN4fndMlDU0T
oiJxtnpL4XyF4Nw/RZSVMZg4I/dT5UDxULCm/YWnewoJZDtCcs/PDMQq4tE5GxPJW9acrvokNdY4
KWrNy479EUho89aadJwSWqtCP2L8zlNUgvlV+D+OQB3Rr6bHdimxHO0FXF6CHuAVcoj4ZVa1NLAX
zT/6KaHBwu/D0t6qxPQeVzV2wZFMR9j5YH2nQAdZk0zWMnjgaJCHadn5pji9kGZecFsoR/ugbqQr
W8LYbVvhO00eP1KTurZhGREPuo/9RMeyqL6r5WCtsDKqcrsQyK6FH+2su1dAz9ldw/UJ/jMZ+Ctc
dcDPC7g5AC8ncOiWLM3c/Vj8vlxiypzFP4hipvel8ecl1yCXM89Jc/t61q5n7+zi/Vs99MJrIF7r
8OfIn07I01XDlX/HT4yoCIbrCJzK0hPAXldCPe62KhHeiRSd5fvNM4F1fSEO9oxk/Ss9XLvMJ71w
JaqizimU3mGa5twOqCyphCTw5EI+M5OdBLSbpxEgh5BunlctzCz/bOg/eeDyvAM3Yl0BMVxdrXf6
sZg6YrO6mA7AbDhewO8s1HXWYE/iyXcK/pOraKrKhRSXawFyZYIN1iRkPJNE8yddSWlO6jpiWLgq
KZy23JsU2ukb1PTemzLWcWou1N/Gkd4m+eqBOtmnlR0pYM9FRlrv+OfbapCj05q6ZpMOX2sG9Ife
EfdIVAsgO05CgRJVbxnrHOLBa8uQKKpTRCfiXcRr6SwR7SHc2DHmoDeNwjlJG3GYtwNV6YbwUIv0
h0UGghy31yIRaELrL/ZGdQJ6ZahjyQ13Ar4AwVk6awzkLkPbd4nIpACatobtU/zWtj84v5tBgB1/
aMZCzQjHa5kSrDfN3Kh9B+YLt+g+t/yTKyXShx9avesdVxo6YByb9Y5aOVFBxdtu0IqxHWFJVcBG
4ek0/0KObOxWgQUD4AaptMQYA2vMPzj5IPevRP4lhulOmMO/1rRFo/T6JZCF2bXrJ9c7DvnOi6AK
vkoDGAiken6e4aEADArM9RcsfWorAS7g7qZIbCLzBxcLdmlTnEvQi5EmOkaWF8K8ZyNvckeP/ari
OYVxGori6vwoVtrSGELbdf0RO86+zCTzu/6ZP/rS6P13ug1ip+7fl7yiOnySBAwRHhkO+mshHnyb
p7Zb7G1Opx1GrGdC+4y9Wjj3qaREm+NkoTnyDYPAcI8H3NYdPXibLss8uyNDTMkB9++YQQ6fQp+S
T33f5iE0pu5NNH/hoNHje05xa2vUnXdcQrLQ6dMGr7VXGQmm/NKhDguOcujW6vbQpElWKR0RmOSx
jlIMxGJ2zbnBAiCmYWHo2EuYKGbdby1MgBPqPHwB8L3pCPrzH0GGtdeoUIBXmIciEOan+dLC2jbB
1FETosR04Mxs4vySOTsBgOv+9ePf/ZDNUGXeRJMWyBd6pStfP835JPXY9W54qQxZg5exICIL/bde
4vrhNMgBMeLVWTeqQoDDo4V5uOKiLwwaOlm0BbRXdVsEQ4ZGP7W+mfehiRfYsRH7hNyuQ2d7NTJH
8m6YYzi9fhNeiaqa/GL/owibZU92N2mT2B+UtugxyC0IKkwoQgsvnlypg5I1gEYOk4YaNXKC2AZ/
q6IroZUxPHsu/CROc6gcdmQpqcbdZo4381fWaMjny3I+K8zVtmr2BM17zbBbfdPtnG7NMduZFa7R
6Adr7DzWql1K0VoRaR0ib3uWMm2GyQq2T8/IIjB7pASjcTSIAlJSmDxaUytmwjtR6ePLhIhhvpeZ
ds3eTiW9vRxpfREReXJL6BWjhtyV+bQkUiXqnMU6maAPhPyzdG4CCb91y4iEbySXwgNZMiMWnVlV
fk8CgtK7CxSYp2Yym2ekKLIWYJU9w76LjlbwgEyo9UNsCbTBRfr3I5HKUOvQZrJUzjtjTlq3Q4wG
bhjhdDO1yZBaezc9NLGz9ZLEhHfIrYqMI3e559HMjsX3qoXywMNzGs8vCe7fSTD4n7ETjSB1rMI1
Qfpa/sQ1wtWRkLn+fxZ+ujtudam0H4dGAddvxhSYHr28Wi6TiUa/rrhog5rnh6kRsi/sTT2IHK5P
ifE9HKTOuoFu3h5aH+nTVFyubUETZ3U7yp2y/IVL4NdGcPky6cQilKGG0of0M/kFnbSvpaFItcl4
6VkeqBOlXzdP/356Pp78gqevhXfsDK0/ZKfJ0yop78XT154qBAfAI6n5RrcKw3YN1E7QUxs+Zikw
fBekvZF5D+dGtJF+U4PwCBpLHRw5diqtNSge+jjH/BM2ifeQmBR8LHeF3NlMNZKUG1KByqxLXhDz
w7mnWcrfm9f/OtzGgTPQosA6CVh5YSzxl8aOm+dtv8f1NNEeidl44vBABq3qJHJEhPZH6vTXgP3T
ZDhHpUe9uvl7Bh/0TCBYtU5zWKBRtWtYZNgDZ64s6c3gS2kFx6ux2BzXzi+vJamYejLEvmIn27FP
cSypCyAfWnKiVmflXi/A/WihVnP3mHqjHUpVUXt4Cn2biIGfKAVokO5aEl0MEtrnsYKYWFMWSaR5
vLABJtzYN72yhOquOs4oyCMEsY7gK+4iZ5ZPf4AXfwIAr0YRrxCD6IYjKbBDOLqyxyNEiDB9+uX8
E2gYyqYzTSasNJs7UxjLvgxyc1jaJa1GCTFE145dQwcEsuJ4959VdNNsohWFA+OsYMu/C7qoFdUt
hSpFAdNm6anfmg/gskauTi0rCy827ejw4mlFy3yR9JXcXUycPkRpqdyEpzisasp0QxCJHguZqSnO
qxetQUERaRfasq2YZ/FqS6yxwxh1fD78rtHjulLN//GkwaYgKSnK9Wcruj3N+qpbVXtwqcysDbvR
3Z1BeeX0uE+RntDGTkBd7rmhX1JQizqWeJdQ9kiCc7F9GvEyRpDcRfglrLXarXpoFPqIGm8vkkNq
dL+pQw9S3aa9f4E1W+luw8IHjQDgfCaUesBtEaPAPLSg9iIP5sa4QzjySsSCYoQYwhGPcWUIGsml
9oPyy8ap/c2NycsMRYqU+TJDjFxELYZbT8IrqHoTXihmhKoqkwjvZ+U9pc2HmWx8fHDJ0GCKk7ty
HHU0TnahDm7QGaCV4HQzOxj3I15tReYPjcTg6LxkSw8bnR75tRy3746U9ighf17CbtlotN8pxAT9
mAU7C6dMSbnIJkfSilv8iCyJnrv+C0tp+oTcUu8k/bhr/eR83GXhVFHw1j7cx2z3sD6VIXoer2qo
6F/fx2lEwi+j4beBgJyVsipcYmIK/PQ3pEg9XFDzte9jddRFKeGuhE+rm31lVCW/15R8aQPPLJCw
/aS9MrZx9FxHEsk93l0LTlYo6rL0eB4UGVY0iRUGfa+2E63Yntk9YHni2ojnXnrI7NDMqSNm+jC+
BFPiU6qnrLBxd45Tkc3FKQujuNTLCN/b1EUN5qMycKZzgTsJzuz7eCrp/ae8HyBrRjFlOl64DTgC
2seO7pgTo+YkJFYglKyp12ZzVfrptMYDTkXrmXF3DQuFwZQFNlg5co1gUyj21tnarBbO8+Kiv+eZ
gVJugXEYn28YBtTUCC5sL5PzSCA9QaAq59BpQvj1zhrBcqmzeD173YmL4sqajRKFHBMDPqoYU5jU
hCIUkvv570MkjsZ4BN6v5HKzUNnEO/Rx2pyRjpxF8qtDFEY67HkUDaOz0a/qBqT8V2wMWV0k1w/t
rEilaz3u5sJIRKq5NO5goFYNzLOGC7InS+YwXAhjTIdBI3gxuQdJrp/vHs07wV8kGvXFnMLAdIUo
GUrehiOkH89AB/h6jOD4DduOO/VervWqqVA2A2bWrEkC9Nb+hSskRdI9ljha59wA4DXWIrDTLPWY
rTV0OYhbxIAdmi6fNxbHp8I93HfbxbweVDxw3Puf6OKOcjP6zxXG02Csr6WNSzQGEM3i//T95MVc
qZrXvJrJ9hRIOzEm/5Yd8Jcjiz3aGc2WITatYMvHJPM3wAVQmBcqTJq5CJmU8gU+mGqk2z+7kFQJ
AJS/HA9AzSzCybTYqFQmj6GkHhtO7Rj7+ZkoJ56ZuX66o3pOGkz9b/GFEPWoY40WSfPrmv6fbpj2
2XE4ElwierQ8xda9bLsD5eqFThc92GPgH4aOMQDaQQJ3uex4ySP5gqmVbgNN3ZAe7VLO4o0npD6X
rAKuC+o3v+yr3G4cmUKEwZbpWrR1PF7eDHWl9LNgD6rCrXScBfxTEk4f9xN8oF+ZYZ32SZr7y+NF
5Sh55vkZyMovXiRvjBLtLLVXwoVhmcTesxc8FpRMtS8OY+KoWvS6V1XAO4hkphl3EBDF8cJF4niF
6LoyVd1WnR6Rf30QnfBe1Ns58szfB75vQFgdlYtB5lBQVmWoDwd7DMfeGf1mF/O4trmrhoLPbxhl
disdzSWrWd1y6JFfaeSy5zjGGieyHR0kJHANq/kv3eT6K8eCEzriqB4PZCu8VKb5l31XW8W8yDnx
rGhCaPwfvNrEXcHk9V5lWX52uvlMh0GQT5E1GVt8eH91ix9Dwpz7sbo+yaADXmC0MoyIWFvb+rej
XsYoJxeUv+Bv2+Y+KE59dKTx+WersC7ckV+36WimPrcY7uCs4WkrTaGZ8Qr9Gi//wDPDe5k6MGl1
peztMFbAcs/1G8oOxiHAGU1Mc2rgpQg1OCPd7dXsI1mC52cYTAkLQfBMv4IhgSo1NbSyPedgFUEu
8wE8BVQHTp3iosg+i/lUQoxtc3UFG4liF/978kN8Bsbnfr//TewqpuBfWfRCmxHRztXCsvZMjvze
KcBX3BHKlg1lFXuwZbCisDxAgoSniW3uI4vMphvd11ycj6sdRmi2uhcvtLwzmo8d5xayICPTEeah
PKORkWcTp/LItlbAdo9SJcd0r0H8Z19DX4PyOeH0hws/Bov+Tnmd+LAHu1Den0mvJ7+flUlSTFv/
WbQrrcjFYizHo+3BDt/6RWyAlKXYPSAO0KDvJHui1wXwYRD+2DCvKgn6LPokAO8jbUtQPIO38sFR
/fiZAmtcBsKOPO73SjWmj9xvRvSk5zxeC3PcOX2q0d1cPKvIPRiA8QDOm05eCPlUAZ2PxJe7Hx8C
rCW3k0PadVIyxyGVipNsfnaESoskg+BljY4J0F/bhGhfyNvRv/clh+absIBZMr0KwTqcqCoEYuIQ
mi5ng+5RPltvvw5/bFLw3fCdCFCsOnhuV0GumreeLQt2u0SYWgIO9/TlS2DbOIjJLZOGZq28bXSg
1u8aaE+W2Zby3aLSVDJ2Is4diL7LKestqRGA1j6ePuK/SQ3geCtqLVVjRPqxT/s3r/IiolW5+q8v
BaHDFy3w5w6iGulb/b8t0YmRu30w1wDPxnWmE3NgKvtKkzkIDpP2LKHzdbwUPFYtYzr73cWsyE8T
uy4qd6Cr+DcJ4NigSqlmLhm+KWlNS18O+bSSn14b2iok72tOrWjWc8kF/ti46FFPt1OXo2Qey7Cm
/G2nPqLiJlqtFf53XqqB9SVCEpX0NjV3LuyiRD258e1mJrmPwEn33H0k9wNBzmJuyHVbyflC21zV
PiW2HEQffKoefcrwjgwR+JEqKclsozpWJPbY00n1NGY9vVEEPEqD6TH2Dyu9o+yhEQvosZm0VXMi
YItt1ykJ2AgTciJS7+vgJv97tA+OQs9PG10+HU6bab/zvOi2AdL1yxxTsuRgktPjV2At+W9fyTvB
mYaT/oqzZBuzNndxX2POQ/SD420iVN4EDCeH4e2f9VBH+m69VGgwCFgJsxbZ0pNyBcSgQFAFHEGe
jpb8Xj9MsDboBD8lS/taKQy53YphxSgeE/N+IuLmDmxzTmFnZA6ThxmQ0WLa79875O7fRJXPw145
2T5F4cnBg1EOacm7SJ0ssWTKLy9HxI64QQQu4G9idOc1qU7HVcW4296hMZko8lfT8XlOi1uzLtDc
wrUP7b8O1pnRETYYZ8grYPcxRrZnhNfAwhHVZi2h+5OCVK9AYpeZdlqLYKsFBq0HLLdYQ9eWJuiW
H493QUJSTgyDt+YmFITXcGarSUuPjh4Hby/Iru80tqivxDQ5XAR5Cc7mlI2TTOiofSH5sC0Z8/pK
/ZkgQI8akGsWzVweCQccuRy0S6zFbOr8FAMivNaibcYcw8bTZFjhQfHuNtl7cPdJKnmE2PtHVNjy
5+YZNVlWEGDSQlD0dRYwPRwxE1hNjOWUXFiaf60A97OSACugWmxdqZu1ILhUXwIDOgY+2bC2mhp6
Rh4lPXpWNlI6krWt3knWXEIKOOf+jKdJlOX21UwHO1aIp95xllFv1vyKQhH2clbgbObCKLwdNOaf
8IRaXgWTHGx+vVEFpOC1m05XG6jluWB1KGHHhPIbwE9+SAxHOSYF3KDeTyWifsqONHW/REhw8UR+
PQDkQluZBspkyrVIXYnP+j8ADWTuBZJfB/B+ucTiKBBQE9Fyb52QEtP7KfUJf3E2IIO9EwlsamtH
s0vcezHvx0e11eHoX6s76BOdDSJWtTEXCPxpR0SzPoi6Fs2R3M9nXyukS3Yue15XkkK2s9Pamlcv
xyaVer2J63lNvr3wYFnIc9JWpaE380MDNMrEyS41GnwDBHUOBSzc+bN814fklKKGCqkDWV+NyUx/
G+HF6y27T5mWa8kuRggUMSDRnhWnwRYhTQUVnDpoOZBLN8oLkrN06jU0Z8Iv08h/esbfnl/dC61x
ASni7ATZz5Yd/FUA4PKyII6G3VnR8K6+6dDKU7mivLgqCWMN1CmC3qyFmQjVk0a2WwFEFcQwb+zD
sYwlqg5UNCovgoiKSZHYAseO9zmUMgHLexb7q3nHsbF6hwhs/0Zs/sYoeMbX0uwkRNT8y58H31oq
U9TYCmSnVlHCOCMXzu0D0y7jNE1elf6Iezlk8cm7K5w/TRySWiP2WdhQ2k1b5TCYcl9zO21PqmXO
T/LnU0CcJ3xBBHz0P51zkcBEMKJ1z+No7DuIoxRt2hjcHduPfOVsRi/9t2FEWdb4SPnN7tfjzD1l
ajSxAIDRzyxDo+esp5EAm5CWqB0zQuvA5vPUglth0atWPq0p+/tf4Yg3ya1Cddg3R8f4yLP0t2MH
vMgswem9W4R8FUM2HsQuZI49FFA4JIgea8/vv/PYoBeJCbNY4jKb3kUizZ2bx/XC4Fe3UQ+DTLfT
oDnok/c4b/WUzExIyFGGIjA9YCrmsH5CyxCCbfbWDL4ksf3gW4EyQpqv/SfY2VLduddaGuzLYlyY
RillOLFoGyEUtHiY4DU5AAY26fBGlVvb617QBBm3xbjGDkKuzEy8nqLjJvNEKRUTt3FHnwnb5oCS
xjd6CtwDgdKI8V1SSt/ExnZoM4kXo1i0ZDg/DQ1cZIIYxgpI2NNucknqpZIPZXnrqzOcqwqJlIvS
oRdPkth1ugr04kJL08dxwqcvpylk35QLdTfjx2JopqHvDX2Ta6EMNfxJRFZzMsobC3GwV1961cHZ
MHa8kifMYUmUw+1wt8tVlY9oz3ExfLrIR41ysemKNDGjU1/CRXwsXANo2rDdWDIhlRvXBpBMjh+0
AI447Yj5YAmTdLV062s4TO1GWOBy6HTE9i2UfYK8foNdngtpdhx3P5l66URm/Vijj8EZBA6TbLOp
sxOq6YDFo1Le9s3Ajr7LoVTKOWARuLAEHuXBA9dLqFjdZsNn1bL6retfgA1Vdvc5pjUCHxei7gVO
Vr1J2iwkjPDEqRFGS5N2woCWfMxlZazQZGodr56ETVMjP1A1P3IsnVfl5wFdIPG/lPQOiulFB0pu
gTqtpc+f6z9j0VHVydXEBz0Z81Gow1yoxKE4m+2esP4kwTqzhVotxGZf+x56Ak63q6zceItFW9I8
Y4A8HZiUjqm652ubziRW7ubylsFswHyqoAAtMxoCB6er3oqDYdvn7snq26/EoVNB+iV7Ych67bfH
rcDU4MA7Kll0QkREUKyU4zdJ9rmQSvXa+Fc+AZ2QEFNeXgpGf5Kcu0Qm3iNdc1wOdQMimmZTjvwS
7ZYO0yyx3sYC28cYlkh66T6/axUQJC5UAroRJGXcUodAWsxyUjPlcwn9vFNpA1GBsfHsy4rG7CHQ
A5dZbsM5T1qS4p41Wt0hpH0Voj05kg3/pU9/PDB4U/IRdhdxwrRqCiDdGUJgZJQupWwzgC6ymqHd
zSpEKiA8xgFVCXphx+KSFoUoP/aLy8BftGTaQt3Hqd1eZtYz9dSDn31YUxvUuy7lcPYOAyzCEqie
pG4C+u/EbeXtcQKc/DyNOBX0yyF0EEMx+mOqKaJ0X48FZ5TMjvdx1KTVbHzghcepr3A0YteNazru
lLuimhVWwY4bTck6xjKinLm+FNBSTI180GJvYBf/Y2P2/53jEj+a9ERWi63l+42ozXQIA6aqNTcU
uJUaSmYwGlI9d4TKspkgElJd+dcE3pJXBWqqbCzd1q9kahJ5gXSZqA5fd89IlS8VCRJCLBz+sAMS
5SMAVWtQcJ+YfzNaKnTgjF08LdZU2mayel1py6x6sNidelBRQnwvhDuRJliwKVuKvsc1EDoOckG6
nmWcu6cSZISg8daRO2RXFZRWGtYxfnFEBWYVlMrr6MecN54sF1hYHRANVN9eAAqFTov3O7bIBvUg
jm5VDGL5zFF6+4JadKeAjp13yP70Ubo7P/By+snpAd8KHNImxGDQdikM3lCR0oINOnwCJac6x4M3
IKNT8ZJfRdPZ0fT+jtfY+zigrzQeXTs9tYLBWBnymBN3XWD7B3h2/pFIFEJi6JT92TJvDJDtfnwh
8HUaGa65JiyH1gI2zgFo0acFmUnclJDh4boCneG+klgtlux+HTzh/u/ekTRvUtTm419cRhRy0avO
6L1sgwINP4UgSYM+WZnj9H4lnTshX/y/Y4scGmV157H3kRuVyo+j5MtukWgSgiKjCB87t0Ivtx/k
EhqhKy1Ict2YdMC0yQIrzwtv3SFFYXx2JWcCpYJbG8UsjPeUsqek0n4KKChCDNWlkwWYLHygW4Nv
bFZcbo8yGQ+67U8sH2z52wt+apqPD7LDm0pqCif3VYjmv0C9LWW7TbufPIQxY7aFDgFhd0mDYYkT
gV5W2syAiQj80yLyXz47iS0y/Zw6MgEuddnDPHYuI34On2+UnZ6uWJrDEmseOtMBELGJ4WTAuSZU
F7CMjrNZpjqwoQEgwEqicaOzbLadZce+Q2GkqoGsiX9BsuJFyUky2zCv6PT+bHL9V9jxE9SHXK9S
lo84HL2Vp229B8xfvf+eAx8bpviyRf3vUtrFUKNJvIzXAUgedhAd9dGRJ8PWec7YYWLxxC199mK9
Jjq/ZRZXv2Hj+eQFdNRnkkxnHHuyPkXIN5gHoCv7f52EoopzvPZxrX5sJWNeV+YH6CmWG/d33h/L
oHe1Fpfp8bwKVOUoHvj+kcOFFMZUTNyfK5WQXw47aS+eAAA8JKwC6xU4Gdt5ZvK2oli1/HIO8VkD
0/fRNjGBQfb805NhjDCGe64kTl8GefVit32Ip6XcHk/S9BqSBeWLSu9MCDpdMutNaIY2vUokVITE
5QJIHBM9LLNCKhGQ4WYZAUEueHj9lEJ63q6C9DOIEGXaaaQPamd/mTeCgINU/89HpIYFACYVTh04
6wYbuezsp2qAHGOm07YlRMAV7BrNZsTUz0//A5mj0iYxp99CEzrgn5UDtUHrbQRntsbjTg7ilCSu
r3rJp/PnlhsGYqnBzSvtcksQUTPVX78H/vCoGFDNi7f5J9tmIAjomdJLPx0Jh4/Jta94LbjgiTLG
uLZmdxrvuWJw2+IzhkU19iZB3gj5KT6Emo2x1Xvp3iev2RpPqw18vkWmrhMI67pk3l8f/G3b95MW
Ga44LLcneU03DqSMg0P2cqqyV57qMzJOmW5B+QoGO3rRtcw/ScbtwYZvbsCXL3bb4DHikQsZ5V3N
y9pXSssNmemsnmkq0KJjc0EWih8ctJ9hmseArMFGCIBzFPz/Mhc4UJaeSmjQt2FU9Cu9f5lDyRrg
ub3lc32rrVKxum5pl+xnYGYE7aHAA9Auta5/u81HgdmxBsM3mwUIgs3GGCNZ47lLOVYcMlmNAqZV
qgEcxdOdn06BOHpEW59If6LdBjITqRkN+nim6eVdL4Lu1Uz0izWadiUK0qUv5ztWNdw/6PNbidb1
kpS6Sgf9EaUO9GZM1rR+8SjV2oDv0mEGVkC8L5Pol9id3EYKTlUZ551VGChpjCMzvbLYlm4lBWew
av+sP1YMu7/4ei6c0mDw4Fes9f8i8VdxKY+skyjOSunBuTlk+1+uSdVx95be+HCo/KYx0zIMaWXV
/5VD+9UXcl7oL8cm1LGFJIBE2RZlN3us/RDTQ4ff+Jl5NAaLTItvwoUE/sxYIpFjajDhYOqVz22s
QacQVR32UQgmCtw+McMQ/+UWA7pxlXvAeJAMw2Rez+N6OdAEyf0X5u9Ntj0yahbqsihv0Z+WB4eM
olJWk77iV5lQa84DmaMrspDy0MF0kzNv1+8Ewmcr88NtNa8s3erM9if3sxY69lVS5h5uV9isFEXx
1zkQeGmlQwDkC8LBjmuSGLgPCwGrVTpFmX899Zw4J14zJGA3l9wy8+Nja1+E3AWQdWlnnZu6tikO
FRG33ZIiC22jn9VqT3FXvrRFKHl0MJvLW/KB7OdFaiJSEmJlMT3xE97vvX2Lz+VryvOuswKgoWa8
zmx1pKPWPQMtVoChwIp+J1UGONGRNS7RZ3UlTFFwkk+RYqsYlQ8MmUMDBaA5u6Dn5o4v1qfeLLqs
CqxxXEVWpdl0ol1eTuf9aNoJMR4ZOkh/9hgf0DCopcBL7S5rdjyDGaYXbxOqf1lNNS6qSk5zEEbZ
cFg4tD7heUyZteN3IbhKL3Dxyvv3gCkiQJRa/fE2iWhY4SmtuQaNaxmc7OR/gG8ZFuL0amQAQEJN
uMsb7rj2p1xsUg01eneMtQvxSAcrsZSLTcs1UR5kyyTXWSjNv1cyQODEBxeXuhJDf/CfPmBxVMy5
OFsDL3XyVbYeDv6LQYbe++05Oey622P1StPXpgYsLzE8A1lnSgux0NKadzxc9TQrSo8KnKoBTPsO
xDaLFUD156OXgm0Q8xaBjmoFX0aa40cF59b0tyPr+REHcU54aCcfNZhQr8yzuXA3hsNpCpNlUQb9
xR2LdSP7VllKQ0WIatgCuRDV10y0ZW5RxR9Z9SQ7qH2l3oz2jvmWyIi9p+pbBJ7yRwmNt/c9/iBG
bpZc7OhiK0WfmY/MAtonRt7TI0Fk2FVl5itrJV/LhwIY0UBX7Q2Zjg57FbbHJUBkwoe9yiBw4d2E
hVzemd7VoFR678PweFHejzbkRKAJZMKr5VoB+8a295CB1J+zzloILmNTylfcbZKc0yeuWEaWqMN3
aecjB2QwDdnskmO7zkHvN8ndzZfyE9O2H9E3x79JVbULLsZ3AJnHZ8DeHrs/Mjtkvlg++rNEfRXn
26Md0M33nRmadWJpU3KVFCJXF9DRsEXkVPgMm24HJv9Cve9do1Z2nlUl768B+RH1l/xaNMiiUmH9
+kX9OXBhtKHoSyyWHes8tidhW4LFl4utNaDsdTTPf5KvV+YbvnxQSwF57Vgy/PLquXdM/6njVIty
kKUUHYsTW5qAb+l9hjXwEMtCDtgwI+fTM/OyjPkQcHGyBKImB0HhMAv11ac//dXjUkNGxOJlryLV
x/Qkq0OwtJiIwyffy3oQtILIpA+BuRfDmbEjJFWvr8CYXaDYWoV6+tTG5GX4QmWvOCgKQ+rMfYKA
3C3dBdsFinofUA8jDWwekn/7CUwWQJX3Rb11k7DOmLFHx+FraimspW+O/cUzzwWBCzVbIQafVRr/
fTURLQ9Y553qIlGW2OuvxBhRUP5fRh3j5ePFBRkl/GA2xnxo2iE+hlLI9MDegfM2J8SRVY/7SDRN
+aeZXkbpWeHE96wbhsorPgk+P6V2yF304f7y2cW8KQaO/+WDKmQHuWcWzbFWJkhMjQb5Vsdpb2ag
Wb0QYkMB3Q0eQLztjvnLqRdA4Ayny5frjVG7743mK3hWeqOBzL8lhwij9Gl37xRxz4D0xfH1BMg4
rWuLaBQaJIL0IK7az65gIthvz4QjbcEhfZYnFL2zmgNG+QjdaDuPbzOTfbIf8fvPbcpNqqgAbKgM
yGMj2GRQy8GFWnEPk9LrJbjYvk+rVmEJ+hd0Yb1oBEu5gU4QIIJc1SdTyLsm1Ye6zqvfuWizSLiP
qVkzvXUHISTu8zZF9UJb2Mt06Pfzzdvmgfd8YYetSsaKiBKa67TmvXt+sCGfPTK/eedyPpr0g8Na
Z9PZoD1dzf590+u53+a0lALVpPuHZUA5+ytZZQo7JxVJqyl6kyrDn4UjXvlNRgSffn/YDLljIjTS
qrqjS69HcaLjHyQASxMzdQTrIEVCAWJRvj8ZXhBS5bYMz5TK+3YTXHtVnv+ePwVrTdYbhNx1oTOU
WcS7z0hDmYP7L8xrQFo0btilSfPJZa6xeypqrfCuzskSdU8EQ37jTVOoHOhRT0JPUTljzDOztiWp
96Swf3Kp48OoJwkekm5++6baKk6du3dX5+V1y6heUIS4psmRSr7T/cuSbUpdmQ+0eFdzzqeIEzQC
SwbKzxKD2Pm/l8zZsZ6X6qbkXTyimiy4vjdmRu8WKmnJY50sgcWRgGn7z6Pv8zIVeJ2MVjzMt17A
djNvuj+jMZZBZSbsqH5vp0gF17FaFtNCtFYEiBANrRH/494rP3w1eOlRIQuVVpugbnHug8Ewk9NT
ZP9AwRc8fwwDeSDsoTtuMI1Cu40TEs9SNN9nFskzJkn+QukcQIByvmMdiakeAH+Vhgg5+bmCj5du
EUu/FQS48wxzjOIDxh3i1LwZudvjZIiZoK4HDyMj1aR+ovRx6wh9chHG1gEbyY53IKAPORb+CBTh
sUVpZqX9nfxE2Vhjd0T/XcJfhYAbEhrCYjyblqiTr7RNQoKPoWgesjp6bAbiwvKYDJ+X5AhKV+zn
lWgJYDMdpMooBK8Uj6U7oyI9MNT14MDxg40bfp7kKePZMBW/8Mi/ZQ7u6/lx62+z1EeQyn/VRcyL
YKYZcF7OI4iwzowmFIRNvpLRDYryV/2NNjtnNOSyWabEEWHpcMtaSji3GeMrGoqVeQN3I7aCKLNy
ColJhBz57xpQWZCoJOOjRzrqghtZf4N618QfukE50HfQfp0kVRrNvpZqTlSTqAAOLskHPIZ/DrFx
2cCbFIHjkFX/Yl+xgFiWrC4EoujFWlcfirmEi6xMsD+fUOV6VGK95wONFlhpHKuoGLLsoKgMQ9ds
/Yb3ka7iPcQOvrVwiQCqB6fo/MnZH05UoKQ206qjzhIGcNWWj+brjGOvrr/u5RsZOH3RdwMhvXk/
ZHfx+tfXt5jA8bK7SBSDMoaBUGnJbkw5joJ2Ox7pQ5SWaeiIY1I0vdP0bx8xtOPuaKu4JV29EcCd
5+d+lorNYlTCi5Mxg1xelcpqflbc2ZB+ZiQyZRM4/OfqOkXaTlk4+G4T54f9kbCmH6vV/tWgkomH
t25j6jJX5GZzhplHX+tBz/Lvy/vqY0UZbKCPZUisvUsAj6/hFRlysDXShGNniAMVNvj6rGvkLPsu
eT/t0STRTMmUITBddFHo5QXtn7owYzzaF0eF3iaXb7HJO9/RRPLJB9ZuD+H69XclGJxprbEv0ywj
Rp+ce2OUHO7x7ln5E9Gp7KcMKTGF1GSIvnLYPDe5cXqJCi5yYtRXLqlJTQ1/YWFdcsS60uFkn2Ad
dtTrISr7HWwX1InSUHiSBLZ+QNxxHrzgYz9XnwTOyKQ/Dl7V8PaH6jPur7QFPnAF2kCmIko/9grk
VXoKkwZ5ZZaHFFWq3GBW34Ntj2GjorAEn1cpuQfueI5UxlUvAPma3gm4Kyy3tFcDcKdCuU70BwT7
h3gnG/UPN+A4J74X4TewbIRumCVtrBlgsxQEG500J+QHWQqRx4kR5DKYPok1vcdWBox81WIAIq9/
kLTGlWjQrFaFPNGQrGpC29y5EEoI357X6JSA+ph91FTc8oPada4zhvRf6zOb2o/1owIsI9caLFri
VExyWLruBduiH9RMBfIXHpwYXGn+zuDBd9ejk6P+b3ttXyDvouBQKfQp+4xMWCr1Ikh80wVQRm+s
IkagMZ9/F32sKYBEyPplETGPbcPSLXAI8nWbxhdZWYxEIl6HsKkv6YlbXaKfSYGKZ/Y4pH/TMpGN
OlSaWFDPhfjVd7V1VK64VeWsyyqP9aGJhqP+k8kmLHnoxKt5zxlyoy2PYB1y1LV+Rg5vOIiWxDIL
bZaLYnpNx/0a6xDjT2P0lTqMDCepkuMVzlM2CxpDpLfROBHW8PNVFufolq0KpJP57PhBQgf1EpKX
GI/9pJCtYPvstXE6iuL/k9bOK6TtMHI7shJNM5m0P/CkGvZZHu/Nz1DqL+txHvTUZrBciTUGYXkT
mCcf4NjorOHm1eUtsayHf3FAO3dWq/obHPz7C/FSiSSiXBnbmhFXLoSPw/0haIl57vuFWXTwInfS
C/jGgmaVlEGJLM5I083y1EA6wAmNcV4TJbNuarjT+oyQt5CxhQr1FC39lc1acoTY+H9ZZxeJiXww
dI7OAl7WZ5eVEGsDKey7cTk2gMK7z4jY8FqGwhQUHVvsmTJyBnFYAkQxs0hh1j8WLDw19/SPsxOo
EpmO3QN6ivyo1mvtYwfnoLdNCXGlBPXuNUwEWKCKnec3vpE9LrdzUEHsQcEZIPVUqyGSx4i0Ggch
eeoP6e6B8TZXFaO44XYM+QVNoc1tVPrzkB0pCRJM1zqW4jO3KTkyTq5IQPplps4KcJMjS88EBRYp
J6BOsMWi4g5GCZY3R2uu/78zpA9PS2LZ4Ts6vEsT44GMcTJP6B1QUtWrENXaU/S8yCz4TOoKgvyj
JRRXRLC+uNM2BHolfMStCdrc7ok7co0UCOuslvJfVE5cFqKVrYu0ip+VjUcsR3chzU2TP7diFqAY
vB/zEBElEcoeqy8nnalHPfjJs9Rk8lQ5/3So/vrYJfjC0I8FVvQUMGLG/Tq9Pg7rIvbYVImdJB6l
N7+XGQY4hK/Fo0Nqew98xF8tPar19hG5WkV7Ajsj94qtZKggG+1TZJ8PiChA+K7Lk2c9Xkivk2Gz
THmy7StE9PqL8oIvO9gRls4HPgxEk62awxQWNChiR+geXgCaUkKaD///1k/TvHVkjt2x6RPpbsE4
DotTloqRQK5D5419WmgRAlrIuWb8Svvrl9/NmxfhcUJ8rSHdfPSPaCyJhFaLwgq3Gmeq1rJ3gDHQ
ELwPCH6njTnLp3nJ/F5hifGqTpQ2QUbC1/jZ2Zu3RWvfgnGk5AgoHRIAkDkumo2G6lxg6hj7wXDC
uzjbRbFHQ+AwXjl8WX/wrIPip31K1f0dXpEnhju8XmtT638nFTvbiW1cjpZKCX64iF6rcyaU2ex9
63wA+g9Wx1gqpfCX22YmNOvOy1a2zRy+uRVl5jG2AagqaMLv/Q0WOKwtIDbcbnXskOnOKQFycaw8
xH7AgZx7FybUbBImzV97MiVE6NAtias/n3s2O6HriVhI5EUUF2bGn7cBbCytG5L43tjVTJaF7q5z
2V+Q5nMcpuSTvJPPDoVWEyfUZ7sZu0hxjRZpZif0zvcwyQZSF722lG9q9Zch7oEmmstGGZ4OQuI7
sD7IjS6KqDbmuaMQT1hO9u045fdc27zvNiijurfZBjSihxzu2QeDW2v/f1KMXWOGgsAOwZTJa/+V
6fG7VZMPW7q/ru6T22IodLEkoRqN6S4WduOcJDd5swYGD6UyLBXBEWH2tCbgxcoStmpDeuZzUiSk
u+k+a/31BHPkHyVowe/B+Dq/sO33ZoR72GZWQE/6JFtDI/fBWHcnUP5SCSaPHl2i2HZEEF/JVDfE
QS9LSwu9GMDX55nKC3by7Cgmw7IP/JzX/XSkE3xuYwzUgfdue/IokV73g8Ph76brwBxD/7M2O0N5
b9PtjT4tgJJzZdYT+DPr1kyYLCAE0PytFtGg/ePNrTBf2HI74mrpdzZWVPDhuFyFyjLS7AnrH6r8
Q/fJG7fshs74qGGzz7dLCwjukJF9tGmtQx/Xa49Bz3T6+P6o3YBRkLWyK4G5OHyhWyj8+7Az7UL7
g895Bj6B2A9qkxkUwTeFKNASQ4yE8ogNtFPdWDv+bP2UEBCHJkqfP6WOLFI3SwpnTaRhmaOprKpn
kRYMO+XNWBY1wY1w8cGQkvcOpktb3Kg9nKc/Qr3fMvrZplA5x4Q5ZkhULwdD1ZtKDt4Gn/AOdBKJ
y9S6owNRVKULnRawZ/T+YFdzT3Cuoq7BNzkm65wsmb2Z0oJGjVqp81nPU5ZzbWHXo/E5w3LpXv0f
mW8qeNQd832JO9XS0O1ryR0Xfk+cGLLATnaYnOc2W+dhzL3SCz8KltSyeAuL1Dl+0NOOz3aA32Pa
6S8y652dWv7wKLaEW6RSl5VQVJNtLEZikyyoi6Dtzolj6oDT0zImBIVfNC1Mcem+sAL3lzqavh+k
Qlhz5XEv1fD3QOFfKVzFZcFtH2XRTLg1ewAtRYX0abF9L37+TQTzpxGS9L1XbZheev0OaLv3hNgN
YT2sju0slirZ0K+Z/dGenyiWO06clGsM0qj16ZFcn8BoaXoSKkdL5m48wri2CYioVcIrLAql+CU2
ceLKElK4ZUVA6x46zF/mJ9cf8v0A1eY+jroGC/M87M9O+TydurylLd07DWMuOg5Y0601eXP9fSP5
KZfyM+UqDR7nTWi6RIuwZHurJvvx7jYC9joJaEb7qAKddzgaZ3zFyjrCEKtpW2FK8f8evMFx9F0g
I42V17nq0qMNghSCfq2lXIuUsCKcFJvBEj9lFApCBCdgBIzTOF8NW0CkcTuQjAHjMVBQ3Z0l5MsR
4GwQTOIIqC0H8RlGvA+BVnMjEoWliPd3wK8B8ZgQsIMJZ6lfqaZ/UiQnZqA3W+95qvw4n4zz8DQJ
ZuGkxSavyJI/zbkgXyiNRrvzP2c8HKTJZRjlPIQroNCnVXGp7UMwWrXxQ6jk0KFaJPlnYyzeb+EG
dELl9TnDoptDPn8G145Brrf9yp0ozz9ut4sJhgWdQrnytgixUp1k7HrgBiPQmL+hmPaCZh9wl6Pj
oqYE8q8Lx7mIQodFfQqxiEdyGHxNQSGICaqKbCRIjrYcrDWTS2/3RtKuP/Px3A6kNRoWscM2IGko
0JZ92vvg2glo688PXIvMpu+5pFg5LFmo5olvTcHrMGt9xahpnll0n5aLHCy7Yf5SO766P301O7We
0H5j2dSsOCY76m7BS8EoewTj5VQa+w712NwTpK3+iCRb71/ofUHx+vEsRISzMtaVc7U1waaQHLrS
G0E5KdOcbLvg0bEdr5stJ+NTDj+t7UC5T0AMDpLuldOrwKadQQULtBni6/xorp45rohqBF+J3cla
B0DUdMtz7SYsJY1CeVurP2Tf1mW5yOk1e6JA9SGVMhEYKhHVsZVA0PIx6tQEMah32NC5dzlgp/tA
BpfZcc96CewMYA+Mo8WacSsWghtlzAoUc+eXZJgLxnkCSjaPHA1Dv/cgqBFezHgcCOwhrhQJjQMU
GiYQo1fuedpFe0ifEMwoQa1ORmmrHQV3ABJlh9DuhE2hDPWKG+aF+PuAMG9sJkhIcrDWpYriVoLm
e+DQRwq2+XIvfC28ROLGjd78lIo48ncfWq6/42kt7q8mzUsMRmiQT5/2Uo6j0c+7Qq+Llt5AUekn
LStvUGIJ5F55FOkkIarEidi7QKu6hhSinqovb8h6nVavqUQugbOR/mzsXZCh7SCnedk7ShQNj0WJ
oAE8g9/sKgQ+wdzAWvNqVzXYM/nQ0kxbAVrhFh42JpVuQZP9FTrRNqIJwcvCG3h3Hnaw7K7Q2NuK
hr1EzX3a3C46YYZ/9Za4cKfKftzMyWh8DLKeW9Ef0ZXud5XZbOTsUBhKTFjNzt5Q0kLcQ9nEZ9Ae
FbL7dXoMDcfZ6z0EkgwB5wvRnAs0gRp0i82WtwmE00RP/sjag4jjGoJvzaZKzYcbiHSTgz9HbESw
PX0pBQh68+NdpwyJq7rZkDWNJfg1fxHqLq0UGZmzL3pp172znGvN95BYPbg5rekGWxhtMhIlm8rx
hPYNrUdn4C7M/vBSMPOafzkyWrfn9t22eXrBgo27pQY7OrjeMHE3aZ245a9iJacTr3Ibmy2HxEz4
oVorbXGAsIVeowEG54Yy9c4n1RtLCJSIJ3TmTyvSu0QxFr/78XAL1lSefZ6FfBLlQ1vz03DKAVJc
TP7zXLg2TFeVKP/sOIbwtwovdSYdUjsivl7wYiSL0xYfa+zyMd91HxxKzauS8s51XjI67t7QiQfM
f/HBaR9bNWLxRjHnYHgqJyVRoK56z4I4OSk9UpRbormv08eNr8xyZs1B0LG8Mjgh8Tmx3foPXGtk
x9XaOAKQDNBCFjjIY77bi8rFOSNzTmW7AJRcUVfEajD7O0++W2yk5tJq8t2I/JVMdTy794kq8sW6
aUlA5yFeo4+MN696M3JO6BFI0X15B9LKt2J4hB9s1zZUzpoffoJqF2NLJ/bVFeEu8mKu+8IQApRx
tLk91gUK1Cfo3mAgbisWSZnk71W7lsjrY2MdtsMfjdncGBRrmOCmhf31fIvfVhFnTiCTIZBfWgbl
R8ZjfyVI/jw0YQ1cWeJhICouiqOpUsS5v79+Evf3yBqjLJTtvOrgfjJCJoar2PdZNwKT7rCzlHJ3
D4JZClUvacDAHzlwKGCx4WZe1IJHa04V740JwWnW4CtL+IC861CDgoFaOpVoIIkXVPpXGqA4WqUU
hEqOlwrlQZufup8NNnS/WMD1S4ixqO74L5yEZbpIWhQllMbc1Mmgi2QwJfUufCVwfJHNaYYP2c7T
wivNZrPIARh97CJHWEqVpi9qmIooHn/aJkUjhPOjJmat7c7eAoILYU1fLtBlPeChAru3E8NIH6Zb
Nzl+X7ucWRaeHzcr0iR+BY6MaVcttND2/26+4Opxo+uTGiwRq1zv59tKBI0QKqviTtmbTD0Pv/gl
vp/zeQHucnEU3CmgK1TSxoWNXWsQ2viVZK7ChGNjgzLujQvwWuFxA4LlQwPNcxPEswxUoVshiu2t
rGCdbtvQCKz+0Bv97Y+n4hs+EsGt0i4zX2Dy9ZrmwsBSXpuQzFG0EJy6jsGjjMNiCzQp+4roAP8/
IwdIZqBGNGousoRQDIXPhhSdJtHSetN2qkKmMQVewi9xY04d5Dbm28AdQKTOvqXZ1VrCGWTNy5Kk
fXgewuJXMI4SbGEpcPRmp1srj0SglglkUi+YStGqxiDOQCAC5cvnUyd8CVKD6l1ZQq4obvQl9Vt8
NerznMOkSlchQN8+NSAXYh/BkKUbWJp8B4gLxI4wkg18JOJ5SuO6qTHdbeE1lJZLAHku4iVjPvkY
1XXIdOhW4Fl77gbkrLrqy6RYZm2gqid1cfJ8bsi/g4rulRhgMFVcdgOQ3kWn75VFfh3jx+cW1z2k
uRqI/Faw/5BIlcqviwpisxYZqxU+xj/pybzoqC19Br4ITZXdfZLtEnDigxSD5Q2S7t2RjbEW+tN2
1t/ryE6xRavmouE0jEBZ3FT7Wfx4RQPK/Z5nkw84zerJCUwjcIaQMtlZ3eA4dDXAz1Ay7KXH+Mli
BVHgHmdUtiI64FGVpr9N4JLhpetHGvgt90iGQnfCRwLj5HSNsIwgYATJpYon3/oeJrVvi5vdrSCX
NQ12QikRfL9pNZ4JUNdTsXVr8vM77TNWL30cqnvoLTS+ueukGu+wVzNSZ4s+TqFD3miWa6+RkGPP
jEOas7hnxpQQuxw8IaC80x6OI3pkKVlXNr56BzOe18gyR89MqDj0J7L0dg94vy8WjGSr5Ghc1Fbe
l3s7C/ANuypMASdS4b/9XBNQ8dpf2uf5b7lPc1R1BGVT/t8+8E8ZJ3Vj18xd66rmfYJkHa4KQtJp
VH9hYVSlmkWEKQUYKKGLtX97GzWhINtJuS2ddwnEyOgYhNhoN4NpTqgPB6tz1XCLODeqCPjD2s02
exucXLS3nf+QRyXRRZuZmJyXpyuy73tsvjn9VuSZ5yFV/R4Ms2iI6qacapHhafZqseGP2DcWii5t
uzuXVA88CEFaPr2Rh4qE7RyuwKtS3KviDuSk47dNQou12UiGMV7DIWwCygUFi+ybwMVA4fXh5sk2
I4R7WanepfYkeZui/PWpgh67WiQHvx73po6SaWqlJhhA8dWaHTQy6orS4aH6NByiKor6zh7BSYWt
RcpU/QkCxBSO+CMf3xGPfxlrw79JVKZb8gZdmqNZAvHeM4hz+oNJUBEdU/OjQ3KKUIfrjPXGD/u8
KduPNVMo7M+KpeKfeOlXeUzR6R0Mje+um3jUnqzPsCbQXAzr7ogaEMemeP16jsPJz+wyuIrkgbxl
QB9CHub0U8pRuK+dDg6LZpSo0QhuLnCgraVhy3BZDo69uEkYxyZ7Jxs2X5dJAUGcXS5xCWN0+nL6
s/wQw22uAwj3BfL0bBRffwr/gXbU6NA1qx2Fx+fgU3Amx2QDkkn2AGiotu4JFnhPls8QxoJ2NAby
9b5zGSpuxCp18U6PX0Rn59AMzbixL2li3gP1Pi4+RTfKr9pkjLJP39UyPsfB7lTGZ3n/R8X6h5mv
QyU+eUSEAfhoTX1r280zFd/QdChC5SJRiqwoolLCEpgnup0ZBPfI4fD9K7QL5aVZMZi4zHt8uMdY
2qJlpCiEdi+9TOX4gZ843vnzdMyGqTIjuSm0YJ7ldeXlK411STXcIGQOuITmxIqjIhGts+TNyFsH
atp1zxKESkt3F5kbcBYilyGkCD+ltNShKLzvLLqgG6GaIBjUU2KjwMxrFr7vEt8uufIULhSALTrB
kGZrWF5y2C38UoQ72Erjlc3qRzZJZkHt/hYV9S2/UucNIPf7VJ7VoMgqIwf0v0P6PmgosFB9EYlD
Ly5i4uwD9S9i/0pymLGbZxfE0wZbGPVTyCTEJFuNIdOfTylmbE26Oafu8mHeZx5+Z/c40QtEQhxm
1kkSGODbn7tCLQCZVqszSGP1jea0IDd4pzdNlNwZWmaGbv6dJnC32hSYJKHtTC23e+GJrFrGGBk8
lbaQaZxj/Cxyt7yboo3zesCv9ksxN0k6lw1sx2DwkadwBLEcj3F45UhCUb8nswTc/HMmAkBqMjEz
NCknM6AdVhmtwOQIWqx6PTQE9oo/AKiwp9WIcbRAFkivDpndyBne9BzQfzTTXZYoCN4Uj57YaSvu
NIMDSQ/EA3XTXeV9/RFqZ3tbeT4nyZYLZmTzM/MBTDQB2MNB2PWRUMT8eTos1VhSvc2gK7ATA669
43rNSSHQTCu16EudSGznzHF6LGD3lQslhfxity8ytrqbx3KfgVr0FvJ/t6agPaTg2YC7enWof4Lg
ZgEdZ7koGVGqTh/LT51YU96ny0zPUu0pGqYkmCVQSnztitlTOyTv1d+65MIwo4d9FrnlWqdKhSxP
dD3lzU+ApH9uhaeZB9GHGf27Yg9crw1TPyZ+D3yI+gh6yKDAHffb+t+mUB/BEIqV7Bsrxh7AR5j0
DyR+XL8hYBFZRZH3O8M4x5aWRg/p4jqo4WLP/a/mwApbyqlaCeaoRARkmBH0KWxSdIXBMfcS4OkU
yM3xbfwmMDzRpAvXgeSrbMFZR9bzFtE675YM1g6vWXjW09r1HjsTL4U8IS2hxqDNQuk6JqdZ4Q2i
3fg19OplK67sNqqqhl1A/ZmIHpuK2zTjCbka1sWJ6H5Cq237G6CYTKRhc7mGbjc6VhAmPASk8gjg
cET1T1dAVbVRHbmLdW40SXW8yArArX0nvORgsIkiSgZ6XN1T7JxrpzraWopSDRDXPZYxmwG/jLUt
FgRUdbW//m8VVBwQeVCg/sUM1o9z8CDbNREzFDrfq/RGC+kF60Rv5L2FTJrT0emSCQi9Du1CH+B3
R0X/Xu8wMNwpLDVtmg3vBtoJ7ekTcoFXWKYw2QIN5zoR0BKzYCqBqtjigMhZtxWXcB735v0HOgvD
il2CuY46xhCQGTaUMsY3J68ZxZ01P6x3/jY97E0H7pj70W9FHhGRcXKNEepBckr0pzyVBWvR1+Ut
4hfAUc0jbkJy1NSjbgt6XxvU3MvgqT3RrerrQ4tS+eKEiy79nlAvJZalwQAK/YBE2pwoPNpS2mtV
DxtCX/1g4SuecXEBupSNIunaG8KRtsQ6nQDQJfZ93jJyGMoRQ89v8KR+w+9Wty+9Ppf4RwHLXJPi
RICONIq+d1aqM/6T9sevXR/edO4q1VkIVW0ymZ2LkzB7rPL2G2TAwcaOq2m1tny0f3Vxy9gy7uqq
UaS6ypzL1RD6VuyVgjdccH8tbjlZr3x0E6RJjRN7Ui1CFUGe8Rt5iiXyEV8ya+RPzGD0unXSI20d
yXlCpLT+tyFPb026EET7ouwyMdR+SSWl1DFRao/EAF6mdbLDB8qrO4yLLqohJ+jMGFK8dmrXpR7R
vvOCXsS5qdmp9mnxJDthA7hfAjaEd2n/BiNlWLuTPlFkDqyohbEu57Y6R9j/t+UX7BoOnXfc4vaN
shulMAtVfFPV2oflSyHXbsP3PUEDStlzUEfI0X9ZPEUwx7hLuoZnFzaKDVp2DX2REznYg1LrlNW5
iltdKSHinYn21PRIlMusj2iy6WgqSA1EzQ60H0Fy+BP413P+9WvRYalBgCFEjlG8Ljf88Rxb/ByQ
YqvhYxU+rtldiG70DhrWTOPA38GJRzy9MqMSA+L32UAMjSt9ZA/5iXBszGIj/F30cOSaAgDNU8Le
S4LL9hoMjqdjA8oNP1bdBNQfIoOEfP4IOMufCwnAwyQ7z0ihAgaxPQs+IphXMPc0DgokUlLdvZ20
d51jkhzdF2TkGv6iYLILcM7OaO0AL10kfZh4vx00nAPabIeJ9uQWdWG/lL3Mf5O5RxuI3QQFRlf+
6F06xybSnPSVV6qXqMAdROYQLpgm6MFyX1sj5hHZyf8C29Wlx+RF+d/BK4Xa6W1RnihuL3s3B6uB
vS4NWq1RZ0LhnA1bzUUl8SCqKGVBJ9sXL3sLVSfvb50QvjI1RWIvpbibwaQNrhXLE1/tvGv/fynY
gWVtbdwRRGAQ9Z/+bawX0waqF6uhd9aXHfml5LRhchf4BWQua+DQVAP74z7ntmjBGp9YXcbf4ItE
UoE5gEirgWgvuJ3XJuCFL2NhmH/z3tcoWswTRxZsoe/y+P3NauR13SLKlgr6MAgparwpzxMGp0AL
NxAtyHx3hBkpcvZyFV87zTo6xgssmt9YiJn3r1iXoTch/1brKRYiZvveU8Tgk/iykZulSKJadShj
LcGtY+ej2vI90xbeRpVWahoMijAUyF5RYDVwKOV5+q6g0XO5nYQxK7m4++gUnHvK9QdO1Ic/Qx4s
ChvtBykPH1S/VQ23xBxH40KNIUOBv8/csJrcTDid1159DHMsjfrWazFOtpOEXxNy7DdZo+YvfHAA
YW9eBGfZ42N0FPp//wLWniV5Lc0yWmRE2WXLQn5sQZ0nd71T7xr8QLM83nmAGu9fWezjPL5nCSP0
QkiTMuxWzZ1Y2EurZbMUItvJ4q+AFPgzf7bapavhn0qq+cnfU96WlkX0vhSA2AGrntBRDsMnbVpf
B/S6bqjE9eoBsibeZFI1ZDlw0ry5U6ttYDMaBJ0FvT61wHgjJFKbCh+3koBD482qvDDfSIwy9Hj+
e5jFu+gPrAGFY1eTnq4/YqbuaLTl0M/mTM5lhU6EH5136IaqmjgHhVZ4iq/ZrCGcw2ufoqTM20Vk
3SdB4o9PRJT/Je3Tj+ODl2sKqp/sQots5gFZ/Naosm40SLtao0fBsxVDEAezf2JfMYsVXh8mdSt3
2qELMgx0EM0ZRj/cN9p0ab6Aoj4yKYnV2KtGXvF8MX43jxUEKOls96BfH/eWBj06vjQIRcSEhjX3
pc5mxVTJeCaNvyzpEpQMtRtyWdaSyWB7CeNVn/g95+/xUxqVdHHzBU+hRNPuYyLquWI/ocSqUBCV
kmcduP+vDXv/pz4pPGxxH2rNnq2dSkWyOdeR8MW5HyJzWGf1zK+CQLb89ORNXlaa2iHJ1Ju7C9Cn
nidmR5LPOpuXtUTff2nL7IikZhPKHvhKIIcKxJ6HUhDQmJxoT33O93I3GXUkonBzH1ZbmjpHtMvs
zTfnhikfSdh70xpc4Kf5tFkIcGGcydZOQ3MiEcQ0gy33oSP4djYSfH4LuW1HxZpn4aqNzTZpUYPK
rU1wHKBCD1y9DiehijP36acaUks//ZCLzL/erC/Bo2xo6c0aUmW1xZ2qaAtUIZK9y1t6TEfG8nN0
RI5Xxm18Y/UrYhKJ8m9Og7M9Y8Q22cwgs5mv0O0I0279PB3TGYOdcsF3E4LNFmzcsjkJRt77b5rG
C9zicUgKR8a5BxNE/XsMfXtbHpXplOGbPD8MyEgUhKOpDg743HUj3hfrtqPgN1/0ht0YDZhnV6Zs
kTCNwo364dO4smuerTVQL1xOlxRcAsBjpwMsOpXAPy3LktRM81foDsIR8E1m+ryiK9Kfo2MwdZr0
XwGzA4//N/2nwfEtTmqocl158rz4ntuAxKXSPNxwhmfvyh0umGyriOLVU2WDneBOrb1635YTnZ+l
jU/q4f7VgnHBEebFbitTgB7+22w6e/I1ZZq6imEIbOO1JoANVWlgRU4VCZiw+hcRBudc2ntkEcB3
7oke2OouEVJBwJJg5+ZtDvv3skG1nT6gm5XW0zR/0FR4AyURvkE5Y49KCzmRKflShgEk00jSZteh
IoKKjTSKFrpH1SSSM9ZL+IbZeb829b2T7yrXc2ZXlwGEcobN/XnKTD5JxfIAF/VZRFhPFUEvMV9J
Q91kcp5WPMnMzmBt2ZpIYNIhyhMQV20LTJ1uTti3diFzZ3WAdkT4ROSpvUSSeFQHnz2kU+WhtHsb
kc9ZxLyAldZmSkPpTCHXIq5hqV7PMbQrWONum6M8UX16Sczl8yhIAUnbXkGqsV+jzI4RrDHQkjSt
7oPDkLMFSovlxjlCFOQLxEPCClXY1Xkqe9mtMjkG2uwYfYoP4Y4KlGS75vQ3MEQ3W4avh3J1f5rG
22drC4/5mv+fAWOQTgpskHikDKwFISaJ+8HNA7hTzpt9hQv30K2nWglcpjBM8jU4p8NhOcTCMYq1
RhbHhXINiXD/Or27Cy8yBO6OkIkVJ1IijlErBwkaKO/yMTJDNU5JHUJTAKiApNARqWm+ZChjqU0J
OQqHZB6ALuC5Ol2mgKxnICemXfwmNR7g4crvhMcn6DWUMpvnygGm9RMglP6UuXVbtg3FUowCXXFO
VxDXbtqRLsvk2fchv7m+3O9AVDEwUq89Xu4ViF0I5OBbIvdjbMvBy7bqxHlIenmIi2WMZO1DFuzL
ZgT19ruEbFoZ8iTUFFCqzxOpUJ6VtvLD6929GP3YzsH/cxMXHWNcPpK9TB7DVY5Ieu6J9qCNCuB2
DmmcZlDkYOwupuFrkXMXiEAFosIog69dkBgdSHeGgJiJUWfN81aNHpFCLBolSz8r7LzZDAPnUaUo
wRjR3YxkHWFho9RVV4Z2fYH6kNiLtzCFAbMhYpl0UecnwaM2EBu7SgrSmWRrtQt92Gn4JU9qsHL5
u0/Z0D1cAUce9BL/Bo7RMKFPXlBG2So77hZEF/E785TSirHY9cFS4btXcDbv4nkwqzhRahaj61CP
fEYA+Yhn9tU/RP0oMcWnDtvpJ1FRmLV5qAyFhW+CTh/wjZKewWrh0H5Z9Y0lpzVrc/W05FKfyqX5
0kfPyXlm6NxVTe89OgqdBe6IjlygCT3rbncT/X8HkLLroufeQOJjgpuVL3yQzzr3rY2lxoxOm97C
Z2swzsuXDBJ02u+gsGdsawePflqZtwSnMKdJCBmFCmaYOFuqYtwYEXGNt2/kpiKdSKWeNJ/7mnwo
jeoZHaWJMBQT+x2ANW+Tgh1vA5r861RHXyU5cPJZJIh9ftP5gnlFN8MBM7MRBlPBBKGdYGipRpdo
qTLTQJ9ykq/C8C03dhwhluDVumuWyV6cv6uvhqDo12v/AHDDj6+lggiwU++hlqfta0tw1b2nGGlr
dI9QUNgvK34+16AfSQmKK+f6e1aS7fvM2SA/W6GtLpO+Uw28MRWzA2P1hlBPKvsF4bClo1CCP0TT
Ods8fZA/JHBkvBZckSDcwsoJWqkqqbrpvBNN3tT1KYoYA63tSDMEyZVjNAYDHJKo8JZoMWfLPp9v
YFBol6DVL6vJ7RJcMbfHCvUdnz+ThEZf87Z3GHwHd9MJz6AYM0LTbByCFK71wnazkXcG4+SiOZKC
ZFkicmd10hEbB9JDWD8Kij3PVXxRiZ/0cHg5wmxx7YU4BdrZwKEZsP//JBkx0gSzh3yYXlCk3ROQ
Fi5pTYRGUiJNkRmaTjkSjMLUpCglEFFKBWGO+jZwVhdxToW+INfUcMZzEKDN1qt0YYHd4hE0q7X9
RzXm4wD4wvqXmVtpuY6fds/QnmrYZntOyo3cbrVY/7YeEvhES6foIfUW2e7D8/VOAt//noFbZH7y
JJXutVAHr4XM2r6gO6MJgWpOQkG1M0OINaH3VKSQurCqCyLDfZF2Wk5mP/vPlZTy3rlu8X0NtGl7
tfv6GO/Rd0vf+/7dzER1Nlfic9RNtYFRCUuNCJcHxHefTTR0sJ5jhdZWog9ZUw0gRAWM/7Q9cNPW
HPLoWOaUl4jR9LLrAOxQoBd6204jW28yaEF2DZB5XHyU/xpQ5LXJuB07SXNlshMnrBojFNb4wgY0
eZeaAnT0n12hL//I49jRwXuEREDLEY4nnPX/Bn09Q2A6w7cu5KWWpz7jwWi8tyyDefH7Eg6mWgF6
JnsIv2RAlShs1lg3Rb5s2/02HZvlsmvuyWtNvvBO9r/cR/FOp/lELZ2z4bOhk0ZqZKRw5VPeq90P
o+02pPKIY8DwbPBpbbGnlTVOW1R+/E08qsVOBdp1yjq5cXj3WIalWV2H+6k41yJrPUQ7I8GxkBwm
G1G4ZF6DKunyM2sCr/XtKDf3HUddCMtgIPOyJNGyFGzXRKy60/hF8mukKr8TKMm/VR64iONqFtEb
lbkQPI9flsUH96P3t7bJWaCu3YHfu8bhrz91RxUewzAXS15oaQfVSmM04YZ7D3JpP6SZJEsppaZM
UKBn2AVwD8W356nYxhZnGuFdbNds/jeOxYPTrAfEck8RYCIFtox0Z783Hg9YRNy5FEZxuiPspR6Z
i8SONR7pjU6VN+VCd4IYt2ll+0HDvMJM6l9iS0atLflpdkrkbJQZe2pMrrF252zbaB53Pnnsw0If
Kq7Hrw97TlrAmAu+wxf5jnsip57AyNZBVtlE7ZYzA6XfILLm/qU/eR5QFFbLwwPeTnM8eHt9Djxm
ESQHxwQBNnwrUY9pRXdKZ91FxNKf+Y1xOLt86J5vzp0USGwALUdZ1flE3lvl/ALmyv6ZIR7wK/Gm
XigFjgfcxCSQKdW7PQD1+hErpnDRn2JicyTI0w3UeqRBX0467Fj06GVplTrc2rHZVXZebtgsbQyz
kiqgQzIojrHezwQlETHsC1TQeoNtjQftCmDln6FRvGRvlw6KM0h4wlM/HH9z5PK7AtWOb+oboDSQ
u9c81OZiKSx7NHjyJpTFr+/IrDi14/P1CnNcZab66cDR4ciy8lnAchYMe5LOguUGsMpZ5MiFuKjc
HpIAXFKla4CWm0k82QZqv+G+OJ5S1t9OM5i0/0DR6tcoxVSrdfb7dPXlFpjn1UD5qYXBYXtTAmr/
p3YUlyejv1qlfnz0n2oAb7rWa2FyjHMtmt82+WfRwZs8hLbv88L19HIdrcGL35CQpMonlaB/3HVA
kqdr5TJZop/WNpMQevFokBp1/qMfixW7I3U4Adc+2i5tKMb5Y6nlqMlRwMWwZhIqQi34JT9kx4cY
IRmCN5iYnt09l+nMhrC+ol8I4QV6pVkmCoPfaaaAN2W/2iC9/UgcSVzEQddbCIYb3c1ppvCZVvaR
6zpwtfzkHTHuVYwWyoWvb+t4YVEJ2qcY4Q+CqXb7fM/lbTb1SiDaKbIENWTsLUQZ94tI/NvDqp4f
2jjcG7hmXtJanqUD3SjOz8zCRhcSTo5N0AzJub1Hj6kLw1+o7H3KNEZxkBlrFIhh4H4SAbjf3iNB
ROFdznH8ktyZhv+L7wJ+bHvAYgX4lGvYdyAhY+XBWcp3Epz6Lmb4eHBosccrviynqKjA5B7UHEng
W4Y+F40sow5X6XT5oBvnezTzejJqmF3XueKONHEfaJmiD1YzkjfZVvavoyXNKcPvKEj4WFJXQZ9w
Z04kjgAkdRSK3knDJmE4n5QZYkMZmb9Kqcf+Q5Y2PqDjkl36S4QRcYEv0nu1cLafTOxsxpQ2fHnj
7f2q//EKjJY5uSrj4MYqbf8q0dGLwv4OpNYq35oE5u/Vq33aoBS5qQ/RMXZ9TpQ29xwthiRTxgrU
CV2K8E9u7WPT6pgIX6w2zfj/ks02jthnWp1p0zBav8j2vBV6CIRgdJKpag6aSsbi/y5mF401+PDi
YiU5fN7Hv6mi0+lgsQBFtUmP2uCLyKNChkKNr64ER5t7Bje3O2vl3em2YneGEo6iTZqAARGnxYGu
DMY2TqnCMfh4pM38rvgqLiZ/qCYzi4Uc7TMn1NYZj9XIexPOMVW6idLTJpSfD6C23xPDVRLsK3sI
3OV6dzzuiZ7KZjpjVZNsx45frBdKw1OAacC6JxWzz3+JqPDicDCpeBfZwsyGsPTCkj+pElCs/8Xu
fLNav46yxEY2hCQhOEEfpShEVB/3doNTBzAA0rqEoxbpbIvwUQMLbFwiyDXL8UUdomGzzdnTri7w
PS/xaJt8rd9wrSwQynk55WIKezYQ7nnpv8ALkw76dP4HJ28zKqlTm12tP7F8ESvmSBRDmzbnCxEO
lRfS6lFnE/RFtBl95bWVKR0NabHn64nK8dCjhEDkHSu/gz+DVnpIZGNIyjISP8mc1+INH6nFhn1J
yoGgqbZUWSPi+cysWRZ1YdrjFP3F1CMIjUeDEuIHBw2UZ/ySP6ZrSN6TOLIfT3DpXwsde74LlhxB
o+cNgoorDFxyb3qLxlNpsyt+ndGH6erEhVofiPQr8KJa07ydnZqgQmFu/vTFCh3ljLmk5MxgeDy4
mbUXOayIPThUuZdW3wU7yDboJ6wp91RynlQiK7uzn/B2NWlF7Wr6T4yVL3QFn3P1StLTBOiXWysq
C2CgER3rdIRy2m15baCnHGJIAnsZC6/+ROb7nDqU6WbDaCGbaI+Yl0qORcVmQ+qA5Hr9gfT3Rdlc
8iTWZZCScU5/wE7U79brUtSRruBlEQxSNVIbQbajAPwMHX3A+RxLLB+HgCAi9QVmBOy7w03pIFLS
67bz1acHahsWKJFlaJ2K0e1fAV6EMi/HM3xgToBDTUh4WtuLMCfM+Ui3lZtMpO+U6tqdjqiG/2Tp
WwXF+uc7rE/ZsMop7Hb+aqHHaakV//XL/CJhMQRlCWvYd3Uh1FAgexn6uWv/QysduBiv0Y+dXvXj
WANARLPiKVA98bGHMDdKILHilgqEdl3pQ4Ry0B1ccMKZoKHZjgWAtz/D+mobDFDzbkFGnyC+Rp5n
6OAnJwCmpw5gMQ+XxJTS2wSmqEybG1Kjv0XQqE8QRllTC3gjGLywVoza/dS29LI4rnYM462Dnlfy
M1/Tc6qzxYFDeJjYpYxbGZUQ2M+hDQd2AIm21DX0CEL8SDO3jNEpzciIWsYyzydJ1LQ+0Lg0Ac4e
hucXjnQTUvV5oovMRK/aMwi+eN1Vcyjq68enfgveloBuhLnE5aslf4TcpHcGHXaNfxl7+UI5+Dn7
l0KBTZ+tERzPyvwXHl1MOvYkRgqazdqbxpZoj2qRU3j6kBBUetDkf7B105DSrDJ9AsO/PMNxzGtq
53nyTSPD8SdQ2JsYdkJIA6pGbAo2S4C32kdoFvSW9BZ79BS5OVDnGMd+MFwOi5+S33WGWyacNwIQ
rGQOpPC39hkPJ3zIUgomWHSsy249ypeG2na3d8MOUzEpHKQ9qEvdt1MRImWLQdsULqWQBYPGU/NS
XC1vJUJ8RQ/3yP5lNNZNGqzIPl0kNOzkBOHZ8PktUWdmN/GKtZLPbTxRk6oXD9++cAgRlJGs5uYw
2JRqK2FjOMgTZPIovNAJ3mlgveD/d5i4Fbut6kuZyUlDuAJAWwJ1yNShej14WE9WR9BLKDU+4PcI
YBOv+1tSGD1PG8LwWic7DEP8jMPfq8YiUOXViaJjpRFKUYm9dAZSHaFw8wuFqQh3vBf3hjPU3tHB
XtW02qRLE7uOIARY67rdjCprX8oueev82urqTPUmVHJ2vRjkbZTqYZZFQOeoxvXR98ccTr4yUA9u
JavSt77J7OjoizpWOnk6Ve+zpufTwMNGbAfI7YDOo66oDcsvWkVdQ2zpLgqJN5SS2eKVsq180jba
7G2FqzZ5pCvtl/408cVPuXUPdCSNBFtWZ98PfHVQwjacIQibt+Nq56SEVWmv7cP9YZwNah8liFHT
TWGQDxeo/XGYGlb7bWQdYwhetprhQy1jRN1EtCpAds0bIjx78d6Ir4XuOFGGnjZmgAgPX3qLFydZ
P9j1x9xIZVbERCiddz6OrGqsQYRxdH0zj/VUxyDXQMvjRT2sxiDcgiV5iyIwxTeJ74j/6MreE7NI
UztSwLlUQwPYwdPb6Lh0C3QYvHQecNe7VGdZ3m7aQQfe9u9njzlMaVviND+F9OKDFW+XVUdCl6T+
m0eNvknvL3towDDykgdEyIWbAHbcf6q0NW/hHt5PsIZxIrNUR00TcavdYKzkg0Og88acjqDlzHsA
CrYrqb6fp4Y8ceBuHq6Aqr1tvvWOuh3CV/uKs0b9kdwJqCiZqgZwfVLeA1VnDv1AL84nCjG95OD3
ikSyPXithg34MGHgGclPn4gemLZIwnOgftuJ/cgo4mfvzWUbxt+7+8GjmM+ppkcEcw87Gp43gKQw
wLyW/i6vq2Koxwyk+CBofFsY7J3abocZNzqY2j93EZdz00tM6RYFE8VyAGlFfnQBYmKV4NrCP/9G
I3enGKVPX8xZza0fHMIaEe2uY0PzAyTn7lbaN6EVMrxVw9mvV9NFn1v9h0nCqtSpZ/CunF42hy6N
47eUMvIc07ccbp7OZMCgG7wtiJP4kfj45qIU5m1KdsOpbBeMs+sWEuETeHqIDIoJuew4SzLGnDXK
7AtCWJf3NdJ91n4idG8TcjU4iLxgLVbPMrn9eFy1rVc6qRhq5xRG5wG7kUmNBou/xhzrHaKOXEjG
uHEKwy0On0kX1rDwNpLlI5Z7NaJNbbQ2w/4tRPBHQsqlOSPlEOpA3LBVLu/z9t23yLdPUEtxj34s
OiIePXCxz9Qh7T+ABso4zQ9fW8+vakZi2aAEpMsqdxLtTMXJRx8P3rClMXg2MvyZCfueUsLOLuPR
SjROMX5zTk34n7KUKQDrnoMPg378Y1A13k1FtQmmNNn9jUgQhOvxvV86AjfGz4ndVLmzxMm31Dzb
ylZCtAtBTCDm/r1zGvuJy9aS0Qne2D4Hm6kHmwp4hgjWU9KVG80wg6tb1NwEwUKZDP8ji2klwBGA
tDUtYKoTpptzwpkyz2FP2AzKN+HMzNTKbwoJXvT78a4QQhb8828g3Xas3huF6oeMPQMXVeS5v7T5
mEJuDhG2/MprTaW+N7Of28NIyyASkr+54lY6TUeo4SY0apGe54+4G8wxMaiC7mVNElDMZvFixECZ
dJsT5jCwZMFHOQYOQ4u84cW31vDOP4gZa6xVxi+Vs75h0Hyxhs16BuGnCsIkcZaIOAW/ALZrIIna
JgUEdhDqXQrI2ksmrftLdQqKvlwQpykg35nfjy9+tHbWWIIopzlGOH90vqNKK6MZ6ehsWXIn76NO
gGEOvh7KWsLj6Ws5n53v3lMlyXYMnRgd4JXwyNhBmUM16rkqws0a9zIpOjBZqAjNoYZl15gy0cIm
+NUaRaN+R6VhIF0WtArsAv35TG4z49GiY10yANYOAcMIfx7dljLSvXyFnmd1zI5rcYh+aXQ2B+vF
ESsKgbZtuM0F3RbrdCFl6LmszApDsVpJq0lhuLfpSBSSjH4K7QpGc97VXFPduBlRE/TIl/SjQIqq
1oKzaClFSGn1fWL7q7aGHg+LZp6XUANDJ+w+rEZqs8mBjLCAEIBSToSg8f1ncfWM11SAhjxo6q+A
ZTGdUZI6Z7Dor6Gw7I17cxkdx8gkI0I2ZijMd8i4njUhng0jhRcvn04PxvzxX7Eh/RsV9zIHDSfS
R/PAuDu9lVR23S7vfsmqNO+J1egb/QePqhgpj88WVDS5qnIoyXpQjKYo74pWlpmm/L6sJAsWXFUA
U3JsfnvWNsPm+UK/gc8d3skEPcLlqTVfv360ONg65kcQRhii6cjzGv7n/LtOSkwJNQLVXJnP0QAr
vNmaOYG6jK5uaA0PyPt+3R28rXxQtVRiLNRSbQy0P+NzY7V8HKFLRhmV+8cdFgxRJz56SHlUY9y3
3+f3brKkjp2IBeCbKx5EG3LBfi0QocK83QCuku28nDIZvco4V7o+WrCLBBqOiNwy/b4Yl9kGZTl/
j+UXuanAMEqMIWKv65bExMtYG5u+AzP10DnZIzNIUeJi2DdWL1UM4lU2Lqr/tMwLAW4scKpopbLc
BQGsCrK50+I0bAxdyjdR/YB1DZdemJWzP8ROTrM0T85SlCoyct9eqYUTbezkevnvXHARKoe7VQRa
wnSTHtkQ3RnJVOqZWeVuMBoQODZXwaFAHzlNxjZalILor/PBeP2jZljti05LHfDsn5wHjtMOcXef
k3rw9KWoQo4dx9T7kne96CYUBBlVqj75+cUJCM6P3ukc4YXJL3/SKS7DHY2kN3kFrAbSUqs1ANqN
9DE1oaIBPoHRZMAyG/eEfYAGZEjbiVXCG/BuGl21uGJT3IkusKBoGEhsanN+ETF5JHd7X4+wQS7E
EfeXh9KwZEUolet77ExOiL+CUcdVHXgyuB1UtdlNOtQndBp4suzgoPn/bXpHZ3X4hGT54hTcDjyx
oJFj4hjKSTxKzhoR3aFIerOQgVawSldLMl2HTh8+7t6l88Yb62n9du1WxlQo9b06MPf3bCnX5Q/c
OJeqIbRG0slpNXtNsPt74AwycmNko/mruIGXs5b2YVl7QsGbohElXrbxOUtYQ420OwlJ+1585/2S
PBzqUsDUrSV1H/XfRaTWw8snUcV4xoIyHFBxKspWJ0tknlM9ge5K7ORnCS0LcyRctvhyp2N5oNjQ
nRGjaAfxdln0l9/HJvI+KazTez8NubWbluaLl4YuOqKDPyjWIrpwwzJ9wGXFtBFEl2XZ/5UL0/iX
qf3jmMG4u2/ydByiRZO4j8DMWVFNGw05gth5k1XDJ9oH0Dtp7nk32rTloZn4M0msYIeQxy+WvFyS
y8ZaGrhlw5hqxz2/LUG/lL4W8XLOnRsh+k1M12l8boWfg+QwUqp6Wxi+bzXBpOtfqYICE8WLmZjg
yTYxac5EJ/qlQe6SS9+OPbVoPYPvcfA9ieA9tKbCzaXOAcO7AHKhqXXZAZay4rFZuZRT5zpcslCM
C/SeCgiLNOkIxPMuTnCT73CzxHHiUo/AH8a9NC1/tTdBuBJItopXQovTdXZLTeSB6QN1uJ4O38cG
Nc0DPAEPBlQGVov342T86RgymxHSb+GOpjZEkSfROWZZaDqAnAWuWhgDg70n73sVcUfWcdHhMBaW
FVM9b+W98vlBgetIcjq2U/NUYmhpzK3Gt8DIAeUmPafCXns9096sc6iGUEz/5vQwjMfUANV86qVB
HQVXhueHDgHM3XGoWM9ib/xi9/AjJWE9q57panJt1J0bEnlHC6lbj7cjoL1jmlwzwqKVfI2iB1kF
NLoQng/jCrKTAbL9tiYfOo0UFwdOZwHs+AnZuuXP6ldPVH4Uo4phNtb8vCTsDccdNRWy01iaNBIb
xIV2/U1GWrBKO5CfaqkqDgVnNx8FX4pISx80QwNXSBBQFmqA5jLUu5xLSmreZtdAR3x4rP9WPMDp
eCP2AuPiPG+pWWnWXEyQXsgtHV9sj+9GrpfGtrWyzIwwhSx0igKc/x9jN7rrfesZ4jIZ0vpz88xB
iPK//TLOzAuSZVeM5Ax5JUJxs/sfAWjUoXPFcCTZgbSUpwl4HDdp2gLeRhKg7eJmaXLsXbWes7f9
EblzykUakooSJH4+IWOmj73PvKRAK5Z/O9KJ6ca/zBZbjdgQG3yu4QlkVd9t8hBOrK2/5kXt0T2o
aaOEIvIpj5rKFdncN3OAWC8iUMNRAf+7/gOu/OzQVEMWqF17H7IvArJR74l83oFhh1+ZRAT5QEoZ
xELsAQyb89RqUIhQOqMuBHlc8D4UX2CheABftQGlocMaU8Fwjn9kuxqHBepfN2m3iQ9hcstGrndj
LFybiUhaRtjBd+u4HT/Pk825zegQ2175JqhAVSuS6Uk7v3WulmHsMmg9n8OovFd5s0nNG8+yhPZE
zSkVB/HkuE2fMuLwyeH18IoHUayz709oJDgFkpTmqv/NO3h6ao2KGyVm2rgKbIzCkl3YOXV1mFlc
fMCJkn1G58mdULI7TNTKTgkBSRiE+8l2t/8uyrkyfHnJIzeI8a0zOGMSXIzuXbMJZz+O9zafwd66
lMWVKec+SVVbH5o9onXBpsNGnp4AT4iiFKKnuozcoTfXzFIjaFYP1K6T954spJLOtYRP/Yp1iJS+
brjpbbYasN6VY57UQsSwZ4T10ZfOTKX8YJg/EyE+z3RvFrmpjjawH24ru9FW7qZS/xqpvvCcx7ET
v4Xe8PA4B25/KUvsqPQDz+zX6B5Cesgu24Ee9rlUjLZyqEfGy8bRITR4rbjPK2Ndg5o7mlSoE5iO
fx+VwZmDEKDfVKvKCEoxxde9MZW/V27KxSQxgdcO+JjxPoxKe4KiSZ5ja912Ul5xnh8PubOJpR6s
6haZ+iii3jrzVGVnkUms6G6q9lg8O6Z2rWiZErWW9RywstDxTDZiM7jHSkrKzLBhp/yl99QmENbH
4hqKiXlchFEWyepQaIM5+VNFrYUQzA/5TngUDprEZfr1U+1fhiNwFVjVMl+jQnQ1+jJ/FYCdWjxI
ApIlJsJ1SsUqoHlNQ9vO3W0HkV335dJ/UPdsf8Co2UVZDYCZNQREjq8P2xo+aX6PAlOVhwwDwbbP
XSxllRmHfUErPv+5ZGtf1xgNRgklYimPzF58ok19/cxrk7f32j3Y66vzBeyMGovyHGmKwyr4ngiw
A+4K0kG97BFy7aaiV+A/j1guTnQpzxrsagpd8SXavsFN1NTj0Z9ElH4GTuD/Q3ydhb/mlfZd0G1O
+K/9nCYyMakqfLYgWI9g3DOW4fYrVQLFBhKEvDe175Vv4uPhBwL31JrOuCpfAc/OQk3MjZth6iAO
PSJ/I56tl9noOkkZbNdG6SB7Y2kkjqjxTCJRCctqiPLxQB3ixtSmSL74cvVxa9UQbVsXoVyJCd9T
nf49CSdMifNqCe+Iln008/u3aWi07rEckKL1fmMfRzXrwX6Cp6Rd6gWu5ZtQvxICNk75sqMOW3lP
S+icKh+Or6MDdknhvnQgfy77Ca+5EcSAlB3rZxHXknpRjg3NvoK4EbE0HDgiaqJza4IJvHziBbvH
V3epJAETW48c0aB9bpbO52Be1aV3x6B/deg8ZOaPaZ6hAcsYeHJwd1B0KReNg7ptpjXeKlZs7IWA
jk3S01mSjAhNL8HldMs44gba2wl4OkgE5HykiDhJlKztkMxymhDxfWzcZBcthRl4b+ANbZ93QCpl
En5tyQhclH4NBQ9biWWmIVJEPxTQN8HirJ27uaj5XoSNKwxwkmh65t821X6wR3T+H0aRwrBcAVEL
iG2VF5xogqc9GWNrvlT7U79S3zUKYwIMe2ikn0K7arMU83PE+w9JoTObjXYN/hb1a77m1+i6KFWw
wMcWI0u8HmOmlQlHkQbY/ZpTFRuYFMEGFgt6Q7TDXBD166fpJYi6uhUDWCrfTBJIlYQgERcPSPQ4
b3X1Rz8j6JtL3JM8ZUlJw0wjlKapUOc39cevy9S3/1UrKCDTeyXapxQTA5lhmZnq8jUEXJ0a19mF
FYFdNFZG0+WMi/hB7bXZL0wZVpBoew6xbPQjjrWk0qrshVE59RXSvSUYR96aCOpOJ99Rbg0fgZdQ
petJsjrarsNlGF/e4c7+oxxWysQeDkbahfrEeEFU00TnmZO1TGmhUnaammvEUR5SRp/vJ5Kh2ng0
ViHvlyAYd3sTiZn7XljTCSTM7CaMQRNrwo4VUkii84u22my+Vs7pyNvCmdF+Mor7iTEhVlEuo4n7
GSfcgeGBi1QWsYRmcHaJ23lhjRxr4/2oC+qishUABZDWv2wn0IretI0VJr6/NCHHmSh4YQXvopfh
wEV6U3w0fKfSzgN6noyxe5LM/zjQKI5ViY3+q7Sg8HxlRtvbzvrhnCPyVVK6sgMa7Dzf75dcMBU9
M0swgxb+w0N9yoTEMzPRxio+FjBAozutiBPGGgbkBkXRAwnfKZBbvnDOX3InWG9a/dAKFWHCHexC
37kzXJ3NIpfNF0yhZxHbXcBjHsZg6AnZxLgx5moe7Stj+QFNp34Kr6IRS6IbQge0pqFeTQ/Xck6b
r/XGcPAQAffcdHF32mQTRKUs7DYJiI1JenBDXaa2/ycr+hBT2NTdX0HK3FA2GIaBySSZ7Wc4Ns48
7vAFkiHa+e8NUg++muQrFeDvd3Kar0Pybwpwaa7rx9+o4rX2VFtV6wn7ZKHYcFO2nEl9xbj1WYQI
4xalvBeluKkYZVrUnL1YUJZTAtMk054WBxYG4e104OJK3yKQQ9srhSA+wzrDHm0pE+S50nEisH0Y
FKIQRN8yMWg9gsKhf6RQ+0Yken+DIbMG6smSxVHZFXe+uFZDujBfxXQdNWMTXfM2WN3mMjOhtR6J
pIJbRI2KZL5wsA2i057JMPPoFcfCp0SZrJ7aaltQcg2jvi3ZUOxP45VFdjXJClXRCBkJRdAjRVby
GKiyr0UxNO01Z7AtZZu81AXuBaPChHCGDA29YmaWfKOQMH+nsXrAr87Iye490W9LbLkEoRW8sBV+
h3K6Qh0Azil3vF6y3tX5vFJdJBYC1ZWBAjV02AAJFhGLluuFCeEXjqBWlx8AVT95GzIs7XsCu2QC
OloSmUs/DduTHSjHn5VilamsG2P4hnjyk0vEwxqpEeEhnYyo4Yra4QP/CJaEsY3HSSl4EZednFi/
gSPTvscap7IlrOCdwjeMH6LH1pDb57f7wgZlALdec3fyl17YwHXKKQCnhtR+WGKmp5u0eeeBJeyw
GcD19qIuGk4dWgw1viLJnLuk7u3y3wOmg7WHcX9bqGqohXiSvKhNpZtv86VNgSgwm1sJOP1INOxS
ldAOkVRSTWz7QMuudjLrp6XmbTa+/5dqlCKrrDVjq5+9kK5ZF9vVG0yB5z5aJZY310gOk0gx2Uyz
p5OUgzU5fyTcCN60ejvHQ0rkIfHKXx/W609mBAbjJ4We6VVPDdYtRFP5nVJPmfyuuTml2F52sVY/
lVgdsPX9UiKjSbVnzDYZzyG+iJFEOVaD8FiPuPXhjYClgI6OpBI2WczGI7MT/pr6AgoqPt/Gm+CT
itlGjM2azvViaWN6ER+xMBFIzK6RXJ1ji5V7kCo/wiOthLBKhjE7RZPMXXWYccUKZQ4gPg9K4+O8
E9qCtUkBWseslkF3+KzMjHZGI2O/2+8jyY3npwUZSqlyaJGTh9ET7IbGcqbuHGKrlesuFnNPtjhS
C8poz18IkRd/679Flb5CaTbvl5irVHNodHznwhDrdG/HVkZwQfdJkUIIz99TPvj0fmw33nH5uTAy
6vM7l4435rlKL+dP/45IGxS7uOXP0C4PZqgKtd8055/KIaZQyYW+xdig3F1y4urwlzQJgeXUZ5xI
36YK2Co4M8p2ZgRonXG10j7PF52bkYYXz4VdY6jflfcUqlzGS3QMEnCYtNN0ApGO5er9nuShD/10
ZnsPV4b7GZvZeXNSTv7xNe3ZhZhxFo5JnQD/wBR9Ds0al86HTE6TWs/FMLGormIN9NZtmc7xhtP+
zM6Pgf7fj3k/6WrSdU1jGjSzPGGiHcFPTaysmUGSlkK4+JlNSrvOBhYFCyyPnvxpJzWEAna3Y7j/
ReAZggM5CQnnkChFcxeLT3R5lK4Jq6kMTgFrChTtRbcEgwWIxhcUkOzhrF5DtZjwcpqcxz2m/B9U
7gvS0TnARL7SR/5E/aLw3zl+oEGY+TgjRjLaYPigXebzqJdI9O8ulSx/U7in55aMozH1iv7jzQd8
AORSovmIry/aZloaIX4JUuPQAo5C0SQwG7tmBk/R9+NWkHVAdFPv7Y/uboBclERFuQJ8Y1SQ0EMO
D7jevxZPaY3Fzf3Q5VbQh1ao3DEjcO+rP6VO7Gp9tiuZ90txbHTzGB+HTGv7oq5Cz4I+NeW0i8rl
RpStDR/EkIJhUOa9AtRx0ZP5H671UoWqIiT6erR5xtqpLYHuqr8HbnGuJjzItfQw51d8yKS0PRs1
aAryQw6sJVMOKSDvgX5ZYUSZmnpFuNEWE8kV1UmAN+IL9AgQ/HlH2M1SGv9alb567CwYquvBzKZ6
DkWOGMFIU/aEuw+ceKrhZfnOG0C0QB9dOoHiOvcPtbZ8QZa49kjUR920pYMyYRL+FOuToeq52wag
ToZ0EKVeqLHgvQlfoG/IBagi5V3lQj9dQV0LVIxGStR3qP8vqeuRA0E/PdkRcy8CAWqPP6uGw6AT
EQw26celRvh10tgnbv3ULe1E07pBLK2XUPUlto6tKxJJaPjeGzNeKTrochISs97tMDFEFPw8E0Ri
zugQy/dfun4EF7EtnrNPI/5n3lx2gcEsTUWw3sxQ4xWcA6BqgalGNtmABa8P0PoQcqKKglblzPiD
rrdIjyqUZDbo7mKWEi5YohNurlH6z9VXPse7BOdkpNwHcp8Owkbhq8lJeVYGi+lhbGeiUKwUpiov
ni9eGkXoQFny7XOwKLY6pjckd49mNvC1H5NYJpJq8q5bvSWNbkzKQdXAhSggG/NL5V820lT9xdb1
PKbVzmgUcYoxDDr+vAN1Zk1YiRHRmCyFLJN5sNqsN0rMzka1siB/aR0DWPuXx6D0ErV13RBs+jH3
YHPXBxsD++192+GtT6bHoepj7sHPfflD1qf3DUUuLPVUnoYjYg2ydimaRvmBtSoQGlQ51YjgKDMy
dveFXMaksy2Zom5Fh1fiVqfR1Mwm4C03rC4IDpvHoW6Xgknon3p+z2e74ryZ3iYGHbioEBzpOnjD
fbZut7ANM4PgXkV8iTp4aQJS+LqwqJ0dQnmat/DMOlDNrMS7QtBxI3394yGX3vRWq2qL0//3CVwv
xoxN6OeIcJPn4w4Fqf0MtLo8zVDM7jHnIValT1Gn4/YKKTm6ZLO/Yf9kOtRIPYmhdc5OeJUDcG/v
Hj1eWBerIV2q5S4RnqWTXT/rpvmr1mHcWaGM1TaL2aCvtwYYMuuKo01ISGHj4V18na1df17H3hSF
RNOkp7aRKDh1WdXjZX+f22IGhIpBnulRc6rALbePkefVBEQIJJwm3u6nVolBV/yAJ/2SzGm0x7vv
6cb/dh4lEO69DeS5b2yn+HXpzJqz8Yja2MJnmn8P4exNo5SSZhjgMEMhncP1kzMD+PkR8EJqiFXA
k6RlvIWt5WxkQ0LLaj8GtePOHO5qjnPnQv23qjAAVlBWYzh7PPD/NzZq+CGnZPMVKPLcLn23+abH
tuXg5kbVQbRta64VqHpXeqpSOwXoTD8bP9ejLwVJ3fFYIAmfyA+xAezCjeGkra64DTU/7oRZQ85v
P0iH/Jn1X+35Yw1MhNNsfwiG+OWrGVbIC6ga9sWTQd1OirxpTyCRfNmIsNvY/JLJFmywrOsxgA8B
+OHc4cJsF3rEV4Srty+dT00dj7f+DDyJhVMHcqW+EPQim13vrRmBoie0n5LaTZi6jO6NSGYfDqM0
Te6pKZRCwM4va7MhK8QPLyqdyo3XBcIToIeE9of/ZgROoCK+DGT6RQDj9ymbbpDrUfh7Tg6zUDlt
2S80GIjX1k2rEdarnCSUm0VccuMsGD9XcKi9Y6lQDDc2SMF+DRDh1r++1itxKgXO8c3Dzkw/mTlp
lDx1bQGQEQD0zqRNuRXfCBrYvY3j7Pqz1h+83nxWKMVHQOyaPikeJtoX3x+pAKM7cWj/48WiC/ck
FvWo/TGDpp6voP00dgId3jutpUl6BDtqIXyMTKl2Ks9CJ48wvcrMOeVhNfBgrvzVb3y3J+VuKZvs
KUsN7KgCdkgzc7U9s281EBiE8Kv+rEM3GvQgCinhpQmzSth0Chi8tLjocP2YCPWH9IVfspmYzwmD
gY1mQGJLFgxy9nBVLr1NOsjqZtYagqkuzI2Vswn7s1+FfbwdctJCqYn4gVqqK8gZLrMV9LzvO1OL
O4J9Y1l95zRgWyD1KyoimAjpxw52wRTeWwk+Ka0ouTixBE/DBLIhiOKQf0oXFPqUgc/omQcWg2e4
B3ZE3SZ5tNnj2sfjtBiwZr1tCls4MU65tf3wrpWm/jU4MA5YXovs3/t1T1EC4d8kwOfEEbyawv5v
KLStrBkYYnGFS2zukJoePyh5THKzHilWGZshek0Mluaz5zpUaqOFS+4F4H8E5inrnsbNUjlZSSWC
iudX8PBJvHBxVXEVb30SSNuTAoa7JkWdc5Iry48WSx5FW4QJLfROb/cj4D2N4ycqLfkT6PFJJf8h
zKjS7i8Il8f5FDz+ZL84O+UoAf6huKYq4sg02vOWYKjTzr00Gx8SXOq5LxaCf0qR2D0hNzs2ewox
OkCrywZtIYbsRFleJdeq9IFNMBAJMm5diECP17bypoV/Azhm0YtTJr/BqmBTmRSXbiIlhTgZOh6L
PjEknORL4ATrQUMKXUhZPLmxi+hpVozfDjgwtZ3e2uk5Ce0LrQQbVhDUVyB0pmqBaLsKU4tyxVvT
Hy+Ub/w5vnAgTfiVs3HYnhNE8mCl+iirHHkB7BT3VoW0cXrisEf9227IFTqsJn+rWVnd7jkSc2CI
vO+xqEN5iyA6g9LmnWa5biSQlNYSmrJ2AW2nzLyKjpee3Ssr//HwzCShY8j1EYhKOhVEVWDe2xJG
U5fiwr/NtfKewrNRgWKRRW1l5JwHraK2DICR0+a/+vIlRIiSnz7ObL5F9THvhnwnG0DggmScgwMO
y+2g9V9Djm9n81ucS19SEQ7x4h3oQqVm7VPW3T2sy7v38Bz98PqqLwSEetJJwlqKsGsye2EpuL0B
l5qGfnVvmMzDjF4AoJKbznzcIizLY+kM8lchAuiWpL1VGDOW8z2wasTZciRb9zBe5+mr+QeLtqHQ
OWhUsP0Juz1/Wmmp4CakIQafhY0Wb1SEC46KCCQlZ0oeXWYLVrNyNrxQR73h/HYySKJOQgBjlvTp
E8/SvuVA7mv6BuDOC0HGlK1RfAU4sp2PL547fnup4SH8tl1zY6qQB81AT5SfSeOiqt8TSUWArcx4
5sdrNskdWDOLGOuJY0QKIDRhxXMhcPWNQ0nzyGx7J7OaIFB9w6cdHwK6VEcB4/64bqb2DC2n7vSi
v1sKi7SJXtKVWYXNTpu+IdvbqGZqPhWA4M6A+8/oxWBMVYxehDNJUH+KTb3e4mts2BvB5cyduuLn
WlAI+H8NE5O8ZCA1OcUy2hnD2nDzGnLMLRrvwNR1Uxf92PyPpWnzVWouHhdE5kHJXZtc6NwgYsGS
r8s78qdWrqgzBTsCSewS+4u5DnCXWMu8U0U0OvEGbe9VTmYcaIE7+nTw0004fTggq1alGV3hZ0AO
flkh5UuyZTbgvDP16+T6HAYhouigBGQtieXX8+X8poF/W1xVD6cFEiXEKpsK4PjFIkOWvCbJd+Ul
p+0P6F3kNtU/lPUnd2lzSkF8O+Ga9UgAJL92aQMGs/HUkMAZzudHQYta2+xe/ig8gR+0+ckrqOB5
fF3J/8cv8x30ZEpOJtA5rkqVfDqKc+d5DWYdEpVw2SkDXtZTfHkbPCEQaqn9OiDLxJjr9wfFmjbW
wlufihgeMnaZwk6Bm1J4eGITOLRUto3ltq/QWYqS61J7jNrUxfbKspERCjVTiDbP1MNuQGRqOCCZ
eCtDILULSXh6SIhGM2ibkoMWWSe7S5FE7rqmoQJCThBJ2KoyrdSGf+8Tp8oB/e1QgYImucsrq85y
dTciOBz6SvO1ScQn8vNF4MOtdyT/uviucJp5ZX6Yt6Su9vq1U2rfJU8egMvFMSpxSYzRlYRmflWy
9ZMYmKZPhyNVwdvujg8nXSF67WvwuxmWrRWTncIYC+zWYpETRoHgcGAWeUDJnMVa4GvjreOvK1+b
ymBkoKmhfArQPc4SyqHJLQ6rdEuqSeTTq3V1VYKE/qLochmoQVpzYB/xQhlP125tn6KoK/3YDEhW
C05AKlcOFUSkfwqBfjrShlb8s7dnZZX6YD4hemqtBuEetLyTn2of8rzfgA1HTMU1uRneTkf5L+OR
c2gLVqqaYGv+YF0GuOxQIksKDOYQwHboPNPcT43NKPxjYuvIGqxr9fpE6MmWV4xDv2Fg05v1012t
HP/JtI3+S+wjaUyPyJHL0L2PmT1bbqP51XFs8u9JsUQSl2w7x0ygzskpLK/eJCDbp7onB0sWN3+6
CmKM/QCvTlHEA7FkhMKN4yRCSyPry+Mf0qt8tG8IhN5KCLeqB6Zrq4EPNRoXSJEJCPrWyQ6aPpbv
TtWyBPDjmhZhSjuTSw2XVMMIvkHz9ZGH/cPsuObTp9dsWC0xuopqVi4DsmRHn2kevC8m2qh7rLTG
3XJv/iY/tF/Vn3QAyGk1UHh3pKVRu1qv4oDNvuvNVZEFLylhF2XsVFuJ6+PKsXVZPpKvz5wLitHt
7XYJ0PhFmj+OXSsnwkDZB5pYrIZ01vvFY32skufGbfB1jwQj/6EdEdXXLwSlHHmuJ0U0dPA3nkLu
m/U8+hmBPyIDaq88u2LzHtujGAs89BX/mfK/r5alQirmeRsSLwebMDsQVnXuUEVicet7gxs+Ui5T
9zomA2AAhYrtPRvRl8N7mTB0YE5ycolEBXaTf7TYm7t6s8pL7oYKS2qYMBVXUHvrpdrIhRPvQQb3
rtcRGjfcrb2ScnEL9wvP6gjh0/QLA6nvN+qWV/xU2Ga+i4RCq/KfQdoOJwYf5+bxryvAnFKgvydv
U7q9onJVLIqTSXvrPsl+c3yTmbip7E+5+5jjDIQbmRTYOdXFHm0ieZu9JkDuB6iZBctESlwcIca0
QIq07+RPIi2JhCusB7iCcVve7Qkz6AWFb/Kswwi0tgZ1/pju6qsjHK26ix4kLs9lmTWmfsdsna9S
hokDL6fUy77T56fWzPmQoXps0sgw9q8PItAHT6lmqWp6ykglzcF+12y23l7kvK2RHV/I9w3rdY58
bwWVJDQtJ1uwqBvJcTB1ysm+eIxGtpFvPi8L+dGC8uiH37ZAwAb28MPCrA9rI2aaZjv0gtiGtW5K
G0npoDxOQFyG1QtYm/uGf6NR/uBbjrYoCQ3+VOwy5HJY4BDRtmh0AK5N8c+B4TBR+p80pyqXOEO1
zFgY8LVtqcNXN+h1eJIPBwGvhPyVLqJAH3Y5chOzCnJqUECV97cxX8Zp6raW93GzzOShy12sUfKC
NqJ/VYA2ON/9mTP3NxzIABKEC+ak4b6x+AwkNecA1V9dGz4ht8c2cCgV5JLIMuspd2cJEvp3PvZF
SfG9xdJWo0+3nPONVP8h0eTNTAgeGYILZsHtIcOkGlaDDcdJ8vNS2cI+lEepydMU4cxHwHUbYFWK
0m0jfcfeUfQPqKF250TxBBE/d1PVmnNdF4P9ANDW9hzm0CwRDDncc5tSG+s14yLdWgRZHRw+fNNM
jFoQYVuQgbsYGeXc14IFxgOuUOQ9SXqntiDMeajJ8JZCCuv5Xlw47+ar4KjS858D8ggjhddKWqFK
DyZu/kySmVW8pOcgJ6vyRSDpXWRSd57VooG9u+qRZ205C5m/1rp9UNi/fS9oTqT0SUk+p3o2mlXt
07uj/79XZ4aBDKwzxbMEd1fXV7iZvnNEQWPNyZY6YL4LMq0VaTOOTimEWe8JrJ+EI4eu9onj1Te8
OiUGZOXD6Dre/h1MBtEnjNO2HfT5JvcnVloqjNdM0a55tcsvUqXQkpHGWN1P3qDw17wKZ6BH0eSq
5dCM3KgL52uwY3lYsgnKLtZmJJgLf97L8L3g2Kgt64tXLG/KTW7PKJT8kuOp44s18PQ+q1GhjRRy
Q9auk/Mepw64t/Ftl/xtcnfgMqUDUOMU4Nsbflitu7ykbxGhAiagSOih0S0SkfxCDlFV21zwB22V
Tdf2Ni8EtNoMhSYRCnUHFP3u24M8qNhjU/3o/lBeToBRFr6LElcfjF9eFu3bM7jpgbMHlqcAtr19
izcSuVHtRFUMiUefyvCih5+CU3L5h6xHO5LGiVpPtG9y8S1VyvOrkVM8ZRVcQ4FN2MiMGrBYViD+
oNzmGu7p1UHlBdLlS1DjbTWaqKtip3ICEirZ0WlZLCQ1/kYRQu6Tu2XqBlbf7oLUuQy1V5nP8pp+
kEIAgSsM9FbtSHeL3zI/quhFboGZ9auoUlEo4AMaqdrzqpqClusN0B1nDJIvIif94vfSCfuSArgH
SCS6cbxPvozT+X5jXB+b4d8/Eo9oDLWRSP+8AFLD8KdTyF2SCBfwH9xLnAbD/0dAZo4jkkkSrurY
/R8CO1znU+tIbhrnHWZDrcrPUSBnovQ89Sa0y4UZaee00hwewBcXB7J9nToWJVWuquciViBPVfO8
Eva2sY0wVR/3T1mqo8mJsPjyAwENM64JOnn5nFPtlClaZewWc5hiS7qay9+L7/fdsFcwQ4DlCI7O
SgIPPzbw5fAqgx4yOb4jKL7Fo6r8A1LuqGsbjGboXRmyTyY5/HbPpNs94s9+ZJF50Zfhnom4fCEe
nlRaecNOqtJK0Nlp0xS7RBRV6eLCLB0hmHpozI48MF8OnMpPgJtWAqEl7z9se10728fyfpdt6IFP
7/PeuXoXw5XQzbraa36jaOHmLSvFFxQ4a59nuGu5V3ealNQaPcuXv/zC52klD8Kvu7ZrWeA62yaq
43YeWcshZkQEvef9HQL/Ah0bg+broB/DJJvX0dpGWS37O+WLmSboUwhQErKw/tbgLMFZU3waV8ob
ULMedpmRY0HnSPz8jmoXGUkhzQju0SwJu5SzoI90nPA00AQzD4gtlOD5IVsMDBos/8RYCCbBnyoE
H4VoHWyznI6+YVUql84U0s+SEXnSXNtR7yzglskyO2pN6FPe7auey9InNZ6P5yWiyFv/6LG8gt/l
NqOA6hOcaNraeQdNF2765Jcjqbyl6OfeA8uXK4a5XUsrBdAuylcB9lTcFi+io1unBKK2giF4NgjS
lpfULsN1j3s7RbiowenrfA7eDPo/onwAILOWFbqPtpq5UovN7rpVO9gIDQ0JW3D5M8wl9+J9NtnI
cavXvdauobr/6/xyTKcZ1Vel2CTQKq37fb0zde3ojWocxlF+FMUjiRkErmf1QLaSgAj3UdRzYuFG
cTDEovl/pLnj9ZvsZqxMK0yfujSzL9DCHGkBaZyh3gUAWLyZpk/DbdnB/Gp9RAyfvSSV1VnJ59GR
YV0om+/wu7TaaLSFfKvgIPD+7hMJPHJYhO2pMtmJ2cVa1Ev1Bb0uRFzTz7kryPucf3mJeAsV+OOv
661T3uE80acz3mW/IH6XeN+yeks3X2nqtM+/Zg5RtQfjRl4boOiHD6ayAcvDlQt18KkJyjWfQw0y
SaCe72q8nJEmRCHX5kHO9pZ2uHmAxP3EpjuiaVB4gusjrRLTZBb4WjEH8b4pEn9f7djj/PWDLarN
HyS5D3NXVVXBavnPXmTKAXhPIQdPCz47IohLsxgyxktLHYDSZdCy8Y9hT2C7aqkZHcQkX4Nte0/b
yAJkjOV/qMJmSx/8bb2Did8yN+cbXsuDgEjaHEnl4q1Uvpq9PQ3BqZO78GFu3LftSTiT+K/NCWbt
iTyopxB4C+9SmVLL8oBKtpfHuvG0G1MNhD4C+7KRPNhpbw6MrKV8RVe0NJvHPg0Hc5jwcnVGbZyN
M2Hez7QmjOF16IKHuoMFbk351gYPeoa4/yQNC4d+xxcc6dgcbv4DEf4VKn/p5UOSc9hJoWhBfq2+
nHIf2lvTC/BHFHrzVaUJyKmFHey2/1pjA6JR58w2q1GKrBG95edhXVVgq9se7Onzs3IVOgmC1UxA
7Wi9Vmiio1Gs2Cy92NqXnWYVbkfamcHa3ud6+G3YZtVvUe9eiLLoeKB3Po8pJ6Osj0OciNtAYuQh
fHAdyrZG0yETk3A2K9NATrIFSaIBByLdJ+YJnisL/DiL6Hc8P0caYDOSVfWk3v61vo1VZ0Bt/K8v
MagycPbQEV/Vy7LlnUYRxqzC7LStT/feW8W1lqA1QpyQiUx0qfAFapmWO3WSwEB1rBl+PBg7MqV3
gmIjlI4zZ3UiId6L9Ny5p61ibc/484ghJO52s+R8Y59GmQVAEABO6sxCDsIr9UJureGxBAIaiyrO
CsWUB2gEZv2u/r52YpIf9Uj461W3ZllQNy1LHTC9wxxXvv5OLWIpmGj9s85QHPjpLHl5hLk68+Yj
UedcBOcDNe8/f5YmO8kPM2XTgldbCEnXw3K0tAKkFQ1L0UEWOOsQwLsIEz3S8BBkqj9TuzTB63bo
Le6M3N26kvJhkhsXoMoWYsYmk+3cPVbZ0VlpJkIuDXwx5aNdsiJ5XjJoDsal7o9NueDfH9ChVmvl
62KVjN3lzDZDtzZsELVeEeYAMiMi0FYF9jWIwEFGzPFzIJE2gQ5qh1QWKwqig7puldfJ/Y8+pLbU
Kv4pFh/Q1xTe9NMdv3L/D3IR2A+kQRvuiIoiFghyD5Mz50xdRTgt8lSzOWuKlGt4xa0C1oT75mn8
JO4wIzuJgvL7ss3chT0qOrcwQk+d9b8OJxe/qw5/KzGeXKn5qHw/ys76eg6D+6m/whO74mI9JCTo
KfgS2aNapJRdCKa0P1CtXgmXKVxMBLBe4fNvkgGrQ2+DRGq0CrnJ4YS2XQ0ZVDCNIyP0iPQHmRuN
3wtOby6Be71HcWg6Fkh5VIlVFDZA0dpyncKDPL2TK2Og6YklLQJ9IqkoKfZZ+BkkK4lbTHUZ0sYs
rmJsALUMj3i8KKl3nkhXJft/N64P5JkP8x5l02aV5QIRN1+RGkdilI730jJ3hUuX8+lENUVAjD/t
/WZg6MtPBWcrdgprtFIJXqm2as15FV1MmqNcPMakptQ+IvDgc3YsNlX/9vjUa4jsFUTdDvqfqF6v
cjrHj+WuvixNzDarFvMNx5J/DeBabqaUj2U98eulC/jTzRPiQC+GUfF9Lg9zHaF+NM2OYl2e9TXL
3tuwtn3B+hzl61ZWUfl0/7wG2cJvE/yMw1DgjpdFkY3YGJsHCSNeEWoh1f5O1jGDj65QsXCOj+1G
yLwmooHDF6cfZwZFtHQrUkS50+ZQ+JYNV680DYLsJBwoXI3nX9z6fVJnqH31Y56BPLEkJgEwOloW
0kiyy6XqJcWHBRsI++B1tcFKV3ohUs8ZxM1thN0Q3Hb/MjyLKDrPt2+hyePSiGTf2ZAZ6jO3Lt2/
x1HQkvgAPTyoTlFnpu1IXzqfzlI+cUGn4R+baluyv39VsLap9oKEH737ScI9pT8eLUlZ5mbIsqj2
K4rFopV1sLIlQk00jKytTdiOz5qbnpIt/rB84E3mKHgDPl/Fy5PwDu8WuyfR0tg9193V7YEndQEe
yj1mTmrtB85hyaLer3IBfihAUdOcNdN4TS3eTurweo3lHPmxTQ0zjFRCq8oPuyk6NSYmLra5JJv4
nLWmj8S0TJgzBGTruUjGhDgn5tdfec69Cshg8wmhyxlOfBKZfgTtHjOLGkyNgGP8B/bvdtVCD1rW
m5T5IEGYahYulCUeeynyw9/ru5OFsbMgLtCtxkXxpDob5bbNQRlphQ1k6JYEMYVfqCn4zQxAv0Zh
BqOFZ/EvNp5C9PrLcEAtdKSVXhqQRCeUnk9/uoiZfi9TscmJPA9cLIgWbgeQX6cHxgAlXhJfuwwb
QU6LDHmYtLywYvNKxg+2SgK+s77m7GXQBozEbeEJDnnqilTsOxSN9uckxFr0NQgparIISGIi47ET
lxTZfZf8hwITsXlPmvfqCiLNhHVtqHeqSpYrjRouvy5NCg31PaYBZuHCgz4G4kcqPgX6XPlS70CK
CzYxMCnOpB+Bdm5Qgeqo/8p5/tQ0i2z+FxSnLkkQ+LQJCf+b7CNmv2xCiL4m1jZj+gspGdxeVwhA
jAOh0fVLdWihPag0HEybdq/wqnHWnEKA5S9/dY2coiEDF8qtb2ZoLZL3W2ri4jZfS1Se/yVeYu++
y8/4JsFxr6UfXdM+FSkmAoP5x4xviPQ47nlXMaQuyYg6HKs9XgRyQklVUhcJ6PyuEDbuhjp1gJF0
JmyJbW7JR3i8XqGtz0Sk6o7+Wc+GWL7UK9bgCWQ1mtL9nFyDNJeRErxrRASE+74iw6IN76M5VA6a
NDVr0WAZ5SUAk2lCWVxn9JIvwERvF94IDAdQrJRRvaZQGEfqn/t+gGw+QjC00pQbD4/nmmnSyt/T
GFFVpEpv16uYU4juOGD5y30HopdAmKOZqyO/GNhA8VbQKUi9ohYQ9NNYx8lfUvW4dn67jVbai/Tb
/h0+zpF2VAfNiPi7WqL6pcJBSIEvFXsAcxSWue2mLJTSnE004sIRJvcAaXv3F7Un0yHEwE7nqzo6
ZTPZOEVD/Ax842sIAqBAxmIu+wubRXpmZsYSu7Cla+YMAhXDnlQDILyE928whnbYzSgbWsArF9oj
ec+OUhxQATVSBdoMLTOuxgA+Ju3InpraVOH6+VBOWlm9bVlbT/i6V+nzmroQzvWtGh4BmnYC6ldB
ej54AlCK+w7Wyt+rr4oo3yZMbzB5VkyLAsjz35IhKoDGXfd6fsm7Yxg/4eobOTeDllGtsK5X9Wb7
8FDngPKJnisxcnv8TIlfW7l1+mhNaRXaB2dW+UnWUwkKRj2oi8ksmnZTK4+N0GT1zACFlU4XQyh4
S9hf2oSYjg38XsJhBSo3sKnZEyWi9FzV8II8S3ksb/Dt/CVmkqZnaDBkzOAS6eym984bAs8jg2D/
7+4bL8cYnm4nj1p1Nx1j28qjL1J1cx11ttdzMLmZRs1hrrhjmrstZ9Xp493Pw7L2mTbNkaXARMdl
CEP9BTxjZVlbCLhZyVvBlnZFwmLnKvADvcMODiRtJWm7ShzANS9rbyPr/nJVdgkYCaTGlyCvjU7l
OQ/HAEBGvaCK2cXmnLxp6Emb/4pZZ/aqNpfJ1d0tc7AM0aPTUmFLqPmr1Oi4LG2N7WtnD36FOGNp
lHwXUCIfHTy+RKfPTPCpYWK8TubUxC/0coaB8KV4dEFuI8KS1B1UMSu7YbGIyfXNnSQZ++XFfrhw
P0OMhPf7GFk473KADead5DtnhocRXPkpm0ak/qzjjQJysQ4JIOidqrdJzgGB2/VcpNuf1Wy2+CaZ
35LnZmhhsWOXMfTGjXXI1XQ3i4aEPiYOfv661/NAyIvVW7v+enGaQ+KNERYdCISsaPq8EnBOn0Mf
JtxaWlgoQfEORYIPi+qUSd2yOHDot/8EUkPvfl6cMNzvRSwBwOUuX6hU+PbE1KIfAABkOL/cj4S3
iD087AravlLDzMYJX7jz6IZ1wL+Ml5f9/150ZgFzAwEd/OhfRKxd5FqXqzw0/im98PYCvQk/s5k0
8EniH8x0Pk86GIKCy+lRRXuoxc7LRL1cEvRSSzp10f7sbSwF2jWGXOSzk8HWKcn4Zkk2BLx64wa8
ocAXX2qSNx+fBf63cN6SSOXrqmRv+p3hIJIpeUktaCkkZ2z9VgYJzeAtEzw0yzqCzv1DY7ewWTAn
lc4/7ewK/LWvd/cFjzWi8uq2kUXtbuL0sUa2f4cYOedJSBGat7QpoIb+YJPHksuau9yuSxkduuns
SGIxEKe8G/r1iMkdRMPwHvSXDlkzROzCimn/teUWB1tqX/uv2KyGgEbGjTz9ep7Sbzub+2whGXp2
URkxiZMcdLBFn4lWDI5JxS1/AN8tn1/gx3s8Csp0EyJLVZYluR621bwejWyOOfS6hU0yVIwjwADf
9vcnxfLjB4WSnz7bHm2neC3CczyZ2NtmgRRZuGkYySKAGwDXchqfUAB/Zcy8TEUI+pyVhBoVy/6v
ItftXTZtuVGSy3oUm4pmdQezCdtoKdzKCbbwrnYehWAIHCSSufNsPPGUA7/WfmyQwNQ29X0MCM2P
sjogxvefyyUKmkD9QU3cGFEARz6ow8EhNbL/1nWdAZFgldkPkzsAQZxZIMxy1RXTfg2oh+PaK/n1
ABwxn2jxgwqRcaWGyess9oQDZmEayGawc+L4MC1KRkVk7W1r6N5YJs6RMIRkPQpMyGnMr/Plw3RF
U4txXIhdUHAGBYiOXf63CPbqRIe3ys+B4/AXbVMqi63Y+MA8xpJk2veM1qAF9qAOtAT37iqeXu/t
D8r9pMFWVAKnM/LXkIB6EXQ1LUTQnreMUy5LE25gS6oB+2FgSUZAC2HagCVaDTX/RTmCftUnMkxb
1q11YZJQEMuuZxtflmKZavpYv8yGEMD/Ha7KG8HIWZvbb3XC3PK3r4RO1gmEJff7BVTZ73CzxO2W
EOiKDtAbmETS+qtdbAhI34nJjZDOP3hxiM57FX5JoxM1Y7GuAiig3djrRP2MuWzzDDixlqdZA1Db
tvxWuvf+Iemg4oNule9IZXzkFCPuXHHpfkXOUWXPxqvsJ3zrHsp6S+B6EGt1YgcxjyWe921vf2pC
hdUfQzANuA+DDnmeWFcQ/NI6LofVVWxYB0Dl3Qr9nm8B/1JB0ajSTgSRoZxrwNC6+Q1AxIo9XiDg
y+V1SxF8xqKwVS38iB2zBzzWACnGBkBhb6m2ySyL11Wqa3o1qCUoPnF+WBd9OtPTm7tL5w+9NAB6
JZIqQMuQkYoK/qsvfoQRawpztjIldeXM+JPQtKll/0VvBaCECOvzlxsZHdUFJLzsFmFUVRHeZSh5
V1qK6jIuV8n3Duh6t7Tbavm3W4jt3NZyJEQRlJsE/eu0UuoUeeT5dLhKQ9SuwvVC8EvqRPvgUO/M
lfUV6mitGbPAWISCj1WuHyecBqB2MrXhCEYb+D1nvxAa2OSV1T/hgL5Jr+ON8hCY33rxiuwQL7MI
15vFgsCsUuiitQ/hz5t0udznhs0fl4l7RfdaafXjJP+GiZ77vZmoUtTnQp/bbN0zOLAnI06Nq0J9
+LyeWGp1Cc5zuOnylEi63uRtka7wuE1mtqiyeoiOR0r+Kbqa7rcMeNGOBUMg/VzsUNyjwFJQAAON
tEjpaB/fm+ETjZ/r4PKKy3NmDWw5j0LIkGTjOWuAYcS0RecwusTh60g5HVd1tvj4aPa2/xGsPN/X
hvf90xPZNX7Nm2qnHXuwmktUk3hNnV/NcZ3w38okIb3qXcHCtp+5fLNiCKHDOdk93rRQEfI0z7KR
KRohAUHBX0dtLAaSLWyfU/Ao5wc6dxkWSO+W8i/gUSeoluDemMDGzr8dYtKCQfBtxY45Xt3oTsgD
o1jyCCYgGb5SXqxSyJhFEO+1JL0UWrXqe7scAujzXyEIGIQNsUvJtWGToE08ild7lPSnKazQ/7uJ
hENl6Es5JmaQabrKJiC55BpZveyz2/2v+1G79wP7JBmjx+62P9e22Pfx8Ycv4AAypkMpsoTcy7fv
gaVe2k8RO9LZqh8BWnvgMWybAD2TNzaW2JuZ0IjKU9sUiE27eX3QJLOkQcDsjOun1zm3ukqrsQvp
2etti6rvea4+sR2a4C/a7xeVg0dHegJjA2vdIkqVEj3hRyLBGqthaHXvs+IxlEYcNsB6gLcmBrAT
efFSsDTJhfixz0Wona5WnDvlywuGi5BHHm69zlzF3qJE7R2F4CNQdl7TECuoJ2gtHAPXmn0HU7eA
CYQS2k5wJQ3jjPYU0oUSE2oXTOcOW5yLyDGp/5QaD+b+TXPM1ASmTsD3PmYRwHXKgDrRaPSz81G2
WgtsRqHlcrI8Klt1ZaZGMDdk3qp1caQTe9gFDf4sQmZDVmlk9AnTnuRsAl3m0Qf+BLp7uTd3Vlu9
9odHmi9rARlD15TOSjbrroxlgcxJKKuRdt/KjEhVzADyLd5hbdFQ5OUHooTtQlMcQeSGldz5HCAf
RxG1Qkyc9qbZ1+1Jil2kRUzR9WhpfOSUWUJIg6hDoEmIwkfhogKo4WYDUg2whbBMv4ntJarRYYNZ
4zjVARssf/COcSJC/uPY+1QjRD87PI0RLPdfyIA+RFy4VwFbe4I0sXHQBHmc5HdVYcV73muJ5eTg
Ez7Jl8nrmEqxa6zULSID+CCnfLQvVbr7fERGgfo73H1yLUTPaKmAEJoVn5eoon/OlZ8GivbOs9Td
NnrjtRTdRa1ckol2kkafq1TpOFt9uvYSUSnH4HZjZY0oLTFyMcNQf5KqurSxLfLIRK4ZITMTof6w
TISNCq36uY68B37QeokVx7u0/3LCXZTka2qhs7WekPdnJ14uWg3N7eVWYdyqw5432s5KEuxS2Zbe
TXo3hLbZB7L3s6bevDAitbvhZNznZlYvAHnrXplROkSD06fKBX8NJuz0TykSpVYxpNrcZSEijty2
ivUYXdqPdmoWkV7xp0qrmbYeeF9vIGSksibnxkKrdV+z91yj5lEyRGrcZZOkjT7yquum1yx8kZAU
PSdtIF3wnUGOKICy1aUzs2UewN3eyVUToIdS6dIafRCtzXmkUIvuoo4x7a1tTHovtQaRW6/WuJiC
4uzM2lQqe9KUviSX3ZbB84/fJ0Z2DUPctHNSF9mP5ev8EGSnjFm89ib9CyJKae6vO35Txn7gH7qe
A+UQubBDqN4TKlUuEn/zXKyjqT66WBPMi8yXLZ3bxIKJgMWPeOaUQvv963eEgjshRlCdQ5Iu2Gkk
LiAg0gqR0da2FUu4VMD3Socx/MS3ihIJXUb4H2BD7yIBxR9WBHEvsm7zCdRPRyJXQDzEtcyq2y4N
oWdtPk9WmXkMMjVUn/97kdacvfnrrvj2CRuUNAnFvc4UgL04MvxKEwGY8CT4MwtsfNm4fBGRaNwq
yYVduwPF/SnT0uDu7Nq0M6hMkDyK4JhaOTnHjNE0POiybtKJvYaMs4N8uHzPy4G0PodpFu9A/8gm
IzNI6+bsCm2l/rZNctGuJxWDMMs5L7wjORv/3o3vLnceoFBZzy15Ha+bVA4xbY8oosu2nrmjAD3F
gTF7agPiIWcrxgurnMMaVPR1nK6OhHudG4LT+cac/kteRwQelPrmA1dwqg/zwvRkiAWfBE+hGE32
8XlEVMpCa491TQ7CfzSE4gryt1mJIK7DliKjZPNGifKuy13FdJbEJ3zfe5WmPHCB0MgC4q9BPfgo
+4wdfSlhRD4oBRU6mCpqhTq+lmLqrS/3EJSVcQOP1nNKXaFnvSuFm8/g1tKurfLKwi6Nhrm0Gns4
TWgmcBc3YoLfHfMsWqPSjNZMgHfg2JhGsKLtGlBKH+Qy3qaxeoSAPUaS3HUGvv78gdr4OEsZDXr7
iIE5TqzIqg07SCx85sBVFI1yHJM2QEe95BcsfNMhDUS9lppIDQeDc7XwpL9I5FhuCU1kYla7D97h
tv4U3aVhCX28ToMWrA4qdhGs4q5gtgreCAV1jMIelC7eO1m0K7fF+3dlab/OY50ds8vYrpqPiSbf
LdsI25wbUWLLVCUbMLgeQ5D3bbnyCnv73hKWpAgbo/m0QfjfG4pk0pTYmgzYdzhF8iVDIaL/jz48
fbEbL3cb2YwsMoId3OWxKTayKe9tywhVpmAlyYpLdrNAo3dU8N9aH5+fwma62SjPQhQxoLClhSsM
8aJJRviPMbYKsRBJmeqDP+fIhyDIv8AdpGD2qxyYJ+N4E1z/Zs+vB2XA3SzuBUOB8inKV+Rke/dg
S8irk3hy4HICUFnKCsEYv+Ct2PdNnXqPrcv2MLixWHDcdVK5JzthTcH1PGC0fymIBm+uMBktV4Dw
EOIFce/ZKdVy0AwyLNxieKZ0TY+i5a+tvv+hMP4zR050EEGFv0zbtBTbUnGRXmYh0xiiuITCx/oS
ZEAwMrmFt/FkdyipEmYnLlwJBNfI5cERlcVfHZjtWtYHc0W/Lramdla+uqI9q0GcH9JI7rbPyUy7
bhi6coAAL+P78Ar6kf8AXxGHrcxce+spk6LnA3TUBeWyKCPfLBz3oi3EZ+qJ3+jfvZ11XcBbEi4O
VtZrK8w6APfc+8gaXuCpGwt+uSdekP0Hyxyn/g3Ziv9eS1dEwuwlpKaurHXbPSYzGEee7i30Zqhp
NAOgCVahP+kBkc2jmsKxv+gfn0JCD2bVQ2zlQmflhG5SYduR08RQCOIqML0NVM+lxlbPCoaM+RAj
ReO3A+X1IVIkuiit0T76x7oCBFqJehM545qNRzkU1HwP40TQnYTVeOj11kmqhhOxZMctYTrbvDSY
D7uiw4srmRFtiMYQSUFRs7EREUB0rdWngCHxjhCcHyEPUpUMIhhj51Q3t3MXj0HohJyvV8tNPjgY
42PQG2zeAu1JO9EuGvsBy7m8Xao/L5D8CBUVszCUmYV1WhRHb97PIdmplhmRoYdepX7x4lUYcgmT
rIfRQyvG5QZRrPwH96e3jBqhq/bPfDWjuspvQGuEV4wsELixUd4rIYOZX7LaKeB29cr9w5BK+HmX
7RmIZTmwIB6vR++l8fmYXvxBIGhEvU45k7MVjfAUXdt/KePEXw3hRdruP+2f9OG3FSiLlxmrpGXE
hIId75MR8toyaw6oojf54EoJo4SQuzpPM9hTV5R03RRn0Uq3AtHZCUkxDPcbIqGJSBYY1BA9Ex09
jKH7xroLiG2bhgnYyNZOs2eN2lKUr/Xx+VZHB4cBDj9fyj4LY43CV8zdq1GDuPYv5bdbo0I1IuNy
05Q2ubnO3bBdbSMekEaD718mg7BTFE7oTRhWA+Xjob+007Bbdb1OUH6vF3JbTBegxJuEIulDeOl9
fMV5MuDQJ3sVcWuMzNVbWvS112jpnoIH2GhWz9vjz6JP26ap/lLokgn92WnkVA+qr6i1F4ZmNXuy
uHnVdPtCENIlO21xR3oP2rwxynrr4d4iW3AMFR1Wp6b8C7kwHYy8d6av6ZdnJgiL4769C5IJKkJS
RQ2M++/eTJTCNFfJ4SxddAHcyougMRDpCxb3tUGwgAnfuc4w46pGxflosZI5AFg7kH1t80gls/j+
xIICeWtGaYPo6jbrR8gYsP/7ZPfCEuyrCabMrZK9vy5JD5tyvGo9a3SiwiPpXRxuIvFDy3JPAxIj
8mM2gpXtNAzCLxelTYNX5n84QphHMSYLMe4KGna2EFFtYUHThEBojMTDBUGVsTEtqBgfm49Ap7BS
MrTmggHxXjSGI2JIo+UN/tSTKf51/9PxDcsaCJeHqLE3MzFe6qT3RudsAqk+4lrEdWc85iSMdsx6
dXnb986eKPy2CO7j4mU/WumnYvOHqeN6qm0Y3RWda03FiNG+oU2eOVH0osmLebNti8MAfZm8iMXy
gMTxU+vIHBbJ3y9nLxO59F+ijaSGmgp+IblkrTpibhykorPeS+B+PhkTEeRdihmvc6HqZ0Gok89x
VuQatExvIXGfFoSN6GhZ0K+1D6ik7KK6jyZtybwAK6xUUew1dSm1aNy/DDyRb/jOow2vli9qVg5v
yZ6Qito1P/KHXWp8PiitXwmWse+ztKoiXB7x1mhiDHc048qpOMBnszxSx/sJYXkfzOL5MWyhw5/4
Rcn1AJ02FZ8OkoaefhUodR8gHk6ZRw/eToPcb2HX1PysvB2GQoqor+DjLyBxpECi6Ix6SUqk+fw+
Wp2ubxBY1MjNOjb1baTTQQJCS0dRpoA1sqsKv7gh45uGKQQMwDf/IuzcyESP6vDQ/t1Doosz8unF
gKsgpir2F6E47z4zcZU7AaASafDQvbCjdZWvrSdc1IOj8YmrDIoFku+LUEqIeBDEywD5B0AcMuzy
OmcRdz+FzJImJlyIgLYZINEO6uu5AaMuNRO/ToRh518keAMes2a2d6Vbsxn/1m0k7EdeG4CsftXK
hdLdHFPhcfIazXFdrNYJ5jym+eU8Y2sQlNI1KtJb59OkH8v/Iw20ZlrFgM9tk2Ly8gERnNnQhkXY
xWLrZdGFFublxDGbjgBK1ct4q+adznRdNUOaA6SUP4KDqmTInQiS9kW30SSp5NATqokYW51g9Gzr
hh6vY/I1yzIzNanWrUacmE4H8I9FHGwwQ/e+08wgJUFSgFz+0US0oGACaCcEEuZ088Acv5nOuUh5
mh7WtQNnba3uAxBgP7RAW5NxIkcFTZSGdlOd10iaaXrmn0kD272/ACpKFD2pzfDQHwEoCbIbEKuU
QgxhS4ik34awTxP84ZVHlu/v5dp76qUnYhhk2YzlBlj74/lxD995EN9x+4sBmpTwF2148K9izVF4
bipdVVndJCX7BppOXDGchWRb5+Ju8qjolOHZWhawCFVYD3eWggY5IOwa6Z20nMsvgOoGCvHY/+3U
jBlSrQBUBEbPZxk3xSniuKNE6h+OLmslwx7q8LtYg8cJidRqtegwW+k2OtH1kwJWVvX36xWtryTb
txTnmhj6hb9Qqreh9iNBjBM9W1Rp+7fxx4knZ8AOKmluORVe/hU57zMmF9iBu7MojrPYRSkqFoMZ
vFKNK2Z3McqrteEq6Q2nb/xvqYDS4uZl47YDzACw00us/pDNDB+p3J2ZSSBk7dQsXTAKPQfs4B6I
5yyLnVSnrxMU45qTnGIHm+JpQqBMFq2a+weBy3kQy6aH3tae4i9vaicjvn5yEfR8dQEyeStw4/BS
2uxCcsaICDwuFDELYvMxZCoPs5Ux1QR/hOUn8C6+jOysJai4xqh4d3iLX17vn0ZgQlxrHXspRg9z
D5Scl1dGL8NSIUHxMqCQRZZFZCmSngFtVCSOyhbsrjeE7cZe9vy/HegCUrt+hCmIcTd8YYdUwyoz
dwuyA/8an9eDDecTwEbr5ptbwzKhH14L8hNJ20SvvBRmBKX7bPAgrY+qF7FEaQxPzpbilNoVnTex
mqrn1tIYgpKmVVnFLwNlHD5sqm3BsVML4G52z/kdVojFsttq55jgkmYUZ5rgSwGXxEec3BCe7wXv
8FblXYug0GZLcdhuRxCOeVaqS1qPx86nSVPtCI5v2PXuHeNVx0Xi7gY6qE0gpxXrGjtXhuZQeIjA
tIK2SBEEkXbn/XkWfrCaWBZYmrRyA4/EqKHmQo58AUigSJiJoY6NrDTNoQWOBKJm9eRQtxat/Tlr
aPCj/AfepCX53EeqoVPZY2+5bRYZVz2jSsQ/OTzD+sE7tjJ9jRNvSq19HKpld2qCmCq2Nt50398M
G2Efqdj/4SW/9jRby7nlDIgQYbnj2cPH+D0RUowkCmIZF3e0qgYfrdUK/B12GTFL668AgufS3eut
OOQgAxGsnYdJAzr/h55+fVGV83W5JSqjT1ILXFelp+MzzJEuAbkGX80HicEzVOgS5qErO8r3zEi6
ytRz950OE6FzEmdoAG2LEBrbIoX12pikfVP/YM1eTwqjvVJQ5w4oho9bzkCEaMku6GX5nqtzNWWd
UkCD8V3XrJJwX60p+xZtwcbQ6mNDnYyNH0KDOB8KB9Wb8Rv9bGZqpmIek39sKUE3laXFshr3uhkp
6a7ePLCru5lGiGwU59lwmaiV+F7hmlIjZpb7ipoeH19u2t+vdu8EWm6/HTN7DvQm7SBy7SVXXNBH
ybNZInnPi4jiNMW9ciTCmfTtTq0B1g+x/uOf6HhxxIXxKfS23AKajzx/h+timkVOwRok4IiKEgcW
Nvr7HmYYzcvKPsfjSJZtf6UFfYJJsZZi34zkvkP4WcYl0o2/I/hPtbmrt5hsyC6FwtSG+Fon+cl+
3aTvHy0KPyCRHjRuQIFituTlA4BB0gTtCKXbEcnMmZk/OuQyrjxP3W5X5PA+2W9IIDRDGJxiqsBq
7axP3kkyLMHsTWUj/mjH2iESkpySmjMTGKTsbnikh4NI6RvromBv32X0mPF/rsEM2t+OwmCDIBG8
KnvKHsvMUOVvmACQQ9YWM8LjXDAXgRTfl2kVvoie1/27bJLeFRLp0Sv4/nInqDHpGQkwZPEtlJlU
W1z5348cQcZhltVfWa9ux77TmSRq/8GTYKeBIxlgaMlgPadmVxkHLtqcI+ly4RrKvO8OP7EFM0cu
U1IpaCJMcX9LmHNXSLqoRWXXwzMVR6Iq+ttl7fnVwWHjBQe3u5cOd12AMGPHKcgfXxE+YFhSzyqw
xFIOryuk5HEN2gxpjmlcckuHmUlyAfDSE8SCIdlv2M7Jx8lJe5I7/5PkvrJiv+BGxa7pUMnGQxH+
f/zRGdN1dLebstXvmMPMw5rOKhQxKBst/tsSb55xB8qmz0QqYxsE0iiCtb7HGvlFTDRDLiIeS9yQ
LqD3lnGiK9gvG5Lo9pK4x0bC135RL8YPE7NDycO95Qqeb5TujkVJIH/fZcuiOCNQlE6G6XbL2mql
uyJQ9T3CXIVKRm/DxZgynUUVgnaQEpWjgEoGAzZDel+wln9srP+OWuA0BxpVgYWXpxXy0LNv/yft
quANEQ5/qhQ3z2dPTNEzMtKoRofF75f+Ad+Ufc55j/8olkN/yXhpmd+AgLTZfLWA9cp8KxUtucqs
lBByfkoqEAVvh48Ir62LYgpGfthq2h9FRmIUA/0bbeBzFXkS9RAb9/VytxhY8WC2d4f3KgrMEnm2
KXZ5WP90kRzSqWz2gHaARbsVfyHwPaypdP2F0RGwb+UVG3pr4H4NaskY4j21SQIaz1AU+yZr9ap4
nCTz/l2//9YctFSA4Tl0EFytKTBcaZCEcaAkx0OjGisrusAjdPmFiVVShhXyx78sawAHScsIBEgO
O53TBbhU9d2+3OuVc4E2c9EcEpIhrY4HSu+H7Gab/SFTcpjEp7gW2Z2yvik87wJYnBVKH53CJqHT
knj28GpUO5f6OM3QcyNsj/BhHDdPu/kIZM6xWmrpt7iaW7Y5i7sOqWHIjOXWnHMekM/oQfRjSZkd
H4HUqCU4/mA+2pv2lrpLI2A5MkeqsY6VHWu+WoX2Ay4Q/F1lHk+aKBNOHjC6DbxnAlo2514ZekEd
iZjk7BRbIsp3fr8cw5JxXkXtdpYpOQNgFbp3zV8EBMcM7pAqAibTF9SjtX0/bFc84Y8j65oSuuAm
dGkYjFIBxm4ubbZ9H9RW+jBkjFyEjqBgKo6PHE/HRWrZA/mC2CNtnXqz6uZTtAwRO0T/IUTLA1zr
CEE1ZfKky55COCsLpnHqkK0r0UFX5VfTwClRZToCifXIyLTi0kY+9AecirfEdLZoQGL9M6nJSUqL
h4qrEk5Yc6JgcArMEL9Q/ABymXqUOICf1qtAqBtqsb4SBDmU7YpjeAaUn9yHsE6GAnmHr1132IVm
B+LkObchlYlqdEr+zrW0YkAb1Yz1v/Aoz/s5N5/saSstYfJizs1rF64wg7klTOdYxAD4WfzGYTc4
YAO9OqBPb8GOC2R0dcdr3YS+/82M6+SImy/4ZVz0+LArUK1t35OneyOgia1Dx2cduy2AjE2o84Y4
gMpZf4UmMcoisyN3TxHrKmWQw4q4ze/uW61KxgU9Np+lTGti2uZ9/HFsLO4Qbhf+GSF/4Rspic6K
VtXpqftAUgAgMvvcvjIITyBXMDgXjhvPdUcsrivZgZlKWKIKCxsILZ2R4M1PvAKv6gFzcTJ5VCps
bDKAYpVtSxcYjhaRmG5l7dK0TBJKC34Rsi3JrdII4AS43tv98u6T8p2vJqSP7UXuaMZiJDReCuIY
MFgzF+jD7KQuM8qkhGYfBjt8roIaBt8ruoD0ZXNwkOf+XP7PmvNROb3puvj4ihz4koJyiLrRkUYY
qv+fyPJWawQ8R/WS/xsC5N8Rg0lOuhNmAW9ChLKYCzJrXWSmzQGkkiZzHGNSGBL+7NP1E76xaGRo
3ehcnz4oid1hIfT7wm8EDGZrJtVOJ4g9IEH4a8iPf1AfLHrDJI1pt+Gn7ySUYtMIlU/rAFTR3fen
+sjQK7N8WcxtoijFqAhdCaaTJnZ+VVR1fsfpxHZc8MphaZQch+eWkskuaUSWWUKLertIpnVvQ0D8
bOZ2nvIT27p8LdzQNjIb+uv6RgwxD2McrfXlVnjIVtfRo7qyc3KD93O3nn5FrP92ND8Chi2Qp+47
bdMZb0xaB5E9574mkG8sTpgHPS72TUOrwcfxZ/KOP4TM6LoNTR51IlHYYSPsXgudVJqGSZmRvX8a
COsBq6l/zAuFsANljbNoZeFCRLExaPK/+zOWF+IgOwE9UCk57msZMz+pDmhDlEnSrUlOrkcNkcJJ
SdsS/oBBA9kr58JcJfnNKFe/KFpkmd9qr5uSCU2DNeidxu4K58if9ZtpUbRRoJCtCA9ugfOUQEVw
mMAa1wiOoiHK+URfWJ5pjw+bJC6aJTW3H0dUaLRzPSzap4KaJHJJarQG/cjsY6jJ93URluZrCniX
/86GOB8VsWqBUviHurkOe5mzlqaL5fdm09GhBf6VjrGrkCxQMXvWcgYLJd96W4ZoK8cH9o3VNTMP
4gkJc/IKNNHOiVQUXjj+9fwkvDYq7G+sSybm9/doV2HQY3FSMCvNt+muiBDczcS4CtsbRYj8NSft
BcJyq/AT2/gPE2/eUDEHCHESnAj012kJ5Vm1xRcgxwh3VTjgnSqhIdVHof5H74htc4lbNZWBjiRH
XxEgoz5m4ZzP1jyI+tEuE4VntnbdlWTh4k6r7DkxicQsiuaGXbWEgvwozrUPh7vZ1HI2r40D1For
V5QHnKoGuAY4vNzEND4nIkh6vN/kicTufxI3+9/kvWpXabQxJSk/Q9VDp5gce7qpS1CoKHm7QUNK
1YQYZswgG20m1d9QBU/zxXcejNi4ahqQ3U6oeLy1hQzm25xvTTdy+V8Z9RAxmeg8RzNyjQAivraR
1jZeH8/1h4B/NZObzD3K8to92WLP0N5iukzkDOMHNUHVMswkZcyDcrteRM+1B1zyhCJCvmaJa7hT
wc8Zms441pCIWrh4OyXtlNYX2LdxWxln3R+OxYmKTf6zWQUdXyecWinf+w+55DJx0ncwGpkdZpU9
5qQKrWtTIacvwmgJeIXO96vGawkzuD4DXrRMY6oY5HItIBcxTrlL6fiDDfuSGoihOpbdD1Fj55Cj
BPWKotkofuuhSi1KqppyLTJkgYPJQaAFb/FGQTtKqw7fXHtzU2VnNpPPKDVsiQur21pws1ZzSMXV
HPMzXmMCzJ+mt+Rzdt6HEKf7QJMpMqK1vfHlZH7tVs38YBxSgq6q9TRwAYLZ/4feqNCsB/BdfJxr
/8Xaa1dSH5pxGxwpMeb2ryHrnZTPG0He2c4WMJTJux6IWPcFrH59LVAxYeL6B8rWk0ASkknfukjP
sKyqU5qDtD3lK8eBS14PqfddgHMcLy7H9w/mSiGIyY/VH09+HaD09mC4zHLU/1HcsmRVrEVOwWNd
lPoWG7kPpeGCjR5TdxLFxOjHYFMSLmrfgHklAxpxZVwUwWTYepW5A0/j38hAjJ5EuVJwnVyEmlaN
KqDwrZSlKpowl9bDlx9Wx+wDYQ0IADuMp8S1pLIKhm7r2JFJsCuqHF/UQKXCZDkerIhkmM0YGsDO
0qe0Ug5a747I2cLvCPyJZiEolVedKQWDM/b6mg+rCuWl4VhrHQSQIK4zyB7vuA52yNqUhrMBGIbp
Ccre8NbwlhTC3a+jgnX2bLJI2lmXNyMgfW/JVbgQjbvRMmzYFBq32MxEdilLQ3X+/lnV3ABDvDzY
5prFe/r/z9JFrwb7glktftdHabWfhsLdk9P3SgrsEVXCKG45MmksOz4OiKuFdaTlMXTyJJxZ+3le
NuPYzNW7I/qmG54g1RXpaOPT2XL32+pagGf21nuYYwv8NjON0QVjGmOe4MV179nFv1I36HTqNQy9
D0xnszhxe4RwAE3rCrVd4Qke/FzYT/ChUn/RyMmm9vRVhcKftJxKJBdOb98ItxPWuoEgt6gvHMfK
c3ePkQIPAmIyIqZzXKytZjgRD22aNuaMgfV0RNJae554NMaDSK9p7wJlqX9Hd3aUquLzzxeoVb6j
DOYYZoISAlPugyXKIO1SYfcLIqReV7OD/RfzuPg9wUY7eplt/0XbcPPezTU1FT51mhreSx+SVMUr
NbBO6G1QDTLFHnjWy7lPUFH7ypsXChQlMjmM0Hvh6kdjuvWTJILrtjGsd0X97miuIsJ7V7hkTJgg
2iVO5rCmtr1OvjktT4mhO7Es5fTNv+GjghlXwH2T1F+eVtENJkzRtlgCAdZTLX6tMa3Wa/fZwamo
5mO2lgCUCAVb/iY09fabNpjrw6XxPHeF0/tRUEBFDEXBUOo6IEXSN+G7xwYA/SLo2jpLzTBGcB5n
WDQaxRo6695WK+52FVzI4uSJG42Wi+RwFGvyjuiqTqORQcFH9T7Uq3pDHN9fGkV4OQtWl8RNf80M
Iv9cgB9utIRPUpt2CCG7zQbvOjtemx9BNP+IjlzpPyTUYPFPs3NxkL+MsD3EgrUZn+USTCLMksMa
7MgjMiI545sxYqgAdrjDC5ORNMDNSWeAGlw0QPRdsy3/D/J2lh0jjIYOpAZfv2ZDqYUIhWeL8eCd
JrICySUDBYGgUl8YWFPQwSDqdit+dwih6yGP53V0Bw4iW/FsTq7loTJ73NB/Or6AUYO7jEQOM/A3
KBuXe8guoFK0D4rzov3eJbMndKnMPS/dskBmzKdpBUQa6aogaNNuOdxPav/TTokMkFERQZ8gf5b6
mdm7VxHtLAJDR8WV9+dHZLVs0XgGiHgxsJcJaTQ8XBfa53RVnBVt3t7XSutaE3WBIbEr/vH8oUfj
4W4dVXjCdPYvOEgo9Ly1wn/seXEhC/+uL4mpt+dhFEfyTzfbylJzhsEflHnDMQaMo+cac7IzmzEX
2Uo+52C9uOZy6RQmzmMknT48TU8z+y3vrcvjXKzj+O4UWEw0N4zhvIoD2qbSvu5reZ/L+VuHS+VR
lb5AXbcbl7t4Ly+7YEu39daOjArGFZaR7pYnkjXFvD89oROEvoMemU0ntrwUurt53TQXF6B5Dhf6
MM907bWOXwaHsteSjiMHwTVeVLyuQZFjogspagtSkrCxWeT5c89CVTcre3Vnnjh8yCXhnn9wJU3A
3P7T28b8y3CPhIrZa4w52uieky2Rh1e3P/bBOPV4fh3EnQrrME8FZNviy14aoUoH2gyDI0DEPxpA
GhWIdV0tL8iY8O1Zg040KMtzVL4UwFsxhw46CetZRLUbuo5H/TIH7NYAj/pOumDZOGdaE2gTwHiA
DSsrgNm7bReqVu/N0pF2+higQmJCWmGe3QtLWHXxAqh0/JVYTihFHbcsXWVLtBb0el2yJYRtkA3n
dYzCfD7i4c8QSLcHiasDBMmybr/XByoZQpSth2eEuyG3QRn124inFAaE3RGA5W6m6CIZ64akqZ0G
BH/XErtbwC4txGY+RFVksCqyrR45r8cJAU9qBF6w1fbXDWMcUVz1RoErhcQuK63C+0UKxRcGxugq
BuMMV2mCaXja+2b9zINs0KikR4FiQj1mqKDxIpNGllFcMPG6ADV5yBawJXGIGVmuFZuBmzC53dJA
QeRhVDMkghopVMGfyCHgJT7cmqESsUDQguDt632aIlFKwKJuK56hHQZeFcb8TAsU+P4SbNceT8y1
fnAq6MWKkzyUMlcJ4siwSWtfmxJcxYbqgUvsAMh+gWFEMU00Q+Bzki21gOLQVYahPfjZkyG4iFsT
ItaCqhqcBNoIpRI6mblkiLw1hxnwcyxnPlDC64DlOqB8j4VmO+Ig0dK1qhQqKbvxWJQpep83fi2z
tcvb/r6bWBmo7LXjDrvtA3xHDte9xQLSbPKPt0JjYBjhbn7BWep2Txhv0V72w6D+oATeYpgEbdJX
uQtuL7VDGcUPNOIVxUditOzT6gF7vgmF46sSMWn0zD2azoe6TxPniEvkIIdmOqsrqaWqmjW3zy7r
pMwFBIgA/gp7cOxWplfbdpV2X/CC2e0pWuUcnbJmgylDawzbdGVOr2lT12q4+VnfQ+hVSh+Dtlfu
l4hsY3atM1yXfYtZ9w883ToVkf2E+Kue878bTG9KWzuYMFoyAU8buGXS6kJ88AQhFEXGgozwuMLH
PKTQSCzWPPT//AeCZvpSdBCSutPH9qBhbwGGYx/gX/oR/Usvov12FRkvt9Y7VKLWmQ9WgsulXuB0
ckkPLDJmf4a3DGE5eaqx8SflT+y9RvqFXtkUJrWC/km7ubsKoON+zDB+mVJIHgBbVEstCn85T1ur
5lOsVEMazpPAUU5RDNZzBCbl2Fl4nlVCIg2xj9667SNhjH95ivBBl+PCNShxsRH+dWd/OG6o5Xjq
nc7i6NXLTU26J5fXaVkXoALZ1jEz9+rLZx9f2yVwVorS5B7fAc04I1s6dQr4syoTj26qXG7N9U2N
289Vmxqw2hDsfXtp+PW+SXN04lwOOhFXGf7dj40/rvIR9cQN44Y0IfuTjuPeYeEqy0gF+2qP1WS5
nHNZIIP4k7vGvFl6H8oY6gjmsq/O2XcwwY9ufI6qk/m22z07jZSpFvo4Zz4gtzgjp8awbgQkRs0T
6ACFvrs/GaocdYDHZmBDOxNF+K0i+RYbYy02bcRmwDFCBSP43APo4EG4LfAqtzAg+Tz7mX5ZofQw
qaz3l/NYMuGrtQSjYGYkBTx6nac4RtNEIl9iJA2KJEUYIT+kN/dT4h4HwS50i7RwzgqeCKRuuClI
rydoBd7XtiNZGRt4IlHep0sU9ICM10KjdlWHtKJ4j3qHmc7Rradiux74o++CX/8r2HBZ/ghelkr8
okCeN46usPHfkqPRF8wpgY/EzUwShuXrrbpxBTSrWbSbRNfLxclAW+8QGy4T4X5ooTH14fb284xu
JuLT+FMF6i6OO3hUpDDHI7JVfuuspTX0FfDnWpYEAIIfqKEfJwD2LfYQmOTyYW/scChnF+K/J9B9
AXBlHFlX9K2KZsS84ATFPeRuREHYCOAw5YikxyMBf6efA9487tdof/9OR2kC9f/vv9J8rasJNmEa
QCFNLPC5nTobWULOFj20WQWweFyUdNNLQ/QEpx43vx+EqHVrWXOsSdw9PIyopJVJudsMEwVpfTJL
LgxcjEV+7gsUdfWF5CayOKzKCAeaRHgZ36VTkLAfVdWp9hQ44AR/SDl88sxPmYy282VlRQB0EVO+
MjPKN1BC57uFLCfuHSjnW1syoT8X3SmuJwCYdxtJxRPUT7bivfWrrI6KNwFoXE3zd3rXi4GHHn7/
7SVys5PlYe3Qv4fWybKsEEmAUL2REMoKqKWC0Elenckgxud1skccg+rKVP8ehJ8HQImURddCdUSQ
DKRM5LUVuouc1K/cUs18EtnU9fNhxy1eEPP6lFJpw8izo11xBmMAuYYEDTJygrIizZ4Xgb/Iqo8X
smMaKPFuz3hcFjhiZ7YF0BwQSZdpQdAtMJRyZJfp8eM/Mf53R8qcetoucDktghZ0LK+53SNN+h6A
0hPWrRXi9dVJXlSE5K736EzeBCErrfxav2f64rj12DJvVNNdzHlxhmXAVrxFvBJVf/NrWIwrIO8H
EEUdfAd6t2KITnzQpdRza2DHYsJunqD/jZuYKprdTiaCNDnuedY5LHf42eb/R/EoXIN1TKrIgEnl
GV94DRKKBgfnqUGega8gF0q9O4Eq0OBmfiSw0/EPTPQ4T7h4UWwKTnsKtTNk7pH54DImk3NRcEP3
VF386o6bLw1jpSrV3kL/BL+AlHWe3gH6zizSVHDfaUAggNLkeciMmwVhhyghcyJuGD+KCDfSoBa5
MM4wiZKy/v+Z+9N2vENErlOoNZg54X0j8Y6ytuoTMn6IHuBLpab/wgr59iJZpoh+x4tK0nyp6Y/i
T1BKkHtfsqG684LhfqZxQnI5GsfC+EoK8s8cEVn0chC4EIqBxbbaTBq+1rDNYIOqFnuFP8CrP/o6
ozMExugwdDZ4iBKV+vtldaRQG38XYeRzIAOMVkYlUcQx+ktQOPLkfTXgfy69k90bwYwILlGIhlGR
k8JXeIF2kyVqeL/pT9wQDqlE53/G/Jm8Ff6j88xAnVrM/9dRUwC+SyJYfuyyp+2eFE60pnxrmj8z
OrWtSvX2/ItYien+evQaPws0OqlCHJjyh9t8ML842qWqvZvxHALgdq/QS+wjsM1vQkXOmsJfld+8
UpgYE5tN1yY8CBt33jeO5VvslsEN5M296WlF/jtYPMYux+tO3B2h7v/DUE1gYxTf8I7lwPEOgu83
qrje7s9RmZ3BPhtCcfUc+bZ64TkKGwbUuv71NGuYhXFN7gZdRF1Emfj+dt/s3ii59fPWZqb8dnws
qLNIofMZBCyKuTRpC25J8uPz/WCNhaA4x156bagvDkV2TeSwvo474GX7+cSizlZZVaiT782k4diT
5ZC0GZ2nZ84JsLAJZNZoG6aHhxQONFOyFVeueENK4G8VyBQGmigJVlEaSrBhZa6DK7NF9IYUNJEu
5S5qIwlNLDVzhui0Lj1N+Y1VlPSqPoyIAanMr6agsx47wlWB56/QFZVwWrH9EtZrplVkHifjx9ms
SgRVmMdROYsQ0MBldDJsYnkjoh4IqjohvMFVzmVutQWMhyX+5i0vXM4o0VWZHDOYvZJAuH1jNDs2
IbwaPtn5xWyrAx3Sd8gdiIKNOjjsHrCojM4gaUV0jVt99WZKZlDqSuWFumbFBMfkLgnyQeCj/bmI
F6GMMbqX2Ing5uN49112plXRBPwkXgQebpIg0Waq0BshtM3m6bw2vql5cJ0cesUGti8F9bY/wGfv
SdVY9KEoWe364Sern+k3CSqi+ukq1D5+laxU8BwM9SZW7jupcjDjKsZi9/4sESqYw71+qBBQ8/5P
HVf9XUCKrYXdk1Rg7Bkqhr0REelFr0J55IXO3A4g+qkDwS0M973bd7RQ18ZQpWBniTH2sKVorHSz
V2gwIWK1Twxh/cz2pvniR0sx1wmhsHE/9KvtZ5fxfoYT0Bp6ilJr4/LTDWLdfdctptby5g32tK5g
mgYri6FFwpvpHSkyoi8NOnzkJTtLI82ta+E99/eQOvlUeqE3Bw0clU8YHy3s8tbPlylE+tX2pvTo
bI32P9KatDmNQ5hNlhzM96zXxf5tzg+fkxeD0mEKnZXLCj1CoufEKttRuvdRPeGcMMbvj91Os7md
HlOGoMNNhSzDnZS7hrLko6APsYqIfj1dFuUgN7m1+hnudAfX6Qyl54OWXMuUlh36ixi6hWTTk0un
TsgohHtmx8NyIfij6zjyeX1mjZkXj1oz6UGLGv3i5+VvtPBD1bj4KGaDCQaXvQgAJJwynemvCmGx
zCCq+UdXmNN01Kr8WNXpnHjyoNE61LX98pdVODFcaZ87N2zRLCmmVvWz1SQNGPu36B/9KQiBI1w3
6MaK9mVs52GjjAKMRjVHpmLPXPS7BRH4VIC8E029TWgwRpYPn6plT21o2mnRC+8e0unOqjbddrSW
ergUTbAe70ihOr/GqCEq3XaSse+RcBiqkorvmD4LfPoWMO2tuNoyvJOSnSTwaufG/WE5DVHQ1pxi
h51WlLx+G4nOQrkO5gv3M+xsMC1ThrmRteFMIo06Cc1Gt4Sla6jlTkcHNxadu0MRjr4AFz8mJ2Gj
e9UGSsD7aSeJ6UQsFIaauFJ+wOipOGwdybCDj1xh/B4w9RNbkb5i01f6VeEZxRuFdNTFoj+NkGHF
JN8/TBNfcwHNjku5/3FJJW8FXVDitn3/HjTaGXmLGUd6D/8eNQ/GHCz5st9P2etCcaHOJ+1SVOlm
xovnQqzmUQuhXjsjwsAqt9ffKRikRFWpzcYgNWxJgPVIMgJRbxb7NX94f9ld5vkVZ1OQmLANB0Fe
VB2ar4oXAZ/Y/+lMU+cSF06c29o9Hi1lx6dEDPnj0Uy0737ajluB+vXaiD0S1pNPGfgGhm/D5mbL
hMZYPFyXSbaYgDPSDDJyn4UctWxW3MCMetCj9HdzduoBHF9q4r6UfUjuLzcFgeKubNzlFmw1emFb
m0Y3lfdnYNm1IJ96NfznD8MSMCMNjSjnO9+H7FlEoKcVG6VKBzPZPTYfqc0dZzwN6yeUrQ86Iuck
UasikVXrZh/6Q1uU/X3kL6r2Qu4ygAwc8bD9iGIpq78lB4PsmAc1+rKkd89kjnyiJl2rT6C60DLc
HwHD0Fq8Rt/P/P+j3BWp+ttynPzAEhiaZ+7rCm3ZdXqkrx/SGX0sfaI7ueogkQ8zopt6RnTxVXNo
Z9MtyUUhk+RQyK7HeSMWK2Dp3ppbrlK7e/DopvnT8haMLtuySFV93STWEikeoJc4t282Vcbq1KaU
cyYBB/4de8UZn4FKe+eukTQ4c78s92aEYPqUst3jAbmPWB+xkuP5MClAs6ce48o/cOJy1zTTsZJX
8hw0yItD602Cl2E9ak6mYAseRitT1dGFnS0R87CAIVOiQ7nTrjmRao5/ova0dxe261/t6ocmqq2x
GrBSTx3kVoCrAHBU4HV1peupRK3QhTb2QHetsFJ7vOXXUUfwC7+ZEAmfr0p194yWX66VcZPnjLG9
zoLiAu99w/9QlpkSVd+e7N6kZF7Y3ZVgYjhKlHSeklFziZ3vGSU+rQUpDGAonhJkY+svvAetweA+
quv6bNndJHbFeWBGGsywAIdNMxFx3iEsl9oBOcYIKKqBcN+smrbFAbI4IG1xcplmr7Q2FzLGD4R+
3ZIjqP9qYqTLqu+kHuhz0eIPt9QFq27B+ZraVprxGumzaw8zGL+/LnWJ+C3iFtwFefZz9s9ogR/q
IwSAFcooLLZLooJI57G0vJLY5rvSlVF0Pncy55cLckzDATtT8Y7l+K5RIQRXnI+n4ibDTmlMc3BR
vq+SVp4/TX+g7nlaEglI1kW/L2QLFgs03FSLBHaAmRUYJMnoMydj17oJGirVXXaSeSE5LZ8xQKHi
NCx1wxQhj3aIK6DOm3WuKW+S5wrz3uGN0fwYbtwzjQffJdIZdBJ8bqNfn14/EPtK9zpmASthW+vd
rHoDoS2fsShHWAz+Q70acF7FHqv38/xbX86hlaYwJh3i8KZa0vEpBZFQdYvEEEu5b5ZjusW/sXeN
vokEfPncOu2WHbqwUHgb2bCZWzFItrbmSdYIVyt59T/3BEh0LM+n4QE3OGR10rIXTGgarErzWRnj
0rTr1Ym3tND6QOOk5VcD1Gl9JSzIVzS47Q0W8ImIJvx4q1uLJQuqVgB02Gv4Z0pPq2JcNUpw1c3K
MdUKqcu+Wd0ztsy/DPxYq553Decf7Pp3UYLYD5kChIcd3xBtrQVLvpXVguVIZv4FYSgnkPMLHKIg
Or72WCy7/BplKoZyhoD/X1nZc+eVj9UMq3CUtjJ9SyQZcz4RrOmaV7bolHkGOrYgwuPgOWPgiwUt
kOuJIEOWVAu67Au1GJBHoEMnuMlXITX/2K6eWXeWGEB4JpLeyvQMeVMcPZdlWLqkaQLHp/R3bS6V
bPrdIxoiU/5wW/0TOYJ8dUwYWsPPZvssJqgUG9T1fwSks17I8WixhyTsUhTH4ks5HNUkSu01Gn/3
73o20gmZCSJZ4dBVkHk6WE54RkvPQjWGQ3JBiU7F/bVhXGvu687BeRquRhE58FeRZUIAl6UM/FLm
kR/ZQ+opgVtYX4CiZmXDjHf6NzTfvPlS+aHdbsaDap+NzcEn8ZxofDQqIZcbur6v49DD3AWR1zkN
8FFDzBzo4O/SU+R3HIOPIj1Mey1A7UYNeOtoRVOcf1fxzDZjXOfNFdx+a1I+7Jzva1om2064ADuV
n6/7oymg3Mi3IzzqWTnH8RI/GmT6jYpMpHD1BPoqsGJji2wg3QLEERqIdMcqhBe/KfTXu7ySoJFz
o6NMr22WG+YMxbdLYgWcelBSVD8jhNj2WJKdJdQa9fCE3l0VcF2MeQGtF4hkpSbaauO2hAjeUb9F
ZHtB4BGuejsAd1XwknuMstflV3ttNMaskjJGftHapRObiWtIF22yoW2COpIPOSMRekV9XqZe18Ko
ltLYFMAQt7aYp67dHX35sBNr9Jl9FPt3ninZI4COgAzuWFezEmBTCclCfLuX4sCng3m3JC2OMKKa
UUzDYOfnGGIXeFOb0XGw9BAIZqMdaLD/3MUV1YB7M95deJ7gotwyESeghcD4bcjhQPCgdK4wq+Iw
od9aMYtks6QJQuuV8+yaYYTktxls9/C24Xnlk3FADmqdiMF6M7k34IOnYJWgIyWB0hkL9IdMi1VK
2iZeUhueQCzU1zPPi5H9PKwxaHEkyuZQuRPOJN+Y2oVH+0Erqz5SKvVvEBpRMnTqoG6u4/m/Wd7j
J1k4Vl0Tz4Ci8f650MnHDZ7AmIp1+QchGvsvcZNqnQLnRzBraVFhaRo6KxdqotH+PQkigp/6XHIG
aROpwEPJqO3ORnHro5RSk9ln9GQGKGqkq3O63myjbCwWV3+BjkPDAMTpvSoshUOgDOzIAAqwp6eb
+57qwlV7Shslco4ZgAL5c1wGVyOAbC/DJtsHB2T7BgForB4lnkt9W+ih9rfauMWP6ploYGPyM9TT
lQJE+9RsBZS9CP10Xxt/i8v4xoYKtSo+erriJCcUyeQlQujmILt5OiXs5uq+L12MsOQEMV/+NcsN
BCgKeK0+3xTKZhMWQRoOkAwQH3/U3GyhIzg6EXd4seOlyg/8NyiXDKUJxhpNIM6awXA6CLQEwjlG
NntaZnh8EyD1Cx72A+/yLKHT9wBW6c2tHa1BXz9zLK+Hq/XPczd+KWubvV1ZmLW9YeP9ZsVI9W+l
8aLgLj8Ogx62gS3QRh+VSERIiEKXD4ZIeBVZxvS5bPCgQYXCEr6YIprPuG7BOWlXOQ1FM0NhgDVq
IiDDPwcLgkh7HxB3oGEQ7o9yDCg2Ys+13cTpFfcV2V/tAkxF9aM6FfKlZewpVzr+3JUYAv7Jvhau
HNjblIWPDdmqqI8zqma+krtMA5U8pYunwUAN5HgKMc+6RytYHmW06hklz17Hgrv8eB6LOJOZtFxm
7EqWwLyEI6vdGT6t8BEdEXNuN19zq1CGpB6u9vXlnj0MbsaLlLiu2HdKx4HhsN9RFJX/1m012YFX
6LLGsaFkts7ty2d8elUkA4rJGHSroSv96pd5BqljUSl3rpPg+KQF2mZC8TD/bQ63ZoDp35pa8+rx
oFS34uhyPKMr+oB6xcGSI0IJI0ZVroecxq/CSg7Ik4IFNHtxSDwsdRgmK1Bwc6R59F2L1DpHcBTv
lYAEYkPeQqCZMt8vwwgi5W2oYgla4DKhFPthYIWVZd1X3sYPIrbkPdB/1sNrA+WkV1u9TgWJQd0Z
jYZLePyAdmJdlAR2RmMy6tmNGkRb5VI6cMyc8kOMRLu/tfttWuqK1LG5jHd4ns29kg9qun3SXuDW
ASzPdlplyrG54ID2ohwWReZOSm6fUEZDdryioKU7BQ79mzN3Z1TcJyH/SyoD8nJ25L8VlSLyh5qN
GgV1D6D7L1YB9hVGumKyBKXPNdksbDKwjfG7IS3tC/LteOZlf5lCf2O2KRwHvPUoIUkRLZ1Wbi0B
FlmYu8Tm229uqF+HA3ZQRZq+RUUoq2WgxBLvSImNcoGoEU9CRRhbxBnRltjFWiw0xjQcOQAuLhQG
KwHu0FnNvtbSAqIPsjtGt58jVwt+FuitSqHizRB9KF87AbqbLQRdm1QUzi0w/a18ED+P30/BUXKf
4AIIYGfREUcMOjLy1guzbySQot3OGvqomA3KEZDZZ9nH0jbPkmamk4tcXu35SkDBmoca5horqfq6
i/M6kV1nzm63CRB6etIyRtcEnl0IVWtXZ93eAdDDL1lkPN0LCSC4ic5SHx3RyZ40jizkuy1iZyjL
n67XLPIA72pBQMXdakGYYndR8ws03miy8xn3ZpLy46nO6goEghrHIFs1x1tPgv48JaY4CaJJK9MS
KNNxd9ZYAXM0nvXq4Qwt1HhbCZNnxIFvVo6f9EojLbo3skxxNg4Nnc8O7oMipJH23MILy1twrLuO
yhwxcUYuKhyn4WJmuVSC+ER6Jo1bWVC9iNnx+l5kHuEjFvs3z3ZRX2FUDSxNAl7pKv2CMUmmg9BC
hx/n6/5zJReQ2XcG7D7zuY2BbQwhYW2zAFUUWOaUYILVJ3cIsFG7MiLNTn/arOo/Xsm0f1SKi796
nffCsQS+aFsnAu/tMHRyHtNcxrsPrNJPEWjybFnHDcRNrsK/XILYY3MtGykx3ssGamRgi34MfOv/
hHGrxoakVrHuCuk/LwN6aIsDxr+kUWO7iSFpUSevp5kNbmq6Na/GTfpFo/A21LgQo/Qvle/vFgKL
Z2IOIDxXl94rH1SwiIAkf8l0/aW1rhxIYbbrB3/vqkD0Hs809LKd/kIpxtOufPaPRFAfl14shcOu
R5PrTrlJXYkI3PSDwH96VMv/Ns/id1VGJUwkAqgQcwybxyA0T0H7SyVwWXvYk3kibt7MgQ+bpSaO
1Ul0ICYO5VPHo1L8H6Ld85TpMC1elGbBcQ7MiTt6RFsl/guKoqk2bWi8aAyXyEgSotKrW9qahymk
7Cqq0fHeyDcRkUKFHFR/1lVe0dPgKycfe4rLEZE/wDEnn9oOM6643Woa91zD3MCKhGfuvWL+tk4j
BCLhTuwSovXjGYfRUjJARPuM3SBC/Cxg6pZXQP45JsKy8P6sggo6/5i/Vrdu0b+JR3RlNa+KQJRS
1q2oko4Naieoqt0C7cjG2qt1Xw4MCgYkqwJ5ss1zP/IYDDTxX54hdrzYqLhQHwHBn9q7e03SkZgd
3fnq9nfx7SYVYWJpg8vNxtpuRRLo4nHmb8cxakvo8kjwamGOL+kP9LHHJzBnR4xw/PZ/vWLWreK9
RsagJuvvXU1yTq4WwPxSxe24Q+HU/WiL8omQAx55tZIh4L0WiXXM4JgCZBdzewvAW9o9ZYSG+0I5
RE4JM+qn5fjqD7QHSHoXB/n5sSLgTMMHaxoS9+ZkwiLZt17nZbJlwa1ejtsOKiAebTKa6IhnoCXS
FLqJgawiHw60uA21I9TP7i7vD78MPoTZ+XVhwrRUK1GPmfWG+HlXdIwxXj4g82lhgoqVsj3lPECH
UgcR04uFWJQDMSL02NcejbkE+wD7ZwSIzgLFW3rfzty1S/quMlkYt9S7DOMkm+xlW8v4gwXaRw34
1ACphfobYf11UilGLKChxUwyluO/Z/+l/40Jgi+2EuHfjyUvIpl4skfL5k7GtjUFx/cB82vZeMk+
N8x9Dkl89pf0yCbRaOnudktzcYGzIFAbhrb8V+xYPm+vFy2Yqi5ZH4rpOocvfYM8nRoNHJM5FbCV
Fw0bh6vKI3135nCCIAZY2QVf2oni76vM/A/PF1QC7JPWTnxovJuZiB30z0cF9R0gY/y3xVcbsDqR
nxOFFOMyWNdld9/bxjw3g9FxRs8d4baqKt+f+dvfR1OeQNdmwSO7x9tSrndxE6DfImdj7xQft4yK
2thCAIBaPdsGyMSWIxByvRwMvkUzCjHdf51J0kWf1KnXplRHsC60FifaFZFUiQ2w20Ymc8IyWcIl
ggH6FOmsPqKBOvVxO+8Na/LNQ/oXSGmxb8KPl3CYo2HYcflNaadL2OR5MrBI8ZUilNJhjVufi3MY
J08gDUmLvp3BQ3JdOKSJrIGA+lui+Aln7XBnguquoTOJzsBYicEv1V9QP5mO3MPni29U5/JKZVhf
g1aXjsmtyybfJsrwpsXv/Gq29XPmtDSTCQO7h2MBirRSuxCP6bBObQAUgTL+VL+NkZerDzz6LwmS
AM/LOFt4TH4/4VA6TlhSX97rRlwneAAnO/LizkOnJ9Kj06WxFPc1UMYSAYfCmm1KwgcFSr9ypKO5
U3bW0lH7kHNd4+BayxmCfBxXu2V8VXnJwV+HjEUXVdqI7G8LBUUBgH6GsB9l1+vULyyKfJuxbzKA
GoaEaJIJblPp6bJ+sEa/MdPt12d/2aguB8F04avzRvz1LhDLkr5I0R1n6IYHkvHz2YhsQhZV6HGZ
f9P9d6D0Xe2GJqdgWa/V1whhQdgnoKmcmMj7wwkP4MMnZ7xmTpxfWIVCgyreXyC2R2EuV1jVhbpS
rYa+mBWIC192FyIDWZfRoAnnu4yqQavn0C75pKmYrg+60DudOVJhEFXmYhUYQ8xG/d8IQHDCaQ+H
LgA8MNFI5WBRW/vQVtxw1dxmRn/69UNd4E0szwSTdXBUOhIfpj2CQHQ7F32q6MowNMeWPbcbmpqA
UWuGocqvRpDokxKdRbtSClSQ6zFjWhGRn3z555wgfOp3/9ij6OfNVW4VYFDabjkrUQ4mlP8ZGQb/
CSw8dB8dzHbrWAL6gSYoea+6R2mWjv7/z1q5cTAg+MAU7P5vNGl8oBYmE/TjlAXyt7AK6zOXD3Ay
gVVm66qAIuQ292zUwWxEa+7vihnCFq65LMH4ILpTq8CeYK7Z2XI8sgtYY2eU4uvTTP/tmahl5OAM
t46IBFCRaWULpGfNZOaMpiiZBjMj5sV+qJTL6/8diQtyfzRTCuqi6/MGb3DauyfYYhWhk75yIaGd
g6K6jkaNvxDKl2wuA5Xd7i3jbUF9KHWc7RiiL5lyq/bbtyasyvTh6edhr7hxlB1XQIasSYuJ/Aji
AuAT4bnceceYrHfSgxruyov1aL0QYb7Te6DqtP83TABRnH19lKvsba1pCdZhsRANE6wo8ce8Hg6W
7VgKjzNi/uWjpZi2nxMwKH74F3aVZFBKVERBuz+2+OkuER1cbJfUA2fSz+/xtN60Pf9ONvZ+sHMf
yzSLyZymOnAFJmkeWYjpg04E4Ma7q8ebpWDslYnAXp5QdRjw9yaIWC3B4ZyuyRAFI7ZdvyYKjK2Q
vkMapXOc6R8ZySVYCGNaIspUUNO+FQQDETTiMIr1QgmaynhCCKev9oDo7l6OQ2DTDljQi2s50obI
b/5VlMzyuOhmzqJ/khKAv8pNlnPiNQUpHxUf4pNlHOBNkh7QOKXc1YrCJe2UC1K5hXzR4rtKUf0R
UPLT1sWcBc9W53SUJiqo7Zi3Jf0WNPdGMKjN2X1c8YhwgB5U4dfDmWy4eu/eKgcl6LT9ALVeYV4I
Sk/t34M+oJ+nSRefEFjGcoJ7hJp1Sgw7BvEmElVO6KsZOprKuzdlgtmiIkTom1UQhKQ2ofLbMDmt
lOZZt1KJMe/d3nayZPW8TovoVtGDcNWOp7vUuV4zBcnCGLQm4sjpehXPmeMacsiZdr9pUTjxkX8T
FxsPWmbTEuhDG/X4pF+ImbpMWgt5BOZrD8gYZDzjeNeJwkiYcQF5Av3Z1y893eMAS4z5+YDJIJG3
4uehbFF2nFF18DrB9r1cyqYsIIBQzFDxSxUVdPe61kdSswqrlLzMUjh+Z8zy9iqYua2gfMZl1A2C
wG7++1gw6V4YhoNAcXn+9fWLq2Y8DHfTr4aQ3Ry39ENIHRtRo2leO3fVOLiEK1sGLlbIiDImqn9a
Ook7edYDDHChjBVea/xuHySf8oHJeLO+MO3B+6oCBxuLalxtUIU4yFNUo5+Xcx7pS02f4kcPgjE8
6s2mFtYoK3DfsKKntwnAIGv0SwcQSytL+aoOreQnxj1VDqP4e67Qjd633jr//swZZ7ZBmZOCpmqI
FXWyeIY3L0uBXqZTHatehyWRfIhIRgX/FTOKBb9Eq0FYCNgFyD2NMycDZ9hAHp6vwnjzyxQwU2VP
vYeISxjr6Npmb3FTj06PNkBxvcW0FWJeXC0vAr50VxzZmHs3NdQkxf5jHDrCu7Hgv3JBRBzg7B0f
wqidHzPRa/B6JaOkv6xMXPVgX1r1m90v0rusM/lUjeEOlTib4qElJnZIe8e+8NJoapJVOJMMTSKB
kAJIR66qLLtmErkLFQLjC4xW/ZoPl90XGL2u7l+RGCmYrhEH64rg5FBnA2lovYxrcvsHw4EAca5T
7f3qiQrXwmQIIEM+tzQ4rw/Lp2bDyU2WTDunWyJaoGs22p6Lf5OBZfLepiaXYyeyv5mAo+FRsHOC
DeSqRJi/eF+OnhYEPJhtM4xbIy2duhijR+CUNW2P7oA2kx2e+c6D+Jl2RrotDwuZbJcjNL5BE25w
9VDlGMKerGnWtsRIjGkWBsdIyeeQB7ds53995OCPkglPyQQ21Fymop3IQPOncys55InhCeEkj7ll
R8jJCTVyQ8TsublFIb4nDMPCe/alOD/pIleidUMURCA/RBfxGG4TMa9wqP2m8a3CutqM1LLIteWU
JHelgdHlZ4nUnyq4NxSPkP4BBxpa5wTc12pknkKZXn3S2JtE0/5YHsP0TTHsAhChQwcBy/TTMj47
M/UOVQ8VV9HKg6VvIVLQVqoLQhKpUpjOTA0Gh29ZE+lSYyixZqMAYAEOGM+LQ0MM+9J6gs0FiYrE
ed0ZW8UKyJHggH1Mg+tbp7gfZdCpqKqp88/Ayq7o5hFUd3pkeGdkDt4Ft1ekk9ur7Pcp5H5R4Z4j
0aAKuRhHCWFnviS6Hlc0OZiJmD7u61h4cQhm71J9Oyw8WccEQvRFf8nPxRkLznLxtMI3UTD+p+s6
2o1IS2DsnX0bff4Q1eWs+tO46I86mp6kNjj2zij6UtvSF9rmEmJ0qSmlgpDgChhUZXYd8xFEaVyc
GjismLRole04+SDPKIYE670XnhUqSIjeMKabfCgzGN34m78HhY1gtjMl7TSPVWGldyBOfyQ7zlxS
p+g/Rgc5ARWCkgdv18/8qH4RrmCJD4lFZ/O8cZY+mfHc7c0Wr0edd0hCAxKAEPgUMPYlEb0teDPz
4Cmq0f8AdKvGW8GVjMSZucnBLkiMtX/sbdyMJhBoTKFDVa4VMRk2GuKnjBJSon0R9FOxPEzhQh6u
zgRvZRAPJS9XVbByQLUGaX693mx8OtjmX+u6FlnYNTYniMtSxTFrV8UZvmT3Wba3tSKRk8gDQTC8
5KUqJbgdM95vjA+Bd9PpGya3WuVTlY0704oVEH6ZOH+BwMWCcK4+KuVGeB3n/0LCDHYcNo/UdA8p
CTEdMOR7N3WCcynjPie5SjlW6RleiawB71G/YTu0AauBeKkQHl9a6WXdlCsCWXsAnzx3pNbFe2oN
OzQV7TNrPQyJRXX+JWL4uFpbNksPSRBvIFhrnjEHrEabJ2py9bmqNHobsrZkwyGXBG9LE+eoImJ7
Db6SdDV6Ii8ePkTdyKfo+mKHAg0FUeqFByt/sPH76FiwwKJzzkJlJg6eHOnRxFKLQTU2N+U1AVbH
HuejKc0dT7wCTDeJt9LEcPyxzGcSl3sRi/s/mu1Ofmv2qspUUAWga719G7XUG1mwQIzpTgebXFEZ
5lJ2hnJ28APRmgCxqRKid5BQCnhDWANnfRWoJge++WsMIpJDA1FqmAuVWB5E3xtTn2o+oAFkIS9p
Bp/nU0HfsklHP7mejW7XA+RTOhCt2idtUtm+3N8eG2Zk9wJ7wuAZtka/WTLDIE+WxmvFdWCk6IL2
iZwDzhODtunULzieU23LhbS2aXtef1gphuujOlRyvUKjM6M6/7QrAy0m7SgFo0ldQdxIkz7dCbRS
jGyAhyI8J4svOy+i2szKlCv3kLbxSRAOTmu3CoxhwhyMoFnMQkr8iM9F9JMFU6Wy7dhhIFSh7Tpq
g3A9P1vFk3gFVF1Z7hEevfzj0b4HjldNCoCXtebI7O16m5F4VP9u2D2VNf1crhXonRZngOibOdOb
EWVoRaDG7n/d0wNEuxfsuwOSopWrEogh1SEbKpWjKXjkeVu6wmbcjGNC/mnimyooR5fHJ2NmreTM
K0y2R8JRFL5NF9FULmf4eIVolJnHoq3J681FSNtTWNN7IatClYDSMbvsfU0kLCQBu47ULtydn2dM
oGjUCd68zIcJeRjGWFplfi6G+Mk431c0a7lqtenizv1+Eiuv5cbprSllsNYKpquO5AA4t/uMo4sH
tvd+RL8556yxLzQh1JEwZISQm+1IHjKVVQ1jOD+81KvnUR5me5G7pliuNlzW0fhsEj8asPineleb
wXPGHfqvd34UyX8SocWnIFzEY8EKzm+mDlEPvkfX8Fd/3M312d0BCyZ8989bPI/xQx53eejiZ+aR
EDgwTb6YLOLCCXy2kL4be5n/YoeqwSzMuSrS2LWHBgwIhhLFEr6A574nEjgWQ1ztsB39GM2nq2mW
/6sfDjHhmvCFHu4IQzWxzGFKnsFFLaV1U8kKNquB0WAQkxDiwrPVAt5x8Q6H8NrVdecJAY6ITZgt
daGKDuc2GGmsGZGhYTE5nObeCHIVM25n+qqHc0jf6T1Oq6TEuV3v22FcsdfmNQk6BPrf4amPkWXs
yUVKKOlQsm6J0maIA+xC1AnbdJ09nwNxbBHy5jJng6LnPdLyu9NSp2x+HDjT2vA2+4m0HY98gpOL
AGfq7qTD0CYHrmMTYL2uiwiD5I+BONAhMhGrq4Ou/eUfAC2LvC5GQBbpOPzNB/DK1Ii5p1eZyCGD
EQyaOidaKWAX7AZo9b9eIZx9UNRy64pQcJElVJxE8DlDJmw8DFsfUsUfmGKoC7vr88619YKVpt3E
/FDcRTz3esps2E5MkJfJm+2D+sOACAw6O7bcGIDDrrp16GuyLIBR1dJgElipdeZSUzJVOszYdPpy
4SmawESGslQN25XB3Kk1kp4G4sT/KyhLlOyXH/8NX/feYXQMT3VmIB7aznzsloAseOnvDCsbYoWx
U6U3lYRuezr9I6GGRm6co+Kh6naDvyfAPwxcRtwItX8+N8iKljEXfN2CjTpJ2z+lrlMgc+kSwd2n
wYl/bCxUjBE+hDdfotRVB8vJhD0zB/2/0RctaMithGW6eXKC9mGrxIxql38KASSbTEgxrfmtN0cU
3Ejui5hzrSTlCJ0qnybnBkJB1OHZJJKKKUvN9j4oSfBpSBlj9SVm/chRsrjWuWIZZzFiZcYKeaVx
b3DjRLlIED/dvSUgwwLHAmTbdR+Tflz6oj5fZUlv6taiK08tAUq1ZnsSMzw7VQbzXVfVNV3YwUzI
a1o4amwoLbMGIjJxq7iHFd6tpXuj2oO0u0VsrDFXyRXedpsP5aWSxYF8zxqAbJenajOgjC3yd4dA
dYKMeBbTm3njQKPqnQP3a7/55fZ5wtSQCD5mIQn/QUBVM7Qg6nzKsLI+FcqyTGcOtdUB/3DhLuEO
AFHwqDIFKQBWfUUPyJx55xf2pgoLsdOIiiIPIYmk+UuqepaRVZ5XZF+qXpIkZ/WwKvNGHV+xuulP
yCRj/D5KtzjANM4H8wuwFeVely5VA+Is2f5sL/yiqAJ0wjlAju7NUnAuww1CW2ypco2B2ndNwoyP
Y8EZXba3i1Ls/EkXsrOtd70sUozyDBALC04UoNu5uEMJs/15GbbV01uuNZcCDdIoGbhU5DS3yWYT
ZNlXeRebE7CUi0R21R6RdFyIHk9WXe8XwFcplpGfIutXykQLZ1iaZwtQfx8MfA7j2IG6UlttDsUd
+N8TY6ruQOGqWLOnEJ/6bwL6Lq5GT8SB0U6kyM7I/EOZkxEmYFwU1GxhXo4yZruy8/jF8OnP0WAE
4g42UMju7kL58BCX8b/hvXkU5VYUorsXujCePzLc7JXhAJDWC7a0AEDkbJd3NE4sbRCB/vJYy5Es
/9sjMvdU5Juv2zREy1fDx6xnkQ0bhKn0m3Rsdcl3z9sFc6HIofc8dYyc0iT80NGx1khxc5rylHDM
mVCZHg9TJFBA/mdX1XXJZIDw/rZJTKuzgcOn3ybfibBA8Q0D9TN8WhfncXiEOT48edxT61x8c70V
kcifPi0e5UY1rcvKETm8HzZ9jkv0dW+Jpisel3oqjk2jzLl6lI3Qujvyitx+oWG+ruwMSbakwW2m
vj9v2A5IbXMLa+XdNzSR8qAUX1ZFLEvFLAkUtW/ZiPTMeKXY/v5bWIeuBRYCPscOHhVEdvSU+cKL
Knn8T06Dxkpv3iAPyHtLaJ1p9XkuvqSlNKFjF9IcMZldaymGx2253Iv41v1IwQtWHJChuJqXRM+K
5V4DIn71SfA9LmQeUdF3TtBbW5FwmEVE8yUUltbdqIP+OdEobAJhFTcbmop2sE0bnrGV76itAsyV
3GKrxpfKhmPklByXjnw9V7fsTNRwCUkrWvNZYbWuBDBxirB9i5SapSG9cq/iMz5eY3i5eLjiUJR3
Gd1cJw4lOM4St/5uIXbdyfVQyRFSSYatUoWpoTwTLkSGWDl2jmJEpVNE1+/Cu5fOsH4Qsj9O2Rh8
Nbihjn1QeQMZmnkoE+2kJVLIZRA7eIMbbJp+JSB4jBgBvrh2jK0XrQJHa4fABYNIHJBAQm1g9N8j
ya6nGPwk6RYmkY23LXDiEOyQyeLI2q8JqUbK8GUO0sTw48xWDGHzhkT9aRKxqBzAQnAjkiag9SXO
yuO4k0gHMLxUSFh/nVcNIhlUnQmW95xzP/s2owwjTJ368ciwUJUG9RHFQGfZfQnPMByS4SDXm7kP
iZQHFgK0Qw18zs3VzaU9dKWPMMTvti6vd8Hx1Rl9XqdZPTMhjXHpfc4QSemGhX6qeTrtjTOuNcZG
jRF9NPFCKn27rdQApulVervvmh4p/96VfPn7Sl4SsMKdcKsXkNPlskTueDselUu3YnqKDQUqVFQV
QwPIkABZDJxbfewEaYTSaYyUx5kAKrE2pzQhB2P7ctd2/kuelDheELpalrMH64cKMmNNKd/T0V0x
+In/TONS/RxertfRZoou8DZyuCEAXRelZEzBAMu+QE99DqT7em2dqoPI+RJgpUWzJM5PMA7J+4sG
MdFW448vAJE2wW51wahDSJDK2dyL/4p+xAMqyvnF4IZq3SiLAvdWAiSlG+W84Jy4dzzbjB94BCn0
lCc2WrSzQugQ8W+pwNBfoIn8g07+kYjJlNmy90x+XFMfLn0iw91/QWxSj9tCmsRWJ3g0Xyh+iJ4p
Ls4PV7TxNu45s9sP5/pWcGT0gl3fLqNRsCDddjcnsJStcayEiBy17zPAQrwt7dHTFUuil5+GddV+
5mj8YoBXr4Mtta9BhsSyvFihGecqHAHo1vgG0ayvV/bEJkzMKGg1d9jQr2wKQqqvmPr6a+KTHcog
BvIBvgzmkU9gPR++J3msL2OMsKgixt+gnyn5l8obcKPn7cCzqUdIg3vYQHpe/w7Pt4EAjJuqmr8u
gLkuB0oebGdCGAVdtywvFhtfX++mkc916h4dHxnQd2/62fghGaRZv2A8lDZHqlQMMNplrxoEwqiq
yU945iPHBxE27b5p6P0oPDdF7a1BkUsF0/XfHSNQXTgubCNL8rrDz0WEJfT2IxFTPbU+50owrtyS
4vq9HWGKmzUdvgT9lYjRTsmDgFkSnic1FB37HHnJkUTr4KYgIz/6mWwaSfAneaEo9ZqhoRaPDVkz
wmxnXdGkYqO8vmRps9PSt7/mOnIQpcMrN7IOeRdP9sfIRe32BHxdC20NNHERWeus2KFYmoPEs5Ej
MsBj4K/D9xwFMRzCOphyhzAGREh00sXWxO+/a+khUI6D0aS+kRRtg2GKMdFInAywOyDMBfsluWoB
wHDoSV/3zolrDnWq1BVYcme7FDetFVS4be0o9YeVw/BA8k65v+0fjJJZkWFvvwHcESSyUI/Gzaqh
bP9800/U7J4NWTprgM4vlTDOB5vW2AJptnY2kSJl4XtReOL2W6KqebSqWtzsDLrHlqAaZC48uIFo
z1LSRRSTicMno5OVL0KQjsxuZNvJylXVejUFixlu980noyksuh+TFTbdrQe1tiAcneo4BKLKrXcI
K4GVVDy8PiggzOafJfypwSynUQ1IRRkGxmZ06P8zFMDtQ1E0qd1gdilkJH1Ea+KhHfJHSnzkocmj
EV55eDNvR3Nr/XnL7tqLfrIh02ARVgkurMhgFCz+Uuv3AGp0eo9N9dQmtm9XlzQB+lxTQyLm7LXv
LVa3satCb6cZaOGrD3Bv5a+vhjk/MliP17m23pavyTu3s6V7/2KOzNfmBy38+Gft5rvBcJAINZCM
jLI4KrooqtwquBNZtNXMDT4/m3FnyN10m+p5nT6q3YXTUvHM/b8dV8OUd6SHML5gs3Zhq0yO0/+n
9SaPFXUReyDjutKkEyOtLTQHxY+gCFc0fE6KWz/pkBveCKcTOzEP3+bC4gKKK8APJKayzgent08C
3X6sJFh4y90Fo0+8BmEBo38wE0EFafmzWEAiKqNdgFetwCBSBF2bpglkJ79md/5v+wPyIDr0LugO
Sd1+SUasp3vEGTAD20hWi2GuZjtLLod16sZd6ktz7LMYSgt+aoCReG9oq4g1y8KW3KmIU6r105rO
RrCkJJ7rPWdS3Jx0mLEl1kkY0UgvnVyJA4HVdvp2y9n2w75lTPY67O/PeTa+rynlUTb6PBHZ/zpj
QXujDqne7AhtAv6fOoGM9Dwp4MBVeafRJ3vxWsUg9MlgmjxIZx0AJQx4Y3IHF7R5Xwuxrd+lkxJH
GA75fLk++fcpxZOdtskOQGyFIHXR5niLYYhYiKNfwCPhUHqHHWJ069mmhOmBFudy44MWznkWPjTb
qQ4ReoNWAdS5WHneOl7xJewS0G3KW8wkruUv3F3BOzIOPk6SNSIiNh6BGzAEHsJjiRLuzPHxSCoL
Dd9KlXtgxzTnkZlEKy/6/FhTN9xblZiPOnBzxP3w+JchWow0pQArrXGNon39nwMAJBZPD6zeWQrr
5SdsmO+HaGcGKm2d6H4U0otV/I0F2Nn/jj5mYNQZq7pICttIsyp8gDO7CcYjU98a75u/H2xTgT2w
wwC0wFr88qJyIfsb8+/IcNYsm7mYwY/bvfCb3A+8w+X8d+53jttFn2S0fJJIciFQgiQGueZ+WtNb
eTOF5EBY1Z7x6Fbf+xA5x5hRW4Hn6wQm4uOOXDtav2JfptioCmpN8aSg6McL5snbdz+0qOBTnHWz
30860L27n/jkZ/JufT/Dljj6hLYdx1OWSdt8zMfTPNQoRVyv8Khd2IPpac+CYOMXdCeV+liN27ug
JhJLS2QFTvSHNMbiKVVfTIjkzQtPKtjowJO7YSA2T3wRr6f5WLQcacBvxbZKKFxJYT+8Hh4YIXxf
1Isr0gXTxwSkfJKAsL2xVgQhXkkXpk0WzphewrTwldNXyrkaTsc1VCo22JwirdS36RlIBOrNZlmz
nu1S0aytHw4lsUqtGIViomxU/3+rlvR5Mk9GQS9SdgLpBWAjeK+NaHjJtkM6IlZF+Niy+A5lmsQJ
DzS46RMMWrx0UNI7aP6EHvSMdzB8SN2m0kslRlusiWrfYNo1EgnBgpJh3MriCErnJIrYaZmfiAyX
jpZVCLOEs8f4W5ZabZyrBOFN84PnQKy14APjIj/ObbMOW5PVBk8MOuoYfLl7aomK+T7XFjl0Zk3u
UGHEU/pTCB9uLavFqsqQUQE7Wc4HFrxBOXmQW/UrR0a91MLnCMppnV5dN0f/IoScC5WF6eKY4vLj
1H9x0277xIdQiDbvItUX8502MhL8OxXKVcvLWYEo1XIBCSMXvGDwnv79Zh00c2rtiQOWpYKT7gFZ
j+BK60k0yAvylItKFUjGRTZ+/whvtexeDfhESGOjHxD/OjzeetAx6px5m49pf5OPw8PNXaVkcX7L
u17wbmzyL2PRDHOwg4PLrilPYcE+ioFShIpvzbbhatQ/LtXXrqROTTuUdHZdXRn49A7hhMOilhsu
RJkd7EMx/NX4Q0GA4Hbg1eAkGwNeNMsZgZ9euq13ND1illHmf4tAtMMIvQwHoVUxcQbSdlomtkjc
Hl7CLrccRt0ifgOs7tcxYDJ9d99AZ45AiZ6VIGFg6pacuxfD8TxwoUKMLzhkU48ndTZNZA5ciB5e
HoOerAqAl755mQVx+wx9aHhnaU29VuNRcggmmyh6BbIJVizZRG3z2XGTEJtNKcw9TWN1RwzLr/6M
5gJNbJpKHzUG1R01/XgCqUgeHDwIPoqUP7Amd78Tkmn2JwMPNy9729M2/vEBCGNaI7Xv2+9QARgw
Rxfwm76JlCQ2vEThICjQ4itzHYT89AsHT+s0jZoEVFmfVIw+m4YKRTC1L8itZsDQcMMr8vS2tvBt
nn5OfgJrpjm7j+oAsNocEtjOoWXnTrTUthdQqnSLxutn8xc4Rg0czVohJi0Sz6DbAsqYNaZklO5b
OPNb/7IQ/3MwX9D9/W17/yxk/iM0pahsPp0nVA0tV/eUK29fF1Hzmz+xowJnCvmYqwELTo7ZfU+c
7lgmaZlHUJl/+yLP0pnXGB0y6rKDPVgkG0JE4KMr4LOEAdYM1qv4iB91OlmQY21Z7OxkhDw47COm
Rv1DQxEReJQZIHFTa9P5NkWuzNJH3Y3+4URK8qRV2LZymv38M5LA0a9Mh3Aj/2Fgg7o5BDtdat3a
RM428bYGZDq7aXXzbXJ8stQke0NAsW7KaPXDM/oitMHg3oz7sCW7Tv0pG7QVrSST4nAqH0FWk7Ul
8LIRZRigrXFAPLroQiAuNKAHXjU2igc1o3E9HsapiUIApwu6srHyy7ENy3bArwH36MsA4VAsSY+9
KxqyMdAbqUrcZp3QEWnO/xgKSHHdMySyYCmX0a2vjOQEOcwsQ4HnucuylWfpkcqtCI3fXdPaNmhy
v+Cueuxzeplw3o0S//66m8o3EY95PyYR1bIStjtMYZbuIYe6fgGyaiEhkc6E1HUK8fx5dNmwY/2w
k3rOxUyLjcv+zJbNat9HROYW+z/Mmf+QsAIEQH7zj/ino+Aw0OZqFP2tYkLO/1x3EIHHRzBLedqD
jf6VwoE6cpTAC9IdFzpdxj+50i4BSASwt8+UQ1r9R2z+cgzVy1y2wnoIA9H2qnEsb6s2tssDdr6j
4mBfHqorXx2YO5mnVit0BX0Vkgih0cB1yH5CVjQwcJRWib1fnjp/U+9QCwAU34DZBDmF6nmO76jL
vZvgxmpXklFiDj5zRuwOnWl9FFVym2zunmcDcddgaO8vJhHYMeD1QndB8IB2jpmTL3tg5NaR/WW8
o02qLpTqxcbq6LXOH2f0S1Rd/FrldRInjmnJVIdZCW+tRMYUoAOqj6Gj8xq04CkfIPjuzojTdUql
5EIYe7D/qyBCkQ6xNTWIrE4sAhpP6IuU7oQeQa2zjRIFiA+Xc0kjF9hHcXI64zXIk29n3iML2P+w
ijclBMfE89L8sCZSdTeggeEghbO5lDjo40XI6bXkeMXn+fPliv+h+27bOlq3AT8uYqnDjHdndxzt
AZuogeuJuxg/pNkS+6CgsUhckUcbrShI2jcqcGopb6IbCNEaXnYBdC/K4n18qnwA64o9E3tKyl+/
NYkQcOVzkcv4Bb2W6L+fLVg6X+TbaUQ6/Cp+g7E6mKb5IuxnLs3/jzwanjzYHVcftOB1yR9sTVDI
Ta369mGgk+dJ7tBGF1PtnRvJpGqmVvghtVc1TqifBJFJnou40m/aU3Fmd+6glUAbI+ZCCwGP6Riq
2Q8loFWkE1iJnlA3MbtZB0afCBr/o+9jJQHiUQK3SLu+5VYcLLSoApDvelb+qauaNB4pbvKzJv6r
vgyBgVtWTu8zSpNxiKARhTWZ9HmIS51Z5raRbGEMjC9FTI7J4P4lK9ZzOKNaDm9gcQmTWH1zUUqT
MYouhvm4HM4Ke0xt2jsvi0vIYtrsKQiRqfYTQ/SOF5gzlzu5tyoetm/sZpXk7kV/JgyJ0WR74qFz
lSHvBzr2D7+VKOc6L99L36QndP1IG7BZgI6XcLoPDS+EROacOE6crlM3FCzIxS3AC4t377NcGh26
BTGdtj9Ijv4KI6MgGbAgth3Xbyg0YW3zW7vWYdBNuUES0R4xYGJwMxVL4SEcFx6Z/OBWa04Oub11
G4RLZymypbHs/0olqVz5wOJHAFqSXB0Q3FPMIIz1ZSLMdAUoSPacsB8db2rS7CqLSh1/gxOzJHXA
bV0bXz4Fjq9/h0Bbzr1GlUbgr9b20Q4JDTSHZzMMH7hqHpvKuFb76FATu/8RdJ8GfUXpMNlCSgr6
7S7mrg3ubGGriAAuYKzrd3rCms8COvfQJLAMVHowTeuDbLSO8eftVrwW7+4Hz9Q0I5e/zTrfAxBv
vyC+peEOgZ8FGZR64agP/Ft03nd8nNgHu5EkMy1y5Qx8PaoQZRQNROGv6IocRsVDJUZ/RpKOdZ22
Uze8MGf4XsgghWRzo8zgXN333Y0GPle4Ctk1rSAD64aQiZFzK3nVU/1B7VLnSipNFiPXOGKztpBw
4DECoIxnNGm1ojoeRk1cdz+QqyEYeZE8k3/EgKWA1c2iJpjx+VOVeqV1Z59PC1tNHATTDI04P2UP
UhBUjFP2K4Kjh7S/XAe1o998uqGEwIkFg+FGMP67Ntary/Dcm/aaUShz/olwIGezT8lq4PBPzEgI
9flSatgITDt9L9Y9UQDTkACQ1EJughI0QXTce/eG8u0KZOl3CrIVVYXoWikXmtPmT3l5w5wuOyD6
CZJacavwWs3MNc1V5qqpLaACCghbR7qFFmXRqUhSuw+oMlOmx92wsubZUf+UYD7mBq26Ha0kl5sS
jJDJzgcSpAaGN8LjyDHszpEjiFs9ZgwbjTMZhZkARe/ionjfCxOik8mAv5XlbtFgja4dACod09ty
8DLgs60JzXeJSivdrq56mqgAktL65cb6ngl0s3Eof5HBH9kJ8VXxJ3UOoLdm3RkNocJmLby9/0Xv
ZdOCaoale2V2Nd4XxxjnIWjl3qZgITpjYSXD+Rle7rHfBzJVASObzOq+MZHlKPEAl8vdn7Ip740p
tHMBxtVCJvZDbu3cSn88Ln6sxl0eKqPOedcKk57m9/7JL2HJaWTcYykMSwDsI8jYWIYrItTeJHbF
p4E89pjD661zTSvgtTrWmWoAPjgGhSCnXMYu1z8oVHWhCkqsxeVLMbSD7P7eI7EHMms9YsppDIN9
/9PFTKOFC9PtCpFiG7D96zIWgYWrCooYcafu222xFhlaaHL6hfRUePll/WH+tLLiAzDKuTjWVQwS
Hdu09KqL5ZkD6GxOQC+BMmNAN5F5JiZoNk09Vr5lcXUNdAIydhlofRMIZR4stYmr4S7cmr/m/CQp
4in5mOnZ5gREHgTCP1CNdXODYXV4MM3jSwcuriadY6wkAUbG+2l3mPjtF/fXrW8ClSHZRKXmoFJS
zgFCL+0vdp2/YnvGerm79rZ3sBLcefYQnWswWFqqSI2IXJQE2qhj8EjHL19Mwp8Gmnod9ZNH5OOB
nnXCao/wVtdERHW+D2Ay94np/W0HHLapXGbO0rH4i9X9upjXFFIXcSZRg6+HvSdKjiXpVj6KpeKI
Vy7zuzWEud5RTqnwmTspU2e2lAG3wheFvjW+vAXeslEln7SUkqKXRKy37Cyh1HJwtAWCscPbIvJ4
CEHP8ASgc5vg1WYw236bm4NcJF038qlg0/CxA4SfUy79805f9mREUuwqBq7FjtL6x3wajDiPHOX2
Q3XZDFz9ZQjTeOo6m/u9BEm57b2/2Ajp2uxurGgoNdnRk4ZU71jm//glhIyD/vXfEDQZI5G2oqty
XUTzY71ZhrdTtBeK1TZkGO3P4uRCL3c/kpQWFXf4fHuztZDZz6MUBqRkZP4hQlEEEGczFb6TsQ/4
vnWUT6/O/ZYX64AilcoPxSANk2JPkI/XRHtIX7aPTHLDnF2frdmqKJ45wlkrLJCc3e4UU63N3MTr
1f7DesVKjZHYSVBKuCA29BRQ46B1WCXPU9muA3iZLQfoStFOt/QOZqByR8trMlFFuOc2lrsktqgR
J7RrOFvXkGNxvWSdMjrsWi3c/SlrJcolf8eH9nFssX/pM+1MY5sNvPVdn/22HUtTFX7/eTP3q+O6
b35hR3JkNHge6FxBQAaQlGI/l3VhGCXPwyL048JAy/eUjakOJ6G6y4fNakgrLUv1z2P0VHbv8WkZ
jjbS2aZUb8R1sYQKjXdmYJzL/s5/+rnj8blBPFTWainRsJKnFeT5zVUFDh9IeUfig4vDSUsqBP3C
Lgq8BW1+IQmJ+LoYqKxdzRrQe1569Wpc2IdemjfY8Eb7g+Chtuiazs3FJgx4dBgPj3VSfpczq+Dm
Zt2eH2DqCg+ONH25zkfbj7D40SJEIaAwtCWJ+PTMsKCb1yGfZLq3z4oG1B9l+biAojocSBm34AUM
zUrh4PdfT6XBXc7l3qoESa2neu/Mv3uiUjWOqH5T3/BT4iw2MgCtAfon8nwDp6d8MbLH28bOeIKZ
oMs0VtOO+kFstmDocW4NGwgoBrJYKhWYIFq/dNOv9UAWxMsJHeMzBpJg/h36yClMf7Hsm9vPGlGR
pNmbYNm/A1Fj4btbwksZS3+rtaysbnr/3OPZWSuCdORMCzmxaBEX78HN1dqrnd50Z1ELvlvVZhLy
gSYPIgkYQpOwJBSKsXf84ADXUU2tmacQwUddgCpDr2Tw+tpIolnn0DGskWS1RPKKY3kW5iCC/Sb/
krStm0fKqQ2kTXpZO/Y0tyGJHTGBq8ds/wofC7T4N/UyEU59R8sEillW4EQb7O3NrwiL7vQo9mHy
fKzFa0PHa/GcmjL9unhCNHgE8D0z9xffjNWt7qYCsmC1AUps0RFcs/JhVM3BvQ1JDKQ2i9R8lMrd
4sUme4W3VQvjR+BvNywbTV8pryfYeRQ+8T04wBAkSEg2j43Xjsl4y3PeedYTEV8GKXeGonrhNgW1
wRUecdI8UzyAVqrvMEfAoFmAPqmURGsb/lmiCwU1pRNn9iQ/ZPQPiu9fbBDskKyvvgBv0XI3E54k
OpJfxDKGiaRLVrlEjxz1VM9kwfZNRPkirbTWotKePtRSQOzI58V4TFJUhTQwwVLKj13Zaplk2zSp
xKqCkn/M1Y/CKI9yys1dzevFChvFoTna144xk3lsiyBEM+OpUgpkcCRCp3pFFR/WVnT3zg5BWunU
fDJJYcsRRzWtZzizIXCDFcexST7DNMe/B9MqZNuvrVkPjwFW2FUf4IYdbQe1SJeRFtW+F4NlXrFb
I9Dv+3olXq63AmWTLCnDJ8uJTB3f7vaIUp2ELmrtTh/S9r7I5kfMiB+SfWYsRU8bxbSqQeSgbya3
E+Rg+HirWc/HNbOnDnF5mFPI7rEg8OpMGpaLJOy0g1M0OFrCeDzK046mL4iLAc55h0wUsXH0vtdk
nPk2vcmeSLKadiSV6oee2C1MmN/bYEK2K9oSbMSxeLka7SaVYhWzA5YUz+9A5eCiakblJTBiKhMI
X1WNw04zwJtI3YeKrYBiPoSXQwxO5w5qnbBFEO0A1pSk+lmCDVckxQZ8Gi5AP3Nn1YRv/3p5jyxz
yE/8GYOjUe3NrS2KN4eS/+M/ieNWX741Ex+ob+2BpBpUOOyP9plB5xfMo5eSeFuzn7mmHhjEAfNg
CvRk+IBS0J8k9fQ9YbzYn2/mIejTq5chktHpRgVPArt2ssS6CVo2UtF+JAQewimBP9E5OhHct8rS
bj0EKJnGWdpQw5g8npUb1vs6jUH7R6+rKWThh4lMABDZQecarbWibenJ54u7Q0+UBJEWeD+/81jG
q/rcYDhDOKeDOFMYXOhltNUvyStjT5BWC8vp9Xj4R8CrwiZRL+h7E1o57RhCng8r+SdfbYg4mVPW
YYp4ecyG+MGQ0Clo9OPxhOxHUArohRkRRhKnaCWP9HbdSh1VPQoI4vgezu6yYRNay50tt/uHk6hD
ocm04o+5OU/LIHxyNnAx8XEjgEir6wuAyoMfBwiNcr8Jm6W8hGj+kCCXz50dzlGsjMcBuo49qOHj
WVufJzauiObMqqnLWbVMZOG2wicUReYtyeYe3wA+93dx6NtT+w6Bq6jK5G5U3f/q7XMmLfVPhCf2
DzVtPW8tcCBY36240ujnIBIyBklGxm+PxOMR4UIv7XIMnfNddeYqDzjZl1BLAyaJqZM4MDHx/EqE
re21OgkqHOhzqtMNvsqKo2G2aKu0+ON7y3YffWFzCevNTD3kf0uHqLCVb6+hq/L89KfLgc+osfOf
RaXI4Skg/q/BxkLak1fzlglinHWD/+l0V2qsITfibau6YY5JobnLaege97boM6QJdlhReG+Kv/fV
gicCM/GeXRLc2UdpON386vvwlTi9s1LF0Te4HBBHb5yi7aom/uXOUIp6YRTcwm1J6xNIbCzPP/fl
R9HwhD943OLLN3ij2SPk3FvSBCTGphXZ4kXPCvJk8WLY2tNiwscm1mH5ApfJ+Pjy4ymOqip/8sAa
9tjND3HDdPtBV30Qofrg3jx3CLnJrIa2T3MfhUkRGRJ+uEY4SKrfwt3330x3doXwlhpLbue6Gagh
ETs7eXjFRCOXVCWHgpqyuiQiP8Qcbd0YOp3d8r7EsMSk41ahdwxI8tbU+APEeCQXbpNw/Qyeh6wf
C2sxKU+cFzjKbQkF1VtNWts1GYh5Zo8Gxfr27QTJ7o99qEiVx3qM7k+sVXn4cAjuLBQyk2o6xheD
r0ZPfdfidMFIXzpXzEdu1UZV0/SmT1BTKBrALX70MBwbwQcamAac/kqhW3uMg5rZpj30Xu4Vh5EQ
y2Ep7TFB1WCfb34/WgQ9C0F3GQURtCQ0OdWRb9xSF8Fsh2i6xrwWTSBBikOmjiy0Grlm3r0ciHt+
AfUvp//XVIs8T6P/ZERdECJjUeC/g66rAQrGDQaHSPz6lt2CJZh9aVx9BuypT4Ue4/J761OVekdR
Dvu8aN7IF++egqMn7ib7Yf4mK657hoL+DOeV2itXS/0n+/zn0/1XXgma2ctSqblHCjSdLBj6p+n5
eZnUW9V5lIR+HYR7wXAOoEeL8gv9FtmNPWfl1byLnpEO+h9eWQRfovaJckARoOEzISbaxpD5kU/8
yybuGyjd9wlu1hgZysnWhQca2JE9OxAZX7vrkUSdfzVOd+oSAXQQ5p1aVbH1Go7LW5gi4+sPHCOS
jOHFB5zU/11koXO8kb8G0WfJ09H4yyMbqI/HtVJluovYL+E+x0IT3CaUtybevDfUtfQfoz69jZqr
ssVHvySa/x7Ysz11kYpL6CQklAXlfDv7AMOT/oBbIxAEM/2OVMg1OvPkb16ZMhs+3/dxYQtHxZvX
CUedhf5EM+FfUZOaEFrHI6FGpWYY6jIMah7KeOpwXBszundq8L24f8/HmiGwfpfiU/gXnaCf1dCy
x+i4G0cum0YpvzEnbACYKIhEsM1+NisCaCCk1fHOsUed/0aqshnxZk9vH2QMdShdV7J4sbQc3R9M
jy9vsn0GV+AZBPoBIjWLdegpTpd82jCRl6jrhs7DyG+7FdfzxKlfEhpC8ivwoyGNzs04wpkieGrH
REBUpoRAKijG66D7QQrv1ItWSBDgCHIUbUWn1vOWBCGP2FnvszEFaw6+ZcmroJJy8UEVXCbbsHHB
jTzhKZKMqYgmbniiX6aWbXz9thzxEuAbeaHNz3WMbTsQr2/QsCzAR3+/tfiTyVODUrhlBuMKY/xE
rZHfZYMuOelx/hPfvm3WOpfqfyaED1KS+6T6ifHO2BtOpRNxnMZmTQ8m6HpbdppCfNHA4NdS/8CJ
RQj5gxPDYBSdED+7vWoDnGuMooAIHYrueKw3f9BZgllDBP0wlguXSwnzwphvNJmswhNZTZMfSFH0
2xnm6RwN8H1gB290bNRRdzZYn77QcDAjzjgO3fjKnLidpOiyeATXFup2hr4icTWHy67DP5ihBs2q
DEpq/oTpwa65SCWbrlcy6SLVvkarmBnRIy/yhjYJs1iGG3zV2gnaYbp0LV1DYsP+suj3ZmuaZKG1
rHkUN/nC8OH//BbPSpqXSWWclKlat++OciQMw2DhvwZoREPTJhU48xKPuJ9NzY3cAw5Un46uUBf9
iDFVbtpobfWvfBvZU888BigvJX9bEfjFvLJwuW4/cuW7NjRfEyyHGxcsPIgurj8TxEVshFl/Fj8b
oqSs5HJGFICsWO0vaIZZdVqhmhOoi88CuD5Ox0F8j3VV06VEIc02x5h4N5wLwfEf+g1ZG4lDb6sF
CgSSHhMfJyVH9tptM1mP0afW9PQBgamypG9Rct4Pb2iB2hiukFUcW5B1g1wjA69WnUrDTMX9RjzP
Jx9McOSI0QgRnwP35+Jqz+L1x3OfUQWEojwawDviAcrlpRiKy3zc8yWMgE87ueC8pgbtyPcaJUg+
3x0kQz+sw6MRBCpw0mC/bPbprAT6/KPWUw/74ZbjJkNV9C9kNV0ZNzMS41I3YXztI/8bV7dm+DqP
umWsnAim8S6HsU1vPOd/F83WCZdEjOptu6GCbjwj6jfBkUfQpgfirmi2jgAdrV6cjxuYak/wYR1W
4aWc7B85wYB9JByecA2vqGRUxw0Mee4bG8TXfwKHUFXxBUVD3wuC+weEkT4qK6DOHxqR90m6Vmeq
6fCSMC4bkPwZ1rflsBDkfy41kdQGFlEooZGG+Id48BiIlUQn9gCwWoB/TPnYaIGtyrlHOOp/L711
r03Lns52i3R53WlJi7kIPDsvh9G4iFniHIqPSe32aa/9Uyj8+rSqn1UwuuzminUSwUzR6lLi9fxX
JmGgAU4Ry0KIcZkgZa0U3N4xqhFwbeeY36/SJGWMA6ZWWgWTJp0VaUHjgp3P7aFtwad2KT6qY/Ro
FozoBgpNvFRVRE86gi05hF8p2eeFexRNEIBtT3ISzODssX45zxkPvregqGQOI4uvzL0YAGH3SwKU
7XlxKCJL+D5ymyXQTDYJf1gNqRy4qSMSN01GuV0wstMs00kiGiD+VNJesDbK/Y8fCT2za2gNMnei
/jeQYt21Vv10DMziTLXcfEYFZLRoMelh6b7KxXyzMRkNnwYLclYVQkwJMFoJBXAFAa8FCBsrYOyl
XZs91QF38ILiTFGzBfyEyVELCgJYcqhZfN6CPRbpWZXPNoc3qM85vkfNxzeDLecU3AtWWObHsd7Q
w6Ppb7O0R9zinzds7UXJyJl4jxC6vtVZXtiwfm59IZEkwe1kZ/5kr519dV5ScJzzTTGbLSGfytoK
LLsG3/6Uj9Niz6ZhIxRLavHa1FN/tKgu+5gvh0DsicbLLlC8Vay2j2UQJja1u3XzGwsWnr5twBLq
Vcbty64hobIWAOBt7/yhOgLtX6L62fr8FcQZb1iXH4WUCqmJjO9mqQet7NcWr3RGwMNBjc+fuJMr
PixZ2ulupPn49CRuwSoxLbRTVdoh7TA725ytL2tltrX9tRVKhUPi/U9m88U8kzbV0KJC6qjWS4GV
x9Chw1iUvSQ3FTRXjDu5lfFkMUIwMUGxxERa/EmJLV3nccJ2bIhdCBKLpa1C+UuOAhDB5EQz13fX
GmavRF7jQRkCz90yEJRJj5iLSg4nOYsjZFOow20Xxp+DN/BCxmSE4HUUhj2Ki26PsJlxpjRfw8Qn
pth9cQZBl4Xe4pyaFElYQVaw/TJR0OlunzmVmo6Q/TTK0O6vvSB7M4cAq0TLRwK2N9SY1997nilV
xV6Yg98eivbJhAisqdxOP4AqD3Kifp73oQSqe69MwfrwPMLyJ5rb50tKt8F3Uu0OLMqjY6DNy5Hn
XEhx3VIgL/Wbl0uX5UXBZbzbz88oYlyuE+YgUE64bZaUat4egFUFD3vSK8Z0Azz4bkJAsKmLEzSH
SXVXDOQpPnEGVvocJwT29HWknIaDRBovTFYsOQbRrY4wqIo2xUcXvvkp7ThQNNcdCgmJdGX+Npsl
vp9cw+LsuFMvR7ZxO0SO6wCCGXZCnCnKuqnuXbd7nmT972cRUklMGGrTGwHS72MKintaZMNyTBOS
N7GzmDdNrIy5TD8u3SZKmMu1getkeiHMY8pW8qqFuWHBcWrcqoLsM01oHpU599CSm6A3VQfZcy/n
CGpGewhJDPnIbesLLEWm2WBlvc8BD9DfGRYAZMLJpO2Pe220AdjO+WolBtEbhq0Y2MpxsgdRlikd
eUHoDbf/h2vvQjQpiF4D4UjezglbyzKqxxps+jyjBNTSkrhzZpwaqx25p0krAd8cXyYHrRQOOsQa
Qd68YaF/vLyDsdfFaWhVTs64QYwoN6i16ZHhk1vV0q6PmDaYQjrG2dmMm/PMo/rEA207CzC7bD+N
eCdhvO3bevf8I/549X0svBOW+vLDojBOVFARsZGyyfjXoh7bIgCqYrFUmrb7gYRBJSQXVkMQl9ck
wwISPAREp/QYzMBljnwaGihvPvbOQ5UAnpZtC7Lyg4jSXZ2TBBliCvWFYKZ3LfKqXtwEGDeVXubG
PJTrbJu2NUIJ0S0VBs4Iy8FmhG+T+8j4B1LOi9AMexEtTHSLXPsCd85QjjbH1omq66MaVTT7c8I8
24tBq3Dhfj50JXDvVCH5T+bwgX6mW0TmDnz5mhRkdB7WBOdSZgqY34+xD+6ZmjQy4IBf78RMOuq8
67S6uh7jAqz8TyVoby4+LhVt+HMO71GBYV8aBul/RHXpnqB/g8DNkGOFW5Gr/Jhkmb4aNgw+CcKt
eY/yscd/8+AjJnENEVwyaWsVVEITwNCNGtBmkIkKU6Nu0nlLHuFprhEQyAtFb8c7cqF5l+K1y3+u
ZJMd6wu2KqZN6O9rRdJz5l1pQUc0xsvRyDehOy/pxhfUfYLXxyJ2W1aeX2mre2baMveCDH6SQqRN
QdTmOCi2YVdBSX9C5pNXj9cTI/LLT4Ab7HDXGpRAWmID8tSwVX46A3sbULMQTyq7DqsbAUD3L3oK
StoRks932qaXkTS2XX0g/zkhhr0NtUoxdEdQpCcCbWN9sH9FEEau1v4i70NBRLM7rkIKQOVJTHiQ
f+rbUf54zPU2ced1PIigBna6xoAMfW96G1FOf9QqQaYTn1O3LmyqkY0f7q29tlKLRIRzjQteRSER
zsfj7CS3wi1zDW3W3DFXdE83/QVKDf1wEOvnWicx+Svi4rvTa6P3vmcx1CXvMtzMn+fHvINc9dYA
nWxPCX/WOSIiX3SuNfZ+nCPY+hyNT+aWs0rnqT/e4EmMqfY4gDSpf+j8rRXUCE6GXRGW1MH2b171
P/zzw3pK1kq5/tOnCJjtU31sPwy3nGNlgzEZCtwJWTaoDZ2cbhmcVw4dqrqsiTrJT/fAhAW8+0DT
X0ImiFUZc/0ScGRGz3udMKh3IchAI69u1ZZvGwWLsie8wmYzR1Rpm6UezqnELo8DNfn/cQi2wWjz
VevZUnkXWTY8f4hNB0j0Z16b/zTa46ZwUcGPgpdqlKJL7cE89K0xdc7q174xTBPaVzh+O8VhsWSo
auHf+Xh2MAyhU9ENb7wwQ2sXzeTASgW4SD9iAsNdPL45wvbIkNo3ghlcSDa6aReMdJ1Pyiubj6sv
ORb1jju10CNZT51/rOZoY2LkOxDxJuzR/7IvthMMtsWHkYzuck0x9ij0MFFIckkmgWFkg5/e2wMz
r3CW8ujJMbLJJmXZ+qrFxHp6xk0bapfmpc98m/ZgzUFdQpixMDJmGLe+1PoYhe83KzyclpCkNWaJ
GMOQAyNRAk6/EeRJEsI/oK3DAGqC7CxldBy9LbRRVXvjX9vwjfmRlR/nsvRPsy9omusUC1L/nfog
mh/w16DslCHZNU2MYzkc6V8Cb964kdDXR+qVny50M3+ybBG62VdMjS7NUBAWqzQKfYQTu4zZ7PfN
oDgbW1jeajHApnpTQS9h4Cxy8F/FIGAT6fRqRWey7s6mSvjnMoQf0WE8INrIL8GU5vdDaE4W8Gzx
WsZf/BH/VUaLFUxuJJ3+GfS6q1wOo2gF7djbHbIGuXR6e8LXtU4KjRWFy37CAUL6QlwR0oKITpTx
vEicGe+6rA8b03Wlcn76fjta1KlWk6DC0KKfNQrR9pvLHKw/mhUmffzvls9QFgAn37pQQvFvEhIB
xAC63jd/7lps+/UFgxkuAoYzJ9svFqiwP6c6SdP2Qg9HeIqjJVnV9o44GwGigskizKBAMvy5bPTe
LzUIh2wAofp7Ys2dWiFMWgjY3Y2tiAwRnrhW7zBtzKM/wTLNncKlZHoSg4SSEcAMR7OSkCLnffVq
qMhQIAQFS+Dr4uPIyCbu05l3ZYpVuDycMHbLpqS00irjcxFO+4+UktrIWThA6hGSGtdxMuE+vtcY
vUUtfJuk0vGD4s8lC/pOOIuaMrOPfbvTTAj2JXz8Q0uz7YCDDRSBVP/Te9uczgBWsABxMuNrTMum
de2uNaQOW352Zx5uhhRbR39TmmRiRZpbCfFB3xRbbDVnC/UGKeHGidgRJ8+/lAmBdrbpPhh5Cu14
jqWps/oCQ5kRxCyAW6E85SKx41dD3WIQ8hKfIxW8gPirDkhvsKcMuPndQPCcVw7IbtvZf+VvL+vh
ehe6X7CgOtPw/gaw+Wqlq+F55+JwaZJzG+WgTaP9Lg5Wv4/qMSKfRSq/Zx/ViQ15C2bbhXAGr22d
kQoiycCej770pmQqIPo1ovIGrSH22pgAR9rZAOCSRWP5BP2zotOfImbcDergt8QM98ZWa7hfoZ0n
s4E8CawTY5eBKby9ufK03EwbSww+q/aYm4DrETN9uNJSFd2t048LimoYb3vVA+mBHZFsz/WFwbRI
7VDZLLFii4ZrK7nPDD+KduJfKjbAko3aYXY6xtu98Of7zVa/Zk+IS0xXHtu0j24HpN+hNi1HoM7N
zcz2LImpYaKSsEBrYxT6lPGaz1Lpd5uji1hFESwHwIa5PrnvNgSfJOZvYqsn8VYpK2c1diY2KEYQ
GbcCHB+37qKybVJzEkJ0M6WpVV8ezf0IP6Mvf/wIYISMel460Nz/ooGCHYUwDqlKhStzsn7J5AaK
Tt599NX4yhOekM3AzC1WsijSmZjd6+wBpXelc8xEAPDltgJooX+M5mwJZVlngr1CLdE5kaV3kIyh
UjuR9PFYLCjnHF0U6mDPH/bTlZ46WrynQOlyCbKrZzIrxKTY9QLUNlZB1a1PdxAmnOWJtkOf4Vl7
i3zROSEpDqsP+8aLzSQI3s30Sx/g3bKSKE4X5u4miQtxY+w+ffZc/xHbQXUTEQDIjTBNPXbyQz2e
r+h6XWQPQewuTuukY/qYU7LH8YY+vZPHoGPK6t7mtcB2840eBNxNZLGjlQf5eBctjwfNvNYz4fM+
yuH5AETR8skXMQkAvc0O0KKY5mDFcEqdTRg5kSE7mq6IoRVbjEsj96NbzcytTEaomdcc0VWLwCfm
a9BFfdL+MrD3RhhntYUjp6BtTvURSNsbcPhqx+6fvNG9hAhXQYpxGC6I9pnHn79IRiO/xjJ/k27V
fBs3bMEwbvrpXOPeXAXMYzn61dt+EtT69uaXlVsz0GGKQ1Wx9k2XBfhG4ZL08KHdBcFWOkvIqr99
W3fNrjmrobcjrGzBbvCTBgJt+HVcFZLLqg5eq66+UhCNQWFCNrsRyLi1c9scLkKw6UJuO8HCs82d
x2K93b0xzv2JcY6IPSUvjWmexJnIyulLRWDDPE3t5A/vio6qTCQmhX1VXydD3J2B0Bvv/gXSbDUZ
TKiDpQmwn3j4clNJDLwyOO84M2t2SD2cKE2VyiN8m+E6EQhaSrepygHz19/PRqf2sabWdn8De19H
NQdT8BCblXb/BmFOYS5kqfEvO3/5h1I+zgtuXCMlP+DE7NT8j64iAvRx9BkPfsyevL1f/7p6rpFv
nKx6WKoBbfGOBHtd/leIp02DFRw1650EnAu1SYshVB0/drFs09QKpirdTYFNJkcuazlJPXWaWDKm
PcB8nBL2OmJg0VmLz228FTINJThR0O89+x3ZwOawExjZFAUjmIRYzwJ2Ji4/Xki2ePppiXsAW6e/
lrOisB8XcrhT2VlWHeY3UnvCk6gzfPr/8zluwV6CNuhOIh1amUwmS1lRMB5Nj0CX63GWijYF4cWv
l2R4IqMJ+Bw4yuLfBYunTkzwxUaZRjcgKi5bDmXM+hZxyNRrvxG2hrOObX1Cjg67yTgIJLw+AD5N
cptbqVmTRA5bRhcUA4agIvaGmXRdfyVePPec0anKUARbInm1EXa34M4hIAxilv/rwMinjG08oKGE
z02tdKABrJdw2twRPwfHwhAOqFCfLx5GWTXmN3lM/M/LN9utfo7J5G4yXLj1Y+ZN/3Lfc3EJsrzy
XQFnUg6jfeIkWhbEcyCJ7C04+UcoCuK3Okqqd3GHeuowhx3Aat/Icta3rQ2JltGmQgQIkeOWnzJ8
H2ukuEUSNClhFIFiyAYFvkNRpZF7Yj8n9lUJ8sqBcQv8SMQz62rd0nBR9fwkshrtyweazN56NW/b
Xz71e7s8jYvf12OUAEKZW0UsqIhOcspifxh0eAXIMX5Viw4QJ21F5f7nKwt5wnloJob6z+NmUzSS
GQHROJYpeYu3AI+u9Uv7NKI3gvzXu6j/fa9a/KYByhhuNVhfp542R/GsU4RWT8igPXoH+h3WCV9J
TDoQbuc3+zdVtQCERnV2dvdya6BZc9kp5SAE0CjnEIyxcNSzIsZBFv+7S3cbiSgVPHAnRZUy2PRJ
j5phLkP9DHvlYeBW0BZB6R/xnr9jKx+spjlQRna22sNOniSt43i06Xcd+AYkOClVj+teCM8q/SUS
67gYc7wgOtTwh4Oaxf67cHF5fPG5VGVQmjAdHphEMqcPFZEPXGYXa6ur8ikFuVeBA+uK+FnLDd5x
uP6PILsDkn0Vm/nCebVaZJNFEADoBHwz55MnBCy5y8DouVOa1xLk4mfeHb/qnbTNjD8KSx/rOJU/
6PrqHjxtRRqvpNYuhhnHyGmpXCvcHEGpeIoSPls47Lu2TfwCPKq8BeO8HlWH7NsCITGtBa76PzMp
KS8qMFoWIFXEEKXukIvc3NMFZlTsmepC7ShP0n+0r7V8RvQTzY/PJij5pgOAwIgGedYKk/Lg6v1Y
J8+oRrUiS3rh1EkUkVHPJBMNYjD8n6s1ZnYzw7WwAk2sImmO04nGz/ymqD/x5wnmYZ/+ZbkI5jTx
9ESCxqccDJp02m++PIIyH7YXJ7cO490/nfiG2iFK/E6lgHxTKL7C7k/Mb0Eq/raz5TdW5/65s3D9
Nv40PgD6jpaUrqH2P8g523Ay3IvljjU+4ej7lJ0j5CehLRMbpDB6jJKEiD1pG80f+TWSludrUOBn
Qi6Cm0xRmfzcDZFZx28DA2TlrLOIUg5Oc363qylK2V3zK9ILCx59RuF4d+Q8Yxi827/Le9eeh7mi
2//WAlIGyUDJj9rUHIuLuoAHL24hWnbzC5FQi5HUPnNcl11S5bU5DA3mAsWOZ38XrpnbBY4LJB1v
4XpYlagipuIJ6v7dC45Q/iulqQw4y73IcJGVYgs51PPBLvaFW983Cyy3iZvqQzmnrbHnEKChhcN4
wM0arpUp+q/gDG/xsgWh/Io+rMzSc4e12s2Nmaq7oNKwNKrrOrBreukDicFDflpBQjK4Brg=
`protect end_protected

