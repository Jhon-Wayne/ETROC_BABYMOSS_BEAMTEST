

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cQDd3XIPPlgRDhqULvYHvwCty2ZrVwzfefmANvx1dZIylIMC/SlAcj88wfYJOEUSOPC1U3p3rRJH
cF/G+RPdfg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hcwXqOGXIKp1yMXglvtwKNDD2csTguI/218BbAfP1Qe5YaY7t7J14bh3PN4/sY8v5SUfs5PPhYYF
AVoQ7+Y8KyIAkFOjVjl8Q3cizlaMAyaX6UCc4wmflvCCOjy7mkT0VJKPELyiFH5OE1gTiKu4NfqY
cLpas2QiSAVn/xZw83g=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JJiSVarYWytdLFzHp3wkrD5+jxEb6zxCxwIxMuHES7X4vO/81ppoMZmSB67P59pBX5Chyu0EswKT
bCRha6XDZljqkcBWrrqj3cLRE57UCaEr1RVpDNBMw7hjNrwCb9eTELEwb3X0mZPKBqVrRNroBMN5
Mb9o7SPJ2GKhIDEDF5Q=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
x9rjekK3vn0E248BFQkRU8rm2REs1XV6NiMfscimCVnt3moe1QOgVJzTLPCcPYvThLcZJXwVyFUX
J1k2lVxuHKaC3FNNToKLX7girUcVANbS6jS2AjaAfdpYmQXF6epSjXy+KOWM7AfrGv2r7XNIcV6T
P4He3ZDDIABlWanBaDiVD6NYtB9SspFXaifjJ2faT9Et8gWmYJogYQ4BjXl960BUcxWS5faBudWm
MidcfsfVFpzH5bJ9L+thBkdIh/P3Rjr9ssCSzEagp+1l0DsZGX583KqMaKiaZiIsR+KyQ8Hrld0H
vh5k+kh3k9z7ewkJNwM0LCpa2Y0qGSJOxIauzg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bMGW+/GNxe7XIGxZQsPwYg9NhBUySelE4d3DawPwcsMkcAefxMJ1JdlslSvSp+VjxIobQhkauqfs
plGQEEjRkhr+3m8iz7uiwT6s+TtBZQ509t+m12KAHsziCshi0m7JEPgqnpkYUxS5ZbKQCRgudms0
J1TIIpIIdBJiHjiJWPFKhl2FSk46olekE0MQ/LvS36IE6UC8sP+H2MLZpAxpzqHuZ9TNFvVcyr9C
pc7viw1i7pElJF0USsLWRjDFrkLdXdznJwKPhjmDvq2WWhH0UZss4B7FZEDrUrjB/HO8EjVy2Hj1
fpw3eQ84VC/StEBHWhh2/ovbE1xsoAsXeBE8Tw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pp8HZNaXt/evJqKzoiOa8A1cmkUh/1mQf/2Vkpam3N+hCoX7wAAqGU/zZVMPYP16RpMjeC5zeSin
YvUeVcdgv5x+e+joKUcjexTi2LwQorDqPIl0bCwYx4LccUexnWG6I9/pSM85Q6QNP03F3dTfZ+nY
q8I48HLVTNxhG5xD9+JTBp8D7rjXe9TJGi+hVikOsYhuY2PrwtvuAWhuicAfJnsIE23LJrp0i1cL
6oyVsfKsx+68L6qOWniySUGZ5yDe5zDF3WoQ1oHIZl8/tfnTJcGPsIRyeo3fpk/6/w5zWnz1pHuZ
HvGPaU9zIF3KNoE/3qKTDNhAcVbvP4+ohJfKxw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69472)
`protect data_block
IysePaxxzJCAR6tJ0yqBu4rBvb8nIRXT22NxNY01QJBjghSvDSHincBfGNDjCNTWk7AWhhT1YxGp
0f5l+k/yXWroVfj2d3K7Kp7WIp0Lh1P5Vu9fJnKbf54oIiDRwe5mM8WfL2q7GIkeGC4A1PIZutOu
1DK+p+UVPRgHcR3zqY0EBuWCguegi9cr+x2+L2xCSpShmaxkSUdkKs3iAXuE+hfFZerT3cgzjGAU
zY5+fsNsdzu6ORTVXKQfz9FAHihuUr9ERnwamBp6m/ied/DM7chCz14cSvl8/KRpbxIuvuO9HupR
g0tor66ixrOuH9hfSwvIOHszDWwVB4FEPRfYdxKLbmxUAxtMk8CO1OaXa/1ZEuGGfPW+A6BZLPgk
nQY2kmOA73OQ40m2EnP5OdUJ48vgl0BxfAGUl8kDpsef6jmhhpeGqMaJO67yE/i1VqXqzAKMXmyn
HH12hY1gaEKwcJcuClCOrjv4Xmp83XlAX439FVOi1ppTltj/h5HMiTrIXNNNI24k/2HbmWK9CsXG
+aEjPDWpilGWy/Nrd0ZsReQtLEaOH473cqQLYaYOve70byHerAel2SPHfOkbKHIIevwDvn3Eo6za
GvWWqSVAg1ugf+7MRfyLAJghUXXXxW24peYPkrm37zAw5OoeBHT0pElLuQNlooCaL5+SYIMaI8Nh
434y08IEaW48fGQAUoHv6MUkGx0MQOIFwD3+O1qjgtc6C9WNI5dB/IcDhZOn/s/fr0pH7EeWZe/X
7+Y4gO7cl9fZcW4tcCYf1KJVi5KhsLSd3Nrr0sZYkHCnwKemhAfCLBJM4p/ilxujyR2vvkukFPhT
Q1KP3dvXvr6dPZ/DvimlDt8YorVs3k7GdoU18m5WZY974n0ey6o0OwgLVCKnI0TRBB8k69C1kPg7
OKXAkQHpLeOMwX5aX9kFwSh09JqMY/3fZtopW4PAzPvloTN1KIzs3VJilp4faC9xnL47Mdf2zvCM
ajag0gGTmVR4AsNl5uR3N6OxtEmRv+s7HQx1xBzp2dziRl8BYeIhaWpSN3UZCNGfTDHVr4Ip3/BS
FckAfAs7D3mkVZyMG/SRzheub7k5wBhnVD5XwZOhxVHfZAp+Pdm964JkOItQCOX550cN/P3orDTY
/XKMy+nip7Eh/R3b0ZxcHJE3y5nSR4sgPJwSSJLQEPvu+PMU1gaES3GFpYG4aAVWUKRFKvbXlnfr
P2OE8BNjXMOvSxlzfydAo+ppu+eHJurDiAOAEfJymNjme6GuPEkifDDZRRonq3/J/2mkzSj5ekmT
3O9NqPtXyBoxoEZMSEKDMZay2m4mUZQ9yCl2eM5oedioLO2PAB0rz2qooO4wriBdv1wiiyzmSS+q
KKS0o+cojsUH+BAMVw6VFI9kUng3VLddGHdKOZ6Gqyv8UvdXfcUwmiBR6L2yBSM/sLHagQBQ9++C
TZdTdN/qT/WZFPAU49belmuPdpl28/ojtHvd/e42Xfabe+KvRTGKnBbn1c/Q32t7MUcVFZ28hwGn
fUbE8CQ60Tufzsz+WJ/kcYVGXa+cADEy/NgV1X4RrmeIH7v9z0bNBYM3zKetRxy6uUlepfwaNMgs
m7R46EeU7NwxtIjLFLbvLHgFCpAUE/8w9KikhdZ/oWaaN5FFiNp5Zbb5o3iMGH+1cB/1kESwzpjl
t7D4kBBSDeGFVgpJPyHhov2h4RYKs9MIpYAvwyGtMIh5xOdbtfymWEWjOEYqJNhUKLJbcX2LkZ+z
O2FAFJIVFDjiEAQpJv2jxGr1BLambUcmaGzS87GsiyV1+0PqEJpgIWc87Z1HMxexTl6iQbTxhAh/
Wf9YPdbLlCE7+2XqHPAJAyEHpmDUijDdp34mdAouKHOYnJTBlg8d02baoMqDWYHvRwwgWCQshAnd
nvZFMiSITeyx44vbRxoMC8N0KD9UPlJ33vaBGtruRDf2Yl9vyfb7bFxsxqxWvWvOImRk0y7joHqP
A8heVSPC4nyLotaUaykOW3YBU5tJmdyOFZ+biJuxuI4e4Hm99lgp01MQ6RUH44neqU3qn4A8fHZs
uJBZq0LIWmJ+Exiho7OQq8ZaB+qTl0bjle0O2dU8Yf7CDUAzEYTykz03/qUbI5RWSWuLqbJok0q4
uwl2MnBpmeUr14j8kQ6fX2+G8x9Tj9M2IBbeg5eGyGIBLWts6RMuDvE39+e3HKF92o5rtQn/DwcV
L8XO0urhXQnsq9xPea8mbtrdxyDTT4Yxrk5tJGytSYkc73F4eLrbAKwbnOZxFMtj/+CXvzYj0Lvy
PIcgPs7kvgnBzdfo6hrrz+VggkSbXICAuIWOBpbXJ2Pnk3m7VcfpfrKRTIzzP/qrKyCs24X5Ezt+
+ylyRFO6mHUGdYzBngY95SazcRScatxETxK/vCD0dV5c0BhuYj7gV8mmuXEIo9YCf/CWQ2FkeGB5
w1lAVaDbFqexBgXB1Z6C8pwS+xlqdtVLpZ9VFlp5WJfE3x/P2mDL+8XGJNVj28zNhXnvd+pacD3h
o7GAu4cE+/Eg+XYBo/Izq3hNLoYfhfuaqRjYkRhyVCykngUgHPpe0BdcKIYiXqbuxjz56HvZQn/m
1M8aWCbcdNHygPp6FcPBmmcHT6Htmjq44m0YaNeYL4EcV3G+sHnZ0acFk6ka1alSclUPPkJlIJ01
PuY1AYC8VEYSxOBAbGuossHpG+N70jgQIL0GUIChpuLWFy/D++GDvq58rMWhe7CI/iRKJS345pLj
r7mCrSNjpF5A8sDvf/6YsRH38B49GDDzy7Jo9hhr/MLOOsHBcB9EQpHOdnOFZxjoSvh6qdAx2xVb
pAxA790f2tIj1IUOXMwAMH9wrDYYyy48hrVttWUkbeyYxCXuv7tK4c/kEaJ9PTJC+DewTQozCHhr
FXUXyCRU0BTZJl+KqPBtSXq2JQd6oYICmP0YKtSW9H9Ondeb7Egcl3dIKxDfe/u5qE8wzx/lTXQK
l1y13r5xSOdpW1PdZ7+fYeGFvcPCSRzLSn+VhIepwRcLq0voRIAZIhWBY5F6VfiLHJWfxCLjmVRe
lyR2iD8oThTyiCNOQiH1IP5Ema3+7UPfHQqa85Sb/WdiLVQeLdT8hfJ0Y33sx3ucX2eNFK3w/5sY
Ni/gyJpq7MSKmTNHZDUDPO9YvnL6WGuGYoeYBCIZhK/T3qi0+eAFEQl+GMRkz+H7NUQfKSctWeK0
4G9kPrSSe7W2+u/aecgJ6BhECENCf5SqBVQcqPogZ29TYVH44+35wtZlP8hrxIYcRhsryJkEeH8/
F6evWdz9Kgg+IOW89V1fU+cA6Bo6m6CPSMjpgn74NRxZbikwJhaa6uKCOx4n2ezEvd2fU4QNtMp2
qRCkZ8E1saEPDWeKpBk9rNwOjqgCzuTxmSLk+ejXNswpxuNHzHuzrOSszV0IkcWYzerHvGQAUP4f
oidTRscN69YER1BPJEGyKtkgZFyIYZAhr6knKPZ03yeVxfzeBVVdzfxLfhNAJMfzb3IyMYyi3+oF
JWdrMWwDP5trfrqlCAhGtPJgZtDeOy+KwkBTkT3EOXl1857npjikd2G+epDpDdynYnZmvbd53+/2
E2E93Wv6fw0KPDBGN8QAMhrUxfwfFSqSNG8dYX122/ULFBUG//ghoeGFlmlyqGzimhfVr3O+fBGo
533vkS7tbNojQKmnUgVYJcjkTeWwLYzyq+Tlg6dGGnFGw8RQOLvbyY2hqt9yfkQmpnnI08wmDBiM
GqsPwIlIrFcQFggltwfw7EWndLIBwWytOqmE9t5cbjfJ4TBsXlqCFOCsuuiccjirdKErv88IDxa+
MYUcxrz4W6P8O83IwrXnuWz8vpXFiT+vSV8qAIUrGDrB1Z4TOw6gZZPvqudEwbSoaxL0VK4EVs6C
0triB3G2TcnmAocw7VVnf5E6wd7YuSX39/nuTlrrSV+yAc08rH01OT+uuHYzWIRRbgc7SrmHvwNh
YOgpj34e++nH9di30d8BrbrX17X8B2g2xHEHeyoDjdLc8jRzHYbAJRodKuxYaJb359WCFBeyvRyk
aCSFUIVYwtwJuOXyD7bVVVBkN3bJW1+EsDSyc5U8zYzr1l8zOgNGbCpL+qQZDOtxf353xPrK9WC1
U3aoNr6YLxwqwGjBE6lRjeE2Qbe8BwvI0Twq/GdPqkdiNNHauX+xITFWLCtbsMVyCz1CRgxttN2H
vrWlbzl2Aoa6267aTsDdf/wE2yp7tad36aOixy86uLIDSoZSBqeEbthawoEHszBBCW3EaCHy3qwv
1i9j86ScPizUOD98sKCUZ4Zyb5gRBimsC20vq3Md9RYTHZLVt9xb+CcKK2g4Ig9a3wrsVFOuiLEh
0EV0GSTVOdVmc2vFKJBOPrVoZjx0ryuR79wqdD2HhgpluHddKZjvRxJrqGRaXzElU+B5/GSX3RnP
Gpyrmpdif6wWQYL6CQAAwtrx2Ec0ETGptDKOJxPZIpdAnZgQ97KJJ+0WSPIPEJM7YfK7bhIT1eqq
m/V70RtapIl2MOzAqYCcnooKexNtGQ32Edy1pP4XnO/yjJHo85QUq700l7RbUA7lyZW2+mJW/ZKX
5reYA+MhCx8ApkrIFEnVFABuw/5xqaVZBICFUIddD7MEiMomv46PAyq00hoCFPr85BGBnsBornFt
q1TXag6JwiRwgNrgRoqVggiIkvUGiQaVyxEgZJF43bwczMvF1IJ+vEdp0kXZx/Y4NDBnP9NccUo4
Wz0xr8XYZazq4bIZAAiRk12IP7IbV1OEYmIxP+oPiRL1yFUDBOQK3YLelWmbhh6Ce9CFBc8NJEtC
Bb4y/Y1zQgYjv4hZyBFUs7tIWPNR51D2Tn+4SZ7z/U8K7Z4Fc0c2p2fMcIyxdSnZEovnCxVExAZD
Bk/Jnyxe2LZup3gcJsuadk7eEka5Ww/JfARKcMkBpTBF9JR3kFPnKgSWcwQhvoMCaooGk5nzlkaa
rNsvatNByBaIbm5q3XdVP8DZLiCb+HgLHGRNYWi4jzqYlZ1Y5IRIxFsrVISaIP1HArzeQO/aayKt
v19GxnS8Z9dTfU/AMl18XiJGZ9rqazBxvrLGCoRYpcwgRj0E4FiRRqPtaZx3KEhWNUyychGD+kz6
VgeuW9dCJGuwGNVdHSfiX0/8OpN5tDoFw6CF5ucJSzUyS/YevYU8QaFz7HE9spkjArF7XfG1tMcw
RGHXJw+4XWph8sj/zt0RKbBHaZpky5InsKeWyQjNeAid128ZQ2UERbljhoUQaHs8qAha6SbTplJv
KEKhpQ2Rw1oeuGaArDqvjR4pPiQD75rxrzR06bXT59yDaFPoiUbMQe5uKHq0AJUOQueav5RwvSwk
JpmIXo9YMLZ/wnCXiXIctEBiRgBrJhBTvcWelATiG8LqWdgDH1hMTMoR06xTPUBZI1vORFtMiAd2
yZX/NB7IWIMlGW1uKqEb45FYY51joNTwZnTlhF8GMHakMpnyDJQceMkLBvbOp3ySRP3x9HwYSWgt
jF//LO52V9XeRERPudCUe+w2tuRWNbTheFVv9VI2cEdEFub6LHNP8Vuwgxgt+dSrI1M8N+pL3NUp
j/Yv/hzUBG5EPJmJ8lqKiveDeS4e2NN4tQI6t+eBPYQhJ5ZXd5rTTW4Vh1pKRFW/+F0aeN16m6CM
JlkhPI+0GT5wUuYaOH3pFUUtbehpOZ+5yUMevAfS6QSBGrkISenATsRDrZaEA1z6aJdr/wgPV3Vd
Nrxhg1W8iApi3F9C6jWv6BZyF6YT615oMQEUdlpiPzl50ydW+/hqdnbh+hD3HAtoM/yqaS74jbhW
H/nEaM1S946zsaGIgy/BPPIl78HsCzQ3MmPDCHecFB7YhkRM9l1cCgrAvdGWb5KCepml60UYysvE
FJj0KMJbAuQ0d86oM+3jsRw+vJORPCQ4JYXjCKXnI4gwZ0V6gVZb6CNDYrwpVhs8UAH8riGWqHkm
0MJ0uTPBWoNRWE9QODw7xFoSmqwtz4FzmtQ0NXjP3n/CtkQBB6ZEG3dLVAmL6626UMlDEbuDWlXN
VYT+jHXSVSWE2ggAqnozo1C6zPytNVBkZEYZUzEQdHcDAxlrt/GGOuti2Cua9pYw+6bUILoTAYCB
lnq0y6LWJECKkMkFDybkuYMYJPQHZjaZHk2WQUGEuF6zq6kYoOaM0gC+87OQy6cqT19IakLyEKCg
b/HkalSc1rEhl4XW8b63Tkehs3T0zJEOSXI5kdaOMt2o/sgyptkNT/WIO7YiyBRcf3LaGND1diOp
j0K+X8uAbEjRbJSSiqwN/RWVv+Hi1997Ewqgvdry3SzOLQx6jnEIr/Crq467Z+4Ln/RXLx8i7p7T
JvSPfTM8R33RA+5Hfja1+BxtTWnzWNElu/prr98bO0hPBdZW2ksZ5atMVm5TIBRNHeKHsxn1g+L+
byr/ZYLw6G7h6xI/qZnCxjPPN74J8gzsfFxut9j/KpGf/W/G1+EX3swo784i4pKEp0IjU3jJbqqb
7jd5L9JKERjjJVqpfNmihpQ/YesM7eMe8B4dhVTIxAuSc+OlVBX6LFVk01/ImwptDdDVWWUflHR/
OTmYJoH7W1NojkdWKsw2bpfyB0CHg2vq22EmmZrLqibxo7GodUPr/JLq/rYtxAb9T3Hw4YNTc4/x
LHScYp1qTt7GouuTmQuSt4U/NJb8FKyQZwkv770y/XypG3aK6lQH7NfKTP+Ti5jdHdKllaiIDHU8
MaH2wIGawlu7E6rFOcXbGx0H/UxJi6ch8pptAqHwXL1fypqoPfpt5w+IqQEGvJfNHihdpK4wz7XM
Nt6bf7ep0OamteXEWnNZvzN/2kIGsOOzVUE66w6jA7xSopexXUqzRFWeMVtsSCQfkET7cuD78wzk
U+g0IQt1EetnaeQVnaLguVZ+y5qkw6cmRbqf1Ua02VC2ecOtylU7HnDCRlfwzTLmukiNiY56RyBa
eK1oXKyayh/02FB7e7f7BAgEOQt2aRUahLUggwxwhr2DnS53+cQNQz+vKKcBzlfIKPB9XoixW2QX
M0a6dqtebopm1IjgK1rBdoDZfnMS/rOmmPddt/JvWuhA7g6yDnaRd7EgAkjKSQrd/lr7panCeBCK
lw7xQL7+CQyB0mwiVgQ/qeebtXnm+kUPhLesqnbZ8Ji8BHjR0Gj0S+vDdzumBN1T+Of6Dnq+Dy/0
kqbHSPB/5fjjeC+tVTUVvsXUn41WRwD6F8fKXIwP3gzD4FFVhHuOgAWLXC+ZgKfXxyReqkCo8kPz
OtHd+bH7LP/so2irmxksnc9F9M4Eo1krr2m1Lo/AUSj/eODK9Md96K3ouE/mO4DP74rdnedV7oLJ
zBYxUtdqJnMjFfkzfBlhfC0c9MepyPUfVESHeZtacXmLP827PF06VCzbVF17BdC/NlPuxbI+jgDd
ijhWr6fxwEpgNS3EBHVNlXNwlWEqQrhIlqlzJQaVe7x5+kI7BGLKLiMCbC9+yq9H/o2Cvom8QHYD
spLGbrdbS0+s+cMSgEKqMgsRNxZ+lIvimfbdqZ1J/DCzBZVBVkWZeagdvJgNYYmSDtz3BbVNtXP8
rU4cqg4a3GF+2BDcPFYERYO5HmJatetGaQ26HeE6l3lF9ueVDM4Qn1Dqg9otnUBTSY9s2MSMKQk9
/afVmn9LKi8JuZE51t4Wi3JOFfh9stc9esncyzShToFxpM+2eNfMiInVomvn+fQoBwYsyjV74PXM
Pwq3Nle8cJTaNpIO4LXcgW9opHP9wLUcoODli8NOCnAkIOpPskgKLGId815zR6dUL6TNWSKkIZN6
7hjLnJvHMSz9EahAUTe6v+rn4xU3XNqvEFPZV+cIvjqCGbPvZehd48rgomsWhtOsZrGO+Q2Cc2So
jO4ryzQjrSmT0fc3Y1gV/JlUjvfolb/BraR0mDsY04SHfE2TJKshZyb7L7llYS8+tF3FBLO56XcV
QdWWCyjuzEt0zZUmah2xMpnG0EPKYtWalpYeLEH0KWFrMmvpkZnyRm3WrpaAbq6yi2LZI40TFY3t
4fZZyOHtl8NbEJi5bEApuCH9axsgwu3YvqBWRLv2lLZKHw2zWZAc6QGT5PbDTr6mFVV9aprDV4LY
86WuJ7H4LB/2zFPrG9YDy+GmkFzazfHtXXN8j/c1qP9ZcF/LiCsPfJahwlDORnFl9HV6vWHXFNzW
C3a/Du6MN50s+w5vQWapBPKQ46ZkPAKXE14Q4uKhykysX41TSrjvy8GhPKzkm7k6ZcNvAu9vZAZc
u6HhpuQq1SCQVsfnc9GhJZ7rEMj0UszhNg1z0RFYAkEnF9dtrWiYpiOkVVVcZPTJanM2ixkdeQtk
rnXOA+8HDpELMTPGZaa15iHcduMIX7mXEZ1vhZ7usRxEsX+/cDcYrsn6UGZvjnhLoB3E4QtjjMd8
pmGZfhN9PrCMGyVHeSrYYF+LQ4xWLUxCTsJuOaOY/TvUpXcq7fEizWvK20gRI3SYQTfD1kO9fOYS
cb8B6piKd/PcMctg5DIA5nrpzO158oDzHEfXHLDwj6El7bKp9/VsmE+lxU/S2YgcuqSe90ndlkG8
iy7Pgl1jgg858n4/Eh7APa32dVHL783QvVFb31+kIBUxlpD44s0bqqiSjZMbsDGGyX9+UdGY3+uJ
FgZk30QBfFPGB/bVopxz/0W9tGRHu2VFulkyBGPRUFEio1VyY/xukY99HMPRIu8XR7sy3S2rQllQ
aWhoVBu57oBoP5iegG7Of01hl3/Yuj6HlshupIWiM5fNlIeQY1sI4AiEKWAbt9s6d37/ptGUUfz9
C28zYNiYHCBGP6l632HiIXj/bsADC9rKLg+ALzW7v++yHZKepODn07TfJ//QQxvl3bTnKV8hQeIb
bwxmFuIqtj4v4JHrtb5hvt2qqwlPoBxMyUQGpnqmWf8Go8o9UkWzbDgKPLmNGIM6PiipkyL/i+sR
ZwuZfBWEgCjIHAvtUXvE/n0tcpEkgyWiyi/OY/ersyhvjPNieIeJwdpyuvSUUxIbeK508Olk8TGD
bjwx9Lfp9Ww3XeH3ebe2eo5/yFximpxgk4NSvnEuy30Q+bU/b3TejZvSc1FWoKmMjufCHZZmDyau
+fStBznPNIkuIzJ+akhF886DTtj/CR267IUWdFvJcxkHZMKOjFmTDDuSCFuOpG0hSERahAFfXsed
zeAOlBWdWb1IGi99XZCnqcHZkY1H9wzI6Nz9ziejdtadE7Q6NK7S/xaltrODhIxDPdKnSz1UTQIn
D1/fVzBiZtVVDQ0sJ8fNp8ia3E8vTvMUj0HPKq9vHwj4mBgNcc5/O50xID4tTh5dcyL8PftxN2FD
GbYwVmP7aEX9wUuQMbBnLFyF1T03TQRnlQfz2XKOrt+FuIHcZnBh76Npft/94NMGe50KAZxZ0MaK
cFQ2sjuyHYJ5ri1jHOimMAfyhOEkOoBJM26RrfjehaBNnrKOJCyrjvAFinPd04+x3ujFa88urwFJ
SW1zLAlZdsZjIs9VLrJ5znWqb46SC0gt4ZwNlqMsdFyDGnI+dhw7tsT7iGoYfLDyFwiz2JslUloz
Z78ePgXQoyOMDIq6QyIzKO6KX7CVNDFYw5mEo+QfXCwfENNXyMtSYhJOl6DYC3TNsTHDuzLgF3Sh
IoAIfl8U7d6dkcc/+X/h0jf86QHBLl4hZ8/cRwFG/Rg3gYdtb8M84ptHu5jIV5VpuHIJhB6TYCtM
5SOUlB71zxXx9HiiKkw6MuswNI7HeGABtYVYffK3Jut5euLu+V1J93aaLAC96oyVbwZM6K4VyS+h
/fWPDbdE8sX8CfVEpOnskqKWiIT/5BMR4DEXTmlRKtuoa0Sv6moP6IAfjue+IG6BVf77BR8rfTX5
XpNsfKKCZABgMEpTP1B0ub8WS9jV0wVvjgCqHsBdI1veND6rmK6nO949AvCQSqh/ez33DCBKyimy
wbLGO5nHhaID+ajPEXwbge8sOI9QbxUlHWZ+9JEpz4Gp45QYCY+L1I4cYax+j2iTSA2HLkTgRU1K
KdDDNIMGxOJf7Qjxkr7OPiBmow9oOyhEC/cpvZx3Mm8VKVEpxwf8FyJIgYvcFQojcmAUSWKJZssJ
COBVHnL1Bscogj9c2qJd+auLQp4cwRnvWQq7ewTZTeZoPXvZTR+iNf0/HG6MDt0Ep0N6Ooc31yQS
I0AzObGIcCAWnn0T65Rb80OCuLwqbuEyIYS6jLThFLLQo90b1FsdbqwXLeOT5nE4wAgG9t0YFlye
j6K0XWOtQqtDJX8UjwItsyygjq6A9ETfEilTjjAxHvoLmzCFVATwuYiIVSQr2g5wak7mFhLXxSJ/
/aHc6MFnCEpn52axjDLhqjUsLXv40ZkLqFVOjwxw5/arwE0BLudOiMXncwaeaV4csvYAHbyzbzH+
SyeADewy/PUUOQQwcqgLDpXmKt24pW6DYHpkiLwWQNQP380b4NVT3aAvPg3WwHgM7qn/rqAmE+P+
qsIAsoLmgQHG55pXMCMpqMCNiRih7Lk0OHZsbMuA2Dm6zrSdjYOv1XGA3qD1n8SaucJfWSnZ4aQD
+3SWIp4ZSvbsN8EaHZivLoTcbxFL+m/wOxsaXpEKMhwRKQ6XOLb4HNjSt9Q5hWJClJW76Zn7kWTA
qrnrAtqc/qhbQ3JwUY6zfdL2L82+HhxqJgf3xSTqdpXMUh4IoPkpy50EDr1aOuzKieim34Cth+Rr
2LKmR4feClgL7x/piOcYrFrRXarC2dFL9B2pvp7kJFgBFOkaDAlXzZJ1reudAdkjsD4mceEFOFe+
5XvK6H/ra1/zOJEkAAI5v6ehuNzW7aLvYPJcCmoVgAZCYKo9hfhK1HwAVrPnLOKxd9jkROBGe/l5
jWeJ9jBwOZ1+PFiLuKbMFozTiphfvaeZWbbjiYU2y9FcnUn6NOnJYVCPTltqainA2ubgyhio8xnF
rCHCnqF+DPwsyVcoUA3j7i5jOzCL4ZRpaKSSTxXHZEtDKyjX69NKMiHq5RnwPzgVqt58yK81v/mc
b6y6+8np2rTtKAjzLF3LSR7i6BOHfkj/Mdf+1DMOERoLC8ZrsyDtSctC/MqBxbqvqlDdmIXJildv
mxPBRt5fkLiDJAXK6x1pEc2VP8n+XNdtjpmjnUjvXDHhk3dnUQHMqp4xCuZzj+r9BRaS9kSZdZI7
QmD223WBocK1mbQifEUmrQU1t+tCUouhaS6uZjhwcAEEthok6LLRN1uNH9WrD3rTkE/zGXEIf93h
9C6sjl0o3wMCc22X5WjlUkgCnKXmfRL7GY7T7aFQIMO91Qmyjc/14wgNlslB0jIa9f82f9nsjgGf
vC+ZLQq49NyhH2Nsxw/swo0J1vGOU/YUNU6B5QPDIWdaydxK8FLN13sfSiRZQuHXEMI4SWcKFY7i
1sLvGJV112XJxAhykCfaPRJG0Wdk6jVgXjnzwg2zdUAAtA+tFBo4+kRm9IRZlNbLyOuOCv9Y1DXJ
LjE8FEZWayD0fy//jPX/YT1elc8OYJF97OwJfRYbYk3Qko3tbo9pkirSYrfyYsW3NwUQmAx8r7IC
hU7ngKL3vMAR9lFZS4PfPsGk+3yEinBKzjx5wrQVFSih/iKRrQslLRmpT76Dnl4LzNs19+KG+JiT
DzDWvrTqNqen+9xOW9HoCpEXV6amBMMrHCA3VAQ8xAGQ8evcB5jAxUy2gCIJWZNmZFlOa8cN52yR
tpaD5t6ubB7WOhkDWuTJQ+9IAXerh1KOKKiyQZ7uucl26y6/JUl2BTa+W4UBqlyzg+zqkgk7RUy7
1AaLdhWK+X9Fs3etX56T+M6/Mz/cU8o0EDOjN9ZAysV/jOPdbMA5F+RpW9NiTnq+rAu5wEp933BH
nGBPNdX+pxiF61RKBUuE8vVJNVlWLnb5TSOlwSZphC9wJltX4SmegI8LlSfMDimuy6wpT5dUKmuy
5TlWP4dZbCDmFS+WxqNwA5IyGVOQoXqSq6a9dpZ74l+GWPUTZPpTPUiYBXWD9BRt0Pc1PKO1PTYA
lKmpXQG6dHkCn6OLbzNAigOOti3yuylk3pt6EuWAu2IQ9xNVNFOsW4nxjnDLFBsoY2QnXW1Z0X8N
SeUj6K4g1Ipy6EG2A4hbAoqPcBZYqkzFN2lnvS6rfL8g67rNHtZP3itmJ1oqpmYgnJF4Maja/rZE
Vt8bTX3hJ9+QGE5raiXedvVK6ny3HVT6j7VemIVRdhuV2Qy7IAejujP7tXx/GuhrBKW0jILnh7de
SDDnKh5I/geA/KMIi/3OLuHrQnWcHahpGwAIkTqstwmsEB9Z/v0ltAd7/1AHGqXZZmy4IuRu7SpR
xNwqpFnySknOp4PqI+HAkafl3bW0+nhrfk1SQcKTmJwzRGWKZfEWXLuF9kb7n+oAj4IzLvQ7rGMN
UoX3qm8Tdkmr6dSMarXwpBP3zxcwFXqf4uB2R8eJPB9KwbpUv6gtDcMHr5RINLnmVDTAHrRomAe+
6zfU+CLk0uf35xhhv8zz9Wo5e7CRVGM9OL/t4cVm/Ou1GZ74AymCn4xD/ocAdcIVmTbvNOEHaWTy
rWWvco1oan5pIyvHmxasi0T5q99eCChynBtRHN5yhJSVeGI+XPaQ9s81bpLZ1pNBwIwBVE2RMPTt
Pzu9MW7K6iLuZgdE9E+MC45u1h2kqYF53GO1YSjyeVf0Sa9TdLwBkTv60r7Coe23asJcqHc0gvfi
OIKjZ9h8q19tBs9EyFNIkOR286uGcsoyN9xMFGAgoTT/gey0LzjsnOI7WtN2jW7JKCUitf9Dd1bc
MSq/IcItwuAZZsoIwZSHhI2R/qvIVVX+5axH2gK3E9lMx1A/T83s+c/wKt3y/G/i47kLD6qQoqCw
Lovwh9FYgL8zSS87Szivg0ojO4xFzWzpZwIwbffkxehOQGbUrUdD8MBFTAzhn29xYndvsgqvRhY7
/gQ2Fk8ML6t2RFiGinJIDzztyGUq11sfRZw33VJM9JL8m/2EuXZ5x2JtRib/1q78Xu+yu5rX0bWl
Xs+PUGpA6HxZ1X4eCf34CK/xHNR7R5pVmuFFP5g4NpUONTITRjbVbapYRytBVHbGlGFzEsWg86U/
yY5SaESRoe6QkCw5odyAft5K+N4KsSbruszB6BL8t+rAWctI35Eh8TBgjiAuUQNPUvHFhYStaAv8
oPp5PRRYrlNJh3AKKa0hs1Oe20oUu8r17NaoddfbP3JuKfpCMlweCsNAFbWpPv5r1hyfla2aR1eC
QL3oOFcXFxTRzSU5E/n0N3yFq3H+XrjhPW4+l6GMEMTRRAcQnerR4gi2+r5sQgZ78G7fFwzszMe5
Nk/DX9TWsVECi4CLc82rC2x+nCmm/geXUIi49WPCBzWpzTF6w9sf6CDcoZrpYjoTfFdXgDQs6uPA
9la0FlZWC4j0OG9ekPSnrvnER7qfpAnwcYJ60muDJBNX3eEnkf3uVqowsr7t9SNTYLs+bhKpzLnO
awX8PBj8v5hWBXdX5H7haGP0q4nAOLjZqzHKDxxW/Y5idP5gj3thzvwTvNeSzfkwLzXmqFoclreQ
O6xvNXYpJeVux9jA3i+AVrJdKmqR1tfin2muduJXDPedHv//D7qFeXMcj31H/Nod2PiPPIddonPI
3tPxBWj9Jr8rbnpZEbcr+6S/Ucw1AighX5Syg9N0OFLK9lHPTbsouYvMsBMB6yl8wO+t4doL9mcw
YkUZgu2M4hk5KwWcmgESkcnCUnuBCHhjCr64aR9TCbalmftqUMp55UY7jaMujGnnm9ZTrnJT6xW6
SxPeORHZSYgQ/urwfVgUNnBhkiv2uNMRDHUSeve//ymdLnLFiBjBnxxul8cin38+iBpLV+geaz9D
Sg3IRXRZL/ldZzSk9WJvKOlYMmBJxYlXewBMJi2q8zD+zcB+wP0FCQjtmFA0Na0+rw/sYwW53ZZl
nquihlAyH2tmjwZrn0yeCjcM8y+G6xq2YFGG7UbQgJbowqhHPEbgni/ZQQaxqv5Wz2vZfPJww3Hp
tLQl3zmwFWM9O4oMPToHTX8bPSx96X4GERx0EVrpfD78kN1RYdIZtMGUq3UdI8BmQzlrrcCwaGdZ
9fqMbUZUf4Tp0WHSTlqMeOVU3/oMgsaRttKom1mRHptZSbOfFfdCIjFOo74LV7W8aAxVdh46CLjV
BlA1NkSnsEx6NTt9+6U2IojUu2qRleDswOFCnpitbzdfhdhUHs3lBAA6Lvc/H03DoErs02UZlqOZ
XLn9NY+CVmiBQpzpbiGFkkaz+a3FwsnH8//RFq49rHQNfixKE/iLCVo3dokmTyMjH55qrozTSpoR
LuOzboWRCm1cPP8+MSUZDMSPxUw4gDctzcZM7wnqdMwlIQOap5cFJQ/xZunVNUdQ6grPBKWLaWpK
Hfk4v+qKbJT47neMPnpyFfuYLTEYgH7+pM9SKFU1VAxec3xz6fJW3snaIOOUIsjuV2hhFIaY7gjI
LjtLnWS103sUNoAznW5xnBDQWX6H7rYVfJse0DNmPPUiT901fUoJchd4mKnn5i6OLvf7mMN75zTu
O4mcCMHbIrzlqerX6arKGT+tHnVtrZzpp+iISPUsneAaH7OjiPC0r8aYUOaXEvryFx9bUSmR5io1
t6IwfYveT+LVXxsPDGjo0bpcvv+7c7P+/ae+mmEx6CUGpY5IU5XyC8wTQx+kgY2+2csppzycGDZr
JjOHDYqrSNckKWjLWTS+hDVQBuqK6UiJG5XiQvXXCO/LMgVqWEUq2dnYezS8mJYyOVZoN002mPd0
12xY35bsgGCyu2ZNW7uXriyrrE7GLeJu8aebLBCX4eBFJJYA14QFZmJ0EWlcA6W6pZ63rku99fzT
5YIk0S6q819g2G0239iYCagEXm+M8C0zXnXPVPB1qT7OPfZ5kZnaIFpSFaxeuuuGlV1keVkP1iD9
/CQgwmN6945AFb58bGQ3NAbZ75apbksgc4Pl0ct5PXlRmA5N3kt0TH/mlaxCAFs++aFsC8K9pvT9
eK37IVfoRzErgTXtoaLdUfH3dJhDAc8GaCpvwHIVdwvhD1CGYB5cOhuSv2z866/UgisXUlzqHVKm
toqvnb7wO0FDCZ3QkoA2b3zuysNcPZ+Ji5QCTYKqlZT06nN72aiaR/jDHd3V5C/QTLWy+/J7hKRE
X+rsObg6rRfqGZ+XZahgwvKNBoK1k95HLK38OhNuowFBCwUI8kVWCTuefIoTnQ+6KpDl+7BmOtVh
Fj2kEb3J2uWub6PwuDEbndX3BIfqJ4oMNED20h0kxyL4Splo30vEAAxWy/iwuIafaXy+2PmKCp4b
xMl07mSe+GSDylyQ3JqyAlkGZr9yTHF4Ol/R07JxxoQB6HxmqDAji4IAc85AIpnIII/mMEgmLeZz
ovJeCsphuWMgR55ES5grPAibeQp5DyDwzbvZE9HMixhTAUNxwCTl9eSRUkdzGRN4LJR+vwCT1yp+
z0CkufM9B8LR4SVtyijWiV8x/9m3ZK6fBwCQeMb7GY3waBQ0OGjq9FgNY414ob39JMumOraK50o0
tL66+75SJtr0l7tVgpQx2aydRfqdoAfPmYupDeTRrRZlB6YnfEkxsWYmVjpPCTUJ9Bc+Gl3Q1iJf
WSQqbnvxEl/C4OYLpS8tOO2tB96MDj01XJ2YMve/fIYnex85BDhgbZqbxAtCld8ep9rL2W9BIIj+
Np4TLLhSpOGVjs1lgywDrfqZMrxsObYV4TKC+8Pw6tX9m9sch08AdlX+a7BmejKUdTtQ8zSS4g56
PNKSvs1/UFMQqof0NFO4gfuIxzZEMereiG7Jbtj1tpzYkFhw355mZ32adqi+LWYASVXuhrAAHVen
fTi3aZJ/HXFMZo5ZxmB/4e7gtkuHu8Pi/mIcT992TqAclIWX5Hb8TbTG72par32gcPYScz6PoNLP
R+4+1aSzh6roTYrnHzHnFuUvzo2jI9arnqsOHoVP2BpppkmKqL8LuTAh4eyoLngi8uVwvnKFbObn
KEiVHvQX5uiQ3U868cz59lmRs6oA3FG5EykgnJ5a4JQ+Ub7y4hm6ZOnhkfDqsuZ3EkqjFLNJstPe
maWb/fYFwyH7TPkVxkuSbfQeXV+ogvEifvOsyuQy9s1Kx/gHrrLDbiELqhhh2Lb9aCq/4GaebSj1
xLk+yLZY/WTZatXMS8+CtUdIOmqWZi7MTIcjpG6cuOGIFuRISXb9ukVcJur2tXQs/YpRCt5p4W9J
504ppzf1y1hczfgldsHTjLl8EGLAgYJzDEGOcpxeAA7iQfIlkvSokmCg8GR319NgfYqceFCwKDK/
vN+Zb1jK1aqev0r4LE+/jz2RWw1GSCfldaM/02WRUDVAEFkgqe+joO+RuIppTjPxms6W65931Vxo
yLZcbucT9MKrJ4R8/q7e4j6WSzn3o0ST7xqBRMkHccmdvsZks1z4z1TzlL1z31TqkGvpB7KjCB0z
b/e/qUZe/Dvf4+jbEPNoq+ZYW4xXvIzo8LfZKwyeBfAcgts8O8KnPlAHOCNFLi7wII38QhN06d3r
E/5WiFlv5WXEUxLNLXyiBjnoKRN5XCLK014d5VNFD1sfR4gJJXV5fkTnZ/rU54fMDBeCMiCeeZmk
GpDsiphENvZMQ67NfOrBrDYG1ZRwgkp2JiE0fNfqqKXC0BknuNgX6d+YHsVsM3Yl6V3PyIgK8Id9
fjdqNwN1lw9whf5EJIKd7YxMwVgQjmwwrb+RzniT7V4GgyDAnK8eN5jsmiuKIlP4F5abVwjTxvPZ
qy4wNsSkXzz3PuL33LIolVpLvWm5TL4r3FhmuhnI+DNgbq/a4+e/HWNlcjFlcN6wYQC4mpwqLl8W
XGoWd6aH3b2CmPHQ4DLPePs7WYTSR+RXLQsmEQt+nmJoTfU46VNahUM0PTGJif8BWhlM5A1MLmIT
YA3C96H1iJNEhZKlYCICyRyUn2ctxSwb+SFYeg2U7FQZpskSH7fPZy5WvFBYem95ofpFJSGTfo+s
Y6Q4jkTNmaqfaGapuogmAlMMyxlrPbS+LF+3PsN5lgHRsj9QbK5KwAllyZaQFDXf3V9JR6zvdIY0
2Wl4y3UFbAIm7S7v/0KyAan3rjBKb0q7jSFl2UhMjSZfg6jxKOrcbEDSIrE+7mCLLElrpinFgZN0
7JlXwT0KviNvW6tg9oinwSYH48e5GXWJRl8x7PGFktoF0wBhyUUdeScH/Gw5dejpcYyA50Nr2RLr
0YYlIYq0E249V9eNc57vl+US2GyJcQrxN9bEaAXg+mhxFi4FhSwdah62xo5/CKV2L633n6mWlR1w
tPRlmY9Hxsq5det1MRmKvzoiL2xxLJ8pKwtMAzI9r24XgOMplE2g5wb59hhnsD2lyELWzOiQtam4
iVDfrARzJl8XV2n1hQtfMcFa/edvwNVC8wcFHf8uD8arAJ2ktFPJShyGbjCSSsgwzBqQBmGe91YC
Ruq8hejJKNFPr3TKQoB4UH6D9j1HqPbl/bo4KLiSKLDTQ2zgnlIdG6EONJGg2TSWLS6X5s7lrVt4
qIM2qqahKZgEOvWocPW3tvspEgwQjCHy5iX99QwcjIjwt6WDJLcL4VRX/Zzim8t+yMeC5ZzUEzQj
NnvQlJyEjmHHYmbxHVz1bk+P3sK9BKfoG5zCnAio1dGQrIyJfqcLUeVXdXjQi+mdKBpz8M23NYuO
icIu4oTvk9fxmWx3Wz0NOI4Eqy7dMIY2aXUjaMmeoOQnWLrw1ZypVGqyr0nnVnSlvqhtxap4DeVL
JY5Sk3B1wOjXLz4ZStH7+mkNwxJZmyLw0+yu1Lz7ifcZgI7FcG7HOwnUSjgvCg6hUriofAj2aUy3
CtgKzd3wBwQ39IqKOLevT4S9CSK0EyRaZg0CG8O+5yV+8zgg/SHjAjJy/Rjkcn5Rkby8yZHQKC1v
XBDitd99P0x8UaUzm/7rsA2/GhrAYchIcL8ofq+nCgHVVVTtj3Clb3nnhx0bOyEhNwSXwhI2fvER
0tKuV7kXXFPcYwppNS8HfDC15Aq68MAfCe4MZjR7dnmnq/M8+ciPVs3lRE4MToRQCiGu4lGnFwtX
iJjjV5lyWxTkR/xdOmOPStepEYeDJB+ZkaqCEkik8CYgsCurFw+ZV2KTH9hmwJtuvN1Fif2W9OTe
UwGFyZ7ahnWFd2r0ENvwx+b9oUiAtHyxemGTvw9EsVGZHNB8x5kDwjSla2RaxCHIQMP/qRHdaIfs
56ySvr5T2i+knbuwSTYgyrj1QJBpeJLLHVF0R9uP7BnpJExLfD8APeI1eMR+W7gKuwaEahE4A3wi
amk+JBavvqmRsgHVEPK2yiRdW88DGpEYOR0PXKSg3aD4dhgG6h/+1L/O2BeAqt/NA3HS8NNeBFR8
DcJuZ5N7YBy2dy8kHwEas+uFUjESL0IEHozRJor7mGNq5Awv2jmxuKDHHESapvZsAeL11xyGa+MW
ruu8M65KWRofVQHCoi10ZDAnHOUnsK/ygH/rVhBD305IXOhLGjF+RUsLe0U7rQ6sE8RvhzG4hVPS
pdDrtyb+csXgZyL2Hc5mW5ypFDpGo258LYx+RYSlOPIRkC1x4OFStAcwI5l4zaoz55Gb4g4F0zQ9
pVWQZ/b0NqB82HIqWNCsC9reLHtedgss71IDN9dkqJmc9r5OLQuefvAwk1dBlnNXNoFE7ozFkyG0
ejkMPbDrbLloQjHgGOEAWDHs8fsAhNIq0v3csIg+UNxRaadJmjc88DH+Mq8ssAurfJ59ALuNkutD
vAtWCl6OX15ArH2HPhu+ZxdxyVr3LgtZeo8VxMgve0QdnMKDX1Jt5qDU7jG/65jc9P5qOfHSKzra
eKXYiImcFKslNsPCmUFBZry+X1X7/XDXgfxnGhjWdOzHaFj+sa47yQfgWf6Td1TLv7UtVPU9bhEj
nBjSaeVGLBGevk5oBbCeIz7GTH8Zknjizp3J1O767+S5tJVvM1jJWn131KrGLQMQMO57rkFKCopB
xKtPl039FDoutP808Yra/Xpw9rRRs3tWLHVghqOJ6wAMeaxIXvGc3qI5pCb1CeUxYa3OPJsPwlnc
ffV7gTP9dAcmVuxY4L9AYNmzlR0try1xIrtLaEudROvboOD9q2Q/PBSk3H66gB/NqDG/Y8JyAtqn
+GwHYCuepk91qebCG8jSQAua8nxb8+d3lY50Y7CF6vTITEo6XUdIJTu+wj+/AYoJ4K0IavgQbeq/
hPAUBPJ5mfGOxiX5P/MJWSJvQnA+eHx1OcnXYgagjQwSTrjeHNNj582vDsjSrznjeCMIVp8Xz419
HKRgTu6UmEzpPQvROz/QbOFBAlS0//BV2X+xCBcvq7UeJfxTqBhwxipACf2PDjhuinWhQ0BuBmsZ
oN0le3ilRhDhio9Zzf8h2iwPLY9v6mUtIN8PdiM3QxFLAhUoOVFnASytxslQouHAKQUBO9b0+neb
UJGVNHtJES6UF6u7vPxrmnFo06GveXH7RuohodSu3dCEZ09BNEs3hATZsQf8l7NfoBk/gIjPZad3
YdZmE3SRH8bJSoyMy1hr+7bX/TWcKSZCTpuXQJrrdRbsFOeu9mJXf7lxF+5FIDcMOPI+pKBLQHDX
9J2N/RnTlB48fYk8kvdvoziDVMbR0R2yLXTIj/6MD0qxegyX6OwM2eAToWHu2RhS12TgjZTFHh2u
NObtMaUIDIprPAA8wUDrHAvChPkxputIh0dnsI9a1+Cf8I1Sk2keC7IbleRICT1JGZgrubZfJHrV
QEo0haaq6NpVFHqaDuUg8OG6yNMafWG73ItwSSHGBT9K9NnLnTPM7gVR/h0rnjmfLuTwmZkJXIOJ
OMiBCi462gkOzqC8PRMx1eXbvrmMTeHt0blT/vSc/i7TRSjzBBKgl2xVdrpEYz1PixO+fTIBXiqX
U/hOk5jF8ZbRxPsLpcL/WeZVSgGebWHY1oTpoZvW2xJmVy/pDwPN4AJKE49rqycxh+u3xm3RZTjP
3HwUxR6RbBZV9L6r+xh2+YUZTNbCroTJ5raJjQqXB2C03Efu3SG0N8ZlOpY12rHWFyncpGoyfduk
JA9R8qQvEUkU42rNzSiVLyl2OdpxvQEbEv2t+812Bq+pG/IuYMjz5Fu81Voxxi4DZ6mWzN+GxJAM
y4lP3mJABAd+lrRlzs176VSeCAyRHtZtHCqRqDvIVxoyfUwmZtrPvRgHa8e1TseNe8nIqdfaGsEB
YygQaE6l9eUeSA6JYRZqXbwAxKM18g4tjzHgA2+Waad4bS5XjVsvgwTg3dQXTwY2MXHFrKuQ/Yc9
HB7va6FmllIicu2s9fO6tvH9rfOGMydOt1af5b0Zad25n3DaaBXjMh3IHU3kRbCLDCi7eKrEKDxq
yuCDTLgGv4Zu1CTvhWRMWlIwWkYA+rfW6k2NDxQiJRh6aJUo9n3dIaDcsZRoP6Cnu+qfiwN3sCdG
E+gU1kjj/a9upWk+Mlp2PfNB2bOZLixopQ9EX8ofXjF+NWZBIRaB5EFcf9MYrz0A8i3/3V9fLs6O
Yq09oaw/wHvTfQ8uzHcytsxsAQYBtTlEfgntkkjgdBlyq4T7DI7xFVN9XIJ76kDXnX08/hxQCbzj
7NC/2vSqUrDNUAznSyWff9C7tvW4xDx+0mBGX2PIKmrwDoNUhlB9wEjmBXVICv3K8hsGg3V+g7ve
3GWL9nrcelKJi/XxgHiMOwLwnSabMi0YzfqKgej2IVTEEfmwdlsXnM2Tm+tGedEOFjv/qveRNKhh
jxc2RYf99+ZIMJ6QAEtDyzhZ13wiwEMfLiSAgRUgbp+CwSxwwPQiK0OsOBdgUfzsU6KxcgmRAExm
0LD/23EHdh/QWo7h7XpVAocLOlOtn572zxiVEokNNi3kxs412DFRhf8TuBLZy/fwBYUFs83pUVQr
XtE417eaSuuBmlFzZ84/xAgIDWbxoNIHJCmn1DZXEX4c7fp22G45tPtA0pV3nGzk3ZoPvCqi18vJ
lv9wQNCMJCYVlVZhLA5xwQW7F3TMBH7nExdB/fGrVYL/ETiJJtL3n6z7vGWCfTcm9ggbfHO9aJfY
yUX5GqwyIR02ysG2WasbirX+7alXIhgaX/dORNCQG77+RE1R5qVMm5GW7BLrVOv0tlHkrfhckfEz
KY+iUb9PuRoP0XRJDRr3WLr5EFGnBLwC4QZgIWqCORCmei3sARaxisnq1ug3OeFwrW/0TR73zBaX
9lEIXk2kislG+B2r7kispCOQfgBeTkJX+mMxGxufwqyFD2CPIt2noEWcVj6VJ+QQF6dHqouOnc0N
28O4/e9OyQxvfOxYF/6rXVCUOOpV2ZsU37h/5iLRDg8wlrzpx8GEzlMWmiGuvvrNxmTyMzjCKBPx
Mua3qJArAmPUfsaB2d08raF0qnzR7JfqJljC95tVPFkspq2+0kBbI67GcyrMybunAYr7MIEPMVSw
ItvEj4FYkGrofWSlamcBEB3hIoUN0eFd8uTwrFMyg4h6Or6nTdG//73Df5ttxOy1AXs0lGgNIDLr
ciszKhJl3g0sCLxyDBTX0IOS3eg7X5koUWM5RpXdUn9fJhHeztzgD69vu20uUm2wEegmLoxuxsfD
VW62JBdfg++nARD0zDSqo5OXNYZzZku497TgxZ3hoZTPJ8RLEEXkAPETB2cIK6oCVw4kwzdE+Er5
yv+GGR5C+fZD+tj5zLIvOLhr9cLVAoNotNlV/yrzL2Veo4mfIugUq7XuWECX2UIbayxqXaJJCnAX
KImq72IE36V05ld2VeqorPpg+t0EWENHlzFvckbrfhXK6s2dNe1AB8kZ++23YBR5GbDq7YKBxCS4
9CgwmFgjixhZ/+YKuJhmRTshiqDdQN5Uu0u5cwXEVmtuWorQgK9sL6FW+cH9I+ewHYgJMizBa0Ou
TCzUjq9dI5HplGH79AszWaD397nHZ8jHmzKbGizZIVGVHNm2ymEVSp4+VArnOx+GugueisFjcp1s
B3gGa8uPsZtHuIpD4SRc8pyhnKQ2rnn+QmeVcQpLQqyjpUOBCh+SY1TanP6HO31FkdUKupBuvAYy
EClPeReLzIs3t0692KaJkeSlu+WPum8hvgCDu1TRlWJ3lpNJobMAHiZFXXD/Z9OsjwzCq/Usxiim
6wSIfnPcTvSvtDLgHSl9v8Z7cftojIDmvX8vRo/qTJeqFioRG3ONN6lYRjQIAEQ/LkmeTqES9vrx
fnP5+rAx56/NKysnBSh0h+/7yywZfW8Ckrz6E5CNP4hs/8vCdpEHZSF/3ox5FZTzzpecWHnSRQUm
T2qwJa8CpTe3egD/3XoqChVbzeaqiaXw25bPovMwBAhcA8LGVFfWIk17Awq9ECfEAlIaenfr2tdo
CNGWEKw9mU6kFULtLmXKtOHFvIQfM3f+Jztgd0ShVCN9OiR9vzieRgT2JujoDWHU7x6xh/bgSHmE
V7QIkwabJyoX9k09WGfj9q0k9+6OiXWfTuoUezYOHt+rP5aMUjvew4FEgFkAyp+BnZ2THaNarfBg
OgMvV7SbchUrvxMQ6NyB3iYHtO18emH4wrVgmIgPFECQYpDKdyoFqWx2FNH0RPM/1xaApXuVvoNU
jip+DH6eZElavt/YOzr0g64PcRtR9cWERc4SrieTGhd4/D95dOlv1RTato8fXnzdryMxwC6psRqT
NMwyMXsL6ppUZjLgamW3fDqlnwdowYkRI/6Wgxf6X5NUMxlJNvYQT8vlj1reyiLioQHJw2YV7elE
C10eJPcWl48WnzxN7dRYO8nZHFYcnsuCynnWxmXyqZEXxhji/hjCdByZZL401yDqR5+F4PQzrWgq
v42RvLIRItTg90dTZSosQ98l0fRbsbSvz+cPX4jQDiQTrGhvnIR3ZmZ/zrN4A5WeutLA0aPfS8ad
KMtwJIOUTT23akKFyBFI8kVZXgNxl1oVZdawsd/vfs0t+a7fHaDagdkuAOIu5deuOs+MrLN3hug8
fVhEO4ZIAlL6U4N5lC/Sgka79ZOCvwjEMukKsYbg9ulJZruW8vcyH1jHYzsM1rmbYL0unyDiMsaL
MD5rkV1glj1qGdfVD36e55GC3mLgCCJaadyDuEfe4DQAqWEIsBROC4R0pjCxoAeGlNUhvii8Gxc0
XiBlm8NgjyCY6hteP1mUJRWlzuW+tmQMUcfM6lhxNx2mfTs4R3s3h4QO9kJac+XdPpQGCd667vJC
jruv0v07sSSrK2PA9mlSyNp9Y141Cy5k+4XzQfgRI9pzPiglLbPyzPb+FxP7ntyLGkw1z0958WVr
yIkCxRaA7TFJelKhYSX15cUi4HMtkzHihQVOBmUsJmuMLmad+u9IM38XMx76SsDwLxDeM3Xzjmt0
powuMdATnxlQwF1ZCytS+elr3Pkqn4roZnUE8UtNW4vNDL+yQp40R5HgfK5E0BT7hQTIEQeclW1N
X4emRG+fTWmVyaDuqOMK4yZg6TCv5BBr/gPAe9WZGLjXQ3KDJWFc0Xt7dntEnjO10gMkv80P2dw5
5ThRSlD+Q1DWWlVtNRoSMDH7pLd1rW5k1SGG8LTPcRSMQasFQ/m9qE+E8yFRIv0z84zl03NKpQQA
zLb2FIcoawA0++Ttiu7hnucqKpLZSYtGG+ADGg7mokvDY2h2/KKpw4KhCa5q/HkGd2477WDu3ewo
a8hayJSgXeJSSlZjSsayVUj9FiOSehXBpZ/+hC1ftblHlfP+0HqwfpZzqSnbvVR6xLHz9QTQ4b4t
7zXlF/H3jEaFoSjVf0sxLcQuUUcjGeNUKUJiIegk8WwCNivg4Puu4K40MYVAQG54FMqli8d1P2nL
tI3BkQq63LwyO1KTtaHWRVokKRRuwzypzTCWgCa/AsGdq9UJwFYXuAWlTyTJ4/Hzwuuh/us47tw0
UOBw5OHttzAUvnEd7VkiN2KdP4sglGV2y5kUDZzlb8FJdhNQFkXlQTsa7IBd2mJz5mQ1gvl2phyy
wvnYdzkxC+AAvrRywFccbSKvUvYp7HjxP5w34RVV0iYAV1hHfq6tc1QYQKoPtg9CXFZycq2b1Fat
Q0AEanVoPXrT2KwQRV2DDqKzYoEVJjbsvqWfpTJD0H5CwrDtjqo66Zsv0Yw2ik9jYOMhtROJCJMB
FWaRpXFuQjx3XYa6b5Tk91Md9xz6/iW/XTrglVgyNPbuTlmiQlPGUh49uArMLjXP3Y53odSRt6rB
UVZkiMOLdPCl453Zv2OyHiPIHSXLYcrALlo7hrj/FBCX0kQ6NxfTb6vn+mb7TgYEIeF3HKzkXDvc
xggSP074k15y0VO703VtMEiB02lItsHUUpQLsrmUUc0vlmwOoyFEJ4S8i5Fx2pP6PiPkhV2p8hpA
zXT+q+H+9+DB8tLxEoLBKDwbUkSfEANdw81OxtoZh6M6DeExhWDd57LgMvPYLRxOh5s6FR5aA472
bNwTQy7H3Eewzw3flRGitTmi6JpWMwS8SeLO6479/dFq1TFvgrIZY57YwaRgs7zsx1mlzwTzsi0B
3FeokIXvNEdT6ZlHFPJNRDJKvkLcqW0e2Fb5z+ADWqkpnA3m3A+BvEPGML6dQnv8xx4nQD1QzV4m
tQ8lyzMlLjN4q/hUFvKVoPq7XySUgcLaIrEZIw49M6ejF1zgulC00i+6WE3WsfRHxntkpAbGz+lx
fbDlm9EymgUVTH7fGaIyRftGI7tHQUsXzcsXPhCUNaT6Cr85LaZv1eJAnJFTyboDiIiD2B7Ixxkz
wk+c75XxyzPdP1qZJbOhoyMbfdnLQuZ/AIHUGw5/fBJU02+/SQgUpuIITNTl7v6xHw7RxjYtMwYB
7cRNnMnnia85oz1B1BKXilcMVK8j1mmENLdEPRELImitbZOrZicN+NKHGrJUBzEur1MS+iaziIN8
EYOJPbeYOQIHZ4gbTfSk99U0EJmeCim5hnQpxQlnIfjp9OV7tIfVPsGrI+YD/Jc7WrFej4cw+Uhl
4xPB7W0GMoZI/lYZNKHETIvmKXShVjDVbNTaJQUwvfd0IQpnIFzv5RZM4bUN0Ra30t+p5uAugLh5
6tkLCVipT2KPoJkWQgkwUagfkFmbv05U2LHWSmWprj0DtkTsmlHDWeRg83KCAnHs9VQOqcK+WTqK
RsRIX23dPzr3G9lEAN3eAzO8Zv6/jVi2VcdEIa9Ui+t3IXyEb31GpUJ6EbU3K/Aozvw0ExVdAD7p
ZB8ySJzc+KzEEfde+TLsuTECZlmgcArqG+CdjG9rxP8Rv3jqvnODKB1N9founRswNPAWtWgJKmeh
UZ8yNyJHmkqjmQNHlGokoOCfwuUjkN5Mb4FJ3sZ1cVapX7yWhQH0ho29RvURaTFzlfZ12RW/wuIU
MTRMao5wiOSmtv4ZIQ3MVuY9DFtq8NhF5pKxk4KYh6meIYwFDMDXsXmmyHEvZV7X3cd0ghWbaTSS
fxW3LcJTaAOyFxGW+qdWSgfPFAYobHl7N7gc4feGO9A/yeqkHRyjmHL4IGfUuGpbqa77qYtH5/u8
JPZXIZuC7rIevd7OamVOj8yqrFRDJkYWTAXyilOkF4kchvWnIwHZlJSQn1G7BMp0tWoMN9/UfW1r
ZTpJ24ip+GiJJaCD3mnCnhxS3Y1jpkbgSxy/IkyGMmgHZuM0UXm0Qx4RbMl9TTRmfTTj1fMrm59V
0JIAUdRrhJ5CCTrGOm3OolK82Me+7t+A4MmlGbPqG0TZzmujW4X984hSGYTO1icqFfsdkyVVg6hQ
j80yEgRSPfe20aRZ81LLH0Znkl9C7XGyBMRFhHfuG1TUwbQACo4oEjQjSJtKziSQvgrkx/VkvPAr
/GUiV/H4mzbClM49mDC/wkM8cwJfGViQdawoyjayGwcTw6hQXTVW2zOz+/IOT9sNyQgy6bS3OPOq
LPmhk91UYMSR5m4pIZZnlXtqIDAK9z15h3FED5FEa/+uOmHJI+BZJfJgKMHXYDUG7l/gcIOWOVVm
rWuz14cGPZJdDxlCSU9+Nfn83TYDus03Aq3MO2C87KPfL7JX+f3VBlCVMPu59TXDPcZEES+6uO/7
lqE1xvWF0V+vdHajgIJFZ3BcGS9IxeSX1nYCEmQwLBv1XqAX0C0ItM9mTLJStx7JB2iL65orjuLq
KcWoiZNmnItrGXb6W96b/0596+5cORVsbk8mLQCry2nIYL5D3P1VfzTcin19nktxreZytmxSN4yN
MZ9cfJwPqVzd3wuWcPD8Uog3RYH7agnsWx2AQWRgKhQeyEgbd+oCJfkRTobdM8AbSpSXP3lNPGWO
kyRA6WjHlyDji8jUV81y0MxGhxRHmRZgU4pM9dBNzQI8e780BlxoJ+WS530rz9AYbPsLcN1vVmNJ
T6j2WJ+hSbun+gPxRyuwxqm62Q5/D9wjCMX7wZhEFoUxSjuR5jGhZZyuwAlHEZWnokt8zqYtJGKG
j2/wsVVq4W623XqPDdCFn6j/dOT6P3qNbW5DfPaQiW4MI/LFJ5eB2hQ2BjmwaOAuCBXZQczXId2x
GCCeB+hBAsqjiTL4jwkGrCRoLfJCG5tDBpWmF1jBvzVU532l9XGueAOkDDZjIKNN2j8Z3sqNs2Uf
i/3dgyCIe9YpGVzXeYI+Wp1i8jyUihyxDrKwj4rf9tC5N43zrQty025xsT6WTI5NLXmIa/PC/z7Q
nol+JCmiPMJJR9v3/fWTl4WMyIPToWuCrtbP9+6MpvZcbJ0MxZC1VIpGY3SXnr9XBmk1rc4cRd+m
sotshnQA5vAKu59Z++S2qgVd+ZTKTDZ1g92ChrlSnzk1hTe7byYzcTSlWLQqKoUJ2u6scTuRIXs9
eNJN3r4jcWVsB9ymXdJkf4QE62RVnXAgmD197PMxuvx3HAxzfEA48b9LMzks7mJ2AQUVe9LSyufb
CiXjA/ByTUikEv0CqE3sQDIDJarhU+VWEpHD7IAQrWDBIEIJ+wTHAHWB7a8TGTpV101w7ivFpBJH
UbgqGw3VzDEVX7NPz9Gt/QLAvhuwFgXvt5INKpm+HIWZ8ABf6IK/olYhQLcH1Lkv26SjfxLtW3gJ
qJs5Uznz8wRuj6tr5oZpWKHgPbwbLNxu59zh2PFIC6nsWU5MAu4L/DsejzaXiffpI6VhSp3yVTax
pvXu3hJpjqgzxZaLHNzUNGQmQFdVuLoWbHH1t6YqMSdolzFLoSL/FNF+wI5xPm+1l6oFPbFgGjUb
V3+53oYvTOml76JzmJz7p7Am5siOluQSLfj3ztIlIxjjzaai3Qnk+VffzAR344NkEgw6SEVwjwn3
8SQg8KYoo18ktX8YPnkzFHmsvuCQYeKP0pbktWsaVubzr5ltBdVOHpqsAqvTNmnVfeZ9ccGvQe1T
5KYLBuj+LHvnkkcqo+LQ8ITLGksqTJDbtu7VVcUkJReQp+lf9HEGtt9Iad1B6LlzNCGKfQdrDtmQ
G/3WkQcG4XrQRcoBkd4jJ1GECq12cKv+OD+lsZRcRC9HRRUMPpf6N3880aX7G6bnpxJL5Vqi9M20
wbo+maFODTmEnFYu0buR46bc8led1adWPskL92A7/fD5YZ+hixZf0y+906HwB4FWkYXVd/rEMAWB
5PSi9d4pw+sZd0UTwH3Ar8YXAta9CSSkXrUysf6+OZnd845ieV9BelliKIt/lImPFEFtwPZZEa9C
pGg+XdjNfWgzWdWPx3QjjZ0iaRWruFxhvtDpGdAVf8ALMwAgpqWKtX3y0+whb0aCXU+t+rmJw7io
r6JKxKlAANzVH0sI6w1MLyO0gabnMzEKXoBRqQEwk9MAnSE2bsoDa9pspCPHqjZag0oWtqzD8+kt
v7mg0aqOCunkNRHE5BGp9Pys4MTXHY8lmySeDkaEq7kAVx7UIiGDPVovdePFtn93fgALIxEEQQIw
TPWSrUnRZ/mP4S/1WNeFASmIX7DoOg43tUQjQxxrGrfw1w0GJpv2EvDWBCcBAfnFcT07x9HnyPOl
8ZdGgeEJdjKGjVqBp5FzAo/gDg3vKt/d3mr3hE4VMi9G3ZYpe9mTuPo2H3U7uLZflbYFLQJ0u+pQ
Ik8oE7jsus5cwAyDhicWFdjdu4QHOd20zxTdQDi1jnyIdW5w5gLZwtrusk5yBYlbuhYkXbImrUJc
1+xlO95IdRdEOeaA6hNEs2EPCGN9mbCmeWDpEHkdtq2oJRiLLXyzxYfVxx+Hzn6+c7S1f2+MoxWe
QAzD6PCwPoegE6b4sBrLkafwF5Yy1a0KzTvtmnxDl+767Yo9Xci2RqkZrnduca8xfNgmvAtXUbuR
bGZRvSHzNTJav35dj+fghhuGcwXVAHu4sp37XgTpE+5diR4YgVp8+Ol98OAMgYN18aOlD076a3tz
5CjcQRUZAfOnSPBu0sqzZlR5ChZ6KK4m34wKhWlG18snb32wlpQJBlU5FU+aYl20h3CiCYp87BrO
eENQ6jZXPYcWl6Oqa2Dc2+RII3UujyNGJL7CWAt6la8w912tjqlc10v16F/n5oVHMefDoISDir1S
WUfBqRJTp6rLlnPMNAxQBWB/vGorHxM62pFusWmS8scJyfmumnWVg6pnuc0xv6fjsg9+Ew1zgjqY
wQvK1fwvUN2iBI3wsbCeN4JQlpKOyqVj4zE7EVMZ1ZqS7yqmpmvVSLMwQdRRYAu+aLaXflZP9AwQ
Ct7P2ciOox0Brfpso+P3P69RyOySsoU3apcegz2o6/18acM+dMhhrdBvYwalFVEFHbFKLM8cSiYr
LEEb/RDw4K/R/cizebCdAPv1+z4zDfp1oNwJ3jhlsyGeTyoADLSmW1b+PFaWwsSR7DoWx/vNcfuO
PEcWefiN9kt1GKHwvfS9fZqn8BwpfMfJv1CV5IHMjbznkZBngkq7ne2pumOIx8Q0o3slccpSeXJP
p6pVYnAk3LTjXgGdGJX5fEZEm10IV1s8WAlHD6T5D8G5dXtZE5q0Mm9cOB+GJwyp50uOacWIb1Bp
vZDg6mC9zPfdNJXQrXdZX/XldP5fxatEKmA9pqspkWDdaxrxwrbZsDyttNyVf1+CNQstfpx7zP+W
qWt9uvwh4f7eXjC3VDA7A8xlYsi30R1tb4/G4FqTmo/Uxlh9+EPdkB7VLxKLzn711U2puL1CD53W
Yv7AAQel8TdsTxCmBLHxuaPVEHQ9igL2uBpI/VJIVpT6nX3Gdvf22wf0nD2QqydqZ7lYfie/N2FZ
MCsw+JbuLjMu6r58/+biHe+0oABPQD8Um3cLrRAO1T5Duu8fPod1sois8R8vSgQAMQesm2nIrdkA
aZALI0LiVR3T5oMaS6J/ohUwfbYa0CQhcnJZcmlnVHsQbLZo35Ve79plWqoeui9ewLld3oyAfvVH
oRphHRAcLpUQEF0zhMjv96F+zgzLVjdz3bw4/aQqmBEsmQlrxNRlP8sRkLbWMY/qRSCjmYP4XXWC
qO+DBhU6FbRfMHj5LGjpcvAqs+ZdW6S8xENV2iWzjFeaCZnYkAlHWrrY17d11chwQPPRvmX63K5A
JgpXrOsJU4LnZzxzjlUERyCzl6aElFVIji5bUG7+JdjmXRCnEMpHDZQOwQruyaxsVriuOuen4s2x
uxjwTXvs11xKzAKxFyNhuYm4K/NQgBJHZ61kGutTZ2IIOeHJ7z8j1QZI8ZsytBeK+CleVgp3rDjF
wVbaZFSdtZRSWytREHIplgDUvjKU8qZXT+703EvDonww8PAivo7RvhVdrhrpr1VCr4nIp8p/ztP5
TsLrrWCNFTkU2GkrVOUqIsXVMxJXtAgXEzZiYc8JpVgwNPgrOm1j9nnWk5ekcwVas1BYdiZQLWjO
kbQNSv6roi3j1Fs4Y9XTCG2Fd7ACGVfZNpzbFyD/ouW94FVZz+lQ6CVVqdu1VmKqV0zSoOY4clt0
maipIZDu1JLyiD8UskninlgD1T4SFMRs/iW7jMY6jsnisQcfm06aOiHFYRdNDWyN1sdCbbkiPJsE
d9X+w8TiurlyGo3AGPYuzz10smoqv4W+VGJzXBLDT+g8MQICjz7pD9BNOctiwoq1CmDd71NZfcUD
aENX/j9CFWuZHgmkULuYe+qC6s3KoQq9P9ZpTGtXlkwhf/U/HijpDTruoSlQ2Q31eS/O9sKQLxdy
h2pO8MgzCjVYevIqTdmFl+0NWZXANu+GYQjYEabGW9z7fz4PyJfAXp2whpDgmYWI3+sBF7nPn1pG
MNSsNpYxPxADjW6re4vTVcPzSrvhDh3yZ1jpSpIsKeEOm30psfgCkYyr0Gs+JjZ5ploe2yCiCyGo
qYNXrJjL61qMptfylEnuZq2vDy4Z0VeEUVYUW0rXjv0UiDVPgXxMv/KZ6KcHkXiebJ2l0oFtm+O1
tLQ8PjyilBh3h9o/RL3m+lrvVbWjsbaC5LMS7fMKFZIi8MjCOVM30w8TuHLD7T3uj3I9jOGouQea
Mgg2jwrTz99QOOoysg12q6wgII8NJjAZ2biqqO7XGpJ9Ag5zT5bF5V/eJ83KhXheTpYMrRBPACvW
4/D/sP70YeLyLeiclUD7MZwK3BpYDkp9snAgkSHOxpbvhoWuJgECLiTTZk5dZ23OKOLHDk49AmxS
MJtQuzIsxj0GhF4ayJJnz3ybOt+RSi+FT+vPXhcsCYHnDYEN+35uiZH5xhkSFulUhzSKTHubEjoP
PH+clIZoMKUFxP3ISMgsQQ1MIlZSSe1fpNXp9jaGVj9l563T80bS6xgSJMhHFDfKLv9qWSyt+AVE
Vl9yFjoa3axpFkQ/E60YW9BoUQPs26xp447/jo1EKBt9C0NzxGf9IIun4+zO+XF7qHU+QmLhnppq
6DNT0nzhhfz4O9iJcAc1gz7K05OJvzAAwvD2SXvA2QKfnz6m9Zv26QLh5BrRJdJKB/0CBif4ARan
J04qsej1sRBAfXYvs+XBme5IMlQ6PHOdWqY6jo9nxnuBmHLKoLmiRnXlyOZ5uKjv1GOFKHl3YiYG
IqTf25m7B4xnPADCYa5ExE09K4mCD4ZumpmqEmeuwCub1YJTmXhnHriBUJslJ7Jb2z5xs1DAzotd
RzsT7KQL88J2xDJ5E6aJlWxNVUA+acKV2CayXejHNYIGnlalxIQrOoBl6VAowkJsc+5b4JrTTgEQ
Q0tAd8UOwbBlTem5iql/R1Igvui1n2WL7cMGf1OSD8Z7diBYuVgumUhPhIWFKzN8wT5wlKY4+rWE
+MrNR3d3Zz/6BEHstnD8suWWr+H9fSl3rsvzLvRgBlGNd0WX4+FnNpoQkrHKJxAbbqaAQ5nRecSx
Z8tGrdU0gvh5+c4a7qxqw+f9eqNbk7nnFAbvUGlU7+LeaagjyAwIVFWa7/ZKlunvfRxH+pb+UwSM
eh/4IbJCGP7REtnLmdLp7xhpWfaiLIYI26XSXDq5VtVH1taKUNtvAPGOcDP0EIKqfPgwo1py9Hlh
T1CBIrZhxcNEwL+jOpIfRPuHfKwf6JM3N8EkAHIyld+C1icfzlg4WKsUhQk2MpVeysat6bgB0Vrs
8pC+eNMp694yMPZqTzALd+eAOYF6wAQRsO1VcOPHsxqOWNQd+vx4g/X0oUrw7DkxuMqio2PG03i7
OF8JKy/QmCP5w3IVckdcNVFNEs3kgfBIzdp1GHxMqZUA4Jupyx8X0hItfh4pMEjFihlZLK0dfZk5
el6M7+S7g8G6wW7VViZ89AIj6sM8zHNVCPMr7BGu2LlnRjgqzungRPsrhiJQVMP3kHOVF/eb4iVB
g3Rmb5r0owft4wpZOdxbPYXhDVSm8B+YH4hjo1hmdBw16eEDTb7BF8iAnIF9ATOS7u5ewGxS8+SP
3PLACyJFD273CSXng9VcfYkD+t17RxxYqMpsAxGJSWo6wPB9HQ+8VZ2XuSxVaa0qtecEwE8ES+9I
gaHb3/2eaxra+KzjU1h3/YFi6prXp6o/EPdyQQlnVIedZeDWozK6y9jpUR+Y+PDN8Jvs7n5krqIH
dBxyn68DyeI3NkZUFud2iyhVQ7T4c3dX8UWnWvfw6RXBtonm7ys1t9lrQ6wPIQMGVW2k7UHzjqHn
4XOTWSpI8ETGYJuuhiVxe0pUlTaDn3Gsj/5bXy5sCsqXZ/Xad5DAtyEKqxXpW/NBdWccBEb6UqOH
TBfShU8kEOyVw+hIW6T9dl5WT8rHvtxy81CuxoE/k+kfygFgLcVd39c7e22XSC2FDliFLqWAut1m
gDE1XB88pAQe0z9NgPthZxYmfMBQ8TScKS7p4NhTJMIsbAnIMiHlXB98soyXM+ChZLvU8T5inPxs
WJA90wvYWoM+YWB2GN7L9bQSjarSWx48hLFKD0D7+KGQv2eKZhbONMeKr+E6LAO+buLLwU/Sleo3
zEwUUBHk5dbAS5VZPOiXindgmkU1DAa/P9HCOu6LjTLZ+S+VvoaYnGcnD/3WVkZkjLan9SnMsgyQ
PSLnzHJV9Ui6Nu7pokvd13+A/6BumtF541/i5/q0R65u293wxmgpPMCNMBWnVXl0gNknqlwwADpE
UquaABWuEOmpoVPbPvv/12wMWgttzit2fxOeyTD5jSsZlZol4WwVzeg/YtuQpWd+qT+sWw9H4ovc
yErqMnh7POh1iUhwrq2+5jCwR9dK7aEfuu6ltrXgYvBNSJ0iBoHf7v7rSwYEGQZYi6ydMtZN4pyW
hngs7I39yA6C6/h0LUP0FlpQGcu4b5pr6uZGPbnYzdr0Q8Oabz6APDSH0nT7zl+HXafyU6Ep4moP
wjOt1wLkT5jusOa6C1O5sxOUaCo71tjFRicbrSD8YTUat82WpMC6R22lS8R5qIIj9lWfNhQNLQ64
UEi3zL1N1mDIfkt4dgYzSixryczxZcg8RGvEtKsZ6sF2epUaj49znQYgakyalwQVMK3ynQxJRUWg
cPhekrehs/vlNd49g5Q/IJAGLMuCQetHCzX4YBNEBoeoDyIAoUF0oKpIbofk/0Fa+j3rwICgNlEH
xft9cCdkdyLzfVbR8JgVwPrjvUfLu9jVtRapyJf2gr9VWK4Ygiqd93yLKyEIKD+NhKElAvWz/RPy
EyWgxtjjBjLefPHGQwvKM8NVaWx2GGrfRwrk8pUCpoZB/4K+wyduHX/mAV/3GT7BEcFqztT6DtP5
grxK83U00paUS73B0BHipicip91wHR4TvotSLM4wXop0fy0O6PI1Xdd//Hm78+am4vK/j5o53Z8k
Goub1mpntLLLRew44TC8TgytKAAhT8+2UmAyMP4+hsFJbXj4V2iXHjLQVvAQ3SMuH+OHfKi6E/D0
3i+I3OBF/OE9sjIH9WcMJaEWRgACxNW9JWnlRacmy6Ysz9TPJWa8WvJT3lDPtPkPIvSiGMXdm3tn
m0jUxysstlCQOdWg5bYb1X6SU/wOZw9t4a5MZIRw4KSoWVYMm5qS85FhSPQujkQ/L6XihAt9nXUc
B3iE1a4ednL6oEdvCixyFPTqAi0bpwUN580w4FJFzhAT2m5OaPgqEMthN5qjQ89k+94jDfowCVKY
8QSGcUq+7gD1psMVfWFcSelJv+mawb7FIa5sCwap3Ub0PSrWG8BpJtEfZsMAXWDvwjbeiaDK03/q
2PHFqc5rNPP6EgT4QEKNmPC2SgF1mtTpH4/+ZU8wWdfycMTmPoF5m4hugnNNb7k8FhlrdGYPc3Aq
mcplEc4wTeC/TdKMO7nJ4jL6DbOmesjxafsLDVCoea6L6LxcjUIRQqg8ziFZ1De81dQcajwkXbB8
jpI68HqDtHloTml0K8U5CRyyTTW6UQYGtE6ZCh3hzqOWDNdcTM5Rju0fGNGPEbGpSJor95a+JYVd
dZiVCqgEYyxuSavR0BitfAqT5EwTAwQujHsKoofanhMe+Ij/t3quKfGDSB/AIjy2S02uV21YxVvg
jGcsRUohvBOLK93y7OC8nK3+hHjLGTWA/tvy7nLTJBm4rSmoJ6CmMjQGUYl+19T3q1UYfpAehviB
gCBXg4kiqf2h+Hkp5x9DMW5PGps7KVKdXnwnOWD6olEHDoCGWwr08xXWxwALFt/yARLHYK+lrKhe
5ejKtSaaj1TspVIDu1Eq/ZKQBypXUsnLmpZYq7uHm+BqKjFAmKz4fgsyhqzBjPbixPxMhcDueWTp
lRP0bLow3/xaCSfT0qv/JXEoAF2MSN8/FYs7ibLUEMnfnBJu8npYb8WP+afMPoopwYytHHacw82K
F/+qT2NxM3hzOOxl6Qw8G+D5ZUkS8+hJQOHFXmuqKgPOjVJzeTqvc1o0S80dFP298LtC0cBHjqU+
hwdfjFzXPT718t09vXn0+TXUitY6vQ9oByh41YKTZWmMa+tdWJsItsYHgOxiEeRZdLhmDwTF6LK6
/2uy+c01tEwmraEvnkfepAo4EVngYz1XfFivJ6JFArV3ROvlLD49TEL28nFn4o2Q1F28jobviea2
2QgYMRnxawPDjDMPcReS7Jxkwj7sd/CMNsOD1I0hqISj3R/fhHaVNaxSamCYXF3OMvQA+8AOXjgG
ekzuikVpSgqXEvakRLYXog4hRcKAJ64iroir+lCFMTyzPerU76yx8pPTbKBabpDcCG2+c3Py3olJ
73rMWX7RdNKyYHSU7666S8+ewqyC4GxgcI1Gml3JGNlO5SGKYiNwcTr8tqnLQ4GA0EEV0UDn8xC8
gVcr/xg0jTJV4TaBFjWkHaGVwOurH8krpJJ+7TIXqdAQPt+b5UpfumHeU8m7EZztK5gGbqq1jAHh
mIayheZSqJE1xQf8FRnLbZWlenSH2pDvzjmrPg4Fhe5+EXl7Gi/jqET7m2Vh09OVMwCuBR6Jvft9
rOaBW+RJAXo9+xO6JsaB+G93QpphYUaG4D2ZUEkrTuzCtIUEy5iwCYfu6MEqVCNzdlazxDUkkA7R
N80WgXTNoqegV84gT9JPA1815fKZm6O5MCg2vPxEMv6POS7CZ3zTIqRB4/iqte/J3uJ3TxT4rGmR
kgcgCCAYj/TMSaqMzN4O4H95sZjtJMO1oX6GBHjCK6ik8JDCA2b+1xWm+9n9GJNAcxdNeTjsPnNG
oKOq13L9ahnGRBB3vUksq2XOKccPb6Rlvx3OPFizdl/arx2Yc0e4enxWvlt9OozCAY7zcRZPvR9n
gPNAGRmeugslppNX8ss6bDMoen35OOyuUH44aQ2819XMWT0DwtmhlypTpEbHHuwqVgk+DvACncuw
2tGeS+1K51z/Fh09hXxDpxQopiTBhjk/0yjuG9gtwWhRInb8y32tEx0rR6j1m2QQ7n63azy3/Zit
eVORc7E5pNuPsoBEYPIDyKqIKu5nmMNtGhAXNKlpaXqyKeZCIX4q4rYfpq7cOrTID7J5DdgykMB6
D3SiqYKDjrto/ZO6B//1VL/c2GPjmfVGFPd5FtETkaIyusJa01tt/4++JG5YfEDX6EF3iIhyP97h
oD5S697YmhgKOACPh5e8pHG9PswzibSeo/vwBK/xS2A6aqE3LoVpbVw4a/QIwgLxNgXa2CkAP4aZ
wv0RCAS73BLryGvs6VJ1FLODndy+YSk6rzEnKMAylPSrOU/rvYzuiPF4OmbQ+hgI1l7ajTtHAU3C
IZvdkfGjqBEs1DfWoQa54zH2rBlP36ZWG51Gti/UsPytHDwJZOjxMphbbss6gL3JhT1/4vDeLha3
4jOCbbheV6cGtwpbS1vJOLxViBDTRuRjRNlKSb0+qRaI6oIg0jG1ndNz8/zvKGTXxnFwhtwAZ0Xv
vLCg3fo97u08rKAXEvCh2TF3IVQ+zFUXf8AERyOi6ng8NDHKapDy10sT2jinUVGWVQlOSFohje3/
QdS5/knUJOEw3n6ru7xhjFNaYXh2Qq5KFdI+YVHXi5lSUdFZaXqIvmtHNDcVX7AOH0oQXN7VZNnN
4+rCNvEowIyoMa/f98ek1xxe4FN/fyQSUF+2pEns5DuO/QueJMnVlUCixuYYAH8eUUS5MFZ1XwA2
ZBXFgCl1bjx+xeBd3vT2JIqsJxQg1/Voppzhbk/rX+TWv3DidtQXlKFivY/V3ELXgbDpAcxcz7Am
CSVWEqq+PGJiLIAy1Dct89QEYnZ0hrJ3K/mA5DhxVwOPOgSQ4W4rNCrgga7jZMzCil7cuFqLax3e
VHLkEgyZkKaY/+88izOfiK0SPcU4DC2R4QXO2JwWESSJ7EO1MjxfoNYU7LOf0SCgEKcHXoHZb+EL
n74vKT5r60fPj4rM39TcKjlFfdUWpZ7R/bkJf4i6754uL00Y3sh9UkpXohxtObtle8Geo/qyNtTl
/DBNPj04SMkq0bc40XpJn9r+gKn83P4zG8twRzRcu2sW+Mc20lL7lfcNtIaSbv1ECeaIm+Rk5K7U
DCuGzfFGn2s0wG/2elBQ5mLXipDugIAWrIJBVFTw3oJ83HogszCiQ4jEyyVNg/4RTEEPaf/86dNG
dSh78xzNHYrkIh82vtIvOF7rNGqYcm+WbRtwhUrYIxU7R8+ZFqotNX2pZWZnLWwjvvdGd6KJNVHl
/og1bEjuTIN15AUX3dvRk/9YI0UaiFPCLOkRqE7e+3L/EQ3/G2kpnT/moIk/JNK9uKfCe/LID/ul
nUTyvU2a1Wvp/Zaly1+BxVlWA+MJuz4+wP63hsQ8MYbSbln8w12bVGo6CTZRcwKD4QV9LjEDSe+N
7uMmzWqiXMl9djUWFRkVgNN7Ns2JP/Q9v6tSO3apJysSfiJrlYEr8uFPTd2cTRHhUR7lpYsCRAM8
u3QTeg9dGo3BIwICOpnyku+qEj3BEQ2AEt4QfO5kDfhALxO2RXYS8SK//GyJZUIkF/s19yFIyiZj
+h6qvFeCY7ajX/kIZjGL4PBulCSaYuDIzinHgvlJ5fhMZwDCCnb2PWjhdS9NMu/F5A7bV6gZDKOT
dma3haCabiQekE4Zf7G0lqrOm5VdNxh6tHKm23+k72QCm+Ek+c4mk2JTPZhWF/cEE7hYcmvdw8nB
EixNIICIbC6Xs7NbUEZ6ojmkOjBE8rd4NqRu3gvZWu8D4wiOFilln7qOr0fcpH/tbUGFJLegW2zY
ywlCth2J+tevPTGBcRbhHDeSOwO3vcbQYzkPSabZLGZ2Gdqi+zPN2s8g7iamQ5xho5dKkUG/xxNs
0UcbtGcLVXcF//LCI/1SnDMwgRMrOOpCAEF8jH2k6rxa0uId7Tn+TJooH75vTY44EtoFGQ2rPXZX
Ln7b9JNZuhJrafTxwodvBqfKrMmvelY6ypPjoKSw3QR6E5rB6Yzgi+P7AUG57w8Da8VRtdlGLPS9
XyiTxH2ocsQNy8pg+vUyilGUt30iSgdtjTsTzGDpgNxFuLcF1W35JkgLTGV4qf6sgigsA44i2rM7
O565UEcyNHTIl3ltrdS7gDjQEhJG5MBnaDPNkh2pZIOUi8aR8I9+qKkYW1GoVJvnNY89+HEB/YyD
lCZW4wW1PqdKRKW8g90WV5u4ukE/sm++J0CTqKaQE3kMwWZFJOeBRD8Ms5iEUIFDgti4JgL1vsk/
QdyqOw2GOi+F0qKDYWqGQzALuDUiXeexsNZ/6YyPXmg2iRpjImT0WQyQOAC5VbtMMWTXYGs7cwxM
q4WqmJx787naCwr2kPDQQEkq685zspfY3EEae3oapdTYRvGGqPlIi8p+e25TRpRpYJZDrYQS/ATM
m5u/UmS4qgYfAYtqo4sXItRacNV2PiiaG4JG/Sx9kkX6tbxLLRbBZxCS6Fv94CPvz6fa61G0QuB6
OlhLDYlSSD4kOfePWVFaEQHUpEOMrhXx1iHtgS9qRc/1WhQLPdKb7DjvHJQhLlrmnP8r0LqKNTMp
3xptygITbvIRAkPo3GODwd2HYrwGS6s8Mzh9tpedcHpKIgea8vtpfXFrEtBDs24IYMyYw/XkPdi1
DvuKAcoXutQMTkFe/aS90j2xGuvPTpWmHeSp7vBAQ2jPGSI7nUjA9RKIZcOStSCt7TWPdSfNf3oh
TMo8hiTvU27zS0nCw3WBMEiZt3st5/jGfaFQ3FYxplPPVN2t2mG+NeNUSOMLkdBKocBUiaadn22I
TcWyjhSyn5BjAAkKKPNCQ3mU337E+SKFlXG3wyR9Dm3EltJACW6LSIRoomEN/p1XXFChKSol9Urb
STtnN3f+OHjJ9UQNF7OhWi0xBlscyQCz99dTyYAvSN2hZzI0jFcVv9xy0Z4bVAU6Y6+neBqstMAp
/hAsBREDRrlOTZhQ2m+nuCp7Z8IkatQRGeGiyI8AuxgPe+FzZUsR+gQJOFKMqFdn3r+RQ65KtRXn
ZfjLbIUtWZJmDt8WUoxY6gl1ic7aGcCnCJDtrS+fU6iPmIoJbA4tBYLVL6feJmxfsFIIXU0kAsti
CJcK3Wtq9K6bduBcN9Gq1xCjcWK9qoOX4IQ1sdnmwsfJBiPxeRSzKEJbVixdiaJvL/UkG/RYWqmI
qhH68+eLeYrtrZLpxzwBysOZJNIkDmEs0vMVpgPcmCKtNgg6npu73egtC+GBy0WZvg5Cn4Pt0BI0
HPd7tS003FAuecl9t6s4k2T+ZQODv2z36LthgvX4zQDXXtsQWHfXdfCIgYpaiSmxESi0+7Z2LdaM
bMHbVuNG06+hz+VnsbHWCKrYBdxDg5Uy0AEcLy6c1j5LBh4NrDhSHrcMJjGWWjVo+gwGktasjA+F
BYcBSPW6LFwkghB7K1M5jiVVr967qbO9VwAmSPehXkCFZEbL6abZP2kBNY2noHmHimfWsaSUtCKN
uhBVcDRQVj64miRZoMAVEjBBSS/g6a7qorm2DuSD4BoyMGwfXRllyfwkPvBiwKkH2AY4lcJfracq
1Enx2ACyyxFtuOf+YzpjEguRUgY3lVkFVpACvU4aU1JyngN1uLTJC4J8dEU51E9h5SUunjkBaTwt
Wp8ue8/i/fW0C/yKXNaRkpKaTG2jI8X9f2juO9LNoaqYq0HYkFOeEqg30v4ltPjvUhEnASreXZ3+
DphVVTHR45jCpRXqnSVH6TtbgSmSKx9xlwSsS7jpFQEG1z+wvfPeK3O6xCEVXrjFsQ1cgzB3VYxc
zsi//1cpo9cCD+UYTF/pbCzf6bOSJXFIHMji8SeDJAF+IEHa2vFE3Eh1BKXb/lLef/+pw+ysF5Bw
d/TlKM+fSJXt9ml1jFlPIocQxAfKTPzD1ZniyPNsj6j/E8gZdN3RnfEAUYKJapFN9gGIgBZfNg9X
9hjL7q0knU6xJDTxq/EveJh0liQKMsMMy4kTipgBSpC8MXVi+QD6kujoFmGzrj6+Gnczxv2vu/F7
hKN057nKQQuWbN7ZwhuXzrWubN7VUnKSm70uzNOSTdahe16Gfb6dye5uZP00Om/si9wLThJt/12D
KIkAft6rvIuUfHk0T7jQ7Oc8gOadgn7CZi+kq2JL8NCtwrb1sg1EUxbroq7x/2QARP1PWebA473R
8E77HnUv6A0S93sXEedv5CxpAtBocoY2lDIdtXXFMz0vTyO9eqhEMEabr6+BX+Jl4rjntYCdBTpk
/EfTHldoHMuDbeb8IHb99/7AcSTkdWgedt2xpJ+GUGFiUCy8KxFAF0ig+w5bTR/U6tQ9REXf6+nD
59w2ksfqt2br9+lAbqH0VJUPYQRlmRrl+MC7JeQEtLVps7e5q37myb356PW9XLCAuoDejQ7fi88h
ldtquw2XzEvZ/Q3x7Ku2HMzri3qyUR9mxwqzOf8vmDnXwr1b5VXY3yAnYrSMMLfc/4dYmZ4rqNTq
oKqovmRputR2YbnjB8Ekbvx6PtDKEtXrRVVopyMXonT2Ylv9wke0dGGN/qzVc8nJavaBskOnjkTV
bR/wHq34Wf34BFAKWajFCLroS845eMgOSDISSochJBK2X8ZIOQySHdYIdPTaVxTXuK/SiRYVyQVh
L++FYRV2mHTdNKzUfaHPH2dEeJyCbh4o47wk/Qc6XK04UjKClpepaXorYzdLVkcRQK1jgzHl9OEa
eGzadfGygubnugXkEMCAOHdtRS6SGtxNlpUj51iBx3akZfm/wsV6dUfkU91nAf0spfd1Cj+FtWDJ
LW6p8VgyPjLbCg/7HB1GlyEYMDpkNN+jpsLjNi1oLxtv9wnSLrVa7aGgUTK2Rxixn7NL3Ktq4ec8
q/rkz1LsWNitD6f3KENQsCltShVdbaOtZKo/zF3mbP24oZazDFXeLCc8y5YL0M8Qhp8gPAlCpGgT
/raoQEirPmrT4pnfX0l9bhvcm1MJGYVPc+Kb4sRhFRpog9oqa8mm5TG2rtHC9tpnOgI95X/DtB4K
/roc8vdAyj0HOvO2eS4Xz93C8dCh3dxtMOLcfFKJAD144eNYU7XKCawYhqHbC2viwUOaZS0ezOfz
RYMjfiCaOCTHaJa87G0VIwRinOIGY2IuvqFB7BiUnnp6+Lm4RzYUXAErLmE7BIkZB/PB5XPTK6OR
gn55yjAvppoCGcGwuGXpGMyagF73GxGMqNzXE/97Lextia+wFPPzdPn1jKpRRPe1XopdMfH7z9g4
N/CBLzJYN7XryQTWXMApwnEYdHJRdbUYfa5GJLlA3GePfgBnQRweagMKEJoywsl9601lLqsdir0c
19O/3vwfi3kLMDxlaLd8M6fNDZtKWjuDXKzjRn3P84cCqA87JaD8BvNSzkHjpxX/zTfgPzwKNZjA
v6+oojlAn6NCdFb5cZ9mGFExeIwHAnEI8CRM1qD28RO6k3rXnSb4kUVrnbbIXI3QgVoVsI1Fmhgt
+9Pm+ulI1wUGz5p7FrPUB/YMjuNzWE8H2SGvP2scjlG5l62hUxsbsBmnGhhU3l7cUVbsyae+RqCy
ag57MwxoK9wQLhveEPQgIWV5Kab85SjuBOccpRW+6bcbgN48hkYYKL0jvKEhdISZ/OUZWFsGZNwH
EQbsdF0S0mrTDAvm+xBDp1t+SbBKdsRPMk0qqLC37ta+yYgtjv9tt6Kvls6DYjFxzJsyT40tAYL+
GIK3AmgOxyQee+ShcQYjDXq/We/Qo7HzZxZA/1sk73UplE/RjUeRY/a7GEkX3RTf2QpUnlcfwb0U
aaXuluouKo7YHyTbCWZ4LJLsDgtfcKDGRtZPXSzxJFcVZEalNrNYEzr7dyXRekZdFJsOyGBCtfNQ
kXnB6gQOb2wxp8vUxU05xmqw8iMDgk8VtkkbZZZb/CZp+KgNgRM/T1ZbMXJ2pIikKTnBOCuheEIL
KoDwKTG1FGgZB5E7GT9NVQejAWc/hGWRR40Sk0He5VWUjGT1w6ejbS94zfriSyrCapSOoGClUKqJ
pBHrz8ciweKiwTn0xTH2zub1nqmHxPfyicYCel8c+68NpS3yFw0mz5A6FbJC/BpSewSuIrFa4Faa
wEzeSHFd4mZtyHuEYQa+l/xBpPa99GdaI8OCa54jcVm8Kv4lsqnEIB+sALOitNM7HObhKR8dMq+8
Ymscw94jKn+A/iVCanqA5l0arNRlUrTv7nUh60/rqPDAEYuf2M0VXpe9/3UbpQJDG6g2HdMxfJHU
nnR+Dn1/KRf0YyCL6Juroscsb5ruBvEs596TukgjxMxlosgFKlMOJ85vbn/Tzw98lm4V8IgyUQ+S
mDfUjilQz1MYkwNNYVSJvZdWzEr+ihlDcTLJwb/Qo1vjG4sp5zneR0XVhpJRF35HOseOFoo8Aj1X
eOw+SDhpq+8mr6GYSLA/FUXSG2iVf3xp1WAQlWLYYYD4ZbatmA3DFn9+d4xBSMuUV7Ux504kjrj9
aWp6CNssHXorTC/s5AhCccOlLUrlbzNR+f+DOWtdfiUo+oej9c86E5c3gUn4ByrWqW0LK7PaUMu6
ay6IPc6uiOGr8i/WLcBAruDRrnIG29/k2cJQvguTDgsCoF66cvk8XCblwzwqSDFuJ4HH6nsS2d+S
Ly5lZ6V0PXaQl7OjavCOsDzs0j3TMZ63XEB65iEjiw+OuRvLStz599peYNUzJ/ZhpR/jV+UiWcES
3ARO1m7IEj4XQvjqBFsGK6LpaC+g4eOG41gvE8XO1pj9TvWNJBtIHT4MWCfOJ+HyAWtyXkdXDcqJ
sODkM5jYih7zcuQznRbT4eDkqpfpId2mfgdWlepQMNgOROavMxo0s9AJKx22VJUQ/j8Y+3gTh3JA
9dGqfw5cYU0AlRhnc5YdJOnGAdzBEQvUwLrsP3ci5njAtTaPulTTtvJERjxDWu1AL4K/g4quo8Hq
7rO5Vj45ZlFGL/deKSFSFOiVkwlavag2ye+AXdXQO3okKAvEA+QRks+BLPPcE1Ktf9X/TtSHemDu
66Tk1p83mMcybx97HUrbgQQK8RrG2Tnl90Ua2Uf1OiDmAXIglOMrX1Ns9lxIgRS+VBgVYffa/5eZ
yHe91wsHrRb4Q6ZJPcXntGO5A8wkJqriKeFv44cTynFnd6muQFnLPMHuFIMRzJp0EIbSrPGMoHtd
mKYvKGpuqEGGZX0FxAw8kyaLfQKxzppZ03390mJ6/R/EdxQVOeWSZutN6P79QxifbMKXqpsQNKcv
UegEvEOM3R/dwGZFRtBVvXR3mVnpBsoqodSDDx7d3D50acbZwuB8JzQjJewY2ofRYyx01RHwM8PB
AYj1yfEZknhaITEt6UDXm+buzcM/l9o/SgfBLGRrw2QfaDGTd7sP4GnjiJ0H+35a2akCh8Hegbnr
lhqX7YudAg5/O15gP8j1vF6913nn8tvhUCf3p0jzTeAWZpsJ4V5MkHt+Y/3lMjyC87WeDSE/YbOP
j+r+fzEBaCkpKMrX9QwcBD+kNFc++AJZI4T8cuSz7MjrcJ1O8dnlDZ8LOj9Gf4l4q+a/VQDlKaG3
OUBDt0hvu8ml7QRyzsT1JnMCZwLd+fxsDffjkSN/SGPLjW8JAj4Sn7KzTloTl3T9QwutqkpFh4mq
4995+0zdbX8z6XCTnpuuzCayMufYW5U1AO/tbyU5T1WdM0mo23yUahAQza+xfGMfEUdvzE/BJNYA
WZiEaYh+arVuWNp2YsDfiEpShi0BAdazUtgQG8hNQMSgNIwRiMN91ZBvFjbjd8yIF/z+dSpJaP+v
WQtD1Uv35/JW3YmfDypiOjANROf4+fY9bQ2litpEqczCj2JuB1b310vlLW2f9QgR9Rq4Q7q2I0Tg
+NkEVOpccxUx/JLq2qp27Adzst6sIiCseWfSCS8njp53FHC2ChwYixiiQb21TyBvUkRE1e4PCYLq
fNIUwNCsY2Q0b1F0eGy1Rv6Lf0c6EKVvfhqaWD0fMcyuJJCxoyPUmhsNYe15ZjJV4KZsb6mhOxex
9ZlWBr+vtraPAgHob1ldygRE/TEh5axnLrhKw1d8VzBtT4o+k/50Bg2p0zTALCd5GrM1hl4tTTKq
WjLzOHe7C93czmPb3IRHrbFxcXzfTbjrNM3UWulS/s25/aWZauibJWVTVp0CIM2iQp6IP4Cv2mBV
/kafuAGDYARuGBefAFxiQBB6CY2X3EMO6+s+RlRp2f8wEpoAufnRCluTQ5toURaROX/H+MapGxEt
flT4f56LLI12IHqRxgQ8RxaZnX+vQMkKUtgILYjO9LtDD6CjgoI/qT/FoTaTLExTEUDUhXuClcpd
ooV8v3j2xNNvsnNfaS9NHHq+DhI/wPoHUHecltrZzrTCfPiZCGVbWLpggQduFGAFGHrGEflxe0mE
mVApd9hHO8iCOGCrKFMzWdJwPUnwy/d4Qj+aKCe4IiLwPe1K2waOEegu+7E+xFUSOP/pNovy5iGf
wG0nyc0/asrj70I4Ze/QQm7assf1BrknAWBNfipFtfqZoDGt4qsSzkBzwwImd+WIMRTjeZw8YFWf
CmjaImfAJFAtO1/7Sg20sOo9WFbQZQnbTt5gToemiVIsLDAYZJpNaSAdOtPgrViip24MAOOcaSzU
VccMMSQDYeVxYOKyAuJ2GCrcMnkbKz33lHkBGqx5trPkfQ474pkj3nUqrI78JuQkHcCLIlaDlx4A
zHwNWNPyAYDFcxg8YzNgyhNS2HZOPVg1qrQDLSP0Fbp+UVP9PO3Te+8vAhPGqTKSeJMfAnzo4Av+
fS9eFi6wSqBNsVHVW3tGX5wApoWubKAXDRmbK+EIytS5IcTvYpb504Ni5Rm5goUDQgSCbHdugwtu
2GYpmrf64jCb6RFK4mlcp2PCw/Sp9ZmvF3cAMhT1jpRQGVkm/KzYQrya5OipQLRHtZRtoEpNt80W
gEkFZbkMlld9Peoy1N3HUu7A9fJMn5zboO26NteoqdIeuZljgYytAE6XqsMJP/oiGhsi9DS6gFWS
ikIcYOIzHMLcG3JE5D6tZIoVymtWM+i/VuG/UisPnM+H/xdStlP/mMWetbCC9hALnmMIVC4XO6Vn
zH2j7HlAAPFumKcr9dznthBcXxAm45EfnTQS+NVJV3vJTm58EMW8Zr/6gMU0RJonJ33fUqzczRFw
47N5jHj7O/BhJs2T7JLGaOQOFZ8wlbbGRR+I21AuBd73qGnzlrj+OnWOtSUGdCJ+aOj6syJUXCSH
IJg81z7DJ+fW0KgfcYJhJtYsoOO9bwboQdLIc4Tc2Jgnnrr20l1nuGGyRai6R/+gCOn8sMQiEpsE
qMx56fstCyl507YcOaRF7yi0vwIMkQLcqS6peIJLExZQaJmUxIpeSyLY+IeF8A3wci4cUiCkqu4l
uue+KcjCxTKdz78nRW4xjC1xZtgU43qQR+QURFZROZfk5bN1P4vxQmBDC3Lhpooe6I4HsZyLtMxa
o9olhdmbY2GmgVALCxoEDfN2mWpcgjAYqnRDDR4kdjd4e2eB3LvUqaCfWKcHq/o/hoGtib0r3dgg
SVdQBdmCvDFHo1zvmGBFp96ySMsS/FtBxawLLYDgTKu31EjqSyhUXPazR1iNPVLlEDLLo4+7U+hO
S44ftVHrqcGrQbYnzAJuddwbBAXNoTsIe54BaoN8UjjBTf00DUu9Cp0mMMn07PSvxE/v6OkvMyhK
Rmr5YRpgZgOzWOnZBCDzo/fdZeaRolGNjTue7M10e9vk31EofYRDHBj6JNeIKXbGxoU6nK4LEv8h
CuCX4/pRNyZtBOsd310/yRcB6hDMVstBf1pj6TzeOQda9ivl9luOVPXQrc75VOO/uQTsVe8FNE7+
acTj9whZaONihbW6ilrXnMsWa6ezWF+NsItM50SwBDMN0eWGqEgLCkj1kOn8ILyT0cyI8RhDgpgb
ng43jbHD0LOAeF16iWLHCM+UnMc85QUPbA/nz1UI8eSvqF8GaKQKIs4Hi2SIBnWKm0TPSGLFmsmA
cjwtKmMU3mto4i5czqyCLDLWEyO7+XdQuoxszzT0o2lx0fk8GoQ5yV5s7fuISBPyCrv6MI6QGWbg
R7hJe3KF2hz1aV4aIOxMpY6OF5FXGD+oiZhaMdJZ3FHQTfvSSeO8wtOwSIMZrBFvQfHr3C9UaGwV
slm3lpxsuVfXP5wnfjmMSbpSdHT3DDlbqiSLEa0fNJmQSXXSN+Nu2knrWcTF1Lm9Ot9dkzpJHsHN
EpKMB4HSXvUddDME/36IdavJbrl7x0CUU55mkZww2UzUEcM3YtmcMjq5E7zzZ8ujn29l2BEdlKu7
QBo7gj1qzdJ9O71gsKK7YCaaVUdGZu5H8AnYVLEbK2fV8lhvy7zQdRqV1d+4Q7HdGO44siWPJ/ra
/xoQT03AIj+yVEqwBwmyQeBoZKS3DB5VmSWUwMWSoN9262/sRMejhP+v5XpZ/ZrlBP5BJ50AZ5vR
S/p7nqM2gxavAXjEbqe/68MQjNYhMV4nr9oPWt/Xy0peabRhKwua/g2z2Gz2tQKYXh7lIZjONie7
ldGda0hnQ5Ip0tP8jCTphe/qLCCxu/0Akt6cEUoQEbkK2RVn9yXDr/qWw8l+CFeMEz+o4B6PPcJn
ELfGM/+wK5W4AgaOu0WnMq0keLLE1to2ylzMKIHTp9AgCLhFceJp2fzvn+RQYN21tNB3eWZvpIsP
EZNj7am5Gjxs0qWNZScM/OfGp/zx8Opy9jdE7U+nC+L1KJ3Is3wwlc67cK380JVIQShUi6C4KmWX
KEf2wbxaRE+cNGqpREWwte5ozoyC/RDY2FbuvrCYhPaUGrPN5SOXa4g3mp+MjfNheSfQxlI2MQYH
tSXbSOurP+7n++k4XZpzkwAIYhufM05MY0nNDV9lKvQFGHgKhmCd5FFtELDLzZkVO4cQb4r5huG4
aJP15N/nnfYyC2iXCoh70Z/SJf9ltIc2WjxaL19ELQwtcqUN5L3praR/vDYBhqG7sGQw3URJmMSc
uGiGGlnYKI1Wd9YwOySDhAvitnFdlkRIp2t3Nv5VW4gJT/s1cWHI6i07Nt51Dtoy5Dz8P1lz9S6A
x5OmV1+yBafEZTRX5ta4IbQlDM8w17YBRdevaxLQ53sRFgX56458P5PhwFf7AKWTDy+HOeyT7WH6
KbzWi21ETZ0uLr2+6h4dUgqt7B4Go7kOndXZpkYSckZWrXRG+o4dDngU7tPNKANoF1KprbHd6WUD
mrbTpSwXK8IElRJzqEXWmZk9GZOgeTzbAWmvEKcORsczJdOLbO7LO7mlKfgOQmyz+LYiwCBrbXZL
9tr55Dlh0huHFwIaJ9lTPN6sXpG4pinl45HDK0aCwR4P8XaWy40DWWWK1sa0W17clZBkQxnIOIi1
Exitl0wt+3vXT5WPrUWgfjVLe8dWH0lhom+SzFFBqayv04z/3SVjXd226jIm1dwooY5vIpRSkKCw
wyuRV9pVw4rju97rxabYw9qydvfWDk6iLM53jrlv/RPUDL19DuMdnnsYvYqDksL8tCOi3efqToHV
Db8zDpC0AjHpYjnUWdu5FndcdvPY36cNw2Om7n25F4KQCVOqEObzhOnHxbHdErd+F52F4n1CHIcd
eO+d5hgymOFX3b3vbzemPR7khmknzcxIyKgNdcP3+v/A3ADxMVFpeyBTE3FbSy8YfLdspFgAvYnX
I6rZLeAr9W9KljCtTP0Xl1XOncXOOXudcjPy1wlPBbBJeVgZ9gHXV89b6RhwOgC744+MIgsb3X9f
F8CjmnCseIomcauHpDjPRB07QFYI/oEnvmFIpGSRvsxwwzIucgGk7YWoH/bjQ6itcUHgpMO9Kutg
1Jg7eOyyRta1gzsSuWTsWVgpP02GhgrPP5U7uWmAE5/yI4sBWyBK9MsMQCn4dHv3B6Jw0BlDdOtq
dhPMn+wZDjb+KabnaHbw75ssmj+IwsfwUQCHmKU0Uv7kTcpFfxXbHxckYNAqs560DPeDzgulZALX
UGfdLuDFGrlYa8js47MB0ebkdW7T7AGSQqyP8QisEU6CkJFINWkIhIPupr7YeLKeNX8tjTiFb+X1
PzkAaLFay3z37p0Yqz2OuQZhdrvC+sekX5mnGgqY5xdjDIg4AYEKGaVRptsAz6SLYgFATOcFKZ+y
QIAZDY1u/oW+oNzBhku4vAjAT6YKBWQ+RJiojO/qU3sc38UU/jmYSPwhR5D67kBWMSssg1s2jBz2
mTZNzMpbeLxOF7GpxtPjLFVNC9al3569X4ZtfLl5jvaIfd0Qx8r9pDN8PmSN2XUKjdhQp9xJROMn
6Q9b7bnz6YXG/8iKxxEzvatQQd/dg+WmAKAb8tJlOWDjyJcedmnZ43x0eSub+6032gE8TNhjpKSl
dxTtJDEQY8ZKkrEV5xFdeq2Mw69X7+G8I8wAybCtmratB8ENwDIXjhaS/NgTPTa2qQ3lfk7WgyHu
riZ1ICS/EqWYkErZXWcmxqMaBrIZXLDAIJKdtCDeEgiHKtzvqksE47QKhKc0R5htcMF3YFKor1oc
TYItB3xfMYU2ZtYPDLTtpjrwrPjvXAwpq18st1pMWPIn3kFg6GaP1IT4vVafeVyb8D/pny7A/SfU
lIUZ/Gu+HwQHKrYnBRU2rX3aMVBT14XoGesVSdY3lSZ3kc3oUEL8i6TqBFPIpdjp5ew+TNtde0DB
Ya5w7i5PbqU6HGmnk8+we6ttYsXGmo2j6QW6ICLXQ+lkk/pZsq+trYkyAqyaFiD1RE6ERs/wrlvP
VKjXj1R8yr68WJRVhiqfx6iP3Ih4sXp8USFTCpJRQ1wsOoVlVTMnSo6rjSNq2kDFoI46PJKsI7dI
DGasmDPD+Dj6V/Nsa0M1B1CSYLRE/4zT8KCqsO5Q69WgnBBdC6EPUHMR54p1FMCGhkA8k/n2h55y
4ws/wH2RNnwhMNfGBIq+sG1I3iOCvo7WzPLkdSrjNgyJchwAWyLyCtfXsqcsVnfdPGg3OjlRZIZQ
tce0BcJxNZ329CyTuKd9A3+NTZIrrq57R0gM3fcN2mrH87391QdRfnqwhTk+mliczJcvejLwi1KV
ZiSPC3P8imMaVqH1sXVqaUzyUdVc9my5LEq7ec57GOPrODn1+smMNeVa6tjLbHf97QFrPBaEAZ5a
yD+Cq4vsB3Nlc50drelxbm103q+KP8ny0t+Z+i7Vbeb1WhDPWEj6FiI4fE8xbQWX7aQqeGWeXkU8
ZuNke1MRpvd9z1tVRBrH12IusPSmjcgfAJsY4zmN3xW7gwqIzj+xgVc1xv9uC8+5fNGDtFLPsITU
EDhnOjGm0Vsbmn+WcnFgAzFam+kqPWFsLdHP6x++StGPPkDbIqAhWXZ+S+MLS6cwIh1NTNPVm1Fw
paXJSGlvXdSYCe+C/Ityj0YXntpkAqaa/irhcxpEyiw5dyrO+jRjvhM1+Y24FYQpGhyp2i/NerZo
oxQE+sPutn2IVWZjNXWdKYx4sinIwnrkx3J/uqOJTHYBsxq0Y46EyfoQ/TU5KY/ka2LaMtSbCi2O
dm2UCTfcqA7WLp+bGC3bR+jfkRi6oMBsjbZedLr/KV5LZuJbZiKc23jSmUJcskdVVgAASoQTUifK
WLCeFjGKmJA8pGJsN+sc/LtUsbbDoUbLz5Ax8kOzsFzQS7iVZChttUCSAu+WYCTPRqb6pRayP2l8
8+pxX4/WhQ6TgY1vgQYNq9oCEoVmJvs7CMWHfiuLwLYQT3uNDSXQW+BQWtmdxhNy1ai9DoS2naI6
lLphmki9y8N2h7syFo2rbXibTXZuizcOHC2Ac8zGnVFJAjsfKe6e7HL9rvdCXfm3YpXUMfthtDh+
7loZPJnpvgeh3Zh6fxWnlTevUL3ZEVAQ9OsxLbIQBHOOfLGSk/47rwPI295MF+QoUnAP9Ekl/VlD
yttM2om1BS6ILpV4L938gLF3YHpcGA7WHqzx6A5LHBI2c0gaNMzKJT89XtkinRFdqCvCqp8OKMlu
oBLJwXUZcCPadxtJMAG1Oo07uYKHaGOn5bviGRkZSotfW/gdOPtzgVzFvq5pB0Pc/vVsdDZr+hTb
Jn2Mlvr/uJOyhmStq9yUghygGhes2EesvUT0bInM4C+R2tZcGP56y5R+LCSelWtWqebA0JzF4Lbi
24T4gqAQSbyN4dNNRSGpvP5w961M55p17eT+Mwisy7sCewSiUwH3J3JfYSbvw0bmeZZIZdV6ha1b
+LVCjJR0il58+T+Fxjye84FlHGrvMtAS/6hRgXsI1tCqAFF7FFttEBtntKgSOkG4dhrMfLPY/DnY
F28Q/5eCVLQ9qbUk8PKzy1Yw8Lwm7ya+jIwE14aZVF2cd80zkZwHuKuyNJ/4Ub9DujAzVO4Qr37G
PKZD6FYOTNE6UFj/MZY0uj6Z30uCKAz3pePihTVeFuTNUvhGasqNspM9e39K8lisfQoK9OolqYCB
kEtna7aP5Nps8nW9fSmvwk9NcteMdTVc+athkIqFqCWe6ikKuQrpriayA4LGvP7f0p5Ea3LYTtfy
+If3ai6vFqXrzbauGLCuGlTbzcJ49iqF7eVVFUWjnqEkos9W5gHkgJeyxnJg1FQXN58w/cp635hf
ZegSzhVQOKVB7rf088anwti2PTQKSDBHwtVFN/6Zj0U5TtcR0rSxzjTUWH/0AklcH1FmX0feN7mQ
dmf94vs4wvGyoztK4dNAEf70Koe398BgcuX+XlkGySivrc2GjGowgVsL4siKypamb9WZ9QrvPkNE
HVF2GsnAbbQIAkVtmrvlq86MeaMGwzS9czxpt3inO8ulSoWrNX2JK0IyXuE5QP0cYiFwhqyt1ML/
gXkV93Qx4SeqV9Ft76IINaePUIUXl9sB0t9kyfbfg7jl4C/l0tXD3Nai51XEHHhPvM0xmhFc0YFf
xghwN8XQVGs8qypYyoMiMsA/vV3QCHURHqvhn3iPVU80Z8OT/qMk3zrAqirwPct0JT4jd64nBiPv
+8VqPY+1Pwox0aIQSorgH1Wsak2yo06CdGk34m2LJZfpvT17b6ixvGVCszMIyC4n3OMlmIxCg+dP
ClNUShxSCKpuwj1Lcaq0Np1TvyVD266H8K/KRixITj2Kr1K0AQeYIKFGWWUh60HbHzuFL0JWsgxh
WVmZ6L3aUkf4gqHg0BACZ/AcXiH2f+yhC3zqlLpezVRwIZjo42Kf5FSj6GDulWNdhBLevvXYW3vJ
4+7Xi8lfDTVcBbPcq0gu1iGMmkpdfR2imvLo5n5GKHfc4KC3qMabivjhuoXJjkfRH9CLKOhC9Acz
mjN6RjmZiicfx8MjRgl6/K5QICMKcesiDOy0aaROa5pL+KVn0/c67hHS2rgEVuEUWk+STPD6Cr0n
4zANONJUU0ATnWTd2dTCvFGxeluDRkD+wk7fajEIPW5Akk405E6KjxkqOzRQm+5PHlG36I/Ev6LE
BRPWEBRWB5A6PmmnUg7eNHRpa7GIWv3ZMIZsxefZI/vG7M1BJiE1KjVOB4fRYUvfEQVmdUASbSGq
ohkLpWKCSCN0b+OwUC1z/88+i4mQysWdCUqfLNMkCyp3FH7dTm8ly5VOq8+LxaUqIKlkvVrUvaiO
6jG31bUSQAw+6iSdmFVbyKEcFhxNp5QakBlkB7Xx0kBqJiIPRVQyNiaAnV3P6Lf/PTlTS5GVazdJ
2AjeglZ+uzEASkZ2LO/7PFgq7fighm/vv04fMz6SWb7fx7mnsbxCdrqe0UmHP+B+5r5Aqq5jfMDJ
asSiPW9D4L/KxmW7ZqUuUyKAm8oNuLW8G+w/Lbi5+scmNkmbqnoNbjJg4gEQuu/ibUCFYy3Fqged
O5f1a02Mb21vUK/oo9njMc+pnuMysvZYB/fUYIGzp2h/LgGqMkNdmv0R7PObl7dx+pNWPGjrdF4P
jBVncQ0+5AbEM5W34EkBPbL0bhRyEbN8NhlNlf5l/c2psHTror2bNsyNW93oyv+iQGBNmqgpPEBC
kMHxsF4jISp9XhyHipRHLUm96SGJnrCauL8ittBIyjvEQdPvCkWYIuCWZp+jURdMsjCViMyC3uXr
58xrli9u+oysae+9N1K5/EwfJpcM0BjyaZRN8sdVtZlXhxIXFLM3nDtg816m/wjAVNfr+/VxYt/U
YeQf4tax1z0gh5oJYhU7X6nC4OLx7lBZiv3fV+VdMOIxrKPU9uPSot/TNRB9C8TMXkU6V0M2P/A7
HxmAi4hR1vhIplxGqp69SPdUd5VVJp/c4nsm4mgqeZyQ32iiSS/Vm0KkaKpYbQvaBLV8l6yZzYyX
B2iJiHu5P86UgLRBL+flUUZs72Z4vyW0bLrea5vUoCY0pUylZgS7vRq3U4kKt3NQ0ia7KOfbx49i
wtz3y51Od90VVZ84OQBQoS2c51DpDNnJi30rBGjq3yxjV58q7xoKjVkcIaXngk0z95Ay0ePQtiv0
NlDZQZNxIlzkXA/hYRtlAtVXejVBjo9KKoEfUurun7Fdu7yhL6nZsnGjzLNRj9kxjbtANmfNBaFl
Vx9fqhCIueTMwvFQE44bgu5PX2xpNRyytmIWn8hiBqRzWslEDLkufFFAJn+6qJ4ZaWJEMjzywNM9
k6pztEgqH32H1lJuhU/4gKqTmxrQ7QczbVwZVyNaq5OIBtI+mv5GpZXiwfoMNxmowKx/5HrS4zUb
0Ny0Yw0dqDYvLP3rmBVfeNozkFaTyZM+pxHccjHkjp9dGB8buiWi1TOhkN3T88zXxrFzMn28DP0E
3SUEeb4g5RTp7WMAGpUvLo13gm0AAitQn7hKRgBac42nuKeJIrH04KPW37puj7yZCVwUihYQLJCe
PF+Oy28QBBLXSqHUvu9I7NxcBArzx4LD4Nr1ZioCSfOHUyIbVWPxICwuXH7gRcDxS0rqBOyjpgff
zkrb4doFTwUGwjm3OfMEdVRgNEyyHahbRWiWyZDg0YjP1+pevjgV50Yz6OQk4/A37amS9Go9auVZ
QM2KAqlApryIwtlwuOEnACfq+WzHuh72zfRAInWtT679E47rG8JOO0rl6tzXe4dIxvTrsXJrK+SK
l3C9TKAgLj13LfvaSCLjhLZO31CCcxPEcc9nZL0nfMpdsKIatDBOVshC/TydQnJRxn2jG5y3ZEtQ
FBumjMdaqJjCNkZgvN5vjhvvxytot7FCs7XTvs+nyMBjQCPiP9kfOL4P1U2dhCgJPx5M4ouP3T/o
uHoVpB0vZcwmJGkxNeWnETg3/mKD78uyq81pFLYuSZ35j30pJWYnXetOB3RcXp0qc8fNSB3YmABj
vEYFFh77fYRMPKkoiReStMJnI1y1ws7To9+m017pQrN6XbOeIUedn8d0ZZnQ5lxWlgF1yu+BqGbR
l/fWn+K9cMytnDsnZ1vPY7XGvNpl/8D4PO99MK5BAd9yVx+2Zjx2mynlyFwurpIvulU07W4yqMwX
ianJzQSP0RL1UVXPd8un3vewVFrb6M76TmHRl+bIvsG1eQC8x8TgR04VYsiq+GWsuwPB3+m8HOcH
Z8pQeOUQKFFaHqKZdBEjtkTlVcscKOJVJ8ISWWA3gWocXO2XREGxx/Cp1EF8/oRj18pZpW+OFSIK
L48sJhA1hkiYe5GN0GXMXEjHE/fk+PgAcxh2bvc9l36v2C7Ra2Taqb2kv3Ox/JFqMm/HxBJExhQf
2+tN3fGNkVHYFGcHBTrVANP3yvRBMHZJcEUD2Z7yG9tdNiM7uaXnWljQoIW+0z8ev47VQTZDptyd
e/JkxWcGA+OyI9D+EHs3dHJDn2Dt4/VrZp4J0p1vokvY5LXP58II0d4VFx1yRB52UWvgYfrSiMxo
eQYySN3yOeKSrUhhp+UEpB/AuoAcjc0IGeMbQjaWhxnjKhDXX585xIjTadiCNlqfXkI9RgHpOC3P
HD7zMVsP/R3IsHV0g5j3X7K2CjE1rAaxR041u5rzXaDNGJOHPTdQxeGs/1dhqjV7vpH7Md+dr3y7
Q3ER8Yn3XeqrMsuXBvdDC1NqkmOZ1gfnYoxthgW2idDO/YBNZM8zEbVNo0yrqkvFLNLIFKrXpmeB
EyXs2lZ1gxmK57NAPKV7pb1pJ4eeb5ySKJ5N7iyY+fiscHcGyQ5NS/MtGjPwPq88oTMp6DFPDp31
qWM5/iep3GRAosQ7NS3pp7R7rx4cDcDrn4q+HFQQGhKdBUIfptUosqIjghGUZ+CmrDfQvRbf7R7B
2r14AByf23w1xad7BdS8igXWkhXKB1O3fyIL0iJ8hrngm71PRif4C20asYwaR051okGuqeF4PnyO
jtkNmfy3+uSiPEtz6+gSah6WQZ+BJXaHVAcd43qWMC+e3yQgTdRr1aiw0u9nuZl9nWjls+e4qhaz
skieDVGUPNPLSLCJFpuPhSL9UjXtIs+0tkfDbW2UrTyREKTIcR6VqSAJwO5xOGRWMsC4zXwX7d4b
oozK2W/0Zk0ePwW+obmZdHcEc9emEyOZ7MIKgWmqD8I+YsNLskoFDjVCuDppQ60q62sjLYmbCEKT
/Cs1qWTqOCISN2ceQ1TKmp/CxqDoOxGbNRZL32AMxsPV8LC2cUahq9uY07a2Tq5Q4iJJTHQu2RzG
v6eWttCMmhNKPpac1bzGpImgwNXw3DQRT8vWP3iqpFs5UEGORD5r95UGeTSulT4+pENrj0wmJKqn
3la4R5qVDH6U24jVfB36zE/1zp6W7jtvGtOH3S3KlY4hrpouNUdLhbz3HO3pI2ruK4kxwHgb9urz
lWmPiue9ozN0T2GFD35nbLefaK0HhKnSps/sJe+omFUggi+I0MsWy46M1BTE5PZpBstvyX3DgHl4
uivm2Ny/WGSw+qDxMb8SjHiWkv4nXBONm64ErWlvr+zOr98CYQvGHUJgFD40nWLWsPEvcSe8H358
S1yxjzEcuoqE2nrLkUhI3ZStdJvMnqp3SxUlYVW//5t0Uvh/1jo6z6yD4Ex82lNlK6djnycUXbYI
5xFNjnb8QGxShJUC6gE5lDOQ9v0rtFn/YHtP1fCI1DOjVSG4CxW3opeJKolZMdXadG9gV6i/AYqL
3cBfuT7ej94UJ3qVwQ9s0GPas371AD266HgxGy6XDRTjFwl0BVrGnqr3c0HxJYopVxK2tvZNm/Aj
C1iGy/Qfz1OnbVMuz41QtO6PdVAJuDX2eOu2rCxO3UO4fjvtAuQn1E7nEANslhM82a5wptZvABbN
uG4rjEJEketu3X8Te1kiShQ1ITf0yTafN+YjFjuqmuOOssSrwHOSRc5GOk14OFqFiEOt0NdHAJhJ
VFi466nrNB+pKrWVBJKm6c7/y1X18HKge9bWh5+ljh+8jPUMaIdE3RdtR83jfdr5yjXl+UDNt6T4
wJrkXgiKjnPVuGZ7CxuKiUAGjVKBxYYbAAAASCU+SdyoKEu4TZmgWHz5inMM4clBQwgLddOzXRWh
GLmkTFdzgBSmr1fR1tMNc008u0MZHil3kGAehSqbAcYZM/H/z3JxBvMh7PEEmsawt6ODc4OnmHzx
E0Z2Beeo4fqopL/chUA52HxevWkVxwxq7+J5LWBlaBd0WSFN/GVlK/LEFJtaI3d0gg9F13WZm2u6
TNHiwm5KqV1rg9ESMiZmcZVeRSDMIFY6ZmKXDiMwVZwz82rflQanVWQgpu+DZWdSlFRcxhYiA/nk
xwZ14FzfSB99ntYYkKSViVKEwG8KKS7negBPXGlz4rcILV68KnTwS4YUjcX7hrab3fgoBdPKz3mA
rGb+jlCjy6RGgvmbfAuLXSmjzJdFQ5GklY0W7n1JGWZGG/XUk/tBannsNpVDKqxX+OJTvQ1z4q0q
c5hHBl9Qqfem7/SVLr0CLr1QB8YCZ4CtxNY2oi64UaQBjnZsuFtTiAwL8/eC9Yned0/AafRZjlUx
X36cRxTVQWmEfEeAkPOimr8ATjJ4oRun9BdPyn0ZJy7wChNdEvuzZOK63AhmdxFIO5s/ijmZsooc
bLkQSdoskNuTkixisp5OP/nKeed0CDXReevyGdBOuJyxI0s5cHoHWMPeX2vzqkGbk4k0gFgf/n8d
NGw1UfDaEHrsrXXsfVTB2gTGB/yypY3Pj/jJ7CcwEfYP3nvphOCrdKcwP2+rLqUBg7iMNAUGYh65
XW5zrag8ySjWv1h21WcZJXB6dFE5AGqqDFTjL96Nd0a3Lv3yHK2xR7+6KVfmVJKOuC4BbfXhKKJw
5v3HDvTF2wknYuUfBI2iJ6g4hCKWjilVWhlkUiuAa3OV1z/xba7iR7mpVpWr8ostY5ZPB1YC0Wzf
7lOzmOins3L/RSpOp99nO+mk8+CZJ4D1xicD5Ayhjqw713Y8rABMKFtBeP71qfnop1thrkWbpD3p
cEWpIwyEwP5Xsblp3sMjQdw9NAPPRHGujrQ5rzKN9hGw94YYCV7f5JY3t2v3GggjpKV3+sxHjwvg
gE/GWuZocPlmwuIFwLAxTxiTrgAbfoC419QrhP0grxL3nrlM13ezXu9LsoGGqK0kdOq+6F2XMjS8
vPCM+6feYI2d9URwVTFRvkLRKeknlOeU7WU/aakStgZO4fsj3WNIw0Ai4FFrcLIQlagVx2EF0VN0
Ngm0OFwA2vYcuplWISe7+ctMy8M6NX+2zJoYKmKOR0ygSSD02I7a2zCg+fhy1S0N7wCUUxv0VCyf
XPIzAcYKiZyV1416osnuAoy06ncEfeYdM0xK7hPdDxEF33utNQJauNxLNuYH0Ps2rYEQZ0jXGLRd
eL+kNK7mjMiF+YtK39liqKhNQgvD2w2xlGkczBpENcw7y80m8AHDxYzajv+TnaMLxjSRqHUn7+BK
JagHeslI6nqcMrfuVdADh9PVVThPZtwfPHgrPyOlYq+QXfoTGPeq5Iz4m5Yyc2lRXeLJeB1nz61p
rNmedetEWmVOS2fxE8IHyA/TxrmD6Iwm04r6osmuKjKKQnSRYOnQLgYpeZARtasGv9RWheVZ/JSO
SF49ZZ9q8aI0+owa0/kzfkO2Gj28VvpYmVYc4EAVve751ST33Lg/2e/D/74FEhij4sp3YMEcnU6l
Q+XhxlPnXtIxzzpswR7CFaLOu9ESDXVacucqSbfSL8jddOY2INCn20s9IC2lDF4hGNllpkDWK1Lj
y9zqmyOg0qtQvRZGHtvY6Ul5ca1f7OKKo8tg2FqjBAYQojQ3a75VSK20SgyQLkE9H/BZIK5z+6tl
zdt2z3AhPQ66Gs5IbvZswZFImXvjDQJdcr1T1kn88MYWtvyrcOU/WKySxuGjTy48IFcVMvxAn13c
A8iathHcVGQ5memq99Hlq+rq7vHzLsTQ438WgECo04BSUlxUD4gCbU/tUsfSE0S8kVDRMrpuPiCw
Mw4FJgcGl7I9fwG9HF2r+wwWr8811shaiYoBVCSwQUsRsO37S1QyXr9SGUXY8VgxZqRzjnDDAVlx
lr9GkZI5QD+A+jQwu9zyxcSeWV6kFayIVgRcI78QjxQJTLLT9D0GzWS1FQ3liXGJsyWTtV7sqLjo
RKVjhjc53zVSX5E00brRO9mi9/Mg+ge6j40W9hViB+v86ghAmy19lm63R1CTWFFRwN982IBgOsfQ
DUtmhDoiKcW+qecwqlkiyrGJDbZHYOn7I622NFfvoP8MI4JtEuhfYdP45oN6pGsd8ueaQmf23Ucc
iIEZE03RoNi7syW5Sh1EGrw4zCCRROQus8gV5X+cSMAqJ+FkluWttdnrA1tkWBI6/Z8t+Vo8A/fx
s/UDLqFcLBfNR4mPz7vutQl28MNOTdu/XS+Y6hz76jCAViIWEDV1kBiPl4+ACbTxBbTMQJ8fUk8E
GDm09P4aJ102HF3QXnUCKB7QKpWtL7o/T5j2fbcBpDyBX5oU0PArMHIUYo01tKfoQ/+HJhYhiUTr
ltmAxhPckWaY4hB35Si6SDgsjh+aa2EOqZq+gD+PLq1fVE7CvRmG/84sY76u3JRPUjSIXeihLSqW
S97BS7A82E9pWrolE4WAbCg7QBRH3+GncERjw3+bSSOspDK/xykN7HCfbygMHkYv0VF/nUNEFtl2
h358UyL0MuMxm+n0OCKeP2VPIrayJcT7v2LBjioRuBU6WgIexj7dv4gLASSXszriU6lgPcGOrGBP
x5/Zs+vyxLqbxrr6hb8u3z/mk2zjtSPSsst1TB8xF21O6qa6M9MeJE5Rc50bJcfT836fmrvUf11y
HvIOPFwFbDWr8VZh/uQkBa8tiAKkB71js8F/HJ+ck/Rhp6rdACgFjmPQafagZ11BsK+t5zgC+Tgf
F4PFVV4S1UcqE3CLstp6Cbf0lKbnM+0Evb5/s5VgR3Wn2gdjR0wSHTKAwNlClRhGnoRr+1Hb25gV
FwJe+glJm8lGN9foHa5qYUxkvXu3nwWVAmysXpyBFb75pn1dibh1dGklkfPi5SesQuxD8Opqjmtr
Xkh6dS4Qy/a4GhvPzjzDFRGqFKAEX9nd4+ZflvmXvQRtRVVxp4crV2AtKH9FT60NceN031ZcLwtS
xjQ6zGdUO7UFAll7sCUuhD0eN2vbzohCQMWJQj/1n8AF3ZaUThaFAaCn4R82CfNYrMUCvjYwTUjQ
k4U7xoj+uxzhCfjmCfpXCCD1cg/F9GxEPl8LRLnt0Gx5cqt52jmVh5jrXGGJxTUb/+tgyGzceAcs
QJeKXPpYVQuGRipUrej90y+ebpgIrsIKS1U9JyzCHZccMwDSSB0Mfnonx8ZTKlOE6U/fARPc8cA7
Pdh842we6yl66fuLr/2c6wesesqC4QCguBM+AiuTBRc1eeDn4bItGGomghAWdvNEDYyGq0FuGwEO
PhlGoZzCCGvjZfKFDS6fiJcglGxcEkGKPFdiIVFaSDadzHgNVW1o9fU8oA1IFh0Caoohmtcc/o52
UVW5g+IzaFNXeY4LXUr04E/UIQ0OWiHQzyLta1E41wHmpqOfyNZKPECvlHL8Rw3RWeCYQPslyguS
qhCu0/hjh/KuD5++jG8mfd2ZZGUq4iuwjZaflJyrIJAAfQvFv5DDtKawz+P7p8num8L6Lpzq6UH6
5UKrAHrr24QhsP45GeyBC/+vmgHU/MQOJM7nExHLwXCDLcY7j/vFYqg4pEEKJn5y2bmMIdH9pu+F
kCv4lA41WunqZLEnbxYteIzVMuarVWmfUxwQBwyZlLyzcMKF0VxQ0n90VG1mJkHiNAfLAY+TU2zX
kS24pe24lvyZcD+ORjVc9EW0bvPKeqOOaO1nQqrjZ+5IGyqJjFbBpaY7ex9vht0c0haAPMG+mJKA
vYSBh1uwwMA6hqk2YdfPjCXrMW9PrxrNJgMS6mYUlp044df94XrUQukKgYL72aNiPMWA3o5YgsUL
RjBJE+OLJl3sJITXl/eEOwqVk9qvvbJcvMkQDzQuxvBUAqRK6jGVRKY+uooGh62xgP2Fgvii1Yst
yUyD1Ajo0wy/y7SgDMFBjUg3u2ZdZt8E/OhVRGDkdsNkN/qqr5Uvlz+cm2k2OQJa4J1je97g96x9
70VcFd/kT6TFe9VwQtpLctYFjaHyAXv6Coi6F53o27Lt46B3pDOCRjvpV+tmEYOK9PwJymFqrlIK
ufXDtoUlDFFZS9z/GpOR88u1UEtKuLkMZmLMVadu/p+k2ctB4H6i5tdT8f965VPBMhqDsc94pFLi
2g1uzU5WJDaiKmDuwhfOuNe8kpmf7g6JrG/v2x7Htk2tXHaNLlrV1V8R9T/IgRFGksWTeKWbp6Sr
DizNtSpxECWbkzTnk36WqorjEde85cGNTdftbXpxqYohBWY40gzy2EyMt1wxYQ8weB+nwAlbPsyZ
3tD+ZtMXD7rwL3PZQiqnsyyYOqWUiNIb/Pe/s2K8v9DQdnw9b+g+J1/zK+fAv+itbbd35yLkCJYJ
3xWgaJ7wkKt86aFeiGNoEQgeda0OVL73BTmONGWCKlnlLpYBChHWoOAMfmjNLsEpZMRwAHaoACBu
I5KJt+RM9FuvFjX+Ypf44GzaGfDRh6a0X6qgUFvCwZb+TwMFjP3ty/4cE7yxcP78CFq+hiXkkBIO
f4NCP3RPKbe6QOKUMmtA5w50wKtZ/kr0fclZABt9fjhF3ypFXlF9fK1Fur2VznTzl20vy1P/O1aV
LGzVSz9lK3VyzWECy0plfAn+9LmRY+1fhX2dvRpbtQV0bu3ZjuLRg1nowbd7i5XeVsbQlP8VkcPR
Svs+jWSw3ii2JHGTURmFmGf5dAvJ6748kJ3QCl/1HgYqUujVbVCEArN7CfIyQfaAyftkpiepOMhV
QOwyvDc9qiEUXiaxJuv8sGx0mE6wU3nN/Heqx8kF/D8eHLqdbVCaC5LZ6cCO9ovrYzs5qeLaO0pZ
181wMeUJawj0thEpoq1K+Wu/TbCIK8UPJG69AV3f/WFDdE4IlinOkPnGlMYqrN6jAvtxwykl3mgi
aCXTc5t6+GvEUE2pQGRFbra2GlM3R/FIpJRrZBCkSwwefof0l7NiJHh5BvdSjpcQjCFVnwRv93Pk
r89L1cnpl0sHIclAIEFkN4PLmh0P33AZADJMWWgfykmwscCkvNjKaRtKvY0Hm9ASARSjOaAuadKW
Te7lwBkAOlnCzvV55gjN7ChAr6dYnzSe3UZI5FKNsTgvOZSOr8jLj8tTCyBNn2a1tsIJG/sQSW+b
5ixmRH+6J/3TvFx2xF4qcwIs1X6kUBRc7x7sRl/spq5ZmQ7BsuU23gi9VeGiqoH2FFOzHq6gGrF9
ZdcPhJrvlDehUSwlscrOiFDDpgh6k4YGwN+0dzWHuZ7NOVjF4n7lfh6Tn8nzMNIZwzoKJapQa6Sn
MLYPqR8PvJn1FXrOqXqeD+3JcVjufqEgM+XPdVXzV1GWKBnYaSDKJnokYuhzsjM4KRTFP2w/ffRP
yPhPiSqgsLjJ0Elqc48KyovQbHN5VJfT8flhD9DU8ho34bC0CEEbhHl3WJGE6QwRL2yCwP6jxI5/
x08j0oBqiXqoW9ZnLEemwTWKyy516P47kvZ3X8ssluRHJ9XxHWoHtov0bss6rbfcYWHnGkqZ9/Em
LRIhj6Nzz01SFaI8YimmhzZTwH6/qv9ETGR5OnEKCTmP7bhE7wRmnb7EH+jzHfbUoCcGJXwIYQ6h
Y+AlJvXM1Lp0jsQGmeHP3HzfSPWHFAe0vGvtOWDA7RvXLlmv5sd+vMqL9zeZxdecqJ17zQw16W0H
EbFIkq6gQgpf3yt1yuC5DbNI0D3X5Sqa06G0NbMTl7wegkyG1Uk+dK0ORlzNDhS+vj2sDCk1vPQQ
uN4qg4GEiUJG39yR7RMT7W+t061P0sXnmsrYvYCdsjOfiRCjnOLB701yPk8DRxqJiTJsuRfK344V
mG0cCgDnuU4V/oilqOWhLuTslubW3t+ytapRRkZcQdaDBcl2jaF1k9n8UL7WzwDncBljSQrlvA0a
kRYxXVPxqkVJmEnepmELOrJRTYK/K/THf1GSkPG02rDsaylX2Rt81iBzip/0eLNkF/LgKSOBboWe
Dk1mGzyTVIBiEQCTPs2Kdzh/tvRxPUCU1WQt7/rdjgg7LGM2VWoCvuaUg4pLMKLSutvKwXbc8FnI
lLcSbf/f2AK9CEQOnXp+7PGwi7rGxQvvPaWovyUeiXVmBdqTgPDJEja/WWR7YennOJQukIIzNmYc
ZF+t/FZXpQXVcpj57PkPZqiutDarQ2Jb3Doaxdb9+JIwttgRbYQ3dIXokzQKAsK16RokmwqsnTKb
x3foFwe63CzpR2EFXDeCJGufcATgyfZZ7a225jo5ZbyP4o+IsaSPCxoEs5BvNp6vXFzw8Ff+xVz0
MBK5iGEAl0iTw0f8vULy3We3pak6FNfTE8sUBFmWo9n9SrFB0d4N0yYOKMFU4Oxy7Ch1Go5fnBnM
DoKKRKN0WLmvXuulCpfm8i1rfWQAmNSwKpJ+71rAXNm393Pk0B0JUG7KSbFme2x/kGlkT/K3dJ3a
b/0mUD8OudJ0xRmKsgpYpgnHY/7KwoB/XyltdNQ+nMOz7HA1jMP7xkOOehaUJV8rvIT8zKorG8La
dylOEoxTY3wrC/3uYH41BlBhQa1cH/IRntXb1Q2n2G7GcIuwAbgELxwVehcdw2NLnpcZQbRK2tLj
m1omSt+NAcYY3GAidIdnO0gWBRr6pfWRzmP/SZHqJukCT8H8ZO4z4N0szdpkPA6YK8JdfHI78lij
kmu8hULpb2dp01JwXLhUcp1q+EQIceb7A+5E4Y673lvuNFynDBXWfSmGS0LOmESmZ5RaJ/jWY8Ux
iSSjkhIy1KBOLAwb0jDOJ+4jgeFKupu3p+BiCUBzdTHh4a/6f8IdJqcOs1b9tHFsCXrMTKDjP6Lm
7usLFyRmSuKGagptR+CYS53TQn5AAg1RL5S6TmHCoL77YMk66YA3Y6f8Qd2+ueVc6cu0wAN+RgJ5
P6Jqsnl6zGKNwj7Z3RthnrmR8W3gs0k7skPzbVj3ysHu3uScLPHa+bd2RWz2d4bSiL1n1g+Y3xTf
S8Jbr/y+CJGuyf/yTttKd5Z974uMVBMJE5EY1AgiXSERl4QujFpn1wVytbQlr5NOrenRkA8PvUr2
RndlyddOYpdVb8cSzDjSRaVIUBOpQOGJvA8BZiP+oErfB2GYZEj/sAHC8JUhU/4p6Us/eD3eJlwO
LSsPS7ch6f+2c+rXM3lyHMvinHSRY47AOYfN1B3gYysp7gJ5H4Cob5cGx++2+UdXOkFK1KfuoTfX
LK1yMjpfRucUb4wItU7AUHrcZXn6eA6fxdMAhr7xJRUeKMfClIV3kRH67iXYntujboYv8c9RIaXY
dQ6RJ7MI9yRqFVhEMFkmUkFD8tt/0o5+x6H2cMHwFlvGKAHvjK2CCuQh8xqNaACAHVTt+NpXNOpu
PRuCwvwMUr1qi1bR8CfF/klZJARr1P9SAy0Wm94JN6BSR2iaZnq7l6zvz2PVW36b55JUNFOZIvja
bEuzb1BWeBg8ohjrvTr7ZjaBtIBaMJ/eUXF8zrBnISq9Y5fFFuq+FEQhQW1sCeapo4aSW8gOrUf+
DTd2KMgmOGpqXcFf7NJiGILLScWDs3Ayg25aisJgS2uhg3WKv5HuJ565ZEmEVpUUhVms2iAHw3wd
X/G7UCALW4Pjf0YVsUBZA2tGRgUNYAqLPDvpe634if6CJT9gRMUl7Dep+uHjpPtNOAKVFnKPzqIY
HqPzerUdVDjALHOl74oh+F+hmvfd3bPI37ncboWdNruTIXNuceLuo6OvuY0C22Jl8H9XJTDbsW1f
Uo+wS+VGsns4Q2qO82etJg8hE8udgHXJSa179hdKLxPErvKS16z49rvEwWvoGoFaDSJ10GdUnJ5s
yyDhULEqYa5q/Jlzz/TAYuskDCZqyIVpT4y4Cul2xMpNJY3GFHT+nA22mVFWoF/S6Hai7UQx/X1f
WbCIfEwwbwrSPIEGGZ8jvJgxGDsXZpoTCnTz5m5qpsoRUv9/euGP5UXKPOYpecLm2/guI65hH3Jg
K4exRNgWvQmuygzLdvUcSyExnKnpCEWz8nXabyxFxNMvBJTV47aOvbk8BTql5klGaNlHEjmdKddZ
edicH9IZFxTgZJyBw81p/H4aaf2sRCWdwMbB/E0huHmllhRlAf9jhDPGd21ZtJgluFsz0h8qZwyO
Cq7DL/8tZ8767MOWqBq0UNd/uLThL0aV0EVLzmZFjyB6oGUuUaXu25F4kpLlHW9qNd1jvWJojBRo
hq10BBvyWJ86ezh2oqN3jTaNypHEJfK6OZMkR8wCu2o6KOu8cgY4OdAf9u131lYdeND0tm2ZWVaO
kJE0AWqda1ZnQ9FsCRF58VumUcJxuz5vKPyVT/LUb4O/+dVMEaHrHR/tsDiaSGUcvW7CXSSn7NV5
xOjqzPl8urZSSPG1nslVsc5xjBbVBkT1BjetLzpR0Khd+u1TzC0ar2D210lmU3IjbwONr7G4cvHQ
8l4fraNuF3BGTsv9AFUQc8phG7q1sQXS0N1nDfMHkeJms0zIqOz0+CImh4nhakEKvZG4/PEWEhhT
ZSadiL6+OZQySXW8SdE7heLmcGTIUedOZ2PDz8Q5kxOXK2Lv2CEQ8dhG/U8AhasJpDAfOG0+xc6t
AkV4lf38xL1y10Bbgk77Ew+xTOmOUqHAM86+LrMTicOQIYxdlIBa1WedzGsKKGocTg0O3iVlxxzv
Pg1IaxEzPWNxG8vvXJTn4EksH2VyZajPVGNQ1Da8vxBl7d5TENguxyO78sicegLnlxsLq3+6uQ9X
TrDOguoqStjQz24w+5wOoagskOVPkBJP03gayCMUFzU/R7Zo9u0JahOWFycBMRHKjrynT2CtIxpc
96kFIVHF66X2vC4iFEpy1b1wlxgCq2lsvpWxZ+hC/pWZgJ3VuWvvsZa0dIBlSkUHe7i5xUzA0oQT
KpKpUdjlgkDk5nZe7UHUg66dHmP5Iv2l5JIlrwqTSL9zE1EyGEqeIupEwHwIu69SW6yvxQXrdx2n
BvNnIN8x9DoMgf+HG6tYOBSq9zV4D5w0xCoqQFyP/p/08MmNcCi4P4pp1iWsyIrkGvsw8lMbKknP
lCkjjmW0MxbNmFJ/PU7F+4TU7vMyJzvtRNdl/QeFvV4xJSsgRCchjG3b5oJQJmOODwTjmbn8lrZW
fYZhxT2ICYUC2qNj1LOZcSFt8yKTNPoHZXN0Rc6P/5PNU/XSZCou7EMwzsaYLLHBLZ5Wiv52xPWV
5ZlnxBOEyDMtlBpPdJj9oc6pW/kuJxCjH9Tc1HUv7fNgFjQrcWZ/nqdK1ZVmDaw6L865k4l1VeQC
KiXBjdIxr5LHa2gZnU67Za1OFMp9Tg6Lsgc1tjaQtPlrvaUmcT27A97ItSxPU9x0h3xpz5DmHT4u
mZa7/B8QNPuDBdAlI9hFBQJzscJ98pL6e5DCRNWavRjrNpoPw3anWz5wqn7ydwpW7M/uM9CaE0vx
c2a1NIALa3FcO0oA4jfH5S53CVhGerGMKhn+mXHfmTSIJYdGbNus8rBmxhDc5x/VbBpTolcAnb7M
4ZrpKJjqIODK521X3MOBcXpdMBqItiH6wJkuDqqsi55b4GxZvHfU1DSXIKKrdSxgGmge20bIvRjk
UcvblivnP1rNrzzL0Cs6sVn8YD1zGAq9VO6LJTD4lZFFUq5pk1EQgpIpSHsANMzKB3SLy0pDzQ44
m3uXR8VzU4LcTpvfLYKz8jzHofiZJq+U3iD+vrR3CZVvfVg8t8luZtWRGjIKzqXl4Mp63y5fty0V
WJCWssEUtrm0FD4alxd0YP2AgmAApRm5Jr6PhIbRF1xei4UOEkMblFBeSTPOPJ8T4YRrxIa13ZKT
JN6/bawFsgwD0rhIsy6ZRo8UkI1FW3s108zDwjr3zE7rZfOnyM3xgBi2o+oFPdpgS8IuK7nGnccK
HROCSPyDLHOB3QciXuDWXTSTEeyeUsTWQgog9MckYt9R1TuW+VI4DskL2UkIIaD5WXfS0zRyuLSq
yZO1qPh3D+zsLKz5hwWTBtzdSSA4FG80LlKnKn+EA1r4/UyiMEf1abvWotyrPhpuf0lCz4cdDLaJ
/UV+DqaaF/hyZkGqAPvSeAjoGwH/qvpV6qGxxa2iAn3cI7fOb4vVbZQEBpnOxAU3p2brs3IDb7z3
pGtXeISTMS84WhEiNb1a3EAa++rDNoI3bnlSr1o/of4dKMB5KXOF+0XsjJVgEONDGAZUpumFkbie
knPrwyqSQsPec+Lo0NfutsyRNNJJwA00Hp+XYhqNNDeFKnKoL+J8BYrO4qcccyyQQZU3GGzdiL/p
F9D64kqtwyhmCm4XHQBcOIwyxl6qpfr3ONpphsKVcrknzeBM6F9uPomQC1birv4ih2g9UyHhc/TD
MYaKOyHsSssccil0FumLPB3Sto1y2h1a95auW++U+wJcPGFUmNxcHLE4F4iYJiZVdLNwTwt3Nw4B
5DWAHpm15/bBR6HWaC/agwUQ4qnB23KGJCO5hprhO8Q0nV06V21nhRQenX7+tzLLq+f1WlrKrCkn
pH9TWXKxsdGGZH/939yA8A+EDiNQmj7sjexku+HgdHHiQFU8AeG+Rpnlaze67qMRPkrZHeObqC8C
CBuYZ+K5iCziiiqPlaCRzwXzzXWtSyKMC1SbbDjl6hKq4J6W+t1tRP0QP8izcAmj6twywW0zUoB8
086sNCK7XAJdjsRvSKE+zgutbW1NONt00vO2HYkFWUSCv+GXjVNt1j2wi0BqkeA/QYcKR/yXy/2u
b+XclQZqb8vYk9rgOaFRPkiTUMvUW3lOnTwJHR+lLgmOO9Ormk2DeGuGmI9rWQXLO+27cd3Mxmxb
UzFXp1XIkYR44CDeoz5bQzZfS4P8YkNE89wiTWSUBnHCtdBLvVDW0naNdZQt0YZaJogH+C4y5o9+
jN9u7InrmjZri5whIHA1odoEe9OwLAprcMS2SCKAzknmsuUqydT8AUjC3HeNVV8mNlIbl8LI3hXg
QGECCTmcCb5ExjAwGkPl9Mtn7VAED9/vbHUjmTYnE6SxgQl7VxJIfIcnNuz5QCwX6YicjrzuSffG
0O5NHnIJv0qdjE27fhLOzgzbc52QYJsBvM/ScW8J03UFQm0y9WGy8/e1It7pZ5xuePVKFMbJuS+E
/w7Bg55Kak1y80MHmqW/pILTldNHju2mD029gvZWjbHg3mZmOZUjtYLblxQTdPJEX3k1ZLm/j1sj
OnDnfeKhNXCiCKcMv0BcwP2cNMCfCo5JTDauVf72WIK16TWDBiM2lUFwFwqXCYBUqL//kL7Xrwb5
sgmo3vnGpbx5SVuxNhgNEmJVVhsEKtRWgB56se3da+RJPKWHaeBXuP8JI4yQSzzCPFy2Hkp/UtNX
YwbbiiVHcPKYIbmiTkDABfkz/jV3Y3gq0cNDO4i6L72JgDrFcxOAfBmrRY6tizDyOp/EuFLXaKHf
2SucNjOV0egod6it6N7RAd7Vv9BBfiAOFiNIKERSfyHQFn3+2yq67jALQ/CgP6v/T6LiUtPc45Eg
DP+XLEqDlu8TOsBNG8itC8VhF6dv5kR3qpkJAioD79DE+oPqbvn87gKIomYfndKrnk6Y1CfygPwR
Yfvv8lbgu5+4wAeMZ088WLqGDCkYqIGRVMXgGZOIjgSHFv58YYi6dHdd9m6eyYN7qDbdyB1UDDjm
v3bZ24iNxv07aZX9UOoZXqAh8wrldihfnOoNYC8pJYmcMkJbH1M1bM6rysuudIMFiREj+AEWD5ll
7+k8Kr7E3iHXwBAdNWmeT1Z2fdu7/Nf9yt+cZgwX4UE7VgPb73rM9oOjlkPOWnLarS27A68TjY7x
9vF/2KKM8RavnPriW8oLe7rf6jnkdBXK9CJZQOOFrG8gnvmmE35/49y1HinBnPTVCT4eXTptGoZG
xnQShPG5OFSfTxkSpWlDTNwDaLVP4NBbcQex/PwXIW0lyfF1/8kAIchoRxRwFUjxkHfMoy6hh7+Q
k0xd0x88pbUHhMZKhoMrItb2goyNh+BZDlIqa/wWoCkt7DWLZsidxi5Zm+pPzsSzak7dyQWjz5Pb
b0VhXZCWNWOCD8gFTi8TMC6nYVK6sJRseUZjvxyHwIF7kq5Th93RIEJn6fAmRu+eua3wL0oMDzNl
uJ9v/w0lCvfpgyU6VZ37gpyC58RYMTWIZIFixUNnBqN0Fd6XXxvCVIyQSKxVFjCBC6I0s6beeVlI
06v5DRc7UX3ly/o2g0ZqKwUxo4ijE+8JW8odToJhYGxZiis5LprvFmh1O1GxVaLflQoylU4EMO74
K0+qu5i7T4jXIS/2lgopXzWa3PJ4mrgm0d7SIFim2mCbbYUAuIFD/PvdwPS8HxAsVB1iQbubDBFu
Ug9mctb7WMg8dFpZc3Fevyu+fosdTa9LJJ4UrK1SYYq1QWSt5KNdzo2/KDItkAWIE+EWMUeBJ4hi
84p91JkQIsfW9vRva6S+pipTPWoDeFgBgkONIOPLUvcFlcFpZaP6PBAsmHefz2f5nwq3tmomfGMa
a2YVXiSrg4GxrbhBjiyJE5AixQ8JQDEo2H4u/VQwlAJ5twgMfssLdLsB8Xl2oebhbouPMtXdwlhi
TkZyzikBEKU7qICRV6+HrvR6l/TfKxOL2cYg5KbEwyK2A7HQJzryQ7Qts7RSrz8SfgkgceYEgedI
4GnwH0KmTqCd5vYhWoykSUP0Pz5CKfxLAzUo2z3k0j8akxQ8kC4halOLAXalTbtRPYZr5WCcSRcw
R0uxCjWybjLcMtVn0AObjR8B6hufI/a+e/bnWrhHXZUAeLKTp/l5ORiZYSi99EKU4oCdvUvDPLlp
fyJYsYyTBxq+OTxET1/EVW4FSM4kThL0uFoZ8zo02m0GejHwPj65T/lWup06atwXEY+QRVym7lfB
2knWwZkErfzN9zT5Aldq0JpRrLjDm13/PwxeyQwi/FtQkDqGuhnylOcQg+JLnHXjTUVVx5EE8Enq
Lvl2U1jUJmW0eyCC26UG3iJOr2e0UqdhX1v2rR2BCSZZUPvsarKYNYaElCRM+b5wCGasmD/QVIxi
THtjisKLhV9nUu1mfHa1H4DLQiQ3NfyI0Adi3iXwpFKu5RSdl8uUBBCI842txe33NNCXJ+aGQ+B2
W7aVU8cUQ0vfceoaBRHzOXLrxPY5UnV+kXojRjmH9N2mVEzRxU7iZJ25JzBSdFWm5bS723HHu/vu
H344yQJASeedBWq5RXvBl9bJp1QIfz8OdBLeLFVKxrgpPTRMDTSkjX6De54wAYFbMroSOX5lGIit
1vuRvH8iBDsPoBKkVvGGBEjy7d+f4xFl+V6FownmGw4wD823U2x+2LAXTmS/OVfEwm7SGkMJ3hho
BbsSiuwJw6U1ybRe77OpvkIrmrcHpc9PhQk9ZEmGMOqSp3K3rWotKyWA9AOYEIyzvpEL406sSDVj
0iD2Ts3R8qTpfYslQlxKWco61cFSrriYiKHdoPIFE0G4buVgohFVfFZVEkTzUIWQSoUsWHXgveKH
wWy+J6bLZSJEoWOnGY0MD8IdqIKY8tlske2bu7cd8pct+TJuA+6aU/yQU4V74r2DL5qOXZDgbvp+
1RpNhLy4WRq2foBI8wzU7I50S+421QyU+UR8xutmhhPpN7AkvlIZPoYBn/CUd7Rz7q1MU53ysI9B
PHEU0IiMIsqGiFXjCGaMA7VH6JMS7+m494cKe3K7TE1gEnoploDnRRPnvvmtfO/CknBrB0fnf+FG
3bifBK/ZqWlbJIvH/aL8/eEyNoXOerI6Pis+qlW3rsa5OzseKFL8sjU7uAXuAvXnzqmbAbBHukFB
92voyk41TL3ggcOGvpgAZnNQ9z/SyFgh3Vg8YqqYfq+RPHAS3QL/dzAXGiHCFyas9utekrJMSlKe
1Xndo6MrhiXCoeLPetfOgGf0I3favEssyA5BjviL4iYodKh4Kno7BlwcbDHFes2PB49N10Xum0UF
g86Sy0x3jDqKBPjc2RsNHOeapYn2mUdXITO+MlX/pjJ/+jr5HpDXYq6TNuVE+9Da/9o3+s+61zF1
4OC9LqBaeGluFIqkh2EUyxHopgLqJSnoKx/HMCP7G3CgAR7s6gtc6Tp5Uc5VEUPzTk0g2XyQdiba
t59F1oLmludbeewPB3lIdD2vqqQmgTYp2lex0gPtm1O4gVM+8xDtAmBTv0ZTnbmnIs7Yf6aU+EIF
9to/8jMpVozTVaOPfRw2SX3StRsmEqgnt3j8G/sfxUPTG7yAPyRVho83SgIFL2HkudinDJJNmWNa
m4+Ifgpi5TYcnVQNgEyDQmlheQrKWPmFYu5aA7edN8g24lMdyrdBAlr4Uu0yJC9Yk14O4EZ0d72L
hKhvqUH+1i4QEfyscn7nLJHUIV9k3vv9qmkCSB0LAaVWeYGfVQ8ktqwzj8hRf5IqP5wHqU+UXnKE
Eu2xwqtSwPYAPy9Wh6Oz2eQkMsK2EhWxfI4O8ckXUMBXRmGwoaxXnhch/oHnJ6n13s8y44mbZobL
fikAT9UC+fZD6dqawa7WAgjgzFwZWtIPLIRdsLSw1Y4qd4jaKWBn8jXrB62/8Mv1eYJbyZGrIb13
xSN5sNhLt4TPx7eIbFsTT2vhbR3QYVif51W6/A0NxMCexesOdW0v/jg1RGXcLh+RcyB56+V/fLrS
TAJJyrY+uARELkSh3DRsLtB5n4y4e84Qe61SZHwoTMlGVq2lo6C7OEpArcEGvfvVNLpeF/wZHZ8+
oA+3VMHtCEMI58zgO4fPKsK5026/OqpasuqqF+CIARL3XfCbg47JDlDnZlnbwlKjqx41Aompsn3S
HHKiRZJPvNZnLlsDmg/7TLXcU8CWqt7+ujr/3GFxiwXkssKPq3e1EcCe7+r8oVAe6LK5StPh+hwu
3SrmPwBIvD4qA3s2rCZIPcZJ1xPySCeqrmJlG0X9qvD52SXEa7/qe4EWZbNp5RnXB0fTqmcpOZBc
pKc6qt9pM28j6AYLdLdLjkX2g+kX03M8kFVMzPNquSTb4eOQYBnodAN7g0oCXRAD0UzNUsXHEX3i
553ZigsurmFn1sIKsqgBHEe0UTLwoj5U2NoQBWUKytgRIzSXb4jSWJruAuCW1mawLJWo4TFh/PHC
hPPSTMEvnCuYB1eXch60qLQT9EUeJu6Wx7vlZ/yhm61AC6z6MoCnUsWgYGRhezKR0UYLyHApYdjh
ur1u0kQldQaYlLFX0FLiFjde4keHvyvLn7pEesqIB1RFFUn7siC7ywzRfQawzT3w+x7cvjoI9xMh
30A9zELMZeidvCAXMbPXi7oNq8A1BoRg/G8Eyfenju6xNMbT3/Gx5Uq70EJt9O15zxv3/gge+U1w
AtdRHe9yWL1s5IQ6Y2RPWL58+AmWlnwMeBDJqVj//Z1pppo34Dyj0xr6NbSf8281THqau9+VXUQ7
N50Js7Q/6iIV3TWSe5Lao7bbekhjLqowIMZVoyAW4tj6ylMbWUoGlzrora2crBGRVjZaKQ8Hfcl7
g+aP7f7uGiKuWKHAbOBbWY2ykegQOSxZCKY1xrZSLMEqDmtHr/dSROvzW73Vh26ESL92QEvnoefC
L7m1a9jc0o8A/uIkdYRp+EcZpm+uB1vArKWwsYW2vdmZaXtjNCFFhX8+y9/zDToa7wB4kB7D9oMi
Wr1aLscc2ydv5qdeiLLJ63sBH2gZQMFcwu7oqZEc9o43n7jC8XSYDnQ9BqqQCrtV+IZb1pXzG6Hp
DpFZXY/sbNGgRFOhuGXZz2NOCi+ttqQlsab6AHf5D1Cmfy4lpTN/+d9+av3jYp2H6xKMFlu29PoK
OzJQ9TNieZp0VxvyAiP8dvROiw7n7Cr+/DnTOiBDz42kaRqU/4bPHaazlmL5QIKJ/mId59mPL12e
Kn7+5xfyoSKqywPzvaXjW3REaFU/ilBl7Pglt8cyBcEPl+5WPpQ5NeReOUfwievmAN0QHk3dnjyO
eVO0t03Zsf4rAY9CWMqLobYQ8P17bRTKiojQQc71Ef6CM/L1VWTp3D2xI2unk+X+FyOh9yt/IYZM
HTZr18LDLzAhz5PvlITxQGxYCKyYmBBSVM+YRttWMAvQ1eKy1nIxDo5ZnW3ZEtzIu0EbbCcTXCqN
npl6jYSwJpmLlbOQey4SZx8wPWwWYoMy4ZW8D04LgC0RS7R6pIGu4+TUH1IfylVNr+A+B0BHPJix
UwjzLoL37y7PLLOlTu+iV9VDiKlH/1yZX+7KoMxkJUuBYHXa1NUIo59F1cJKpN3BVsMDfKSJ9EwL
X6npJVicnu8chrKslLuXd32JSw6Y29vRcXDXLT7R37L3EifT3cixtvn/zXY/wiRlPTAWPmiwdByD
gnqjRGR/PKojD79w7U/y42cd+fv5LgAbgsPhjmTj5vbl6TTVGsOkr3VgwLJbfmbJHtsUJ0q9sh4J
6QytEq3L2wcopHh6uzf7BwdvIYXc7yNicluArbjtez649MZerrncb3wr7hSRSroH65zrJL6l5O+E
QTa+V9zpnJylH5YeoGL4kk9gp0soUukVa+xBp+GHI216A0wQkm+u4eUHjRj6KU2OD8QSLuv0+Ld3
zaQhunmkaJKbs7LVNx7H+QntoGx5ri8ZOd5GzmiWVdLxM4axNnoLUtpa58CyJKfI30cPobkfhueU
/2/dJLbHwJBAAgg2smwjMhC+9Qwtx9rOMt1yP59zmcgTTcVj8APni+m/9ScfqJVM9VRdaobWlwIJ
K0rfC+cOuo45RvWpj1DcFJGzPIxUT4NZbesVhu65BVOSB3NEg0GI+ix8Dy1Yxm+HkPtJFt2KXAsA
FzW0wKn+7nplzjAXqnACOeggHGXLQ1V8JbfiQzqsVJTR0ugCTGk0+bOX9u+xpFsnCUaH/Q3fi7i6
dcsGdLz5ZCKdWvz75KDhDvPudqucUSDuKJsxee5rIaMDGhlPWKW04RvJlJx8N/cSB0gQWz0+qsZW
eHX8qp01eK50X+/ZdsGT+bmIYAN7ia+CYKmTE5Axic+8kCkEWfi5F+cP3vm3RWjCzxCH/Mv2JDmm
g/pML9b7z2Iv1mbnhRjm6Gd8v961SsbpOd4GICDGUNlmPi/Tpg5TZJEA7GUqz/mofBKneTgV4cya
1LztduRc5VjWfLjVfJd4LCL1JlhCTp93D/6xUr+K1BqI4Md+lh8We1Z7FAJY/UM+XUYSl86vUf5Y
RiymDY0YKtEzN/IrH9r6N0esPGdp2ET4nc7Rr7nAjuCcYOdMr5shvknjOTJKXXEteFOYQ7m5FMTb
HGwPpoe+blBgCwLvgWjUEKKSCrns0WpJKtg3xGGNNFnjG+8refB+vRKsuClnQFBXnrQRwro4oGz2
bGPwV7wwIsTXf6hbD1f3rsliGsC/+im1i+NmvsLz851LiqUez2ADC8aP0Wdb/+w+vRksDIU/dyFG
Tbr6/3mY5xngH8tISJjErjs5nFgtgl8Xa8RKd2GjU/CBCWEmWzG/et66ztUKYtKhD5+O4FWepqB9
gKJacJSBLsRn/oKWeN3SzbXp4ZpEmA2uJOAGlraionCrj+x/MySKmeMkxzO3iWlrjGpqyScyRbWp
0YQHJ1SVAVsdEl5CL5djSxPquAzvvSbbnBBtiBNdwZuNor3bd6+xHUrhntr2UDeiEX/zBN+XHNjv
e5UOQipNwU3MfaQSzMQCUZaXyiUJTQVPTDGdoVlr+yrwB0csu4rheIGjYQd20ruW6e6pIeLnicRd
okmAMnnEDKujEmw597tLiSvdwvspvf+CqYsdCmNj6XpDwpH0IgZs1qhgIln38qiRwnThcG5Ttycb
L1tdjla/dqpI4OgmRFBF//UckMKBYJUH5+Q+BNLMw6ah/wn85uYUNZ+ZrIm10qsXaxplLXa832yH
qSTn/vjau9H5j6PVMW3peBnGadZ9SZECX3yxrVGPzxO+60dqSCywHgsn8Yrbx4lL+5PjRYKFoatt
rhUpCjSaC9D5HUFuZ9TJZsHTLnGNRub4ORwnRrbLb1p1F1U7q63ibVaPGPnaayjCEuHcvq2H31WT
N0d04K74of215EGrC1wBqGNjMwl+WFUV+5eJU/pFS0QOFO3vyfA+Fso9afdvNWxGD0gmvpPFiJz/
kMC64IUg5i1QPHVuuY+X3OGFh1n/Dqs6LvMypZocC+yJfz/2fOcFrS0H3zxXLI3DdVzFwEpfwtzb
gYbBRugQsh5s6nWGfDNc2vO6vgq6S+c1sISXWAwPXsnJX0Thwm0AJg7RaxJdgDCBFSTj88LXGoj1
yphGfqxRf/Q7nJPOYumwmzg3Kv1G39BD7hh8tLO4lct5EmUi6jbpsu2IqS3uC/RTORfwiQh46wLJ
8b+8Qj+9h6Kk18OVk8fCj1xgfaiCZzGLoCIzuwzbiqirjVVNS0C58ofJ44M8LTz6L1jAjP51oXjQ
gl1tfMvKcuQDs0ng/gM+/6x3zvpP2CQCtKcl7om05PubegZn/+P/JbGL+K/oz/6i4gzX6QmVfORx
RpcDY9DTJD/nVnhU0N8qKGz4exlzFz8SoMr7eAq7k3OugnWinjpwZN1M9Y/1Wy2H2AcYZopJor/V
v0bD9zeggGENQV0GixyWkY94jM0omMEHUo1vtfIsbhR6rfpXkgtpeGmOnkrtuMjbc+w6pK3YgpdV
N57vaLvzCMf6OT9Dx60A4VW4b4Jg2BRxb0k4cqOFsdeWl1yw0JqQ9PAXNw0rtpygulvDr9WL4Qrq
XKIPePe+HcC3jQenaf1paI4n2Pnm89kf67l+qd6FFGvjTZpGOPOO5XtozQ03PuYW5LqnrjNVxAmy
Aoa/8aFop1BUMWk/P+ErsRGy8a8wWI1hZP/A3TAFa3ghHXVRVDpkN3SL+hbo3TJ6fsEdWIpdiiuB
QQ9YAUk/zIciy81op/Hhihpc8vGFJZsL8G77qVFUS1LTJSX5ZbzdozfpDnciE70Ia6EIqbmhtsrX
FuXLsPbl7pw4WAaMHYjfJ8S9/8bg/o8AgAwrYfMJOupbadoPitFpF8n9vYxYyPaF2go9vVv7eBRB
2KPecC6LKF8q9TdJvgXbPLx3Dr8VHjdVbY+V+Uaz5kF+qOuVtzyl3QKRG7cEe66pEhBJxIya56Wh
cthqw5jUsXwuS3fjIWM+/h0O34TelLX173qvsZtff5ts+MaYsj36g72LBPV21N6NO8/EXQlRdExh
KFUwmI2g399JvPKRA+cZhPqSbSmMwUszwPt2BE7x6U8WSUKJCLmhtELFe5LuzU1gIgc5fH47eAy3
K1W3Gd6DEE+rqE6M0Ikkk+nntooILz4itbeXCuyfUl0H+4iC9C3pJ2KDcwTGtR3cIZYXe0kK4Zoi
POMQa+mw+z8sQ3m36R1GUh3HlP1O2bzbOiN1UbYwkXQxz2lx0BEKS1GD37oYsikL0z70QpvodTcb
dSOjRql2KfuhYhVLcr8sgFJIoKq3YQ65AVGCWyZ1zx8VDtAjjESWEnB5TclK6eMQQBx+UCwsQVZr
4jG/7zjMXj/05qeRCIjz7AFLfxtd9YAv/UguSeOpG0CH758wPQPbJq0R9/HSoQ+MYTjyYKjS12B8
dhe1EUZvBOaIQE/r3K6Me56FIa1Wx03D6nhVdRM2y4SOonJ4O6W3gmuMwvmkrgvyQO8SDfMjGesn
K8axW5ZidGaWEBocHaJWJ7M60BiroT5UjmS6oZUeBt9m3G6qb6MUsotMJGrp2NGXuWXVfp/Y5hUQ
XD+uNALulqyOm71Fcth4eAHzUS7zFfsgnHrtJMuJOFw0j0Gfjmra8H4IsB9G7d/853qlVbTxTfY6
Xoh5BJFrDTYqYjagARXx4YhwbArhZk9lTycfJn2v5X900eNAADT4OkeyRvbX2j/soCH2WQADAdIR
UU/yAx490YHoM/HqVQVjEOQhF6xrNpdSfiekWW7ir5YyWn222A1/TkSn1/0dIROFSEU1S4rgamBr
R1TWFiksxatR1AoFl9mrB5W5UCezU+3g8THnfQSHDdHpFJcD1jegBgM+hLZL5CfwCXhp0gqjepG7
wDkwOY9lQCizccdh+hOP+kAxNiXdJMF0vfgbzE2SsdITFpHic3mrnX0r3vNo5j9p5bzSCliPhACD
EuIuOto46Oyn8ejHljNW2YR4XRsABQ9ETLHdprj8Oda4PBp8WD7S4wr5GwQ4bseD5mo0TASf1Wtt
WQgXbZVHnbYHgxL1+oKodvpXijTY3aNF3kPWS41aBS5hwrIBNA/wtzLaY/UQibgGjbR8zNO7HNAt
J6heXvNBwBC+ncBZ7uGKWP5wQCZyuoNQ8LUkSilDEsXR//3HWIsib1IXdIurES50TV4LnqhiZpvf
u+eYw2GkkN0fz0B6j6SL70sXr2h5xuAFcrWgj4gv+HsEkh4ZYECpR0lYMbGpDqk34dzm6071HgbA
fYD/UvIQF/0qOCxTl4tsM4ZCQnw/f8S9n6Gj3AW+XEpdlHy1+akdXQx2OXIK8Enmy4fsS5hb/P1O
nGCNgmuonoFExj/+xXLT6aBs/6lX2Dd+I2VWlPYi6gTsm8IOQoDdy4T098dbMH5PAnf3BXv5hkR4
BSAMYp1N4/e3S9c33fAnrvbb6UnF+DBCS7rCK/2uy5bmp9aN7UopOmOHY1PuJCoLBWlf7ECFUJ4R
zul35wxoVekM/oXyOw/7qcQ2kcWPvUMZAMNKHCr+7vDvewFgvl5XOgUjxbGvJmtRGpfVOu9DD0m5
937xgq6rPbHAIC5ZYYgoof9KywOVo7syrktoKbgZjSh45XzUsg2whaYBocERWVf8VgHGz0NT/cQI
KmaeqzolgLPfLpfAFLso+UNCUCWAsz+W1gKy/nTbGTtoAzioImLGWIeS4l2XjNuiQZezYzUnK0yi
JlxaAC9BHc+3f3Cy5i0BavtETJvw2vuUe8Lc9f5Re3SDrGvrZ04bah1EMujinE89Q742QKOXNd3D
hCmKA31g1XQcTQyQLS8Por/ocUmGkmNkJsWw+gXd2sU4E/3a1eXICNoorCoCDdOpnPIdMTNmVbbb
gv07MxDXxPxZoOe/63hbnORzryBp/QCg7NQIaQl8cmF5Q58ZO+dnVaQwF/VM0k5wsf1FtKlCZvm0
QijPOQbe30L2+jEebntvD0/7lykDP1hA0emP85K8JAz8SAN0jFkCKsHoxMvw8tbB7QK6pqb0P2DE
PIYJ08P59eu36qI1TuY9QJeHlVWloDrHu9lLx8/z0i/WG+zlUiSFeH+8WE+obeMhvm4zOKqm2Wga
40usX3GiSiiIUZAX+qe53SCsnxipeGxVJ48ZQV0XzZFnqEccYT6RDc5kQxquKA888cO3yT+O8sZG
wx2HGOUSfmVIZVKpBze8bLNjw56QvKutsFJ8blN9G9VIrkaWsR6Eq9dE3UzsC9u4fzDKF5bPpdnn
n4BL9Sgt+mPn1KcXEHan4tpeAP/lXJfkjUqHs7DpVzOebQwYjlcRkFVygZIB3kiLZ/8rl7c5QG3p
2P2JcQPc+NT18lgThd7yRRaefiVUKZsCcast5o66ukmGIoJEvQ6Rg1GJrU4jwtsVGTte/bI9SF3t
OCJ0jyIdqtgf7/P65M3zolnDTQi4Uc/+QSC1p7KRFmgS9oj31puxBiLa5Druq+OklMYrrpVddEuF
tH20X2EGUclkZGXS4LKeeiiKN7vLc8XQImb+JJjR7WB00PG3Yj5+CrvdL9PXiqfyJebsL9vTed/+
cRECf5w9kc8epsa/f/FLBCp/z4WTNDGZeOClNZsLFe7AAfid4jMbG/gCUEeGV28Za80iZGMhAeMA
M4M70IX/kxNrmo7Nz4b+VOC/z2FCuFFRZ4juAK9/wMdx6oBNfqYHZ5ZxM6HnzJnXnq6F3Yi4ep+t
Hh0NIlxVjRKJUZ8BrVSL+UDtnhLkldKuQjFoghPZASJycUawIVnIDjHJzFozs7ZhEY1iX7A6Dahs
RdxnZbnuuumtaEWSs1p3y7Qn/z+DqfP2ZgdmqVy19Z/LxfbKhFZK6fC9bptBi7FIVDx61RsqvcfV
PKzq8PuqK2Qi1UuNy7HEKijqstDei3U2getm0LW5CoNJHUqOe0pS4gNtMyCWdGHT2lZ+EUt03oHc
UFi5k5aJjIdsYh0n2xlqOgxFc1MoooNkCjgN1i5n32SIEjfPEEbHMBeRo8FNe3EfYtGQdNqjnZn4
gFnWeYYu61N/bFBhjYYnChxjA33/3iBNFXHLcFiduyw6sY0cKimEx3fzgRbW0AJq9xxUrISfXVcJ
/Q9N4IPAAc/UMAfBxVBGIW7svoAP1YZpSiVH1Sx5WeuG1J/DqI9OMB0JntO2WI6xngdWx1WzfNxj
rnQIiSA++IA+dZXokOUGSZEapBFg1qILYpSpTtf+96Bxouz8qXapxAsUefcPyuH9limgh5uIGxeM
WGFgsj8Zg5etbYkb/tyiNUxoxrMoAynVEku/RXi3qQi8vtn/6qpxE9LxfrWHW2nQoLvAAbbjUS0p
trua3BLTHWfCLttbs9j6H/QB7nP7r7smSUazwwfJ6Gzr884wcMgiunJfANXChQM/7kFiPhlcs8Md
15A4/VvwgytPVE8F9tjMizh6kUwhGEmUZePWBhb0HDkrPs/4BcW7dIgfcFFDzbzPjf4K/NSGOHDy
WW34D50BJ1S7FoWeYHV9zUiztJmLocb1dBc1TyHbcJ7670oJc3YcbgI4RyOJTifcQORO+skRRqCh
yGybABylBw88gC8hyCfJ7fAzc/ubYXV1h0Xf7XzySqp+CJaY4ojpzzftb9sYkHYgQxW6khvtRiYm
Wep+KURw+dNTJvTXjhbCrzvLwq0hcCrKTfDrP9NKqyuBapbO2TOYf08YHz0Xd8Ef+Kr3nyFhapcz
N/pbxcBmIphj0DxNsThcXLjjD3aUGG51nhcz69/YaXWdkzYlk/tvDY3YKU2J6nbMq3tV2DmUFcmw
Y5GIaaxk8aLBw0pB5Ig7HOVdMKcr+ADWqoU9WTIo3WT7GxlM4gvx1y4338Dr8OfL/LtfAyUMg2np
gqbYFkBUNpkw8QuZO4huiiDWZabnyqJNRh0Twgfl9ivbxg0n4ZUHctcy688m7EXrTs1AGJjaCtLZ
j6L5lCanEhm77e2xcmaOVf8KSr4dEiFQGwM9FKxYFChvp53eRfV1/N9k84RfhRXbR4o28Wl/6jFy
f0XbXvSLzGLR30UNtQ74/ORyEx+GBR5u3GDRrjpnu8oGsHC3LCmZG4+JpvzVg9fltlbHHIEIIt3g
D8vGdtdIou+LgwszgfbWD6hFtxGMOnRRfneM6WhbYE+kSCn4Kf1ZTqoUNL7M7bi7g9RadRNrWKOk
rzEsajEb6iSdrgQyvlYQTIS1srPiWg+C/rhscyWIstFLo4PB2xUlHNb4WFaGYwaFjQJY6lj3y3GY
T9pY9MtxP1zn0fvdGCu/0DBApsjLXbkTbhMTROPVWa8l1WOJYh1vGzuRGqpSTaBRFQG/Z+kcFeO7
Z0V3i03B9cMNuxiJeejuo0X+LdT6kEWDwR1I5SxkpCh90ALErzh7w8MAAorfiwo9TX2xZRh9UelR
CZ9bsDEqUGEoEA8/LfS7vve4kdHNenvvPZYPXRAA6HyPc8thhr6nhSFtmyo1UsxAmNTe9aBTT/7j
tcz8umh8iOZHENX8tRZvbKYpiB0c2VtaTOF/T24Ch9R6GerC4Rx+m3xgWeCrQagthE8++EqJu35Y
Qr3qDAH+axIpd6+Jt1gM/Lf/wVwdOojFoetVRjkOtJ2m+DeuIsabF7efAXLPWlg8h4p7b2+eOWIl
LrtJT50Wi7wapYook654HM0vbNETPGqNd7S5vTWXTtzJOHz/ywmQx3mKkKy6oSl6AKLmGVc4dckC
hGHuBa9da94LXez8NG9Fz0WP2ufuZT4zvPynuRo7EeCDeb5RB4hVm/C7h5JVksZalYP3EXSxsMvc
cYKYJTctRBprm6MeiCnEgWfngeTXmblsETw6JJ9tO7jA8afk7a32a274Toof83ZAYdPjQ+0GPw5d
B00tgtIuPqX3wwPUsbKTP2VgyzDF8hcfgDnHMYNP1hyldCWXZCyQLHMv9qZN8ZWi9GRO5KuuYulX
B8FsHJqLqGSgcdxuInUrkCYMBLqQuFj+zE6ClSYmUEBfCDMKobhYHNP2wV/4dg7Kmq9IzDTckufA
WgHmFNNZarKdd9bh2zuAVZ72MQ5/lmw/lnEZrG9opm9/FU46vYJm0CGAuR31Fn3tBufvHjKgrSVw
9AM5YPG74H1bNlsF1tldvGCM7ssq0hXHBcgFZub6pReZ0Vyu4hCIFseF+jqrm7C+OKXnIuGEBxUb
UnnRc37hlmv7/9QVf/f8rPRrD8Z4NzCiacQTgkSKjhSXDfG0VbbRgK0X8GHu6kuuo3gu2oXcSxjW
XuXbg7jwF4Bvn9d1FR1aaHXm/kEyB2p4PHATx/RGa00Z08uBJt6SyA1h+HMQo7ZW8vuMtchCup0R
rGjnykNf5SH2V3nnp7lUfY5CggjPhrrQEmZ1z3mEIL0z+iQgDr3q4N/YJkU3QGr3MR8f3h6rwydR
yV+RCLgXUkoVC9h2tYKaTpbZQwnvh0xyN2a6cXchJe1b8iw/xbm6rIYbUEAOCCSyLb4CoiWSUTip
52Gc4Ixv/DmG4WaR1nRbhsOm5hPEfBSuqDF8SATOl+fm/9/Axqi0kmdRJKbN70uulvN4pbyZB9PQ
83GepjNKZTwreJsm+V7cJTYNeAjR0on5dQMYebs4Jhp42AweQwM+5YGK+6RBx3OtQ0KvJ29yVabH
9GCW3wCR1lSgBgFdApJhMDyGOuSenfq5Lny3MHFX7KqGlO1r8uCkD11UBRYUeuAH1X59GHNhqDiR
UR7oLTGz55b2E77lVZ0hchzVl26jcPGM4euANY+T55Cow8Ds6YLCwG8IZjBkZCdLv05iAwHqRVSa
Z7EkdlRblMdNOfRCQPGHCphz1GVw3Hr6xklH0qz39lD1JZp8XxDh398CcjFUc7pMuz5Ok4VBQa95
cjYsaaJbD9Dt0+abi+4fJB82FHu+UEUs2pwRp48K/2c3kED4n31vawu75l0/tuKzYK/ze3cP8n+Q
GDu3+ZZgc8qKaTkPQR1ZNvmFUOXM6/w7BbsTDRrU4LwedNckJvMn19Hz/z9UAfhEXLrg3whcfJfD
5DTL+FdyEj5NSePcjJWb4ALJne4TzROcTGEWLL+2489+8jXzeUlPlGdh+N/zzD8yfymrz+dA7bIV
isMnk+1tvXf3DuCtl2YLBx/IEy8hkSFkeRx6+kALPKcTw9Vh18PnaKi5j0vyAbE9UAKfktz+E1mS
oX5PiEMszbEZs5Vp96xxlkBlOS7T1nyvkxE40TJFmtALzq4LKb6FZ2/EjH5xQRcVd3Il+wq/t115
BRydA9DR/SA2vwiknxRoNbvYDNnhQdovWO0jyVzgCRaSCgl9dYmmMU0IKo5dWYYvGedDXskvBUcl
P5CbCi2QAZuC40qrkiy83VPKefXxg3zyad025gZvUeaDIe6ad2x/MmbiPs1qN4DN879vN9msKjpn
VwQf1U9PfBMVl10LWR/CxkTNLyuYE8pUOF7U0jvM3k8y3cPHL2K9g6A5uVny5MVzaQUUGzFl686l
rUP4njDKegL3l7WFRKRVhewZrK3RyZTENQZqJ5IjCiMAJ7XUckuGvwbxJexdwaMmOhoSri+hB0gM
ikAP1NJjvvjodZXk1aY6sV+L3QfGP83EhWJLFsm2AQ92JhLh7nhgOrnGJ6+UTCmf/yUUW5dDm7zZ
dhLtYFBU8W/ZboMtC7Txx4TQJi5iD/vTMO0j+J0u6sUuw/GumtuTl9v0FdqvcN+9frYMiPsHbN7V
WBy4CtqKcs+EaZ2DEdagHqb3pzXsTDpKMXjlEgUrdNxuir8PqNdPj7lRF8ZS5NMHpQmuk5hL7Fxj
ko6eAn5cH9bBNHD92MXx//miGvw3HnJvOjfh2hEpVuhoTMz6kDrUt3jZgAWAfhwiB6tQkoWJy+2F
yKqD3NqlaD9b5TqrrOco4Bta/1++khmm5fFLrjppInIoDmArtXpD3ak7ltUbKwEJ21bEEbq4Pzdc
b20uMlCnwwjGiU7+34a+XhM3kkuPHMRbvMXfbFTzl/R5oZq+yi0kPmIyEigBxwW3veK4yYAXbn2L
O/Po7UgHhXYf0tq9/bAENQ7K6/9OyZ+RJZeEQLgtqa1fI+J9McjtrthoT/lwcnDOwoqCu+cLw+Hw
PZxZHUtb97/5RZZmL+1o5uJHNT68pKCRV2s7LHFfAbK8h8cB/odvPt+UMT3tdbq2OwLdHU6/k1yp
jlFEQP7x4Tp2QaY91bnVMh1rmLJBreHy8tzKMMzursvXw0uiJAvwO4hKHC6KJePoMqk/Cr0oBzE+
P6xBxnOLqMu1GopMooKsds1q3xqxp6tMwS8ZLpFLyyarm/SrYu2/daalFN/g+JfjgWaTRtO7LEnQ
G3BGYc6hp/nDWd8mx/XNmZBr3mRWhhLorMj5asudIS+S2z6ZxGvNPx3+miNMFQj62l1oxAyL7COk
j8pA0sUtWGM7XOs43zLeVaX7k1TeTUdMpdZg1EelYzJeOxvLrVMoFKfDUVTLylZ1anlYwenKeqcZ
2xZDRdPxq6Mqrkjrf33qu1TA2zXA7a9je8GG9k1+VaNNeTviBWrIeqPXh7ytt6lKY/3IZHMYISJI
taCCvjxIDSqYZM0stlkGWtuGKvUGQyHe8jJkHxa16yHrxFP6ylrUgWsbxRCAmQxAUuGaeh1zdL3g
Lj4D9T3PUb7g+Q/lJv+dsAKMgPsjh+rvW0zaZl0GGBId6pBFXhsA4A3qiQ+JNoGbvBzK3yx+4GGz
umq5wXcZD19cRFvnvebkEif+Dlm0IFQ96ytO0JjritGF6L7uwk8I7v+bRVuWHUKH1kfrzftK1prB
5Qq/wjPAJowkG5++BfX8bx+cJwMvqc5NzJoUUTcv7rOkavMFYJ0pJ8t7IsZw1jhntx068+cIpu3A
Bftbb+9MIIpHFVkt+Pa4ZGnd8tmfLG4uES7qF0LhQAwm5++BDk8t0P4lOaV4lrVfKQ8wHfMgliuL
FtCKBrOZ+IhOu1Zjox1u+DRv6cas/vogBctqIh7Q4LPoXLy1E5rQhyvwCYoY7I6uR7QMPHwjgYZ8
ji75WjlVwTT3g3UnBDVDaXTx/dqyS8iaXJpWpLzTWOcNeqBy0fSuunrwIoqsTL6eztoyJFz3eXs7
TnW9PczBht/yiaU5UnM54To9W/Qdm2NT8bJaJO65108t/kzFMoyQeV1kU6EVOyJoWFWgwDhk1Jgk
9tB+w1r32GD5gL+SWTIXXk5WkWVMpANhu+ItydE9Pr3NX/CWXZZfjt5yEZyl606pBwO+fNFkp87t
OOa8xOOCLmZdQfgFRb+v04IC3oZZHfhpbTlbFf28yPQ1caSBv+ox7j3ZAMtLo7qzlJDrG4KDljvf
zMxVj7wtBuMmdcqPgm3iQsYm7YN36Ug5s29H1hPOdrRp+8yfo3xgMKMIWBYPlAMu4caqs0om2rBb
QPROCHu55eeOaBZpqvNtHKuSJDX8rvshHMJa/rNe2s6YLGsJuPgv3nsLjmwb4BSNTP+I+SQGpqns
NgkJ+gFkURMOzNprhBY5pXyKi5yYc2zjxTRo5z7zxPWX2mY+zvGX3EblnupiC2lJxbd53BWDCcvQ
UzblgzgT2bsto44pewS3vGacyIr+CwiiGEqQ78fc1Mk4avkpRov+jLd33ntv3joe/q2wEasWoCzp
7gD5nYFE8VQqsMFYKoAlUS4oiznP3Lud9GEzO9mjVzYtzSbIvLB1/2loqD0CKGbWzMnak69VQiml
BhRPsHjGeAqyaMHBpAMuxxQ7pnimQ0HeQVHVgQTTCjaKlP8RaACeVvmBZCFwpGwiBgKeHLMfhk6j
fRktZUz/u8J5IOk5hgTHDP3qLO8892SRkMnyr1Wbxwf8mWaKQ2D8YHCJgH7ZuRC/Av8ievXZErG4
Kkofsv3s9LB0KoCwWEh97N7VmaPCyBuKvM9AolAbvG4S7jsRk0rKrovpoSqf2XO7jJi5f0Nap0Jl
7FCFcc5e7KCLCIGhNFnyO1u2iZwuk4ldyQC2Rfce0ZSB/NKjH2Sk5xRttmUEiiP8TxcJvuRDGi6n
Mgo5BSAKsdhkPp3jXrhhNZXYeVeA05k4gCjL9o4PSYaV2vHoVOc6TlK7xRjyEe7q5iKdy+C0Q5ev
//zB/ZKoq9rmiHPGlAbiu6PKhyP75msryczk2boov8VmD2ECA/LHlNJbklpNpQuTeI8ZAQ1IG87i
dq5Ge4RdILvC2XXVwT9SKD4sFkP0aA2iforyuKNoEhkwdFZsXVYRmyKn8Yl+5UGe/MJXEUXcLHmL
NBpzmpamEDc1cNEA51194EwhftBO79vNAnxIOvN0VdcjLyDiko6S8/tlBCKkzZS000CHwgJ2HoPh
xS/GZhRkn9zDGY6LXseaVyLySOM0GlD+pF2v5+RlJ+gZ/7xdzoCRjIAVzFRuSOLiocuA63Os2in6
h8jphsbJKYuPfdFHS8dCKE8C7+rI1EdMzlkG7evfqddSlSoujVaIReeWkMnmD7CBQYPBv9iUBSgW
dbqNbaUQ1Efmw/EW1Cq6PID12z5u39npit976pnGHKYpQokX4jB9zfofaDcX8qkPHFJTiYar15iJ
fULa6zOcJn/i+gh4NXQByPBRyOBJwhyMp9NuRdeAI5oOBrf6eIeYYJm+bdP3XieSqW6g2iSiGTW2
WZrLprk0V/51n1wLAsvGesXqNfWGup7NO9PiGUBrB8XAy8GbsgsmsVg/2V4x5eHHxYd4kn9vYNWB
TpsiWqNCG7BbbvW0ix3mkNuP9ONlJfz+fkRhyiyrmkVAYvaeYWS3LKB6RqW93ViZZXh6pguNxla2
9EpkVXXjDi+3CssgbIoJrfwgHVjF5MOTyOWU8FObqQFPUmeb8X0O6ab4UJh+yrpLNJtB0gZQbP7b
CDntJWCgVzXn6v18D0mOrByXoAcqUhKLX3LpAwLxPXvSx9IDvvbtXHOlBgeMmq/I9AbuPti61P74
RMg78zbhYU17r3OZuS9cJvV5a6UN0BqJNozsHlkKZ23M0nW/sPW9ZFITDHeOrnMXvTbM9mlxJF7y
Z/iB2dbrXmCJbdHZft3aUsx/J5YyLv46KRfkHTlxjmPLGx9iHgE6CQH98kBi8htZhQL+7GX1lHmt
YXR8ezsr/VXvPrkhVskIePe4tFMJsyn8G9n7JGz5Grz+yAoQzUHdVIr8oGUOH/YVx4+mlIl2ep6b
+wnq9HQ+s3XK+l3ekPghYKZ0ivn3zu0z0egui4hdlb7n24dn5ibBT4hMfuoG1+3E+zflkdbOfbSL
6il8A5qeVv+xhmpCOseZb7nmyDKaYyPELTGKZNIn+CFA6Ro31xPc0UwoYRvpqvAdfzjYuoE7H9mr
ItesuZdAT5t32WT90WbAl3vtFlNQdfKWFXtSnO33nEtaj5RF+VyDnx/u410llYCA+AXphKN+zK1K
vrDx4lDRN+L3/2QBGkL/5GTl7RAv8gsgD0rIiryK/SxbMkwrwvCuJnNnPHy6Az9y09nnKx5/5Of9
/LRW4xFGk/tZoN7HM+0P/uwc/pzz0d4n+hJXhOwOPCcelJlB8wNptp2nkURK98Z41CoD3tJSFE3o
BGbcS3ho08YhlKzVliBIMfC1jSswv5KDEEuTkq4gQDs0JA40F3/83WI93zxK++8j/uGheeuGQB8H
GNm3s2Gw7z1qMFDHRAGwT61ijYnvjkvS9z/qVL2OiDFLAnV8tMsXDobCyFHmRt4h+XIcYxtaGVJu
bSf+AtHpW+LOCv+J54NsqXfgZNKYj06iGzILmlgSk7TfhkSKppqiolRi3ZLjPIUTpoqis6sL9bzm
3Hjh6eJxt5kENKaT4uM0v4cqO5h7P9myy7k5Gd03jKS8yBKZGdKVYnSNiF4luYIkSDXSVhGGZouh
T7O60qMz7Dbtv6N4ZRo/m/CSebbcBL0LqipzzZyGVyZAT3qvWK5yJ4BNgdKuDKd/61GCOCXMR/vV
r9cuEeKv9KOe6QUWp33Z6Fi6S+wLttmLjBV4M8Va12ohS36KmGBRasUOjwXcUplVC+licOqGB7O1
aJY9B+j/tuZZvmA4iP/x+nWqBMn67LybInADGDiwA2IrNh4Wz9puRg6uo3PylaKus8Li/HkaT0Er
v8zvO7NGb3kxhHMVBCfbh69weXwbrh053fhuikj4B0+ZrR84i/4k34uGggHgGsQWsJ8f4Ouye2Pk
+P8Sb727fvaRJygRbwZxqe+noGnqOFk6AH50zPsbWksDaCKMwfLEhxHVp+UXJxUmhlHx/aEzFWad
Du5ylHl9q/CnkBQsqofUbxBmrJpQrH2biDfk1ZRjPNCSV4drZM+dmEbpUYHH7jBb1fPhpIUPaRys
N36cm0RBzwBtrUeekviny18BXYgQEGHC0e5Ns5c6AoREHvzAPYzEqx2cLVHpaXn4xBovrsU1Fwnz
BUcKHwjhPVSEDJqdWySyfzdSc4p3b1U9+tKSTf19dImKIp9cPSXha5eHKXsiIjUFdZeScGasJzfw
aNm8/T1v2jAsSdUP7VX3ob4EstStLRciJ41Ie5zzuJxwZ1gT0AYuSp8lMtPb/Rofn8yhkah4EGVW
uT8JKCgp4pXmQtfnPvWhY2og9wAZcMK6uJMa2iso8nCTb6erTlhGzqdNL/F2/bO2a1TY//blk0lD
hkQ1o/G5tk4TV7zyOxSdO3gQ2QQ5PxKHZDKaA4j5XZBtLGN3/u49eMeIIMPd+QUHFOSOSTsZaOMj
8XMl8Wx/kEKZ+thQp4DklY52zNpqhjj/DfIWTb0H3ECOhzC2or92LWLi0FDYpJKXebwHSIfkiIce
GASWukC/FakHSXILQUJ2WTGhehRYUy+FiTh/Fb6ghPNoV7uzsHJQaw48Yeir057ZvF5+m0+Lp/8I
2AJ+AbX5L9xi1lQylv6bN5FM8QyezgUE7XvjYgydkCJax34lHyqC63uUapoF3fIrKTILPuK+R6eW
olGwgkFq1JsioJU2Ub7AO+Sa0XlRxDsgwa3/caPiLnLokCktTKhltNDCMDtbBN/qVHfIwE1Qx05J
mUqYb48pVLBBod9t/n8AC2EXiMdgpcLqRMpY7pTsTazAH4qCo47C4pU8GN5Nm8utcb4wphSV9pru
impRxAbcRcUP1U4jBPsVtzngzaOVUQXM/ZNey8uEnJmbqfvH+2g7gPwsutDPhapbLAT0Z0fp+upw
Vq6xIG9793u73f+4xAEu4rJfrnI+7BTLuqbicyS7QAeryokXbbvpGObEoGNrZUqa3yMXdjttPAa0
HYhPlpe0ZeJ2VMmShPG0mo58rLdx0XLZ1Nsr6wI8hlw4YIcrQ6RKiTFj5x+cuLZFrEzy4fVD1SPN
NgTcsxsvTMDIDnGgs2f+JS5lGDy4HwFsE262TH/yPTv7tclEnry1kFBDF6JhkvzlQARZDvSwS7mY
Y7rx55Tib95V8Ii/AcierJv//oJvc4x9FJy8M9gmVMJhM5rSZpUUWDAnDcBTdO0MZOAl0yQXU1kw
0HvhF1XzjwHxQyhH0gmaVJEXjcQ7mC6+FjtZQh1KNGLH7/MreemG/8Lb9k7DpAOuUuHWFdYgHkrn
wSUS3Hx/ZorHbCFv6lLdmc2fgZvi7EMFjHHaefgpa576YA3NRJv0N74UGniUORpP752FMMEAmDVm
o84OC5gQZuEf5ggTvRnoTzJDqasqvuIsMza7qSatwsKnZuLzAb3ZxgTEtWlEj7g0tBwVcVZqvItI
fRSi0293jaknAO9R4OUz8RX4LhR3AKTbBWADfBHUbT0HitE/k7gNETkNIbOn4c01RV/0IbKh38W9
9Ws5Iza+2+T4qkdnBzEBfjcDzxPZcqWTs3Gv0lsJ2eWknp5ECrGPI6OWUEK+TNuTzXPh295es6/+
MR234bwI27eDwetm+2hJ+AzY4Bux0RxAAxrxUy5wB+ggD2bY0YuxyhedOzXoJma3NASU/KYQwi7N
Ro2s2DYM5DpWUjS4qsdJc5vkQWZhXaswbXXPb1CqaSdlz5mkpU5Fi1hF1/cNrtdDoqHrz+ke6BCV
R0sxQlcvABNWCEEYXhduTUmOqtOunEU/0Ve475i6XStX7wi/sWksPKnbl6Iywzgb/SCBsksVT81e
/pqv/zmRK6GMcFaYUJ0/7//uI0y0N08CfnlWBFnN+vGtu2jofvi9DOX2I2kDg50SEeQpqcgkRxOx
Dt2ItEmiASo+gd06cZYsNlG4GLi58l+CQ2Fb+ZsTBmrIxp5SFVkGCZu77q0EIUCC45LxmDxI7oaB
FT3RMwT+o1LogkLjPllV2VeTMtOeYPBVUZcLDwpuRYUXlSwwgdyrl/U2xwKVX85dSmVJ+cgaQ8iP
hC9xcJRGI1YU7AAnLf88F/8wr+lZl/9qkxdPXLVt7zmdCDJ4MsVJ1DTe8LdNlxMxD1GoR1M79nPV
kXYEyArbgsNXoaKI/bnNwxCDWr8hQ8MzHKW8yzsQ3DMFxflz2mR7pJyk3KxN0nsRGPJaFYv3VUu8
blIvrpk53Km0osCAGb0loFCdIsOtPGw76o7LtOGNUAyXnqeoWPTkfM0mduRUfyRJCZOsILzKn9yV
H3g34NDkOW9DYCQQxl6BBcDJ80bJt/hAYzLMCkm5nAuQ/+smSckQp/mC3LZTP4vfEJA+cP0Vkxhn
7rebcu0QJh3OjUZdxov2TtdQnTCvfsxr7qgD2EhN5XafR+tXbNXiJst4mmfNHVXU8Gc7KHlkXjeX
g0yGvOfXu8FaoyCIZuxOVlcI6EzS40AvuoeTNgg0OXWGeVtLzfAMGFyL1q325Wssp6iuu5gd8P7m
DpEFePbVMDCFpcBrDYMLEAniW2E6lTCC1mh60z0hs2ibGhRV0BPZ3CxBswbDWBN2GtV7t3DTGTz+
VQcghWX41WrFo+/7DgCzhRKo4XVZSYp8tHFsalDA9Acw/nD0mArswgUWgJ72F0jocDWUJwZzFeu8
7pvr8u2TPkNXsePCNyQq5R6nEK6zhrcjBSytFFVUQ3hMLUI+F7U4LcdiWuqBs42/9Z0EdrvMxlS8
pklSL4ZD0Q2sdm9F5Qffi5eR7ZXgc1SBXhAWIzo2nbx9h9sQHRUCnF36K/jVTicFCatfj6a/f98w
riLyqpnUgy9BQHNsZnjDF+mnT+AsarTh33r6DH6S8geCfVis5/d9deYBMYfHJzHpmD5KMT+ze8Xo
mVfMCNGZKV/ImKIJmx6ad0Nz9yAYvrDFk7MiRe5K3JNDVOMz5bSEMDITRMfIj4v4b0mF7A2r30LR
iWOij+ZPgGWgrlDzD7BL8Ou8P9Kx274VBTPA9aDEwESGpbs0Xgy5Z/uKaOkeOVoAx87iQBy1G6Ky
gW2Q2QbkETE28ZcA9NoDdEUwfEmzBJCE1q8lQf72pAzqna5v0/tLzmbaCqxkqndAapPNdsP/Ofp8
fOSD/CWkyztugFmn/gIVaaw74ELmbLDPGkgBPpHBhtvoHCweMvkIpyUGHl1Jr4Fu1BlB0DI3DRcH
KmJXfIJcENz2g6ME2LQTn3fVWOQi4OHe+e61vI7B8KZp8xZx1GrdpEHuK4AB0CgMuNVMhepsKOWj
frqGkMYq9FGbD0U61REvcbBSq/nMHTJDugoRvi8DNlfkwrL0s9cD4dZWExgTJLOn+9urGVo7bFz1
i2B81/ZwRoRxwICIW0Vi/jd04sCfPF9xmgbdQgGU81j/c1jIX7TdqQlgmk16bCj7JJWvpqt/ts8l
hb5w1DD2GwQW7KmZ8UYRyR9iFNKaK4NFDNumpfyDXwDtCVOtE/oQNA/Zv6C8Rse3pPdg8GFVDKfb
ANxKuuy8okZ/MYAEZKMSTbjVwcm/R1Lz5ynpl8PNSNnPesi1QBYy7Dlt44YYeYC7xVoYjYs/GoKx
kfkaVgd5f8mV2J7XcqofHzzWdyHzlPK/d/HjufbW8SnaIzoQ/O1k7ECuIu5m+D3KvKYElrVluHIe
1eVFzuRZeZC7c+02TZoiq5N0C93FcqsPRtjuoiglcLXSUIWJuEYYLe0NEQQQwKUkUekBL74aSZpR
e/7MUrwJblPxZ7Ss5+z0HS9kUl9dD7uMWSDvtvjHk+9JoPfZ/mDdGRVLvjc+oCFfAqQoFP88H3Oq
dTgCSvL9RqPqGqrpeoad9KGEbVSUSveW2X/zabzwkQDA7kFU8JyMBopBKBACiRISJ0NBgvYpmE5J
xcYYeOwCvsJmmaCgoiU0mf6g+7YsW1Q0Yr5SctEHTQ7E1OT28XKJkh887irpXJUOfa1PKhQLQRlK
cL/a8woZAe84wlIzNJAnTE2PSxrZ9HLKT1fgyB9XtFlB9Ss8wjJmCjfpAagSpzFqYRGPFZUW6I0j
IUhb1pEtR+3ltbvKLmCMe2kPXLOfMIk6fUDHXaz6QLx9INFqPCZgHmdwH7jiefiyMlRobBzAsQqu
ACuuPqqlv1d65FSQ3CqGU67BFYUgMww9tgG62tbyRRZnVw60Yt5xK36nXQtpCkcpEVke9mMm5iIG
/ZWJXp5+0Bqi8Am9eJtVyEQsoSVCkxz99k4K4YF7WAWbWw+P+PcgDVtIYNtzbWfGRjLfbmaZEl4u
NAVCG5oUbVXiNquAlk/a0OL97Run0/qEQ3R+ViTvuA3i7Zifkbpa5dqWrspHBNIRlVLviBijlcas
3VJSjXmgTBMQTII2SfiMpqjcRxvdtunVs1/903zEE87LWolbWtjmvc47kbUtmFY/3spWR8o+lhDX
Wg8fTG/RATXF73hrspSCqvuo7dV4XTXgmDshyrYNqcfdZuzGYg/vjQgYw6Bnzqs9OlFNkoWikTZX
Al+BFzlojvEHvTC4KqGg/mxiVO3DLaTTIiLHOm6LdEM3KpjJuBGlLB+5C/A+rwoCCWcXALVZa14s
dbJd7JgjWxUUstuyyURT+L/Je5SmxfiScxeIE4KZTerFAUEED3BzAjpCbGXmzjFHaCEE9LLFIABP
BSh9lkh6lsbnkBE84mJGmrEC67PWspwkuXNdOqSZ/aaWjXrSgKmOOwVPUC3P+KGErt6R9tHtvE1E
qYwXfy1IekuSCHeBXiOnmwqj7JCLGBQakyXJmhmxaY889ztbJTfZv0fwWpaPGv29n/N4w//t5smQ
fw2NHOsdRS8/cerTzxfjG6iWgmzyvSIxu80RCWqFDHRPA/Wpuk+xgvP11ZHAN34+Lmq+UEIqVFZ6
WQWVIPDPAql00Xe9dRxVsYtYKede0JOzGdsou4quaNTxqWjrC7vgOzaBE9+NlFb8Uc4Sg7ZDTcBs
rL4CyH8n0Z20kebyDfoi/9ccM75ZRALsVHYsQpCjPzGz6VgMhK9/+fFqge4SJq8cdT+V+/d2SHfC
vCbIj/XZO6AlbeOkD1V7y2GXTA3JVtN5zRckTTwcGUM4RyAuXohQ/eVWpRmjWfhGZZwe0OaxqSjl
x1ohS5OnSpclS1Tmi6eS1lr4cdsj38VUjDUm4RxfESg0XZLTBfdSchgFXJ2RlGxBcI8/GSm7NBgW
sQ1FcJ6l+VE2TSBu7spd+oPOVJedlEO3Y7s0DS0xj1HdY540aUhZ/lVYFz73WPisEe8RbHGSL0C1
5p6gZ5Rm4xae+udqImcNExYGrTsvAICWi6UIuddd8nJaZPCQEHXC7qHpcN8caYq7OckDEs3dprdK
EjgriNpmMYIxQwkcr6iw63QTl2SHEWtEjKD66kPgjfOAuX2U+ccE+lRayo8aE5YqT3RJxHI0texM
m2JTFF8oCnxngkwBl1U6DPlqb8s3CuLZHHiiaB30IPmKW2Tf6Dx8jycPTF7oNVqlHRdg3oCdLnSD
as6vWTcr6IuwEaI3NjFmgou98YhlLTzyLhrv6Qhp9r58Fof4rMU2xadFIvCZfAzzbs7qJSQy+1O5
BamrzoYYUJbzO5HHkrHVvXrAlN8ZMFcaRnqTNF/DJ0ZV4+WeXBXir9y7R9wHTWZ/+PkezJM95yOh
v3hfqb6gPrY8PYRKfQ80UvfBpiXA9QRYjyl3TFtdXCCsujkZJc8Mldw5zJB8PLkoX16o+OSfM4V+
Jik0xgMc4rIIxo4lK2t31gLNe6keyMqVB+Ix6xFf7+4awFhQKOiAeRE7eRhHD/13obXj5J6Uugee
MI7AGq1H4loXGJzVDoJmTG4zGz5OHy/UO5YpcQJCvOobGiUHRX7YaJ0A09WBecWudeZIEWmNUS/V
foMnudIesYpYC6QXUtSl7htW8iya5JAC5pKn+JPDRqu+sCjJtBfDhwQL29CNnpmFdHgvXvDGaN06
SB2uLwnDkLJBS5WhB5sVXkblYSeKJU3fQYHn8uPsm8oBKVdDMEsgHxgR/DSNn2HzYLyYgxv9raVJ
QfmY1v5Bn2tjwi2Qq6QDJ1O/GnFGAKJby371qNOXLKE68h9AdV+sXDq/z3mpkXmpfnfkA0gyNQ1T
7imYekqPPB/Tarnk3Qm/vSaCdcSJringCK6hA3marEHQs2j3K3fDUXMwo/WUfvlN36mYO3n0h088
sCW1dGH5qGANTSNvKhv4u6zhpaSxt5jExkcQZqpHLEr6dJWSACj6pRT/KGNOoz9aqE5Z5XwTQTyB
oeRZxP+/j0Ea0cUXcp3s+d/cfMcYbmzxN+5FQDeNp3G2KpC0ICd6dHWNwQwu6g12Ln0AmJ1JbBty
ZGDuQz9PajdezUm8YvrekrAlRgwJz/QTnpQS2IAEp7gG5r068jf6yy9gdp0/u/nofkyTd24jksRN
tNwLqwwbFmKvW7XzSPW3t0LJEx46Q61mScMhv18QbLb3OCg489GXtx5UXMFcXNIY1JK0rt3Lm9qg
/QwBfzLbDaxh/+WvwYpBycLSZPnYdTl8AVyukC9x8i3bXeuEWz47oy43zACUcCkJ/Q8/5CUSfa/i
+npjUjG49UdADS/P3TsvT2jPG3Zh8AhMmuTLeSjnHSm5iskdLd96VDKM26bc3YwiE7WEi3u202ek
9oz64ElvbuipC/+/Qq0dWaABpwFWMO6VHFsKG1sstdzIY6EiS17tFRioO0ZvJ3hJm2oFc67r/4i5
pDQmwoN2tuLUeu34EB5M2Iyl0BexelogiD4+DttLF2gUw0pL6RT9pABjhOFxZ8WaL5Wl9+xnXyXy
6KR9jql9nmSV6E+a4xD/TuGcnGO0OEHO5Tnj96h0WtBvVE1ic6C84J2nYze5cLW0u4cpb+qMaZVf
EOUQ4l3+okVWiwjzJLZ3tWy7pRLV1q0cyXQzKCMYUv4Ck8m7c1f0V//VGhR6YHu7DPiRPFm3O89G
yyrwwRYTyF81EzefAam48Zav1a5cAcZCjOWRRhgaONcfxUA3asPVlYd0/Zh2pSTdO28kjDO1X33x
8mXTJJWaQhYeoRqQhkeNDz7L2c/m12Bom4mm5hYnSTsCJD77yJJgOyXtlsy6ZnjLihkpi/hcCZ5J
W6LmgPZ0Kp0kSVAW/tJx09v4+xf058Ny9QmzVYV7oOamRzUjtHLgBs/0OixatG4pNY3kb37EbouW
pkknhL+vntsCqfkNHnwhVAGtHEX01nWYDbY3zvHOvlmgz9XS/FG7uYfGWlQId+wCSGia2u+ilUYP
XU7XFXbrOXq7kj6KOWIG+dFHMd7b8CO5o5vbtj5r0XI99DdmKb9j0RZGo6eUILxrT/TZhvGUPAgF
m5ZYuNGUGaoL56t1emloB+2HWf2fHQQI5wDhKTgogYazML4ny16BKDhk7KtXfJQsw6V4RoYEk4xA
AlS6NsougJaT+RIuQ2CpyxkS5a5xxHdrKDfiGYyFSb3e9x2UEO6TKeN2fuqcZXpExuTitK47ZM7c
Vvk8YfHC2DJ2xg4/HFUpPmDjhFM//qqfSuSUsDxAvxhudckh2cX6/mqrq5WNLP1p69W8wvXoa0n0
ENbC9HJ+82ig6QqCKC8DuAKFPnBrvFLrc2a5XXCtcIg8I8gxENeoQLH2NLWm2M/F3PuUgPjXHJ3C
njZPNB4muFUfmYSQ7d1jLjQpUu5U8OeKXnjqjBh9wIWNEfn7r/lOwWU5pZVc3OtFRiPqw0KOkWQd
tTusQW/Mx4tC7oypO9CBNth6/xltpLzXonGOLsc8w6XU+pJRD5GXgWv4YaGBkKCAWLHnkFs3K+Cd
qijREBBn02qorTJq68A9q0kxi8bboT+Y7/FLmGUheiD+SnIgWxMpPqOshDjjtbDFfE5njy39B7m0
7YnxDvYSGCkjR3YA0GtcWCz4H8zzFvrbzrGzKcY/wR64bfv6eiRQc7jlZHm/udRb44MT3SCwD1qE
zV9Iiu/rwpHbyd7+RGBDiMlJLLt0xZYvMwFg0jTXCJzC4J9Cugz/Iwf3u4DYp42Ru53CL/m6VuuM
qW8LdR4KGvnqDkh8Tjn1gjRZahNDGXAjyNpZz7kwv305NItF9abLck6AxIG7xYOSxWkjmdaa5Xtn
eZNW5ud4ZppgGnL80JXPerO/VhX5UynNZKG4N4tIJsKRCuqfd+68n0JkstF8kTGVnNT9Jv4ma6tz
bvukzN2m7LRPB4awobFI1yy93sT55Xtk/CKCZHzIafQ4m6apYxg5cKkCPIFdbMMHTxx4s2TyaL9T
KC0Fnxkx3BiKUmlFs7MrjlzElGwzuoahztcMDbZ0DbCbl5I06xlqjtYHwzsEeg==
`protect end_protected

